module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2478, n2426, n2670,
         n2671, n2669, n2685, n2686, n2684, n2718, n2719, n2717, n2982, g2124,
         n2981, n2985, g1430, n2984, n2988, g744, n2987, n2991, g56, n2990,
         n3742, n3741, n8104, g16802, n8103, DFF_1_n1, g16823, n8102, g2950,
         n4423, n4274, g2883, n4330, g22026, g2888, g23358, g2896, n4431,
         g24473, g2892, g25201, g2903, n4305, g26037, g2900, n4291, g26798,
         g2908, n4355, n4273, g2912, n4482, g23357, g2917, n4479, g24476,
         g2924, n4349, g25199, g2920, n4280, DFF_15_n1, n4281, n8099,
         DFF_16_n1, n8098, DFF_18_n1, n4279, g2879, n4351, g2934, g2935, g2938,
         g2941, g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2969, g2972,
         g2975, g2978, g2981, g2874, g18754, g1506, n4288, g18781, g1501,
         n4565, g18803, g1496, n4557, g18821, g1491, n4326, g18835, g1486,
         n4390, g18852, g1481, n4320, g18866, g1476, n4374, g18883, g1471,
         n4378, g21880, g2877, g19154, g813, n4289, g19163, g809, n4567,
         g19173, g805, n4559, g19184, g801, n4327, g20310, g797, n4391, g20343,
         g793, n4321, g20376, g789, n4375, g20417, g785, n4379, g21878, g2873,
         g19153, g125, n4290, g19162, g121, n4569, g19172, g117, n4561, g19144,
         g113, n4328, g19149, g109, n4392, g19157, g105, n4322, g19167, g101,
         n4376, g19178, g97, n4380, g20874, g2857, g18885, g2200, n4287,
         g18975, g2195, n4563, g18968, g2190, n4555, g18942, g2185, n4325,
         g18906, g2180, n4389, g18867, g2175, n4319, g18836, g2170, n4373,
         g18957, g2165, n4377, g21882, g2878, n4598, n4382, n4383, g3109,
         n4494, g18669, g18719, g3211, g18782, g3084, n4445, g17222, g3085,
         g17225, g3086, g17234, g3087, n4344, g17224, g3091, n4448, g17228,
         g3092, n4451, g17246, g3093, g17226, g3094, g17235, g3095, g17269,
         g3096, g25450, g3097, g25451, g3098, n4434, g25452, g3099, n4443,
         g28420, g3100, g28421, g28425, g3102, n4343, g29936, g3103, n4447,
         g29939, g3104, n4452, g29941, g3105, g30796, g3106, n4438, g30798,
         g3107, g30801, g3108, g17229, g3155, g17247, g3158, g17302, g3161,
         n4444, g17236, g3164, g17270, g3167, g17340, g3170, n4441, g17248,
         g3173, n4338, g17303, g3176, n4450, g17383, g17271, g3182, g17341,
         g3185, g17429, g3088, n8090, DFF_131_n1, n8089, DFF_132_n1, g3197,
         n8088, DFF_134_n1, g3201, n4406, g3204, g3207, n4329, g3188, n4405,
         g3133, n8087, g3128, n8086, n8084, DFF_144_n1, g3124, n8083,
         DFF_146_n1, n8082, n8081, n8080, DFF_149_n1, g3112, g3110, g3111,
         n8079, n8078, n8077, DFF_155_n1, n8076, DFF_156_n1, g3151, n4424,
         g3142, n4301, g185, n4384, n4318, n4512, g165, n4369, g22100, g130,
         g22122, g131, g22141, g129, g22123, g133, g22142, g134, g22161, g132,
         g22025, g142, g22027, g143, g22030, g141, g22028, g145, g22031, g146,
         g22037, g22032, g148, g22038, g149, g22047, g147, g22039, g151,
         g22048, g152, g22063, g150, g22049, g154, g22064, g155, g22079, g153,
         g22065, g157, g22080, g158, g22101, g156, g22081, g160, g22102, g161,
         g22124, g159, g22103, g22125, g164, g22143, g162, g25204, g169,
         g25206, g170, g25211, g168, g25207, g172, g25212, g173, g25218, g171,
         g25213, g175, g25219, g176, g25228, g174, g25220, g178, g25229, g179,
         g25239, g177, g30261, g186, g30267, g30275, g192, g30637, g231,
         g30640, g234, g30645, g237, g30668, g195, g30674, g198, g30680, g201,
         g30641, g240, g30646, g243, g30653, g246, g30276, g204, g30284, g207,
         g30292, g210, g30254, g249, g30257, g252, g30262, g30245, g213,
         g30246, g216, g30248, g219, g30258, g258, g30263, g261, g30268, g264,
         g30635, g222, g30636, g225, g30639, g228, g30661, g267, g30669, g270,
         g30675, g273, g25027, g92, g25932, g88, g26529, g83, g27120, g27594,
         g74, g28145, g70, g28634, g65, g29109, g61, g29353, g29579, g52,
         g13110, g180, g181, n4506, g309, n4388, g27253, g354, g27255, g343,
         g27258, g27256, g369, g27259, g358, g27265, g361, g27260, g384,
         g27266, g373, g27277, g376, g27267, g398, g27278, g388, g27293, g391,
         g28732, g408, g28735, g411, g28744, g414, g29194, g417, g29197, g420,
         g29201, g423, g28736, g28745, g428, g28754, g426, g26803, g429,
         g26804, g432, g26807, g435, g26805, g438, g26808, g441, g26812, g444,
         g27759, g448, g27760, g449, g27762, g447, g29606, g312, g29608, g313,
         g29611, g314, g30699, g315, g30700, g30702, g317, g30455, g318,
         g30468, g319, g30482, g320, g29167, g322, g29169, g323, g29172, g321,
         g26655, g403, g26659, g404, g26664, g402, g450, n8066, DFF_299_n1,
         g452, n8065, DFF_301_n1, g454, DFF_303_n1, g280, n8062, DFF_305_n1,
         g282, n8061, DFF_307_n1, g284, n8060, DFF_309_n1, g286, n8059,
         DFF_311_n1, g288, n8058, DFF_313_n1, g290, n8057, n4485, n4282, n8056,
         g21346, g305, n4278, n8055, DFF_328_n1, g349, g350, g351, g352, g353,
         g357, g364, g365, g366, g367, g368, g372, g379, g380, g381, g383,
         g387, g394, g395, g396, g397, g324, g337, n4298, n4372, g550, n4313,
         g21842, g554, g18678, g557, n4360, g18726, g513, g523, g524, g455,
         g564, g569, g458, g570, g571, g461, g572, g573, g465, g574, g565,
         g566, g567, g471, g568, g489, n4461, g485, n4466, g23067, g486,
         g23093, g487, g23117, g488, g23385, g23399, g24174, g24178, g477,
         g24207, g478, g24216, g479, g23092, g480, g23000, g484, g23022, g464,
         g24206, g24215, g24228, g528, g535, g542, g13149, g543, g544, g21851,
         g548, g13111, g549, g499, n4541, g13160, g558, g559, g27261, g576,
         g27268, g577, g27279, g575, g27269, g579, g27280, g27294, g578,
         g27281, g582, g27295, g583, g27311, g581, g27296, g585, g27312, g586,
         g27327, g584, g24491, g587, g24498, g590, g24507, g593, g24499, g596,
         g24508, g599, g24519, g602, g28345, g614, g28349, g617, g28353,
         g28342, g605, g28344, g608, g28348, g611, g26541, g490, g26545, g493,
         g26553, g496, g506, n4570, g22578, n4571, g525, n8047, DFF_444_n1,
         n8046, DFF_445_n1, n8045, DFF_446_n1, n8044, DFF_447_n1, n8043,
         DFF_448_n1, DFF_449_n1, g536, g537, g24059, g538, n4492, n8040, n4359,
         g629, n4295, g16654, g630, g20314, g659, g20682, g640, n4404, g23136,
         g633, n4478, g23324, g653, n4422, g24426, g646, n4414, g25185, g660,
         n4403, g26660, g672, n4413, g26776, g27672, g679, n4477, g28199, g686,
         n4396, g28668, g692, n4418, g20875, g699, g20879, g700, g20891, g698,
         g20880, g702, g20892, g703, g20901, g701, g20893, g705, g20902, g706,
         g20921, g704, g20903, g708, g20922, g709, g20944, g707, g20923,
         g20945, g712, g20966, g710, g20946, g714, g20967, g715, g20989, g713,
         g20968, g717, g20990, g718, g21009, g716, g20991, g720, g21010, g721,
         g21031, g719, g21011, g723, g21032, g724, g21051, g722, g20876, g726,
         g20881, g20894, g725, g20924, g729, g20947, g730, g20969, g728,
         g20948, g732, g20970, g733, g20992, g731, g25260, g735, g25262, g736,
         g25266, g734, g22218, g738, g22231, g739, g22242, g737, n4323, n4312,
         g22126, g818, g22145, g819, g22162, g817, g22146, g821, g22163, g822,
         g22177, g820, g22029, g830, g22033, g831, g22040, g829, g22034, g833,
         g22041, g834, g22054, g832, g22042, g836, g22055, g837, g22066, g835,
         g22056, g22067, g840, g22087, g838, g22068, g842, g22088, g843,
         g22104, g841, g22089, g845, g22105, g846, g22127, g844, g22106, g848,
         g22128, g849, g22147, g847, g22129, g851, g22148, g852, g22164, g850,
         g25209, g857, g25214, g25221, g856, g25215, g860, g25222, g861,
         g25230, g859, g25223, g863, g25231, g864, g25240, g862, g25232, g866,
         g25241, g867, g25248, g865, g30269, g873, g30277, g876, g30285, g879,
         g30643, g918, g30648, g921, g30654, g30676, g882, g30681, g885,
         g30687, g888, g30649, g927, g30655, g930, g30662, g933, g30286, g891,
         g30293, g894, g30298, g897, g30259, g936, g30264, g939, g30270, g942,
         g30247, g900, g30249, g903, g30251, g906, g30265, g30271, g948,
         g30278, g951, g30638, g909, g30642, g912, g30647, g915, g30670, g954,
         g30677, g957, g30682, g960, g25042, g780, g25935, g776, g26530, g771,
         g27123, g767, g27603, g762, g28146, g758, g28635, g753, g29110,
         g29354, g29580, g740, g868, g869, n4363, n4364, g1088, n4381, g996,
         n4387, g27257, g1041, g27262, g1030, g27270, g1033, g27263, g1056,
         g27271, g1045, g27282, g1048, g27272, g27283, g1060, g27297, g1063,
         g27284, g1085, g27298, g1075, g27313, g1078, g28738, g1095, g28746,
         g1098, g28758, g1101, g29198, g1104, g29204, g1107, g29209, g1110,
         g28747, g1114, g28759, g1115, g28767, g1113, g26806, g1116, g26809,
         g26813, g1122, g26810, g1125, g26814, g1128, g26818, g1131, g27761,
         g1135, g27763, g1136, g27765, g1134, g29609, g999, g29612, g1000,
         g29616, g1001, g30701, g1002, g30703, g1003, g30705, g1004, g30470,
         g1005, g30485, g1006, g30500, g29170, g1009, g29173, g1010, g29179,
         g1008, g26661, g1090, g26665, g1091, g26669, g1089, g1137, n8027,
         DFF_649_n1, g1139, n8026, DFF_651_n1, g1141, n8025, DFF_653_n1, g967,
         n8024, DFF_655_n1, g969, DFF_657_n1, g971, n8021, DFF_659_n1, g973,
         n8020, DFF_661_n1, g975, n8019, DFF_663_n1, g977, n8018, n4486, n4283,
         g986, n4432, g26183, g992, n4277, n8017, g1029, g1036, g1037, g1038,
         g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067,
         g1068, g1069, g1070, g1074, g1081, g1083, g1084, g1011, g1024, n4371,
         n4316, g1236, n4300, g21843, g1240, g18707, g1243, n4353, g18763,
         g1196, n4304, g1199, g1209, g1210, g1142, g1255, g1145, g1256, g1257,
         g1148, g1258, g1259, g1152, g1260, g1251, g1155, g1252, g1253, g1158,
         g1254, g1176, n4460, n4459, g1172, n4465, g23081, g1173, g23111,
         g23126, g1175, g23392, g23406, g24179, g24181, g1164, g24213, g1165,
         g24223, g1166, g23110, g1167, g23014, g1171, g23039, g1151, g24212,
         g24222, g24235, g1214, g1221, g13155, g1229, n4549, n4361, g13124,
         g1235, g1186, n4548, g13171, g1244, g1245, g27273, g1262, g27285,
         g1263, g27299, g1261, g27286, g1265, g27300, g1266, g27314, g1264,
         g27301, g1268, g27315, g1269, g27328, g27316, g1271, g27329, g1272,
         g27339, g1270, g24501, g1273, g24510, g1276, g24521, g1279, g24511,
         g1282, g24522, g1285, g24532, g1288, g28351, g1300, g28355, g1303,
         g28360, g1306, g28346, g1291, g28350, g1294, g28354, g1297, g26547,
         g26557, g1180, g26569, g1183, g1192, n4454, g22615, n8009, DFF_783_n1,
         DFF_792_n1, g1211, n8008, DFF_794_n1, n8007, DFF_795_n1, n8006,
         DFF_796_n1, n8005, DFF_797_n1, n8004, DFF_798_n1, n8003, DFF_799_n1,
         g1222, g1223, g24072, g1224, n4489, n4358, g1315, n4294, g16671,
         g1316, g20333, g1345, n4428, g20717, g1326, n4402, g21969, g1319,
         n4476, g23329, g1339, n4421, g24430, g1332, n4412, g25189, g1346,
         n4401, g26666, g1358, n4411, g26781, g1352, n4469, g27678, g1365,
         n4475, g27718, g1372, n4395, g28321, g1378, n4417, g20882, g20896,
         g1386, g20910, g1384, g20897, g1388, g20911, g1389, g20925, g1387,
         g20912, g1391, g20926, g1392, g20949, g1390, g20927, g1394, g20950,
         g1395, g20972, g1393, g20951, g1397, g20973, g1398, g20993, g1396,
         g20974, g1400, g20994, g21015, g1399, g20995, g1403, g21016, g1404,
         g21033, g1402, g21017, g1406, g21034, g1407, g21052, g1405, g21035,
         g1409, g21053, g1410, g21070, g1408, g20883, g1412, g20898, g1413,
         g20913, g1411, g20952, g1415, g20975, g1416, g20996, g20976, g1418,
         g20997, g1419, g21018, g1417, g25263, g1421, g25267, g1422, g25270,
         g1420, g22234, g1424, g22247, g1425, g22263, g1423, n4317, n4515,
         g1547, n4368, g22149, g1512, g22166, g1513, g22178, g1511, g22167,
         g22179, g1516, g22191, g1514, g22035, g1524, g22043, g1525, g22057,
         g1523, g22044, g1527, g22058, g1528, g22073, g1526, g22059, g1530,
         g22074, g1531, g22090, g1529, g22075, g1533, g22091, g1534, g22112,
         g1532, g22092, g1536, g22113, g22130, g1535, g22114, g1539, g22131,
         g1540, g22150, g1538, g22132, g1542, g22151, g1543, g22168, g1541,
         g22152, g1545, g22169, g1546, g22180, g1544, g25217, g1551, g25224,
         g1552, g25233, g1550, g25225, g1554, g25234, g1555, g25242, g25235,
         g1557, g25243, g1558, g25249, g1556, g25244, g1560, g25250, g1561,
         g25255, g1559, g30279, g1567, g30287, g1570, g30294, g1573, g30651,
         g1612, g30657, g1615, g30663, g1618, g30683, g1576, g30688, g1579,
         g30692, g1582, g30658, g30664, g1624, g30671, g1627, g30295, g1585,
         g30299, g1588, g30302, g1591, g30266, g1630, g30272, g1633, g30280,
         g1636, g30250, g1594, g30252, g1597, g30255, g1600, g30273, g1639,
         g30281, g1642, g30288, g1645, g30644, g1603, g30650, g30656, g1609,
         g30678, g1648, g30684, g1651, g30689, g1654, g25056, g1466, g25938,
         g1462, g26531, g1457, g27129, g1453, g27612, g1448, g28147, g1444,
         g28636, g1439, g29111, g1435, g29355, g29581, g1426, g1562, g1563,
         n4518, g1690, n4386, g27264, g1735, g27274, g1724, g27287, g1727,
         g27275, g1750, g27288, g1739, g27302, g1742, g27289, g1765, g27303,
         g1754, g27317, g1757, g27304, g1779, g27318, g27330, g1772, g28749,
         g1789, g28760, g1792, g28771, g1795, g29205, g1798, g29212, g1801,
         g29218, g1804, g28761, g1808, g28772, g1809, g28778, g1807, g26811,
         g1810, g26815, g1813, g26820, g1816, g26816, g1819, g26821, g1822,
         g26824, g27764, g1829, g27766, g1830, g27768, g1828, g29613, g1693,
         g29617, g1694, g29620, g1695, g30704, g1696, g30706, g1697, g30708,
         g1698, g30487, g1699, g30503, g1700, g30338, g1701, g29178, g1703,
         g29181, g1704, g29184, g1702, g26667, g26670, g1785, g26675, g1783,
         g1831, n7988, DFF_999_n1, g1833, n7987, DFF_1001_n1, g1835, n7986,
         DFF_1003_n1, g1661, n7985, DFF_1005_n1, g1663, n7984, DFF_1007_n1,
         g1665, n7983, DFF_1009_n1, g1667, DFF_1011_n1, g1669, n7980,
         DFF_1013_n1, g1671, n7979, n4484, n4284, g1680, n4488, g28903, g1686,
         n4276, n7978, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745,
         g1747, g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768,
         g1775, g1776, g1777, g1778, g1705, g1718, n4296, n4315, g1930, n4366,
         g21845, g1934, g18743, g1937, n4311, g18794, g1890, n4297, g1893,
         g1903, g1904, g1836, g1944, g1949, g1950, g1951, g1842, g1953, g1846,
         g1954, g1945, g1849, g1946, g1947, g1852, g1948, g1870, n4458, n4457,
         g1866, n4464, g23097, g1867, g23124, g1868, g23137, g1869, g23400,
         g23413, g24182, g24208, g1858, g24219, g1859, g24231, g1860, g23123,
         g1861, g23030, g1865, g23058, g1845, g24218, g24230, g24243, g1908,
         g1915, g1922, g13164, g1923, DFF_1099_n1, n7971, g13135, g1929, g1880,
         n4545, g13182, g1938, g1939, g27290, g1956, g27305, g1957, g27319,
         g1955, g27306, g1959, g27320, g1960, g27331, g1958, g27321, g1962,
         g27332, g1963, g27340, g1961, g27333, g27341, g1966, g27346, g1964,
         g24513, g1967, g24524, g1970, g24534, g1973, g24525, g1976, g24535,
         g1979, g24545, g1982, g28357, g1994, g28362, g1997, g28366, g2000,
         g28352, g1985, g28356, g1988, g28361, g1991, g26559, g26573, g1874,
         g26592, g1877, g1886, n4493, g22651, n7968, DFF_1133_n1, g28990,
         DFF_1142_n1, g1905, n7967, DFF_1144_n1, n7966, DFF_1145_n1, n7965,
         DFF_1146_n1, n7964, DFF_1147_n1, n7963, DFF_1148_n1, n7962,
         DFF_1149_n1, g1916, g1917, g24083, n7960, n4357, g2009, n4293, g16692,
         g2010, g20353, g2039, n4427, g20752, g2020, n4400, g21972, g2013,
         n4474, g23339, g2033, n4420, g24434, g2026, n4410, g25194, g2040,
         n4399, g26671, g2052, n4409, g26789, g2046, n4468, g27682, g2059,
         n4473, g27722, g28325, g2072, n4416, g20899, g2079, g20915, g2080,
         g20934, g2078, g20916, g2082, g20935, g2083, g20953, g2081, g20936,
         g2085, g20954, g2086, g20977, g2084, g20955, g2088, g20978, g2089,
         g20999, g2087, g20979, g2091, g21000, g21019, g2090, g21001, g2094,
         g21020, g2095, g21039, g2093, g21021, g2097, g21040, g2098, g21054,
         g2096, g21041, g2100, g21055, g2101, g21071, g2099, g21056, g2103,
         g21072, g2104, g21080, g2102, g20900, g2106, g20917, g20937, g2105,
         g20980, g2109, g21002, g2110, g21022, g2108, g21003, g2112, g21023,
         g2113, g21042, g2111, g25268, g2115, g25271, g2116, g25279, g2114,
         g22249, g2118, g22267, g2119, g22280, g2117, n4324, g2241, n4367,
         g22170, g2206, g22182, g2207, g22192, g2205, g22183, g2209, g22193,
         g2210, g22200, g2208, g22045, g2218, g22060, g2219, g22076, g2217,
         g22061, g2221, g22077, g2222, g22097, g2220, g22078, g2224, g22098,
         g22115, g2223, g22099, g2227, g22116, g2228, g22138, g2226, g22117,
         g2230, g22139, g2231, g22153, g2229, g22140, g2233, g22154, g2234,
         g22171, g2232, g22155, g2236, g22172, g2237, g22184, g2235, g22173,
         g2239, g22185, g22194, g2238, g25227, g2245, g25236, g2246, g25245,
         g2244, g25237, g2248, g25246, g2249, g25251, g2247, g25247, g2251,
         g25252, g2252, g25256, g2250, g25253, g2254, g25257, g2255, g25259,
         g2253, g30289, g2261, g30296, g30300, g2267, g30660, g2306, g30666,
         g2309, g30672, g2312, g30690, g2270, g30693, g2273, g30695, g2276,
         g30667, g2315, g30673, g2318, g30679, g2321, g30301, g2279, g30303,
         g2282, g30304, g2285, g30274, g2324, g30282, g30290, g2330, g30253,
         g2288, g30256, g2291, g30260, g2294, g30283, g2333, g30291, g2336,
         g30297, g2339, g30652, g2297, g30659, g2300, g30665, g2303, g30686,
         g2342, g30691, g2345, g30694, g2348, g25067, g2160, g25940, g26532,
         g2151, g27131, g2147, g27621, g2142, g28148, g2138, g28637, g2133,
         g29112, g2129, g29357, g29582, g2120, g2256, g2257, n4516, g27276,
         g2429, g27291, g2418, g27307, g2421, g27292, g2444, g27308, g2433,
         g27322, g2436, g27309, g2459, g27323, g2448, g27334, g2451, g27324,
         g2473, g27335, g2463, g27342, g2466, g28763, g2483, g28773, g2486,
         g28782, g29213, g2492, g29221, g2495, g29226, g2498, g28774, g2502,
         g28783, g2503, g28788, g2501, g26817, g2504, g26822, g2507, g26825,
         g2510, g26823, g2513, g26826, g2516, g26827, g2519, g27767, g2523,
         g27769, g2524, g27771, g29618, g2387, g29621, g2388, g29623, g2389,
         g30707, g2390, g30709, g2391, g30566, g2392, g30505, g2393, g30341,
         g2394, g30356, g2395, g29182, g2397, g29185, g2398, g29187, g2396,
         g26672, g2478, g26676, g2479, g26025, g2525, n7946, DFF_1349_n1,
         g2527, n7945, DFF_1351_n1, g2529, n7944, DFF_1353_n1, g2355, n7943,
         DFF_1355_n1, g2357, n7942, DFF_1357_n1, g2359, n7941, DFF_1359_n1,
         g2361, n7940, DFF_1361_n1, n7938, DFF_1363_n1, g2365, n7937, n4483,
         n4285, g2374, n4487, g30055, g2380, n4275, n7936, DFF_1378_n1, g2417,
         g2424, g2425, g2426, g2427, g2428, g2432, g2439, g2441, g2442, g2443,
         g2447, g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471,
         g2472, g2412, n4314, n4370, g2624, n4299, g21847, g2628, g18780,
         g2631, n4352, g18820, g2584, n4303, g2587, g2597, g2598, g2530, g2638,
         g2643, g2533, g2645, g2536, g2646, g2647, g2540, g2648, g2639, g2543,
         g2640, g2641, g2546, g2642, g2564, n4456, n4455, g2560, n4463, g23114,
         g2561, g23133, g2562, g21970, g23407, g23418, g24209, g24214, g2552,
         g24226, g2553, g24238, g2554, g23132, g2555, g23047, g2559, g23076,
         g2539, g24225, g24237, g24250, g2602, g2609, g13175, g2617, n7930,
         g30072, n7929, g13143, g2623, g2574, n4543, g13194, g2632, g2633,
         g27310, g2650, g27325, g2651, g27336, g2649, g27326, g2653, g27337,
         g2654, g27343, g2652, g27338, g2656, g27344, g27347, g2655, g27345,
         g2659, g27348, g2660, g27354, g2658, g24527, g2661, g24537, g2664,
         g24547, g2667, g24538, g2670, g24548, g2673, g24557, g2676, g28364,
         g2688, g28368, g2691, g28371, g2694, g28358, g2679, g28363, g28367,
         g2685, g26575, g2565, g26596, g2568, g26616, g2571, g2580, g22687,
         n7926, g30061, g2599, n7925, DFF_1494_n1, n7924, DFF_1495_n1, n7923,
         DFF_1496_n1, n7922, DFF_1497_n1, n7921, DFF_1498_n1, n7920,
         DFF_1499_n1, g2611, g24092, g2612, n4490, n7918, n4356, g2703, n4292,
         g16718, g2704, g20375, g2733, g20789, g2714, n4398, g21974, g2707,
         n4472, g23348, g2727, n4419, g24438, g2720, n4408, g25197, g2734,
         n4397, g26677, g2746, n4407, g26795, g27243, g2753, n4471, g27724,
         g2760, n4393, g28328, g2766, n4415, g20918, g2773, g20939, g2774,
         g20962, g2772, g20940, g2776, g20963, g2777, g20981, g2775, g20964,
         g2779, g20982, g2780, g21004, g2778, g20983, g2782, g21005, g2783,
         g21025, g21006, g2785, g21026, g2786, g21043, g2784, g21027, g2788,
         g21044, g2789, g21060, g2787, g21045, g2791, g21061, g2792, g21073,
         g2790, g21062, g2794, g21074, g2795, g21081, g2793, g21075, g2797,
         g21082, g2798, g21094, g20919, g2800, g20941, g2801, g20965, g2799,
         g21007, g2803, g21028, g2804, g21046, g2802, g21029, g2806, g21047,
         g2807, g21063, g2805, g25272, g2809, g25280, g2810, g25288, g2808,
         g22269, g2812, g22284, g2813, g22299, g20877, n7913, DFF_1561_n1,
         g20884, n7912, DFF_1562_n1, n4263_Tj_Payload, n4269, g3043, n4268,
         g3044, n4267, g3045, n4266, g3046, n4265, g3047, n4272, g3048, n4271,
         g3049, n4270, g3050, n4259, g3051, n4236, g3052, n4239, g3053, n4237,
         n4234, g3056, n4233, g3057, n4238, g3058, n4235, g3059, n4240, g3060,
         n4232, g3061, n4245, g3062, n4248, g3063, n4246, g3064, n4243, g3065,
         n4242, g3066, n4247, g3067, n4244, g3068, n4249, g3069, n4241, n4254,
         g3071, n4257, g3072, n4255, g3073, n4252, g3074, n4251, g3075, n4256,
         g3076, n4253, g3077, n4258, g3078, n4250, g2997, g25265, g2993,
         g26048, n7909, g23330, g3006, g24445, g3002, g25191, g3013, g26031,
         g26786, g3024, n4262, g3018, n4481, g23359, g3028, n4350, g24446,
         g3036, n4480, g25202, g3032, n7907, DFF_1612_n1, g2987, n4365, g16824,
         g16844, g16853, g16860, g16803, g16835, g16851, g16857, g16866, g3083,
         n4261, N995, n4577, g16845, g16854, g16861, g16880, g18755, g18804,
         g18837, g18868, g18907, g2990, N690, n4578, n4260, n4309, n4308,
         n4307, n4306, n4524, n4525, n4511, n4509, n4499, n4520, n3683, n3887,
         n3686, n3890, n3692, n3896, n4513, n3897, n3424, n3427, n3433, n4529,
         n4530, n4522, n4523, n4521, n3171, n3159, n3163, n3893, n3690, n3689,
         n3431, n3430, n3168, n3160, n3164, n3172, n4527, n4528, n4526, n2313,
         n3167, n3894, n3888, n3891, n2302, n2289, n2303, n2275, n4066, n4065,
         n4606, n4618, n4640, n2351, n2430, n2792, n2632, n3936, n3253, n3252,
         n3254, n4102, n3038, n3070, n3102, n3130, n3036, n3068, n3065, n3128,
         n2800, n2798, n2616, n2594, n3940, n3705, n3933, n3939, n3016, n3000,
         n3008, n3023, n3700, n4058, n4123, n4101, n3938, n4182, n3944, n4073,
         n3749, n3751, n3758, n3788, n4057, n4122, n4263, Tj_OUT1, Tj_OUT2,
         Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8,
         Tj_OUT5678, Tj_Trigger, n19, n63, n129, n138, n144, n167, n257, n264,
         n265, n266, n335, n433, n440, n509, n598, n605, n673, n758, n765,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6681, n6682, n6706,
         n6707, n6708, n6709, n6710, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6834, n6836, n6837, n6838, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6969, n6970, n6971, n6972, n6973, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7041, n7042,
         n7043, n7044, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7908, n7910,
         n7911, n7914, n7915, n7916, n7917, n7919, n7927, n7928, n7931, n7932,
         n7933, n7934, n7935, n7939, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7961, n7969, n7970,
         n7972, n7973, n7974, n7975, n7976, n7977, n7981, n7982, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8022,
         n8023, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8041, n8042, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8063, n8064, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8085, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8100, n8101, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, U4467_n1, U4904_n1, U4930_n1, U5128_n1, U5141_n1, U5749_n1,
         U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1,
         U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1,
         U5764_n1, U5882_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U6140_n1,
         U6460_n1, U6470_n1, U6562_n1, U6563_n1, U6718_n1, U7116_n1, U7118_n1,
         U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n7277), .CLK(n7464), .Q(
        n8104), .QN(n13231) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n7277), .CLK(n7464), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n7277), .CLK(n7464), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n7277), .CLK(n7464), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n7278), .CLK(n7465), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n7278), .CLK(n7465), .Q(
        g2888), .QN(n7049) );
  SDFFX1 DFF_6_Q_reg ( .D(g23358), .SI(g2888), .SE(n7278), .CLK(n7465), .Q(
        g2896), .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n7278), .CLK(n7465), .Q(
        g2892), .QN(n7048) );
  SDFFX1 DFF_8_Q_reg ( .D(g25201), .SI(g2892), .SE(n7278), .CLK(n7465), .Q(
        g2903), .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n7278), .CLK(n7465), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n7278), .CLK(n7465), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n7278), .CLK(n7465), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n7278), .CLK(n7465), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n7278), .CLK(n7465), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n7278), .CLK(n7465), .Q(
        g2920), .QN(n6995) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n7278), .CLK(n7465), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n7275), .CLK(n7462), .Q(
        n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n7275), .CLK(n7462), .Q(g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n7275), .CLK(n7462), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n7275), .CLK(n7462), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n7275), .CLK(n7462), .Q(
        g2934), .QN(n7262) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n7275), .CLK(n7462), .Q(
        g2935), .QN(n7243) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n7276), .CLK(n7463), .Q(
        g2938), .QN(n7244) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n7276), .CLK(n7463), .Q(
        g2941), .QN(n7241) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n7276), .CLK(n7463), .Q(
        g2944) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n7276), .CLK(n7463), .Q(
        g2947), .QN(n7245) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n7276), .CLK(n7463), .Q(
        g2953), .QN(n7246) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n7276), .CLK(n7463), .Q(
        g2956), .QN(n7248) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n7276), .CLK(n7463), .Q(
        g2959), .QN(n7242) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n7276), .CLK(n7463), .Q(
        g2962), .QN(n7260) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n7276), .CLK(n7463), .Q(
        g2963), .QN(n7251) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n7276), .CLK(n7463), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n7275), .CLK(n7462), .Q(
        g2969), .QN(n7254) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n7275), .CLK(n7462), .Q(
        g2972), .QN(n7252) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n7275), .CLK(n7462), .Q(
        g2975), .QN(n7253) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n7275), .CLK(n7462), .Q(
        g2978), .QN(n7249) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n7275), .CLK(n7462), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n7275), .CLK(n7462), .Q(
        g2874), .QN(n7250) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n7276), .CLK(n7463), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n7276), .CLK(n7463), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n7277), .CLK(n7464), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n7277), .CLK(n7464), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n7277), .CLK(n7464), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n7277), .CLK(n7464), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n7277), .CLK(n7464), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n7277), .CLK(n7464), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n7285), .CLK(n7472), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n7285), .CLK(n7472), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n7285), .CLK(n7472), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n7285), .CLK(n7472), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n7285), .CLK(n7472), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n7285), .CLK(n7472), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n7285), .CLK(n7472), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n7285), .CLK(n7472), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n7286), .CLK(n7473), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n7286), .CLK(n7473), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n7286), .CLK(n7473), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n7286), .CLK(n7473), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n7286), .CLK(n7473), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n7286), .CLK(n7473), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n7286), .CLK(n7473), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n7286), .CLK(n7473), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n7286), .CLK(n7473), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n7299), .CLK(n7486), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n7299), .CLK(n7486), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n7301), .CLK(n7488), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n7301), .CLK(n7488), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n7302), .CLK(n7489), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n7302), .CLK(n7489), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n7302), .CLK(n7489), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n7302), .CLK(n7489), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n7302), .CLK(n7489), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n7302), .CLK(n7489), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n7302), .CLK(n7489), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n7302), .CLK(n7489), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n7302), .CLK(n7489), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n7302), .CLK(n7489), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n7302), .CLK(n7489), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n7302), .CLK(n7489), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n7303), .CLK(n7490), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n7303), .CLK(n7490), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n7303), .CLK(n7490), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n7303), .CLK(n7490), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n7303), .CLK(n7490), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n7303), .CLK(n7490), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n7303), .CLK(n7490), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n7303), .CLK(n7490), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n7303), .CLK(n7490), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n7303), .CLK(n7490), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n7303), .CLK(n7490), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n7303), .CLK(n7490), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n7318), .CLK(n7505), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n7401), .CLK(n7588), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n7401), .CLK(n7588), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n7401), .CLK(n7588), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n7402), .CLK(n7589), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n7402), .CLK(n7589), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n7402), .CLK(n7589), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n7403), .CLK(n7590), .Q(
        g3085) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n7404), .CLK(n7591), .Q(
        g3086) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n7404), .CLK(n7591), .Q(
        g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n7404), .CLK(n7591), .Q(
        g3091), .QN(n4448) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n7404), .CLK(n7591), .Q(
        g3092), .QN(n4451) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n7404), .CLK(n7591), .Q(
        g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n7404), .CLK(n7591), .Q(
        g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n7404), .CLK(n7591), .Q(
        g3095) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n7404), .CLK(n7591), .Q(
        g3096) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n7404), .CLK(n7591), .Q(
        g3097) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n7404), .CLK(n7591), .Q(
        g3098), .QN(n4434) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n7404), .CLK(n7591), .Q(
        g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n7404), .CLK(n7591), .Q(
        g3100) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n7405), .CLK(n7592), .Q(
        test_so7) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n7402), .CLK(n7589), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n7402), .CLK(n7589), .Q(
        g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n7402), .CLK(n7589), .Q(
        g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n7402), .CLK(n7589), .Q(
        g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n7402), .CLK(n7589), .Q(
        g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n7403), .CLK(n7590), .Q(
        g3107) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n7403), .CLK(n7590), .Q(
        g3108) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n7403), .CLK(n7590), .Q(
        g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n7403), .CLK(n7590), .Q(
        g3158) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n7403), .CLK(n7590), .Q(
        g3161), .QN(n4444) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n7403), .CLK(n7590), .Q(
        g3164) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n7403), .CLK(n7590), .Q(
        g3167) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n7403), .CLK(n7590), .Q(
        g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n7403), .CLK(n7590), .Q(
        g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n7403), .CLK(n7590), .Q(
        g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n7403), .CLK(n7590), .Q(
        test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n7402), .CLK(n7589), 
        .Q(g3182) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n7402), .CLK(n7589), .Q(
        g3185) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n7402), .CLK(n7589), .Q(
        g3088) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n7402), .CLK(n7589), .Q(
        n8090), .QN(DFF_131_n1) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n7283), .CLK(n7470), .Q(
        n8089), .QN(DFF_132_n1) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n7405), .CLK(n7592), .Q(
        g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n7405), .CLK(n7592), .Q(
        n8088), .QN(DFF_134_n1) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n7283), .CLK(n7470), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n7283), .CLK(n7470), .Q(
        g3204) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n7283), .CLK(n7470), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n7282), .CLK(n7469), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n19), .SI(g3188), .SE(n7283), .CLK(n7470), .Q(
        g3133), .QN(n6707) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n7283), .CLK(n7470), .Q(
        n8087) );
  SDFFX1 DFF_141_Q_reg ( .D(n129), .SI(n8087), .SE(n7283), .CLK(n7470), .Q(
        g3128), .QN(n6894) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n7283), .CLK(n7470), .Q(
        n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n7284), .CLK(n7471), .Q(
        test_so9) );
  SDFFX1 DFF_144_Q_reg ( .D(n138), .SI(test_si10), .SE(n7283), .CLK(n7470), 
        .Q(n8084), .QN(DFF_144_n1) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n7283), .CLK(n7470), .Q(
        g3124) );
  SDFFX1 DFF_146_Q_reg ( .D(n144), .SI(g3124), .SE(n7283), .CLK(n7470), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n7283), .CLK(n7470), .Q(
        n8082) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n7284), .CLK(n7471), .Q(
        n8081) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n7284), .CLK(n7471), .Q(
        n8080), .QN(DFF_149_n1) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n7284), .CLK(n7471), .Q(
        g3112) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n7284), .CLK(n7471), .Q(
        g3110) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n7284), .CLK(n7471), .Q(
        g3111) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n7284), .CLK(n7471), .Q(
        n8079), .QN(n13232) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n7284), .CLK(n7471), .Q(
        n8078), .QN(n13233) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n7284), .CLK(n7471), .Q(
        n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n7284), .CLK(n7471), .Q(
        n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n7284), .CLK(n7471), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n7284), .CLK(n7471), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n7285), .CLK(n7472), .Q(
        test_so10), .QN(n7274) );
  SDFFX1 DFF_160_Q_reg ( .D(n19), .SI(test_si11), .SE(n7281), .CLK(n7468), .Q(
        g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n7281), .CLK(n7468), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n7281), .CLK(n7468), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n7282), .CLK(n7469), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n7305), .CLK(n7492), .Q(
        g130), .QN(n7225) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n7305), .CLK(n7492), .Q(
        g131), .QN(n7224) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n7305), .CLK(n7492), .Q(
        g129), .QN(n6831) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n7305), .CLK(n7492), .Q(
        g133), .QN(n7223) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n7305), .CLK(n7492), .Q(
        g134), .QN(n7222) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n7305), .CLK(n7492), .Q(
        g132), .QN(n6830) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n7305), .CLK(n7492), .Q(
        g142), .QN(n7221) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n7306), .CLK(n7493), .Q(
        g143), .QN(n7220) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n7306), .CLK(n7493), .Q(
        g141), .QN(n6829) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n7306), .CLK(n7493), .Q(
        g145), .QN(n7219) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n7306), .CLK(n7493), .Q(
        g146), .QN(n7218) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n7306), .CLK(n7493), .Q(
        test_so11) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n7306), .CLK(n7493), 
        .Q(g148), .QN(n7217) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n7306), .CLK(n7493), .Q(
        g149), .QN(n7216) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n7306), .CLK(n7493), .Q(
        g147), .QN(n6828) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n7307), .CLK(n7494), .Q(
        g151), .QN(n7215) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n7308), .CLK(n7495), .Q(
        g152), .QN(n7214) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n7308), .CLK(n7495), .Q(
        g150), .QN(n6827) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n7308), .CLK(n7495), .Q(
        g154), .QN(n7213) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n7308), .CLK(n7495), .Q(
        g155), .QN(n7212) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n7308), .CLK(n7495), .Q(
        g153), .QN(n6826) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n7309), .CLK(n7496), .Q(
        g157), .QN(n7211) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n7309), .CLK(n7496), .Q(
        g158), .QN(n7210) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n7309), .CLK(n7496), .Q(
        g156), .QN(n6825) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n7309), .CLK(n7496), .Q(
        g160), .QN(n6787) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n7309), .CLK(n7496), .Q(
        g161), .QN(n6786) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n7310), .CLK(n7497), .Q(
        g159), .QN(n6785) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n7310), .CLK(n7497), .Q(
        test_so12) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n7309), .CLK(n7496), 
        .Q(g164), .QN(n6824) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n7309), .CLK(n7496), .Q(
        g162), .QN(n6823) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n7309), .CLK(n7496), .Q(
        g169), .QN(n6893) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n7309), .CLK(n7496), .Q(
        g170), .QN(n6892) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n7308), .CLK(n7495), .Q(
        g168), .QN(n6891) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n7308), .CLK(n7495), .Q(
        g172), .QN(n6890) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n7308), .CLK(n7495), .Q(
        g173), .QN(n6889) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n7308), .CLK(n7495), .Q(
        g171), .QN(n6888) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n7308), .CLK(n7495), .Q(
        g175), .QN(n6887) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n7308), .CLK(n7495), .Q(
        g176), .QN(n6886) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n7308), .CLK(n7495), .Q(
        g174), .QN(n6885) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n7309), .CLK(n7496), .Q(
        g178), .QN(n6884) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n7309), .CLK(n7496), .Q(
        g179), .QN(n6883) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n7309), .CLK(n7496), .Q(
        g177), .QN(n6882) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n7316), .CLK(n7503), .Q(
        g186) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n7317), .CLK(n7504), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n7317), .CLK(n7504), 
        .Q(g192) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n7317), .CLK(n7504), .Q(
        g231) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n7317), .CLK(n7504), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n7317), .CLK(n7504), .Q(
        g237) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n7317), .CLK(n7504), .Q(
        g195) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n7317), .CLK(n7504), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n7310), .CLK(n7497), .Q(
        g201) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n7310), .CLK(n7497), .Q(
        g240) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n7310), .CLK(n7497), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n7310), .CLK(n7497), .Q(
        g246) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n7310), .CLK(n7497), .Q(
        g204) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n7310), .CLK(n7497), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n7310), .CLK(n7497), .Q(
        g210) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n7310), .CLK(n7497), .Q(
        g249) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n7310), .CLK(n7497), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n7310), .CLK(n7497), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n7311), .CLK(n7498), 
        .Q(g213) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n7311), .CLK(n7498), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n7311), .CLK(n7498), .Q(
        g219) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n7311), .CLK(n7498), .Q(
        g258) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n7311), .CLK(n7498), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n7311), .CLK(n7498), .Q(
        g264) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n7311), .CLK(n7498), .Q(
        g222) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n7311), .CLK(n7498), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n7311), .CLK(n7498), .Q(
        g228) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n7311), .CLK(n7498), .Q(
        g267) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n7311), .CLK(n7498), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n7279), .CLK(n7466), .Q(
        g273) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n7282), .CLK(n7469), .Q(
        g92), .QN(n6994) );
  SDFFX1 DFF_237_Q_reg ( .D(g25932), .SI(g92), .SE(n7282), .CLK(n7469), .Q(g88), .QN(n6977) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n7282), .CLK(n7469), .Q(g83), .QN(n6993) );
  SDFFX1 DFF_239_Q_reg ( .D(g27120), .SI(g83), .SE(n7282), .CLK(n7469), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n7282), .CLK(n7469), 
        .Q(g74), .QN(n6992) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n7282), .CLK(n7469), .Q(g70), .QN(n6975) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n7282), .CLK(n7469), .Q(g65), .QN(n6991) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n7282), .CLK(n7469), .Q(g61), .QN(n6971) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n7282), .CLK(n7469), .Q(g56), .QN(n6600) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n7282), .CLK(n7469), .Q(g52), .QN(n6439) );
  SDFFX1 DFF_246_Q_reg ( .D(g13110), .SI(g52), .SE(n7279), .CLK(n7466), .Q(
        g180) );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n7279), .CLK(n7466), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n7279), .CLK(n7466), .Q(
        g181), .QN(n7001) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n7279), .CLK(n7466), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n7279), .CLK(n7466), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n7314), .CLK(n7501), .Q(
        g354), .QN(n6935) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n7315), .CLK(n7502), .Q(
        g343), .QN(n6934) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n7312), .CLK(n7499), .Q(
        test_so16) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n7314), .CLK(n7501), 
        .Q(g369), .QN(n6913) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n7314), .CLK(n7501), .Q(
        g358), .QN(n6912) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n7314), .CLK(n7501), .Q(
        g361), .QN(n6911) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n7314), .CLK(n7501), .Q(
        g384), .QN(n6654) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n7314), .CLK(n7501), .Q(
        g373), .QN(n6656) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n7314), .CLK(n7501), .Q(
        g376), .QN(n6655) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n7314), .CLK(n7501), .Q(
        g398), .QN(n6924) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n7314), .CLK(n7501), .Q(
        g388), .QN(n6923) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n7312), .CLK(n7499), .Q(
        g391), .QN(n6922) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n7312), .CLK(n7499), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n7313), .CLK(n7500), .Q(
        g411) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n7313), .CLK(n7500), .Q(
        g414) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n7313), .CLK(n7500), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n7313), .CLK(n7500), .Q(
        g420) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n7312), .CLK(n7499), .Q(
        g423) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n7312), .CLK(n7499), .Q(
        test_so17) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n7312), .CLK(n7499), 
        .Q(g428), .QN(n6967) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n7312), .CLK(n7499), .Q(
        g426), .QN(n6966) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n7312), .CLK(n7499), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n7312), .CLK(n7499), .Q(
        g432) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n7312), .CLK(n7499), .Q(
        g435) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n7313), .CLK(n7500), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n7313), .CLK(n7500), .Q(
        g441) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n7313), .CLK(n7500), .Q(
        g444) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n7313), .CLK(n7500), .Q(
        g448), .QN(n6965) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n7313), .CLK(n7500), .Q(
        g449), .QN(n6964) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n7313), .CLK(n7500), .Q(
        g447), .QN(n6963) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n7313), .CLK(n7500), .Q(
        g312), .QN(n6564) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n7313), .CLK(n7500), .Q(
        g313), .QN(n6563) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n7311), .CLK(n7498), .Q(
        g314), .QN(n6562) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n7312), .CLK(n7499), .Q(
        g315), .QN(n6561) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n7312), .CLK(n7499), .Q(
        test_so18) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n7279), .CLK(n7466), 
        .Q(g317), .QN(n6560) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n7279), .CLK(n7466), .Q(
        g318), .QN(n6559) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n7279), .CLK(n7466), .Q(
        g319), .QN(n6558) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n7279), .CLK(n7466), .Q(
        g320), .QN(n6557) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n7317), .CLK(n7504), .Q(
        g322), .QN(n6596) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n7317), .CLK(n7504), .Q(
        g323), .QN(n6595) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n7317), .CLK(n7504), .Q(
        g321), .QN(n6594) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n7317), .CLK(n7504), .Q(
        g403), .QN(n6962) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n7317), .CLK(n7504), .Q(
        g404), .QN(n6961) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n7318), .CLK(n7505), .Q(
        g402), .QN(n6960) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n7318), .CLK(n7505), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n7318), .CLK(n7505), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n7318), .CLK(n7505), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n7318), .CLK(n7505), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n7318), .CLK(n7505), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n7318), .CLK(n7505), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n7306), .CLK(n7493), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n7306), .CLK(n7493), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n7306), .CLK(n7493), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n7306), .CLK(n7493), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n7307), .CLK(n7494), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n7307), .CLK(n7494), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n7307), .CLK(n7494), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n7307), .CLK(n7494), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n7307), .CLK(n7494), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n7307), .CLK(n7494), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n7307), .CLK(n7494), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n7307), .CLK(n7494), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n7314), .CLK(n7501), .Q(
        n8056), .QN(n13234) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n7280), .CLK(n7467), .Q(
        g305), .QN(n6710) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n7280), .CLK(n7467), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n7314), .CLK(n7501), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n7314), .CLK(n7501), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n7315), .CLK(n7502), .Q(g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n7315), .CLK(n7502), .Q(g351) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n7315), .CLK(n7502), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n7315), .CLK(n7502), .Q(g353) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n7315), .CLK(n7502), .Q(g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n7315), .CLK(n7502), .Q(g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n7315), .CLK(n7502), .Q(g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n7315), .CLK(n7502), .Q(g366) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n7315), .CLK(n7502), .Q(g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n7315), .CLK(n7502), .Q(g368) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n7315), .CLK(n7502), .Q(g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n7316), .CLK(n7503), .Q(g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n7316), .CLK(n7503), .Q(g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n7316), .CLK(n7503), .Q(g381) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n7316), .CLK(n7503), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n7316), .CLK(n7503), .Q(g383) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n7316), .CLK(n7503), .Q(g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n7316), .CLK(n7503), .Q(g394) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n7316), .CLK(n7503), .Q(g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n7316), .CLK(n7503), .Q(g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n7316), .CLK(n7503), .Q(g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n7316), .CLK(n7503), .Q(g324) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n7325), .CLK(n7512), .Q(
        g5629) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n7325), .CLK(n7512), .Q(
        g5648) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n7325), .CLK(n7512), .Q(
        g337) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n7326), .CLK(n7513), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n7326), .CLK(n7513), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n7326), .CLK(n7513), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(g21842), .SI(g550), .SE(n7326), .CLK(n7513), .Q(
        g554), .QN(n7236) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n7326), .CLK(n7513), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n7326), .CLK(n7513), .Q(
        test_so22), .QN(n7271) );
  SDFFX1 DFF_362_Q_reg ( .D(n266), .SI(test_si23), .SE(n7326), .CLK(n7513), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n7326), .CLK(n7513), .Q(g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n7326), .CLK(n7513), .Q(g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n7326), .CLK(n7513), .Q(g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n7326), .CLK(n7513), .Q(g569) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n7327), .CLK(n7514), .Q(g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n7327), .CLK(n7514), .Q(g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n7327), .CLK(n7514), .Q(g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n7327), .CLK(n7514), .Q(g573) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n7327), .CLK(n7514), .Q(g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n7327), .CLK(n7514), .Q(g565) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n7327), .CLK(n7514), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n7327), .CLK(n7514), .Q(g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n7327), .CLK(n7514), .Q(g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n7327), .CLK(n7514), .Q(g489) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n7327), .CLK(n7514), .Q(
        test_so23), .QN(n7268) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n7327), .CLK(n7514), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n7328), .CLK(n7515), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n7328), .CLK(n7515), .Q(
        g486) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n7328), .CLK(n7515), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n7328), .CLK(n7515), .Q(
        g488) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n7328), .CLK(n7515), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n7328), .CLK(n7515), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n7328), .CLK(n7515), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n7328), .CLK(n7515), .Q(
        g477) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n7328), .CLK(n7515), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n7328), .CLK(n7515), .Q(
        g479) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n7328), .CLK(n7515), .Q(
        g480) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n7329), .CLK(n7516), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n7329), .CLK(n7516), .Q(
        g464) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n7329), .CLK(n7516), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n7329), .CLK(n7516), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n7328), .CLK(n7515), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n257), .SI(g471), .SE(n7329), .CLK(n7516), .Q(g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n7329), .CLK(n7516), .Q(g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n7329), .CLK(n7516), .Q(g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n7329), .CLK(n7516), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n7329), .CLK(n7516), .Q(g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n7330), .CLK(n7517), .Q(
        g548) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n7329), .CLK(n7516), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n7329), .CLK(n7516), .Q(g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n7329), .CLK(n7516), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n7330), .CLK(n7517), .Q(g559) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n7340), .CLK(n7527), .Q(
        g576), .QN(n6610) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n7340), .CLK(n7527), .Q(
        g577), .QN(n6612) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n7340), .CLK(n7527), .Q(
        g575), .QN(n6611) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n7340), .CLK(n7527), .Q(
        g579), .QN(n6622) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n7340), .CLK(n7527), .Q(
        test_so25) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n7340), .CLK(n7527), 
        .Q(g578), .QN(n6623) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n7340), .CLK(n7527), .Q(
        g582), .QN(n6447) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n7340), .CLK(n7527), .Q(
        g583), .QN(n6449) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n7340), .CLK(n7527), .Q(
        g581), .QN(n6448) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n7340), .CLK(n7527), .Q(
        g585), .QN(n6632) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n7340), .CLK(n7527), .Q(
        g586), .QN(n6634) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n7341), .CLK(n7528), .Q(
        g584), .QN(n6633) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n7341), .CLK(n7528), .Q(
        g587) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n7341), .CLK(n7528), .Q(
        g590) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n7341), .CLK(n7528), .Q(
        g593) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n7341), .CLK(n7528), .Q(
        g596) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n7341), .CLK(n7528), .Q(
        g599) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n7341), .CLK(n7528), .Q(
        g602) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n7341), .CLK(n7528), .Q(
        g614) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n7341), .CLK(n7528), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n7342), .CLK(n7529), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n7341), .CLK(n7528), 
        .Q(g605) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n7341), .CLK(n7528), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n7341), .CLK(n7528), .Q(
        g611) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n7343), .CLK(n7530), .Q(
        g490) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n7343), .CLK(n7530), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n7343), .CLK(n7530), .Q(
        g496) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n7343), .CLK(n7530), .Q(g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n7343), .CLK(n7530), .Q(
        n4571), .QN(n6681) );
  SDFFX1 DFF_442_Q_reg ( .D(n265), .SI(n4571), .SE(n7343), .CLK(n7530), .Q(
        g16297), .QN(n6682) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n7343), .CLK(n7530), .Q(
        g525), .QN(n7005) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n7343), .CLK(n7530), 
        .Q(n8047), .QN(DFF_444_n1) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n7343), .CLK(n7530), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n7343), .CLK(n7530), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n7343), .CLK(n7530), 
        .Q(n8044), .QN(DFF_447_n1) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n7343), .CLK(n7530), 
        .Q(n8043), .QN(DFF_448_n1) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n7344), .CLK(n7531), 
        .Q(test_so27), .QN(DFF_449_n1) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n7307), .CLK(
        n7494), .Q(g536), .QN(n6409) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n7307), .CLK(n7494), 
        .Q(g537), .QN(n6408) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n7280), .CLK(n7467), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n7307), .CLK(n7494), .Q(
        n8040), .QN(n13227) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n7321), .CLK(n7508), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n7321), .CLK(n7508), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n7326), .CLK(n7513), .Q(
        g630), .QN(n7044) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n7332), .CLK(n7519), .Q(
        g659) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n7332), .CLK(n7519), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(n7332), .CLK(n7519), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n7332), .CLK(n7519), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n7332), .CLK(n7519), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n7332), .CLK(n7519), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(n7332), .CLK(n7519), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n7332), .CLK(n7519), .Q(
        test_so28), .QN(n7270) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n7333), .CLK(n7520), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(g28199), .SI(g679), .SE(n7333), .CLK(n7520), .Q(
        g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n7333), .CLK(n7520), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n7333), .CLK(n7520), .Q(
        g699), .QN(n7123) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n7333), .CLK(n7520), .Q(
        g700), .QN(n7122) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n7333), .CLK(n7520), .Q(
        g698), .QN(n7161) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n7333), .CLK(n7520), .Q(
        g702), .QN(n7121) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n7333), .CLK(n7520), .Q(
        g703), .QN(n7120) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n7333), .CLK(n7520), .Q(
        g701), .QN(n7160) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n7333), .CLK(n7520), .Q(
        g705), .QN(n7119) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n7333), .CLK(n7520), .Q(
        g706), .QN(n7118) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n7333), .CLK(n7520), .Q(
        g704), .QN(n7159) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n7335), .CLK(n7522), .Q(
        g708), .QN(n7117) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n7335), .CLK(n7522), .Q(
        g709), .QN(n7116) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n7335), .CLK(n7522), .Q(
        g707), .QN(n7158) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n7335), .CLK(n7522), .Q(
        test_so29) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n7332), .CLK(n7519), 
        .Q(g712), .QN(n7115) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n7332), .CLK(n7519), .Q(
        g710), .QN(n7157) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n7334), .CLK(n7521), .Q(
        g714), .QN(n7114) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n7334), .CLK(n7521), .Q(
        g715), .QN(n7113) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n7334), .CLK(n7521), .Q(
        g713), .QN(n7156) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n7334), .CLK(n7521), .Q(
        g717), .QN(n7112) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n7334), .CLK(n7521), .Q(
        g718), .QN(n7111) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n7334), .CLK(n7521), .Q(
        g716), .QN(n7155) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n7334), .CLK(n7521), .Q(
        g720), .QN(n7110) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n7334), .CLK(n7521), .Q(
        g721), .QN(n7109) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n7334), .CLK(n7521), .Q(
        g719), .QN(n7154) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n7334), .CLK(n7521), .Q(
        g723), .QN(n7108) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n7334), .CLK(n7521), .Q(
        g724), .QN(n7107) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n7335), .CLK(n7522), .Q(
        g722), .QN(n7153) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n7335), .CLK(n7522), .Q(
        g726), .QN(n7106) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n7335), .CLK(n7522), .Q(
        test_so30) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n7334), .CLK(n7521), 
        .Q(g725), .QN(n7152) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n7342), .CLK(n7529), .Q(
        g729), .QN(n6847) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n7342), .CLK(n7529), .Q(
        g730) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n7342), .CLK(n7529), .Q(
        g728), .QN(n6901) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n7342), .CLK(n7529), .Q(
        g732), .QN(n6846) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n7342), .CLK(n7529), .Q(
        g733), .QN(n6838) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n7342), .CLK(n7529), .Q(
        g731), .QN(n6900) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n7342), .CLK(n7529), .Q(
        g735), .QN(n6774) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n7342), .CLK(n7529), .Q(
        g736), .QN(n6773) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n7342), .CLK(n7529), .Q(
        g734), .QN(n6778) );
  SDFFX1 DFF_508_Q_reg ( .D(g22218), .SI(g734), .SE(n7342), .CLK(n7529), .Q(
        g738), .QN(n7165) );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(n7342), .CLK(n7529), .Q(
        g739), .QN(n7229) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n7280), .CLK(n7467), .Q(
        g737), .QN(n7232) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n7280), .CLK(n7467), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n7280), .CLK(n7467), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n7280), .CLK(n7467), .Q(
        test_so31), .QN(n7267) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n7291), .CLK(n7478), 
        .Q(g818), .QN(n7209) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n7291), .CLK(n7478), .Q(
        g819), .QN(n7208) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n7291), .CLK(n7478), .Q(
        g817), .QN(n6822) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n7291), .CLK(n7478), .Q(
        g821), .QN(n7207) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n7291), .CLK(n7478), .Q(
        g822), .QN(n7206) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n7291), .CLK(n7478), .Q(
        g820), .QN(n6821) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n7291), .CLK(n7478), .Q(
        g830), .QN(n7205) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n7292), .CLK(n7479), .Q(
        g831), .QN(n7204) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n7292), .CLK(n7479), .Q(
        g829), .QN(n6820) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n7292), .CLK(n7479), .Q(
        g833), .QN(n7203) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n7292), .CLK(n7479), .Q(
        g834), .QN(n7202) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n7292), .CLK(n7479), .Q(
        g832), .QN(n6819) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n7292), .CLK(n7479), .Q(
        g836), .QN(n7201) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n7292), .CLK(n7479), .Q(
        g837), .QN(n7200) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n7292), .CLK(n7479), .Q(
        g835), .QN(n6818) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n7292), .CLK(n7479), .Q(
        test_so32) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n7290), .CLK(n7477), 
        .Q(g840), .QN(n7199) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n7290), .CLK(n7477), .Q(
        g838), .QN(n6817) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n7290), .CLK(n7477), .Q(
        g842), .QN(n7198) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n7290), .CLK(n7477), .Q(
        g843), .QN(n7197) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n7290), .CLK(n7477), .Q(
        g841), .QN(n6816) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n7288), .CLK(n7475), .Q(
        g845), .QN(n7196) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n7290), .CLK(n7477), .Q(
        g846), .QN(n7195) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n7290), .CLK(n7477), .Q(
        g844), .QN(n6815) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n7290), .CLK(n7477), .Q(
        g848), .QN(n6814) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n7290), .CLK(n7477), .Q(
        g849), .QN(n6813) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n7290), .CLK(n7477), .Q(
        g847), .QN(n6812) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n7291), .CLK(n7478), .Q(
        g851), .QN(n6811) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n7291), .CLK(n7478), .Q(
        g852), .QN(n6810) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n7291), .CLK(n7478), .Q(
        g850), .QN(n6809) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n7291), .CLK(n7478), .Q(
        g857), .QN(n6881) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n7291), .CLK(n7478), .Q(
        test_so33) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n7287), .CLK(n7474), 
        .Q(g856), .QN(n6880) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n7287), .CLK(n7474), .Q(
        g860), .QN(n6879) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n7287), .CLK(n7474), .Q(
        g861), .QN(n6878) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n7287), .CLK(n7474), .Q(
        g859), .QN(n6877) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n7287), .CLK(n7474), .Q(
        g863), .QN(n6876) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n7287), .CLK(n7474), .Q(
        g864), .QN(n6875) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n7287), .CLK(n7474), .Q(
        g862), .QN(n6874) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n7287), .CLK(n7474), .Q(
        g866), .QN(n6873) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n7287), .CLK(n7474), .Q(
        g867), .QN(n6872) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n7288), .CLK(n7475), .Q(
        g865), .QN(n6871) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n7297), .CLK(n7484), .Q(
        g873) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n7297), .CLK(n7484), .Q(
        g876) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n7297), .CLK(n7484), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n7297), .CLK(n7484), .Q(
        g918) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n7297), .CLK(n7484), .Q(
        g921) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n7297), .CLK(n7484), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n7292), .CLK(n7479), 
        .Q(g882) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n7292), .CLK(n7479), .Q(
        g885) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n7292), .CLK(n7479), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n7293), .CLK(n7480), .Q(
        g927) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n7293), .CLK(n7480), .Q(
        g930) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n7293), .CLK(n7480), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n7293), .CLK(n7480), .Q(
        g891) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n7293), .CLK(n7480), .Q(
        g894) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n7293), .CLK(n7480), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n7293), .CLK(n7480), .Q(
        g936) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n7293), .CLK(n7480), .Q(
        g939) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n7293), .CLK(n7480), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n7296), .CLK(n7483), .Q(
        g900) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n7296), .CLK(n7483), .Q(
        g903) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n7296), .CLK(n7483), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n7297), .CLK(n7484), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n7297), .CLK(n7484), 
        .Q(g948) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n7297), .CLK(n7484), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n7297), .CLK(n7484), .Q(
        g909) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n7297), .CLK(n7484), .Q(
        g912) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n7293), .CLK(n7480), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n7293), .CLK(n7480), .Q(
        g954) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n7293), .CLK(n7480), .Q(
        g957) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n7288), .CLK(n7475), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n7288), .CLK(n7475), .Q(
        g780), .QN(n6990) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n7288), .CLK(n7475), .Q(
        g776), .QN(n6978) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n7288), .CLK(n7475), .Q(
        g771), .QN(n6989) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n7288), .CLK(n7475), .Q(
        g767), .QN(n6435) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n7288), .CLK(n7475), .Q(
        g762), .QN(n6988) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n7288), .CLK(n7475), .Q(
        g758) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n7288), .CLK(n7475), .Q(
        g753), .QN(n6987) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n7289), .CLK(n7476), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n7289), .CLK(n7476), 
        .Q(g744), .QN(n6599) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n7289), .CLK(n7476), .Q(
        g740), .QN(n6438) );
  SDFFX1 DFF_596_Q_reg ( .D(g13110), .SI(g740), .SE(n7289), .CLK(n7476), .Q(
        g868) );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n7289), .CLK(n7476), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n7289), .CLK(n7476), .Q(
        g869), .QN(n7000) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n7289), .CLK(n7476), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n7289), .CLK(n7476), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n7289), .CLK(n7476), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n7289), .CLK(n7476), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n7296), .CLK(n7483), .Q(
        g1041), .QN(n6933) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n7296), .CLK(n7483), .Q(
        g1030), .QN(n6932) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n7296), .CLK(n7483), .Q(
        g1033), .QN(n6931) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n7296), .CLK(n7483), .Q(
        g1056), .QN(n6910) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n7296), .CLK(n7483), .Q(
        g1045), .QN(n6909) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n7296), .CLK(n7483), .Q(
        g1048), .QN(n6908) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n7296), .CLK(n7483), .Q(
        test_so37) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n7295), .CLK(n7482), 
        .Q(g1060), .QN(n6652) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n7295), .CLK(n7482), .Q(
        g1063), .QN(n6653) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n7296), .CLK(n7483), .Q(
        g1085), .QN(n6921) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n7296), .CLK(n7483), .Q(
        g1075), .QN(n6920) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n7294), .CLK(n7481), .Q(
        g1078), .QN(n6919) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n7294), .CLK(n7481), .Q(
        g1095) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n7295), .CLK(n7482), .Q(
        g1098) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n7295), .CLK(n7482), .Q(
        g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n7295), .CLK(n7482), .Q(
        g1104) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n7295), .CLK(n7482), .Q(
        g1107) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n7294), .CLK(n7481), .Q(
        g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n7294), .CLK(n7481), .Q(
        g1114), .QN(n6959) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n7294), .CLK(n7481), .Q(
        g1115), .QN(n6944) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n7294), .CLK(n7481), .Q(
        g1113), .QN(n6958) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n7294), .CLK(n7481), .Q(
        g1116) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n7294), .CLK(n7481), .Q(
        test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n7294), .CLK(n7481), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n7295), .CLK(n7482), .Q(
        g1125) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n7295), .CLK(n7482), .Q(
        g1128) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n7295), .CLK(n7482), .Q(
        g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n7295), .CLK(n7482), .Q(
        g1135), .QN(n6957) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n7295), .CLK(n7482), .Q(
        g1136), .QN(n6943) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n7294), .CLK(n7481), .Q(
        g1134), .QN(n6956) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n7294), .CLK(n7481), .Q(
        g999), .QN(n6556) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n7295), .CLK(n7482), .Q(
        g1000), .QN(n6539) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n7294), .CLK(n7481), .Q(
        g1001), .QN(n6555) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n7288), .CLK(n7475), .Q(
        g1002), .QN(n6554) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n7290), .CLK(n7477), .Q(
        g1003), .QN(n6538) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n7290), .CLK(n7477), .Q(
        g1004), .QN(n6553) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n7288), .CLK(n7475), .Q(
        g1005), .QN(n6552) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n7289), .CLK(n7476), .Q(
        g1006), .QN(n6537) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n7289), .CLK(n7476), .Q(
        test_so39) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n7297), .CLK(n7484), 
        .Q(g1009), .QN(n6593) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n7298), .CLK(n7485), .Q(
        g1010), .QN(n6587) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n7298), .CLK(n7485), .Q(
        g1008), .QN(n6592) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n7298), .CLK(n7485), .Q(
        g1090), .QN(n6955) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n7298), .CLK(n7485), .Q(
        g1091), .QN(n6942) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n7298), .CLK(n7485), .Q(
        g1089), .QN(n6954) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n7298), .CLK(n7485), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n7298), .CLK(n7485), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n7298), .CLK(n7485), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n7298), .CLK(n7485), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n7298), .CLK(n7485), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n7298), .CLK(n7485), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n7298), .CLK(n7485), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n7299), .CLK(n7486), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n7299), .CLK(n7486), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n7299), .CLK(n7486), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n7286), .CLK(n7473), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n7286), .CLK(n7473), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n7286), .CLK(n7473), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n7287), .CLK(n7474), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n7287), .CLK(n7474), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n7287), .CLK(n7474), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n7299), .CLK(n7486), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n7299), .CLK(n7486), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n7299), .CLK(n7486), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(g26183), .SI(g986), .SE(n7299), .CLK(n7486), .Q(
        g992), .QN(n6997) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n7299), .CLK(n7486), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n7299), .CLK(n7486), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n7299), .CLK(n7486), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n7300), .CLK(n7487), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n7300), .CLK(n7487), .Q(
        g1038) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n7300), .CLK(n7487), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n7300), .CLK(n7487), .Q(g1040) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n7300), .CLK(n7487), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n7300), .CLK(n7487), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n7300), .CLK(n7487), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n7300), .CLK(n7487), .Q(
        g1053) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n7300), .CLK(n7487), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n7300), .CLK(n7487), .Q(
        g1055) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n7300), .CLK(n7487), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n7300), .CLK(n7487), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n7301), .CLK(n7488), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n7301), .CLK(n7488), .Q(
        g1068) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n7301), .CLK(n7488), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n7301), .CLK(n7488), .Q(
        g1070) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n7301), .CLK(n7488), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n7301), .CLK(n7488), .Q(
        g1081) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n7301), .CLK(n7488), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n7301), .CLK(n7488), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n7301), .CLK(n7488), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n7301), .CLK(n7488), .Q(
        g1011) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n7321), .CLK(n7508), .Q(
        g5657) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n7321), .CLK(n7508), .Q(
        g5686) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n7321), .CLK(n7508), .Q(
        g1024) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n7322), .CLK(n7509), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n7322), .CLK(n7509), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n7322), .CLK(n7509), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(g21843), .SI(g1236), .SE(n7322), .CLK(n7509), .Q(
        g1240), .QN(n7235) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n7322), .CLK(n7509), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n7322), .CLK(n7509), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n433), .SI(g1196), .SE(n7322), .CLK(n7509), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n7322), .CLK(n7509), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n7322), .CLK(n7509), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n7322), .CLK(n7509), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n7322), .CLK(n7509), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n7323), .CLK(n7510), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n7323), .CLK(n7510), .Q(
        g1257) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n7323), .CLK(n7510), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n7323), .CLK(n7510), .Q(
        g1259) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n7323), .CLK(n7510), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n7323), .CLK(n7510), .Q(
        g1251) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n7323), .CLK(n7510), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n7323), .CLK(n7510), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n7323), .CLK(n7510), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n7323), .CLK(n7510), .Q(
        g1176) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n7323), .CLK(n7510), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n7323), .CLK(n7510), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n7324), .CLK(n7511), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n7324), .CLK(n7511), .Q(
        g1173) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n7324), .CLK(n7511), .Q(
        test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n7324), .CLK(n7511), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n7324), .CLK(n7511), .Q(
        g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n7324), .CLK(n7511), .Q(
        g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n7324), .CLK(n7511), .Q(
        g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n7324), .CLK(n7511), .Q(
        g1164) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n7324), .CLK(n7511), .Q(
        g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n7324), .CLK(n7511), .Q(
        g1166) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n7324), .CLK(n7511), .Q(
        g1167) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n7324), .CLK(n7511), .Q(
        g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n7325), .CLK(n7512), .Q(
        g1151) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n7325), .CLK(n7512), .Q(
        g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n7325), .CLK(n7512), .Q(
        g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n7325), .CLK(n7512), .Q(
        g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n440), .SI(g1158), .SE(n7325), .CLK(n7512), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n7325), .CLK(n7512), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n7325), .CLK(n7512), .Q(
        test_so45) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n7325), .CLK(n7512), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n7325), .CLK(n7512), .Q(
        n4549), .QN(n6407) );
  SDFFX1 DFF_750_Q_reg ( .D(n7265), .SI(n4549), .SE(n7330), .CLK(n7517), .Q(
        n4361) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n7330), .CLK(n7517), .Q(
        g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n7330), .CLK(n7517), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n7330), .CLK(n7517), .Q(
        g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n7330), .CLK(n7517), .Q(
        g1245) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n7344), .CLK(n7531), .Q(
        g1262), .QN(n6607) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n7344), .CLK(n7531), .Q(
        g1263), .QN(n6609) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n7344), .CLK(n7531), .Q(
        g1261), .QN(n6608) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n7344), .CLK(n7531), .Q(
        g1265), .QN(n6619) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n7344), .CLK(n7531), .Q(
        g1266), .QN(n6621) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n7344), .CLK(n7531), .Q(
        g1264), .QN(n6620) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n7344), .CLK(n7531), .Q(
        g1268), .QN(n6445) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n7344), .CLK(n7531), .Q(
        g1269), .QN(n6446) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n7344), .CLK(n7531), .Q(
        test_so46) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n7344), .CLK(n7531), 
        .Q(g1271), .QN(n6629) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n7344), .CLK(n7531), .Q(
        g1272), .QN(n6631) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n7345), .CLK(n7532), .Q(
        g1270), .QN(n6630) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n7345), .CLK(n7532), .Q(
        g1273) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n7345), .CLK(n7532), .Q(
        g1276) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n7345), .CLK(n7532), .Q(
        g1279) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n7345), .CLK(n7532), .Q(
        g1282) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n7345), .CLK(n7532), .Q(
        g1285) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n7345), .CLK(n7532), .Q(
        g1288) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n7345), .CLK(n7532), .Q(
        g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n7345), .CLK(n7532), .Q(
        g1303) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n7345), .CLK(n7532), .Q(
        g1306) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n7345), .CLK(n7532), .Q(
        g1291) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n7346), .CLK(n7533), .Q(
        g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n7346), .CLK(n7533), .Q(
        g1297) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n7346), .CLK(n7533), .Q(
        test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n7346), .CLK(n7533), 
        .Q(g1180) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n7346), .CLK(n7533), .Q(
        g1183) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n7346), .CLK(n7533), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n7346), .CLK(n7533), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n264), .SI(n8009), .SE(n7346), .CLK(n7533), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n7346), .CLK(n7533), .Q(
        g1211), .QN(n7004) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n7346), .CLK(n7533), 
        .Q(n8008), .QN(DFF_794_n1) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n7347), .CLK(n7534), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n7347), .CLK(n7534), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n7347), .CLK(n7534), 
        .Q(n8005), .QN(DFF_797_n1) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n7347), .CLK(n7534), 
        .Q(n8004), .QN(DFF_798_n1) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n7347), .CLK(n7534), 
        .Q(n8003), .QN(DFF_799_n1) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n7347), .CLK(n7534), 
        .Q(g1222), .QN(n6415) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n7347), .CLK(n7534), 
        .Q(g1223), .QN(n6414) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n7347), .CLK(n7534), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n7347), .CLK(n7534), .Q(
        test_so48), .QN(n13230) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n7321), .CLK(n7508), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n7321), .CLK(n7508), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n7322), .CLK(n7509), .Q(
        g1316), .QN(n7043) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n7335), .CLK(n7522), .Q(
        g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n7335), .CLK(n7522), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(n7335), .CLK(n7522), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n7335), .CLK(n7522), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n7335), .CLK(n7522), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n7336), .CLK(n7523), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(n7336), .CLK(n7523), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n7336), .CLK(n7523), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n7336), .CLK(n7523), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n7336), .CLK(n7523), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n7336), .CLK(n7523), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n7347), .CLK(n7534), .Q(
        test_so49) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n7348), .CLK(n7535), 
        .Q(g1386), .QN(n7105) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n7348), .CLK(n7535), .Q(
        g1384), .QN(n7151) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n7348), .CLK(n7535), .Q(
        g1388), .QN(n7104) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n7348), .CLK(n7535), .Q(
        g1389), .QN(n7103) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n7348), .CLK(n7535), .Q(
        g1387), .QN(n7150) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n7348), .CLK(n7535), .Q(
        g1391), .QN(n7102) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n7348), .CLK(n7535), .Q(
        g1392), .QN(n7101) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n7348), .CLK(n7535), .Q(
        g1390), .QN(n7149) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n7348), .CLK(n7535), .Q(
        g1394), .QN(n7100) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n7348), .CLK(n7535), .Q(
        g1395), .QN(n7099) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n7348), .CLK(n7535), .Q(
        g1393), .QN(n7148) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n7348), .CLK(n7535), .Q(
        g1397), .QN(n7098) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n7349), .CLK(n7536), .Q(
        g1398), .QN(n7097) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n7349), .CLK(n7536), .Q(
        g1396), .QN(n7147) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n7349), .CLK(n7536), .Q(
        g1400), .QN(n7096) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n7350), .CLK(n7537), .Q(
        test_so50) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n7347), .CLK(n7534), 
        .Q(g1399), .QN(n7146) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n7347), .CLK(n7534), .Q(
        g1403), .QN(n7095) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n7349), .CLK(n7536), .Q(
        g1404), .QN(n7094) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n7349), .CLK(n7536), .Q(
        g1402), .QN(n7145) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n7349), .CLK(n7536), .Q(
        g1406), .QN(n7093) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n7349), .CLK(n7536), .Q(
        g1407), .QN(n7092) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n7349), .CLK(n7536), .Q(
        g1405), .QN(n7144) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n7349), .CLK(n7536), .Q(
        g1409), .QN(n7091) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n7349), .CLK(n7536), .Q(
        g1410), .QN(n7090) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n7349), .CLK(n7536), .Q(
        g1408), .QN(n7143) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n7349), .CLK(n7536), .Q(
        g1412), .QN(n7089) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n7350), .CLK(n7537), .Q(
        g1413), .QN(n7088) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n7350), .CLK(n7537), .Q(
        g1411), .QN(n7142) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n7350), .CLK(n7537), .Q(
        g1415), .QN(n6845) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n7350), .CLK(n7537), .Q(
        g1416), .QN(n6837) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n7350), .CLK(n7537), .Q(
        test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n7345), .CLK(n7532), 
        .Q(g1418), .QN(n6844) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n7346), .CLK(n7533), .Q(
        g1419), .QN(n6836) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n7346), .CLK(n7533), .Q(
        g1417), .QN(n6899) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n7350), .CLK(n7537), .Q(
        g1421), .QN(n6772) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n7350), .CLK(n7537), .Q(
        g1422), .QN(n6771) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n7350), .CLK(n7537), .Q(
        g1420), .QN(n6777) );
  SDFFX1 DFF_858_Q_reg ( .D(g22234), .SI(g1420), .SE(n7350), .CLK(n7537), .Q(
        g1424), .QN(n7164) );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(n7350), .CLK(n7537), .Q(
        g1425), .QN(n7228) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n7350), .CLK(n7537), .Q(
        g1423), .QN(n7231) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n7351), .CLK(n7538), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n7351), .CLK(n7538), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n7351), .CLK(n7538), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n7352), .CLK(n7539), .Q(
        g1512), .QN(n7194) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n7353), .CLK(n7540), .Q(
        g1513), .QN(n7193) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n7353), .CLK(n7540), .Q(
        g1511), .QN(n6808) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n7353), .CLK(n7540), .Q(
        test_so52) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n7354), .CLK(n7541), 
        .Q(g1516), .QN(n7192) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n7354), .CLK(n7541), .Q(
        g1514), .QN(n6807) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n7354), .CLK(n7541), .Q(
        g1524), .QN(n7191) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n7354), .CLK(n7541), .Q(
        g1525), .QN(n7190) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n7354), .CLK(n7541), .Q(
        g1523), .QN(n6806) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n7354), .CLK(n7541), .Q(
        g1527), .QN(n7189) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n7354), .CLK(n7541), .Q(
        g1528), .QN(n7188) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n7354), .CLK(n7541), .Q(
        g1526), .QN(n6805) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n7354), .CLK(n7541), .Q(
        g1530), .QN(n7187) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n7355), .CLK(n7542), .Q(
        g1531), .QN(n7186) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n7355), .CLK(n7542), .Q(
        g1529), .QN(n6804) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n7355), .CLK(n7542), .Q(
        g1533), .QN(n7185) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n7355), .CLK(n7542), .Q(
        g1534), .QN(n7184) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n7355), .CLK(n7542), .Q(
        g1532), .QN(n6803) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n7355), .CLK(n7542), .Q(
        g1536), .QN(n7183) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n7355), .CLK(n7542), .Q(
        test_so53) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n7351), .CLK(n7538), 
        .Q(g1535), .QN(n6802) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n7352), .CLK(n7539), .Q(
        g1539), .QN(n7182) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n7352), .CLK(n7539), .Q(
        g1540), .QN(n7181) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n7352), .CLK(n7539), .Q(
        g1538), .QN(n6801) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n7353), .CLK(n7540), .Q(
        g1542), .QN(n6784) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n7353), .CLK(n7540), .Q(
        g1543), .QN(n6783) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n7353), .CLK(n7540), .Q(
        g1541), .QN(n6782) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n7354), .CLK(n7541), .Q(
        g1545), .QN(n6800) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n7353), .CLK(n7540), .Q(
        g1546), .QN(n6799) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n7353), .CLK(n7540), .Q(
        g1544), .QN(n6798) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n7353), .CLK(n7540), .Q(
        g1551), .QN(n6870) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n7353), .CLK(n7540), .Q(
        g1552), .QN(n6869) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n7353), .CLK(n7540), .Q(
        g1550), .QN(n6868) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n7353), .CLK(n7540), .Q(
        g1554), .QN(n6867) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n7354), .CLK(n7541), .Q(
        g1555), .QN(n6866) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n7354), .CLK(n7541), .Q(
        test_so54) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n7351), .CLK(n7538), 
        .Q(g1557), .QN(n6865) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n7351), .CLK(n7538), .Q(
        g1558), .QN(n6864) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n7351), .CLK(n7538), .Q(
        g1556), .QN(n6863) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n7351), .CLK(n7538), .Q(
        g1560), .QN(n6862) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n7351), .CLK(n7538), .Q(
        g1561), .QN(n6861) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n7351), .CLK(n7538), .Q(
        g1559), .QN(n6860) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n7362), .CLK(n7549), .Q(
        g1567) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n7362), .CLK(n7549), .Q(
        g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n7362), .CLK(n7549), .Q(
        g1573) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n7362), .CLK(n7549), .Q(
        g1612) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n7362), .CLK(n7549), .Q(
        g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n7362), .CLK(n7549), .Q(
        g1618) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n7362), .CLK(n7549), .Q(
        g1576) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n7363), .CLK(n7550), .Q(
        g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n7356), .CLK(n7543), .Q(
        g1582) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n7356), .CLK(n7543), .Q(
        test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n7356), .CLK(n7543), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n7356), .CLK(n7543), .Q(
        g1627) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n7356), .CLK(n7543), .Q(
        g1585) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n7357), .CLK(n7544), .Q(
        g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n7357), .CLK(n7544), .Q(
        g1591) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n7357), .CLK(n7544), .Q(
        g1630) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n7357), .CLK(n7544), .Q(
        g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n7357), .CLK(n7544), .Q(
        g1636) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n7362), .CLK(n7549), .Q(
        g1594) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n7362), .CLK(n7549), .Q(
        g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n7362), .CLK(n7549), .Q(
        g1600) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n7363), .CLK(n7550), .Q(
        g1639) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n7363), .CLK(n7550), .Q(
        g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n7363), .CLK(n7550), .Q(
        g1645) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n7363), .CLK(n7550), .Q(
        g1603) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n7363), .CLK(n7550), .Q(
        test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n7357), .CLK(n7544), 
        .Q(g1609) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n7357), .CLK(n7544), .Q(
        g1648) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n7357), .CLK(n7544), .Q(
        g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n7355), .CLK(n7542), .Q(
        g1654) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n7356), .CLK(n7543), .Q(
        g1466), .QN(n6986) );
  SDFFX1 DFF_937_Q_reg ( .D(g25938), .SI(g1466), .SE(n7356), .CLK(n7543), .Q(
        g1462), .QN(n6976) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n7356), .CLK(n7543), .Q(
        g1457), .QN(n6985) );
  SDFFX1 DFF_939_Q_reg ( .D(g27129), .SI(g1457), .SE(n7356), .CLK(n7543), .Q(
        g1453), .QN(n6434) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n7356), .CLK(n7543), .Q(
        g1448), .QN(n6984) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n7356), .CLK(n7543), .Q(
        g1444), .QN(n6973) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n7356), .CLK(n7543), .Q(
        g1439), .QN(n6983) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n7351), .CLK(n7538), .Q(
        g1435), .QN(n6970) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n7351), .CLK(n7538), .Q(
        g1430), .QN(n6598) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n7352), .CLK(n7539), .Q(
        g1426), .QN(n6437) );
  SDFFX1 DFF_946_Q_reg ( .D(g13110), .SI(g1426), .SE(n7352), .CLK(n7539), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n7352), .CLK(n7539), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n7352), .CLK(n7539), .Q(g1563), .QN(n6999) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n7352), .CLK(n7539), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n7352), .CLK(n7539), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n7360), .CLK(n7547), .Q(
        g1735), .QN(n6930) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n7360), .CLK(n7547), .Q(
        g1724), .QN(n6929) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n7360), .CLK(n7547), .Q(
        g1727), .QN(n6928) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n7360), .CLK(n7547), .Q(
        g1750), .QN(n6907) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n7360), .CLK(n7547), .Q(
        g1739), .QN(n6906) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n7359), .CLK(n7546), .Q(
        g1742), .QN(n6905) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n7359), .CLK(n7546), .Q(
        g1765), .QN(n6649) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n7360), .CLK(n7547), .Q(
        g1754), .QN(n6651) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n7359), .CLK(n7546), .Q(
        g1757), .QN(n6650) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n7360), .CLK(n7547), .Q(
        g1779), .QN(n6918) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n7360), .CLK(n7547), .Q(
        test_so58) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n7357), .CLK(n7544), 
        .Q(g1772), .QN(n6917) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n7358), .CLK(n7545), .Q(
        g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n7359), .CLK(n7546), .Q(
        g1792) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n7359), .CLK(n7546), .Q(
        g1795) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n7359), .CLK(n7546), .Q(
        g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n7359), .CLK(n7546), .Q(
        g1801) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n7358), .CLK(n7545), .Q(
        g1804) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n7358), .CLK(n7545), .Q(
        g1808), .QN(n6953) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n7358), .CLK(n7545), .Q(
        g1809), .QN(n6941) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n7358), .CLK(n7545), .Q(
        g1807), .QN(n6952) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n7358), .CLK(n7545), .Q(
        g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n7358), .CLK(n7545), .Q(
        g1813) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n7358), .CLK(n7545), .Q(
        g1816) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n7359), .CLK(n7546), .Q(
        g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n7359), .CLK(n7546), .Q(
        g1822) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n7359), .CLK(n7546), .Q(
        test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n7358), .CLK(n7545), 
        .Q(g1829), .QN(n6951) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n7359), .CLK(n7546), .Q(
        g1830), .QN(n6940) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n7358), .CLK(n7545), .Q(
        g1828), .QN(n6950) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n7358), .CLK(n7545), .Q(
        g1693), .QN(n6551) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n7358), .CLK(n7545), .Q(
        g1694), .QN(n6536) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n7357), .CLK(n7544), .Q(
        g1695), .QN(n6550) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n7357), .CLK(n7544), .Q(
        g1696), .QN(n6549) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n7357), .CLK(n7544), .Q(
        g1697), .QN(n6535) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n7355), .CLK(n7542), .Q(
        g1698), .QN(n6548) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n7355), .CLK(n7542), .Q(
        g1699), .QN(n6547) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n7355), .CLK(n7542), .Q(
        g1700), .QN(n6534) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n7355), .CLK(n7542), .Q(
        g1701), .QN(n6546) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n7363), .CLK(n7550), .Q(
        g1703), .QN(n6591) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n7363), .CLK(n7550), .Q(
        g1704), .QN(n6586) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n7360), .CLK(n7547), .Q(
        g1702), .QN(n6590) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n7360), .CLK(n7547), .Q(
        test_so60) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n7360), .CLK(n7547), 
        .Q(g1785), .QN(n6939) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n7360), .CLK(n7547), .Q(
        g1783), .QN(n6949) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n7361), .CLK(n7548), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n7361), .CLK(n7548), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n7361), .CLK(n7548), .Q(
        g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n7361), .CLK(n7548), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n7361), .CLK(n7548), .Q(
        g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n7361), .CLK(n7548), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n7361), .CLK(n7548), .Q(
        g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n7361), .CLK(n7548), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n7361), .CLK(n7548), .Q(
        g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n7361), .CLK(n7548), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n7361), .CLK(n7548), .Q(
        g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n7361), .CLK(n7548), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n7362), .CLK(n7549), .Q(
        g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n7362), .CLK(n7549), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n7277), .CLK(n7464), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n7277), .CLK(n7464), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n7285), .CLK(n7472), .Q(
        g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n7285), .CLK(n7472), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n7359), .CLK(n7546), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(g28903), .SI(g1680), .SE(n7363), .CLK(n7550), .Q(
        g1686) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n7363), .CLK(n7550), .Q(
        n7978) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n7363), .CLK(n7550), .Q(
        g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n7363), .CLK(n7550), .Q(
        g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n7364), .CLK(n7551), .Q(
        g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n7364), .CLK(n7551), .Q(
        g1732) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n7364), .CLK(n7551), .Q(
        g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n7364), .CLK(n7551), .Q(
        g1734) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n7364), .CLK(n7551), .Q(
        g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n7364), .CLK(n7551), .Q(
        g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n7364), .CLK(n7551), .Q(
        test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n7364), .CLK(
        n7551), .Q(g1747) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n7364), .CLK(n7551), .Q(
        g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n7364), .CLK(n7551), .Q(
        g1749) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n7364), .CLK(n7551), .Q(
        g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n7364), .CLK(n7551), .Q(
        g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n7365), .CLK(n7552), .Q(
        g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n7365), .CLK(n7552), .Q(
        g1762) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n7365), .CLK(n7552), .Q(
        g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n7365), .CLK(n7552), .Q(
        g1764) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n7365), .CLK(n7552), .Q(
        g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n7365), .CLK(n7552), .Q(
        g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n7365), .CLK(n7552), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n7365), .CLK(n7552), .Q(
        g1777) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n7365), .CLK(n7552), .Q(
        g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n7365), .CLK(n7552), .Q(
        g1705) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n7365), .CLK(n7552), .Q(
        test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n7365), .CLK(
        n7552), .Q(g5738) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n7366), .CLK(n7553), .Q(
        g1718) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n7366), .CLK(n7553), .Q(
        g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n7366), .CLK(n7553), .Q(
        g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n7366), .CLK(n7553), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(g21845), .SI(g1930), .SE(n7366), .CLK(n7553), .Q(
        g1934), .QN(n7234) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n7366), .CLK(n7553), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n7366), .CLK(n7553), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n605), .SI(g1890), .SE(n7367), .CLK(n7554), .Q(
        g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n7367), .CLK(n7554), .Q(
        g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n7367), .CLK(n7554), .Q(
        g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n7367), .CLK(n7554), .Q(
        g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n7367), .CLK(n7554), .Q(
        g1949) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n7368), .CLK(n7555), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n7368), .CLK(n7555), .Q(
        g1951) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n7368), .CLK(n7555), .Q(
        test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n7368), .CLK(
        n7555), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n7368), .CLK(n7555), .Q(
        g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n7368), .CLK(n7555), .Q(
        g1945) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n7368), .CLK(n7555), .Q(
        g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n7368), .CLK(n7555), .Q(
        g1947) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n7368), .CLK(n7555), .Q(
        g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n7368), .CLK(n7555), .Q(
        g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n7368), .CLK(n7555), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n7368), .CLK(n7555), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n7369), .CLK(n7556), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n7369), .CLK(n7556), .Q(
        g1867) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n7369), .CLK(n7556), .Q(
        g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n7369), .CLK(n7556), .Q(
        g1869) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n7369), .CLK(n7556), .Q(
        g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n7369), .CLK(n7556), .Q(
        test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n7369), .CLK(n7556), 
        .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n7369), .CLK(n7556), .Q(
        g1858) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n7369), .CLK(n7556), .Q(
        g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n7369), .CLK(n7556), .Q(
        g1860) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n7369), .CLK(n7556), .Q(
        g1861) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n7369), .CLK(n7556), .Q(
        g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n7370), .CLK(n7557), .Q(
        g1845) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n7370), .CLK(n7557), .Q(
        g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n7370), .CLK(n7557), .Q(
        g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n7370), .CLK(n7557), .Q(
        g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n598), .SI(g1852), .SE(n7370), .CLK(n7557), .Q(
        g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n7370), .CLK(n7557), .Q(
        g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n7370), .CLK(n7557), .Q(
        g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n7370), .CLK(n7557), .Q(
        g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n7370), .CLK(n7557), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n7264), .SI(test_si67), .SE(n7371), .CLK(n7558), 
        .Q(n7971) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n7370), .CLK(n7557), .Q(
        g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n7370), .CLK(n7557), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n7370), .CLK(n7557), .Q(
        g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n7371), .CLK(n7558), .Q(
        g1939) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n7372), .CLK(n7559), .Q(
        g1956), .QN(n6604) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n7372), .CLK(n7559), .Q(
        g1957), .QN(n6606) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n7372), .CLK(n7559), .Q(
        g1955), .QN(n6605) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n7372), .CLK(n7559), .Q(
        g1959), .QN(n6616) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n7372), .CLK(n7559), .Q(
        g1960), .QN(n6618) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n7371), .CLK(n7558), .Q(
        g1958), .QN(n6617) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n7371), .CLK(n7558), .Q(
        g1962), .QN(n6442) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n7372), .CLK(n7559), .Q(
        g1963), .QN(n6444) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n7371), .CLK(n7558), .Q(
        g1961), .QN(n6443) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n7371), .CLK(n7558), .Q(
        test_so67) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n7372), .CLK(n7559), 
        .Q(g1966), .QN(n6628) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n7372), .CLK(n7559), .Q(
        g1964), .QN(n6627) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n7372), .CLK(n7559), .Q(
        g1967) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n7372), .CLK(n7559), .Q(
        g1970) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n7372), .CLK(n7559), .Q(
        g1973) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n7372), .CLK(n7559), .Q(
        g1976) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n7373), .CLK(n7560), .Q(
        g1979) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n7373), .CLK(n7560), .Q(
        g1982) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n7373), .CLK(n7560), .Q(
        g1994) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n7373), .CLK(n7560), .Q(
        g1997) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n7373), .CLK(n7560), .Q(
        g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n7373), .CLK(n7560), .Q(
        g1985) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n7373), .CLK(n7560), .Q(
        g1988) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n7373), .CLK(n7560), .Q(
        g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n7373), .CLK(n7560), .Q(
        test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n7373), .CLK(n7560), 
        .Q(g1874) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n7373), .CLK(n7560), .Q(
        g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n7373), .CLK(n7560), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n7374), .CLK(n7561), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(g28990), .SI(n7968), .SE(n7374), .CLK(n7561), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n7374), .CLK(n7561), 
        .Q(g1905), .QN(n7003) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n7374), .CLK(n7561), 
        .Q(n7967), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n7374), .CLK(n7561), 
        .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n7374), .CLK(n7561), 
        .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n7374), .CLK(n7561), 
        .Q(n7964), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n7374), .CLK(n7561), 
        .Q(n7963), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n7374), .CLK(n7561), 
        .Q(n7962), .QN(DFF_1149_n1) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n7374), .CLK(n7561), 
        .Q(g1916), .QN(n6413) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n7374), .CLK(n7561), 
        .Q(g1917), .QN(n6412) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n7374), .CLK(n7561), .Q(
        test_so69) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n7285), .CLK(n7472), 
        .Q(n7960), .QN(n13229) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n7321), .CLK(n7508), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n7321), .CLK(n7508), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n7366), .CLK(n7553), .Q(
        g2010), .QN(n7042) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n7366), .CLK(n7553), .Q(
        g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n7366), .CLK(n7553), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(n7366), .CLK(n7553), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n7366), .CLK(n7553), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n7367), .CLK(n7554), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n7367), .CLK(n7554), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(n7367), .CLK(n7554), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n7367), .CLK(n7554), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n7367), .CLK(n7554), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n7367), .CLK(n7554), .Q(
        test_so70), .QN(n7272) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n7367), .CLK(n7554), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n7375), .CLK(n7562), .Q(
        g2079), .QN(n7087) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n7375), .CLK(n7562), .Q(
        g2080), .QN(n7086) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n7375), .CLK(n7562), .Q(
        g2078), .QN(n7141) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n7375), .CLK(n7562), .Q(
        g2082), .QN(n7085) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n7375), .CLK(n7562), .Q(
        g2083), .QN(n7084) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n7376), .CLK(n7563), .Q(
        g2081), .QN(n7140) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n7376), .CLK(n7563), .Q(
        g2085), .QN(n7083) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n7376), .CLK(n7563), .Q(
        g2086), .QN(n7082) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n7376), .CLK(n7563), .Q(
        g2084), .QN(n7139) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n7376), .CLK(n7563), .Q(
        g2088), .QN(n7081) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n7376), .CLK(n7563), .Q(
        g2089), .QN(n7080) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n7376), .CLK(n7563), .Q(
        g2087), .QN(n7138) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n7376), .CLK(n7563), .Q(
        g2091), .QN(n7079) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n7376), .CLK(n7563), .Q(
        test_so71) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n7376), .CLK(n7563), 
        .Q(g2090), .QN(n7137) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n7376), .CLK(n7563), .Q(
        g2094), .QN(n7078) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n7376), .CLK(n7563), .Q(
        g2095), .QN(n7077) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n7377), .CLK(n7564), .Q(
        g2093), .QN(n7136) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n7377), .CLK(n7564), .Q(
        g2097), .QN(n7076) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n7377), .CLK(n7564), .Q(
        g2098), .QN(n7075) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n7377), .CLK(n7564), .Q(
        g2096), .QN(n7135) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n7377), .CLK(n7564), .Q(
        g2100), .QN(n7074) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n7377), .CLK(n7564), .Q(
        g2101), .QN(n7073) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n7377), .CLK(n7564), .Q(
        g2099), .QN(n7134) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n7377), .CLK(n7564), .Q(
        g2103), .QN(n7072) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n7377), .CLK(n7564), .Q(
        g2104), .QN(n7071) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n7377), .CLK(n7564), .Q(
        g2102), .QN(n7133) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n7377), .CLK(n7564), .Q(
        g2106), .QN(n7070) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n7377), .CLK(n7564), .Q(
        test_so72) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n7375), .CLK(n7562), 
        .Q(g2105), .QN(n7132) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n7375), .CLK(n7562), .Q(
        g2109), .QN(n6843) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n7375), .CLK(n7562), .Q(
        g2110) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n7375), .CLK(n7562), .Q(
        g2108), .QN(n6898) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n7375), .CLK(n7562), .Q(
        g2112), .QN(n6842) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n7375), .CLK(n7562), .Q(
        g2113), .QN(n6834) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n7375), .CLK(n7562), .Q(
        g2111), .QN(n6897) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n7378), .CLK(n7565), .Q(
        g2115), .QN(n6770) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n7378), .CLK(n7565), .Q(
        g2116), .QN(n6769) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n7378), .CLK(n7565), .Q(
        g2114), .QN(n6776) );
  SDFFX1 DFF_1208_Q_reg ( .D(g22249), .SI(g2114), .SE(n7378), .CLK(n7565), .Q(
        g2118), .QN(n7163) );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(n7378), .CLK(n7565), .Q(
        g2119), .QN(n7227) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n7378), .CLK(n7565), .Q(
        g2117), .QN(n7230) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n7378), .CLK(n7565), .Q(
        g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n7378), .CLK(n7565), .Q(
        test_so73), .QN(n7266) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n7378), .CLK(
        n7565), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n7378), .CLK(n7565), .Q(
        g2206), .QN(n7180) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n7383), .CLK(n7570), .Q(
        g2207), .QN(n7179) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n7383), .CLK(n7570), .Q(
        g2205), .QN(n6797) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n7378), .CLK(n7565), .Q(
        g2209), .QN(n7178) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n7383), .CLK(n7570), .Q(
        g2210), .QN(n7177) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n7383), .CLK(n7570), .Q(
        g2208), .QN(n6796) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n7383), .CLK(n7570), .Q(
        g2218), .QN(n7176) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n7383), .CLK(n7570), .Q(
        g2219), .QN(n7175) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n7383), .CLK(n7570), .Q(
        g2217), .QN(n6795) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n7383), .CLK(n7570), .Q(
        g2221), .QN(n7174) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n7383), .CLK(n7570), .Q(
        g2222), .QN(n7173) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n7383), .CLK(n7570), .Q(
        g2220), .QN(n6794) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n7383), .CLK(n7570), .Q(
        g2224), .QN(n7172) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n7384), .CLK(n7571), .Q(
        test_so74) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n7380), .CLK(n7567), 
        .Q(g2223), .QN(n6793) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n7380), .CLK(n7567), .Q(
        g2227), .QN(n7171) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n7382), .CLK(n7569), .Q(
        g2228), .QN(n7170) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n7382), .CLK(n7569), .Q(
        g2226), .QN(n6792) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n7382), .CLK(n7569), .Q(
        g2230), .QN(n7169) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n7382), .CLK(n7569), .Q(
        g2231), .QN(n7168) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n7382), .CLK(n7569), .Q(
        g2229), .QN(n6791) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n7382), .CLK(n7569), .Q(
        g2233), .QN(n7167) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n7382), .CLK(n7569), .Q(
        g2234), .QN(n7166) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n7382), .CLK(n7569), .Q(
        g2232), .QN(n6790) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n7382), .CLK(n7569), .Q(
        g2236), .QN(n6781) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n7382), .CLK(n7569), .Q(
        g2237), .QN(n6780) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n7382), .CLK(n7569), .Q(
        g2235), .QN(n6779) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n7383), .CLK(n7570), .Q(
        g2239), .QN(n6789) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n7384), .CLK(n7571), .Q(
        test_so75) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n7381), .CLK(n7568), 
        .Q(g2238), .QN(n6788) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n7381), .CLK(n7568), .Q(
        g2245), .QN(n6859) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n7381), .CLK(n7568), .Q(
        g2246), .QN(n6858) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n7381), .CLK(n7568), .Q(
        g2244), .QN(n6857) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n7381), .CLK(n7568), .Q(
        g2248), .QN(n6856) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n7381), .CLK(n7568), .Q(
        g2249), .QN(n6855) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n7381), .CLK(n7568), .Q(
        g2247), .QN(n6854) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n7381), .CLK(n7568), .Q(
        g2251), .QN(n6853) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n7381), .CLK(n7568), .Q(
        g2252), .QN(n6852) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n7381), .CLK(n7568), .Q(
        g2250), .QN(n6851) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n7381), .CLK(n7568), .Q(
        g2254), .QN(n6850) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n7381), .CLK(n7568), .Q(
        g2255), .QN(n6849) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n7382), .CLK(n7569), .Q(
        g2253), .QN(n6848) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n7394), .CLK(n7581), .Q(
        g2261) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n7394), .CLK(n7581), .Q(
        test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n7394), .CLK(n7581), 
        .Q(g2267) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n7394), .CLK(n7581), .Q(
        g2306) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n7394), .CLK(n7581), .Q(
        g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n7394), .CLK(n7581), .Q(
        g2312) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n7394), .CLK(n7581), .Q(
        g2270) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n7394), .CLK(n7581), .Q(
        g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n7384), .CLK(n7571), .Q(
        g2276) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n7384), .CLK(n7571), .Q(
        g2315) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n7384), .CLK(n7571), .Q(
        g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n7384), .CLK(n7571), .Q(
        g2321) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n7384), .CLK(n7571), .Q(
        g2279) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n7384), .CLK(n7571), .Q(
        g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n7384), .CLK(n7571), .Q(
        g2285) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n7384), .CLK(n7571), .Q(
        g2324) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n7384), .CLK(n7571), .Q(
        test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n7384), .CLK(n7571), 
        .Q(g2330) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n7393), .CLK(n7580), .Q(
        g2288) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n7393), .CLK(n7580), .Q(
        g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n7394), .CLK(n7581), .Q(
        g2294) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n7394), .CLK(n7581), .Q(
        g2333) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n7394), .CLK(n7581), .Q(
        g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n7394), .CLK(n7581), .Q(
        g2339) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n7395), .CLK(n7582), .Q(
        g2297) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n7395), .CLK(n7582), .Q(
        g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n7385), .CLK(n7572), .Q(
        g2303) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n7385), .CLK(n7572), .Q(
        g2342) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n7385), .CLK(n7572), .Q(
        g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n7379), .CLK(n7566), .Q(
        g2348) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n7379), .CLK(n7566), .Q(
        g2160), .QN(n6982) );
  SDFFX1 DFF_1287_Q_reg ( .D(g25940), .SI(g2160), .SE(n7379), .CLK(n7566), .Q(
        test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n7379), .CLK(n7566), 
        .Q(g2151), .QN(n6981) );
  SDFFX1 DFF_1289_Q_reg ( .D(g27131), .SI(g2151), .SE(n7379), .CLK(n7566), .Q(
        g2147), .QN(n6433) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n7379), .CLK(n7566), .Q(
        g2142), .QN(n6980) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n7379), .CLK(n7566), .Q(
        g2138), .QN(n6972) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n7379), .CLK(n7566), .Q(
        g2133), .QN(n6979) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n7379), .CLK(n7566), .Q(
        g2129), .QN(n6969) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n7379), .CLK(n7566), .Q(
        g2124), .QN(n6597) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n7379), .CLK(n7566), .Q(
        g2120), .QN(n6436) );
  SDFFX1 DFF_1296_Q_reg ( .D(g13110), .SI(g2120), .SE(n7380), .CLK(n7567), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n7380), .CLK(n7567), .Q(
        g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n7380), .CLK(n7567), .Q(
        g2257), .QN(n6998) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n7380), .CLK(n7567), .Q(
        g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n7380), .CLK(n7567), .Q(
        test_so79) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n7392), .CLK(n7579), 
        .Q(g2429), .QN(n6927) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n7393), .CLK(n7580), .Q(
        g2418), .QN(n6926) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n7393), .CLK(n7580), .Q(
        g2421), .QN(n6925) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n7393), .CLK(n7580), .Q(
        g2444), .QN(n6904) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n7393), .CLK(n7580), .Q(
        g2433), .QN(n6903) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n7392), .CLK(n7579), .Q(
        g2436), .QN(n6902) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n7392), .CLK(n7579), .Q(
        g2459), .QN(n6646) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n7392), .CLK(n7579), .Q(
        g2448), .QN(n6648) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n7392), .CLK(n7579), .Q(
        g2451), .QN(n6647) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n7393), .CLK(n7580), .Q(
        g2473), .QN(n6916) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n7393), .CLK(n7580), .Q(
        g2463), .QN(n6915) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n7385), .CLK(n7572), .Q(
        g2466), .QN(n6914) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n7385), .CLK(n7572), .Q(
        g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n7392), .CLK(n7579), .Q(
        g2486) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n7392), .CLK(n7579), .Q(
        test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n7385), .CLK(n7572), 
        .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n7385), .CLK(n7572), .Q(
        g2495) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n7385), .CLK(n7572), .Q(
        g2498) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n7389), .CLK(n7576), .Q(
        g2502), .QN(n6948) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n7389), .CLK(n7576), .Q(
        g2503), .QN(n6938) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n7389), .CLK(n7576), .Q(
        g2501), .QN(n6947) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n7389), .CLK(n7576), .Q(
        g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n7389), .CLK(n7576), .Q(
        g2507) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n7389), .CLK(n7576), .Q(
        g2510) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n7389), .CLK(n7576), .Q(
        g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n7390), .CLK(n7577), .Q(
        g2516) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n7390), .CLK(n7577), .Q(
        g2519) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n7390), .CLK(n7577), .Q(
        g2523), .QN(n6946) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n7389), .CLK(n7576), .Q(
        g2524), .QN(n6937) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n7389), .CLK(n7576), .Q(
        test_so81) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n7385), .CLK(n7572), 
        .Q(g2387), .QN(n6545) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n7385), .CLK(n7572), .Q(
        g2388), .QN(n6533) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n7385), .CLK(n7572), .Q(
        g2389), .QN(n6544) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n7385), .CLK(n7572), .Q(
        g2390), .QN(n6543) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n7378), .CLK(n7565), .Q(
        g2391), .QN(n6532) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n7380), .CLK(n7567), .Q(
        g2392), .QN(n6542) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n7379), .CLK(n7566), .Q(
        g2393), .QN(n6541) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n7380), .CLK(n7567), .Q(
        g2394), .QN(n6531) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n7380), .CLK(n7567), .Q(
        g2395), .QN(n6540) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n7395), .CLK(n7582), .Q(
        g2397), .QN(n6589) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n7395), .CLK(n7582), .Q(
        g2398), .QN(n6585) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n7393), .CLK(n7580), .Q(
        g2396), .QN(n6588) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n7393), .CLK(n7580), .Q(
        g2478), .QN(n6945) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n7393), .CLK(n7580), .Q(
        g2479), .QN(n6936) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n7393), .CLK(n7580), .Q(
        test_so82) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n7304), .CLK(n7491), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n7304), .CLK(n7491), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n7304), .CLK(n7491), .Q(
        g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n7304), .CLK(n7491), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n7304), .CLK(n7491), .Q(
        g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n7304), .CLK(n7491), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n7304), .CLK(n7491), .Q(
        g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n7304), .CLK(n7491), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n7304), .CLK(n7491), .Q(
        g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n7304), .CLK(n7491), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n7304), .CLK(n7491), .Q(
        g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n7304), .CLK(n7491), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n7305), .CLK(n7492), .Q(
        g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n7305), .CLK(n7492), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n7305), .CLK(n7492), .Q(
        test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n7305), .CLK(
        n7492), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n7318), .CLK(n7505), .Q(
        g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n7318), .CLK(n7505), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n7392), .CLK(n7579), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n7398), .CLK(n7585), .Q(
        g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n7395), .CLK(n7582), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n7395), .CLK(n7582), .Q(
        g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n7395), .CLK(n7582), .Q(
        g2424) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n7395), .CLK(n7582), .Q(
        g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n7395), .CLK(n7582), .Q(
        g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n7395), .CLK(n7582), .Q(
        g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n7395), .CLK(n7582), .Q(
        g2428) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n7395), .CLK(n7582), .Q(
        g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n7396), .CLK(n7583), .Q(
        g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n7396), .CLK(n7583), .Q(
        test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n7396), .CLK(
        n7583), .Q(g2441) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n7396), .CLK(n7583), .Q(
        g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n7396), .CLK(n7583), .Q(
        g2443) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n7396), .CLK(n7583), .Q(
        g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n7396), .CLK(n7583), .Q(
        g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n7396), .CLK(n7583), .Q(
        g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n7396), .CLK(n7583), .Q(
        g2456) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n7396), .CLK(n7583), .Q(
        g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n7396), .CLK(n7583), .Q(
        g2458) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n7396), .CLK(n7583), .Q(
        g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n7397), .CLK(n7584), .Q(
        g2469) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n7397), .CLK(n7584), .Q(
        g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n7397), .CLK(n7584), .Q(
        g2471) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n7397), .CLK(n7584), .Q(
        g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n7397), .CLK(n7584), .Q(
        test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n7330), .CLK(n7517), 
        .Q(g5747) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n7330), .CLK(n7517), .Q(
        g5796) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n7330), .CLK(n7517), .Q(
        g2412) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n7330), .CLK(n7517), .Q(
        g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n7330), .CLK(n7517), .Q(
        g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n7331), .CLK(n7518), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(g21847), .SI(g2624), .SE(n7331), .CLK(n7518), .Q(
        g2628), .QN(n7233) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n7331), .CLK(n7518), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n7331), .CLK(n7518), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n765), .SI(g2584), .SE(n7388), .CLK(n7575), .Q(
        g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n7388), .CLK(n7575), .Q(
        g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n7388), .CLK(n7575), .Q(
        g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n7387), .CLK(n7574), .Q(
        g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n7387), .CLK(n7574), .Q(
        g2643) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n7387), .CLK(n7574), .Q(
        test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n7388), .CLK(
        n7575), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n7388), .CLK(n7575), .Q(
        g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n7388), .CLK(n7575), .Q(
        g2647) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n7386), .CLK(n7573), .Q(
        g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n7386), .CLK(n7573), .Q(
        g2639) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n7386), .CLK(n7573), .Q(
        g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n7386), .CLK(n7573), .Q(
        g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n7386), .CLK(n7573), .Q(
        g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n7386), .CLK(n7573), .Q(
        g2564) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n7386), .CLK(n7573), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n7386), .CLK(n7573), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n7387), .CLK(n7574), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n7390), .CLK(n7577), .Q(
        g2561) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n7390), .CLK(n7577), .Q(
        g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n7390), .CLK(n7577), .Q(
        test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n7387), .CLK(n7574), 
        .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n7387), .CLK(n7574), .Q(
        g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n7387), .CLK(n7574), .Q(
        g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n7388), .CLK(n7575), .Q(
        g2552) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n7388), .CLK(n7575), .Q(
        g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n7388), .CLK(n7575), .Q(
        g2554) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n7386), .CLK(n7573), .Q(
        g2555) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n7386), .CLK(n7573), .Q(
        g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n7386), .CLK(n7573), .Q(
        g2539) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n7386), .CLK(n7573), .Q(
        g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n7387), .CLK(n7574), .Q(
        g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n7387), .CLK(n7574), .Q(
        g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n758), .SI(g2546), .SE(n7387), .CLK(n7574), .Q(
        g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n7387), .CLK(n7574), .Q(
        g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n7387), .CLK(n7574), .Q(
        test_so88) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n7388), .CLK(n7575), 
        .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n7388), .CLK(n7575), .Q(
        n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n7389), .CLK(n7576), .Q(
        n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n7388), .CLK(n7575), .Q(
        g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n7389), .CLK(n7576), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n7390), .CLK(n7577), .Q(
        g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n7390), .CLK(n7577), .Q(
        g2633) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n7390), .CLK(n7577), .Q(
        g2650), .QN(n6601) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n7391), .CLK(n7578), .Q(
        g2651), .QN(n6603) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n7391), .CLK(n7578), .Q(
        g2649), .QN(n6602) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n7391), .CLK(n7578), .Q(
        g2653), .QN(n6613) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n7392), .CLK(n7579), .Q(
        g2654), .QN(n6615) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n7392), .CLK(n7579), .Q(
        g2652), .QN(n6614) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n7392), .CLK(n7579), .Q(
        g2656), .QN(n6440) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n7392), .CLK(n7579), .Q(
        test_so89) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n7391), .CLK(n7578), 
        .Q(g2655), .QN(n6441) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n7391), .CLK(n7578), .Q(
        g2659), .QN(n6624) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n7391), .CLK(n7578), .Q(
        g2660), .QN(n6626) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n7390), .CLK(n7577), .Q(
        g2658), .QN(n6625) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n7390), .CLK(n7577), .Q(
        g2661) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n7390), .CLK(n7577), .Q(
        g2664) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n7391), .CLK(n7578), .Q(
        g2667) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n7391), .CLK(n7578), .Q(
        g2670) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n7391), .CLK(n7578), .Q(
        g2673) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n7391), .CLK(n7578), .Q(
        g2676) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n7391), .CLK(n7578), .Q(
        g2688) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n7391), .CLK(n7578), .Q(
        g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n7319), .CLK(n7506), .Q(
        g2694) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n7397), .CLK(n7584), .Q(
        g2679) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n7397), .CLK(n7584), .Q(
        test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n7397), .CLK(n7584), 
        .Q(g2685) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n7397), .CLK(n7584), .Q(
        g2565) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n7397), .CLK(n7584), .Q(
        g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n7319), .CLK(n7506), .Q(
        g2571) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n7389), .CLK(n7576), .Q(
        g2580), .QN(n6766) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n7319), .CLK(n7506), .Q(
        n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n7319), .CLK(n7506), .Q(
        g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n7320), .CLK(n7507), 
        .Q(g2599), .QN(n7002) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n7320), .CLK(n7507), 
        .Q(n7925), .QN(DFF_1494_n1) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n7320), .CLK(n7507), 
        .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n7320), .CLK(n7507), 
        .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n7320), .CLK(n7507), 
        .Q(n7922), .QN(DFF_1497_n1) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n7320), .CLK(n7507), 
        .Q(n7921), .QN(DFF_1498_n1) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n7320), .CLK(n7507), 
        .Q(n7920), .QN(DFF_1499_n1) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n7320), .CLK(n7507), 
        .Q(test_so91), .QN(n6411) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n7305), .CLK(
        n7492), .Q(g2611), .QN(n6410) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n7398), .CLK(n7585), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n7318), .CLK(n7505), .Q(
        n7918), .QN(n13228) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n7331), .CLK(n7518), .Q(
        g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n7331), .CLK(n7518), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n7331), .CLK(n7518), .Q(
        g2704), .QN(n7041) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n7336), .CLK(n7523), .Q(
        g2733) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n7336), .CLK(n7523), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(n7336), .CLK(n7523), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n7336), .CLK(n7523), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n7336), .CLK(n7523), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n7336), .CLK(n7523), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(n7337), .CLK(n7524), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n7337), .CLK(n7524), .Q(
        test_so92), .QN(n7269) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n7337), .CLK(n7524), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(g27724), .SI(g2753), .SE(n7337), .CLK(n7524), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n7337), .CLK(n7524), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n7337), .CLK(n7524), .Q(
        g2773), .QN(n7069) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n7337), .CLK(n7524), .Q(
        g2774), .QN(n7068) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n7337), .CLK(n7524), .Q(
        g2772), .QN(n7131) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n7337), .CLK(n7524), .Q(
        g2776), .QN(n7067) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n7338), .CLK(n7525), .Q(
        g2777), .QN(n7066) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n7338), .CLK(n7525), .Q(
        g2775), .QN(n7130) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n7338), .CLK(n7525), .Q(
        g2779), .QN(n7065) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n7338), .CLK(n7525), .Q(
        g2780), .QN(n7064) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n7338), .CLK(n7525), .Q(
        g2778), .QN(n7129) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n7339), .CLK(n7526), .Q(
        g2782), .QN(n7063) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n7339), .CLK(n7526), .Q(
        g2783), .QN(n7062) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n7340), .CLK(n7527), .Q(
        test_so93) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n7337), .CLK(n7524), 
        .Q(g2785), .QN(n7061) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n7337), .CLK(n7524), .Q(
        g2786), .QN(n7060) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n7337), .CLK(n7524), .Q(
        g2784), .QN(n7128) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n7338), .CLK(n7525), .Q(
        g2788), .QN(n7059) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n7339), .CLK(n7526), .Q(
        g2789), .QN(n7058) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n7339), .CLK(n7526), .Q(
        g2787), .QN(n7127) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n7339), .CLK(n7526), .Q(
        g2791), .QN(n7057) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n7339), .CLK(n7526), .Q(
        g2792), .QN(n7056) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n7339), .CLK(n7526), .Q(
        g2790), .QN(n7126) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n7339), .CLK(n7526), .Q(
        g2794), .QN(n7055) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n7339), .CLK(n7526), .Q(
        g2795), .QN(n7054) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n7339), .CLK(n7526), .Q(
        g2793), .QN(n7125) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n7339), .CLK(n7526), .Q(
        g2797), .QN(n7053) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n7339), .CLK(n7526), .Q(
        g2798), .QN(n7052) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n7320), .CLK(n7507), .Q(
        test_so94) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n7338), .CLK(n7525), 
        .Q(g2800), .QN(n7051) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n7338), .CLK(n7525), .Q(
        g2801), .QN(n7050) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n7338), .CLK(n7525), .Q(
        g2799), .QN(n7124) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n7338), .CLK(n7525), .Q(
        g2803), .QN(n6841) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n7338), .CLK(n7525), .Q(
        g2804) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n7338), .CLK(n7525), .Q(
        g2802), .QN(n6896) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n7397), .CLK(n7584), .Q(
        g2806), .QN(n6840) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n7397), .CLK(n7584), .Q(
        g2807), .QN(n6832) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n7398), .CLK(n7585), .Q(
        g2805), .QN(n6895) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n7398), .CLK(n7585), .Q(
        g2809), .QN(n6768) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n7398), .CLK(n7585), .Q(
        g2810), .QN(n6767) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n7398), .CLK(n7585), .Q(
        g2808), .QN(n6775) );
  SDFFX1 DFF_1558_Q_reg ( .D(g22269), .SI(g2808), .SE(n7398), .CLK(n7585), .Q(
        g2812), .QN(n7162) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n7398), .CLK(n7585), .Q(
        g2813), .QN(n7226) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n7398), .CLK(n7585), .Q(
        test_so95) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n7320), .CLK(n7507), 
        .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n7320), .CLK(n7507), .Q(
        n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263_Tj_Payload), .SI(n7912), .SE(n7320), .CLK(
        n7507), .Q(n4598), .QN(n6431) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n7280), .CLK(n7467), .Q(
        g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n7280), .CLK(n7467), .Q(
        g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n7280), .CLK(n7467), .Q(
        g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n7280), .CLK(n7467), .Q(
        g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n7280), .CLK(n7467), .Q(
        g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n7281), .CLK(n7468), .Q(
        g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n7281), .CLK(n7468), .Q(
        g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n7281), .CLK(n7468), .Q(
        g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n7281), .CLK(n7468), .Q(
        g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n7281), .CLK(n7468), .Q(
        g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n7281), .CLK(n7468), .Q(
        g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n7281), .CLK(n7468), .Q(
        test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n7371), .CLK(n7558), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n7371), .CLK(n7558), .Q(
        g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n7371), .CLK(n7558), .Q(
        g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n7371), .CLK(n7558), .Q(
        g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n7371), .CLK(n7558), .Q(
        g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n7371), .CLK(n7558), .Q(
        g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n7398), .CLK(n7585), .Q(
        g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n7398), .CLK(n7585), .Q(
        g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n7399), .CLK(n7586), .Q(
        g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n7399), .CLK(n7586), .Q(
        g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n7399), .CLK(n7586), .Q(
        g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n7399), .CLK(n7586), .Q(
        g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n7399), .CLK(n7586), .Q(
        g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n7399), .CLK(n7586), .Q(
        g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n7400), .CLK(n7587), .Q(
        test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n7400), .CLK(n7587), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n7400), .CLK(n7587), .Q(
        g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n7400), .CLK(n7587), .Q(
        g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n7400), .CLK(n7587), .Q(
        g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n7401), .CLK(n7588), .Q(
        g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n7401), .CLK(n7588), .Q(
        g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n7401), .CLK(n7588), .Q(
        g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n7401), .CLK(n7588), .Q(
        g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n7318), .CLK(n7505), .Q(
        g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n7319), .CLK(n7506), .Q(
        g2993), .QN(n6432) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n7331), .CLK(n7518), .Q(
        n7909), .QN(n13235) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(n7331), .CLK(n7518), .Q(
        g3006), .QN(n6428) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n7331), .CLK(n7518), .Q(
        g3002), .QN(n6430) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n7331), .CLK(n7518), .Q(
        g3013), .QN(n6427) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n7332), .CLK(n7519), .Q(
        test_so98), .QN(n7273) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n7332), .CLK(n7519), 
        .Q(g3024), .QN(n6429) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n7319), .CLK(n7506), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(n7319), .CLK(n7506), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n7319), .CLK(n7506), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n7319), .CLK(n7506), .Q(
        g3032), .QN(n6706) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n7319), .CLK(n7506), .Q(
        g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n7319), .CLK(n7506), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n7319), .CLK(n7506), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n7398), .CLK(n7585), .Q(
        g8275) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n7399), .CLK(n7586), .Q(
        g8274), .QN(n7257) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n7399), .CLK(n7586), .Q(
        g8273), .QN(n13238) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n7399), .CLK(n7586), .Q(
        g8272), .QN(n13237) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n7399), .CLK(n7586), .Q(
        g8268), .QN(n13236) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n7399), .CLK(n7586), .Q(
        g8269), .QN(n7258) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n7399), .CLK(n7586), .Q(
        test_so99) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n7400), .CLK(n7587), 
        .Q(g8271), .QN(n7256) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n7400), .CLK(n7587), .Q(
        g3083), .QN(n7261) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n7400), .CLK(n7587), .Q(
        g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n7400), .CLK(n7587), .Q(
        n4577), .QN(n6709) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n7400), .CLK(n7587), .Q(
        g8266), .QN(n13241) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n7400), .CLK(n7587), .Q(
        g8265), .QN(n13240) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n7281), .CLK(n7468), .Q(
        g8264), .QN(n7239) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n7400), .CLK(n7587), .Q(
        g8262) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n7401), .CLK(n7588), .Q(
        g8263), .QN(n7240) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n7401), .CLK(n7588), .Q(
        g8260), .QN(n7237) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n7401), .CLK(n7588), .Q(
        g8261), .QN(n13239) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n7401), .CLK(n7588), .Q(
        g8259), .QN(n7238) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n7401), .CLK(n7588), .Q(
        g2990), .QN(n7259) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n7281), .CLK(n7468), .Q(
        n4578), .QN(n6708) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n7405), .CLK(n7592), .Q(
        test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n7321), .CLK(n7508), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n7321), .CLK(n7508), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n7321), .CLK(n7508), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n7331), .CLK(n7518), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n7380), .CLK(n7567), .Q(
        g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n7352), .CLK(n7539), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n7352), .CLK(n7539), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n7380), .CLK(n7567), .Q(
        n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n7279), .CLK(n7466), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n7279), .CLK(n7466), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n3065), .IN2(n3016), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n3023), .IN2(n3000), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n3008), .IN2(n3068), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n3128), .IN2(n3036), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(n3758), .IN2(n3788), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n3751), .IN2(n3749), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n2792), .IN2(n2632), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n2351), .IN2(n2430), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(n4263), .Q(n4263_Tj_Payload)
         );
  NBUFFX2 U7253 ( .INP(n7449), .Z(n7276) );
  NBUFFX2 U7254 ( .INP(n7449), .Z(n7275) );
  NBUFFX2 U7255 ( .INP(n7407), .Z(n7400) );
  NBUFFX2 U7256 ( .INP(n7408), .Z(n7399) );
  NBUFFX2 U7257 ( .INP(n7428), .Z(n7339) );
  NBUFFX2 U7258 ( .INP(n7428), .Z(n7338) );
  NBUFFX2 U7259 ( .INP(n7428), .Z(n7337) );
  NBUFFX2 U7260 ( .INP(n7434), .Z(n7320) );
  NBUFFX2 U7261 ( .INP(n7434), .Z(n7319) );
  NBUFFX2 U7262 ( .INP(n7410), .Z(n7391) );
  NBUFFX2 U7263 ( .INP(n7412), .Z(n7386) );
  NBUFFX2 U7264 ( .INP(n7412), .Z(n7387) );
  NBUFFX2 U7265 ( .INP(n7411), .Z(n7388) );
  NBUFFX2 U7266 ( .INP(n7430), .Z(n7331) );
  NBUFFX2 U7267 ( .INP(n7408), .Z(n7397) );
  NBUFFX2 U7268 ( .INP(n7409), .Z(n7396) );
  NBUFFX2 U7269 ( .INP(n7408), .Z(n7398) );
  NBUFFX2 U7270 ( .INP(n7439), .Z(n7304) );
  NBUFFX2 U7271 ( .INP(n7411), .Z(n7390) );
  NBUFFX2 U7272 ( .INP(n7411), .Z(n7389) );
  NBUFFX2 U7273 ( .INP(n7410), .Z(n7392) );
  NBUFFX2 U7274 ( .INP(n7414), .Z(n7379) );
  NBUFFX2 U7275 ( .INP(n7412), .Z(n7385) );
  NBUFFX2 U7276 ( .INP(n7409), .Z(n7395) );
  NBUFFX2 U7277 ( .INP(n7410), .Z(n7393) );
  NBUFFX2 U7278 ( .INP(n7409), .Z(n7394) );
  NBUFFX2 U7279 ( .INP(n7414), .Z(n7381) );
  NBUFFX2 U7280 ( .INP(n7413), .Z(n7382) );
  NBUFFX2 U7281 ( .INP(n7414), .Z(n7380) );
  NBUFFX2 U7282 ( .INP(n7413), .Z(n7384) );
  NBUFFX2 U7283 ( .INP(n7413), .Z(n7383) );
  NBUFFX2 U7284 ( .INP(n7415), .Z(n7378) );
  NBUFFX2 U7285 ( .INP(n7415), .Z(n7377) );
  NBUFFX2 U7286 ( .INP(n7415), .Z(n7376) );
  NBUFFX2 U7287 ( .INP(n7416), .Z(n7375) );
  NBUFFX2 U7288 ( .INP(n7416), .Z(n7374) );
  NBUFFX2 U7289 ( .INP(n7416), .Z(n7373) );
  NBUFFX2 U7290 ( .INP(n7417), .Z(n7372) );
  NBUFFX2 U7291 ( .INP(n7417), .Z(n7371) );
  NBUFFX2 U7292 ( .INP(n7417), .Z(n7370) );
  NBUFFX2 U7294 ( .INP(n7418), .Z(n7369) );
  NBUFFX2 U7295 ( .INP(n7418), .Z(n7368) );
  NBUFFX2 U7296 ( .INP(n7418), .Z(n7367) );
  NBUFFX2 U7297 ( .INP(n7419), .Z(n7366) );
  NBUFFX2 U7298 ( .INP(n7419), .Z(n7365) );
  NBUFFX2 U7299 ( .INP(n7419), .Z(n7364) );
  NBUFFX2 U7300 ( .INP(n7420), .Z(n7361) );
  NBUFFX2 U7301 ( .INP(n7421), .Z(n7358) );
  NBUFFX2 U7302 ( .INP(n7421), .Z(n7359) );
  NBUFFX2 U7303 ( .INP(n7421), .Z(n7360) );
  NBUFFX2 U7304 ( .INP(n7422), .Z(n7357) );
  NBUFFX2 U7305 ( .INP(n7422), .Z(n7356) );
  NBUFFX2 U7306 ( .INP(n7420), .Z(n7363) );
  NBUFFX2 U7307 ( .INP(n7420), .Z(n7362) );
  NBUFFX2 U7308 ( .INP(n7422), .Z(n7355) );
  NBUFFX2 U7309 ( .INP(n7423), .Z(n7354) );
  NBUFFX2 U7310 ( .INP(n7423), .Z(n7353) );
  NBUFFX2 U7311 ( .INP(n7423), .Z(n7352) );
  NBUFFX2 U7312 ( .INP(n7424), .Z(n7351) );
  NBUFFX2 U7313 ( .INP(n7424), .Z(n7350) );
  NBUFFX2 U7314 ( .INP(n7424), .Z(n7349) );
  NBUFFX2 U7315 ( .INP(n7425), .Z(n7348) );
  NBUFFX2 U7316 ( .INP(n7429), .Z(n7336) );
  NBUFFX2 U7317 ( .INP(n7425), .Z(n7347) );
  NBUFFX2 U7318 ( .INP(n7425), .Z(n7346) );
  NBUFFX2 U7319 ( .INP(n7426), .Z(n7345) );
  NBUFFX2 U7320 ( .INP(n7433), .Z(n7324) );
  NBUFFX2 U7321 ( .INP(n7433), .Z(n7323) );
  NBUFFX2 U7322 ( .INP(n7433), .Z(n7322) );
  NBUFFX2 U7323 ( .INP(n7441), .Z(n7300) );
  NBUFFX2 U7324 ( .INP(n7441), .Z(n7298) );
  NBUFFX2 U7325 ( .INP(n7443), .Z(n7294) );
  NBUFFX2 U7326 ( .INP(n7442), .Z(n7295) );
  NBUFFX2 U7327 ( .INP(n7444), .Z(n7289) );
  NBUFFX2 U7328 ( .INP(n7442), .Z(n7296) );
  NBUFFX2 U7329 ( .INP(n7443), .Z(n7293) );
  NBUFFX2 U7330 ( .INP(n7442), .Z(n7297) );
  NBUFFX2 U7331 ( .INP(n7445), .Z(n7287) );
  NBUFFX2 U7332 ( .INP(n7445), .Z(n7288) );
  NBUFFX2 U7333 ( .INP(n7444), .Z(n7290) );
  NBUFFX2 U7334 ( .INP(n7443), .Z(n7292) );
  NBUFFX2 U7335 ( .INP(n7444), .Z(n7291) );
  NBUFFX2 U7336 ( .INP(n7429), .Z(n7334) );
  NBUFFX2 U7337 ( .INP(n7429), .Z(n7335) );
  NBUFFX2 U7338 ( .INP(n7430), .Z(n7333) );
  NBUFFX2 U7339 ( .INP(n7430), .Z(n7332) );
  NBUFFX2 U7340 ( .INP(n7434), .Z(n7321) );
  NBUFFX2 U7341 ( .INP(n7426), .Z(n7344) );
  NBUFFX2 U7342 ( .INP(n7426), .Z(n7343) );
  NBUFFX2 U7343 ( .INP(n7427), .Z(n7342) );
  NBUFFX2 U7344 ( .INP(n7427), .Z(n7341) );
  NBUFFX2 U7345 ( .INP(n7427), .Z(n7340) );
  NBUFFX2 U7346 ( .INP(n7431), .Z(n7330) );
  NBUFFX2 U7347 ( .INP(n7431), .Z(n7329) );
  NBUFFX2 U7348 ( .INP(n7431), .Z(n7328) );
  NBUFFX2 U7349 ( .INP(n7432), .Z(n7327) );
  NBUFFX2 U7350 ( .INP(n7432), .Z(n7326) );
  NBUFFX2 U7351 ( .INP(n7432), .Z(n7325) );
  NBUFFX2 U7352 ( .INP(n7447), .Z(n7280) );
  NBUFFX2 U7353 ( .INP(n7436), .Z(n7313) );
  NBUFFX2 U7354 ( .INP(n7437), .Z(n7312) );
  NBUFFX2 U7355 ( .INP(n7436), .Z(n7315) );
  NBUFFX2 U7356 ( .INP(n7436), .Z(n7314) );
  NBUFFX2 U7357 ( .INP(n7448), .Z(n7279) );
  NBUFFX2 U7358 ( .INP(n7437), .Z(n7311) );
  NBUFFX2 U7359 ( .INP(n7435), .Z(n7317) );
  NBUFFX2 U7360 ( .INP(n7435), .Z(n7316) );
  NBUFFX2 U7361 ( .INP(n7437), .Z(n7310) );
  NBUFFX2 U7362 ( .INP(n7438), .Z(n7309) );
  NBUFFX2 U7363 ( .INP(n7438), .Z(n7308) );
  NBUFFX2 U7364 ( .INP(n7438), .Z(n7307) );
  NBUFFX2 U7365 ( .INP(n7439), .Z(n7306) );
  NBUFFX2 U7366 ( .INP(n7439), .Z(n7305) );
  NBUFFX2 U7367 ( .INP(n7447), .Z(n7281) );
  NBUFFX2 U7368 ( .INP(n7446), .Z(n7284) );
  NBUFFX2 U7369 ( .INP(n7447), .Z(n7282) );
  NBUFFX2 U7370 ( .INP(n7446), .Z(n7283) );
  NBUFFX2 U7371 ( .INP(n7406), .Z(n7404) );
  NBUFFX2 U7372 ( .INP(n7406), .Z(n7403) );
  NBUFFX2 U7373 ( .INP(n7407), .Z(n7402) );
  NBUFFX2 U7374 ( .INP(n7407), .Z(n7401) );
  NBUFFX2 U7375 ( .INP(n7435), .Z(n7318) );
  NBUFFX2 U7376 ( .INP(n7440), .Z(n7303) );
  NBUFFX2 U7377 ( .INP(n7440), .Z(n7302) );
  NBUFFX2 U7378 ( .INP(n7440), .Z(n7301) );
  NBUFFX2 U7379 ( .INP(n7441), .Z(n7299) );
  NBUFFX2 U7380 ( .INP(n7445), .Z(n7286) );
  NBUFFX2 U7381 ( .INP(n7446), .Z(n7285) );
  NBUFFX2 U7382 ( .INP(n7448), .Z(n7278) );
  NBUFFX2 U7383 ( .INP(n7448), .Z(n7277) );
  NBUFFX2 U7384 ( .INP(n7636), .Z(n7463) );
  NBUFFX2 U7385 ( .INP(n7636), .Z(n7462) );
  NBUFFX2 U7386 ( .INP(n7594), .Z(n7587) );
  NBUFFX2 U7387 ( .INP(n7595), .Z(n7586) );
  NBUFFX2 U7388 ( .INP(n7615), .Z(n7526) );
  NBUFFX2 U7389 ( .INP(n7615), .Z(n7525) );
  NBUFFX2 U7390 ( .INP(n7615), .Z(n7524) );
  NBUFFX2 U7391 ( .INP(n7621), .Z(n7507) );
  NBUFFX2 U7392 ( .INP(n7621), .Z(n7506) );
  NBUFFX2 U7393 ( .INP(n7597), .Z(n7578) );
  NBUFFX2 U7394 ( .INP(n7599), .Z(n7573) );
  NBUFFX2 U7395 ( .INP(n7599), .Z(n7574) );
  NBUFFX2 U7396 ( .INP(n7598), .Z(n7575) );
  NBUFFX2 U7397 ( .INP(n7617), .Z(n7518) );
  NBUFFX2 U7398 ( .INP(n7595), .Z(n7584) );
  NBUFFX2 U7399 ( .INP(n7596), .Z(n7583) );
  NBUFFX2 U7400 ( .INP(n7595), .Z(n7585) );
  NBUFFX2 U7401 ( .INP(n7626), .Z(n7491) );
  NBUFFX2 U7402 ( .INP(n7598), .Z(n7577) );
  NBUFFX2 U7403 ( .INP(n7598), .Z(n7576) );
  NBUFFX2 U7404 ( .INP(n7597), .Z(n7579) );
  NBUFFX2 U7405 ( .INP(n7601), .Z(n7566) );
  NBUFFX2 U7406 ( .INP(n7599), .Z(n7572) );
  NBUFFX2 U7407 ( .INP(n7596), .Z(n7582) );
  NBUFFX2 U7408 ( .INP(n7597), .Z(n7580) );
  NBUFFX2 U7409 ( .INP(n7596), .Z(n7581) );
  NBUFFX2 U7410 ( .INP(n7601), .Z(n7568) );
  NBUFFX2 U7411 ( .INP(n7600), .Z(n7569) );
  NBUFFX2 U7412 ( .INP(n7601), .Z(n7567) );
  NBUFFX2 U7413 ( .INP(n7600), .Z(n7571) );
  NBUFFX2 U7414 ( .INP(n7600), .Z(n7570) );
  NBUFFX2 U7415 ( .INP(n7602), .Z(n7565) );
  NBUFFX2 U7416 ( .INP(n7602), .Z(n7564) );
  NBUFFX2 U7417 ( .INP(n7602), .Z(n7563) );
  NBUFFX2 U7418 ( .INP(n7603), .Z(n7562) );
  NBUFFX2 U7419 ( .INP(n7603), .Z(n7561) );
  NBUFFX2 U7420 ( .INP(n7603), .Z(n7560) );
  NBUFFX2 U7421 ( .INP(n7604), .Z(n7559) );
  NBUFFX2 U7422 ( .INP(n7604), .Z(n7558) );
  NBUFFX2 U7423 ( .INP(n7604), .Z(n7557) );
  NBUFFX2 U7424 ( .INP(n7605), .Z(n7556) );
  NBUFFX2 U7425 ( .INP(n7605), .Z(n7555) );
  NBUFFX2 U7426 ( .INP(n7605), .Z(n7554) );
  NBUFFX2 U7427 ( .INP(n7606), .Z(n7553) );
  NBUFFX2 U7428 ( .INP(n7606), .Z(n7552) );
  NBUFFX2 U7429 ( .INP(n7606), .Z(n7551) );
  NBUFFX2 U7430 ( .INP(n7607), .Z(n7548) );
  NBUFFX2 U7431 ( .INP(n7608), .Z(n7545) );
  NBUFFX2 U7432 ( .INP(n7608), .Z(n7546) );
  NBUFFX2 U7433 ( .INP(n7608), .Z(n7547) );
  NBUFFX2 U7434 ( .INP(n7609), .Z(n7544) );
  NBUFFX2 U7435 ( .INP(n7609), .Z(n7543) );
  NBUFFX2 U7436 ( .INP(n7607), .Z(n7550) );
  NBUFFX2 U7437 ( .INP(n7607), .Z(n7549) );
  NBUFFX2 U7438 ( .INP(n7609), .Z(n7542) );
  NBUFFX2 U7439 ( .INP(n7610), .Z(n7541) );
  NBUFFX2 U7440 ( .INP(n7610), .Z(n7540) );
  NBUFFX2 U7441 ( .INP(n7610), .Z(n7539) );
  NBUFFX2 U7442 ( .INP(n7611), .Z(n7538) );
  NBUFFX2 U7443 ( .INP(n7611), .Z(n7537) );
  NBUFFX2 U7444 ( .INP(n7611), .Z(n7536) );
  NBUFFX2 U7445 ( .INP(n7612), .Z(n7535) );
  NBUFFX2 U7446 ( .INP(n7616), .Z(n7523) );
  NBUFFX2 U7447 ( .INP(n7612), .Z(n7534) );
  NBUFFX2 U7448 ( .INP(n7612), .Z(n7533) );
  NBUFFX2 U7449 ( .INP(n7613), .Z(n7532) );
  NBUFFX2 U7450 ( .INP(n7620), .Z(n7511) );
  NBUFFX2 U7451 ( .INP(n7620), .Z(n7510) );
  NBUFFX2 U7452 ( .INP(n7620), .Z(n7509) );
  NBUFFX2 U7453 ( .INP(n7628), .Z(n7487) );
  NBUFFX2 U7454 ( .INP(n7628), .Z(n7485) );
  NBUFFX2 U7455 ( .INP(n7630), .Z(n7481) );
  NBUFFX2 U7456 ( .INP(n7629), .Z(n7482) );
  NBUFFX2 U7457 ( .INP(n7631), .Z(n7476) );
  NBUFFX2 U7458 ( .INP(n7629), .Z(n7483) );
  NBUFFX2 U7459 ( .INP(n7630), .Z(n7480) );
  NBUFFX2 U7460 ( .INP(n7629), .Z(n7484) );
  NBUFFX2 U7461 ( .INP(n7632), .Z(n7474) );
  NBUFFX2 U7462 ( .INP(n7632), .Z(n7475) );
  NBUFFX2 U7463 ( .INP(n7631), .Z(n7477) );
  NBUFFX2 U7464 ( .INP(n7630), .Z(n7479) );
  NBUFFX2 U7465 ( .INP(n7631), .Z(n7478) );
  NBUFFX2 U7466 ( .INP(n7616), .Z(n7521) );
  NBUFFX2 U7467 ( .INP(n7616), .Z(n7522) );
  NBUFFX2 U7468 ( .INP(n7617), .Z(n7520) );
  NBUFFX2 U7469 ( .INP(n7617), .Z(n7519) );
  NBUFFX2 U7470 ( .INP(n7621), .Z(n7508) );
  NBUFFX2 U7471 ( .INP(n7613), .Z(n7531) );
  NBUFFX2 U7472 ( .INP(n7613), .Z(n7530) );
  NBUFFX2 U7473 ( .INP(n7614), .Z(n7529) );
  NBUFFX2 U7474 ( .INP(n7614), .Z(n7528) );
  NBUFFX2 U7475 ( .INP(n7614), .Z(n7527) );
  NBUFFX2 U7476 ( .INP(n7618), .Z(n7517) );
  NBUFFX2 U7477 ( .INP(n7618), .Z(n7516) );
  NBUFFX2 U7478 ( .INP(n7618), .Z(n7515) );
  NBUFFX2 U7479 ( .INP(n7619), .Z(n7514) );
  NBUFFX2 U7480 ( .INP(n7619), .Z(n7513) );
  NBUFFX2 U7481 ( .INP(n7619), .Z(n7512) );
  NBUFFX2 U7482 ( .INP(n7634), .Z(n7467) );
  NBUFFX2 U7483 ( .INP(n7623), .Z(n7500) );
  NBUFFX2 U7484 ( .INP(n7624), .Z(n7499) );
  NBUFFX2 U7485 ( .INP(n7623), .Z(n7502) );
  NBUFFX2 U7486 ( .INP(n7623), .Z(n7501) );
  NBUFFX2 U7487 ( .INP(n7635), .Z(n7466) );
  NBUFFX2 U7488 ( .INP(n7624), .Z(n7498) );
  NBUFFX2 U7489 ( .INP(n7622), .Z(n7504) );
  NBUFFX2 U7490 ( .INP(n7622), .Z(n7503) );
  NBUFFX2 U7491 ( .INP(n7624), .Z(n7497) );
  NBUFFX2 U7492 ( .INP(n7625), .Z(n7496) );
  NBUFFX2 U7493 ( .INP(n7625), .Z(n7495) );
  NBUFFX2 U7494 ( .INP(n7625), .Z(n7494) );
  NBUFFX2 U7495 ( .INP(n7626), .Z(n7493) );
  NBUFFX2 U7496 ( .INP(n7626), .Z(n7492) );
  NBUFFX2 U7497 ( .INP(n7634), .Z(n7468) );
  NBUFFX2 U7498 ( .INP(n7633), .Z(n7471) );
  NBUFFX2 U7499 ( .INP(n7634), .Z(n7469) );
  NBUFFX2 U7500 ( .INP(n7633), .Z(n7470) );
  NBUFFX2 U7501 ( .INP(n7593), .Z(n7591) );
  NBUFFX2 U7502 ( .INP(n7593), .Z(n7590) );
  NBUFFX2 U7503 ( .INP(n7594), .Z(n7589) );
  NBUFFX2 U7504 ( .INP(n7594), .Z(n7588) );
  NBUFFX2 U7505 ( .INP(n7622), .Z(n7505) );
  NBUFFX2 U7506 ( .INP(n7627), .Z(n7490) );
  NBUFFX2 U7507 ( .INP(n7627), .Z(n7489) );
  NBUFFX2 U7508 ( .INP(n7627), .Z(n7488) );
  NBUFFX2 U7509 ( .INP(n7628), .Z(n7486) );
  NBUFFX2 U7510 ( .INP(n7632), .Z(n7473) );
  NBUFFX2 U7511 ( .INP(n7633), .Z(n7472) );
  NBUFFX2 U7512 ( .INP(n7635), .Z(n7465) );
  NBUFFX2 U7513 ( .INP(n7635), .Z(n7464) );
  NBUFFX2 U7514 ( .INP(n7406), .Z(n7405) );
  NBUFFX2 U7515 ( .INP(n7593), .Z(n7592) );
  NBUFFX2 U7516 ( .INP(n7645), .Z(n7595) );
  NBUFFX2 U7517 ( .INP(n7458), .Z(n7408) );
  NBUFFX2 U7518 ( .INP(n7645), .Z(n7596) );
  NBUFFX2 U7519 ( .INP(n7458), .Z(n7409) );
  NBUFFX2 U7520 ( .INP(n7645), .Z(n7593) );
  NBUFFX2 U7521 ( .INP(n7458), .Z(n7406) );
  NBUFFX2 U7522 ( .INP(n7645), .Z(n7594) );
  NBUFFX2 U7523 ( .INP(n7458), .Z(n7407) );
  NBUFFX2 U7524 ( .INP(n7641), .Z(n7615) );
  NBUFFX2 U7525 ( .INP(n7454), .Z(n7428) );
  NBUFFX2 U7526 ( .INP(n7644), .Z(n7598) );
  NBUFFX2 U7527 ( .INP(n7457), .Z(n7411) );
  NBUFFX2 U7528 ( .INP(n7644), .Z(n7599) );
  NBUFFX2 U7529 ( .INP(n7457), .Z(n7412) );
  NBUFFX2 U7530 ( .INP(n7644), .Z(n7597) );
  NBUFFX2 U7531 ( .INP(n7457), .Z(n7410) );
  NBUFFX2 U7532 ( .INP(n7644), .Z(n7601) );
  NBUFFX2 U7533 ( .INP(n7457), .Z(n7414) );
  NBUFFX2 U7534 ( .INP(n7644), .Z(n7600) );
  NBUFFX2 U7535 ( .INP(n7457), .Z(n7413) );
  NBUFFX2 U7536 ( .INP(n7643), .Z(n7602) );
  NBUFFX2 U7537 ( .INP(n7456), .Z(n7415) );
  NBUFFX2 U7538 ( .INP(n7643), .Z(n7603) );
  NBUFFX2 U7539 ( .INP(n7456), .Z(n7416) );
  NBUFFX2 U7540 ( .INP(n7643), .Z(n7604) );
  NBUFFX2 U7541 ( .INP(n7456), .Z(n7417) );
  NBUFFX2 U7542 ( .INP(n7643), .Z(n7605) );
  NBUFFX2 U7543 ( .INP(n7456), .Z(n7418) );
  NBUFFX2 U7544 ( .INP(n7643), .Z(n7606) );
  NBUFFX2 U7545 ( .INP(n7456), .Z(n7419) );
  NBUFFX2 U7546 ( .INP(n7642), .Z(n7608) );
  NBUFFX2 U7547 ( .INP(n7455), .Z(n7421) );
  NBUFFX2 U7548 ( .INP(n7642), .Z(n7607) );
  NBUFFX2 U7549 ( .INP(n7455), .Z(n7420) );
  NBUFFX2 U7550 ( .INP(n7642), .Z(n7609) );
  NBUFFX2 U7551 ( .INP(n7455), .Z(n7422) );
  NBUFFX2 U7552 ( .INP(n7642), .Z(n7610) );
  NBUFFX2 U7553 ( .INP(n7455), .Z(n7423) );
  NBUFFX2 U7554 ( .INP(n7642), .Z(n7611) );
  NBUFFX2 U7555 ( .INP(n7455), .Z(n7424) );
  NBUFFX2 U7556 ( .INP(n7641), .Z(n7612) );
  NBUFFX2 U7557 ( .INP(n7454), .Z(n7425) );
  NBUFFX2 U7558 ( .INP(n7640), .Z(n7620) );
  NBUFFX2 U7559 ( .INP(n7453), .Z(n7433) );
  NBUFFX2 U7560 ( .INP(n7638), .Z(n7629) );
  NBUFFX2 U7561 ( .INP(n7451), .Z(n7442) );
  NBUFFX2 U7562 ( .INP(n7638), .Z(n7630) );
  NBUFFX2 U7563 ( .INP(n7451), .Z(n7443) );
  NBUFFX2 U7564 ( .INP(n7638), .Z(n7631) );
  NBUFFX2 U7565 ( .INP(n7451), .Z(n7444) );
  NBUFFX2 U7566 ( .INP(n7641), .Z(n7616) );
  NBUFFX2 U7567 ( .INP(n7454), .Z(n7429) );
  NBUFFX2 U7568 ( .INP(n7640), .Z(n7617) );
  NBUFFX2 U7569 ( .INP(n7453), .Z(n7430) );
  NBUFFX2 U7570 ( .INP(n7640), .Z(n7621) );
  NBUFFX2 U7571 ( .INP(n7453), .Z(n7434) );
  NBUFFX2 U7572 ( .INP(n7641), .Z(n7613) );
  NBUFFX2 U7573 ( .INP(n7454), .Z(n7426) );
  NBUFFX2 U7574 ( .INP(n7641), .Z(n7614) );
  NBUFFX2 U7575 ( .INP(n7454), .Z(n7427) );
  NBUFFX2 U7576 ( .INP(n7640), .Z(n7618) );
  NBUFFX2 U7577 ( .INP(n7453), .Z(n7431) );
  NBUFFX2 U7578 ( .INP(n7640), .Z(n7619) );
  NBUFFX2 U7579 ( .INP(n7453), .Z(n7432) );
  NBUFFX2 U7580 ( .INP(n7639), .Z(n7623) );
  NBUFFX2 U7581 ( .INP(n7452), .Z(n7436) );
  NBUFFX2 U7582 ( .INP(n7639), .Z(n7624) );
  NBUFFX2 U7583 ( .INP(n7452), .Z(n7437) );
  NBUFFX2 U7584 ( .INP(n7639), .Z(n7625) );
  NBUFFX2 U7585 ( .INP(n7452), .Z(n7438) );
  NBUFFX2 U7586 ( .INP(n7639), .Z(n7626) );
  NBUFFX2 U7587 ( .INP(n7452), .Z(n7439) );
  NBUFFX2 U7588 ( .INP(n7637), .Z(n7634) );
  NBUFFX2 U7589 ( .INP(n7450), .Z(n7447) );
  NBUFFX2 U7590 ( .INP(n7639), .Z(n7622) );
  NBUFFX2 U7591 ( .INP(n7452), .Z(n7435) );
  NBUFFX2 U7592 ( .INP(n7638), .Z(n7627) );
  NBUFFX2 U7593 ( .INP(n7451), .Z(n7440) );
  NBUFFX2 U7594 ( .INP(n7638), .Z(n7628) );
  NBUFFX2 U7595 ( .INP(n7451), .Z(n7441) );
  NBUFFX2 U7596 ( .INP(n7637), .Z(n7632) );
  NBUFFX2 U7597 ( .INP(n7450), .Z(n7445) );
  NBUFFX2 U7598 ( .INP(n7637), .Z(n7633) );
  NBUFFX2 U7599 ( .INP(n7450), .Z(n7446) );
  NBUFFX2 U7600 ( .INP(n7637), .Z(n7635) );
  NBUFFX2 U7601 ( .INP(n7450), .Z(n7448) );
  NBUFFX2 U7602 ( .INP(n7637), .Z(n7636) );
  NBUFFX2 U7603 ( .INP(n7450), .Z(n7449) );
  NBUFFX2 U7604 ( .INP(n7461), .Z(n7450) );
  NBUFFX2 U7605 ( .INP(n7461), .Z(n7451) );
  NBUFFX2 U7606 ( .INP(n7461), .Z(n7452) );
  NBUFFX2 U7607 ( .INP(n7460), .Z(n7453) );
  NBUFFX2 U7608 ( .INP(n7460), .Z(n7454) );
  NBUFFX2 U7609 ( .INP(n7460), .Z(n7455) );
  NBUFFX2 U7610 ( .INP(n7459), .Z(n7456) );
  NBUFFX2 U7611 ( .INP(n7459), .Z(n7457) );
  NBUFFX2 U7612 ( .INP(n7459), .Z(n7458) );
  NBUFFX2 U7613 ( .INP(test_se), .Z(n7459) );
  NBUFFX2 U7614 ( .INP(test_se), .Z(n7460) );
  NBUFFX2 U7615 ( .INP(test_se), .Z(n7461) );
  NBUFFX2 U7616 ( .INP(n7648), .Z(n7637) );
  NBUFFX2 U7617 ( .INP(n7648), .Z(n7638) );
  NBUFFX2 U7618 ( .INP(n7648), .Z(n7639) );
  NBUFFX2 U7619 ( .INP(n7647), .Z(n7640) );
  NBUFFX2 U7620 ( .INP(n7647), .Z(n7641) );
  NBUFFX2 U7621 ( .INP(n7647), .Z(n7642) );
  NBUFFX2 U7622 ( .INP(n7646), .Z(n7643) );
  NBUFFX2 U7623 ( .INP(n7646), .Z(n7644) );
  NBUFFX2 U7624 ( .INP(n7646), .Z(n7645) );
  NBUFFX2 U7625 ( .INP(CK), .Z(n7646) );
  NBUFFX2 U7626 ( .INP(CK), .Z(n7647) );
  NBUFFX2 U7627 ( .INP(CK), .Z(n7648) );
  INVX0 U7628 ( .INP(n7649), .ZN(n765) );
  INVX0 U7629 ( .INP(n7650), .ZN(n758) );
  INVX0 U7630 ( .INP(n7651), .ZN(n63) );
  INVX0 U7631 ( .INP(n7652), .ZN(n605) );
  INVX0 U7632 ( .INP(n7653), .ZN(n598) );
  INVX0 U7633 ( .INP(n7654), .ZN(n440) );
  INVX0 U7634 ( .INP(n7655), .ZN(n433) );
  XNOR2X1 U7635 ( .IN1(n7260), .IN2(n7656), .Q(n4281) );
  XOR2X1 U7636 ( .IN1(n7657), .IN2(n7262), .Q(n4280) );
  NAND2X0 U7637 ( .IN1(g2879), .IN2(n7658), .QN(n4279) );
  NAND2X0 U7638 ( .IN1(DFF_18_n1), .IN2(g8021), .QN(n7658) );
  NOR2X0 U7639 ( .IN1(n7659), .IN2(n7660), .QN(n4278) );
  NOR2X0 U7640 ( .IN1(n7661), .IN2(n7662), .QN(n7660) );
  NOR2X0 U7641 ( .IN1(n7663), .IN2(n7664), .QN(n7659) );
  NAND4X0 U7642 ( .IN1(n7665), .IN2(n7666), .IN3(n7667), .IN4(n7668), .QN(
        n7664) );
  NOR3X0 U7643 ( .IN1(n7669), .IN2(n7670), .IN3(n7671), .QN(n7668) );
  XOR2X1 U7644 ( .IN1(n6991), .IN2(n7672), .Q(n7671) );
  XNOR2X1 U7645 ( .IN1(n6971), .IN2(n7673), .Q(n7670) );
  XOR2X1 U7646 ( .IN1(n6977), .IN2(n7674), .Q(n7669) );
  XOR2X1 U7647 ( .IN1(n6975), .IN2(n7675), .Q(n7667) );
  XNOR2X1 U7648 ( .IN1(n6994), .IN2(n4513), .Q(n7666) );
  XNOR2X1 U7649 ( .IN1(n6439), .IN2(n7676), .Q(n7665) );
  NAND4X0 U7650 ( .IN1(n7677), .IN2(n7678), .IN3(n7679), .IN4(n7680), .QN(
        n7663) );
  NOR3X0 U7651 ( .IN1(n7681), .IN2(n7682), .IN3(n7683), .QN(n7680) );
  XOR2X1 U7652 ( .IN1(n6992), .IN2(n7684), .Q(n7683) );
  XOR2X1 U7653 ( .IN1(n6600), .IN2(n7685), .Q(n7682) );
  XOR2X1 U7654 ( .IN1(n6993), .IN2(n7686), .Q(n7681) );
  XOR2X1 U7655 ( .IN1(test_so15), .IN2(n7687), .Q(n7679) );
  NOR2X0 U7656 ( .IN1(n7688), .IN2(n7689), .QN(n4277) );
  NOR2X0 U7657 ( .IN1(n7690), .IN2(n7691), .QN(n7689) );
  NOR4X0 U7658 ( .IN1(n7692), .IN2(n7693), .IN3(n7694), .IN4(n7695), .QN(n7688) );
  NAND3X0 U7659 ( .IN1(n7696), .IN2(n7697), .IN3(n7698), .QN(n7695) );
  XNOR2X1 U7660 ( .IN1(n7699), .IN2(n6989), .Q(n7698) );
  XOR2X1 U7661 ( .IN1(n7700), .IN2(n6599), .Q(n7697) );
  XOR2X1 U7662 ( .IN1(n7701), .IN2(n6438), .Q(n7696) );
  NAND3X0 U7663 ( .IN1(n7702), .IN2(n7703), .IN3(n7704), .QN(n7694) );
  XOR2X1 U7664 ( .IN1(n7705), .IN2(g758), .Q(n7704) );
  XOR2X1 U7665 ( .IN1(n7706), .IN2(n6988), .Q(n7703) );
  XOR2X1 U7666 ( .IN1(n7707), .IN2(n6987), .Q(n7702) );
  NAND3X0 U7667 ( .IN1(n7708), .IN2(n7709), .IN3(n7710), .QN(n7693) );
  XOR2X1 U7668 ( .IN1(n7711), .IN2(n6990), .Q(n7710) );
  XOR2X1 U7669 ( .IN1(n7712), .IN2(n6978), .Q(n7709) );
  XOR2X1 U7670 ( .IN1(n7713), .IN2(n6435), .Q(n7708) );
  NAND3X0 U7671 ( .IN1(n7714), .IN2(n7678), .IN3(n7715), .QN(n7692) );
  XNOR2X1 U7672 ( .IN1(test_so36), .IN2(n7716), .Q(n7715) );
  NOR2X0 U7673 ( .IN1(n7717), .IN2(n7718), .QN(n4276) );
  NOR2X0 U7674 ( .IN1(n7719), .IN2(n7720), .QN(n7718) );
  NOR2X0 U7675 ( .IN1(n7721), .IN2(n7722), .QN(n7717) );
  NAND4X0 U7676 ( .IN1(n7723), .IN2(n7724), .IN3(n7725), .IN4(n7726), .QN(
        n7722) );
  NOR3X0 U7677 ( .IN1(n7727), .IN2(n7728), .IN3(n7729), .QN(n7726) );
  XOR2X1 U7678 ( .IN1(n6983), .IN2(n7730), .Q(n7729) );
  XNOR2X1 U7679 ( .IN1(n6970), .IN2(n7731), .Q(n7728) );
  XOR2X1 U7680 ( .IN1(n6976), .IN2(n7732), .Q(n7727) );
  XOR2X1 U7681 ( .IN1(n6434), .IN2(n7733), .Q(n7725) );
  XOR2X1 U7682 ( .IN1(n6973), .IN2(n7734), .Q(n7724) );
  XNOR2X1 U7683 ( .IN1(n6437), .IN2(n7735), .Q(n7723) );
  NAND4X0 U7684 ( .IN1(n7736), .IN2(n7678), .IN3(n7737), .IN4(n7738), .QN(
        n7721) );
  NOR3X0 U7685 ( .IN1(n7739), .IN2(n7740), .IN3(n7741), .QN(n7738) );
  XOR2X1 U7686 ( .IN1(n6985), .IN2(n7742), .Q(n7741) );
  XNOR2X1 U7687 ( .IN1(n6986), .IN2(n7743), .Q(n7740) );
  XOR2X1 U7688 ( .IN1(n6598), .IN2(n7744), .Q(n7739) );
  XOR2X1 U7689 ( .IN1(n6984), .IN2(n7745), .Q(n7737) );
  NOR2X0 U7690 ( .IN1(n7746), .IN2(n7747), .QN(n4275) );
  NOR2X0 U7691 ( .IN1(n7748), .IN2(n7749), .QN(n7747) );
  NOR4X0 U7692 ( .IN1(n7750), .IN2(n7751), .IN3(n7752), .IN4(n7753), .QN(n7746) );
  NAND3X0 U7693 ( .IN1(n7754), .IN2(n7755), .IN3(n7756), .QN(n7753) );
  XOR2X1 U7694 ( .IN1(n7757), .IN2(n6433), .Q(n7756) );
  XOR2X1 U7695 ( .IN1(n7758), .IN2(n6972), .Q(n7755) );
  XNOR2X1 U7696 ( .IN1(n7759), .IN2(n6436), .Q(n7754) );
  NAND3X0 U7697 ( .IN1(n7760), .IN2(n7761), .IN3(n7762), .QN(n7752) );
  XOR2X1 U7698 ( .IN1(n7763), .IN2(n6979), .Q(n7762) );
  XOR2X1 U7699 ( .IN1(n7764), .IN2(n6969), .Q(n7761) );
  XNOR2X1 U7700 ( .IN1(n7765), .IN2(n6982), .Q(n7760) );
  NAND3X0 U7701 ( .IN1(n7766), .IN2(n7767), .IN3(n7768), .QN(n7751) );
  XOR2X1 U7702 ( .IN1(n7769), .IN2(n6981), .Q(n7768) );
  XOR2X1 U7703 ( .IN1(n7770), .IN2(n6597), .Q(n7767) );
  XOR2X1 U7704 ( .IN1(n7771), .IN2(n6980), .Q(n7766) );
  NAND3X0 U7705 ( .IN1(n7772), .IN2(n7678), .IN3(n7773), .QN(n7750) );
  XOR2X1 U7706 ( .IN1(test_so78), .IN2(n7774), .Q(n7773) );
  NAND2X0 U7707 ( .IN1(n7775), .IN2(n7776), .QN(n4274) );
  INVX0 U7708 ( .INP(n7777), .ZN(n7776) );
  XNOR2X1 U7709 ( .IN1(n4330), .IN2(n4423), .Q(n7775) );
  NAND2X0 U7710 ( .IN1(n7778), .IN2(n7779), .QN(n4273) );
  NAND2X0 U7711 ( .IN1(n7780), .IN2(n7781), .QN(n7779) );
  NAND2X0 U7712 ( .IN1(n4482), .IN2(n7782), .QN(n7780) );
  NAND2X0 U7713 ( .IN1(n2426), .IN2(n7783), .QN(n4272) );
  NAND3X0 U7714 ( .IN1(n7784), .IN2(n7785), .IN3(n7786), .QN(n7783) );
  OR2X1 U7715 ( .IN1(n7787), .IN2(n7788), .Q(n7785) );
  NAND2X0 U7716 ( .IN1(n7789), .IN2(DFF_449_n1), .QN(n7784) );
  NAND2X0 U7717 ( .IN1(n7790), .IN2(n7791), .QN(n4271) );
  NAND2X0 U7718 ( .IN1(n2446), .IN2(n7792), .QN(n7791) );
  NAND3X0 U7719 ( .IN1(n7793), .IN2(n7794), .IN3(n7786), .QN(n7790) );
  OR2X1 U7720 ( .IN1(n7795), .IN2(n7788), .Q(n7794) );
  NAND2X0 U7721 ( .IN1(n6409), .IN2(n7789), .QN(n7793) );
  NAND2X0 U7722 ( .IN1(n7796), .IN2(n7797), .QN(n4270) );
  NAND2X0 U7723 ( .IN1(n2446), .IN2(n7798), .QN(n7797) );
  NAND3X0 U7724 ( .IN1(n7799), .IN2(n7800), .IN3(n7786), .QN(n7796) );
  NAND2X0 U7725 ( .IN1(n7801), .IN2(n7802), .QN(n7800) );
  NAND2X0 U7726 ( .IN1(n6408), .IN2(n7789), .QN(n7799) );
  NAND2X0 U7727 ( .IN1(n7803), .IN2(n7804), .QN(n4269) );
  NAND3X0 U7728 ( .IN1(n7805), .IN2(n7806), .IN3(n7786), .QN(n7804) );
  OR2X1 U7729 ( .IN1(n7807), .IN2(n7788), .Q(n7806) );
  NAND2X0 U7730 ( .IN1(n7789), .IN2(DFF_444_n1), .QN(n7805) );
  NAND3X0 U7731 ( .IN1(n2426), .IN2(n7808), .IN3(n2440), .QN(n4268) );
  NAND3X0 U7732 ( .IN1(n7809), .IN2(n7810), .IN3(n7786), .QN(n7808) );
  OR2X1 U7733 ( .IN1(n7811), .IN2(n7788), .Q(n7810) );
  NAND2X0 U7734 ( .IN1(n7789), .IN2(DFF_445_n1), .QN(n7809) );
  NAND3X0 U7735 ( .IN1(n2426), .IN2(n7812), .IN3(n2440), .QN(n4267) );
  NAND3X0 U7736 ( .IN1(n7813), .IN2(n7814), .IN3(n7786), .QN(n7812) );
  OR2X1 U7737 ( .IN1(n7815), .IN2(n7788), .Q(n7814) );
  NAND2X0 U7738 ( .IN1(n7789), .IN2(DFF_446_n1), .QN(n7813) );
  NAND2X0 U7739 ( .IN1(n7803), .IN2(n7816), .QN(n4266) );
  NAND3X0 U7740 ( .IN1(n7817), .IN2(n7818), .IN3(n7786), .QN(n7816) );
  NAND2X0 U7741 ( .IN1(n7819), .IN2(n7802), .QN(n7818) );
  NAND2X0 U7742 ( .IN1(n7789), .IN2(DFF_447_n1), .QN(n7817) );
  AND2X1 U7743 ( .IN1(n2426), .IN2(n7820), .Q(n7803) );
  NAND2X0 U7744 ( .IN1(n2446), .IN2(n2445), .QN(n7820) );
  NAND2X0 U7745 ( .IN1(n2426), .IN2(n7821), .QN(n4265) );
  NAND3X0 U7746 ( .IN1(n7822), .IN2(n7823), .IN3(n7786), .QN(n7821) );
  OR2X1 U7747 ( .IN1(n7824), .IN2(n7788), .Q(n7823) );
  NAND2X0 U7748 ( .IN1(n7789), .IN2(DFF_448_n1), .QN(n7822) );
  NAND2X0 U7749 ( .IN1(DFF_1562_n1), .IN2(n7825), .QN(n4263) );
  NAND2X0 U7750 ( .IN1(n7826), .IN2(n7827), .QN(n4262) );
  XOR2X1 U7751 ( .IN1(n4481), .IN2(n7828), .Q(n7826) );
  XNOR2X1 U7752 ( .IN1(n7829), .IN2(n7830), .Q(n4261) );
  XOR2X1 U7753 ( .IN1(n7830), .IN2(n7831), .Q(n4260) );
  INVX0 U7754 ( .INP(n7832), .ZN(n7831) );
  NOR2X0 U7755 ( .IN1(g3231), .IN2(n13233), .QN(n7830) );
  NAND3X0 U7756 ( .IN1(n7833), .IN2(n7834), .IN3(n7835), .QN(n4259) );
  NAND2X0 U7757 ( .IN1(test_so22), .IN2(n7836), .QN(n7835) );
  XOR2X1 U7758 ( .IN1(n7837), .IN2(n7838), .Q(n7836) );
  XOR3X1 U7759 ( .IN1(n7795), .IN2(n7787), .IN3(n7839), .Q(n7838) );
  XOR2X1 U7760 ( .IN1(n7824), .IN2(n7801), .Q(n7839) );
  AND3X1 U7761 ( .IN1(n7840), .IN2(n7841), .IN3(n7842), .Q(n7801) );
  NAND2X0 U7762 ( .IN1(n7843), .IN2(n7844), .QN(n7841) );
  NAND2X0 U7763 ( .IN1(n7845), .IN2(n7846), .QN(n7840) );
  NAND3X0 U7764 ( .IN1(n7847), .IN2(n7848), .IN3(n7849), .QN(n7824) );
  NAND2X0 U7765 ( .IN1(n7850), .IN2(n7851), .QN(n7848) );
  NAND2X0 U7766 ( .IN1(n7852), .IN2(n7853), .QN(n7847) );
  NAND3X0 U7767 ( .IN1(n7854), .IN2(n7855), .IN3(n7856), .QN(n7787) );
  NAND2X0 U7768 ( .IN1(n7857), .IN2(n7844), .QN(n7855) );
  NAND2X0 U7769 ( .IN1(n7845), .IN2(n7858), .QN(n7854) );
  NAND3X0 U7770 ( .IN1(n7859), .IN2(n7860), .IN3(n7849), .QN(n7795) );
  NAND2X0 U7771 ( .IN1(n7861), .IN2(n7851), .QN(n7860) );
  NAND2X0 U7772 ( .IN1(n7852), .IN2(n7862), .QN(n7859) );
  XOR3X1 U7773 ( .IN1(n7815), .IN2(n7807), .IN3(n7863), .Q(n7837) );
  XOR2X1 U7774 ( .IN1(n7811), .IN2(n7819), .Q(n7863) );
  AND3X1 U7775 ( .IN1(n7864), .IN2(n7865), .IN3(n7842), .Q(n7819) );
  NAND2X0 U7776 ( .IN1(n7866), .IN2(n7844), .QN(n7865) );
  NAND2X0 U7777 ( .IN1(n7845), .IN2(n7867), .QN(n7864) );
  NAND3X0 U7778 ( .IN1(n7868), .IN2(n7869), .IN3(n7842), .QN(n7811) );
  NAND2X0 U7779 ( .IN1(n7870), .IN2(n7844), .QN(n7869) );
  NAND2X0 U7780 ( .IN1(n7845), .IN2(n7871), .QN(n7868) );
  NAND3X0 U7781 ( .IN1(n7872), .IN2(n7873), .IN3(n7842), .QN(n7807) );
  NAND2X0 U7782 ( .IN1(n7874), .IN2(n7851), .QN(n7873) );
  NAND2X0 U7783 ( .IN1(n7852), .IN2(n7875), .QN(n7872) );
  NAND3X0 U7784 ( .IN1(n7876), .IN2(n7877), .IN3(n7842), .QN(n7815) );
  NAND2X0 U7785 ( .IN1(n7878), .IN2(n7851), .QN(n7877) );
  NAND2X0 U7786 ( .IN1(n7852), .IN2(n7879), .QN(n7876) );
  NAND4X0 U7787 ( .IN1(n7786), .IN2(n7789), .IN3(n7880), .IN4(n7881), .QN(
        n7834) );
  NAND2X0 U7788 ( .IN1(n13227), .IN2(n7882), .QN(n7881) );
  NAND2X0 U7789 ( .IN1(n4492), .IN2(g3229), .QN(n7880) );
  AND2X1 U7790 ( .IN1(n7788), .IN2(n2478), .Q(n7789) );
  INVX0 U7791 ( .INP(n7802), .ZN(n7788) );
  NAND2X0 U7792 ( .IN1(n7883), .IN2(g557), .QN(n7833) );
  XOR2X1 U7793 ( .IN1(n7792), .IN2(n7798), .Q(n7883) );
  NAND3X0 U7794 ( .IN1(n7884), .IN2(n7885), .IN3(n7856), .QN(n7798) );
  AND2X1 U7795 ( .IN1(n7842), .IN2(n7886), .Q(n7856) );
  NAND2X0 U7796 ( .IN1(n7887), .IN2(n7844), .QN(n7886) );
  NAND2X0 U7797 ( .IN1(n7888), .IN2(n7844), .QN(n7885) );
  NAND2X0 U7798 ( .IN1(n7845), .IN2(n7889), .QN(n7884) );
  NOR2X0 U7799 ( .IN1(n7844), .IN2(n7887), .QN(n7845) );
  NAND3X0 U7800 ( .IN1(n7890), .IN2(n7891), .IN3(n7849), .QN(n7792) );
  AND2X1 U7801 ( .IN1(n7842), .IN2(n2430), .Q(n7849) );
  AND2X1 U7802 ( .IN1(n2478), .IN2(g499), .Q(n7842) );
  NAND2X0 U7803 ( .IN1(n7892), .IN2(n7851), .QN(n7891) );
  NAND2X0 U7804 ( .IN1(n7852), .IN2(n7893), .QN(n7890) );
  NOR2X0 U7805 ( .IN1(n7851), .IN2(n7887), .QN(n7852) );
  NAND2X0 U7806 ( .IN1(n7894), .IN2(n7895), .QN(n4258) );
  NAND2X0 U7807 ( .IN1(n2361), .IN2(n7896), .QN(n7895) );
  NAND3X0 U7808 ( .IN1(n7897), .IN2(n7898), .IN3(n7899), .QN(n7894) );
  NAND2X0 U7809 ( .IN1(n7900), .IN2(n7901), .QN(n7898) );
  NAND2X0 U7810 ( .IN1(n6410), .IN2(n7902), .QN(n7897) );
  NAND3X0 U7811 ( .IN1(n7903), .IN2(n7904), .IN3(n2375), .QN(n4257) );
  NAND3X0 U7812 ( .IN1(n7905), .IN2(n7906), .IN3(n7899), .QN(n7903) );
  NAND2X0 U7813 ( .IN1(n7908), .IN2(n7901), .QN(n7906) );
  NAND2X0 U7814 ( .IN1(n7902), .IN2(DFF_1495_n1), .QN(n7905) );
  NAND2X0 U7815 ( .IN1(n7904), .IN2(n7910), .QN(n4256) );
  NAND3X0 U7816 ( .IN1(n7911), .IN2(n7914), .IN3(n7899), .QN(n7910) );
  NAND2X0 U7817 ( .IN1(n7915), .IN2(n7901), .QN(n7914) );
  NAND2X0 U7818 ( .IN1(n7902), .IN2(DFF_1499_n1), .QN(n7911) );
  NAND3X0 U7819 ( .IN1(n7916), .IN2(n7904), .IN3(n2375), .QN(n4255) );
  NAND3X0 U7820 ( .IN1(n7917), .IN2(n7919), .IN3(n7899), .QN(n7916) );
  NAND2X0 U7821 ( .IN1(n7927), .IN2(n7901), .QN(n7919) );
  NAND2X0 U7822 ( .IN1(n7902), .IN2(DFF_1496_n1), .QN(n7917) );
  NAND2X0 U7823 ( .IN1(n7928), .IN2(n7931), .QN(n4254) );
  NAND3X0 U7824 ( .IN1(n7932), .IN2(n7933), .IN3(n7899), .QN(n7931) );
  NAND2X0 U7825 ( .IN1(n7934), .IN2(n7901), .QN(n7933) );
  NAND2X0 U7826 ( .IN1(n7902), .IN2(DFF_1494_n1), .QN(n7932) );
  NAND2X0 U7827 ( .IN1(n7935), .IN2(n7939), .QN(n4253) );
  NAND2X0 U7828 ( .IN1(n2361), .IN2(n7947), .QN(n7939) );
  NAND3X0 U7829 ( .IN1(n7948), .IN2(n7949), .IN3(n7899), .QN(n7935) );
  NAND2X0 U7830 ( .IN1(n7950), .IN2(n7901), .QN(n7949) );
  NAND2X0 U7831 ( .IN1(n7902), .IN2(n6411), .QN(n7948) );
  NAND2X0 U7832 ( .IN1(n7928), .IN2(n7951), .QN(n4252) );
  NAND3X0 U7833 ( .IN1(n7952), .IN2(n7953), .IN3(n7899), .QN(n7951) );
  NAND2X0 U7834 ( .IN1(n7954), .IN2(n7901), .QN(n7953) );
  NAND2X0 U7835 ( .IN1(n7902), .IN2(DFF_1497_n1), .QN(n7952) );
  AND2X1 U7836 ( .IN1(n7904), .IN2(n7955), .Q(n7928) );
  NAND2X0 U7837 ( .IN1(n2361), .IN2(n2374), .QN(n7955) );
  NAND2X0 U7838 ( .IN1(n7904), .IN2(n7956), .QN(n4251) );
  NAND3X0 U7839 ( .IN1(n7957), .IN2(n7958), .IN3(n7899), .QN(n7956) );
  NAND2X0 U7840 ( .IN1(n7959), .IN2(n7901), .QN(n7958) );
  NAND2X0 U7841 ( .IN1(n7902), .IN2(DFF_1498_n1), .QN(n7957) );
  NAND2X0 U7842 ( .IN1(n2361), .IN2(n7961), .QN(n7904) );
  NAND3X0 U7843 ( .IN1(n7969), .IN2(n7970), .IN3(n7972), .QN(n4250) );
  NAND2X0 U7844 ( .IN1(n7973), .IN2(g2631), .QN(n7972) );
  XOR2X1 U7845 ( .IN1(n7896), .IN2(n7947), .Q(n7973) );
  NAND4X0 U7846 ( .IN1(n7974), .IN2(n2351), .IN3(n7975), .IN4(n7976), .QN(
        n7947) );
  NAND2X0 U7847 ( .IN1(n7977), .IN2(n7981), .QN(n7976) );
  NAND2X0 U7848 ( .IN1(n7982), .IN2(n7989), .QN(n7975) );
  NAND4X0 U7849 ( .IN1(n7974), .IN2(n7990), .IN3(n7991), .IN4(n7992), .QN(
        n7896) );
  NAND2X0 U7850 ( .IN1(n7993), .IN2(n7994), .QN(n7992) );
  NAND2X0 U7851 ( .IN1(n7995), .IN2(n7996), .QN(n7991) );
  NAND4X0 U7852 ( .IN1(n7899), .IN2(n7902), .IN3(n7997), .IN4(n7998), .QN(
        n7970) );
  NAND2X0 U7853 ( .IN1(n13228), .IN2(n7882), .QN(n7998) );
  NAND2X0 U7854 ( .IN1(n4490), .IN2(g3229), .QN(n7997) );
  NOR2X0 U7855 ( .IN1(n7961), .IN2(n7901), .QN(n7902) );
  NAND2X0 U7856 ( .IN1(n7999), .IN2(g2584), .QN(n7969) );
  XOR2X1 U7857 ( .IN1(n8000), .IN2(n8001), .Q(n7999) );
  XNOR3X1 U7858 ( .IN1(n7934), .IN2(n7959), .IN3(n8002), .Q(n8001) );
  XNOR2X1 U7859 ( .IN1(n7915), .IN2(n7927), .Q(n8002) );
  AND3X1 U7860 ( .IN1(n8010), .IN2(n8011), .IN3(n7974), .Q(n7927) );
  NAND2X0 U7861 ( .IN1(n8012), .IN2(n7981), .QN(n8011) );
  NAND2X0 U7862 ( .IN1(n7982), .IN2(n8013), .QN(n8010) );
  AND4X1 U7863 ( .IN1(n7974), .IN2(n7990), .IN3(n8014), .IN4(n8015), .Q(n7915)
         );
  NAND2X0 U7864 ( .IN1(n8016), .IN2(n7994), .QN(n8015) );
  NAND2X0 U7865 ( .IN1(n7995), .IN2(n8022), .QN(n8014) );
  NAND2X0 U7866 ( .IN1(n8023), .IN2(n7994), .QN(n7990) );
  AND4X1 U7867 ( .IN1(n7974), .IN2(n2351), .IN3(n8028), .IN4(n8029), .Q(n7959)
         );
  NAND2X0 U7868 ( .IN1(n8030), .IN2(n7981), .QN(n8029) );
  NAND2X0 U7869 ( .IN1(n7982), .IN2(n8031), .QN(n8028) );
  AND3X1 U7870 ( .IN1(n8032), .IN2(n8033), .IN3(n7974), .Q(n7934) );
  NAND2X0 U7871 ( .IN1(n8034), .IN2(n7981), .QN(n8033) );
  NAND2X0 U7872 ( .IN1(n7982), .IN2(n8035), .QN(n8032) );
  XOR3X1 U7873 ( .IN1(n7908), .IN2(n7954), .IN3(n8036), .Q(n8000) );
  XOR2X1 U7874 ( .IN1(n7950), .IN2(n7900), .Q(n8036) );
  NAND2X0 U7875 ( .IN1(n8037), .IN2(n8038), .QN(n7900) );
  NAND2X0 U7876 ( .IN1(n8039), .IN2(n8041), .QN(n8038) );
  NAND2X0 U7877 ( .IN1(n8042), .IN2(n8048), .QN(n8037) );
  AND4X1 U7878 ( .IN1(n7974), .IN2(n2351), .IN3(n8049), .IN4(n8050), .Q(n7950)
         );
  NAND2X0 U7879 ( .IN1(n8051), .IN2(n7981), .QN(n8050) );
  NAND2X0 U7880 ( .IN1(n7982), .IN2(n8052), .QN(n8049) );
  NOR2X0 U7881 ( .IN1(n7981), .IN2(n8023), .QN(n7982) );
  NAND2X0 U7882 ( .IN1(n8053), .IN2(n8054), .QN(n7954) );
  NAND2X0 U7883 ( .IN1(n8039), .IN2(n8063), .QN(n8054) );
  NAND2X0 U7884 ( .IN1(n8042), .IN2(n8064), .QN(n8053) );
  NAND2X0 U7885 ( .IN1(n8067), .IN2(n8068), .QN(n7908) );
  NAND2X0 U7886 ( .IN1(n8039), .IN2(n8069), .QN(n8068) );
  NOR2X0 U7887 ( .IN1(n8070), .IN2(n7995), .QN(n8039) );
  NOR2X0 U7888 ( .IN1(n7994), .IN2(n8023), .QN(n7995) );
  NAND2X0 U7889 ( .IN1(n8042), .IN2(n8071), .QN(n8067) );
  NOR2X0 U7890 ( .IN1(n8070), .IN2(n7994), .QN(n8042) );
  INVX0 U7891 ( .INP(n7974), .ZN(n8070) );
  NOR2X0 U7892 ( .IN1(n7961), .IN2(n4543), .QN(n7974) );
  OR3X1 U7893 ( .IN1(g2637), .IN2(g30072), .IN3(g2633), .Q(n7961) );
  NAND2X0 U7894 ( .IN1(n8072), .IN2(n8073), .QN(n4249) );
  NAND2X0 U7895 ( .IN1(n2289), .IN2(n8074), .QN(n8073) );
  NAND3X0 U7896 ( .IN1(n8075), .IN2(n8085), .IN3(n8091), .QN(n8072) );
  NAND2X0 U7897 ( .IN1(n8092), .IN2(n8093), .QN(n8085) );
  NAND2X0 U7898 ( .IN1(n6412), .IN2(n8094), .QN(n8075) );
  NAND3X0 U7899 ( .IN1(n2275), .IN2(n8095), .IN3(n2303), .QN(n4248) );
  NAND3X0 U7900 ( .IN1(n8096), .IN2(n8097), .IN3(n8091), .QN(n8095) );
  NAND2X0 U7901 ( .IN1(n8100), .IN2(n8093), .QN(n8097) );
  NAND2X0 U7902 ( .IN1(n8094), .IN2(DFF_1145_n1), .QN(n8096) );
  NAND2X0 U7903 ( .IN1(n2275), .IN2(n8101), .QN(n4247) );
  NAND3X0 U7904 ( .IN1(n8105), .IN2(n8106), .IN3(n8091), .QN(n8101) );
  NAND2X0 U7905 ( .IN1(n8107), .IN2(n8093), .QN(n8106) );
  NAND2X0 U7906 ( .IN1(n8094), .IN2(DFF_1149_n1), .QN(n8105) );
  NAND3X0 U7907 ( .IN1(n2275), .IN2(n8108), .IN3(n2303), .QN(n4246) );
  NAND3X0 U7908 ( .IN1(n8109), .IN2(n8110), .IN3(n8091), .QN(n8108) );
  NAND2X0 U7909 ( .IN1(n8111), .IN2(n8093), .QN(n8110) );
  NAND2X0 U7910 ( .IN1(n8094), .IN2(DFF_1146_n1), .QN(n8109) );
  NAND2X0 U7911 ( .IN1(n8112), .IN2(n8113), .QN(n4245) );
  NAND3X0 U7912 ( .IN1(n8114), .IN2(n8115), .IN3(n8091), .QN(n8113) );
  NAND2X0 U7913 ( .IN1(n8116), .IN2(n8093), .QN(n8115) );
  NAND2X0 U7914 ( .IN1(n8094), .IN2(DFF_1144_n1), .QN(n8114) );
  NAND2X0 U7915 ( .IN1(n8117), .IN2(n8118), .QN(n4244) );
  NAND2X0 U7916 ( .IN1(n2289), .IN2(n8119), .QN(n8118) );
  NAND3X0 U7917 ( .IN1(n8120), .IN2(n8121), .IN3(n8091), .QN(n8117) );
  OR2X1 U7918 ( .IN1(n8122), .IN2(n8123), .Q(n8121) );
  NAND2X0 U7919 ( .IN1(n6413), .IN2(n8094), .QN(n8120) );
  NAND2X0 U7920 ( .IN1(n8112), .IN2(n8124), .QN(n4243) );
  NAND3X0 U7921 ( .IN1(n8125), .IN2(n8126), .IN3(n8091), .QN(n8124) );
  NAND2X0 U7922 ( .IN1(n8127), .IN2(n8093), .QN(n8126) );
  NAND2X0 U7923 ( .IN1(n8094), .IN2(DFF_1147_n1), .QN(n8125) );
  AND2X1 U7924 ( .IN1(n2275), .IN2(n8128), .Q(n8112) );
  NAND2X0 U7925 ( .IN1(n2289), .IN2(n2302), .QN(n8128) );
  NAND2X0 U7926 ( .IN1(n2275), .IN2(n8129), .QN(n4242) );
  NAND3X0 U7927 ( .IN1(n8130), .IN2(n8131), .IN3(n8091), .QN(n8129) );
  NAND2X0 U7928 ( .IN1(n8132), .IN2(n8093), .QN(n8131) );
  NAND2X0 U7929 ( .IN1(n8094), .IN2(DFF_1148_n1), .QN(n8130) );
  NAND3X0 U7930 ( .IN1(n8133), .IN2(n8134), .IN3(n8135), .QN(n4241) );
  NAND2X0 U7931 ( .IN1(n8136), .IN2(g1890), .QN(n8135) );
  XOR2X1 U7932 ( .IN1(n8137), .IN2(n8138), .Q(n8136) );
  XOR3X1 U7933 ( .IN1(n8116), .IN2(n8127), .IN3(n8139), .Q(n8138) );
  XOR2X1 U7934 ( .IN1(n8100), .IN2(n8111), .Q(n8139) );
  NAND2X0 U7935 ( .IN1(n8140), .IN2(n8141), .QN(n8111) );
  NAND3X0 U7936 ( .IN1(n8142), .IN2(n8143), .IN3(n8144), .QN(n8141) );
  NAND2X0 U7937 ( .IN1(n8145), .IN2(n8146), .QN(n8140) );
  NAND2X0 U7938 ( .IN1(n8147), .IN2(n8148), .QN(n8100) );
  NAND2X0 U7939 ( .IN1(n8149), .IN2(n8150), .QN(n8148) );
  NAND2X0 U7940 ( .IN1(n8151), .IN2(n8152), .QN(n8147) );
  NAND2X0 U7941 ( .IN1(n8153), .IN2(n8154), .QN(n8127) );
  NAND2X0 U7942 ( .IN1(n8149), .IN2(n8155), .QN(n8154) );
  NAND2X0 U7943 ( .IN1(n8151), .IN2(n8156), .QN(n8153) );
  NAND2X0 U7944 ( .IN1(n8157), .IN2(n8158), .QN(n8116) );
  NAND3X0 U7945 ( .IN1(n8142), .IN2(n8143), .IN3(n8159), .QN(n8158) );
  NAND2X0 U7946 ( .IN1(n8145), .IN2(n8160), .QN(n8157) );
  INVX0 U7947 ( .INP(n8161), .ZN(n8145) );
  XNOR3X1 U7948 ( .IN1(n8132), .IN2(n8092), .IN3(n8162), .Q(n8137) );
  XOR2X1 U7949 ( .IN1(n8122), .IN2(n8107), .Q(n8162) );
  AND4X1 U7950 ( .IN1(n8142), .IN2(n8163), .IN3(n8164), .IN4(n8165), .Q(n8107)
         );
  OR2X1 U7951 ( .IN1(n8166), .IN2(n8167), .Q(n8165) );
  NAND2X0 U7952 ( .IN1(n8168), .IN2(n8166), .QN(n8164) );
  NAND3X0 U7953 ( .IN1(n8169), .IN2(n8170), .IN3(n8171), .QN(n8122) );
  NAND2X0 U7954 ( .IN1(n8172), .IN2(n8173), .QN(n8170) );
  NAND2X0 U7955 ( .IN1(n8174), .IN2(n8175), .QN(n8169) );
  NAND2X0 U7956 ( .IN1(n8176), .IN2(n8177), .QN(n8092) );
  NAND2X0 U7957 ( .IN1(n8149), .IN2(n8178), .QN(n8177) );
  NOR2X0 U7958 ( .IN1(n8179), .IN2(n8168), .QN(n8149) );
  NAND2X0 U7959 ( .IN1(n8151), .IN2(n8180), .QN(n8176) );
  NOR2X0 U7960 ( .IN1(n8179), .IN2(n8181), .QN(n8151) );
  AND3X1 U7961 ( .IN1(n8182), .IN2(n8183), .IN3(n8171), .Q(n8132) );
  NAND2X0 U7962 ( .IN1(n8184), .IN2(n8173), .QN(n8183) );
  NAND2X0 U7963 ( .IN1(n8174), .IN2(n8185), .QN(n8182) );
  NAND4X0 U7964 ( .IN1(n8091), .IN2(n8094), .IN3(n8186), .IN4(n8187), .QN(
        n8134) );
  OR2X1 U7965 ( .IN1(n7882), .IN2(test_so69), .Q(n8187) );
  NAND2X0 U7966 ( .IN1(n13229), .IN2(n7882), .QN(n8186) );
  AND2X1 U7967 ( .IN1(n2313), .IN2(n8123), .Q(n8094) );
  INVX0 U7968 ( .INP(n8093), .ZN(n8123) );
  NAND2X0 U7969 ( .IN1(n8188), .IN2(g1937), .QN(n8133) );
  XOR2X1 U7970 ( .IN1(n8074), .IN2(n8119), .Q(n8188) );
  NAND3X0 U7971 ( .IN1(n8189), .IN2(n8190), .IN3(n8171), .QN(n8119) );
  NAND2X0 U7972 ( .IN1(n8161), .IN2(n8191), .QN(n8171) );
  NAND2X0 U7973 ( .IN1(n8142), .IN2(n8192), .QN(n8191) );
  NAND2X0 U7974 ( .IN1(n8193), .IN2(n8142), .QN(n8161) );
  NAND2X0 U7975 ( .IN1(n8194), .IN2(n8173), .QN(n8190) );
  NAND2X0 U7976 ( .IN1(n8174), .IN2(n8195), .QN(n8189) );
  INVX0 U7977 ( .INP(n8143), .ZN(n8174) );
  NAND2X0 U7978 ( .IN1(n8193), .IN2(n8192), .QN(n8143) );
  NAND4X0 U7979 ( .IN1(n8142), .IN2(n8163), .IN3(n8196), .IN4(n8197), .QN(
        n8074) );
  NAND2X0 U7980 ( .IN1(n8198), .IN2(n8181), .QN(n8197) );
  NAND2X0 U7981 ( .IN1(n8168), .IN2(n8199), .QN(n8196) );
  NOR2X0 U7982 ( .IN1(n8181), .IN2(n8200), .QN(n8168) );
  NAND2X0 U7983 ( .IN1(n8200), .IN2(n8181), .QN(n8163) );
  INVX0 U7984 ( .INP(n8192), .ZN(n8200) );
  INVX0 U7985 ( .INP(n8179), .ZN(n8142) );
  NAND2X0 U7986 ( .IN1(n2313), .IN2(g1880), .QN(n8179) );
  NAND2X0 U7987 ( .IN1(n8201), .IN2(n8202), .QN(n4240) );
  NAND2X0 U7988 ( .IN1(n2217), .IN2(n8203), .QN(n8202) );
  NAND3X0 U7989 ( .IN1(n8204), .IN2(n8205), .IN3(n8206), .QN(n8201) );
  NAND2X0 U7990 ( .IN1(n8207), .IN2(n8208), .QN(n8205) );
  NAND2X0 U7991 ( .IN1(n6414), .IN2(n8209), .QN(n8204) );
  NAND3X0 U7992 ( .IN1(n8210), .IN2(n8211), .IN3(n2231), .QN(n4239) );
  NAND3X0 U7993 ( .IN1(n8212), .IN2(n8213), .IN3(n8206), .QN(n8210) );
  NAND2X0 U7994 ( .IN1(n8214), .IN2(n8208), .QN(n8213) );
  NAND2X0 U7995 ( .IN1(n8209), .IN2(DFF_795_n1), .QN(n8212) );
  NAND2X0 U7996 ( .IN1(n8211), .IN2(n8215), .QN(n4238) );
  NAND3X0 U7997 ( .IN1(n8216), .IN2(n8217), .IN3(n8206), .QN(n8215) );
  NAND2X0 U7998 ( .IN1(n8218), .IN2(n8208), .QN(n8217) );
  NAND2X0 U7999 ( .IN1(n8209), .IN2(DFF_799_n1), .QN(n8216) );
  NAND3X0 U8000 ( .IN1(n8219), .IN2(n8211), .IN3(n2231), .QN(n4237) );
  NAND3X0 U8001 ( .IN1(n8220), .IN2(n8221), .IN3(n8206), .QN(n8219) );
  NAND2X0 U8002 ( .IN1(n8222), .IN2(n8208), .QN(n8221) );
  NAND2X0 U8003 ( .IN1(n8209), .IN2(DFF_796_n1), .QN(n8220) );
  NAND2X0 U8004 ( .IN1(n8223), .IN2(n8224), .QN(n4236) );
  NAND3X0 U8005 ( .IN1(n8225), .IN2(n8226), .IN3(n8206), .QN(n8224) );
  NAND2X0 U8006 ( .IN1(n8227), .IN2(n8208), .QN(n8226) );
  NAND2X0 U8007 ( .IN1(n8209), .IN2(DFF_794_n1), .QN(n8225) );
  NAND2X0 U8008 ( .IN1(n8228), .IN2(n8229), .QN(n4235) );
  NAND2X0 U8009 ( .IN1(n2217), .IN2(n8230), .QN(n8229) );
  NAND3X0 U8010 ( .IN1(n8231), .IN2(n8232), .IN3(n8206), .QN(n8228) );
  NAND2X0 U8011 ( .IN1(n8233), .IN2(n8208), .QN(n8232) );
  NAND2X0 U8012 ( .IN1(n6415), .IN2(n8209), .QN(n8231) );
  NAND2X0 U8013 ( .IN1(n8223), .IN2(n8234), .QN(n4234) );
  NAND3X0 U8014 ( .IN1(n8235), .IN2(n8236), .IN3(n8206), .QN(n8234) );
  NAND2X0 U8015 ( .IN1(n8237), .IN2(n8208), .QN(n8236) );
  NAND2X0 U8016 ( .IN1(n8209), .IN2(DFF_797_n1), .QN(n8235) );
  AND2X1 U8017 ( .IN1(n8211), .IN2(n8238), .Q(n8223) );
  NAND2X0 U8018 ( .IN1(n2217), .IN2(n2230), .QN(n8238) );
  NAND2X0 U8019 ( .IN1(n8211), .IN2(n8239), .QN(n4233) );
  NAND3X0 U8020 ( .IN1(n8240), .IN2(n8241), .IN3(n8206), .QN(n8239) );
  NAND2X0 U8021 ( .IN1(n8242), .IN2(n8208), .QN(n8241) );
  NAND2X0 U8022 ( .IN1(n8209), .IN2(DFF_798_n1), .QN(n8240) );
  NAND2X0 U8023 ( .IN1(n2217), .IN2(n8243), .QN(n8211) );
  NAND3X0 U8024 ( .IN1(n8244), .IN2(n8245), .IN3(n8246), .QN(n4232) );
  NAND2X0 U8025 ( .IN1(n8247), .IN2(g1196), .QN(n8246) );
  XOR2X1 U8026 ( .IN1(n8248), .IN2(n8249), .Q(n8247) );
  XOR3X1 U8027 ( .IN1(n8227), .IN2(n8237), .IN3(n8250), .Q(n8249) );
  XOR2X1 U8028 ( .IN1(n8214), .IN2(n8222), .Q(n8250) );
  NAND2X0 U8029 ( .IN1(n8251), .IN2(n8252), .QN(n8222) );
  NAND3X0 U8030 ( .IN1(n8253), .IN2(n8254), .IN3(n8255), .QN(n8252) );
  NAND2X0 U8031 ( .IN1(n8256), .IN2(n8257), .QN(n8251) );
  NAND2X0 U8032 ( .IN1(n8258), .IN2(n8259), .QN(n8214) );
  NAND2X0 U8033 ( .IN1(n8260), .IN2(n8261), .QN(n8259) );
  NAND2X0 U8034 ( .IN1(n8262), .IN2(n8263), .QN(n8258) );
  INVX0 U8035 ( .INP(n8261), .ZN(n8263) );
  NAND2X0 U8036 ( .IN1(n8264), .IN2(n8265), .QN(n8237) );
  NAND2X0 U8037 ( .IN1(n8260), .IN2(n8266), .QN(n8265) );
  NAND2X0 U8038 ( .IN1(n8262), .IN2(n8267), .QN(n8264) );
  NAND2X0 U8039 ( .IN1(n8268), .IN2(n8269), .QN(n8227) );
  NAND3X0 U8040 ( .IN1(n8253), .IN2(n8254), .IN3(n8270), .QN(n8269) );
  NAND2X0 U8041 ( .IN1(n8256), .IN2(n8271), .QN(n8268) );
  INVX0 U8042 ( .INP(n8272), .ZN(n8256) );
  XNOR3X1 U8043 ( .IN1(n8242), .IN2(n8207), .IN3(n8273), .Q(n8248) );
  XNOR2X1 U8044 ( .IN1(n8233), .IN2(n8218), .Q(n8273) );
  AND4X1 U8045 ( .IN1(n8253), .IN2(n8274), .IN3(n8275), .IN4(n8276), .Q(n8218)
         );
  NAND2X0 U8046 ( .IN1(n8277), .IN2(n8278), .QN(n8276) );
  NAND2X0 U8047 ( .IN1(n8279), .IN2(n8280), .QN(n8275) );
  AND3X1 U8048 ( .IN1(n8281), .IN2(n8282), .IN3(n8283), .Q(n8233) );
  NAND2X0 U8049 ( .IN1(n8284), .IN2(n8285), .QN(n8282) );
  NAND2X0 U8050 ( .IN1(n8286), .IN2(n8287), .QN(n8281) );
  NAND2X0 U8051 ( .IN1(n8288), .IN2(n8289), .QN(n8207) );
  NAND2X0 U8052 ( .IN1(n8260), .IN2(n8290), .QN(n8289) );
  NOR2X0 U8053 ( .IN1(n8291), .IN2(n8279), .QN(n8260) );
  NAND2X0 U8054 ( .IN1(n8262), .IN2(n8292), .QN(n8288) );
  NOR2X0 U8055 ( .IN1(n8291), .IN2(n8278), .QN(n8262) );
  INVX0 U8056 ( .INP(n8253), .ZN(n8291) );
  AND3X1 U8057 ( .IN1(n8293), .IN2(n8294), .IN3(n8283), .Q(n8242) );
  NAND2X0 U8058 ( .IN1(n8295), .IN2(n8285), .QN(n8294) );
  NAND2X0 U8059 ( .IN1(n8286), .IN2(n8296), .QN(n8293) );
  NAND4X0 U8060 ( .IN1(n8206), .IN2(n8209), .IN3(n8297), .IN4(n8298), .QN(
        n8245) );
  NAND2X0 U8061 ( .IN1(n4489), .IN2(g3229), .QN(n8298) );
  NAND2X0 U8062 ( .IN1(n7882), .IN2(n13230), .QN(n8297) );
  NOR2X0 U8063 ( .IN1(n8243), .IN2(n8208), .QN(n8209) );
  NAND2X0 U8064 ( .IN1(n8299), .IN2(g1243), .QN(n8244) );
  XOR2X1 U8065 ( .IN1(n8203), .IN2(n8230), .Q(n8299) );
  NAND3X0 U8066 ( .IN1(n8300), .IN2(n8301), .IN3(n8283), .QN(n8230) );
  NAND2X0 U8067 ( .IN1(n8272), .IN2(n8302), .QN(n8283) );
  NAND2X0 U8068 ( .IN1(n8253), .IN2(n8303), .QN(n8302) );
  NAND2X0 U8069 ( .IN1(n8304), .IN2(n8253), .QN(n8272) );
  NAND2X0 U8070 ( .IN1(n8305), .IN2(n8285), .QN(n8301) );
  NAND2X0 U8071 ( .IN1(n8286), .IN2(n8306), .QN(n8300) );
  INVX0 U8072 ( .INP(n8254), .ZN(n8286) );
  NAND2X0 U8073 ( .IN1(n8304), .IN2(n8303), .QN(n8254) );
  NAND4X0 U8074 ( .IN1(n8253), .IN2(n8274), .IN3(n8307), .IN4(n8308), .QN(
        n8203) );
  NAND2X0 U8075 ( .IN1(n8309), .IN2(n8278), .QN(n8308) );
  NAND2X0 U8076 ( .IN1(n8279), .IN2(n8310), .QN(n8307) );
  NOR2X0 U8077 ( .IN1(n8278), .IN2(n8311), .QN(n8279) );
  NAND2X0 U8078 ( .IN1(n8311), .IN2(n8278), .QN(n8274) );
  INVX0 U8079 ( .INP(n8303), .ZN(n8311) );
  NOR2X0 U8080 ( .IN1(n8243), .IN2(n4548), .QN(n8253) );
  OR3X1 U8081 ( .IN1(g1249), .IN2(n7265), .IN3(g1245), .Q(n8243) );
  NAND2X0 U8082 ( .IN1(n3896), .IN2(g88), .QN(n4528) );
  NAND2X0 U8083 ( .IN1(n3890), .IN2(g1462), .QN(n4527) );
  NAND2X0 U8084 ( .IN1(n3887), .IN2(test_so78), .QN(n4526) );
  NAND2X0 U8085 ( .IN1(n3692), .IN2(test_so15), .QN(n4521) );
  OR2X1 U8086 ( .IN1(n8312), .IN2(n6434), .Q(n4523) );
  OR2X1 U8087 ( .IN1(n8313), .IN2(n6433), .Q(n4522) );
  NAND2X0 U8088 ( .IN1(n8314), .IN2(n8315), .QN(n3254) );
  NAND2X0 U8089 ( .IN1(n8316), .IN2(n8317), .QN(n8314) );
  INVX0 U8090 ( .INP(n8318), .ZN(n8316) );
  NAND4X0 U8091 ( .IN1(n8319), .IN2(n8320), .IN3(n8321), .IN4(g309), .QN(n3023) );
  NAND4X0 U8092 ( .IN1(n8322), .IN2(n8323), .IN3(n8324), .IN4(g996), .QN(n3016) );
  NAND4X0 U8093 ( .IN1(n8325), .IN2(n8326), .IN3(n8327), .IN4(g1690), .QN(
        n3008) );
  NAND4X0 U8094 ( .IN1(n8328), .IN2(n8329), .IN3(n8330), .IN4(test_so79), .QN(
        n3000) );
  XOR2X1 U8095 ( .IN1(n8331), .IN2(n8332), .Q(n2800) );
  NAND2X0 U8096 ( .IN1(n8333), .IN2(n8334), .QN(n8331) );
  NAND2X0 U8097 ( .IN1(n8332), .IN2(n8335), .QN(n8334) );
  NAND3X0 U8098 ( .IN1(n8336), .IN2(n8337), .IN3(n8338), .QN(n8335) );
  NAND2X0 U8099 ( .IN1(n8339), .IN2(n8340), .QN(n8337) );
  NAND3X0 U8100 ( .IN1(n8341), .IN2(g996), .IN3(n8342), .QN(n8336) );
  NAND3X0 U8101 ( .IN1(n8343), .IN2(n8338), .IN3(n8344), .QN(n8333) );
  XOR2X1 U8102 ( .IN1(n8345), .IN2(n8346), .Q(n2719) );
  XOR2X1 U8103 ( .IN1(n8347), .IN2(n8348), .Q(n2686) );
  XOR2X1 U8104 ( .IN1(n8349), .IN2(n7770), .Q(n2671) );
  INVX0 U8105 ( .INP(n8350), .ZN(n2670) );
  INVX0 U8106 ( .INP(n8351), .ZN(n266) );
  INVX0 U8107 ( .INP(n8352), .ZN(n265) );
  INVX0 U8108 ( .INP(n8353), .ZN(n264) );
  XOR2X1 U8109 ( .IN1(n8340), .IN2(n8354), .Q(n2616) );
  NAND2X0 U8110 ( .IN1(n8355), .IN2(n8356), .QN(n8354) );
  NAND2X0 U8111 ( .IN1(n8357), .IN2(n8358), .QN(n8356) );
  NAND4X0 U8112 ( .IN1(n8359), .IN2(n8360), .IN3(n8361), .IN4(n8338), .QN(
        n8355) );
  NAND3X0 U8113 ( .IN1(n8332), .IN2(n8362), .IN3(n8343), .QN(n8361) );
  AND3X1 U8114 ( .IN1(n8363), .IN2(n8340), .IN3(n3102), .Q(n8343) );
  OR2X1 U8115 ( .IN1(n8364), .IN2(n8342), .Q(n8360) );
  NAND2X0 U8116 ( .IN1(n8365), .IN2(n8342), .QN(n8359) );
  NAND2X0 U8117 ( .IN1(n8366), .IN2(n8367), .QN(n8365) );
  NAND2X0 U8118 ( .IN1(n8332), .IN2(n8368), .QN(n8367) );
  NAND3X0 U8119 ( .IN1(n8369), .IN2(n8362), .IN3(n8370), .QN(n8368) );
  INVX0 U8120 ( .INP(n8339), .ZN(n8370) );
  NAND2X0 U8121 ( .IN1(n8371), .IN2(n8372), .QN(n8339) );
  NAND2X0 U8122 ( .IN1(n8373), .IN2(n3102), .QN(n8372) );
  INVX0 U8123 ( .INP(n8363), .ZN(n8373) );
  NAND2X0 U8124 ( .IN1(n8364), .IN2(n8374), .QN(n8369) );
  NAND2X0 U8125 ( .IN1(n8375), .IN2(n8344), .QN(n8366) );
  NAND2X0 U8126 ( .IN1(n2632), .IN2(n8371), .QN(n8375) );
  INVX0 U8127 ( .INP(n8376), .ZN(n257) );
  NOR4X0 U8128 ( .IN1(g559), .IN2(g21851), .IN3(g563), .IN4(n8377), .QN(n2478)
         );
  NOR2X0 U8129 ( .IN1(n4298), .IN2(g499), .QN(n8377) );
  NOR2X0 U8130 ( .IN1(n7802), .IN2(n7786), .QN(n2446) );
  AND2X1 U8131 ( .IN1(n4360), .IN2(n8378), .Q(n7786) );
  NAND2X0 U8132 ( .IN1(n7005), .IN2(n7271), .QN(n8378) );
  NAND2X0 U8133 ( .IN1(n7271), .IN2(n8379), .QN(n7802) );
  NAND2X0 U8134 ( .IN1(n4360), .IN2(n7005), .QN(n8379) );
  NAND2X0 U8135 ( .IN1(g499), .IN2(n8380), .QN(n2445) );
  NAND4X0 U8136 ( .IN1(n8381), .IN2(n8382), .IN3(n8383), .IN4(n8384), .QN(
        n8380) );
  NAND2X0 U8137 ( .IN1(n6778), .IN2(g629), .QN(n8383) );
  NAND2X0 U8138 ( .IN1(n6774), .IN2(g6677), .QN(n8382) );
  NAND2X0 U8139 ( .IN1(n6773), .IN2(g6911), .QN(n8381) );
  NAND2X0 U8140 ( .IN1(n7887), .IN2(n7851), .QN(n2430) );
  INVX0 U8141 ( .INP(n8384), .ZN(n7887) );
  NAND4X0 U8142 ( .IN1(n8385), .IN2(n8386), .IN3(n8387), .IN4(n8388), .QN(
        n8384) );
  NOR4X0 U8143 ( .IN1(n8389), .IN2(n7867), .IN3(n7875), .IN4(n7846), .QN(n8388) );
  NAND3X0 U8144 ( .IN1(n7870), .IN2(n8390), .IN3(n7878), .QN(n8389) );
  NAND3X0 U8145 ( .IN1(n8391), .IN2(n8392), .IN3(n8393), .QN(n8390) );
  NAND2X0 U8146 ( .IN1(n7229), .IN2(g6911), .QN(n8393) );
  NAND2X0 U8147 ( .IN1(n7232), .IN2(g629), .QN(n8392) );
  NAND2X0 U8148 ( .IN1(n7165), .IN2(g6677), .QN(n8391) );
  NOR3X0 U8149 ( .IN1(n7850), .IN2(n7857), .IN3(n7861), .QN(n8387) );
  NOR2X0 U8150 ( .IN1(n7888), .IN2(n7892), .QN(n8385) );
  INVX0 U8151 ( .INP(n7893), .ZN(n7892) );
  NAND2X0 U8152 ( .IN1(g2574), .IN2(n8394), .QN(n2374) );
  NAND4X0 U8153 ( .IN1(n8395), .IN2(n8396), .IN3(n8397), .IN4(n8398), .QN(
        n8394) );
  NAND2X0 U8154 ( .IN1(n6775), .IN2(g2703), .QN(n8397) );
  NAND2X0 U8155 ( .IN1(n6768), .IN2(g7425), .QN(n8396) );
  NAND2X0 U8156 ( .IN1(n6767), .IN2(g7487), .QN(n8395) );
  NOR2X0 U8157 ( .IN1(n7901), .IN2(n7899), .QN(n2361) );
  AND2X1 U8158 ( .IN1(n4352), .IN2(n8399), .Q(n7899) );
  NAND2X0 U8159 ( .IN1(n7002), .IN2(n4303), .QN(n8399) );
  NAND2X0 U8160 ( .IN1(n4303), .IN2(n8400), .QN(n7901) );
  NAND2X0 U8161 ( .IN1(n4352), .IN2(n7002), .QN(n8400) );
  NAND2X0 U8162 ( .IN1(n8023), .IN2(n7981), .QN(n2351) );
  INVX0 U8163 ( .INP(n8398), .ZN(n8023) );
  NAND4X0 U8164 ( .IN1(n8401), .IN2(n8402), .IN3(n8403), .IN4(n8404), .QN(
        n8398) );
  NOR4X0 U8165 ( .IN1(n8405), .IN2(n8063), .IN3(n8035), .IN4(n8041), .QN(n8404) );
  NAND3X0 U8166 ( .IN1(n8071), .IN2(n8406), .IN3(n8012), .QN(n8405) );
  NAND3X0 U8167 ( .IN1(n8407), .IN2(n8408), .IN3(n8409), .QN(n8406) );
  NAND2X0 U8168 ( .IN1(n7226), .IN2(g7487), .QN(n8409) );
  OR2X1 U8169 ( .IN1(n4292), .IN2(test_so95), .Q(n8408) );
  NAND2X0 U8170 ( .IN1(n7162), .IN2(g7425), .QN(n8407) );
  NOR3X0 U8171 ( .IN1(n8051), .IN2(n7993), .IN3(n8016), .QN(n8403) );
  NOR2X0 U8172 ( .IN1(n8030), .IN2(n7977), .QN(n8401) );
  INVX0 U8173 ( .INP(n7989), .ZN(n7977) );
  NOR3X0 U8174 ( .IN1(g1943), .IN2(n7264), .IN3(g1939), .QN(n2313) );
  NAND2X0 U8175 ( .IN1(g1880), .IN2(n8410), .QN(n2302) );
  NAND4X0 U8176 ( .IN1(n8411), .IN2(n8412), .IN3(n8413), .IN4(n8192), .QN(
        n8410) );
  NAND4X0 U8177 ( .IN1(n8414), .IN2(n8415), .IN3(n8416), .IN4(n8417), .QN(
        n8192) );
  NOR4X0 U8178 ( .IN1(n8418), .IN2(n8150), .IN3(n8155), .IN4(n8159), .QN(n8417) );
  NAND3X0 U8179 ( .IN1(n8146), .IN2(n8419), .IN3(n8180), .QN(n8418) );
  NAND3X0 U8180 ( .IN1(n8420), .IN2(n8421), .IN3(n8422), .QN(n8419) );
  NAND2X0 U8181 ( .IN1(n7227), .IN2(g7357), .QN(n8422) );
  NAND2X0 U8182 ( .IN1(n7230), .IN2(g2009), .QN(n8421) );
  NAND2X0 U8183 ( .IN1(n7163), .IN2(g7229), .QN(n8420) );
  AND3X1 U8184 ( .IN1(n8175), .IN2(n8199), .IN3(n8166), .Q(n8416) );
  NOR2X0 U8185 ( .IN1(n8184), .IN2(n8194), .QN(n8414) );
  INVX0 U8186 ( .INP(n8195), .ZN(n8194) );
  NAND2X0 U8187 ( .IN1(n6776), .IN2(g2009), .QN(n8413) );
  NAND2X0 U8188 ( .IN1(n6770), .IN2(g7229), .QN(n8412) );
  NAND2X0 U8189 ( .IN1(n6769), .IN2(g7357), .QN(n8411) );
  NOR2X0 U8190 ( .IN1(n8093), .IN2(n8091), .QN(n2289) );
  AND2X1 U8191 ( .IN1(n4311), .IN2(n8423), .Q(n8091) );
  NAND2X0 U8192 ( .IN1(n7003), .IN2(n4297), .QN(n8423) );
  NAND2X0 U8193 ( .IN1(n4297), .IN2(n8424), .QN(n8093) );
  NAND2X0 U8194 ( .IN1(n4311), .IN2(n7003), .QN(n8424) );
  NAND2X0 U8195 ( .IN1(g1186), .IN2(n8425), .QN(n2230) );
  NAND4X0 U8196 ( .IN1(n8426), .IN2(n8427), .IN3(n8428), .IN4(n8303), .QN(
        n8425) );
  NAND4X0 U8197 ( .IN1(n8429), .IN2(n8430), .IN3(n8431), .IN4(n8432), .QN(
        n8303) );
  NOR4X0 U8198 ( .IN1(n8433), .IN2(n8261), .IN3(n8266), .IN4(n8270), .QN(n8432) );
  NAND3X0 U8199 ( .IN1(n8257), .IN2(n8434), .IN3(n8292), .QN(n8433) );
  INVX0 U8200 ( .INP(n8290), .ZN(n8292) );
  NAND3X0 U8201 ( .IN1(n8435), .IN2(n8436), .IN3(n8437), .QN(n8434) );
  NAND2X0 U8202 ( .IN1(n7228), .IN2(g7161), .QN(n8437) );
  NAND2X0 U8203 ( .IN1(n7231), .IN2(g1315), .QN(n8436) );
  NAND2X0 U8204 ( .IN1(n7164), .IN2(g6979), .QN(n8435) );
  NOR3X0 U8205 ( .IN1(n8284), .IN2(n8309), .IN3(n8277), .QN(n8431) );
  NOR2X0 U8206 ( .IN1(n8295), .IN2(n8305), .QN(n8429) );
  INVX0 U8207 ( .INP(n8306), .ZN(n8305) );
  NAND2X0 U8208 ( .IN1(n6777), .IN2(g1315), .QN(n8428) );
  NAND2X0 U8209 ( .IN1(n6772), .IN2(g6979), .QN(n8427) );
  NAND2X0 U8210 ( .IN1(n6771), .IN2(g7161), .QN(n8426) );
  NOR2X0 U8211 ( .IN1(n8208), .IN2(n8206), .QN(n2217) );
  AND2X1 U8212 ( .IN1(n4353), .IN2(n8438), .Q(n8206) );
  NAND2X0 U8213 ( .IN1(n7004), .IN2(n4304), .QN(n8438) );
  NAND2X0 U8214 ( .IN1(n4304), .IN2(n8439), .QN(n8208) );
  NAND2X0 U8215 ( .IN1(n4353), .IN2(n7004), .QN(n8439) );
  INVX0 U8216 ( .INP(g27380), .ZN(n19) );
  INVX0 U8217 ( .INP(g24734), .ZN(n144) );
  INVX0 U8218 ( .INP(g25435), .ZN(n138) );
  INVX0 U8219 ( .INP(g26135), .ZN(n129) );
  NAND2X0 U8220 ( .IN1(n8440), .IN2(n8441), .QN(g30801) );
  NAND2X0 U8221 ( .IN1(n4494), .IN2(g3108), .QN(n8441) );
  NAND2X0 U8222 ( .IN1(g30072), .IN2(g3109), .QN(n8440) );
  NAND2X0 U8223 ( .IN1(n8442), .IN2(n8443), .QN(g30798) );
  NAND2X0 U8224 ( .IN1(n4383), .IN2(g3107), .QN(n8443) );
  NAND2X0 U8225 ( .IN1(g30072), .IN2(g8030), .QN(n8442) );
  NAND2X0 U8226 ( .IN1(n8444), .IN2(n8445), .QN(g30796) );
  OR2X1 U8227 ( .IN1(g8106), .IN2(n4438), .Q(n8445) );
  NAND2X0 U8228 ( .IN1(g30072), .IN2(g8106), .QN(n8444) );
  NAND2X0 U8229 ( .IN1(n8446), .IN2(n8447), .QN(g30709) );
  NAND2X0 U8230 ( .IN1(n8448), .IN2(g7264), .QN(n8447) );
  OR2X1 U8231 ( .IN1(n8449), .IN2(n6532), .Q(n8446) );
  NAND2X0 U8232 ( .IN1(n8450), .IN2(n8451), .QN(g30708) );
  NAND2X0 U8233 ( .IN1(n8452), .IN2(n4618), .QN(n8451) );
  OR2X1 U8234 ( .IN1(n8453), .IN2(n6548), .Q(n8450) );
  NAND2X0 U8235 ( .IN1(n8454), .IN2(n8455), .QN(g30707) );
  NAND2X0 U8236 ( .IN1(n8448), .IN2(g5555), .QN(n8455) );
  OR2X1 U8237 ( .IN1(n8456), .IN2(n6543), .Q(n8454) );
  NAND2X0 U8238 ( .IN1(n8457), .IN2(n8458), .QN(g30706) );
  NAND2X0 U8239 ( .IN1(n8452), .IN2(g7014), .QN(n8458) );
  OR2X1 U8240 ( .IN1(n8459), .IN2(n6535), .Q(n8457) );
  NAND2X0 U8241 ( .IN1(n8460), .IN2(n8461), .QN(g30705) );
  OR2X1 U8242 ( .IN1(g1088), .IN2(n6553), .Q(n8461) );
  NAND2X0 U8243 ( .IN1(n2594), .IN2(g1088), .QN(n8460) );
  NAND2X0 U8244 ( .IN1(n8462), .IN2(n8463), .QN(g30704) );
  NAND2X0 U8245 ( .IN1(n8452), .IN2(g5511), .QN(n8463) );
  AND2X1 U8246 ( .IN1(n8464), .IN2(n8465), .Q(n8452) );
  XOR2X1 U8247 ( .IN1(n8466), .IN2(n8467), .Q(n8464) );
  NAND2X0 U8248 ( .IN1(n8468), .IN2(n8469), .QN(n8467) );
  NAND2X0 U8249 ( .IN1(n8470), .IN2(n8471), .QN(n8469) );
  NAND4X0 U8250 ( .IN1(n8472), .IN2(n8473), .IN3(n8474), .IN4(n8475), .QN(
        n8468) );
  NAND3X0 U8251 ( .IN1(n8476), .IN2(n8477), .IN3(n8478), .QN(n8474) );
  OR2X1 U8252 ( .IN1(n8479), .IN2(n8480), .Q(n8473) );
  NAND2X0 U8253 ( .IN1(n8481), .IN2(n8480), .QN(n8472) );
  NAND2X0 U8254 ( .IN1(n8482), .IN2(n8483), .QN(n8481) );
  NAND2X0 U8255 ( .IN1(n8476), .IN2(n8484), .QN(n8483) );
  NAND3X0 U8256 ( .IN1(n8485), .IN2(n8477), .IN3(n8486), .QN(n8484) );
  INVX0 U8257 ( .INP(n8487), .ZN(n8486) );
  NAND3X0 U8258 ( .IN1(n8488), .IN2(n8479), .IN3(n8489), .QN(n8485) );
  NAND2X0 U8259 ( .IN1(n8490), .IN2(n8491), .QN(n8482) );
  NAND2X0 U8260 ( .IN1(n8492), .IN2(n8493), .QN(n8490) );
  NAND2X0 U8261 ( .IN1(n8489), .IN2(n8488), .QN(n8492) );
  OR2X1 U8262 ( .IN1(n8494), .IN2(n6549), .Q(n8462) );
  NAND2X0 U8263 ( .IN1(n8495), .IN2(n8496), .QN(g30703) );
  OR2X1 U8264 ( .IN1(g6712), .IN2(n6538), .Q(n8496) );
  NAND2X0 U8265 ( .IN1(n2594), .IN2(g6712), .QN(n8495) );
  NAND2X0 U8266 ( .IN1(n8497), .IN2(n8498), .QN(g30702) );
  NAND2X0 U8267 ( .IN1(n8499), .IN2(n4640), .QN(n8498) );
  OR2X1 U8268 ( .IN1(n8500), .IN2(n6560), .Q(n8497) );
  NAND2X0 U8269 ( .IN1(n8501), .IN2(n8502), .QN(g30701) );
  OR2X1 U8270 ( .IN1(g5472), .IN2(n6554), .Q(n8502) );
  NAND2X0 U8271 ( .IN1(n2594), .IN2(g5472), .QN(n8501) );
  NAND2X0 U8272 ( .IN1(n8503), .IN2(n8504), .QN(g30700) );
  NAND2X0 U8273 ( .IN1(n8499), .IN2(g6447), .QN(n8504) );
  NAND2X0 U8274 ( .IN1(test_so18), .IN2(n4499), .QN(n8503) );
  NAND2X0 U8275 ( .IN1(n8505), .IN2(n8506), .QN(g30699) );
  NAND2X0 U8276 ( .IN1(n8499), .IN2(g5437), .QN(n8506) );
  AND2X1 U8277 ( .IN1(n8507), .IN2(n8508), .Q(n8499) );
  XOR2X1 U8278 ( .IN1(n8509), .IN2(n8510), .Q(n8507) );
  NAND2X0 U8279 ( .IN1(n8511), .IN2(n8512), .QN(n8510) );
  NAND2X0 U8280 ( .IN1(n8513), .IN2(n8514), .QN(n8512) );
  NAND4X0 U8281 ( .IN1(n8515), .IN2(n8516), .IN3(n8517), .IN4(n8518), .QN(
        n8511) );
  NAND3X0 U8282 ( .IN1(n8519), .IN2(n8520), .IN3(n8521), .QN(n8517) );
  OR2X1 U8283 ( .IN1(n8522), .IN2(n8523), .Q(n8516) );
  NAND2X0 U8284 ( .IN1(n8524), .IN2(n8523), .QN(n8515) );
  NAND2X0 U8285 ( .IN1(n8525), .IN2(n8526), .QN(n8524) );
  NAND2X0 U8286 ( .IN1(n8519), .IN2(n8527), .QN(n8526) );
  NAND3X0 U8287 ( .IN1(n8528), .IN2(n8520), .IN3(n8529), .QN(n8527) );
  INVX0 U8288 ( .INP(n8530), .ZN(n8529) );
  NAND3X0 U8289 ( .IN1(n8531), .IN2(n8522), .IN3(n8532), .QN(n8528) );
  NAND2X0 U8290 ( .IN1(n8533), .IN2(n8534), .QN(n8525) );
  NAND2X0 U8291 ( .IN1(n8535), .IN2(n8536), .QN(n8533) );
  NAND2X0 U8292 ( .IN1(n8532), .IN2(n8531), .QN(n8535) );
  OR2X1 U8293 ( .IN1(n8537), .IN2(n6561), .Q(n8505) );
  NAND2X0 U8294 ( .IN1(n8538), .IN2(n8539), .QN(g30695) );
  NAND2X0 U8295 ( .IN1(n4367), .IN2(g2276), .QN(n8539) );
  NAND2X0 U8296 ( .IN1(n8540), .IN2(g2241), .QN(n8538) );
  NAND2X0 U8297 ( .IN1(n8541), .IN2(n8542), .QN(g30694) );
  NAND2X0 U8298 ( .IN1(n4367), .IN2(g2348), .QN(n8542) );
  NAND2X0 U8299 ( .IN1(n8543), .IN2(g2241), .QN(n8541) );
  NAND2X0 U8300 ( .IN1(n8544), .IN2(n8545), .QN(g30693) );
  NAND2X0 U8301 ( .IN1(g2273), .IN2(n7266), .QN(n8545) );
  NAND2X0 U8302 ( .IN1(test_so73), .IN2(n8540), .QN(n8544) );
  NAND2X0 U8303 ( .IN1(n8546), .IN2(n8547), .QN(g30692) );
  NAND2X0 U8304 ( .IN1(n4368), .IN2(g1582), .QN(n8547) );
  NAND2X0 U8305 ( .IN1(n8548), .IN2(g1547), .QN(n8546) );
  NAND2X0 U8306 ( .IN1(n8549), .IN2(n8550), .QN(g30691) );
  NAND2X0 U8307 ( .IN1(g2345), .IN2(n7266), .QN(n8550) );
  NAND2X0 U8308 ( .IN1(n8543), .IN2(test_so73), .QN(n8549) );
  NAND2X0 U8309 ( .IN1(n8551), .IN2(n8552), .QN(g30690) );
  NAND2X0 U8310 ( .IN1(n4324), .IN2(g2270), .QN(n8552) );
  NAND2X0 U8311 ( .IN1(n8540), .IN2(g6837), .QN(n8551) );
  NAND3X0 U8312 ( .IN1(n8553), .IN2(n8554), .IN3(n8555), .QN(n8540) );
  NAND2X0 U8313 ( .IN1(n8556), .IN2(n8557), .QN(n8554) );
  XOR2X1 U8314 ( .IN1(n8558), .IN2(n7769), .Q(n8556) );
  NAND2X0 U8315 ( .IN1(n8559), .IN2(g2175), .QN(n8553) );
  NAND2X0 U8316 ( .IN1(n8560), .IN2(n8561), .QN(g30689) );
  NAND2X0 U8317 ( .IN1(n4368), .IN2(g1654), .QN(n8561) );
  NAND2X0 U8318 ( .IN1(n8562), .IN2(g1547), .QN(n8560) );
  NAND2X0 U8319 ( .IN1(n8563), .IN2(n8564), .QN(g30688) );
  NAND2X0 U8320 ( .IN1(n4515), .IN2(g1579), .QN(n8564) );
  NAND2X0 U8321 ( .IN1(n8548), .IN2(g6782), .QN(n8563) );
  NAND2X0 U8322 ( .IN1(n8565), .IN2(n8566), .QN(g30687) );
  NAND2X0 U8323 ( .IN1(g888), .IN2(n7267), .QN(n8566) );
  NAND2X0 U8324 ( .IN1(test_so31), .IN2(n8567), .QN(n8565) );
  NAND2X0 U8325 ( .IN1(n8568), .IN2(n8569), .QN(g30686) );
  NAND2X0 U8326 ( .IN1(n4324), .IN2(g2342), .QN(n8569) );
  NAND2X0 U8327 ( .IN1(n8543), .IN2(g6837), .QN(n8568) );
  AND3X1 U8328 ( .IN1(n8570), .IN2(n8571), .IN3(n8572), .Q(n8543) );
  NAND2X0 U8329 ( .IN1(n8559), .IN2(n8573), .QN(n8572) );
  NAND2X0 U8330 ( .IN1(n8574), .IN2(n8557), .QN(n8570) );
  XNOR2X1 U8331 ( .IN1(n7759), .IN2(n2669), .Q(n8574) );
  NAND2X0 U8332 ( .IN1(n8575), .IN2(n8576), .QN(g30684) );
  NAND2X0 U8333 ( .IN1(n4515), .IN2(g1651), .QN(n8576) );
  NAND2X0 U8334 ( .IN1(n8562), .IN2(g6782), .QN(n8575) );
  NAND2X0 U8335 ( .IN1(n8577), .IN2(n8578), .QN(g30683) );
  NAND2X0 U8336 ( .IN1(n4317), .IN2(g1576), .QN(n8578) );
  NAND2X0 U8337 ( .IN1(n8548), .IN2(g6573), .QN(n8577) );
  NAND3X0 U8338 ( .IN1(n8579), .IN2(n8580), .IN3(n8581), .QN(n8548) );
  NAND2X0 U8339 ( .IN1(n8582), .IN2(n8583), .QN(n8580) );
  XOR2X1 U8340 ( .IN1(n8584), .IN2(n8585), .Q(n8582) );
  NAND2X0 U8341 ( .IN1(n8586), .IN2(g1481), .QN(n8579) );
  NAND2X0 U8342 ( .IN1(n8587), .IN2(n8588), .QN(g30682) );
  NAND2X0 U8343 ( .IN1(g960), .IN2(n7267), .QN(n8588) );
  NAND2X0 U8344 ( .IN1(n8589), .IN2(test_so31), .QN(n8587) );
  NAND2X0 U8345 ( .IN1(n8590), .IN2(n8591), .QN(g30681) );
  NAND2X0 U8346 ( .IN1(n4312), .IN2(g885), .QN(n8591) );
  NAND2X0 U8347 ( .IN1(n8567), .IN2(g6518), .QN(n8590) );
  NAND2X0 U8348 ( .IN1(n8592), .IN2(n8593), .QN(g30680) );
  NAND2X0 U8349 ( .IN1(n4369), .IN2(g201), .QN(n8593) );
  NAND2X0 U8350 ( .IN1(n8594), .IN2(g165), .QN(n8592) );
  NAND2X0 U8351 ( .IN1(n8595), .IN2(n8596), .QN(g30679) );
  NAND2X0 U8352 ( .IN1(n4367), .IN2(g2321), .QN(n8596) );
  NAND2X0 U8353 ( .IN1(n8597), .IN2(g2241), .QN(n8595) );
  NAND2X0 U8354 ( .IN1(n8598), .IN2(n8599), .QN(g30678) );
  NAND2X0 U8355 ( .IN1(n4317), .IN2(g1648), .QN(n8599) );
  NAND2X0 U8356 ( .IN1(n8562), .IN2(g6573), .QN(n8598) );
  AND3X1 U8357 ( .IN1(n8600), .IN2(n8601), .IN3(n8602), .Q(n8562) );
  NAND2X0 U8358 ( .IN1(n8586), .IN2(n8603), .QN(n8602) );
  NAND2X0 U8359 ( .IN1(n8604), .IN2(n8583), .QN(n8600) );
  XNOR2X1 U8360 ( .IN1(n7735), .IN2(n2684), .Q(n8604) );
  NAND2X0 U8361 ( .IN1(n8605), .IN2(n8606), .QN(g30677) );
  NAND2X0 U8362 ( .IN1(n4312), .IN2(g957), .QN(n8606) );
  NAND2X0 U8363 ( .IN1(n8589), .IN2(g6518), .QN(n8605) );
  NAND2X0 U8364 ( .IN1(n8607), .IN2(n8608), .QN(g30676) );
  NAND2X0 U8365 ( .IN1(n4323), .IN2(g882), .QN(n8608) );
  NAND2X0 U8366 ( .IN1(n8567), .IN2(g6368), .QN(n8607) );
  NAND3X0 U8367 ( .IN1(n8609), .IN2(n8610), .IN3(n8611), .QN(n8567) );
  NAND2X0 U8368 ( .IN1(n8612), .IN2(n8613), .QN(n8610) );
  XNOR2X1 U8369 ( .IN1(n7699), .IN2(n8614), .Q(n8612) );
  NAND2X0 U8370 ( .IN1(n8615), .IN2(g793), .QN(n8609) );
  NAND2X0 U8371 ( .IN1(n8616), .IN2(n8617), .QN(g30675) );
  NAND2X0 U8372 ( .IN1(n4369), .IN2(g273), .QN(n8617) );
  NAND2X0 U8373 ( .IN1(n8618), .IN2(g165), .QN(n8616) );
  NAND2X0 U8374 ( .IN1(n8619), .IN2(n8620), .QN(g30674) );
  NAND2X0 U8375 ( .IN1(n4512), .IN2(g198), .QN(n8620) );
  NAND2X0 U8376 ( .IN1(n8594), .IN2(g6313), .QN(n8619) );
  NAND2X0 U8377 ( .IN1(n8621), .IN2(n8622), .QN(g30673) );
  NAND2X0 U8378 ( .IN1(g2318), .IN2(n7266), .QN(n8622) );
  NAND2X0 U8379 ( .IN1(n8597), .IN2(test_so73), .QN(n8621) );
  NAND2X0 U8380 ( .IN1(n8623), .IN2(n8624), .QN(g30672) );
  NAND2X0 U8381 ( .IN1(n4367), .IN2(g2312), .QN(n8624) );
  NAND2X0 U8382 ( .IN1(n8625), .IN2(g2241), .QN(n8623) );
  NAND2X0 U8383 ( .IN1(n8626), .IN2(n8627), .QN(g30671) );
  NAND2X0 U8384 ( .IN1(n4368), .IN2(g1627), .QN(n8627) );
  NAND2X0 U8385 ( .IN1(n8628), .IN2(g1547), .QN(n8626) );
  NAND2X0 U8386 ( .IN1(n8629), .IN2(n8630), .QN(g30670) );
  NAND2X0 U8387 ( .IN1(n4323), .IN2(g954), .QN(n8630) );
  NAND2X0 U8388 ( .IN1(n8589), .IN2(g6368), .QN(n8629) );
  AND3X1 U8389 ( .IN1(n8631), .IN2(n8632), .IN3(n8633), .Q(n8589) );
  NAND2X0 U8390 ( .IN1(n8615), .IN2(n8634), .QN(n8633) );
  NAND2X0 U8391 ( .IN1(n8613), .IN2(n8635), .QN(n8631) );
  XOR2X1 U8392 ( .IN1(n8636), .IN2(n8637), .Q(n8635) );
  NOR2X0 U8393 ( .IN1(n8638), .IN2(n8639), .QN(n8637) );
  XOR2X1 U8394 ( .IN1(n8640), .IN2(n8641), .Q(n8638) );
  NAND2X0 U8395 ( .IN1(n8642), .IN2(n8643), .QN(g30669) );
  NAND2X0 U8396 ( .IN1(n4512), .IN2(g270), .QN(n8643) );
  NAND2X0 U8397 ( .IN1(n8618), .IN2(g6313), .QN(n8642) );
  NAND2X0 U8398 ( .IN1(n8644), .IN2(n8645), .QN(g30668) );
  NAND2X0 U8399 ( .IN1(n4318), .IN2(g195), .QN(n8645) );
  NAND2X0 U8400 ( .IN1(n8594), .IN2(g6231), .QN(n8644) );
  NAND3X0 U8401 ( .IN1(n8646), .IN2(n8647), .IN3(n8648), .QN(n8594) );
  NAND2X0 U8402 ( .IN1(n8649), .IN2(n8650), .QN(n8647) );
  XOR2X1 U8403 ( .IN1(n8651), .IN2(n8652), .Q(n8649) );
  NAND2X0 U8404 ( .IN1(n8653), .IN2(g105), .QN(n8646) );
  NAND2X0 U8405 ( .IN1(n8654), .IN2(n8655), .QN(g30667) );
  NAND2X0 U8406 ( .IN1(n4324), .IN2(g2315), .QN(n8655) );
  NAND2X0 U8407 ( .IN1(n8597), .IN2(g6837), .QN(n8654) );
  AND3X1 U8408 ( .IN1(n8656), .IN2(n8571), .IN3(n8657), .Q(n8597) );
  NAND2X0 U8409 ( .IN1(n8559), .IN2(n4389), .QN(n8657) );
  NAND2X0 U8410 ( .IN1(n8557), .IN2(n8658), .QN(n8656) );
  XOR2X1 U8411 ( .IN1(n8659), .IN2(n8660), .Q(n8658) );
  AND2X1 U8412 ( .IN1(n8661), .IN2(n8558), .Q(n8660) );
  NAND2X0 U8413 ( .IN1(n8662), .IN2(n8663), .QN(g30666) );
  NAND2X0 U8414 ( .IN1(g2309), .IN2(n7266), .QN(n8663) );
  NAND2X0 U8415 ( .IN1(n8625), .IN2(test_so73), .QN(n8662) );
  NAND2X0 U8416 ( .IN1(n8664), .IN2(n8665), .QN(g30665) );
  NAND2X0 U8417 ( .IN1(n4367), .IN2(g2303), .QN(n8665) );
  NAND2X0 U8418 ( .IN1(n8666), .IN2(g2241), .QN(n8664) );
  NAND2X0 U8419 ( .IN1(n8667), .IN2(n8668), .QN(g30664) );
  NAND2X0 U8420 ( .IN1(n4515), .IN2(g1624), .QN(n8668) );
  NAND2X0 U8421 ( .IN1(n8628), .IN2(g6782), .QN(n8667) );
  NAND2X0 U8422 ( .IN1(n8669), .IN2(n8670), .QN(g30663) );
  NAND2X0 U8423 ( .IN1(n4368), .IN2(g1618), .QN(n8670) );
  NAND2X0 U8424 ( .IN1(n8671), .IN2(g1547), .QN(n8669) );
  NAND2X0 U8425 ( .IN1(n8672), .IN2(n8673), .QN(g30662) );
  NAND2X0 U8426 ( .IN1(g933), .IN2(n7267), .QN(n8673) );
  NAND2X0 U8427 ( .IN1(n8674), .IN2(test_so31), .QN(n8672) );
  NAND2X0 U8428 ( .IN1(n8675), .IN2(n8676), .QN(g30661) );
  NAND2X0 U8429 ( .IN1(n4318), .IN2(g267), .QN(n8676) );
  NAND2X0 U8430 ( .IN1(n8618), .IN2(g6231), .QN(n8675) );
  AND3X1 U8431 ( .IN1(n8677), .IN2(n8678), .IN3(n8679), .Q(n8618) );
  NAND2X0 U8432 ( .IN1(n8653), .IN2(n8680), .QN(n8679) );
  NAND2X0 U8433 ( .IN1(n8681), .IN2(n8650), .QN(n8677) );
  XNOR2X1 U8434 ( .IN1(n7676), .IN2(n2717), .Q(n8681) );
  NAND2X0 U8435 ( .IN1(n8682), .IN2(n8683), .QN(g30660) );
  NAND2X0 U8436 ( .IN1(n4324), .IN2(g2306), .QN(n8683) );
  NAND2X0 U8437 ( .IN1(n8625), .IN2(g6837), .QN(n8682) );
  AND3X1 U8438 ( .IN1(n8684), .IN2(n8571), .IN3(n8685), .Q(n8625) );
  NAND2X0 U8439 ( .IN1(n8559), .IN2(n4373), .QN(n8685) );
  NAND2X0 U8440 ( .IN1(n8686), .IN2(n4529), .QN(n8571) );
  NAND2X0 U8441 ( .IN1(n8557), .IN2(n8687), .QN(n8684) );
  XOR2X1 U8442 ( .IN1(n7774), .IN2(n8688), .Q(n8687) );
  NAND2X0 U8443 ( .IN1(n8689), .IN2(n8690), .QN(g30659) );
  NAND2X0 U8444 ( .IN1(g2300), .IN2(n7266), .QN(n8690) );
  NAND2X0 U8445 ( .IN1(test_so73), .IN2(n8666), .QN(n8689) );
  NAND2X0 U8446 ( .IN1(n8691), .IN2(n8692), .QN(g30658) );
  NAND2X0 U8447 ( .IN1(n8628), .IN2(g6573), .QN(n8692) );
  AND3X1 U8448 ( .IN1(n8693), .IN2(n8601), .IN3(n8694), .Q(n8628) );
  NAND2X0 U8449 ( .IN1(n8586), .IN2(n4390), .QN(n8694) );
  NAND2X0 U8450 ( .IN1(n8583), .IN2(n8695), .QN(n8693) );
  XOR2X1 U8451 ( .IN1(n7733), .IN2(n8696), .Q(n8695) );
  NAND2X0 U8452 ( .IN1(n8585), .IN2(n8697), .QN(n8696) );
  NAND2X0 U8453 ( .IN1(test_so55), .IN2(n4317), .QN(n8691) );
  NAND2X0 U8454 ( .IN1(n8698), .IN2(n8699), .QN(g30657) );
  NAND2X0 U8455 ( .IN1(n4515), .IN2(g1615), .QN(n8699) );
  NAND2X0 U8456 ( .IN1(n8671), .IN2(g6782), .QN(n8698) );
  NAND2X0 U8457 ( .IN1(n8700), .IN2(n8701), .QN(g30656) );
  NAND2X0 U8458 ( .IN1(n4368), .IN2(g1609), .QN(n8701) );
  NAND2X0 U8459 ( .IN1(n8702), .IN2(g1547), .QN(n8700) );
  NAND2X0 U8460 ( .IN1(n8703), .IN2(n8704), .QN(g30655) );
  NAND2X0 U8461 ( .IN1(n4312), .IN2(g930), .QN(n8704) );
  NAND2X0 U8462 ( .IN1(n8674), .IN2(g6518), .QN(n8703) );
  NAND2X0 U8463 ( .IN1(n8705), .IN2(n8706), .QN(g30654) );
  NAND2X0 U8464 ( .IN1(test_so34), .IN2(n7267), .QN(n8706) );
  NAND2X0 U8465 ( .IN1(n8707), .IN2(test_so31), .QN(n8705) );
  NAND2X0 U8466 ( .IN1(n8708), .IN2(n8709), .QN(g30653) );
  NAND2X0 U8467 ( .IN1(n4369), .IN2(g246), .QN(n8709) );
  NAND2X0 U8468 ( .IN1(n8710), .IN2(g165), .QN(n8708) );
  NAND2X0 U8469 ( .IN1(n8711), .IN2(n8712), .QN(g30652) );
  NAND2X0 U8470 ( .IN1(n4324), .IN2(g2297), .QN(n8712) );
  NAND2X0 U8471 ( .IN1(n8666), .IN2(g6837), .QN(n8711) );
  NAND3X0 U8472 ( .IN1(n8713), .IN2(n8714), .IN3(n8555), .QN(n8666) );
  NAND2X0 U8473 ( .IN1(n8686), .IN2(n8715), .QN(n8555) );
  INVX0 U8474 ( .INP(n4529), .ZN(n8715) );
  NAND2X0 U8475 ( .IN1(n8716), .IN2(n8557), .QN(n8714) );
  XOR2X1 U8476 ( .IN1(n7770), .IN2(n8350), .Q(n8716) );
  NOR2X0 U8477 ( .IN1(n8717), .IN2(n8718), .QN(n8350) );
  XOR2X1 U8478 ( .IN1(n4529), .IN2(n7764), .Q(n8718) );
  NAND2X0 U8479 ( .IN1(n8559), .IN2(n8719), .QN(n8713) );
  NAND2X0 U8480 ( .IN1(n8720), .IN2(n8721), .QN(g30651) );
  NAND2X0 U8481 ( .IN1(n4317), .IN2(g1612), .QN(n8721) );
  NAND2X0 U8482 ( .IN1(n8671), .IN2(g6573), .QN(n8720) );
  AND3X1 U8483 ( .IN1(n8722), .IN2(n8601), .IN3(n8723), .Q(n8671) );
  NAND2X0 U8484 ( .IN1(n8586), .IN2(n4374), .QN(n8723) );
  NAND2X0 U8485 ( .IN1(n8724), .IN2(n4530), .QN(n8601) );
  NAND2X0 U8486 ( .IN1(n8583), .IN2(n8725), .QN(n8722) );
  XOR2X1 U8487 ( .IN1(n7732), .IN2(n8726), .Q(n8725) );
  AND2X1 U8488 ( .IN1(n8727), .IN2(n8728), .Q(n8726) );
  NAND2X0 U8489 ( .IN1(n8729), .IN2(n8730), .QN(g30650) );
  NAND2X0 U8490 ( .IN1(test_so56), .IN2(n4515), .QN(n8730) );
  NAND2X0 U8491 ( .IN1(n8702), .IN2(g6782), .QN(n8729) );
  NAND2X0 U8492 ( .IN1(n8731), .IN2(n8732), .QN(g30649) );
  NAND2X0 U8493 ( .IN1(n4323), .IN2(g927), .QN(n8732) );
  NAND2X0 U8494 ( .IN1(n8674), .IN2(g6368), .QN(n8731) );
  AND3X1 U8495 ( .IN1(n8733), .IN2(n8632), .IN3(n8734), .Q(n8674) );
  NAND2X0 U8496 ( .IN1(n8615), .IN2(n4391), .QN(n8734) );
  NAND2X0 U8497 ( .IN1(n8613), .IN2(n8735), .QN(n8733) );
  XOR2X1 U8498 ( .IN1(n7713), .IN2(n8736), .Q(n8735) );
  NAND2X0 U8499 ( .IN1(n8614), .IN2(n8737), .QN(n8736) );
  NAND2X0 U8500 ( .IN1(n8738), .IN2(n8739), .QN(g30648) );
  NAND2X0 U8501 ( .IN1(n4312), .IN2(g921), .QN(n8739) );
  NAND2X0 U8502 ( .IN1(n8707), .IN2(g6518), .QN(n8738) );
  NAND2X0 U8503 ( .IN1(n8740), .IN2(n8741), .QN(g30647) );
  NAND2X0 U8504 ( .IN1(g915), .IN2(n7267), .QN(n8741) );
  NAND2X0 U8505 ( .IN1(test_so31), .IN2(n8742), .QN(n8740) );
  NAND2X0 U8506 ( .IN1(n8743), .IN2(n8744), .QN(g30646) );
  NAND2X0 U8507 ( .IN1(n4512), .IN2(g243), .QN(n8744) );
  NAND2X0 U8508 ( .IN1(n8710), .IN2(g6313), .QN(n8743) );
  NAND2X0 U8509 ( .IN1(n8745), .IN2(n8746), .QN(g30645) );
  NAND2X0 U8510 ( .IN1(n4369), .IN2(g237), .QN(n8746) );
  NAND2X0 U8511 ( .IN1(n8747), .IN2(g165), .QN(n8745) );
  NAND2X0 U8512 ( .IN1(n8748), .IN2(n8749), .QN(g30644) );
  NAND2X0 U8513 ( .IN1(n4317), .IN2(g1603), .QN(n8749) );
  NAND2X0 U8514 ( .IN1(n8702), .IN2(g6573), .QN(n8748) );
  NAND3X0 U8515 ( .IN1(n8750), .IN2(n8751), .IN3(n8581), .QN(n8702) );
  NAND2X0 U8516 ( .IN1(n8724), .IN2(n8752), .QN(n8581) );
  INVX0 U8517 ( .INP(n4530), .ZN(n8752) );
  NAND2X0 U8518 ( .IN1(n8753), .IN2(n8583), .QN(n8751) );
  XOR2X1 U8519 ( .IN1(n2685), .IN2(n7744), .Q(n8753) );
  NAND2X0 U8520 ( .IN1(n8754), .IN2(n8755), .QN(n2685) );
  XOR2X1 U8521 ( .IN1(n8347), .IN2(n7731), .Q(n8755) );
  NAND2X0 U8522 ( .IN1(n8586), .IN2(n8756), .QN(n8750) );
  NAND2X0 U8523 ( .IN1(n8757), .IN2(n8758), .QN(g30643) );
  NAND2X0 U8524 ( .IN1(n4323), .IN2(g918), .QN(n8758) );
  NAND2X0 U8525 ( .IN1(n8707), .IN2(g6368), .QN(n8757) );
  AND3X1 U8526 ( .IN1(n8759), .IN2(n8632), .IN3(n8760), .Q(n8707) );
  NAND2X0 U8527 ( .IN1(n8615), .IN2(n4375), .QN(n8760) );
  NAND2X0 U8528 ( .IN1(n8761), .IN2(n8762), .QN(n8632) );
  NAND2X0 U8529 ( .IN1(n8613), .IN2(n8763), .QN(n8759) );
  XOR2X1 U8530 ( .IN1(n8764), .IN2(n8765), .Q(n8763) );
  AND2X1 U8531 ( .IN1(n8766), .IN2(n8767), .Q(n8765) );
  NAND2X0 U8532 ( .IN1(n8768), .IN2(n8769), .QN(g30642) );
  NAND2X0 U8533 ( .IN1(n4312), .IN2(g912), .QN(n8769) );
  NAND2X0 U8534 ( .IN1(n8742), .IN2(g6518), .QN(n8768) );
  NAND2X0 U8535 ( .IN1(n8770), .IN2(n8771), .QN(g30641) );
  NAND2X0 U8536 ( .IN1(n4318), .IN2(g240), .QN(n8771) );
  NAND2X0 U8537 ( .IN1(n8710), .IN2(g6231), .QN(n8770) );
  AND3X1 U8538 ( .IN1(n8772), .IN2(n8678), .IN3(n8773), .Q(n8710) );
  NAND2X0 U8539 ( .IN1(n8653), .IN2(n4392), .QN(n8773) );
  NAND2X0 U8540 ( .IN1(n8650), .IN2(n8774), .QN(n8772) );
  XOR2X1 U8541 ( .IN1(n8775), .IN2(n8776), .Q(n8774) );
  NAND2X0 U8542 ( .IN1(n8652), .IN2(n8777), .QN(n8776) );
  NAND2X0 U8543 ( .IN1(n8778), .IN2(n8779), .QN(g30640) );
  NAND2X0 U8544 ( .IN1(n4512), .IN2(g234), .QN(n8779) );
  NAND2X0 U8545 ( .IN1(n8747), .IN2(g6313), .QN(n8778) );
  NAND2X0 U8546 ( .IN1(n8780), .IN2(n8781), .QN(g30639) );
  NAND2X0 U8547 ( .IN1(n4369), .IN2(g228), .QN(n8781) );
  NAND2X0 U8548 ( .IN1(n8782), .IN2(g165), .QN(n8780) );
  NAND2X0 U8549 ( .IN1(n8783), .IN2(n8784), .QN(g30638) );
  NAND2X0 U8550 ( .IN1(n4323), .IN2(g909), .QN(n8784) );
  NAND2X0 U8551 ( .IN1(n8742), .IN2(g6368), .QN(n8783) );
  NAND3X0 U8552 ( .IN1(n8785), .IN2(n8786), .IN3(n8611), .QN(n8742) );
  NAND2X0 U8553 ( .IN1(n8761), .IN2(n8640), .QN(n8611) );
  NAND2X0 U8554 ( .IN1(n8787), .IN2(n8613), .QN(n8786) );
  XOR2X1 U8555 ( .IN1(n8639), .IN2(n8641), .Q(n8787) );
  NAND2X0 U8556 ( .IN1(n8788), .IN2(n8789), .QN(n8639) );
  XOR2X1 U8557 ( .IN1(n7716), .IN2(n8640), .Q(n8789) );
  NAND2X0 U8558 ( .IN1(n8615), .IN2(n8790), .QN(n8785) );
  NAND2X0 U8559 ( .IN1(n8791), .IN2(n8792), .QN(g30637) );
  NAND2X0 U8560 ( .IN1(n4318), .IN2(g231), .QN(n8792) );
  NAND2X0 U8561 ( .IN1(n8747), .IN2(g6231), .QN(n8791) );
  AND3X1 U8562 ( .IN1(n8793), .IN2(n8678), .IN3(n8794), .Q(n8747) );
  NAND2X0 U8563 ( .IN1(n8653), .IN2(n4376), .QN(n8794) );
  NAND2X0 U8564 ( .IN1(n8795), .IN2(n8796), .QN(n8678) );
  NAND2X0 U8565 ( .IN1(n8650), .IN2(n8797), .QN(n8793) );
  XOR2X1 U8566 ( .IN1(n7674), .IN2(n8798), .Q(n8797) );
  AND2X1 U8567 ( .IN1(n8799), .IN2(n8800), .Q(n8798) );
  NAND2X0 U8568 ( .IN1(n8801), .IN2(n8802), .QN(g30636) );
  NAND2X0 U8569 ( .IN1(n4512), .IN2(g225), .QN(n8802) );
  NAND2X0 U8570 ( .IN1(n8782), .IN2(g6313), .QN(n8801) );
  NAND2X0 U8571 ( .IN1(n8803), .IN2(n8804), .QN(g30635) );
  NAND2X0 U8572 ( .IN1(n4318), .IN2(g222), .QN(n8804) );
  NAND2X0 U8573 ( .IN1(n8782), .IN2(g6231), .QN(n8803) );
  NAND3X0 U8574 ( .IN1(n8805), .IN2(n8806), .IN3(n8648), .QN(n8782) );
  NAND2X0 U8575 ( .IN1(n8795), .IN2(n8346), .QN(n8648) );
  NAND2X0 U8576 ( .IN1(n8807), .IN2(n8650), .QN(n8806) );
  XOR2X1 U8577 ( .IN1(n2718), .IN2(n7685), .Q(n8807) );
  NAND2X0 U8578 ( .IN1(n8808), .IN2(n8809), .QN(n2718) );
  XOR2X1 U8579 ( .IN1(n7673), .IN2(n8346), .Q(n8809) );
  NAND2X0 U8580 ( .IN1(n8653), .IN2(n8810), .QN(n8805) );
  NAND2X0 U8581 ( .IN1(n8811), .IN2(n8812), .QN(g30566) );
  NAND2X0 U8582 ( .IN1(n8448), .IN2(n4606), .QN(n8812) );
  AND2X1 U8583 ( .IN1(n8813), .IN2(n8814), .Q(n8448) );
  XOR2X1 U8584 ( .IN1(n8815), .IN2(n8816), .Q(n8813) );
  NAND2X0 U8585 ( .IN1(n8817), .IN2(n8818), .QN(n8816) );
  NAND2X0 U8586 ( .IN1(n8819), .IN2(n8820), .QN(n8818) );
  NAND4X0 U8587 ( .IN1(n8821), .IN2(n8822), .IN3(n8823), .IN4(n8824), .QN(
        n8817) );
  NAND3X0 U8588 ( .IN1(n8825), .IN2(n8826), .IN3(n8827), .QN(n8823) );
  OR2X1 U8589 ( .IN1(n8828), .IN2(n8829), .Q(n8822) );
  NAND2X0 U8590 ( .IN1(n8830), .IN2(n8829), .QN(n8821) );
  NAND2X0 U8591 ( .IN1(n8831), .IN2(n8832), .QN(n8830) );
  NAND2X0 U8592 ( .IN1(n8825), .IN2(n8833), .QN(n8832) );
  NAND3X0 U8593 ( .IN1(n8834), .IN2(n8826), .IN3(n8835), .QN(n8833) );
  INVX0 U8594 ( .INP(n8836), .ZN(n8835) );
  NAND2X0 U8595 ( .IN1(n8828), .IN2(n8837), .QN(n8834) );
  NAND2X0 U8596 ( .IN1(n8838), .IN2(n8839), .QN(n8831) );
  NAND2X0 U8597 ( .IN1(n2792), .IN2(n8840), .QN(n8838) );
  OR2X1 U8598 ( .IN1(n8841), .IN2(n6542), .Q(n8811) );
  NAND2X0 U8599 ( .IN1(n8842), .IN2(n8843), .QN(g30505) );
  NAND2X0 U8600 ( .IN1(n8844), .IN2(g5555), .QN(n8843) );
  OR2X1 U8601 ( .IN1(n8456), .IN2(n6541), .Q(n8842) );
  NAND2X0 U8602 ( .IN1(n8845), .IN2(n8846), .QN(g30503) );
  NAND2X0 U8603 ( .IN1(n8847), .IN2(g7014), .QN(n8846) );
  OR2X1 U8604 ( .IN1(n8459), .IN2(n6534), .Q(n8845) );
  NAND2X0 U8605 ( .IN1(n8848), .IN2(n8849), .QN(g30500) );
  NAND2X0 U8606 ( .IN1(n2798), .IN2(g1088), .QN(n8849) );
  NAND2X0 U8607 ( .IN1(test_so39), .IN2(n4381), .QN(n8848) );
  NAND2X0 U8608 ( .IN1(n8850), .IN2(n8851), .QN(g30487) );
  NAND2X0 U8609 ( .IN1(n8847), .IN2(g5511), .QN(n8851) );
  OR2X1 U8610 ( .IN1(n8494), .IN2(n6547), .Q(n8850) );
  NAND2X0 U8611 ( .IN1(n8852), .IN2(n8853), .QN(g30485) );
  OR2X1 U8612 ( .IN1(g6712), .IN2(n6537), .Q(n8853) );
  NAND2X0 U8613 ( .IN1(n2798), .IN2(g6712), .QN(n8852) );
  NAND2X0 U8614 ( .IN1(n8854), .IN2(n8855), .QN(g30482) );
  NAND2X0 U8615 ( .IN1(n8856), .IN2(n4640), .QN(n8855) );
  OR2X1 U8616 ( .IN1(n8500), .IN2(n6557), .Q(n8854) );
  NAND2X0 U8617 ( .IN1(n8857), .IN2(n8858), .QN(g30470) );
  OR2X1 U8618 ( .IN1(g5472), .IN2(n6552), .Q(n8858) );
  NAND2X0 U8619 ( .IN1(n2798), .IN2(g5472), .QN(n8857) );
  NAND2X0 U8620 ( .IN1(n8859), .IN2(n8860), .QN(g30468) );
  NAND2X0 U8621 ( .IN1(n8856), .IN2(g6447), .QN(n8860) );
  OR2X1 U8622 ( .IN1(n8861), .IN2(n6558), .Q(n8859) );
  NAND2X0 U8623 ( .IN1(n8862), .IN2(n8863), .QN(g30455) );
  NAND2X0 U8624 ( .IN1(n8856), .IN2(g5437), .QN(n8863) );
  AND2X1 U8625 ( .IN1(n8864), .IN2(n8508), .Q(n8856) );
  XOR2X1 U8626 ( .IN1(n8865), .IN2(n8519), .Q(n8864) );
  NAND2X0 U8627 ( .IN1(n8866), .IN2(n8867), .QN(n8865) );
  NAND2X0 U8628 ( .IN1(n8519), .IN2(n8868), .QN(n8867) );
  NAND3X0 U8629 ( .IN1(n8869), .IN2(n8870), .IN3(n8518), .QN(n8868) );
  NAND2X0 U8630 ( .IN1(n8530), .IN2(n8509), .QN(n8870) );
  NAND2X0 U8631 ( .IN1(n8536), .IN2(n8871), .QN(n8530) );
  OR2X1 U8632 ( .IN1(n8872), .IN2(n8873), .Q(n8871) );
  NAND3X0 U8633 ( .IN1(n8874), .IN2(g309), .IN3(n8523), .QN(n8869) );
  NAND3X0 U8634 ( .IN1(n8521), .IN2(n8518), .IN3(n8534), .QN(n8866) );
  AND3X1 U8635 ( .IN1(n8872), .IN2(n8509), .IN3(n3130), .Q(n8521) );
  OR2X1 U8636 ( .IN1(n8537), .IN2(n6559), .Q(n8862) );
  NAND2X0 U8637 ( .IN1(n8875), .IN2(n8876), .QN(g30356) );
  NAND2X0 U8638 ( .IN1(n8844), .IN2(n4606), .QN(n8876) );
  OR2X1 U8639 ( .IN1(n8841), .IN2(n6540), .Q(n8875) );
  NAND2X0 U8640 ( .IN1(n8877), .IN2(n8878), .QN(g30341) );
  NAND2X0 U8641 ( .IN1(n8844), .IN2(g7264), .QN(n8878) );
  AND2X1 U8642 ( .IN1(n8879), .IN2(n8814), .Q(n8844) );
  XOR2X1 U8643 ( .IN1(n8880), .IN2(n8825), .Q(n8879) );
  NAND2X0 U8644 ( .IN1(n8881), .IN2(n8882), .QN(n8880) );
  NAND2X0 U8645 ( .IN1(n8825), .IN2(n8883), .QN(n8882) );
  NAND3X0 U8646 ( .IN1(n8884), .IN2(n8885), .IN3(n8824), .QN(n8883) );
  NAND2X0 U8647 ( .IN1(n8836), .IN2(n8815), .QN(n8885) );
  NAND2X0 U8648 ( .IN1(n8840), .IN2(n8886), .QN(n8836) );
  NAND2X0 U8649 ( .IN1(n8887), .IN2(n3038), .QN(n8886) );
  INVX0 U8650 ( .INP(n8888), .ZN(n8887) );
  NAND3X0 U8651 ( .IN1(n8889), .IN2(test_so79), .IN3(n8829), .QN(n8884) );
  NAND3X0 U8652 ( .IN1(n8827), .IN2(n8824), .IN3(n8839), .QN(n8881) );
  AND3X1 U8653 ( .IN1(n8888), .IN2(n8815), .IN3(n3038), .Q(n8827) );
  OR2X1 U8654 ( .IN1(n8449), .IN2(n6531), .Q(n8877) );
  NAND2X0 U8655 ( .IN1(n8890), .IN2(n8891), .QN(g30338) );
  NAND2X0 U8656 ( .IN1(n8847), .IN2(n4618), .QN(n8891) );
  AND2X1 U8657 ( .IN1(n8892), .IN2(n8465), .Q(n8847) );
  XOR2X1 U8658 ( .IN1(n8893), .IN2(n8476), .Q(n8892) );
  NAND2X0 U8659 ( .IN1(n8894), .IN2(n8895), .QN(n8893) );
  NAND2X0 U8660 ( .IN1(n8476), .IN2(n8896), .QN(n8895) );
  NAND3X0 U8661 ( .IN1(n8897), .IN2(n8898), .IN3(n8475), .QN(n8896) );
  NAND2X0 U8662 ( .IN1(n8487), .IN2(n8466), .QN(n8898) );
  NAND2X0 U8663 ( .IN1(n8493), .IN2(n8899), .QN(n8487) );
  OR2X1 U8664 ( .IN1(n8900), .IN2(n8901), .Q(n8899) );
  NAND3X0 U8665 ( .IN1(n8902), .IN2(g1690), .IN3(n8480), .QN(n8897) );
  NAND3X0 U8666 ( .IN1(n8478), .IN2(n8475), .IN3(n8491), .QN(n8894) );
  AND3X1 U8667 ( .IN1(n8900), .IN2(n8466), .IN3(n3070), .Q(n8478) );
  OR2X1 U8668 ( .IN1(n8453), .IN2(n6546), .Q(n8890) );
  NAND2X0 U8669 ( .IN1(n8903), .IN2(n8904), .QN(g30304) );
  NAND2X0 U8670 ( .IN1(n4367), .IN2(g2285), .QN(n8904) );
  NAND2X0 U8671 ( .IN1(n8905), .IN2(g2241), .QN(n8903) );
  NAND2X0 U8672 ( .IN1(n8906), .IN2(n8907), .QN(g30303) );
  NAND2X0 U8673 ( .IN1(g2282), .IN2(n7266), .QN(n8907) );
  NAND2X0 U8674 ( .IN1(test_so73), .IN2(n8905), .QN(n8906) );
  NAND2X0 U8675 ( .IN1(n8908), .IN2(n8909), .QN(g30302) );
  NAND2X0 U8676 ( .IN1(n4368), .IN2(g1591), .QN(n8909) );
  NAND2X0 U8677 ( .IN1(n8910), .IN2(g1547), .QN(n8908) );
  NAND2X0 U8678 ( .IN1(n8911), .IN2(n8912), .QN(g30301) );
  NAND2X0 U8679 ( .IN1(n4324), .IN2(g2279), .QN(n8912) );
  NAND2X0 U8680 ( .IN1(n8905), .IN2(g6837), .QN(n8911) );
  NAND2X0 U8681 ( .IN1(n8913), .IN2(n8914), .QN(n8905) );
  NAND2X0 U8682 ( .IN1(n8915), .IN2(n8557), .QN(n8914) );
  XOR2X1 U8683 ( .IN1(n7771), .IN2(n8916), .Q(n8915) );
  NAND2X0 U8684 ( .IN1(n8559), .IN2(g2185), .QN(n8913) );
  NAND2X0 U8685 ( .IN1(n8917), .IN2(n8918), .QN(g30300) );
  NAND2X0 U8686 ( .IN1(n4367), .IN2(g2267), .QN(n8918) );
  NAND2X0 U8687 ( .IN1(n8919), .IN2(g2241), .QN(n8917) );
  NAND2X0 U8688 ( .IN1(n8920), .IN2(n8921), .QN(g30299) );
  NAND2X0 U8689 ( .IN1(n4515), .IN2(g1588), .QN(n8921) );
  NAND2X0 U8690 ( .IN1(n8910), .IN2(g6782), .QN(n8920) );
  NAND2X0 U8691 ( .IN1(n8922), .IN2(n8923), .QN(g30298) );
  NAND2X0 U8692 ( .IN1(g897), .IN2(n7267), .QN(n8923) );
  NAND2X0 U8693 ( .IN1(test_so31), .IN2(n8924), .QN(n8922) );
  NAND2X0 U8694 ( .IN1(n8925), .IN2(n8926), .QN(g30297) );
  NAND2X0 U8695 ( .IN1(n4367), .IN2(g2339), .QN(n8926) );
  NAND2X0 U8696 ( .IN1(n8927), .IN2(g2241), .QN(n8925) );
  NAND2X0 U8697 ( .IN1(n8928), .IN2(n8929), .QN(g30296) );
  NAND2X0 U8698 ( .IN1(test_so76), .IN2(n7266), .QN(n8929) );
  NAND2X0 U8699 ( .IN1(test_so73), .IN2(n8919), .QN(n8928) );
  NAND2X0 U8700 ( .IN1(n8930), .IN2(n8931), .QN(g30295) );
  NAND2X0 U8701 ( .IN1(n4317), .IN2(g1585), .QN(n8931) );
  NAND2X0 U8702 ( .IN1(n8910), .IN2(g6573), .QN(n8930) );
  NAND2X0 U8703 ( .IN1(n8932), .IN2(n8933), .QN(n8910) );
  NAND2X0 U8704 ( .IN1(n8934), .IN2(n8583), .QN(n8933) );
  XOR2X1 U8705 ( .IN1(n8935), .IN2(n8936), .Q(n8934) );
  NAND2X0 U8706 ( .IN1(n8586), .IN2(g1491), .QN(n8932) );
  NAND2X0 U8707 ( .IN1(n8937), .IN2(n8938), .QN(g30294) );
  NAND2X0 U8708 ( .IN1(n4368), .IN2(g1573), .QN(n8938) );
  NAND2X0 U8709 ( .IN1(n8939), .IN2(g1547), .QN(n8937) );
  NAND2X0 U8710 ( .IN1(n8940), .IN2(n8941), .QN(g30293) );
  NAND2X0 U8711 ( .IN1(n4312), .IN2(g894), .QN(n8941) );
  NAND2X0 U8712 ( .IN1(n8924), .IN2(g6518), .QN(n8940) );
  NAND2X0 U8713 ( .IN1(n8942), .IN2(n8943), .QN(g30292) );
  NAND2X0 U8714 ( .IN1(n4369), .IN2(g210), .QN(n8943) );
  NAND2X0 U8715 ( .IN1(n8944), .IN2(g165), .QN(n8942) );
  NAND2X0 U8716 ( .IN1(n8945), .IN2(n8946), .QN(g30291) );
  NAND2X0 U8717 ( .IN1(g2336), .IN2(n7266), .QN(n8946) );
  NAND2X0 U8718 ( .IN1(test_so73), .IN2(n8927), .QN(n8945) );
  NAND2X0 U8719 ( .IN1(n8947), .IN2(n8948), .QN(g30290) );
  NAND2X0 U8720 ( .IN1(n4367), .IN2(g2330), .QN(n8948) );
  NAND2X0 U8721 ( .IN1(n8949), .IN2(g2241), .QN(n8947) );
  NAND2X0 U8722 ( .IN1(n8950), .IN2(n8951), .QN(g30289) );
  NAND2X0 U8723 ( .IN1(n4324), .IN2(g2261), .QN(n8951) );
  NAND2X0 U8724 ( .IN1(n8919), .IN2(g6837), .QN(n8950) );
  NAND2X0 U8725 ( .IN1(n8952), .IN2(n8953), .QN(n8919) );
  NAND2X0 U8726 ( .IN1(n8557), .IN2(n8954), .QN(n8953) );
  XNOR2X1 U8727 ( .IN1(n7765), .IN2(n8955), .Q(n8954) );
  NAND2X0 U8728 ( .IN1(n8559), .IN2(g2165), .QN(n8952) );
  NAND2X0 U8729 ( .IN1(n8956), .IN2(n8957), .QN(g30288) );
  NAND2X0 U8730 ( .IN1(n4368), .IN2(g1645), .QN(n8957) );
  NAND2X0 U8731 ( .IN1(n8958), .IN2(g1547), .QN(n8956) );
  NAND2X0 U8732 ( .IN1(n8959), .IN2(n8960), .QN(g30287) );
  NAND2X0 U8733 ( .IN1(n4515), .IN2(g1570), .QN(n8960) );
  NAND2X0 U8734 ( .IN1(n8939), .IN2(g6782), .QN(n8959) );
  NAND2X0 U8735 ( .IN1(n8961), .IN2(n8962), .QN(g30286) );
  NAND2X0 U8736 ( .IN1(n4323), .IN2(g891), .QN(n8962) );
  NAND2X0 U8737 ( .IN1(n8924), .IN2(g6368), .QN(n8961) );
  NAND2X0 U8738 ( .IN1(n8963), .IN2(n8964), .QN(n8924) );
  NAND2X0 U8739 ( .IN1(n8965), .IN2(n8613), .QN(n8964) );
  XOR2X1 U8740 ( .IN1(n8966), .IN2(n8967), .Q(n8965) );
  NAND2X0 U8741 ( .IN1(n8615), .IN2(g801), .QN(n8963) );
  NAND2X0 U8742 ( .IN1(n8968), .IN2(n8969), .QN(g30285) );
  NAND2X0 U8743 ( .IN1(g879), .IN2(n7267), .QN(n8969) );
  NAND2X0 U8744 ( .IN1(test_so31), .IN2(n8970), .QN(n8968) );
  NAND2X0 U8745 ( .IN1(n8971), .IN2(n8972), .QN(g30284) );
  NAND2X0 U8746 ( .IN1(n4512), .IN2(g207), .QN(n8972) );
  NAND2X0 U8747 ( .IN1(n8944), .IN2(g6313), .QN(n8971) );
  NAND2X0 U8748 ( .IN1(n8973), .IN2(n8974), .QN(g30283) );
  NAND2X0 U8749 ( .IN1(n4324), .IN2(g2333), .QN(n8974) );
  NAND2X0 U8750 ( .IN1(n8927), .IN2(g6837), .QN(n8973) );
  NAND2X0 U8751 ( .IN1(n8975), .IN2(n8976), .QN(n8927) );
  NAND3X0 U8752 ( .IN1(n8557), .IN2(n8977), .IN3(n8978), .QN(n8976) );
  XNOR2X1 U8753 ( .IN1(n8717), .IN2(n7764), .Q(n8978) );
  NAND2X0 U8754 ( .IN1(n8979), .IN2(n8980), .QN(n8717) );
  XOR2X1 U8755 ( .IN1(n8349), .IN2(n7763), .Q(n8980) );
  NAND2X0 U8756 ( .IN1(n8559), .IN2(g2200), .QN(n8975) );
  NAND2X0 U8757 ( .IN1(n8981), .IN2(n8982), .QN(g30282) );
  NAND2X0 U8758 ( .IN1(test_so77), .IN2(n7266), .QN(n8982) );
  NAND2X0 U8759 ( .IN1(test_so73), .IN2(n8949), .QN(n8981) );
  NAND2X0 U8760 ( .IN1(n8983), .IN2(n8984), .QN(g30281) );
  NAND2X0 U8761 ( .IN1(n4515), .IN2(g1642), .QN(n8984) );
  NAND2X0 U8762 ( .IN1(n8958), .IN2(g6782), .QN(n8983) );
  NAND2X0 U8763 ( .IN1(n8985), .IN2(n8986), .QN(g30280) );
  NAND2X0 U8764 ( .IN1(n4368), .IN2(g1636), .QN(n8986) );
  NAND2X0 U8765 ( .IN1(n8987), .IN2(g1547), .QN(n8985) );
  NAND2X0 U8766 ( .IN1(n8988), .IN2(n8989), .QN(g30279) );
  NAND2X0 U8767 ( .IN1(n4317), .IN2(g1567), .QN(n8989) );
  NAND2X0 U8768 ( .IN1(n8939), .IN2(g6573), .QN(n8988) );
  NAND2X0 U8769 ( .IN1(n8990), .IN2(n8991), .QN(n8939) );
  NAND2X0 U8770 ( .IN1(n8583), .IN2(n8992), .QN(n8991) );
  XOR2X1 U8771 ( .IN1(n7743), .IN2(n8727), .Q(n8992) );
  NAND2X0 U8772 ( .IN1(n8586), .IN2(g1471), .QN(n8990) );
  NAND2X0 U8773 ( .IN1(n8993), .IN2(n8994), .QN(g30278) );
  NAND2X0 U8774 ( .IN1(g951), .IN2(n7267), .QN(n8994) );
  NAND2X0 U8775 ( .IN1(test_so31), .IN2(n8995), .QN(n8993) );
  NAND2X0 U8776 ( .IN1(n8996), .IN2(n8997), .QN(g30277) );
  NAND2X0 U8777 ( .IN1(n4312), .IN2(g876), .QN(n8997) );
  NAND2X0 U8778 ( .IN1(n8970), .IN2(g6518), .QN(n8996) );
  NAND2X0 U8779 ( .IN1(n8998), .IN2(n8999), .QN(g30276) );
  NAND2X0 U8780 ( .IN1(n4318), .IN2(g204), .QN(n8999) );
  NAND2X0 U8781 ( .IN1(n8944), .IN2(g6231), .QN(n8998) );
  NAND2X0 U8782 ( .IN1(n9000), .IN2(n9001), .QN(n8944) );
  NAND2X0 U8783 ( .IN1(n9002), .IN2(n8650), .QN(n9001) );
  XOR2X1 U8784 ( .IN1(n9003), .IN2(n7684), .Q(n9002) );
  NAND2X0 U8785 ( .IN1(n8653), .IN2(g113), .QN(n9000) );
  NAND2X0 U8786 ( .IN1(n9004), .IN2(n9005), .QN(g30275) );
  NAND2X0 U8787 ( .IN1(n4369), .IN2(g192), .QN(n9005) );
  NAND2X0 U8788 ( .IN1(n9006), .IN2(g165), .QN(n9004) );
  NAND2X0 U8789 ( .IN1(n9007), .IN2(n9008), .QN(g30274) );
  NAND2X0 U8790 ( .IN1(n4324), .IN2(g2324), .QN(n9008) );
  NAND2X0 U8791 ( .IN1(n8949), .IN2(g6837), .QN(n9007) );
  NAND2X0 U8792 ( .IN1(n9009), .IN2(n9010), .QN(n8949) );
  NAND3X0 U8793 ( .IN1(n8557), .IN2(n8977), .IN3(n9011), .QN(n9010) );
  XOR2X1 U8794 ( .IN1(n7758), .IN2(n9012), .Q(n9011) );
  NOR2X0 U8795 ( .IN1(n9013), .IN2(n9014), .QN(n9012) );
  NOR2X0 U8796 ( .IN1(n7771), .IN2(n8349), .QN(n9013) );
  NAND2X0 U8797 ( .IN1(n8559), .IN2(g2190), .QN(n9009) );
  NAND2X0 U8798 ( .IN1(n9015), .IN2(n9016), .QN(g30273) );
  NAND2X0 U8799 ( .IN1(n4317), .IN2(g1639), .QN(n9016) );
  NAND2X0 U8800 ( .IN1(n8958), .IN2(g6573), .QN(n9015) );
  NAND2X0 U8801 ( .IN1(n9017), .IN2(n9018), .QN(n8958) );
  NAND3X0 U8802 ( .IN1(n8583), .IN2(n9019), .IN3(n9020), .QN(n9018) );
  XOR2X1 U8803 ( .IN1(n7731), .IN2(n8754), .Q(n9020) );
  NOR2X0 U8804 ( .IN1(n9021), .IN2(n9022), .QN(n8754) );
  XOR2X1 U8805 ( .IN1(n4530), .IN2(n9023), .Q(n9022) );
  NAND2X0 U8806 ( .IN1(n8586), .IN2(g1506), .QN(n9017) );
  NAND2X0 U8807 ( .IN1(n9024), .IN2(n9025), .QN(g30272) );
  NAND2X0 U8808 ( .IN1(n4515), .IN2(g1633), .QN(n9025) );
  NAND2X0 U8809 ( .IN1(n8987), .IN2(g6782), .QN(n9024) );
  NAND2X0 U8810 ( .IN1(n9026), .IN2(n9027), .QN(g30271) );
  NAND2X0 U8811 ( .IN1(n4312), .IN2(g948), .QN(n9027) );
  NAND2X0 U8812 ( .IN1(n8995), .IN2(g6518), .QN(n9026) );
  NAND2X0 U8813 ( .IN1(n9028), .IN2(n9029), .QN(g30270) );
  NAND2X0 U8814 ( .IN1(g942), .IN2(n7267), .QN(n9029) );
  NAND2X0 U8815 ( .IN1(test_so31), .IN2(n9030), .QN(n9028) );
  NAND2X0 U8816 ( .IN1(n9031), .IN2(n9032), .QN(g30269) );
  NAND2X0 U8817 ( .IN1(n4323), .IN2(g873), .QN(n9032) );
  NAND2X0 U8818 ( .IN1(n8970), .IN2(g6368), .QN(n9031) );
  NAND2X0 U8819 ( .IN1(n9033), .IN2(n9034), .QN(n8970) );
  NAND2X0 U8820 ( .IN1(n8613), .IN2(n9035), .QN(n9034) );
  XOR2X1 U8821 ( .IN1(n7711), .IN2(n8766), .Q(n9035) );
  NAND2X0 U8822 ( .IN1(n8615), .IN2(g785), .QN(n9033) );
  NAND2X0 U8823 ( .IN1(n9036), .IN2(n9037), .QN(g30268) );
  NAND2X0 U8824 ( .IN1(n4369), .IN2(g264), .QN(n9037) );
  NAND2X0 U8825 ( .IN1(n9038), .IN2(g165), .QN(n9036) );
  NAND2X0 U8826 ( .IN1(n9039), .IN2(n9040), .QN(g30267) );
  NAND2X0 U8827 ( .IN1(test_so13), .IN2(n4512), .QN(n9040) );
  NAND2X0 U8828 ( .IN1(n9006), .IN2(g6313), .QN(n9039) );
  NAND2X0 U8829 ( .IN1(n9041), .IN2(n9042), .QN(g30266) );
  NAND2X0 U8830 ( .IN1(n4317), .IN2(g1630), .QN(n9042) );
  NAND2X0 U8831 ( .IN1(n8987), .IN2(g6573), .QN(n9041) );
  NAND2X0 U8832 ( .IN1(n9043), .IN2(n9044), .QN(n8987) );
  NAND3X0 U8833 ( .IN1(n8583), .IN2(n9019), .IN3(n9045), .QN(n9044) );
  XNOR2X1 U8834 ( .IN1(n9046), .IN2(n7734), .Q(n9045) );
  NAND2X0 U8835 ( .IN1(n9047), .IN2(n9048), .QN(n9046) );
  NAND2X0 U8836 ( .IN1(n4530), .IN2(n8936), .QN(n9048) );
  NAND2X0 U8837 ( .IN1(n8586), .IN2(g1496), .QN(n9043) );
  NAND2X0 U8838 ( .IN1(n9049), .IN2(n9050), .QN(g30265) );
  NAND2X0 U8839 ( .IN1(test_so35), .IN2(n4323), .QN(n9050) );
  NAND2X0 U8840 ( .IN1(n8995), .IN2(g6368), .QN(n9049) );
  NAND2X0 U8841 ( .IN1(n9051), .IN2(n9052), .QN(n8995) );
  NAND2X0 U8842 ( .IN1(n9053), .IN2(n8613), .QN(n9052) );
  XOR2X1 U8843 ( .IN1(n7716), .IN2(n8788), .Q(n9053) );
  NOR2X0 U8844 ( .IN1(n9054), .IN2(n9055), .QN(n8788) );
  XOR2X1 U8845 ( .IN1(n9056), .IN2(n8640), .Q(n9055) );
  NAND2X0 U8846 ( .IN1(n8615), .IN2(g813), .QN(n9051) );
  NAND2X0 U8847 ( .IN1(n9057), .IN2(n9058), .QN(g30264) );
  NAND2X0 U8848 ( .IN1(n4312), .IN2(g939), .QN(n9058) );
  NAND2X0 U8849 ( .IN1(n9030), .IN2(g6518), .QN(n9057) );
  NAND2X0 U8850 ( .IN1(n9059), .IN2(n9060), .QN(g30263) );
  NAND2X0 U8851 ( .IN1(n4512), .IN2(g261), .QN(n9060) );
  NAND2X0 U8852 ( .IN1(n9038), .IN2(g6313), .QN(n9059) );
  NAND2X0 U8853 ( .IN1(n9061), .IN2(n9062), .QN(g30262) );
  NAND2X0 U8854 ( .IN1(n4369), .IN2(test_so14), .QN(n9062) );
  NAND2X0 U8855 ( .IN1(n9063), .IN2(g165), .QN(n9061) );
  NAND2X0 U8856 ( .IN1(n9064), .IN2(n9065), .QN(g30261) );
  NAND2X0 U8857 ( .IN1(n4318), .IN2(g186), .QN(n9065) );
  NAND2X0 U8858 ( .IN1(n9006), .IN2(g6231), .QN(n9064) );
  NAND2X0 U8859 ( .IN1(n9066), .IN2(n9067), .QN(n9006) );
  NAND2X0 U8860 ( .IN1(n8650), .IN2(n9068), .QN(n9067) );
  XNOR2X1 U8861 ( .IN1(n4513), .IN2(n8799), .Q(n9068) );
  NAND2X0 U8862 ( .IN1(n8653), .IN2(g97), .QN(n9066) );
  NAND2X0 U8863 ( .IN1(n9069), .IN2(n9070), .QN(g30260) );
  NAND2X0 U8864 ( .IN1(n4367), .IN2(g2294), .QN(n9070) );
  NAND2X0 U8865 ( .IN1(n9071), .IN2(g2241), .QN(n9069) );
  NAND2X0 U8866 ( .IN1(n9072), .IN2(n9073), .QN(g30259) );
  NAND2X0 U8867 ( .IN1(n4323), .IN2(g936), .QN(n9073) );
  NAND2X0 U8868 ( .IN1(n9030), .IN2(g6368), .QN(n9072) );
  NAND2X0 U8869 ( .IN1(n9074), .IN2(n9075), .QN(n9030) );
  NAND2X0 U8870 ( .IN1(n9076), .IN2(n8613), .QN(n9075) );
  XNOR2X1 U8871 ( .IN1(n7705), .IN2(n9077), .Q(n9076) );
  NAND2X0 U8872 ( .IN1(n8615), .IN2(g805), .QN(n9074) );
  NAND2X0 U8873 ( .IN1(n9078), .IN2(n9079), .QN(g30258) );
  NAND2X0 U8874 ( .IN1(n4318), .IN2(g258), .QN(n9079) );
  NAND2X0 U8875 ( .IN1(n9038), .IN2(g6231), .QN(n9078) );
  NAND2X0 U8876 ( .IN1(n9080), .IN2(n9081), .QN(n9038) );
  NAND2X0 U8877 ( .IN1(n9082), .IN2(n8650), .QN(n9081) );
  XOR2X1 U8878 ( .IN1(n7673), .IN2(n8808), .Q(n9082) );
  NOR2X0 U8879 ( .IN1(n9083), .IN2(n9084), .QN(n8808) );
  XOR2X1 U8880 ( .IN1(n7672), .IN2(n8346), .Q(n9084) );
  NAND2X0 U8881 ( .IN1(n8653), .IN2(g125), .QN(n9080) );
  NAND2X0 U8882 ( .IN1(n9085), .IN2(n9086), .QN(g30257) );
  NAND2X0 U8883 ( .IN1(n4512), .IN2(g252), .QN(n9086) );
  NAND2X0 U8884 ( .IN1(n9063), .IN2(g6313), .QN(n9085) );
  NAND2X0 U8885 ( .IN1(n9087), .IN2(n9088), .QN(g30256) );
  NAND2X0 U8886 ( .IN1(g2291), .IN2(n7266), .QN(n9088) );
  NAND2X0 U8887 ( .IN1(test_so73), .IN2(n9071), .QN(n9087) );
  NAND2X0 U8888 ( .IN1(n9089), .IN2(n9090), .QN(g30255) );
  NAND2X0 U8889 ( .IN1(n4368), .IN2(g1600), .QN(n9090) );
  NAND2X0 U8890 ( .IN1(n9091), .IN2(g1547), .QN(n9089) );
  NAND2X0 U8891 ( .IN1(n9092), .IN2(n9093), .QN(g30254) );
  NAND2X0 U8892 ( .IN1(n4318), .IN2(g249), .QN(n9093) );
  NAND2X0 U8893 ( .IN1(n9063), .IN2(g6231), .QN(n9092) );
  NAND2X0 U8894 ( .IN1(n9094), .IN2(n9095), .QN(n9063) );
  NAND2X0 U8895 ( .IN1(n9096), .IN2(n8650), .QN(n9095) );
  XOR2X1 U8896 ( .IN1(n9097), .IN2(n9098), .Q(n9096) );
  NAND2X0 U8897 ( .IN1(n9099), .IN2(n9100), .QN(n9097) );
  NAND2X0 U8898 ( .IN1(n8796), .IN2(n7684), .QN(n9100) );
  NAND2X0 U8899 ( .IN1(n8653), .IN2(g117), .QN(n9094) );
  NAND2X0 U8900 ( .IN1(n9101), .IN2(n9102), .QN(g30253) );
  NAND2X0 U8901 ( .IN1(n4324), .IN2(g2288), .QN(n9102) );
  NAND2X0 U8902 ( .IN1(n9071), .IN2(g6837), .QN(n9101) );
  NAND2X0 U8903 ( .IN1(n9103), .IN2(n9104), .QN(n9071) );
  NAND2X0 U8904 ( .IN1(n9105), .IN2(n8557), .QN(n9104) );
  XOR2X1 U8905 ( .IN1(n7763), .IN2(n8979), .Q(n9105) );
  AND3X1 U8906 ( .IN1(n9106), .IN2(n9107), .IN3(n9108), .Q(n8979) );
  INVX0 U8907 ( .INP(n9014), .ZN(n9108) );
  NAND2X0 U8908 ( .IN1(n8916), .IN2(n9109), .QN(n9014) );
  NAND2X0 U8909 ( .IN1(n8349), .IN2(n7771), .QN(n9109) );
  AND3X1 U8910 ( .IN1(n9110), .IN2(n8661), .IN3(n8558), .Q(n8916) );
  AND2X1 U8911 ( .IN1(n8688), .IN2(n9111), .Q(n8558) );
  XOR2X1 U8912 ( .IN1(n8349), .IN2(n9112), .Q(n9111) );
  AND2X1 U8913 ( .IN1(n9113), .IN2(n8955), .Q(n8688) );
  XOR2X1 U8914 ( .IN1(n7765), .IN2(n4529), .Q(n9113) );
  XOR2X1 U8915 ( .IN1(n8349), .IN2(n7769), .Q(n8661) );
  XOR2X1 U8916 ( .IN1(n8349), .IN2(n7757), .Q(n9110) );
  NAND2X0 U8917 ( .IN1(n9114), .IN2(n7758), .QN(n9107) );
  INVX0 U8918 ( .INP(n7771), .ZN(n9114) );
  NAND2X0 U8919 ( .IN1(n4529), .IN2(n9115), .QN(n9106) );
  INVX0 U8920 ( .INP(n8349), .ZN(n4529) );
  NAND2X0 U8921 ( .IN1(n8559), .IN2(g2195), .QN(n9103) );
  NOR2X0 U8922 ( .IN1(n8686), .IN2(n8557), .QN(n8559) );
  AND4X1 U8923 ( .IN1(n9116), .IN2(n9117), .IN3(n9118), .IN4(n8814), .Q(n8557)
         );
  NAND2X0 U8924 ( .IN1(n8824), .IN2(n9119), .QN(n9118) );
  NAND2X0 U8925 ( .IN1(n9120), .IN2(n8840), .QN(n9119) );
  NAND3X0 U8926 ( .IN1(n8829), .IN2(n8837), .IN3(n8889), .QN(n9120) );
  INVX0 U8927 ( .INP(n2792), .ZN(n8837) );
  NAND2X0 U8928 ( .IN1(n9121), .IN2(n9122), .QN(n2792) );
  NAND2X0 U8929 ( .IN1(n9123), .IN2(n9124), .QN(n9117) );
  NAND2X0 U8930 ( .IN1(n4529), .IN2(n9125), .QN(n9124) );
  NAND2X0 U8931 ( .IN1(n9122), .IN2(n9126), .QN(n9116) );
  INVX0 U8932 ( .INP(n3036), .ZN(n9126) );
  NAND2X0 U8933 ( .IN1(n9127), .IN2(n9121), .QN(n3036) );
  NAND3X0 U8934 ( .IN1(n9128), .IN2(n9129), .IN3(n9130), .QN(n9122) );
  NAND2X0 U8935 ( .IN1(n6585), .IN2(n8449), .QN(n9130) );
  NAND2X0 U8936 ( .IN1(n6588), .IN2(n8841), .QN(n9129) );
  NAND2X0 U8937 ( .IN1(n6589), .IN2(n8456), .QN(n9128) );
  INVX0 U8938 ( .INP(n8977), .ZN(n8686) );
  NAND2X0 U8939 ( .IN1(n9123), .IN2(n8814), .QN(n8977) );
  AND2X1 U8940 ( .IN1(n8955), .IN2(n9131), .Q(n9123) );
  NAND2X0 U8941 ( .IN1(n9125), .IN2(n7748), .QN(n9131) );
  NAND4X0 U8942 ( .IN1(n8659), .IN2(n7759), .IN3(n9132), .IN4(n9133), .QN(
        n7748) );
  NOR3X0 U8943 ( .IN1(n7769), .IN2(n9112), .IN3(n7770), .QN(n9133) );
  NAND4X0 U8944 ( .IN1(n9132), .IN2(n7769), .IN3(n4529), .IN4(n9134), .QN(
        n9125) );
  NOR4X0 U8945 ( .IN1(n7759), .IN2(n8659), .IN3(n7774), .IN4(n9135), .QN(n9134) );
  INVX0 U8946 ( .INP(n7770), .ZN(n9135) );
  INVX0 U8947 ( .INP(n9112), .ZN(n7774) );
  INVX0 U8948 ( .INP(n7757), .ZN(n8659) );
  AND4X1 U8949 ( .IN1(n9115), .IN2(n9136), .IN3(n9137), .IN4(n7765), .Q(n9132)
         );
  NOR2X0 U8950 ( .IN1(n7771), .IN2(n7764), .QN(n9137) );
  INVX0 U8951 ( .INP(n7758), .ZN(n9115) );
  NAND2X0 U8952 ( .IN1(n7749), .IN2(n8349), .QN(n8955) );
  NAND2X0 U8953 ( .IN1(n9138), .IN2(n9139), .QN(g30252) );
  NAND2X0 U8954 ( .IN1(n4515), .IN2(g1597), .QN(n9139) );
  NAND2X0 U8955 ( .IN1(n9091), .IN2(g6782), .QN(n9138) );
  NAND2X0 U8956 ( .IN1(n9140), .IN2(n9141), .QN(g30251) );
  NAND2X0 U8957 ( .IN1(g906), .IN2(n7267), .QN(n9141) );
  NAND2X0 U8958 ( .IN1(test_so31), .IN2(n9142), .QN(n9140) );
  NAND2X0 U8959 ( .IN1(n9143), .IN2(n9144), .QN(g30250) );
  NAND2X0 U8960 ( .IN1(n4317), .IN2(g1594), .QN(n9144) );
  NAND2X0 U8961 ( .IN1(n9091), .IN2(g6573), .QN(n9143) );
  NAND2X0 U8962 ( .IN1(n9145), .IN2(n9146), .QN(n9091) );
  NAND2X0 U8963 ( .IN1(n9147), .IN2(n8583), .QN(n9146) );
  XOR2X1 U8964 ( .IN1(n9021), .IN2(n7730), .Q(n9147) );
  NAND3X0 U8965 ( .IN1(n9148), .IN2(n9149), .IN3(n9047), .QN(n9021) );
  NOR2X0 U8966 ( .IN1(n8935), .IN2(n9150), .QN(n9047) );
  NOR2X0 U8967 ( .IN1(n8936), .IN2(n4530), .QN(n9150) );
  NAND3X0 U8968 ( .IN1(n9151), .IN2(n8697), .IN3(n8585), .QN(n8935) );
  AND3X1 U8969 ( .IN1(n9152), .IN2(n8727), .IN3(n8728), .Q(n8585) );
  XOR2X1 U8970 ( .IN1(n8347), .IN2(n7743), .Q(n8728) );
  XOR2X1 U8971 ( .IN1(n8347), .IN2(n9153), .Q(n9152) );
  XOR2X1 U8972 ( .IN1(n4530), .IN2(n7742), .Q(n8697) );
  INVX0 U8973 ( .INP(n8347), .ZN(n4530) );
  XOR2X1 U8974 ( .IN1(n8347), .IN2(n7733), .Q(n9151) );
  NAND2X0 U8975 ( .IN1(n8936), .IN2(n7734), .QN(n9149) );
  OR2X1 U8976 ( .IN1(n8347), .IN2(n7734), .Q(n9148) );
  NAND2X0 U8977 ( .IN1(n8586), .IN2(g1501), .QN(n9145) );
  NOR2X0 U8978 ( .IN1(n8724), .IN2(n8583), .QN(n8586) );
  AND4X1 U8979 ( .IN1(n9154), .IN2(n9155), .IN3(n9156), .IN4(n8465), .Q(n8583)
         );
  NAND2X0 U8980 ( .IN1(n8475), .IN2(n9157), .QN(n9156) );
  NAND2X0 U8981 ( .IN1(n9158), .IN2(n8493), .QN(n9157) );
  NAND4X0 U8982 ( .IN1(n8902), .IN2(n8489), .IN3(n8480), .IN4(n8488), .QN(
        n9158) );
  NAND2X0 U8983 ( .IN1(n9159), .IN2(n9160), .QN(n9155) );
  NAND2X0 U8984 ( .IN1(n4530), .IN2(n9161), .QN(n9160) );
  NAND2X0 U8985 ( .IN1(n8488), .IN2(n9162), .QN(n9154) );
  INVX0 U8986 ( .INP(n3068), .ZN(n9162) );
  NAND2X0 U8987 ( .IN1(n9163), .IN2(n8489), .QN(n3068) );
  NAND3X0 U8988 ( .IN1(n9164), .IN2(n9165), .IN3(n9166), .QN(n8488) );
  NAND2X0 U8989 ( .IN1(n6586), .IN2(n8459), .QN(n9166) );
  NAND2X0 U8990 ( .IN1(n6590), .IN2(n8453), .QN(n9165) );
  NAND2X0 U8991 ( .IN1(n6591), .IN2(n8494), .QN(n9164) );
  INVX0 U8992 ( .INP(n9019), .ZN(n8724) );
  NAND2X0 U8993 ( .IN1(n9159), .IN2(n8465), .QN(n9019) );
  AND2X1 U8994 ( .IN1(n8727), .IN2(n9167), .Q(n9159) );
  NAND2X0 U8995 ( .IN1(n9161), .IN2(n7719), .QN(n9167) );
  NAND4X0 U8996 ( .IN1(n9168), .IN2(n7735), .IN3(n9169), .IN4(n9170), .QN(
        n7719) );
  AND3X1 U8997 ( .IN1(n7744), .IN2(n7742), .IN3(n7732), .Q(n9170) );
  NAND4X0 U8998 ( .IN1(n9169), .IN2(n8584), .IN3(n4530), .IN4(n9171), .QN(
        n9161) );
  NOR4X0 U8999 ( .IN1(n7735), .IN2(n9168), .IN3(n7732), .IN4(n7744), .QN(n9171) );
  INVX0 U9000 ( .INP(n7733), .ZN(n9168) );
  NOR4X0 U9001 ( .IN1(n7734), .IN2(n9023), .IN3(n9172), .IN4(n7731), .QN(n9169) );
  OR2X1 U9002 ( .IN1(n7745), .IN2(n7743), .Q(n9172) );
  NAND2X0 U9003 ( .IN1(n7720), .IN2(n8347), .QN(n8727) );
  NAND2X0 U9004 ( .IN1(n9173), .IN2(n9174), .QN(g30249) );
  NAND2X0 U9005 ( .IN1(n4312), .IN2(g903), .QN(n9174) );
  NAND2X0 U9006 ( .IN1(n9142), .IN2(g6518), .QN(n9173) );
  NAND2X0 U9007 ( .IN1(n9175), .IN2(n9176), .QN(g30248) );
  NAND2X0 U9008 ( .IN1(n4369), .IN2(g219), .QN(n9176) );
  NAND2X0 U9009 ( .IN1(n9177), .IN2(g165), .QN(n9175) );
  NAND2X0 U9010 ( .IN1(n9178), .IN2(n9179), .QN(g30247) );
  NAND2X0 U9011 ( .IN1(n4323), .IN2(g900), .QN(n9179) );
  NAND2X0 U9012 ( .IN1(n9142), .IN2(g6368), .QN(n9178) );
  NAND2X0 U9013 ( .IN1(n9180), .IN2(n9181), .QN(n9142) );
  NAND2X0 U9014 ( .IN1(n9182), .IN2(n8613), .QN(n9181) );
  XOR2X1 U9015 ( .IN1(n9054), .IN2(n9056), .Q(n9182) );
  NAND2X0 U9016 ( .IN1(n9077), .IN2(n9183), .QN(n9054) );
  XOR2X1 U9017 ( .IN1(n7705), .IN2(n8762), .Q(n9183) );
  NOR2X0 U9018 ( .IN1(n8966), .IN2(n9184), .QN(n9077) );
  XOR2X1 U9019 ( .IN1(n8967), .IN2(n8640), .Q(n9184) );
  NAND3X0 U9020 ( .IN1(n8737), .IN2(n9185), .IN3(n8614), .QN(n8966) );
  AND3X1 U9021 ( .IN1(n9186), .IN2(n8766), .IN3(n8767), .Q(n8614) );
  XOR2X1 U9022 ( .IN1(n8640), .IN2(n7711), .Q(n8767) );
  XOR2X1 U9023 ( .IN1(n7712), .IN2(n8640), .Q(n9186) );
  XOR2X1 U9024 ( .IN1(n7713), .IN2(n8640), .Q(n9185) );
  XOR2X1 U9025 ( .IN1(n8762), .IN2(n7699), .Q(n8737) );
  NAND2X0 U9026 ( .IN1(n8615), .IN2(g809), .QN(n9180) );
  NOR2X0 U9027 ( .IN1(n8761), .IN2(n8613), .QN(n8615) );
  AND2X1 U9028 ( .IN1(n9187), .IN2(n9188), .Q(n8613) );
  NAND3X0 U9029 ( .IN1(n9189), .IN2(n8766), .IN3(n9190), .QN(n9188) );
  NAND2X0 U9030 ( .IN1(n8762), .IN2(n9191), .QN(n9190) );
  AND3X1 U9031 ( .IN1(n9189), .IN2(n8766), .IN3(n9187), .Q(n8761) );
  AND3X1 U9032 ( .IN1(n9192), .IN2(n7651), .IN3(n9193), .Q(n9187) );
  NAND2X0 U9033 ( .IN1(n9194), .IN2(n8374), .QN(n9193) );
  NAND2X0 U9034 ( .IN1(n8338), .IN2(n9195), .QN(n9192) );
  NAND2X0 U9035 ( .IN1(n9196), .IN2(n8371), .QN(n9195) );
  NAND3X0 U9036 ( .IN1(n8342), .IN2(n8374), .IN3(n8341), .QN(n9196) );
  INVX0 U9037 ( .INP(n2632), .ZN(n8374) );
  NAND2X0 U9038 ( .IN1(n9197), .IN2(n9198), .QN(n2632) );
  NAND3X0 U9039 ( .IN1(n9199), .IN2(n9200), .IN3(n9201), .QN(n9198) );
  NAND2X0 U9040 ( .IN1(n6592), .IN2(g1088), .QN(n9201) );
  NAND2X0 U9041 ( .IN1(n6593), .IN2(g5472), .QN(n9200) );
  NAND2X0 U9042 ( .IN1(n6587), .IN2(g6712), .QN(n9199) );
  NAND2X0 U9043 ( .IN1(n7691), .IN2(n8640), .QN(n8766) );
  NAND2X0 U9044 ( .IN1(n9191), .IN2(n7690), .QN(n9189) );
  NAND4X0 U9045 ( .IN1(n7699), .IN2(n8636), .IN3(n9202), .IN4(n9203), .QN(
        n7690) );
  NOR3X0 U9046 ( .IN1(n7700), .IN2(n7712), .IN3(n7713), .QN(n9203) );
  NAND4X0 U9047 ( .IN1(n9202), .IN2(n7713), .IN3(n8762), .IN4(n9204), .QN(
        n9191) );
  NOR4X0 U9048 ( .IN1(n8641), .IN2(n8636), .IN3(n7699), .IN4(n8764), .QN(n9204) );
  INVX0 U9049 ( .INP(n7712), .ZN(n8764) );
  INVX0 U9050 ( .INP(n7701), .ZN(n8636) );
  INVX0 U9051 ( .INP(n7700), .ZN(n8641) );
  INVX0 U9052 ( .INP(n8640), .ZN(n8762) );
  AND4X1 U9053 ( .IN1(n7705), .IN2(n9056), .IN3(n9205), .IN4(n8967), .Q(n9202)
         );
  INVX0 U9054 ( .INP(n7706), .ZN(n8967) );
  NOR2X0 U9055 ( .IN1(n7716), .IN2(n7711), .QN(n9205) );
  NAND2X0 U9056 ( .IN1(n9206), .IN2(n9207), .QN(g30246) );
  NAND2X0 U9057 ( .IN1(n4512), .IN2(g216), .QN(n9207) );
  NAND2X0 U9058 ( .IN1(n9177), .IN2(g6313), .QN(n9206) );
  NAND2X0 U9059 ( .IN1(n9208), .IN2(n9209), .QN(g30245) );
  NAND2X0 U9060 ( .IN1(n4318), .IN2(g213), .QN(n9209) );
  NAND2X0 U9061 ( .IN1(n9177), .IN2(g6231), .QN(n9208) );
  NAND2X0 U9062 ( .IN1(n9210), .IN2(n9211), .QN(n9177) );
  NAND2X0 U9063 ( .IN1(n9212), .IN2(n8650), .QN(n9211) );
  XOR2X1 U9064 ( .IN1(n9083), .IN2(n7672), .Q(n9212) );
  NAND3X0 U9065 ( .IN1(n9213), .IN2(n9214), .IN3(n9099), .QN(n9083) );
  NOR2X0 U9066 ( .IN1(n9003), .IN2(n9215), .QN(n9099) );
  NOR2X0 U9067 ( .IN1(n8796), .IN2(n7684), .QN(n9215) );
  NAND3X0 U9068 ( .IN1(n9216), .IN2(n8777), .IN3(n8652), .QN(n9003) );
  AND3X1 U9069 ( .IN1(n9217), .IN2(n8799), .IN3(n8800), .Q(n8652) );
  XNOR2X1 U9070 ( .IN1(n8346), .IN2(n4513), .Q(n8800) );
  AND3X1 U9071 ( .IN1(n9218), .IN2(n9219), .IN3(n9220), .Q(n4513) );
  NAND2X0 U9072 ( .IN1(g186), .IN2(g6231), .QN(n9220) );
  NAND2X0 U9073 ( .IN1(test_so13), .IN2(g6313), .QN(n9219) );
  NAND2X0 U9074 ( .IN1(g192), .IN2(g165), .QN(n9218) );
  XOR2X1 U9075 ( .IN1(n9221), .IN2(n8346), .Q(n9217) );
  XOR2X1 U9076 ( .IN1(n8796), .IN2(n7686), .Q(n8777) );
  XOR2X1 U9077 ( .IN1(n8775), .IN2(n8346), .Q(n9216) );
  NAND2X0 U9078 ( .IN1(n7684), .IN2(n7675), .QN(n9214) );
  NAND2X0 U9079 ( .IN1(n8796), .IN2(n9098), .QN(n9213) );
  NAND2X0 U9080 ( .IN1(n8653), .IN2(g121), .QN(n9210) );
  NOR2X0 U9081 ( .IN1(n8795), .IN2(n8650), .QN(n8653) );
  AND2X1 U9082 ( .IN1(n9222), .IN2(n9223), .Q(n8650) );
  NAND3X0 U9083 ( .IN1(n9224), .IN2(n8799), .IN3(n9225), .QN(n9223) );
  NAND2X0 U9084 ( .IN1(n8796), .IN2(n9226), .QN(n9225) );
  AND3X1 U9085 ( .IN1(n9224), .IN2(n8799), .IN3(n9222), .Q(n8795) );
  AND3X1 U9086 ( .IN1(n9227), .IN2(n8508), .IN3(n9228), .Q(n9222) );
  NAND2X0 U9087 ( .IN1(n8531), .IN2(n9229), .QN(n9228) );
  INVX0 U9088 ( .INP(n3128), .ZN(n9229) );
  NAND2X0 U9089 ( .IN1(n9230), .IN2(n8532), .QN(n3128) );
  NAND2X0 U9090 ( .IN1(n8518), .IN2(n9231), .QN(n9227) );
  NAND2X0 U9091 ( .IN1(n9232), .IN2(n8536), .QN(n9231) );
  NAND4X0 U9092 ( .IN1(n8874), .IN2(n8532), .IN3(n8523), .IN4(n8531), .QN(
        n9232) );
  NAND3X0 U9093 ( .IN1(n9233), .IN2(n9234), .IN3(n9235), .QN(n8531) );
  NAND2X0 U9094 ( .IN1(n6596), .IN2(n8537), .QN(n9235) );
  NAND2X0 U9095 ( .IN1(n6595), .IN2(n8861), .QN(n9234) );
  NAND2X0 U9096 ( .IN1(n6594), .IN2(n8500), .QN(n9233) );
  NAND2X0 U9097 ( .IN1(n7662), .IN2(n8346), .QN(n8799) );
  NAND2X0 U9098 ( .IN1(n9226), .IN2(n7661), .QN(n9224) );
  NAND4X0 U9099 ( .IN1(n7676), .IN2(n7674), .IN3(n9236), .IN4(n9237), .QN(
        n7661) );
  AND3X1 U9100 ( .IN1(n7685), .IN2(n7687), .IN3(n7686), .Q(n9237) );
  NAND4X0 U9101 ( .IN1(n9236), .IN2(n8651), .IN3(n8796), .IN4(n9238), .QN(
        n9226) );
  NOR4X0 U9102 ( .IN1(n7676), .IN2(n7687), .IN3(n7674), .IN4(n7685), .QN(n9238) );
  INVX0 U9103 ( .INP(n8775), .ZN(n7687) );
  INVX0 U9104 ( .INP(n8346), .ZN(n8796) );
  AND4X1 U9105 ( .IN1(n4513), .IN2(n9098), .IN3(n9239), .IN4(n7672), .Q(n9236)
         );
  NOR2X0 U9106 ( .IN1(n9240), .IN2(n7673), .QN(n9239) );
  NAND2X0 U9107 ( .IN1(n9241), .IN2(n9242), .QN(g30072) );
  NAND2X0 U9108 ( .IN1(g2574), .IN2(n7930), .QN(n9242) );
  NAND2X0 U9109 ( .IN1(n4543), .IN2(n9243), .QN(n9241) );
  NAND2X0 U9110 ( .IN1(n9244), .IN2(n9245), .QN(n9243) );
  NAND2X0 U9111 ( .IN1(n7264), .IN2(n9246), .QN(n9245) );
  NAND2X0 U9112 ( .IN1(n9247), .IN2(n7929), .QN(n9244) );
  INVX0 U9113 ( .INP(g7302), .ZN(n9247) );
  NAND2X0 U9114 ( .IN1(n9248), .IN2(n9249), .QN(g30061) );
  NAND2X0 U9115 ( .IN1(g2580), .IN2(n7926), .QN(n9249) );
  NAND2X0 U9116 ( .IN1(n6766), .IN2(n9250), .QN(n9248) );
  NAND2X0 U9117 ( .IN1(n9251), .IN2(n9252), .QN(n9250) );
  NAND2X0 U9118 ( .IN1(n4370), .IN2(g16437), .QN(n9252) );
  NAND2X0 U9119 ( .IN1(g28990), .IN2(g7390), .QN(n9251) );
  NAND2X0 U9120 ( .IN1(n9253), .IN2(n9254), .QN(g30055) );
  NAND2X0 U9121 ( .IN1(n4487), .IN2(DFF_1378_n1), .QN(n9254) );
  NAND2X0 U9122 ( .IN1(n9255), .IN2(g2374), .QN(n9253) );
  NAND2X0 U9123 ( .IN1(n9256), .IN2(n9257), .QN(n9255) );
  NAND2X0 U9124 ( .IN1(g28903), .IN2(g7264), .QN(n9257) );
  NAND2X0 U9125 ( .IN1(n4524), .IN2(g2380), .QN(n9256) );
  NAND2X0 U9126 ( .IN1(n9258), .IN2(n9259), .QN(g29941) );
  NAND2X0 U9127 ( .IN1(n4494), .IN2(g3105), .QN(n9259) );
  NAND2X0 U9128 ( .IN1(n7264), .IN2(g3109), .QN(n9258) );
  NAND2X0 U9129 ( .IN1(n9260), .IN2(n9261), .QN(g29939) );
  OR2X1 U9130 ( .IN1(g8030), .IN2(n4452), .Q(n9261) );
  NAND2X0 U9131 ( .IN1(n7264), .IN2(g8030), .QN(n9260) );
  NAND2X0 U9132 ( .IN1(n9262), .IN2(n9263), .QN(g29936) );
  OR2X1 U9133 ( .IN1(g8106), .IN2(n4447), .Q(n9263) );
  NAND2X0 U9134 ( .IN1(n7264), .IN2(g8106), .QN(n9262) );
  AND2X1 U9135 ( .IN1(n9264), .IN2(n9265), .Q(n7264) );
  NAND2X0 U9136 ( .IN1(g1880), .IN2(DFF_1099_n1), .QN(n9265) );
  NAND3X0 U9137 ( .IN1(n9266), .IN2(n9267), .IN3(n4545), .QN(n9264) );
  NAND2X0 U9138 ( .IN1(n7265), .IN2(n9268), .QN(n9267) );
  NAND2X0 U9139 ( .IN1(n9269), .IN2(n7971), .QN(n9266) );
  INVX0 U9140 ( .INP(g7052), .ZN(n9269) );
  NAND2X0 U9141 ( .IN1(n9270), .IN2(n9271), .QN(g29623) );
  NAND2X0 U9142 ( .IN1(n9272), .IN2(n4606), .QN(n9271) );
  OR2X1 U9143 ( .IN1(n8841), .IN2(n6544), .Q(n9270) );
  NAND2X0 U9144 ( .IN1(n9273), .IN2(n9274), .QN(g29621) );
  NAND2X0 U9145 ( .IN1(n9272), .IN2(g7264), .QN(n9274) );
  OR2X1 U9146 ( .IN1(n8449), .IN2(n6533), .Q(n9273) );
  NAND2X0 U9147 ( .IN1(n9275), .IN2(n9276), .QN(g29620) );
  NAND2X0 U9148 ( .IN1(n9277), .IN2(n4618), .QN(n9276) );
  OR2X1 U9149 ( .IN1(n8453), .IN2(n6550), .Q(n9275) );
  NAND2X0 U9150 ( .IN1(n9278), .IN2(n9279), .QN(g29618) );
  NAND2X0 U9151 ( .IN1(n9272), .IN2(g5555), .QN(n9279) );
  AND2X1 U9152 ( .IN1(n9280), .IN2(n8814), .Q(n9272) );
  NAND2X0 U9153 ( .IN1(n9121), .IN2(n9281), .QN(n8814) );
  NAND2X0 U9154 ( .IN1(n8349), .IN2(n9282), .QN(n9280) );
  NAND3X0 U9155 ( .IN1(n9283), .IN2(n8824), .IN3(n9284), .QN(n9282) );
  NAND3X0 U9156 ( .IN1(n8819), .IN2(n8815), .IN3(n8825), .QN(n8349) );
  OR2X1 U9157 ( .IN1(n8456), .IN2(n6545), .Q(n9278) );
  NAND2X0 U9158 ( .IN1(n9285), .IN2(n9286), .QN(g29617) );
  NAND2X0 U9159 ( .IN1(n9277), .IN2(g7014), .QN(n9286) );
  OR2X1 U9160 ( .IN1(n8459), .IN2(n6536), .Q(n9285) );
  NAND2X0 U9161 ( .IN1(n9287), .IN2(n9288), .QN(g29616) );
  OR2X1 U9162 ( .IN1(g1088), .IN2(n6555), .Q(n9288) );
  NAND2X0 U9163 ( .IN1(n9289), .IN2(g1088), .QN(n9287) );
  NAND2X0 U9164 ( .IN1(n9290), .IN2(n9291), .QN(g29613) );
  NAND2X0 U9165 ( .IN1(n9277), .IN2(g5511), .QN(n9291) );
  AND2X1 U9166 ( .IN1(n9292), .IN2(n8465), .Q(n9277) );
  NAND2X0 U9167 ( .IN1(n8489), .IN2(n9293), .QN(n8465) );
  NAND2X0 U9168 ( .IN1(n8347), .IN2(n9294), .QN(n9292) );
  NAND3X0 U9169 ( .IN1(n9295), .IN2(n8475), .IN3(n9296), .QN(n9294) );
  NAND3X0 U9170 ( .IN1(n8470), .IN2(n8466), .IN3(n8476), .QN(n8347) );
  OR2X1 U9171 ( .IN1(n8494), .IN2(n6551), .Q(n9290) );
  NAND2X0 U9172 ( .IN1(n9297), .IN2(n9298), .QN(g29612) );
  OR2X1 U9173 ( .IN1(g6712), .IN2(n6539), .Q(n9298) );
  NAND2X0 U9174 ( .IN1(n9289), .IN2(g6712), .QN(n9297) );
  NAND2X0 U9175 ( .IN1(n9299), .IN2(n9300), .QN(g29611) );
  NAND2X0 U9176 ( .IN1(n9301), .IN2(n4640), .QN(n9300) );
  OR2X1 U9177 ( .IN1(n8500), .IN2(n6562), .Q(n9299) );
  NAND2X0 U9178 ( .IN1(n9302), .IN2(n9303), .QN(g29609) );
  OR2X1 U9179 ( .IN1(g5472), .IN2(n6556), .Q(n9303) );
  NAND2X0 U9180 ( .IN1(n9289), .IN2(g5472), .QN(n9302) );
  AND2X1 U9181 ( .IN1(n9304), .IN2(n7651), .Q(n9289) );
  NAND2X0 U9182 ( .IN1(n9197), .IN2(n9305), .QN(n7651) );
  NAND2X0 U9183 ( .IN1(n8640), .IN2(n9306), .QN(n9304) );
  NAND3X0 U9184 ( .IN1(n9307), .IN2(n8338), .IN3(n9308), .QN(n9306) );
  NAND3X0 U9185 ( .IN1(n8357), .IN2(n8340), .IN3(n8332), .QN(n8640) );
  NAND2X0 U9186 ( .IN1(n9309), .IN2(n9310), .QN(g29608) );
  NAND2X0 U9187 ( .IN1(n9301), .IN2(g6447), .QN(n9310) );
  OR2X1 U9188 ( .IN1(n8861), .IN2(n6563), .Q(n9309) );
  NAND2X0 U9189 ( .IN1(n9311), .IN2(n9312), .QN(g29606) );
  NAND2X0 U9190 ( .IN1(n9301), .IN2(g5437), .QN(n9312) );
  AND2X1 U9191 ( .IN1(n9313), .IN2(n8508), .Q(n9301) );
  NAND2X0 U9192 ( .IN1(n8532), .IN2(n9314), .QN(n8508) );
  NAND2X0 U9193 ( .IN1(n8346), .IN2(n9315), .QN(n9313) );
  NAND3X0 U9194 ( .IN1(n9316), .IN2(n8518), .IN3(n9317), .QN(n9315) );
  NAND3X0 U9195 ( .IN1(n8513), .IN2(n8509), .IN3(n8519), .QN(n8346) );
  OR2X1 U9196 ( .IN1(n8537), .IN2(n6564), .Q(n9311) );
  NOR2X0 U9197 ( .IN1(n9318), .IN2(n9319), .QN(g29582) );
  XNOR2X1 U9198 ( .IN1(n6436), .IN2(n2981), .Q(n9319) );
  NOR2X0 U9199 ( .IN1(n9320), .IN2(n9321), .QN(g29581) );
  XNOR2X1 U9200 ( .IN1(n6437), .IN2(n2984), .Q(n9321) );
  NOR2X0 U9201 ( .IN1(n9322), .IN2(n9323), .QN(g29580) );
  XNOR2X1 U9202 ( .IN1(n6438), .IN2(n2987), .Q(n9323) );
  NOR2X0 U9203 ( .IN1(n9324), .IN2(n9325), .QN(g29579) );
  XNOR2X1 U9204 ( .IN1(n6439), .IN2(n2990), .Q(n9325) );
  NOR2X0 U9205 ( .IN1(n9318), .IN2(n9326), .QN(g29357) );
  XNOR2X1 U9206 ( .IN1(n6597), .IN2(n2982), .Q(n9326) );
  NOR2X0 U9207 ( .IN1(n9320), .IN2(n9327), .QN(g29355) );
  XNOR2X1 U9208 ( .IN1(n6598), .IN2(n2985), .Q(n9327) );
  NOR2X0 U9209 ( .IN1(n9322), .IN2(n9328), .QN(g29354) );
  XOR2X1 U9210 ( .IN1(n6599), .IN2(n9329), .Q(n9328) );
  NOR2X0 U9211 ( .IN1(n9324), .IN2(n9330), .QN(g29353) );
  XNOR2X1 U9212 ( .IN1(n6600), .IN2(n2991), .Q(n9330) );
  NAND2X0 U9213 ( .IN1(n9331), .IN2(n9332), .QN(g29226) );
  NAND2X0 U9214 ( .IN1(n9333), .IN2(n4606), .QN(n9332) );
  NAND2X0 U9215 ( .IN1(n4509), .IN2(g2498), .QN(n9331) );
  NAND2X0 U9216 ( .IN1(n9334), .IN2(n9335), .QN(g29221) );
  NAND2X0 U9217 ( .IN1(n9333), .IN2(g7264), .QN(n9335) );
  NAND2X0 U9218 ( .IN1(n4524), .IN2(g2495), .QN(n9334) );
  NAND2X0 U9219 ( .IN1(n9336), .IN2(n9337), .QN(g29218) );
  NAND2X0 U9220 ( .IN1(n9338), .IN2(n4618), .QN(n9337) );
  NAND2X0 U9221 ( .IN1(n4511), .IN2(g1804), .QN(n9336) );
  NAND2X0 U9222 ( .IN1(n9339), .IN2(n9340), .QN(g29213) );
  NAND2X0 U9223 ( .IN1(n9333), .IN2(g5555), .QN(n9340) );
  XOR2X1 U9224 ( .IN1(n9341), .IN2(n9342), .Q(n9333) );
  NAND3X0 U9225 ( .IN1(test_so79), .IN2(n9343), .IN3(n9344), .QN(n9341) );
  XOR2X1 U9226 ( .IN1(n9345), .IN2(n9342), .Q(n9344) );
  NAND2X0 U9227 ( .IN1(n9346), .IN2(n9347), .QN(n9343) );
  INVX0 U9228 ( .INP(n8330), .ZN(n9347) );
  NOR2X0 U9229 ( .IN1(n8840), .IN2(n4285), .QN(n8330) );
  NAND2X0 U9230 ( .IN1(n9348), .IN2(n9349), .QN(n9346) );
  NAND2X0 U9231 ( .IN1(n4516), .IN2(g2492), .QN(n9339) );
  NAND2X0 U9232 ( .IN1(n9350), .IN2(n9351), .QN(g29212) );
  NAND2X0 U9233 ( .IN1(n9338), .IN2(g7014), .QN(n9351) );
  NAND2X0 U9234 ( .IN1(n4525), .IN2(g1801), .QN(n9350) );
  NAND2X0 U9235 ( .IN1(n9352), .IN2(n9353), .QN(g29209) );
  NAND2X0 U9236 ( .IN1(n4381), .IN2(g1110), .QN(n9353) );
  NAND2X0 U9237 ( .IN1(n9354), .IN2(g1088), .QN(n9352) );
  NAND2X0 U9238 ( .IN1(n9355), .IN2(n9356), .QN(g29205) );
  NAND2X0 U9239 ( .IN1(n9338), .IN2(g5511), .QN(n9356) );
  XOR2X1 U9240 ( .IN1(n9357), .IN2(n9358), .Q(n9338) );
  NAND3X0 U9241 ( .IN1(n9359), .IN2(g1690), .IN3(n9360), .QN(n9357) );
  XOR2X1 U9242 ( .IN1(n4284), .IN2(n8325), .Q(n9360) );
  NAND2X0 U9243 ( .IN1(n9361), .IN2(n9362), .QN(n9359) );
  INVX0 U9244 ( .INP(n8327), .ZN(n9362) );
  NOR2X0 U9245 ( .IN1(n8493), .IN2(n4284), .QN(n8327) );
  NAND2X0 U9246 ( .IN1(n9363), .IN2(n9364), .QN(n9361) );
  NAND2X0 U9247 ( .IN1(n4518), .IN2(g1798), .QN(n9355) );
  NAND2X0 U9248 ( .IN1(n9365), .IN2(n9366), .QN(g29204) );
  NAND2X0 U9249 ( .IN1(n4364), .IN2(g1107), .QN(n9366) );
  NAND2X0 U9250 ( .IN1(n9354), .IN2(g6712), .QN(n9365) );
  NAND2X0 U9251 ( .IN1(n9367), .IN2(n9368), .QN(g29201) );
  NAND2X0 U9252 ( .IN1(n9369), .IN2(n4640), .QN(n9368) );
  NAND2X0 U9253 ( .IN1(n4506), .IN2(g423), .QN(n9367) );
  NAND2X0 U9254 ( .IN1(n9370), .IN2(n9371), .QN(g29198) );
  NAND2X0 U9255 ( .IN1(n4363), .IN2(g1104), .QN(n9371) );
  NAND2X0 U9256 ( .IN1(n9354), .IN2(g5472), .QN(n9370) );
  XOR2X1 U9257 ( .IN1(n9372), .IN2(n9373), .Q(n9354) );
  NAND3X0 U9258 ( .IN1(n9374), .IN2(g996), .IN3(n9375), .QN(n9372) );
  XOR2X1 U9259 ( .IN1(n9376), .IN2(n9373), .Q(n9375) );
  NAND2X0 U9260 ( .IN1(n9377), .IN2(n9378), .QN(n9374) );
  INVX0 U9261 ( .INP(n8324), .ZN(n9378) );
  NOR2X0 U9262 ( .IN1(n8371), .IN2(n4283), .QN(n8324) );
  NAND2X0 U9263 ( .IN1(n9379), .IN2(n9380), .QN(n9377) );
  NAND2X0 U9264 ( .IN1(n9381), .IN2(n9382), .QN(g29197) );
  NAND2X0 U9265 ( .IN1(n9369), .IN2(g6447), .QN(n9382) );
  NAND2X0 U9266 ( .IN1(n4499), .IN2(g420), .QN(n9381) );
  NAND2X0 U9267 ( .IN1(n9383), .IN2(n9384), .QN(g29194) );
  NAND2X0 U9268 ( .IN1(n9369), .IN2(g5437), .QN(n9384) );
  XOR2X1 U9269 ( .IN1(n9385), .IN2(n9386), .Q(n9369) );
  NAND3X0 U9270 ( .IN1(n9387), .IN2(g309), .IN3(n9388), .QN(n9385) );
  XOR2X1 U9271 ( .IN1(n4282), .IN2(n8319), .Q(n9388) );
  NAND2X0 U9272 ( .IN1(n9389), .IN2(n9390), .QN(n9387) );
  INVX0 U9273 ( .INP(n8321), .ZN(n9390) );
  NOR2X0 U9274 ( .IN1(n8536), .IN2(n4282), .QN(n8321) );
  NAND2X0 U9275 ( .IN1(n9391), .IN2(n9392), .QN(n9389) );
  NAND2X0 U9276 ( .IN1(n4520), .IN2(g417), .QN(n9383) );
  NAND2X0 U9277 ( .IN1(n9393), .IN2(n9394), .QN(g29187) );
  NAND2X0 U9278 ( .IN1(n9395), .IN2(g2396), .QN(n9394) );
  NAND2X0 U9279 ( .IN1(n9396), .IN2(n8841), .QN(n9395) );
  NAND2X0 U9280 ( .IN1(n9397), .IN2(n8841), .QN(n9393) );
  NAND2X0 U9281 ( .IN1(n9398), .IN2(n9399), .QN(g29185) );
  NAND2X0 U9282 ( .IN1(n9400), .IN2(g2398), .QN(n9399) );
  NAND2X0 U9283 ( .IN1(n9396), .IN2(n8449), .QN(n9400) );
  NAND2X0 U9284 ( .IN1(n9397), .IN2(n8449), .QN(n9398) );
  NAND2X0 U9285 ( .IN1(n9401), .IN2(n9402), .QN(g29184) );
  NAND2X0 U9286 ( .IN1(n9403), .IN2(g1702), .QN(n9402) );
  NAND2X0 U9287 ( .IN1(n9404), .IN2(n8453), .QN(n9403) );
  NAND2X0 U9288 ( .IN1(n9405), .IN2(n8453), .QN(n9401) );
  NAND2X0 U9289 ( .IN1(n9406), .IN2(n9407), .QN(g29182) );
  NAND2X0 U9290 ( .IN1(n9408), .IN2(g2397), .QN(n9407) );
  NAND2X0 U9291 ( .IN1(n9396), .IN2(n8456), .QN(n9408) );
  INVX0 U9292 ( .INP(n9409), .ZN(n9396) );
  NAND2X0 U9293 ( .IN1(n9397), .IN2(n8456), .QN(n9406) );
  AND2X1 U9294 ( .IN1(n9410), .IN2(n9409), .Q(n9397) );
  NAND3X0 U9295 ( .IN1(n9410), .IN2(n9411), .IN3(n9121), .QN(n9409) );
  NAND2X0 U9296 ( .IN1(n9412), .IN2(n9283), .QN(n9411) );
  NAND3X0 U9297 ( .IN1(n8825), .IN2(n8824), .IN3(n8889), .QN(n9412) );
  INVX0 U9298 ( .INP(n9284), .ZN(n8889) );
  NAND2X0 U9299 ( .IN1(n8826), .IN2(n8828), .QN(n9284) );
  NAND2X0 U9300 ( .IN1(n3038), .IN2(n9413), .QN(n8828) );
  NAND3X0 U9301 ( .IN1(n9414), .IN2(n9415), .IN3(n9416), .QN(n9413) );
  NAND3X0 U9302 ( .IN1(n9417), .IN2(n9418), .IN3(n9419), .QN(n9416) );
  NAND2X0 U9303 ( .IN1(n9420), .IN2(n9421), .QN(n9418) );
  NAND2X0 U9304 ( .IN1(n9422), .IN2(n9423), .QN(n9417) );
  NAND3X0 U9305 ( .IN1(n9424), .IN2(n9425), .IN3(n9426), .QN(n9415) );
  NAND2X0 U9306 ( .IN1(n9422), .IN2(n9421), .QN(n9425) );
  NAND2X0 U9307 ( .IN1(n9427), .IN2(n9423), .QN(n9424) );
  NAND3X0 U9308 ( .IN1(n9428), .IN2(n9429), .IN3(n9430), .QN(n9414) );
  NAND2X0 U9309 ( .IN1(n9420), .IN2(n9423), .QN(n9429) );
  NAND2X0 U9310 ( .IN1(n9421), .IN2(n9427), .QN(n9428) );
  NAND2X0 U9311 ( .IN1(n3038), .IN2(n9431), .QN(n8826) );
  NAND3X0 U9312 ( .IN1(n9432), .IN2(n9433), .IN3(n9434), .QN(n9431) );
  NAND3X0 U9313 ( .IN1(n9435), .IN2(n9436), .IN3(n9437), .QN(n9434) );
  NAND2X0 U9314 ( .IN1(n9438), .IN2(n9439), .QN(n9435) );
  NAND3X0 U9315 ( .IN1(n9440), .IN2(n9441), .IN3(n9442), .QN(n9433) );
  NAND2X0 U9316 ( .IN1(n9443), .IN2(n9444), .QN(n9441) );
  NAND2X0 U9317 ( .IN1(n9445), .IN2(n9438), .QN(n9440) );
  NAND3X0 U9318 ( .IN1(n9446), .IN2(n9447), .IN3(n9448), .QN(n9432) );
  NAND2X0 U9319 ( .IN1(n9444), .IN2(n9438), .QN(n9447) );
  INVX0 U9320 ( .INP(n9449), .ZN(n9438) );
  INVX0 U9321 ( .INP(n9437), .ZN(n9444) );
  NAND2X0 U9322 ( .IN1(n9443), .IN2(n9439), .QN(n9446) );
  INVX0 U9323 ( .INP(n9442), .ZN(n9439) );
  NAND2X0 U9324 ( .IN1(n9450), .IN2(n9451), .QN(n9410) );
  NAND3X0 U9325 ( .IN1(n3038), .IN2(n8888), .IN3(n9283), .QN(n9451) );
  NAND4X0 U9326 ( .IN1(n9422), .IN2(n9420), .IN3(n9452), .IN4(n9453), .QN(
        n8888) );
  NOR4X0 U9327 ( .IN1(n9436), .IN2(n9437), .IN3(n9449), .IN4(n9442), .QN(n9453) );
  XNOR2X1 U9328 ( .IN1(n7758), .IN2(n4555), .Q(n9442) );
  NAND3X0 U9329 ( .IN1(n9454), .IN2(n9455), .IN3(n9456), .QN(n7758) );
  NAND2X0 U9330 ( .IN1(test_so77), .IN2(test_so73), .QN(n9456) );
  NAND2X0 U9331 ( .IN1(g6837), .IN2(g2324), .QN(n9455) );
  NAND2X0 U9332 ( .IN1(g2241), .IN2(g2330), .QN(n9454) );
  XNOR2X1 U9333 ( .IN1(n7757), .IN2(n4389), .Q(n9449) );
  NAND3X0 U9334 ( .IN1(n9457), .IN2(n9458), .IN3(n9459), .QN(n7757) );
  NAND2X0 U9335 ( .IN1(test_so73), .IN2(g2318), .QN(n9459) );
  NAND2X0 U9336 ( .IN1(g6837), .IN2(g2315), .QN(n9458) );
  NAND2X0 U9337 ( .IN1(g2241), .IN2(g2321), .QN(n9457) );
  XNOR2X1 U9338 ( .IN1(n9112), .IN2(n4373), .Q(n9437) );
  NAND3X0 U9339 ( .IN1(n9460), .IN2(n9461), .IN3(n9462), .QN(n9112) );
  NAND2X0 U9340 ( .IN1(test_so73), .IN2(g2309), .QN(n9462) );
  NAND2X0 U9341 ( .IN1(g6837), .IN2(g2306), .QN(n9461) );
  NAND2X0 U9342 ( .IN1(g2241), .IN2(g2312), .QN(n9460) );
  NAND2X0 U9343 ( .IN1(n9445), .IN2(n9443), .QN(n9436) );
  XOR2X1 U9344 ( .IN1(n7764), .IN2(n4287), .Q(n9443) );
  NAND3X0 U9345 ( .IN1(n9463), .IN2(n9464), .IN3(n9465), .QN(n7764) );
  NAND2X0 U9346 ( .IN1(test_so73), .IN2(g2336), .QN(n9465) );
  NAND2X0 U9347 ( .IN1(g6837), .IN2(g2333), .QN(n9464) );
  NAND2X0 U9348 ( .IN1(g2241), .IN2(g2339), .QN(n9463) );
  INVX0 U9349 ( .INP(n9448), .ZN(n9445) );
  XOR2X1 U9350 ( .IN1(n7759), .IN2(n8573), .Q(n9448) );
  AND3X1 U9351 ( .IN1(n9466), .IN2(n9467), .IN3(n9468), .Q(n7759) );
  NAND2X0 U9352 ( .IN1(g2348), .IN2(g2241), .QN(n9468) );
  NAND2X0 U9353 ( .IN1(g2342), .IN2(g6837), .QN(n9467) );
  NAND2X0 U9354 ( .IN1(test_so73), .IN2(g2345), .QN(n9466) );
  AND3X1 U9355 ( .IN1(n9421), .IN2(n9423), .IN3(n9427), .Q(n9452) );
  INVX0 U9356 ( .INP(n9419), .ZN(n9427) );
  XOR2X1 U9357 ( .IN1(n7765), .IN2(n4377), .Q(n9419) );
  AND3X1 U9358 ( .IN1(n9469), .IN2(n9470), .IN3(n9471), .Q(n7765) );
  NAND2X0 U9359 ( .IN1(g2261), .IN2(g6837), .QN(n9471) );
  NAND2X0 U9360 ( .IN1(test_so76), .IN2(test_so73), .QN(n9470) );
  NAND2X0 U9361 ( .IN1(g2267), .IN2(g2241), .QN(n9469) );
  XOR2X1 U9362 ( .IN1(n9136), .IN2(g2195), .Q(n9423) );
  INVX0 U9363 ( .INP(n7763), .ZN(n9136) );
  NAND3X0 U9364 ( .IN1(n9472), .IN2(n9473), .IN3(n9474), .QN(n7763) );
  NAND2X0 U9365 ( .IN1(test_so73), .IN2(g2291), .QN(n9474) );
  NAND2X0 U9366 ( .IN1(g6837), .IN2(g2288), .QN(n9473) );
  NAND2X0 U9367 ( .IN1(g2241), .IN2(g2294), .QN(n9472) );
  XOR2X1 U9368 ( .IN1(n9475), .IN2(g2175), .Q(n9421) );
  INVX0 U9369 ( .INP(n7769), .ZN(n9475) );
  NAND3X0 U9370 ( .IN1(n9476), .IN2(n9477), .IN3(n9478), .QN(n7769) );
  NAND2X0 U9371 ( .IN1(test_so73), .IN2(g2273), .QN(n9478) );
  NAND2X0 U9372 ( .IN1(g6837), .IN2(g2270), .QN(n9477) );
  NAND2X0 U9373 ( .IN1(g2241), .IN2(g2276), .QN(n9476) );
  INVX0 U9374 ( .INP(n9426), .ZN(n9420) );
  XNOR2X1 U9375 ( .IN1(n7771), .IN2(n4325), .Q(n9426) );
  NAND3X0 U9376 ( .IN1(n9479), .IN2(n9480), .IN3(n9481), .QN(n7771) );
  NAND2X0 U9377 ( .IN1(g2279), .IN2(g6837), .QN(n9481) );
  NAND2X0 U9378 ( .IN1(g2285), .IN2(g2241), .QN(n9480) );
  NAND2X0 U9379 ( .IN1(test_so73), .IN2(g2282), .QN(n9479) );
  INVX0 U9380 ( .INP(n9430), .ZN(n9422) );
  XNOR2X1 U9381 ( .IN1(n7770), .IN2(n9482), .Q(n9430) );
  NAND3X0 U9382 ( .IN1(n9483), .IN2(n9484), .IN3(n9485), .QN(n7770) );
  NAND2X0 U9383 ( .IN1(test_so73), .IN2(g2300), .QN(n9485) );
  NAND2X0 U9384 ( .IN1(g6837), .IN2(g2297), .QN(n9484) );
  NAND2X0 U9385 ( .IN1(g2241), .IN2(g2303), .QN(n9483) );
  NAND2X0 U9386 ( .IN1(n9127), .IN2(test_so79), .QN(n9450) );
  NAND2X0 U9387 ( .IN1(n9486), .IN2(n9487), .QN(g29181) );
  NAND2X0 U9388 ( .IN1(n9488), .IN2(g1704), .QN(n9487) );
  NAND2X0 U9389 ( .IN1(n9404), .IN2(n8459), .QN(n9488) );
  NAND2X0 U9390 ( .IN1(n9405), .IN2(n8459), .QN(n9486) );
  NAND2X0 U9391 ( .IN1(n9489), .IN2(n9490), .QN(g29179) );
  NAND2X0 U9392 ( .IN1(n9491), .IN2(g1008), .QN(n9490) );
  NAND2X0 U9393 ( .IN1(n9492), .IN2(g1088), .QN(n9491) );
  NAND2X0 U9394 ( .IN1(n9493), .IN2(g1088), .QN(n9489) );
  NAND2X0 U9395 ( .IN1(n9494), .IN2(n9495), .QN(g29178) );
  NAND2X0 U9396 ( .IN1(n9496), .IN2(g1703), .QN(n9495) );
  NAND2X0 U9397 ( .IN1(n9404), .IN2(n8494), .QN(n9496) );
  INVX0 U9398 ( .INP(n9497), .ZN(n9404) );
  NAND2X0 U9399 ( .IN1(n9405), .IN2(n8494), .QN(n9494) );
  AND2X1 U9400 ( .IN1(n9498), .IN2(n9497), .Q(n9405) );
  NAND3X0 U9401 ( .IN1(n9498), .IN2(n9499), .IN3(n8489), .QN(n9497) );
  NAND2X0 U9402 ( .IN1(n9500), .IN2(n9295), .QN(n9499) );
  NAND3X0 U9403 ( .IN1(n8476), .IN2(n8475), .IN3(n8902), .QN(n9500) );
  INVX0 U9404 ( .INP(n9296), .ZN(n8902) );
  NAND2X0 U9405 ( .IN1(n8477), .IN2(n8479), .QN(n9296) );
  NAND2X0 U9406 ( .IN1(n3070), .IN2(n9501), .QN(n8479) );
  NAND3X0 U9407 ( .IN1(n9502), .IN2(n9503), .IN3(n9504), .QN(n9501) );
  NAND3X0 U9408 ( .IN1(n9505), .IN2(n9506), .IN3(n9507), .QN(n9504) );
  NAND2X0 U9409 ( .IN1(n9508), .IN2(n9509), .QN(n9506) );
  NAND2X0 U9410 ( .IN1(n9510), .IN2(n9511), .QN(n9505) );
  NAND3X0 U9411 ( .IN1(n9512), .IN2(n9513), .IN3(n9514), .QN(n9503) );
  NAND2X0 U9412 ( .IN1(n9510), .IN2(n9509), .QN(n9513) );
  INVX0 U9413 ( .INP(n9515), .ZN(n9510) );
  NAND3X0 U9414 ( .IN1(n9516), .IN2(n9517), .IN3(n9515), .QN(n9502) );
  NAND2X0 U9415 ( .IN1(n9508), .IN2(n9511), .QN(n9517) );
  INVX0 U9416 ( .INP(n9514), .ZN(n9508) );
  NAND2X0 U9417 ( .IN1(n9509), .IN2(n9518), .QN(n9516) );
  INVX0 U9418 ( .INP(n9519), .ZN(n9509) );
  NAND2X0 U9419 ( .IN1(n3070), .IN2(n9520), .QN(n8477) );
  NAND3X0 U9420 ( .IN1(n9521), .IN2(n9522), .IN3(n9523), .QN(n9520) );
  NAND3X0 U9421 ( .IN1(n9524), .IN2(n9525), .IN3(n9526), .QN(n9523) );
  NAND2X0 U9422 ( .IN1(n9527), .IN2(n9528), .QN(n9525) );
  NAND2X0 U9423 ( .IN1(n9529), .IN2(n9530), .QN(n9524) );
  NAND3X0 U9424 ( .IN1(n9531), .IN2(n9532), .IN3(n9533), .QN(n9522) );
  NAND2X0 U9425 ( .IN1(n9534), .IN2(n9528), .QN(n9532) );
  NAND2X0 U9426 ( .IN1(n9527), .IN2(n9529), .QN(n9531) );
  NAND3X0 U9427 ( .IN1(n9535), .IN2(n9536), .IN3(n9537), .QN(n9521) );
  NAND2X0 U9428 ( .IN1(n9534), .IN2(n9529), .QN(n9536) );
  NAND2X0 U9429 ( .IN1(n9528), .IN2(n9530), .QN(n9535) );
  NAND2X0 U9430 ( .IN1(n9538), .IN2(n9539), .QN(n9498) );
  NAND2X0 U9431 ( .IN1(n9163), .IN2(g1690), .QN(n9539) );
  NAND3X0 U9432 ( .IN1(n3070), .IN2(n8900), .IN3(n9295), .QN(n9538) );
  NAND4X0 U9433 ( .IN1(n9527), .IN2(n9534), .IN3(n9540), .IN4(n9541), .QN(
        n8900) );
  NOR4X0 U9434 ( .IN1(n9519), .IN2(n9512), .IN3(n9514), .IN4(n9515), .QN(n9541) );
  XNOR2X1 U9435 ( .IN1(n8756), .IN2(n7744), .Q(n9515) );
  INVX0 U9436 ( .INP(n8348), .ZN(n7744) );
  NAND3X0 U9437 ( .IN1(n9542), .IN2(n9543), .IN3(n9544), .QN(n8348) );
  NAND2X0 U9438 ( .IN1(test_so56), .IN2(g6782), .QN(n9544) );
  NAND2X0 U9439 ( .IN1(g6573), .IN2(g1603), .QN(n9543) );
  NAND2X0 U9440 ( .IN1(g1547), .IN2(g1609), .QN(n9542) );
  XNOR2X1 U9441 ( .IN1(g1491), .IN2(n8936), .Q(n9514) );
  INVX0 U9442 ( .INP(n7745), .ZN(n8936) );
  NAND3X0 U9443 ( .IN1(n9545), .IN2(n9546), .IN3(n9547), .QN(n7745) );
  NAND2X0 U9444 ( .IN1(g6782), .IN2(g1588), .QN(n9547) );
  NAND2X0 U9445 ( .IN1(g6573), .IN2(g1585), .QN(n9546) );
  NAND2X0 U9446 ( .IN1(g1547), .IN2(g1591), .QN(n9545) );
  NAND2X0 U9447 ( .IN1(n9518), .IN2(n9511), .QN(n9512) );
  XOR2X1 U9448 ( .IN1(g1501), .IN2(n7730), .Q(n9511) );
  INVX0 U9449 ( .INP(n9023), .ZN(n7730) );
  NAND3X0 U9450 ( .IN1(n9548), .IN2(n9549), .IN3(n9550), .QN(n9023) );
  NAND2X0 U9451 ( .IN1(g6782), .IN2(g1597), .QN(n9550) );
  NAND2X0 U9452 ( .IN1(g6573), .IN2(g1594), .QN(n9549) );
  NAND2X0 U9453 ( .IN1(g1547), .IN2(g1600), .QN(n9548) );
  INVX0 U9454 ( .INP(n9507), .ZN(n9518) );
  XOR2X1 U9455 ( .IN1(g1471), .IN2(n7743), .Q(n9507) );
  NAND3X0 U9456 ( .IN1(n9551), .IN2(n9552), .IN3(n9553), .QN(n7743) );
  NAND2X0 U9457 ( .IN1(g6782), .IN2(g1570), .QN(n9553) );
  NAND2X0 U9458 ( .IN1(g6573), .IN2(g1567), .QN(n9552) );
  NAND2X0 U9459 ( .IN1(g1547), .IN2(g1573), .QN(n9551) );
  XNOR2X1 U9460 ( .IN1(g1481), .IN2(n7742), .Q(n9519) );
  INVX0 U9461 ( .INP(n8584), .ZN(n7742) );
  NAND3X0 U9462 ( .IN1(n9554), .IN2(n9555), .IN3(n9556), .QN(n8584) );
  NAND2X0 U9463 ( .IN1(g6782), .IN2(g1579), .QN(n9556) );
  NAND2X0 U9464 ( .IN1(g6573), .IN2(g1576), .QN(n9555) );
  NAND2X0 U9465 ( .IN1(g1547), .IN2(g1582), .QN(n9554) );
  AND3X1 U9466 ( .IN1(n9528), .IN2(n9529), .IN3(n9530), .Q(n9540) );
  INVX0 U9467 ( .INP(n9533), .ZN(n9530) );
  XOR2X1 U9468 ( .IN1(g1496), .IN2(n7734), .Q(n9533) );
  NAND3X0 U9469 ( .IN1(n9557), .IN2(n9558), .IN3(n9559), .QN(n7734) );
  NAND2X0 U9470 ( .IN1(g6782), .IN2(g1633), .QN(n9559) );
  NAND2X0 U9471 ( .IN1(g6573), .IN2(g1630), .QN(n9558) );
  NAND2X0 U9472 ( .IN1(g1547), .IN2(g1636), .QN(n9557) );
  XOR2X1 U9473 ( .IN1(n4390), .IN2(n7733), .Q(n9529) );
  NAND3X0 U9474 ( .IN1(n9560), .IN2(n9561), .IN3(n9562), .QN(n7733) );
  NAND2X0 U9475 ( .IN1(g6782), .IN2(g1624), .QN(n9562) );
  NAND2X0 U9476 ( .IN1(test_so55), .IN2(g6573), .QN(n9561) );
  NAND2X0 U9477 ( .IN1(g1547), .IN2(g1627), .QN(n9560) );
  XOR2X1 U9478 ( .IN1(n4288), .IN2(n7731), .Q(n9528) );
  NAND3X0 U9479 ( .IN1(n9563), .IN2(n9564), .IN3(n9565), .QN(n7731) );
  NAND2X0 U9480 ( .IN1(g6782), .IN2(g1642), .QN(n9565) );
  NAND2X0 U9481 ( .IN1(g6573), .IN2(g1639), .QN(n9564) );
  NAND2X0 U9482 ( .IN1(g1547), .IN2(g1645), .QN(n9563) );
  INVX0 U9483 ( .INP(n9526), .ZN(n9534) );
  XNOR2X1 U9484 ( .IN1(g1476), .IN2(n7732), .Q(n9526) );
  INVX0 U9485 ( .INP(n9153), .ZN(n7732) );
  NAND3X0 U9486 ( .IN1(n9566), .IN2(n9567), .IN3(n9568), .QN(n9153) );
  NAND2X0 U9487 ( .IN1(g6782), .IN2(g1615), .QN(n9568) );
  NAND2X0 U9488 ( .IN1(g6573), .IN2(g1612), .QN(n9567) );
  NAND2X0 U9489 ( .IN1(g1547), .IN2(g1618), .QN(n9566) );
  INVX0 U9490 ( .INP(n9537), .ZN(n9527) );
  XOR2X1 U9491 ( .IN1(n7735), .IN2(n8603), .Q(n9537) );
  AND3X1 U9492 ( .IN1(n9569), .IN2(n9570), .IN3(n9571), .Q(n7735) );
  NAND2X0 U9493 ( .IN1(g1648), .IN2(g6573), .QN(n9571) );
  NAND2X0 U9494 ( .IN1(g1651), .IN2(g6782), .QN(n9570) );
  NAND2X0 U9495 ( .IN1(g1654), .IN2(g1547), .QN(n9569) );
  NAND2X0 U9496 ( .IN1(n9572), .IN2(n9573), .QN(g29173) );
  NAND2X0 U9497 ( .IN1(n9574), .IN2(g1010), .QN(n9573) );
  NAND2X0 U9498 ( .IN1(n9492), .IN2(g6712), .QN(n9574) );
  NAND2X0 U9499 ( .IN1(n9493), .IN2(g6712), .QN(n9572) );
  NAND2X0 U9500 ( .IN1(n9575), .IN2(n9576), .QN(g29172) );
  NAND2X0 U9501 ( .IN1(n9577), .IN2(g321), .QN(n9576) );
  NAND2X0 U9502 ( .IN1(n9578), .IN2(n8500), .QN(n9577) );
  NAND2X0 U9503 ( .IN1(n9579), .IN2(n8500), .QN(n9575) );
  NAND2X0 U9504 ( .IN1(n9580), .IN2(n9581), .QN(g29170) );
  NAND2X0 U9505 ( .IN1(n9582), .IN2(g1009), .QN(n9581) );
  NAND2X0 U9506 ( .IN1(n9492), .IN2(g5472), .QN(n9582) );
  INVX0 U9507 ( .INP(n3065), .ZN(n9492) );
  NAND2X0 U9508 ( .IN1(n9493), .IN2(g5472), .QN(n9580) );
  AND2X1 U9509 ( .IN1(n9583), .IN2(n3065), .Q(n9493) );
  NAND3X0 U9510 ( .IN1(n9583), .IN2(n9584), .IN3(n9197), .QN(n3065) );
  NAND2X0 U9511 ( .IN1(n9585), .IN2(n9307), .QN(n9584) );
  NAND3X0 U9512 ( .IN1(n8332), .IN2(n8338), .IN3(n8341), .QN(n9585) );
  INVX0 U9513 ( .INP(n9308), .ZN(n8341) );
  NAND2X0 U9514 ( .IN1(n8362), .IN2(n8364), .QN(n9308) );
  NAND2X0 U9515 ( .IN1(n3102), .IN2(n9586), .QN(n8364) );
  NAND3X0 U9516 ( .IN1(n9587), .IN2(n9588), .IN3(n9589), .QN(n9586) );
  NAND3X0 U9517 ( .IN1(n9590), .IN2(n9591), .IN3(n9592), .QN(n9589) );
  INVX0 U9518 ( .INP(n9593), .ZN(n9592) );
  NAND2X0 U9519 ( .IN1(n9594), .IN2(n9595), .QN(n9591) );
  NAND2X0 U9520 ( .IN1(n9596), .IN2(n9597), .QN(n9590) );
  NAND3X0 U9521 ( .IN1(n9598), .IN2(n9599), .IN3(n9600), .QN(n9588) );
  NAND2X0 U9522 ( .IN1(n9593), .IN2(n9595), .QN(n9599) );
  NAND2X0 U9523 ( .IN1(n9594), .IN2(n9597), .QN(n9598) );
  NAND3X0 U9524 ( .IN1(n9601), .IN2(n9602), .IN3(n9603), .QN(n9587) );
  NAND2X0 U9525 ( .IN1(n9597), .IN2(n9593), .QN(n9602) );
  NAND2X0 U9526 ( .IN1(n9596), .IN2(n9595), .QN(n9601) );
  NAND2X0 U9527 ( .IN1(n3102), .IN2(n9604), .QN(n8362) );
  NAND3X0 U9528 ( .IN1(n9605), .IN2(n9606), .IN3(n9607), .QN(n9604) );
  NAND3X0 U9529 ( .IN1(n9608), .IN2(n9609), .IN3(n9610), .QN(n9607) );
  NAND2X0 U9530 ( .IN1(n9611), .IN2(n9612), .QN(n9609) );
  NAND2X0 U9531 ( .IN1(n9613), .IN2(n9614), .QN(n9608) );
  NAND3X0 U9532 ( .IN1(n9615), .IN2(n9616), .IN3(n9617), .QN(n9606) );
  NAND2X0 U9533 ( .IN1(n9612), .IN2(n9614), .QN(n9616) );
  NAND2X0 U9534 ( .IN1(n9618), .IN2(n9613), .QN(n9615) );
  NAND3X0 U9535 ( .IN1(n9619), .IN2(n9620), .IN3(n9621), .QN(n9605) );
  NAND2X0 U9536 ( .IN1(n9618), .IN2(n9612), .QN(n9620) );
  NAND2X0 U9537 ( .IN1(n9611), .IN2(n9613), .QN(n9619) );
  INVX0 U9538 ( .INP(n9617), .ZN(n9611) );
  NAND2X0 U9539 ( .IN1(n9622), .IN2(n9623), .QN(n9583) );
  NAND2X0 U9540 ( .IN1(n9194), .IN2(g996), .QN(n9623) );
  NAND3X0 U9541 ( .IN1(n3102), .IN2(n8363), .IN3(n9307), .QN(n9622) );
  NAND4X0 U9542 ( .IN1(n9596), .IN2(n9594), .IN3(n9624), .IN4(n9625), .QN(
        n8363) );
  AND4X1 U9543 ( .IN1(n9626), .IN2(n9613), .IN3(n9614), .IN4(n9612), .Q(n9625)
         );
  XOR2X1 U9544 ( .IN1(n7713), .IN2(n4391), .Q(n9612) );
  NAND3X0 U9545 ( .IN1(n9627), .IN2(n9628), .IN3(n9629), .QN(n7713) );
  NAND2X0 U9546 ( .IN1(test_so31), .IN2(g933), .QN(n9629) );
  NAND2X0 U9547 ( .IN1(g6518), .IN2(g930), .QN(n9628) );
  NAND2X0 U9548 ( .IN1(g6368), .IN2(g927), .QN(n9627) );
  INVX0 U9549 ( .INP(n9621), .ZN(n9614) );
  XNOR2X1 U9550 ( .IN1(n7701), .IN2(n8634), .Q(n9621) );
  NAND3X0 U9551 ( .IN1(n9630), .IN2(n9631), .IN3(n9632), .QN(n7701) );
  NAND2X0 U9552 ( .IN1(g954), .IN2(g6368), .QN(n9632) );
  NAND2X0 U9553 ( .IN1(g957), .IN2(g6518), .QN(n9631) );
  NAND2X0 U9554 ( .IN1(test_so31), .IN2(g960), .QN(n9630) );
  XOR2X1 U9555 ( .IN1(n7716), .IN2(n4289), .Q(n9613) );
  NAND3X0 U9556 ( .IN1(n9633), .IN2(n9634), .IN3(n9635), .QN(n7716) );
  NAND2X0 U9557 ( .IN1(test_so31), .IN2(g951), .QN(n9635) );
  NAND2X0 U9558 ( .IN1(g6518), .IN2(g948), .QN(n9634) );
  NAND2X0 U9559 ( .IN1(test_so35), .IN2(g6368), .QN(n9633) );
  NOR2X0 U9560 ( .IN1(n9617), .IN2(n9610), .QN(n9626) );
  INVX0 U9561 ( .INP(n9618), .ZN(n9610) );
  XOR2X1 U9562 ( .IN1(n7712), .IN2(n4375), .Q(n9618) );
  NAND3X0 U9563 ( .IN1(n9636), .IN2(n9637), .IN3(n9638), .QN(n7712) );
  NAND2X0 U9564 ( .IN1(test_so34), .IN2(test_so31), .QN(n9638) );
  NAND2X0 U9565 ( .IN1(g6518), .IN2(g921), .QN(n9637) );
  NAND2X0 U9566 ( .IN1(g6368), .IN2(g918), .QN(n9636) );
  XOR2X1 U9567 ( .IN1(n7705), .IN2(n4559), .Q(n9617) );
  AND3X1 U9568 ( .IN1(n9639), .IN2(n9640), .IN3(n9641), .Q(n7705) );
  NAND2X0 U9569 ( .IN1(test_so31), .IN2(g942), .QN(n9641) );
  NAND2X0 U9570 ( .IN1(g6518), .IN2(g939), .QN(n9640) );
  NAND2X0 U9571 ( .IN1(g6368), .IN2(g936), .QN(n9639) );
  AND3X1 U9572 ( .IN1(n9597), .IN2(n9595), .IN3(n9593), .Q(n9624) );
  XOR2X1 U9573 ( .IN1(n7711), .IN2(n4379), .Q(n9593) );
  NAND3X0 U9574 ( .IN1(n9642), .IN2(n9643), .IN3(n9644), .QN(n7711) );
  NAND2X0 U9575 ( .IN1(test_so31), .IN2(g879), .QN(n9644) );
  NAND2X0 U9576 ( .IN1(g6518), .IN2(g876), .QN(n9643) );
  NAND2X0 U9577 ( .IN1(g6368), .IN2(g873), .QN(n9642) );
  XOR2X1 U9578 ( .IN1(n9056), .IN2(g809), .Q(n9595) );
  INVX0 U9579 ( .INP(n7707), .ZN(n9056) );
  NAND3X0 U9580 ( .IN1(n9645), .IN2(n9646), .IN3(n9647), .QN(n7707) );
  NAND2X0 U9581 ( .IN1(test_so31), .IN2(g906), .QN(n9647) );
  NAND2X0 U9582 ( .IN1(g6518), .IN2(g903), .QN(n9646) );
  NAND2X0 U9583 ( .IN1(g6368), .IN2(g900), .QN(n9645) );
  XOR2X1 U9584 ( .IN1(n7699), .IN2(g793), .Q(n9597) );
  AND3X1 U9585 ( .IN1(n9648), .IN2(n9649), .IN3(n9650), .Q(n7699) );
  NAND2X0 U9586 ( .IN1(test_so31), .IN2(g888), .QN(n9650) );
  NAND2X0 U9587 ( .IN1(g6518), .IN2(g885), .QN(n9649) );
  NAND2X0 U9588 ( .IN1(g6368), .IN2(g882), .QN(n9648) );
  INVX0 U9589 ( .INP(n9603), .ZN(n9594) );
  XNOR2X1 U9590 ( .IN1(n7700), .IN2(n9651), .Q(n9603) );
  NAND3X0 U9591 ( .IN1(n9652), .IN2(n9653), .IN3(n9654), .QN(n7700) );
  NAND2X0 U9592 ( .IN1(g909), .IN2(g6368), .QN(n9654) );
  NAND2X0 U9593 ( .IN1(g912), .IN2(g6518), .QN(n9653) );
  NAND2X0 U9594 ( .IN1(test_so31), .IN2(g915), .QN(n9652) );
  INVX0 U9595 ( .INP(n9600), .ZN(n9596) );
  XNOR2X1 U9596 ( .IN1(n7706), .IN2(n4327), .Q(n9600) );
  NAND3X0 U9597 ( .IN1(n9655), .IN2(n9656), .IN3(n9657), .QN(n7706) );
  NAND2X0 U9598 ( .IN1(test_so31), .IN2(g897), .QN(n9657) );
  NAND2X0 U9599 ( .IN1(g6518), .IN2(g894), .QN(n9656) );
  NAND2X0 U9600 ( .IN1(g6368), .IN2(g891), .QN(n9655) );
  NAND2X0 U9601 ( .IN1(n9658), .IN2(n9659), .QN(g29169) );
  NAND2X0 U9602 ( .IN1(n9660), .IN2(g323), .QN(n9659) );
  NAND2X0 U9603 ( .IN1(n9578), .IN2(n8861), .QN(n9660) );
  NAND2X0 U9604 ( .IN1(n9579), .IN2(n8861), .QN(n9658) );
  NAND2X0 U9605 ( .IN1(n9661), .IN2(n9662), .QN(g29167) );
  NAND2X0 U9606 ( .IN1(n9663), .IN2(g322), .QN(n9662) );
  NAND2X0 U9607 ( .IN1(n9578), .IN2(n8537), .QN(n9663) );
  INVX0 U9608 ( .INP(n9664), .ZN(n9578) );
  NAND2X0 U9609 ( .IN1(n9579), .IN2(n8537), .QN(n9661) );
  AND2X1 U9610 ( .IN1(n9665), .IN2(n9664), .Q(n9579) );
  NAND3X0 U9611 ( .IN1(n9665), .IN2(n9666), .IN3(n8532), .QN(n9664) );
  NAND2X0 U9612 ( .IN1(n9667), .IN2(n9316), .QN(n9666) );
  NAND3X0 U9613 ( .IN1(n8519), .IN2(n8518), .IN3(n8874), .QN(n9667) );
  INVX0 U9614 ( .INP(n9317), .ZN(n8874) );
  NAND2X0 U9615 ( .IN1(n8520), .IN2(n8522), .QN(n9317) );
  NAND2X0 U9616 ( .IN1(n3130), .IN2(n9668), .QN(n8522) );
  NAND3X0 U9617 ( .IN1(n9669), .IN2(n9670), .IN3(n9671), .QN(n9668) );
  NAND3X0 U9618 ( .IN1(n9672), .IN2(n9673), .IN3(n9674), .QN(n9671) );
  NAND2X0 U9619 ( .IN1(n9675), .IN2(n9676), .QN(n9673) );
  NAND2X0 U9620 ( .IN1(n9677), .IN2(n9678), .QN(n9672) );
  NAND3X0 U9621 ( .IN1(n9679), .IN2(n9680), .IN3(n9681), .QN(n9670) );
  NAND2X0 U9622 ( .IN1(n9677), .IN2(n9676), .QN(n9680) );
  INVX0 U9623 ( .INP(n9682), .ZN(n9677) );
  NAND3X0 U9624 ( .IN1(n9683), .IN2(n9684), .IN3(n9682), .QN(n9669) );
  NAND2X0 U9625 ( .IN1(n9675), .IN2(n9678), .QN(n9684) );
  INVX0 U9626 ( .INP(n9681), .ZN(n9675) );
  NAND2X0 U9627 ( .IN1(n9676), .IN2(n9685), .QN(n9683) );
  INVX0 U9628 ( .INP(n9686), .ZN(n9676) );
  NAND2X0 U9629 ( .IN1(n3130), .IN2(n9687), .QN(n8520) );
  NAND3X0 U9630 ( .IN1(n9688), .IN2(n9689), .IN3(n9690), .QN(n9687) );
  NAND3X0 U9631 ( .IN1(n9691), .IN2(n9692), .IN3(n9693), .QN(n9690) );
  NAND2X0 U9632 ( .IN1(n9694), .IN2(n9695), .QN(n9692) );
  NAND2X0 U9633 ( .IN1(n9696), .IN2(n9697), .QN(n9691) );
  NAND3X0 U9634 ( .IN1(n9698), .IN2(n9699), .IN3(n9700), .QN(n9689) );
  NAND2X0 U9635 ( .IN1(n9701), .IN2(n9695), .QN(n9699) );
  NAND2X0 U9636 ( .IN1(n9694), .IN2(n9696), .QN(n9698) );
  NAND3X0 U9637 ( .IN1(n9702), .IN2(n9703), .IN3(n9704), .QN(n9688) );
  NAND2X0 U9638 ( .IN1(n9701), .IN2(n9696), .QN(n9703) );
  NAND2X0 U9639 ( .IN1(n9695), .IN2(n9697), .QN(n9702) );
  NAND2X0 U9640 ( .IN1(n9705), .IN2(n9706), .QN(n9665) );
  NAND2X0 U9641 ( .IN1(n9230), .IN2(g309), .QN(n9706) );
  NAND3X0 U9642 ( .IN1(n3130), .IN2(n8872), .IN3(n9316), .QN(n9705) );
  NAND4X0 U9643 ( .IN1(n9694), .IN2(n9701), .IN3(n9707), .IN4(n9708), .QN(
        n8872) );
  NOR4X0 U9644 ( .IN1(n9686), .IN2(n9679), .IN3(n9681), .IN4(n9682), .QN(n9708) );
  XNOR2X1 U9645 ( .IN1(n8810), .IN2(n7685), .Q(n9682) );
  INVX0 U9646 ( .INP(n8345), .ZN(n7685) );
  NAND3X0 U9647 ( .IN1(n9709), .IN2(n9710), .IN3(n9711), .QN(n8345) );
  NAND2X0 U9648 ( .IN1(g6313), .IN2(g225), .QN(n9711) );
  NAND2X0 U9649 ( .IN1(g6231), .IN2(g222), .QN(n9710) );
  NAND2X0 U9650 ( .IN1(g165), .IN2(g228), .QN(n9709) );
  XNOR2X1 U9651 ( .IN1(g113), .IN2(n7684), .Q(n9681) );
  INVX0 U9652 ( .INP(n9240), .ZN(n7684) );
  NAND3X0 U9653 ( .IN1(n9712), .IN2(n9713), .IN3(n9714), .QN(n9240) );
  NAND2X0 U9654 ( .IN1(g6313), .IN2(g207), .QN(n9714) );
  NAND2X0 U9655 ( .IN1(g6231), .IN2(g204), .QN(n9713) );
  NAND2X0 U9656 ( .IN1(g165), .IN2(g210), .QN(n9712) );
  NAND2X0 U9657 ( .IN1(n9685), .IN2(n9678), .QN(n9679) );
  XOR2X1 U9658 ( .IN1(g121), .IN2(n7672), .Q(n9678) );
  AND3X1 U9659 ( .IN1(n9715), .IN2(n9716), .IN3(n9717), .Q(n7672) );
  NAND2X0 U9660 ( .IN1(g213), .IN2(g6231), .QN(n9717) );
  NAND2X0 U9661 ( .IN1(g216), .IN2(g6313), .QN(n9716) );
  NAND2X0 U9662 ( .IN1(g219), .IN2(g165), .QN(n9715) );
  INVX0 U9663 ( .INP(n9674), .ZN(n9685) );
  XOR2X1 U9664 ( .IN1(n4513), .IN2(n4380), .Q(n9674) );
  XNOR2X1 U9665 ( .IN1(g105), .IN2(n7686), .Q(n9686) );
  INVX0 U9666 ( .INP(n8651), .ZN(n7686) );
  NAND3X0 U9667 ( .IN1(n9718), .IN2(n9719), .IN3(n9720), .QN(n8651) );
  NAND2X0 U9668 ( .IN1(g6313), .IN2(g198), .QN(n9720) );
  NAND2X0 U9669 ( .IN1(g6231), .IN2(g195), .QN(n9719) );
  NAND2X0 U9670 ( .IN1(g165), .IN2(g201), .QN(n9718) );
  AND3X1 U9671 ( .IN1(n9695), .IN2(n9696), .IN3(n9697), .Q(n9707) );
  INVX0 U9672 ( .INP(n9700), .ZN(n9697) );
  XNOR2X1 U9673 ( .IN1(g117), .IN2(n9098), .Q(n9700) );
  INVX0 U9674 ( .INP(n7675), .ZN(n9098) );
  NAND3X0 U9675 ( .IN1(n9721), .IN2(n9722), .IN3(n9723), .QN(n7675) );
  NAND2X0 U9676 ( .IN1(g6313), .IN2(g252), .QN(n9723) );
  NAND2X0 U9677 ( .IN1(g6231), .IN2(g249), .QN(n9722) );
  NAND2X0 U9678 ( .IN1(test_so14), .IN2(g165), .QN(n9721) );
  XOR2X1 U9679 ( .IN1(n4392), .IN2(n8775), .Q(n9696) );
  NAND3X0 U9680 ( .IN1(n9724), .IN2(n9725), .IN3(n9726), .QN(n8775) );
  NAND2X0 U9681 ( .IN1(g6313), .IN2(g243), .QN(n9726) );
  NAND2X0 U9682 ( .IN1(g6231), .IN2(g240), .QN(n9725) );
  NAND2X0 U9683 ( .IN1(g165), .IN2(g246), .QN(n9724) );
  XOR2X1 U9684 ( .IN1(n4290), .IN2(n7673), .Q(n9695) );
  NAND3X0 U9685 ( .IN1(n9727), .IN2(n9728), .IN3(n9729), .QN(n7673) );
  NAND2X0 U9686 ( .IN1(g6313), .IN2(g261), .QN(n9729) );
  NAND2X0 U9687 ( .IN1(g6231), .IN2(g258), .QN(n9728) );
  NAND2X0 U9688 ( .IN1(g165), .IN2(g264), .QN(n9727) );
  INVX0 U9689 ( .INP(n9693), .ZN(n9701) );
  XOR2X1 U9690 ( .IN1(n4376), .IN2(n7674), .Q(n9693) );
  INVX0 U9691 ( .INP(n9221), .ZN(n7674) );
  NAND3X0 U9692 ( .IN1(n9730), .IN2(n9731), .IN3(n9732), .QN(n9221) );
  NAND2X0 U9693 ( .IN1(g6313), .IN2(g234), .QN(n9732) );
  NAND2X0 U9694 ( .IN1(g6231), .IN2(g231), .QN(n9731) );
  NAND2X0 U9695 ( .IN1(g165), .IN2(g237), .QN(n9730) );
  INVX0 U9696 ( .INP(n9704), .ZN(n9694) );
  XOR2X1 U9697 ( .IN1(n7676), .IN2(n8680), .Q(n9704) );
  AND3X1 U9698 ( .IN1(n9733), .IN2(n9734), .IN3(n9735), .Q(n7676) );
  NAND2X0 U9699 ( .IN1(g267), .IN2(g6231), .QN(n9735) );
  NAND2X0 U9700 ( .IN1(g270), .IN2(g6313), .QN(n9734) );
  NAND2X0 U9701 ( .IN1(g273), .IN2(g165), .QN(n9733) );
  AND3X1 U9702 ( .IN1(n9736), .IN2(n2982), .IN3(n9737), .Q(g29112) );
  NAND2X0 U9703 ( .IN1(n6969), .IN2(n9738), .QN(n9737) );
  OR2X1 U9704 ( .IN1(n9738), .IN2(n6969), .Q(n2982) );
  INVX0 U9705 ( .INP(n3159), .ZN(n9738) );
  AND3X1 U9706 ( .IN1(n9739), .IN2(n2985), .IN3(n9740), .Q(g29111) );
  NAND2X0 U9707 ( .IN1(n6970), .IN2(n9741), .QN(n9740) );
  OR2X1 U9708 ( .IN1(n9741), .IN2(n6970), .Q(n2985) );
  INVX0 U9709 ( .INP(n3163), .ZN(n9741) );
  NOR3X0 U9710 ( .IN1(n9742), .IN2(n9322), .IN3(n9329), .QN(g29110) );
  INVX0 U9711 ( .INP(n2988), .ZN(n9329) );
  NAND2X0 U9712 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NOR2X0 U9713 ( .IN1(n3167), .IN2(test_so36), .QN(n9742) );
  AND3X1 U9714 ( .IN1(n9743), .IN2(n2991), .IN3(n9744), .Q(g29109) );
  NAND2X0 U9715 ( .IN1(n6971), .IN2(n9745), .QN(n9744) );
  OR2X1 U9716 ( .IN1(n9745), .IN2(n6971), .Q(n2991) );
  INVX0 U9717 ( .INP(n3171), .ZN(n9745) );
  AND2X1 U9718 ( .IN1(n9746), .IN2(n9747), .Q(g28990) );
  NAND2X0 U9719 ( .IN1(g1886), .IN2(DFF_1133_n1), .QN(n9747) );
  NAND2X0 U9720 ( .IN1(n4493), .IN2(n9748), .QN(n9746) );
  NAND2X0 U9721 ( .IN1(n9749), .IN2(n9750), .QN(n9748) );
  NAND2X0 U9722 ( .IN1(n4315), .IN2(DFF_1142_n1), .QN(n9750) );
  NAND2X0 U9723 ( .IN1(n8353), .IN2(g7194), .QN(n9749) );
  NAND2X0 U9724 ( .IN1(n9751), .IN2(n9752), .QN(n8353) );
  NAND2X0 U9725 ( .IN1(g1192), .IN2(DFF_783_n1), .QN(n9752) );
  NAND2X0 U9726 ( .IN1(n4454), .IN2(n9753), .QN(n9751) );
  NAND2X0 U9727 ( .IN1(n9754), .IN2(n9755), .QN(n9753) );
  NAND2X0 U9728 ( .IN1(n4316), .IN2(DFF_792_n1), .QN(n9755) );
  NAND2X0 U9729 ( .IN1(n8352), .IN2(g6944), .QN(n9754) );
  NAND2X0 U9730 ( .IN1(n9756), .IN2(n9757), .QN(n8352) );
  NAND2X0 U9731 ( .IN1(n6681), .IN2(g506), .QN(n9757) );
  NAND3X0 U9732 ( .IN1(n6682), .IN2(n4372), .IN3(n4570), .QN(n9756) );
  AND2X1 U9733 ( .IN1(n9758), .IN2(n9759), .Q(g28903) );
  NAND2X0 U9734 ( .IN1(n4488), .IN2(n7978), .QN(n9759) );
  NAND3X0 U9735 ( .IN1(n9760), .IN2(n9761), .IN3(g1680), .QN(n9758) );
  NAND2X0 U9736 ( .IN1(g26183), .IN2(g7014), .QN(n9761) );
  NAND2X0 U9737 ( .IN1(n4525), .IN2(g1686), .QN(n9760) );
  NAND2X0 U9738 ( .IN1(n9762), .IN2(n9763), .QN(g28788) );
  NAND2X0 U9739 ( .IN1(n9764), .IN2(g2501), .QN(n9763) );
  NAND2X0 U9740 ( .IN1(n9765), .IN2(n8841), .QN(n9764) );
  NAND2X0 U9741 ( .IN1(n9766), .IN2(n8841), .QN(n9762) );
  NAND2X0 U9742 ( .IN1(n9767), .IN2(n9768), .QN(g28783) );
  NAND2X0 U9743 ( .IN1(n9769), .IN2(g2503), .QN(n9768) );
  NAND2X0 U9744 ( .IN1(n9765), .IN2(n8449), .QN(n9769) );
  NAND2X0 U9745 ( .IN1(n9766), .IN2(n8449), .QN(n9767) );
  NAND2X0 U9746 ( .IN1(n9770), .IN2(n9771), .QN(g28782) );
  NAND2X0 U9747 ( .IN1(n4606), .IN2(n9772), .QN(n9771) );
  NAND2X0 U9748 ( .IN1(n4509), .IN2(test_so80), .QN(n9770) );
  NAND2X0 U9749 ( .IN1(n9773), .IN2(n9774), .QN(g28778) );
  NAND2X0 U9750 ( .IN1(n9775), .IN2(g1807), .QN(n9774) );
  NAND2X0 U9751 ( .IN1(n9776), .IN2(n8453), .QN(n9775) );
  NAND2X0 U9752 ( .IN1(n9777), .IN2(n8453), .QN(n9773) );
  NAND2X0 U9753 ( .IN1(n9778), .IN2(n9779), .QN(g28774) );
  NAND2X0 U9754 ( .IN1(n9780), .IN2(g2502), .QN(n9779) );
  NAND2X0 U9755 ( .IN1(n9765), .IN2(n8456), .QN(n9780) );
  AND3X1 U9756 ( .IN1(test_so79), .IN2(n9781), .IN3(n9782), .Q(n9765) );
  NAND2X0 U9757 ( .IN1(n9766), .IN2(n8456), .QN(n9778) );
  INVX0 U9758 ( .INP(n9783), .ZN(n9766) );
  NAND2X0 U9759 ( .IN1(n9784), .IN2(n9785), .QN(g28773) );
  NAND2X0 U9760 ( .IN1(g7264), .IN2(n9772), .QN(n9785) );
  NAND2X0 U9761 ( .IN1(n4524), .IN2(g2486), .QN(n9784) );
  NAND2X0 U9762 ( .IN1(n9786), .IN2(n9787), .QN(g28772) );
  NAND2X0 U9763 ( .IN1(n9788), .IN2(g1809), .QN(n9787) );
  NAND2X0 U9764 ( .IN1(n9776), .IN2(n8459), .QN(n9788) );
  NAND2X0 U9765 ( .IN1(n9777), .IN2(n8459), .QN(n9786) );
  NAND2X0 U9766 ( .IN1(n9789), .IN2(n9790), .QN(g28771) );
  NAND2X0 U9767 ( .IN1(n4618), .IN2(n9791), .QN(n9790) );
  NAND2X0 U9768 ( .IN1(n4511), .IN2(g1795), .QN(n9789) );
  NAND2X0 U9769 ( .IN1(n9792), .IN2(n9793), .QN(g28767) );
  NAND2X0 U9770 ( .IN1(n9794), .IN2(g1113), .QN(n9793) );
  NAND2X0 U9771 ( .IN1(n9795), .IN2(g1088), .QN(n9794) );
  NAND2X0 U9772 ( .IN1(n9796), .IN2(g1088), .QN(n9792) );
  NAND2X0 U9773 ( .IN1(n9797), .IN2(n9798), .QN(g28763) );
  NAND2X0 U9774 ( .IN1(g5555), .IN2(n9772), .QN(n9798) );
  NAND2X0 U9775 ( .IN1(n9783), .IN2(n9799), .QN(n9772) );
  NAND2X0 U9776 ( .IN1(n9800), .IN2(n9349), .QN(n9799) );
  NAND2X0 U9777 ( .IN1(test_so79), .IN2(n9801), .QN(n9800) );
  NAND2X0 U9778 ( .IN1(n9782), .IN2(n9781), .QN(n9801) );
  INVX0 U9779 ( .INP(n9348), .ZN(n9782) );
  NAND3X0 U9780 ( .IN1(n9802), .IN2(n9803), .IN3(n9804), .QN(n9348) );
  NAND2X0 U9781 ( .IN1(n6938), .IN2(n8449), .QN(n9804) );
  NAND2X0 U9782 ( .IN1(n6947), .IN2(n8841), .QN(n9803) );
  NAND2X0 U9783 ( .IN1(n6948), .IN2(n8456), .QN(n9802) );
  NAND3X0 U9784 ( .IN1(test_so79), .IN2(n9781), .IN3(n8329), .QN(n9783) );
  INVX0 U9785 ( .INP(n9349), .ZN(n8329) );
  NAND3X0 U9786 ( .IN1(n9805), .IN2(n9806), .IN3(n9807), .QN(n9349) );
  NAND2X0 U9787 ( .IN1(g5555), .IN2(g2483), .QN(n9807) );
  NAND2X0 U9788 ( .IN1(test_so80), .IN2(n4606), .QN(n9806) );
  NAND2X0 U9789 ( .IN1(g7264), .IN2(g2486), .QN(n9805) );
  NAND2X0 U9790 ( .IN1(n9808), .IN2(n9809), .QN(n9781) );
  NAND2X0 U9791 ( .IN1(n9345), .IN2(n4285), .QN(n9809) );
  NAND3X0 U9792 ( .IN1(n8328), .IN2(n8840), .IN3(n9342), .QN(n9808) );
  NAND2X0 U9793 ( .IN1(n673), .IN2(g2257), .QN(n8840) );
  AND3X1 U9794 ( .IN1(n9810), .IN2(n9811), .IN3(n9812), .Q(n673) );
  NAND2X0 U9795 ( .IN1(test_so73), .IN2(n6858), .QN(n9812) );
  NAND2X0 U9796 ( .IN1(n6859), .IN2(g6837), .QN(n9811) );
  NAND2X0 U9797 ( .IN1(n6857), .IN2(g2241), .QN(n9810) );
  INVX0 U9798 ( .INP(n9345), .ZN(n8328) );
  NAND3X0 U9799 ( .IN1(n8719), .IN2(n9813), .IN3(n9814), .QN(n9345) );
  NAND2X0 U9800 ( .IN1(n4516), .IN2(g2483), .QN(n9797) );
  NAND2X0 U9801 ( .IN1(n9815), .IN2(n9816), .QN(g28761) );
  NAND2X0 U9802 ( .IN1(n9817), .IN2(g1808), .QN(n9816) );
  NAND2X0 U9803 ( .IN1(n9776), .IN2(n8494), .QN(n9817) );
  AND3X1 U9804 ( .IN1(n9818), .IN2(g1690), .IN3(n9819), .Q(n9776) );
  NAND2X0 U9805 ( .IN1(n9777), .IN2(n8494), .QN(n9815) );
  INVX0 U9806 ( .INP(n9820), .ZN(n9777) );
  NAND2X0 U9807 ( .IN1(n9821), .IN2(n9822), .QN(g28760) );
  NAND2X0 U9808 ( .IN1(g7014), .IN2(n9791), .QN(n9822) );
  NAND2X0 U9809 ( .IN1(n4525), .IN2(g1792), .QN(n9821) );
  NAND2X0 U9810 ( .IN1(n9823), .IN2(n9824), .QN(g28759) );
  NAND2X0 U9811 ( .IN1(n9825), .IN2(g1115), .QN(n9824) );
  NAND2X0 U9812 ( .IN1(n9795), .IN2(g6712), .QN(n9825) );
  NAND2X0 U9813 ( .IN1(n9796), .IN2(g6712), .QN(n9823) );
  NAND2X0 U9814 ( .IN1(n9826), .IN2(n9827), .QN(g28758) );
  NAND2X0 U9815 ( .IN1(n4381), .IN2(g1101), .QN(n9827) );
  NAND2X0 U9816 ( .IN1(n9828), .IN2(g1088), .QN(n9826) );
  NAND2X0 U9817 ( .IN1(n9829), .IN2(n9830), .QN(g28754) );
  NAND2X0 U9818 ( .IN1(n9831), .IN2(g426), .QN(n9830) );
  NAND2X0 U9819 ( .IN1(n9832), .IN2(n8500), .QN(n9831) );
  NAND2X0 U9820 ( .IN1(n9833), .IN2(n8500), .QN(n9829) );
  NAND2X0 U9821 ( .IN1(n9834), .IN2(n9835), .QN(g28749) );
  NAND2X0 U9822 ( .IN1(g5511), .IN2(n9791), .QN(n9835) );
  NAND2X0 U9823 ( .IN1(n9820), .IN2(n9836), .QN(n9791) );
  NAND2X0 U9824 ( .IN1(n9837), .IN2(n9364), .QN(n9836) );
  NAND2X0 U9825 ( .IN1(g1690), .IN2(n9838), .QN(n9837) );
  NAND2X0 U9826 ( .IN1(n9819), .IN2(n9818), .QN(n9838) );
  INVX0 U9827 ( .INP(n9363), .ZN(n9819) );
  NAND3X0 U9828 ( .IN1(n9839), .IN2(n9840), .IN3(n9841), .QN(n9363) );
  NAND2X0 U9829 ( .IN1(n6941), .IN2(n8459), .QN(n9841) );
  NAND2X0 U9830 ( .IN1(n6952), .IN2(n8453), .QN(n9840) );
  NAND2X0 U9831 ( .IN1(n6953), .IN2(n8494), .QN(n9839) );
  NAND3X0 U9832 ( .IN1(n9818), .IN2(g1690), .IN3(n8326), .QN(n9820) );
  INVX0 U9833 ( .INP(n9364), .ZN(n8326) );
  NAND3X0 U9834 ( .IN1(n9842), .IN2(n9843), .IN3(n9844), .QN(n9364) );
  NAND2X0 U9835 ( .IN1(g5511), .IN2(g1789), .QN(n9844) );
  NAND2X0 U9836 ( .IN1(n4618), .IN2(g1795), .QN(n9843) );
  NAND2X0 U9837 ( .IN1(g7014), .IN2(g1792), .QN(n9842) );
  NAND2X0 U9838 ( .IN1(n9845), .IN2(n9846), .QN(n9818) );
  NAND2X0 U9839 ( .IN1(n9847), .IN2(n4284), .QN(n9846) );
  NAND3X0 U9840 ( .IN1(n8325), .IN2(n8493), .IN3(n9358), .QN(n9845) );
  NAND2X0 U9841 ( .IN1(n509), .IN2(g1563), .QN(n8493) );
  AND3X1 U9842 ( .IN1(n9848), .IN2(n9849), .IN3(n9850), .Q(n509) );
  NAND2X0 U9843 ( .IN1(n6869), .IN2(g6782), .QN(n9850) );
  NAND2X0 U9844 ( .IN1(n6870), .IN2(g6573), .QN(n9849) );
  NAND2X0 U9845 ( .IN1(n6868), .IN2(g1547), .QN(n9848) );
  INVX0 U9846 ( .INP(n9847), .ZN(n8325) );
  NAND3X0 U9847 ( .IN1(n9851), .IN2(n8756), .IN3(n9852), .QN(n9847) );
  NAND2X0 U9848 ( .IN1(n4518), .IN2(g1789), .QN(n9834) );
  NAND2X0 U9849 ( .IN1(n9853), .IN2(n9854), .QN(g28747) );
  NAND2X0 U9850 ( .IN1(n9855), .IN2(g1114), .QN(n9854) );
  NAND2X0 U9851 ( .IN1(n9795), .IN2(g5472), .QN(n9855) );
  AND3X1 U9852 ( .IN1(n9856), .IN2(g996), .IN3(n9857), .Q(n9795) );
  NAND2X0 U9853 ( .IN1(n9796), .IN2(g5472), .QN(n9853) );
  INVX0 U9854 ( .INP(n9858), .ZN(n9796) );
  NAND2X0 U9855 ( .IN1(n9859), .IN2(n9860), .QN(g28746) );
  NAND2X0 U9856 ( .IN1(n4364), .IN2(g1098), .QN(n9860) );
  NAND2X0 U9857 ( .IN1(n9828), .IN2(g6712), .QN(n9859) );
  NAND2X0 U9858 ( .IN1(n9861), .IN2(n9862), .QN(g28745) );
  NAND2X0 U9859 ( .IN1(n9863), .IN2(g428), .QN(n9862) );
  NAND2X0 U9860 ( .IN1(n9832), .IN2(n8861), .QN(n9863) );
  NAND2X0 U9861 ( .IN1(n9833), .IN2(n8861), .QN(n9861) );
  NAND2X0 U9862 ( .IN1(n9864), .IN2(n9865), .QN(g28744) );
  NAND2X0 U9863 ( .IN1(n4640), .IN2(n9866), .QN(n9865) );
  NAND2X0 U9864 ( .IN1(n4506), .IN2(g414), .QN(n9864) );
  NAND2X0 U9865 ( .IN1(n9867), .IN2(n9868), .QN(g28738) );
  NAND2X0 U9866 ( .IN1(n4363), .IN2(g1095), .QN(n9868) );
  NAND2X0 U9867 ( .IN1(n9828), .IN2(g5472), .QN(n9867) );
  NAND2X0 U9868 ( .IN1(n9858), .IN2(n9869), .QN(n9828) );
  NAND2X0 U9869 ( .IN1(n9870), .IN2(n9380), .QN(n9869) );
  NAND2X0 U9870 ( .IN1(g996), .IN2(n9871), .QN(n9870) );
  NAND2X0 U9871 ( .IN1(n9857), .IN2(n9856), .QN(n9871) );
  INVX0 U9872 ( .INP(n9379), .ZN(n9857) );
  NAND3X0 U9873 ( .IN1(n9872), .IN2(n9873), .IN3(n9874), .QN(n9379) );
  NAND2X0 U9874 ( .IN1(n6958), .IN2(g1088), .QN(n9874) );
  NAND2X0 U9875 ( .IN1(n6959), .IN2(g5472), .QN(n9873) );
  NAND2X0 U9876 ( .IN1(n6944), .IN2(g6712), .QN(n9872) );
  NAND3X0 U9877 ( .IN1(n9856), .IN2(g996), .IN3(n8323), .QN(n9858) );
  INVX0 U9878 ( .INP(n9380), .ZN(n8323) );
  NAND3X0 U9879 ( .IN1(n9875), .IN2(n9876), .IN3(n9877), .QN(n9380) );
  NAND2X0 U9880 ( .IN1(g1088), .IN2(g1101), .QN(n9877) );
  NAND2X0 U9881 ( .IN1(g5472), .IN2(g1095), .QN(n9876) );
  NAND2X0 U9882 ( .IN1(g6712), .IN2(g1098), .QN(n9875) );
  NAND2X0 U9883 ( .IN1(n9878), .IN2(n9879), .QN(n9856) );
  NAND2X0 U9884 ( .IN1(n9376), .IN2(n4283), .QN(n9879) );
  NAND3X0 U9885 ( .IN1(n8322), .IN2(n8371), .IN3(n9373), .QN(n9878) );
  NAND2X0 U9886 ( .IN1(n335), .IN2(g869), .QN(n8371) );
  AND3X1 U9887 ( .IN1(n9880), .IN2(n9881), .IN3(n9882), .Q(n335) );
  NAND2X0 U9888 ( .IN1(n6880), .IN2(test_so31), .QN(n9882) );
  OR2X1 U9889 ( .IN1(n4312), .IN2(test_so33), .Q(n9881) );
  NAND2X0 U9890 ( .IN1(n6881), .IN2(g6368), .QN(n9880) );
  INVX0 U9891 ( .INP(n9376), .ZN(n8322) );
  NAND3X0 U9892 ( .IN1(n8790), .IN2(n9883), .IN3(n9884), .QN(n9376) );
  NAND2X0 U9893 ( .IN1(n9885), .IN2(n9886), .QN(g28736) );
  NAND2X0 U9894 ( .IN1(test_so17), .IN2(n9887), .QN(n9886) );
  NAND2X0 U9895 ( .IN1(n9832), .IN2(n8537), .QN(n9887) );
  AND3X1 U9896 ( .IN1(n9888), .IN2(g309), .IN3(n9889), .Q(n9832) );
  NAND2X0 U9897 ( .IN1(n9833), .IN2(n8537), .QN(n9885) );
  INVX0 U9898 ( .INP(n9890), .ZN(n9833) );
  NAND2X0 U9899 ( .IN1(n9891), .IN2(n9892), .QN(g28735) );
  NAND2X0 U9900 ( .IN1(g6447), .IN2(n9866), .QN(n9892) );
  NAND2X0 U9901 ( .IN1(n4499), .IN2(g411), .QN(n9891) );
  NAND2X0 U9902 ( .IN1(n9893), .IN2(n9894), .QN(g28732) );
  NAND2X0 U9903 ( .IN1(g5437), .IN2(n9866), .QN(n9894) );
  NAND2X0 U9904 ( .IN1(n9890), .IN2(n9895), .QN(n9866) );
  NAND2X0 U9905 ( .IN1(n9896), .IN2(n9392), .QN(n9895) );
  NAND2X0 U9906 ( .IN1(g309), .IN2(n9897), .QN(n9896) );
  NAND2X0 U9907 ( .IN1(n9889), .IN2(n9888), .QN(n9897) );
  INVX0 U9908 ( .INP(n9391), .ZN(n9889) );
  NAND3X0 U9909 ( .IN1(n9898), .IN2(n9899), .IN3(n9900), .QN(n9391) );
  OR2X1 U9910 ( .IN1(n4520), .IN2(test_so17), .Q(n9900) );
  NAND2X0 U9911 ( .IN1(n6967), .IN2(n8861), .QN(n9899) );
  NAND2X0 U9912 ( .IN1(n6966), .IN2(n8500), .QN(n9898) );
  NAND3X0 U9913 ( .IN1(n9888), .IN2(g309), .IN3(n8320), .QN(n9890) );
  INVX0 U9914 ( .INP(n9392), .ZN(n8320) );
  NAND3X0 U9915 ( .IN1(n9901), .IN2(n9902), .IN3(n9903), .QN(n9392) );
  NAND2X0 U9916 ( .IN1(g5437), .IN2(g408), .QN(n9903) );
  NAND2X0 U9917 ( .IN1(n4640), .IN2(g414), .QN(n9902) );
  NAND2X0 U9918 ( .IN1(g6447), .IN2(g411), .QN(n9901) );
  NAND2X0 U9919 ( .IN1(n9904), .IN2(n9905), .QN(n9888) );
  NAND2X0 U9920 ( .IN1(n9906), .IN2(n4282), .QN(n9905) );
  NAND3X0 U9921 ( .IN1(n8319), .IN2(n8536), .IN3(n9386), .QN(n9904) );
  NAND2X0 U9922 ( .IN1(n167), .IN2(g181), .QN(n8536) );
  AND3X1 U9923 ( .IN1(n9907), .IN2(n9908), .IN3(n9909), .Q(n167) );
  NAND2X0 U9924 ( .IN1(n6892), .IN2(g6313), .QN(n9909) );
  NAND2X0 U9925 ( .IN1(n6893), .IN2(g6231), .QN(n9908) );
  NAND2X0 U9926 ( .IN1(n6891), .IN2(g165), .QN(n9907) );
  INVX0 U9927 ( .INP(n9906), .ZN(n8319) );
  NAND3X0 U9928 ( .IN1(n8810), .IN2(n9910), .IN3(n9911), .QN(n9906) );
  NAND2X0 U9929 ( .IN1(n4520), .IN2(g408), .QN(n9893) );
  NOR2X0 U9930 ( .IN1(n9912), .IN2(n9913), .QN(g28668) );
  XOR2X1 U9931 ( .IN1(n4418), .IN2(n9914), .Q(n9913) );
  NOR2X0 U9932 ( .IN1(n4396), .IN2(n9915), .QN(n9914) );
  NOR2X0 U9933 ( .IN1(n9318), .IN2(n9916), .QN(g28637) );
  XNOR2X1 U9934 ( .IN1(n6979), .IN2(n3160), .Q(n9916) );
  NOR2X0 U9935 ( .IN1(n9320), .IN2(n9917), .QN(g28636) );
  XNOR2X1 U9936 ( .IN1(n6983), .IN2(n3164), .Q(n9917) );
  NOR2X0 U9937 ( .IN1(n9322), .IN2(n9918), .QN(g28635) );
  XOR2X1 U9938 ( .IN1(n6987), .IN2(n9919), .Q(n9918) );
  NOR2X0 U9939 ( .IN1(n9324), .IN2(n9920), .QN(g28634) );
  XNOR2X1 U9940 ( .IN1(n6991), .IN2(n3172), .Q(n9920) );
  NAND2X0 U9941 ( .IN1(n9921), .IN2(n9922), .QN(g28425) );
  OR2X1 U9942 ( .IN1(g3109), .IN2(n4343), .Q(n9922) );
  NAND2X0 U9943 ( .IN1(n7265), .IN2(g3109), .QN(n9921) );
  NAND2X0 U9944 ( .IN1(n9923), .IN2(n9924), .QN(g28421) );
  NAND2X0 U9945 ( .IN1(n4383), .IN2(test_so7), .QN(n9924) );
  NAND2X0 U9946 ( .IN1(n7265), .IN2(g8030), .QN(n9923) );
  NAND2X0 U9947 ( .IN1(n9925), .IN2(n9926), .QN(g28420) );
  NAND2X0 U9948 ( .IN1(n4382), .IN2(g3100), .QN(n9926) );
  NAND2X0 U9949 ( .IN1(n7265), .IN2(g8106), .QN(n9925) );
  AND2X1 U9950 ( .IN1(n9927), .IN2(n9928), .Q(n7265) );
  NAND2X0 U9951 ( .IN1(n6407), .IN2(g1186), .QN(n9928) );
  NAND3X0 U9952 ( .IN1(n9929), .IN2(n9930), .IN3(n4548), .QN(n9927) );
  NAND2X0 U9953 ( .IN1(g6750), .IN2(g21851), .QN(n9930) );
  NAND2X0 U9954 ( .IN1(n4371), .IN2(n4361), .QN(n9929) );
  NAND2X0 U9955 ( .IN1(n9931), .IN2(n9932), .QN(g28371) );
  NAND2X0 U9956 ( .IN1(n4299), .IN2(g2694), .QN(n9932) );
  NAND2X0 U9957 ( .IN1(n9933), .IN2(g2624), .QN(n9931) );
  NAND2X0 U9958 ( .IN1(n9934), .IN2(n9935), .QN(g28368) );
  NAND2X0 U9959 ( .IN1(n4370), .IN2(g2691), .QN(n9935) );
  NAND2X0 U9960 ( .IN1(n9933), .IN2(g7390), .QN(n9934) );
  NAND2X0 U9961 ( .IN1(n9936), .IN2(n9937), .QN(g28367) );
  NAND2X0 U9962 ( .IN1(n4299), .IN2(g2685), .QN(n9937) );
  NAND2X0 U9963 ( .IN1(n9938), .IN2(g2624), .QN(n9936) );
  NAND2X0 U9964 ( .IN1(n9939), .IN2(n9940), .QN(g28366) );
  NAND2X0 U9965 ( .IN1(n4366), .IN2(g2000), .QN(n9940) );
  NAND2X0 U9966 ( .IN1(n9941), .IN2(g1930), .QN(n9939) );
  NAND2X0 U9967 ( .IN1(n9942), .IN2(n9943), .QN(g28364) );
  NAND2X0 U9968 ( .IN1(n4314), .IN2(g2688), .QN(n9943) );
  NAND2X0 U9969 ( .IN1(n9933), .IN2(n9246), .QN(n9942) );
  NAND2X0 U9970 ( .IN1(n9944), .IN2(n9945), .QN(n9933) );
  NAND2X0 U9971 ( .IN1(n3252), .IN2(n9946), .QN(n9945) );
  NAND2X0 U9972 ( .IN1(n9947), .IN2(n7994), .QN(n9944) );
  NAND2X0 U9973 ( .IN1(n9948), .IN2(n9949), .QN(g28363) );
  NAND2X0 U9974 ( .IN1(n9938), .IN2(g7390), .QN(n9949) );
  NAND2X0 U9975 ( .IN1(n4370), .IN2(test_so90), .QN(n9948) );
  NAND2X0 U9976 ( .IN1(n9950), .IN2(n9951), .QN(g28362) );
  NAND2X0 U9977 ( .IN1(n4315), .IN2(g1997), .QN(n9951) );
  NAND2X0 U9978 ( .IN1(n9941), .IN2(g7194), .QN(n9950) );
  NAND2X0 U9979 ( .IN1(n9952), .IN2(n9953), .QN(g28361) );
  NAND2X0 U9980 ( .IN1(n4366), .IN2(g1991), .QN(n9953) );
  NAND2X0 U9981 ( .IN1(n9954), .IN2(g1930), .QN(n9952) );
  NAND2X0 U9982 ( .IN1(n9955), .IN2(n9956), .QN(g28360) );
  NAND2X0 U9983 ( .IN1(n4300), .IN2(g1306), .QN(n9956) );
  NAND2X0 U9984 ( .IN1(n9957), .IN2(g1236), .QN(n9955) );
  NAND2X0 U9985 ( .IN1(n9958), .IN2(n9959), .QN(g28358) );
  NAND2X0 U9986 ( .IN1(g7302), .IN2(n9938), .QN(n9959) );
  NAND2X0 U9987 ( .IN1(n9960), .IN2(n9961), .QN(n9938) );
  NAND2X0 U9988 ( .IN1(n9947), .IN2(n7981), .QN(n9961) );
  NAND4X0 U9989 ( .IN1(n8315), .IN2(n9962), .IN3(n8317), .IN4(n9946), .QN(
        n9960) );
  AND4X1 U9990 ( .IN1(n9963), .IN2(n9964), .IN3(n9965), .IN4(n9966), .Q(n8317)
         );
  NAND4X0 U9991 ( .IN1(n9967), .IN2(n9968), .IN3(n9969), .IN4(n9970), .QN(
        n9966) );
  OR2X1 U9992 ( .IN1(n9971), .IN2(n9972), .Q(n9969) );
  NAND2X0 U9993 ( .IN1(n9973), .IN2(n9974), .QN(n9967) );
  NAND2X0 U9994 ( .IN1(n9975), .IN2(n9976), .QN(n9973) );
  NAND4X0 U9995 ( .IN1(n9977), .IN2(n9978), .IN3(n9979), .IN4(n9980), .QN(
        n9965) );
  NAND2X0 U9996 ( .IN1(n9981), .IN2(n9974), .QN(n9979) );
  NAND2X0 U9997 ( .IN1(n9982), .IN2(n9983), .QN(n9977) );
  NAND3X0 U9998 ( .IN1(n9972), .IN2(n9971), .IN3(n9984), .QN(n9983) );
  NOR2X0 U9999 ( .IN1(n9974), .IN2(n9985), .QN(n9972) );
  NAND2X0 U10000 ( .IN1(n9986), .IN2(n9987), .QN(n9964) );
  NAND2X0 U10001 ( .IN1(n9988), .IN2(n9989), .QN(n9987) );
  NAND4X0 U10002 ( .IN1(n9971), .IN2(n9974), .IN3(n9990), .IN4(n9991), .QN(
        n9989) );
  NAND2X0 U10003 ( .IN1(n9980), .IN2(n9968), .QN(n9991) );
  NAND2X0 U10004 ( .IN1(n9975), .IN2(n9970), .QN(n9990) );
  NAND2X0 U10005 ( .IN1(n9981), .IN2(n9992), .QN(n9988) );
  NAND2X0 U10006 ( .IN1(n9975), .IN2(n9993), .QN(n9992) );
  NAND2X0 U10007 ( .IN1(n9982), .IN2(n9970), .QN(n9993) );
  NAND4X0 U10008 ( .IN1(n9994), .IN2(n9995), .IN3(n9996), .IN4(n9997), .QN(
        n9963) );
  NOR2X0 U10009 ( .IN1(n9998), .IN2(n9999), .QN(n9994) );
  NOR2X0 U10010 ( .IN1(n9970), .IN2(n10000), .QN(n9999) );
  NOR3X0 U10011 ( .IN1(n9985), .IN2(n10001), .IN3(n9980), .QN(n9998) );
  NAND2X0 U10012 ( .IN1(n3253), .IN2(n10002), .QN(n9962) );
  INVX0 U10013 ( .INP(n10003), .ZN(n10002) );
  AND3X1 U10014 ( .IN1(n10004), .IN2(n10005), .IN3(n10006), .Q(n3253) );
  NAND2X0 U10015 ( .IN1(n9970), .IN2(n10007), .QN(n10006) );
  NAND2X0 U10016 ( .IN1(n10008), .IN2(n10009), .QN(n10007) );
  NAND3X0 U10017 ( .IN1(n9974), .IN2(n10010), .IN3(n9971), .QN(n10009) );
  NAND2X0 U10018 ( .IN1(n9986), .IN2(n10011), .QN(n10008) );
  NAND2X0 U10019 ( .IN1(n10012), .IN2(n10013), .QN(n10011) );
  NAND2X0 U10020 ( .IN1(n9984), .IN2(n10014), .QN(n10013) );
  NAND2X0 U10021 ( .IN1(n10015), .IN2(n10016), .QN(n10014) );
  NAND3X0 U10022 ( .IN1(n9971), .IN2(n9976), .IN3(n9975), .QN(n10016) );
  NAND2X0 U10023 ( .IN1(n9982), .IN2(n10017), .QN(n10015) );
  NAND2X0 U10024 ( .IN1(n9996), .IN2(n9985), .QN(n10012) );
  NAND3X0 U10025 ( .IN1(n10018), .IN2(n9968), .IN3(n9996), .QN(n10005) );
  INVX0 U10026 ( .INP(n9971), .ZN(n9996) );
  NAND2X0 U10027 ( .IN1(n10019), .IN2(n9978), .QN(n10018) );
  NAND2X0 U10028 ( .IN1(n9986), .IN2(n9974), .QN(n9978) );
  NAND2X0 U10029 ( .IN1(n9980), .IN2(n9975), .QN(n10019) );
  NAND2X0 U10030 ( .IN1(n9997), .IN2(n10020), .QN(n10004) );
  NAND3X0 U10031 ( .IN1(n10021), .IN2(n9995), .IN3(n10022), .QN(n10020) );
  NAND3X0 U10032 ( .IN1(n9984), .IN2(n9975), .IN3(n9981), .QN(n10022) );
  INVX0 U10033 ( .INP(n9976), .ZN(n9981) );
  NAND3X0 U10034 ( .IN1(n10017), .IN2(n9968), .IN3(n9980), .QN(n9995) );
  NAND3X0 U10035 ( .IN1(n10023), .IN2(n9971), .IN3(n9980), .QN(n10021) );
  INVX0 U10036 ( .INP(n9970), .ZN(n9980) );
  NAND3X0 U10037 ( .IN1(n10024), .IN2(n10025), .IN3(n10026), .QN(n9970) );
  NAND2X0 U10038 ( .IN1(g5796), .IN2(g2426), .QN(n10026) );
  NAND2X0 U10039 ( .IN1(g5747), .IN2(g2424), .QN(n10025) );
  NAND2X0 U10040 ( .IN1(g2412), .IN2(g2428), .QN(n10024) );
  NAND3X0 U10041 ( .IN1(n10027), .IN2(n10028), .IN3(n10029), .QN(n9971) );
  NAND2X0 U10042 ( .IN1(g5796), .IN2(g2441), .QN(n10029) );
  NAND2X0 U10043 ( .IN1(g5747), .IN2(g2439), .QN(n10028) );
  NAND2X0 U10044 ( .IN1(g2412), .IN2(g2443), .QN(n10027) );
  NAND2X0 U10045 ( .IN1(n10030), .IN2(n10031), .QN(n10023) );
  NAND2X0 U10046 ( .IN1(n10001), .IN2(n9984), .QN(n10031) );
  NOR2X0 U10047 ( .IN1(n10010), .IN2(n10017), .QN(n10001) );
  INVX0 U10048 ( .INP(n9974), .ZN(n10017) );
  NAND3X0 U10049 ( .IN1(n10032), .IN2(n10033), .IN3(n10034), .QN(n9974) );
  NAND2X0 U10050 ( .IN1(g5796), .IN2(g2456), .QN(n10034) );
  NAND2X0 U10051 ( .IN1(g5747), .IN2(g2454), .QN(n10033) );
  NAND2X0 U10052 ( .IN1(g2412), .IN2(g2458), .QN(n10032) );
  NAND2X0 U10053 ( .IN1(n9985), .IN2(n9976), .QN(n10030) );
  NAND3X0 U10054 ( .IN1(n10035), .IN2(n10036), .IN3(n10037), .QN(n9976) );
  NAND2X0 U10055 ( .IN1(g5796), .IN2(g2471), .QN(n10037) );
  NAND2X0 U10056 ( .IN1(g5747), .IN2(g2469), .QN(n10036) );
  NAND2X0 U10057 ( .IN1(test_so85), .IN2(g2412), .QN(n10035) );
  NAND2X0 U10058 ( .IN1(n8318), .IN2(n10003), .QN(n8315) );
  NAND2X0 U10059 ( .IN1(n4314), .IN2(g2679), .QN(n9958) );
  NAND2X0 U10060 ( .IN1(n10038), .IN2(n10039), .QN(g28357) );
  NAND2X0 U10061 ( .IN1(n4296), .IN2(g1994), .QN(n10039) );
  NAND2X0 U10062 ( .IN1(n9941), .IN2(n9268), .QN(n10038) );
  NAND2X0 U10063 ( .IN1(n10040), .IN2(n10041), .QN(n9941) );
  NAND2X0 U10064 ( .IN1(n9947), .IN2(n8181), .QN(n10041) );
  NAND4X0 U10065 ( .IN1(n10042), .IN2(n10043), .IN3(n10044), .IN4(n9946), .QN(
        n10040) );
  NAND2X0 U10066 ( .IN1(n10045), .IN2(n10046), .QN(n10042) );
  INVX0 U10067 ( .INP(n10047), .ZN(n10045) );
  NAND2X0 U10068 ( .IN1(n10048), .IN2(n10049), .QN(g28356) );
  NAND2X0 U10069 ( .IN1(n4315), .IN2(g1988), .QN(n10049) );
  NAND2X0 U10070 ( .IN1(n9954), .IN2(g7194), .QN(n10048) );
  NAND2X0 U10071 ( .IN1(n10050), .IN2(n10051), .QN(g28355) );
  NAND2X0 U10072 ( .IN1(n4316), .IN2(g1303), .QN(n10051) );
  NAND2X0 U10073 ( .IN1(n9957), .IN2(g6944), .QN(n10050) );
  NAND2X0 U10074 ( .IN1(n10052), .IN2(n10053), .QN(g28354) );
  NAND2X0 U10075 ( .IN1(n4300), .IN2(g1297), .QN(n10053) );
  NAND2X0 U10076 ( .IN1(n10054), .IN2(g1236), .QN(n10052) );
  NAND2X0 U10077 ( .IN1(n10055), .IN2(n10056), .QN(g28353) );
  NAND2X0 U10078 ( .IN1(n10057), .IN2(g550), .QN(n10056) );
  NAND2X0 U10079 ( .IN1(n4313), .IN2(test_so26), .QN(n10055) );
  NAND2X0 U10080 ( .IN1(n10058), .IN2(n10059), .QN(g28352) );
  NAND2X0 U10081 ( .IN1(g7052), .IN2(n9954), .QN(n10059) );
  NAND2X0 U10082 ( .IN1(n10060), .IN2(n10061), .QN(n9954) );
  NAND2X0 U10083 ( .IN1(n9947), .IN2(n8173), .QN(n10061) );
  NAND4X0 U10084 ( .IN1(n10043), .IN2(n10062), .IN3(n10046), .IN4(n9946), .QN(
        n10060) );
  AND4X1 U10085 ( .IN1(n10063), .IN2(n10064), .IN3(n10065), .IN4(n10066), .Q(
        n10046) );
  NAND2X0 U10086 ( .IN1(n10067), .IN2(n10068), .QN(n10066) );
  NAND2X0 U10087 ( .IN1(n10069), .IN2(n10070), .QN(n10067) );
  NAND3X0 U10088 ( .IN1(n10071), .IN2(n10072), .IN3(n10073), .QN(n10070) );
  NAND2X0 U10089 ( .IN1(n10074), .IN2(n10075), .QN(n10069) );
  NAND2X0 U10090 ( .IN1(n10076), .IN2(n10077), .QN(n10075) );
  NAND2X0 U10091 ( .IN1(n10078), .IN2(n10079), .QN(n10077) );
  INVX0 U10092 ( .INP(n10080), .ZN(n10076) );
  NAND2X0 U10093 ( .IN1(n10081), .IN2(n10082), .QN(n10065) );
  NAND2X0 U10094 ( .IN1(n10083), .IN2(n10084), .QN(n10082) );
  NAND3X0 U10095 ( .IN1(n10085), .IN2(n10079), .IN3(n10080), .QN(n10084) );
  NAND2X0 U10096 ( .IN1(n10086), .IN2(n10087), .QN(n10080) );
  NAND2X0 U10097 ( .IN1(n10088), .IN2(n10089), .QN(n10087) );
  NAND2X0 U10098 ( .IN1(n10090), .IN2(n10073), .QN(n10086) );
  NAND2X0 U10099 ( .IN1(n10091), .IN2(n10078), .QN(n10083) );
  NAND2X0 U10100 ( .IN1(n10092), .IN2(n10093), .QN(n10078) );
  NAND2X0 U10101 ( .IN1(n10094), .IN2(n10089), .QN(n10093) );
  NAND3X0 U10102 ( .IN1(n10095), .IN2(n10071), .IN3(n10096), .QN(n10064) );
  NAND2X0 U10103 ( .IN1(n10097), .IN2(n10098), .QN(n10063) );
  NAND3X0 U10104 ( .IN1(n10099), .IN2(n10100), .IN3(n10101), .QN(n10098) );
  NAND2X0 U10105 ( .IN1(n10095), .IN2(n10102), .QN(n10101) );
  NAND2X0 U10106 ( .IN1(n10096), .IN2(n10089), .QN(n10100) );
  NAND2X0 U10107 ( .IN1(n10073), .IN2(n10103), .QN(n10099) );
  NAND2X0 U10108 ( .IN1(n10094), .IN2(n10104), .QN(n10103) );
  NAND2X0 U10109 ( .IN1(n10105), .IN2(n10085), .QN(n10104) );
  NAND2X0 U10110 ( .IN1(n10106), .IN2(n10044), .QN(n10062) );
  AND4X1 U10111 ( .IN1(n10107), .IN2(n10108), .IN3(n10109), .IN4(n10110), .Q(
        n10044) );
  NAND2X0 U10112 ( .IN1(n10111), .IN2(n10068), .QN(n10110) );
  NAND2X0 U10113 ( .IN1(n10112), .IN2(n10113), .QN(n10111) );
  NAND2X0 U10114 ( .IN1(n10091), .IN2(n10105), .QN(n10113) );
  INVX0 U10115 ( .INP(n10071), .ZN(n10091) );
  NAND2X0 U10116 ( .IN1(n10073), .IN2(n10114), .QN(n10112) );
  NAND2X0 U10117 ( .IN1(n10115), .IN2(n10116), .QN(n10114) );
  NAND2X0 U10118 ( .IN1(n10117), .IN2(n10085), .QN(n10116) );
  NAND2X0 U10119 ( .IN1(n10118), .IN2(n10119), .QN(n10117) );
  NAND3X0 U10120 ( .IN1(n10090), .IN2(n10079), .IN3(n10094), .QN(n10119) );
  NAND2X0 U10121 ( .IN1(n10071), .IN2(n10088), .QN(n10118) );
  NAND2X0 U10122 ( .IN1(n10097), .IN2(n10102), .QN(n10115) );
  NAND2X0 U10123 ( .IN1(n10081), .IN2(n10120), .QN(n10109) );
  NAND2X0 U10124 ( .IN1(n10121), .IN2(n10122), .QN(n10120) );
  NAND3X0 U10125 ( .IN1(n10102), .IN2(n10079), .IN3(n10074), .QN(n10122) );
  NAND2X0 U10126 ( .IN1(n10123), .IN2(n10089), .QN(n10121) );
  NAND3X0 U10127 ( .IN1(n10124), .IN2(n10125), .IN3(n10126), .QN(n10123) );
  NAND3X0 U10128 ( .IN1(n10097), .IN2(n10090), .IN3(n10094), .QN(n10126) );
  INVX0 U10129 ( .INP(n10079), .ZN(n10097) );
  NAND2X0 U10130 ( .IN1(n10074), .IN2(n10088), .QN(n10125) );
  NAND3X0 U10131 ( .IN1(n10105), .IN2(n10071), .IN3(n10085), .QN(n10124) );
  NAND3X0 U10132 ( .IN1(n10127), .IN2(n10128), .IN3(n10129), .QN(n10071) );
  NAND2X0 U10133 ( .IN1(test_so63), .IN2(g1775), .QN(n10129) );
  NAND2X0 U10134 ( .IN1(g1718), .IN2(g1705), .QN(n10128) );
  NAND2X0 U10135 ( .IN1(g5738), .IN2(g1777), .QN(n10127) );
  NAND3X0 U10136 ( .IN1(n10079), .IN2(n10072), .IN3(n10095), .QN(n10108) );
  NOR2X0 U10137 ( .IN1(n10074), .IN2(n10073), .QN(n10095) );
  NAND3X0 U10138 ( .IN1(n10130), .IN2(n10131), .IN3(n10132), .QN(n10079) );
  NAND2X0 U10139 ( .IN1(test_so63), .IN2(g1760), .QN(n10132) );
  NAND2X0 U10140 ( .IN1(g1718), .IN2(g1764), .QN(n10131) );
  NAND2X0 U10141 ( .IN1(g5738), .IN2(g1762), .QN(n10130) );
  NAND3X0 U10142 ( .IN1(n10074), .IN2(n10096), .IN3(n10073), .QN(n10107) );
  INVX0 U10143 ( .INP(n10089), .ZN(n10073) );
  NAND3X0 U10144 ( .IN1(n10133), .IN2(n10134), .IN3(n10135), .QN(n10089) );
  NAND2X0 U10145 ( .IN1(test_so63), .IN2(g1730), .QN(n10135) );
  NAND2X0 U10146 ( .IN1(g1718), .IN2(g1734), .QN(n10134) );
  NAND2X0 U10147 ( .IN1(g5738), .IN2(g1732), .QN(n10133) );
  INVX0 U10148 ( .INP(n10085), .ZN(n10074) );
  NAND3X0 U10149 ( .IN1(n10136), .IN2(n10137), .IN3(n10138), .QN(n10085) );
  NAND2X0 U10150 ( .IN1(test_so63), .IN2(g1745), .QN(n10138) );
  NAND2X0 U10151 ( .IN1(g1718), .IN2(g1749), .QN(n10137) );
  NAND2X0 U10152 ( .IN1(g5738), .IN2(g1747), .QN(n10136) );
  INVX0 U10153 ( .INP(n10139), .ZN(n10106) );
  NAND2X0 U10154 ( .IN1(n10047), .IN2(n10139), .QN(n10043) );
  NAND2X0 U10155 ( .IN1(n4296), .IN2(g1985), .QN(n10058) );
  NAND2X0 U10156 ( .IN1(n10140), .IN2(n10141), .QN(g28351) );
  NAND2X0 U10157 ( .IN1(n4371), .IN2(g1300), .QN(n10141) );
  NAND2X0 U10158 ( .IN1(n9957), .IN2(n10142), .QN(n10140) );
  NAND2X0 U10159 ( .IN1(n10143), .IN2(n10144), .QN(n9957) );
  NAND2X0 U10160 ( .IN1(n9947), .IN2(n8278), .QN(n10144) );
  NAND4X0 U10161 ( .IN1(n10145), .IN2(n10146), .IN3(n10147), .IN4(n9946), .QN(
        n10143) );
  NAND2X0 U10162 ( .IN1(n10148), .IN2(n10149), .QN(n10145) );
  INVX0 U10163 ( .INP(n10150), .ZN(n10148) );
  NAND2X0 U10164 ( .IN1(n10151), .IN2(n10152), .QN(g28350) );
  NAND2X0 U10165 ( .IN1(n4316), .IN2(g1294), .QN(n10152) );
  NAND2X0 U10166 ( .IN1(n10054), .IN2(g6944), .QN(n10151) );
  NAND2X0 U10167 ( .IN1(n10153), .IN2(n10154), .QN(g28349) );
  NAND2X0 U10168 ( .IN1(n4372), .IN2(g617), .QN(n10154) );
  NAND2X0 U10169 ( .IN1(n10057), .IN2(g6642), .QN(n10153) );
  NAND2X0 U10170 ( .IN1(n10155), .IN2(n10156), .QN(g28348) );
  NAND2X0 U10171 ( .IN1(n4313), .IN2(g611), .QN(n10156) );
  NAND2X0 U10172 ( .IN1(n10157), .IN2(g550), .QN(n10155) );
  NAND2X0 U10173 ( .IN1(n10158), .IN2(n10159), .QN(g28346) );
  NAND2X0 U10174 ( .IN1(g6750), .IN2(n10054), .QN(n10159) );
  NAND2X0 U10175 ( .IN1(n10160), .IN2(n10161), .QN(n10054) );
  NAND2X0 U10176 ( .IN1(n9947), .IN2(n8285), .QN(n10161) );
  NAND4X0 U10177 ( .IN1(n10146), .IN2(n10162), .IN3(n10149), .IN4(n9946), .QN(
        n10160) );
  AND4X1 U10178 ( .IN1(n10163), .IN2(n10164), .IN3(n10165), .IN4(n10166), .Q(
        n10149) );
  NAND2X0 U10179 ( .IN1(n10167), .IN2(n10168), .QN(n10166) );
  NAND2X0 U10180 ( .IN1(n10169), .IN2(n10170), .QN(n10167) );
  NAND3X0 U10181 ( .IN1(n10171), .IN2(n10172), .IN3(n10173), .QN(n10170) );
  NAND2X0 U10182 ( .IN1(n10174), .IN2(n10175), .QN(n10169) );
  NAND2X0 U10183 ( .IN1(n10176), .IN2(n10177), .QN(n10175) );
  NAND2X0 U10184 ( .IN1(n10178), .IN2(n10179), .QN(n10177) );
  INVX0 U10185 ( .INP(n10180), .ZN(n10176) );
  NAND2X0 U10186 ( .IN1(n10181), .IN2(n10182), .QN(n10165) );
  NAND2X0 U10187 ( .IN1(n10183), .IN2(n10184), .QN(n10182) );
  NAND3X0 U10188 ( .IN1(n10185), .IN2(n10179), .IN3(n10180), .QN(n10184) );
  NAND2X0 U10189 ( .IN1(n10186), .IN2(n10187), .QN(n10180) );
  NAND2X0 U10190 ( .IN1(n10188), .IN2(n10189), .QN(n10187) );
  NAND2X0 U10191 ( .IN1(n10190), .IN2(n10173), .QN(n10186) );
  NAND2X0 U10192 ( .IN1(n10191), .IN2(n10178), .QN(n10183) );
  NAND2X0 U10193 ( .IN1(n10192), .IN2(n10193), .QN(n10178) );
  NAND2X0 U10194 ( .IN1(n10194), .IN2(n10189), .QN(n10193) );
  NAND3X0 U10195 ( .IN1(n10195), .IN2(n10171), .IN3(n10196), .QN(n10164) );
  NAND2X0 U10196 ( .IN1(n10197), .IN2(n10198), .QN(n10163) );
  NAND3X0 U10197 ( .IN1(n10199), .IN2(n10200), .IN3(n10201), .QN(n10198) );
  NAND2X0 U10198 ( .IN1(n10195), .IN2(n10202), .QN(n10201) );
  NAND2X0 U10199 ( .IN1(n10196), .IN2(n10189), .QN(n10200) );
  NAND2X0 U10200 ( .IN1(n10173), .IN2(n10203), .QN(n10199) );
  NAND2X0 U10201 ( .IN1(n10194), .IN2(n10204), .QN(n10203) );
  NAND2X0 U10202 ( .IN1(n10205), .IN2(n10185), .QN(n10204) );
  NAND2X0 U10203 ( .IN1(n10206), .IN2(n10147), .QN(n10162) );
  AND4X1 U10204 ( .IN1(n10207), .IN2(n10208), .IN3(n10209), .IN4(n10210), .Q(
        n10147) );
  NAND2X0 U10205 ( .IN1(n10211), .IN2(n10168), .QN(n10210) );
  NAND2X0 U10206 ( .IN1(n10212), .IN2(n10213), .QN(n10211) );
  NAND2X0 U10207 ( .IN1(n10191), .IN2(n10205), .QN(n10213) );
  INVX0 U10208 ( .INP(n10171), .ZN(n10191) );
  NAND2X0 U10209 ( .IN1(n10173), .IN2(n10214), .QN(n10212) );
  NAND2X0 U10210 ( .IN1(n10215), .IN2(n10216), .QN(n10214) );
  NAND2X0 U10211 ( .IN1(n10217), .IN2(n10185), .QN(n10216) );
  NAND2X0 U10212 ( .IN1(n10218), .IN2(n10219), .QN(n10217) );
  NAND3X0 U10213 ( .IN1(n10190), .IN2(n10179), .IN3(n10194), .QN(n10219) );
  NAND2X0 U10214 ( .IN1(n10171), .IN2(n10188), .QN(n10218) );
  NAND2X0 U10215 ( .IN1(n10197), .IN2(n10202), .QN(n10215) );
  NAND2X0 U10216 ( .IN1(n10181), .IN2(n10220), .QN(n10209) );
  NAND2X0 U10217 ( .IN1(n10221), .IN2(n10222), .QN(n10220) );
  NAND3X0 U10218 ( .IN1(n10202), .IN2(n10179), .IN3(n10174), .QN(n10222) );
  NAND2X0 U10219 ( .IN1(n10223), .IN2(n10189), .QN(n10221) );
  NAND3X0 U10220 ( .IN1(n10224), .IN2(n10225), .IN3(n10226), .QN(n10223) );
  NAND3X0 U10221 ( .IN1(n10197), .IN2(n10190), .IN3(n10194), .QN(n10226) );
  INVX0 U10222 ( .INP(n10179), .ZN(n10197) );
  NAND2X0 U10223 ( .IN1(n10174), .IN2(n10188), .QN(n10225) );
  NAND3X0 U10224 ( .IN1(n10205), .IN2(n10171), .IN3(n10185), .QN(n10224) );
  NAND3X0 U10225 ( .IN1(n10227), .IN2(n10228), .IN3(n10229), .QN(n10171) );
  NAND2X0 U10226 ( .IN1(g5686), .IN2(g1083), .QN(n10229) );
  NAND2X0 U10227 ( .IN1(g5657), .IN2(g1081), .QN(n10228) );
  NAND2X0 U10228 ( .IN1(g1024), .IN2(g1011), .QN(n10227) );
  NAND3X0 U10229 ( .IN1(n10179), .IN2(n10172), .IN3(n10195), .QN(n10208) );
  NOR2X0 U10230 ( .IN1(n10174), .IN2(n10173), .QN(n10195) );
  NAND3X0 U10231 ( .IN1(n10230), .IN2(n10231), .IN3(n10232), .QN(n10179) );
  NAND2X0 U10232 ( .IN1(g5686), .IN2(g1068), .QN(n10232) );
  NAND2X0 U10233 ( .IN1(g5657), .IN2(g1066), .QN(n10231) );
  NAND2X0 U10234 ( .IN1(g1024), .IN2(g1070), .QN(n10230) );
  NAND3X0 U10235 ( .IN1(n10174), .IN2(n10196), .IN3(n10173), .QN(n10207) );
  INVX0 U10236 ( .INP(n10189), .ZN(n10173) );
  NAND3X0 U10237 ( .IN1(n10233), .IN2(n10234), .IN3(n10235), .QN(n10189) );
  NAND2X0 U10238 ( .IN1(g5686), .IN2(g1038), .QN(n10235) );
  NAND2X0 U10239 ( .IN1(g5657), .IN2(g1036), .QN(n10234) );
  NAND2X0 U10240 ( .IN1(g1024), .IN2(g1040), .QN(n10233) );
  INVX0 U10241 ( .INP(n10185), .ZN(n10174) );
  NAND3X0 U10242 ( .IN1(n10236), .IN2(n10237), .IN3(n10238), .QN(n10185) );
  NAND2X0 U10243 ( .IN1(g5686), .IN2(g1053), .QN(n10238) );
  NAND2X0 U10244 ( .IN1(g5657), .IN2(g1051), .QN(n10237) );
  NAND2X0 U10245 ( .IN1(g1024), .IN2(g1055), .QN(n10236) );
  INVX0 U10246 ( .INP(n10239), .ZN(n10206) );
  NAND2X0 U10247 ( .IN1(n10150), .IN2(n10239), .QN(n10146) );
  NAND2X0 U10248 ( .IN1(n4371), .IN2(g1291), .QN(n10158) );
  NAND2X0 U10249 ( .IN1(n10240), .IN2(n10241), .QN(g28345) );
  NAND2X0 U10250 ( .IN1(n4298), .IN2(g614), .QN(n10241) );
  NAND2X0 U10251 ( .IN1(n10057), .IN2(n10242), .QN(n10240) );
  NAND2X0 U10252 ( .IN1(n10243), .IN2(n10244), .QN(n10057) );
  NAND2X0 U10253 ( .IN1(n9947), .IN2(n7844), .QN(n10244) );
  NAND4X0 U10254 ( .IN1(n10245), .IN2(n10246), .IN3(n10247), .IN4(n9946), .QN(
        n10243) );
  NAND2X0 U10255 ( .IN1(n10248), .IN2(n10249), .QN(n10245) );
  INVX0 U10256 ( .INP(n10250), .ZN(n10248) );
  NAND2X0 U10257 ( .IN1(n10251), .IN2(n10252), .QN(g28344) );
  NAND2X0 U10258 ( .IN1(n4372), .IN2(g608), .QN(n10252) );
  NAND2X0 U10259 ( .IN1(n10157), .IN2(g6642), .QN(n10251) );
  NAND2X0 U10260 ( .IN1(n10253), .IN2(n10254), .QN(g28342) );
  NAND2X0 U10261 ( .IN1(g6485), .IN2(n10157), .QN(n10254) );
  NAND2X0 U10262 ( .IN1(n10255), .IN2(n10256), .QN(n10157) );
  NAND2X0 U10263 ( .IN1(n9947), .IN2(n7851), .QN(n10256) );
  NAND4X0 U10264 ( .IN1(n10246), .IN2(n10257), .IN3(n10249), .IN4(n9946), .QN(
        n10255) );
  INVX0 U10265 ( .INP(n9947), .ZN(n9946) );
  AND4X1 U10266 ( .IN1(n10258), .IN2(n10259), .IN3(n10260), .IN4(n10261), .Q(
        n10249) );
  NAND2X0 U10267 ( .IN1(n10262), .IN2(n10263), .QN(n10261) );
  NAND2X0 U10268 ( .IN1(n10264), .IN2(n10265), .QN(n10262) );
  NAND3X0 U10269 ( .IN1(n10266), .IN2(n10267), .IN3(n10268), .QN(n10265) );
  NAND2X0 U10270 ( .IN1(n10269), .IN2(n10270), .QN(n10264) );
  NAND2X0 U10271 ( .IN1(n10271), .IN2(n10272), .QN(n10270) );
  NAND2X0 U10272 ( .IN1(n10273), .IN2(n10274), .QN(n10272) );
  INVX0 U10273 ( .INP(n10275), .ZN(n10271) );
  NAND2X0 U10274 ( .IN1(n10276), .IN2(n10277), .QN(n10260) );
  NAND2X0 U10275 ( .IN1(n10278), .IN2(n10279), .QN(n10277) );
  NAND3X0 U10276 ( .IN1(n10280), .IN2(n10274), .IN3(n10275), .QN(n10279) );
  NAND2X0 U10277 ( .IN1(n10281), .IN2(n10282), .QN(n10275) );
  NAND2X0 U10278 ( .IN1(n10283), .IN2(n10284), .QN(n10282) );
  NAND2X0 U10279 ( .IN1(n10285), .IN2(n10268), .QN(n10281) );
  NAND2X0 U10280 ( .IN1(n10286), .IN2(n10273), .QN(n10278) );
  NAND2X0 U10281 ( .IN1(n10287), .IN2(n10288), .QN(n10273) );
  NAND2X0 U10282 ( .IN1(n10289), .IN2(n10284), .QN(n10288) );
  NAND3X0 U10283 ( .IN1(n10290), .IN2(n10266), .IN3(n10291), .QN(n10259) );
  NAND2X0 U10284 ( .IN1(n10292), .IN2(n10293), .QN(n10258) );
  NAND3X0 U10285 ( .IN1(n10294), .IN2(n10295), .IN3(n10296), .QN(n10293) );
  NAND2X0 U10286 ( .IN1(n10290), .IN2(n10297), .QN(n10296) );
  NAND2X0 U10287 ( .IN1(n10291), .IN2(n10284), .QN(n10295) );
  NAND2X0 U10288 ( .IN1(n10268), .IN2(n10298), .QN(n10294) );
  NAND2X0 U10289 ( .IN1(n10289), .IN2(n10299), .QN(n10298) );
  NAND2X0 U10290 ( .IN1(n10300), .IN2(n10280), .QN(n10299) );
  NAND2X0 U10291 ( .IN1(n10301), .IN2(n10247), .QN(n10257) );
  AND4X1 U10292 ( .IN1(n10302), .IN2(n10303), .IN3(n10304), .IN4(n10305), .Q(
        n10247) );
  NAND2X0 U10293 ( .IN1(n10306), .IN2(n10263), .QN(n10305) );
  NAND2X0 U10294 ( .IN1(n10307), .IN2(n10308), .QN(n10306) );
  NAND2X0 U10295 ( .IN1(n10286), .IN2(n10300), .QN(n10308) );
  INVX0 U10296 ( .INP(n10266), .ZN(n10286) );
  NAND2X0 U10297 ( .IN1(n10268), .IN2(n10309), .QN(n10307) );
  NAND2X0 U10298 ( .IN1(n10310), .IN2(n10311), .QN(n10309) );
  NAND2X0 U10299 ( .IN1(n10312), .IN2(n10280), .QN(n10311) );
  NAND2X0 U10300 ( .IN1(n10313), .IN2(n10314), .QN(n10312) );
  NAND3X0 U10301 ( .IN1(n10285), .IN2(n10274), .IN3(n10289), .QN(n10314) );
  NAND2X0 U10302 ( .IN1(n10266), .IN2(n10283), .QN(n10313) );
  NAND2X0 U10303 ( .IN1(n10292), .IN2(n10297), .QN(n10310) );
  NAND2X0 U10304 ( .IN1(n10276), .IN2(n10315), .QN(n10304) );
  NAND2X0 U10305 ( .IN1(n10316), .IN2(n10317), .QN(n10315) );
  NAND3X0 U10306 ( .IN1(n10297), .IN2(n10274), .IN3(n10269), .QN(n10317) );
  NAND2X0 U10307 ( .IN1(n10318), .IN2(n10284), .QN(n10316) );
  NAND3X0 U10308 ( .IN1(n10319), .IN2(n10320), .IN3(n10321), .QN(n10318) );
  NAND3X0 U10309 ( .IN1(n10292), .IN2(n10285), .IN3(n10289), .QN(n10321) );
  INVX0 U10310 ( .INP(n10274), .ZN(n10292) );
  NAND2X0 U10311 ( .IN1(n10269), .IN2(n10283), .QN(n10320) );
  NAND3X0 U10312 ( .IN1(n10300), .IN2(n10266), .IN3(n10280), .QN(n10319) );
  NAND3X0 U10313 ( .IN1(n10322), .IN2(n10323), .IN3(n10324), .QN(n10266) );
  NAND2X0 U10314 ( .IN1(g5648), .IN2(g396), .QN(n10324) );
  NAND2X0 U10315 ( .IN1(g5629), .IN2(g394), .QN(n10323) );
  NAND2X0 U10316 ( .IN1(g337), .IN2(g324), .QN(n10322) );
  NAND3X0 U10317 ( .IN1(n10274), .IN2(n10267), .IN3(n10290), .QN(n10303) );
  NOR2X0 U10318 ( .IN1(n10269), .IN2(n10268), .QN(n10290) );
  NAND3X0 U10319 ( .IN1(n10325), .IN2(n10326), .IN3(n10327), .QN(n10274) );
  NAND2X0 U10320 ( .IN1(g5648), .IN2(g381), .QN(n10327) );
  NAND2X0 U10321 ( .IN1(g5629), .IN2(g379), .QN(n10326) );
  NAND2X0 U10322 ( .IN1(g337), .IN2(g383), .QN(n10325) );
  NAND3X0 U10323 ( .IN1(n10269), .IN2(n10291), .IN3(n10268), .QN(n10302) );
  INVX0 U10324 ( .INP(n10284), .ZN(n10268) );
  NAND3X0 U10325 ( .IN1(n10328), .IN2(n10329), .IN3(n10330), .QN(n10284) );
  NAND2X0 U10326 ( .IN1(g5648), .IN2(g351), .QN(n10330) );
  NAND2X0 U10327 ( .IN1(g5629), .IN2(g349), .QN(n10329) );
  NAND2X0 U10328 ( .IN1(g337), .IN2(g353), .QN(n10328) );
  INVX0 U10329 ( .INP(n10280), .ZN(n10269) );
  NAND3X0 U10330 ( .IN1(n10331), .IN2(n10332), .IN3(n10333), .QN(n10280) );
  NAND2X0 U10331 ( .IN1(g5648), .IN2(g366), .QN(n10333) );
  NAND2X0 U10332 ( .IN1(g5629), .IN2(g364), .QN(n10332) );
  NAND2X0 U10333 ( .IN1(g337), .IN2(g368), .QN(n10331) );
  INVX0 U10334 ( .INP(n10334), .ZN(n10301) );
  NAND2X0 U10335 ( .IN1(n10250), .IN2(n10334), .QN(n10246) );
  NAND2X0 U10336 ( .IN1(n4298), .IN2(g605), .QN(n10253) );
  NOR2X0 U10337 ( .IN1(n10335), .IN2(n10336), .QN(g28328) );
  XOR2X1 U10338 ( .IN1(n4415), .IN2(n10337), .Q(n10336) );
  NOR2X0 U10339 ( .IN1(n4393), .IN2(n10338), .QN(n10337) );
  NOR2X0 U10340 ( .IN1(n10339), .IN2(n10340), .QN(g28325) );
  XNOR2X1 U10341 ( .IN1(n4416), .IN2(n10341), .Q(n10340) );
  NAND2X0 U10342 ( .IN1(test_so70), .IN2(n10342), .QN(n10341) );
  NOR2X0 U10343 ( .IN1(n10343), .IN2(n10344), .QN(g28321) );
  XNOR2X1 U10344 ( .IN1(n4417), .IN2(n10345), .Q(n10344) );
  NAND2X0 U10345 ( .IN1(n10346), .IN2(g1372), .QN(n10345) );
  NOR2X0 U10346 ( .IN1(n9912), .IN2(n10347), .QN(g28199) );
  XNOR2X1 U10347 ( .IN1(n4396), .IN2(n9915), .Q(n10347) );
  AND3X1 U10348 ( .IN1(n9736), .IN2(n3160), .IN3(n10348), .Q(g28148) );
  NAND2X0 U10349 ( .IN1(n6972), .IN2(n10349), .QN(n10348) );
  OR2X1 U10350 ( .IN1(n10349), .IN2(n6972), .Q(n3160) );
  INVX0 U10351 ( .INP(n3424), .ZN(n10349) );
  AND3X1 U10352 ( .IN1(n9739), .IN2(n3164), .IN3(n10350), .Q(g28147) );
  NAND2X0 U10353 ( .IN1(n6973), .IN2(n10351), .QN(n10350) );
  OR2X1 U10354 ( .IN1(n10351), .IN2(n6973), .Q(n3164) );
  INVX0 U10355 ( .INP(n3427), .ZN(n10351) );
  NOR3X0 U10356 ( .IN1(n10352), .IN2(n9322), .IN3(n9919), .QN(g28146) );
  INVX0 U10357 ( .INP(n3168), .ZN(n9919) );
  NAND2X0 U10358 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NOR2X0 U10359 ( .IN1(n3430), .IN2(g758), .QN(n10352) );
  AND3X1 U10360 ( .IN1(n9743), .IN2(n3172), .IN3(n10353), .Q(g28145) );
  NAND2X0 U10361 ( .IN1(n6975), .IN2(n10354), .QN(n10353) );
  OR2X1 U10362 ( .IN1(n10354), .IN2(n6975), .Q(n3172) );
  INVX0 U10363 ( .INP(n3433), .ZN(n10354) );
  NAND2X0 U10364 ( .IN1(n10355), .IN2(n10356), .QN(g27771) );
  NAND2X0 U10365 ( .IN1(test_so81), .IN2(n10357), .QN(n10356) );
  NAND2X0 U10366 ( .IN1(n10358), .IN2(n8841), .QN(n10357) );
  NAND2X0 U10367 ( .IN1(n10359), .IN2(n8841), .QN(n10355) );
  NAND2X0 U10368 ( .IN1(n10360), .IN2(n10361), .QN(g27769) );
  NAND2X0 U10369 ( .IN1(n10362), .IN2(g2524), .QN(n10361) );
  NAND2X0 U10370 ( .IN1(n10358), .IN2(n8449), .QN(n10362) );
  NAND2X0 U10371 ( .IN1(n10359), .IN2(n8449), .QN(n10360) );
  NAND2X0 U10372 ( .IN1(n10363), .IN2(n10364), .QN(g27768) );
  NAND2X0 U10373 ( .IN1(n10365), .IN2(g1828), .QN(n10364) );
  NAND2X0 U10374 ( .IN1(n10366), .IN2(n8453), .QN(n10365) );
  NAND2X0 U10375 ( .IN1(n10367), .IN2(n8453), .QN(n10363) );
  NAND2X0 U10376 ( .IN1(n10368), .IN2(n10369), .QN(g27767) );
  NAND2X0 U10377 ( .IN1(n10370), .IN2(g2523), .QN(n10369) );
  NAND2X0 U10378 ( .IN1(n10358), .IN2(n8456), .QN(n10370) );
  AND4X1 U10379 ( .IN1(n10371), .IN2(test_so79), .IN3(n10372), .IN4(n10373), 
        .Q(n10358) );
  NAND2X0 U10380 ( .IN1(n10359), .IN2(n8456), .QN(n10368) );
  AND3X1 U10381 ( .IN1(n10374), .IN2(n10375), .IN3(test_so79), .Q(n10359) );
  NAND2X0 U10382 ( .IN1(n10376), .IN2(n10377), .QN(n10375) );
  NAND2X0 U10383 ( .IN1(n10378), .IN2(n10379), .QN(n10377) );
  NAND2X0 U10384 ( .IN1(n10380), .IN2(n10381), .QN(n10374) );
  NAND2X0 U10385 ( .IN1(n10382), .IN2(n10383), .QN(n10380) );
  NAND2X0 U10386 ( .IN1(n10384), .IN2(n10385), .QN(g27766) );
  NAND2X0 U10387 ( .IN1(n10386), .IN2(g1830), .QN(n10385) );
  NAND2X0 U10388 ( .IN1(n10366), .IN2(n8459), .QN(n10386) );
  NAND2X0 U10389 ( .IN1(n10367), .IN2(n8459), .QN(n10384) );
  NAND2X0 U10390 ( .IN1(n10387), .IN2(n10388), .QN(g27765) );
  NAND2X0 U10391 ( .IN1(n10389), .IN2(g1134), .QN(n10388) );
  NAND2X0 U10392 ( .IN1(n10390), .IN2(g1088), .QN(n10389) );
  NAND2X0 U10393 ( .IN1(n10391), .IN2(g1088), .QN(n10387) );
  NAND2X0 U10394 ( .IN1(n10392), .IN2(n10393), .QN(g27764) );
  NAND2X0 U10395 ( .IN1(n10394), .IN2(g1829), .QN(n10393) );
  NAND2X0 U10396 ( .IN1(n10366), .IN2(n8494), .QN(n10394) );
  AND4X1 U10397 ( .IN1(n10395), .IN2(n10396), .IN3(n10397), .IN4(g1690), .Q(
        n10366) );
  NAND2X0 U10398 ( .IN1(n10367), .IN2(n8494), .QN(n10392) );
  AND3X1 U10399 ( .IN1(n10398), .IN2(n10399), .IN3(g1690), .Q(n10367) );
  NAND2X0 U10400 ( .IN1(n10400), .IN2(n10401), .QN(n10399) );
  NAND2X0 U10401 ( .IN1(n10402), .IN2(n10403), .QN(n10401) );
  NAND2X0 U10402 ( .IN1(n10404), .IN2(n10405), .QN(n10398) );
  NAND2X0 U10403 ( .IN1(n10406), .IN2(n10407), .QN(n10404) );
  NAND2X0 U10404 ( .IN1(n10408), .IN2(n10409), .QN(g27763) );
  NAND2X0 U10405 ( .IN1(n10410), .IN2(g1136), .QN(n10409) );
  NAND2X0 U10406 ( .IN1(n10390), .IN2(g6712), .QN(n10410) );
  NAND2X0 U10407 ( .IN1(n10391), .IN2(g6712), .QN(n10408) );
  NAND2X0 U10408 ( .IN1(n10411), .IN2(n10412), .QN(g27762) );
  NAND2X0 U10409 ( .IN1(n10413), .IN2(g447), .QN(n10412) );
  NAND2X0 U10410 ( .IN1(n10414), .IN2(n8500), .QN(n10413) );
  NAND2X0 U10411 ( .IN1(n10415), .IN2(n8500), .QN(n10411) );
  NAND2X0 U10412 ( .IN1(n10416), .IN2(n10417), .QN(g27761) );
  NAND2X0 U10413 ( .IN1(n10418), .IN2(g1135), .QN(n10417) );
  NAND2X0 U10414 ( .IN1(n10390), .IN2(g5472), .QN(n10418) );
  AND4X1 U10415 ( .IN1(n10419), .IN2(n10420), .IN3(n10421), .IN4(g996), .Q(
        n10390) );
  NAND2X0 U10416 ( .IN1(n10391), .IN2(g5472), .QN(n10416) );
  AND3X1 U10417 ( .IN1(n10422), .IN2(n10423), .IN3(g996), .Q(n10391) );
  NAND2X0 U10418 ( .IN1(n10424), .IN2(n10425), .QN(n10423) );
  NAND2X0 U10419 ( .IN1(n10426), .IN2(n10427), .QN(n10425) );
  NAND2X0 U10420 ( .IN1(n10428), .IN2(n10429), .QN(n10422) );
  NAND2X0 U10421 ( .IN1(n10430), .IN2(n10431), .QN(n10428) );
  NAND2X0 U10422 ( .IN1(n10432), .IN2(n10433), .QN(g27760) );
  NAND2X0 U10423 ( .IN1(n10434), .IN2(g449), .QN(n10433) );
  NAND2X0 U10424 ( .IN1(n10414), .IN2(n8861), .QN(n10434) );
  NAND2X0 U10425 ( .IN1(n10415), .IN2(n8861), .QN(n10432) );
  NAND2X0 U10426 ( .IN1(n10435), .IN2(n10436), .QN(g27759) );
  NAND2X0 U10427 ( .IN1(n10437), .IN2(g448), .QN(n10436) );
  NAND2X0 U10428 ( .IN1(n10414), .IN2(n8537), .QN(n10437) );
  AND4X1 U10429 ( .IN1(n10438), .IN2(n10439), .IN3(n10440), .IN4(g309), .Q(
        n10414) );
  NAND2X0 U10430 ( .IN1(n10415), .IN2(n8537), .QN(n10435) );
  AND3X1 U10431 ( .IN1(n10441), .IN2(n10442), .IN3(g309), .Q(n10415) );
  NAND2X0 U10432 ( .IN1(n10443), .IN2(n10444), .QN(n10442) );
  NAND2X0 U10433 ( .IN1(n10445), .IN2(n10446), .QN(n10444) );
  NAND2X0 U10434 ( .IN1(n10447), .IN2(n10448), .QN(n10441) );
  NAND2X0 U10435 ( .IN1(n10449), .IN2(n10450), .QN(n10447) );
  NOR2X0 U10436 ( .IN1(n10335), .IN2(n10451), .QN(g27724) );
  XNOR2X1 U10437 ( .IN1(n4393), .IN2(n10338), .Q(n10451) );
  NOR2X0 U10438 ( .IN1(n10339), .IN2(n10452), .QN(g27722) );
  XOR2X1 U10439 ( .IN1(n7272), .IN2(n10342), .Q(n10452) );
  NOR2X0 U10440 ( .IN1(n10343), .IN2(n10453), .QN(g27718) );
  XOR2X1 U10441 ( .IN1(n4395), .IN2(n10346), .Q(n10453) );
  NOR3X0 U10442 ( .IN1(n10454), .IN2(n10339), .IN3(n10342), .QN(g27682) );
  NOR3X0 U10443 ( .IN1(n4468), .IN2(n4473), .IN3(n10455), .QN(n10342) );
  NOR2X0 U10444 ( .IN1(n10456), .IN2(g2059), .QN(n10454) );
  NOR2X0 U10445 ( .IN1(n4468), .IN2(n10455), .QN(n10456) );
  NOR3X0 U10446 ( .IN1(n10457), .IN2(n10343), .IN3(n10346), .QN(g27678) );
  NOR3X0 U10447 ( .IN1(n4469), .IN2(n4475), .IN3(n10458), .QN(n10346) );
  NOR2X0 U10448 ( .IN1(n10459), .IN2(g1365), .QN(n10457) );
  NOR2X0 U10449 ( .IN1(n4469), .IN2(n10458), .QN(n10459) );
  AND3X1 U10450 ( .IN1(n10460), .IN2(n10461), .IN3(n9915), .Q(g27672) );
  NAND3X0 U10451 ( .IN1(n10462), .IN2(g679), .IN3(test_so28), .QN(n9915) );
  OR2X1 U10452 ( .IN1(n10463), .IN2(g679), .Q(n10460) );
  NOR2X0 U10453 ( .IN1(n10464), .IN2(n7270), .QN(n10463) );
  NOR2X0 U10454 ( .IN1(n9318), .IN2(n10465), .QN(g27621) );
  XNOR2X1 U10455 ( .IN1(n4522), .IN2(n6980), .Q(n10465) );
  NOR2X0 U10456 ( .IN1(n9320), .IN2(n10466), .QN(g27612) );
  XNOR2X1 U10457 ( .IN1(n4523), .IN2(n6984), .Q(n10466) );
  NOR2X0 U10458 ( .IN1(n9322), .IN2(n10467), .QN(g27603) );
  XOR2X1 U10459 ( .IN1(n6988), .IN2(n10468), .Q(n10467) );
  NOR2X0 U10460 ( .IN1(n9324), .IN2(n10469), .QN(g27594) );
  XNOR2X1 U10461 ( .IN1(n4521), .IN2(n6992), .Q(n10469) );
  NAND4X0 U10462 ( .IN1(n10470), .IN2(n10471), .IN3(n3700), .IN4(n10472), .QN(
        g27380) );
  AND4X1 U10463 ( .IN1(n10473), .IN2(n10474), .IN3(n10475), .IN4(n10476), .Q(
        n10472) );
  NAND4X0 U10464 ( .IN1(n10477), .IN2(n10478), .IN3(n10479), .IN4(n10480), 
        .QN(n10475) );
  NAND2X0 U10465 ( .IN1(n10481), .IN2(n8082), .QN(n10480) );
  NAND2X0 U10466 ( .IN1(n10482), .IN2(n8081), .QN(n10479) );
  NAND2X0 U10467 ( .IN1(n10483), .IN2(n10484), .QN(n10474) );
  NAND2X0 U10468 ( .IN1(n10485), .IN2(n10486), .QN(n10484) );
  NAND3X0 U10469 ( .IN1(n10477), .IN2(g3188), .IN3(n4384), .QN(n10486) );
  INVX0 U10470 ( .INP(n3705), .ZN(n10485) );
  NAND2X0 U10471 ( .IN1(n10487), .IN2(g3151), .QN(n10473) );
  OR2X1 U10472 ( .IN1(n10488), .IN2(n13232), .Q(n10471) );
  NAND2X0 U10473 ( .IN1(n6707), .IN2(n10489), .QN(n10470) );
  NAND2X0 U10474 ( .IN1(n10490), .IN2(n10491), .QN(g27354) );
  OR2X1 U10475 ( .IN1(n10492), .IN2(n6625), .Q(n10491) );
  NAND2X0 U10476 ( .IN1(n10492), .IN2(n10493), .QN(n10490) );
  NAND2X0 U10477 ( .IN1(n10494), .IN2(n10495), .QN(g27348) );
  NAND2X0 U10478 ( .IN1(n10496), .IN2(n10493), .QN(n10495) );
  OR2X1 U10479 ( .IN1(n10496), .IN2(n6626), .Q(n10494) );
  NAND2X0 U10480 ( .IN1(n10497), .IN2(n10498), .QN(g27347) );
  OR2X1 U10481 ( .IN1(n10492), .IN2(n6441), .Q(n10498) );
  NAND2X0 U10482 ( .IN1(n10499), .IN2(n10492), .QN(n10497) );
  NAND2X0 U10483 ( .IN1(n10500), .IN2(n10501), .QN(g27346) );
  OR2X1 U10484 ( .IN1(n10502), .IN2(n6627), .Q(n10501) );
  NAND2X0 U10485 ( .IN1(n10502), .IN2(n10503), .QN(n10500) );
  NAND2X0 U10486 ( .IN1(n10504), .IN2(n10505), .QN(g27345) );
  OR2X1 U10487 ( .IN1(n10506), .IN2(n6624), .Q(n10505) );
  NAND2X0 U10488 ( .IN1(n10506), .IN2(n10493), .QN(n10504) );
  NAND3X0 U10489 ( .IN1(n9984), .IN2(n9975), .IN3(n10507), .QN(n10493) );
  NAND2X0 U10490 ( .IN1(n10508), .IN2(n10509), .QN(g27344) );
  NAND2X0 U10491 ( .IN1(test_so89), .IN2(n10510), .QN(n10509) );
  NAND2X0 U10492 ( .IN1(n10499), .IN2(n10496), .QN(n10508) );
  NAND2X0 U10493 ( .IN1(n10511), .IN2(n10512), .QN(g27343) );
  OR2X1 U10494 ( .IN1(n10492), .IN2(n6614), .Q(n10512) );
  NAND2X0 U10495 ( .IN1(n10513), .IN2(n10492), .QN(n10511) );
  NAND2X0 U10496 ( .IN1(n10514), .IN2(n10515), .QN(g27342) );
  OR2X1 U10497 ( .IN1(n10516), .IN2(n6914), .Q(n10515) );
  NAND2X0 U10498 ( .IN1(n10516), .IN2(n10517), .QN(n10514) );
  NAND2X0 U10499 ( .IN1(n10518), .IN2(n10519), .QN(g27341) );
  OR2X1 U10500 ( .IN1(n10520), .IN2(n6628), .Q(n10519) );
  NAND2X0 U10501 ( .IN1(n10520), .IN2(n10503), .QN(n10518) );
  NAND2X0 U10502 ( .IN1(n10521), .IN2(n10522), .QN(g27340) );
  OR2X1 U10503 ( .IN1(n10502), .IN2(n6443), .Q(n10522) );
  NAND2X0 U10504 ( .IN1(n10523), .IN2(n10502), .QN(n10521) );
  NAND2X0 U10505 ( .IN1(n10524), .IN2(n10525), .QN(g27339) );
  OR2X1 U10506 ( .IN1(n10526), .IN2(n6630), .Q(n10525) );
  NAND2X0 U10507 ( .IN1(n10526), .IN2(n10527), .QN(n10524) );
  NAND2X0 U10508 ( .IN1(n10528), .IN2(n10529), .QN(g27338) );
  OR2X1 U10509 ( .IN1(n10506), .IN2(n6440), .Q(n10529) );
  NAND2X0 U10510 ( .IN1(n10506), .IN2(n10499), .QN(n10528) );
  AND3X1 U10511 ( .IN1(n10530), .IN2(n10531), .IN3(n10532), .Q(n10499) );
  NAND2X0 U10512 ( .IN1(n10507), .IN2(n9968), .QN(n10531) );
  XOR2X1 U10513 ( .IN1(n9997), .IN2(g3229), .Q(n10507) );
  NAND4X0 U10514 ( .IN1(n9986), .IN2(n7882), .IN3(n9982), .IN4(n9984), .QN(
        n10530) );
  INVX0 U10515 ( .INP(n9968), .ZN(n9984) );
  NAND2X0 U10516 ( .IN1(n10533), .IN2(n10534), .QN(g27337) );
  NAND2X0 U10517 ( .IN1(n10513), .IN2(n10496), .QN(n10534) );
  OR2X1 U10518 ( .IN1(n10496), .IN2(n6615), .Q(n10533) );
  NAND2X0 U10519 ( .IN1(n10535), .IN2(n10536), .QN(g27336) );
  NAND2X0 U10520 ( .IN1(n10537), .IN2(n10492), .QN(n10536) );
  OR2X1 U10521 ( .IN1(n10492), .IN2(n6602), .Q(n10535) );
  AND2X1 U10522 ( .IN1(g22687), .IN2(g2624), .Q(n10492) );
  NAND2X0 U10523 ( .IN1(n10538), .IN2(n10539), .QN(g27335) );
  OR2X1 U10524 ( .IN1(n10540), .IN2(n6915), .Q(n10539) );
  NAND2X0 U10525 ( .IN1(n10540), .IN2(n10517), .QN(n10538) );
  NAND2X0 U10526 ( .IN1(n10541), .IN2(n10542), .QN(g27334) );
  OR2X1 U10527 ( .IN1(n10516), .IN2(n6647), .Q(n10542) );
  NAND2X0 U10528 ( .IN1(n10543), .IN2(n10516), .QN(n10541) );
  NAND2X0 U10529 ( .IN1(n10544), .IN2(n10545), .QN(g27333) );
  NAND2X0 U10530 ( .IN1(n10546), .IN2(n10503), .QN(n10545) );
  NAND2X0 U10531 ( .IN1(n10547), .IN2(n10105), .QN(n10503) );
  NOR2X0 U10532 ( .IN1(n10102), .IN2(n10088), .QN(n10105) );
  NAND2X0 U10533 ( .IN1(test_so67), .IN2(n10548), .QN(n10544) );
  NAND2X0 U10534 ( .IN1(n10549), .IN2(n10550), .QN(g27332) );
  OR2X1 U10535 ( .IN1(n10520), .IN2(n6444), .Q(n10550) );
  NAND2X0 U10536 ( .IN1(n10523), .IN2(n10520), .QN(n10549) );
  NAND2X0 U10537 ( .IN1(n10551), .IN2(n10552), .QN(g27331) );
  OR2X1 U10538 ( .IN1(n10502), .IN2(n6617), .Q(n10552) );
  NAND2X0 U10539 ( .IN1(n10553), .IN2(n10502), .QN(n10551) );
  NAND2X0 U10540 ( .IN1(n10554), .IN2(n10555), .QN(g27330) );
  OR2X1 U10541 ( .IN1(n10556), .IN2(n6917), .Q(n10555) );
  NAND2X0 U10542 ( .IN1(n10556), .IN2(n10557), .QN(n10554) );
  NAND2X0 U10543 ( .IN1(n10558), .IN2(n10559), .QN(g27329) );
  OR2X1 U10544 ( .IN1(n10560), .IN2(n6631), .Q(n10559) );
  NAND2X0 U10545 ( .IN1(n10560), .IN2(n10527), .QN(n10558) );
  NAND2X0 U10546 ( .IN1(n10561), .IN2(n10562), .QN(g27328) );
  NAND2X0 U10547 ( .IN1(test_so46), .IN2(n10563), .QN(n10562) );
  NAND2X0 U10548 ( .IN1(n10564), .IN2(n10526), .QN(n10561) );
  NAND2X0 U10549 ( .IN1(n10565), .IN2(n10566), .QN(g27327) );
  OR2X1 U10550 ( .IN1(n10567), .IN2(n6633), .Q(n10566) );
  NAND2X0 U10551 ( .IN1(n10567), .IN2(n10568), .QN(n10565) );
  NAND2X0 U10552 ( .IN1(n10569), .IN2(n10570), .QN(g27326) );
  OR2X1 U10553 ( .IN1(n10506), .IN2(n6613), .Q(n10570) );
  NAND2X0 U10554 ( .IN1(n10513), .IN2(n10506), .QN(n10569) );
  AND3X1 U10555 ( .IN1(n10571), .IN2(n10000), .IN3(n10572), .Q(n10513) );
  NAND3X0 U10556 ( .IN1(n9985), .IN2(n7882), .IN3(n9986), .QN(n10572) );
  INVX0 U10557 ( .INP(n9997), .ZN(n9986) );
  NAND2X0 U10558 ( .IN1(n10573), .IN2(n10574), .QN(g27325) );
  NAND2X0 U10559 ( .IN1(n10537), .IN2(n10496), .QN(n10574) );
  OR2X1 U10560 ( .IN1(n10496), .IN2(n6603), .Q(n10573) );
  INVX0 U10561 ( .INP(n10510), .ZN(n10496) );
  NAND2X0 U10562 ( .IN1(g7390), .IN2(g22687), .QN(n10510) );
  NAND2X0 U10563 ( .IN1(n10575), .IN2(n10576), .QN(g27324) );
  OR2X1 U10564 ( .IN1(n10577), .IN2(n6916), .Q(n10576) );
  NAND2X0 U10565 ( .IN1(n10577), .IN2(n10517), .QN(n10575) );
  NAND3X0 U10566 ( .IN1(n10578), .IN2(n10579), .IN3(n10580), .QN(n10517) );
  NAND2X0 U10567 ( .IN1(n10581), .IN2(n10582), .QN(g27323) );
  OR2X1 U10568 ( .IN1(n10540), .IN2(n6648), .Q(n10582) );
  NAND2X0 U10569 ( .IN1(n10543), .IN2(n10540), .QN(n10581) );
  NAND2X0 U10570 ( .IN1(n10583), .IN2(n10584), .QN(g27322) );
  OR2X1 U10571 ( .IN1(n10516), .IN2(n6902), .Q(n10584) );
  NAND2X0 U10572 ( .IN1(n10585), .IN2(n10516), .QN(n10583) );
  NAND2X0 U10573 ( .IN1(n10586), .IN2(n10587), .QN(g27321) );
  NAND2X0 U10574 ( .IN1(n10546), .IN2(n10523), .QN(n10587) );
  AND3X1 U10575 ( .IN1(n10588), .IN2(n10589), .IN3(n10590), .Q(n10523) );
  NAND2X0 U10576 ( .IN1(n10547), .IN2(n10102), .QN(n10589) );
  XOR2X1 U10577 ( .IN1(n10068), .IN2(g3229), .Q(n10547) );
  NAND4X0 U10578 ( .IN1(n10094), .IN2(n7882), .IN3(n10081), .IN4(n10090), .QN(
        n10588) );
  INVX0 U10579 ( .INP(n10072), .ZN(n10094) );
  OR2X1 U10580 ( .IN1(n10546), .IN2(n6442), .Q(n10586) );
  NAND2X0 U10581 ( .IN1(n10591), .IN2(n10592), .QN(g27320) );
  OR2X1 U10582 ( .IN1(n10520), .IN2(n6618), .Q(n10592) );
  NAND2X0 U10583 ( .IN1(n10553), .IN2(n10520), .QN(n10591) );
  NAND2X0 U10584 ( .IN1(n10593), .IN2(n10594), .QN(g27319) );
  NAND2X0 U10585 ( .IN1(n10595), .IN2(n10502), .QN(n10594) );
  OR2X1 U10586 ( .IN1(n10502), .IN2(n6605), .Q(n10593) );
  AND2X1 U10587 ( .IN1(g22651), .IN2(g1930), .Q(n10502) );
  NAND2X0 U10588 ( .IN1(n10596), .IN2(n10597), .QN(g27318) );
  NAND2X0 U10589 ( .IN1(n10598), .IN2(n10557), .QN(n10597) );
  NAND2X0 U10590 ( .IN1(test_so58), .IN2(n10599), .QN(n10596) );
  NAND2X0 U10591 ( .IN1(n10600), .IN2(n10601), .QN(g27317) );
  OR2X1 U10592 ( .IN1(n10556), .IN2(n6650), .Q(n10601) );
  NAND2X0 U10593 ( .IN1(n10602), .IN2(n10556), .QN(n10600) );
  NAND2X0 U10594 ( .IN1(n10603), .IN2(n10604), .QN(g27316) );
  OR2X1 U10595 ( .IN1(n10605), .IN2(n6629), .Q(n10604) );
  NAND2X0 U10596 ( .IN1(n10605), .IN2(n10527), .QN(n10603) );
  NAND2X0 U10597 ( .IN1(n10606), .IN2(n10205), .QN(n10527) );
  NOR2X0 U10598 ( .IN1(n10202), .IN2(n10188), .QN(n10205) );
  NAND2X0 U10599 ( .IN1(n10607), .IN2(n10608), .QN(g27315) );
  OR2X1 U10600 ( .IN1(n10560), .IN2(n6446), .Q(n10608) );
  NAND2X0 U10601 ( .IN1(n10564), .IN2(n10560), .QN(n10607) );
  NAND2X0 U10602 ( .IN1(n10609), .IN2(n10610), .QN(g27314) );
  NAND2X0 U10603 ( .IN1(n10611), .IN2(n10526), .QN(n10610) );
  OR2X1 U10604 ( .IN1(n10526), .IN2(n6620), .Q(n10609) );
  NAND2X0 U10605 ( .IN1(n10612), .IN2(n10613), .QN(g27313) );
  OR2X1 U10606 ( .IN1(n10614), .IN2(n6919), .Q(n10613) );
  NAND2X0 U10607 ( .IN1(n10614), .IN2(n10615), .QN(n10612) );
  NAND2X0 U10608 ( .IN1(n10616), .IN2(n10617), .QN(g27312) );
  NAND2X0 U10609 ( .IN1(n10618), .IN2(n10568), .QN(n10617) );
  OR2X1 U10610 ( .IN1(n10618), .IN2(n6634), .Q(n10616) );
  NAND2X0 U10611 ( .IN1(n10619), .IN2(n10620), .QN(g27311) );
  OR2X1 U10612 ( .IN1(n10567), .IN2(n6448), .Q(n10620) );
  NAND2X0 U10613 ( .IN1(n10621), .IN2(n10567), .QN(n10619) );
  NAND2X0 U10614 ( .IN1(n10622), .IN2(n10623), .QN(g27310) );
  OR2X1 U10615 ( .IN1(n10506), .IN2(n6601), .Q(n10623) );
  NAND2X0 U10616 ( .IN1(n10537), .IN2(n10506), .QN(n10622) );
  AND2X1 U10617 ( .IN1(g7302), .IN2(g22687), .Q(n10506) );
  AND4X1 U10618 ( .IN1(n10571), .IN2(n10532), .IN3(n10624), .IN4(n10625), .Q(
        n10537) );
  NAND2X0 U10619 ( .IN1(g3229), .IN2(n10010), .QN(n10625) );
  NAND2X0 U10620 ( .IN1(n10626), .IN2(n7882), .QN(n10624) );
  NAND2X0 U10621 ( .IN1(n10627), .IN2(n10000), .QN(n10626) );
  NAND2X0 U10622 ( .IN1(n9975), .IN2(n9968), .QN(n10000) );
  INVX0 U10623 ( .INP(n9985), .ZN(n9975) );
  OR3X1 U10624 ( .IN1(n9968), .IN2(n7882), .IN3(n10627), .Q(n10532) );
  NAND2X0 U10625 ( .IN1(n9982), .IN2(n9997), .QN(n10627) );
  INVX0 U10626 ( .INP(n10010), .ZN(n9982) );
  NAND3X0 U10627 ( .IN1(n10628), .IN2(n10629), .IN3(n10630), .QN(n10010) );
  NAND2X0 U10628 ( .IN1(n6626), .IN2(g7390), .QN(n10630) );
  NAND2X0 U10629 ( .IN1(n6625), .IN2(g2624), .QN(n10629) );
  NAND2X0 U10630 ( .IN1(n6624), .IN2(n9246), .QN(n10628) );
  NAND3X0 U10631 ( .IN1(n10631), .IN2(n10632), .IN3(n10633), .QN(n9968) );
  NAND2X0 U10632 ( .IN1(n6615), .IN2(g7390), .QN(n10633) );
  NAND2X0 U10633 ( .IN1(n6614), .IN2(g2624), .QN(n10632) );
  NAND2X0 U10634 ( .IN1(n6613), .IN2(n9246), .QN(n10631) );
  NAND3X0 U10635 ( .IN1(n9985), .IN2(n9997), .IN3(g3229), .QN(n10571) );
  NAND3X0 U10636 ( .IN1(n10634), .IN2(n10635), .IN3(n10636), .QN(n9997) );
  NAND2X0 U10637 ( .IN1(n6603), .IN2(g7390), .QN(n10636) );
  NAND2X0 U10638 ( .IN1(n6602), .IN2(g2624), .QN(n10635) );
  NAND2X0 U10639 ( .IN1(n6601), .IN2(n9246), .QN(n10634) );
  NAND3X0 U10640 ( .IN1(n10637), .IN2(n10638), .IN3(n10639), .QN(n9985) );
  OR2X1 U10641 ( .IN1(n4370), .IN2(test_so89), .Q(n10639) );
  NAND2X0 U10642 ( .IN1(n6441), .IN2(g2624), .QN(n10638) );
  NAND2X0 U10643 ( .IN1(n6440), .IN2(n9246), .QN(n10637) );
  NAND2X0 U10644 ( .IN1(n10640), .IN2(n10641), .QN(g27309) );
  OR2X1 U10645 ( .IN1(n10577), .IN2(n6646), .Q(n10641) );
  NAND2X0 U10646 ( .IN1(n10577), .IN2(n10543), .QN(n10640) );
  AND3X1 U10647 ( .IN1(n10642), .IN2(n10643), .IN3(n10644), .Q(n10543) );
  NAND2X0 U10648 ( .IN1(n10578), .IN2(n10645), .QN(n10643) );
  XOR2X1 U10649 ( .IN1(n10646), .IN2(g3229), .Q(n10578) );
  OR4X1 U10650 ( .IN1(n10646), .IN2(g3229), .IN3(n10647), .IN4(n10645), .Q(
        n10642) );
  NAND2X0 U10651 ( .IN1(n10648), .IN2(n10649), .QN(g27308) );
  OR2X1 U10652 ( .IN1(n10540), .IN2(n6903), .Q(n10649) );
  NAND2X0 U10653 ( .IN1(n10585), .IN2(n10540), .QN(n10648) );
  NAND2X0 U10654 ( .IN1(n10650), .IN2(n10651), .QN(g27307) );
  NAND2X0 U10655 ( .IN1(n10652), .IN2(n10516), .QN(n10651) );
  OR2X1 U10656 ( .IN1(n10516), .IN2(n6925), .Q(n10650) );
  AND2X1 U10657 ( .IN1(n10653), .IN2(n8841), .Q(n10516) );
  NAND2X0 U10658 ( .IN1(n10654), .IN2(n10655), .QN(g27306) );
  NAND2X0 U10659 ( .IN1(n10553), .IN2(n10546), .QN(n10655) );
  AND3X1 U10660 ( .IN1(n10656), .IN2(n10657), .IN3(n10658), .Q(n10553) );
  NAND3X0 U10661 ( .IN1(n10088), .IN2(n7882), .IN3(n10081), .QN(n10658) );
  OR2X1 U10662 ( .IN1(n10546), .IN2(n6616), .Q(n10654) );
  NAND2X0 U10663 ( .IN1(n10659), .IN2(n10660), .QN(g27305) );
  NAND2X0 U10664 ( .IN1(n10595), .IN2(n10520), .QN(n10660) );
  OR2X1 U10665 ( .IN1(n10520), .IN2(n6606), .Q(n10659) );
  AND2X1 U10666 ( .IN1(g22651), .IN2(g7194), .Q(n10520) );
  NAND2X0 U10667 ( .IN1(n10661), .IN2(n10662), .QN(g27304) );
  OR2X1 U10668 ( .IN1(n10663), .IN2(n6918), .Q(n10662) );
  NAND2X0 U10669 ( .IN1(n10663), .IN2(n10557), .QN(n10661) );
  NAND3X0 U10670 ( .IN1(n10664), .IN2(n10665), .IN3(n10666), .QN(n10557) );
  NAND2X0 U10671 ( .IN1(n10667), .IN2(n10668), .QN(g27303) );
  NAND2X0 U10672 ( .IN1(n10602), .IN2(n10598), .QN(n10668) );
  OR2X1 U10673 ( .IN1(n10598), .IN2(n6651), .Q(n10667) );
  NAND2X0 U10674 ( .IN1(n10669), .IN2(n10670), .QN(g27302) );
  OR2X1 U10675 ( .IN1(n10556), .IN2(n6905), .Q(n10670) );
  NAND2X0 U10676 ( .IN1(n10671), .IN2(n10556), .QN(n10669) );
  NAND2X0 U10677 ( .IN1(n10672), .IN2(n10673), .QN(g27301) );
  OR2X1 U10678 ( .IN1(n10605), .IN2(n6445), .Q(n10673) );
  NAND2X0 U10679 ( .IN1(n10605), .IN2(n10564), .QN(n10672) );
  AND3X1 U10680 ( .IN1(n10674), .IN2(n10675), .IN3(n10676), .Q(n10564) );
  NAND2X0 U10681 ( .IN1(n10606), .IN2(n10202), .QN(n10675) );
  XOR2X1 U10682 ( .IN1(n10168), .IN2(g3229), .Q(n10606) );
  NAND4X0 U10683 ( .IN1(n10194), .IN2(n7882), .IN3(n10181), .IN4(n10190), .QN(
        n10674) );
  INVX0 U10684 ( .INP(n10172), .ZN(n10194) );
  NAND2X0 U10685 ( .IN1(n10677), .IN2(n10678), .QN(g27300) );
  OR2X1 U10686 ( .IN1(n10560), .IN2(n6621), .Q(n10678) );
  NAND2X0 U10687 ( .IN1(n10611), .IN2(n10560), .QN(n10677) );
  NAND2X0 U10688 ( .IN1(n10679), .IN2(n10680), .QN(g27299) );
  NAND2X0 U10689 ( .IN1(n10681), .IN2(n10526), .QN(n10680) );
  OR2X1 U10690 ( .IN1(n10526), .IN2(n6608), .Q(n10679) );
  INVX0 U10691 ( .INP(n10563), .ZN(n10526) );
  NAND2X0 U10692 ( .IN1(g1236), .IN2(g22615), .QN(n10563) );
  NAND2X0 U10693 ( .IN1(n10682), .IN2(n10683), .QN(g27298) );
  OR2X1 U10694 ( .IN1(n10684), .IN2(n6920), .Q(n10683) );
  NAND2X0 U10695 ( .IN1(n10684), .IN2(n10615), .QN(n10682) );
  NAND2X0 U10696 ( .IN1(n10685), .IN2(n10686), .QN(g27297) );
  OR2X1 U10697 ( .IN1(n10614), .IN2(n6653), .Q(n10686) );
  NAND2X0 U10698 ( .IN1(n10687), .IN2(n10614), .QN(n10685) );
  NAND2X0 U10699 ( .IN1(n10688), .IN2(n10689), .QN(g27296) );
  OR2X1 U10700 ( .IN1(n10690), .IN2(n6632), .Q(n10689) );
  NAND2X0 U10701 ( .IN1(n10690), .IN2(n10568), .QN(n10688) );
  NAND2X0 U10702 ( .IN1(n10691), .IN2(n10300), .QN(n10568) );
  NOR2X0 U10703 ( .IN1(n10297), .IN2(n10283), .QN(n10300) );
  NAND2X0 U10704 ( .IN1(n10692), .IN2(n10693), .QN(g27295) );
  NAND2X0 U10705 ( .IN1(n10621), .IN2(n10618), .QN(n10693) );
  OR2X1 U10706 ( .IN1(n10618), .IN2(n6449), .Q(n10692) );
  NAND2X0 U10707 ( .IN1(n10694), .IN2(n10695), .QN(g27294) );
  OR2X1 U10708 ( .IN1(n10567), .IN2(n6623), .Q(n10695) );
  NAND2X0 U10709 ( .IN1(n10696), .IN2(n10567), .QN(n10694) );
  NAND2X0 U10710 ( .IN1(n10697), .IN2(n10698), .QN(g27293) );
  OR2X1 U10711 ( .IN1(n10699), .IN2(n6922), .Q(n10698) );
  NAND2X0 U10712 ( .IN1(n10699), .IN2(n10700), .QN(n10697) );
  NAND2X0 U10713 ( .IN1(n10701), .IN2(n10702), .QN(g27292) );
  OR2X1 U10714 ( .IN1(n10577), .IN2(n6904), .Q(n10702) );
  NAND2X0 U10715 ( .IN1(n10585), .IN2(n10577), .QN(n10701) );
  AND3X1 U10716 ( .IN1(n10703), .IN2(n10704), .IN3(n10705), .Q(n10585) );
  NAND3X0 U10717 ( .IN1(n10706), .IN2(n7882), .IN3(n10707), .QN(n10703) );
  NAND2X0 U10718 ( .IN1(n10708), .IN2(n10709), .QN(g27291) );
  NAND2X0 U10719 ( .IN1(n10652), .IN2(n10540), .QN(n10709) );
  OR2X1 U10720 ( .IN1(n10540), .IN2(n6926), .Q(n10708) );
  AND2X1 U10721 ( .IN1(n10653), .IN2(g7264), .Q(n10540) );
  NAND2X0 U10722 ( .IN1(n10710), .IN2(n10711), .QN(g27290) );
  NAND2X0 U10723 ( .IN1(n10595), .IN2(n10546), .QN(n10711) );
  AND4X1 U10724 ( .IN1(n10656), .IN2(n10590), .IN3(n10712), .IN4(n10713), .Q(
        n10595) );
  NAND2X0 U10725 ( .IN1(g3229), .IN2(n10072), .QN(n10713) );
  NAND2X0 U10726 ( .IN1(n10714), .IN2(n7882), .QN(n10712) );
  OR2X1 U10727 ( .IN1(n10715), .IN2(n10096), .Q(n10714) );
  INVX0 U10728 ( .INP(n10657), .ZN(n10096) );
  NAND2X0 U10729 ( .IN1(n10092), .IN2(n10102), .QN(n10657) );
  INVX0 U10730 ( .INP(n10088), .ZN(n10092) );
  NAND3X0 U10731 ( .IN1(n10090), .IN2(g3229), .IN3(n10715), .QN(n10590) );
  NOR2X0 U10732 ( .IN1(n10072), .IN2(n10081), .QN(n10715) );
  INVX0 U10733 ( .INP(n10068), .ZN(n10081) );
  NAND3X0 U10734 ( .IN1(n10716), .IN2(n10717), .IN3(n10718), .QN(n10072) );
  NAND2X0 U10735 ( .IN1(n6627), .IN2(g1930), .QN(n10718) );
  OR2X1 U10736 ( .IN1(n4296), .IN2(test_so67), .Q(n10717) );
  NAND2X0 U10737 ( .IN1(n6628), .IN2(g7194), .QN(n10716) );
  INVX0 U10738 ( .INP(n10102), .ZN(n10090) );
  NAND3X0 U10739 ( .IN1(n10719), .IN2(n10720), .IN3(n10721), .QN(n10102) );
  NAND2X0 U10740 ( .IN1(n6617), .IN2(g1930), .QN(n10721) );
  NAND2X0 U10741 ( .IN1(n6616), .IN2(n9268), .QN(n10720) );
  NAND2X0 U10742 ( .IN1(n6618), .IN2(g7194), .QN(n10719) );
  NAND3X0 U10743 ( .IN1(n10088), .IN2(n10068), .IN3(g3229), .QN(n10656) );
  NAND3X0 U10744 ( .IN1(n10722), .IN2(n10723), .IN3(n10724), .QN(n10068) );
  NAND2X0 U10745 ( .IN1(n6605), .IN2(g1930), .QN(n10724) );
  NAND2X0 U10746 ( .IN1(n6604), .IN2(n9268), .QN(n10723) );
  NAND2X0 U10747 ( .IN1(n6606), .IN2(g7194), .QN(n10722) );
  NAND3X0 U10748 ( .IN1(n10725), .IN2(n10726), .IN3(n10727), .QN(n10088) );
  NAND2X0 U10749 ( .IN1(n6443), .IN2(g1930), .QN(n10727) );
  NAND2X0 U10750 ( .IN1(n6442), .IN2(n9268), .QN(n10726) );
  NAND2X0 U10751 ( .IN1(n6444), .IN2(g7194), .QN(n10725) );
  OR2X1 U10752 ( .IN1(n10546), .IN2(n6604), .Q(n10710) );
  INVX0 U10753 ( .INP(n10548), .ZN(n10546) );
  NAND2X0 U10754 ( .IN1(g7052), .IN2(g22651), .QN(n10548) );
  NAND2X0 U10755 ( .IN1(n10728), .IN2(n10729), .QN(g27289) );
  OR2X1 U10756 ( .IN1(n10663), .IN2(n6649), .Q(n10729) );
  NAND2X0 U10757 ( .IN1(n10663), .IN2(n10602), .QN(n10728) );
  AND3X1 U10758 ( .IN1(n10730), .IN2(n10731), .IN3(n10732), .Q(n10602) );
  NAND2X0 U10759 ( .IN1(n10664), .IN2(n10733), .QN(n10731) );
  XOR2X1 U10760 ( .IN1(n10734), .IN2(g3229), .Q(n10664) );
  OR4X1 U10761 ( .IN1(n10734), .IN2(g3229), .IN3(n10735), .IN4(n10733), .Q(
        n10730) );
  NAND2X0 U10762 ( .IN1(n10736), .IN2(n10737), .QN(g27288) );
  NAND2X0 U10763 ( .IN1(n10671), .IN2(n10598), .QN(n10737) );
  OR2X1 U10764 ( .IN1(n10598), .IN2(n6906), .Q(n10736) );
  NAND2X0 U10765 ( .IN1(n10738), .IN2(n10739), .QN(g27287) );
  NAND2X0 U10766 ( .IN1(n10740), .IN2(n10556), .QN(n10739) );
  OR2X1 U10767 ( .IN1(n10556), .IN2(n6928), .Q(n10738) );
  AND2X1 U10768 ( .IN1(n10741), .IN2(n8453), .Q(n10556) );
  NAND2X0 U10769 ( .IN1(n10742), .IN2(n10743), .QN(g27286) );
  OR2X1 U10770 ( .IN1(n10605), .IN2(n6619), .Q(n10743) );
  NAND2X0 U10771 ( .IN1(n10611), .IN2(n10605), .QN(n10742) );
  AND3X1 U10772 ( .IN1(n10744), .IN2(n10745), .IN3(n10746), .Q(n10611) );
  NAND3X0 U10773 ( .IN1(n10188), .IN2(n7882), .IN3(n10181), .QN(n10746) );
  NAND2X0 U10774 ( .IN1(n10747), .IN2(n10748), .QN(g27285) );
  NAND2X0 U10775 ( .IN1(n10681), .IN2(n10560), .QN(n10748) );
  OR2X1 U10776 ( .IN1(n10560), .IN2(n6609), .Q(n10747) );
  AND2X1 U10777 ( .IN1(g22615), .IN2(g6944), .Q(n10560) );
  NAND2X0 U10778 ( .IN1(n10749), .IN2(n10750), .QN(g27284) );
  NAND2X0 U10779 ( .IN1(n10751), .IN2(n10615), .QN(n10750) );
  NAND3X0 U10780 ( .IN1(n10752), .IN2(n10753), .IN3(n10754), .QN(n10615) );
  OR2X1 U10781 ( .IN1(n10751), .IN2(n6921), .Q(n10749) );
  NAND2X0 U10782 ( .IN1(n10755), .IN2(n10756), .QN(g27283) );
  OR2X1 U10783 ( .IN1(n10684), .IN2(n6652), .Q(n10756) );
  NAND2X0 U10784 ( .IN1(n10687), .IN2(n10684), .QN(n10755) );
  NAND2X0 U10785 ( .IN1(n10757), .IN2(n10758), .QN(g27282) );
  OR2X1 U10786 ( .IN1(n10614), .IN2(n6908), .Q(n10758) );
  NAND2X0 U10787 ( .IN1(n10759), .IN2(n10614), .QN(n10757) );
  NAND2X0 U10788 ( .IN1(n10760), .IN2(n10761), .QN(g27281) );
  OR2X1 U10789 ( .IN1(n10690), .IN2(n6447), .Q(n10761) );
  NAND2X0 U10790 ( .IN1(n10690), .IN2(n10621), .QN(n10760) );
  AND3X1 U10791 ( .IN1(n10762), .IN2(n10763), .IN3(n10764), .Q(n10621) );
  NAND2X0 U10792 ( .IN1(n10691), .IN2(n10297), .QN(n10763) );
  XOR2X1 U10793 ( .IN1(n10263), .IN2(g3229), .Q(n10691) );
  NAND4X0 U10794 ( .IN1(n10289), .IN2(n7882), .IN3(n10276), .IN4(n10285), .QN(
        n10762) );
  INVX0 U10795 ( .INP(n10267), .ZN(n10289) );
  NAND2X0 U10796 ( .IN1(n10765), .IN2(n10766), .QN(g27280) );
  NAND2X0 U10797 ( .IN1(test_so25), .IN2(n10767), .QN(n10766) );
  NAND2X0 U10798 ( .IN1(n10696), .IN2(n10618), .QN(n10765) );
  NAND2X0 U10799 ( .IN1(n10768), .IN2(n10769), .QN(g27279) );
  NAND2X0 U10800 ( .IN1(n10770), .IN2(n10567), .QN(n10769) );
  OR2X1 U10801 ( .IN1(n10567), .IN2(n6611), .Q(n10768) );
  AND2X1 U10802 ( .IN1(g22578), .IN2(g550), .Q(n10567) );
  NAND2X0 U10803 ( .IN1(n10771), .IN2(n10772), .QN(g27278) );
  OR2X1 U10804 ( .IN1(n10773), .IN2(n6923), .Q(n10772) );
  NAND2X0 U10805 ( .IN1(n10773), .IN2(n10700), .QN(n10771) );
  NAND2X0 U10806 ( .IN1(n10774), .IN2(n10775), .QN(g27277) );
  NAND2X0 U10807 ( .IN1(n10776), .IN2(n10699), .QN(n10775) );
  OR2X1 U10808 ( .IN1(n10699), .IN2(n6655), .Q(n10774) );
  NAND2X0 U10809 ( .IN1(n10777), .IN2(n10778), .QN(g27276) );
  OR2X1 U10810 ( .IN1(n10577), .IN2(n6927), .Q(n10778) );
  NAND2X0 U10811 ( .IN1(n10652), .IN2(n10577), .QN(n10777) );
  AND2X1 U10812 ( .IN1(n10653), .IN2(g5555), .Q(n10577) );
  AND2X1 U10813 ( .IN1(n10779), .IN2(n7772), .Q(n10653) );
  NAND2X0 U10814 ( .IN1(n10780), .IN2(n7749), .QN(n10779) );
  INVX0 U10815 ( .INP(n10781), .ZN(n7749) );
  AND4X1 U10816 ( .IN1(n10704), .IN2(n10644), .IN3(n10782), .IN4(n10783), .Q(
        n10652) );
  NAND2X0 U10817 ( .IN1(g3229), .IN2(n10647), .QN(n10783) );
  NAND2X0 U10818 ( .IN1(n10784), .IN2(n7882), .QN(n10782) );
  NAND2X0 U10819 ( .IN1(n10705), .IN2(n10785), .QN(n10784) );
  INVX0 U10820 ( .INP(n10786), .ZN(n10785) );
  NAND2X0 U10821 ( .IN1(n10580), .IN2(n10645), .QN(n10705) );
  INVX0 U10822 ( .INP(n10706), .ZN(n10580) );
  NAND3X0 U10823 ( .IN1(n10579), .IN2(g3229), .IN3(n10786), .QN(n10644) );
  NOR2X0 U10824 ( .IN1(n10647), .IN2(n10707), .QN(n10786) );
  INVX0 U10825 ( .INP(n10646), .ZN(n10707) );
  NAND3X0 U10826 ( .IN1(n10787), .IN2(n10788), .IN3(n10789), .QN(n10647) );
  NAND2X0 U10827 ( .IN1(n6915), .IN2(n8449), .QN(n10789) );
  NAND2X0 U10828 ( .IN1(n6914), .IN2(n8841), .QN(n10788) );
  NAND2X0 U10829 ( .IN1(n6916), .IN2(n8456), .QN(n10787) );
  INVX0 U10830 ( .INP(n10645), .ZN(n10579) );
  NAND3X0 U10831 ( .IN1(n10790), .IN2(n10791), .IN3(n10792), .QN(n10645) );
  NAND2X0 U10832 ( .IN1(n6903), .IN2(n8449), .QN(n10792) );
  NAND2X0 U10833 ( .IN1(n6902), .IN2(n8841), .QN(n10791) );
  NAND2X0 U10834 ( .IN1(n6904), .IN2(n8456), .QN(n10790) );
  NAND3X0 U10835 ( .IN1(n10646), .IN2(n10706), .IN3(g3229), .QN(n10704) );
  NAND3X0 U10836 ( .IN1(n10793), .IN2(n10794), .IN3(n10795), .QN(n10706) );
  NAND2X0 U10837 ( .IN1(n6648), .IN2(n8449), .QN(n10795) );
  NAND2X0 U10838 ( .IN1(n6647), .IN2(n8841), .QN(n10794) );
  NAND2X0 U10839 ( .IN1(n6646), .IN2(n8456), .QN(n10793) );
  NAND3X0 U10840 ( .IN1(n10796), .IN2(n10797), .IN3(n10798), .QN(n10646) );
  NAND2X0 U10841 ( .IN1(n6926), .IN2(n8449), .QN(n10798) );
  NAND2X0 U10842 ( .IN1(n6925), .IN2(n8841), .QN(n10797) );
  NAND2X0 U10843 ( .IN1(n6927), .IN2(n8456), .QN(n10796) );
  NAND2X0 U10844 ( .IN1(n10799), .IN2(n10800), .QN(g27275) );
  OR2X1 U10845 ( .IN1(n10663), .IN2(n6907), .Q(n10800) );
  NAND2X0 U10846 ( .IN1(n10671), .IN2(n10663), .QN(n10799) );
  AND3X1 U10847 ( .IN1(n10801), .IN2(n10802), .IN3(n10803), .Q(n10671) );
  NAND3X0 U10848 ( .IN1(n10804), .IN2(n7882), .IN3(n10805), .QN(n10801) );
  NAND2X0 U10849 ( .IN1(n10806), .IN2(n10807), .QN(g27274) );
  NAND2X0 U10850 ( .IN1(n10740), .IN2(n10598), .QN(n10807) );
  OR2X1 U10851 ( .IN1(n10598), .IN2(n6929), .Q(n10806) );
  INVX0 U10852 ( .INP(n10599), .ZN(n10598) );
  NAND2X0 U10853 ( .IN1(n10741), .IN2(g7014), .QN(n10599) );
  NAND2X0 U10854 ( .IN1(n10808), .IN2(n10809), .QN(g27273) );
  OR2X1 U10855 ( .IN1(n10605), .IN2(n6607), .Q(n10809) );
  NAND2X0 U10856 ( .IN1(n10681), .IN2(n10605), .QN(n10808) );
  AND2X1 U10857 ( .IN1(g6750), .IN2(g22615), .Q(n10605) );
  AND4X1 U10858 ( .IN1(n10744), .IN2(n10676), .IN3(n10810), .IN4(n10811), .Q(
        n10681) );
  NAND2X0 U10859 ( .IN1(g3229), .IN2(n10172), .QN(n10811) );
  NAND2X0 U10860 ( .IN1(n10812), .IN2(n7882), .QN(n10810) );
  OR2X1 U10861 ( .IN1(n10813), .IN2(n10196), .Q(n10812) );
  INVX0 U10862 ( .INP(n10745), .ZN(n10196) );
  NAND2X0 U10863 ( .IN1(n10192), .IN2(n10202), .QN(n10745) );
  INVX0 U10864 ( .INP(n10188), .ZN(n10192) );
  NAND3X0 U10865 ( .IN1(n10190), .IN2(g3229), .IN3(n10813), .QN(n10676) );
  NOR2X0 U10866 ( .IN1(n10172), .IN2(n10181), .QN(n10813) );
  INVX0 U10867 ( .INP(n10168), .ZN(n10181) );
  NAND3X0 U10868 ( .IN1(n10814), .IN2(n10815), .IN3(n10816), .QN(n10172) );
  NAND2X0 U10869 ( .IN1(n6629), .IN2(n10142), .QN(n10816) );
  NAND2X0 U10870 ( .IN1(n6630), .IN2(g1236), .QN(n10815) );
  NAND2X0 U10871 ( .IN1(n6631), .IN2(g6944), .QN(n10814) );
  INVX0 U10872 ( .INP(n10202), .ZN(n10190) );
  NAND3X0 U10873 ( .IN1(n10817), .IN2(n10818), .IN3(n10819), .QN(n10202) );
  NAND2X0 U10874 ( .IN1(n6619), .IN2(n10142), .QN(n10819) );
  NAND2X0 U10875 ( .IN1(n6620), .IN2(g1236), .QN(n10818) );
  NAND2X0 U10876 ( .IN1(n6621), .IN2(g6944), .QN(n10817) );
  NAND3X0 U10877 ( .IN1(n10188), .IN2(n10168), .IN3(g3229), .QN(n10744) );
  NAND3X0 U10878 ( .IN1(n10820), .IN2(n10821), .IN3(n10822), .QN(n10168) );
  NAND2X0 U10879 ( .IN1(n6607), .IN2(n10142), .QN(n10822) );
  NAND2X0 U10880 ( .IN1(n6608), .IN2(g1236), .QN(n10821) );
  NAND2X0 U10881 ( .IN1(n6609), .IN2(g6944), .QN(n10820) );
  NAND3X0 U10882 ( .IN1(n10823), .IN2(n10824), .IN3(n10825), .QN(n10188) );
  NAND2X0 U10883 ( .IN1(n6445), .IN2(n10142), .QN(n10825) );
  OR2X1 U10884 ( .IN1(n4300), .IN2(test_so46), .Q(n10824) );
  NAND2X0 U10885 ( .IN1(n6446), .IN2(g6944), .QN(n10823) );
  NAND2X0 U10886 ( .IN1(n10826), .IN2(n10827), .QN(g27272) );
  NAND2X0 U10887 ( .IN1(test_so37), .IN2(n10828), .QN(n10827) );
  NAND2X0 U10888 ( .IN1(n10751), .IN2(n10687), .QN(n10826) );
  AND3X1 U10889 ( .IN1(n10829), .IN2(n10830), .IN3(n10831), .Q(n10687) );
  NAND2X0 U10890 ( .IN1(n10752), .IN2(n10832), .QN(n10830) );
  XOR2X1 U10891 ( .IN1(n10833), .IN2(g3229), .Q(n10752) );
  OR4X1 U10892 ( .IN1(n10833), .IN2(g3229), .IN3(n10834), .IN4(n10832), .Q(
        n10829) );
  NAND2X0 U10893 ( .IN1(n10835), .IN2(n10836), .QN(g27271) );
  OR2X1 U10894 ( .IN1(n10684), .IN2(n6909), .Q(n10836) );
  NAND2X0 U10895 ( .IN1(n10759), .IN2(n10684), .QN(n10835) );
  NAND2X0 U10896 ( .IN1(n10837), .IN2(n10838), .QN(g27270) );
  NAND2X0 U10897 ( .IN1(n10839), .IN2(n10614), .QN(n10838) );
  OR2X1 U10898 ( .IN1(n10614), .IN2(n6931), .Q(n10837) );
  AND2X1 U10899 ( .IN1(n10840), .IN2(g1088), .Q(n10614) );
  NAND2X0 U10900 ( .IN1(n10841), .IN2(n10842), .QN(g27269) );
  OR2X1 U10901 ( .IN1(n10690), .IN2(n6622), .Q(n10842) );
  NAND2X0 U10902 ( .IN1(n10696), .IN2(n10690), .QN(n10841) );
  AND3X1 U10903 ( .IN1(n10843), .IN2(n10844), .IN3(n10845), .Q(n10696) );
  NAND3X0 U10904 ( .IN1(n10283), .IN2(n7882), .IN3(n10276), .QN(n10845) );
  NAND2X0 U10905 ( .IN1(n10846), .IN2(n10847), .QN(g27268) );
  NAND2X0 U10906 ( .IN1(n10770), .IN2(n10618), .QN(n10847) );
  OR2X1 U10907 ( .IN1(n10618), .IN2(n6612), .Q(n10846) );
  INVX0 U10908 ( .INP(n10767), .ZN(n10618) );
  NAND2X0 U10909 ( .IN1(g6642), .IN2(g22578), .QN(n10767) );
  NAND2X0 U10910 ( .IN1(n10848), .IN2(n10849), .QN(g27267) );
  OR2X1 U10911 ( .IN1(n10850), .IN2(n6924), .Q(n10849) );
  NAND2X0 U10912 ( .IN1(n10850), .IN2(n10700), .QN(n10848) );
  NAND3X0 U10913 ( .IN1(n10851), .IN2(n10852), .IN3(n10853), .QN(n10700) );
  NAND2X0 U10914 ( .IN1(n10854), .IN2(n10855), .QN(g27266) );
  OR2X1 U10915 ( .IN1(n10773), .IN2(n6656), .Q(n10855) );
  NAND2X0 U10916 ( .IN1(n10776), .IN2(n10773), .QN(n10854) );
  NAND2X0 U10917 ( .IN1(n10856), .IN2(n10857), .QN(g27265) );
  NAND2X0 U10918 ( .IN1(n10858), .IN2(n10699), .QN(n10857) );
  OR2X1 U10919 ( .IN1(n10699), .IN2(n6911), .Q(n10856) );
  NAND2X0 U10920 ( .IN1(n10859), .IN2(n10860), .QN(g27264) );
  OR2X1 U10921 ( .IN1(n10663), .IN2(n6930), .Q(n10860) );
  NAND2X0 U10922 ( .IN1(n10740), .IN2(n10663), .QN(n10859) );
  AND2X1 U10923 ( .IN1(n10741), .IN2(g5511), .Q(n10663) );
  AND2X1 U10924 ( .IN1(n10861), .IN2(n7736), .Q(n10741) );
  NAND2X0 U10925 ( .IN1(n10780), .IN2(n7720), .QN(n10861) );
  INVX0 U10926 ( .INP(n10862), .ZN(n7720) );
  AND4X1 U10927 ( .IN1(n10802), .IN2(n10732), .IN3(n10863), .IN4(n10864), .Q(
        n10740) );
  NAND2X0 U10928 ( .IN1(g3229), .IN2(n10735), .QN(n10864) );
  NAND2X0 U10929 ( .IN1(n10865), .IN2(n7882), .QN(n10863) );
  NAND2X0 U10930 ( .IN1(n10803), .IN2(n10866), .QN(n10865) );
  INVX0 U10931 ( .INP(n10867), .ZN(n10866) );
  NAND2X0 U10932 ( .IN1(n10666), .IN2(n10733), .QN(n10803) );
  INVX0 U10933 ( .INP(n10804), .ZN(n10666) );
  NAND3X0 U10934 ( .IN1(n10665), .IN2(g3229), .IN3(n10867), .QN(n10732) );
  NOR2X0 U10935 ( .IN1(n10735), .IN2(n10805), .QN(n10867) );
  INVX0 U10936 ( .INP(n10734), .ZN(n10805) );
  NAND3X0 U10937 ( .IN1(n10868), .IN2(n10869), .IN3(n10870), .QN(n10735) );
  OR2X1 U10938 ( .IN1(n4525), .IN2(test_so58), .Q(n10870) );
  NAND2X0 U10939 ( .IN1(n6917), .IN2(n8453), .QN(n10869) );
  NAND2X0 U10940 ( .IN1(n6918), .IN2(n8494), .QN(n10868) );
  INVX0 U10941 ( .INP(n10733), .ZN(n10665) );
  NAND3X0 U10942 ( .IN1(n10871), .IN2(n10872), .IN3(n10873), .QN(n10733) );
  NAND2X0 U10943 ( .IN1(n6906), .IN2(n8459), .QN(n10873) );
  NAND2X0 U10944 ( .IN1(n6905), .IN2(n8453), .QN(n10872) );
  NAND2X0 U10945 ( .IN1(n6907), .IN2(n8494), .QN(n10871) );
  NAND3X0 U10946 ( .IN1(n10734), .IN2(n10804), .IN3(g3229), .QN(n10802) );
  NAND3X0 U10947 ( .IN1(n10874), .IN2(n10875), .IN3(n10876), .QN(n10804) );
  NAND2X0 U10948 ( .IN1(n6651), .IN2(n8459), .QN(n10876) );
  NAND2X0 U10949 ( .IN1(n6650), .IN2(n8453), .QN(n10875) );
  NAND2X0 U10950 ( .IN1(n6649), .IN2(n8494), .QN(n10874) );
  NAND3X0 U10951 ( .IN1(n10877), .IN2(n10878), .IN3(n10879), .QN(n10734) );
  NAND2X0 U10952 ( .IN1(n6929), .IN2(n8459), .QN(n10879) );
  NAND2X0 U10953 ( .IN1(n6928), .IN2(n8453), .QN(n10878) );
  NAND2X0 U10954 ( .IN1(n6930), .IN2(n8494), .QN(n10877) );
  NAND2X0 U10955 ( .IN1(n10880), .IN2(n10881), .QN(g27263) );
  NAND2X0 U10956 ( .IN1(n10759), .IN2(n10751), .QN(n10881) );
  AND3X1 U10957 ( .IN1(n10882), .IN2(n10883), .IN3(n10884), .Q(n10759) );
  NAND3X0 U10958 ( .IN1(n10885), .IN2(n7882), .IN3(n10886), .QN(n10882) );
  OR2X1 U10959 ( .IN1(n10751), .IN2(n6910), .Q(n10880) );
  NAND2X0 U10960 ( .IN1(n10887), .IN2(n10888), .QN(g27262) );
  NAND2X0 U10961 ( .IN1(n10839), .IN2(n10684), .QN(n10888) );
  OR2X1 U10962 ( .IN1(n10684), .IN2(n6932), .Q(n10887) );
  AND2X1 U10963 ( .IN1(n10840), .IN2(g6712), .Q(n10684) );
  NAND2X0 U10964 ( .IN1(n10889), .IN2(n10890), .QN(g27261) );
  OR2X1 U10965 ( .IN1(n10690), .IN2(n6610), .Q(n10890) );
  NAND2X0 U10966 ( .IN1(n10770), .IN2(n10690), .QN(n10889) );
  AND2X1 U10967 ( .IN1(g6485), .IN2(g22578), .Q(n10690) );
  AND4X1 U10968 ( .IN1(n10843), .IN2(n10764), .IN3(n10891), .IN4(n10892), .Q(
        n10770) );
  NAND2X0 U10969 ( .IN1(g3229), .IN2(n10267), .QN(n10892) );
  NAND2X0 U10970 ( .IN1(n10893), .IN2(n7882), .QN(n10891) );
  OR2X1 U10971 ( .IN1(n10894), .IN2(n10291), .Q(n10893) );
  INVX0 U10972 ( .INP(n10844), .ZN(n10291) );
  NAND2X0 U10973 ( .IN1(n10287), .IN2(n10297), .QN(n10844) );
  INVX0 U10974 ( .INP(n10283), .ZN(n10287) );
  NAND3X0 U10975 ( .IN1(n10285), .IN2(g3229), .IN3(n10894), .QN(n10764) );
  NOR2X0 U10976 ( .IN1(n10267), .IN2(n10276), .QN(n10894) );
  INVX0 U10977 ( .INP(n10263), .ZN(n10276) );
  NAND3X0 U10978 ( .IN1(n10895), .IN2(n10896), .IN3(n10897), .QN(n10267) );
  NAND2X0 U10979 ( .IN1(n6634), .IN2(g6642), .QN(n10897) );
  NAND2X0 U10980 ( .IN1(n6632), .IN2(n10242), .QN(n10896) );
  NAND2X0 U10981 ( .IN1(n6633), .IN2(g550), .QN(n10895) );
  INVX0 U10982 ( .INP(n10297), .ZN(n10285) );
  NAND3X0 U10983 ( .IN1(n10898), .IN2(n10899), .IN3(n10900), .QN(n10297) );
  OR2X1 U10984 ( .IN1(n4372), .IN2(test_so25), .Q(n10900) );
  NAND2X0 U10985 ( .IN1(n6622), .IN2(n10242), .QN(n10899) );
  NAND2X0 U10986 ( .IN1(n6623), .IN2(g550), .QN(n10898) );
  NAND3X0 U10987 ( .IN1(n10283), .IN2(n10263), .IN3(g3229), .QN(n10843) );
  NAND3X0 U10988 ( .IN1(n10901), .IN2(n10902), .IN3(n10903), .QN(n10263) );
  NAND2X0 U10989 ( .IN1(n6612), .IN2(g6642), .QN(n10903) );
  NAND2X0 U10990 ( .IN1(n6610), .IN2(n10242), .QN(n10902) );
  NAND2X0 U10991 ( .IN1(n6611), .IN2(g550), .QN(n10901) );
  NAND3X0 U10992 ( .IN1(n10904), .IN2(n10905), .IN3(n10906), .QN(n10283) );
  NAND2X0 U10993 ( .IN1(n6449), .IN2(g6642), .QN(n10906) );
  NAND2X0 U10994 ( .IN1(n6447), .IN2(n10242), .QN(n10905) );
  NAND2X0 U10995 ( .IN1(n6448), .IN2(g550), .QN(n10904) );
  NAND2X0 U10996 ( .IN1(n10907), .IN2(n10908), .QN(g27260) );
  OR2X1 U10997 ( .IN1(n10850), .IN2(n6654), .Q(n10908) );
  NAND2X0 U10998 ( .IN1(n10850), .IN2(n10776), .QN(n10907) );
  AND3X1 U10999 ( .IN1(n10909), .IN2(n10910), .IN3(n10911), .Q(n10776) );
  NAND2X0 U11000 ( .IN1(n10851), .IN2(n10912), .QN(n10910) );
  XOR2X1 U11001 ( .IN1(n10913), .IN2(g3229), .Q(n10851) );
  OR4X1 U11002 ( .IN1(n10913), .IN2(g3229), .IN3(n10914), .IN4(n10912), .Q(
        n10909) );
  NAND2X0 U11003 ( .IN1(n10915), .IN2(n10916), .QN(g27259) );
  OR2X1 U11004 ( .IN1(n10773), .IN2(n6912), .Q(n10916) );
  NAND2X0 U11005 ( .IN1(n10858), .IN2(n10773), .QN(n10915) );
  NAND2X0 U11006 ( .IN1(n10917), .IN2(n10918), .QN(g27258) );
  NAND2X0 U11007 ( .IN1(test_so16), .IN2(n10919), .QN(n10918) );
  NAND2X0 U11008 ( .IN1(n10920), .IN2(n10699), .QN(n10917) );
  INVX0 U11009 ( .INP(n10919), .ZN(n10699) );
  NAND2X0 U11010 ( .IN1(n10921), .IN2(n8500), .QN(n10919) );
  NAND2X0 U11011 ( .IN1(n10922), .IN2(n10923), .QN(g27257) );
  NAND2X0 U11012 ( .IN1(n10839), .IN2(n10751), .QN(n10923) );
  AND4X1 U11013 ( .IN1(n10883), .IN2(n10831), .IN3(n10924), .IN4(n10925), .Q(
        n10839) );
  NAND2X0 U11014 ( .IN1(g3229), .IN2(n10834), .QN(n10925) );
  NAND2X0 U11015 ( .IN1(n10926), .IN2(n7882), .QN(n10924) );
  NAND2X0 U11016 ( .IN1(n10884), .IN2(n10927), .QN(n10926) );
  INVX0 U11017 ( .INP(n10928), .ZN(n10927) );
  NAND2X0 U11018 ( .IN1(n10754), .IN2(n10832), .QN(n10884) );
  INVX0 U11019 ( .INP(n10885), .ZN(n10754) );
  NAND3X0 U11020 ( .IN1(n10753), .IN2(g3229), .IN3(n10928), .QN(n10831) );
  NOR2X0 U11021 ( .IN1(n10834), .IN2(n10886), .QN(n10928) );
  INVX0 U11022 ( .INP(n10833), .ZN(n10886) );
  NAND3X0 U11023 ( .IN1(n10929), .IN2(n10930), .IN3(n10931), .QN(n10834) );
  NAND2X0 U11024 ( .IN1(n6919), .IN2(g1088), .QN(n10931) );
  NAND2X0 U11025 ( .IN1(n6921), .IN2(g5472), .QN(n10930) );
  NAND2X0 U11026 ( .IN1(n6920), .IN2(g6712), .QN(n10929) );
  INVX0 U11027 ( .INP(n10832), .ZN(n10753) );
  NAND3X0 U11028 ( .IN1(n10932), .IN2(n10933), .IN3(n10934), .QN(n10832) );
  NAND2X0 U11029 ( .IN1(n6908), .IN2(g1088), .QN(n10934) );
  NAND2X0 U11030 ( .IN1(n6910), .IN2(g5472), .QN(n10933) );
  NAND2X0 U11031 ( .IN1(n6909), .IN2(g6712), .QN(n10932) );
  NAND3X0 U11032 ( .IN1(n10833), .IN2(n10885), .IN3(g3229), .QN(n10883) );
  NAND3X0 U11033 ( .IN1(n10935), .IN2(n10936), .IN3(n10937), .QN(n10885) );
  NAND2X0 U11034 ( .IN1(n6653), .IN2(g1088), .QN(n10937) );
  OR2X1 U11035 ( .IN1(n4363), .IN2(test_so37), .Q(n10936) );
  NAND2X0 U11036 ( .IN1(n6652), .IN2(g6712), .QN(n10935) );
  NAND3X0 U11037 ( .IN1(n10938), .IN2(n10939), .IN3(n10940), .QN(n10833) );
  NAND2X0 U11038 ( .IN1(n6931), .IN2(g1088), .QN(n10940) );
  NAND2X0 U11039 ( .IN1(n6933), .IN2(g5472), .QN(n10939) );
  NAND2X0 U11040 ( .IN1(n6932), .IN2(g6712), .QN(n10938) );
  OR2X1 U11041 ( .IN1(n10751), .IN2(n6933), .Q(n10922) );
  INVX0 U11042 ( .INP(n10828), .ZN(n10751) );
  NAND2X0 U11043 ( .IN1(n10840), .IN2(g5472), .QN(n10828) );
  AND2X1 U11044 ( .IN1(n10941), .IN2(n7714), .Q(n10840) );
  NAND2X0 U11045 ( .IN1(n10780), .IN2(n7691), .QN(n10941) );
  INVX0 U11046 ( .INP(n10942), .ZN(n7691) );
  NAND2X0 U11047 ( .IN1(n10943), .IN2(n10944), .QN(g27256) );
  OR2X1 U11048 ( .IN1(n10850), .IN2(n6913), .Q(n10944) );
  NAND2X0 U11049 ( .IN1(n10858), .IN2(n10850), .QN(n10943) );
  AND3X1 U11050 ( .IN1(n10945), .IN2(n10946), .IN3(n10947), .Q(n10858) );
  NAND3X0 U11051 ( .IN1(n10948), .IN2(n7882), .IN3(n10949), .QN(n10945) );
  NAND2X0 U11052 ( .IN1(n10950), .IN2(n10951), .QN(g27255) );
  NAND2X0 U11053 ( .IN1(n10920), .IN2(n10773), .QN(n10951) );
  OR2X1 U11054 ( .IN1(n10773), .IN2(n6934), .Q(n10950) );
  AND2X1 U11055 ( .IN1(n10921), .IN2(g6447), .Q(n10773) );
  NAND2X0 U11056 ( .IN1(n10952), .IN2(n10953), .QN(g27253) );
  OR2X1 U11057 ( .IN1(n10850), .IN2(n6935), .Q(n10953) );
  NAND2X0 U11058 ( .IN1(n10920), .IN2(n10850), .QN(n10952) );
  AND2X1 U11059 ( .IN1(n10921), .IN2(g5437), .Q(n10850) );
  AND2X1 U11060 ( .IN1(n10954), .IN2(n7677), .Q(n10921) );
  NAND2X0 U11061 ( .IN1(n10780), .IN2(n7662), .QN(n10954) );
  INVX0 U11062 ( .INP(n10955), .ZN(n7662) );
  AND4X1 U11063 ( .IN1(n10946), .IN2(n10911), .IN3(n10956), .IN4(n10957), .Q(
        n10920) );
  NAND2X0 U11064 ( .IN1(g3229), .IN2(n10914), .QN(n10957) );
  NAND2X0 U11065 ( .IN1(n10958), .IN2(n7882), .QN(n10956) );
  NAND2X0 U11066 ( .IN1(n10947), .IN2(n10959), .QN(n10958) );
  INVX0 U11067 ( .INP(n10960), .ZN(n10959) );
  NAND2X0 U11068 ( .IN1(n10853), .IN2(n10912), .QN(n10947) );
  INVX0 U11069 ( .INP(n10948), .ZN(n10853) );
  NAND3X0 U11070 ( .IN1(n10852), .IN2(g3229), .IN3(n10960), .QN(n10911) );
  NOR2X0 U11071 ( .IN1(n10914), .IN2(n10949), .QN(n10960) );
  INVX0 U11072 ( .INP(n10913), .ZN(n10949) );
  NAND3X0 U11073 ( .IN1(n10961), .IN2(n10962), .IN3(n10963), .QN(n10914) );
  NAND2X0 U11074 ( .IN1(n6924), .IN2(n8537), .QN(n10963) );
  NAND2X0 U11075 ( .IN1(n6923), .IN2(n8861), .QN(n10962) );
  NAND2X0 U11076 ( .IN1(n6922), .IN2(n8500), .QN(n10961) );
  INVX0 U11077 ( .INP(n10912), .ZN(n10852) );
  NAND3X0 U11078 ( .IN1(n10964), .IN2(n10965), .IN3(n10966), .QN(n10912) );
  NAND2X0 U11079 ( .IN1(n6913), .IN2(n8537), .QN(n10966) );
  NAND2X0 U11080 ( .IN1(n6912), .IN2(n8861), .QN(n10965) );
  NAND2X0 U11081 ( .IN1(n6911), .IN2(n8500), .QN(n10964) );
  NAND3X0 U11082 ( .IN1(n10913), .IN2(n10948), .IN3(g3229), .QN(n10946) );
  NAND3X0 U11083 ( .IN1(n10967), .IN2(n10968), .IN3(n10969), .QN(n10948) );
  NAND2X0 U11084 ( .IN1(n6654), .IN2(n8537), .QN(n10969) );
  NAND2X0 U11085 ( .IN1(n6656), .IN2(n8861), .QN(n10968) );
  NAND2X0 U11086 ( .IN1(n6655), .IN2(n8500), .QN(n10967) );
  NAND3X0 U11087 ( .IN1(n10970), .IN2(n10971), .IN3(n10972), .QN(n10913) );
  NAND2X0 U11088 ( .IN1(n6935), .IN2(n8537), .QN(n10972) );
  NAND2X0 U11089 ( .IN1(n6934), .IN2(n8861), .QN(n10971) );
  OR2X1 U11090 ( .IN1(n4506), .IN2(test_so16), .Q(n10970) );
  AND3X1 U11091 ( .IN1(n10973), .IN2(n10974), .IN3(n10338), .Q(g27243) );
  NAND3X0 U11092 ( .IN1(n10975), .IN2(g2753), .IN3(test_so92), .QN(n10338) );
  OR2X1 U11093 ( .IN1(n10976), .IN2(g2753), .Q(n10973) );
  NOR2X0 U11094 ( .IN1(n10977), .IN2(n7269), .QN(n10976) );
  AND3X1 U11095 ( .IN1(n10978), .IN2(n9736), .IN3(n4522), .Q(g27131) );
  NAND2X0 U11096 ( .IN1(n6433), .IN2(n8313), .QN(n10978) );
  INVX0 U11097 ( .INP(n3683), .ZN(n8313) );
  AND3X1 U11098 ( .IN1(n10979), .IN2(n9739), .IN3(n4523), .Q(g27129) );
  NAND2X0 U11099 ( .IN1(n6434), .IN2(n8312), .QN(n10979) );
  INVX0 U11100 ( .INP(n3686), .ZN(n8312) );
  NOR3X0 U11101 ( .IN1(n10980), .IN2(n9322), .IN3(n10468), .QN(g27123) );
  INVX0 U11102 ( .INP(n3431), .ZN(n10468) );
  NAND2X0 U11103 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NOR2X0 U11104 ( .IN1(n3689), .IN2(g767), .QN(n10980) );
  AND3X1 U11105 ( .IN1(n10981), .IN2(n9743), .IN3(n4521), .Q(g27120) );
  OR2X1 U11106 ( .IN1(test_so15), .IN2(n3692), .Q(n10981) );
  NAND2X0 U11107 ( .IN1(n10982), .IN2(n10983), .QN(g26827) );
  NAND2X0 U11108 ( .IN1(n10984), .IN2(n4606), .QN(n10983) );
  NAND2X0 U11109 ( .IN1(n4509), .IN2(g2519), .QN(n10982) );
  NAND2X0 U11110 ( .IN1(n10985), .IN2(n10986), .QN(g26826) );
  NAND2X0 U11111 ( .IN1(n10984), .IN2(g7264), .QN(n10986) );
  NAND2X0 U11112 ( .IN1(n4524), .IN2(g2516), .QN(n10985) );
  NAND2X0 U11113 ( .IN1(n10987), .IN2(n10988), .QN(g26825) );
  NAND2X0 U11114 ( .IN1(n4606), .IN2(n10989), .QN(n10988) );
  NAND2X0 U11115 ( .IN1(n4509), .IN2(g2510), .QN(n10987) );
  NAND2X0 U11116 ( .IN1(n10990), .IN2(n10991), .QN(g26824) );
  NAND2X0 U11117 ( .IN1(n10992), .IN2(n4618), .QN(n10991) );
  NAND2X0 U11118 ( .IN1(test_so59), .IN2(n4511), .QN(n10990) );
  NAND2X0 U11119 ( .IN1(n10993), .IN2(n10994), .QN(g26823) );
  NAND2X0 U11120 ( .IN1(n10984), .IN2(g5555), .QN(n10994) );
  XOR2X1 U11121 ( .IN1(n10995), .IN2(n10376), .Q(n10984) );
  NAND3X0 U11122 ( .IN1(n10372), .IN2(n10996), .IN3(test_so79), .QN(n10995) );
  NAND2X0 U11123 ( .IN1(n10371), .IN2(n10373), .QN(n10996) );
  OR2X1 U11124 ( .IN1(test_so81), .IN2(n4509), .Q(n10373) );
  AND2X1 U11125 ( .IN1(n10997), .IN2(n10998), .Q(n10371) );
  NAND2X0 U11126 ( .IN1(n6937), .IN2(n8449), .QN(n10998) );
  NAND2X0 U11127 ( .IN1(n6946), .IN2(n8456), .QN(n10997) );
  NAND2X0 U11128 ( .IN1(n10999), .IN2(n11000), .QN(n10372) );
  NAND3X0 U11129 ( .IN1(n10376), .IN2(n10378), .IN3(n10383), .QN(n11000) );
  INVX0 U11130 ( .INP(n10381), .ZN(n10376) );
  NAND3X0 U11131 ( .IN1(n10382), .IN2(n10381), .IN3(n10379), .QN(n10999) );
  NAND2X0 U11132 ( .IN1(n4516), .IN2(g2513), .QN(n10993) );
  NAND2X0 U11133 ( .IN1(n11001), .IN2(n11002), .QN(g26822) );
  NAND2X0 U11134 ( .IN1(g7264), .IN2(n10989), .QN(n11002) );
  NAND2X0 U11135 ( .IN1(n4524), .IN2(g2507), .QN(n11001) );
  NAND2X0 U11136 ( .IN1(n11003), .IN2(n11004), .QN(g26821) );
  NAND2X0 U11137 ( .IN1(n10992), .IN2(g7014), .QN(n11004) );
  NAND2X0 U11138 ( .IN1(n4525), .IN2(g1822), .QN(n11003) );
  NAND2X0 U11139 ( .IN1(n11005), .IN2(n11006), .QN(g26820) );
  NAND2X0 U11140 ( .IN1(n4618), .IN2(n11007), .QN(n11006) );
  NAND2X0 U11141 ( .IN1(n4511), .IN2(g1816), .QN(n11005) );
  NAND2X0 U11142 ( .IN1(n11008), .IN2(n11009), .QN(g26818) );
  NAND2X0 U11143 ( .IN1(n4381), .IN2(g1131), .QN(n11009) );
  NAND2X0 U11144 ( .IN1(n11010), .IN2(g1088), .QN(n11008) );
  NAND2X0 U11145 ( .IN1(n11011), .IN2(n11012), .QN(g26817) );
  NAND2X0 U11146 ( .IN1(g5555), .IN2(n10989), .QN(n11012) );
  NAND2X0 U11147 ( .IN1(n11013), .IN2(n11014), .QN(n10989) );
  OR2X1 U11148 ( .IN1(n10379), .IN2(test_so79), .Q(n11014) );
  INVX0 U11149 ( .INP(n10383), .ZN(n10379) );
  NAND3X0 U11150 ( .IN1(n11015), .IN2(n11016), .IN3(n11017), .QN(n10383) );
  NAND2X0 U11151 ( .IN1(g5555), .IN2(g2504), .QN(n11017) );
  NAND2X0 U11152 ( .IN1(n4606), .IN2(g2510), .QN(n11016) );
  NAND2X0 U11153 ( .IN1(g7264), .IN2(g2507), .QN(n11015) );
  NAND2X0 U11154 ( .IN1(n10378), .IN2(test_so79), .QN(n11013) );
  INVX0 U11155 ( .INP(n10382), .ZN(n10378) );
  NAND2X0 U11156 ( .IN1(n9814), .IN2(n11018), .QN(n10382) );
  NAND3X0 U11157 ( .IN1(n11019), .IN2(n11020), .IN3(n11021), .QN(n11018) );
  NAND2X0 U11158 ( .IN1(n6849), .IN2(test_so73), .QN(n11021) );
  NAND2X0 U11159 ( .IN1(n6850), .IN2(g6837), .QN(n11020) );
  NAND2X0 U11160 ( .IN1(n6848), .IN2(g2241), .QN(n11019) );
  INVX0 U11161 ( .INP(n11022), .ZN(n9814) );
  NAND2X0 U11162 ( .IN1(n4516), .IN2(g2504), .QN(n11011) );
  NAND2X0 U11163 ( .IN1(n11023), .IN2(n11024), .QN(g26816) );
  NAND2X0 U11164 ( .IN1(n10992), .IN2(g5511), .QN(n11024) );
  XOR2X1 U11165 ( .IN1(n11025), .IN2(n10400), .Q(n10992) );
  NAND3X0 U11166 ( .IN1(n11026), .IN2(g1690), .IN3(n10396), .QN(n11025) );
  NAND2X0 U11167 ( .IN1(n11027), .IN2(n11028), .QN(n10396) );
  NAND3X0 U11168 ( .IN1(n10400), .IN2(n10402), .IN3(n10407), .QN(n11028) );
  INVX0 U11169 ( .INP(n10405), .ZN(n10400) );
  NAND3X0 U11170 ( .IN1(n10406), .IN2(n10405), .IN3(n10403), .QN(n11027) );
  INVX0 U11171 ( .INP(n10407), .ZN(n10403) );
  NAND2X0 U11172 ( .IN1(n10395), .IN2(n10397), .QN(n11026) );
  NAND2X0 U11173 ( .IN1(n6940), .IN2(n8459), .QN(n10397) );
  AND2X1 U11174 ( .IN1(n11029), .IN2(n11030), .Q(n10395) );
  NAND2X0 U11175 ( .IN1(n6950), .IN2(n8453), .QN(n11030) );
  NAND2X0 U11176 ( .IN1(n6951), .IN2(n8494), .QN(n11029) );
  NAND2X0 U11177 ( .IN1(n4518), .IN2(g1819), .QN(n11023) );
  NAND2X0 U11178 ( .IN1(n11031), .IN2(n11032), .QN(g26815) );
  NAND2X0 U11179 ( .IN1(g7014), .IN2(n11007), .QN(n11032) );
  NAND2X0 U11180 ( .IN1(n4525), .IN2(g1813), .QN(n11031) );
  NAND2X0 U11181 ( .IN1(n11033), .IN2(n11034), .QN(g26814) );
  NAND2X0 U11182 ( .IN1(n4364), .IN2(g1128), .QN(n11034) );
  NAND2X0 U11183 ( .IN1(n11010), .IN2(g6712), .QN(n11033) );
  NAND2X0 U11184 ( .IN1(n11035), .IN2(n11036), .QN(g26813) );
  NAND2X0 U11185 ( .IN1(n4381), .IN2(g1122), .QN(n11036) );
  NAND2X0 U11186 ( .IN1(n11037), .IN2(g1088), .QN(n11035) );
  NAND2X0 U11187 ( .IN1(n11038), .IN2(n11039), .QN(g26812) );
  NAND2X0 U11188 ( .IN1(n11040), .IN2(n4640), .QN(n11039) );
  NAND2X0 U11189 ( .IN1(n4506), .IN2(g444), .QN(n11038) );
  NAND2X0 U11190 ( .IN1(n11041), .IN2(n11042), .QN(g26811) );
  NAND2X0 U11191 ( .IN1(g5511), .IN2(n11007), .QN(n11042) );
  NAND2X0 U11192 ( .IN1(n11043), .IN2(n11044), .QN(n11007) );
  NAND2X0 U11193 ( .IN1(n4386), .IN2(n10407), .QN(n11044) );
  NAND3X0 U11194 ( .IN1(n11045), .IN2(n11046), .IN3(n11047), .QN(n10407) );
  NAND2X0 U11195 ( .IN1(g5511), .IN2(g1810), .QN(n11047) );
  NAND2X0 U11196 ( .IN1(n4618), .IN2(g1816), .QN(n11046) );
  NAND2X0 U11197 ( .IN1(g7014), .IN2(g1813), .QN(n11045) );
  NAND2X0 U11198 ( .IN1(n10402), .IN2(g1690), .QN(n11043) );
  INVX0 U11199 ( .INP(n10406), .ZN(n10402) );
  NAND2X0 U11200 ( .IN1(n9852), .IN2(n11048), .QN(n10406) );
  NAND3X0 U11201 ( .IN1(n11049), .IN2(n11050), .IN3(n11051), .QN(n11048) );
  NAND2X0 U11202 ( .IN1(n6861), .IN2(g6782), .QN(n11051) );
  NAND2X0 U11203 ( .IN1(n6862), .IN2(g6573), .QN(n11050) );
  NAND2X0 U11204 ( .IN1(n6860), .IN2(g1547), .QN(n11049) );
  INVX0 U11205 ( .INP(n11052), .ZN(n9852) );
  NAND2X0 U11206 ( .IN1(n4518), .IN2(g1810), .QN(n11041) );
  NAND2X0 U11207 ( .IN1(n11053), .IN2(n11054), .QN(g26810) );
  NAND2X0 U11208 ( .IN1(n4363), .IN2(g1125), .QN(n11054) );
  NAND2X0 U11209 ( .IN1(n11010), .IN2(g5472), .QN(n11053) );
  XOR2X1 U11210 ( .IN1(n11055), .IN2(n10424), .Q(n11010) );
  NAND3X0 U11211 ( .IN1(n11056), .IN2(g996), .IN3(n10420), .QN(n11055) );
  NAND2X0 U11212 ( .IN1(n11057), .IN2(n11058), .QN(n10420) );
  NAND3X0 U11213 ( .IN1(n10424), .IN2(n10426), .IN3(n10431), .QN(n11058) );
  INVX0 U11214 ( .INP(n10429), .ZN(n10424) );
  NAND3X0 U11215 ( .IN1(n10430), .IN2(n10429), .IN3(n10427), .QN(n11057) );
  INVX0 U11216 ( .INP(n10431), .ZN(n10427) );
  NAND2X0 U11217 ( .IN1(n10419), .IN2(n10421), .QN(n11056) );
  NAND2X0 U11218 ( .IN1(n6943), .IN2(g6712), .QN(n10421) );
  AND2X1 U11219 ( .IN1(n11059), .IN2(n11060), .Q(n10419) );
  NAND2X0 U11220 ( .IN1(n6956), .IN2(g1088), .QN(n11060) );
  NAND2X0 U11221 ( .IN1(n6957), .IN2(g5472), .QN(n11059) );
  NAND2X0 U11222 ( .IN1(n11061), .IN2(n11062), .QN(g26809) );
  NAND2X0 U11223 ( .IN1(n11037), .IN2(g6712), .QN(n11062) );
  NAND2X0 U11224 ( .IN1(n4364), .IN2(test_so38), .QN(n11061) );
  NAND2X0 U11225 ( .IN1(n11063), .IN2(n11064), .QN(g26808) );
  NAND2X0 U11226 ( .IN1(n11040), .IN2(g6447), .QN(n11064) );
  NAND2X0 U11227 ( .IN1(n4499), .IN2(g441), .QN(n11063) );
  NAND2X0 U11228 ( .IN1(n11065), .IN2(n11066), .QN(g26807) );
  NAND2X0 U11229 ( .IN1(n4640), .IN2(n11067), .QN(n11066) );
  NAND2X0 U11230 ( .IN1(n4506), .IN2(g435), .QN(n11065) );
  NAND2X0 U11231 ( .IN1(n11068), .IN2(n11069), .QN(g26806) );
  NAND2X0 U11232 ( .IN1(n4363), .IN2(g1116), .QN(n11069) );
  NAND2X0 U11233 ( .IN1(n11037), .IN2(g5472), .QN(n11068) );
  NAND2X0 U11234 ( .IN1(n11070), .IN2(n11071), .QN(n11037) );
  NAND2X0 U11235 ( .IN1(n4387), .IN2(n10431), .QN(n11071) );
  NAND3X0 U11236 ( .IN1(n11072), .IN2(n11073), .IN3(n11074), .QN(n10431) );
  NAND2X0 U11237 ( .IN1(g1088), .IN2(g1122), .QN(n11074) );
  NAND2X0 U11238 ( .IN1(g5472), .IN2(g1116), .QN(n11073) );
  NAND2X0 U11239 ( .IN1(test_so38), .IN2(g6712), .QN(n11072) );
  NAND2X0 U11240 ( .IN1(n10426), .IN2(g996), .QN(n11070) );
  INVX0 U11241 ( .INP(n10430), .ZN(n10426) );
  NAND2X0 U11242 ( .IN1(n9884), .IN2(n11075), .QN(n10430) );
  NAND3X0 U11243 ( .IN1(n11076), .IN2(n11077), .IN3(n11078), .QN(n11075) );
  NAND2X0 U11244 ( .IN1(n6871), .IN2(test_so31), .QN(n11078) );
  NAND2X0 U11245 ( .IN1(n6872), .IN2(g6518), .QN(n11077) );
  NAND2X0 U11246 ( .IN1(n6873), .IN2(g6368), .QN(n11076) );
  INVX0 U11247 ( .INP(n11079), .ZN(n9884) );
  NAND2X0 U11248 ( .IN1(n11080), .IN2(n11081), .QN(g26805) );
  NAND2X0 U11249 ( .IN1(n11040), .IN2(g5437), .QN(n11081) );
  XOR2X1 U11250 ( .IN1(n11082), .IN2(n10443), .Q(n11040) );
  NAND3X0 U11251 ( .IN1(n11083), .IN2(g309), .IN3(n10439), .QN(n11082) );
  NAND2X0 U11252 ( .IN1(n11084), .IN2(n11085), .QN(n10439) );
  NAND3X0 U11253 ( .IN1(n10443), .IN2(n10445), .IN3(n10450), .QN(n11085) );
  INVX0 U11254 ( .INP(n10448), .ZN(n10443) );
  NAND3X0 U11255 ( .IN1(n10449), .IN2(n10448), .IN3(n10446), .QN(n11084) );
  INVX0 U11256 ( .INP(n10450), .ZN(n10446) );
  NAND2X0 U11257 ( .IN1(n10438), .IN2(n10440), .QN(n11083) );
  NAND2X0 U11258 ( .IN1(n6963), .IN2(n8500), .QN(n10440) );
  AND2X1 U11259 ( .IN1(n11086), .IN2(n11087), .Q(n10438) );
  NAND2X0 U11260 ( .IN1(n6964), .IN2(n8861), .QN(n11087) );
  NAND2X0 U11261 ( .IN1(n6965), .IN2(n8537), .QN(n11086) );
  NAND2X0 U11262 ( .IN1(n4520), .IN2(g438), .QN(n11080) );
  NAND2X0 U11263 ( .IN1(n11088), .IN2(n11089), .QN(g26804) );
  NAND2X0 U11264 ( .IN1(g6447), .IN2(n11067), .QN(n11089) );
  NAND2X0 U11265 ( .IN1(n4499), .IN2(g432), .QN(n11088) );
  NAND2X0 U11266 ( .IN1(n11090), .IN2(n11091), .QN(g26803) );
  NAND2X0 U11267 ( .IN1(g5437), .IN2(n11067), .QN(n11091) );
  NAND2X0 U11268 ( .IN1(n11092), .IN2(n11093), .QN(n11067) );
  NAND2X0 U11269 ( .IN1(n4388), .IN2(n10450), .QN(n11093) );
  NAND3X0 U11270 ( .IN1(n11094), .IN2(n11095), .IN3(n11096), .QN(n10450) );
  NAND2X0 U11271 ( .IN1(g5437), .IN2(g429), .QN(n11096) );
  NAND2X0 U11272 ( .IN1(n4640), .IN2(g435), .QN(n11095) );
  NAND2X0 U11273 ( .IN1(g6447), .IN2(g432), .QN(n11094) );
  NAND2X0 U11274 ( .IN1(n10445), .IN2(g309), .QN(n11092) );
  INVX0 U11275 ( .INP(n10449), .ZN(n10445) );
  NAND2X0 U11276 ( .IN1(n9911), .IN2(n11097), .QN(n10449) );
  NAND3X0 U11277 ( .IN1(n11098), .IN2(n11099), .IN3(n11100), .QN(n11097) );
  NAND2X0 U11278 ( .IN1(n6883), .IN2(g6313), .QN(n11100) );
  NAND2X0 U11279 ( .IN1(n6884), .IN2(g6231), .QN(n11099) );
  NAND2X0 U11280 ( .IN1(n6882), .IN2(g165), .QN(n11098) );
  INVX0 U11281 ( .INP(n11101), .ZN(n9911) );
  NAND2X0 U11282 ( .IN1(n4520), .IN2(g429), .QN(n11090) );
  NOR2X0 U11283 ( .IN1(n7777), .IN2(n11102), .QN(g26798) );
  XNOR2X1 U11284 ( .IN1(n4355), .IN2(n11103), .Q(n11102) );
  NAND2X0 U11285 ( .IN1(n11104), .IN2(g2900), .QN(n11103) );
  NOR2X0 U11286 ( .IN1(n10335), .IN2(n11105), .QN(g26795) );
  XOR2X1 U11287 ( .IN1(n10977), .IN2(test_so92), .Q(n11105) );
  NOR2X0 U11288 ( .IN1(n10339), .IN2(n11106), .QN(g26789) );
  XOR2X1 U11289 ( .IN1(g2046), .IN2(n10455), .Q(n11106) );
  INVX0 U11290 ( .INP(n11107), .ZN(n10455) );
  NOR2X0 U11291 ( .IN1(n11108), .IN2(n11109), .QN(g26786) );
  XNOR2X1 U11292 ( .IN1(n6429), .IN2(n3741), .Q(n11108) );
  NOR2X0 U11293 ( .IN1(n10343), .IN2(n11110), .QN(g26781) );
  XNOR2X1 U11294 ( .IN1(n4469), .IN2(n10458), .Q(n11110) );
  NOR2X0 U11295 ( .IN1(n9912), .IN2(n11111), .QN(g26776) );
  XOR2X1 U11296 ( .IN1(n10464), .IN2(test_so28), .Q(n11111) );
  NOR3X0 U11297 ( .IN1(n11112), .IN2(n10335), .IN3(n10975), .QN(g26677) );
  INVX0 U11298 ( .INP(n10977), .ZN(n10975) );
  NAND3X0 U11299 ( .IN1(g2734), .IN2(g2746), .IN3(n11113), .QN(n10977) );
  NOR2X0 U11300 ( .IN1(n11114), .IN2(g2746), .QN(n11112) );
  NOR2X0 U11301 ( .IN1(n4397), .IN2(n11115), .QN(n11114) );
  NAND2X0 U11302 ( .IN1(n11116), .IN2(n11117), .QN(g26676) );
  NAND2X0 U11303 ( .IN1(n11118), .IN2(g2479), .QN(n11117) );
  NAND2X0 U11304 ( .IN1(n11119), .IN2(n8449), .QN(n11118) );
  NAND2X0 U11305 ( .IN1(n11120), .IN2(n8449), .QN(n11116) );
  NAND2X0 U11306 ( .IN1(n11121), .IN2(n11122), .QN(g26675) );
  NAND2X0 U11307 ( .IN1(n11123), .IN2(g1783), .QN(n11122) );
  NAND2X0 U11308 ( .IN1(n11124), .IN2(n8453), .QN(n11123) );
  NAND2X0 U11309 ( .IN1(n11125), .IN2(n8453), .QN(n11121) );
  NAND2X0 U11310 ( .IN1(n11126), .IN2(n11127), .QN(g26672) );
  NAND2X0 U11311 ( .IN1(n11128), .IN2(g2478), .QN(n11127) );
  NAND2X0 U11312 ( .IN1(n11119), .IN2(n8456), .QN(n11128) );
  NAND2X0 U11313 ( .IN1(n11120), .IN2(n8456), .QN(n11126) );
  NOR3X0 U11314 ( .IN1(n11129), .IN2(n10339), .IN3(n11107), .QN(g26671) );
  NOR3X0 U11315 ( .IN1(n4399), .IN2(n4409), .IN3(n11130), .QN(n11107) );
  NOR2X0 U11316 ( .IN1(n11131), .IN2(g2052), .QN(n11129) );
  NOR2X0 U11317 ( .IN1(n4399), .IN2(n11130), .QN(n11131) );
  INVX0 U11318 ( .INP(n11132), .ZN(n11130) );
  NAND2X0 U11319 ( .IN1(n11133), .IN2(n11134), .QN(g26670) );
  NAND2X0 U11320 ( .IN1(n11135), .IN2(g1785), .QN(n11134) );
  NAND2X0 U11321 ( .IN1(n11124), .IN2(n8459), .QN(n11135) );
  NAND2X0 U11322 ( .IN1(n11125), .IN2(n8459), .QN(n11133) );
  NAND2X0 U11323 ( .IN1(n11136), .IN2(n11137), .QN(g26669) );
  NAND2X0 U11324 ( .IN1(n11138), .IN2(g1089), .QN(n11137) );
  NAND2X0 U11325 ( .IN1(n11139), .IN2(g1088), .QN(n11138) );
  NAND2X0 U11326 ( .IN1(n11140), .IN2(g1088), .QN(n11136) );
  NAND2X0 U11327 ( .IN1(n11141), .IN2(n11142), .QN(g26667) );
  NAND2X0 U11328 ( .IN1(test_so60), .IN2(n11143), .QN(n11142) );
  NAND2X0 U11329 ( .IN1(n11124), .IN2(n8494), .QN(n11143) );
  NAND2X0 U11330 ( .IN1(n11125), .IN2(n8494), .QN(n11141) );
  NOR2X0 U11331 ( .IN1(n11124), .IN2(n4386), .QN(n11125) );
  INVX0 U11332 ( .INP(n3751), .ZN(n11124) );
  NAND3X0 U11333 ( .IN1(n11144), .IN2(g1690), .IN3(n8489), .QN(n3751) );
  AND4X1 U11334 ( .IN1(n11145), .IN2(n11146), .IN3(n11147), .IN4(n11148), .Q(
        n8489) );
  NOR4X0 U11335 ( .IN1(n11149), .IN2(n11150), .IN3(n8901), .IN4(n11151), .QN(
        n11148) );
  XOR2X1 U11336 ( .IN1(g1496), .IN2(n11152), .Q(n11151) );
  NAND3X0 U11337 ( .IN1(n11153), .IN2(n11154), .IN3(n11155), .QN(n11152) );
  NAND2X0 U11338 ( .IN1(n7184), .IN2(g6782), .QN(n11155) );
  NAND2X0 U11339 ( .IN1(n7185), .IN2(g6573), .QN(n11154) );
  NAND2X0 U11340 ( .IN1(n6803), .IN2(g1547), .QN(n11153) );
  INVX0 U11341 ( .INP(n3070), .ZN(n8901) );
  XOR2X1 U11342 ( .IN1(g1506), .IN2(n11156), .Q(n11150) );
  NAND3X0 U11343 ( .IN1(n11157), .IN2(n11158), .IN3(n11159), .QN(n11156) );
  NAND2X0 U11344 ( .IN1(n7181), .IN2(g6782), .QN(n11159) );
  NAND2X0 U11345 ( .IN1(n7182), .IN2(g6573), .QN(n11158) );
  NAND2X0 U11346 ( .IN1(n6801), .IN2(g1547), .QN(n11157) );
  NAND3X0 U11347 ( .IN1(n11160), .IN2(n11161), .IN3(n11162), .QN(n11149) );
  XOR2X1 U11348 ( .IN1(n11163), .IN2(n4326), .Q(n11162) );
  NAND3X0 U11349 ( .IN1(n11164), .IN2(n11165), .IN3(n11166), .QN(n11163) );
  NAND2X0 U11350 ( .IN1(n7186), .IN2(g6782), .QN(n11166) );
  NAND2X0 U11351 ( .IN1(n7187), .IN2(g6573), .QN(n11165) );
  NAND2X0 U11352 ( .IN1(n6804), .IN2(g1547), .QN(n11164) );
  XOR2X1 U11353 ( .IN1(n11167), .IN2(n4390), .Q(n11161) );
  NAND3X0 U11354 ( .IN1(n11168), .IN2(n11169), .IN3(n11170), .QN(n11167) );
  NAND2X0 U11355 ( .IN1(n7188), .IN2(g6782), .QN(n11170) );
  NAND2X0 U11356 ( .IN1(n7189), .IN2(g6573), .QN(n11169) );
  NAND2X0 U11357 ( .IN1(n6805), .IN2(g1547), .QN(n11168) );
  XOR2X1 U11358 ( .IN1(n11171), .IN2(n4374), .Q(n11160) );
  NAND3X0 U11359 ( .IN1(n11172), .IN2(n11173), .IN3(n11174), .QN(n11171) );
  NAND2X0 U11360 ( .IN1(n7192), .IN2(g6782), .QN(n11174) );
  OR2X1 U11361 ( .IN1(n4317), .IN2(test_so52), .Q(n11173) );
  NAND2X0 U11362 ( .IN1(n6807), .IN2(g1547), .QN(n11172) );
  NOR3X0 U11363 ( .IN1(n11175), .IN2(n11176), .IN3(n11177), .QN(n11147) );
  XOR2X1 U11364 ( .IN1(g1501), .IN2(n11178), .Q(n11177) );
  NAND3X0 U11365 ( .IN1(n11179), .IN2(n11180), .IN3(n11181), .QN(n11178) );
  OR2X1 U11366 ( .IN1(n4515), .IN2(test_so53), .Q(n11181) );
  NAND2X0 U11367 ( .IN1(n7183), .IN2(g6573), .QN(n11180) );
  NAND2X0 U11368 ( .IN1(n6802), .IN2(g1547), .QN(n11179) );
  XOR2X1 U11369 ( .IN1(g1481), .IN2(n11182), .Q(n11176) );
  NAND3X0 U11370 ( .IN1(n11183), .IN2(n11184), .IN3(n11185), .QN(n11182) );
  NAND2X0 U11371 ( .IN1(n7190), .IN2(g6782), .QN(n11185) );
  NAND2X0 U11372 ( .IN1(n7191), .IN2(g6573), .QN(n11184) );
  NAND2X0 U11373 ( .IN1(n6806), .IN2(g1547), .QN(n11183) );
  XOR2X1 U11374 ( .IN1(n8756), .IN2(n11186), .Q(n11175) );
  NAND3X0 U11375 ( .IN1(n11187), .IN2(n11188), .IN3(n11189), .QN(n11186) );
  NAND2X0 U11376 ( .IN1(n6783), .IN2(g6782), .QN(n11189) );
  NAND2X0 U11377 ( .IN1(n6784), .IN2(g6573), .QN(n11188) );
  NAND2X0 U11378 ( .IN1(n6782), .IN2(g1547), .QN(n11187) );
  XOR2X1 U11379 ( .IN1(n11190), .IN2(n8603), .Q(n11146) );
  NAND3X0 U11380 ( .IN1(n11191), .IN2(n11192), .IN3(n11193), .QN(n11190) );
  NAND2X0 U11381 ( .IN1(n6799), .IN2(g6782), .QN(n11193) );
  NAND2X0 U11382 ( .IN1(n6800), .IN2(g6573), .QN(n11192) );
  NAND2X0 U11383 ( .IN1(n6798), .IN2(g1547), .QN(n11191) );
  XOR2X1 U11384 ( .IN1(n11194), .IN2(n4378), .Q(n11145) );
  NAND3X0 U11385 ( .IN1(n11195), .IN2(n11196), .IN3(n11197), .QN(n11194) );
  NAND2X0 U11386 ( .IN1(n7193), .IN2(g6782), .QN(n11197) );
  NAND2X0 U11387 ( .IN1(n7194), .IN2(g6573), .QN(n11196) );
  NAND2X0 U11388 ( .IN1(n6808), .IN2(g1547), .QN(n11195) );
  INVX0 U11389 ( .INP(n9293), .ZN(n11144) );
  NAND3X0 U11390 ( .IN1(n11198), .IN2(n11199), .IN3(n11200), .QN(n9293) );
  NAND2X0 U11391 ( .IN1(n6939), .IN2(n8459), .QN(n11200) );
  NAND2X0 U11392 ( .IN1(n6949), .IN2(n8453), .QN(n11199) );
  OR2X1 U11393 ( .IN1(n4518), .IN2(test_so60), .Q(n11198) );
  AND3X1 U11394 ( .IN1(n11201), .IN2(n11202), .IN3(n10458), .Q(g26666) );
  NAND3X0 U11395 ( .IN1(g1346), .IN2(g1358), .IN3(n11203), .QN(n10458) );
  OR2X1 U11396 ( .IN1(n11204), .IN2(g1358), .Q(n11201) );
  AND2X1 U11397 ( .IN1(g1346), .IN2(n11203), .Q(n11204) );
  NAND2X0 U11398 ( .IN1(n11205), .IN2(n11206), .QN(g26665) );
  NAND2X0 U11399 ( .IN1(n11207), .IN2(g1091), .QN(n11206) );
  NAND2X0 U11400 ( .IN1(n11139), .IN2(g6712), .QN(n11207) );
  NAND2X0 U11401 ( .IN1(n11140), .IN2(g6712), .QN(n11205) );
  NAND2X0 U11402 ( .IN1(n11208), .IN2(n11209), .QN(g26664) );
  NAND2X0 U11403 ( .IN1(n11210), .IN2(g402), .QN(n11209) );
  NAND2X0 U11404 ( .IN1(n11211), .IN2(n8500), .QN(n11210) );
  NAND2X0 U11405 ( .IN1(n11212), .IN2(n8500), .QN(n11208) );
  NAND2X0 U11406 ( .IN1(n11213), .IN2(n11214), .QN(g26661) );
  NAND2X0 U11407 ( .IN1(n11215), .IN2(g1090), .QN(n11214) );
  NAND2X0 U11408 ( .IN1(n11139), .IN2(g5472), .QN(n11215) );
  NAND2X0 U11409 ( .IN1(n11140), .IN2(g5472), .QN(n11213) );
  NOR2X0 U11410 ( .IN1(n11139), .IN2(n4387), .QN(n11140) );
  INVX0 U11411 ( .INP(n3758), .ZN(n11139) );
  NAND3X0 U11412 ( .IN1(n9197), .IN2(g996), .IN3(n11216), .QN(n3758) );
  INVX0 U11413 ( .INP(n9305), .ZN(n11216) );
  NAND3X0 U11414 ( .IN1(n11217), .IN2(n11218), .IN3(n11219), .QN(n9305) );
  NAND2X0 U11415 ( .IN1(n6954), .IN2(g1088), .QN(n11219) );
  NAND2X0 U11416 ( .IN1(n6955), .IN2(g5472), .QN(n11218) );
  NAND2X0 U11417 ( .IN1(n6942), .IN2(g6712), .QN(n11217) );
  AND4X1 U11418 ( .IN1(n11220), .IN2(n11221), .IN3(n11222), .IN4(n11223), .Q(
        n9197) );
  NOR4X0 U11419 ( .IN1(n11224), .IN2(n11225), .IN3(n11226), .IN4(n11227), .QN(
        n11223) );
  XOR2X1 U11420 ( .IN1(n8790), .IN2(n11228), .Q(n11227) );
  NAND3X0 U11421 ( .IN1(n11229), .IN2(n11230), .IN3(n11231), .QN(n11228) );
  NAND2X0 U11422 ( .IN1(n6812), .IN2(test_so31), .QN(n11231) );
  NAND2X0 U11423 ( .IN1(n6813), .IN2(g6518), .QN(n11230) );
  NAND2X0 U11424 ( .IN1(n6814), .IN2(g6368), .QN(n11229) );
  XNOR2X1 U11425 ( .IN1(n4391), .IN2(n11232), .Q(n11226) );
  NAND3X0 U11426 ( .IN1(n11233), .IN2(n11234), .IN3(n11235), .QN(n11232) );
  NAND2X0 U11427 ( .IN1(n6819), .IN2(test_so31), .QN(n11235) );
  NAND2X0 U11428 ( .IN1(n7202), .IN2(g6518), .QN(n11234) );
  NAND2X0 U11429 ( .IN1(n7203), .IN2(g6368), .QN(n11233) );
  XOR2X1 U11430 ( .IN1(g801), .IN2(n11236), .Q(n11225) );
  NAND3X0 U11431 ( .IN1(n11237), .IN2(n11238), .IN3(n11239), .QN(n11236) );
  NAND2X0 U11432 ( .IN1(n6818), .IN2(test_so31), .QN(n11239) );
  NAND2X0 U11433 ( .IN1(n7200), .IN2(g6518), .QN(n11238) );
  NAND2X0 U11434 ( .IN1(n7201), .IN2(g6368), .QN(n11237) );
  NAND3X0 U11435 ( .IN1(n11240), .IN2(n3102), .IN3(n11241), .QN(n11224) );
  XOR2X1 U11436 ( .IN1(n11242), .IN2(n4289), .Q(n11241) );
  NAND3X0 U11437 ( .IN1(n11243), .IN2(n11244), .IN3(n11245), .QN(n11242) );
  NAND2X0 U11438 ( .IN1(n6815), .IN2(test_so31), .QN(n11245) );
  NAND2X0 U11439 ( .IN1(n7195), .IN2(g6518), .QN(n11244) );
  NAND2X0 U11440 ( .IN1(n7196), .IN2(g6368), .QN(n11243) );
  XOR2X1 U11441 ( .IN1(n11246), .IN2(n4559), .Q(n11240) );
  NAND3X0 U11442 ( .IN1(n11247), .IN2(n11248), .IN3(n11249), .QN(n11246) );
  NAND2X0 U11443 ( .IN1(test_so31), .IN2(n6817), .QN(n11249) );
  NAND2X0 U11444 ( .IN1(n7199), .IN2(g6518), .QN(n11248) );
  OR2X1 U11445 ( .IN1(n4323), .IN2(test_so32), .Q(n11247) );
  NOR3X0 U11446 ( .IN1(n11250), .IN2(n11251), .IN3(n11252), .QN(n11222) );
  XOR2X1 U11447 ( .IN1(g809), .IN2(n11253), .Q(n11252) );
  NAND3X0 U11448 ( .IN1(n11254), .IN2(n11255), .IN3(n11256), .QN(n11253) );
  NAND2X0 U11449 ( .IN1(n6816), .IN2(test_so31), .QN(n11256) );
  NAND2X0 U11450 ( .IN1(n7197), .IN2(g6518), .QN(n11255) );
  NAND2X0 U11451 ( .IN1(n7198), .IN2(g6368), .QN(n11254) );
  XOR2X1 U11452 ( .IN1(n9883), .IN2(n11257), .Q(n11251) );
  NAND3X0 U11453 ( .IN1(n11258), .IN2(n11259), .IN3(n11260), .QN(n11257) );
  NAND2X0 U11454 ( .IN1(n6809), .IN2(test_so31), .QN(n11260) );
  NAND2X0 U11455 ( .IN1(n6810), .IN2(g6518), .QN(n11259) );
  NAND2X0 U11456 ( .IN1(n6811), .IN2(g6368), .QN(n11258) );
  XNOR2X1 U11457 ( .IN1(n4375), .IN2(n11261), .Q(n11250) );
  NAND3X0 U11458 ( .IN1(n11262), .IN2(n11263), .IN3(n11264), .QN(n11261) );
  NAND2X0 U11459 ( .IN1(n6821), .IN2(test_so31), .QN(n11264) );
  NAND2X0 U11460 ( .IN1(n7206), .IN2(g6518), .QN(n11263) );
  NAND2X0 U11461 ( .IN1(n7207), .IN2(g6368), .QN(n11262) );
  XOR2X1 U11462 ( .IN1(n11265), .IN2(n4379), .Q(n11221) );
  NAND3X0 U11463 ( .IN1(n11266), .IN2(n11267), .IN3(n11268), .QN(n11265) );
  NAND2X0 U11464 ( .IN1(n6822), .IN2(test_so31), .QN(n11268) );
  NAND2X0 U11465 ( .IN1(n7208), .IN2(g6518), .QN(n11267) );
  NAND2X0 U11466 ( .IN1(n7209), .IN2(g6368), .QN(n11266) );
  XOR2X1 U11467 ( .IN1(n11269), .IN2(n4321), .Q(n11220) );
  NAND3X0 U11468 ( .IN1(n11270), .IN2(n11271), .IN3(n11272), .QN(n11269) );
  NAND2X0 U11469 ( .IN1(n6820), .IN2(test_so31), .QN(n11272) );
  NAND2X0 U11470 ( .IN1(n7204), .IN2(g6518), .QN(n11271) );
  NAND2X0 U11471 ( .IN1(n7205), .IN2(g6368), .QN(n11270) );
  NOR3X0 U11472 ( .IN1(n11273), .IN2(n9912), .IN3(n10462), .QN(g26660) );
  INVX0 U11473 ( .INP(n10464), .ZN(n10462) );
  NAND3X0 U11474 ( .IN1(g660), .IN2(g672), .IN3(n11274), .QN(n10464) );
  NOR2X0 U11475 ( .IN1(n11275), .IN2(g672), .QN(n11273) );
  NOR2X0 U11476 ( .IN1(n4403), .IN2(n11276), .QN(n11275) );
  NAND2X0 U11477 ( .IN1(n11277), .IN2(n11278), .QN(g26659) );
  NAND2X0 U11478 ( .IN1(n11279), .IN2(g404), .QN(n11278) );
  NAND2X0 U11479 ( .IN1(n11211), .IN2(n8861), .QN(n11279) );
  NAND2X0 U11480 ( .IN1(n11212), .IN2(n8861), .QN(n11277) );
  NAND2X0 U11481 ( .IN1(n11280), .IN2(n11281), .QN(g26655) );
  NAND2X0 U11482 ( .IN1(n11282), .IN2(g403), .QN(n11281) );
  NAND2X0 U11483 ( .IN1(n11211), .IN2(n8537), .QN(n11282) );
  NAND2X0 U11484 ( .IN1(n11212), .IN2(n8537), .QN(n11280) );
  NOR2X0 U11485 ( .IN1(n11211), .IN2(n4388), .QN(n11212) );
  INVX0 U11486 ( .INP(n3788), .ZN(n11211) );
  NAND3X0 U11487 ( .IN1(n11283), .IN2(g309), .IN3(n8532), .QN(n3788) );
  AND4X1 U11488 ( .IN1(n11284), .IN2(n11285), .IN3(n11286), .IN4(n11287), .Q(
        n8532) );
  NOR4X0 U11489 ( .IN1(n11288), .IN2(n11289), .IN3(n8873), .IN4(n11290), .QN(
        n11287) );
  XOR2X1 U11490 ( .IN1(g117), .IN2(n11291), .Q(n11290) );
  NAND3X0 U11491 ( .IN1(n11292), .IN2(n11293), .IN3(n11294), .QN(n11291) );
  NAND2X0 U11492 ( .IN1(n7214), .IN2(g6313), .QN(n11294) );
  NAND2X0 U11493 ( .IN1(n7215), .IN2(g6231), .QN(n11293) );
  NAND2X0 U11494 ( .IN1(n6827), .IN2(g165), .QN(n11292) );
  INVX0 U11495 ( .INP(n3130), .ZN(n8873) );
  XOR2X1 U11496 ( .IN1(g125), .IN2(n11295), .Q(n11289) );
  NAND3X0 U11497 ( .IN1(n11296), .IN2(n11297), .IN3(n11298), .QN(n11295) );
  NAND2X0 U11498 ( .IN1(n7210), .IN2(g6313), .QN(n11298) );
  NAND2X0 U11499 ( .IN1(n7211), .IN2(g6231), .QN(n11297) );
  NAND2X0 U11500 ( .IN1(n6825), .IN2(g165), .QN(n11296) );
  NAND3X0 U11501 ( .IN1(n11299), .IN2(n11300), .IN3(n11301), .QN(n11288) );
  XOR2X1 U11502 ( .IN1(n11302), .IN2(n4328), .Q(n11301) );
  NAND3X0 U11503 ( .IN1(n11303), .IN2(n11304), .IN3(n11305), .QN(n11302) );
  NAND2X0 U11504 ( .IN1(n7216), .IN2(g6313), .QN(n11305) );
  NAND2X0 U11505 ( .IN1(n7217), .IN2(g6231), .QN(n11304) );
  NAND2X0 U11506 ( .IN1(n6828), .IN2(g165), .QN(n11303) );
  XOR2X1 U11507 ( .IN1(n11306), .IN2(n4392), .Q(n11300) );
  NAND3X0 U11508 ( .IN1(n11307), .IN2(n11308), .IN3(n11309), .QN(n11306) );
  NAND2X0 U11509 ( .IN1(n7218), .IN2(g6313), .QN(n11309) );
  NAND2X0 U11510 ( .IN1(n7219), .IN2(g6231), .QN(n11308) );
  OR2X1 U11511 ( .IN1(n4369), .IN2(test_so11), .Q(n11307) );
  XOR2X1 U11512 ( .IN1(n11310), .IN2(n11311), .Q(n11299) );
  NAND3X0 U11513 ( .IN1(n11312), .IN2(n11313), .IN3(n11314), .QN(n11310) );
  NAND2X0 U11514 ( .IN1(n6786), .IN2(g6313), .QN(n11314) );
  NAND2X0 U11515 ( .IN1(n6787), .IN2(g6231), .QN(n11313) );
  NAND2X0 U11516 ( .IN1(n6785), .IN2(g165), .QN(n11312) );
  NOR3X0 U11517 ( .IN1(n11315), .IN2(n11316), .IN3(n11317), .QN(n11286) );
  XOR2X1 U11518 ( .IN1(g121), .IN2(n11318), .Q(n11317) );
  NAND3X0 U11519 ( .IN1(n11319), .IN2(n11320), .IN3(n11321), .QN(n11318) );
  NAND2X0 U11520 ( .IN1(n7212), .IN2(g6313), .QN(n11321) );
  NAND2X0 U11521 ( .IN1(n7213), .IN2(g6231), .QN(n11320) );
  NAND2X0 U11522 ( .IN1(n6826), .IN2(g165), .QN(n11319) );
  XOR2X1 U11523 ( .IN1(n9910), .IN2(n11322), .Q(n11316) );
  NAND3X0 U11524 ( .IN1(n11323), .IN2(n11324), .IN3(n11325), .QN(n11322) );
  NAND2X0 U11525 ( .IN1(n6824), .IN2(g6313), .QN(n11325) );
  OR2X1 U11526 ( .IN1(n4318), .IN2(test_so12), .Q(n11324) );
  NAND2X0 U11527 ( .IN1(n6823), .IN2(g165), .QN(n11323) );
  XNOR2X1 U11528 ( .IN1(n4376), .IN2(n11326), .Q(n11315) );
  NAND3X0 U11529 ( .IN1(n11327), .IN2(n11328), .IN3(n11329), .QN(n11326) );
  NAND2X0 U11530 ( .IN1(n7222), .IN2(g6313), .QN(n11329) );
  NAND2X0 U11531 ( .IN1(n7223), .IN2(g6231), .QN(n11328) );
  NAND2X0 U11532 ( .IN1(n6830), .IN2(g165), .QN(n11327) );
  XOR2X1 U11533 ( .IN1(n11330), .IN2(n4380), .Q(n11285) );
  NAND3X0 U11534 ( .IN1(n11331), .IN2(n11332), .IN3(n11333), .QN(n11330) );
  NAND2X0 U11535 ( .IN1(n7224), .IN2(g6313), .QN(n11333) );
  NAND2X0 U11536 ( .IN1(n7225), .IN2(g6231), .QN(n11332) );
  NAND2X0 U11537 ( .IN1(n6831), .IN2(g165), .QN(n11331) );
  XOR2X1 U11538 ( .IN1(n11334), .IN2(n4322), .Q(n11284) );
  NAND3X0 U11539 ( .IN1(n11335), .IN2(n11336), .IN3(n11337), .QN(n11334) );
  NAND2X0 U11540 ( .IN1(n7220), .IN2(g6313), .QN(n11337) );
  NAND2X0 U11541 ( .IN1(n7221), .IN2(g6231), .QN(n11336) );
  NAND2X0 U11542 ( .IN1(n6829), .IN2(g165), .QN(n11335) );
  INVX0 U11543 ( .INP(n9314), .ZN(n11283) );
  NAND3X0 U11544 ( .IN1(n11338), .IN2(n11339), .IN3(n11340), .QN(n9314) );
  NAND2X0 U11545 ( .IN1(n6962), .IN2(n8537), .QN(n11340) );
  NAND2X0 U11546 ( .IN1(n6961), .IN2(n8861), .QN(n11339) );
  NAND2X0 U11547 ( .IN1(n6960), .IN2(n8500), .QN(n11338) );
  NAND2X0 U11548 ( .IN1(n11341), .IN2(n11342), .QN(g26616) );
  NAND2X0 U11549 ( .IN1(n4299), .IN2(g2571), .QN(n11342) );
  NAND2X0 U11550 ( .IN1(n11343), .IN2(g2624), .QN(n11341) );
  NAND2X0 U11551 ( .IN1(n11344), .IN2(n11345), .QN(g26596) );
  NAND2X0 U11552 ( .IN1(n4370), .IN2(g2568), .QN(n11345) );
  NAND2X0 U11553 ( .IN1(n11343), .IN2(g7390), .QN(n11344) );
  NAND2X0 U11554 ( .IN1(n11346), .IN2(n11347), .QN(g26592) );
  NAND2X0 U11555 ( .IN1(n4366), .IN2(g1877), .QN(n11347) );
  NAND2X0 U11556 ( .IN1(n11348), .IN2(g1930), .QN(n11346) );
  NAND2X0 U11557 ( .IN1(n11349), .IN2(n11350), .QN(g26575) );
  NAND2X0 U11558 ( .IN1(n4314), .IN2(g2565), .QN(n11350) );
  NAND2X0 U11559 ( .IN1(n11343), .IN2(n9246), .QN(n11349) );
  NOR3X0 U11560 ( .IN1(n7994), .IN2(n4303), .IN3(n11351), .QN(n11343) );
  NAND2X0 U11561 ( .IN1(n11352), .IN2(n11353), .QN(g26573) );
  NAND2X0 U11562 ( .IN1(n4315), .IN2(g1874), .QN(n11353) );
  NAND2X0 U11563 ( .IN1(n11348), .IN2(g7194), .QN(n11352) );
  NAND2X0 U11564 ( .IN1(n11354), .IN2(n11355), .QN(g26569) );
  NAND2X0 U11565 ( .IN1(n4300), .IN2(g1183), .QN(n11355) );
  NAND2X0 U11566 ( .IN1(n11356), .IN2(g1236), .QN(n11354) );
  NAND2X0 U11567 ( .IN1(n11357), .IN2(n11358), .QN(g26559) );
  NAND2X0 U11568 ( .IN1(n11348), .IN2(n9268), .QN(n11358) );
  NOR3X0 U11569 ( .IN1(n8181), .IN2(n4297), .IN3(n11359), .QN(n11348) );
  NAND2X0 U11570 ( .IN1(test_so68), .IN2(n4296), .QN(n11357) );
  NAND2X0 U11571 ( .IN1(n11360), .IN2(n11361), .QN(g26557) );
  NAND2X0 U11572 ( .IN1(n4316), .IN2(g1180), .QN(n11361) );
  NAND2X0 U11573 ( .IN1(n11356), .IN2(g6944), .QN(n11360) );
  NAND2X0 U11574 ( .IN1(n11362), .IN2(n11363), .QN(g26553) );
  NAND2X0 U11575 ( .IN1(n4313), .IN2(g496), .QN(n11363) );
  NAND2X0 U11576 ( .IN1(n11364), .IN2(g550), .QN(n11362) );
  NAND2X0 U11577 ( .IN1(n11365), .IN2(n11366), .QN(g26547) );
  NAND2X0 U11578 ( .IN1(n11356), .IN2(n10142), .QN(n11366) );
  NOR3X0 U11579 ( .IN1(n8278), .IN2(n4304), .IN3(n11367), .QN(n11356) );
  NAND2X0 U11580 ( .IN1(test_so47), .IN2(n4371), .QN(n11365) );
  NAND2X0 U11581 ( .IN1(n11368), .IN2(n11369), .QN(g26545) );
  NAND2X0 U11582 ( .IN1(n4372), .IN2(g493), .QN(n11369) );
  NAND2X0 U11583 ( .IN1(n11364), .IN2(g6642), .QN(n11368) );
  NAND2X0 U11584 ( .IN1(n11370), .IN2(n11371), .QN(g26541) );
  NAND2X0 U11585 ( .IN1(n4298), .IN2(g490), .QN(n11371) );
  NAND2X0 U11586 ( .IN1(n11364), .IN2(n10242), .QN(n11370) );
  NOR3X0 U11587 ( .IN1(n7271), .IN2(n7844), .IN3(n11372), .QN(n11364) );
  NOR2X0 U11588 ( .IN1(n9318), .IN2(n11373), .QN(g26532) );
  XNOR2X1 U11589 ( .IN1(n4526), .IN2(n6981), .Q(n11373) );
  NOR2X0 U11590 ( .IN1(n9320), .IN2(n11374), .QN(g26531) );
  XNOR2X1 U11591 ( .IN1(n4527), .IN2(n6985), .Q(n11374) );
  NOR2X0 U11592 ( .IN1(n9322), .IN2(n11375), .QN(g26530) );
  XOR2X1 U11593 ( .IN1(n6989), .IN2(n11376), .Q(n11375) );
  NOR2X0 U11594 ( .IN1(n9324), .IN2(n11377), .QN(g26529) );
  XNOR2X1 U11595 ( .IN1(n4528), .IN2(n6993), .Q(n11377) );
  AND2X1 U11596 ( .IN1(n11378), .IN2(n11379), .Q(g26183) );
  NAND2X0 U11597 ( .IN1(n4432), .IN2(n8017), .QN(n11379) );
  NAND2X0 U11598 ( .IN1(n11380), .IN2(g986), .QN(n11378) );
  NAND2X0 U11599 ( .IN1(n11381), .IN2(n11382), .QN(n11380) );
  NAND2X0 U11600 ( .IN1(n4364), .IN2(n6997), .QN(n11382) );
  OR2X1 U11601 ( .IN1(g21346), .IN2(n4364), .Q(n11381) );
  NAND4X0 U11602 ( .IN1(n3700), .IN2(n11383), .IN3(n11384), .IN4(n11385), .QN(
        g26149) );
  NOR4X0 U11603 ( .IN1(n11386), .IN2(n11387), .IN3(n11388), .IN4(n11389), .QN(
        n11385) );
  NOR2X0 U11604 ( .IN1(n4441), .IN2(n11390), .QN(n11389) );
  NOR2X0 U11605 ( .IN1(n4338), .IN2(n11391), .QN(n11388) );
  NOR2X0 U11606 ( .IN1(n10488), .IN2(DFF_156_n1), .QN(n11387) );
  NAND3X0 U11607 ( .IN1(n11392), .IN2(n11393), .IN3(n11394), .QN(n11386) );
  NAND2X0 U11608 ( .IN1(n3936), .IN2(n11395), .QN(n11394) );
  NAND4X0 U11609 ( .IN1(n11396), .IN2(n11397), .IN3(n11398), .IN4(n11399), 
        .QN(n11395) );
  NAND2X0 U11610 ( .IN1(n11400), .IN2(g3088), .QN(n11399) );
  NAND2X0 U11611 ( .IN1(n11401), .IN2(g3164), .QN(n11398) );
  NAND2X0 U11612 ( .IN1(n11402), .IN2(g3158), .QN(n11397) );
  NAND2X0 U11613 ( .IN1(n10483), .IN2(g3182), .QN(n11396) );
  NAND2X0 U11614 ( .IN1(n11403), .IN2(g3167), .QN(n11393) );
  NAND2X0 U11615 ( .IN1(n3939), .IN2(n11404), .QN(n11392) );
  NAND3X0 U11616 ( .IN1(n11405), .IN2(n11406), .IN3(n11407), .QN(n11404) );
  NAND2X0 U11617 ( .IN1(n3940), .IN2(g3185), .QN(n11407) );
  NAND2X0 U11618 ( .IN1(test_so8), .IN2(n10478), .QN(n11406) );
  NAND2X0 U11619 ( .IN1(n11408), .IN2(g3155), .QN(n11405) );
  NOR3X0 U11620 ( .IN1(n11409), .IN2(n11410), .IN3(n11411), .QN(n11384) );
  NOR2X0 U11621 ( .IN1(n4444), .IN2(n11412), .QN(n11411) );
  NOR2X0 U11622 ( .IN1(n4450), .IN2(n11413), .QN(n11410) );
  NOR2X0 U11623 ( .IN1(n11414), .IN2(DFF_149_n1), .QN(n11409) );
  NAND2X0 U11624 ( .IN1(n10489), .IN2(n8086), .QN(n11383) );
  NAND2X0 U11625 ( .IN1(n11415), .IN2(n11416), .QN(g26135) );
  NOR4X0 U11626 ( .IN1(n11417), .IN2(n11418), .IN3(n11419), .IN4(n11420), .QN(
        n11416) );
  NOR2X0 U11627 ( .IN1(n4447), .IN2(n11391), .QN(n11420) );
  NOR2X0 U11628 ( .IN1(n11421), .IN2(n11422), .QN(n11419) );
  INVX0 U11629 ( .INP(n3936), .ZN(n11422) );
  NOR4X0 U11630 ( .IN1(n11423), .IN2(n11424), .IN3(n11425), .IN4(n11426), .QN(
        n11421) );
  NOR2X0 U11631 ( .IN1(n4438), .IN2(n11427), .QN(n11426) );
  NOR2X0 U11632 ( .IN1(n4434), .IN2(n11428), .QN(n11425) );
  AND2X1 U11633 ( .IN1(g3100), .IN2(n11401), .Q(n11424) );
  AND2X1 U11634 ( .IN1(g3108), .IN2(n11400), .Q(n11423) );
  NOR2X0 U11635 ( .IN1(n4343), .IN2(n11390), .QN(n11418) );
  NAND4X0 U11636 ( .IN1(n11429), .IN2(n11430), .IN3(n11431), .IN4(n11432), 
        .QN(n11417) );
  NAND2X0 U11637 ( .IN1(test_so10), .IN2(n10487), .QN(n11432) );
  NAND2X0 U11638 ( .IN1(test_so7), .IN2(n11403), .QN(n11431) );
  OR2X1 U11639 ( .IN1(n10476), .IN2(n11433), .Q(n11430) );
  NAND2X0 U11640 ( .IN1(n3939), .IN2(n11434), .QN(n11429) );
  NAND3X0 U11641 ( .IN1(n11435), .IN2(n11436), .IN3(n11437), .QN(n11434) );
  NAND2X0 U11642 ( .IN1(n3940), .IN2(g3107), .QN(n11437) );
  NAND2X0 U11643 ( .IN1(n10478), .IN2(g3105), .QN(n11436) );
  NAND2X0 U11644 ( .IN1(n11408), .IN2(g3097), .QN(n11435) );
  NOR4X0 U11645 ( .IN1(n11438), .IN2(n11439), .IN3(n11440), .IN4(n11441), .QN(
        n11415) );
  NOR2X0 U11646 ( .IN1(n4452), .IN2(n11413), .QN(n11441) );
  NOR2X0 U11647 ( .IN1(n10488), .IN2(DFF_155_n1), .QN(n11440) );
  NOR2X0 U11648 ( .IN1(n4443), .IN2(n11412), .QN(n11439) );
  NAND3X0 U11649 ( .IN1(n11442), .IN2(n11443), .IN3(n3700), .QN(n11438) );
  NAND2X0 U11650 ( .IN1(n11444), .IN2(n8081), .QN(n11443) );
  NAND2X0 U11651 ( .IN1(n6894), .IN2(n10489), .QN(n11442) );
  NAND2X0 U11652 ( .IN1(n11445), .IN2(n11446), .QN(g26104) );
  NOR4X0 U11653 ( .IN1(n11447), .IN2(n11448), .IN3(n11449), .IN4(n11450), .QN(
        n11446) );
  NOR2X0 U11654 ( .IN1(n4448), .IN2(n11391), .QN(n11450) );
  NAND3X0 U11655 ( .IN1(n10477), .IN2(n4406), .IN3(n3933), .QN(n11391) );
  NOR2X0 U11656 ( .IN1(n11451), .IN2(n10476), .QN(n11449) );
  NAND2X0 U11657 ( .IN1(n3705), .IN2(n11408), .QN(n10476) );
  INVX0 U11658 ( .INP(n10481), .ZN(n11451) );
  NOR2X0 U11659 ( .IN1(n4344), .IN2(n11390), .QN(n11448) );
  NAND2X0 U11660 ( .IN1(n11452), .IN2(n4329), .QN(n11390) );
  NAND4X0 U11661 ( .IN1(n11453), .IN2(n11454), .IN3(n11455), .IN4(n11456), 
        .QN(n11447) );
  NAND2X0 U11662 ( .IN1(n10487), .IN2(g3142), .QN(n11456) );
  AND3X1 U11663 ( .IN1(n3940), .IN2(g3204), .IN3(n4073), .Q(n10487) );
  NAND2X0 U11664 ( .IN1(n11403), .IN2(g3086), .QN(n11455) );
  AND2X1 U11665 ( .IN1(n10477), .IN2(n11408), .Q(n11403) );
  NAND2X0 U11666 ( .IN1(n3939), .IN2(n11457), .QN(n11454) );
  NAND3X0 U11667 ( .IN1(n11458), .IN2(n11459), .IN3(n11460), .QN(n11457) );
  NAND2X0 U11668 ( .IN1(n3940), .IN2(g3095), .QN(n11460) );
  NAND2X0 U11669 ( .IN1(n10478), .IN2(g3093), .QN(n11459) );
  NAND2X0 U11670 ( .IN1(test_so6), .IN2(n11408), .QN(n11458) );
  NAND2X0 U11671 ( .IN1(n3936), .IN2(n11461), .QN(n11453) );
  NAND4X0 U11672 ( .IN1(n11462), .IN2(n11463), .IN3(n11464), .IN4(n11465), 
        .QN(n11461) );
  NAND2X0 U11673 ( .IN1(n11400), .IN2(g3096), .QN(n11465) );
  NOR2X0 U11674 ( .IN1(n4329), .IN2(n4406), .QN(n11400) );
  NAND2X0 U11675 ( .IN1(n11401), .IN2(g3085), .QN(n11464) );
  NOR2X0 U11676 ( .IN1(g3201), .IN2(n4329), .QN(n11401) );
  NAND2X0 U11677 ( .IN1(n11402), .IN2(g3211), .QN(n11463) );
  INVX0 U11678 ( .INP(n11428), .ZN(n11402) );
  NAND2X0 U11679 ( .IN1(n10483), .IN2(g3094), .QN(n11462) );
  INVX0 U11680 ( .INP(n11427), .ZN(n10483) );
  NOR4X0 U11681 ( .IN1(n11466), .IN2(n11467), .IN3(n11468), .IN4(n11469), .QN(
        n11445) );
  NOR2X0 U11682 ( .IN1(n4451), .IN2(n11413), .QN(n11469) );
  NAND2X0 U11683 ( .IN1(n11452), .IN2(g3207), .QN(n11413) );
  AND3X1 U11684 ( .IN1(n4406), .IN2(g3188), .IN3(n10477), .Q(n11452) );
  AND2X1 U11685 ( .IN1(n3938), .IN2(g3204), .Q(n10477) );
  AND2X1 U11686 ( .IN1(n3944), .IN2(g3197), .Q(n3938) );
  AND3X1 U11687 ( .IN1(DFF_132_n1), .IN2(DFF_131_n1), .IN3(DFF_134_n1), .Q(
        n3944) );
  NOR2X0 U11688 ( .IN1(n13233), .IN2(n10488), .QN(n11468) );
  NAND3X0 U11689 ( .IN1(n10478), .IN2(g3204), .IN3(n4073), .QN(n10488) );
  NOR2X0 U11690 ( .IN1(n11427), .IN2(g3188), .QN(n10478) );
  NAND2X0 U11691 ( .IN1(n4329), .IN2(g3201), .QN(n11427) );
  NOR2X0 U11692 ( .IN1(n4445), .IN2(n11412), .QN(n11467) );
  NAND3X0 U11693 ( .IN1(n3939), .IN2(n4406), .IN3(n3933), .QN(n11412) );
  NOR2X0 U11694 ( .IN1(g3188), .IN2(n4329), .QN(n3933) );
  NAND3X0 U11695 ( .IN1(n11470), .IN2(n11471), .IN3(n3700), .QN(n11466) );
  NAND2X0 U11696 ( .IN1(n11444), .IN2(n8082), .QN(n11471) );
  NAND2X0 U11697 ( .IN1(n10489), .IN2(n8087), .QN(n11470) );
  NAND2X0 U11698 ( .IN1(n7825), .IN2(n11472), .QN(g26048) );
  NAND2X0 U11699 ( .IN1(n11473), .IN2(n11474), .QN(n11472) );
  XOR2X1 U11700 ( .IN1(n7909), .IN2(n11475), .Q(n11473) );
  NOR2X0 U11701 ( .IN1(n7777), .IN2(n11476), .QN(g26037) );
  XOR2X1 U11702 ( .IN1(n4291), .IN2(n11104), .Q(n11476) );
  NOR2X0 U11703 ( .IN1(n11477), .IN2(n11109), .QN(g26031) );
  XOR2X1 U11704 ( .IN1(test_so98), .IN2(n3742), .Q(n11477) );
  NAND2X0 U11705 ( .IN1(n11478), .IN2(n11479), .QN(g26025) );
  NAND2X0 U11706 ( .IN1(test_so82), .IN2(n11480), .QN(n11479) );
  NAND2X0 U11707 ( .IN1(n11119), .IN2(n8841), .QN(n11480) );
  INVX0 U11708 ( .INP(n3749), .ZN(n11119) );
  NAND2X0 U11709 ( .IN1(n11120), .IN2(n8841), .QN(n11478) );
  AND2X1 U11710 ( .IN1(test_so79), .IN2(n3749), .Q(n11120) );
  NAND3X0 U11711 ( .IN1(n9121), .IN2(n11481), .IN3(test_so79), .QN(n3749) );
  INVX0 U11712 ( .INP(n9281), .ZN(n11481) );
  NAND3X0 U11713 ( .IN1(n11482), .IN2(n11483), .IN3(n11484), .QN(n9281) );
  NAND2X0 U11714 ( .IN1(n6936), .IN2(n8449), .QN(n11484) );
  OR2X1 U11715 ( .IN1(n4509), .IN2(test_so82), .Q(n11483) );
  NAND2X0 U11716 ( .IN1(n6945), .IN2(n8456), .QN(n11482) );
  AND4X1 U11717 ( .IN1(n11485), .IN2(n11486), .IN3(n11487), .IN4(n11488), .Q(
        n9121) );
  NOR4X0 U11718 ( .IN1(n11489), .IN2(n11490), .IN3(n11491), .IN4(n11492), .QN(
        n11488) );
  XOR2X1 U11719 ( .IN1(n8719), .IN2(n11493), .Q(n11492) );
  NAND3X0 U11720 ( .IN1(n11494), .IN2(n11495), .IN3(n11496), .QN(n11493) );
  NAND2X0 U11721 ( .IN1(n6780), .IN2(test_so73), .QN(n11496) );
  NAND2X0 U11722 ( .IN1(n6781), .IN2(g6837), .QN(n11495) );
  NAND2X0 U11723 ( .IN1(n6779), .IN2(g2241), .QN(n11494) );
  XOR2X1 U11724 ( .IN1(g2180), .IN2(n11497), .Q(n11491) );
  NAND3X0 U11725 ( .IN1(n11498), .IN2(n11499), .IN3(n11500), .QN(n11497) );
  NAND2X0 U11726 ( .IN1(n7173), .IN2(test_so73), .QN(n11500) );
  NAND2X0 U11727 ( .IN1(n7174), .IN2(g6837), .QN(n11499) );
  NAND2X0 U11728 ( .IN1(n6794), .IN2(g2241), .QN(n11498) );
  XOR2X1 U11729 ( .IN1(g2185), .IN2(n11501), .Q(n11490) );
  NAND3X0 U11730 ( .IN1(n11502), .IN2(n11503), .IN3(n11504), .QN(n11501) );
  OR2X1 U11731 ( .IN1(n7266), .IN2(test_so74), .Q(n11504) );
  NAND2X0 U11732 ( .IN1(n7172), .IN2(g6837), .QN(n11503) );
  NAND2X0 U11733 ( .IN1(n6793), .IN2(g2241), .QN(n11502) );
  NAND3X0 U11734 ( .IN1(n11505), .IN2(n3038), .IN3(n11506), .QN(n11489) );
  XOR2X1 U11735 ( .IN1(n11507), .IN2(n4287), .Q(n11506) );
  NAND3X0 U11736 ( .IN1(n11508), .IN2(n11509), .IN3(n11510), .QN(n11507) );
  NAND2X0 U11737 ( .IN1(n7166), .IN2(test_so73), .QN(n11510) );
  NAND2X0 U11738 ( .IN1(n7167), .IN2(g6837), .QN(n11509) );
  NAND2X0 U11739 ( .IN1(n6790), .IN2(g2241), .QN(n11508) );
  XOR2X1 U11740 ( .IN1(n11511), .IN2(n4555), .Q(n11505) );
  NAND3X0 U11741 ( .IN1(n11512), .IN2(n11513), .IN3(n11514), .QN(n11511) );
  NAND2X0 U11742 ( .IN1(n7170), .IN2(test_so73), .QN(n11514) );
  NAND2X0 U11743 ( .IN1(n7171), .IN2(g6837), .QN(n11513) );
  NAND2X0 U11744 ( .IN1(n6792), .IN2(g2241), .QN(n11512) );
  NOR3X0 U11745 ( .IN1(n11515), .IN2(n11516), .IN3(n11517), .QN(n11487) );
  XOR2X1 U11746 ( .IN1(g2195), .IN2(n11518), .Q(n11517) );
  NAND3X0 U11747 ( .IN1(n11519), .IN2(n11520), .IN3(n11521), .QN(n11518) );
  NAND2X0 U11748 ( .IN1(n7168), .IN2(test_so73), .QN(n11521) );
  NAND2X0 U11749 ( .IN1(n7169), .IN2(g6837), .QN(n11520) );
  NAND2X0 U11750 ( .IN1(n6791), .IN2(g2241), .QN(n11519) );
  XOR2X1 U11751 ( .IN1(n9813), .IN2(n11522), .Q(n11516) );
  NAND3X0 U11752 ( .IN1(n11523), .IN2(n11524), .IN3(n11525), .QN(n11522) );
  OR2X1 U11753 ( .IN1(n7266), .IN2(test_so75), .Q(n11525) );
  NAND2X0 U11754 ( .IN1(n6789), .IN2(g6837), .QN(n11524) );
  NAND2X0 U11755 ( .IN1(n6788), .IN2(g2241), .QN(n11523) );
  XOR2X1 U11756 ( .IN1(g2170), .IN2(n11526), .Q(n11515) );
  NAND3X0 U11757 ( .IN1(n11527), .IN2(n11528), .IN3(n11529), .QN(n11526) );
  NAND2X0 U11758 ( .IN1(n7177), .IN2(test_so73), .QN(n11529) );
  NAND2X0 U11759 ( .IN1(n7178), .IN2(g6837), .QN(n11528) );
  NAND2X0 U11760 ( .IN1(n6796), .IN2(g2241), .QN(n11527) );
  XOR2X1 U11761 ( .IN1(n11530), .IN2(n4377), .Q(n11486) );
  NAND3X0 U11762 ( .IN1(n11531), .IN2(n11532), .IN3(n11533), .QN(n11530) );
  NAND2X0 U11763 ( .IN1(n7179), .IN2(test_so73), .QN(n11533) );
  NAND2X0 U11764 ( .IN1(n7180), .IN2(g6837), .QN(n11532) );
  NAND2X0 U11765 ( .IN1(n6797), .IN2(g2241), .QN(n11531) );
  XOR2X1 U11766 ( .IN1(n11534), .IN2(n4319), .Q(n11485) );
  NAND3X0 U11767 ( .IN1(n11535), .IN2(n11536), .IN3(n11537), .QN(n11534) );
  NAND2X0 U11768 ( .IN1(n7175), .IN2(test_so73), .QN(n11537) );
  NAND2X0 U11769 ( .IN1(n7176), .IN2(g6837), .QN(n11536) );
  NAND2X0 U11770 ( .IN1(n6795), .IN2(g2241), .QN(n11535) );
  AND3X1 U11771 ( .IN1(n11538), .IN2(n9736), .IN3(n4526), .Q(g25940) );
  OR2X1 U11772 ( .IN1(test_so78), .IN2(n3887), .Q(n11538) );
  AND3X1 U11773 ( .IN1(n11539), .IN2(n9739), .IN3(n4527), .Q(g25938) );
  OR2X1 U11774 ( .IN1(g1462), .IN2(n3890), .Q(n11539) );
  NOR3X0 U11775 ( .IN1(n11540), .IN2(n9322), .IN3(n11376), .QN(g25935) );
  INVX0 U11776 ( .INP(n3690), .ZN(n11376) );
  NAND2X0 U11777 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NOR2X0 U11778 ( .IN1(n3893), .IN2(g776), .QN(n11540) );
  AND3X1 U11779 ( .IN1(n11541), .IN2(n9743), .IN3(n4528), .Q(g25932) );
  OR2X1 U11780 ( .IN1(g88), .IN2(n3896), .Q(n11541) );
  NAND2X0 U11781 ( .IN1(n11542), .IN2(n11543), .QN(g25489) );
  NAND2X0 U11782 ( .IN1(n11544), .IN2(n7274), .QN(n11543) );
  NAND2X0 U11783 ( .IN1(n11545), .IN2(n11546), .QN(n11544) );
  NAND2X0 U11784 ( .IN1(n4424), .IN2(n11547), .QN(n11546) );
  NAND2X0 U11785 ( .IN1(n11433), .IN2(g3142), .QN(n11547) );
  INVX0 U11786 ( .INP(n10482), .ZN(n11433) );
  NAND2X0 U11787 ( .IN1(n6709), .IN2(n6708), .QN(n10482) );
  NAND2X0 U11788 ( .IN1(n4301), .IN2(n10481), .QN(n11545) );
  NAND2X0 U11789 ( .IN1(DFF_15_n1), .IN2(DFF_16_n1), .QN(n10481) );
  NAND4X0 U11790 ( .IN1(g3151), .IN2(g3097), .IN3(g3142), .IN4(test_so10), 
        .QN(n11542) );
  NAND2X0 U11791 ( .IN1(n11548), .IN2(n11549), .QN(g25452) );
  OR2X1 U11792 ( .IN1(g3109), .IN2(n4443), .Q(n11549) );
  NAND2X0 U11793 ( .IN1(g21851), .IN2(g3109), .QN(n11548) );
  NAND2X0 U11794 ( .IN1(n11550), .IN2(n11551), .QN(g25451) );
  OR2X1 U11795 ( .IN1(g8030), .IN2(n4434), .Q(n11551) );
  NAND2X0 U11796 ( .IN1(g21851), .IN2(g8030), .QN(n11550) );
  NAND2X0 U11797 ( .IN1(n11552), .IN2(n11553), .QN(g25450) );
  NAND2X0 U11798 ( .IN1(n4382), .IN2(g3097), .QN(n11553) );
  NAND2X0 U11799 ( .IN1(g21851), .IN2(g8106), .QN(n11552) );
  NAND3X0 U11800 ( .IN1(n11554), .IN2(n11555), .IN3(n3700), .QN(g25442) );
  NAND2X0 U11801 ( .IN1(n11444), .IN2(g3111), .QN(n11555) );
  NAND2X0 U11802 ( .IN1(n10489), .IN2(g3124), .QN(n11554) );
  NAND3X0 U11803 ( .IN1(n11556), .IN2(n11557), .IN3(n3700), .QN(g25435) );
  NAND2X0 U11804 ( .IN1(n11444), .IN2(g3110), .QN(n11557) );
  NAND2X0 U11805 ( .IN1(n10489), .IN2(DFF_144_n1), .QN(n11556) );
  NAND3X0 U11806 ( .IN1(n11558), .IN2(n11559), .IN3(n3700), .QN(g25420) );
  NAND2X0 U11807 ( .IN1(n11444), .IN2(g3112), .QN(n11559) );
  INVX0 U11808 ( .INP(n11414), .ZN(n11444) );
  NAND3X0 U11809 ( .IN1(n11408), .IN2(g3204), .IN3(n4073), .QN(n11414) );
  NOR2X0 U11810 ( .IN1(n11428), .IN2(g3188), .QN(n11408) );
  NAND2X0 U11811 ( .IN1(n4406), .IN2(n4329), .QN(n11428) );
  NAND2X0 U11812 ( .IN1(test_so9), .IN2(n10489), .QN(n11558) );
  NAND2X0 U11813 ( .IN1(n11560), .IN2(n11561), .QN(g25288) );
  NAND2X0 U11814 ( .IN1(n11562), .IN2(n11563), .QN(n11561) );
  OR2X1 U11815 ( .IN1(n11563), .IN2(n6775), .Q(n11560) );
  NAND2X0 U11816 ( .IN1(n11564), .IN2(n11565), .QN(g25280) );
  NAND2X0 U11817 ( .IN1(n11566), .IN2(n11562), .QN(n11565) );
  OR2X1 U11818 ( .IN1(n11566), .IN2(n6767), .Q(n11564) );
  NAND2X0 U11819 ( .IN1(n11567), .IN2(n11568), .QN(g25279) );
  NAND2X0 U11820 ( .IN1(n11569), .IN2(n11570), .QN(n11568) );
  OR2X1 U11821 ( .IN1(n11570), .IN2(n6776), .Q(n11567) );
  NAND2X0 U11822 ( .IN1(n11571), .IN2(n11572), .QN(g25272) );
  NAND2X0 U11823 ( .IN1(n11573), .IN2(n11562), .QN(n11572) );
  AND4X1 U11824 ( .IN1(n11574), .IN2(n11575), .IN3(n11576), .IN4(n11577), .Q(
        n11562) );
  NAND2X0 U11825 ( .IN1(n6896), .IN2(g2703), .QN(n11577) );
  NOR2X0 U11826 ( .IN1(n11578), .IN2(n11579), .QN(n11576) );
  NOR4X0 U11827 ( .IN1(n11580), .IN2(n11581), .IN3(n11582), .IN4(n11583), .QN(
        n11579) );
  XOR2X1 U11828 ( .IN1(n4419), .IN2(n8016), .Q(n11583) );
  INVX0 U11829 ( .INP(n8022), .ZN(n8016) );
  NAND3X0 U11830 ( .IN1(n11584), .IN2(n11585), .IN3(n11586), .QN(n8022) );
  NAND2X0 U11831 ( .IN1(n7064), .IN2(g7487), .QN(n11586) );
  NAND2X0 U11832 ( .IN1(n7129), .IN2(g2703), .QN(n11585) );
  NAND2X0 U11833 ( .IN1(n7065), .IN2(g7425), .QN(n11584) );
  XOR2X1 U11834 ( .IN1(n4472), .IN2(n8051), .Q(n11582) );
  INVX0 U11835 ( .INP(n8052), .ZN(n8051) );
  NAND3X0 U11836 ( .IN1(n11587), .IN2(n11588), .IN3(n11589), .QN(n8052) );
  NAND2X0 U11837 ( .IN1(n7066), .IN2(g7487), .QN(n11589) );
  NAND2X0 U11838 ( .IN1(n7130), .IN2(g2703), .QN(n11588) );
  NAND2X0 U11839 ( .IN1(n7067), .IN2(g7425), .QN(n11587) );
  NAND3X0 U11840 ( .IN1(n11590), .IN2(n11591), .IN3(n11592), .QN(n11581) );
  XOR2X1 U11841 ( .IN1(g2714), .IN2(n8048), .Q(n11592) );
  INVX0 U11842 ( .INP(n8041), .ZN(n8048) );
  NAND3X0 U11843 ( .IN1(n11593), .IN2(n11594), .IN3(n11595), .QN(n8041) );
  NAND2X0 U11844 ( .IN1(n7068), .IN2(g7487), .QN(n11595) );
  NAND2X0 U11845 ( .IN1(n7131), .IN2(g2703), .QN(n11594) );
  NAND2X0 U11846 ( .IN1(n7069), .IN2(g7425), .QN(n11593) );
  XOR2X1 U11847 ( .IN1(g2734), .IN2(n8064), .Q(n11591) );
  INVX0 U11848 ( .INP(n8063), .ZN(n8064) );
  NAND3X0 U11849 ( .IN1(n11596), .IN2(n11597), .IN3(n11598), .QN(n8063) );
  NAND2X0 U11850 ( .IN1(n7060), .IN2(g7487), .QN(n11598) );
  NAND2X0 U11851 ( .IN1(n7128), .IN2(g2703), .QN(n11597) );
  NAND2X0 U11852 ( .IN1(n7061), .IN2(g7425), .QN(n11596) );
  XOR2X1 U11853 ( .IN1(g2753), .IN2(n8034), .Q(n11590) );
  INVX0 U11854 ( .INP(n8035), .ZN(n8034) );
  NAND3X0 U11855 ( .IN1(n11599), .IN2(n11600), .IN3(n11601), .QN(n8035) );
  NAND2X0 U11856 ( .IN1(n7054), .IN2(g7487), .QN(n11601) );
  NAND2X0 U11857 ( .IN1(n7125), .IN2(g2703), .QN(n11600) );
  NAND2X0 U11858 ( .IN1(n7055), .IN2(g7425), .QN(n11599) );
  NAND4X0 U11859 ( .IN1(n11602), .IN2(n11603), .IN3(n11604), .IN4(n11605), 
        .QN(n11580) );
  XOR2X1 U11860 ( .IN1(n4415), .IN2(n7989), .Q(n11605) );
  NAND3X0 U11861 ( .IN1(n11606), .IN2(n11607), .IN3(n11608), .QN(n7989) );
  NAND2X0 U11862 ( .IN1(n7050), .IN2(g7487), .QN(n11608) );
  NAND2X0 U11863 ( .IN1(n7124), .IN2(g2703), .QN(n11607) );
  NAND2X0 U11864 ( .IN1(n7051), .IN2(g7425), .QN(n11606) );
  NOR2X0 U11865 ( .IN1(n11609), .IN2(n11610), .QN(n11604) );
  XOR2X1 U11866 ( .IN1(n4393), .IN2(n7993), .Q(n11610) );
  INVX0 U11867 ( .INP(n7996), .ZN(n7993) );
  NAND3X0 U11868 ( .IN1(n11611), .IN2(n11612), .IN3(n11613), .QN(n7996) );
  NAND2X0 U11869 ( .IN1(n7052), .IN2(g7487), .QN(n11613) );
  OR2X1 U11870 ( .IN1(n4292), .IN2(test_so94), .Q(n11612) );
  NAND2X0 U11871 ( .IN1(n7053), .IN2(g7425), .QN(n11611) );
  XOR2X1 U11872 ( .IN1(n7269), .IN2(n8071), .Q(n11609) );
  INVX0 U11873 ( .INP(n8069), .ZN(n8071) );
  NAND3X0 U11874 ( .IN1(n11614), .IN2(n11615), .IN3(n11616), .QN(n8069) );
  NAND2X0 U11875 ( .IN1(n7056), .IN2(g7487), .QN(n11616) );
  NAND2X0 U11876 ( .IN1(n7126), .IN2(g2703), .QN(n11615) );
  NAND2X0 U11877 ( .IN1(n7057), .IN2(g7425), .QN(n11614) );
  XOR2X1 U11878 ( .IN1(g2746), .IN2(n8012), .Q(n11603) );
  INVX0 U11879 ( .INP(n8013), .ZN(n8012) );
  NAND3X0 U11880 ( .IN1(n11617), .IN2(n11618), .IN3(n11619), .QN(n8013) );
  NAND2X0 U11881 ( .IN1(n7058), .IN2(g7487), .QN(n11619) );
  NAND2X0 U11882 ( .IN1(n7127), .IN2(g2703), .QN(n11618) );
  NAND2X0 U11883 ( .IN1(n7059), .IN2(g7425), .QN(n11617) );
  XOR2X1 U11884 ( .IN1(g2720), .IN2(n8030), .Q(n11602) );
  INVX0 U11885 ( .INP(n8031), .ZN(n8030) );
  NAND3X0 U11886 ( .IN1(n11620), .IN2(n11621), .IN3(n11622), .QN(n8031) );
  NAND2X0 U11887 ( .IN1(n7062), .IN2(g7487), .QN(n11622) );
  OR2X1 U11888 ( .IN1(n4292), .IN2(test_so93), .Q(n11621) );
  NAND2X0 U11889 ( .IN1(n7063), .IN2(g7425), .QN(n11620) );
  NOR2X0 U11890 ( .IN1(n4356), .IN2(g2804), .QN(n11578) );
  NAND2X0 U11891 ( .IN1(n6841), .IN2(g7425), .QN(n11575) );
  INVX0 U11892 ( .INP(n8402), .ZN(n11574) );
  NAND3X0 U11893 ( .IN1(n11623), .IN2(n11624), .IN3(n11625), .QN(n8402) );
  NAND2X0 U11894 ( .IN1(n6832), .IN2(g7487), .QN(n11625) );
  NAND2X0 U11895 ( .IN1(n6895), .IN2(g2703), .QN(n11624) );
  NAND2X0 U11896 ( .IN1(n6840), .IN2(g7425), .QN(n11623) );
  OR2X1 U11897 ( .IN1(n11573), .IN2(n6768), .Q(n11571) );
  NAND2X0 U11898 ( .IN1(n11626), .IN2(n11627), .QN(g25271) );
  NAND2X0 U11899 ( .IN1(n11628), .IN2(n11569), .QN(n11627) );
  OR2X1 U11900 ( .IN1(n11628), .IN2(n6769), .Q(n11626) );
  NAND2X0 U11901 ( .IN1(n11629), .IN2(n11630), .QN(g25270) );
  NAND2X0 U11902 ( .IN1(n11631), .IN2(n11632), .QN(n11630) );
  OR2X1 U11903 ( .IN1(n11632), .IN2(n6777), .Q(n11629) );
  NAND2X0 U11904 ( .IN1(n11633), .IN2(n11634), .QN(g25268) );
  NAND2X0 U11905 ( .IN1(n11635), .IN2(n11569), .QN(n11634) );
  AND4X1 U11906 ( .IN1(n11636), .IN2(n11637), .IN3(n11638), .IN4(n11639), .Q(
        n11569) );
  NAND2X0 U11907 ( .IN1(n6898), .IN2(g2009), .QN(n11639) );
  NOR2X0 U11908 ( .IN1(n11640), .IN2(n11641), .QN(n11638) );
  NOR4X0 U11909 ( .IN1(n11642), .IN2(n11643), .IN3(n11644), .IN4(n11645), .QN(
        n11641) );
  XOR2X1 U11910 ( .IN1(n4400), .IN2(n8180), .Q(n11645) );
  INVX0 U11911 ( .INP(n8178), .ZN(n8180) );
  NAND3X0 U11912 ( .IN1(n11646), .IN2(n11647), .IN3(n11648), .QN(n8178) );
  NAND2X0 U11913 ( .IN1(n7086), .IN2(g7357), .QN(n11648) );
  NAND2X0 U11914 ( .IN1(n7141), .IN2(g2009), .QN(n11647) );
  NAND2X0 U11915 ( .IN1(n7087), .IN2(g7229), .QN(n11646) );
  XOR2X1 U11916 ( .IN1(n4410), .IN2(n8184), .Q(n11644) );
  INVX0 U11917 ( .INP(n8185), .ZN(n8184) );
  NAND3X0 U11918 ( .IN1(n11649), .IN2(n11650), .IN3(n11651), .QN(n8185) );
  NAND2X0 U11919 ( .IN1(n7080), .IN2(g7357), .QN(n11651) );
  NAND2X0 U11920 ( .IN1(n7138), .IN2(g2009), .QN(n11650) );
  NAND2X0 U11921 ( .IN1(n7081), .IN2(g7229), .QN(n11649) );
  NAND3X0 U11922 ( .IN1(n11652), .IN2(n11653), .IN3(n11654), .QN(n11643) );
  XOR2X1 U11923 ( .IN1(n4416), .IN2(n8195), .Q(n11654) );
  NAND3X0 U11924 ( .IN1(n11655), .IN2(n11656), .IN3(n11657), .QN(n8195) );
  OR2X1 U11925 ( .IN1(n4357), .IN2(test_so72), .Q(n11657) );
  NAND2X0 U11926 ( .IN1(n7132), .IN2(g2009), .QN(n11656) );
  NAND2X0 U11927 ( .IN1(n7070), .IN2(g7229), .QN(n11655) );
  XOR2X1 U11928 ( .IN1(test_so70), .IN2(n8198), .Q(n11653) );
  INVX0 U11929 ( .INP(n8199), .ZN(n8198) );
  NAND3X0 U11930 ( .IN1(n11658), .IN2(n11659), .IN3(n11660), .QN(n8199) );
  NAND2X0 U11931 ( .IN1(n7071), .IN2(g7357), .QN(n11660) );
  NAND2X0 U11932 ( .IN1(n7133), .IN2(g2009), .QN(n11659) );
  NAND2X0 U11933 ( .IN1(n7072), .IN2(g7229), .QN(n11658) );
  XOR2X1 U11934 ( .IN1(g2052), .IN2(n8146), .Q(n11652) );
  INVX0 U11935 ( .INP(n8144), .ZN(n8146) );
  NAND3X0 U11936 ( .IN1(n11661), .IN2(n11662), .IN3(n11663), .QN(n8144) );
  NAND2X0 U11937 ( .IN1(n7077), .IN2(g7357), .QN(n11663) );
  NAND2X0 U11938 ( .IN1(n7136), .IN2(g2009), .QN(n11662) );
  NAND2X0 U11939 ( .IN1(n7078), .IN2(g7229), .QN(n11661) );
  NAND4X0 U11940 ( .IN1(n11664), .IN2(n11665), .IN3(n11666), .IN4(n11667), 
        .QN(n11642) );
  XOR2X1 U11941 ( .IN1(g2059), .IN2(n8160), .Q(n11667) );
  INVX0 U11942 ( .INP(n8159), .ZN(n8160) );
  NAND3X0 U11943 ( .IN1(n11668), .IN2(n11669), .IN3(n11670), .QN(n8159) );
  NAND2X0 U11944 ( .IN1(n7073), .IN2(g7357), .QN(n11670) );
  NAND2X0 U11945 ( .IN1(n7134), .IN2(g2009), .QN(n11669) );
  NAND2X0 U11946 ( .IN1(n7074), .IN2(g7229), .QN(n11668) );
  NOR2X0 U11947 ( .IN1(n11671), .IN2(n11672), .QN(n11666) );
  XOR2X1 U11948 ( .IN1(n4399), .IN2(n8156), .Q(n11672) );
  INVX0 U11949 ( .INP(n8155), .ZN(n8156) );
  NAND3X0 U11950 ( .IN1(n11673), .IN2(n11674), .IN3(n11675), .QN(n8155) );
  OR2X1 U11951 ( .IN1(n4357), .IN2(test_so71), .Q(n11675) );
  NAND2X0 U11952 ( .IN1(n7137), .IN2(g2009), .QN(n11674) );
  NAND2X0 U11953 ( .IN1(n7079), .IN2(g7229), .QN(n11673) );
  XOR2X1 U11954 ( .IN1(n4468), .IN2(n8152), .Q(n11671) );
  INVX0 U11955 ( .INP(n8150), .ZN(n8152) );
  NAND3X0 U11956 ( .IN1(n11676), .IN2(n11677), .IN3(n11678), .QN(n8150) );
  NAND2X0 U11957 ( .IN1(n7075), .IN2(g7357), .QN(n11678) );
  NAND2X0 U11958 ( .IN1(n7135), .IN2(g2009), .QN(n11677) );
  NAND2X0 U11959 ( .IN1(n7076), .IN2(g7229), .QN(n11676) );
  XOR2X1 U11960 ( .IN1(g2013), .IN2(n8172), .Q(n11665) );
  INVX0 U11961 ( .INP(n8175), .ZN(n8172) );
  NAND3X0 U11962 ( .IN1(n11679), .IN2(n11680), .IN3(n11681), .QN(n8175) );
  NAND2X0 U11963 ( .IN1(n7084), .IN2(g7357), .QN(n11681) );
  NAND2X0 U11964 ( .IN1(n7140), .IN2(g2009), .QN(n11680) );
  NAND2X0 U11965 ( .IN1(n7085), .IN2(g7229), .QN(n11679) );
  XOR2X1 U11966 ( .IN1(n4420), .IN2(n8166), .Q(n11664) );
  NAND3X0 U11967 ( .IN1(n11682), .IN2(n11683), .IN3(n11684), .QN(n8166) );
  NAND2X0 U11968 ( .IN1(n7082), .IN2(g7357), .QN(n11684) );
  NAND2X0 U11969 ( .IN1(n7139), .IN2(g2009), .QN(n11683) );
  NAND2X0 U11970 ( .IN1(n7083), .IN2(g7229), .QN(n11682) );
  NOR2X0 U11971 ( .IN1(n4357), .IN2(g2110), .QN(n11640) );
  NAND2X0 U11972 ( .IN1(n6843), .IN2(g7229), .QN(n11637) );
  INVX0 U11973 ( .INP(n8415), .ZN(n11636) );
  NAND3X0 U11974 ( .IN1(n11685), .IN2(n11686), .IN3(n11687), .QN(n8415) );
  NAND2X0 U11975 ( .IN1(n6834), .IN2(g7357), .QN(n11687) );
  NAND2X0 U11976 ( .IN1(n6897), .IN2(g2009), .QN(n11686) );
  NAND2X0 U11977 ( .IN1(n6842), .IN2(g7229), .QN(n11685) );
  OR2X1 U11978 ( .IN1(n11635), .IN2(n6770), .Q(n11633) );
  NAND2X0 U11979 ( .IN1(n11688), .IN2(n11689), .QN(g25267) );
  NAND2X0 U11980 ( .IN1(n11690), .IN2(n11631), .QN(n11689) );
  OR2X1 U11981 ( .IN1(n11690), .IN2(n6771), .Q(n11688) );
  NAND2X0 U11982 ( .IN1(n11691), .IN2(n11692), .QN(g25266) );
  NAND2X0 U11983 ( .IN1(n11693), .IN2(n11694), .QN(n11692) );
  OR2X1 U11984 ( .IN1(n11694), .IN2(n6778), .Q(n11691) );
  NAND2X0 U11985 ( .IN1(n11695), .IN2(n11696), .QN(g25265) );
  NAND2X0 U11986 ( .IN1(n11109), .IN2(n7825), .QN(n11696) );
  NAND2X0 U11987 ( .IN1(n11697), .IN2(n11474), .QN(n11695) );
  XOR2X1 U11988 ( .IN1(n6432), .IN2(n6431), .Q(n11697) );
  NAND2X0 U11989 ( .IN1(n11698), .IN2(n11699), .QN(g25263) );
  NAND2X0 U11990 ( .IN1(n11700), .IN2(n11631), .QN(n11699) );
  AND4X1 U11991 ( .IN1(n11701), .IN2(n11702), .IN3(n11703), .IN4(n11704), .Q(
        n11631) );
  NAND2X0 U11992 ( .IN1(n6837), .IN2(g7161), .QN(n11704) );
  NOR2X0 U11993 ( .IN1(n11705), .IN2(n11706), .QN(n11703) );
  NOR4X0 U11994 ( .IN1(n11707), .IN2(n11708), .IN3(n11709), .IN4(n11710), .QN(
        n11706) );
  XOR2X1 U11995 ( .IN1(n4421), .IN2(n8277), .Q(n11710) );
  INVX0 U11996 ( .INP(n8280), .ZN(n8277) );
  NAND3X0 U11997 ( .IN1(n11711), .IN2(n11712), .IN3(n11713), .QN(n8280) );
  NAND2X0 U11998 ( .IN1(n7101), .IN2(g7161), .QN(n11713) );
  NAND2X0 U11999 ( .IN1(n7149), .IN2(g1315), .QN(n11712) );
  NAND2X0 U12000 ( .IN1(n7102), .IN2(g6979), .QN(n11711) );
  XOR2X1 U12001 ( .IN1(n4476), .IN2(n8284), .Q(n11709) );
  INVX0 U12002 ( .INP(n8287), .ZN(n8284) );
  NAND3X0 U12003 ( .IN1(n11714), .IN2(n11715), .IN3(n11716), .QN(n8287) );
  NAND2X0 U12004 ( .IN1(n7103), .IN2(g7161), .QN(n11716) );
  NAND2X0 U12005 ( .IN1(n7150), .IN2(g1315), .QN(n11715) );
  NAND2X0 U12006 ( .IN1(n7104), .IN2(g6979), .QN(n11714) );
  NAND3X0 U12007 ( .IN1(n11717), .IN2(n11718), .IN3(n11719), .QN(n11708) );
  XOR2X1 U12008 ( .IN1(g1365), .IN2(n8271), .Q(n11719) );
  INVX0 U12009 ( .INP(n8270), .ZN(n8271) );
  NAND3X0 U12010 ( .IN1(n11720), .IN2(n11721), .IN3(n11722), .QN(n8270) );
  NAND2X0 U12011 ( .IN1(n7092), .IN2(g7161), .QN(n11722) );
  NAND2X0 U12012 ( .IN1(n7144), .IN2(g1315), .QN(n11721) );
  NAND2X0 U12013 ( .IN1(n7093), .IN2(g6979), .QN(n11720) );
  XOR2X1 U12014 ( .IN1(n4469), .IN2(n8261), .Q(n11718) );
  NAND3X0 U12015 ( .IN1(n11723), .IN2(n11724), .IN3(n11725), .QN(n8261) );
  NAND2X0 U12016 ( .IN1(n7094), .IN2(g7161), .QN(n11725) );
  NAND2X0 U12017 ( .IN1(n7145), .IN2(g1315), .QN(n11724) );
  NAND2X0 U12018 ( .IN1(n7095), .IN2(g6979), .QN(n11723) );
  XOR2X1 U12019 ( .IN1(g1346), .IN2(n8267), .Q(n11717) );
  INVX0 U12020 ( .INP(n8266), .ZN(n8267) );
  NAND3X0 U12021 ( .IN1(n11726), .IN2(n11727), .IN3(n11728), .QN(n8266) );
  NAND2X0 U12022 ( .IN1(n7097), .IN2(g7161), .QN(n11728) );
  NAND2X0 U12023 ( .IN1(n7147), .IN2(g1315), .QN(n11727) );
  NAND2X0 U12024 ( .IN1(n7098), .IN2(g6979), .QN(n11726) );
  NAND4X0 U12025 ( .IN1(n11729), .IN2(n11730), .IN3(n11731), .IN4(n11732), 
        .QN(n11707) );
  XOR2X1 U12026 ( .IN1(n4417), .IN2(n8306), .Q(n11732) );
  NAND3X0 U12027 ( .IN1(n11733), .IN2(n11734), .IN3(n11735), .QN(n8306) );
  NAND2X0 U12028 ( .IN1(n7088), .IN2(g7161), .QN(n11735) );
  NAND2X0 U12029 ( .IN1(n7142), .IN2(g1315), .QN(n11734) );
  NAND2X0 U12030 ( .IN1(n7089), .IN2(g6979), .QN(n11733) );
  NOR2X0 U12031 ( .IN1(n11736), .IN2(n11737), .QN(n11731) );
  XOR2X1 U12032 ( .IN1(n4395), .IN2(n8309), .Q(n11737) );
  INVX0 U12033 ( .INP(n8310), .ZN(n8309) );
  NAND3X0 U12034 ( .IN1(n11738), .IN2(n11739), .IN3(n11740), .QN(n8310) );
  NAND2X0 U12035 ( .IN1(n7090), .IN2(g7161), .QN(n11740) );
  NAND2X0 U12036 ( .IN1(n7143), .IN2(g1315), .QN(n11739) );
  NAND2X0 U12037 ( .IN1(n7091), .IN2(g6979), .QN(n11738) );
  XOR2X1 U12038 ( .IN1(n4411), .IN2(n8257), .Q(n11736) );
  INVX0 U12039 ( .INP(n8255), .ZN(n8257) );
  NAND3X0 U12040 ( .IN1(n11741), .IN2(n11742), .IN3(n11743), .QN(n8255) );
  OR2X1 U12041 ( .IN1(n4358), .IN2(test_so50), .Q(n11743) );
  NAND2X0 U12042 ( .IN1(n7146), .IN2(g1315), .QN(n11742) );
  NAND2X0 U12043 ( .IN1(n7096), .IN2(g6979), .QN(n11741) );
  XOR2X1 U12044 ( .IN1(g1332), .IN2(n8295), .Q(n11730) );
  INVX0 U12045 ( .INP(n8296), .ZN(n8295) );
  NAND3X0 U12046 ( .IN1(n11744), .IN2(n11745), .IN3(n11746), .QN(n8296) );
  NAND2X0 U12047 ( .IN1(n7099), .IN2(g7161), .QN(n11746) );
  NAND2X0 U12048 ( .IN1(n7148), .IN2(g1315), .QN(n11745) );
  NAND2X0 U12049 ( .IN1(n7100), .IN2(g6979), .QN(n11744) );
  XOR2X1 U12050 ( .IN1(n4402), .IN2(n8290), .Q(n11729) );
  NAND3X0 U12051 ( .IN1(n11747), .IN2(n11748), .IN3(n11749), .QN(n8290) );
  NAND2X0 U12052 ( .IN1(n7105), .IN2(g7161), .QN(n11749) );
  NAND2X0 U12053 ( .IN1(n7151), .IN2(g1315), .QN(n11748) );
  OR2X1 U12054 ( .IN1(n4308), .IN2(test_so49), .Q(n11747) );
  NOR2X0 U12055 ( .IN1(n4294), .IN2(test_so51), .QN(n11705) );
  NAND2X0 U12056 ( .IN1(n6845), .IN2(g6979), .QN(n11702) );
  INVX0 U12057 ( .INP(n8430), .ZN(n11701) );
  NAND3X0 U12058 ( .IN1(n11750), .IN2(n11751), .IN3(n11752), .QN(n8430) );
  NAND2X0 U12059 ( .IN1(n6836), .IN2(g7161), .QN(n11752) );
  NAND2X0 U12060 ( .IN1(n6899), .IN2(g1315), .QN(n11751) );
  NAND2X0 U12061 ( .IN1(n6844), .IN2(g6979), .QN(n11750) );
  OR2X1 U12062 ( .IN1(n11700), .IN2(n6772), .Q(n11698) );
  NAND2X0 U12063 ( .IN1(n11753), .IN2(n11754), .QN(g25262) );
  NAND2X0 U12064 ( .IN1(n11755), .IN2(n11693), .QN(n11754) );
  OR2X1 U12065 ( .IN1(n11755), .IN2(n6773), .Q(n11753) );
  NAND2X0 U12066 ( .IN1(n11756), .IN2(n11757), .QN(g25260) );
  NAND2X0 U12067 ( .IN1(n11758), .IN2(n11693), .QN(n11757) );
  AND4X1 U12068 ( .IN1(n11759), .IN2(n11760), .IN3(n11761), .IN4(n11762), .Q(
        n11693) );
  NAND2X0 U12069 ( .IN1(n6901), .IN2(g629), .QN(n11762) );
  NOR2X0 U12070 ( .IN1(n11763), .IN2(n11764), .QN(n11761) );
  NOR4X0 U12071 ( .IN1(n11765), .IN2(n11766), .IN3(n11767), .IN4(n11768), .QN(
        n11764) );
  XOR2X1 U12072 ( .IN1(n4422), .IN2(n7857), .Q(n11768) );
  INVX0 U12073 ( .INP(n7858), .ZN(n7857) );
  NAND3X0 U12074 ( .IN1(n11769), .IN2(n11770), .IN3(n11771), .QN(n7858) );
  NAND2X0 U12075 ( .IN1(n7118), .IN2(g6911), .QN(n11771) );
  NAND2X0 U12076 ( .IN1(n7159), .IN2(g629), .QN(n11770) );
  NAND2X0 U12077 ( .IN1(n7119), .IN2(g6677), .QN(n11769) );
  XOR2X1 U12078 ( .IN1(n4478), .IN2(n7861), .Q(n11767) );
  INVX0 U12079 ( .INP(n7862), .ZN(n7861) );
  NAND3X0 U12080 ( .IN1(n11772), .IN2(n11773), .IN3(n11774), .QN(n7862) );
  NAND2X0 U12081 ( .IN1(n7120), .IN2(g6911), .QN(n11774) );
  NAND2X0 U12082 ( .IN1(n7160), .IN2(g629), .QN(n11773) );
  NAND2X0 U12083 ( .IN1(n7121), .IN2(g6677), .QN(n11772) );
  NAND3X0 U12084 ( .IN1(n11775), .IN2(n11776), .IN3(n11777), .QN(n11766) );
  XOR2X1 U12085 ( .IN1(g640), .IN2(n7843), .Q(n11777) );
  INVX0 U12086 ( .INP(n7846), .ZN(n7843) );
  NAND3X0 U12087 ( .IN1(n11778), .IN2(n11779), .IN3(n11780), .QN(n7846) );
  NAND2X0 U12088 ( .IN1(n7122), .IN2(g6911), .QN(n11780) );
  NAND2X0 U12089 ( .IN1(n7161), .IN2(g629), .QN(n11779) );
  NAND2X0 U12090 ( .IN1(n7123), .IN2(g6677), .QN(n11778) );
  XOR2X1 U12091 ( .IN1(g660), .IN2(n7866), .Q(n11776) );
  INVX0 U12092 ( .INP(n7867), .ZN(n7866) );
  NAND3X0 U12093 ( .IN1(n11781), .IN2(n11782), .IN3(n11783), .QN(n7867) );
  NAND2X0 U12094 ( .IN1(n7115), .IN2(g6911), .QN(n11783) );
  NAND2X0 U12095 ( .IN1(n7157), .IN2(g629), .QN(n11782) );
  OR2X1 U12096 ( .IN1(n4309), .IN2(test_so29), .Q(n11781) );
  XOR2X1 U12097 ( .IN1(g679), .IN2(n7874), .Q(n11775) );
  INVX0 U12098 ( .INP(n7875), .ZN(n7874) );
  NAND3X0 U12099 ( .IN1(n11784), .IN2(n11785), .IN3(n11786), .QN(n7875) );
  NAND2X0 U12100 ( .IN1(n7109), .IN2(g6911), .QN(n11786) );
  NAND2X0 U12101 ( .IN1(n7154), .IN2(g629), .QN(n11785) );
  NAND2X0 U12102 ( .IN1(n7110), .IN2(g6677), .QN(n11784) );
  NAND4X0 U12103 ( .IN1(n11787), .IN2(n11788), .IN3(n11789), .IN4(n11790), 
        .QN(n11765) );
  XOR2X1 U12104 ( .IN1(n4418), .IN2(n7893), .Q(n11790) );
  NAND3X0 U12105 ( .IN1(n11791), .IN2(n11792), .IN3(n11793), .QN(n7893) );
  OR2X1 U12106 ( .IN1(n4359), .IN2(test_so30), .Q(n11793) );
  NAND2X0 U12107 ( .IN1(n7152), .IN2(g629), .QN(n11792) );
  NAND2X0 U12108 ( .IN1(n7106), .IN2(g6677), .QN(n11791) );
  NOR2X0 U12109 ( .IN1(n11794), .IN2(n11795), .QN(n11789) );
  XOR2X1 U12110 ( .IN1(n4396), .IN2(n7888), .Q(n11795) );
  INVX0 U12111 ( .INP(n7889), .ZN(n7888) );
  NAND3X0 U12112 ( .IN1(n11796), .IN2(n11797), .IN3(n11798), .QN(n7889) );
  NAND2X0 U12113 ( .IN1(n7107), .IN2(g6911), .QN(n11798) );
  NAND2X0 U12114 ( .IN1(n7153), .IN2(g629), .QN(n11797) );
  NAND2X0 U12115 ( .IN1(n7108), .IN2(g6677), .QN(n11796) );
  XOR2X1 U12116 ( .IN1(n7270), .IN2(n7870), .Q(n11794) );
  INVX0 U12117 ( .INP(n7871), .ZN(n7870) );
  NAND3X0 U12118 ( .IN1(n11799), .IN2(n11800), .IN3(n11801), .QN(n7871) );
  NAND2X0 U12119 ( .IN1(n7111), .IN2(g6911), .QN(n11801) );
  NAND2X0 U12120 ( .IN1(n7155), .IN2(g629), .QN(n11800) );
  NAND2X0 U12121 ( .IN1(n7112), .IN2(g6677), .QN(n11799) );
  XOR2X1 U12122 ( .IN1(g672), .IN2(n7878), .Q(n11788) );
  INVX0 U12123 ( .INP(n7879), .ZN(n7878) );
  NAND3X0 U12124 ( .IN1(n11802), .IN2(n11803), .IN3(n11804), .QN(n7879) );
  NAND2X0 U12125 ( .IN1(n7113), .IN2(g6911), .QN(n11804) );
  NAND2X0 U12126 ( .IN1(n7156), .IN2(g629), .QN(n11803) );
  NAND2X0 U12127 ( .IN1(n7114), .IN2(g6677), .QN(n11802) );
  XOR2X1 U12128 ( .IN1(g646), .IN2(n7850), .Q(n11787) );
  INVX0 U12129 ( .INP(n7853), .ZN(n7850) );
  NAND3X0 U12130 ( .IN1(n11805), .IN2(n11806), .IN3(n11807), .QN(n7853) );
  NAND2X0 U12131 ( .IN1(n7116), .IN2(g6911), .QN(n11807) );
  NAND2X0 U12132 ( .IN1(n7158), .IN2(g629), .QN(n11806) );
  NAND2X0 U12133 ( .IN1(n7117), .IN2(g6677), .QN(n11805) );
  NOR2X0 U12134 ( .IN1(n4359), .IN2(g730), .QN(n11763) );
  NAND2X0 U12135 ( .IN1(n6847), .IN2(g6677), .QN(n11760) );
  INVX0 U12136 ( .INP(n8386), .ZN(n11759) );
  NAND3X0 U12137 ( .IN1(n11808), .IN2(n11809), .IN3(n11810), .QN(n8386) );
  NAND2X0 U12138 ( .IN1(n6838), .IN2(g6911), .QN(n11810) );
  NAND2X0 U12139 ( .IN1(n6900), .IN2(g629), .QN(n11809) );
  NAND2X0 U12140 ( .IN1(n6846), .IN2(g6677), .QN(n11808) );
  OR2X1 U12141 ( .IN1(n11758), .IN2(n6774), .Q(n11756) );
  NAND2X0 U12142 ( .IN1(n11811), .IN2(n11812), .QN(g25259) );
  OR2X1 U12143 ( .IN1(n11813), .IN2(n6848), .Q(n11812) );
  NAND2X0 U12144 ( .IN1(n11813), .IN2(n11022), .QN(n11811) );
  NAND2X0 U12145 ( .IN1(n11814), .IN2(n11815), .QN(g25257) );
  OR2X1 U12146 ( .IN1(n11816), .IN2(n6849), .Q(n11815) );
  NAND2X0 U12147 ( .IN1(n11816), .IN2(n11022), .QN(n11814) );
  NAND2X0 U12148 ( .IN1(n11817), .IN2(n11818), .QN(g25256) );
  NAND2X0 U12149 ( .IN1(n11813), .IN2(n4377), .QN(n11818) );
  OR2X1 U12150 ( .IN1(n11813), .IN2(n6851), .Q(n11817) );
  NAND2X0 U12151 ( .IN1(n11819), .IN2(n11820), .QN(g25255) );
  NAND2X0 U12152 ( .IN1(n11821), .IN2(n11052), .QN(n11820) );
  OR2X1 U12153 ( .IN1(n11821), .IN2(n6860), .Q(n11819) );
  NAND2X0 U12154 ( .IN1(n11822), .IN2(n11823), .QN(g25253) );
  OR2X1 U12155 ( .IN1(n11824), .IN2(n6850), .Q(n11823) );
  NAND2X0 U12156 ( .IN1(n11824), .IN2(n11022), .QN(n11822) );
  NAND4X0 U12157 ( .IN1(g2200), .IN2(g2175), .IN3(n11825), .IN4(n11826), .QN(
        n11022) );
  NOR4X0 U12158 ( .IN1(n4563), .IN2(n4555), .IN3(n4389), .IN4(n4377), .QN(
        n11826) );
  NOR2X0 U12159 ( .IN1(n4373), .IN2(n4325), .QN(n11825) );
  NAND2X0 U12160 ( .IN1(n11827), .IN2(n11828), .QN(g25252) );
  NAND2X0 U12161 ( .IN1(n11816), .IN2(n4377), .QN(n11828) );
  OR2X1 U12162 ( .IN1(n11816), .IN2(n6852), .Q(n11827) );
  NAND2X0 U12163 ( .IN1(n11829), .IN2(n11830), .QN(g25251) );
  NAND2X0 U12164 ( .IN1(n11813), .IN2(n4373), .QN(n11830) );
  OR2X1 U12165 ( .IN1(n11813), .IN2(n6854), .Q(n11829) );
  NAND2X0 U12166 ( .IN1(n11831), .IN2(n11832), .QN(g25250) );
  OR2X1 U12167 ( .IN1(n11833), .IN2(n6861), .Q(n11832) );
  NAND2X0 U12168 ( .IN1(n11833), .IN2(n11052), .QN(n11831) );
  NAND2X0 U12169 ( .IN1(n11834), .IN2(n11835), .QN(g25249) );
  NAND2X0 U12170 ( .IN1(n11821), .IN2(n4378), .QN(n11835) );
  OR2X1 U12171 ( .IN1(n11821), .IN2(n6863), .Q(n11834) );
  NAND2X0 U12172 ( .IN1(n11836), .IN2(n11837), .QN(g25248) );
  OR2X1 U12173 ( .IN1(n11838), .IN2(n6871), .Q(n11837) );
  NAND2X0 U12174 ( .IN1(n11838), .IN2(n11079), .QN(n11836) );
  NAND2X0 U12175 ( .IN1(n11839), .IN2(n11840), .QN(g25247) );
  NAND2X0 U12176 ( .IN1(n11824), .IN2(n4377), .QN(n11840) );
  OR2X1 U12177 ( .IN1(n11824), .IN2(n6853), .Q(n11839) );
  NAND2X0 U12178 ( .IN1(n11841), .IN2(n11842), .QN(g25246) );
  NAND2X0 U12179 ( .IN1(n11816), .IN2(n4373), .QN(n11842) );
  OR2X1 U12180 ( .IN1(n11816), .IN2(n6855), .Q(n11841) );
  NAND2X0 U12181 ( .IN1(n11843), .IN2(n11844), .QN(g25245) );
  NAND2X0 U12182 ( .IN1(n11845), .IN2(n11813), .QN(n11844) );
  OR2X1 U12183 ( .IN1(n11813), .IN2(n6857), .Q(n11843) );
  AND2X1 U12184 ( .IN1(g13110), .IN2(g2241), .Q(n11813) );
  NAND2X0 U12185 ( .IN1(n11846), .IN2(n11847), .QN(g25244) );
  OR2X1 U12186 ( .IN1(n11848), .IN2(n6862), .Q(n11847) );
  NAND2X0 U12187 ( .IN1(n11848), .IN2(n11052), .QN(n11846) );
  NAND4X0 U12188 ( .IN1(g1506), .IN2(g1481), .IN3(n11849), .IN4(n11850), .QN(
        n11052) );
  NOR4X0 U12189 ( .IN1(n4565), .IN2(n4557), .IN3(n4390), .IN4(n4378), .QN(
        n11850) );
  NOR2X0 U12190 ( .IN1(n4374), .IN2(n4326), .QN(n11849) );
  NAND2X0 U12191 ( .IN1(n11851), .IN2(n11852), .QN(g25243) );
  NAND2X0 U12192 ( .IN1(n11833), .IN2(n4378), .QN(n11852) );
  OR2X1 U12193 ( .IN1(n11833), .IN2(n6864), .Q(n11851) );
  NAND2X0 U12194 ( .IN1(n11853), .IN2(n11854), .QN(g25242) );
  NAND2X0 U12195 ( .IN1(test_so54), .IN2(n11855), .QN(n11854) );
  NAND2X0 U12196 ( .IN1(n11821), .IN2(n4374), .QN(n11853) );
  NAND2X0 U12197 ( .IN1(n11856), .IN2(n11857), .QN(g25241) );
  NAND2X0 U12198 ( .IN1(n11858), .IN2(n11079), .QN(n11857) );
  OR2X1 U12199 ( .IN1(n11858), .IN2(n6872), .Q(n11856) );
  NAND2X0 U12200 ( .IN1(n11859), .IN2(n11860), .QN(g25240) );
  NAND2X0 U12201 ( .IN1(n4379), .IN2(n11838), .QN(n11860) );
  OR2X1 U12202 ( .IN1(n11838), .IN2(n6874), .Q(n11859) );
  NAND2X0 U12203 ( .IN1(n11861), .IN2(n11862), .QN(g25239) );
  OR2X1 U12204 ( .IN1(n11863), .IN2(n6882), .Q(n11862) );
  NAND2X0 U12205 ( .IN1(n11863), .IN2(n11101), .QN(n11861) );
  NAND2X0 U12206 ( .IN1(n11864), .IN2(n11865), .QN(g25237) );
  NAND2X0 U12207 ( .IN1(n11824), .IN2(n4373), .QN(n11865) );
  OR2X1 U12208 ( .IN1(n11824), .IN2(n6856), .Q(n11864) );
  NAND2X0 U12209 ( .IN1(n11866), .IN2(n11867), .QN(g25236) );
  NAND2X0 U12210 ( .IN1(n11845), .IN2(n11816), .QN(n11867) );
  OR2X1 U12211 ( .IN1(n11816), .IN2(n6858), .Q(n11866) );
  AND2X1 U12212 ( .IN1(g13110), .IN2(test_so73), .Q(n11816) );
  NAND2X0 U12213 ( .IN1(n11868), .IN2(n11869), .QN(g25235) );
  NAND2X0 U12214 ( .IN1(n11848), .IN2(n4378), .QN(n11869) );
  OR2X1 U12215 ( .IN1(n11848), .IN2(n6865), .Q(n11868) );
  NAND2X0 U12216 ( .IN1(n11870), .IN2(n11871), .QN(g25234) );
  NAND2X0 U12217 ( .IN1(n11833), .IN2(n4374), .QN(n11871) );
  OR2X1 U12218 ( .IN1(n11833), .IN2(n6866), .Q(n11870) );
  NAND2X0 U12219 ( .IN1(n11872), .IN2(n11873), .QN(g25233) );
  NAND2X0 U12220 ( .IN1(n11874), .IN2(n11821), .QN(n11873) );
  OR2X1 U12221 ( .IN1(n11821), .IN2(n6868), .Q(n11872) );
  INVX0 U12222 ( .INP(n11855), .ZN(n11821) );
  NAND2X0 U12223 ( .IN1(g13110), .IN2(g1547), .QN(n11855) );
  NAND2X0 U12224 ( .IN1(n11875), .IN2(n11876), .QN(g25232) );
  OR2X1 U12225 ( .IN1(n11877), .IN2(n6873), .Q(n11876) );
  NAND2X0 U12226 ( .IN1(n11877), .IN2(n11079), .QN(n11875) );
  NAND4X0 U12227 ( .IN1(g813), .IN2(g793), .IN3(n11878), .IN4(n11879), .QN(
        n11079) );
  NOR4X0 U12228 ( .IN1(n4567), .IN2(n4559), .IN3(n4391), .IN4(n4379), .QN(
        n11879) );
  NOR2X0 U12229 ( .IN1(n4375), .IN2(n4327), .QN(n11878) );
  NAND2X0 U12230 ( .IN1(n11880), .IN2(n11881), .QN(g25231) );
  NAND2X0 U12231 ( .IN1(n4379), .IN2(n11858), .QN(n11881) );
  OR2X1 U12232 ( .IN1(n11858), .IN2(n6875), .Q(n11880) );
  NAND2X0 U12233 ( .IN1(n11882), .IN2(n11883), .QN(g25230) );
  NAND2X0 U12234 ( .IN1(n11838), .IN2(n4375), .QN(n11883) );
  OR2X1 U12235 ( .IN1(n11838), .IN2(n6877), .Q(n11882) );
  NAND2X0 U12236 ( .IN1(n11884), .IN2(n11885), .QN(g25229) );
  OR2X1 U12237 ( .IN1(n11886), .IN2(n6883), .Q(n11885) );
  NAND2X0 U12238 ( .IN1(n11886), .IN2(n11101), .QN(n11884) );
  NAND2X0 U12239 ( .IN1(n11887), .IN2(n11888), .QN(g25228) );
  NAND2X0 U12240 ( .IN1(n4380), .IN2(n11863), .QN(n11888) );
  OR2X1 U12241 ( .IN1(n11863), .IN2(n6885), .Q(n11887) );
  NAND2X0 U12242 ( .IN1(n11889), .IN2(n11890), .QN(g25227) );
  OR2X1 U12243 ( .IN1(n11824), .IN2(n6859), .Q(n11890) );
  NAND2X0 U12244 ( .IN1(n11845), .IN2(n11824), .QN(n11889) );
  AND2X1 U12245 ( .IN1(g13110), .IN2(g6837), .Q(n11824) );
  NOR4X0 U12246 ( .IN1(g2195), .IN2(g2190), .IN3(n4287), .IN4(n4325), .QN(
        n11845) );
  NAND2X0 U12247 ( .IN1(n11891), .IN2(n11892), .QN(g25225) );
  NAND2X0 U12248 ( .IN1(n11848), .IN2(n4374), .QN(n11892) );
  OR2X1 U12249 ( .IN1(n11848), .IN2(n6867), .Q(n11891) );
  NAND2X0 U12250 ( .IN1(n11893), .IN2(n11894), .QN(g25224) );
  NAND2X0 U12251 ( .IN1(n11874), .IN2(n11833), .QN(n11894) );
  OR2X1 U12252 ( .IN1(n11833), .IN2(n6869), .Q(n11893) );
  AND2X1 U12253 ( .IN1(g13110), .IN2(g6782), .Q(n11833) );
  NAND2X0 U12254 ( .IN1(n11895), .IN2(n11896), .QN(g25223) );
  NAND2X0 U12255 ( .IN1(n11877), .IN2(n4379), .QN(n11896) );
  OR2X1 U12256 ( .IN1(n11877), .IN2(n6876), .Q(n11895) );
  NAND2X0 U12257 ( .IN1(n11897), .IN2(n11898), .QN(g25222) );
  NAND2X0 U12258 ( .IN1(n11858), .IN2(n4375), .QN(n11898) );
  OR2X1 U12259 ( .IN1(n11858), .IN2(n6878), .Q(n11897) );
  NAND2X0 U12260 ( .IN1(n11899), .IN2(n11900), .QN(g25221) );
  NAND2X0 U12261 ( .IN1(n11901), .IN2(n11838), .QN(n11900) );
  OR2X1 U12262 ( .IN1(n11838), .IN2(n6880), .Q(n11899) );
  AND2X1 U12263 ( .IN1(g13110), .IN2(test_so31), .Q(n11838) );
  NAND2X0 U12264 ( .IN1(n11902), .IN2(n11903), .QN(g25220) );
  OR2X1 U12265 ( .IN1(n11904), .IN2(n6884), .Q(n11903) );
  NAND2X0 U12266 ( .IN1(n11904), .IN2(n11101), .QN(n11902) );
  NAND4X0 U12267 ( .IN1(g125), .IN2(g105), .IN3(n11905), .IN4(n11906), .QN(
        n11101) );
  NOR4X0 U12268 ( .IN1(n4569), .IN2(n4561), .IN3(n4392), .IN4(n4380), .QN(
        n11906) );
  NOR2X0 U12269 ( .IN1(n4376), .IN2(n4328), .QN(n11905) );
  NAND2X0 U12270 ( .IN1(n11907), .IN2(n11908), .QN(g25219) );
  NAND2X0 U12271 ( .IN1(n4380), .IN2(n11886), .QN(n11908) );
  OR2X1 U12272 ( .IN1(n11886), .IN2(n6886), .Q(n11907) );
  NAND2X0 U12273 ( .IN1(n11909), .IN2(n11910), .QN(g25218) );
  NAND2X0 U12274 ( .IN1(n11863), .IN2(n4376), .QN(n11910) );
  OR2X1 U12275 ( .IN1(n11863), .IN2(n6888), .Q(n11909) );
  NAND2X0 U12276 ( .IN1(n11911), .IN2(n11912), .QN(g25217) );
  OR2X1 U12277 ( .IN1(n11848), .IN2(n6870), .Q(n11912) );
  NAND2X0 U12278 ( .IN1(n11874), .IN2(n11848), .QN(n11911) );
  AND2X1 U12279 ( .IN1(g13110), .IN2(g6573), .Q(n11848) );
  NOR4X0 U12280 ( .IN1(g1501), .IN2(g1496), .IN3(n4288), .IN4(n4326), .QN(
        n11874) );
  NAND2X0 U12281 ( .IN1(n11913), .IN2(n11914), .QN(g25215) );
  NAND2X0 U12282 ( .IN1(n11877), .IN2(n4375), .QN(n11914) );
  OR2X1 U12283 ( .IN1(n11877), .IN2(n6879), .Q(n11913) );
  NAND2X0 U12284 ( .IN1(n11915), .IN2(n11916), .QN(g25214) );
  NAND2X0 U12285 ( .IN1(test_so33), .IN2(n11917), .QN(n11916) );
  NAND2X0 U12286 ( .IN1(n11901), .IN2(n11858), .QN(n11915) );
  INVX0 U12287 ( .INP(n11917), .ZN(n11858) );
  NAND2X0 U12288 ( .IN1(g13110), .IN2(g6518), .QN(n11917) );
  NAND2X0 U12289 ( .IN1(n11918), .IN2(n11919), .QN(g25213) );
  NAND2X0 U12290 ( .IN1(n11904), .IN2(n4380), .QN(n11919) );
  OR2X1 U12291 ( .IN1(n11904), .IN2(n6887), .Q(n11918) );
  NAND2X0 U12292 ( .IN1(n11920), .IN2(n11921), .QN(g25212) );
  NAND2X0 U12293 ( .IN1(n11886), .IN2(n4376), .QN(n11921) );
  OR2X1 U12294 ( .IN1(n11886), .IN2(n6889), .Q(n11920) );
  NAND2X0 U12295 ( .IN1(n11922), .IN2(n11923), .QN(g25211) );
  NAND2X0 U12296 ( .IN1(n11924), .IN2(n11863), .QN(n11923) );
  OR2X1 U12297 ( .IN1(n11863), .IN2(n6891), .Q(n11922) );
  AND2X1 U12298 ( .IN1(g13110), .IN2(g165), .Q(n11863) );
  NAND2X0 U12299 ( .IN1(n11925), .IN2(n11926), .QN(g25209) );
  OR2X1 U12300 ( .IN1(n11877), .IN2(n6881), .Q(n11926) );
  NAND2X0 U12301 ( .IN1(n11901), .IN2(n11877), .QN(n11925) );
  AND2X1 U12302 ( .IN1(g13110), .IN2(g6368), .Q(n11877) );
  NOR4X0 U12303 ( .IN1(g809), .IN2(g805), .IN3(n4289), .IN4(n4327), .QN(n11901) );
  NAND2X0 U12304 ( .IN1(n11927), .IN2(n11928), .QN(g25207) );
  NAND2X0 U12305 ( .IN1(n11904), .IN2(n4376), .QN(n11928) );
  OR2X1 U12306 ( .IN1(n11904), .IN2(n6890), .Q(n11927) );
  NAND2X0 U12307 ( .IN1(n11929), .IN2(n11930), .QN(g25206) );
  NAND2X0 U12308 ( .IN1(n11924), .IN2(n11886), .QN(n11930) );
  OR2X1 U12309 ( .IN1(n11886), .IN2(n6892), .Q(n11929) );
  AND2X1 U12310 ( .IN1(g13110), .IN2(g6313), .Q(n11886) );
  NAND2X0 U12311 ( .IN1(n11931), .IN2(n11932), .QN(g25204) );
  OR2X1 U12312 ( .IN1(n11904), .IN2(n6893), .Q(n11932) );
  NAND2X0 U12313 ( .IN1(n11924), .IN2(n11904), .QN(n11931) );
  AND2X1 U12314 ( .IN1(g13110), .IN2(g6231), .Q(n11904) );
  NOR4X0 U12315 ( .IN1(g121), .IN2(g117), .IN3(n4290), .IN4(n4328), .QN(n11924) );
  NOR2X0 U12316 ( .IN1(n11933), .IN2(n11934), .QN(g25202) );
  XOR2X1 U12317 ( .IN1(n6706), .IN2(n11935), .Q(n11934) );
  NOR3X0 U12318 ( .IN1(n7777), .IN2(n4057), .IN3(n11104), .QN(g25201) );
  NOR2X0 U12319 ( .IN1(n4058), .IN2(n4305), .QN(n11104) );
  NAND2X0 U12320 ( .IN1(n11936), .IN2(g2892), .QN(n4058) );
  NOR2X0 U12321 ( .IN1(n11937), .IN2(n11938), .QN(g25199) );
  XNOR2X1 U12322 ( .IN1(n6995), .IN2(n11939), .Q(n11938) );
  NOR2X0 U12323 ( .IN1(n10335), .IN2(n11940), .QN(g25197) );
  XOR2X1 U12324 ( .IN1(n4397), .IN2(n11113), .Q(n11940) );
  NOR2X0 U12325 ( .IN1(n10339), .IN2(n11941), .QN(g25194) );
  XOR2X1 U12326 ( .IN1(n4399), .IN2(n11132), .Q(n11941) );
  AND3X1 U12327 ( .IN1(n11942), .IN2(n3742), .IN3(n11474), .Q(g25191) );
  NAND2X0 U12328 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  OR2X1 U12329 ( .IN1(g3013), .IN2(n4065), .Q(n11942) );
  NOR2X0 U12330 ( .IN1(n10343), .IN2(n11943), .QN(g25189) );
  XOR2X1 U12331 ( .IN1(n4401), .IN2(n11203), .Q(n11943) );
  NOR2X0 U12332 ( .IN1(n9912), .IN2(n11944), .QN(g25185) );
  XOR2X1 U12333 ( .IN1(n4403), .IN2(n11274), .Q(n11944) );
  NOR2X0 U12334 ( .IN1(n9318), .IN2(n11945), .QN(g25067) );
  XNOR2X1 U12335 ( .IN1(n6982), .IN2(n3888), .Q(n11945) );
  NAND2X0 U12336 ( .IN1(g2241), .IN2(n7678), .QN(n3888) );
  INVX0 U12337 ( .INP(n9736), .ZN(n9318) );
  NAND2X0 U12338 ( .IN1(n11946), .IN2(n10780), .QN(n9736) );
  NOR2X0 U12339 ( .IN1(n9320), .IN2(n11947), .QN(g25056) );
  XNOR2X1 U12340 ( .IN1(n6986), .IN2(n3891), .Q(n11947) );
  NAND2X0 U12341 ( .IN1(g1547), .IN2(n7678), .QN(n3891) );
  INVX0 U12342 ( .INP(n9739), .ZN(n9320) );
  NAND2X0 U12343 ( .IN1(n11948), .IN2(n10780), .QN(n9739) );
  NOR2X0 U12344 ( .IN1(n9322), .IN2(n11949), .QN(g25042) );
  XNOR2X1 U12345 ( .IN1(n6990), .IN2(n3894), .Q(n11949) );
  NAND2X0 U12346 ( .IN1(test_so31), .IN2(n7678), .QN(n3894) );
  AND2X1 U12347 ( .IN1(n11950), .IN2(n10780), .Q(n9322) );
  NOR2X0 U12348 ( .IN1(n9324), .IN2(n11951), .QN(g25027) );
  XNOR2X1 U12349 ( .IN1(n6994), .IN2(n3897), .Q(n11951) );
  NAND2X0 U12350 ( .IN1(g165), .IN2(n7678), .QN(n3897) );
  INVX0 U12351 ( .INP(n9743), .ZN(n9324) );
  NAND2X0 U12352 ( .IN1(n11952), .IN2(n10780), .QN(n9743) );
  NAND2X0 U12353 ( .IN1(n3700), .IN2(n11953), .QN(g24734) );
  NAND2X0 U12354 ( .IN1(n10489), .IN2(DFF_146_n1), .QN(n11953) );
  AND2X1 U12355 ( .IN1(n3940), .IN2(n3705), .Q(n10489) );
  NAND2X0 U12356 ( .IN1(n11954), .IN2(n11955), .QN(g24557) );
  NAND2X0 U12357 ( .IN1(n11956), .IN2(n8318), .QN(n11955) );
  NAND2X0 U12358 ( .IN1(n4299), .IN2(g2676), .QN(n11954) );
  NAND2X0 U12359 ( .IN1(n11957), .IN2(n11958), .QN(g24548) );
  NAND2X0 U12360 ( .IN1(n4370), .IN2(g2673), .QN(n11958) );
  NAND3X0 U12361 ( .IN1(n9947), .IN2(n8318), .IN3(g7390), .QN(n11957) );
  NAND2X0 U12362 ( .IN1(n11959), .IN2(n11960), .QN(g24547) );
  NAND2X0 U12363 ( .IN1(n11956), .IN2(n10003), .QN(n11960) );
  INVX0 U12364 ( .INP(n11961), .ZN(n11956) );
  NAND2X0 U12365 ( .IN1(n4299), .IN2(g2667), .QN(n11959) );
  NAND2X0 U12366 ( .IN1(n11962), .IN2(n11963), .QN(g24545) );
  NAND2X0 U12367 ( .IN1(n11964), .IN2(n10047), .QN(n11963) );
  NAND2X0 U12368 ( .IN1(n4366), .IN2(g1982), .QN(n11962) );
  NAND2X0 U12369 ( .IN1(n11965), .IN2(n11966), .QN(g24538) );
  NAND3X0 U12370 ( .IN1(n9947), .IN2(n8318), .IN3(g7302), .QN(n11966) );
  NAND4X0 U12371 ( .IN1(n11967), .IN2(n11968), .IN3(n11969), .IN4(n11970), 
        .QN(n8318) );
  NAND3X0 U12372 ( .IN1(n7650), .IN2(g185), .IN3(test_so88), .QN(n11970) );
  NAND3X0 U12373 ( .IN1(n11971), .IN2(n11972), .IN3(n11973), .QN(n7650) );
  NAND2X0 U12374 ( .IN1(g7390), .IN2(g2641), .QN(n11973) );
  NAND2X0 U12375 ( .IN1(g2624), .IN2(g2564), .QN(n11972) );
  NAND2X0 U12376 ( .IN1(n9246), .IN2(g2639), .QN(n11971) );
  NAND2X0 U12377 ( .IN1(g2624), .IN2(g2676), .QN(n11969) );
  NAND2X0 U12378 ( .IN1(n9246), .IN2(g2670), .QN(n11968) );
  NAND2X0 U12379 ( .IN1(g7390), .IN2(g2673), .QN(n11967) );
  NAND2X0 U12380 ( .IN1(n4314), .IN2(g2670), .QN(n11965) );
  NAND2X0 U12381 ( .IN1(n11974), .IN2(n11975), .QN(g24537) );
  NAND2X0 U12382 ( .IN1(n4370), .IN2(g2664), .QN(n11975) );
  NAND3X0 U12383 ( .IN1(n9947), .IN2(n10003), .IN3(g7390), .QN(n11974) );
  NAND2X0 U12384 ( .IN1(n11976), .IN2(n11977), .QN(g24535) );
  NAND2X0 U12385 ( .IN1(n4315), .IN2(g1979), .QN(n11977) );
  NAND3X0 U12386 ( .IN1(n10047), .IN2(n9947), .IN3(g7194), .QN(n11976) );
  NAND2X0 U12387 ( .IN1(n11978), .IN2(n11979), .QN(g24534) );
  NAND2X0 U12388 ( .IN1(n11964), .IN2(n10139), .QN(n11979) );
  INVX0 U12389 ( .INP(n11980), .ZN(n11964) );
  NAND2X0 U12390 ( .IN1(n4366), .IN2(g1973), .QN(n11978) );
  NAND2X0 U12391 ( .IN1(n11981), .IN2(n11982), .QN(g24532) );
  NAND2X0 U12392 ( .IN1(n11983), .IN2(n10150), .QN(n11982) );
  NAND2X0 U12393 ( .IN1(n4300), .IN2(g1288), .QN(n11981) );
  NAND2X0 U12394 ( .IN1(n11984), .IN2(n11985), .QN(g24527) );
  NAND2X0 U12395 ( .IN1(n4314), .IN2(g2661), .QN(n11985) );
  NAND3X0 U12396 ( .IN1(n9947), .IN2(n10003), .IN3(n9246), .QN(n11984) );
  NAND4X0 U12397 ( .IN1(n11986), .IN2(n11987), .IN3(n11988), .IN4(n11989), 
        .QN(n10003) );
  NAND3X0 U12398 ( .IN1(g185), .IN2(g2598), .IN3(n7649), .QN(n11989) );
  NAND3X0 U12399 ( .IN1(n11990), .IN2(n11991), .IN3(n11992), .QN(n7649) );
  NAND2X0 U12400 ( .IN1(g7390), .IN2(g2645), .QN(n11992) );
  NAND2X0 U12401 ( .IN1(g7302), .IN2(g2643), .QN(n11991) );
  NAND2X0 U12402 ( .IN1(g2624), .IN2(g2647), .QN(n11990) );
  NAND2X0 U12403 ( .IN1(g7302), .IN2(g2661), .QN(n11988) );
  NAND2X0 U12404 ( .IN1(g2624), .IN2(g2667), .QN(n11987) );
  NAND2X0 U12405 ( .IN1(g7390), .IN2(g2664), .QN(n11986) );
  NAND2X0 U12406 ( .IN1(n11993), .IN2(n11994), .QN(g24525) );
  NAND3X0 U12407 ( .IN1(n10047), .IN2(n9947), .IN3(g7052), .QN(n11994) );
  NAND4X0 U12408 ( .IN1(n11995), .IN2(n11996), .IN3(n11997), .IN4(n11998), 
        .QN(n10047) );
  NAND3X0 U12409 ( .IN1(g185), .IN2(g1922), .IN3(n7653), .QN(n11998) );
  NAND3X0 U12410 ( .IN1(n11999), .IN2(n12000), .IN3(n12001), .QN(n7653) );
  NAND2X0 U12411 ( .IN1(g1930), .IN2(g1870), .QN(n12001) );
  NAND2X0 U12412 ( .IN1(n9268), .IN2(g1945), .QN(n12000) );
  NAND2X0 U12413 ( .IN1(g7194), .IN2(g1947), .QN(n11999) );
  NAND2X0 U12414 ( .IN1(n9268), .IN2(g1976), .QN(n11997) );
  NAND2X0 U12415 ( .IN1(g7194), .IN2(g1979), .QN(n11996) );
  NAND2X0 U12416 ( .IN1(g1930), .IN2(g1982), .QN(n11995) );
  NAND2X0 U12417 ( .IN1(n4296), .IN2(g1976), .QN(n11993) );
  NAND2X0 U12418 ( .IN1(n12002), .IN2(n12003), .QN(g24524) );
  NAND2X0 U12419 ( .IN1(n4315), .IN2(g1970), .QN(n12003) );
  NAND3X0 U12420 ( .IN1(n10139), .IN2(n9947), .IN3(g7194), .QN(n12002) );
  NAND2X0 U12421 ( .IN1(n12004), .IN2(n12005), .QN(g24522) );
  NAND2X0 U12422 ( .IN1(n4316), .IN2(g1285), .QN(n12005) );
  NAND3X0 U12423 ( .IN1(n10150), .IN2(n9947), .IN3(g6944), .QN(n12004) );
  NAND2X0 U12424 ( .IN1(n12006), .IN2(n12007), .QN(g24521) );
  NAND2X0 U12425 ( .IN1(n11983), .IN2(n10239), .QN(n12007) );
  INVX0 U12426 ( .INP(n12008), .ZN(n11983) );
  NAND2X0 U12427 ( .IN1(n4300), .IN2(g1279), .QN(n12006) );
  NAND2X0 U12428 ( .IN1(n12009), .IN2(n12010), .QN(g24519) );
  NAND2X0 U12429 ( .IN1(n12011), .IN2(n10250), .QN(n12010) );
  NAND2X0 U12430 ( .IN1(n4313), .IN2(g602), .QN(n12009) );
  NAND2X0 U12431 ( .IN1(n12012), .IN2(n12013), .QN(g24513) );
  NAND2X0 U12432 ( .IN1(n4296), .IN2(g1967), .QN(n12013) );
  NAND3X0 U12433 ( .IN1(n10139), .IN2(n9947), .IN3(n9268), .QN(n12012) );
  NAND4X0 U12434 ( .IN1(n12014), .IN2(n12015), .IN3(n12016), .IN4(n12017), 
        .QN(n10139) );
  NAND3X0 U12435 ( .IN1(g185), .IN2(g1904), .IN3(n7652), .QN(n12017) );
  NAND3X0 U12436 ( .IN1(n12018), .IN2(n12019), .IN3(n12020), .QN(n7652) );
  NAND2X0 U12437 ( .IN1(g1930), .IN2(g1953), .QN(n12020) );
  NAND2X0 U12438 ( .IN1(g7052), .IN2(g1949), .QN(n12019) );
  NAND2X0 U12439 ( .IN1(g7194), .IN2(g1951), .QN(n12018) );
  NAND2X0 U12440 ( .IN1(g7052), .IN2(g1967), .QN(n12016) );
  NAND2X0 U12441 ( .IN1(g7194), .IN2(g1970), .QN(n12015) );
  NAND2X0 U12442 ( .IN1(g1930), .IN2(g1973), .QN(n12014) );
  NAND2X0 U12443 ( .IN1(n12021), .IN2(n12022), .QN(g24511) );
  NAND3X0 U12444 ( .IN1(n10150), .IN2(n9947), .IN3(g6750), .QN(n12022) );
  NAND4X0 U12445 ( .IN1(n12023), .IN2(n12024), .IN3(n12025), .IN4(n12026), 
        .QN(n10150) );
  NAND3X0 U12446 ( .IN1(n7654), .IN2(g185), .IN3(test_so45), .QN(n12026) );
  NAND3X0 U12447 ( .IN1(n12027), .IN2(n12028), .IN3(n12029), .QN(n7654) );
  NAND2X0 U12448 ( .IN1(g6944), .IN2(g1253), .QN(n12029) );
  NAND2X0 U12449 ( .IN1(g6750), .IN2(g1251), .QN(n12028) );
  NAND2X0 U12450 ( .IN1(g1236), .IN2(g1176), .QN(n12027) );
  NAND2X0 U12451 ( .IN1(g1236), .IN2(g1288), .QN(n12025) );
  NAND2X0 U12452 ( .IN1(g6944), .IN2(g1285), .QN(n12024) );
  NAND2X0 U12453 ( .IN1(n10142), .IN2(g1282), .QN(n12023) );
  NAND2X0 U12454 ( .IN1(n4371), .IN2(g1282), .QN(n12021) );
  NAND2X0 U12455 ( .IN1(n12030), .IN2(n12031), .QN(g24510) );
  NAND2X0 U12456 ( .IN1(n4316), .IN2(g1276), .QN(n12031) );
  NAND3X0 U12457 ( .IN1(n10239), .IN2(n9947), .IN3(g6944), .QN(n12030) );
  NAND2X0 U12458 ( .IN1(n12032), .IN2(n12033), .QN(g24508) );
  NAND2X0 U12459 ( .IN1(n4372), .IN2(g599), .QN(n12033) );
  NAND3X0 U12460 ( .IN1(n10250), .IN2(n9947), .IN3(g6642), .QN(n12032) );
  NAND2X0 U12461 ( .IN1(n12034), .IN2(n12035), .QN(g24507) );
  NAND2X0 U12462 ( .IN1(n12011), .IN2(n10334), .QN(n12035) );
  INVX0 U12463 ( .INP(n12036), .ZN(n12011) );
  NAND2X0 U12464 ( .IN1(n4313), .IN2(g593), .QN(n12034) );
  NAND2X0 U12465 ( .IN1(n12037), .IN2(n12038), .QN(g24501) );
  NAND2X0 U12466 ( .IN1(n4371), .IN2(g1273), .QN(n12038) );
  NAND3X0 U12467 ( .IN1(n10239), .IN2(n9947), .IN3(n10142), .QN(n12037) );
  NAND4X0 U12468 ( .IN1(n12039), .IN2(n12040), .IN3(n12041), .IN4(n12042), 
        .QN(n10239) );
  NAND3X0 U12469 ( .IN1(g185), .IN2(g1210), .IN3(n7655), .QN(n12042) );
  NAND3X0 U12470 ( .IN1(n12043), .IN2(n12044), .IN3(n12045), .QN(n7655) );
  NAND2X0 U12471 ( .IN1(n10142), .IN2(g1255), .QN(n12045) );
  NAND2X0 U12472 ( .IN1(g1236), .IN2(g1259), .QN(n12044) );
  NAND2X0 U12473 ( .IN1(g6944), .IN2(g1257), .QN(n12043) );
  NAND2X0 U12474 ( .IN1(g6750), .IN2(g1273), .QN(n12041) );
  NAND2X0 U12475 ( .IN1(g1236), .IN2(g1279), .QN(n12040) );
  NAND2X0 U12476 ( .IN1(g6944), .IN2(g1276), .QN(n12039) );
  NAND2X0 U12477 ( .IN1(n12046), .IN2(n12047), .QN(g24499) );
  NAND3X0 U12478 ( .IN1(n10250), .IN2(n9947), .IN3(g6485), .QN(n12047) );
  NAND4X0 U12479 ( .IN1(n12048), .IN2(n12049), .IN3(n12050), .IN4(n12051), 
        .QN(n10250) );
  NAND3X0 U12480 ( .IN1(g185), .IN2(g542), .IN3(n8376), .QN(n12051) );
  NAND3X0 U12481 ( .IN1(n12052), .IN2(n12053), .IN3(n12054), .QN(n8376) );
  NAND2X0 U12482 ( .IN1(g6642), .IN2(g567), .QN(n12054) );
  NAND2X0 U12483 ( .IN1(n10242), .IN2(g565), .QN(n12053) );
  NAND2X0 U12484 ( .IN1(g550), .IN2(g489), .QN(n12052) );
  NAND2X0 U12485 ( .IN1(g6485), .IN2(g596), .QN(n12050) );
  NAND2X0 U12486 ( .IN1(g550), .IN2(g602), .QN(n12049) );
  NAND2X0 U12487 ( .IN1(g6642), .IN2(g599), .QN(n12048) );
  NAND2X0 U12488 ( .IN1(n4298), .IN2(g596), .QN(n12046) );
  NAND2X0 U12489 ( .IN1(n12055), .IN2(n12056), .QN(g24498) );
  NAND2X0 U12490 ( .IN1(n4372), .IN2(g590), .QN(n12056) );
  NAND3X0 U12491 ( .IN1(n10334), .IN2(n9947), .IN3(g6642), .QN(n12055) );
  NAND2X0 U12492 ( .IN1(n12057), .IN2(n12058), .QN(g24491) );
  NAND2X0 U12493 ( .IN1(n4298), .IN2(g587), .QN(n12058) );
  NAND3X0 U12494 ( .IN1(n10334), .IN2(n9947), .IN3(n10242), .QN(n12057) );
  NAND4X0 U12495 ( .IN1(n12059), .IN2(n12060), .IN3(n12061), .IN4(n12062), 
        .QN(n10334) );
  NAND3X0 U12496 ( .IN1(g185), .IN2(g524), .IN3(n8351), .QN(n12062) );
  NAND3X0 U12497 ( .IN1(n12063), .IN2(n12064), .IN3(n12065), .QN(n8351) );
  NAND2X0 U12498 ( .IN1(g6642), .IN2(g571), .QN(n12065) );
  NAND2X0 U12499 ( .IN1(g6485), .IN2(g569), .QN(n12064) );
  NAND2X0 U12500 ( .IN1(g550), .IN2(g573), .QN(n12063) );
  NAND2X0 U12501 ( .IN1(n10242), .IN2(g587), .QN(n12061) );
  NAND2X0 U12502 ( .IN1(g550), .IN2(g593), .QN(n12060) );
  NAND2X0 U12503 ( .IN1(g6642), .IN2(g590), .QN(n12059) );
  AND3X1 U12504 ( .IN1(n12066), .IN2(n7778), .IN3(n11939), .Q(g24476) );
  NAND3X0 U12505 ( .IN1(g2924), .IN2(g2917), .IN3(n12067), .QN(n11939) );
  OR2X1 U12506 ( .IN1(n12068), .IN2(g2924), .Q(n12066) );
  NOR2X0 U12507 ( .IN1(n4479), .IN2(n7781), .QN(n12068) );
  INVX0 U12508 ( .INP(n12067), .ZN(n7781) );
  NOR2X0 U12509 ( .IN1(n7777), .IN2(n12069), .QN(g24473) );
  XOR2X1 U12510 ( .IN1(n7048), .IN2(n11936), .Q(n12069) );
  NOR3X0 U12511 ( .IN1(n11933), .IN2(n4101), .IN3(n11935), .QN(g24446) );
  NOR2X0 U12512 ( .IN1(n4102), .IN2(n4480), .QN(n11935) );
  OR2X1 U12513 ( .IN1(n12070), .IN2(n4350), .Q(n4102) );
  NOR2X0 U12514 ( .IN1(n11109), .IN2(n12071), .QN(g24445) );
  XNOR2X1 U12515 ( .IN1(n6430), .IN2(n4066), .Q(n12071) );
  NOR3X0 U12516 ( .IN1(n12072), .IN2(n10335), .IN3(n11113), .QN(g24438) );
  INVX0 U12517 ( .INP(n11115), .ZN(n11113) );
  NAND3X0 U12518 ( .IN1(g2720), .IN2(g2727), .IN3(n12073), .QN(n11115) );
  NOR2X0 U12519 ( .IN1(n12074), .IN2(g2720), .QN(n12072) );
  NOR2X0 U12520 ( .IN1(n4419), .IN2(n12075), .QN(n12074) );
  NOR3X0 U12521 ( .IN1(n12076), .IN2(n10339), .IN3(n11132), .QN(g24434) );
  NOR3X0 U12522 ( .IN1(n4410), .IN2(n4420), .IN3(n12077), .QN(n11132) );
  NOR2X0 U12523 ( .IN1(n12078), .IN2(g2026), .QN(n12076) );
  NOR2X0 U12524 ( .IN1(n4420), .IN2(n12077), .QN(n12078) );
  NOR3X0 U12525 ( .IN1(n12079), .IN2(n10343), .IN3(n11203), .QN(g24430) );
  NOR3X0 U12526 ( .IN1(n4412), .IN2(n4421), .IN3(n12080), .QN(n11203) );
  NOR2X0 U12527 ( .IN1(n12081), .IN2(g1332), .QN(n12079) );
  NOR2X0 U12528 ( .IN1(n4421), .IN2(n12080), .QN(n12081) );
  NOR3X0 U12529 ( .IN1(n12082), .IN2(n9912), .IN3(n11274), .QN(g24426) );
  INVX0 U12530 ( .INP(n11276), .ZN(n11274) );
  NAND3X0 U12531 ( .IN1(g646), .IN2(g653), .IN3(n12083), .QN(n11276) );
  NOR2X0 U12532 ( .IN1(n12084), .IN2(g646), .QN(n12082) );
  NOR2X0 U12533 ( .IN1(n4422), .IN2(n12085), .QN(n12084) );
  NAND2X0 U12534 ( .IN1(n12086), .IN2(n12087), .QN(g24250) );
  NAND2X0 U12535 ( .IN1(n4463), .IN2(g2546), .QN(n12087) );
  NAND2X0 U12536 ( .IN1(n10781), .IN2(g2560), .QN(n12086) );
  NAND2X0 U12537 ( .IN1(n12088), .IN2(n12089), .QN(g24243) );
  NAND2X0 U12538 ( .IN1(n4464), .IN2(g1852), .QN(n12089) );
  NAND2X0 U12539 ( .IN1(n10862), .IN2(g1866), .QN(n12088) );
  NAND2X0 U12540 ( .IN1(n12090), .IN2(n12091), .QN(g24238) );
  NAND2X0 U12541 ( .IN1(n4463), .IN2(g2554), .QN(n12091) );
  NAND2X0 U12542 ( .IN1(n9127), .IN2(g2560), .QN(n12090) );
  NAND2X0 U12543 ( .IN1(n12092), .IN2(n12093), .QN(g24237) );
  NAND2X0 U12544 ( .IN1(n4455), .IN2(g2543), .QN(n12093) );
  NAND2X0 U12545 ( .IN1(n10781), .IN2(g8167), .QN(n12092) );
  NAND2X0 U12546 ( .IN1(n12094), .IN2(n12095), .QN(g24235) );
  NAND2X0 U12547 ( .IN1(n4465), .IN2(g1158), .QN(n12095) );
  NAND2X0 U12548 ( .IN1(n10942), .IN2(g1172), .QN(n12094) );
  NAND2X0 U12549 ( .IN1(n12096), .IN2(n12097), .QN(g24231) );
  NAND2X0 U12550 ( .IN1(n4464), .IN2(g1860), .QN(n12097) );
  NAND2X0 U12551 ( .IN1(n9163), .IN2(g1866), .QN(n12096) );
  NAND2X0 U12552 ( .IN1(n12098), .IN2(n12099), .QN(g24230) );
  NAND2X0 U12553 ( .IN1(n4457), .IN2(g1849), .QN(n12099) );
  NAND2X0 U12554 ( .IN1(n10862), .IN2(g8082), .QN(n12098) );
  NAND2X0 U12555 ( .IN1(n12100), .IN2(n12101), .QN(g24228) );
  NAND2X0 U12556 ( .IN1(n4466), .IN2(g471), .QN(n12101) );
  NAND2X0 U12557 ( .IN1(n10955), .IN2(g485), .QN(n12100) );
  NAND2X0 U12558 ( .IN1(n12102), .IN2(n12103), .QN(g24226) );
  NAND2X0 U12559 ( .IN1(n4455), .IN2(g2553), .QN(n12103) );
  NAND2X0 U12560 ( .IN1(n9127), .IN2(g8167), .QN(n12102) );
  NAND2X0 U12561 ( .IN1(n12104), .IN2(n12105), .QN(g24225) );
  NAND2X0 U12562 ( .IN1(n4456), .IN2(g2540), .QN(n12105) );
  NAND2X0 U12563 ( .IN1(n10781), .IN2(g8087), .QN(n12104) );
  NOR2X0 U12564 ( .IN1(n8820), .IN2(n8824), .QN(n10781) );
  NAND2X0 U12565 ( .IN1(n8829), .IN2(n8825), .QN(n8820) );
  INVX0 U12566 ( .INP(n8839), .ZN(n8825) );
  NAND2X0 U12567 ( .IN1(n12106), .IN2(n12107), .QN(g24223) );
  NAND2X0 U12568 ( .IN1(n4465), .IN2(g1166), .QN(n12107) );
  NAND2X0 U12569 ( .IN1(n9194), .IN2(g1172), .QN(n12106) );
  NAND2X0 U12570 ( .IN1(n12108), .IN2(n12109), .QN(g24222) );
  NAND2X0 U12571 ( .IN1(n4459), .IN2(g1155), .QN(n12109) );
  NAND2X0 U12572 ( .IN1(n10942), .IN2(g8007), .QN(n12108) );
  NAND2X0 U12573 ( .IN1(n12110), .IN2(n12111), .QN(g24219) );
  NAND2X0 U12574 ( .IN1(n4457), .IN2(g1859), .QN(n12111) );
  NAND2X0 U12575 ( .IN1(n9163), .IN2(g8082), .QN(n12110) );
  NAND2X0 U12576 ( .IN1(n12112), .IN2(n12113), .QN(g24218) );
  NAND2X0 U12577 ( .IN1(n4458), .IN2(g1846), .QN(n12113) );
  NAND2X0 U12578 ( .IN1(n10862), .IN2(g8012), .QN(n12112) );
  NOR2X0 U12579 ( .IN1(n8471), .IN2(n8475), .QN(n10862) );
  NAND2X0 U12580 ( .IN1(n8480), .IN2(n8476), .QN(n8471) );
  INVX0 U12581 ( .INP(n8491), .ZN(n8476) );
  NAND2X0 U12582 ( .IN1(n12114), .IN2(n12115), .QN(g24216) );
  NAND2X0 U12583 ( .IN1(n4466), .IN2(g479), .QN(n12115) );
  NAND2X0 U12584 ( .IN1(n9230), .IN2(g485), .QN(n12114) );
  NAND2X0 U12585 ( .IN1(n12116), .IN2(n12117), .QN(g24215) );
  NAND2X0 U12586 ( .IN1(n10955), .IN2(g7956), .QN(n12117) );
  NAND2X0 U12587 ( .IN1(test_so24), .IN2(n4461), .QN(n12116) );
  NAND2X0 U12588 ( .IN1(n12118), .IN2(n12119), .QN(g24214) );
  NAND2X0 U12589 ( .IN1(n4456), .IN2(g2552), .QN(n12119) );
  NAND2X0 U12590 ( .IN1(n9127), .IN2(g8087), .QN(n12118) );
  INVX0 U12591 ( .INP(n9283), .ZN(n9127) );
  NAND3X0 U12592 ( .IN1(n8824), .IN2(n8839), .IN3(n8829), .QN(n9283) );
  INVX0 U12593 ( .INP(n8815), .ZN(n8829) );
  NAND2X0 U12594 ( .IN1(n12120), .IN2(n12121), .QN(g24213) );
  NAND2X0 U12595 ( .IN1(n4459), .IN2(g1165), .QN(n12121) );
  NAND2X0 U12596 ( .IN1(n9194), .IN2(g8007), .QN(n12120) );
  NAND2X0 U12597 ( .IN1(n12122), .IN2(n12123), .QN(g24212) );
  NAND2X0 U12598 ( .IN1(n4460), .IN2(g1152), .QN(n12123) );
  NAND2X0 U12599 ( .IN1(n10942), .IN2(g7961), .QN(n12122) );
  NOR2X0 U12600 ( .IN1(n8358), .IN2(n8338), .QN(n10942) );
  NAND2X0 U12601 ( .IN1(n8332), .IN2(n8342), .QN(n8358) );
  INVX0 U12602 ( .INP(n8344), .ZN(n8332) );
  NAND2X0 U12603 ( .IN1(n12124), .IN2(n12125), .QN(g24209) );
  NAND2X0 U12604 ( .IN1(n4463), .IN2(g2536), .QN(n12125) );
  NAND2X0 U12605 ( .IN1(n12126), .IN2(g2560), .QN(n12124) );
  NAND2X0 U12606 ( .IN1(n12127), .IN2(n12128), .QN(g24208) );
  NAND2X0 U12607 ( .IN1(n4458), .IN2(g1858), .QN(n12128) );
  NAND2X0 U12608 ( .IN1(n9163), .IN2(g8012), .QN(n12127) );
  INVX0 U12609 ( .INP(n9295), .ZN(n9163) );
  NAND3X0 U12610 ( .IN1(n8475), .IN2(n8491), .IN3(n8480), .QN(n9295) );
  INVX0 U12611 ( .INP(n8466), .ZN(n8480) );
  NAND2X0 U12612 ( .IN1(n12129), .IN2(n12130), .QN(g24207) );
  NAND2X0 U12613 ( .IN1(n4461), .IN2(g478), .QN(n12130) );
  NAND2X0 U12614 ( .IN1(n9230), .IN2(g7956), .QN(n12129) );
  NAND2X0 U12615 ( .IN1(n12131), .IN2(n12132), .QN(g24206) );
  NAND2X0 U12616 ( .IN1(g465), .IN2(n7268), .QN(n12132) );
  NAND2X0 U12617 ( .IN1(test_so23), .IN2(n10955), .QN(n12131) );
  NOR2X0 U12618 ( .IN1(n8514), .IN2(n8518), .QN(n10955) );
  NAND2X0 U12619 ( .IN1(n8519), .IN2(n8523), .QN(n8514) );
  INVX0 U12620 ( .INP(n8534), .ZN(n8519) );
  NAND2X0 U12621 ( .IN1(n12133), .IN2(n12134), .QN(g24182) );
  NAND2X0 U12622 ( .IN1(n4464), .IN2(g1842), .QN(n12134) );
  NAND2X0 U12623 ( .IN1(n12135), .IN2(g1866), .QN(n12133) );
  NAND2X0 U12624 ( .IN1(n12136), .IN2(n12137), .QN(g24181) );
  NAND2X0 U12625 ( .IN1(n4460), .IN2(g1164), .QN(n12137) );
  NAND2X0 U12626 ( .IN1(n9194), .IN2(g7961), .QN(n12136) );
  INVX0 U12627 ( .INP(n9307), .ZN(n9194) );
  NAND3X0 U12628 ( .IN1(n8338), .IN2(n8344), .IN3(n8342), .QN(n9307) );
  INVX0 U12629 ( .INP(n8340), .ZN(n8342) );
  NAND2X0 U12630 ( .IN1(n12138), .IN2(n12139), .QN(g24179) );
  NAND2X0 U12631 ( .IN1(n4465), .IN2(g1148), .QN(n12139) );
  NAND2X0 U12632 ( .IN1(n12140), .IN2(g1172), .QN(n12138) );
  NAND2X0 U12633 ( .IN1(n12141), .IN2(n12142), .QN(g24178) );
  NAND2X0 U12634 ( .IN1(g477), .IN2(n7268), .QN(n12142) );
  NAND2X0 U12635 ( .IN1(test_so23), .IN2(n9230), .QN(n12141) );
  INVX0 U12636 ( .INP(n9316), .ZN(n9230) );
  NAND3X0 U12637 ( .IN1(n8518), .IN2(n8534), .IN3(n8523), .QN(n9316) );
  INVX0 U12638 ( .INP(n8509), .ZN(n8523) );
  NAND2X0 U12639 ( .IN1(n12143), .IN2(n12144), .QN(g24174) );
  NAND2X0 U12640 ( .IN1(n4466), .IN2(g461), .QN(n12144) );
  NAND2X0 U12641 ( .IN1(n12145), .IN2(g485), .QN(n12143) );
  NAND2X0 U12642 ( .IN1(n12146), .IN2(n12147), .QN(g24092) );
  NAND2X0 U12643 ( .IN1(g3229), .IN2(n4483), .QN(n12147) );
  NAND2X0 U12644 ( .IN1(n7882), .IN2(g2380), .QN(n12146) );
  NAND2X0 U12645 ( .IN1(n12148), .IN2(n12149), .QN(g24083) );
  NAND2X0 U12646 ( .IN1(g3229), .IN2(n4484), .QN(n12149) );
  NAND2X0 U12647 ( .IN1(n7882), .IN2(g1686), .QN(n12148) );
  INVX0 U12648 ( .INP(g3229), .ZN(n7882) );
  NAND2X0 U12649 ( .IN1(n12150), .IN2(n12151), .QN(g24072) );
  NAND2X0 U12650 ( .IN1(g3229), .IN2(n4486), .QN(n12151) );
  OR2X1 U12651 ( .IN1(g3229), .IN2(n6997), .Q(n12150) );
  NAND2X0 U12652 ( .IN1(n12152), .IN2(n12153), .QN(g24059) );
  NAND2X0 U12653 ( .IN1(g3229), .IN2(n4485), .QN(n12153) );
  OR2X1 U12654 ( .IN1(g3229), .IN2(n6710), .Q(n12152) );
  NAND2X0 U12655 ( .IN1(n12154), .IN2(n12155), .QN(g23418) );
  NAND2X0 U12656 ( .IN1(n4455), .IN2(g2533), .QN(n12155) );
  NAND2X0 U12657 ( .IN1(n12126), .IN2(g8167), .QN(n12154) );
  NAND2X0 U12658 ( .IN1(n12156), .IN2(n12157), .QN(g23413) );
  NAND2X0 U12659 ( .IN1(n12135), .IN2(g8082), .QN(n12157) );
  NAND2X0 U12660 ( .IN1(test_so65), .IN2(n4457), .QN(n12156) );
  NAND2X0 U12661 ( .IN1(n12158), .IN2(n12159), .QN(g23407) );
  NAND2X0 U12662 ( .IN1(n4456), .IN2(g2530), .QN(n12159) );
  NAND2X0 U12663 ( .IN1(n12126), .IN2(g8087), .QN(n12158) );
  INVX0 U12664 ( .INP(n7772), .ZN(n12126) );
  NAND3X0 U12665 ( .IN1(n8815), .IN2(n8839), .IN3(n8819), .QN(n7772) );
  INVX0 U12666 ( .INP(n8824), .ZN(n8819) );
  NAND3X0 U12667 ( .IN1(n12160), .IN2(n12161), .IN3(n12162), .QN(n8824) );
  NAND2X0 U12668 ( .IN1(n6533), .IN2(n8449), .QN(n12162) );
  NAND2X0 U12669 ( .IN1(n6544), .IN2(n8841), .QN(n12161) );
  NAND2X0 U12670 ( .IN1(n6545), .IN2(n8456), .QN(n12160) );
  NAND3X0 U12671 ( .IN1(n12163), .IN2(n12164), .IN3(n12165), .QN(n8839) );
  NAND2X0 U12672 ( .IN1(n6531), .IN2(n8449), .QN(n12165) );
  NAND2X0 U12673 ( .IN1(n6540), .IN2(n8841), .QN(n12164) );
  NAND2X0 U12674 ( .IN1(n6541), .IN2(n8456), .QN(n12163) );
  NAND3X0 U12675 ( .IN1(n12166), .IN2(n12167), .IN3(n12168), .QN(n8815) );
  NAND2X0 U12676 ( .IN1(n6532), .IN2(n8449), .QN(n12168) );
  INVX0 U12677 ( .INP(n4524), .ZN(n8449) );
  NAND2X0 U12678 ( .IN1(n6542), .IN2(n8841), .QN(n12167) );
  INVX0 U12679 ( .INP(n4509), .ZN(n8841) );
  NAND2X0 U12680 ( .IN1(n6543), .IN2(n8456), .QN(n12166) );
  INVX0 U12681 ( .INP(n4516), .ZN(n8456) );
  NAND2X0 U12682 ( .IN1(n12169), .IN2(n12170), .QN(g23406) );
  NAND2X0 U12683 ( .IN1(n4459), .IN2(g1145), .QN(n12170) );
  NAND2X0 U12684 ( .IN1(n12140), .IN2(g8007), .QN(n12169) );
  NAND2X0 U12685 ( .IN1(n12171), .IN2(n12172), .QN(g23400) );
  NAND2X0 U12686 ( .IN1(n4458), .IN2(g1836), .QN(n12172) );
  NAND2X0 U12687 ( .IN1(n12135), .IN2(g8012), .QN(n12171) );
  INVX0 U12688 ( .INP(n7736), .ZN(n12135) );
  NAND3X0 U12689 ( .IN1(n8466), .IN2(n8491), .IN3(n8470), .QN(n7736) );
  INVX0 U12690 ( .INP(n8475), .ZN(n8470) );
  NAND3X0 U12691 ( .IN1(n12173), .IN2(n12174), .IN3(n12175), .QN(n8475) );
  NAND2X0 U12692 ( .IN1(n6536), .IN2(n8459), .QN(n12175) );
  NAND2X0 U12693 ( .IN1(n6550), .IN2(n8453), .QN(n12174) );
  NAND2X0 U12694 ( .IN1(n6551), .IN2(n8494), .QN(n12173) );
  NAND3X0 U12695 ( .IN1(n12176), .IN2(n12177), .IN3(n12178), .QN(n8491) );
  NAND2X0 U12696 ( .IN1(n6534), .IN2(n8459), .QN(n12178) );
  NAND2X0 U12697 ( .IN1(n6546), .IN2(n8453), .QN(n12177) );
  NAND2X0 U12698 ( .IN1(n6547), .IN2(n8494), .QN(n12176) );
  NAND3X0 U12699 ( .IN1(n12179), .IN2(n12180), .IN3(n12181), .QN(n8466) );
  NAND2X0 U12700 ( .IN1(n6535), .IN2(n8459), .QN(n12181) );
  INVX0 U12701 ( .INP(n4525), .ZN(n8459) );
  NAND2X0 U12702 ( .IN1(n6548), .IN2(n8453), .QN(n12180) );
  INVX0 U12703 ( .INP(n4511), .ZN(n8453) );
  NAND2X0 U12704 ( .IN1(n6549), .IN2(n8494), .QN(n12179) );
  INVX0 U12705 ( .INP(n4518), .ZN(n8494) );
  NAND2X0 U12706 ( .IN1(n12182), .IN2(n12183), .QN(g23399) );
  NAND2X0 U12707 ( .IN1(n4461), .IN2(g458), .QN(n12183) );
  NAND2X0 U12708 ( .IN1(n12145), .IN2(g7956), .QN(n12182) );
  NAND2X0 U12709 ( .IN1(n12184), .IN2(n12185), .QN(g23392) );
  NAND2X0 U12710 ( .IN1(n4460), .IN2(g1142), .QN(n12185) );
  NAND2X0 U12711 ( .IN1(n12140), .IN2(g7961), .QN(n12184) );
  INVX0 U12712 ( .INP(n7714), .ZN(n12140) );
  NAND3X0 U12713 ( .IN1(n8340), .IN2(n8344), .IN3(n8357), .QN(n7714) );
  INVX0 U12714 ( .INP(n8338), .ZN(n8357) );
  NAND3X0 U12715 ( .IN1(n12186), .IN2(n12187), .IN3(n12188), .QN(n8338) );
  NAND2X0 U12716 ( .IN1(n6555), .IN2(g1088), .QN(n12188) );
  NAND2X0 U12717 ( .IN1(n6556), .IN2(g5472), .QN(n12187) );
  NAND2X0 U12718 ( .IN1(n6539), .IN2(g6712), .QN(n12186) );
  NAND3X0 U12719 ( .IN1(n12189), .IN2(n12190), .IN3(n12191), .QN(n8344) );
  OR2X1 U12720 ( .IN1(n4381), .IN2(test_so39), .Q(n12191) );
  NAND2X0 U12721 ( .IN1(n6552), .IN2(g5472), .QN(n12190) );
  NAND2X0 U12722 ( .IN1(n6537), .IN2(g6712), .QN(n12189) );
  NAND3X0 U12723 ( .IN1(n12192), .IN2(n12193), .IN3(n12194), .QN(n8340) );
  NAND2X0 U12724 ( .IN1(n6553), .IN2(g1088), .QN(n12194) );
  NAND2X0 U12725 ( .IN1(n6554), .IN2(g5472), .QN(n12193) );
  NAND2X0 U12726 ( .IN1(n6538), .IN2(g6712), .QN(n12192) );
  NAND2X0 U12727 ( .IN1(n12195), .IN2(n12196), .QN(g23385) );
  NAND2X0 U12728 ( .IN1(g455), .IN2(n7268), .QN(n12196) );
  NAND2X0 U12729 ( .IN1(n12145), .IN2(test_so23), .QN(n12195) );
  INVX0 U12730 ( .INP(n7677), .ZN(n12145) );
  NAND3X0 U12731 ( .IN1(n8509), .IN2(n8534), .IN3(n8513), .QN(n7677) );
  INVX0 U12732 ( .INP(n8518), .ZN(n8513) );
  NAND3X0 U12733 ( .IN1(n12197), .IN2(n12198), .IN3(n12199), .QN(n8518) );
  NAND2X0 U12734 ( .IN1(n6564), .IN2(n8537), .QN(n12199) );
  NAND2X0 U12735 ( .IN1(n6563), .IN2(n8861), .QN(n12198) );
  NAND2X0 U12736 ( .IN1(n6562), .IN2(n8500), .QN(n12197) );
  NAND3X0 U12737 ( .IN1(n12200), .IN2(n12201), .IN3(n12202), .QN(n8534) );
  NAND2X0 U12738 ( .IN1(n6559), .IN2(n8537), .QN(n12202) );
  NAND2X0 U12739 ( .IN1(n6558), .IN2(n8861), .QN(n12201) );
  INVX0 U12740 ( .INP(n4499), .ZN(n8861) );
  NAND2X0 U12741 ( .IN1(n6557), .IN2(n8500), .QN(n12200) );
  NAND3X0 U12742 ( .IN1(n12203), .IN2(n12204), .IN3(n12205), .QN(n8509) );
  NAND2X0 U12743 ( .IN1(n6561), .IN2(n8537), .QN(n12205) );
  INVX0 U12744 ( .INP(n4520), .ZN(n8537) );
  OR2X1 U12745 ( .IN1(n4499), .IN2(test_so18), .Q(n12204) );
  NAND2X0 U12746 ( .IN1(n6560), .IN2(n8500), .QN(n12203) );
  INVX0 U12747 ( .INP(n4506), .ZN(n8500) );
  NOR2X0 U12748 ( .IN1(n11933), .IN2(n12206), .QN(g23359) );
  XNOR2X1 U12749 ( .IN1(n4350), .IN2(n12070), .Q(n12206) );
  NAND2X0 U12750 ( .IN1(n7828), .IN2(g3018), .QN(n12070) );
  INVX0 U12751 ( .INP(n7827), .ZN(n11933) );
  NAND2X0 U12752 ( .IN1(n11109), .IN2(n12207), .QN(n7827) );
  NAND2X0 U12753 ( .IN1(n12208), .IN2(n7825), .QN(n12207) );
  INVX0 U12754 ( .INP(g3234), .ZN(n7825) );
  NAND4X0 U12755 ( .IN1(n4480), .IN2(n4350), .IN3(g3018), .IN4(g3032), .QN(
        n12208) );
  INVX0 U12756 ( .INP(n11474), .ZN(n11109) );
  NOR3X0 U12757 ( .IN1(n7777), .IN2(n4122), .IN3(n11936), .QN(g23358) );
  NOR2X0 U12758 ( .IN1(n4123), .IN2(n4431), .QN(n11936) );
  OR2X1 U12759 ( .IN1(n12209), .IN2(n7049), .Q(n4123) );
  NOR2X0 U12760 ( .IN1(n11937), .IN2(n12210), .QN(g23357) );
  XOR2X1 U12761 ( .IN1(n4479), .IN2(n12067), .Q(n12210) );
  NOR2X0 U12762 ( .IN1(n7782), .IN2(n4482), .QN(n12067) );
  INVX0 U12763 ( .INP(n7778), .ZN(n11937) );
  NAND2X0 U12764 ( .IN1(n7777), .IN2(n12211), .QN(n7778) );
  NAND2X0 U12765 ( .IN1(n13231), .IN2(n12212), .QN(n12211) );
  OR4X1 U12766 ( .IN1(g2917), .IN2(g2924), .IN3(n4482), .IN4(n6995), .Q(n12212) );
  NOR2X0 U12767 ( .IN1(n10335), .IN2(n12213), .QN(g23348) );
  XOR2X1 U12768 ( .IN1(g2727), .IN2(n12075), .Q(n12213) );
  NOR2X0 U12769 ( .IN1(n10339), .IN2(n12214), .QN(g23339) );
  XNOR2X1 U12770 ( .IN1(n4420), .IN2(n12077), .Q(n12214) );
  AND3X1 U12771 ( .IN1(n12215), .IN2(n4066), .IN3(n11474), .Q(g23330) );
  NOR2X0 U12772 ( .IN1(g3234), .IN2(n7828), .QN(n11474) );
  NOR2X0 U12773 ( .IN1(n12216), .IN2(n6431), .QN(n7828) );
  NAND3X0 U12774 ( .IN1(g3006), .IN2(n7909), .IN3(n11475), .QN(n4066) );
  NAND2X0 U12775 ( .IN1(n6428), .IN2(n12217), .QN(n12215) );
  NAND2X0 U12776 ( .IN1(n11475), .IN2(n7909), .QN(n12217) );
  NOR2X0 U12777 ( .IN1(n6432), .IN2(n6431), .QN(n11475) );
  NOR2X0 U12778 ( .IN1(n10343), .IN2(n12218), .QN(g23329) );
  XNOR2X1 U12779 ( .IN1(n4421), .IN2(n12080), .Q(n12218) );
  NOR2X0 U12780 ( .IN1(n9912), .IN2(n12219), .QN(g23324) );
  XOR2X1 U12781 ( .IN1(g653), .IN2(n12085), .Q(n12219) );
  NAND2X0 U12782 ( .IN1(n12220), .IN2(n12221), .QN(g23137) );
  NAND2X0 U12783 ( .IN1(n4464), .IN2(g1869), .QN(n12221) );
  NAND2X0 U12784 ( .IN1(n10405), .IN2(g1866), .QN(n12220) );
  NOR3X0 U12785 ( .IN1(n12222), .IN2(n9912), .IN3(n12083), .QN(g23136) );
  INVX0 U12786 ( .INP(n12085), .ZN(n12083) );
  NAND3X0 U12787 ( .IN1(g640), .IN2(g633), .IN3(n12223), .QN(n12085) );
  NOR2X0 U12788 ( .IN1(n12224), .IN2(g633), .QN(n12222) );
  AND2X1 U12789 ( .IN1(g640), .IN2(n12223), .Q(n12224) );
  NAND2X0 U12790 ( .IN1(n12225), .IN2(n12226), .QN(g23133) );
  NAND2X0 U12791 ( .IN1(n4455), .IN2(g2562), .QN(n12226) );
  NAND2X0 U12792 ( .IN1(n10381), .IN2(g8167), .QN(n12225) );
  NAND2X0 U12793 ( .IN1(n12227), .IN2(n12228), .QN(g23132) );
  NAND2X0 U12794 ( .IN1(n4456), .IN2(g2555), .QN(n12228) );
  NAND2X0 U12795 ( .IN1(n9342), .IN2(g8087), .QN(n12227) );
  NAND2X0 U12796 ( .IN1(n12229), .IN2(n12230), .QN(g23126) );
  NAND2X0 U12797 ( .IN1(n4465), .IN2(g1175), .QN(n12230) );
  NAND2X0 U12798 ( .IN1(n10429), .IN2(g1172), .QN(n12229) );
  NAND2X0 U12799 ( .IN1(n12231), .IN2(n12232), .QN(g23124) );
  NAND2X0 U12800 ( .IN1(n4457), .IN2(g1868), .QN(n12232) );
  NAND2X0 U12801 ( .IN1(n10405), .IN2(g8082), .QN(n12231) );
  NAND2X0 U12802 ( .IN1(n12233), .IN2(n12234), .QN(g23123) );
  NAND2X0 U12803 ( .IN1(n4458), .IN2(g1861), .QN(n12234) );
  NAND2X0 U12804 ( .IN1(n9358), .IN2(g8012), .QN(n12233) );
  NAND2X0 U12805 ( .IN1(n12235), .IN2(n12236), .QN(g23117) );
  NAND2X0 U12806 ( .IN1(n4466), .IN2(g488), .QN(n12236) );
  NAND2X0 U12807 ( .IN1(n10448), .IN2(g485), .QN(n12235) );
  NAND2X0 U12808 ( .IN1(n12237), .IN2(n12238), .QN(g23114) );
  NAND2X0 U12809 ( .IN1(n4456), .IN2(g2561), .QN(n12238) );
  NAND2X0 U12810 ( .IN1(n10381), .IN2(g8087), .QN(n12237) );
  NAND2X0 U12811 ( .IN1(n12239), .IN2(n12240), .QN(g23111) );
  NAND2X0 U12812 ( .IN1(test_so44), .IN2(n4459), .QN(n12240) );
  NAND2X0 U12813 ( .IN1(n10429), .IN2(g8007), .QN(n12239) );
  NAND2X0 U12814 ( .IN1(n12241), .IN2(n12242), .QN(g23110) );
  NAND2X0 U12815 ( .IN1(n4460), .IN2(g1167), .QN(n12242) );
  NAND2X0 U12816 ( .IN1(n9373), .IN2(g7961), .QN(n12241) );
  NAND2X0 U12817 ( .IN1(n12243), .IN2(n12244), .QN(g23097) );
  NAND2X0 U12818 ( .IN1(n4458), .IN2(g1867), .QN(n12244) );
  NAND2X0 U12819 ( .IN1(n10405), .IN2(g8012), .QN(n12243) );
  NAND3X0 U12820 ( .IN1(n12245), .IN2(n12246), .IN3(n12247), .QN(n10405) );
  NAND2X0 U12821 ( .IN1(g5511), .IN2(g1819), .QN(n12247) );
  NAND2X0 U12822 ( .IN1(test_so59), .IN2(n4618), .QN(n12246) );
  NAND2X0 U12823 ( .IN1(g7014), .IN2(g1822), .QN(n12245) );
  NAND2X0 U12824 ( .IN1(n12248), .IN2(n12249), .QN(g23093) );
  NAND2X0 U12825 ( .IN1(n4461), .IN2(g487), .QN(n12249) );
  NAND2X0 U12826 ( .IN1(n10448), .IN2(g7956), .QN(n12248) );
  NAND2X0 U12827 ( .IN1(n12250), .IN2(n12251), .QN(g23092) );
  NAND2X0 U12828 ( .IN1(g480), .IN2(n7268), .QN(n12251) );
  NAND2X0 U12829 ( .IN1(test_so23), .IN2(n9386), .QN(n12250) );
  NAND2X0 U12830 ( .IN1(n12252), .IN2(n12253), .QN(g23081) );
  NAND2X0 U12831 ( .IN1(n4460), .IN2(g1173), .QN(n12253) );
  NAND2X0 U12832 ( .IN1(n10429), .IN2(g7961), .QN(n12252) );
  NAND3X0 U12833 ( .IN1(n12254), .IN2(n12255), .IN3(n12256), .QN(n10429) );
  NAND2X0 U12834 ( .IN1(g1088), .IN2(g1131), .QN(n12256) );
  NAND2X0 U12835 ( .IN1(g5472), .IN2(g1125), .QN(n12255) );
  NAND2X0 U12836 ( .IN1(g6712), .IN2(g1128), .QN(n12254) );
  NAND2X0 U12837 ( .IN1(n12257), .IN2(n12258), .QN(g23076) );
  NAND2X0 U12838 ( .IN1(n4463), .IN2(g2539), .QN(n12258) );
  NAND2X0 U12839 ( .IN1(n9342), .IN2(g2560), .QN(n12257) );
  NAND2X0 U12840 ( .IN1(n12259), .IN2(n12260), .QN(g23067) );
  NAND2X0 U12841 ( .IN1(g486), .IN2(n7268), .QN(n12260) );
  NAND2X0 U12842 ( .IN1(test_so23), .IN2(n10448), .QN(n12259) );
  NAND3X0 U12843 ( .IN1(n12261), .IN2(n12262), .IN3(n12263), .QN(n10448) );
  NAND2X0 U12844 ( .IN1(g5437), .IN2(g438), .QN(n12263) );
  NAND2X0 U12845 ( .IN1(n4640), .IN2(g444), .QN(n12262) );
  NAND2X0 U12846 ( .IN1(g6447), .IN2(g441), .QN(n12261) );
  NAND2X0 U12847 ( .IN1(n12264), .IN2(n12265), .QN(g23058) );
  NAND2X0 U12848 ( .IN1(n4464), .IN2(g1845), .QN(n12265) );
  NAND2X0 U12849 ( .IN1(n9358), .IN2(g1866), .QN(n12264) );
  NAND2X0 U12850 ( .IN1(n12266), .IN2(n12267), .QN(g23047) );
  NAND2X0 U12851 ( .IN1(n4455), .IN2(g2559), .QN(n12267) );
  NAND2X0 U12852 ( .IN1(n9342), .IN2(g8167), .QN(n12266) );
  INVX0 U12853 ( .INP(n4285), .ZN(n9342) );
  NAND3X0 U12854 ( .IN1(n12268), .IN2(n12269), .IN3(n12270), .QN(n4285) );
  NAND2X0 U12855 ( .IN1(g5555), .IN2(g2492), .QN(n12270) );
  NAND2X0 U12856 ( .IN1(n4606), .IN2(g2498), .QN(n12269) );
  NAND2X0 U12857 ( .IN1(g7264), .IN2(g2495), .QN(n12268) );
  NAND2X0 U12858 ( .IN1(n12271), .IN2(n12272), .QN(g23039) );
  NAND2X0 U12859 ( .IN1(n4465), .IN2(g1151), .QN(n12272) );
  NAND2X0 U12860 ( .IN1(n9373), .IN2(g1172), .QN(n12271) );
  NAND2X0 U12861 ( .IN1(n12273), .IN2(n12274), .QN(g23030) );
  NAND2X0 U12862 ( .IN1(n4457), .IN2(g1865), .QN(n12274) );
  NAND2X0 U12863 ( .IN1(n9358), .IN2(g8082), .QN(n12273) );
  INVX0 U12864 ( .INP(n4284), .ZN(n9358) );
  NAND3X0 U12865 ( .IN1(n12275), .IN2(n12276), .IN3(n12277), .QN(n4284) );
  NAND2X0 U12866 ( .IN1(g5511), .IN2(g1798), .QN(n12277) );
  NAND2X0 U12867 ( .IN1(n4618), .IN2(g1804), .QN(n12276) );
  NAND2X0 U12868 ( .IN1(g7014), .IN2(g1801), .QN(n12275) );
  NAND2X0 U12869 ( .IN1(n12278), .IN2(n12279), .QN(g23022) );
  NAND2X0 U12870 ( .IN1(n4466), .IN2(g464), .QN(n12279) );
  NAND2X0 U12871 ( .IN1(n9386), .IN2(g485), .QN(n12278) );
  NAND2X0 U12872 ( .IN1(n12280), .IN2(n12281), .QN(g23014) );
  NAND2X0 U12873 ( .IN1(n4459), .IN2(g1171), .QN(n12281) );
  NAND2X0 U12874 ( .IN1(n9373), .IN2(g8007), .QN(n12280) );
  INVX0 U12875 ( .INP(n4283), .ZN(n9373) );
  NAND3X0 U12876 ( .IN1(n12282), .IN2(n12283), .IN3(n12284), .QN(n4283) );
  NAND2X0 U12877 ( .IN1(g1088), .IN2(g1110), .QN(n12284) );
  NAND2X0 U12878 ( .IN1(g5472), .IN2(g1104), .QN(n12283) );
  NAND2X0 U12879 ( .IN1(g6712), .IN2(g1107), .QN(n12282) );
  NAND2X0 U12880 ( .IN1(n12285), .IN2(n12286), .QN(g23000) );
  NAND2X0 U12881 ( .IN1(n4461), .IN2(g484), .QN(n12286) );
  NAND2X0 U12882 ( .IN1(n9386), .IN2(g7956), .QN(n12285) );
  INVX0 U12883 ( .INP(n4282), .ZN(n9386) );
  NAND3X0 U12884 ( .IN1(n12287), .IN2(n12288), .IN3(n12289), .QN(n4282) );
  NAND2X0 U12885 ( .IN1(g5437), .IN2(g417), .QN(n12289) );
  NAND2X0 U12886 ( .IN1(n4640), .IN2(g423), .QN(n12288) );
  NAND2X0 U12887 ( .IN1(g6447), .IN2(g420), .QN(n12287) );
  NAND2X0 U12888 ( .IN1(n12290), .IN2(n12291), .QN(g22687) );
  OR3X1 U12889 ( .IN1(n12292), .IN2(n4303), .IN3(n11351), .Q(n12291) );
  NAND2X0 U12890 ( .IN1(n12293), .IN2(n12294), .QN(n12290) );
  NAND2X0 U12891 ( .IN1(n7981), .IN2(n11351), .QN(n12293) );
  NAND3X0 U12892 ( .IN1(n12295), .IN2(n12296), .IN3(n12297), .QN(n11351) );
  NAND2X0 U12893 ( .IN1(g7390), .IN2(g2568), .QN(n12297) );
  NAND2X0 U12894 ( .IN1(g2624), .IN2(g2571), .QN(n12296) );
  NAND2X0 U12895 ( .IN1(n9246), .IN2(g2565), .QN(n12295) );
  NAND2X0 U12896 ( .IN1(n12298), .IN2(n12299), .QN(g22651) );
  OR3X1 U12897 ( .IN1(n8167), .IN2(n4297), .IN3(n11359), .Q(n12299) );
  NAND2X0 U12898 ( .IN1(n12300), .IN2(n12294), .QN(n12298) );
  NAND2X0 U12899 ( .IN1(n8173), .IN2(n11359), .QN(n12300) );
  NAND3X0 U12900 ( .IN1(n12301), .IN2(n12302), .IN3(n12303), .QN(n11359) );
  NAND2X0 U12901 ( .IN1(g1930), .IN2(g1877), .QN(n12303) );
  NAND2X0 U12902 ( .IN1(test_so68), .IN2(n9268), .QN(n12302) );
  NAND2X0 U12903 ( .IN1(g7194), .IN2(g1874), .QN(n12301) );
  NAND2X0 U12904 ( .IN1(n12304), .IN2(n12305), .QN(g22615) );
  OR3X1 U12905 ( .IN1(n12306), .IN2(n4304), .IN3(n11367), .Q(n12305) );
  NAND2X0 U12906 ( .IN1(n12307), .IN2(n12294), .QN(n12304) );
  NAND2X0 U12907 ( .IN1(n8285), .IN2(n11367), .QN(n12307) );
  NAND3X0 U12908 ( .IN1(n12308), .IN2(n12309), .IN3(n12310), .QN(n11367) );
  NAND2X0 U12909 ( .IN1(test_so47), .IN2(n10142), .QN(n12310) );
  NAND2X0 U12910 ( .IN1(g1236), .IN2(g1183), .QN(n12309) );
  NAND2X0 U12911 ( .IN1(g6944), .IN2(g1180), .QN(n12308) );
  NAND2X0 U12912 ( .IN1(n12311), .IN2(n12312), .QN(g22578) );
  OR3X1 U12913 ( .IN1(n7271), .IN2(n12313), .IN3(n11372), .Q(n12312) );
  NAND2X0 U12914 ( .IN1(n12314), .IN2(n12294), .QN(n12311) );
  NAND2X0 U12915 ( .IN1(n7851), .IN2(n11372), .QN(n12314) );
  NAND3X0 U12916 ( .IN1(n12315), .IN2(n12316), .IN3(n12317), .QN(n11372) );
  NAND2X0 U12917 ( .IN1(g6642), .IN2(g493), .QN(n12317) );
  NAND2X0 U12918 ( .IN1(g6485), .IN2(g490), .QN(n12316) );
  NAND2X0 U12919 ( .IN1(g550), .IN2(g496), .QN(n12315) );
  NOR2X0 U12920 ( .IN1(n12318), .IN2(n12319), .QN(g22299) );
  NOR2X0 U12921 ( .IN1(n11563), .IN2(test_so95), .QN(n12319) );
  NOR2X0 U12922 ( .IN1(n10335), .IN2(n12320), .QN(g22284) );
  AND2X1 U12923 ( .IN1(n12321), .IN2(n7226), .Q(n12320) );
  NOR2X0 U12924 ( .IN1(n12322), .IN2(n12323), .QN(g22280) );
  AND2X1 U12925 ( .IN1(n12324), .IN2(n7230), .Q(n12323) );
  NOR2X0 U12926 ( .IN1(n12325), .IN2(n12326), .QN(g22269) );
  AND2X1 U12927 ( .IN1(n12327), .IN2(n7162), .Q(n12326) );
  NOR2X0 U12928 ( .IN1(n10339), .IN2(n12328), .QN(g22267) );
  AND2X1 U12929 ( .IN1(n12329), .IN2(n7227), .Q(n12328) );
  NOR2X0 U12930 ( .IN1(n12330), .IN2(n12331), .QN(g22263) );
  NOR2X0 U12931 ( .IN1(n11632), .IN2(g1423), .QN(n12331) );
  NOR2X0 U12932 ( .IN1(n12332), .IN2(n12333), .QN(g22249) );
  AND2X1 U12933 ( .IN1(n12334), .IN2(n7163), .Q(n12333) );
  NOR2X0 U12934 ( .IN1(n10343), .IN2(n12335), .QN(g22247) );
  AND2X1 U12935 ( .IN1(n12336), .IN2(n7228), .Q(n12335) );
  NOR2X0 U12936 ( .IN1(n12337), .IN2(n12338), .QN(g22242) );
  AND2X1 U12937 ( .IN1(n12339), .IN2(n7232), .Q(n12338) );
  NOR2X0 U12938 ( .IN1(n12340), .IN2(n12341), .QN(g22234) );
  AND2X1 U12939 ( .IN1(n12342), .IN2(n7164), .Q(n12341) );
  NOR2X0 U12940 ( .IN1(n9912), .IN2(n12343), .QN(g22231) );
  AND2X1 U12941 ( .IN1(n12344), .IN2(n7229), .Q(n12343) );
  NOR2X0 U12942 ( .IN1(n12345), .IN2(n12346), .QN(g22218) );
  AND2X1 U12943 ( .IN1(n12347), .IN2(n7165), .Q(n12346) );
  NAND2X0 U12944 ( .IN1(n12348), .IN2(n12349), .QN(g22200) );
  NAND2X0 U12945 ( .IN1(n11946), .IN2(n4373), .QN(n12349) );
  OR2X1 U12946 ( .IN1(n11946), .IN2(n6796), .Q(n12348) );
  NAND2X0 U12947 ( .IN1(n12350), .IN2(n12351), .QN(g22194) );
  OR2X1 U12948 ( .IN1(n11946), .IN2(n6788), .Q(n12351) );
  NAND2X0 U12949 ( .IN1(n11946), .IN2(n8573), .QN(n12350) );
  NAND2X0 U12950 ( .IN1(n12352), .IN2(n12353), .QN(g22193) );
  NAND2X0 U12951 ( .IN1(n12354), .IN2(n4373), .QN(n12353) );
  OR2X1 U12952 ( .IN1(n12354), .IN2(n7177), .Q(n12352) );
  NAND2X0 U12953 ( .IN1(n12355), .IN2(n12356), .QN(g22192) );
  NAND2X0 U12954 ( .IN1(n11946), .IN2(n4377), .QN(n12356) );
  OR2X1 U12955 ( .IN1(n11946), .IN2(n6797), .Q(n12355) );
  NAND2X0 U12956 ( .IN1(n12357), .IN2(n12358), .QN(g22191) );
  NAND2X0 U12957 ( .IN1(n11948), .IN2(n4374), .QN(n12358) );
  OR2X1 U12958 ( .IN1(n11948), .IN2(n6807), .Q(n12357) );
  NAND2X0 U12959 ( .IN1(n12359), .IN2(n12360), .QN(g22185) );
  NAND2X0 U12960 ( .IN1(test_so75), .IN2(n12361), .QN(n12360) );
  NAND2X0 U12961 ( .IN1(n12354), .IN2(n8573), .QN(n12359) );
  NAND2X0 U12962 ( .IN1(n12362), .IN2(n12363), .QN(g22184) );
  OR2X1 U12963 ( .IN1(n11946), .IN2(n6779), .Q(n12363) );
  NAND2X0 U12964 ( .IN1(n9482), .IN2(n11946), .QN(n12362) );
  NAND2X0 U12965 ( .IN1(n12364), .IN2(n12365), .QN(g22183) );
  NAND2X0 U12966 ( .IN1(n12366), .IN2(n4373), .QN(n12365) );
  OR2X1 U12967 ( .IN1(n12366), .IN2(n7178), .Q(n12364) );
  NAND2X0 U12968 ( .IN1(n12367), .IN2(n12368), .QN(g22182) );
  NAND2X0 U12969 ( .IN1(n12354), .IN2(n4377), .QN(n12368) );
  OR2X1 U12970 ( .IN1(n12354), .IN2(n7179), .Q(n12367) );
  NAND2X0 U12971 ( .IN1(n12369), .IN2(n12370), .QN(g22180) );
  OR2X1 U12972 ( .IN1(n11948), .IN2(n6798), .Q(n12370) );
  NAND2X0 U12973 ( .IN1(n11948), .IN2(n8603), .QN(n12369) );
  NAND2X0 U12974 ( .IN1(n12371), .IN2(n12372), .QN(g22179) );
  NAND2X0 U12975 ( .IN1(n12373), .IN2(n4374), .QN(n12372) );
  OR2X1 U12976 ( .IN1(n12373), .IN2(n7192), .Q(n12371) );
  NAND2X0 U12977 ( .IN1(n12374), .IN2(n12375), .QN(g22178) );
  NAND2X0 U12978 ( .IN1(n11948), .IN2(n4378), .QN(n12375) );
  OR2X1 U12979 ( .IN1(n11948), .IN2(n6808), .Q(n12374) );
  NAND2X0 U12980 ( .IN1(n12376), .IN2(n12377), .QN(g22177) );
  NAND2X0 U12981 ( .IN1(n11950), .IN2(n4375), .QN(n12377) );
  OR2X1 U12982 ( .IN1(n11950), .IN2(n6821), .Q(n12376) );
  NAND2X0 U12983 ( .IN1(n12378), .IN2(n12379), .QN(g22173) );
  OR2X1 U12984 ( .IN1(n12366), .IN2(n6789), .Q(n12379) );
  NAND2X0 U12985 ( .IN1(n12366), .IN2(n8573), .QN(n12378) );
  INVX0 U12986 ( .INP(n9813), .ZN(n8573) );
  NAND3X0 U12987 ( .IN1(n12380), .IN2(n12381), .IN3(n12382), .QN(n9813) );
  NAND2X0 U12988 ( .IN1(n6855), .IN2(test_so73), .QN(n12382) );
  NAND2X0 U12989 ( .IN1(n6856), .IN2(g6837), .QN(n12381) );
  NAND2X0 U12990 ( .IN1(n6854), .IN2(g2241), .QN(n12380) );
  NAND2X0 U12991 ( .IN1(n12383), .IN2(n12384), .QN(g22172) );
  OR2X1 U12992 ( .IN1(n12354), .IN2(n6780), .Q(n12384) );
  NAND2X0 U12993 ( .IN1(n9482), .IN2(n12354), .QN(n12383) );
  NAND2X0 U12994 ( .IN1(n12385), .IN2(n12386), .QN(g22171) );
  NAND2X0 U12995 ( .IN1(n11946), .IN2(n4287), .QN(n12386) );
  OR2X1 U12996 ( .IN1(n11946), .IN2(n6790), .Q(n12385) );
  NAND2X0 U12997 ( .IN1(n12387), .IN2(n12388), .QN(g22170) );
  NAND2X0 U12998 ( .IN1(n12366), .IN2(n4377), .QN(n12388) );
  OR2X1 U12999 ( .IN1(n12366), .IN2(n7180), .Q(n12387) );
  NAND2X0 U13000 ( .IN1(n12389), .IN2(n12390), .QN(g22169) );
  OR2X1 U13001 ( .IN1(n12373), .IN2(n6799), .Q(n12390) );
  NAND2X0 U13002 ( .IN1(n12373), .IN2(n8603), .QN(n12389) );
  NAND2X0 U13003 ( .IN1(n12391), .IN2(n12392), .QN(g22168) );
  OR2X1 U13004 ( .IN1(n11948), .IN2(n6782), .Q(n12392) );
  NAND2X0 U13005 ( .IN1(n12393), .IN2(n11948), .QN(n12391) );
  NAND2X0 U13006 ( .IN1(n12394), .IN2(n12395), .QN(g22167) );
  NAND2X0 U13007 ( .IN1(test_so52), .IN2(n12396), .QN(n12395) );
  NAND2X0 U13008 ( .IN1(n12397), .IN2(n4374), .QN(n12394) );
  NAND2X0 U13009 ( .IN1(n12398), .IN2(n12399), .QN(g22166) );
  NAND2X0 U13010 ( .IN1(n12373), .IN2(n4378), .QN(n12399) );
  OR2X1 U13011 ( .IN1(n12373), .IN2(n7193), .Q(n12398) );
  NAND2X0 U13012 ( .IN1(n12400), .IN2(n12401), .QN(g22164) );
  OR2X1 U13013 ( .IN1(n11950), .IN2(n6809), .Q(n12401) );
  NAND2X0 U13014 ( .IN1(n11950), .IN2(n8634), .QN(n12400) );
  NAND2X0 U13015 ( .IN1(n12402), .IN2(n12403), .QN(g22163) );
  NAND2X0 U13016 ( .IN1(n12404), .IN2(n4375), .QN(n12403) );
  OR2X1 U13017 ( .IN1(n12404), .IN2(n7206), .Q(n12402) );
  NAND2X0 U13018 ( .IN1(n12405), .IN2(n12406), .QN(g22162) );
  NAND2X0 U13019 ( .IN1(n4379), .IN2(n11950), .QN(n12406) );
  OR2X1 U13020 ( .IN1(n11950), .IN2(n6822), .Q(n12405) );
  NAND2X0 U13021 ( .IN1(n12407), .IN2(n12408), .QN(g22161) );
  NAND2X0 U13022 ( .IN1(n11952), .IN2(n4376), .QN(n12408) );
  OR2X1 U13023 ( .IN1(n11952), .IN2(n6830), .Q(n12407) );
  NAND2X0 U13024 ( .IN1(n12409), .IN2(n12410), .QN(g22155) );
  OR2X1 U13025 ( .IN1(n12366), .IN2(n6781), .Q(n12410) );
  NAND2X0 U13026 ( .IN1(n12366), .IN2(n9482), .QN(n12409) );
  INVX0 U13027 ( .INP(n8719), .ZN(n9482) );
  NAND3X0 U13028 ( .IN1(n12411), .IN2(n12412), .IN3(n12413), .QN(n8719) );
  NAND2X0 U13029 ( .IN1(n6852), .IN2(test_so73), .QN(n12413) );
  NAND2X0 U13030 ( .IN1(n6853), .IN2(g6837), .QN(n12412) );
  NAND2X0 U13031 ( .IN1(n6851), .IN2(g2241), .QN(n12411) );
  NAND2X0 U13032 ( .IN1(n12414), .IN2(n12415), .QN(g22154) );
  NAND2X0 U13033 ( .IN1(n12354), .IN2(n4287), .QN(n12415) );
  OR2X1 U13034 ( .IN1(n12354), .IN2(n7166), .Q(n12414) );
  NAND2X0 U13035 ( .IN1(n12416), .IN2(n12417), .QN(g22153) );
  NAND2X0 U13036 ( .IN1(n11946), .IN2(n4563), .QN(n12417) );
  OR2X1 U13037 ( .IN1(n11946), .IN2(n6791), .Q(n12416) );
  NAND2X0 U13038 ( .IN1(n12418), .IN2(n12419), .QN(g22152) );
  OR2X1 U13039 ( .IN1(n12397), .IN2(n6800), .Q(n12419) );
  NAND2X0 U13040 ( .IN1(n12397), .IN2(n8603), .QN(n12418) );
  INVX0 U13041 ( .INP(n9851), .ZN(n8603) );
  NAND3X0 U13042 ( .IN1(n12420), .IN2(n12421), .IN3(n12422), .QN(n9851) );
  NAND2X0 U13043 ( .IN1(n6866), .IN2(g6782), .QN(n12422) );
  NAND2X0 U13044 ( .IN1(n6867), .IN2(g6573), .QN(n12421) );
  OR2X1 U13045 ( .IN1(n4368), .IN2(test_so54), .Q(n12420) );
  NAND2X0 U13046 ( .IN1(n12423), .IN2(n12424), .QN(g22151) );
  OR2X1 U13047 ( .IN1(n12373), .IN2(n6783), .Q(n12424) );
  NAND2X0 U13048 ( .IN1(n12393), .IN2(n12373), .QN(n12423) );
  NAND2X0 U13049 ( .IN1(n12425), .IN2(n12426), .QN(g22150) );
  NAND2X0 U13050 ( .IN1(n11948), .IN2(n4288), .QN(n12426) );
  OR2X1 U13051 ( .IN1(n11948), .IN2(n6801), .Q(n12425) );
  NAND2X0 U13052 ( .IN1(n12427), .IN2(n12428), .QN(g22149) );
  NAND2X0 U13053 ( .IN1(n12397), .IN2(n4378), .QN(n12428) );
  OR2X1 U13054 ( .IN1(n12397), .IN2(n7194), .Q(n12427) );
  NAND2X0 U13055 ( .IN1(n12429), .IN2(n12430), .QN(g22148) );
  OR2X1 U13056 ( .IN1(n12404), .IN2(n6810), .Q(n12430) );
  NAND2X0 U13057 ( .IN1(n12404), .IN2(n8634), .QN(n12429) );
  NAND2X0 U13058 ( .IN1(n12431), .IN2(n12432), .QN(g22147) );
  OR2X1 U13059 ( .IN1(n11950), .IN2(n6812), .Q(n12432) );
  NAND2X0 U13060 ( .IN1(n9651), .IN2(n11950), .QN(n12431) );
  NAND2X0 U13061 ( .IN1(n12433), .IN2(n12434), .QN(g22146) );
  NAND2X0 U13062 ( .IN1(n12435), .IN2(n4375), .QN(n12434) );
  OR2X1 U13063 ( .IN1(n12435), .IN2(n7207), .Q(n12433) );
  NAND2X0 U13064 ( .IN1(n12436), .IN2(n12437), .QN(g22145) );
  NAND2X0 U13065 ( .IN1(n12404), .IN2(n4379), .QN(n12437) );
  OR2X1 U13066 ( .IN1(n12404), .IN2(n7208), .Q(n12436) );
  NAND2X0 U13067 ( .IN1(n12438), .IN2(n12439), .QN(g22143) );
  OR2X1 U13068 ( .IN1(n11952), .IN2(n6823), .Q(n12439) );
  NAND2X0 U13069 ( .IN1(n11952), .IN2(n8680), .QN(n12438) );
  NAND2X0 U13070 ( .IN1(n12440), .IN2(n12441), .QN(g22142) );
  NAND2X0 U13071 ( .IN1(n12442), .IN2(n4376), .QN(n12441) );
  OR2X1 U13072 ( .IN1(n12442), .IN2(n7222), .Q(n12440) );
  NAND2X0 U13073 ( .IN1(n12443), .IN2(n12444), .QN(g22141) );
  NAND2X0 U13074 ( .IN1(n4380), .IN2(n11952), .QN(n12444) );
  OR2X1 U13075 ( .IN1(n11952), .IN2(n6831), .Q(n12443) );
  NAND2X0 U13076 ( .IN1(n12445), .IN2(n12446), .QN(g22140) );
  NAND2X0 U13077 ( .IN1(n12366), .IN2(n4287), .QN(n12446) );
  OR2X1 U13078 ( .IN1(n12366), .IN2(n7167), .Q(n12445) );
  NAND2X0 U13079 ( .IN1(n12447), .IN2(n12448), .QN(g22139) );
  NAND2X0 U13080 ( .IN1(n12354), .IN2(n4563), .QN(n12448) );
  OR2X1 U13081 ( .IN1(n12354), .IN2(n7168), .Q(n12447) );
  NAND2X0 U13082 ( .IN1(n12449), .IN2(n12450), .QN(g22138) );
  NAND2X0 U13083 ( .IN1(n11946), .IN2(n4555), .QN(n12450) );
  OR2X1 U13084 ( .IN1(n11946), .IN2(n6792), .Q(n12449) );
  NAND2X0 U13085 ( .IN1(n12451), .IN2(n12452), .QN(g22132) );
  OR2X1 U13086 ( .IN1(n12397), .IN2(n6784), .Q(n12452) );
  NAND2X0 U13087 ( .IN1(n12397), .IN2(n12393), .QN(n12451) );
  INVX0 U13088 ( .INP(n8756), .ZN(n12393) );
  NAND3X0 U13089 ( .IN1(n12453), .IN2(n12454), .IN3(n12455), .QN(n8756) );
  NAND2X0 U13090 ( .IN1(n6864), .IN2(g6782), .QN(n12455) );
  NAND2X0 U13091 ( .IN1(n6865), .IN2(g6573), .QN(n12454) );
  NAND2X0 U13092 ( .IN1(n6863), .IN2(g1547), .QN(n12453) );
  NAND2X0 U13093 ( .IN1(n12456), .IN2(n12457), .QN(g22131) );
  NAND2X0 U13094 ( .IN1(n12373), .IN2(n4288), .QN(n12457) );
  OR2X1 U13095 ( .IN1(n12373), .IN2(n7181), .Q(n12456) );
  NAND2X0 U13096 ( .IN1(n12458), .IN2(n12459), .QN(g22130) );
  NAND2X0 U13097 ( .IN1(n11948), .IN2(n4565), .QN(n12459) );
  OR2X1 U13098 ( .IN1(n11948), .IN2(n6802), .Q(n12458) );
  NAND2X0 U13099 ( .IN1(n12460), .IN2(n12461), .QN(g22129) );
  OR2X1 U13100 ( .IN1(n12435), .IN2(n6811), .Q(n12461) );
  NAND2X0 U13101 ( .IN1(n12435), .IN2(n8634), .QN(n12460) );
  INVX0 U13102 ( .INP(n9883), .ZN(n8634) );
  NAND3X0 U13103 ( .IN1(n12462), .IN2(n12463), .IN3(n12464), .QN(n9883) );
  NAND2X0 U13104 ( .IN1(n6877), .IN2(test_so31), .QN(n12464) );
  NAND2X0 U13105 ( .IN1(n6878), .IN2(g6518), .QN(n12463) );
  NAND2X0 U13106 ( .IN1(n6879), .IN2(g6368), .QN(n12462) );
  NAND2X0 U13107 ( .IN1(n12465), .IN2(n12466), .QN(g22128) );
  OR2X1 U13108 ( .IN1(n12404), .IN2(n6813), .Q(n12466) );
  NAND2X0 U13109 ( .IN1(n9651), .IN2(n12404), .QN(n12465) );
  NAND2X0 U13110 ( .IN1(n12467), .IN2(n12468), .QN(g22127) );
  NAND2X0 U13111 ( .IN1(n4289), .IN2(n11950), .QN(n12468) );
  OR2X1 U13112 ( .IN1(n11950), .IN2(n6815), .Q(n12467) );
  NAND2X0 U13113 ( .IN1(n12469), .IN2(n12470), .QN(g22126) );
  NAND2X0 U13114 ( .IN1(n12435), .IN2(n4379), .QN(n12470) );
  OR2X1 U13115 ( .IN1(n12435), .IN2(n7209), .Q(n12469) );
  NAND2X0 U13116 ( .IN1(n12471), .IN2(n12472), .QN(g22125) );
  OR2X1 U13117 ( .IN1(n12442), .IN2(n6824), .Q(n12472) );
  NAND2X0 U13118 ( .IN1(n12442), .IN2(n8680), .QN(n12471) );
  NAND2X0 U13119 ( .IN1(n12473), .IN2(n12474), .QN(g22124) );
  OR2X1 U13120 ( .IN1(n11952), .IN2(n6785), .Q(n12474) );
  NAND2X0 U13121 ( .IN1(n11311), .IN2(n11952), .QN(n12473) );
  NAND2X0 U13122 ( .IN1(n12475), .IN2(n12476), .QN(g22123) );
  NAND2X0 U13123 ( .IN1(n12477), .IN2(n4376), .QN(n12476) );
  OR2X1 U13124 ( .IN1(n12477), .IN2(n7223), .Q(n12475) );
  NAND2X0 U13125 ( .IN1(n12478), .IN2(n12479), .QN(g22122) );
  NAND2X0 U13126 ( .IN1(n12442), .IN2(n4380), .QN(n12479) );
  OR2X1 U13127 ( .IN1(n12442), .IN2(n7224), .Q(n12478) );
  NAND2X0 U13128 ( .IN1(n12480), .IN2(n12481), .QN(g22117) );
  NAND2X0 U13129 ( .IN1(n12366), .IN2(n4563), .QN(n12481) );
  OR2X1 U13130 ( .IN1(n12366), .IN2(n7169), .Q(n12480) );
  NAND2X0 U13131 ( .IN1(n12482), .IN2(n12483), .QN(g22116) );
  NAND2X0 U13132 ( .IN1(n12354), .IN2(n4555), .QN(n12483) );
  OR2X1 U13133 ( .IN1(n12354), .IN2(n7170), .Q(n12482) );
  NAND2X0 U13134 ( .IN1(n12484), .IN2(n12485), .QN(g22115) );
  NAND2X0 U13135 ( .IN1(n11946), .IN2(n4325), .QN(n12485) );
  OR2X1 U13136 ( .IN1(n11946), .IN2(n6793), .Q(n12484) );
  NAND2X0 U13137 ( .IN1(n12486), .IN2(n12487), .QN(g22114) );
  NAND2X0 U13138 ( .IN1(n12397), .IN2(n4288), .QN(n12487) );
  OR2X1 U13139 ( .IN1(n12397), .IN2(n7182), .Q(n12486) );
  NAND2X0 U13140 ( .IN1(n12488), .IN2(n12489), .QN(g22113) );
  NAND2X0 U13141 ( .IN1(test_so53), .IN2(n12490), .QN(n12489) );
  NAND2X0 U13142 ( .IN1(n12373), .IN2(n4565), .QN(n12488) );
  NAND2X0 U13143 ( .IN1(n12491), .IN2(n12492), .QN(g22112) );
  NAND2X0 U13144 ( .IN1(n11948), .IN2(n4557), .QN(n12492) );
  OR2X1 U13145 ( .IN1(n11948), .IN2(n6803), .Q(n12491) );
  NAND2X0 U13146 ( .IN1(n12493), .IN2(n12494), .QN(g22106) );
  OR2X1 U13147 ( .IN1(n12435), .IN2(n6814), .Q(n12494) );
  NAND2X0 U13148 ( .IN1(n12435), .IN2(n9651), .QN(n12493) );
  INVX0 U13149 ( .INP(n8790), .ZN(n9651) );
  NAND3X0 U13150 ( .IN1(n12495), .IN2(n12496), .IN3(n12497), .QN(n8790) );
  NAND2X0 U13151 ( .IN1(n6874), .IN2(test_so31), .QN(n12497) );
  NAND2X0 U13152 ( .IN1(n6875), .IN2(g6518), .QN(n12496) );
  NAND2X0 U13153 ( .IN1(n6876), .IN2(g6368), .QN(n12495) );
  NAND2X0 U13154 ( .IN1(n12498), .IN2(n12499), .QN(g22105) );
  NAND2X0 U13155 ( .IN1(n4289), .IN2(n12404), .QN(n12499) );
  OR2X1 U13156 ( .IN1(n12404), .IN2(n7195), .Q(n12498) );
  NAND2X0 U13157 ( .IN1(n12500), .IN2(n12501), .QN(g22104) );
  NAND2X0 U13158 ( .IN1(n11950), .IN2(n4567), .QN(n12501) );
  OR2X1 U13159 ( .IN1(n11950), .IN2(n6816), .Q(n12500) );
  NAND2X0 U13160 ( .IN1(n12502), .IN2(n12503), .QN(g22103) );
  NAND2X0 U13161 ( .IN1(test_so12), .IN2(n12504), .QN(n12503) );
  NAND2X0 U13162 ( .IN1(n12477), .IN2(n8680), .QN(n12502) );
  INVX0 U13163 ( .INP(n9910), .ZN(n8680) );
  NAND3X0 U13164 ( .IN1(n12505), .IN2(n12506), .IN3(n12507), .QN(n9910) );
  NAND2X0 U13165 ( .IN1(n6889), .IN2(g6313), .QN(n12507) );
  NAND2X0 U13166 ( .IN1(n6890), .IN2(g6231), .QN(n12506) );
  NAND2X0 U13167 ( .IN1(n6888), .IN2(g165), .QN(n12505) );
  NAND2X0 U13168 ( .IN1(n12508), .IN2(n12509), .QN(g22102) );
  OR2X1 U13169 ( .IN1(n12442), .IN2(n6786), .Q(n12509) );
  NAND2X0 U13170 ( .IN1(n11311), .IN2(n12442), .QN(n12508) );
  NAND2X0 U13171 ( .IN1(n12510), .IN2(n12511), .QN(g22101) );
  NAND2X0 U13172 ( .IN1(n4290), .IN2(n11952), .QN(n12511) );
  OR2X1 U13173 ( .IN1(n11952), .IN2(n6825), .Q(n12510) );
  NAND2X0 U13174 ( .IN1(n12512), .IN2(n12513), .QN(g22100) );
  NAND2X0 U13175 ( .IN1(n12477), .IN2(n4380), .QN(n12513) );
  OR2X1 U13176 ( .IN1(n12477), .IN2(n7225), .Q(n12512) );
  NAND2X0 U13177 ( .IN1(n12514), .IN2(n12515), .QN(g22099) );
  NAND2X0 U13178 ( .IN1(n12366), .IN2(n4555), .QN(n12515) );
  OR2X1 U13179 ( .IN1(n12366), .IN2(n7171), .Q(n12514) );
  NAND2X0 U13180 ( .IN1(n12516), .IN2(n12517), .QN(g22098) );
  NAND2X0 U13181 ( .IN1(test_so74), .IN2(n12361), .QN(n12517) );
  NAND2X0 U13182 ( .IN1(n12354), .IN2(n4325), .QN(n12516) );
  NAND2X0 U13183 ( .IN1(n12518), .IN2(n12519), .QN(g22097) );
  NAND2X0 U13184 ( .IN1(n11946), .IN2(n4389), .QN(n12519) );
  OR2X1 U13185 ( .IN1(n11946), .IN2(n6794), .Q(n12518) );
  NAND2X0 U13186 ( .IN1(n12520), .IN2(n12521), .QN(g22092) );
  NAND2X0 U13187 ( .IN1(n12397), .IN2(n4565), .QN(n12521) );
  OR2X1 U13188 ( .IN1(n12397), .IN2(n7183), .Q(n12520) );
  NAND2X0 U13189 ( .IN1(n12522), .IN2(n12523), .QN(g22091) );
  NAND2X0 U13190 ( .IN1(n12373), .IN2(n4557), .QN(n12523) );
  OR2X1 U13191 ( .IN1(n12373), .IN2(n7184), .Q(n12522) );
  NAND2X0 U13192 ( .IN1(n12524), .IN2(n12525), .QN(g22090) );
  NAND2X0 U13193 ( .IN1(n11948), .IN2(n4326), .QN(n12525) );
  OR2X1 U13194 ( .IN1(n11948), .IN2(n6804), .Q(n12524) );
  NAND2X0 U13195 ( .IN1(n12526), .IN2(n12527), .QN(g22089) );
  NAND2X0 U13196 ( .IN1(n4289), .IN2(n12435), .QN(n12527) );
  OR2X1 U13197 ( .IN1(n12435), .IN2(n7196), .Q(n12526) );
  NAND2X0 U13198 ( .IN1(n12528), .IN2(n12529), .QN(g22088) );
  NAND2X0 U13199 ( .IN1(n12404), .IN2(n4567), .QN(n12529) );
  OR2X1 U13200 ( .IN1(n12404), .IN2(n7197), .Q(n12528) );
  NAND2X0 U13201 ( .IN1(n12530), .IN2(n12531), .QN(g22087) );
  NAND2X0 U13202 ( .IN1(n11950), .IN2(n4559), .QN(n12531) );
  OR2X1 U13203 ( .IN1(n11950), .IN2(n6817), .Q(n12530) );
  NAND2X0 U13204 ( .IN1(n12532), .IN2(n12533), .QN(g22081) );
  OR2X1 U13205 ( .IN1(n12477), .IN2(n6787), .Q(n12533) );
  NAND2X0 U13206 ( .IN1(n12477), .IN2(n11311), .QN(n12532) );
  INVX0 U13207 ( .INP(n8810), .ZN(n11311) );
  NAND3X0 U13208 ( .IN1(n12534), .IN2(n12535), .IN3(n12536), .QN(n8810) );
  NAND2X0 U13209 ( .IN1(n6886), .IN2(g6313), .QN(n12536) );
  NAND2X0 U13210 ( .IN1(n6887), .IN2(g6231), .QN(n12535) );
  NAND2X0 U13211 ( .IN1(n6885), .IN2(g165), .QN(n12534) );
  NAND2X0 U13212 ( .IN1(n12537), .IN2(n12538), .QN(g22080) );
  NAND2X0 U13213 ( .IN1(n4290), .IN2(n12442), .QN(n12538) );
  OR2X1 U13214 ( .IN1(n12442), .IN2(n7210), .Q(n12537) );
  NAND2X0 U13215 ( .IN1(n12539), .IN2(n12540), .QN(g22079) );
  NAND2X0 U13216 ( .IN1(n11952), .IN2(n4569), .QN(n12540) );
  OR2X1 U13217 ( .IN1(n11952), .IN2(n6826), .Q(n12539) );
  NAND2X0 U13218 ( .IN1(n12541), .IN2(n12542), .QN(g22078) );
  NAND2X0 U13219 ( .IN1(n12366), .IN2(n4325), .QN(n12542) );
  OR2X1 U13220 ( .IN1(n12366), .IN2(n7172), .Q(n12541) );
  NAND2X0 U13221 ( .IN1(n12543), .IN2(n12544), .QN(g22077) );
  NAND2X0 U13222 ( .IN1(n12354), .IN2(n4389), .QN(n12544) );
  OR2X1 U13223 ( .IN1(n12354), .IN2(n7173), .Q(n12543) );
  NAND2X0 U13224 ( .IN1(n12545), .IN2(n12546), .QN(g22076) );
  NAND2X0 U13225 ( .IN1(n11946), .IN2(n4319), .QN(n12546) );
  OR2X1 U13226 ( .IN1(n11946), .IN2(n6795), .Q(n12545) );
  NOR2X0 U13227 ( .IN1(n4367), .IN2(n6998), .QN(n11946) );
  NAND2X0 U13228 ( .IN1(n12547), .IN2(n12548), .QN(g22075) );
  NAND2X0 U13229 ( .IN1(n12397), .IN2(n4557), .QN(n12548) );
  OR2X1 U13230 ( .IN1(n12397), .IN2(n7185), .Q(n12547) );
  NAND2X0 U13231 ( .IN1(n12549), .IN2(n12550), .QN(g22074) );
  NAND2X0 U13232 ( .IN1(n12373), .IN2(n4326), .QN(n12550) );
  OR2X1 U13233 ( .IN1(n12373), .IN2(n7186), .Q(n12549) );
  NAND2X0 U13234 ( .IN1(n12551), .IN2(n12552), .QN(g22073) );
  NAND2X0 U13235 ( .IN1(n11948), .IN2(n4390), .QN(n12552) );
  OR2X1 U13236 ( .IN1(n11948), .IN2(n6805), .Q(n12551) );
  NAND2X0 U13237 ( .IN1(n12553), .IN2(n12554), .QN(g22068) );
  NAND2X0 U13238 ( .IN1(n12435), .IN2(n4567), .QN(n12554) );
  OR2X1 U13239 ( .IN1(n12435), .IN2(n7198), .Q(n12553) );
  NAND2X0 U13240 ( .IN1(n12555), .IN2(n12556), .QN(g22067) );
  NAND2X0 U13241 ( .IN1(n12404), .IN2(n4559), .QN(n12556) );
  OR2X1 U13242 ( .IN1(n12404), .IN2(n7199), .Q(n12555) );
  NAND2X0 U13243 ( .IN1(n12557), .IN2(n12558), .QN(g22066) );
  NAND2X0 U13244 ( .IN1(n4327), .IN2(n11950), .QN(n12558) );
  OR2X1 U13245 ( .IN1(n11950), .IN2(n6818), .Q(n12557) );
  NAND2X0 U13246 ( .IN1(n12559), .IN2(n12560), .QN(g22065) );
  NAND2X0 U13247 ( .IN1(n4290), .IN2(n12477), .QN(n12560) );
  OR2X1 U13248 ( .IN1(n12477), .IN2(n7211), .Q(n12559) );
  NAND2X0 U13249 ( .IN1(n12561), .IN2(n12562), .QN(g22064) );
  NAND2X0 U13250 ( .IN1(n12442), .IN2(n4569), .QN(n12562) );
  OR2X1 U13251 ( .IN1(n12442), .IN2(n7212), .Q(n12561) );
  NAND2X0 U13252 ( .IN1(n12563), .IN2(n12564), .QN(g22063) );
  NAND2X0 U13253 ( .IN1(n11952), .IN2(n4561), .QN(n12564) );
  OR2X1 U13254 ( .IN1(n11952), .IN2(n6827), .Q(n12563) );
  NAND2X0 U13255 ( .IN1(n12565), .IN2(n12566), .QN(g22061) );
  NAND2X0 U13256 ( .IN1(n12366), .IN2(n4389), .QN(n12566) );
  OR2X1 U13257 ( .IN1(n12366), .IN2(n7174), .Q(n12565) );
  NAND2X0 U13258 ( .IN1(n12567), .IN2(n12568), .QN(g22060) );
  NAND2X0 U13259 ( .IN1(n12354), .IN2(n4319), .QN(n12568) );
  OR2X1 U13260 ( .IN1(n12354), .IN2(n7175), .Q(n12567) );
  INVX0 U13261 ( .INP(n12361), .ZN(n12354) );
  NAND2X0 U13262 ( .IN1(test_so73), .IN2(g2257), .QN(n12361) );
  NAND2X0 U13263 ( .IN1(n12569), .IN2(n12570), .QN(g22059) );
  NAND2X0 U13264 ( .IN1(n12397), .IN2(n4326), .QN(n12570) );
  OR2X1 U13265 ( .IN1(n12397), .IN2(n7187), .Q(n12569) );
  NAND2X0 U13266 ( .IN1(n12571), .IN2(n12572), .QN(g22058) );
  NAND2X0 U13267 ( .IN1(n12373), .IN2(n4390), .QN(n12572) );
  OR2X1 U13268 ( .IN1(n12373), .IN2(n7188), .Q(n12571) );
  NAND2X0 U13269 ( .IN1(n12573), .IN2(n12574), .QN(g22057) );
  NAND2X0 U13270 ( .IN1(n11948), .IN2(n4320), .QN(n12574) );
  OR2X1 U13271 ( .IN1(n11948), .IN2(n6806), .Q(n12573) );
  NOR2X0 U13272 ( .IN1(n4368), .IN2(n6999), .QN(n11948) );
  NAND2X0 U13273 ( .IN1(n12575), .IN2(n12576), .QN(g22056) );
  NAND2X0 U13274 ( .IN1(test_so32), .IN2(n12577), .QN(n12576) );
  NAND2X0 U13275 ( .IN1(n12435), .IN2(n4559), .QN(n12575) );
  NAND2X0 U13276 ( .IN1(n12578), .IN2(n12579), .QN(g22055) );
  NAND2X0 U13277 ( .IN1(n4327), .IN2(n12404), .QN(n12579) );
  OR2X1 U13278 ( .IN1(n12404), .IN2(n7200), .Q(n12578) );
  NAND2X0 U13279 ( .IN1(n12580), .IN2(n12581), .QN(g22054) );
  NAND2X0 U13280 ( .IN1(n11950), .IN2(n4391), .QN(n12581) );
  OR2X1 U13281 ( .IN1(n11950), .IN2(n6819), .Q(n12580) );
  NAND2X0 U13282 ( .IN1(n12582), .IN2(n12583), .QN(g22049) );
  NAND2X0 U13283 ( .IN1(n12477), .IN2(n4569), .QN(n12583) );
  OR2X1 U13284 ( .IN1(n12477), .IN2(n7213), .Q(n12582) );
  NAND2X0 U13285 ( .IN1(n12584), .IN2(n12585), .QN(g22048) );
  NAND2X0 U13286 ( .IN1(n12442), .IN2(n4561), .QN(n12585) );
  OR2X1 U13287 ( .IN1(n12442), .IN2(n7214), .Q(n12584) );
  NAND2X0 U13288 ( .IN1(n12586), .IN2(n12587), .QN(g22047) );
  NAND2X0 U13289 ( .IN1(n4328), .IN2(n11952), .QN(n12587) );
  OR2X1 U13290 ( .IN1(n11952), .IN2(n6828), .Q(n12586) );
  NAND2X0 U13291 ( .IN1(n12588), .IN2(n12589), .QN(g22045) );
  NAND2X0 U13292 ( .IN1(n12366), .IN2(n4319), .QN(n12589) );
  OR2X1 U13293 ( .IN1(n12366), .IN2(n7176), .Q(n12588) );
  NOR2X0 U13294 ( .IN1(n4324), .IN2(n6998), .QN(n12366) );
  NAND2X0 U13295 ( .IN1(n12590), .IN2(n12591), .QN(g22044) );
  NAND2X0 U13296 ( .IN1(n12397), .IN2(n4390), .QN(n12591) );
  OR2X1 U13297 ( .IN1(n12397), .IN2(n7189), .Q(n12590) );
  NAND2X0 U13298 ( .IN1(n12592), .IN2(n12593), .QN(g22043) );
  NAND2X0 U13299 ( .IN1(n12373), .IN2(n4320), .QN(n12593) );
  OR2X1 U13300 ( .IN1(n12373), .IN2(n7190), .Q(n12592) );
  INVX0 U13301 ( .INP(n12490), .ZN(n12373) );
  NAND2X0 U13302 ( .IN1(g6782), .IN2(g1563), .QN(n12490) );
  NAND2X0 U13303 ( .IN1(n12594), .IN2(n12595), .QN(g22042) );
  NAND2X0 U13304 ( .IN1(n4327), .IN2(n12435), .QN(n12595) );
  OR2X1 U13305 ( .IN1(n12435), .IN2(n7201), .Q(n12594) );
  NAND2X0 U13306 ( .IN1(n12596), .IN2(n12597), .QN(g22041) );
  NAND2X0 U13307 ( .IN1(n12404), .IN2(n4391), .QN(n12597) );
  OR2X1 U13308 ( .IN1(n12404), .IN2(n7202), .Q(n12596) );
  NAND2X0 U13309 ( .IN1(n12598), .IN2(n12599), .QN(g22040) );
  NAND2X0 U13310 ( .IN1(n4321), .IN2(n11950), .QN(n12599) );
  OR2X1 U13311 ( .IN1(n11950), .IN2(n6820), .Q(n12598) );
  NOR2X0 U13312 ( .IN1(n7267), .IN2(n7000), .QN(n11950) );
  NAND2X0 U13313 ( .IN1(n12600), .IN2(n12601), .QN(g22039) );
  NAND2X0 U13314 ( .IN1(n12477), .IN2(n4561), .QN(n12601) );
  OR2X1 U13315 ( .IN1(n12477), .IN2(n7215), .Q(n12600) );
  NAND2X0 U13316 ( .IN1(n12602), .IN2(n12603), .QN(g22038) );
  NAND2X0 U13317 ( .IN1(n4328), .IN2(n12442), .QN(n12603) );
  OR2X1 U13318 ( .IN1(n12442), .IN2(n7216), .Q(n12602) );
  NAND2X0 U13319 ( .IN1(n12604), .IN2(n12605), .QN(g22037) );
  NAND2X0 U13320 ( .IN1(test_so11), .IN2(n12606), .QN(n12605) );
  NAND2X0 U13321 ( .IN1(n11952), .IN2(n4392), .QN(n12604) );
  NAND2X0 U13322 ( .IN1(n12607), .IN2(n12608), .QN(g22035) );
  NAND2X0 U13323 ( .IN1(n12397), .IN2(n4320), .QN(n12608) );
  OR2X1 U13324 ( .IN1(n12397), .IN2(n7191), .Q(n12607) );
  INVX0 U13325 ( .INP(n12396), .ZN(n12397) );
  NAND2X0 U13326 ( .IN1(g6573), .IN2(g1563), .QN(n12396) );
  NAND2X0 U13327 ( .IN1(n12609), .IN2(n12610), .QN(g22034) );
  NAND2X0 U13328 ( .IN1(n12435), .IN2(n4391), .QN(n12610) );
  OR2X1 U13329 ( .IN1(n12435), .IN2(n7203), .Q(n12609) );
  NAND2X0 U13330 ( .IN1(n12611), .IN2(n12612), .QN(g22033) );
  NAND2X0 U13331 ( .IN1(n4321), .IN2(n12404), .QN(n12612) );
  OR2X1 U13332 ( .IN1(n12404), .IN2(n7204), .Q(n12611) );
  NOR2X0 U13333 ( .IN1(n4312), .IN2(n7000), .QN(n12404) );
  NAND2X0 U13334 ( .IN1(n12613), .IN2(n12614), .QN(g22032) );
  NAND2X0 U13335 ( .IN1(n4328), .IN2(n12477), .QN(n12614) );
  OR2X1 U13336 ( .IN1(n12477), .IN2(n7217), .Q(n12613) );
  NAND2X0 U13337 ( .IN1(n12615), .IN2(n12616), .QN(g22031) );
  NAND2X0 U13338 ( .IN1(n12442), .IN2(n4392), .QN(n12616) );
  OR2X1 U13339 ( .IN1(n12442), .IN2(n7218), .Q(n12615) );
  NAND2X0 U13340 ( .IN1(n12617), .IN2(n12618), .QN(g22030) );
  NAND2X0 U13341 ( .IN1(n4322), .IN2(n11952), .QN(n12618) );
  OR2X1 U13342 ( .IN1(n11952), .IN2(n6829), .Q(n12617) );
  INVX0 U13343 ( .INP(n12606), .ZN(n11952) );
  NAND2X0 U13344 ( .IN1(g165), .IN2(g181), .QN(n12606) );
  NAND2X0 U13345 ( .IN1(n12619), .IN2(n12620), .QN(g22029) );
  NAND2X0 U13346 ( .IN1(n4321), .IN2(n12435), .QN(n12620) );
  OR2X1 U13347 ( .IN1(n12435), .IN2(n7205), .Q(n12619) );
  INVX0 U13348 ( .INP(n12577), .ZN(n12435) );
  NAND2X0 U13349 ( .IN1(g6368), .IN2(g869), .QN(n12577) );
  NAND2X0 U13350 ( .IN1(n12621), .IN2(n12622), .QN(g22028) );
  NAND2X0 U13351 ( .IN1(n12477), .IN2(n4392), .QN(n12622) );
  OR2X1 U13352 ( .IN1(n12477), .IN2(n7219), .Q(n12621) );
  NAND2X0 U13353 ( .IN1(n12623), .IN2(n12624), .QN(g22027) );
  NAND2X0 U13354 ( .IN1(n4322), .IN2(n12442), .QN(n12624) );
  OR2X1 U13355 ( .IN1(n12442), .IN2(n7220), .Q(n12623) );
  NOR2X0 U13356 ( .IN1(n4512), .IN2(n7001), .QN(n12442) );
  NOR2X0 U13357 ( .IN1(n7777), .IN2(n12625), .QN(g22026) );
  XNOR2X1 U13358 ( .IN1(n7049), .IN2(n12209), .Q(n12625) );
  OR2X1 U13359 ( .IN1(n4423), .IN2(n4330), .Q(n12209) );
  NAND2X0 U13360 ( .IN1(n13231), .IN2(n7782), .QN(n7777) );
  NAND4X0 U13361 ( .IN1(n4182), .IN2(n4431), .IN3(n4330), .IN4(n12626), .QN(
        n7782) );
  NOR4X0 U13362 ( .IN1(n7049), .IN2(n4423), .IN3(n4355), .IN4(g2900), .QN(
        n12626) );
  NAND2X0 U13363 ( .IN1(n12627), .IN2(n12628), .QN(g22025) );
  NAND2X0 U13364 ( .IN1(n4322), .IN2(n12477), .QN(n12628) );
  OR2X1 U13365 ( .IN1(n12477), .IN2(n7221), .Q(n12627) );
  INVX0 U13366 ( .INP(n12504), .ZN(n12477) );
  NAND2X0 U13367 ( .IN1(g6231), .IN2(g181), .QN(n12504) );
  NOR3X0 U13368 ( .IN1(n12629), .IN2(n10335), .IN3(n12073), .QN(g21974) );
  INVX0 U13369 ( .INP(n12075), .ZN(n12073) );
  NAND3X0 U13370 ( .IN1(g2714), .IN2(g2707), .IN3(n12630), .QN(n12075) );
  NOR2X0 U13371 ( .IN1(n12631), .IN2(g2707), .QN(n12629) );
  AND2X1 U13372 ( .IN1(g2714), .IN2(n12630), .Q(n12631) );
  AND3X1 U13373 ( .IN1(n12077), .IN2(n12632), .IN3(n12633), .Q(g21972) );
  NAND2X0 U13374 ( .IN1(n4474), .IN2(n12634), .QN(n12633) );
  NAND2X0 U13375 ( .IN1(n12635), .IN2(g2020), .QN(n12634) );
  NAND3X0 U13376 ( .IN1(g2020), .IN2(g2013), .IN3(n12635), .QN(n12077) );
  NAND2X0 U13377 ( .IN1(n12636), .IN2(n12637), .QN(g21970) );
  NAND2X0 U13378 ( .IN1(test_so87), .IN2(n4463), .QN(n12637) );
  NAND2X0 U13379 ( .IN1(n10381), .IN2(g2560), .QN(n12636) );
  NAND3X0 U13380 ( .IN1(n12638), .IN2(n12639), .IN3(n12640), .QN(n10381) );
  NAND2X0 U13381 ( .IN1(g5555), .IN2(g2513), .QN(n12640) );
  NAND2X0 U13382 ( .IN1(n4606), .IN2(g2519), .QN(n12639) );
  NAND2X0 U13383 ( .IN1(g7264), .IN2(g2516), .QN(n12638) );
  AND3X1 U13384 ( .IN1(n12080), .IN2(n11202), .IN3(n12641), .Q(g21969) );
  NAND2X0 U13385 ( .IN1(n4476), .IN2(n12642), .QN(n12641) );
  OR2X1 U13386 ( .IN1(n12643), .IN2(n4402), .Q(n12642) );
  INVX0 U13387 ( .INP(n10343), .ZN(n11202) );
  OR3X1 U13388 ( .IN1(n4402), .IN2(n4476), .IN3(n12643), .Q(n12080) );
  NAND2X0 U13389 ( .IN1(n12644), .IN2(n12645), .QN(g21882) );
  NAND2X0 U13390 ( .IN1(n4351), .IN2(g2878), .QN(n12645) );
  NAND2X0 U13391 ( .IN1(n12646), .IN2(g2879), .QN(n12644) );
  NAND2X0 U13392 ( .IN1(n12647), .IN2(n12648), .QN(g21880) );
  NAND2X0 U13393 ( .IN1(n4351), .IN2(g2877), .QN(n12648) );
  NAND2X0 U13394 ( .IN1(n12649), .IN2(g2879), .QN(n12647) );
  NAND2X0 U13395 ( .IN1(n12650), .IN2(n12651), .QN(g21878) );
  NAND2X0 U13396 ( .IN1(test_so4), .IN2(g2879), .QN(n12651) );
  NAND2X0 U13397 ( .IN1(n12646), .IN2(n4351), .QN(n12650) );
  XNOR2X1 U13398 ( .IN1(n7656), .IN2(n12652), .Q(n12646) );
  XOR3X1 U13399 ( .IN1(n12653), .IN2(n12654), .IN3(n12655), .Q(n7656) );
  XOR3X1 U13400 ( .IN1(n7254), .IN2(n7253), .IN3(n12656), .Q(n12655) );
  XOR2X1 U13401 ( .IN1(g2981), .IN2(test_so2), .Q(n12656) );
  XOR2X1 U13402 ( .IN1(n7250), .IN2(n7249), .Q(n12654) );
  XOR2X1 U13403 ( .IN1(n7252), .IN2(n7251), .Q(n12653) );
  NAND2X0 U13404 ( .IN1(n12657), .IN2(n12658), .QN(g21851) );
  NAND2X0 U13405 ( .IN1(g499), .IN2(g544), .QN(n12658) );
  NAND3X0 U13406 ( .IN1(n4298), .IN2(g548), .IN3(n4541), .QN(n12657) );
  NAND2X0 U13407 ( .IN1(n11961), .IN2(n12659), .QN(g21847) );
  OR2X1 U13408 ( .IN1(g2624), .IN2(n7233), .Q(n12659) );
  NAND2X0 U13409 ( .IN1(n9947), .IN2(g2624), .QN(n11961) );
  NAND2X0 U13410 ( .IN1(n11980), .IN2(n12660), .QN(g21845) );
  OR2X1 U13411 ( .IN1(g1930), .IN2(n7234), .Q(n12660) );
  NAND2X0 U13412 ( .IN1(n9947), .IN2(g1930), .QN(n11980) );
  NAND2X0 U13413 ( .IN1(n12008), .IN2(n12661), .QN(g21843) );
  OR2X1 U13414 ( .IN1(g1236), .IN2(n7235), .Q(n12661) );
  NAND2X0 U13415 ( .IN1(n9947), .IN2(g1236), .QN(n12008) );
  NAND2X0 U13416 ( .IN1(n12036), .IN2(n12662), .QN(g21842) );
  OR2X1 U13417 ( .IN1(g550), .IN2(n7236), .Q(n12662) );
  NAND2X0 U13418 ( .IN1(n9947), .IN2(g550), .QN(n12036) );
  NAND4X0 U13419 ( .IN1(n6706), .IN2(n12663), .IN3(n12664), .IN4(n4480), .QN(
        n9947) );
  NOR2X0 U13420 ( .IN1(n4481), .IN2(n4350), .QN(n12664) );
  INVX0 U13421 ( .INP(n12216), .ZN(n12663) );
  NAND4X0 U13422 ( .IN1(n6428), .IN2(g3013), .IN3(n6432), .IN4(n12665), .QN(
        n12216) );
  NOR4X0 U13423 ( .IN1(test_so98), .IN2(n13235), .IN3(n6430), .IN4(n6429), 
        .QN(n12665) );
  NAND2X0 U13424 ( .IN1(n12666), .IN2(n12667), .QN(g21346) );
  NAND2X0 U13425 ( .IN1(n13234), .IN2(DFF_328_n1), .QN(n12667) );
  OR3X1 U13426 ( .IN1(g6447), .IN2(n6710), .IN3(n13234), .Q(n12666) );
  NAND2X0 U13427 ( .IN1(n12668), .IN2(n12669), .QN(g21094) );
  NAND2X0 U13428 ( .IN1(test_so94), .IN2(n12670), .QN(n12669) );
  NAND2X0 U13429 ( .IN1(n4393), .IN2(n11563), .QN(n12668) );
  NAND2X0 U13430 ( .IN1(n12671), .IN2(n12672), .QN(g21082) );
  NAND2X0 U13431 ( .IN1(n4393), .IN2(n11566), .QN(n12672) );
  OR2X1 U13432 ( .IN1(n11566), .IN2(n7052), .Q(n12671) );
  NAND2X0 U13433 ( .IN1(n12673), .IN2(n12674), .QN(g21081) );
  NAND2X0 U13434 ( .IN1(n11563), .IN2(n4471), .QN(n12674) );
  OR2X1 U13435 ( .IN1(n11563), .IN2(n7125), .Q(n12673) );
  NAND2X0 U13436 ( .IN1(n12675), .IN2(n12676), .QN(g21080) );
  NAND2X0 U13437 ( .IN1(n11570), .IN2(n7272), .QN(n12676) );
  OR2X1 U13438 ( .IN1(n11570), .IN2(n7133), .Q(n12675) );
  NAND2X0 U13439 ( .IN1(n12677), .IN2(n12678), .QN(g21075) );
  NAND2X0 U13440 ( .IN1(n4393), .IN2(n11573), .QN(n12678) );
  OR2X1 U13441 ( .IN1(n11573), .IN2(n7053), .Q(n12677) );
  NAND2X0 U13442 ( .IN1(n12679), .IN2(n12680), .QN(g21074) );
  NAND2X0 U13443 ( .IN1(n11566), .IN2(n4471), .QN(n12680) );
  OR2X1 U13444 ( .IN1(n11566), .IN2(n7054), .Q(n12679) );
  NAND2X0 U13445 ( .IN1(n12681), .IN2(n12682), .QN(g21073) );
  NAND2X0 U13446 ( .IN1(n11563), .IN2(n7269), .QN(n12682) );
  OR2X1 U13447 ( .IN1(n11563), .IN2(n7126), .Q(n12681) );
  NAND2X0 U13448 ( .IN1(n12683), .IN2(n12684), .QN(g21072) );
  NAND2X0 U13449 ( .IN1(n11628), .IN2(n7272), .QN(n12684) );
  OR2X1 U13450 ( .IN1(n11628), .IN2(n7071), .Q(n12683) );
  NAND2X0 U13451 ( .IN1(n12685), .IN2(n12686), .QN(g21071) );
  NAND2X0 U13452 ( .IN1(n11570), .IN2(n4473), .QN(n12686) );
  OR2X1 U13453 ( .IN1(n11570), .IN2(n7134), .Q(n12685) );
  NAND2X0 U13454 ( .IN1(n12687), .IN2(n12688), .QN(g21070) );
  NAND2X0 U13455 ( .IN1(n4395), .IN2(n11632), .QN(n12688) );
  OR2X1 U13456 ( .IN1(n11632), .IN2(n7143), .Q(n12687) );
  NAND2X0 U13457 ( .IN1(n12689), .IN2(n12690), .QN(g21063) );
  OR2X1 U13458 ( .IN1(n12318), .IN2(n6895), .Q(n12690) );
  NAND2X0 U13459 ( .IN1(n12318), .IN2(n12691), .QN(n12689) );
  NAND2X0 U13460 ( .IN1(n12692), .IN2(n12693), .QN(g21062) );
  NAND2X0 U13461 ( .IN1(n11573), .IN2(n4471), .QN(n12693) );
  OR2X1 U13462 ( .IN1(n11573), .IN2(n7055), .Q(n12692) );
  NAND2X0 U13463 ( .IN1(n12694), .IN2(n12695), .QN(g21061) );
  NAND2X0 U13464 ( .IN1(n11566), .IN2(n7269), .QN(n12695) );
  OR2X1 U13465 ( .IN1(n11566), .IN2(n7056), .Q(n12694) );
  NAND2X0 U13466 ( .IN1(n12696), .IN2(n12697), .QN(g21060) );
  NAND2X0 U13467 ( .IN1(n11563), .IN2(n4407), .QN(n12697) );
  OR2X1 U13468 ( .IN1(n11563), .IN2(n7127), .Q(n12696) );
  NAND2X0 U13469 ( .IN1(n12698), .IN2(n12699), .QN(g21056) );
  NAND2X0 U13470 ( .IN1(n11635), .IN2(n7272), .QN(n12699) );
  OR2X1 U13471 ( .IN1(n11635), .IN2(n7072), .Q(n12698) );
  NAND2X0 U13472 ( .IN1(n12700), .IN2(n12701), .QN(g21055) );
  NAND2X0 U13473 ( .IN1(n11628), .IN2(n4473), .QN(n12701) );
  OR2X1 U13474 ( .IN1(n11628), .IN2(n7073), .Q(n12700) );
  NAND2X0 U13475 ( .IN1(n12702), .IN2(n12703), .QN(g21054) );
  NAND2X0 U13476 ( .IN1(n4468), .IN2(n11570), .QN(n12703) );
  OR2X1 U13477 ( .IN1(n11570), .IN2(n7135), .Q(n12702) );
  NAND2X0 U13478 ( .IN1(n12704), .IN2(n12705), .QN(g21053) );
  NAND2X0 U13479 ( .IN1(n4395), .IN2(n11690), .QN(n12705) );
  OR2X1 U13480 ( .IN1(n11690), .IN2(n7090), .Q(n12704) );
  NAND2X0 U13481 ( .IN1(n12706), .IN2(n12707), .QN(g21052) );
  NAND2X0 U13482 ( .IN1(n11632), .IN2(n4475), .QN(n12707) );
  OR2X1 U13483 ( .IN1(n11632), .IN2(n7144), .Q(n12706) );
  NAND2X0 U13484 ( .IN1(n12708), .IN2(n12709), .QN(g21051) );
  NAND2X0 U13485 ( .IN1(n4396), .IN2(n11694), .QN(n12709) );
  OR2X1 U13486 ( .IN1(n11694), .IN2(n7153), .Q(n12708) );
  NAND2X0 U13487 ( .IN1(n12710), .IN2(n12711), .QN(g21047) );
  OR2X1 U13488 ( .IN1(n10335), .IN2(n6832), .Q(n12711) );
  NAND2X0 U13489 ( .IN1(n10335), .IN2(n12691), .QN(n12710) );
  NAND2X0 U13490 ( .IN1(n12712), .IN2(n12713), .QN(g21046) );
  OR2X1 U13491 ( .IN1(n12318), .IN2(n6896), .Q(n12713) );
  NAND2X0 U13492 ( .IN1(n12318), .IN2(n12292), .QN(n12712) );
  NOR2X0 U13493 ( .IN1(n4292), .IN2(n7041), .QN(n12318) );
  NAND2X0 U13494 ( .IN1(n12714), .IN2(n12715), .QN(g21045) );
  NAND2X0 U13495 ( .IN1(n11573), .IN2(n7269), .QN(n12715) );
  OR2X1 U13496 ( .IN1(n11573), .IN2(n7057), .Q(n12714) );
  NAND2X0 U13497 ( .IN1(n12716), .IN2(n12717), .QN(g21044) );
  NAND2X0 U13498 ( .IN1(n11566), .IN2(n4407), .QN(n12717) );
  OR2X1 U13499 ( .IN1(n11566), .IN2(n7058), .Q(n12716) );
  NAND2X0 U13500 ( .IN1(n12718), .IN2(n12719), .QN(g21043) );
  NAND2X0 U13501 ( .IN1(n4397), .IN2(n11563), .QN(n12719) );
  OR2X1 U13502 ( .IN1(n11563), .IN2(n7128), .Q(n12718) );
  NAND2X0 U13503 ( .IN1(n12720), .IN2(n12721), .QN(g21042) );
  OR2X1 U13504 ( .IN1(n12322), .IN2(n6897), .Q(n12721) );
  NAND2X0 U13505 ( .IN1(n12322), .IN2(n8193), .QN(n12720) );
  NAND2X0 U13506 ( .IN1(n12722), .IN2(n12723), .QN(g21041) );
  NAND2X0 U13507 ( .IN1(n11635), .IN2(n4473), .QN(n12723) );
  OR2X1 U13508 ( .IN1(n11635), .IN2(n7074), .Q(n12722) );
  NAND2X0 U13509 ( .IN1(n12724), .IN2(n12725), .QN(g21040) );
  NAND2X0 U13510 ( .IN1(n4468), .IN2(n11628), .QN(n12725) );
  OR2X1 U13511 ( .IN1(n11628), .IN2(n7075), .Q(n12724) );
  NAND2X0 U13512 ( .IN1(n12726), .IN2(n12727), .QN(g21039) );
  NAND2X0 U13513 ( .IN1(n11570), .IN2(n4409), .QN(n12727) );
  OR2X1 U13514 ( .IN1(n11570), .IN2(n7136), .Q(n12726) );
  NAND2X0 U13515 ( .IN1(n12728), .IN2(n12729), .QN(g21035) );
  NAND2X0 U13516 ( .IN1(n4395), .IN2(n11700), .QN(n12729) );
  OR2X1 U13517 ( .IN1(n11700), .IN2(n7091), .Q(n12728) );
  NAND2X0 U13518 ( .IN1(n12730), .IN2(n12731), .QN(g21034) );
  NAND2X0 U13519 ( .IN1(n11690), .IN2(n4475), .QN(n12731) );
  OR2X1 U13520 ( .IN1(n11690), .IN2(n7092), .Q(n12730) );
  NAND2X0 U13521 ( .IN1(n12732), .IN2(n12733), .QN(g21033) );
  NAND2X0 U13522 ( .IN1(n4469), .IN2(n11632), .QN(n12733) );
  OR2X1 U13523 ( .IN1(n11632), .IN2(n7145), .Q(n12732) );
  NAND2X0 U13524 ( .IN1(n12734), .IN2(n12735), .QN(g21032) );
  NAND2X0 U13525 ( .IN1(n4396), .IN2(n11755), .QN(n12735) );
  OR2X1 U13526 ( .IN1(n11755), .IN2(n7107), .Q(n12734) );
  NAND2X0 U13527 ( .IN1(n12736), .IN2(n12737), .QN(g21031) );
  NAND2X0 U13528 ( .IN1(n11694), .IN2(n4477), .QN(n12737) );
  OR2X1 U13529 ( .IN1(n11694), .IN2(n7154), .Q(n12736) );
  NAND2X0 U13530 ( .IN1(n12738), .IN2(n12739), .QN(g21029) );
  OR2X1 U13531 ( .IN1(n12325), .IN2(n6840), .Q(n12739) );
  NAND2X0 U13532 ( .IN1(n12325), .IN2(n12691), .QN(n12738) );
  INVX0 U13533 ( .INP(n7981), .ZN(n12691) );
  NAND3X0 U13534 ( .IN1(n12740), .IN2(n12741), .IN3(n12742), .QN(n7981) );
  NAND2X0 U13535 ( .IN1(test_so90), .IN2(g7390), .QN(n12742) );
  NAND2X0 U13536 ( .IN1(g7302), .IN2(g2679), .QN(n12741) );
  NAND2X0 U13537 ( .IN1(g2624), .IN2(g2685), .QN(n12740) );
  NAND2X0 U13538 ( .IN1(n12743), .IN2(n12744), .QN(g21028) );
  NAND2X0 U13539 ( .IN1(n10974), .IN2(g2804), .QN(n12744) );
  INVX0 U13540 ( .INP(n10335), .ZN(n10974) );
  NAND2X0 U13541 ( .IN1(n10335), .IN2(n12292), .QN(n12743) );
  NAND2X0 U13542 ( .IN1(n12745), .IN2(n12746), .QN(g21027) );
  NAND2X0 U13543 ( .IN1(n11573), .IN2(n4407), .QN(n12746) );
  OR2X1 U13544 ( .IN1(n11573), .IN2(n7059), .Q(n12745) );
  NAND2X0 U13545 ( .IN1(n12747), .IN2(n12748), .QN(g21026) );
  NAND2X0 U13546 ( .IN1(n4397), .IN2(n11566), .QN(n12748) );
  OR2X1 U13547 ( .IN1(n11566), .IN2(n7060), .Q(n12747) );
  NAND2X0 U13548 ( .IN1(n12749), .IN2(n12750), .QN(g21025) );
  NAND2X0 U13549 ( .IN1(test_so93), .IN2(n12670), .QN(n12750) );
  NAND2X0 U13550 ( .IN1(n11563), .IN2(n4408), .QN(n12749) );
  NAND2X0 U13551 ( .IN1(n12751), .IN2(n12752), .QN(g21023) );
  OR2X1 U13552 ( .IN1(n10339), .IN2(n6834), .Q(n12752) );
  NAND2X0 U13553 ( .IN1(n10339), .IN2(n8193), .QN(n12751) );
  NAND2X0 U13554 ( .IN1(n12753), .IN2(n12754), .QN(g21022) );
  OR2X1 U13555 ( .IN1(n12322), .IN2(n6898), .Q(n12754) );
  NAND2X0 U13556 ( .IN1(n12322), .IN2(n8167), .QN(n12753) );
  NOR2X0 U13557 ( .IN1(n4293), .IN2(n7042), .QN(n12322) );
  NAND2X0 U13558 ( .IN1(n12755), .IN2(n12756), .QN(g21021) );
  NAND2X0 U13559 ( .IN1(n4468), .IN2(n11635), .QN(n12756) );
  OR2X1 U13560 ( .IN1(n11635), .IN2(n7076), .Q(n12755) );
  NAND2X0 U13561 ( .IN1(n12757), .IN2(n12758), .QN(g21020) );
  NAND2X0 U13562 ( .IN1(n11628), .IN2(n4409), .QN(n12758) );
  OR2X1 U13563 ( .IN1(n11628), .IN2(n7077), .Q(n12757) );
  NAND2X0 U13564 ( .IN1(n12759), .IN2(n12760), .QN(g21019) );
  NAND2X0 U13565 ( .IN1(n4399), .IN2(n11570), .QN(n12760) );
  OR2X1 U13566 ( .IN1(n11570), .IN2(n7137), .Q(n12759) );
  NAND2X0 U13567 ( .IN1(n12761), .IN2(n12762), .QN(g21018) );
  OR2X1 U13568 ( .IN1(n12330), .IN2(n6899), .Q(n12762) );
  NAND2X0 U13569 ( .IN1(n12330), .IN2(n8304), .QN(n12761) );
  NAND2X0 U13570 ( .IN1(n12763), .IN2(n12764), .QN(g21017) );
  NAND2X0 U13571 ( .IN1(n11700), .IN2(n4475), .QN(n12764) );
  OR2X1 U13572 ( .IN1(n11700), .IN2(n7093), .Q(n12763) );
  NAND2X0 U13573 ( .IN1(n12765), .IN2(n12766), .QN(g21016) );
  NAND2X0 U13574 ( .IN1(n4469), .IN2(n11690), .QN(n12766) );
  OR2X1 U13575 ( .IN1(n11690), .IN2(n7094), .Q(n12765) );
  NAND2X0 U13576 ( .IN1(n12767), .IN2(n12768), .QN(g21015) );
  NAND2X0 U13577 ( .IN1(n11632), .IN2(n4411), .QN(n12768) );
  OR2X1 U13578 ( .IN1(n11632), .IN2(n7146), .Q(n12767) );
  NAND2X0 U13579 ( .IN1(n12769), .IN2(n12770), .QN(g21011) );
  NAND2X0 U13580 ( .IN1(n4396), .IN2(n11758), .QN(n12770) );
  OR2X1 U13581 ( .IN1(n11758), .IN2(n7108), .Q(n12769) );
  NAND2X0 U13582 ( .IN1(n12771), .IN2(n12772), .QN(g21010) );
  NAND2X0 U13583 ( .IN1(n11755), .IN2(n4477), .QN(n12772) );
  OR2X1 U13584 ( .IN1(n11755), .IN2(n7109), .Q(n12771) );
  NAND2X0 U13585 ( .IN1(n12773), .IN2(n12774), .QN(g21009) );
  NAND2X0 U13586 ( .IN1(n11694), .IN2(n7270), .QN(n12774) );
  OR2X1 U13587 ( .IN1(n11694), .IN2(n7155), .Q(n12773) );
  NAND2X0 U13588 ( .IN1(n12775), .IN2(n12776), .QN(g21007) );
  OR2X1 U13589 ( .IN1(n12325), .IN2(n6841), .Q(n12776) );
  NAND2X0 U13590 ( .IN1(n12325), .IN2(n12292), .QN(n12775) );
  INVX0 U13591 ( .INP(n7994), .ZN(n12292) );
  NAND3X0 U13592 ( .IN1(n12777), .IN2(n12778), .IN3(n12779), .QN(n7994) );
  NAND2X0 U13593 ( .IN1(g7390), .IN2(g2691), .QN(n12779) );
  NAND2X0 U13594 ( .IN1(g2624), .IN2(g2694), .QN(n12778) );
  NAND2X0 U13595 ( .IN1(n9246), .IN2(g2688), .QN(n12777) );
  INVX0 U13596 ( .INP(n4314), .ZN(n9246) );
  NOR2X0 U13597 ( .IN1(n4306), .IN2(n7041), .QN(n12325) );
  NAND2X0 U13598 ( .IN1(n12780), .IN2(n12781), .QN(g21006) );
  NAND2X0 U13599 ( .IN1(n4397), .IN2(n11573), .QN(n12781) );
  OR2X1 U13600 ( .IN1(n11573), .IN2(n7061), .Q(n12780) );
  NAND2X0 U13601 ( .IN1(n12782), .IN2(n12783), .QN(g21005) );
  NAND2X0 U13602 ( .IN1(n11566), .IN2(n4408), .QN(n12783) );
  OR2X1 U13603 ( .IN1(n11566), .IN2(n7062), .Q(n12782) );
  NAND2X0 U13604 ( .IN1(n12784), .IN2(n12785), .QN(g21004) );
  NAND2X0 U13605 ( .IN1(n4419), .IN2(n11563), .QN(n12785) );
  OR2X1 U13606 ( .IN1(n11563), .IN2(n7129), .Q(n12784) );
  NAND2X0 U13607 ( .IN1(n12786), .IN2(n12787), .QN(g21003) );
  OR2X1 U13608 ( .IN1(n12332), .IN2(n6842), .Q(n12787) );
  NAND2X0 U13609 ( .IN1(n12332), .IN2(n8193), .QN(n12786) );
  INVX0 U13610 ( .INP(n8173), .ZN(n8193) );
  NAND3X0 U13611 ( .IN1(n12788), .IN2(n12789), .IN3(n12790), .QN(n8173) );
  NAND2X0 U13612 ( .IN1(g1930), .IN2(g1991), .QN(n12790) );
  NAND2X0 U13613 ( .IN1(g7052), .IN2(g1985), .QN(n12789) );
  NAND2X0 U13614 ( .IN1(g7194), .IN2(g1988), .QN(n12788) );
  NAND2X0 U13615 ( .IN1(n12791), .IN2(n12792), .QN(g21002) );
  NAND2X0 U13616 ( .IN1(n12632), .IN2(g2110), .QN(n12792) );
  INVX0 U13617 ( .INP(n10339), .ZN(n12632) );
  NAND2X0 U13618 ( .IN1(n10339), .IN2(n8167), .QN(n12791) );
  NAND2X0 U13619 ( .IN1(n12793), .IN2(n12794), .QN(g21001) );
  NAND2X0 U13620 ( .IN1(n11635), .IN2(n4409), .QN(n12794) );
  OR2X1 U13621 ( .IN1(n11635), .IN2(n7078), .Q(n12793) );
  NAND2X0 U13622 ( .IN1(n12795), .IN2(n12796), .QN(g21000) );
  NAND2X0 U13623 ( .IN1(test_so71), .IN2(n12329), .QN(n12796) );
  NAND2X0 U13624 ( .IN1(n4399), .IN2(n11628), .QN(n12795) );
  NAND2X0 U13625 ( .IN1(n12797), .IN2(n12798), .QN(g20999) );
  NAND2X0 U13626 ( .IN1(n11570), .IN2(n4410), .QN(n12798) );
  OR2X1 U13627 ( .IN1(n11570), .IN2(n7138), .Q(n12797) );
  NAND2X0 U13628 ( .IN1(n12799), .IN2(n12800), .QN(g20997) );
  OR2X1 U13629 ( .IN1(n10343), .IN2(n6836), .Q(n12800) );
  NAND2X0 U13630 ( .IN1(n10343), .IN2(n8304), .QN(n12799) );
  NAND2X0 U13631 ( .IN1(n12801), .IN2(n12802), .QN(g20996) );
  NAND2X0 U13632 ( .IN1(test_so51), .IN2(n12803), .QN(n12802) );
  INVX0 U13633 ( .INP(n12330), .ZN(n12803) );
  NAND2X0 U13634 ( .IN1(n12330), .IN2(n12306), .QN(n12801) );
  NOR2X0 U13635 ( .IN1(n4294), .IN2(n7043), .QN(n12330) );
  NAND2X0 U13636 ( .IN1(n12804), .IN2(n12805), .QN(g20995) );
  NAND2X0 U13637 ( .IN1(n4469), .IN2(n11700), .QN(n12805) );
  OR2X1 U13638 ( .IN1(n11700), .IN2(n7095), .Q(n12804) );
  NAND2X0 U13639 ( .IN1(n12806), .IN2(n12807), .QN(g20994) );
  NAND2X0 U13640 ( .IN1(test_so50), .IN2(n12336), .QN(n12807) );
  NAND2X0 U13641 ( .IN1(n11690), .IN2(n4411), .QN(n12806) );
  NAND2X0 U13642 ( .IN1(n12808), .IN2(n12809), .QN(g20993) );
  NAND2X0 U13643 ( .IN1(n4401), .IN2(n11632), .QN(n12809) );
  OR2X1 U13644 ( .IN1(n11632), .IN2(n7147), .Q(n12808) );
  NAND2X0 U13645 ( .IN1(n12810), .IN2(n12811), .QN(g20992) );
  OR2X1 U13646 ( .IN1(n12337), .IN2(n6900), .Q(n12811) );
  NAND2X0 U13647 ( .IN1(n12337), .IN2(n12812), .QN(n12810) );
  NAND2X0 U13648 ( .IN1(n12813), .IN2(n12814), .QN(g20991) );
  NAND2X0 U13649 ( .IN1(n11758), .IN2(n4477), .QN(n12814) );
  OR2X1 U13650 ( .IN1(n11758), .IN2(n7110), .Q(n12813) );
  NAND2X0 U13651 ( .IN1(n12815), .IN2(n12816), .QN(g20990) );
  NAND2X0 U13652 ( .IN1(n11755), .IN2(n7270), .QN(n12816) );
  OR2X1 U13653 ( .IN1(n11755), .IN2(n7111), .Q(n12815) );
  NAND2X0 U13654 ( .IN1(n12817), .IN2(n12818), .QN(g20989) );
  NAND2X0 U13655 ( .IN1(n11694), .IN2(n4413), .QN(n12818) );
  OR2X1 U13656 ( .IN1(n11694), .IN2(n7156), .Q(n12817) );
  NAND2X0 U13657 ( .IN1(n12819), .IN2(n12820), .QN(g20983) );
  NAND2X0 U13658 ( .IN1(n11573), .IN2(n4408), .QN(n12820) );
  OR2X1 U13659 ( .IN1(n11573), .IN2(n7063), .Q(n12819) );
  NAND2X0 U13660 ( .IN1(n12821), .IN2(n12822), .QN(g20982) );
  NAND2X0 U13661 ( .IN1(n4419), .IN2(n11566), .QN(n12822) );
  OR2X1 U13662 ( .IN1(n11566), .IN2(n7064), .Q(n12821) );
  NAND2X0 U13663 ( .IN1(n12823), .IN2(n12824), .QN(g20981) );
  NAND2X0 U13664 ( .IN1(n11563), .IN2(n4472), .QN(n12824) );
  OR2X1 U13665 ( .IN1(n11563), .IN2(n7130), .Q(n12823) );
  NAND2X0 U13666 ( .IN1(n12825), .IN2(n12826), .QN(g20980) );
  OR2X1 U13667 ( .IN1(n12332), .IN2(n6843), .Q(n12826) );
  NAND2X0 U13668 ( .IN1(n12332), .IN2(n8167), .QN(n12825) );
  INVX0 U13669 ( .INP(n8181), .ZN(n8167) );
  NAND3X0 U13670 ( .IN1(n12827), .IN2(n12828), .IN3(n12829), .QN(n8181) );
  NAND2X0 U13671 ( .IN1(g1930), .IN2(g2000), .QN(n12829) );
  NAND2X0 U13672 ( .IN1(n9268), .IN2(g1994), .QN(n12828) );
  INVX0 U13673 ( .INP(n4296), .ZN(n9268) );
  NAND2X0 U13674 ( .IN1(g7194), .IN2(g1997), .QN(n12827) );
  NOR2X0 U13675 ( .IN1(n4307), .IN2(n7042), .QN(n12332) );
  NAND2X0 U13676 ( .IN1(n12830), .IN2(n12831), .QN(g20979) );
  NAND2X0 U13677 ( .IN1(n4399), .IN2(n11635), .QN(n12831) );
  OR2X1 U13678 ( .IN1(n11635), .IN2(n7079), .Q(n12830) );
  NAND2X0 U13679 ( .IN1(n12832), .IN2(n12833), .QN(g20978) );
  NAND2X0 U13680 ( .IN1(n11628), .IN2(n4410), .QN(n12833) );
  OR2X1 U13681 ( .IN1(n11628), .IN2(n7080), .Q(n12832) );
  NAND2X0 U13682 ( .IN1(n12834), .IN2(n12835), .QN(g20977) );
  NAND2X0 U13683 ( .IN1(n4420), .IN2(n11570), .QN(n12835) );
  OR2X1 U13684 ( .IN1(n11570), .IN2(n7139), .Q(n12834) );
  NAND2X0 U13685 ( .IN1(n12836), .IN2(n12837), .QN(g20976) );
  OR2X1 U13686 ( .IN1(n12340), .IN2(n6844), .Q(n12837) );
  NAND2X0 U13687 ( .IN1(n12340), .IN2(n8304), .QN(n12836) );
  INVX0 U13688 ( .INP(n8285), .ZN(n8304) );
  NAND3X0 U13689 ( .IN1(n12838), .IN2(n12839), .IN3(n12840), .QN(n8285) );
  NAND2X0 U13690 ( .IN1(g6944), .IN2(g1294), .QN(n12840) );
  NAND2X0 U13691 ( .IN1(g6750), .IN2(g1291), .QN(n12839) );
  NAND2X0 U13692 ( .IN1(g1236), .IN2(g1297), .QN(n12838) );
  NAND2X0 U13693 ( .IN1(n12841), .IN2(n12842), .QN(g20975) );
  OR2X1 U13694 ( .IN1(n10343), .IN2(n6837), .Q(n12842) );
  NAND2X0 U13695 ( .IN1(n10343), .IN2(n12306), .QN(n12841) );
  NAND2X0 U13696 ( .IN1(n12843), .IN2(n12844), .QN(g20974) );
  NAND2X0 U13697 ( .IN1(n11700), .IN2(n4411), .QN(n12844) );
  OR2X1 U13698 ( .IN1(n11700), .IN2(n7096), .Q(n12843) );
  NAND2X0 U13699 ( .IN1(n12845), .IN2(n12846), .QN(g20973) );
  NAND2X0 U13700 ( .IN1(n4401), .IN2(n11690), .QN(n12846) );
  OR2X1 U13701 ( .IN1(n11690), .IN2(n7097), .Q(n12845) );
  NAND2X0 U13702 ( .IN1(n12847), .IN2(n12848), .QN(g20972) );
  NAND2X0 U13703 ( .IN1(n11632), .IN2(n4412), .QN(n12848) );
  OR2X1 U13704 ( .IN1(n11632), .IN2(n7148), .Q(n12847) );
  NAND2X0 U13705 ( .IN1(n12849), .IN2(n12850), .QN(g20970) );
  OR2X1 U13706 ( .IN1(n9912), .IN2(n6838), .Q(n12850) );
  NAND2X0 U13707 ( .IN1(n9912), .IN2(n12812), .QN(n12849) );
  NAND2X0 U13708 ( .IN1(n12851), .IN2(n12852), .QN(g20969) );
  OR2X1 U13709 ( .IN1(n12337), .IN2(n6901), .Q(n12852) );
  NAND2X0 U13710 ( .IN1(n12337), .IN2(n12313), .QN(n12851) );
  NOR2X0 U13711 ( .IN1(n4295), .IN2(n7044), .QN(n12337) );
  NAND2X0 U13712 ( .IN1(n12853), .IN2(n12854), .QN(g20968) );
  NAND2X0 U13713 ( .IN1(n11758), .IN2(n7270), .QN(n12854) );
  OR2X1 U13714 ( .IN1(n11758), .IN2(n7112), .Q(n12853) );
  NAND2X0 U13715 ( .IN1(n12855), .IN2(n12856), .QN(g20967) );
  NAND2X0 U13716 ( .IN1(n11755), .IN2(n4413), .QN(n12856) );
  OR2X1 U13717 ( .IN1(n11755), .IN2(n7113), .Q(n12855) );
  NAND2X0 U13718 ( .IN1(n12857), .IN2(n12858), .QN(g20966) );
  NAND2X0 U13719 ( .IN1(n4403), .IN2(n11694), .QN(n12858) );
  OR2X1 U13720 ( .IN1(n11694), .IN2(n7157), .Q(n12857) );
  NAND2X0 U13721 ( .IN1(n12859), .IN2(n12860), .QN(g20965) );
  NAND2X0 U13722 ( .IN1(n4415), .IN2(n11563), .QN(n12860) );
  OR2X1 U13723 ( .IN1(n11563), .IN2(n7124), .Q(n12859) );
  NAND2X0 U13724 ( .IN1(n12861), .IN2(n12862), .QN(g20964) );
  NAND2X0 U13725 ( .IN1(n4419), .IN2(n11573), .QN(n12862) );
  OR2X1 U13726 ( .IN1(n11573), .IN2(n7065), .Q(n12861) );
  NAND2X0 U13727 ( .IN1(n12863), .IN2(n12864), .QN(g20963) );
  NAND2X0 U13728 ( .IN1(n11566), .IN2(n4472), .QN(n12864) );
  OR2X1 U13729 ( .IN1(n11566), .IN2(n7066), .Q(n12863) );
  NAND2X0 U13730 ( .IN1(n12865), .IN2(n12866), .QN(g20962) );
  NAND2X0 U13731 ( .IN1(n4398), .IN2(n11563), .QN(n12866) );
  OR2X1 U13732 ( .IN1(n11563), .IN2(n7131), .Q(n12865) );
  INVX0 U13733 ( .INP(n12670), .ZN(n11563) );
  NAND2X0 U13734 ( .IN1(n12867), .IN2(g2703), .QN(n12670) );
  NAND2X0 U13735 ( .IN1(n12868), .IN2(n12869), .QN(g20955) );
  NAND2X0 U13736 ( .IN1(n11635), .IN2(n4410), .QN(n12869) );
  OR2X1 U13737 ( .IN1(n11635), .IN2(n7081), .Q(n12868) );
  NAND2X0 U13738 ( .IN1(n12870), .IN2(n12871), .QN(g20954) );
  NAND2X0 U13739 ( .IN1(n4420), .IN2(n11628), .QN(n12871) );
  OR2X1 U13740 ( .IN1(n11628), .IN2(n7082), .Q(n12870) );
  NAND2X0 U13741 ( .IN1(n12872), .IN2(n12873), .QN(g20953) );
  NAND2X0 U13742 ( .IN1(n11570), .IN2(n4474), .QN(n12873) );
  OR2X1 U13743 ( .IN1(n11570), .IN2(n7140), .Q(n12872) );
  NAND2X0 U13744 ( .IN1(n12874), .IN2(n12875), .QN(g20952) );
  OR2X1 U13745 ( .IN1(n12340), .IN2(n6845), .Q(n12875) );
  NAND2X0 U13746 ( .IN1(n12340), .IN2(n12306), .QN(n12874) );
  INVX0 U13747 ( .INP(n8278), .ZN(n12306) );
  NAND3X0 U13748 ( .IN1(n12876), .IN2(n12877), .IN3(n12878), .QN(n8278) );
  NAND2X0 U13749 ( .IN1(n10142), .IN2(g1300), .QN(n12878) );
  INVX0 U13750 ( .INP(n4371), .ZN(n10142) );
  NAND2X0 U13751 ( .IN1(g1236), .IN2(g1306), .QN(n12877) );
  NAND2X0 U13752 ( .IN1(g6944), .IN2(g1303), .QN(n12876) );
  NOR2X0 U13753 ( .IN1(n4308), .IN2(n7043), .QN(n12340) );
  NAND2X0 U13754 ( .IN1(n12879), .IN2(n12880), .QN(g20951) );
  NAND2X0 U13755 ( .IN1(n4401), .IN2(n11700), .QN(n12880) );
  OR2X1 U13756 ( .IN1(n11700), .IN2(n7098), .Q(n12879) );
  NAND2X0 U13757 ( .IN1(n12881), .IN2(n12882), .QN(g20950) );
  NAND2X0 U13758 ( .IN1(n11690), .IN2(n4412), .QN(n12882) );
  OR2X1 U13759 ( .IN1(n11690), .IN2(n7099), .Q(n12881) );
  NAND2X0 U13760 ( .IN1(n12883), .IN2(n12884), .QN(g20949) );
  NAND2X0 U13761 ( .IN1(n4421), .IN2(n11632), .QN(n12884) );
  OR2X1 U13762 ( .IN1(n11632), .IN2(n7149), .Q(n12883) );
  NAND2X0 U13763 ( .IN1(n12885), .IN2(n12886), .QN(g20948) );
  OR2X1 U13764 ( .IN1(n12345), .IN2(n6846), .Q(n12886) );
  NAND2X0 U13765 ( .IN1(n12345), .IN2(n12812), .QN(n12885) );
  INVX0 U13766 ( .INP(n7851), .ZN(n12812) );
  NAND3X0 U13767 ( .IN1(n12887), .IN2(n12888), .IN3(n12889), .QN(n7851) );
  NAND2X0 U13768 ( .IN1(g6642), .IN2(g608), .QN(n12889) );
  NAND2X0 U13769 ( .IN1(n10242), .IN2(g605), .QN(n12888) );
  INVX0 U13770 ( .INP(n4298), .ZN(n10242) );
  NAND2X0 U13771 ( .IN1(g550), .IN2(g611), .QN(n12887) );
  NAND2X0 U13772 ( .IN1(n12890), .IN2(n12891), .QN(g20947) );
  NAND2X0 U13773 ( .IN1(n10461), .IN2(g730), .QN(n12891) );
  INVX0 U13774 ( .INP(n9912), .ZN(n10461) );
  NAND2X0 U13775 ( .IN1(n9912), .IN2(n12313), .QN(n12890) );
  NAND2X0 U13776 ( .IN1(n12892), .IN2(n12893), .QN(g20946) );
  NAND2X0 U13777 ( .IN1(n11758), .IN2(n4413), .QN(n12893) );
  OR2X1 U13778 ( .IN1(n11758), .IN2(n7114), .Q(n12892) );
  NAND2X0 U13779 ( .IN1(n12894), .IN2(n12895), .QN(g20945) );
  NAND2X0 U13780 ( .IN1(n4403), .IN2(n11755), .QN(n12895) );
  OR2X1 U13781 ( .IN1(n11755), .IN2(n7115), .Q(n12894) );
  NAND2X0 U13782 ( .IN1(n12896), .IN2(n12897), .QN(g20944) );
  NAND2X0 U13783 ( .IN1(n11694), .IN2(n4414), .QN(n12897) );
  OR2X1 U13784 ( .IN1(n11694), .IN2(n7158), .Q(n12896) );
  NAND2X0 U13785 ( .IN1(n12898), .IN2(n12899), .QN(g20941) );
  NAND2X0 U13786 ( .IN1(n4415), .IN2(n11566), .QN(n12899) );
  OR2X1 U13787 ( .IN1(n11566), .IN2(n7050), .Q(n12898) );
  NAND2X0 U13788 ( .IN1(n12900), .IN2(n12901), .QN(g20940) );
  NAND2X0 U13789 ( .IN1(n11573), .IN2(n4472), .QN(n12901) );
  OR2X1 U13790 ( .IN1(n11573), .IN2(n7067), .Q(n12900) );
  NAND2X0 U13791 ( .IN1(n12902), .IN2(n12903), .QN(g20939) );
  NAND2X0 U13792 ( .IN1(n4398), .IN2(n11566), .QN(n12903) );
  OR2X1 U13793 ( .IN1(n11566), .IN2(n7068), .Q(n12902) );
  INVX0 U13794 ( .INP(n12321), .ZN(n11566) );
  NAND2X0 U13795 ( .IN1(n12867), .IN2(g7487), .QN(n12321) );
  NAND2X0 U13796 ( .IN1(n12904), .IN2(n12905), .QN(g20937) );
  NAND2X0 U13797 ( .IN1(n4416), .IN2(n11570), .QN(n12905) );
  OR2X1 U13798 ( .IN1(n11570), .IN2(n7132), .Q(n12904) );
  NAND2X0 U13799 ( .IN1(n12906), .IN2(n12907), .QN(g20936) );
  NAND2X0 U13800 ( .IN1(n4420), .IN2(n11635), .QN(n12907) );
  OR2X1 U13801 ( .IN1(n11635), .IN2(n7083), .Q(n12906) );
  NAND2X0 U13802 ( .IN1(n12908), .IN2(n12909), .QN(g20935) );
  NAND2X0 U13803 ( .IN1(n11628), .IN2(n4474), .QN(n12909) );
  OR2X1 U13804 ( .IN1(n11628), .IN2(n7084), .Q(n12908) );
  NAND2X0 U13805 ( .IN1(n12910), .IN2(n12911), .QN(g20934) );
  NAND2X0 U13806 ( .IN1(n4400), .IN2(n11570), .QN(n12911) );
  OR2X1 U13807 ( .IN1(n11570), .IN2(n7141), .Q(n12910) );
  INVX0 U13808 ( .INP(n12324), .ZN(n11570) );
  NAND3X0 U13809 ( .IN1(n12635), .IN2(g1905), .IN3(test_so69), .QN(n12324) );
  NAND2X0 U13810 ( .IN1(n12912), .IN2(n12913), .QN(g20927) );
  NAND2X0 U13811 ( .IN1(n11700), .IN2(n4412), .QN(n12913) );
  OR2X1 U13812 ( .IN1(n11700), .IN2(n7100), .Q(n12912) );
  NAND2X0 U13813 ( .IN1(n12914), .IN2(n12915), .QN(g20926) );
  NAND2X0 U13814 ( .IN1(n4421), .IN2(n11690), .QN(n12915) );
  OR2X1 U13815 ( .IN1(n11690), .IN2(n7101), .Q(n12914) );
  NAND2X0 U13816 ( .IN1(n12916), .IN2(n12917), .QN(g20925) );
  NAND2X0 U13817 ( .IN1(n11632), .IN2(n4476), .QN(n12917) );
  OR2X1 U13818 ( .IN1(n11632), .IN2(n7150), .Q(n12916) );
  NAND2X0 U13819 ( .IN1(n12918), .IN2(n12919), .QN(g20924) );
  OR2X1 U13820 ( .IN1(n12345), .IN2(n6847), .Q(n12919) );
  NAND2X0 U13821 ( .IN1(n12345), .IN2(n12313), .QN(n12918) );
  INVX0 U13822 ( .INP(n7844), .ZN(n12313) );
  NAND3X0 U13823 ( .IN1(n12920), .IN2(n12921), .IN3(n12922), .QN(n7844) );
  NAND2X0 U13824 ( .IN1(g6642), .IN2(g617), .QN(n12922) );
  NAND2X0 U13825 ( .IN1(g6485), .IN2(g614), .QN(n12921) );
  NAND2X0 U13826 ( .IN1(test_so26), .IN2(g550), .QN(n12920) );
  NOR2X0 U13827 ( .IN1(n4309), .IN2(n7044), .QN(n12345) );
  NAND2X0 U13828 ( .IN1(n12923), .IN2(n12924), .QN(g20923) );
  NAND2X0 U13829 ( .IN1(test_so29), .IN2(n12347), .QN(n12924) );
  NAND2X0 U13830 ( .IN1(n4403), .IN2(n11758), .QN(n12923) );
  NAND2X0 U13831 ( .IN1(n12925), .IN2(n12926), .QN(g20922) );
  NAND2X0 U13832 ( .IN1(n11755), .IN2(n4414), .QN(n12926) );
  OR2X1 U13833 ( .IN1(n11755), .IN2(n7116), .Q(n12925) );
  NAND2X0 U13834 ( .IN1(n12927), .IN2(n12928), .QN(g20921) );
  NAND2X0 U13835 ( .IN1(n4422), .IN2(n11694), .QN(n12928) );
  OR2X1 U13836 ( .IN1(n11694), .IN2(n7159), .Q(n12927) );
  NAND2X0 U13837 ( .IN1(n12929), .IN2(n12930), .QN(g20919) );
  NAND2X0 U13838 ( .IN1(n4415), .IN2(n11573), .QN(n12930) );
  OR2X1 U13839 ( .IN1(n11573), .IN2(n7051), .Q(n12929) );
  NAND2X0 U13840 ( .IN1(n12931), .IN2(n12932), .QN(g20918) );
  NAND2X0 U13841 ( .IN1(n4398), .IN2(n11573), .QN(n12932) );
  OR2X1 U13842 ( .IN1(n11573), .IN2(n7069), .Q(n12931) );
  INVX0 U13843 ( .INP(n12327), .ZN(n11573) );
  NAND2X0 U13844 ( .IN1(n12867), .IN2(g7425), .QN(n12327) );
  NOR3X0 U13845 ( .IN1(n4490), .IN2(n7002), .IN3(g2733), .QN(n12867) );
  NAND2X0 U13846 ( .IN1(n12933), .IN2(n12934), .QN(g20917) );
  NAND2X0 U13847 ( .IN1(test_so72), .IN2(n12329), .QN(n12934) );
  NAND2X0 U13848 ( .IN1(n4416), .IN2(n11628), .QN(n12933) );
  NAND2X0 U13849 ( .IN1(n12935), .IN2(n12936), .QN(g20916) );
  NAND2X0 U13850 ( .IN1(n11635), .IN2(n4474), .QN(n12936) );
  OR2X1 U13851 ( .IN1(n11635), .IN2(n7085), .Q(n12935) );
  NAND2X0 U13852 ( .IN1(n12937), .IN2(n12938), .QN(g20915) );
  NAND2X0 U13853 ( .IN1(n4400), .IN2(n11628), .QN(n12938) );
  OR2X1 U13854 ( .IN1(n11628), .IN2(n7086), .Q(n12937) );
  INVX0 U13855 ( .INP(n12329), .ZN(n11628) );
  NAND2X0 U13856 ( .IN1(n12939), .IN2(g7357), .QN(n12329) );
  NAND2X0 U13857 ( .IN1(n12940), .IN2(n12941), .QN(g20913) );
  NAND2X0 U13858 ( .IN1(n4417), .IN2(n11632), .QN(n12941) );
  OR2X1 U13859 ( .IN1(n11632), .IN2(n7142), .Q(n12940) );
  NAND2X0 U13860 ( .IN1(n12942), .IN2(n12943), .QN(g20912) );
  NAND2X0 U13861 ( .IN1(n4421), .IN2(n11700), .QN(n12943) );
  OR2X1 U13862 ( .IN1(n11700), .IN2(n7102), .Q(n12942) );
  NAND2X0 U13863 ( .IN1(n12944), .IN2(n12945), .QN(g20911) );
  NAND2X0 U13864 ( .IN1(n11690), .IN2(n4476), .QN(n12945) );
  OR2X1 U13865 ( .IN1(n11690), .IN2(n7103), .Q(n12944) );
  NAND2X0 U13866 ( .IN1(n12946), .IN2(n12947), .QN(g20910) );
  NAND2X0 U13867 ( .IN1(n4402), .IN2(n11632), .QN(n12947) );
  OR2X1 U13868 ( .IN1(n11632), .IN2(n7151), .Q(n12946) );
  NOR3X0 U13869 ( .IN1(n4489), .IN2(n7004), .IN3(n12643), .QN(n11632) );
  NAND2X0 U13870 ( .IN1(n12948), .IN2(n12949), .QN(g20903) );
  NAND2X0 U13871 ( .IN1(n11758), .IN2(n4414), .QN(n12949) );
  OR2X1 U13872 ( .IN1(n11758), .IN2(n7117), .Q(n12948) );
  NAND2X0 U13873 ( .IN1(n12950), .IN2(n12951), .QN(g20902) );
  NAND2X0 U13874 ( .IN1(n4422), .IN2(n11755), .QN(n12951) );
  OR2X1 U13875 ( .IN1(n11755), .IN2(n7118), .Q(n12950) );
  NAND2X0 U13876 ( .IN1(n12952), .IN2(n12953), .QN(g20901) );
  NAND2X0 U13877 ( .IN1(n11694), .IN2(n4478), .QN(n12953) );
  OR2X1 U13878 ( .IN1(n11694), .IN2(n7160), .Q(n12952) );
  NAND2X0 U13879 ( .IN1(n12954), .IN2(n12955), .QN(g20900) );
  NAND2X0 U13880 ( .IN1(n4416), .IN2(n11635), .QN(n12955) );
  OR2X1 U13881 ( .IN1(n11635), .IN2(n7070), .Q(n12954) );
  NAND2X0 U13882 ( .IN1(n12956), .IN2(n12957), .QN(g20899) );
  NAND2X0 U13883 ( .IN1(n4400), .IN2(n11635), .QN(n12957) );
  OR2X1 U13884 ( .IN1(n11635), .IN2(n7087), .Q(n12956) );
  INVX0 U13885 ( .INP(n12334), .ZN(n11635) );
  NAND2X0 U13886 ( .IN1(n12939), .IN2(g7229), .QN(n12334) );
  AND3X1 U13887 ( .IN1(n4427), .IN2(g1905), .IN3(test_so69), .Q(n12939) );
  NAND2X0 U13888 ( .IN1(n12958), .IN2(n12959), .QN(g20898) );
  NAND2X0 U13889 ( .IN1(n4417), .IN2(n11690), .QN(n12959) );
  OR2X1 U13890 ( .IN1(n11690), .IN2(n7088), .Q(n12958) );
  NAND2X0 U13891 ( .IN1(n12960), .IN2(n12961), .QN(g20897) );
  NAND2X0 U13892 ( .IN1(n11700), .IN2(n4476), .QN(n12961) );
  OR2X1 U13893 ( .IN1(n11700), .IN2(n7104), .Q(n12960) );
  NAND2X0 U13894 ( .IN1(n12962), .IN2(n12963), .QN(g20896) );
  NAND2X0 U13895 ( .IN1(n4402), .IN2(n11690), .QN(n12963) );
  OR2X1 U13896 ( .IN1(n11690), .IN2(n7105), .Q(n12962) );
  INVX0 U13897 ( .INP(n12336), .ZN(n11690) );
  NAND2X0 U13898 ( .IN1(n12964), .IN2(g7161), .QN(n12336) );
  NAND2X0 U13899 ( .IN1(n12965), .IN2(n12966), .QN(g20894) );
  NAND2X0 U13900 ( .IN1(n4418), .IN2(n11694), .QN(n12966) );
  OR2X1 U13901 ( .IN1(n11694), .IN2(n7152), .Q(n12965) );
  NAND2X0 U13902 ( .IN1(n12967), .IN2(n12968), .QN(g20893) );
  NAND2X0 U13903 ( .IN1(n4422), .IN2(n11758), .QN(n12968) );
  OR2X1 U13904 ( .IN1(n11758), .IN2(n7119), .Q(n12967) );
  NAND2X0 U13905 ( .IN1(n12969), .IN2(n12970), .QN(g20892) );
  NAND2X0 U13906 ( .IN1(n11755), .IN2(n4478), .QN(n12970) );
  OR2X1 U13907 ( .IN1(n11755), .IN2(n7120), .Q(n12969) );
  NAND2X0 U13908 ( .IN1(n12971), .IN2(n12972), .QN(g20891) );
  NAND2X0 U13909 ( .IN1(n4404), .IN2(n11694), .QN(n12972) );
  OR2X1 U13910 ( .IN1(n11694), .IN2(n7161), .Q(n12971) );
  INVX0 U13911 ( .INP(n12339), .ZN(n11694) );
  NAND2X0 U13912 ( .IN1(n12973), .IN2(g629), .QN(n12339) );
  NOR2X0 U13913 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  NAND2X0 U13914 ( .IN1(n12974), .IN2(n12975), .QN(g20883) );
  NAND2X0 U13915 ( .IN1(n4417), .IN2(n11700), .QN(n12975) );
  OR2X1 U13916 ( .IN1(n11700), .IN2(n7089), .Q(n12974) );
  NAND2X0 U13917 ( .IN1(n12976), .IN2(n12977), .QN(g20882) );
  NAND2X0 U13918 ( .IN1(test_so49), .IN2(n12342), .QN(n12977) );
  NAND2X0 U13919 ( .IN1(n4402), .IN2(n11700), .QN(n12976) );
  INVX0 U13920 ( .INP(n12342), .ZN(n11700) );
  NAND2X0 U13921 ( .IN1(n12964), .IN2(g6979), .QN(n12342) );
  NOR3X0 U13922 ( .IN1(n4489), .IN2(n7004), .IN3(g1345), .QN(n12964) );
  NAND2X0 U13923 ( .IN1(n12978), .IN2(n12979), .QN(g20881) );
  NAND2X0 U13924 ( .IN1(test_so30), .IN2(n12344), .QN(n12979) );
  NAND2X0 U13925 ( .IN1(n4418), .IN2(n11755), .QN(n12978) );
  NAND2X0 U13926 ( .IN1(n12980), .IN2(n12981), .QN(g20880) );
  NAND2X0 U13927 ( .IN1(n11758), .IN2(n4478), .QN(n12981) );
  OR2X1 U13928 ( .IN1(n11758), .IN2(n7121), .Q(n12980) );
  NAND2X0 U13929 ( .IN1(n12982), .IN2(n12983), .QN(g20879) );
  NAND2X0 U13930 ( .IN1(n4404), .IN2(n11755), .QN(n12983) );
  OR2X1 U13931 ( .IN1(n11755), .IN2(n7122), .Q(n12982) );
  INVX0 U13932 ( .INP(n12344), .ZN(n11755) );
  NAND2X0 U13933 ( .IN1(n12973), .IN2(g6911), .QN(n12344) );
  NAND2X0 U13934 ( .IN1(n12984), .IN2(n12985), .QN(g20876) );
  NAND2X0 U13935 ( .IN1(n4418), .IN2(n11758), .QN(n12985) );
  OR2X1 U13936 ( .IN1(n11758), .IN2(n7106), .Q(n12984) );
  NAND2X0 U13937 ( .IN1(n12986), .IN2(n12987), .QN(g20875) );
  NAND2X0 U13938 ( .IN1(n4404), .IN2(n11758), .QN(n12987) );
  OR2X1 U13939 ( .IN1(n11758), .IN2(n7123), .Q(n12986) );
  INVX0 U13940 ( .INP(n12347), .ZN(n11758) );
  NAND2X0 U13941 ( .IN1(n12973), .IN2(g6677), .QN(n12347) );
  NOR3X0 U13942 ( .IN1(n4492), .IN2(n7005), .IN3(g659), .QN(n12973) );
  NAND2X0 U13943 ( .IN1(n12988), .IN2(n12989), .QN(g20874) );
  NAND2X0 U13944 ( .IN1(g2879), .IN2(g8096), .QN(n12989) );
  NAND2X0 U13945 ( .IN1(n4351), .IN2(n12649), .QN(n12988) );
  XOR2X1 U13946 ( .IN1(n7657), .IN2(n12652), .Q(n12649) );
  NOR2X0 U13947 ( .IN1(g3231), .IN2(n13232), .QN(n12652) );
  XOR3X1 U13948 ( .IN1(n12990), .IN2(n12991), .IN3(n12992), .Q(n7657) );
  XOR3X1 U13949 ( .IN1(n7246), .IN2(n7245), .IN3(n12993), .Q(n12992) );
  XOR2X1 U13950 ( .IN1(g2944), .IN2(n7248), .Q(n12993) );
  XOR2X1 U13951 ( .IN1(n7242), .IN2(n7241), .Q(n12991) );
  XOR2X1 U13952 ( .IN1(n7244), .IN2(n7243), .Q(n12990) );
  NOR2X0 U13953 ( .IN1(n10335), .IN2(n12994), .QN(g20789) );
  XOR2X1 U13954 ( .IN1(n4398), .IN2(n12630), .Q(n12994) );
  NOR2X0 U13955 ( .IN1(g2733), .IN2(n4292), .QN(n12630) );
  NOR2X0 U13956 ( .IN1(n4356), .IN2(n7041), .QN(n10335) );
  NOR2X0 U13957 ( .IN1(n10339), .IN2(n12995), .QN(g20752) );
  XOR2X1 U13958 ( .IN1(n4400), .IN2(n12635), .Q(n12995) );
  NOR2X0 U13959 ( .IN1(g2039), .IN2(n4293), .QN(n12635) );
  NOR2X0 U13960 ( .IN1(n4357), .IN2(n7042), .QN(n10339) );
  NOR2X0 U13961 ( .IN1(n10343), .IN2(n12996), .QN(g20717) );
  XNOR2X1 U13962 ( .IN1(n4402), .IN2(n12643), .Q(n12996) );
  NAND2X0 U13963 ( .IN1(n4428), .IN2(g1315), .QN(n12643) );
  NOR2X0 U13964 ( .IN1(n4358), .IN2(n7043), .QN(n10343) );
  NOR2X0 U13965 ( .IN1(n9912), .IN2(n12997), .QN(g20682) );
  XOR2X1 U13966 ( .IN1(n4404), .IN2(n12223), .Q(n12997) );
  NOR2X0 U13967 ( .IN1(g659), .IN2(n4295), .QN(n12223) );
  NOR2X0 U13968 ( .IN1(n4359), .IN2(n7044), .QN(n9912) );
  NAND2X0 U13969 ( .IN1(n12998), .IN2(n12999), .QN(g20417) );
  NAND2X0 U13970 ( .IN1(n4351), .IN2(g2963), .QN(n12999) );
  NAND2X0 U13971 ( .IN1(g2879), .IN2(g7334), .QN(n12998) );
  NAND2X0 U13972 ( .IN1(n13000), .IN2(n13001), .QN(g20376) );
  NAND2X0 U13973 ( .IN1(test_so2), .IN2(n4351), .QN(n13001) );
  NAND2X0 U13974 ( .IN1(g2879), .IN2(g6895), .QN(n13000) );
  NAND2X0 U13975 ( .IN1(n13002), .IN2(n13003), .QN(g20375) );
  NAND2X0 U13976 ( .IN1(n4292), .IN2(g2733), .QN(n13003) );
  NAND2X0 U13977 ( .IN1(n13004), .IN2(g2703), .QN(n13002) );
  NAND2X0 U13978 ( .IN1(n13005), .IN2(n13006), .QN(g20353) );
  NAND2X0 U13979 ( .IN1(n4293), .IN2(g2039), .QN(n13006) );
  NAND2X0 U13980 ( .IN1(n13004), .IN2(g2009), .QN(n13005) );
  NAND2X0 U13981 ( .IN1(n13007), .IN2(n13008), .QN(g20343) );
  NAND2X0 U13982 ( .IN1(n4351), .IN2(g2969), .QN(n13008) );
  NAND2X0 U13983 ( .IN1(g2879), .IN2(g6442), .QN(n13007) );
  NAND2X0 U13984 ( .IN1(n13009), .IN2(n13010), .QN(g20333) );
  NAND2X0 U13985 ( .IN1(n4294), .IN2(g1345), .QN(n13010) );
  NAND2X0 U13986 ( .IN1(n13004), .IN2(g1315), .QN(n13009) );
  NAND2X0 U13987 ( .IN1(n13011), .IN2(n13012), .QN(g20314) );
  NAND2X0 U13988 ( .IN1(n4295), .IN2(g659), .QN(n13012) );
  NAND2X0 U13989 ( .IN1(n13004), .IN2(g629), .QN(n13011) );
  INVX0 U13990 ( .INP(n12294), .ZN(n13004) );
  NAND4X0 U13991 ( .IN1(n6428), .IN2(n7273), .IN3(n6427), .IN4(n13013), .QN(
        n12294) );
  AND2X1 U13992 ( .IN1(n6429), .IN2(n6430), .Q(n13013) );
  NAND2X0 U13993 ( .IN1(n13014), .IN2(n13015), .QN(g20310) );
  NAND2X0 U13994 ( .IN1(n4351), .IN2(g2972), .QN(n13015) );
  NAND2X0 U13995 ( .IN1(g2879), .IN2(g6225), .QN(n13014) );
  NAND2X0 U13996 ( .IN1(n13016), .IN2(n13017), .QN(g19184) );
  NAND2X0 U13997 ( .IN1(n4351), .IN2(g2975), .QN(n13017) );
  NAND2X0 U13998 ( .IN1(g2879), .IN2(g4590), .QN(n13016) );
  NAND2X0 U13999 ( .IN1(n13018), .IN2(n13019), .QN(g19178) );
  NAND2X0 U14000 ( .IN1(n4351), .IN2(g2935), .QN(n13019) );
  NAND2X0 U14001 ( .IN1(test_so5), .IN2(g2879), .QN(n13018) );
  NAND2X0 U14002 ( .IN1(n13020), .IN2(n13021), .QN(g19173) );
  NAND2X0 U14003 ( .IN1(n4351), .IN2(g2978), .QN(n13021) );
  NAND2X0 U14004 ( .IN1(g2879), .IN2(g4323), .QN(n13020) );
  NAND2X0 U14005 ( .IN1(n13022), .IN2(n13023), .QN(g19172) );
  NAND2X0 U14006 ( .IN1(n4351), .IN2(g2953), .QN(n13023) );
  NAND2X0 U14007 ( .IN1(g2879), .IN2(g4321), .QN(n13022) );
  NAND2X0 U14008 ( .IN1(n13024), .IN2(n13025), .QN(g19167) );
  NAND2X0 U14009 ( .IN1(n4351), .IN2(g2938), .QN(n13025) );
  NAND2X0 U14010 ( .IN1(g2879), .IN2(g4200), .QN(n13024) );
  NAND2X0 U14011 ( .IN1(n13026), .IN2(n13027), .QN(g19163) );
  NAND2X0 U14012 ( .IN1(n4351), .IN2(g2981), .QN(n13027) );
  NAND2X0 U14013 ( .IN1(g2879), .IN2(g4090), .QN(n13026) );
  NAND2X0 U14014 ( .IN1(n13028), .IN2(n13029), .QN(g19162) );
  NAND2X0 U14015 ( .IN1(n4351), .IN2(g2956), .QN(n13029) );
  NAND2X0 U14016 ( .IN1(g2879), .IN2(g4088), .QN(n13028) );
  NAND2X0 U14017 ( .IN1(n13030), .IN2(n13031), .QN(g19157) );
  NAND2X0 U14018 ( .IN1(n4351), .IN2(g2941), .QN(n13031) );
  NAND2X0 U14019 ( .IN1(g2879), .IN2(g3993), .QN(n13030) );
  NAND2X0 U14020 ( .IN1(n13032), .IN2(n13033), .QN(g19154) );
  NAND2X0 U14021 ( .IN1(n4351), .IN2(g2874), .QN(n13033) );
  NAND2X0 U14022 ( .IN1(test_so3), .IN2(g2879), .QN(n13032) );
  NAND2X0 U14023 ( .IN1(n13034), .IN2(n13035), .QN(g19153) );
  NAND2X0 U14024 ( .IN1(n4351), .IN2(g2959), .QN(n13035) );
  NAND2X0 U14025 ( .IN1(g2879), .IN2(g8249), .QN(n13034) );
  NAND2X0 U14026 ( .IN1(n13036), .IN2(n13037), .QN(g19149) );
  NAND2X0 U14027 ( .IN1(n4351), .IN2(g2944), .QN(n13037) );
  NAND2X0 U14028 ( .IN1(g2879), .IN2(g8175), .QN(n13036) );
  NAND2X0 U14029 ( .IN1(n13038), .IN2(n13039), .QN(g19144) );
  NAND2X0 U14030 ( .IN1(n4351), .IN2(g2947), .QN(n13039) );
  NAND2X0 U14031 ( .IN1(g2879), .IN2(g8023), .QN(n13038) );
  NAND2X0 U14032 ( .IN1(n13040), .IN2(n13041), .QN(g18975) );
  NAND2X0 U14033 ( .IN1(n4351), .IN2(g2195), .QN(n13041) );
  NAND2X0 U14034 ( .IN1(g2879), .IN2(g2981), .QN(n13040) );
  NAND2X0 U14035 ( .IN1(n13042), .IN2(n13043), .QN(g18968) );
  NAND2X0 U14036 ( .IN1(n4351), .IN2(g2190), .QN(n13043) );
  NAND2X0 U14037 ( .IN1(g2879), .IN2(g2978), .QN(n13042) );
  NAND2X0 U14038 ( .IN1(n13044), .IN2(n13045), .QN(g18957) );
  NAND2X0 U14039 ( .IN1(n4351), .IN2(g2165), .QN(n13045) );
  NAND2X0 U14040 ( .IN1(g2879), .IN2(g2963), .QN(n13044) );
  NAND2X0 U14041 ( .IN1(n13046), .IN2(n13047), .QN(g18942) );
  NAND2X0 U14042 ( .IN1(g2879), .IN2(g2975), .QN(n13047) );
  NAND2X0 U14043 ( .IN1(n4351), .IN2(g2185), .QN(n13046) );
  NAND2X0 U14044 ( .IN1(n13048), .IN2(n13049), .QN(g18907) );
  NAND2X0 U14045 ( .IN1(n4365), .IN2(g3061), .QN(n13049) );
  NAND2X0 U14046 ( .IN1(g2987), .IN2(g2997), .QN(n13048) );
  NAND2X0 U14047 ( .IN1(n13050), .IN2(n13051), .QN(g18906) );
  NAND2X0 U14048 ( .IN1(n4351), .IN2(g2180), .QN(n13051) );
  NAND2X0 U14049 ( .IN1(g2879), .IN2(g2972), .QN(n13050) );
  NAND2X0 U14050 ( .IN1(n13052), .IN2(n13053), .QN(g18885) );
  NAND2X0 U14051 ( .IN1(g2879), .IN2(g2874), .QN(n13053) );
  NAND2X0 U14052 ( .IN1(n4351), .IN2(g2200), .QN(n13052) );
  NAND2X0 U14053 ( .IN1(n13054), .IN2(n13055), .QN(g18883) );
  NAND2X0 U14054 ( .IN1(n4351), .IN2(g1471), .QN(n13055) );
  NAND2X0 U14055 ( .IN1(g2879), .IN2(g2935), .QN(n13054) );
  NAND2X0 U14056 ( .IN1(n13056), .IN2(n13057), .QN(g18868) );
  NAND2X0 U14057 ( .IN1(n4365), .IN2(g3060), .QN(n13057) );
  NAND2X0 U14058 ( .IN1(g2987), .IN2(g3078), .QN(n13056) );
  NAND2X0 U14059 ( .IN1(n13058), .IN2(n13059), .QN(g18867) );
  NAND2X0 U14060 ( .IN1(g2879), .IN2(g2969), .QN(n13059) );
  NAND2X0 U14061 ( .IN1(n4351), .IN2(g2175), .QN(n13058) );
  NAND2X0 U14062 ( .IN1(n13060), .IN2(n13061), .QN(g18866) );
  NAND2X0 U14063 ( .IN1(n4351), .IN2(g1476), .QN(n13061) );
  NAND2X0 U14064 ( .IN1(g2879), .IN2(g2938), .QN(n13060) );
  NAND2X0 U14065 ( .IN1(n13062), .IN2(n13063), .QN(g18852) );
  NAND2X0 U14066 ( .IN1(g2879), .IN2(g2941), .QN(n13063) );
  NAND2X0 U14067 ( .IN1(n4351), .IN2(g1481), .QN(n13062) );
  NAND2X0 U14068 ( .IN1(n13064), .IN2(n13065), .QN(g18837) );
  NAND2X0 U14069 ( .IN1(n4365), .IN2(g3059), .QN(n13065) );
  NAND2X0 U14070 ( .IN1(g2987), .IN2(g3077), .QN(n13064) );
  NAND2X0 U14071 ( .IN1(n13066), .IN2(n13067), .QN(g18836) );
  NAND2X0 U14072 ( .IN1(n4351), .IN2(g2170), .QN(n13067) );
  NAND2X0 U14073 ( .IN1(test_so2), .IN2(g2879), .QN(n13066) );
  NAND2X0 U14074 ( .IN1(n13068), .IN2(n13069), .QN(g18835) );
  OR2X1 U14075 ( .IN1(g2879), .IN2(n4390), .Q(n13069) );
  NAND2X0 U14076 ( .IN1(g2879), .IN2(g2944), .QN(n13068) );
  NAND2X0 U14077 ( .IN1(n13070), .IN2(n13071), .QN(g18821) );
  NAND2X0 U14078 ( .IN1(g2879), .IN2(g2947), .QN(n13071) );
  NAND2X0 U14079 ( .IN1(n4351), .IN2(g1491), .QN(n13070) );
  NAND2X0 U14080 ( .IN1(n13072), .IN2(n13073), .QN(g18820) );
  NAND2X0 U14081 ( .IN1(n4299), .IN2(g2584), .QN(n13073) );
  NAND2X0 U14082 ( .IN1(g2624), .IN2(g2631), .QN(n13072) );
  NAND2X0 U14083 ( .IN1(n13074), .IN2(n13075), .QN(g18804) );
  NAND2X0 U14084 ( .IN1(n4365), .IN2(g3058), .QN(n13075) );
  NAND2X0 U14085 ( .IN1(g2987), .IN2(g3076), .QN(n13074) );
  NAND2X0 U14086 ( .IN1(n13076), .IN2(n13077), .QN(g18803) );
  NAND2X0 U14087 ( .IN1(n4351), .IN2(g1496), .QN(n13077) );
  NAND2X0 U14088 ( .IN1(g2879), .IN2(g2953), .QN(n13076) );
  NAND2X0 U14089 ( .IN1(n13078), .IN2(n13079), .QN(g18794) );
  NAND2X0 U14090 ( .IN1(g1937), .IN2(g1930), .QN(n13079) );
  NAND2X0 U14091 ( .IN1(n4366), .IN2(g1890), .QN(n13078) );
  NAND2X0 U14092 ( .IN1(n13080), .IN2(n13081), .QN(g18782) );
  NAND2X0 U14093 ( .IN1(g3109), .IN2(g559), .QN(n13081) );
  OR2X1 U14094 ( .IN1(g3109), .IN2(n4445), .Q(n13080) );
  NAND2X0 U14095 ( .IN1(n13082), .IN2(n13083), .QN(g18781) );
  NAND2X0 U14096 ( .IN1(n4351), .IN2(g1501), .QN(n13083) );
  NAND2X0 U14097 ( .IN1(g2879), .IN2(g2956), .QN(n13082) );
  NAND2X0 U14098 ( .IN1(n13084), .IN2(n13085), .QN(g18780) );
  NAND2X0 U14099 ( .IN1(n4299), .IN2(g2631), .QN(n13085) );
  NAND2X0 U14100 ( .IN1(n7233), .IN2(g2624), .QN(n13084) );
  NAND2X0 U14101 ( .IN1(n13086), .IN2(n13087), .QN(g18763) );
  NAND2X0 U14102 ( .IN1(n4300), .IN2(g1196), .QN(n13087) );
  NAND2X0 U14103 ( .IN1(g1236), .IN2(g1243), .QN(n13086) );
  NAND2X0 U14104 ( .IN1(n13088), .IN2(n13089), .QN(g18755) );
  NAND2X0 U14105 ( .IN1(n4365), .IN2(g3057), .QN(n13089) );
  NAND2X0 U14106 ( .IN1(g2987), .IN2(g3075), .QN(n13088) );
  NAND2X0 U14107 ( .IN1(n13090), .IN2(n13091), .QN(g18754) );
  NAND2X0 U14108 ( .IN1(g2879), .IN2(g2959), .QN(n13091) );
  NAND2X0 U14109 ( .IN1(n4351), .IN2(g1506), .QN(n13090) );
  NAND2X0 U14110 ( .IN1(n13092), .IN2(n13093), .QN(g18743) );
  NAND2X0 U14111 ( .IN1(n7234), .IN2(g1930), .QN(n13093) );
  NAND2X0 U14112 ( .IN1(n4366), .IN2(g1937), .QN(n13092) );
  NAND2X0 U14113 ( .IN1(n13094), .IN2(n13095), .QN(g18726) );
  NAND2X0 U14114 ( .IN1(n4313), .IN2(test_so22), .QN(n13095) );
  NAND2X0 U14115 ( .IN1(g550), .IN2(g557), .QN(n13094) );
  NAND2X0 U14116 ( .IN1(n13096), .IN2(n13097), .QN(g18719) );
  NAND2X0 U14117 ( .IN1(n4383), .IN2(g3211), .QN(n13097) );
  NAND2X0 U14118 ( .IN1(g8030), .IN2(g559), .QN(n13096) );
  NAND2X0 U14119 ( .IN1(n13098), .IN2(n13099), .QN(g18707) );
  NAND2X0 U14120 ( .IN1(n4300), .IN2(g1243), .QN(n13099) );
  NAND2X0 U14121 ( .IN1(n7235), .IN2(g1236), .QN(n13098) );
  NAND2X0 U14122 ( .IN1(n13100), .IN2(n13101), .QN(g18678) );
  NAND2X0 U14123 ( .IN1(n4313), .IN2(g557), .QN(n13101) );
  NAND2X0 U14124 ( .IN1(n7236), .IN2(g550), .QN(n13100) );
  NAND2X0 U14125 ( .IN1(n13102), .IN2(n13103), .QN(g18669) );
  NAND2X0 U14126 ( .IN1(n4382), .IN2(test_so6), .QN(n13103) );
  NAND2X0 U14127 ( .IN1(g8106), .IN2(g559), .QN(n13102) );
  NAND2X0 U14128 ( .IN1(n13104), .IN2(n13105), .QN(g17429) );
  NAND2X0 U14129 ( .IN1(g3109), .IN2(g2574), .QN(n13105) );
  NAND2X0 U14130 ( .IN1(n4494), .IN2(g3088), .QN(n13104) );
  NAND2X0 U14131 ( .IN1(n13106), .IN2(n13107), .QN(g17383) );
  NAND2X0 U14132 ( .IN1(n4494), .IN2(test_so8), .QN(n13107) );
  NAND2X0 U14133 ( .IN1(g3109), .IN2(g1880), .QN(n13106) );
  NAND2X0 U14134 ( .IN1(n13108), .IN2(n13109), .QN(g17341) );
  NAND2X0 U14135 ( .IN1(n4383), .IN2(g3185), .QN(n13109) );
  NAND2X0 U14136 ( .IN1(g8030), .IN2(g2574), .QN(n13108) );
  NAND2X0 U14137 ( .IN1(n13110), .IN2(n13111), .QN(g17340) );
  NAND2X0 U14138 ( .IN1(g3109), .IN2(g1186), .QN(n13111) );
  OR2X1 U14139 ( .IN1(g3109), .IN2(n4441), .Q(n13110) );
  NAND2X0 U14140 ( .IN1(n13112), .IN2(n13113), .QN(g17303) );
  OR2X1 U14141 ( .IN1(g8030), .IN2(n4450), .Q(n13113) );
  NAND2X0 U14142 ( .IN1(g8030), .IN2(g1880), .QN(n13112) );
  NAND2X0 U14143 ( .IN1(n13114), .IN2(n13115), .QN(g17302) );
  NAND2X0 U14144 ( .IN1(g3109), .IN2(g499), .QN(n13115) );
  OR2X1 U14145 ( .IN1(g3109), .IN2(n4444), .Q(n13114) );
  NAND2X0 U14146 ( .IN1(n13116), .IN2(n13117), .QN(g17271) );
  NAND2X0 U14147 ( .IN1(n4382), .IN2(g3182), .QN(n13117) );
  NAND2X0 U14148 ( .IN1(g8106), .IN2(g2574), .QN(n13116) );
  NAND2X0 U14149 ( .IN1(n13118), .IN2(n13119), .QN(g17270) );
  NAND2X0 U14150 ( .IN1(g8030), .IN2(g1186), .QN(n13119) );
  NAND2X0 U14151 ( .IN1(n4383), .IN2(g3167), .QN(n13118) );
  NAND2X0 U14152 ( .IN1(n13120), .IN2(n13121), .QN(g17269) );
  NAND2X0 U14153 ( .IN1(g3109), .IN2(g2633), .QN(n13121) );
  NAND2X0 U14154 ( .IN1(n4494), .IN2(g3096), .QN(n13120) );
  NAND2X0 U14155 ( .IN1(n13122), .IN2(n13123), .QN(g17248) );
  NAND2X0 U14156 ( .IN1(g8106), .IN2(g1880), .QN(n13123) );
  OR2X1 U14157 ( .IN1(g8106), .IN2(n4338), .Q(n13122) );
  NAND2X0 U14158 ( .IN1(n13124), .IN2(n13125), .QN(g17247) );
  NAND2X0 U14159 ( .IN1(n4383), .IN2(g3158), .QN(n13125) );
  NAND2X0 U14160 ( .IN1(g8030), .IN2(g499), .QN(n13124) );
  NAND2X0 U14161 ( .IN1(n13126), .IN2(n13127), .QN(g17246) );
  NAND2X0 U14162 ( .IN1(g3109), .IN2(g1939), .QN(n13127) );
  NAND2X0 U14163 ( .IN1(n4494), .IN2(g3093), .QN(n13126) );
  NAND2X0 U14164 ( .IN1(n13128), .IN2(n13129), .QN(g17236) );
  NAND2X0 U14165 ( .IN1(g8106), .IN2(g1186), .QN(n13129) );
  NAND2X0 U14166 ( .IN1(n4382), .IN2(g3164), .QN(n13128) );
  NAND2X0 U14167 ( .IN1(n13130), .IN2(n13131), .QN(g17235) );
  NAND2X0 U14168 ( .IN1(n4383), .IN2(g3095), .QN(n13131) );
  NAND2X0 U14169 ( .IN1(g8030), .IN2(g2633), .QN(n13130) );
  NAND2X0 U14170 ( .IN1(n13132), .IN2(n13133), .QN(g17234) );
  NAND2X0 U14171 ( .IN1(g3109), .IN2(g1245), .QN(n13133) );
  OR2X1 U14172 ( .IN1(g3109), .IN2(n4344), .Q(n13132) );
  NAND2X0 U14173 ( .IN1(n13134), .IN2(n13135), .QN(g17229) );
  NAND2X0 U14174 ( .IN1(n4382), .IN2(g3155), .QN(n13135) );
  NAND2X0 U14175 ( .IN1(g8106), .IN2(g499), .QN(n13134) );
  NAND2X0 U14176 ( .IN1(n13136), .IN2(n13137), .QN(g17228) );
  OR2X1 U14177 ( .IN1(g8030), .IN2(n4451), .Q(n13137) );
  NAND2X0 U14178 ( .IN1(g8030), .IN2(g1939), .QN(n13136) );
  NAND2X0 U14179 ( .IN1(n13138), .IN2(n13139), .QN(g17226) );
  NAND2X0 U14180 ( .IN1(n4382), .IN2(g3094), .QN(n13139) );
  NAND2X0 U14181 ( .IN1(g8106), .IN2(g2633), .QN(n13138) );
  NAND2X0 U14182 ( .IN1(n13140), .IN2(n13141), .QN(g17225) );
  NAND2X0 U14183 ( .IN1(g8030), .IN2(g1245), .QN(n13141) );
  NAND2X0 U14184 ( .IN1(n4383), .IN2(g3086), .QN(n13140) );
  NAND2X0 U14185 ( .IN1(n13142), .IN2(n13143), .QN(g17224) );
  OR2X1 U14186 ( .IN1(g8106), .IN2(n4448), .Q(n13143) );
  NAND2X0 U14187 ( .IN1(g8106), .IN2(g1939), .QN(n13142) );
  NAND2X0 U14188 ( .IN1(n13144), .IN2(n13145), .QN(g17222) );
  NAND2X0 U14189 ( .IN1(g8106), .IN2(g1245), .QN(n13145) );
  NAND2X0 U14190 ( .IN1(n4382), .IN2(g3085), .QN(n13144) );
  NAND2X0 U14191 ( .IN1(n13146), .IN2(n13147), .QN(g16880) );
  NAND2X0 U14192 ( .IN1(n4365), .IN2(g3056), .QN(n13147) );
  NAND2X0 U14193 ( .IN1(g2987), .IN2(g3074), .QN(n13146) );
  NAND2X0 U14194 ( .IN1(n13148), .IN2(n13149), .QN(g16866) );
  NAND2X0 U14195 ( .IN1(n4365), .IN2(g3051), .QN(n13149) );
  NAND2X0 U14196 ( .IN1(test_so97), .IN2(g2987), .QN(n13148) );
  NAND2X0 U14197 ( .IN1(n13150), .IN2(n13151), .QN(g16861) );
  NAND2X0 U14198 ( .IN1(test_so96), .IN2(n4365), .QN(n13151) );
  NAND2X0 U14199 ( .IN1(g2987), .IN2(g3073), .QN(n13150) );
  NAND2X0 U14200 ( .IN1(n13152), .IN2(n13153), .QN(g16860) );
  NAND2X0 U14201 ( .IN1(n4365), .IN2(g3046), .QN(n13153) );
  NAND2X0 U14202 ( .IN1(g2987), .IN2(g3065), .QN(n13152) );
  NAND2X0 U14203 ( .IN1(n13154), .IN2(n13155), .QN(g16857) );
  NAND2X0 U14204 ( .IN1(n4365), .IN2(g3050), .QN(n13155) );
  NAND2X0 U14205 ( .IN1(g2987), .IN2(g3069), .QN(n13154) );
  NAND2X0 U14206 ( .IN1(n13156), .IN2(n13157), .QN(g16854) );
  NAND2X0 U14207 ( .IN1(n4365), .IN2(g3053), .QN(n13157) );
  NAND2X0 U14208 ( .IN1(g2987), .IN2(g3072), .QN(n13156) );
  NAND2X0 U14209 ( .IN1(n13158), .IN2(n13159), .QN(g16853) );
  NAND2X0 U14210 ( .IN1(n4365), .IN2(g3045), .QN(n13159) );
  NAND2X0 U14211 ( .IN1(g2987), .IN2(g3064), .QN(n13158) );
  NAND2X0 U14212 ( .IN1(n13160), .IN2(n13161), .QN(g16851) );
  NAND2X0 U14213 ( .IN1(n4365), .IN2(g3049), .QN(n13161) );
  NAND2X0 U14214 ( .IN1(g2987), .IN2(g3068), .QN(n13160) );
  NAND2X0 U14215 ( .IN1(n13162), .IN2(n13163), .QN(g16845) );
  NAND2X0 U14216 ( .IN1(n4365), .IN2(g3052), .QN(n13163) );
  NAND2X0 U14217 ( .IN1(g2987), .IN2(g3071), .QN(n13162) );
  NAND2X0 U14218 ( .IN1(n13164), .IN2(n13165), .QN(g16844) );
  NAND2X0 U14219 ( .IN1(n4365), .IN2(g3044), .QN(n13165) );
  NAND2X0 U14220 ( .IN1(g2987), .IN2(g3063), .QN(n13164) );
  NAND2X0 U14221 ( .IN1(n13166), .IN2(n13167), .QN(g16835) );
  NAND2X0 U14222 ( .IN1(n4365), .IN2(g3048), .QN(n13167) );
  NAND2X0 U14223 ( .IN1(g2987), .IN2(g3067), .QN(n13166) );
  NAND2X0 U14224 ( .IN1(n13168), .IN2(n13169), .QN(g16824) );
  NAND2X0 U14225 ( .IN1(n4365), .IN2(g3043), .QN(n13169) );
  NAND2X0 U14226 ( .IN1(g2987), .IN2(g3062), .QN(n13168) );
  NOR2X0 U14227 ( .IN1(g51), .IN2(DFF_1_n1), .QN(g16823) );
  NAND2X0 U14228 ( .IN1(n13170), .IN2(n13171), .QN(g16803) );
  NAND2X0 U14229 ( .IN1(n4365), .IN2(g3047), .QN(n13171) );
  NAND2X0 U14230 ( .IN1(g2987), .IN2(g3066), .QN(n13170) );
  NOR2X0 U14231 ( .IN1(n4423), .IN2(g51), .QN(g16802) );
  NAND2X0 U14232 ( .IN1(n13172), .IN2(n13173), .QN(g16718) );
  OR2X1 U14233 ( .IN1(g2703), .IN2(n7041), .Q(n13173) );
  NAND2X0 U14234 ( .IN1(g2703), .IN2(g2584), .QN(n13172) );
  NAND2X0 U14235 ( .IN1(n13174), .IN2(n13175), .QN(g16692) );
  OR2X1 U14236 ( .IN1(g2009), .IN2(n7042), .Q(n13175) );
  NAND2X0 U14237 ( .IN1(g2009), .IN2(g1890), .QN(n13174) );
  NAND2X0 U14238 ( .IN1(n13176), .IN2(n13177), .QN(g16671) );
  OR2X1 U14239 ( .IN1(g1315), .IN2(n7043), .Q(n13177) );
  NAND2X0 U14240 ( .IN1(g1315), .IN2(g1196), .QN(n13176) );
  NAND2X0 U14241 ( .IN1(n13178), .IN2(n13179), .QN(g16654) );
  OR2X1 U14242 ( .IN1(g629), .IN2(n7044), .Q(n13179) );
  NAND2X0 U14243 ( .IN1(test_so22), .IN2(g629), .QN(n13178) );
  NAND2X0 U14244 ( .IN1(n13180), .IN2(g2987), .QN(g16496) );
  NAND2X0 U14245 ( .IN1(DFF_1612_n1), .IN2(g5388), .QN(n13180) );
  NOR3X0 U14246 ( .IN1(n13181), .IN2(n13182), .IN3(n13183), .QN(g13194) );
  NOR2X0 U14247 ( .IN1(n4314), .IN2(test_so87), .QN(n13183) );
  NOR2X0 U14248 ( .IN1(n4370), .IN2(g2561), .QN(n13182) );
  NOR2X0 U14249 ( .IN1(n4299), .IN2(g2562), .QN(n13181) );
  NOR3X0 U14250 ( .IN1(n13184), .IN2(n13185), .IN3(n13186), .QN(g13182) );
  NOR2X0 U14251 ( .IN1(n4366), .IN2(g1868), .QN(n13186) );
  NOR2X0 U14252 ( .IN1(n4296), .IN2(g1869), .QN(n13185) );
  NOR2X0 U14253 ( .IN1(n4315), .IN2(g1867), .QN(n13184) );
  NOR3X0 U14254 ( .IN1(n13187), .IN2(n13188), .IN3(n13189), .QN(g13175) );
  NOR2X0 U14255 ( .IN1(n4299), .IN2(g2553), .QN(n13189) );
  NOR2X0 U14256 ( .IN1(n4314), .IN2(g2554), .QN(n13188) );
  NOR2X0 U14257 ( .IN1(n4370), .IN2(g2552), .QN(n13187) );
  NOR3X0 U14258 ( .IN1(n13190), .IN2(n13191), .IN3(n13192), .QN(g13171) );
  NOR2X0 U14259 ( .IN1(n4300), .IN2(test_so44), .QN(n13192) );
  NOR2X0 U14260 ( .IN1(n4316), .IN2(g1173), .QN(n13191) );
  NOR2X0 U14261 ( .IN1(n4371), .IN2(g1175), .QN(n13190) );
  NOR3X0 U14262 ( .IN1(n13193), .IN2(n13194), .IN3(n13195), .QN(g13164) );
  NOR2X0 U14263 ( .IN1(n4366), .IN2(g1859), .QN(n13195) );
  NOR2X0 U14264 ( .IN1(n4296), .IN2(g1860), .QN(n13194) );
  NOR2X0 U14265 ( .IN1(n4315), .IN2(g1858), .QN(n13193) );
  NOR3X0 U14266 ( .IN1(n13196), .IN2(n13197), .IN3(n13198), .QN(g13160) );
  NOR2X0 U14267 ( .IN1(n4313), .IN2(g487), .QN(n13198) );
  NOR2X0 U14268 ( .IN1(n4298), .IN2(g488), .QN(n13197) );
  NOR2X0 U14269 ( .IN1(n4372), .IN2(g486), .QN(n13196) );
  NOR3X0 U14270 ( .IN1(n13199), .IN2(n13200), .IN3(n13201), .QN(g13155) );
  NOR2X0 U14271 ( .IN1(n4300), .IN2(g1165), .QN(n13201) );
  NOR2X0 U14272 ( .IN1(n4371), .IN2(g1166), .QN(n13200) );
  NOR2X0 U14273 ( .IN1(n4316), .IN2(g1164), .QN(n13199) );
  NOR3X0 U14274 ( .IN1(n13202), .IN2(n13203), .IN3(n13204), .QN(g13149) );
  NOR2X0 U14275 ( .IN1(n4313), .IN2(g478), .QN(n13204) );
  NOR2X0 U14276 ( .IN1(n4298), .IN2(g479), .QN(n13203) );
  NOR2X0 U14277 ( .IN1(n4372), .IN2(g477), .QN(n13202) );
  NOR3X0 U14278 ( .IN1(n13205), .IN2(n13206), .IN3(n13207), .QN(g13143) );
  NOR2X0 U14279 ( .IN1(n4299), .IN2(g2559), .QN(n13207) );
  NOR2X0 U14280 ( .IN1(n4314), .IN2(g2539), .QN(n13206) );
  NOR2X0 U14281 ( .IN1(n4370), .IN2(g2555), .QN(n13205) );
  NOR3X0 U14282 ( .IN1(n13208), .IN2(n13209), .IN3(n13210), .QN(g13135) );
  NOR2X0 U14283 ( .IN1(n4366), .IN2(g1865), .QN(n13210) );
  NOR2X0 U14284 ( .IN1(n4296), .IN2(g1845), .QN(n13209) );
  NOR2X0 U14285 ( .IN1(n4315), .IN2(g1861), .QN(n13208) );
  NOR3X0 U14286 ( .IN1(n13211), .IN2(n13212), .IN3(n13213), .QN(g13124) );
  NOR2X0 U14287 ( .IN1(n4300), .IN2(g1171), .QN(n13213) );
  NOR2X0 U14288 ( .IN1(n4371), .IN2(g1151), .QN(n13212) );
  NOR2X0 U14289 ( .IN1(n4316), .IN2(g1167), .QN(n13211) );
  NOR3X0 U14290 ( .IN1(n13214), .IN2(n13215), .IN3(n13216), .QN(g13111) );
  NOR2X0 U14291 ( .IN1(n4313), .IN2(g484), .QN(n13216) );
  NOR2X0 U14292 ( .IN1(n4298), .IN2(g464), .QN(n13215) );
  NOR2X0 U14293 ( .IN1(n4372), .IN2(g480), .QN(n13214) );
  AND4X1 U14294 ( .IN1(n6995), .IN2(n10780), .IN3(n7049), .IN4(n13217), .Q(
        g13110) );
  NOR4X0 U14295 ( .IN1(n4349), .IN2(n4330), .IN3(g2912), .IN4(g2917), .QN(
        n13217) );
  INVX0 U14296 ( .INP(n7678), .ZN(n10780) );
  NAND4X0 U14297 ( .IN1(n7048), .IN2(n4431), .IN3(n13218), .IN4(n4355), .QN(
        n7678) );
  AND2X1 U14298 ( .IN1(n4291), .IN2(n4305), .Q(n13218) );
  XOR2X1 U14299 ( .IN1(n7261), .IN2(n7829), .Q(N995) );
  XNOR3X1 U14300 ( .IN1(n13219), .IN2(n13220), .IN3(n13221), .Q(n7829) );
  XOR3X1 U14301 ( .IN1(n13236), .IN2(n13237), .IN3(n13222), .Q(n13221) );
  XOR2X1 U14302 ( .IN1(g8275), .IN2(test_so99), .Q(n13222) );
  XOR2X1 U14303 ( .IN1(n7257), .IN2(n7256), .Q(n13220) );
  XOR2X1 U14304 ( .IN1(n13238), .IN2(n7258), .Q(n13219) );
  XOR2X1 U14305 ( .IN1(n7832), .IN2(n7259), .Q(N690) );
  XOR3X1 U14306 ( .IN1(n13223), .IN2(n13224), .IN3(n13225), .Q(n7832) );
  XOR3X1 U14307 ( .IN1(n13240), .IN2(n13241), .IN3(n13226), .Q(n13225) );
  XOR2X1 U14308 ( .IN1(g8262), .IN2(n13239), .Q(n13226) );
  XOR2X1 U14309 ( .IN1(n7238), .IN2(n7237), .Q(n13224) );
  XOR2X1 U14310 ( .IN1(n7240), .IN2(n7239), .Q(n13223) );
  OR2X1 U3772_U1 ( .IN1(n2230), .IN2(n2217), .Q(n2231) );
  OR2X1 U3776_U1 ( .IN1(n2374), .IN2(n2361), .Q(n2375) );
  OR2X1 U3777_U1 ( .IN1(g51), .IN2(DFF_2_n1), .Q(n4264) );
  OR2X1 U3778_U1 ( .IN1(n2445), .IN2(n2446), .Q(n2440) );
  OR2X1 U3779_U1 ( .IN1(n2478), .IN2(n2446), .Q(n2426) );
  OR2X1 U3780_U1 ( .IN1(n2670), .IN2(n2671), .Q(n2669) );
  OR2X1 U3781_U1 ( .IN1(n2685), .IN2(n2686), .Q(n2684) );
  OR2X1 U3782_U1 ( .IN1(n2718), .IN2(n2719), .Q(n2717) );
  OR2X1 U3783_U1 ( .IN1(n2982), .IN2(g2124), .Q(n2981) );
  OR2X1 U3784_U1 ( .IN1(n2985), .IN2(g1430), .Q(n2984) );
  OR2X1 U3785_U1 ( .IN1(n2988), .IN2(g744), .Q(n2987) );
  OR2X1 U3786_U1 ( .IN1(n2991), .IN2(g56), .Q(n2990) );
  OR2X1 U3787_U1 ( .IN1(n3742), .IN2(test_so98), .Q(n3741) );
  OR2X1 U3901_U1 ( .IN1(n2302), .IN2(n2289), .Q(n2303) );
  OR2X1 U3902_U1 ( .IN1(n2313), .IN2(n2289), .Q(n2275) );
  INVX0 U4467_U2 ( .INP(n3253), .ZN(U4467_n1) );
  NOR2X0 U4467_U1 ( .IN1(n3254), .IN2(U4467_n1), .QN(n3252) );
  INVX0 U4904_U2 ( .INP(n2800), .ZN(U4904_n1) );
  NOR2X0 U4904_U1 ( .IN1(n63), .IN2(U4904_n1), .QN(n2798) );
  INVX0 U4930_U2 ( .INP(n2616), .ZN(U4930_n1) );
  NOR2X0 U4930_U1 ( .IN1(n63), .IN2(U4930_n1), .QN(n2594) );
  INVX0 U5128_U2 ( .INP(n3933), .ZN(U5128_n1) );
  NOR2X0 U5128_U1 ( .IN1(n4406), .IN2(U5128_n1), .QN(n3940) );
  INVX0 U5141_U2 ( .INP(n3939), .ZN(U5141_n1) );
  NOR2X0 U5141_U1 ( .IN1(n4405), .IN2(U5141_n1), .QN(n3936) );
  INVX0 U5749_U2 ( .INP(g2133), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3160), .IN2(U5749_n1), .QN(n3159) );
  INVX0 U5750_U2 ( .INP(g1439), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3164), .IN2(U5750_n1), .QN(n3163) );
  INVX0 U5751_U2 ( .INP(g753), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3168), .IN2(U5751_n1), .QN(n3167) );
  INVX0 U5752_U2 ( .INP(g65), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3172), .IN2(U5752_n1), .QN(n3171) );
  INVX0 U5753_U2 ( .INP(g2142), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4522), .IN2(U5753_n1), .QN(n3424) );
  INVX0 U5754_U2 ( .INP(g2151), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4526), .IN2(U5754_n1), .QN(n3683) );
  INVX0 U5755_U2 ( .INP(g2160), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3888), .IN2(U5755_n1), .QN(n3887) );
  INVX0 U5756_U2 ( .INP(g1448), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4523), .IN2(U5756_n1), .QN(n3427) );
  INVX0 U5757_U2 ( .INP(g1457), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(n3686) );
  INVX0 U5758_U2 ( .INP(g1466), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3891), .IN2(U5758_n1), .QN(n3890) );
  INVX0 U5759_U2 ( .INP(g762), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3431), .IN2(U5759_n1), .QN(n3430) );
  INVX0 U5760_U2 ( .INP(g771), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3690), .IN2(U5760_n1), .QN(n3689) );
  INVX0 U5761_U2 ( .INP(g780), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3894), .IN2(U5761_n1), .QN(n3893) );
  INVX0 U5762_U2 ( .INP(g74), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4521), .IN2(U5762_n1), .QN(n3433) );
  INVX0 U5763_U2 ( .INP(g83), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(n3692) );
  INVX0 U5764_U2 ( .INP(g92), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3897), .IN2(U5764_n1), .QN(n3896) );
  INVX0 U5882_U2 ( .INP(n4102), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(g3036), .IN2(U5882_n1), .QN(n4101) );
  INVX0 U5939_U2 ( .INP(g2257), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n673), .IN2(U5939_n1), .QN(n3038) );
  INVX0 U5940_U2 ( .INP(g1563), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n509), .IN2(U5940_n1), .QN(n3070) );
  INVX0 U5941_U2 ( .INP(g869), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n335), .IN2(U5941_n1), .QN(n3102) );
  INVX0 U5942_U2 ( .INP(g181), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n167), .IN2(U5942_n1), .QN(n3130) );
  INVX0 U6140_U2 ( .INP(g3002), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4066), .IN2(U6140_n1), .QN(n4065) );
  INVX0 U6460_U2 ( .INP(g3233), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(g3230), .IN2(U6460_n1), .QN(n3700) );
  INVX0 U6470_U2 ( .INP(g2892), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4305), .IN2(U6470_n1), .QN(n4182) );
  INVX0 U6562_U2 ( .INP(n3938), .ZN(U6562_n1) );
  NOR2X0 U6562_U1 ( .IN1(g3204), .IN2(U6562_n1), .QN(n3939) );
  INVX0 U6563_U2 ( .INP(n4073), .ZN(U6563_n1) );
  NOR2X0 U6563_U1 ( .IN1(g3204), .IN2(U6563_n1), .QN(n3705) );
  INVX0 U6718_U2 ( .INP(n3944), .ZN(U6718_n1) );
  NOR2X0 U6718_U1 ( .IN1(g3197), .IN2(U6718_n1), .QN(n4073) );
  INVX0 U7116_U2 ( .INP(n4058), .ZN(U7116_n1) );
  NOR2X0 U7116_U1 ( .IN1(g2903), .IN2(U7116_n1), .QN(n4057) );
  INVX0 U7118_U2 ( .INP(n4123), .ZN(U7118_n1) );
  NOR2X0 U7118_U1 ( .IN1(g2896), .IN2(U7118_n1), .QN(n4122) );
  INVX0 U7293_U2 ( .INP(n4598), .ZN(U7293_n1) );
  NOR2X0 U7293_U1 ( .IN1(g3234), .IN2(U7293_n1), .QN(g20877) );
endmodule

