module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n504_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n830_, new_n480_, new_n625_, new_n730_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n837_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_20 );
not g001 ( new_n107_, keyIn_0_5 );
not g002 ( new_n108_, N85 );
and g003 ( new_n109_, new_n108_, N81 );
not g004 ( new_n110_, N81 );
and g005 ( new_n111_, new_n110_, N85 );
or g006 ( new_n112_, new_n109_, new_n111_ );
not g007 ( new_n113_, new_n112_ );
and g008 ( new_n114_, N89, N93 );
not g009 ( new_n115_, new_n114_ );
or g010 ( new_n116_, N89, N93 );
and g011 ( new_n117_, new_n115_, new_n116_ );
or g012 ( new_n118_, new_n113_, new_n117_ );
and g013 ( new_n119_, new_n113_, new_n117_ );
not g014 ( new_n120_, new_n119_ );
and g015 ( new_n121_, new_n120_, new_n118_ );
not g016 ( new_n122_, new_n121_ );
and g017 ( new_n123_, new_n122_, new_n107_ );
and g018 ( new_n124_, new_n121_, keyIn_0_5 );
or g019 ( new_n125_, new_n123_, new_n124_ );
not g020 ( new_n126_, keyIn_0_4 );
and g021 ( new_n127_, N73, N77 );
not g022 ( new_n128_, N73 );
not g023 ( new_n129_, N77 );
and g024 ( new_n130_, new_n128_, new_n129_ );
or g025 ( new_n131_, new_n130_, new_n127_ );
and g026 ( new_n132_, N65, N69 );
not g027 ( new_n133_, N65 );
not g028 ( new_n134_, N69 );
and g029 ( new_n135_, new_n133_, new_n134_ );
or g030 ( new_n136_, new_n135_, new_n132_ );
and g031 ( new_n137_, new_n131_, new_n136_ );
not g032 ( new_n138_, new_n137_ );
or g033 ( new_n139_, new_n131_, new_n136_ );
and g034 ( new_n140_, new_n138_, new_n139_ );
and g035 ( new_n141_, new_n140_, new_n126_ );
not g036 ( new_n142_, new_n140_ );
and g037 ( new_n143_, new_n142_, keyIn_0_4 );
or g038 ( new_n144_, new_n143_, new_n141_ );
and g039 ( new_n145_, new_n125_, new_n144_ );
not g040 ( new_n146_, new_n125_ );
not g041 ( new_n147_, new_n141_ );
or g042 ( new_n148_, new_n140_, new_n126_ );
and g043 ( new_n149_, new_n147_, new_n148_ );
and g044 ( new_n150_, new_n146_, new_n149_ );
or g045 ( new_n151_, new_n150_, new_n145_ );
and g046 ( new_n152_, new_n151_, new_n106_ );
not g047 ( new_n153_, new_n145_ );
or g048 ( new_n154_, new_n125_, new_n144_ );
and g049 ( new_n155_, new_n153_, new_n154_ );
and g050 ( new_n156_, new_n155_, keyIn_0_20 );
or g051 ( new_n157_, new_n152_, new_n156_ );
and g052 ( new_n158_, N129, N137 );
and g053 ( new_n159_, new_n157_, new_n158_ );
or g054 ( new_n160_, new_n155_, keyIn_0_20 );
or g055 ( new_n161_, new_n151_, new_n106_ );
and g056 ( new_n162_, new_n161_, new_n160_ );
not g057 ( new_n163_, new_n158_ );
and g058 ( new_n164_, new_n162_, new_n163_ );
or g059 ( new_n165_, new_n159_, new_n164_ );
and g060 ( new_n166_, new_n165_, keyIn_0_24 );
not g061 ( new_n167_, keyIn_0_24 );
or g062 ( new_n168_, new_n162_, new_n163_ );
or g063 ( new_n169_, new_n157_, new_n158_ );
and g064 ( new_n170_, new_n169_, new_n168_ );
and g065 ( new_n171_, new_n170_, new_n167_ );
or g066 ( new_n172_, new_n166_, new_n171_ );
not g067 ( new_n173_, N17 );
and g068 ( new_n174_, new_n173_, N1 );
not g069 ( new_n175_, N1 );
and g070 ( new_n176_, new_n175_, N17 );
or g071 ( new_n177_, new_n174_, new_n176_ );
and g072 ( new_n178_, N33, N49 );
not g073 ( new_n179_, N33 );
not g074 ( new_n180_, N49 );
and g075 ( new_n181_, new_n179_, new_n180_ );
or g076 ( new_n182_, new_n181_, new_n178_ );
and g077 ( new_n183_, new_n177_, new_n182_ );
not g078 ( new_n184_, new_n183_ );
or g079 ( new_n185_, new_n177_, new_n182_ );
and g080 ( new_n186_, new_n184_, new_n185_ );
not g081 ( new_n187_, new_n186_ );
and g082 ( new_n188_, new_n187_, keyIn_0_8 );
not g083 ( new_n189_, new_n188_ );
or g084 ( new_n190_, new_n187_, keyIn_0_8 );
and g085 ( new_n191_, new_n189_, new_n190_ );
and g086 ( new_n192_, new_n172_, new_n191_ );
or g087 ( new_n193_, new_n170_, new_n167_ );
or g088 ( new_n194_, new_n165_, keyIn_0_24 );
and g089 ( new_n195_, new_n194_, new_n193_ );
not g090 ( new_n196_, new_n191_ );
and g091 ( new_n197_, new_n195_, new_n196_ );
or g092 ( new_n198_, new_n192_, new_n197_ );
not g093 ( new_n199_, keyIn_0_21 );
not g094 ( new_n200_, keyIn_0_7 );
and g095 ( new_n201_, N113, N117 );
not g096 ( new_n202_, N113 );
not g097 ( new_n203_, N117 );
and g098 ( new_n204_, new_n202_, new_n203_ );
or g099 ( new_n205_, new_n204_, new_n201_ );
and g100 ( new_n206_, N121, N125 );
not g101 ( new_n207_, N121 );
not g102 ( new_n208_, N125 );
and g103 ( new_n209_, new_n207_, new_n208_ );
or g104 ( new_n210_, new_n209_, new_n206_ );
and g105 ( new_n211_, new_n205_, new_n210_ );
not g106 ( new_n212_, new_n211_ );
or g107 ( new_n213_, new_n205_, new_n210_ );
and g108 ( new_n214_, new_n212_, new_n213_ );
and g109 ( new_n215_, new_n214_, new_n200_ );
not g110 ( new_n216_, new_n215_ );
or g111 ( new_n217_, new_n214_, new_n200_ );
and g112 ( new_n218_, new_n216_, new_n217_ );
and g113 ( new_n219_, N105, N109 );
not g114 ( new_n220_, N105 );
not g115 ( new_n221_, N109 );
and g116 ( new_n222_, new_n220_, new_n221_ );
or g117 ( new_n223_, new_n222_, new_n219_ );
and g118 ( new_n224_, N97, N101 );
not g119 ( new_n225_, N97 );
not g120 ( new_n226_, N101 );
and g121 ( new_n227_, new_n225_, new_n226_ );
or g122 ( new_n228_, new_n227_, new_n224_ );
and g123 ( new_n229_, new_n223_, new_n228_ );
not g124 ( new_n230_, new_n229_ );
or g125 ( new_n231_, new_n223_, new_n228_ );
and g126 ( new_n232_, new_n230_, new_n231_ );
or g127 ( new_n233_, new_n232_, keyIn_0_6 );
and g128 ( new_n234_, new_n232_, keyIn_0_6 );
not g129 ( new_n235_, new_n234_ );
and g130 ( new_n236_, new_n235_, new_n233_ );
or g131 ( new_n237_, new_n218_, new_n236_ );
and g132 ( new_n238_, new_n218_, new_n236_ );
not g133 ( new_n239_, new_n238_ );
and g134 ( new_n240_, new_n239_, new_n237_ );
or g135 ( new_n241_, new_n240_, new_n199_ );
not g136 ( new_n242_, new_n217_ );
or g137 ( new_n243_, new_n242_, new_n215_ );
not g138 ( new_n244_, keyIn_0_6 );
not g139 ( new_n245_, new_n232_ );
and g140 ( new_n246_, new_n245_, new_n244_ );
or g141 ( new_n247_, new_n246_, new_n234_ );
and g142 ( new_n248_, new_n243_, new_n247_ );
or g143 ( new_n249_, new_n248_, new_n238_ );
or g144 ( new_n250_, new_n249_, keyIn_0_21 );
and g145 ( new_n251_, new_n241_, new_n250_ );
and g146 ( new_n252_, N130, N137 );
or g147 ( new_n253_, new_n251_, new_n252_ );
and g148 ( new_n254_, new_n249_, keyIn_0_21 );
and g149 ( new_n255_, new_n240_, new_n199_ );
or g150 ( new_n256_, new_n255_, new_n254_ );
not g151 ( new_n257_, new_n252_ );
or g152 ( new_n258_, new_n256_, new_n257_ );
and g153 ( new_n259_, new_n258_, new_n253_ );
or g154 ( new_n260_, new_n259_, keyIn_0_25 );
not g155 ( new_n261_, keyIn_0_25 );
and g156 ( new_n262_, new_n256_, new_n257_ );
and g157 ( new_n263_, new_n251_, new_n252_ );
or g158 ( new_n264_, new_n262_, new_n263_ );
or g159 ( new_n265_, new_n264_, new_n261_ );
and g160 ( new_n266_, new_n265_, new_n260_ );
not g161 ( new_n267_, keyIn_0_9 );
not g162 ( new_n268_, N21 );
and g163 ( new_n269_, new_n268_, N5 );
not g164 ( new_n270_, N5 );
and g165 ( new_n271_, new_n270_, N21 );
or g166 ( new_n272_, new_n269_, new_n271_ );
and g167 ( new_n273_, N37, N53 );
not g168 ( new_n274_, N37 );
not g169 ( new_n275_, N53 );
and g170 ( new_n276_, new_n274_, new_n275_ );
or g171 ( new_n277_, new_n276_, new_n273_ );
and g172 ( new_n278_, new_n272_, new_n277_ );
not g173 ( new_n279_, new_n278_ );
or g174 ( new_n280_, new_n272_, new_n277_ );
and g175 ( new_n281_, new_n279_, new_n280_ );
not g176 ( new_n282_, new_n281_ );
and g177 ( new_n283_, new_n282_, new_n267_ );
and g178 ( new_n284_, new_n281_, keyIn_0_9 );
or g179 ( new_n285_, new_n283_, new_n284_ );
or g180 ( new_n286_, new_n266_, new_n285_ );
and g181 ( new_n287_, new_n264_, new_n261_ );
and g182 ( new_n288_, new_n259_, keyIn_0_25 );
or g183 ( new_n289_, new_n287_, new_n288_ );
not g184 ( new_n290_, new_n285_ );
or g185 ( new_n291_, new_n289_, new_n290_ );
and g186 ( new_n292_, new_n291_, new_n286_ );
and g187 ( new_n293_, new_n198_, new_n292_ );
not g188 ( new_n294_, keyIn_0_26 );
or g189 ( new_n295_, new_n149_, new_n236_ );
or g190 ( new_n296_, new_n144_, new_n247_ );
and g191 ( new_n297_, new_n296_, new_n295_ );
or g192 ( new_n298_, new_n297_, keyIn_0_22 );
not g193 ( new_n299_, keyIn_0_22 );
and g194 ( new_n300_, new_n144_, new_n247_ );
and g195 ( new_n301_, new_n149_, new_n236_ );
or g196 ( new_n302_, new_n300_, new_n301_ );
or g197 ( new_n303_, new_n302_, new_n299_ );
and g198 ( new_n304_, new_n298_, new_n303_ );
and g199 ( new_n305_, N131, N137 );
not g200 ( new_n306_, new_n305_ );
or g201 ( new_n307_, new_n304_, new_n306_ );
and g202 ( new_n308_, new_n302_, new_n299_ );
and g203 ( new_n309_, new_n297_, keyIn_0_22 );
or g204 ( new_n310_, new_n309_, new_n308_ );
or g205 ( new_n311_, new_n310_, new_n305_ );
and g206 ( new_n312_, new_n311_, new_n307_ );
or g207 ( new_n313_, new_n312_, new_n294_ );
and g208 ( new_n314_, new_n310_, new_n305_ );
and g209 ( new_n315_, new_n304_, new_n306_ );
or g210 ( new_n316_, new_n314_, new_n315_ );
or g211 ( new_n317_, new_n316_, keyIn_0_26 );
and g212 ( new_n318_, new_n317_, new_n313_ );
not g213 ( new_n319_, N25 );
and g214 ( new_n320_, new_n319_, N9 );
not g215 ( new_n321_, N9 );
and g216 ( new_n322_, new_n321_, N25 );
or g217 ( new_n323_, new_n320_, new_n322_ );
and g218 ( new_n324_, N41, N57 );
not g219 ( new_n325_, N41 );
not g220 ( new_n326_, N57 );
and g221 ( new_n327_, new_n325_, new_n326_ );
or g222 ( new_n328_, new_n327_, new_n324_ );
and g223 ( new_n329_, new_n323_, new_n328_ );
not g224 ( new_n330_, new_n329_ );
or g225 ( new_n331_, new_n323_, new_n328_ );
and g226 ( new_n332_, new_n330_, new_n331_ );
not g227 ( new_n333_, new_n332_ );
and g228 ( new_n334_, new_n333_, keyIn_0_10 );
not g229 ( new_n335_, new_n334_ );
or g230 ( new_n336_, new_n333_, keyIn_0_10 );
and g231 ( new_n337_, new_n335_, new_n336_ );
or g232 ( new_n338_, new_n318_, new_n337_ );
and g233 ( new_n339_, new_n316_, keyIn_0_26 );
and g234 ( new_n340_, new_n312_, new_n294_ );
or g235 ( new_n341_, new_n339_, new_n340_ );
not g236 ( new_n342_, new_n337_ );
or g237 ( new_n343_, new_n341_, new_n342_ );
and g238 ( new_n344_, new_n343_, new_n338_ );
not g239 ( new_n345_, keyIn_0_23 );
and g240 ( new_n346_, new_n125_, new_n243_ );
not g241 ( new_n347_, new_n346_ );
or g242 ( new_n348_, new_n125_, new_n243_ );
and g243 ( new_n349_, new_n347_, new_n348_ );
or g244 ( new_n350_, new_n349_, new_n345_ );
and g245 ( new_n351_, new_n146_, new_n218_ );
or g246 ( new_n352_, new_n351_, new_n346_ );
or g247 ( new_n353_, new_n352_, keyIn_0_23 );
and g248 ( new_n354_, new_n353_, new_n350_ );
and g249 ( new_n355_, N132, N137 );
or g250 ( new_n356_, new_n354_, new_n355_ );
and g251 ( new_n357_, new_n352_, keyIn_0_23 );
and g252 ( new_n358_, new_n349_, new_n345_ );
or g253 ( new_n359_, new_n357_, new_n358_ );
not g254 ( new_n360_, new_n355_ );
or g255 ( new_n361_, new_n359_, new_n360_ );
and g256 ( new_n362_, new_n361_, new_n356_ );
or g257 ( new_n363_, new_n362_, keyIn_0_27 );
not g258 ( new_n364_, keyIn_0_27 );
and g259 ( new_n365_, new_n359_, new_n360_ );
and g260 ( new_n366_, new_n354_, new_n355_ );
or g261 ( new_n367_, new_n365_, new_n366_ );
or g262 ( new_n368_, new_n367_, new_n364_ );
and g263 ( new_n369_, new_n368_, new_n363_ );
not g264 ( new_n370_, keyIn_0_11 );
not g265 ( new_n371_, N29 );
and g266 ( new_n372_, new_n371_, N13 );
not g267 ( new_n373_, N13 );
and g268 ( new_n374_, new_n373_, N29 );
or g269 ( new_n375_, new_n372_, new_n374_ );
and g270 ( new_n376_, N45, N61 );
not g271 ( new_n377_, N45 );
not g272 ( new_n378_, N61 );
and g273 ( new_n379_, new_n377_, new_n378_ );
or g274 ( new_n380_, new_n379_, new_n376_ );
and g275 ( new_n381_, new_n375_, new_n380_ );
not g276 ( new_n382_, new_n381_ );
or g277 ( new_n383_, new_n375_, new_n380_ );
and g278 ( new_n384_, new_n382_, new_n383_ );
not g279 ( new_n385_, new_n384_ );
and g280 ( new_n386_, new_n385_, new_n370_ );
and g281 ( new_n387_, new_n384_, keyIn_0_11 );
or g282 ( new_n388_, new_n386_, new_n387_ );
not g283 ( new_n389_, new_n388_ );
or g284 ( new_n390_, new_n369_, new_n389_ );
and g285 ( new_n391_, new_n367_, new_n364_ );
and g286 ( new_n392_, new_n362_, keyIn_0_27 );
or g287 ( new_n393_, new_n391_, new_n392_ );
or g288 ( new_n394_, new_n393_, new_n388_ );
and g289 ( new_n395_, new_n394_, new_n390_ );
and g290 ( new_n396_, new_n395_, new_n344_ );
and g291 ( new_n397_, new_n293_, new_n396_ );
not g292 ( new_n398_, keyIn_0_16 );
or g293 ( new_n399_, new_n173_, N21 );
or g294 ( new_n400_, new_n268_, N17 );
and g295 ( new_n401_, new_n399_, new_n400_ );
and g296 ( new_n402_, new_n371_, N25 );
and g297 ( new_n403_, new_n319_, N29 );
or g298 ( new_n404_, new_n402_, new_n403_ );
or g299 ( new_n405_, new_n404_, new_n401_ );
and g300 ( new_n406_, new_n268_, N17 );
and g301 ( new_n407_, new_n173_, N21 );
or g302 ( new_n408_, new_n406_, new_n407_ );
or g303 ( new_n409_, new_n319_, N29 );
or g304 ( new_n410_, new_n371_, N25 );
and g305 ( new_n411_, new_n409_, new_n410_ );
or g306 ( new_n412_, new_n408_, new_n411_ );
and g307 ( new_n413_, new_n405_, new_n412_ );
and g308 ( new_n414_, new_n413_, keyIn_0_1 );
not g309 ( new_n415_, keyIn_0_1 );
and g310 ( new_n416_, new_n408_, new_n411_ );
and g311 ( new_n417_, new_n404_, new_n401_ );
or g312 ( new_n418_, new_n416_, new_n417_ );
and g313 ( new_n419_, new_n418_, new_n415_ );
or g314 ( new_n420_, new_n419_, new_n414_ );
not g315 ( new_n421_, keyIn_0_0 );
and g316 ( new_n422_, new_n270_, N1 );
and g317 ( new_n423_, new_n175_, N5 );
or g318 ( new_n424_, new_n422_, new_n423_ );
and g319 ( new_n425_, new_n373_, N9 );
and g320 ( new_n426_, new_n321_, N13 );
or g321 ( new_n427_, new_n425_, new_n426_ );
or g322 ( new_n428_, new_n424_, new_n427_ );
or g323 ( new_n429_, new_n175_, N5 );
or g324 ( new_n430_, new_n270_, N1 );
and g325 ( new_n431_, new_n429_, new_n430_ );
or g326 ( new_n432_, new_n321_, N13 );
or g327 ( new_n433_, new_n373_, N9 );
and g328 ( new_n434_, new_n432_, new_n433_ );
or g329 ( new_n435_, new_n431_, new_n434_ );
and g330 ( new_n436_, new_n428_, new_n435_ );
and g331 ( new_n437_, new_n436_, new_n421_ );
and g332 ( new_n438_, new_n431_, new_n434_ );
and g333 ( new_n439_, new_n424_, new_n427_ );
or g334 ( new_n440_, new_n439_, new_n438_ );
and g335 ( new_n441_, new_n440_, keyIn_0_0 );
or g336 ( new_n442_, new_n437_, new_n441_ );
and g337 ( new_n443_, new_n420_, new_n442_ );
or g338 ( new_n444_, new_n418_, new_n415_ );
or g339 ( new_n445_, new_n413_, keyIn_0_1 );
and g340 ( new_n446_, new_n444_, new_n445_ );
or g341 ( new_n447_, new_n440_, keyIn_0_0 );
or g342 ( new_n448_, new_n436_, new_n421_ );
and g343 ( new_n449_, new_n448_, new_n447_ );
and g344 ( new_n450_, new_n446_, new_n449_ );
or g345 ( new_n451_, new_n443_, new_n450_ );
and g346 ( new_n452_, new_n451_, new_n398_ );
or g347 ( new_n453_, new_n446_, new_n449_ );
or g348 ( new_n454_, new_n420_, new_n442_ );
and g349 ( new_n455_, new_n454_, new_n453_ );
and g350 ( new_n456_, new_n455_, keyIn_0_16 );
or g351 ( new_n457_, new_n456_, new_n452_ );
and g352 ( new_n458_, N133, N137 );
and g353 ( new_n459_, new_n457_, new_n458_ );
or g354 ( new_n460_, new_n455_, keyIn_0_16 );
or g355 ( new_n461_, new_n451_, new_n398_ );
and g356 ( new_n462_, new_n460_, new_n461_ );
not g357 ( new_n463_, new_n458_ );
and g358 ( new_n464_, new_n462_, new_n463_ );
or g359 ( new_n465_, new_n459_, new_n464_ );
and g360 ( new_n466_, new_n465_, keyIn_0_28 );
not g361 ( new_n467_, keyIn_0_28 );
or g362 ( new_n468_, new_n462_, new_n463_ );
or g363 ( new_n469_, new_n457_, new_n458_ );
and g364 ( new_n470_, new_n469_, new_n468_ );
and g365 ( new_n471_, new_n470_, new_n467_ );
or g366 ( new_n472_, new_n466_, new_n471_ );
not g367 ( new_n473_, keyIn_0_12 );
and g368 ( new_n474_, new_n110_, N65 );
and g369 ( new_n475_, new_n133_, N81 );
or g370 ( new_n476_, new_n474_, new_n475_ );
and g371 ( new_n477_, N97, N113 );
and g372 ( new_n478_, new_n225_, new_n202_ );
or g373 ( new_n479_, new_n478_, new_n477_ );
and g374 ( new_n480_, new_n476_, new_n479_ );
not g375 ( new_n481_, new_n480_ );
or g376 ( new_n482_, new_n476_, new_n479_ );
and g377 ( new_n483_, new_n481_, new_n482_ );
not g378 ( new_n484_, new_n483_ );
and g379 ( new_n485_, new_n484_, new_n473_ );
and g380 ( new_n486_, new_n483_, keyIn_0_12 );
or g381 ( new_n487_, new_n485_, new_n486_ );
and g382 ( new_n488_, new_n472_, new_n487_ );
or g383 ( new_n489_, new_n470_, new_n467_ );
or g384 ( new_n490_, new_n465_, keyIn_0_28 );
and g385 ( new_n491_, new_n490_, new_n489_ );
not g386 ( new_n492_, new_n487_ );
and g387 ( new_n493_, new_n491_, new_n492_ );
or g388 ( new_n494_, new_n488_, new_n493_ );
not g389 ( new_n495_, keyIn_0_31 );
and g390 ( new_n496_, new_n275_, N49 );
and g391 ( new_n497_, new_n180_, N53 );
or g392 ( new_n498_, new_n496_, new_n497_ );
and g393 ( new_n499_, new_n378_, N57 );
and g394 ( new_n500_, new_n326_, N61 );
or g395 ( new_n501_, new_n499_, new_n500_ );
or g396 ( new_n502_, new_n498_, new_n501_ );
or g397 ( new_n503_, new_n180_, N53 );
or g398 ( new_n504_, new_n275_, N49 );
and g399 ( new_n505_, new_n503_, new_n504_ );
or g400 ( new_n506_, new_n326_, N61 );
or g401 ( new_n507_, new_n378_, N57 );
and g402 ( new_n508_, new_n506_, new_n507_ );
or g403 ( new_n509_, new_n505_, new_n508_ );
and g404 ( new_n510_, new_n502_, new_n509_ );
and g405 ( new_n511_, new_n510_, keyIn_0_3 );
not g406 ( new_n512_, keyIn_0_3 );
and g407 ( new_n513_, new_n505_, new_n508_ );
and g408 ( new_n514_, new_n498_, new_n501_ );
or g409 ( new_n515_, new_n514_, new_n513_ );
and g410 ( new_n516_, new_n515_, new_n512_ );
or g411 ( new_n517_, new_n511_, new_n516_ );
and g412 ( new_n518_, new_n517_, new_n446_ );
or g413 ( new_n519_, new_n515_, new_n512_ );
or g414 ( new_n520_, new_n510_, keyIn_0_3 );
and g415 ( new_n521_, new_n520_, new_n519_ );
and g416 ( new_n522_, new_n420_, new_n521_ );
or g417 ( new_n523_, new_n518_, new_n522_ );
and g418 ( new_n524_, new_n523_, keyIn_0_19 );
not g419 ( new_n525_, new_n524_ );
or g420 ( new_n526_, new_n523_, keyIn_0_19 );
and g421 ( new_n527_, new_n525_, new_n526_ );
and g422 ( new_n528_, N136, N137 );
or g423 ( new_n529_, new_n527_, new_n528_ );
and g424 ( new_n530_, new_n527_, new_n528_ );
not g425 ( new_n531_, new_n530_ );
and g426 ( new_n532_, new_n531_, new_n529_ );
or g427 ( new_n533_, new_n532_, new_n495_ );
not g428 ( new_n534_, new_n529_ );
or g429 ( new_n535_, new_n534_, new_n530_ );
or g430 ( new_n536_, new_n535_, keyIn_0_31 );
and g431 ( new_n537_, new_n536_, new_n533_ );
not g432 ( new_n538_, N93 );
and g433 ( new_n539_, new_n538_, N77 );
and g434 ( new_n540_, new_n129_, N93 );
or g435 ( new_n541_, new_n539_, new_n540_ );
and g436 ( new_n542_, N109, N125 );
and g437 ( new_n543_, new_n221_, new_n208_ );
or g438 ( new_n544_, new_n543_, new_n542_ );
and g439 ( new_n545_, new_n541_, new_n544_ );
not g440 ( new_n546_, new_n545_ );
or g441 ( new_n547_, new_n541_, new_n544_ );
and g442 ( new_n548_, new_n546_, new_n547_ );
not g443 ( new_n549_, new_n548_ );
and g444 ( new_n550_, new_n549_, keyIn_0_15 );
not g445 ( new_n551_, new_n550_ );
or g446 ( new_n552_, new_n549_, keyIn_0_15 );
and g447 ( new_n553_, new_n551_, new_n552_ );
or g448 ( new_n554_, new_n537_, new_n553_ );
and g449 ( new_n555_, new_n535_, keyIn_0_31 );
and g450 ( new_n556_, new_n532_, new_n495_ );
or g451 ( new_n557_, new_n555_, new_n556_ );
not g452 ( new_n558_, new_n553_ );
or g453 ( new_n559_, new_n557_, new_n558_ );
and g454 ( new_n560_, new_n559_, new_n554_ );
not g455 ( new_n561_, keyIn_0_30 );
not g456 ( new_n562_, keyIn_0_2 );
or g457 ( new_n563_, new_n325_, N45 );
or g458 ( new_n564_, new_n377_, N41 );
and g459 ( new_n565_, new_n563_, new_n564_ );
and g460 ( new_n566_, N33, N37 );
not g461 ( new_n567_, new_n566_ );
or g462 ( new_n568_, N33, N37 );
and g463 ( new_n569_, new_n567_, new_n568_ );
and g464 ( new_n570_, new_n565_, new_n569_ );
and g465 ( new_n571_, new_n377_, N41 );
and g466 ( new_n572_, new_n325_, N45 );
or g467 ( new_n573_, new_n571_, new_n572_ );
and g468 ( new_n574_, new_n179_, new_n274_ );
or g469 ( new_n575_, new_n574_, new_n566_ );
and g470 ( new_n576_, new_n573_, new_n575_ );
or g471 ( new_n577_, new_n576_, new_n570_ );
and g472 ( new_n578_, new_n577_, new_n562_ );
or g473 ( new_n579_, new_n573_, new_n575_ );
or g474 ( new_n580_, new_n565_, new_n569_ );
and g475 ( new_n581_, new_n579_, new_n580_ );
and g476 ( new_n582_, new_n581_, keyIn_0_2 );
or g477 ( new_n583_, new_n578_, new_n582_ );
and g478 ( new_n584_, new_n583_, new_n449_ );
or g479 ( new_n585_, new_n581_, keyIn_0_2 );
or g480 ( new_n586_, new_n577_, new_n562_ );
and g481 ( new_n587_, new_n585_, new_n586_ );
and g482 ( new_n588_, new_n442_, new_n587_ );
or g483 ( new_n589_, new_n588_, new_n584_ );
and g484 ( new_n590_, new_n589_, keyIn_0_18 );
not g485 ( new_n591_, keyIn_0_18 );
or g486 ( new_n592_, new_n442_, new_n587_ );
or g487 ( new_n593_, new_n583_, new_n449_ );
and g488 ( new_n594_, new_n593_, new_n592_ );
and g489 ( new_n595_, new_n594_, new_n591_ );
or g490 ( new_n596_, new_n590_, new_n595_ );
and g491 ( new_n597_, N135, N137 );
or g492 ( new_n598_, new_n596_, new_n597_ );
or g493 ( new_n599_, new_n594_, new_n591_ );
or g494 ( new_n600_, new_n589_, keyIn_0_18 );
and g495 ( new_n601_, new_n600_, new_n599_ );
not g496 ( new_n602_, new_n597_ );
or g497 ( new_n603_, new_n601_, new_n602_ );
and g498 ( new_n604_, new_n598_, new_n603_ );
or g499 ( new_n605_, new_n604_, new_n561_ );
and g500 ( new_n606_, new_n601_, new_n602_ );
and g501 ( new_n607_, new_n596_, new_n597_ );
or g502 ( new_n608_, new_n607_, new_n606_ );
or g503 ( new_n609_, new_n608_, keyIn_0_30 );
and g504 ( new_n610_, new_n609_, new_n605_ );
not g505 ( new_n611_, N89 );
and g506 ( new_n612_, new_n611_, N73 );
and g507 ( new_n613_, new_n128_, N89 );
or g508 ( new_n614_, new_n612_, new_n613_ );
and g509 ( new_n615_, N105, N121 );
and g510 ( new_n616_, new_n220_, new_n207_ );
or g511 ( new_n617_, new_n616_, new_n615_ );
and g512 ( new_n618_, new_n614_, new_n617_ );
not g513 ( new_n619_, new_n618_ );
or g514 ( new_n620_, new_n614_, new_n617_ );
and g515 ( new_n621_, new_n619_, new_n620_ );
not g516 ( new_n622_, new_n621_ );
and g517 ( new_n623_, new_n622_, keyIn_0_14 );
not g518 ( new_n624_, new_n623_ );
or g519 ( new_n625_, new_n622_, keyIn_0_14 );
and g520 ( new_n626_, new_n624_, new_n625_ );
not g521 ( new_n627_, new_n626_ );
or g522 ( new_n628_, new_n610_, new_n627_ );
and g523 ( new_n629_, new_n608_, keyIn_0_30 );
and g524 ( new_n630_, new_n604_, new_n561_ );
or g525 ( new_n631_, new_n629_, new_n630_ );
or g526 ( new_n632_, new_n631_, new_n626_ );
and g527 ( new_n633_, new_n632_, new_n628_ );
not g528 ( new_n634_, new_n633_ );
and g529 ( new_n635_, new_n560_, new_n634_ );
and g530 ( new_n636_, new_n517_, new_n583_ );
and g531 ( new_n637_, new_n521_, new_n587_ );
or g532 ( new_n638_, new_n636_, new_n637_ );
and g533 ( new_n639_, new_n638_, keyIn_0_17 );
not g534 ( new_n640_, keyIn_0_17 );
or g535 ( new_n641_, new_n521_, new_n587_ );
or g536 ( new_n642_, new_n517_, new_n583_ );
and g537 ( new_n643_, new_n642_, new_n641_ );
and g538 ( new_n644_, new_n643_, new_n640_ );
or g539 ( new_n645_, new_n644_, new_n639_ );
and g540 ( new_n646_, N134, N137 );
not g541 ( new_n647_, new_n646_ );
and g542 ( new_n648_, new_n645_, new_n647_ );
or g543 ( new_n649_, new_n643_, new_n640_ );
or g544 ( new_n650_, new_n638_, keyIn_0_17 );
and g545 ( new_n651_, new_n649_, new_n650_ );
and g546 ( new_n652_, new_n651_, new_n646_ );
or g547 ( new_n653_, new_n648_, new_n652_ );
and g548 ( new_n654_, new_n653_, keyIn_0_29 );
not g549 ( new_n655_, keyIn_0_29 );
or g550 ( new_n656_, new_n651_, new_n646_ );
or g551 ( new_n657_, new_n645_, new_n647_ );
and g552 ( new_n658_, new_n657_, new_n656_ );
and g553 ( new_n659_, new_n658_, new_n655_ );
or g554 ( new_n660_, new_n654_, new_n659_ );
not g555 ( new_n661_, keyIn_0_13 );
and g556 ( new_n662_, new_n108_, N69 );
and g557 ( new_n663_, new_n134_, N85 );
or g558 ( new_n664_, new_n662_, new_n663_ );
and g559 ( new_n665_, N101, N117 );
and g560 ( new_n666_, new_n226_, new_n203_ );
or g561 ( new_n667_, new_n666_, new_n665_ );
and g562 ( new_n668_, new_n664_, new_n667_ );
not g563 ( new_n669_, new_n668_ );
or g564 ( new_n670_, new_n664_, new_n667_ );
and g565 ( new_n671_, new_n669_, new_n670_ );
not g566 ( new_n672_, new_n671_ );
and g567 ( new_n673_, new_n672_, new_n661_ );
and g568 ( new_n674_, new_n671_, keyIn_0_13 );
or g569 ( new_n675_, new_n673_, new_n674_ );
not g570 ( new_n676_, new_n675_ );
and g571 ( new_n677_, new_n660_, new_n676_ );
or g572 ( new_n678_, new_n658_, new_n655_ );
or g573 ( new_n679_, new_n653_, keyIn_0_29 );
and g574 ( new_n680_, new_n679_, new_n678_ );
and g575 ( new_n681_, new_n680_, new_n675_ );
or g576 ( new_n682_, new_n677_, new_n681_ );
not g577 ( new_n683_, new_n682_ );
and g578 ( new_n684_, new_n635_, new_n683_ );
and g579 ( new_n685_, new_n684_, new_n494_ );
and g580 ( new_n686_, new_n685_, new_n397_ );
not g581 ( new_n687_, new_n686_ );
and g582 ( new_n688_, new_n687_, N1 );
and g583 ( new_n689_, new_n686_, new_n175_ );
or g584 ( N724, new_n688_, new_n689_ );
or g585 ( new_n691_, new_n195_, new_n196_ );
or g586 ( new_n692_, new_n172_, new_n191_ );
and g587 ( new_n693_, new_n692_, new_n691_ );
not g588 ( new_n694_, new_n292_ );
and g589 ( new_n695_, new_n693_, new_n694_ );
and g590 ( new_n696_, new_n396_, new_n695_ );
and g591 ( new_n697_, new_n685_, new_n696_ );
not g592 ( new_n698_, new_n697_ );
and g593 ( new_n699_, new_n698_, N5 );
and g594 ( new_n700_, new_n697_, new_n270_ );
or g595 ( N725, new_n699_, new_n700_ );
not g596 ( new_n702_, new_n344_ );
and g597 ( new_n703_, new_n395_, new_n702_ );
and g598 ( new_n704_, new_n693_, new_n292_ );
and g599 ( new_n705_, new_n703_, new_n704_ );
and g600 ( new_n706_, new_n685_, new_n705_ );
not g601 ( new_n707_, new_n706_ );
and g602 ( new_n708_, new_n707_, N9 );
and g603 ( new_n709_, new_n706_, new_n321_ );
or g604 ( N726, new_n708_, new_n709_ );
and g605 ( new_n711_, new_n393_, new_n388_ );
and g606 ( new_n712_, new_n369_, new_n389_ );
or g607 ( new_n713_, new_n711_, new_n712_ );
and g608 ( new_n714_, new_n292_, new_n344_ );
and g609 ( new_n715_, new_n714_, new_n713_ );
and g610 ( new_n716_, new_n715_, new_n693_ );
and g611 ( new_n717_, new_n685_, new_n716_ );
not g612 ( new_n718_, new_n717_ );
and g613 ( new_n719_, new_n718_, N13 );
and g614 ( new_n720_, new_n717_, new_n373_ );
or g615 ( N727, new_n719_, new_n720_ );
and g616 ( new_n722_, new_n557_, new_n558_ );
and g617 ( new_n723_, new_n537_, new_n553_ );
or g618 ( new_n724_, new_n722_, new_n723_ );
and g619 ( new_n725_, new_n494_, new_n633_ );
and g620 ( new_n726_, new_n725_, new_n683_ );
and g621 ( new_n727_, new_n726_, new_n724_ );
and g622 ( new_n728_, new_n397_, new_n727_ );
not g623 ( new_n729_, new_n728_ );
and g624 ( new_n730_, new_n729_, N17 );
and g625 ( new_n731_, new_n728_, new_n173_ );
or g626 ( N728, new_n730_, new_n731_ );
and g627 ( new_n733_, new_n696_, new_n727_ );
not g628 ( new_n734_, new_n733_ );
and g629 ( new_n735_, new_n734_, N21 );
and g630 ( new_n736_, new_n733_, new_n268_ );
or g631 ( N729, new_n735_, new_n736_ );
and g632 ( new_n738_, new_n705_, new_n727_ );
not g633 ( new_n739_, new_n738_ );
and g634 ( new_n740_, new_n739_, N25 );
and g635 ( new_n741_, new_n738_, new_n319_ );
or g636 ( N730, new_n740_, new_n741_ );
and g637 ( new_n743_, new_n716_, new_n727_ );
not g638 ( new_n744_, new_n743_ );
and g639 ( new_n745_, new_n744_, N29 );
and g640 ( new_n746_, new_n743_, new_n371_ );
or g641 ( N731, new_n745_, new_n746_ );
or g642 ( new_n748_, new_n491_, new_n492_ );
or g643 ( new_n749_, new_n472_, new_n487_ );
and g644 ( new_n750_, new_n749_, new_n748_ );
and g645 ( new_n751_, new_n750_, new_n682_ );
and g646 ( new_n752_, new_n635_, new_n751_ );
and g647 ( new_n753_, new_n397_, new_n752_ );
not g648 ( new_n754_, new_n753_ );
and g649 ( new_n755_, new_n754_, N33 );
and g650 ( new_n756_, new_n753_, new_n179_ );
or g651 ( N732, new_n755_, new_n756_ );
and g652 ( new_n758_, new_n696_, new_n752_ );
not g653 ( new_n759_, new_n758_ );
and g654 ( new_n760_, new_n759_, N37 );
and g655 ( new_n761_, new_n758_, new_n274_ );
or g656 ( N733, new_n760_, new_n761_ );
and g657 ( new_n763_, new_n705_, new_n752_ );
not g658 ( new_n764_, new_n763_ );
and g659 ( new_n765_, new_n764_, N41 );
and g660 ( new_n766_, new_n763_, new_n325_ );
or g661 ( N734, new_n765_, new_n766_ );
and g662 ( new_n768_, new_n716_, new_n752_ );
not g663 ( new_n769_, new_n768_ );
and g664 ( new_n770_, new_n769_, N45 );
and g665 ( new_n771_, new_n768_, new_n377_ );
or g666 ( N735, new_n770_, new_n771_ );
and g667 ( new_n773_, new_n751_, new_n633_ );
and g668 ( new_n774_, new_n773_, new_n724_ );
and g669 ( new_n775_, new_n397_, new_n774_ );
not g670 ( new_n776_, new_n775_ );
and g671 ( new_n777_, new_n776_, N49 );
and g672 ( new_n778_, new_n775_, new_n180_ );
or g673 ( N736, new_n777_, new_n778_ );
and g674 ( new_n780_, new_n696_, new_n774_ );
not g675 ( new_n781_, new_n780_ );
and g676 ( new_n782_, new_n781_, N53 );
and g677 ( new_n783_, new_n780_, new_n275_ );
or g678 ( N737, new_n782_, new_n783_ );
and g679 ( new_n785_, new_n705_, new_n774_ );
not g680 ( new_n786_, new_n785_ );
and g681 ( new_n787_, new_n786_, N57 );
and g682 ( new_n788_, new_n785_, new_n326_ );
or g683 ( N738, new_n787_, new_n788_ );
and g684 ( new_n790_, new_n716_, new_n774_ );
not g685 ( new_n791_, new_n790_ );
and g686 ( new_n792_, new_n791_, N61 );
and g687 ( new_n793_, new_n790_, new_n378_ );
or g688 ( N739, new_n792_, new_n793_ );
and g689 ( new_n795_, new_n293_, new_n703_ );
and g690 ( new_n796_, new_n726_, new_n560_ );
and g691 ( new_n797_, new_n795_, new_n796_ );
not g692 ( new_n798_, new_n797_ );
and g693 ( new_n799_, new_n798_, N65 );
and g694 ( new_n800_, new_n797_, new_n133_ );
or g695 ( N740, new_n799_, new_n800_ );
and g696 ( new_n802_, new_n773_, new_n560_ );
and g697 ( new_n803_, new_n795_, new_n802_ );
not g698 ( new_n804_, new_n803_ );
and g699 ( new_n805_, new_n804_, N69 );
and g700 ( new_n806_, new_n803_, new_n134_ );
or g701 ( N741, new_n805_, new_n806_ );
and g702 ( new_n808_, new_n684_, new_n750_ );
and g703 ( new_n809_, new_n808_, new_n795_ );
not g704 ( new_n810_, new_n809_ );
and g705 ( new_n811_, new_n810_, N73 );
and g706 ( new_n812_, new_n809_, new_n128_ );
or g707 ( N742, new_n811_, new_n812_ );
or g708 ( new_n814_, new_n726_, new_n773_ );
and g709 ( new_n815_, new_n814_, new_n560_ );
and g710 ( new_n816_, new_n724_, new_n633_ );
or g711 ( new_n817_, new_n816_, new_n635_ );
and g712 ( new_n818_, new_n683_, new_n750_ );
and g713 ( new_n819_, new_n817_, new_n818_ );
or g714 ( new_n820_, new_n815_, new_n819_ );
and g715 ( new_n821_, new_n724_, new_n129_ );
and g716 ( new_n822_, new_n795_, new_n821_ );
and g717 ( new_n823_, new_n820_, new_n822_ );
and g718 ( new_n824_, new_n816_, new_n818_ );
and g719 ( new_n825_, new_n795_, new_n824_ );
not g720 ( new_n826_, new_n825_ );
and g721 ( new_n827_, new_n826_, N77 );
or g722 ( N743, new_n823_, new_n827_ );
and g723 ( new_n829_, new_n715_, new_n198_ );
and g724 ( new_n830_, new_n829_, new_n796_ );
not g725 ( new_n831_, new_n830_ );
and g726 ( new_n832_, new_n831_, N81 );
and g727 ( new_n833_, new_n830_, new_n110_ );
or g728 ( N744, new_n832_, new_n833_ );
and g729 ( new_n835_, new_n829_, new_n802_ );
not g730 ( new_n836_, new_n835_ );
and g731 ( new_n837_, new_n836_, N85 );
and g732 ( new_n838_, new_n835_, new_n108_ );
or g733 ( N745, new_n837_, new_n838_ );
and g734 ( new_n840_, new_n808_, new_n829_ );
not g735 ( new_n841_, new_n840_ );
and g736 ( new_n842_, new_n841_, N89 );
and g737 ( new_n843_, new_n840_, new_n611_ );
or g738 ( N746, new_n842_, new_n843_ );
and g739 ( new_n845_, new_n724_, new_n538_ );
and g740 ( new_n846_, new_n829_, new_n845_ );
and g741 ( new_n847_, new_n820_, new_n846_ );
and g742 ( new_n848_, new_n829_, new_n824_ );
not g743 ( new_n849_, new_n848_ );
and g744 ( new_n850_, new_n849_, N93 );
or g745 ( N747, new_n847_, new_n850_ );
and g746 ( new_n852_, new_n695_, new_n703_ );
and g747 ( new_n853_, new_n852_, new_n796_ );
not g748 ( new_n854_, new_n853_ );
and g749 ( new_n855_, new_n854_, N97 );
and g750 ( new_n856_, new_n853_, new_n225_ );
or g751 ( N748, new_n855_, new_n856_ );
and g752 ( new_n858_, new_n852_, new_n802_ );
not g753 ( new_n859_, new_n858_ );
and g754 ( new_n860_, new_n859_, N101 );
and g755 ( new_n861_, new_n858_, new_n226_ );
or g756 ( N749, new_n860_, new_n861_ );
and g757 ( new_n863_, new_n808_, new_n852_ );
not g758 ( new_n864_, new_n863_ );
and g759 ( new_n865_, new_n864_, N105 );
and g760 ( new_n866_, new_n863_, new_n220_ );
or g761 ( N750, new_n865_, new_n866_ );
and g762 ( new_n868_, new_n724_, new_n221_ );
and g763 ( new_n869_, new_n852_, new_n868_ );
and g764 ( new_n870_, new_n820_, new_n869_ );
and g765 ( new_n871_, new_n852_, new_n824_ );
not g766 ( new_n872_, new_n871_ );
and g767 ( new_n873_, new_n872_, N109 );
or g768 ( N751, new_n870_, new_n873_ );
and g769 ( new_n875_, new_n713_, new_n344_ );
and g770 ( new_n876_, new_n875_, new_n695_ );
and g771 ( new_n877_, new_n876_, new_n796_ );
not g772 ( new_n878_, new_n877_ );
and g773 ( new_n879_, new_n878_, N113 );
and g774 ( new_n880_, new_n877_, new_n202_ );
or g775 ( N752, new_n879_, new_n880_ );
and g776 ( new_n882_, new_n876_, new_n802_ );
not g777 ( new_n883_, new_n882_ );
and g778 ( new_n884_, new_n883_, N117 );
and g779 ( new_n885_, new_n882_, new_n203_ );
or g780 ( N753, new_n884_, new_n885_ );
and g781 ( new_n887_, new_n808_, new_n876_ );
not g782 ( new_n888_, new_n887_ );
and g783 ( new_n889_, new_n888_, N121 );
and g784 ( new_n890_, new_n887_, new_n207_ );
or g785 ( N754, new_n889_, new_n890_ );
and g786 ( new_n892_, new_n724_, new_n208_ );
and g787 ( new_n893_, new_n876_, new_n892_ );
and g788 ( new_n894_, new_n820_, new_n893_ );
and g789 ( new_n895_, new_n876_, new_n824_ );
not g790 ( new_n896_, new_n895_ );
and g791 ( new_n897_, new_n896_, N125 );
or g792 ( N755, new_n894_, new_n897_ );
endmodule