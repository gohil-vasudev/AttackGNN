module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1517_, new_n1575_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n1568_, new_n728_, new_n1479_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n1662_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n1620_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1580_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n1595_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n1640_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1632_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n1647_, new_n324_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n394_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n1657_, new_n1562_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n1576_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n1395_, new_n473_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n1574_, new_n1614_, new_n621_, new_n1423_, new_n1637_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1201_, new_n559_, new_n1282_, new_n1630_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1437_, new_n1598_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n1546_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n1573_, new_n369_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n276_, new_n1032_, new_n1545_, new_n901_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n261_, new_n672_, new_n1496_, new_n1269_, new_n616_, new_n1653_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n1600_, new_n1592_, new_n809_, new_n1631_, new_n1142_, new_n1623_, new_n604_, new_n1461_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1656_, new_n1252_, new_n352_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n1593_, new_n944_, new_n1638_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1625_, new_n993_, new_n1191_, new_n1357_, new_n824_, new_n1628_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1612_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n302_, new_n755_, new_n1040_, new_n1635_, new_n1509_, new_n1559_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1185_, new_n1240_, new_n1510_, new_n354_, new_n968_, new_n1655_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1334_, new_n531_, new_n593_, new_n1543_, new_n1565_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n1660_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1608_, new_n1492_, new_n1619_, new_n278_, new_n304_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n1421_, new_n644_, new_n1594_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n1665_, new_n754_, new_n653_, new_n1659_, new_n905_, new_n377_, new_n1258_, new_n1539_, new_n1643_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n984_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1602_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n1664_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n1567_, new_n1651_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n1597_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1616_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n1644_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1544_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n1646_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n1606_, new_n427_, new_n532_, new_n393_, new_n1617_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1585_, new_n1587_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n966_, new_n351_, new_n1292_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n1560_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1622_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n1618_, new_n1652_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n1611_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1613_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n1584_, new_n1337_, new_n216_, new_n1348_, new_n917_, new_n1555_, new_n1636_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n1601_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n1609_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n1633_, new_n1607_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1582_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1329_, new_n1161_, new_n1648_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1663_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n259_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n222_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1579_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n1621_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n918_, new_n1586_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n253_, new_n825_, new_n1627_, new_n557_, new_n260_, new_n1642_, new_n251_, new_n300_, new_n1503_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n1551_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n1650_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1596_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n1641_, new_n949_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1634_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1649_, new_n1654_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n1571_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1610_, new_n1470_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1604_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1529_, new_n1541_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n1577_, new_n574_, new_n928_, new_n1548_, new_n1578_, new_n319_, new_n1008_, new_n1661_, new_n338_, new_n1615_, new_n707_, new_n740_, new_n957_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n1399_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1589_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1570_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n1583_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n1449_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1605_, new_n464_, new_n1498_, new_n204_, new_n1588_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_43 );
not g0001 ( new_n203_, keyIn_0_32 );
not g0002 ( new_n204_, N69 );
and g0003 ( new_n205_, new_n204_, N65 );
not g0004 ( new_n206_, N65 );
and g0005 ( new_n207_, new_n206_, N69 );
or g0006 ( new_n208_, new_n205_, new_n207_ );
and g0007 ( new_n209_, new_n208_, keyIn_0_8 );
not g0008 ( new_n210_, new_n209_ );
or g0009 ( new_n211_, new_n208_, keyIn_0_8 );
and g0010 ( new_n212_, new_n210_, new_n211_ );
not g0011 ( new_n213_, new_n212_ );
not g0012 ( new_n214_, keyIn_0_9 );
not g0013 ( new_n215_, N77 );
and g0014 ( new_n216_, new_n215_, N73 );
not g0015 ( new_n217_, N73 );
and g0016 ( new_n218_, new_n217_, N77 );
or g0017 ( new_n219_, new_n216_, new_n218_ );
and g0018 ( new_n220_, new_n219_, new_n214_ );
not g0019 ( new_n221_, new_n220_ );
or g0020 ( new_n222_, new_n219_, new_n214_ );
and g0021 ( new_n223_, new_n221_, new_n222_ );
not g0022 ( new_n224_, new_n223_ );
and g0023 ( new_n225_, new_n213_, new_n224_ );
and g0024 ( new_n226_, new_n212_, new_n223_ );
or g0025 ( new_n227_, new_n225_, new_n226_ );
and g0026 ( new_n228_, new_n227_, new_n203_ );
not g0027 ( new_n229_, new_n228_ );
or g0028 ( new_n230_, new_n227_, new_n203_ );
and g0029 ( new_n231_, new_n229_, new_n230_ );
not g0030 ( new_n232_, keyIn_0_10 );
not g0031 ( new_n233_, N85 );
and g0032 ( new_n234_, new_n233_, N81 );
not g0033 ( new_n235_, N81 );
and g0034 ( new_n236_, new_n235_, N85 );
or g0035 ( new_n237_, new_n234_, new_n236_ );
and g0036 ( new_n238_, new_n237_, new_n232_ );
not g0037 ( new_n239_, new_n238_ );
or g0038 ( new_n240_, new_n237_, new_n232_ );
and g0039 ( new_n241_, new_n239_, new_n240_ );
not g0040 ( new_n242_, new_n241_ );
not g0041 ( new_n243_, N93 );
and g0042 ( new_n244_, new_n243_, N89 );
not g0043 ( new_n245_, N89 );
and g0044 ( new_n246_, new_n245_, N93 );
or g0045 ( new_n247_, new_n244_, new_n246_ );
not g0046 ( new_n248_, new_n247_ );
and g0047 ( new_n249_, new_n248_, keyIn_0_11 );
not g0048 ( new_n250_, new_n249_ );
or g0049 ( new_n251_, new_n248_, keyIn_0_11 );
and g0050 ( new_n252_, new_n250_, new_n251_ );
and g0051 ( new_n253_, new_n242_, new_n252_ );
not g0052 ( new_n254_, new_n253_ );
or g0053 ( new_n255_, new_n242_, new_n252_ );
and g0054 ( new_n256_, new_n254_, new_n255_ );
not g0055 ( new_n257_, new_n256_ );
and g0056 ( new_n258_, new_n257_, keyIn_0_33 );
not g0057 ( new_n259_, new_n258_ );
or g0058 ( new_n260_, new_n257_, keyIn_0_33 );
and g0059 ( new_n261_, new_n259_, new_n260_ );
and g0060 ( new_n262_, new_n261_, new_n231_ );
not g0061 ( new_n263_, new_n231_ );
not g0062 ( new_n264_, new_n261_ );
and g0063 ( new_n265_, new_n264_, new_n263_ );
or g0064 ( new_n266_, new_n265_, new_n262_ );
and g0065 ( new_n267_, new_n266_, new_n202_ );
not g0066 ( new_n268_, new_n267_ );
or g0067 ( new_n269_, new_n266_, new_n202_ );
and g0068 ( new_n270_, new_n268_, new_n269_ );
and g0069 ( new_n271_, N129, N137 );
not g0070 ( new_n272_, new_n271_ );
and g0071 ( new_n273_, new_n270_, new_n272_ );
not g0072 ( new_n274_, new_n273_ );
or g0073 ( new_n275_, new_n270_, new_n272_ );
and g0074 ( new_n276_, new_n274_, new_n275_ );
not g0075 ( new_n277_, new_n276_ );
and g0076 ( new_n278_, new_n277_, keyIn_0_47 );
not g0077 ( new_n279_, new_n278_ );
or g0078 ( new_n280_, new_n277_, keyIn_0_47 );
and g0079 ( new_n281_, new_n279_, new_n280_ );
not g0080 ( new_n282_, N17 );
and g0081 ( new_n283_, new_n282_, N1 );
not g0082 ( new_n284_, N1 );
and g0083 ( new_n285_, new_n284_, N17 );
or g0084 ( new_n286_, new_n283_, new_n285_ );
not g0085 ( new_n287_, N49 );
and g0086 ( new_n288_, new_n287_, N33 );
not g0087 ( new_n289_, N33 );
and g0088 ( new_n290_, new_n289_, N49 );
or g0089 ( new_n291_, new_n288_, new_n290_ );
not g0090 ( new_n292_, new_n291_ );
and g0091 ( new_n293_, new_n292_, new_n286_ );
not g0092 ( new_n294_, new_n293_ );
or g0093 ( new_n295_, new_n292_, new_n286_ );
and g0094 ( new_n296_, new_n294_, new_n295_ );
or g0095 ( new_n297_, new_n281_, new_n296_ );
and g0096 ( new_n298_, new_n281_, new_n296_ );
not g0097 ( new_n299_, new_n298_ );
and g0098 ( new_n300_, new_n299_, new_n297_ );
or g0099 ( new_n301_, new_n300_, keyIn_0_55 );
not g0100 ( new_n302_, keyIn_0_55 );
not g0101 ( new_n303_, new_n297_ );
or g0102 ( new_n304_, new_n303_, new_n298_ );
or g0103 ( new_n305_, new_n304_, new_n302_ );
and g0104 ( new_n306_, new_n305_, new_n301_ );
not g0105 ( new_n307_, new_n306_ );
not g0106 ( new_n308_, keyIn_0_57 );
not g0107 ( new_n309_, N101 );
and g0108 ( new_n310_, new_n309_, N97 );
not g0109 ( new_n311_, N97 );
and g0110 ( new_n312_, new_n311_, N101 );
or g0111 ( new_n313_, new_n310_, new_n312_ );
and g0112 ( new_n314_, new_n313_, keyIn_0_12 );
not g0113 ( new_n315_, new_n314_ );
or g0114 ( new_n316_, new_n313_, keyIn_0_12 );
and g0115 ( new_n317_, new_n315_, new_n316_ );
not g0116 ( new_n318_, new_n317_ );
not g0117 ( new_n319_, keyIn_0_13 );
not g0118 ( new_n320_, N109 );
and g0119 ( new_n321_, new_n320_, N105 );
not g0120 ( new_n322_, N105 );
and g0121 ( new_n323_, new_n322_, N109 );
or g0122 ( new_n324_, new_n321_, new_n323_ );
and g0123 ( new_n325_, new_n324_, new_n319_ );
not g0124 ( new_n326_, new_n325_ );
or g0125 ( new_n327_, new_n324_, new_n319_ );
and g0126 ( new_n328_, new_n326_, new_n327_ );
not g0127 ( new_n329_, new_n328_ );
and g0128 ( new_n330_, new_n318_, new_n329_ );
and g0129 ( new_n331_, new_n317_, new_n328_ );
or g0130 ( new_n332_, new_n330_, new_n331_ );
and g0131 ( new_n333_, new_n332_, keyIn_0_34 );
not g0132 ( new_n334_, new_n333_ );
or g0133 ( new_n335_, new_n332_, keyIn_0_34 );
and g0134 ( new_n336_, new_n334_, new_n335_ );
and g0135 ( new_n337_, new_n263_, new_n336_ );
not g0136 ( new_n338_, new_n336_ );
and g0137 ( new_n339_, new_n338_, new_n231_ );
or g0138 ( new_n340_, new_n337_, new_n339_ );
and g0139 ( new_n341_, new_n340_, keyIn_0_45 );
not g0140 ( new_n342_, new_n341_ );
or g0141 ( new_n343_, new_n340_, keyIn_0_45 );
and g0142 ( new_n344_, new_n342_, new_n343_ );
not g0143 ( new_n345_, new_n344_ );
and g0144 ( new_n346_, new_n345_, keyIn_0_16 );
not g0145 ( new_n347_, new_n346_ );
or g0146 ( new_n348_, new_n345_, keyIn_0_16 );
and g0147 ( new_n349_, new_n347_, new_n348_ );
not g0148 ( new_n350_, new_n349_ );
and g0149 ( new_n351_, N131, N137 );
not g0150 ( new_n352_, new_n351_ );
and g0151 ( new_n353_, new_n350_, new_n352_ );
and g0152 ( new_n354_, new_n349_, new_n351_ );
or g0153 ( new_n355_, new_n353_, new_n354_ );
and g0154 ( new_n356_, new_n355_, keyIn_0_49 );
not g0155 ( new_n357_, new_n356_ );
or g0156 ( new_n358_, new_n355_, keyIn_0_49 );
and g0157 ( new_n359_, new_n357_, new_n358_ );
not g0158 ( new_n360_, N25 );
and g0159 ( new_n361_, new_n360_, N9 );
not g0160 ( new_n362_, N9 );
and g0161 ( new_n363_, new_n362_, N25 );
or g0162 ( new_n364_, new_n361_, new_n363_ );
and g0163 ( new_n365_, new_n364_, keyIn_0_21 );
not g0164 ( new_n366_, new_n365_ );
or g0165 ( new_n367_, new_n364_, keyIn_0_21 );
and g0166 ( new_n368_, new_n366_, new_n367_ );
not g0167 ( new_n369_, new_n368_ );
not g0168 ( new_n370_, N57 );
and g0169 ( new_n371_, new_n370_, N41 );
not g0170 ( new_n372_, N41 );
and g0171 ( new_n373_, new_n372_, N57 );
or g0172 ( new_n374_, new_n371_, new_n373_ );
and g0173 ( new_n375_, new_n374_, keyIn_0_22 );
not g0174 ( new_n376_, new_n375_ );
or g0175 ( new_n377_, new_n374_, keyIn_0_22 );
and g0176 ( new_n378_, new_n376_, new_n377_ );
and g0177 ( new_n379_, new_n369_, new_n378_ );
not g0178 ( new_n380_, new_n379_ );
or g0179 ( new_n381_, new_n369_, new_n378_ );
and g0180 ( new_n382_, new_n380_, new_n381_ );
not g0181 ( new_n383_, new_n382_ );
and g0182 ( new_n384_, new_n383_, keyIn_0_36 );
not g0183 ( new_n385_, new_n384_ );
or g0184 ( new_n386_, new_n383_, keyIn_0_36 );
and g0185 ( new_n387_, new_n385_, new_n386_ );
or g0186 ( new_n388_, new_n359_, new_n387_ );
not g0187 ( new_n389_, keyIn_0_49 );
not g0188 ( new_n390_, new_n353_ );
not g0189 ( new_n391_, new_n354_ );
and g0190 ( new_n392_, new_n390_, new_n391_ );
and g0191 ( new_n393_, new_n392_, new_n389_ );
or g0192 ( new_n394_, new_n393_, new_n356_ );
not g0193 ( new_n395_, new_n387_ );
or g0194 ( new_n396_, new_n394_, new_n395_ );
and g0195 ( new_n397_, new_n396_, new_n388_ );
or g0196 ( new_n398_, new_n397_, new_n308_ );
and g0197 ( new_n399_, new_n394_, new_n395_ );
and g0198 ( new_n400_, new_n359_, new_n387_ );
or g0199 ( new_n401_, new_n399_, new_n400_ );
or g0200 ( new_n402_, new_n401_, keyIn_0_57 );
and g0201 ( new_n403_, new_n402_, new_n398_ );
not g0202 ( new_n404_, keyIn_0_50 );
not g0203 ( new_n405_, keyIn_0_46 );
not g0204 ( new_n406_, keyIn_0_35 );
not g0205 ( new_n407_, keyIn_0_14 );
not g0206 ( new_n408_, N117 );
and g0207 ( new_n409_, new_n408_, N113 );
not g0208 ( new_n410_, N113 );
and g0209 ( new_n411_, new_n410_, N117 );
or g0210 ( new_n412_, new_n409_, new_n411_ );
and g0211 ( new_n413_, new_n412_, new_n407_ );
not g0212 ( new_n414_, new_n413_ );
or g0213 ( new_n415_, new_n412_, new_n407_ );
and g0214 ( new_n416_, new_n414_, new_n415_ );
not g0215 ( new_n417_, new_n416_ );
not g0216 ( new_n418_, keyIn_0_15 );
not g0217 ( new_n419_, N125 );
and g0218 ( new_n420_, new_n419_, N121 );
not g0219 ( new_n421_, N121 );
and g0220 ( new_n422_, new_n421_, N125 );
or g0221 ( new_n423_, new_n420_, new_n422_ );
and g0222 ( new_n424_, new_n423_, new_n418_ );
not g0223 ( new_n425_, new_n424_ );
or g0224 ( new_n426_, new_n423_, new_n418_ );
and g0225 ( new_n427_, new_n425_, new_n426_ );
not g0226 ( new_n428_, new_n427_ );
and g0227 ( new_n429_, new_n417_, new_n428_ );
and g0228 ( new_n430_, new_n416_, new_n427_ );
or g0229 ( new_n431_, new_n429_, new_n430_ );
and g0230 ( new_n432_, new_n431_, new_n406_ );
not g0231 ( new_n433_, new_n432_ );
or g0232 ( new_n434_, new_n431_, new_n406_ );
and g0233 ( new_n435_, new_n433_, new_n434_ );
and g0234 ( new_n436_, new_n261_, new_n435_ );
not g0235 ( new_n437_, new_n435_ );
and g0236 ( new_n438_, new_n264_, new_n437_ );
or g0237 ( new_n439_, new_n438_, new_n436_ );
and g0238 ( new_n440_, new_n439_, new_n405_ );
not g0239 ( new_n441_, new_n440_ );
or g0240 ( new_n442_, new_n439_, new_n405_ );
and g0241 ( new_n443_, new_n441_, new_n442_ );
and g0242 ( new_n444_, N132, N137 );
or g0243 ( new_n445_, new_n443_, new_n444_ );
and g0244 ( new_n446_, new_n443_, new_n444_ );
not g0245 ( new_n447_, new_n446_ );
and g0246 ( new_n448_, new_n447_, new_n445_ );
not g0247 ( new_n449_, new_n448_ );
and g0248 ( new_n450_, new_n449_, new_n404_ );
and g0249 ( new_n451_, new_n448_, keyIn_0_50 );
or g0250 ( new_n452_, new_n450_, new_n451_ );
not g0251 ( new_n453_, new_n452_ );
not g0252 ( new_n454_, keyIn_0_23 );
not g0253 ( new_n455_, N29 );
and g0254 ( new_n456_, new_n455_, N13 );
not g0255 ( new_n457_, N13 );
and g0256 ( new_n458_, new_n457_, N29 );
or g0257 ( new_n459_, new_n456_, new_n458_ );
and g0258 ( new_n460_, new_n459_, new_n454_ );
not g0259 ( new_n461_, new_n460_ );
or g0260 ( new_n462_, new_n459_, new_n454_ );
and g0261 ( new_n463_, new_n461_, new_n462_ );
not g0262 ( new_n464_, new_n463_ );
not g0263 ( new_n465_, N61 );
and g0264 ( new_n466_, new_n465_, N45 );
not g0265 ( new_n467_, N45 );
and g0266 ( new_n468_, new_n467_, N61 );
or g0267 ( new_n469_, new_n466_, new_n468_ );
not g0268 ( new_n470_, new_n469_ );
and g0269 ( new_n471_, new_n464_, new_n470_ );
and g0270 ( new_n472_, new_n463_, new_n469_ );
or g0271 ( new_n473_, new_n471_, new_n472_ );
and g0272 ( new_n474_, new_n453_, new_n473_ );
not g0273 ( new_n475_, new_n474_ );
or g0274 ( new_n476_, new_n453_, new_n473_ );
and g0275 ( new_n477_, new_n475_, new_n476_ );
or g0276 ( new_n478_, new_n477_, keyIn_0_58 );
and g0277 ( new_n479_, new_n477_, keyIn_0_58 );
not g0278 ( new_n480_, new_n479_ );
and g0279 ( new_n481_, new_n480_, new_n478_ );
not g0280 ( new_n482_, keyIn_0_56 );
not g0281 ( new_n483_, keyIn_0_48 );
and g0282 ( new_n484_, new_n338_, new_n435_ );
and g0283 ( new_n485_, new_n437_, new_n336_ );
or g0284 ( new_n486_, new_n484_, new_n485_ );
and g0285 ( new_n487_, new_n486_, keyIn_0_44 );
not g0286 ( new_n488_, new_n487_ );
or g0287 ( new_n489_, new_n486_, keyIn_0_44 );
and g0288 ( new_n490_, new_n488_, new_n489_ );
and g0289 ( new_n491_, N130, N137 );
not g0290 ( new_n492_, new_n491_ );
and g0291 ( new_n493_, new_n490_, new_n492_ );
not g0292 ( new_n494_, new_n493_ );
or g0293 ( new_n495_, new_n490_, new_n492_ );
and g0294 ( new_n496_, new_n494_, new_n495_ );
or g0295 ( new_n497_, new_n496_, new_n483_ );
and g0296 ( new_n498_, new_n496_, new_n483_ );
not g0297 ( new_n499_, new_n498_ );
and g0298 ( new_n500_, new_n499_, new_n497_ );
not g0299 ( new_n501_, N21 );
and g0300 ( new_n502_, new_n501_, N5 );
not g0301 ( new_n503_, N5 );
and g0302 ( new_n504_, new_n503_, N21 );
or g0303 ( new_n505_, new_n502_, new_n504_ );
not g0304 ( new_n506_, N53 );
and g0305 ( new_n507_, new_n506_, N37 );
not g0306 ( new_n508_, N37 );
and g0307 ( new_n509_, new_n508_, N53 );
or g0308 ( new_n510_, new_n507_, new_n509_ );
not g0309 ( new_n511_, new_n510_ );
and g0310 ( new_n512_, new_n511_, new_n505_ );
not g0311 ( new_n513_, new_n512_ );
or g0312 ( new_n514_, new_n511_, new_n505_ );
and g0313 ( new_n515_, new_n513_, new_n514_ );
or g0314 ( new_n516_, new_n500_, new_n515_ );
and g0315 ( new_n517_, new_n500_, new_n515_ );
not g0316 ( new_n518_, new_n517_ );
and g0317 ( new_n519_, new_n518_, new_n516_ );
not g0318 ( new_n520_, new_n519_ );
and g0319 ( new_n521_, new_n520_, new_n482_ );
and g0320 ( new_n522_, new_n519_, keyIn_0_56 );
or g0321 ( new_n523_, new_n521_, new_n522_ );
and g0322 ( new_n524_, new_n481_, new_n523_ );
and g0323 ( new_n525_, new_n403_, new_n524_ );
not g0324 ( new_n526_, new_n525_ );
or g0325 ( new_n527_, new_n403_, new_n524_ );
or g0326 ( new_n528_, new_n481_, new_n523_ );
and g0327 ( new_n529_, new_n528_, new_n306_ );
and g0328 ( new_n530_, new_n527_, new_n529_ );
and g0329 ( new_n531_, new_n530_, new_n526_ );
and g0330 ( new_n532_, new_n401_, keyIn_0_57 );
and g0331 ( new_n533_, new_n397_, new_n308_ );
or g0332 ( new_n534_, new_n532_, new_n533_ );
and g0333 ( new_n535_, new_n534_, keyIn_0_63 );
not g0334 ( new_n536_, new_n535_ );
or g0335 ( new_n537_, new_n534_, keyIn_0_63 );
not g0336 ( new_n538_, keyIn_0_58 );
not g0337 ( new_n539_, new_n477_ );
and g0338 ( new_n540_, new_n539_, new_n538_ );
or g0339 ( new_n541_, new_n540_, new_n479_ );
not g0340 ( new_n542_, new_n523_ );
or g0341 ( new_n543_, new_n306_, new_n542_ );
or g0342 ( new_n544_, new_n543_, new_n541_ );
not g0343 ( new_n545_, new_n544_ );
and g0344 ( new_n546_, new_n545_, new_n537_ );
and g0345 ( new_n547_, new_n546_, new_n536_ );
or g0346 ( new_n548_, new_n547_, new_n531_ );
not g0347 ( new_n549_, keyIn_0_28 );
not g0348 ( new_n550_, keyIn_0_0 );
or g0349 ( new_n551_, new_n284_, N5 );
or g0350 ( new_n552_, new_n503_, N1 );
and g0351 ( new_n553_, new_n551_, new_n552_ );
or g0352 ( new_n554_, new_n553_, new_n550_ );
and g0353 ( new_n555_, new_n503_, N1 );
and g0354 ( new_n556_, new_n284_, N5 );
or g0355 ( new_n557_, new_n555_, new_n556_ );
or g0356 ( new_n558_, new_n557_, keyIn_0_0 );
and g0357 ( new_n559_, new_n558_, new_n554_ );
not g0358 ( new_n560_, keyIn_0_1 );
or g0359 ( new_n561_, new_n362_, N13 );
or g0360 ( new_n562_, new_n457_, N9 );
and g0361 ( new_n563_, new_n561_, new_n562_ );
and g0362 ( new_n564_, new_n563_, new_n560_ );
and g0363 ( new_n565_, new_n457_, N9 );
and g0364 ( new_n566_, new_n362_, N13 );
or g0365 ( new_n567_, new_n565_, new_n566_ );
and g0366 ( new_n568_, new_n567_, keyIn_0_1 );
or g0367 ( new_n569_, new_n568_, new_n564_ );
or g0368 ( new_n570_, new_n569_, new_n559_ );
and g0369 ( new_n571_, new_n557_, keyIn_0_0 );
and g0370 ( new_n572_, new_n553_, new_n550_ );
or g0371 ( new_n573_, new_n571_, new_n572_ );
or g0372 ( new_n574_, new_n567_, keyIn_0_1 );
or g0373 ( new_n575_, new_n563_, new_n560_ );
and g0374 ( new_n576_, new_n574_, new_n575_ );
or g0375 ( new_n577_, new_n573_, new_n576_ );
and g0376 ( new_n578_, new_n570_, new_n577_ );
or g0377 ( new_n579_, new_n578_, new_n549_ );
and g0378 ( new_n580_, new_n573_, new_n576_ );
and g0379 ( new_n581_, new_n569_, new_n559_ );
or g0380 ( new_n582_, new_n580_, new_n581_ );
or g0381 ( new_n583_, new_n582_, keyIn_0_28 );
and g0382 ( new_n584_, new_n579_, new_n583_ );
not g0383 ( new_n585_, keyIn_0_29 );
or g0384 ( new_n586_, new_n282_, N21 );
or g0385 ( new_n587_, new_n501_, N17 );
and g0386 ( new_n588_, new_n586_, new_n587_ );
or g0387 ( new_n589_, new_n588_, keyIn_0_2 );
not g0388 ( new_n590_, keyIn_0_2 );
and g0389 ( new_n591_, new_n501_, N17 );
and g0390 ( new_n592_, new_n282_, N21 );
or g0391 ( new_n593_, new_n591_, new_n592_ );
or g0392 ( new_n594_, new_n593_, new_n590_ );
and g0393 ( new_n595_, new_n594_, new_n589_ );
not g0394 ( new_n596_, keyIn_0_3 );
or g0395 ( new_n597_, new_n360_, N29 );
or g0396 ( new_n598_, new_n455_, N25 );
and g0397 ( new_n599_, new_n597_, new_n598_ );
and g0398 ( new_n600_, new_n599_, new_n596_ );
and g0399 ( new_n601_, new_n455_, N25 );
and g0400 ( new_n602_, new_n360_, N29 );
or g0401 ( new_n603_, new_n601_, new_n602_ );
and g0402 ( new_n604_, new_n603_, keyIn_0_3 );
or g0403 ( new_n605_, new_n604_, new_n600_ );
or g0404 ( new_n606_, new_n605_, new_n595_ );
and g0405 ( new_n607_, new_n593_, new_n590_ );
and g0406 ( new_n608_, new_n588_, keyIn_0_2 );
or g0407 ( new_n609_, new_n607_, new_n608_ );
or g0408 ( new_n610_, new_n603_, keyIn_0_3 );
or g0409 ( new_n611_, new_n599_, new_n596_ );
and g0410 ( new_n612_, new_n610_, new_n611_ );
or g0411 ( new_n613_, new_n609_, new_n612_ );
and g0412 ( new_n614_, new_n606_, new_n613_ );
or g0413 ( new_n615_, new_n614_, new_n585_ );
and g0414 ( new_n616_, new_n609_, new_n612_ );
and g0415 ( new_n617_, new_n605_, new_n595_ );
or g0416 ( new_n618_, new_n616_, new_n617_ );
or g0417 ( new_n619_, new_n618_, keyIn_0_29 );
and g0418 ( new_n620_, new_n615_, new_n619_ );
or g0419 ( new_n621_, new_n584_, new_n620_ );
and g0420 ( new_n622_, new_n582_, keyIn_0_28 );
and g0421 ( new_n623_, new_n578_, new_n549_ );
or g0422 ( new_n624_, new_n622_, new_n623_ );
and g0423 ( new_n625_, new_n618_, keyIn_0_29 );
and g0424 ( new_n626_, new_n614_, new_n585_ );
or g0425 ( new_n627_, new_n625_, new_n626_ );
or g0426 ( new_n628_, new_n624_, new_n627_ );
and g0427 ( new_n629_, new_n628_, new_n621_ );
or g0428 ( new_n630_, new_n629_, keyIn_0_39 );
not g0429 ( new_n631_, keyIn_0_39 );
and g0430 ( new_n632_, new_n624_, new_n627_ );
and g0431 ( new_n633_, new_n584_, new_n620_ );
or g0432 ( new_n634_, new_n632_, new_n633_ );
or g0433 ( new_n635_, new_n634_, new_n631_ );
and g0434 ( new_n636_, new_n630_, new_n635_ );
not g0435 ( new_n637_, keyIn_0_17 );
and g0436 ( new_n638_, N133, N137 );
or g0437 ( new_n639_, new_n638_, new_n637_ );
and g0438 ( new_n640_, new_n637_, N133 );
and g0439 ( new_n641_, new_n640_, N137 );
not g0440 ( new_n642_, new_n641_ );
and g0441 ( new_n643_, new_n642_, new_n639_ );
or g0442 ( new_n644_, new_n636_, new_n643_ );
and g0443 ( new_n645_, new_n634_, new_n631_ );
and g0444 ( new_n646_, new_n629_, keyIn_0_39 );
or g0445 ( new_n647_, new_n646_, new_n645_ );
not g0446 ( new_n648_, new_n643_ );
or g0447 ( new_n649_, new_n647_, new_n648_ );
and g0448 ( new_n650_, new_n649_, new_n644_ );
or g0449 ( new_n651_, new_n650_, keyIn_0_51 );
not g0450 ( new_n652_, keyIn_0_51 );
and g0451 ( new_n653_, new_n647_, new_n648_ );
and g0452 ( new_n654_, new_n636_, new_n643_ );
or g0453 ( new_n655_, new_n653_, new_n654_ );
or g0454 ( new_n656_, new_n655_, new_n652_ );
and g0455 ( new_n657_, new_n656_, new_n651_ );
and g0456 ( new_n658_, new_n235_, N65 );
and g0457 ( new_n659_, new_n206_, N81 );
or g0458 ( new_n660_, new_n658_, new_n659_ );
and g0459 ( new_n661_, new_n410_, N97 );
and g0460 ( new_n662_, new_n311_, N113 );
or g0461 ( new_n663_, new_n661_, new_n662_ );
not g0462 ( new_n664_, new_n663_ );
and g0463 ( new_n665_, new_n664_, new_n660_ );
not g0464 ( new_n666_, new_n665_ );
or g0465 ( new_n667_, new_n664_, new_n660_ );
and g0466 ( new_n668_, new_n666_, new_n667_ );
or g0467 ( new_n669_, new_n657_, new_n668_ );
and g0468 ( new_n670_, new_n655_, new_n652_ );
and g0469 ( new_n671_, new_n650_, keyIn_0_51 );
or g0470 ( new_n672_, new_n670_, new_n671_ );
not g0471 ( new_n673_, new_n668_ );
or g0472 ( new_n674_, new_n672_, new_n673_ );
and g0473 ( new_n675_, new_n674_, new_n669_ );
or g0474 ( new_n676_, new_n675_, keyIn_0_59 );
not g0475 ( new_n677_, keyIn_0_59 );
and g0476 ( new_n678_, new_n672_, new_n673_ );
and g0477 ( new_n679_, new_n657_, new_n668_ );
or g0478 ( new_n680_, new_n678_, new_n679_ );
or g0479 ( new_n681_, new_n680_, new_n677_ );
and g0480 ( new_n682_, new_n681_, new_n676_ );
not g0481 ( new_n683_, keyIn_0_61 );
not g0482 ( new_n684_, keyIn_0_53 );
not g0483 ( new_n685_, keyIn_0_41 );
not g0484 ( new_n686_, keyIn_0_30 );
and g0485 ( new_n687_, new_n508_, N33 );
and g0486 ( new_n688_, new_n289_, N37 );
or g0487 ( new_n689_, new_n687_, new_n688_ );
and g0488 ( new_n690_, new_n689_, keyIn_0_4 );
not g0489 ( new_n691_, keyIn_0_4 );
or g0490 ( new_n692_, new_n289_, N37 );
or g0491 ( new_n693_, new_n508_, N33 );
and g0492 ( new_n694_, new_n692_, new_n693_ );
and g0493 ( new_n695_, new_n694_, new_n691_ );
or g0494 ( new_n696_, new_n690_, new_n695_ );
and g0495 ( new_n697_, new_n467_, N41 );
and g0496 ( new_n698_, new_n372_, N45 );
or g0497 ( new_n699_, new_n697_, new_n698_ );
and g0498 ( new_n700_, new_n699_, keyIn_0_5 );
not g0499 ( new_n701_, keyIn_0_5 );
or g0500 ( new_n702_, new_n372_, N45 );
or g0501 ( new_n703_, new_n467_, N41 );
and g0502 ( new_n704_, new_n702_, new_n703_ );
and g0503 ( new_n705_, new_n704_, new_n701_ );
or g0504 ( new_n706_, new_n700_, new_n705_ );
and g0505 ( new_n707_, new_n696_, new_n706_ );
or g0506 ( new_n708_, new_n694_, new_n691_ );
or g0507 ( new_n709_, new_n689_, keyIn_0_4 );
and g0508 ( new_n710_, new_n709_, new_n708_ );
or g0509 ( new_n711_, new_n704_, new_n701_ );
or g0510 ( new_n712_, new_n699_, keyIn_0_5 );
and g0511 ( new_n713_, new_n712_, new_n711_ );
and g0512 ( new_n714_, new_n710_, new_n713_ );
or g0513 ( new_n715_, new_n707_, new_n714_ );
and g0514 ( new_n716_, new_n715_, new_n686_ );
or g0515 ( new_n717_, new_n710_, new_n713_ );
or g0516 ( new_n718_, new_n696_, new_n706_ );
and g0517 ( new_n719_, new_n718_, new_n717_ );
and g0518 ( new_n720_, new_n719_, keyIn_0_30 );
or g0519 ( new_n721_, new_n716_, new_n720_ );
or g0520 ( new_n722_, new_n721_, new_n584_ );
or g0521 ( new_n723_, new_n719_, keyIn_0_30 );
or g0522 ( new_n724_, new_n715_, new_n686_ );
and g0523 ( new_n725_, new_n723_, new_n724_ );
or g0524 ( new_n726_, new_n624_, new_n725_ );
and g0525 ( new_n727_, new_n722_, new_n726_ );
or g0526 ( new_n728_, new_n727_, new_n685_ );
and g0527 ( new_n729_, new_n624_, new_n725_ );
and g0528 ( new_n730_, new_n721_, new_n584_ );
or g0529 ( new_n731_, new_n729_, new_n730_ );
or g0530 ( new_n732_, new_n731_, keyIn_0_41 );
and g0531 ( new_n733_, new_n732_, new_n728_ );
not g0532 ( new_n734_, keyIn_0_19 );
and g0533 ( new_n735_, N135, N137 );
or g0534 ( new_n736_, new_n735_, new_n734_ );
and g0535 ( new_n737_, new_n734_, N135 );
and g0536 ( new_n738_, new_n737_, N137 );
not g0537 ( new_n739_, new_n738_ );
and g0538 ( new_n740_, new_n739_, new_n736_ );
or g0539 ( new_n741_, new_n733_, new_n740_ );
and g0540 ( new_n742_, new_n731_, keyIn_0_41 );
and g0541 ( new_n743_, new_n727_, new_n685_ );
or g0542 ( new_n744_, new_n742_, new_n743_ );
not g0543 ( new_n745_, new_n740_ );
or g0544 ( new_n746_, new_n744_, new_n745_ );
and g0545 ( new_n747_, new_n746_, new_n741_ );
or g0546 ( new_n748_, new_n747_, new_n684_ );
and g0547 ( new_n749_, new_n744_, new_n745_ );
and g0548 ( new_n750_, new_n733_, new_n740_ );
or g0549 ( new_n751_, new_n749_, new_n750_ );
or g0550 ( new_n752_, new_n751_, keyIn_0_53 );
and g0551 ( new_n753_, new_n752_, new_n748_ );
not g0552 ( new_n754_, keyIn_0_26 );
and g0553 ( new_n755_, new_n245_, N73 );
and g0554 ( new_n756_, new_n217_, N89 );
or g0555 ( new_n757_, new_n755_, new_n756_ );
and g0556 ( new_n758_, new_n757_, new_n754_ );
not g0557 ( new_n759_, new_n758_ );
or g0558 ( new_n760_, new_n757_, new_n754_ );
and g0559 ( new_n761_, new_n759_, new_n760_ );
not g0560 ( new_n762_, new_n761_ );
not g0561 ( new_n763_, keyIn_0_27 );
and g0562 ( new_n764_, new_n421_, N105 );
and g0563 ( new_n765_, new_n322_, N121 );
or g0564 ( new_n766_, new_n764_, new_n765_ );
and g0565 ( new_n767_, new_n766_, new_n763_ );
not g0566 ( new_n768_, new_n767_ );
or g0567 ( new_n769_, new_n766_, new_n763_ );
and g0568 ( new_n770_, new_n768_, new_n769_ );
not g0569 ( new_n771_, new_n770_ );
and g0570 ( new_n772_, new_n762_, new_n771_ );
and g0571 ( new_n773_, new_n761_, new_n770_ );
or g0572 ( new_n774_, new_n772_, new_n773_ );
and g0573 ( new_n775_, new_n774_, keyIn_0_38 );
not g0574 ( new_n776_, new_n775_ );
or g0575 ( new_n777_, new_n774_, keyIn_0_38 );
and g0576 ( new_n778_, new_n776_, new_n777_ );
or g0577 ( new_n779_, new_n753_, new_n778_ );
and g0578 ( new_n780_, new_n751_, keyIn_0_53 );
and g0579 ( new_n781_, new_n747_, new_n684_ );
or g0580 ( new_n782_, new_n780_, new_n781_ );
not g0581 ( new_n783_, new_n778_ );
or g0582 ( new_n784_, new_n782_, new_n783_ );
and g0583 ( new_n785_, new_n784_, new_n779_ );
or g0584 ( new_n786_, new_n785_, new_n683_ );
and g0585 ( new_n787_, new_n782_, new_n783_ );
and g0586 ( new_n788_, new_n753_, new_n778_ );
or g0587 ( new_n789_, new_n787_, new_n788_ );
or g0588 ( new_n790_, new_n789_, keyIn_0_61 );
and g0589 ( new_n791_, new_n790_, new_n786_ );
not g0590 ( new_n792_, keyIn_0_31 );
not g0591 ( new_n793_, keyIn_0_6 );
and g0592 ( new_n794_, new_n506_, N49 );
and g0593 ( new_n795_, new_n287_, N53 );
or g0594 ( new_n796_, new_n794_, new_n795_ );
and g0595 ( new_n797_, new_n796_, new_n793_ );
or g0596 ( new_n798_, new_n287_, N53 );
or g0597 ( new_n799_, new_n506_, N49 );
and g0598 ( new_n800_, new_n798_, new_n799_ );
and g0599 ( new_n801_, new_n800_, keyIn_0_6 );
or g0600 ( new_n802_, new_n797_, new_n801_ );
and g0601 ( new_n803_, new_n465_, N57 );
and g0602 ( new_n804_, new_n370_, N61 );
or g0603 ( new_n805_, new_n803_, new_n804_ );
and g0604 ( new_n806_, new_n805_, keyIn_0_7 );
not g0605 ( new_n807_, keyIn_0_7 );
or g0606 ( new_n808_, new_n370_, N61 );
or g0607 ( new_n809_, new_n465_, N57 );
and g0608 ( new_n810_, new_n808_, new_n809_ );
and g0609 ( new_n811_, new_n810_, new_n807_ );
or g0610 ( new_n812_, new_n806_, new_n811_ );
and g0611 ( new_n813_, new_n802_, new_n812_ );
or g0612 ( new_n814_, new_n800_, keyIn_0_6 );
or g0613 ( new_n815_, new_n796_, new_n793_ );
and g0614 ( new_n816_, new_n815_, new_n814_ );
or g0615 ( new_n817_, new_n810_, new_n807_ );
or g0616 ( new_n818_, new_n805_, keyIn_0_7 );
and g0617 ( new_n819_, new_n818_, new_n817_ );
and g0618 ( new_n820_, new_n816_, new_n819_ );
or g0619 ( new_n821_, new_n813_, new_n820_ );
and g0620 ( new_n822_, new_n821_, new_n792_ );
or g0621 ( new_n823_, new_n816_, new_n819_ );
or g0622 ( new_n824_, new_n802_, new_n812_ );
and g0623 ( new_n825_, new_n824_, new_n823_ );
and g0624 ( new_n826_, new_n825_, keyIn_0_31 );
or g0625 ( new_n827_, new_n822_, new_n826_ );
and g0626 ( new_n828_, new_n721_, new_n827_ );
or g0627 ( new_n829_, new_n825_, keyIn_0_31 );
or g0628 ( new_n830_, new_n821_, new_n792_ );
and g0629 ( new_n831_, new_n829_, new_n830_ );
and g0630 ( new_n832_, new_n725_, new_n831_ );
or g0631 ( new_n833_, new_n828_, new_n832_ );
and g0632 ( new_n834_, new_n833_, keyIn_0_40 );
not g0633 ( new_n835_, keyIn_0_40 );
or g0634 ( new_n836_, new_n725_, new_n831_ );
or g0635 ( new_n837_, new_n721_, new_n827_ );
and g0636 ( new_n838_, new_n837_, new_n836_ );
and g0637 ( new_n839_, new_n838_, new_n835_ );
or g0638 ( new_n840_, new_n839_, new_n834_ );
not g0639 ( new_n841_, keyIn_0_18 );
and g0640 ( new_n842_, N134, N137 );
or g0641 ( new_n843_, new_n842_, new_n841_ );
and g0642 ( new_n844_, new_n841_, N134 );
and g0643 ( new_n845_, new_n844_, N137 );
not g0644 ( new_n846_, new_n845_ );
and g0645 ( new_n847_, new_n846_, new_n843_ );
not g0646 ( new_n848_, new_n847_ );
and g0647 ( new_n849_, new_n840_, new_n848_ );
or g0648 ( new_n850_, new_n838_, new_n835_ );
or g0649 ( new_n851_, new_n833_, keyIn_0_40 );
and g0650 ( new_n852_, new_n850_, new_n851_ );
and g0651 ( new_n853_, new_n852_, new_n847_ );
or g0652 ( new_n854_, new_n849_, new_n853_ );
and g0653 ( new_n855_, new_n854_, keyIn_0_52 );
not g0654 ( new_n856_, keyIn_0_52 );
or g0655 ( new_n857_, new_n852_, new_n847_ );
or g0656 ( new_n858_, new_n840_, new_n848_ );
and g0657 ( new_n859_, new_n858_, new_n857_ );
and g0658 ( new_n860_, new_n859_, new_n856_ );
or g0659 ( new_n861_, new_n855_, new_n860_ );
not g0660 ( new_n862_, keyIn_0_37 );
and g0661 ( new_n863_, new_n233_, N69 );
and g0662 ( new_n864_, new_n204_, N85 );
or g0663 ( new_n865_, new_n863_, new_n864_ );
and g0664 ( new_n866_, new_n865_, keyIn_0_24 );
not g0665 ( new_n867_, new_n866_ );
or g0666 ( new_n868_, new_n865_, keyIn_0_24 );
and g0667 ( new_n869_, new_n867_, new_n868_ );
not g0668 ( new_n870_, new_n869_ );
and g0669 ( new_n871_, new_n408_, N101 );
and g0670 ( new_n872_, new_n309_, N117 );
or g0671 ( new_n873_, new_n871_, new_n872_ );
and g0672 ( new_n874_, new_n873_, keyIn_0_25 );
not g0673 ( new_n875_, new_n874_ );
or g0674 ( new_n876_, new_n873_, keyIn_0_25 );
and g0675 ( new_n877_, new_n875_, new_n876_ );
not g0676 ( new_n878_, new_n877_ );
and g0677 ( new_n879_, new_n870_, new_n878_ );
and g0678 ( new_n880_, new_n869_, new_n877_ );
or g0679 ( new_n881_, new_n879_, new_n880_ );
and g0680 ( new_n882_, new_n881_, new_n862_ );
not g0681 ( new_n883_, new_n882_ );
or g0682 ( new_n884_, new_n881_, new_n862_ );
and g0683 ( new_n885_, new_n883_, new_n884_ );
and g0684 ( new_n886_, new_n861_, new_n885_ );
or g0685 ( new_n887_, new_n859_, new_n856_ );
or g0686 ( new_n888_, new_n854_, keyIn_0_52 );
and g0687 ( new_n889_, new_n888_, new_n887_ );
not g0688 ( new_n890_, new_n885_ );
and g0689 ( new_n891_, new_n889_, new_n890_ );
or g0690 ( new_n892_, new_n886_, new_n891_ );
and g0691 ( new_n893_, new_n892_, keyIn_0_60 );
not g0692 ( new_n894_, keyIn_0_60 );
or g0693 ( new_n895_, new_n889_, new_n890_ );
or g0694 ( new_n896_, new_n861_, new_n885_ );
and g0695 ( new_n897_, new_n896_, new_n895_ );
and g0696 ( new_n898_, new_n897_, new_n894_ );
or g0697 ( new_n899_, new_n893_, new_n898_ );
not g0698 ( new_n900_, keyIn_0_62 );
not g0699 ( new_n901_, keyIn_0_42 );
or g0700 ( new_n902_, new_n827_, new_n620_ );
or g0701 ( new_n903_, new_n627_, new_n831_ );
and g0702 ( new_n904_, new_n902_, new_n903_ );
or g0703 ( new_n905_, new_n904_, new_n901_ );
and g0704 ( new_n906_, new_n627_, new_n831_ );
and g0705 ( new_n907_, new_n827_, new_n620_ );
or g0706 ( new_n908_, new_n906_, new_n907_ );
or g0707 ( new_n909_, new_n908_, keyIn_0_42 );
and g0708 ( new_n910_, new_n909_, new_n905_ );
not g0709 ( new_n911_, keyIn_0_20 );
and g0710 ( new_n912_, N136, N137 );
or g0711 ( new_n913_, new_n912_, new_n911_ );
and g0712 ( new_n914_, new_n911_, N136 );
and g0713 ( new_n915_, new_n914_, N137 );
not g0714 ( new_n916_, new_n915_ );
and g0715 ( new_n917_, new_n916_, new_n913_ );
or g0716 ( new_n918_, new_n910_, new_n917_ );
and g0717 ( new_n919_, new_n908_, keyIn_0_42 );
and g0718 ( new_n920_, new_n904_, new_n901_ );
or g0719 ( new_n921_, new_n919_, new_n920_ );
not g0720 ( new_n922_, new_n917_ );
or g0721 ( new_n923_, new_n921_, new_n922_ );
and g0722 ( new_n924_, new_n923_, new_n918_ );
or g0723 ( new_n925_, new_n924_, keyIn_0_54 );
not g0724 ( new_n926_, keyIn_0_54 );
and g0725 ( new_n927_, new_n921_, new_n922_ );
and g0726 ( new_n928_, new_n910_, new_n917_ );
or g0727 ( new_n929_, new_n927_, new_n928_ );
or g0728 ( new_n930_, new_n929_, new_n926_ );
and g0729 ( new_n931_, new_n930_, new_n925_ );
and g0730 ( new_n932_, new_n243_, N77 );
and g0731 ( new_n933_, new_n215_, N93 );
or g0732 ( new_n934_, new_n932_, new_n933_ );
and g0733 ( new_n935_, new_n419_, N109 );
and g0734 ( new_n936_, new_n320_, N125 );
or g0735 ( new_n937_, new_n935_, new_n936_ );
not g0736 ( new_n938_, new_n937_ );
and g0737 ( new_n939_, new_n938_, new_n934_ );
not g0738 ( new_n940_, new_n939_ );
or g0739 ( new_n941_, new_n938_, new_n934_ );
and g0740 ( new_n942_, new_n940_, new_n941_ );
or g0741 ( new_n943_, new_n931_, new_n942_ );
and g0742 ( new_n944_, new_n929_, new_n926_ );
and g0743 ( new_n945_, new_n924_, keyIn_0_54 );
or g0744 ( new_n946_, new_n944_, new_n945_ );
not g0745 ( new_n947_, new_n942_ );
or g0746 ( new_n948_, new_n946_, new_n947_ );
and g0747 ( new_n949_, new_n948_, new_n943_ );
or g0748 ( new_n950_, new_n949_, new_n900_ );
and g0749 ( new_n951_, new_n946_, new_n947_ );
and g0750 ( new_n952_, new_n931_, new_n942_ );
or g0751 ( new_n953_, new_n951_, new_n952_ );
or g0752 ( new_n954_, new_n953_, keyIn_0_62 );
and g0753 ( new_n955_, new_n954_, new_n950_ );
and g0754 ( new_n956_, new_n899_, new_n955_ );
and g0755 ( new_n957_, new_n956_, new_n791_ );
and g0756 ( new_n958_, new_n957_, new_n682_ );
and g0757 ( new_n959_, new_n548_, new_n958_ );
and g0758 ( new_n960_, new_n959_, new_n307_ );
not g0759 ( new_n961_, new_n960_ );
and g0760 ( new_n962_, new_n961_, N1 );
and g0761 ( new_n963_, new_n960_, new_n284_ );
or g0762 ( N724, new_n962_, new_n963_ );
and g0763 ( new_n965_, new_n959_, new_n542_ );
not g0764 ( new_n966_, new_n965_ );
and g0765 ( new_n967_, new_n966_, N5 );
and g0766 ( new_n968_, new_n965_, new_n503_ );
or g0767 ( N725, new_n967_, new_n968_ );
and g0768 ( new_n970_, new_n959_, new_n534_ );
not g0769 ( new_n971_, new_n970_ );
and g0770 ( new_n972_, new_n971_, N9 );
and g0771 ( new_n973_, new_n970_, new_n362_ );
or g0772 ( N726, new_n972_, new_n973_ );
and g0773 ( new_n975_, new_n959_, new_n541_ );
not g0774 ( new_n976_, new_n975_ );
and g0775 ( new_n977_, new_n976_, N13 );
and g0776 ( new_n978_, new_n975_, new_n457_ );
or g0777 ( N727, new_n977_, new_n978_ );
not g0778 ( new_n980_, keyIn_0_105 );
not g0779 ( new_n981_, keyIn_0_82 );
not g0780 ( new_n982_, keyIn_0_76 );
and g0781 ( new_n983_, new_n789_, keyIn_0_61 );
and g0782 ( new_n984_, new_n785_, new_n683_ );
or g0783 ( new_n985_, new_n983_, new_n984_ );
and g0784 ( new_n986_, new_n953_, keyIn_0_62 );
and g0785 ( new_n987_, new_n949_, new_n900_ );
or g0786 ( new_n988_, new_n986_, new_n987_ );
and g0787 ( new_n989_, new_n985_, new_n988_ );
and g0788 ( new_n990_, new_n899_, new_n682_ );
and g0789 ( new_n991_, new_n989_, new_n990_ );
and g0790 ( new_n992_, new_n548_, new_n991_ );
or g0791 ( new_n993_, new_n992_, new_n982_ );
or g0792 ( new_n994_, new_n541_, new_n542_ );
and g0793 ( new_n995_, new_n994_, new_n534_ );
and g0794 ( new_n996_, new_n541_, new_n542_ );
or g0795 ( new_n997_, new_n996_, new_n307_ );
or g0796 ( new_n998_, new_n995_, new_n997_ );
or g0797 ( new_n999_, new_n998_, new_n525_ );
not g0798 ( new_n1000_, keyIn_0_63 );
and g0799 ( new_n1001_, new_n403_, new_n1000_ );
or g0800 ( new_n1002_, new_n1001_, new_n544_ );
or g0801 ( new_n1003_, new_n1002_, new_n535_ );
and g0802 ( new_n1004_, new_n999_, new_n1003_ );
not g0803 ( new_n1005_, new_n991_ );
or g0804 ( new_n1006_, new_n1004_, new_n1005_ );
or g0805 ( new_n1007_, new_n1006_, keyIn_0_76 );
and g0806 ( new_n1008_, new_n1007_, new_n993_ );
and g0807 ( new_n1009_, new_n1008_, new_n307_ );
or g0808 ( new_n1010_, new_n1009_, new_n981_ );
and g0809 ( new_n1011_, new_n1006_, keyIn_0_76 );
and g0810 ( new_n1012_, new_n992_, new_n982_ );
or g0811 ( new_n1013_, new_n1011_, new_n1012_ );
or g0812 ( new_n1014_, new_n1013_, new_n306_ );
or g0813 ( new_n1015_, new_n1014_, keyIn_0_82 );
and g0814 ( new_n1016_, new_n1015_, new_n1010_ );
or g0815 ( new_n1017_, new_n1016_, N17 );
and g0816 ( new_n1018_, new_n1014_, keyIn_0_82 );
and g0817 ( new_n1019_, new_n1009_, new_n981_ );
or g0818 ( new_n1020_, new_n1018_, new_n1019_ );
or g0819 ( new_n1021_, new_n1020_, new_n282_ );
and g0820 ( new_n1022_, new_n1021_, new_n1017_ );
or g0821 ( new_n1023_, new_n1022_, new_n980_ );
and g0822 ( new_n1024_, new_n1020_, new_n282_ );
and g0823 ( new_n1025_, new_n1016_, N17 );
or g0824 ( new_n1026_, new_n1024_, new_n1025_ );
or g0825 ( new_n1027_, new_n1026_, keyIn_0_105 );
and g0826 ( N728, new_n1027_, new_n1023_ );
and g0827 ( new_n1029_, new_n1008_, new_n542_ );
or g0828 ( new_n1030_, new_n1029_, keyIn_0_83 );
not g0829 ( new_n1031_, keyIn_0_83 );
or g0830 ( new_n1032_, new_n1013_, new_n523_ );
or g0831 ( new_n1033_, new_n1032_, new_n1031_ );
and g0832 ( new_n1034_, new_n1033_, new_n1030_ );
or g0833 ( new_n1035_, new_n1034_, new_n501_ );
and g0834 ( new_n1036_, new_n1032_, new_n1031_ );
and g0835 ( new_n1037_, new_n1029_, keyIn_0_83 );
or g0836 ( new_n1038_, new_n1036_, new_n1037_ );
or g0837 ( new_n1039_, new_n1038_, N21 );
and g0838 ( new_n1040_, new_n1039_, new_n1035_ );
or g0839 ( new_n1041_, new_n1040_, keyIn_0_106 );
not g0840 ( new_n1042_, keyIn_0_106 );
and g0841 ( new_n1043_, new_n1038_, N21 );
and g0842 ( new_n1044_, new_n1034_, new_n501_ );
or g0843 ( new_n1045_, new_n1043_, new_n1044_ );
or g0844 ( new_n1046_, new_n1045_, new_n1042_ );
and g0845 ( N729, new_n1046_, new_n1041_ );
and g0846 ( new_n1048_, new_n1008_, new_n534_ );
not g0847 ( new_n1049_, new_n1048_ );
and g0848 ( new_n1050_, new_n1049_, N25 );
and g0849 ( new_n1051_, new_n1048_, new_n360_ );
or g0850 ( N730, new_n1050_, new_n1051_ );
and g0851 ( new_n1053_, new_n1008_, new_n541_ );
or g0852 ( new_n1054_, new_n1053_, keyIn_0_84 );
not g0853 ( new_n1055_, keyIn_0_84 );
or g0854 ( new_n1056_, new_n1013_, new_n481_ );
or g0855 ( new_n1057_, new_n1056_, new_n1055_ );
and g0856 ( new_n1058_, new_n1057_, new_n1054_ );
or g0857 ( new_n1059_, new_n1058_, N29 );
and g0858 ( new_n1060_, new_n1056_, new_n1055_ );
and g0859 ( new_n1061_, new_n1053_, keyIn_0_84 );
or g0860 ( new_n1062_, new_n1060_, new_n1061_ );
or g0861 ( new_n1063_, new_n1062_, new_n455_ );
and g0862 ( new_n1064_, new_n1063_, new_n1059_ );
or g0863 ( new_n1065_, new_n1064_, keyIn_0_107 );
not g0864 ( new_n1066_, keyIn_0_107 );
and g0865 ( new_n1067_, new_n1062_, new_n455_ );
and g0866 ( new_n1068_, new_n1058_, N29 );
or g0867 ( new_n1069_, new_n1067_, new_n1068_ );
or g0868 ( new_n1070_, new_n1069_, new_n1066_ );
and g0869 ( N731, new_n1070_, new_n1065_ );
not g0870 ( new_n1072_, keyIn_0_108 );
not g0871 ( new_n1073_, keyIn_0_77 );
or g0872 ( new_n1074_, new_n897_, new_n894_ );
or g0873 ( new_n1075_, new_n892_, keyIn_0_60 );
and g0874 ( new_n1076_, new_n1075_, new_n1074_ );
and g0875 ( new_n1077_, new_n680_, new_n677_ );
and g0876 ( new_n1078_, new_n675_, keyIn_0_59 );
or g0877 ( new_n1079_, new_n1077_, new_n1078_ );
and g0878 ( new_n1080_, new_n1079_, new_n791_ );
and g0879 ( new_n1081_, new_n1080_, new_n955_ );
and g0880 ( new_n1082_, new_n1081_, new_n1076_ );
and g0881 ( new_n1083_, new_n548_, new_n1082_ );
or g0882 ( new_n1084_, new_n1083_, new_n1073_ );
not g0883 ( new_n1085_, new_n1082_ );
or g0884 ( new_n1086_, new_n1004_, new_n1085_ );
or g0885 ( new_n1087_, new_n1086_, keyIn_0_77 );
and g0886 ( new_n1088_, new_n1087_, new_n1084_ );
and g0887 ( new_n1089_, new_n1088_, new_n307_ );
or g0888 ( new_n1090_, new_n1089_, keyIn_0_85 );
not g0889 ( new_n1091_, keyIn_0_85 );
and g0890 ( new_n1092_, new_n1086_, keyIn_0_77 );
and g0891 ( new_n1093_, new_n1083_, new_n1073_ );
or g0892 ( new_n1094_, new_n1092_, new_n1093_ );
or g0893 ( new_n1095_, new_n1094_, new_n306_ );
or g0894 ( new_n1096_, new_n1095_, new_n1091_ );
and g0895 ( new_n1097_, new_n1096_, new_n1090_ );
or g0896 ( new_n1098_, new_n1097_, new_n289_ );
and g0897 ( new_n1099_, new_n1095_, new_n1091_ );
and g0898 ( new_n1100_, new_n1089_, keyIn_0_85 );
or g0899 ( new_n1101_, new_n1099_, new_n1100_ );
or g0900 ( new_n1102_, new_n1101_, N33 );
and g0901 ( new_n1103_, new_n1102_, new_n1098_ );
or g0902 ( new_n1104_, new_n1103_, new_n1072_ );
and g0903 ( new_n1105_, new_n1101_, N33 );
and g0904 ( new_n1106_, new_n1097_, new_n289_ );
or g0905 ( new_n1107_, new_n1105_, new_n1106_ );
or g0906 ( new_n1108_, new_n1107_, keyIn_0_108 );
and g0907 ( N732, new_n1108_, new_n1104_ );
not g0908 ( new_n1110_, keyIn_0_86 );
and g0909 ( new_n1111_, new_n1088_, new_n542_ );
or g0910 ( new_n1112_, new_n1111_, new_n1110_ );
or g0911 ( new_n1113_, new_n1094_, new_n523_ );
or g0912 ( new_n1114_, new_n1113_, keyIn_0_86 );
and g0913 ( new_n1115_, new_n1114_, new_n1112_ );
or g0914 ( new_n1116_, new_n1115_, new_n508_ );
and g0915 ( new_n1117_, new_n1113_, keyIn_0_86 );
and g0916 ( new_n1118_, new_n1111_, new_n1110_ );
or g0917 ( new_n1119_, new_n1117_, new_n1118_ );
or g0918 ( new_n1120_, new_n1119_, N37 );
and g0919 ( new_n1121_, new_n1120_, new_n1116_ );
or g0920 ( new_n1122_, new_n1121_, keyIn_0_109 );
not g0921 ( new_n1123_, keyIn_0_109 );
and g0922 ( new_n1124_, new_n1119_, N37 );
and g0923 ( new_n1125_, new_n1115_, new_n508_ );
or g0924 ( new_n1126_, new_n1124_, new_n1125_ );
or g0925 ( new_n1127_, new_n1126_, new_n1123_ );
and g0926 ( N733, new_n1127_, new_n1122_ );
not g0927 ( new_n1129_, keyIn_0_110 );
or g0928 ( new_n1130_, new_n1094_, new_n403_ );
and g0929 ( new_n1131_, new_n1130_, keyIn_0_87 );
not g0930 ( new_n1132_, keyIn_0_87 );
and g0931 ( new_n1133_, new_n1088_, new_n534_ );
and g0932 ( new_n1134_, new_n1133_, new_n1132_ );
or g0933 ( new_n1135_, new_n1131_, new_n1134_ );
and g0934 ( new_n1136_, new_n1135_, new_n372_ );
or g0935 ( new_n1137_, new_n1133_, new_n1132_ );
or g0936 ( new_n1138_, new_n1130_, keyIn_0_87 );
and g0937 ( new_n1139_, new_n1138_, new_n1137_ );
and g0938 ( new_n1140_, new_n1139_, N41 );
or g0939 ( new_n1141_, new_n1136_, new_n1140_ );
and g0940 ( new_n1142_, new_n1141_, new_n1129_ );
or g0941 ( new_n1143_, new_n1139_, N41 );
or g0942 ( new_n1144_, new_n1135_, new_n372_ );
and g0943 ( new_n1145_, new_n1144_, new_n1143_ );
and g0944 ( new_n1146_, new_n1145_, keyIn_0_110 );
or g0945 ( N734, new_n1142_, new_n1146_ );
not g0946 ( new_n1148_, keyIn_0_111 );
not g0947 ( new_n1149_, keyIn_0_88 );
and g0948 ( new_n1150_, new_n1088_, new_n541_ );
or g0949 ( new_n1151_, new_n1150_, new_n1149_ );
or g0950 ( new_n1152_, new_n1094_, new_n481_ );
or g0951 ( new_n1153_, new_n1152_, keyIn_0_88 );
and g0952 ( new_n1154_, new_n1153_, new_n1151_ );
or g0953 ( new_n1155_, new_n1154_, N45 );
and g0954 ( new_n1156_, new_n1152_, keyIn_0_88 );
and g0955 ( new_n1157_, new_n1150_, new_n1149_ );
or g0956 ( new_n1158_, new_n1156_, new_n1157_ );
or g0957 ( new_n1159_, new_n1158_, new_n467_ );
and g0958 ( new_n1160_, new_n1159_, new_n1155_ );
or g0959 ( new_n1161_, new_n1160_, new_n1148_ );
and g0960 ( new_n1162_, new_n1158_, new_n467_ );
and g0961 ( new_n1163_, new_n1154_, N45 );
or g0962 ( new_n1164_, new_n1162_, new_n1163_ );
or g0963 ( new_n1165_, new_n1164_, keyIn_0_111 );
and g0964 ( N735, new_n1165_, new_n1161_ );
and g0965 ( new_n1167_, new_n1079_, new_n1076_ );
and g0966 ( new_n1168_, new_n989_, new_n1167_ );
and g0967 ( new_n1169_, new_n548_, new_n1168_ );
and g0968 ( new_n1170_, new_n1169_, new_n307_ );
not g0969 ( new_n1171_, new_n1170_ );
and g0970 ( new_n1172_, new_n1171_, N49 );
and g0971 ( new_n1173_, new_n1170_, new_n287_ );
or g0972 ( N736, new_n1172_, new_n1173_ );
and g0973 ( new_n1175_, new_n1169_, new_n542_ );
not g0974 ( new_n1176_, new_n1175_ );
and g0975 ( new_n1177_, new_n1176_, N53 );
and g0976 ( new_n1178_, new_n1175_, new_n506_ );
or g0977 ( N737, new_n1177_, new_n1178_ );
and g0978 ( new_n1180_, new_n1169_, new_n534_ );
not g0979 ( new_n1181_, new_n1180_ );
and g0980 ( new_n1182_, new_n1181_, N57 );
and g0981 ( new_n1183_, new_n1180_, new_n370_ );
or g0982 ( N738, new_n1182_, new_n1183_ );
and g0983 ( new_n1185_, new_n1169_, new_n541_ );
not g0984 ( new_n1186_, new_n1185_ );
and g0985 ( new_n1187_, new_n1186_, N61 );
and g0986 ( new_n1188_, new_n1185_, new_n465_ );
or g0987 ( N739, new_n1187_, new_n1188_ );
not g0988 ( new_n1190_, keyIn_0_112 );
not g0989 ( new_n1191_, keyIn_0_78 );
not g0990 ( new_n1192_, keyIn_0_75 );
not g0991 ( new_n1193_, keyIn_0_71 );
and g0992 ( new_n1194_, new_n1079_, new_n899_ );
and g0993 ( new_n1195_, new_n1194_, new_n988_ );
or g0994 ( new_n1196_, new_n791_, keyIn_0_64 );
and g0995 ( new_n1197_, new_n791_, keyIn_0_64 );
not g0996 ( new_n1198_, new_n1197_ );
and g0997 ( new_n1199_, new_n1198_, new_n1196_ );
and g0998 ( new_n1200_, new_n1199_, new_n1195_ );
or g0999 ( new_n1201_, new_n1200_, new_n1193_ );
or g1000 ( new_n1202_, new_n682_, new_n1076_ );
or g1001 ( new_n1203_, new_n1202_, new_n955_ );
not g1002 ( new_n1204_, keyIn_0_64 );
and g1003 ( new_n1205_, new_n985_, new_n1204_ );
or g1004 ( new_n1206_, new_n1205_, new_n1197_ );
or g1005 ( new_n1207_, new_n1203_, new_n1206_ );
or g1006 ( new_n1208_, new_n1207_, keyIn_0_71 );
and g1007 ( new_n1209_, new_n1201_, new_n1208_ );
not g1008 ( new_n1210_, keyIn_0_65 );
or g1009 ( new_n1211_, new_n791_, new_n1210_ );
or g1010 ( new_n1212_, new_n985_, keyIn_0_65 );
and g1011 ( new_n1213_, new_n1212_, new_n1211_ );
or g1012 ( new_n1214_, new_n899_, new_n682_ );
or g1013 ( new_n1215_, new_n1214_, new_n988_ );
or g1014 ( new_n1216_, new_n1215_, new_n1213_ );
and g1015 ( new_n1217_, new_n1216_, keyIn_0_73 );
not g1016 ( new_n1218_, keyIn_0_73 );
and g1017 ( new_n1219_, new_n985_, keyIn_0_65 );
and g1018 ( new_n1220_, new_n791_, new_n1210_ );
or g1019 ( new_n1221_, new_n1219_, new_n1220_ );
and g1020 ( new_n1222_, new_n1167_, new_n955_ );
and g1021 ( new_n1223_, new_n1221_, new_n1222_ );
and g1022 ( new_n1224_, new_n1223_, new_n1218_ );
or g1023 ( new_n1225_, new_n1217_, new_n1224_ );
or g1024 ( new_n1226_, new_n1209_, new_n1225_ );
not g1025 ( new_n1227_, keyIn_0_74 );
and g1026 ( new_n1228_, new_n985_, keyIn_0_66 );
not g1027 ( new_n1229_, keyIn_0_66 );
and g1028 ( new_n1230_, new_n791_, new_n1229_ );
or g1029 ( new_n1231_, new_n1228_, new_n1230_ );
and g1030 ( new_n1232_, new_n956_, new_n682_ );
and g1031 ( new_n1233_, new_n1231_, new_n1232_ );
or g1032 ( new_n1234_, new_n1233_, new_n1227_ );
or g1033 ( new_n1235_, new_n791_, new_n1229_ );
or g1034 ( new_n1236_, new_n985_, keyIn_0_66 );
and g1035 ( new_n1237_, new_n1236_, new_n1235_ );
or g1036 ( new_n1238_, new_n988_, new_n1076_ );
or g1037 ( new_n1239_, new_n1238_, new_n1079_ );
or g1038 ( new_n1240_, new_n1239_, new_n1237_ );
or g1039 ( new_n1241_, new_n1240_, keyIn_0_74 );
and g1040 ( new_n1242_, new_n1241_, new_n1234_ );
not g1041 ( new_n1243_, keyIn_0_72 );
and g1042 ( new_n1244_, new_n1079_, new_n1243_ );
and g1043 ( new_n1245_, new_n957_, new_n1244_ );
not g1044 ( new_n1246_, new_n1245_ );
and g1045 ( new_n1247_, new_n1081_, new_n899_ );
or g1046 ( new_n1248_, new_n1247_, new_n1243_ );
and g1047 ( new_n1249_, new_n1248_, new_n1246_ );
or g1048 ( new_n1250_, new_n1242_, new_n1249_ );
or g1049 ( new_n1251_, new_n1226_, new_n1250_ );
and g1050 ( new_n1252_, new_n1251_, new_n1192_ );
and g1051 ( new_n1253_, new_n1207_, keyIn_0_71 );
and g1052 ( new_n1254_, new_n1200_, new_n1193_ );
or g1053 ( new_n1255_, new_n1254_, new_n1253_ );
or g1054 ( new_n1256_, new_n1223_, new_n1218_ );
not g1055 ( new_n1257_, new_n1224_ );
and g1056 ( new_n1258_, new_n1257_, new_n1256_ );
and g1057 ( new_n1259_, new_n1258_, new_n1255_ );
and g1058 ( new_n1260_, new_n1240_, keyIn_0_74 );
and g1059 ( new_n1261_, new_n1233_, new_n1227_ );
or g1060 ( new_n1262_, new_n1260_, new_n1261_ );
not g1061 ( new_n1263_, new_n1249_ );
and g1062 ( new_n1264_, new_n1263_, new_n1262_ );
and g1063 ( new_n1265_, new_n1259_, new_n1264_ );
and g1064 ( new_n1266_, new_n1265_, keyIn_0_75 );
or g1065 ( new_n1267_, new_n1252_, new_n1266_ );
and g1066 ( new_n1268_, new_n542_, keyIn_0_67 );
not g1067 ( new_n1269_, new_n1268_ );
or g1068 ( new_n1270_, new_n542_, keyIn_0_67 );
and g1069 ( new_n1271_, new_n307_, new_n481_ );
and g1070 ( new_n1272_, new_n1271_, new_n1270_ );
and g1071 ( new_n1273_, new_n1272_, new_n1269_ );
and g1072 ( new_n1274_, new_n1273_, new_n534_ );
and g1073 ( new_n1275_, new_n1267_, new_n1274_ );
and g1074 ( new_n1276_, new_n1275_, new_n1191_ );
or g1075 ( new_n1277_, new_n1265_, keyIn_0_75 );
or g1076 ( new_n1278_, new_n1251_, new_n1192_ );
and g1077 ( new_n1279_, new_n1278_, new_n1277_ );
not g1078 ( new_n1280_, new_n1274_ );
or g1079 ( new_n1281_, new_n1279_, new_n1280_ );
and g1080 ( new_n1282_, new_n1281_, keyIn_0_78 );
or g1081 ( new_n1283_, new_n1282_, new_n1079_ );
or g1082 ( new_n1284_, new_n1283_, new_n1276_ );
and g1083 ( new_n1285_, new_n1284_, keyIn_0_89 );
not g1084 ( new_n1286_, keyIn_0_89 );
not g1085 ( new_n1287_, new_n1276_ );
or g1086 ( new_n1288_, new_n1275_, new_n1191_ );
and g1087 ( new_n1289_, new_n1288_, new_n682_ );
and g1088 ( new_n1290_, new_n1289_, new_n1287_ );
and g1089 ( new_n1291_, new_n1290_, new_n1286_ );
or g1090 ( new_n1292_, new_n1285_, new_n1291_ );
and g1091 ( new_n1293_, new_n1292_, new_n206_ );
or g1092 ( new_n1294_, new_n1290_, new_n1286_ );
or g1093 ( new_n1295_, new_n1284_, keyIn_0_89 );
and g1094 ( new_n1296_, new_n1295_, new_n1294_ );
and g1095 ( new_n1297_, new_n1296_, N65 );
or g1096 ( new_n1298_, new_n1293_, new_n1297_ );
and g1097 ( new_n1299_, new_n1298_, new_n1190_ );
or g1098 ( new_n1300_, new_n1296_, N65 );
or g1099 ( new_n1301_, new_n1292_, new_n206_ );
and g1100 ( new_n1302_, new_n1300_, new_n1301_ );
and g1101 ( new_n1303_, new_n1302_, keyIn_0_112 );
or g1102 ( N740, new_n1299_, new_n1303_ );
and g1103 ( new_n1305_, new_n1288_, new_n1076_ );
and g1104 ( new_n1306_, new_n1305_, new_n1287_ );
or g1105 ( new_n1307_, new_n1306_, keyIn_0_90 );
not g1106 ( new_n1308_, keyIn_0_90 );
or g1107 ( new_n1309_, new_n1282_, new_n899_ );
or g1108 ( new_n1310_, new_n1309_, new_n1276_ );
or g1109 ( new_n1311_, new_n1310_, new_n1308_ );
and g1110 ( new_n1312_, new_n1311_, new_n1307_ );
or g1111 ( new_n1313_, new_n1312_, N69 );
and g1112 ( new_n1314_, new_n1310_, new_n1308_ );
and g1113 ( new_n1315_, new_n1306_, keyIn_0_90 );
or g1114 ( new_n1316_, new_n1314_, new_n1315_ );
or g1115 ( new_n1317_, new_n1316_, new_n204_ );
and g1116 ( new_n1318_, new_n1313_, new_n1317_ );
or g1117 ( new_n1319_, new_n1318_, keyIn_0_113 );
not g1118 ( new_n1320_, keyIn_0_113 );
and g1119 ( new_n1321_, new_n1316_, new_n204_ );
and g1120 ( new_n1322_, new_n1312_, N69 );
or g1121 ( new_n1323_, new_n1321_, new_n1322_ );
or g1122 ( new_n1324_, new_n1323_, new_n1320_ );
and g1123 ( N741, new_n1324_, new_n1319_ );
not g1124 ( new_n1326_, keyIn_0_91 );
or g1125 ( new_n1327_, new_n1282_, new_n985_ );
or g1126 ( new_n1328_, new_n1327_, new_n1276_ );
and g1127 ( new_n1329_, new_n1328_, new_n1326_ );
and g1128 ( new_n1330_, new_n1288_, new_n791_ );
and g1129 ( new_n1331_, new_n1330_, new_n1287_ );
and g1130 ( new_n1332_, new_n1331_, keyIn_0_91 );
or g1131 ( new_n1333_, new_n1329_, new_n1332_ );
and g1132 ( new_n1334_, new_n1333_, new_n217_ );
or g1133 ( new_n1335_, new_n1331_, keyIn_0_91 );
or g1134 ( new_n1336_, new_n1328_, new_n1326_ );
and g1135 ( new_n1337_, new_n1336_, new_n1335_ );
and g1136 ( new_n1338_, new_n1337_, N73 );
or g1137 ( new_n1339_, new_n1334_, new_n1338_ );
and g1138 ( new_n1340_, new_n1339_, keyIn_0_114 );
not g1139 ( new_n1341_, keyIn_0_114 );
or g1140 ( new_n1342_, new_n1337_, N73 );
or g1141 ( new_n1343_, new_n1333_, new_n217_ );
and g1142 ( new_n1344_, new_n1342_, new_n1343_ );
and g1143 ( new_n1345_, new_n1344_, new_n1341_ );
or g1144 ( N742, new_n1340_, new_n1345_ );
or g1145 ( new_n1347_, new_n1282_, new_n955_ );
or g1146 ( new_n1348_, new_n1347_, new_n1276_ );
and g1147 ( new_n1349_, new_n1348_, keyIn_0_92 );
not g1148 ( new_n1350_, keyIn_0_92 );
and g1149 ( new_n1351_, new_n1288_, new_n988_ );
and g1150 ( new_n1352_, new_n1351_, new_n1287_ );
and g1151 ( new_n1353_, new_n1352_, new_n1350_ );
or g1152 ( new_n1354_, new_n1349_, new_n1353_ );
and g1153 ( new_n1355_, new_n1354_, new_n215_ );
or g1154 ( new_n1356_, new_n1352_, new_n1350_ );
or g1155 ( new_n1357_, new_n1348_, keyIn_0_92 );
and g1156 ( new_n1358_, new_n1357_, new_n1356_ );
and g1157 ( new_n1359_, new_n1358_, N77 );
or g1158 ( new_n1360_, new_n1355_, new_n1359_ );
and g1159 ( new_n1361_, new_n1360_, keyIn_0_115 );
not g1160 ( new_n1362_, keyIn_0_115 );
or g1161 ( new_n1363_, new_n1358_, N77 );
or g1162 ( new_n1364_, new_n1354_, new_n215_ );
and g1163 ( new_n1365_, new_n1363_, new_n1364_ );
and g1164 ( new_n1366_, new_n1365_, new_n1362_ );
or g1165 ( N743, new_n1361_, new_n1366_ );
not g1166 ( new_n1368_, keyIn_0_68 );
and g1167 ( new_n1369_, new_n534_, new_n1368_ );
not g1168 ( new_n1370_, new_n1369_ );
and g1169 ( new_n1371_, new_n403_, keyIn_0_68 );
not g1170 ( new_n1372_, new_n1371_ );
not g1171 ( new_n1373_, new_n543_ );
and g1172 ( new_n1374_, new_n1373_, new_n541_ );
and g1173 ( new_n1375_, new_n1372_, new_n1374_ );
and g1174 ( new_n1376_, new_n1375_, new_n1370_ );
and g1175 ( new_n1377_, new_n1267_, new_n1376_ );
and g1176 ( new_n1378_, new_n1377_, keyIn_0_79 );
not g1177 ( new_n1379_, new_n1378_ );
or g1178 ( new_n1380_, new_n1377_, keyIn_0_79 );
and g1179 ( new_n1381_, new_n1380_, new_n682_ );
and g1180 ( new_n1382_, new_n1381_, new_n1379_ );
or g1181 ( new_n1383_, new_n1382_, keyIn_0_93 );
not g1182 ( new_n1384_, keyIn_0_93 );
not g1183 ( new_n1385_, keyIn_0_79 );
not g1184 ( new_n1386_, new_n1376_ );
or g1185 ( new_n1387_, new_n1279_, new_n1386_ );
and g1186 ( new_n1388_, new_n1387_, new_n1385_ );
or g1187 ( new_n1389_, new_n1388_, new_n1079_ );
or g1188 ( new_n1390_, new_n1389_, new_n1378_ );
or g1189 ( new_n1391_, new_n1390_, new_n1384_ );
and g1190 ( new_n1392_, new_n1391_, new_n1383_ );
or g1191 ( new_n1393_, new_n1392_, N81 );
and g1192 ( new_n1394_, new_n1390_, new_n1384_ );
and g1193 ( new_n1395_, new_n1382_, keyIn_0_93 );
or g1194 ( new_n1396_, new_n1394_, new_n1395_ );
or g1195 ( new_n1397_, new_n1396_, new_n235_ );
and g1196 ( new_n1398_, new_n1393_, new_n1397_ );
or g1197 ( new_n1399_, new_n1398_, keyIn_0_116 );
not g1198 ( new_n1400_, keyIn_0_116 );
and g1199 ( new_n1401_, new_n1396_, new_n235_ );
and g1200 ( new_n1402_, new_n1392_, N81 );
or g1201 ( new_n1403_, new_n1401_, new_n1402_ );
or g1202 ( new_n1404_, new_n1403_, new_n1400_ );
and g1203 ( N744, new_n1404_, new_n1399_ );
not g1204 ( new_n1406_, keyIn_0_94 );
and g1205 ( new_n1407_, new_n1380_, new_n1076_ );
and g1206 ( new_n1408_, new_n1407_, new_n1379_ );
or g1207 ( new_n1409_, new_n1408_, new_n1406_ );
or g1208 ( new_n1410_, new_n1388_, new_n899_ );
or g1209 ( new_n1411_, new_n1410_, new_n1378_ );
or g1210 ( new_n1412_, new_n1411_, keyIn_0_94 );
and g1211 ( new_n1413_, new_n1412_, new_n1409_ );
or g1212 ( new_n1414_, new_n1413_, N85 );
and g1213 ( new_n1415_, new_n1411_, keyIn_0_94 );
and g1214 ( new_n1416_, new_n1408_, new_n1406_ );
or g1215 ( new_n1417_, new_n1415_, new_n1416_ );
or g1216 ( new_n1418_, new_n1417_, new_n233_ );
and g1217 ( new_n1419_, new_n1414_, new_n1418_ );
or g1218 ( new_n1420_, new_n1419_, keyIn_0_117 );
not g1219 ( new_n1421_, keyIn_0_117 );
and g1220 ( new_n1422_, new_n1417_, new_n233_ );
and g1221 ( new_n1423_, new_n1413_, N85 );
or g1222 ( new_n1424_, new_n1422_, new_n1423_ );
or g1223 ( new_n1425_, new_n1424_, new_n1421_ );
and g1224 ( N745, new_n1425_, new_n1420_ );
not g1225 ( new_n1427_, keyIn_0_95 );
and g1226 ( new_n1428_, new_n1380_, new_n791_ );
and g1227 ( new_n1429_, new_n1428_, new_n1379_ );
or g1228 ( new_n1430_, new_n1429_, new_n1427_ );
or g1229 ( new_n1431_, new_n1388_, new_n985_ );
or g1230 ( new_n1432_, new_n1431_, new_n1378_ );
or g1231 ( new_n1433_, new_n1432_, keyIn_0_95 );
and g1232 ( new_n1434_, new_n1433_, new_n1430_ );
or g1233 ( new_n1435_, new_n1434_, new_n245_ );
and g1234 ( new_n1436_, new_n1432_, keyIn_0_95 );
and g1235 ( new_n1437_, new_n1429_, new_n1427_ );
or g1236 ( new_n1438_, new_n1436_, new_n1437_ );
or g1237 ( new_n1439_, new_n1438_, N89 );
and g1238 ( new_n1440_, new_n1435_, new_n1439_ );
or g1239 ( new_n1441_, new_n1440_, keyIn_0_118 );
not g1240 ( new_n1442_, keyIn_0_118 );
and g1241 ( new_n1443_, new_n1438_, N89 );
and g1242 ( new_n1444_, new_n1434_, new_n245_ );
or g1243 ( new_n1445_, new_n1443_, new_n1444_ );
or g1244 ( new_n1446_, new_n1445_, new_n1442_ );
and g1245 ( N746, new_n1446_, new_n1441_ );
or g1246 ( new_n1448_, new_n1388_, new_n955_ );
or g1247 ( new_n1449_, new_n1448_, new_n1378_ );
and g1248 ( new_n1450_, new_n1449_, keyIn_0_96 );
not g1249 ( new_n1451_, keyIn_0_96 );
and g1250 ( new_n1452_, new_n1380_, new_n988_ );
and g1251 ( new_n1453_, new_n1452_, new_n1379_ );
and g1252 ( new_n1454_, new_n1453_, new_n1451_ );
or g1253 ( new_n1455_, new_n1450_, new_n1454_ );
and g1254 ( new_n1456_, new_n1455_, N93 );
or g1255 ( new_n1457_, new_n1453_, new_n1451_ );
or g1256 ( new_n1458_, new_n1449_, keyIn_0_96 );
and g1257 ( new_n1459_, new_n1458_, new_n1457_ );
and g1258 ( new_n1460_, new_n1459_, new_n243_ );
or g1259 ( new_n1461_, new_n1456_, new_n1460_ );
and g1260 ( new_n1462_, new_n1461_, keyIn_0_119 );
not g1261 ( new_n1463_, keyIn_0_119 );
or g1262 ( new_n1464_, new_n1459_, new_n243_ );
or g1263 ( new_n1465_, new_n1455_, N93 );
and g1264 ( new_n1466_, new_n1464_, new_n1465_ );
and g1265 ( new_n1467_, new_n1466_, new_n1463_ );
or g1266 ( N747, new_n1462_, new_n1467_ );
not g1267 ( new_n1469_, keyIn_0_97 );
not g1268 ( new_n1470_, keyIn_0_80 );
and g1269 ( new_n1471_, new_n481_, new_n306_ );
and g1270 ( new_n1472_, new_n1471_, new_n542_ );
and g1271 ( new_n1473_, new_n1472_, new_n534_ );
and g1272 ( new_n1474_, new_n1267_, new_n1473_ );
and g1273 ( new_n1475_, new_n1474_, new_n1470_ );
not g1274 ( new_n1476_, new_n1473_ );
or g1275 ( new_n1477_, new_n1279_, new_n1476_ );
and g1276 ( new_n1478_, new_n1477_, keyIn_0_80 );
or g1277 ( new_n1479_, new_n1478_, new_n1079_ );
or g1278 ( new_n1480_, new_n1479_, new_n1475_ );
and g1279 ( new_n1481_, new_n1480_, new_n1469_ );
not g1280 ( new_n1482_, new_n1475_ );
or g1281 ( new_n1483_, new_n1474_, new_n1470_ );
and g1282 ( new_n1484_, new_n1483_, new_n682_ );
and g1283 ( new_n1485_, new_n1484_, new_n1482_ );
and g1284 ( new_n1486_, new_n1485_, keyIn_0_97 );
or g1285 ( new_n1487_, new_n1481_, new_n1486_ );
and g1286 ( new_n1488_, new_n1487_, N97 );
or g1287 ( new_n1489_, new_n1485_, keyIn_0_97 );
or g1288 ( new_n1490_, new_n1480_, new_n1469_ );
and g1289 ( new_n1491_, new_n1490_, new_n1489_ );
and g1290 ( new_n1492_, new_n1491_, new_n311_ );
or g1291 ( new_n1493_, new_n1488_, new_n1492_ );
and g1292 ( new_n1494_, new_n1493_, keyIn_0_120 );
not g1293 ( new_n1495_, keyIn_0_120 );
or g1294 ( new_n1496_, new_n1491_, new_n311_ );
or g1295 ( new_n1497_, new_n1487_, N97 );
and g1296 ( new_n1498_, new_n1496_, new_n1497_ );
and g1297 ( new_n1499_, new_n1498_, new_n1495_ );
or g1298 ( N748, new_n1494_, new_n1499_ );
not g1299 ( new_n1501_, keyIn_0_98 );
and g1300 ( new_n1502_, new_n1483_, new_n1076_ );
and g1301 ( new_n1503_, new_n1502_, new_n1482_ );
or g1302 ( new_n1504_, new_n1503_, new_n1501_ );
or g1303 ( new_n1505_, new_n1478_, new_n899_ );
or g1304 ( new_n1506_, new_n1505_, new_n1475_ );
or g1305 ( new_n1507_, new_n1506_, keyIn_0_98 );
and g1306 ( new_n1508_, new_n1507_, new_n1504_ );
or g1307 ( new_n1509_, new_n1508_, N101 );
and g1308 ( new_n1510_, new_n1506_, keyIn_0_98 );
and g1309 ( new_n1511_, new_n1503_, new_n1501_ );
or g1310 ( new_n1512_, new_n1510_, new_n1511_ );
or g1311 ( new_n1513_, new_n1512_, new_n309_ );
and g1312 ( new_n1514_, new_n1509_, new_n1513_ );
or g1313 ( new_n1515_, new_n1514_, keyIn_0_121 );
not g1314 ( new_n1516_, keyIn_0_121 );
and g1315 ( new_n1517_, new_n1512_, new_n309_ );
and g1316 ( new_n1518_, new_n1508_, N101 );
or g1317 ( new_n1519_, new_n1517_, new_n1518_ );
or g1318 ( new_n1520_, new_n1519_, new_n1516_ );
and g1319 ( N749, new_n1520_, new_n1515_ );
not g1320 ( new_n1522_, keyIn_0_122 );
and g1321 ( new_n1523_, new_n1483_, new_n791_ );
and g1322 ( new_n1524_, new_n1523_, new_n1482_ );
or g1323 ( new_n1525_, new_n1524_, keyIn_0_99 );
not g1324 ( new_n1526_, keyIn_0_99 );
or g1325 ( new_n1527_, new_n1478_, new_n985_ );
or g1326 ( new_n1528_, new_n1527_, new_n1475_ );
or g1327 ( new_n1529_, new_n1528_, new_n1526_ );
and g1328 ( new_n1530_, new_n1529_, new_n1525_ );
or g1329 ( new_n1531_, new_n1530_, new_n322_ );
and g1330 ( new_n1532_, new_n1528_, new_n1526_ );
and g1331 ( new_n1533_, new_n1524_, keyIn_0_99 );
or g1332 ( new_n1534_, new_n1532_, new_n1533_ );
or g1333 ( new_n1535_, new_n1534_, N105 );
and g1334 ( new_n1536_, new_n1531_, new_n1535_ );
or g1335 ( new_n1537_, new_n1536_, new_n1522_ );
and g1336 ( new_n1538_, new_n1534_, N105 );
and g1337 ( new_n1539_, new_n1530_, new_n322_ );
or g1338 ( new_n1540_, new_n1538_, new_n1539_ );
or g1339 ( new_n1541_, new_n1540_, keyIn_0_122 );
and g1340 ( N750, new_n1541_, new_n1537_ );
and g1341 ( new_n1543_, new_n1483_, new_n988_ );
and g1342 ( new_n1544_, new_n1543_, new_n1482_ );
or g1343 ( new_n1545_, new_n1544_, keyIn_0_100 );
not g1344 ( new_n1546_, keyIn_0_100 );
or g1345 ( new_n1547_, new_n1478_, new_n955_ );
or g1346 ( new_n1548_, new_n1547_, new_n1475_ );
or g1347 ( new_n1549_, new_n1548_, new_n1546_ );
and g1348 ( new_n1550_, new_n1549_, new_n1545_ );
or g1349 ( new_n1551_, new_n1550_, new_n320_ );
and g1350 ( new_n1552_, new_n1548_, new_n1546_ );
and g1351 ( new_n1553_, new_n1544_, keyIn_0_100 );
or g1352 ( new_n1554_, new_n1552_, new_n1553_ );
or g1353 ( new_n1555_, new_n1554_, N109 );
and g1354 ( new_n1556_, new_n1551_, new_n1555_ );
or g1355 ( new_n1557_, new_n1556_, keyIn_0_123 );
not g1356 ( new_n1558_, keyIn_0_123 );
and g1357 ( new_n1559_, new_n1554_, N109 );
and g1358 ( new_n1560_, new_n1550_, new_n320_ );
or g1359 ( new_n1561_, new_n1559_, new_n1560_ );
or g1360 ( new_n1562_, new_n1561_, new_n1558_ );
and g1361 ( N751, new_n1562_, new_n1557_ );
not g1362 ( new_n1564_, keyIn_0_124 );
not g1363 ( new_n1565_, keyIn_0_81 );
not g1364 ( new_n1566_, keyIn_0_70 );
and g1365 ( new_n1567_, new_n403_, new_n1566_ );
and g1366 ( new_n1568_, new_n534_, keyIn_0_70 );
or g1367 ( new_n1569_, new_n1568_, new_n1567_ );
not g1368 ( new_n1570_, new_n1569_ );
not g1369 ( new_n1571_, keyIn_0_69 );
and g1370 ( new_n1572_, new_n306_, new_n1571_ );
and g1371 ( new_n1573_, new_n307_, keyIn_0_69 );
or g1372 ( new_n1574_, new_n1573_, new_n528_ );
or g1373 ( new_n1575_, new_n1574_, new_n1572_ );
or g1374 ( new_n1576_, new_n1570_, new_n1575_ );
not g1375 ( new_n1577_, new_n1576_ );
and g1376 ( new_n1578_, new_n1267_, new_n1577_ );
and g1377 ( new_n1579_, new_n1578_, new_n1565_ );
not g1378 ( new_n1580_, new_n1579_ );
or g1379 ( new_n1581_, new_n1578_, new_n1565_ );
and g1380 ( new_n1582_, new_n1581_, new_n682_ );
and g1381 ( new_n1583_, new_n1582_, new_n1580_ );
or g1382 ( new_n1584_, new_n1583_, keyIn_0_101 );
not g1383 ( new_n1585_, keyIn_0_101 );
or g1384 ( new_n1586_, new_n1279_, new_n1576_ );
and g1385 ( new_n1587_, new_n1586_, keyIn_0_81 );
or g1386 ( new_n1588_, new_n1587_, new_n1079_ );
or g1387 ( new_n1589_, new_n1588_, new_n1579_ );
or g1388 ( new_n1590_, new_n1589_, new_n1585_ );
and g1389 ( new_n1591_, new_n1590_, new_n1584_ );
or g1390 ( new_n1592_, new_n1591_, N113 );
and g1391 ( new_n1593_, new_n1589_, new_n1585_ );
and g1392 ( new_n1594_, new_n1583_, keyIn_0_101 );
or g1393 ( new_n1595_, new_n1593_, new_n1594_ );
or g1394 ( new_n1596_, new_n1595_, new_n410_ );
and g1395 ( new_n1597_, new_n1592_, new_n1596_ );
or g1396 ( new_n1598_, new_n1597_, new_n1564_ );
and g1397 ( new_n1599_, new_n1595_, new_n410_ );
and g1398 ( new_n1600_, new_n1591_, N113 );
or g1399 ( new_n1601_, new_n1599_, new_n1600_ );
or g1400 ( new_n1602_, new_n1601_, keyIn_0_124 );
and g1401 ( N752, new_n1602_, new_n1598_ );
or g1402 ( new_n1604_, new_n1587_, new_n899_ );
or g1403 ( new_n1605_, new_n1604_, new_n1579_ );
and g1404 ( new_n1606_, new_n1605_, keyIn_0_102 );
not g1405 ( new_n1607_, keyIn_0_102 );
and g1406 ( new_n1608_, new_n1581_, new_n1076_ );
and g1407 ( new_n1609_, new_n1608_, new_n1580_ );
and g1408 ( new_n1610_, new_n1609_, new_n1607_ );
or g1409 ( new_n1611_, new_n1606_, new_n1610_ );
and g1410 ( new_n1612_, new_n1611_, N117 );
or g1411 ( new_n1613_, new_n1609_, new_n1607_ );
or g1412 ( new_n1614_, new_n1605_, keyIn_0_102 );
and g1413 ( new_n1615_, new_n1614_, new_n1613_ );
and g1414 ( new_n1616_, new_n1615_, new_n408_ );
or g1415 ( new_n1617_, new_n1612_, new_n1616_ );
and g1416 ( new_n1618_, new_n1617_, keyIn_0_125 );
not g1417 ( new_n1619_, keyIn_0_125 );
or g1418 ( new_n1620_, new_n1615_, new_n408_ );
or g1419 ( new_n1621_, new_n1611_, N117 );
and g1420 ( new_n1622_, new_n1620_, new_n1621_ );
and g1421 ( new_n1623_, new_n1622_, new_n1619_ );
or g1422 ( N753, new_n1618_, new_n1623_ );
not g1423 ( new_n1625_, keyIn_0_126 );
or g1424 ( new_n1626_, new_n1587_, new_n985_ );
or g1425 ( new_n1627_, new_n1626_, new_n1579_ );
and g1426 ( new_n1628_, new_n1627_, keyIn_0_103 );
not g1427 ( new_n1629_, keyIn_0_103 );
and g1428 ( new_n1630_, new_n1581_, new_n791_ );
and g1429 ( new_n1631_, new_n1630_, new_n1580_ );
and g1430 ( new_n1632_, new_n1631_, new_n1629_ );
or g1431 ( new_n1633_, new_n1628_, new_n1632_ );
and g1432 ( new_n1634_, new_n1633_, new_n421_ );
or g1433 ( new_n1635_, new_n1631_, new_n1629_ );
or g1434 ( new_n1636_, new_n1627_, keyIn_0_103 );
and g1435 ( new_n1637_, new_n1636_, new_n1635_ );
and g1436 ( new_n1638_, new_n1637_, N121 );
or g1437 ( new_n1639_, new_n1634_, new_n1638_ );
and g1438 ( new_n1640_, new_n1639_, new_n1625_ );
or g1439 ( new_n1641_, new_n1637_, N121 );
or g1440 ( new_n1642_, new_n1633_, new_n421_ );
and g1441 ( new_n1643_, new_n1641_, new_n1642_ );
and g1442 ( new_n1644_, new_n1643_, keyIn_0_126 );
or g1443 ( N754, new_n1640_, new_n1644_ );
not g1444 ( new_n1646_, keyIn_0_104 );
and g1445 ( new_n1647_, new_n1581_, new_n988_ );
and g1446 ( new_n1648_, new_n1647_, new_n1580_ );
or g1447 ( new_n1649_, new_n1648_, new_n1646_ );
or g1448 ( new_n1650_, new_n1587_, new_n955_ );
or g1449 ( new_n1651_, new_n1650_, new_n1579_ );
or g1450 ( new_n1652_, new_n1651_, keyIn_0_104 );
and g1451 ( new_n1653_, new_n1652_, new_n1649_ );
or g1452 ( new_n1654_, new_n1653_, new_n419_ );
and g1453 ( new_n1655_, new_n1651_, keyIn_0_104 );
and g1454 ( new_n1656_, new_n1648_, new_n1646_ );
or g1455 ( new_n1657_, new_n1655_, new_n1656_ );
or g1456 ( new_n1658_, new_n1657_, N125 );
and g1457 ( new_n1659_, new_n1654_, new_n1658_ );
or g1458 ( new_n1660_, new_n1659_, keyIn_0_127 );
not g1459 ( new_n1661_, keyIn_0_127 );
and g1460 ( new_n1662_, new_n1657_, N125 );
and g1461 ( new_n1663_, new_n1653_, new_n419_ );
or g1462 ( new_n1664_, new_n1662_, new_n1663_ );
or g1463 ( new_n1665_, new_n1664_, new_n1661_ );
and g1464 ( N755, new_n1665_, new_n1660_ );
endmodule