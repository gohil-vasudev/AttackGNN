module locked_c3540 (  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n143_, new_n144_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1251_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1278_, new_n1279_, new_n1280_;
  NOR2_X1 g0000 ( .A1(G58), .A2(G68), .ZN(new_n137_) );
  INV_X1 g0001 ( .A(new_n137_), .ZN(new_n138_) );
  INV_X1 g0002 ( .A(G50), .ZN(new_n139_) );
  INV_X1 g0003 ( .A(G77), .ZN(new_n140_) );
  NAND2_X1 g0004 ( .A1(new_n139_), .A2(new_n140_), .ZN(new_n141_) );
  NOR2_X1 g0005 ( .A1(new_n138_), .A2(new_n141_), .ZN(G353) );
  NOR2_X1 g0006 ( .A1(G97), .A2(G107), .ZN(new_n143_) );
  INV_X1 g0007 ( .A(new_n143_), .ZN(new_n144_) );
  NAND2_X1 g0008 ( .A1(new_n144_), .A2(G87), .ZN(G355) );
  NAND2_X1 g0009 ( .A1(G1), .A2(G20), .ZN(new_n146_) );
  INV_X1 g0010 ( .A(KEYINPUT49), .ZN(new_n147_) );
  NAND2_X1 g0011 ( .A1(G58), .A2(G232), .ZN(new_n148_) );
  NAND2_X1 g0012 ( .A1(G50), .A2(G226), .ZN(new_n149_) );
  NAND2_X1 g0013 ( .A1(G68), .A2(G238), .ZN(new_n150_) );
  NAND2_X1 g0014 ( .A1(G77), .A2(G244), .ZN(new_n151_) );
  NAND4_X1 g0015 ( .A1(new_n148_), .A2(new_n149_), .A3(new_n150_), .A4(new_n151_), .ZN(new_n152_) );
  NAND2_X1 g0016 ( .A1(new_n152_), .A2(new_n147_), .ZN(new_n153_) );
  NOR2_X1 g0017 ( .A1(new_n152_), .A2(new_n147_), .ZN(new_n154_) );
  NAND2_X1 g0018 ( .A1(G116), .A2(G270), .ZN(new_n155_) );
  NAND2_X1 g0019 ( .A1(G97), .A2(G257), .ZN(new_n156_) );
  NAND2_X1 g0020 ( .A1(G87), .A2(G250), .ZN(new_n157_) );
  NAND3_X1 g0021 ( .A1(new_n155_), .A2(new_n156_), .A3(new_n157_), .ZN(new_n158_) );
  INV_X1 g0022 ( .A(KEYINPUT50), .ZN(new_n159_) );
  NAND2_X1 g0023 ( .A1(G107), .A2(G264), .ZN(new_n160_) );
  NAND2_X1 g0024 ( .A1(new_n160_), .A2(new_n159_), .ZN(new_n161_) );
  NAND3_X1 g0025 ( .A1(G107), .A2(G264), .A3(KEYINPUT50), .ZN(new_n162_) );
  NAND2_X1 g0026 ( .A1(new_n161_), .A2(new_n162_), .ZN(new_n163_) );
  NOR3_X1 g0027 ( .A1(new_n154_), .A2(new_n158_), .A3(new_n163_), .ZN(new_n164_) );
  NAND2_X1 g0028 ( .A1(new_n164_), .A2(new_n153_), .ZN(new_n165_) );
  NAND2_X1 g0029 ( .A1(new_n165_), .A2(new_n146_), .ZN(new_n166_) );
  NOR2_X1 g0030 ( .A1(new_n146_), .A2(G13), .ZN(new_n167_) );
  INV_X1 g0031 ( .A(G257), .ZN(new_n168_) );
  INV_X1 g0032 ( .A(G264), .ZN(new_n169_) );
  NAND2_X1 g0033 ( .A1(new_n168_), .A2(new_n169_), .ZN(new_n170_) );
  NAND3_X1 g0034 ( .A1(new_n167_), .A2(G250), .A3(new_n170_), .ZN(new_n171_) );
  NAND2_X1 g0035 ( .A1(G1), .A2(G13), .ZN(new_n172_) );
  NAND2_X1 g0036 ( .A1(new_n172_), .A2(KEYINPUT2), .ZN(new_n173_) );
  INV_X1 g0037 ( .A(KEYINPUT2), .ZN(new_n174_) );
  NAND3_X1 g0038 ( .A1(new_n174_), .A2(G1), .A3(G13), .ZN(new_n175_) );
  NAND2_X1 g0039 ( .A1(new_n173_), .A2(new_n175_), .ZN(new_n176_) );
  INV_X1 g0040 ( .A(new_n176_), .ZN(new_n177_) );
  NAND2_X1 g0041 ( .A1(new_n177_), .A2(G20), .ZN(new_n178_) );
  INV_X1 g0042 ( .A(new_n178_), .ZN(new_n179_) );
  NOR2_X1 g0043 ( .A1(new_n137_), .A2(new_n139_), .ZN(new_n180_) );
  NAND2_X1 g0044 ( .A1(new_n179_), .A2(new_n180_), .ZN(new_n181_) );
  NAND3_X1 g0045 ( .A1(new_n166_), .A2(new_n171_), .A3(new_n181_), .ZN(new_n182_) );
  INV_X1 g0046 ( .A(new_n182_), .ZN(G361) );
  INV_X1 g0047 ( .A(G238), .ZN(new_n184_) );
  NOR2_X1 g0048 ( .A1(G232), .A2(G244), .ZN(new_n185_) );
  INV_X1 g0049 ( .A(new_n185_), .ZN(new_n186_) );
  NAND2_X1 g0050 ( .A1(G232), .A2(G244), .ZN(new_n187_) );
  NAND2_X1 g0051 ( .A1(new_n186_), .A2(new_n187_), .ZN(new_n188_) );
  NAND2_X1 g0052 ( .A1(new_n188_), .A2(G226), .ZN(new_n189_) );
  INV_X1 g0053 ( .A(new_n189_), .ZN(new_n190_) );
  NOR2_X1 g0054 ( .A1(new_n188_), .A2(G226), .ZN(new_n191_) );
  NOR2_X1 g0055 ( .A1(new_n190_), .A2(new_n191_), .ZN(new_n192_) );
  INV_X1 g0056 ( .A(new_n192_), .ZN(new_n193_) );
  NAND2_X1 g0057 ( .A1(new_n193_), .A2(new_n184_), .ZN(new_n194_) );
  NAND2_X1 g0058 ( .A1(new_n192_), .A2(G238), .ZN(new_n195_) );
  INV_X1 g0059 ( .A(G270), .ZN(new_n196_) );
  NAND2_X1 g0060 ( .A1(new_n169_), .A2(new_n196_), .ZN(new_n197_) );
  NAND2_X1 g0061 ( .A1(G264), .A2(G270), .ZN(new_n198_) );
  NAND2_X1 g0062 ( .A1(new_n197_), .A2(new_n198_), .ZN(new_n199_) );
  INV_X1 g0063 ( .A(G250), .ZN(new_n200_) );
  NAND2_X1 g0064 ( .A1(new_n200_), .A2(new_n168_), .ZN(new_n201_) );
  NAND2_X1 g0065 ( .A1(G250), .A2(G257), .ZN(new_n202_) );
  NAND2_X1 g0066 ( .A1(new_n201_), .A2(new_n202_), .ZN(new_n203_) );
  NAND2_X1 g0067 ( .A1(new_n199_), .A2(new_n203_), .ZN(new_n204_) );
  NAND4_X1 g0068 ( .A1(new_n197_), .A2(new_n201_), .A3(new_n198_), .A4(new_n202_), .ZN(new_n205_) );
  NAND2_X1 g0069 ( .A1(new_n204_), .A2(new_n205_), .ZN(new_n206_) );
  NAND3_X1 g0070 ( .A1(new_n194_), .A2(new_n195_), .A3(new_n206_), .ZN(new_n207_) );
  NAND2_X1 g0071 ( .A1(new_n194_), .A2(new_n195_), .ZN(new_n208_) );
  NAND3_X1 g0072 ( .A1(new_n208_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n209_) );
  NAND2_X1 g0073 ( .A1(new_n209_), .A2(new_n207_), .ZN(G358) );
  INV_X1 g0074 ( .A(KEYINPUT51), .ZN(new_n211_) );
  NAND2_X1 g0075 ( .A1(G97), .A2(G107), .ZN(new_n212_) );
  NAND2_X1 g0076 ( .A1(new_n144_), .A2(new_n212_), .ZN(new_n213_) );
  INV_X1 g0077 ( .A(new_n213_), .ZN(new_n214_) );
  NAND2_X1 g0078 ( .A1(new_n214_), .A2(new_n211_), .ZN(new_n215_) );
  NAND2_X1 g0079 ( .A1(new_n213_), .A2(KEYINPUT51), .ZN(new_n216_) );
  NAND2_X1 g0080 ( .A1(new_n215_), .A2(new_n216_), .ZN(new_n217_) );
  INV_X1 g0081 ( .A(G87), .ZN(new_n218_) );
  NOR2_X1 g0082 ( .A1(new_n218_), .A2(G116), .ZN(new_n219_) );
  INV_X1 g0083 ( .A(G116), .ZN(new_n220_) );
  NOR2_X1 g0084 ( .A1(new_n220_), .A2(G87), .ZN(new_n221_) );
  NOR2_X1 g0085 ( .A1(new_n219_), .A2(new_n221_), .ZN(new_n222_) );
  INV_X1 g0086 ( .A(new_n222_), .ZN(new_n223_) );
  NAND2_X1 g0087 ( .A1(new_n217_), .A2(new_n223_), .ZN(new_n224_) );
  NAND3_X1 g0088 ( .A1(new_n215_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n225_) );
  NAND2_X1 g0089 ( .A1(new_n224_), .A2(new_n225_), .ZN(new_n226_) );
  NAND2_X1 g0090 ( .A1(G58), .A2(G68), .ZN(new_n227_) );
  NAND2_X1 g0091 ( .A1(new_n138_), .A2(new_n227_), .ZN(new_n228_) );
  NAND2_X1 g0092 ( .A1(G50), .A2(G77), .ZN(new_n229_) );
  NAND2_X1 g0093 ( .A1(new_n141_), .A2(new_n229_), .ZN(new_n230_) );
  NAND2_X1 g0094 ( .A1(new_n228_), .A2(new_n230_), .ZN(new_n231_) );
  NAND4_X1 g0095 ( .A1(new_n138_), .A2(new_n141_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n232_) );
  NAND2_X1 g0096 ( .A1(new_n231_), .A2(new_n232_), .ZN(new_n233_) );
  NAND2_X1 g0097 ( .A1(new_n226_), .A2(new_n233_), .ZN(new_n234_) );
  NAND4_X1 g0098 ( .A1(new_n224_), .A2(new_n225_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n235_) );
  NAND2_X1 g0099 ( .A1(new_n234_), .A2(new_n235_), .ZN(G351) );
  INV_X1 g0100 ( .A(KEYINPUT30), .ZN(new_n237_) );
  INV_X1 g0101 ( .A(KEYINPUT3), .ZN(new_n238_) );
  NAND3_X1 g0102 ( .A1(G1), .A2(G20), .A3(G33), .ZN(new_n239_) );
  NAND2_X1 g0103 ( .A1(new_n239_), .A2(new_n238_), .ZN(new_n240_) );
  NAND4_X1 g0104 ( .A1(G1), .A2(G20), .A3(G33), .A4(KEYINPUT3), .ZN(new_n241_) );
  NAND2_X1 g0105 ( .A1(new_n240_), .A2(new_n241_), .ZN(new_n242_) );
  NAND2_X1 g0106 ( .A1(new_n242_), .A2(new_n176_), .ZN(new_n243_) );
  NAND2_X1 g0107 ( .A1(new_n243_), .A2(G20), .ZN(new_n244_) );
  NAND2_X1 g0108 ( .A1(new_n244_), .A2(KEYINPUT4), .ZN(new_n245_) );
  INV_X1 g0109 ( .A(KEYINPUT4), .ZN(new_n246_) );
  NAND3_X1 g0110 ( .A1(new_n243_), .A2(G20), .A3(new_n246_), .ZN(new_n247_) );
  NAND2_X1 g0111 ( .A1(new_n245_), .A2(new_n247_), .ZN(new_n248_) );
  INV_X1 g0112 ( .A(new_n248_), .ZN(new_n249_) );
  NAND2_X1 g0113 ( .A1(new_n249_), .A2(new_n228_), .ZN(new_n250_) );
  INV_X1 g0114 ( .A(new_n243_), .ZN(new_n251_) );
  INV_X1 g0115 ( .A(G1), .ZN(new_n252_) );
  NAND2_X1 g0116 ( .A1(new_n252_), .A2(G20), .ZN(new_n253_) );
  NAND3_X1 g0117 ( .A1(new_n251_), .A2(G58), .A3(new_n253_), .ZN(new_n254_) );
  INV_X1 g0118 ( .A(new_n254_), .ZN(new_n255_) );
  INV_X1 g0119 ( .A(G159), .ZN(new_n256_) );
  INV_X1 g0120 ( .A(G20), .ZN(new_n257_) );
  INV_X1 g0121 ( .A(G33), .ZN(new_n258_) );
  NAND3_X1 g0122 ( .A1(new_n177_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_) );
  NOR2_X1 g0123 ( .A1(new_n259_), .A2(new_n256_), .ZN(new_n260_) );
  INV_X1 g0124 ( .A(G58), .ZN(new_n261_) );
  NAND3_X1 g0125 ( .A1(new_n252_), .A2(G13), .A3(G20), .ZN(new_n262_) );
  INV_X1 g0126 ( .A(new_n262_), .ZN(new_n263_) );
  NAND2_X1 g0127 ( .A1(new_n263_), .A2(new_n261_), .ZN(new_n264_) );
  NOR2_X1 g0128 ( .A1(new_n258_), .A2(G20), .ZN(new_n265_) );
  NAND2_X1 g0129 ( .A1(new_n177_), .A2(new_n265_), .ZN(new_n266_) );
  INV_X1 g0130 ( .A(new_n266_), .ZN(new_n267_) );
  NAND2_X1 g0131 ( .A1(new_n267_), .A2(G68), .ZN(new_n268_) );
  NAND2_X1 g0132 ( .A1(new_n268_), .A2(new_n264_), .ZN(new_n269_) );
  NOR3_X1 g0133 ( .A1(new_n269_), .A2(new_n255_), .A3(new_n260_), .ZN(new_n270_) );
  NAND3_X1 g0134 ( .A1(new_n270_), .A2(new_n250_), .A3(new_n237_), .ZN(new_n271_) );
  NAND2_X1 g0135 ( .A1(new_n270_), .A2(new_n250_), .ZN(new_n272_) );
  NAND2_X1 g0136 ( .A1(new_n272_), .A2(KEYINPUT30), .ZN(new_n273_) );
  NAND2_X1 g0137 ( .A1(new_n273_), .A2(new_n271_), .ZN(new_n274_) );
  NAND4_X1 g0138 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n258_), .A4(G1698), .ZN(new_n275_) );
  INV_X1 g0139 ( .A(new_n275_), .ZN(new_n276_) );
  NAND2_X1 g0140 ( .A1(new_n276_), .A2(G226), .ZN(new_n277_) );
  NAND2_X1 g0141 ( .A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n278_) );
  INV_X1 g0142 ( .A(KEYINPUT32), .ZN(new_n279_) );
  NAND3_X1 g0143 ( .A1(new_n276_), .A2(G226), .A3(new_n279_), .ZN(new_n280_) );
  NAND2_X1 g0144 ( .A1(new_n278_), .A2(new_n280_), .ZN(new_n281_) );
  INV_X1 g0145 ( .A(G1698), .ZN(new_n282_) );
  NAND4_X1 g0146 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n258_), .A4(new_n282_), .ZN(new_n283_) );
  INV_X1 g0147 ( .A(new_n283_), .ZN(new_n284_) );
  NAND2_X1 g0148 ( .A1(new_n284_), .A2(G223), .ZN(new_n285_) );
  NAND2_X1 g0149 ( .A1(new_n281_), .A2(new_n285_), .ZN(new_n286_) );
  NAND2_X1 g0150 ( .A1(new_n286_), .A2(KEYINPUT33), .ZN(new_n287_) );
  INV_X1 g0151 ( .A(KEYINPUT33), .ZN(new_n288_) );
  NAND3_X1 g0152 ( .A1(new_n281_), .A2(new_n288_), .A3(new_n285_), .ZN(new_n289_) );
  NAND2_X1 g0153 ( .A1(new_n287_), .A2(new_n289_), .ZN(new_n290_) );
  INV_X1 g0154 ( .A(G41), .ZN(new_n291_) );
  INV_X1 g0155 ( .A(G45), .ZN(new_n292_) );
  NAND2_X1 g0156 ( .A1(new_n291_), .A2(new_n292_), .ZN(new_n293_) );
  NAND3_X1 g0157 ( .A1(new_n293_), .A2(new_n252_), .A3(G274), .ZN(new_n294_) );
  INV_X1 g0158 ( .A(new_n294_), .ZN(new_n295_) );
  NOR2_X1 g0159 ( .A1(new_n258_), .A2(G41), .ZN(new_n296_) );
  NAND3_X1 g0160 ( .A1(new_n177_), .A2(G87), .A3(new_n296_), .ZN(new_n297_) );
  NOR2_X1 g0161 ( .A1(new_n297_), .A2(KEYINPUT31), .ZN(new_n298_) );
  NAND2_X1 g0162 ( .A1(new_n297_), .A2(KEYINPUT31), .ZN(new_n299_) );
  NAND2_X1 g0163 ( .A1(new_n293_), .A2(new_n252_), .ZN(new_n300_) );
  NAND2_X1 g0164 ( .A1(G33), .A2(G41), .ZN(new_n301_) );
  NAND3_X1 g0165 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n301_), .ZN(new_n302_) );
  NAND2_X1 g0166 ( .A1(new_n302_), .A2(new_n300_), .ZN(new_n303_) );
  INV_X1 g0167 ( .A(new_n303_), .ZN(new_n304_) );
  NAND2_X1 g0168 ( .A1(new_n304_), .A2(G232), .ZN(new_n305_) );
  NAND2_X1 g0169 ( .A1(new_n305_), .A2(new_n299_), .ZN(new_n306_) );
  NOR3_X1 g0170 ( .A1(new_n306_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n307_) );
  NAND3_X1 g0171 ( .A1(new_n290_), .A2(G179), .A3(new_n307_), .ZN(new_n308_) );
  NAND2_X1 g0172 ( .A1(new_n308_), .A2(KEYINPUT34), .ZN(new_n309_) );
  INV_X1 g0173 ( .A(KEYINPUT34), .ZN(new_n310_) );
  NAND4_X1 g0174 ( .A1(new_n290_), .A2(G179), .A3(new_n310_), .A4(new_n307_), .ZN(new_n311_) );
  NAND2_X1 g0175 ( .A1(new_n309_), .A2(new_n311_), .ZN(new_n312_) );
  NAND2_X1 g0176 ( .A1(new_n290_), .A2(new_n307_), .ZN(new_n313_) );
  NAND2_X1 g0177 ( .A1(new_n313_), .A2(G169), .ZN(new_n314_) );
  NAND2_X1 g0178 ( .A1(new_n312_), .A2(new_n314_), .ZN(new_n315_) );
  NAND2_X1 g0179 ( .A1(new_n315_), .A2(new_n274_), .ZN(new_n316_) );
  INV_X1 g0180 ( .A(new_n316_), .ZN(new_n317_) );
  INV_X1 g0181 ( .A(KEYINPUT35), .ZN(new_n318_) );
  NAND2_X1 g0182 ( .A1(new_n313_), .A2(G200), .ZN(new_n319_) );
  NAND2_X1 g0183 ( .A1(new_n319_), .A2(new_n318_), .ZN(new_n320_) );
  NAND3_X1 g0184 ( .A1(new_n313_), .A2(G200), .A3(KEYINPUT35), .ZN(new_n321_) );
  NAND2_X1 g0185 ( .A1(new_n320_), .A2(new_n321_), .ZN(new_n322_) );
  NAND3_X1 g0186 ( .A1(new_n290_), .A2(G190), .A3(new_n307_), .ZN(new_n323_) );
  NAND4_X1 g0187 ( .A1(new_n322_), .A2(new_n271_), .A3(new_n273_), .A4(new_n323_), .ZN(new_n324_) );
  INV_X1 g0188 ( .A(KEYINPUT6), .ZN(new_n325_) );
  NAND2_X1 g0189 ( .A1(new_n276_), .A2(G238), .ZN(new_n326_) );
  NAND2_X1 g0190 ( .A1(new_n326_), .A2(new_n325_), .ZN(new_n327_) );
  NOR3_X1 g0191 ( .A1(new_n275_), .A2(new_n184_), .A3(new_n325_), .ZN(new_n328_) );
  INV_X1 g0192 ( .A(G232), .ZN(new_n329_) );
  NOR2_X1 g0193 ( .A1(new_n283_), .A2(new_n329_), .ZN(new_n330_) );
  NAND4_X1 g0194 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n296_), .A4(G107), .ZN(new_n331_) );
  NAND2_X1 g0195 ( .A1(new_n331_), .A2(new_n294_), .ZN(new_n332_) );
  NOR3_X1 g0196 ( .A1(new_n328_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_) );
  NAND2_X1 g0197 ( .A1(new_n333_), .A2(new_n327_), .ZN(new_n334_) );
  NAND2_X1 g0198 ( .A1(new_n334_), .A2(KEYINPUT7), .ZN(new_n335_) );
  INV_X1 g0199 ( .A(KEYINPUT7), .ZN(new_n336_) );
  NAND3_X1 g0200 ( .A1(new_n333_), .A2(new_n336_), .A3(new_n327_), .ZN(new_n337_) );
  NAND2_X1 g0201 ( .A1(new_n335_), .A2(new_n337_), .ZN(new_n338_) );
  NAND2_X1 g0202 ( .A1(new_n304_), .A2(G244), .ZN(new_n339_) );
  NAND2_X1 g0203 ( .A1(new_n338_), .A2(new_n339_), .ZN(new_n340_) );
  NAND2_X1 g0204 ( .A1(new_n340_), .A2(G169), .ZN(new_n341_) );
  NAND3_X1 g0205 ( .A1(new_n338_), .A2(G179), .A3(new_n339_), .ZN(new_n342_) );
  NAND2_X1 g0206 ( .A1(new_n341_), .A2(new_n342_), .ZN(new_n343_) );
  NAND2_X1 g0207 ( .A1(new_n251_), .A2(new_n253_), .ZN(new_n344_) );
  NAND2_X1 g0208 ( .A1(new_n248_), .A2(new_n344_), .ZN(new_n345_) );
  NAND2_X1 g0209 ( .A1(new_n345_), .A2(G77), .ZN(new_n346_) );
  NOR2_X1 g0210 ( .A1(new_n259_), .A2(new_n261_), .ZN(new_n347_) );
  NAND2_X1 g0211 ( .A1(new_n267_), .A2(G87), .ZN(new_n348_) );
  NAND2_X1 g0212 ( .A1(new_n263_), .A2(new_n140_), .ZN(new_n349_) );
  NAND2_X1 g0213 ( .A1(new_n348_), .A2(new_n349_), .ZN(new_n350_) );
  NOR2_X1 g0214 ( .A1(new_n350_), .A2(new_n347_), .ZN(new_n351_) );
  NAND2_X1 g0215 ( .A1(new_n346_), .A2(new_n351_), .ZN(new_n352_) );
  NAND2_X1 g0216 ( .A1(new_n343_), .A2(new_n352_), .ZN(new_n353_) );
  NAND2_X1 g0217 ( .A1(new_n340_), .A2(G200), .ZN(new_n354_) );
  NAND3_X1 g0218 ( .A1(new_n338_), .A2(G190), .A3(new_n339_), .ZN(new_n355_) );
  NAND4_X1 g0219 ( .A1(new_n354_), .A2(new_n346_), .A3(new_n351_), .A4(new_n355_), .ZN(new_n356_) );
  NAND2_X1 g0220 ( .A1(new_n353_), .A2(new_n356_), .ZN(new_n357_) );
  INV_X1 g0221 ( .A(new_n357_), .ZN(new_n358_) );
  INV_X1 g0222 ( .A(G68), .ZN(new_n359_) );
  NAND2_X1 g0223 ( .A1(new_n248_), .A2(new_n262_), .ZN(new_n360_) );
  NAND2_X1 g0224 ( .A1(new_n360_), .A2(new_n359_), .ZN(new_n361_) );
  NAND3_X1 g0225 ( .A1(new_n251_), .A2(G68), .A3(new_n253_), .ZN(new_n362_) );
  INV_X1 g0226 ( .A(new_n362_), .ZN(new_n363_) );
  NAND2_X1 g0227 ( .A1(new_n267_), .A2(G77), .ZN(new_n364_) );
  INV_X1 g0228 ( .A(new_n364_), .ZN(new_n365_) );
  NOR2_X1 g0229 ( .A1(new_n259_), .A2(new_n139_), .ZN(new_n366_) );
  NOR3_X1 g0230 ( .A1(new_n365_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_) );
  NAND2_X1 g0231 ( .A1(new_n361_), .A2(new_n367_), .ZN(new_n368_) );
  INV_X1 g0232 ( .A(G179), .ZN(new_n369_) );
  NOR2_X1 g0233 ( .A1(new_n275_), .A2(new_n329_), .ZN(new_n370_) );
  NAND3_X1 g0234 ( .A1(new_n177_), .A2(G97), .A3(new_n296_), .ZN(new_n371_) );
  NAND2_X1 g0235 ( .A1(new_n371_), .A2(new_n294_), .ZN(new_n372_) );
  NAND2_X1 g0236 ( .A1(new_n284_), .A2(G226), .ZN(new_n373_) );
  NAND2_X1 g0237 ( .A1(new_n304_), .A2(G238), .ZN(new_n374_) );
  NAND2_X1 g0238 ( .A1(new_n374_), .A2(new_n373_), .ZN(new_n375_) );
  NOR3_X1 g0239 ( .A1(new_n375_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n376_) );
  NAND2_X1 g0240 ( .A1(new_n376_), .A2(new_n369_), .ZN(new_n377_) );
  INV_X1 g0241 ( .A(G169), .ZN(new_n378_) );
  NOR2_X1 g0242 ( .A1(new_n372_), .A2(new_n370_), .ZN(new_n379_) );
  NAND3_X1 g0243 ( .A1(new_n379_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n380_) );
  NAND2_X1 g0244 ( .A1(new_n380_), .A2(new_n378_), .ZN(new_n381_) );
  NAND2_X1 g0245 ( .A1(new_n377_), .A2(new_n381_), .ZN(new_n382_) );
  INV_X1 g0246 ( .A(new_n382_), .ZN(new_n383_) );
  NAND2_X1 g0247 ( .A1(new_n383_), .A2(new_n368_), .ZN(new_n384_) );
  INV_X1 g0248 ( .A(KEYINPUT27), .ZN(new_n385_) );
  NAND2_X1 g0249 ( .A1(new_n380_), .A2(G200), .ZN(new_n386_) );
  NAND2_X1 g0250 ( .A1(new_n386_), .A2(new_n385_), .ZN(new_n387_) );
  NAND3_X1 g0251 ( .A1(new_n380_), .A2(G200), .A3(KEYINPUT27), .ZN(new_n388_) );
  NAND2_X1 g0252 ( .A1(new_n387_), .A2(new_n388_), .ZN(new_n389_) );
  NAND4_X1 g0253 ( .A1(new_n379_), .A2(G190), .A3(new_n373_), .A4(new_n374_), .ZN(new_n390_) );
  NAND2_X1 g0254 ( .A1(new_n390_), .A2(KEYINPUT28), .ZN(new_n391_) );
  INV_X1 g0255 ( .A(KEYINPUT28), .ZN(new_n392_) );
  NAND3_X1 g0256 ( .A1(new_n376_), .A2(G190), .A3(new_n392_), .ZN(new_n393_) );
  NAND2_X1 g0257 ( .A1(new_n393_), .A2(new_n391_), .ZN(new_n394_) );
  NAND4_X1 g0258 ( .A1(new_n389_), .A2(new_n394_), .A3(new_n361_), .A4(new_n367_), .ZN(new_n395_) );
  NAND2_X1 g0259 ( .A1(new_n395_), .A2(new_n384_), .ZN(new_n396_) );
  INV_X1 g0260 ( .A(new_n396_), .ZN(new_n397_) );
  NAND2_X1 g0261 ( .A1(new_n345_), .A2(G50), .ZN(new_n398_) );
  NAND2_X1 g0262 ( .A1(new_n249_), .A2(new_n138_), .ZN(new_n399_) );
  INV_X1 g0263 ( .A(new_n259_), .ZN(new_n400_) );
  NAND2_X1 g0264 ( .A1(new_n400_), .A2(G150), .ZN(new_n401_) );
  NAND2_X1 g0265 ( .A1(new_n263_), .A2(new_n139_), .ZN(new_n402_) );
  NAND2_X1 g0266 ( .A1(new_n267_), .A2(G58), .ZN(new_n403_) );
  NAND4_X1 g0267 ( .A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_) );
  INV_X1 g0268 ( .A(new_n404_), .ZN(new_n405_) );
  NAND2_X1 g0269 ( .A1(new_n405_), .A2(new_n398_), .ZN(new_n406_) );
  INV_X1 g0270 ( .A(G223), .ZN(new_n407_) );
  NOR2_X1 g0271 ( .A1(new_n275_), .A2(new_n407_), .ZN(new_n408_) );
  NAND2_X1 g0272 ( .A1(new_n304_), .A2(G226), .ZN(new_n409_) );
  INV_X1 g0273 ( .A(new_n409_), .ZN(new_n410_) );
  NAND3_X1 g0274 ( .A1(new_n177_), .A2(G77), .A3(new_n296_), .ZN(new_n411_) );
  NAND2_X1 g0275 ( .A1(new_n411_), .A2(new_n294_), .ZN(new_n412_) );
  NOR3_X1 g0276 ( .A1(new_n410_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n413_) );
  INV_X1 g0277 ( .A(KEYINPUT36), .ZN(new_n414_) );
  NAND2_X1 g0278 ( .A1(new_n284_), .A2(G222), .ZN(new_n415_) );
  NAND2_X1 g0279 ( .A1(new_n415_), .A2(new_n414_), .ZN(new_n416_) );
  NAND3_X1 g0280 ( .A1(new_n284_), .A2(G222), .A3(KEYINPUT36), .ZN(new_n417_) );
  NAND3_X1 g0281 ( .A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_) );
  INV_X1 g0282 ( .A(new_n418_), .ZN(new_n419_) );
  NAND2_X1 g0283 ( .A1(new_n419_), .A2(new_n369_), .ZN(new_n420_) );
  NAND2_X1 g0284 ( .A1(new_n418_), .A2(new_n378_), .ZN(new_n421_) );
  NAND3_X1 g0285 ( .A1(new_n406_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_) );
  NAND2_X1 g0286 ( .A1(new_n419_), .A2(G190), .ZN(new_n423_) );
  NAND2_X1 g0287 ( .A1(new_n418_), .A2(G200), .ZN(new_n424_) );
  NAND4_X1 g0288 ( .A1(new_n423_), .A2(new_n405_), .A3(new_n398_), .A4(new_n424_), .ZN(new_n425_) );
  NAND2_X1 g0289 ( .A1(new_n422_), .A2(new_n425_), .ZN(new_n426_) );
  NAND2_X1 g0290 ( .A1(new_n426_), .A2(KEYINPUT37), .ZN(new_n427_) );
  INV_X1 g0291 ( .A(KEYINPUT37), .ZN(new_n428_) );
  NAND3_X1 g0292 ( .A1(new_n422_), .A2(new_n428_), .A3(new_n425_), .ZN(new_n429_) );
  NAND2_X1 g0293 ( .A1(new_n427_), .A2(new_n429_), .ZN(new_n430_) );
  NAND4_X1 g0294 ( .A1(new_n430_), .A2(new_n358_), .A3(new_n324_), .A4(new_n397_), .ZN(new_n431_) );
  NOR2_X1 g0295 ( .A1(new_n431_), .A2(new_n317_), .ZN(new_n432_) );
  INV_X1 g0296 ( .A(new_n432_), .ZN(new_n433_) );
  INV_X1 g0297 ( .A(KEYINPUT0), .ZN(new_n434_) );
  NAND4_X1 g0298 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n296_), .A4(G294), .ZN(new_n435_) );
  NAND2_X1 g0299 ( .A1(new_n435_), .A2(KEYINPUT14), .ZN(new_n436_) );
  INV_X1 g0300 ( .A(new_n436_), .ZN(new_n437_) );
  NOR2_X1 g0301 ( .A1(new_n435_), .A2(KEYINPUT14), .ZN(new_n438_) );
  NOR2_X1 g0302 ( .A1(new_n437_), .A2(new_n438_), .ZN(new_n439_) );
  NAND2_X1 g0303 ( .A1(new_n284_), .A2(G250), .ZN(new_n440_) );
  NAND4_X1 g0304 ( .A1(new_n177_), .A2(new_n258_), .A3(G257), .A4(G1698), .ZN(new_n441_) );
  NOR3_X1 g0305 ( .A1(new_n292_), .A2(G1), .A3(G41), .ZN(new_n442_) );
  NAND2_X1 g0306 ( .A1(new_n442_), .A2(G274), .ZN(new_n443_) );
  INV_X1 g0307 ( .A(new_n442_), .ZN(new_n444_) );
  NAND3_X1 g0308 ( .A1(new_n302_), .A2(G264), .A3(new_n444_), .ZN(new_n445_) );
  NAND4_X1 g0309 ( .A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_) );
  NOR2_X1 g0310 ( .A1(new_n446_), .A2(new_n439_), .ZN(new_n447_) );
  NAND3_X1 g0311 ( .A1(new_n447_), .A2(new_n369_), .A3(KEYINPUT15), .ZN(new_n448_) );
  INV_X1 g0312 ( .A(KEYINPUT15), .ZN(new_n449_) );
  INV_X1 g0313 ( .A(new_n438_), .ZN(new_n450_) );
  NAND2_X1 g0314 ( .A1(new_n450_), .A2(new_n436_), .ZN(new_n451_) );
  NOR2_X1 g0315 ( .A1(new_n275_), .A2(new_n168_), .ZN(new_n452_) );
  NAND2_X1 g0316 ( .A1(new_n445_), .A2(new_n443_), .ZN(new_n453_) );
  NOR2_X1 g0317 ( .A1(new_n453_), .A2(new_n452_), .ZN(new_n454_) );
  NAND4_X1 g0318 ( .A1(new_n454_), .A2(new_n451_), .A3(new_n369_), .A4(new_n440_), .ZN(new_n455_) );
  NAND2_X1 g0319 ( .A1(new_n455_), .A2(new_n449_), .ZN(new_n456_) );
  NAND2_X1 g0320 ( .A1(new_n448_), .A2(new_n456_), .ZN(new_n457_) );
  INV_X1 g0321 ( .A(new_n447_), .ZN(new_n458_) );
  NAND2_X1 g0322 ( .A1(new_n458_), .A2(new_n378_), .ZN(new_n459_) );
  INV_X1 g0323 ( .A(G107), .ZN(new_n460_) );
  NAND2_X1 g0324 ( .A1(new_n360_), .A2(new_n460_), .ZN(new_n461_) );
  NAND2_X1 g0325 ( .A1(new_n400_), .A2(G87), .ZN(new_n462_) );
  NAND4_X1 g0326 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n265_), .A4(G116), .ZN(new_n463_) );
  NAND2_X1 g0327 ( .A1(new_n463_), .A2(KEYINPUT16), .ZN(new_n464_) );
  INV_X1 g0328 ( .A(KEYINPUT16), .ZN(new_n465_) );
  NAND4_X1 g0329 ( .A1(new_n177_), .A2(G116), .A3(new_n465_), .A4(new_n265_), .ZN(new_n466_) );
  NAND2_X1 g0330 ( .A1(new_n466_), .A2(new_n464_), .ZN(new_n467_) );
  NAND2_X1 g0331 ( .A1(new_n252_), .A2(G33), .ZN(new_n468_) );
  NAND2_X1 g0332 ( .A1(new_n262_), .A2(new_n468_), .ZN(new_n469_) );
  INV_X1 g0333 ( .A(new_n469_), .ZN(new_n470_) );
  NAND4_X1 g0334 ( .A1(new_n470_), .A2(G107), .A3(new_n242_), .A4(new_n176_), .ZN(new_n471_) );
  NAND2_X1 g0335 ( .A1(new_n467_), .A2(new_n471_), .ZN(new_n472_) );
  NAND2_X1 g0336 ( .A1(new_n472_), .A2(KEYINPUT17), .ZN(new_n473_) );
  INV_X1 g0337 ( .A(KEYINPUT17), .ZN(new_n474_) );
  NAND3_X1 g0338 ( .A1(new_n467_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_) );
  NAND2_X1 g0339 ( .A1(new_n473_), .A2(new_n475_), .ZN(new_n476_) );
  NAND3_X1 g0340 ( .A1(new_n461_), .A2(new_n476_), .A3(new_n462_), .ZN(new_n477_) );
  NAND3_X1 g0341 ( .A1(new_n477_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n478_) );
  INV_X1 g0342 ( .A(G200), .ZN(new_n479_) );
  NOR2_X1 g0343 ( .A1(new_n447_), .A2(new_n479_), .ZN(new_n480_) );
  INV_X1 g0344 ( .A(G190), .ZN(new_n481_) );
  NOR3_X1 g0345 ( .A1(new_n446_), .A2(new_n439_), .A3(new_n481_), .ZN(new_n482_) );
  NOR2_X1 g0346 ( .A1(new_n480_), .A2(new_n482_), .ZN(new_n483_) );
  NAND4_X1 g0347 ( .A1(new_n483_), .A2(new_n461_), .A3(new_n462_), .A4(new_n476_), .ZN(new_n484_) );
  NAND2_X1 g0348 ( .A1(new_n484_), .A2(new_n478_), .ZN(new_n485_) );
  NAND2_X1 g0349 ( .A1(new_n485_), .A2(new_n434_), .ZN(new_n486_) );
  NAND3_X1 g0350 ( .A1(new_n484_), .A2(new_n478_), .A3(KEYINPUT0), .ZN(new_n487_) );
  NAND2_X1 g0351 ( .A1(new_n486_), .A2(new_n487_), .ZN(new_n488_) );
  INV_X1 g0352 ( .A(new_n488_), .ZN(new_n489_) );
  NOR2_X1 g0353 ( .A1(new_n243_), .A2(new_n469_), .ZN(new_n490_) );
  NAND2_X1 g0354 ( .A1(new_n490_), .A2(G87), .ZN(new_n491_) );
  NAND2_X1 g0355 ( .A1(new_n248_), .A2(new_n491_), .ZN(new_n492_) );
  INV_X1 g0356 ( .A(G97), .ZN(new_n493_) );
  NAND3_X1 g0357 ( .A1(new_n218_), .A2(new_n493_), .A3(new_n460_), .ZN(new_n494_) );
  NAND2_X1 g0358 ( .A1(new_n492_), .A2(new_n494_), .ZN(new_n495_) );
  NAND2_X1 g0359 ( .A1(new_n495_), .A2(KEYINPUT9), .ZN(new_n496_) );
  INV_X1 g0360 ( .A(KEYINPUT9), .ZN(new_n497_) );
  NAND3_X1 g0361 ( .A1(new_n492_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n498_) );
  NOR2_X1 g0362 ( .A1(new_n259_), .A2(new_n359_), .ZN(new_n499_) );
  NAND2_X1 g0363 ( .A1(new_n267_), .A2(G97), .ZN(new_n500_) );
  NAND2_X1 g0364 ( .A1(new_n263_), .A2(new_n218_), .ZN(new_n501_) );
  NAND2_X1 g0365 ( .A1(new_n500_), .A2(new_n501_), .ZN(new_n502_) );
  NOR2_X1 g0366 ( .A1(new_n502_), .A2(new_n499_), .ZN(new_n503_) );
  NAND2_X1 g0367 ( .A1(new_n498_), .A2(new_n503_), .ZN(new_n504_) );
  INV_X1 g0368 ( .A(new_n504_), .ZN(new_n505_) );
  NAND2_X1 g0369 ( .A1(new_n505_), .A2(new_n496_), .ZN(new_n506_) );
  INV_X1 g0370 ( .A(KEYINPUT8), .ZN(new_n507_) );
  INV_X1 g0371 ( .A(G244), .ZN(new_n508_) );
  NOR2_X1 g0372 ( .A1(new_n275_), .A2(new_n508_), .ZN(new_n509_) );
  NOR2_X1 g0373 ( .A1(new_n283_), .A2(new_n184_), .ZN(new_n510_) );
  NOR2_X1 g0374 ( .A1(new_n509_), .A2(new_n510_), .ZN(new_n511_) );
  NAND2_X1 g0375 ( .A1(new_n511_), .A2(new_n507_), .ZN(new_n512_) );
  INV_X1 g0376 ( .A(new_n512_), .ZN(new_n513_) );
  NOR2_X1 g0377 ( .A1(new_n511_), .A2(new_n507_), .ZN(new_n514_) );
  NAND2_X1 g0378 ( .A1(new_n252_), .A2(G45), .ZN(new_n515_) );
  NAND3_X1 g0379 ( .A1(new_n302_), .A2(G250), .A3(new_n515_), .ZN(new_n516_) );
  NAND3_X1 g0380 ( .A1(new_n252_), .A2(G45), .A3(G274), .ZN(new_n517_) );
  NAND3_X1 g0381 ( .A1(new_n177_), .A2(G116), .A3(new_n296_), .ZN(new_n518_) );
  NAND3_X1 g0382 ( .A1(new_n518_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n519_) );
  NOR3_X1 g0383 ( .A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_) );
  INV_X1 g0384 ( .A(new_n520_), .ZN(new_n521_) );
  NAND2_X1 g0385 ( .A1(new_n521_), .A2(G169), .ZN(new_n522_) );
  NAND2_X1 g0386 ( .A1(new_n520_), .A2(G179), .ZN(new_n523_) );
  NAND2_X1 g0387 ( .A1(new_n522_), .A2(new_n523_), .ZN(new_n524_) );
  NAND2_X1 g0388 ( .A1(new_n524_), .A2(new_n506_), .ZN(new_n525_) );
  NAND2_X1 g0389 ( .A1(new_n520_), .A2(G190), .ZN(new_n526_) );
  NAND2_X1 g0390 ( .A1(new_n521_), .A2(G200), .ZN(new_n527_) );
  NAND4_X1 g0391 ( .A1(new_n527_), .A2(new_n505_), .A3(new_n496_), .A4(new_n526_), .ZN(new_n528_) );
  NAND2_X1 g0392 ( .A1(new_n525_), .A2(new_n528_), .ZN(new_n529_) );
  INV_X1 g0393 ( .A(KEYINPUT12), .ZN(new_n530_) );
  NOR2_X1 g0394 ( .A1(new_n275_), .A2(new_n200_), .ZN(new_n531_) );
  INV_X1 g0395 ( .A(new_n531_), .ZN(new_n532_) );
  NOR2_X1 g0396 ( .A1(new_n283_), .A2(new_n508_), .ZN(new_n533_) );
  NAND4_X1 g0397 ( .A1(new_n173_), .A2(new_n175_), .A3(new_n296_), .A4(G283), .ZN(new_n534_) );
  NAND2_X1 g0398 ( .A1(new_n534_), .A2(new_n443_), .ZN(new_n535_) );
  NOR2_X1 g0399 ( .A1(new_n533_), .A2(new_n535_), .ZN(new_n536_) );
  NAND3_X1 g0400 ( .A1(new_n536_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n537_) );
  INV_X1 g0401 ( .A(new_n302_), .ZN(new_n538_) );
  NOR3_X1 g0402 ( .A1(new_n538_), .A2(new_n168_), .A3(new_n442_), .ZN(new_n539_) );
  INV_X1 g0403 ( .A(new_n539_), .ZN(new_n540_) );
  NAND2_X1 g0404 ( .A1(new_n536_), .A2(new_n532_), .ZN(new_n541_) );
  NAND2_X1 g0405 ( .A1(new_n541_), .A2(KEYINPUT12), .ZN(new_n542_) );
  NAND3_X1 g0406 ( .A1(new_n542_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n543_) );
  INV_X1 g0407 ( .A(new_n543_), .ZN(new_n544_) );
  NAND2_X1 g0408 ( .A1(new_n544_), .A2(G190), .ZN(new_n545_) );
  NAND2_X1 g0409 ( .A1(new_n543_), .A2(G200), .ZN(new_n546_) );
  NAND3_X1 g0410 ( .A1(new_n245_), .A2(new_n213_), .A3(new_n247_), .ZN(new_n547_) );
  INV_X1 g0411 ( .A(KEYINPUT13), .ZN(new_n548_) );
  NAND2_X1 g0412 ( .A1(new_n267_), .A2(G107), .ZN(new_n549_) );
  NAND2_X1 g0413 ( .A1(new_n263_), .A2(new_n493_), .ZN(new_n550_) );
  NAND2_X1 g0414 ( .A1(new_n549_), .A2(new_n550_), .ZN(new_n551_) );
  NAND2_X1 g0415 ( .A1(new_n551_), .A2(new_n548_), .ZN(new_n552_) );
  NAND2_X1 g0416 ( .A1(new_n400_), .A2(G77), .ZN(new_n553_) );
  NAND2_X1 g0417 ( .A1(new_n552_), .A2(new_n553_), .ZN(new_n554_) );
  NAND3_X1 g0418 ( .A1(new_n549_), .A2(KEYINPUT13), .A3(new_n550_), .ZN(new_n555_) );
  NAND2_X1 g0419 ( .A1(new_n490_), .A2(G97), .ZN(new_n556_) );
  NAND2_X1 g0420 ( .A1(new_n555_), .A2(new_n556_), .ZN(new_n557_) );
  NOR2_X1 g0421 ( .A1(new_n554_), .A2(new_n557_), .ZN(new_n558_) );
  NAND4_X1 g0422 ( .A1(new_n545_), .A2(new_n546_), .A3(new_n558_), .A4(new_n547_), .ZN(new_n559_) );
  INV_X1 g0423 ( .A(new_n557_), .ZN(new_n560_) );
  NAND4_X1 g0424 ( .A1(new_n560_), .A2(new_n547_), .A3(new_n552_), .A4(new_n553_), .ZN(new_n561_) );
  NAND2_X1 g0425 ( .A1(new_n544_), .A2(new_n369_), .ZN(new_n562_) );
  NAND2_X1 g0426 ( .A1(new_n543_), .A2(new_n378_), .ZN(new_n563_) );
  NAND3_X1 g0427 ( .A1(new_n562_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_) );
  NAND2_X1 g0428 ( .A1(new_n559_), .A2(new_n564_), .ZN(new_n565_) );
  INV_X1 g0429 ( .A(new_n565_), .ZN(new_n566_) );
  INV_X1 g0430 ( .A(KEYINPUT11), .ZN(new_n567_) );
  NAND3_X1 g0431 ( .A1(new_n302_), .A2(G270), .A3(new_n444_), .ZN(new_n568_) );
  NAND2_X1 g0432 ( .A1(new_n568_), .A2(KEYINPUT10), .ZN(new_n569_) );
  INV_X1 g0433 ( .A(KEYINPUT10), .ZN(new_n570_) );
  NAND4_X1 g0434 ( .A1(new_n302_), .A2(new_n444_), .A3(G270), .A4(new_n570_), .ZN(new_n571_) );
  NAND2_X1 g0435 ( .A1(new_n569_), .A2(new_n571_), .ZN(new_n572_) );
  NAND2_X1 g0436 ( .A1(new_n284_), .A2(G257), .ZN(new_n573_) );
  NOR2_X1 g0437 ( .A1(new_n275_), .A2(new_n169_), .ZN(new_n574_) );
  NAND3_X1 g0438 ( .A1(new_n177_), .A2(G303), .A3(new_n296_), .ZN(new_n575_) );
  NAND2_X1 g0439 ( .A1(new_n575_), .A2(new_n443_), .ZN(new_n576_) );
  NOR2_X1 g0440 ( .A1(new_n576_), .A2(new_n574_), .ZN(new_n577_) );
  NAND3_X1 g0441 ( .A1(new_n577_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n578_) );
  NAND2_X1 g0442 ( .A1(new_n578_), .A2(G169), .ZN(new_n579_) );
  NAND4_X1 g0443 ( .A1(new_n577_), .A2(G179), .A3(new_n572_), .A4(new_n573_), .ZN(new_n580_) );
  NAND2_X1 g0444 ( .A1(new_n579_), .A2(new_n580_), .ZN(new_n581_) );
  INV_X1 g0445 ( .A(new_n490_), .ZN(new_n582_) );
  NAND2_X1 g0446 ( .A1(new_n248_), .A2(new_n582_), .ZN(new_n583_) );
  NAND2_X1 g0447 ( .A1(new_n583_), .A2(G116), .ZN(new_n584_) );
  NOR2_X1 g0448 ( .A1(new_n259_), .A2(new_n493_), .ZN(new_n585_) );
  NAND2_X1 g0449 ( .A1(new_n267_), .A2(G283), .ZN(new_n586_) );
  NAND2_X1 g0450 ( .A1(new_n263_), .A2(new_n220_), .ZN(new_n587_) );
  NAND2_X1 g0451 ( .A1(new_n586_), .A2(new_n587_), .ZN(new_n588_) );
  NOR2_X1 g0452 ( .A1(new_n588_), .A2(new_n585_), .ZN(new_n589_) );
  NAND2_X1 g0453 ( .A1(new_n584_), .A2(new_n589_), .ZN(new_n590_) );
  NAND2_X1 g0454 ( .A1(new_n581_), .A2(new_n590_), .ZN(new_n591_) );
  NAND4_X1 g0455 ( .A1(new_n577_), .A2(G190), .A3(new_n572_), .A4(new_n573_), .ZN(new_n592_) );
  NAND2_X1 g0456 ( .A1(new_n578_), .A2(G200), .ZN(new_n593_) );
  NAND4_X1 g0457 ( .A1(new_n593_), .A2(new_n584_), .A3(new_n589_), .A4(new_n592_), .ZN(new_n594_) );
  NAND2_X1 g0458 ( .A1(new_n591_), .A2(new_n594_), .ZN(new_n595_) );
  NAND2_X1 g0459 ( .A1(new_n595_), .A2(new_n567_), .ZN(new_n596_) );
  NAND3_X1 g0460 ( .A1(new_n591_), .A2(KEYINPUT11), .A3(new_n594_), .ZN(new_n597_) );
  NAND3_X1 g0461 ( .A1(new_n566_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_) );
  NOR4_X1 g0462 ( .A1(new_n433_), .A2(new_n489_), .A3(new_n529_), .A4(new_n598_), .ZN(G372) );
  NAND4_X1 g0463 ( .A1(new_n395_), .A2(new_n343_), .A3(new_n352_), .A4(new_n384_), .ZN(new_n600_) );
  NAND2_X1 g0464 ( .A1(new_n600_), .A2(new_n384_), .ZN(new_n601_) );
  NAND2_X1 g0465 ( .A1(new_n324_), .A2(new_n601_), .ZN(new_n602_) );
  NAND2_X1 g0466 ( .A1(new_n602_), .A2(new_n316_), .ZN(new_n603_) );
  NAND2_X1 g0467 ( .A1(new_n603_), .A2(new_n430_), .ZN(new_n604_) );
  NAND2_X1 g0468 ( .A1(new_n604_), .A2(new_n422_), .ZN(new_n605_) );
  INV_X1 g0469 ( .A(new_n605_), .ZN(new_n606_) );
  INV_X1 g0470 ( .A(new_n591_), .ZN(new_n607_) );
  NAND2_X1 g0471 ( .A1(new_n488_), .A2(new_n607_), .ZN(new_n608_) );
  NAND2_X1 g0472 ( .A1(new_n608_), .A2(new_n478_), .ZN(new_n609_) );
  NAND2_X1 g0473 ( .A1(new_n609_), .A2(new_n566_), .ZN(new_n610_) );
  NAND2_X1 g0474 ( .A1(new_n525_), .A2(new_n564_), .ZN(new_n611_) );
  INV_X1 g0475 ( .A(new_n611_), .ZN(new_n612_) );
  NAND2_X1 g0476 ( .A1(new_n610_), .A2(new_n612_), .ZN(new_n613_) );
  NAND3_X1 g0477 ( .A1(new_n432_), .A2(new_n613_), .A3(new_n528_), .ZN(new_n614_) );
  NAND2_X1 g0478 ( .A1(new_n614_), .A2(new_n606_), .ZN(G369) );
  INV_X1 g0479 ( .A(G343), .ZN(new_n616_) );
  NAND4_X1 g0480 ( .A1(new_n252_), .A2(new_n257_), .A3(G13), .A4(G213), .ZN(new_n617_) );
  NOR2_X1 g0481 ( .A1(new_n617_), .A2(new_n616_), .ZN(new_n618_) );
  NAND2_X1 g0482 ( .A1(new_n477_), .A2(new_n618_), .ZN(new_n619_) );
  NAND2_X1 g0483 ( .A1(new_n488_), .A2(new_n619_), .ZN(new_n620_) );
  NAND4_X1 g0484 ( .A1(new_n477_), .A2(new_n457_), .A3(new_n459_), .A4(new_n618_), .ZN(new_n621_) );
  NAND2_X1 g0485 ( .A1(new_n620_), .A2(new_n621_), .ZN(new_n622_) );
  INV_X1 g0486 ( .A(new_n622_), .ZN(new_n623_) );
  NAND2_X1 g0487 ( .A1(new_n590_), .A2(new_n618_), .ZN(new_n624_) );
  NAND3_X1 g0488 ( .A1(new_n596_), .A2(new_n597_), .A3(new_n624_), .ZN(new_n625_) );
  NAND2_X1 g0489 ( .A1(new_n607_), .A2(new_n618_), .ZN(new_n626_) );
  NAND2_X1 g0490 ( .A1(new_n625_), .A2(new_n626_), .ZN(new_n627_) );
  NAND2_X1 g0491 ( .A1(new_n627_), .A2(G330), .ZN(new_n628_) );
  NOR2_X1 g0492 ( .A1(new_n623_), .A2(new_n628_), .ZN(new_n629_) );
  INV_X1 g0493 ( .A(new_n629_), .ZN(new_n630_) );
  INV_X1 g0494 ( .A(new_n618_), .ZN(new_n631_) );
  NAND2_X1 g0495 ( .A1(new_n609_), .A2(new_n631_), .ZN(new_n632_) );
  NAND2_X1 g0496 ( .A1(new_n630_), .A2(new_n632_), .ZN(G399) );
  INV_X1 g0497 ( .A(new_n580_), .ZN(new_n634_) );
  INV_X1 g0498 ( .A(KEYINPUT18), .ZN(new_n635_) );
  NAND2_X1 g0499 ( .A1(new_n544_), .A2(new_n520_), .ZN(new_n636_) );
  NAND2_X1 g0500 ( .A1(new_n636_), .A2(new_n635_), .ZN(new_n637_) );
  NAND3_X1 g0501 ( .A1(new_n544_), .A2(KEYINPUT18), .A3(new_n520_), .ZN(new_n638_) );
  NAND2_X1 g0502 ( .A1(new_n637_), .A2(new_n638_), .ZN(new_n639_) );
  NAND3_X1 g0503 ( .A1(new_n639_), .A2(new_n447_), .A3(new_n634_), .ZN(new_n640_) );
  NAND2_X1 g0504 ( .A1(new_n578_), .A2(new_n369_), .ZN(new_n641_) );
  INV_X1 g0505 ( .A(new_n641_), .ZN(new_n642_) );
  NAND4_X1 g0506 ( .A1(new_n521_), .A2(new_n642_), .A3(new_n458_), .A4(new_n543_), .ZN(new_n643_) );
  NAND2_X1 g0507 ( .A1(new_n640_), .A2(new_n643_), .ZN(new_n644_) );
  NAND2_X1 g0508 ( .A1(new_n644_), .A2(new_n618_), .ZN(new_n645_) );
  NOR2_X1 g0509 ( .A1(new_n598_), .A2(new_n529_), .ZN(new_n646_) );
  NAND3_X1 g0510 ( .A1(new_n646_), .A2(new_n488_), .A3(new_n631_), .ZN(new_n647_) );
  NAND2_X1 g0511 ( .A1(new_n647_), .A2(new_n645_), .ZN(new_n648_) );
  NAND2_X1 g0512 ( .A1(new_n648_), .A2(G330), .ZN(new_n649_) );
  NAND3_X1 g0513 ( .A1(new_n613_), .A2(new_n528_), .A3(new_n631_), .ZN(new_n650_) );
  NAND2_X1 g0514 ( .A1(new_n650_), .A2(new_n649_), .ZN(new_n651_) );
  NAND2_X1 g0515 ( .A1(new_n651_), .A2(new_n252_), .ZN(new_n652_) );
  INV_X1 g0516 ( .A(new_n167_), .ZN(new_n653_) );
  NOR2_X1 g0517 ( .A1(new_n653_), .A2(G41), .ZN(new_n654_) );
  NAND2_X1 g0518 ( .A1(new_n654_), .A2(new_n180_), .ZN(new_n655_) );
  INV_X1 g0519 ( .A(new_n654_), .ZN(new_n656_) );
  NOR2_X1 g0520 ( .A1(new_n494_), .A2(G116), .ZN(new_n657_) );
  NAND3_X1 g0521 ( .A1(new_n656_), .A2(G1), .A3(new_n657_), .ZN(new_n658_) );
  NAND3_X1 g0522 ( .A1(new_n652_), .A2(new_n655_), .A3(new_n658_), .ZN(G364) );
  INV_X1 g0523 ( .A(new_n627_), .ZN(new_n660_) );
  NOR2_X1 g0524 ( .A1(G13), .A2(G33), .ZN(new_n661_) );
  INV_X1 g0525 ( .A(new_n661_), .ZN(new_n662_) );
  NOR2_X1 g0526 ( .A1(new_n662_), .A2(G20), .ZN(new_n663_) );
  NAND3_X1 g0527 ( .A1(new_n660_), .A2(KEYINPUT62), .A3(new_n663_), .ZN(new_n664_) );
  INV_X1 g0528 ( .A(KEYINPUT62), .ZN(new_n665_) );
  NAND2_X1 g0529 ( .A1(new_n660_), .A2(new_n663_), .ZN(new_n666_) );
  NAND2_X1 g0530 ( .A1(new_n666_), .A2(new_n665_), .ZN(new_n667_) );
  INV_X1 g0531 ( .A(KEYINPUT24), .ZN(new_n668_) );
  NAND2_X1 g0532 ( .A1(new_n167_), .A2(G33), .ZN(new_n669_) );
  NAND2_X1 g0533 ( .A1(new_n669_), .A2(new_n668_), .ZN(new_n670_) );
  NAND3_X1 g0534 ( .A1(new_n167_), .A2(G33), .A3(KEYINPUT24), .ZN(new_n671_) );
  NAND2_X1 g0535 ( .A1(new_n670_), .A2(new_n671_), .ZN(new_n672_) );
  NAND2_X1 g0536 ( .A1(new_n180_), .A2(new_n292_), .ZN(new_n673_) );
  NAND2_X1 g0537 ( .A1(new_n233_), .A2(G45), .ZN(new_n674_) );
  NAND3_X1 g0538 ( .A1(new_n674_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n675_) );
  NAND3_X1 g0539 ( .A1(new_n653_), .A2(new_n220_), .A3(KEYINPUT60), .ZN(new_n676_) );
  INV_X1 g0540 ( .A(KEYINPUT60), .ZN(new_n677_) );
  NAND2_X1 g0541 ( .A1(new_n653_), .A2(new_n220_), .ZN(new_n678_) );
  NAND2_X1 g0542 ( .A1(new_n678_), .A2(new_n677_), .ZN(new_n679_) );
  NAND2_X1 g0543 ( .A1(G355), .A2(new_n661_), .ZN(new_n680_) );
  NAND4_X1 g0544 ( .A1(new_n675_), .A2(new_n676_), .A3(new_n679_), .A4(new_n680_), .ZN(new_n681_) );
  INV_X1 g0545 ( .A(new_n663_), .ZN(new_n682_) );
  NAND2_X1 g0546 ( .A1(new_n378_), .A2(G20), .ZN(new_n683_) );
  NAND2_X1 g0547 ( .A1(new_n177_), .A2(new_n683_), .ZN(new_n684_) );
  NAND2_X1 g0548 ( .A1(new_n684_), .A2(new_n682_), .ZN(new_n685_) );
  INV_X1 g0549 ( .A(new_n685_), .ZN(new_n686_) );
  NAND2_X1 g0550 ( .A1(new_n681_), .A2(new_n686_), .ZN(new_n687_) );
  INV_X1 g0551 ( .A(new_n687_), .ZN(new_n688_) );
  NAND2_X1 g0552 ( .A1(G20), .A2(G179), .ZN(new_n689_) );
  NOR3_X1 g0553 ( .A1(new_n689_), .A2(G190), .A3(G200), .ZN(new_n690_) );
  INV_X1 g0554 ( .A(new_n690_), .ZN(new_n691_) );
  NOR2_X1 g0555 ( .A1(new_n691_), .A2(new_n140_), .ZN(new_n692_) );
  NOR2_X1 g0556 ( .A1(new_n257_), .A2(G179), .ZN(new_n693_) );
  NAND3_X1 g0557 ( .A1(new_n693_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n694_) );
  NOR2_X1 g0558 ( .A1(new_n694_), .A2(new_n256_), .ZN(new_n695_) );
  NOR2_X1 g0559 ( .A1(new_n481_), .A2(G200), .ZN(new_n696_) );
  INV_X1 g0560 ( .A(new_n696_), .ZN(new_n697_) );
  NOR2_X1 g0561 ( .A1(new_n697_), .A2(G179), .ZN(new_n698_) );
  NOR2_X1 g0562 ( .A1(new_n698_), .A2(new_n257_), .ZN(new_n699_) );
  NOR2_X1 g0563 ( .A1(new_n699_), .A2(new_n493_), .ZN(new_n700_) );
  NOR3_X1 g0564 ( .A1(new_n689_), .A2(new_n479_), .A3(G190), .ZN(new_n701_) );
  INV_X1 g0565 ( .A(new_n701_), .ZN(new_n702_) );
  NOR2_X1 g0566 ( .A1(new_n702_), .A2(new_n359_), .ZN(new_n703_) );
  NOR4_X1 g0567 ( .A1(new_n700_), .A2(new_n692_), .A3(new_n695_), .A4(new_n703_), .ZN(new_n704_) );
  NAND2_X1 g0568 ( .A1(new_n704_), .A2(KEYINPUT61), .ZN(new_n705_) );
  INV_X1 g0569 ( .A(KEYINPUT61), .ZN(new_n706_) );
  INV_X1 g0570 ( .A(new_n704_), .ZN(new_n707_) );
  NAND2_X1 g0571 ( .A1(new_n707_), .A2(new_n706_), .ZN(new_n708_) );
  INV_X1 g0572 ( .A(new_n684_), .ZN(new_n709_) );
  NAND2_X1 g0573 ( .A1(new_n709_), .A2(new_n258_), .ZN(new_n710_) );
  NAND3_X1 g0574 ( .A1(new_n693_), .A2(new_n481_), .A3(G200), .ZN(new_n711_) );
  NOR2_X1 g0575 ( .A1(new_n711_), .A2(new_n460_), .ZN(new_n712_) );
  NAND2_X1 g0576 ( .A1(G190), .A2(G200), .ZN(new_n713_) );
  NOR2_X1 g0577 ( .A1(new_n689_), .A2(new_n713_), .ZN(new_n714_) );
  NAND2_X1 g0578 ( .A1(new_n714_), .A2(G50), .ZN(new_n715_) );
  NOR3_X1 g0579 ( .A1(new_n713_), .A2(new_n257_), .A3(G179), .ZN(new_n716_) );
  INV_X1 g0580 ( .A(new_n716_), .ZN(new_n717_) );
  NOR2_X1 g0581 ( .A1(new_n717_), .A2(new_n218_), .ZN(new_n718_) );
  INV_X1 g0582 ( .A(new_n718_), .ZN(new_n719_) );
  NOR2_X1 g0583 ( .A1(new_n697_), .A2(new_n689_), .ZN(new_n720_) );
  NAND2_X1 g0584 ( .A1(new_n720_), .A2(G58), .ZN(new_n721_) );
  NAND3_X1 g0585 ( .A1(new_n719_), .A2(new_n715_), .A3(new_n721_), .ZN(new_n722_) );
  NOR3_X1 g0586 ( .A1(new_n722_), .A2(new_n710_), .A3(new_n712_), .ZN(new_n723_) );
  NAND3_X1 g0587 ( .A1(new_n708_), .A2(new_n705_), .A3(new_n723_), .ZN(new_n724_) );
  NAND3_X1 g0588 ( .A1(new_n257_), .A2(G13), .A3(G45), .ZN(new_n725_) );
  NAND2_X1 g0589 ( .A1(new_n725_), .A2(G1), .ZN(new_n726_) );
  NAND2_X1 g0590 ( .A1(new_n726_), .A2(KEYINPUT1), .ZN(new_n727_) );
  INV_X1 g0591 ( .A(KEYINPUT1), .ZN(new_n728_) );
  NAND3_X1 g0592 ( .A1(new_n725_), .A2(G1), .A3(new_n728_), .ZN(new_n729_) );
  NAND2_X1 g0593 ( .A1(new_n727_), .A2(new_n729_), .ZN(new_n730_) );
  NAND2_X1 g0594 ( .A1(new_n656_), .A2(new_n730_), .ZN(new_n731_) );
  INV_X1 g0595 ( .A(new_n731_), .ZN(new_n732_) );
  INV_X1 g0596 ( .A(new_n699_), .ZN(new_n733_) );
  NAND2_X1 g0597 ( .A1(new_n733_), .A2(G294), .ZN(new_n734_) );
  INV_X1 g0598 ( .A(new_n694_), .ZN(new_n735_) );
  NAND2_X1 g0599 ( .A1(new_n735_), .A2(G329), .ZN(new_n736_) );
  NAND2_X1 g0600 ( .A1(new_n690_), .A2(G311), .ZN(new_n737_) );
  NAND2_X1 g0601 ( .A1(new_n709_), .A2(G33), .ZN(new_n738_) );
  NAND2_X1 g0602 ( .A1(new_n716_), .A2(G303), .ZN(new_n739_) );
  NAND2_X1 g0603 ( .A1(new_n714_), .A2(G326), .ZN(new_n740_) );
  NAND2_X1 g0604 ( .A1(new_n720_), .A2(G322), .ZN(new_n741_) );
  NAND3_X1 g0605 ( .A1(new_n741_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n742_) );
  NAND2_X1 g0606 ( .A1(new_n701_), .A2(G317), .ZN(new_n743_) );
  INV_X1 g0607 ( .A(new_n711_), .ZN(new_n744_) );
  NAND2_X1 g0608 ( .A1(new_n744_), .A2(G283), .ZN(new_n745_) );
  NAND2_X1 g0609 ( .A1(new_n745_), .A2(new_n743_), .ZN(new_n746_) );
  NOR3_X1 g0610 ( .A1(new_n738_), .A2(new_n742_), .A3(new_n746_), .ZN(new_n747_) );
  NAND4_X1 g0611 ( .A1(new_n747_), .A2(new_n734_), .A3(new_n736_), .A4(new_n737_), .ZN(new_n748_) );
  NAND3_X1 g0612 ( .A1(new_n724_), .A2(new_n732_), .A3(new_n748_), .ZN(new_n749_) );
  NOR2_X1 g0613 ( .A1(new_n749_), .A2(new_n688_), .ZN(new_n750_) );
  NAND3_X1 g0614 ( .A1(new_n667_), .A2(new_n664_), .A3(new_n750_), .ZN(new_n751_) );
  INV_X1 g0615 ( .A(G330), .ZN(new_n752_) );
  NAND2_X1 g0616 ( .A1(new_n660_), .A2(new_n752_), .ZN(new_n753_) );
  NAND3_X1 g0617 ( .A1(new_n753_), .A2(new_n628_), .A3(new_n731_), .ZN(new_n754_) );
  NAND2_X1 g0618 ( .A1(new_n751_), .A2(new_n754_), .ZN(G396) );
  INV_X1 g0619 ( .A(new_n651_), .ZN(new_n756_) );
  NAND2_X1 g0620 ( .A1(new_n352_), .A2(new_n618_), .ZN(new_n757_) );
  NAND2_X1 g0621 ( .A1(new_n757_), .A2(KEYINPUT5), .ZN(new_n758_) );
  INV_X1 g0622 ( .A(KEYINPUT5), .ZN(new_n759_) );
  NAND3_X1 g0623 ( .A1(new_n352_), .A2(new_n759_), .A3(new_n618_), .ZN(new_n760_) );
  NAND2_X1 g0624 ( .A1(new_n758_), .A2(new_n760_), .ZN(new_n761_) );
  NAND2_X1 g0625 ( .A1(new_n761_), .A2(new_n343_), .ZN(new_n762_) );
  NAND4_X1 g0626 ( .A1(new_n353_), .A2(new_n356_), .A3(new_n758_), .A4(new_n760_), .ZN(new_n763_) );
  NAND2_X1 g0627 ( .A1(new_n763_), .A2(new_n762_), .ZN(new_n764_) );
  NAND2_X1 g0628 ( .A1(new_n756_), .A2(new_n764_), .ZN(new_n765_) );
  INV_X1 g0629 ( .A(new_n764_), .ZN(new_n766_) );
  NAND2_X1 g0630 ( .A1(new_n651_), .A2(new_n766_), .ZN(new_n767_) );
  NAND2_X1 g0631 ( .A1(new_n765_), .A2(new_n767_), .ZN(new_n768_) );
  NAND2_X1 g0632 ( .A1(new_n768_), .A2(new_n731_), .ZN(new_n769_) );
  NAND2_X1 g0633 ( .A1(new_n766_), .A2(new_n661_), .ZN(new_n770_) );
  NAND2_X1 g0634 ( .A1(new_n690_), .A2(G159), .ZN(new_n771_) );
  NAND2_X1 g0635 ( .A1(new_n733_), .A2(G58), .ZN(new_n772_) );
  NAND2_X1 g0636 ( .A1(new_n714_), .A2(G137), .ZN(new_n773_) );
  NAND2_X1 g0637 ( .A1(new_n716_), .A2(G50), .ZN(new_n774_) );
  NAND4_X1 g0638 ( .A1(new_n772_), .A2(new_n771_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_) );
  INV_X1 g0639 ( .A(new_n775_), .ZN(new_n776_) );
  NAND2_X1 g0640 ( .A1(new_n776_), .A2(KEYINPUT20), .ZN(new_n777_) );
  INV_X1 g0641 ( .A(KEYINPUT20), .ZN(new_n778_) );
  NAND2_X1 g0642 ( .A1(new_n775_), .A2(new_n778_), .ZN(new_n779_) );
  NAND2_X1 g0643 ( .A1(new_n777_), .A2(new_n779_), .ZN(new_n780_) );
  NAND2_X1 g0644 ( .A1(new_n744_), .A2(G68), .ZN(new_n781_) );
  NAND2_X1 g0645 ( .A1(new_n701_), .A2(G150), .ZN(new_n782_) );
  NAND2_X1 g0646 ( .A1(new_n720_), .A2(G143), .ZN(new_n783_) );
  NAND3_X1 g0647 ( .A1(new_n781_), .A2(new_n783_), .A3(new_n782_), .ZN(new_n784_) );
  INV_X1 g0648 ( .A(new_n784_), .ZN(new_n785_) );
  NAND2_X1 g0649 ( .A1(new_n735_), .A2(G132), .ZN(new_n786_) );
  NAND2_X1 g0650 ( .A1(new_n786_), .A2(KEYINPUT19), .ZN(new_n787_) );
  NOR2_X1 g0651 ( .A1(new_n786_), .A2(KEYINPUT19), .ZN(new_n788_) );
  NOR2_X1 g0652 ( .A1(new_n710_), .A2(new_n788_), .ZN(new_n789_) );
  NAND4_X1 g0653 ( .A1(new_n780_), .A2(new_n785_), .A3(new_n787_), .A4(new_n789_), .ZN(new_n790_) );
  NAND2_X1 g0654 ( .A1(new_n690_), .A2(G116), .ZN(new_n791_) );
  NAND2_X1 g0655 ( .A1(new_n791_), .A2(KEYINPUT21), .ZN(new_n792_) );
  NOR2_X1 g0656 ( .A1(new_n791_), .A2(KEYINPUT21), .ZN(new_n793_) );
  NAND2_X1 g0657 ( .A1(new_n714_), .A2(G303), .ZN(new_n794_) );
  NAND2_X1 g0658 ( .A1(new_n720_), .A2(G294), .ZN(new_n795_) );
  NAND2_X1 g0659 ( .A1(new_n716_), .A2(G107), .ZN(new_n796_) );
  NAND4_X1 g0660 ( .A1(new_n795_), .A2(new_n796_), .A3(G33), .A4(new_n794_), .ZN(new_n797_) );
  NOR2_X1 g0661 ( .A1(new_n797_), .A2(new_n793_), .ZN(new_n798_) );
  INV_X1 g0662 ( .A(KEYINPUT22), .ZN(new_n799_) );
  NOR2_X1 g0663 ( .A1(new_n711_), .A2(new_n218_), .ZN(new_n800_) );
  NOR2_X1 g0664 ( .A1(new_n800_), .A2(new_n799_), .ZN(new_n801_) );
  NAND2_X1 g0665 ( .A1(new_n800_), .A2(new_n799_), .ZN(new_n802_) );
  INV_X1 g0666 ( .A(new_n802_), .ZN(new_n803_) );
  NOR2_X1 g0667 ( .A1(new_n803_), .A2(new_n801_), .ZN(new_n804_) );
  INV_X1 g0668 ( .A(new_n804_), .ZN(new_n805_) );
  INV_X1 g0669 ( .A(G283), .ZN(new_n806_) );
  NOR2_X1 g0670 ( .A1(new_n702_), .A2(new_n806_), .ZN(new_n807_) );
  INV_X1 g0671 ( .A(G311), .ZN(new_n808_) );
  NOR2_X1 g0672 ( .A1(new_n694_), .A2(new_n808_), .ZN(new_n809_) );
  NOR4_X1 g0673 ( .A1(new_n700_), .A2(new_n684_), .A3(new_n807_), .A4(new_n809_), .ZN(new_n810_) );
  NAND4_X1 g0674 ( .A1(new_n810_), .A2(new_n805_), .A3(new_n792_), .A4(new_n798_), .ZN(new_n811_) );
  NAND2_X1 g0675 ( .A1(new_n684_), .A2(new_n662_), .ZN(new_n812_) );
  INV_X1 g0676 ( .A(new_n812_), .ZN(new_n813_) );
  NAND2_X1 g0677 ( .A1(new_n813_), .A2(new_n140_), .ZN(new_n814_) );
  NAND2_X1 g0678 ( .A1(new_n814_), .A2(new_n732_), .ZN(new_n815_) );
  INV_X1 g0679 ( .A(new_n815_), .ZN(new_n816_) );
  NAND4_X1 g0680 ( .A1(new_n770_), .A2(new_n790_), .A3(new_n811_), .A4(new_n816_), .ZN(new_n817_) );
  NAND2_X1 g0681 ( .A1(new_n769_), .A2(new_n817_), .ZN(G384) );
  NAND2_X1 g0682 ( .A1(new_n317_), .A2(new_n617_), .ZN(new_n819_) );
  NAND2_X1 g0683 ( .A1(new_n368_), .A2(new_n618_), .ZN(new_n820_) );
  NAND3_X1 g0684 ( .A1(new_n395_), .A2(new_n384_), .A3(new_n820_), .ZN(new_n821_) );
  INV_X1 g0685 ( .A(new_n384_), .ZN(new_n822_) );
  NAND2_X1 g0686 ( .A1(new_n822_), .A2(new_n618_), .ZN(new_n823_) );
  NAND2_X1 g0687 ( .A1(new_n821_), .A2(new_n823_), .ZN(new_n824_) );
  NAND2_X1 g0688 ( .A1(new_n824_), .A2(KEYINPUT29), .ZN(new_n825_) );
  INV_X1 g0689 ( .A(KEYINPUT29), .ZN(new_n826_) );
  NAND3_X1 g0690 ( .A1(new_n821_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_) );
  NAND2_X1 g0691 ( .A1(new_n825_), .A2(new_n827_), .ZN(new_n828_) );
  INV_X1 g0692 ( .A(new_n828_), .ZN(new_n829_) );
  NAND2_X1 g0693 ( .A1(new_n356_), .A2(new_n528_), .ZN(new_n830_) );
  INV_X1 g0694 ( .A(new_n830_), .ZN(new_n831_) );
  NAND2_X1 g0695 ( .A1(new_n613_), .A2(new_n831_), .ZN(new_n832_) );
  NAND2_X1 g0696 ( .A1(new_n832_), .A2(new_n353_), .ZN(new_n833_) );
  NAND3_X1 g0697 ( .A1(new_n833_), .A2(new_n631_), .A3(new_n829_), .ZN(new_n834_) );
  NAND2_X1 g0698 ( .A1(new_n822_), .A2(new_n631_), .ZN(new_n835_) );
  NAND2_X1 g0699 ( .A1(new_n834_), .A2(new_n835_), .ZN(new_n836_) );
  INV_X1 g0700 ( .A(new_n617_), .ZN(new_n837_) );
  NAND2_X1 g0701 ( .A1(new_n274_), .A2(new_n837_), .ZN(new_n838_) );
  NAND2_X1 g0702 ( .A1(new_n324_), .A2(new_n838_), .ZN(new_n839_) );
  NAND2_X1 g0703 ( .A1(new_n839_), .A2(new_n316_), .ZN(new_n840_) );
  NAND2_X1 g0704 ( .A1(new_n840_), .A2(new_n819_), .ZN(new_n841_) );
  INV_X1 g0705 ( .A(new_n841_), .ZN(new_n842_) );
  NAND2_X1 g0706 ( .A1(new_n836_), .A2(new_n842_), .ZN(new_n843_) );
  NAND4_X1 g0707 ( .A1(new_n432_), .A2(new_n613_), .A3(new_n528_), .A4(new_n631_), .ZN(new_n844_) );
  NAND2_X1 g0708 ( .A1(new_n844_), .A2(new_n606_), .ZN(new_n845_) );
  NAND3_X1 g0709 ( .A1(new_n843_), .A2(new_n819_), .A3(new_n845_), .ZN(new_n846_) );
  NAND2_X1 g0710 ( .A1(new_n843_), .A2(new_n819_), .ZN(new_n847_) );
  NAND3_X1 g0711 ( .A1(new_n847_), .A2(new_n606_), .A3(new_n844_), .ZN(new_n848_) );
  NAND2_X1 g0712 ( .A1(new_n848_), .A2(new_n846_), .ZN(new_n849_) );
  INV_X1 g0713 ( .A(new_n649_), .ZN(new_n850_) );
  NOR2_X1 g0714 ( .A1(new_n828_), .A2(new_n766_), .ZN(new_n851_) );
  NAND2_X1 g0715 ( .A1(new_n842_), .A2(new_n851_), .ZN(new_n852_) );
  NAND2_X1 g0716 ( .A1(new_n852_), .A2(new_n432_), .ZN(new_n853_) );
  INV_X1 g0717 ( .A(new_n852_), .ZN(new_n854_) );
  NAND2_X1 g0718 ( .A1(new_n854_), .A2(new_n433_), .ZN(new_n855_) );
  NAND2_X1 g0719 ( .A1(new_n855_), .A2(new_n853_), .ZN(new_n856_) );
  NAND2_X1 g0720 ( .A1(new_n856_), .A2(new_n850_), .ZN(new_n857_) );
  NAND2_X1 g0721 ( .A1(new_n849_), .A2(new_n857_), .ZN(new_n858_) );
  NAND4_X1 g0722 ( .A1(new_n848_), .A2(new_n850_), .A3(new_n846_), .A4(new_n856_), .ZN(new_n859_) );
  NAND2_X1 g0723 ( .A1(new_n858_), .A2(new_n859_), .ZN(new_n860_) );
  NAND2_X1 g0724 ( .A1(new_n860_), .A2(new_n178_), .ZN(new_n861_) );
  INV_X1 g0725 ( .A(G13), .ZN(new_n862_) );
  NAND2_X1 g0726 ( .A1(new_n862_), .A2(G1), .ZN(new_n863_) );
  NAND2_X1 g0727 ( .A1(new_n861_), .A2(new_n863_), .ZN(new_n864_) );
  NAND3_X1 g0728 ( .A1(G50), .A2(G58), .A3(G68), .ZN(new_n865_) );
  NAND2_X1 g0729 ( .A1(new_n140_), .A2(G50), .ZN(new_n866_) );
  NAND2_X1 g0730 ( .A1(G50), .A2(G58), .ZN(new_n867_) );
  NAND2_X1 g0731 ( .A1(new_n867_), .A2(new_n359_), .ZN(new_n868_) );
  NAND3_X1 g0732 ( .A1(new_n868_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n869_) );
  NAND3_X1 g0733 ( .A1(new_n869_), .A2(G1), .A3(new_n862_), .ZN(new_n870_) );
  NAND2_X1 g0734 ( .A1(new_n864_), .A2(new_n870_), .ZN(new_n871_) );
  NAND3_X1 g0735 ( .A1(new_n179_), .A2(G116), .A3(new_n214_), .ZN(new_n872_) );
  NAND2_X1 g0736 ( .A1(new_n871_), .A2(new_n872_), .ZN(G367) );
  INV_X1 g0737 ( .A(KEYINPUT55), .ZN(new_n874_) );
  NAND2_X1 g0738 ( .A1(new_n561_), .A2(new_n618_), .ZN(new_n875_) );
  NAND2_X1 g0739 ( .A1(new_n632_), .A2(new_n875_), .ZN(new_n876_) );
  NAND2_X1 g0740 ( .A1(new_n876_), .A2(new_n565_), .ZN(new_n877_) );
  NAND3_X1 g0741 ( .A1(new_n632_), .A2(new_n566_), .A3(new_n875_), .ZN(new_n878_) );
  NAND2_X1 g0742 ( .A1(new_n877_), .A2(new_n878_), .ZN(new_n879_) );
  NAND2_X1 g0743 ( .A1(new_n879_), .A2(new_n630_), .ZN(new_n880_) );
  NAND3_X1 g0744 ( .A1(new_n877_), .A2(new_n629_), .A3(new_n878_), .ZN(new_n881_) );
  NAND2_X1 g0745 ( .A1(new_n880_), .A2(new_n881_), .ZN(new_n882_) );
  NAND2_X1 g0746 ( .A1(new_n607_), .A2(new_n631_), .ZN(new_n883_) );
  NAND3_X1 g0747 ( .A1(new_n488_), .A2(new_n619_), .A3(new_n883_), .ZN(new_n884_) );
  NAND2_X1 g0748 ( .A1(new_n883_), .A2(new_n619_), .ZN(new_n885_) );
  NAND2_X1 g0749 ( .A1(new_n489_), .A2(new_n885_), .ZN(new_n886_) );
  NAND2_X1 g0750 ( .A1(new_n886_), .A2(new_n884_), .ZN(new_n887_) );
  NAND2_X1 g0751 ( .A1(new_n887_), .A2(new_n628_), .ZN(new_n888_) );
  NAND4_X1 g0752 ( .A1(new_n886_), .A2(G330), .A3(new_n627_), .A4(new_n884_), .ZN(new_n889_) );
  NAND2_X1 g0753 ( .A1(new_n888_), .A2(new_n889_), .ZN(new_n890_) );
  NAND2_X1 g0754 ( .A1(new_n882_), .A2(new_n890_), .ZN(new_n891_) );
  NAND2_X1 g0755 ( .A1(new_n891_), .A2(KEYINPUT52), .ZN(new_n892_) );
  INV_X1 g0756 ( .A(KEYINPUT52), .ZN(new_n893_) );
  NAND3_X1 g0757 ( .A1(new_n882_), .A2(new_n893_), .A3(new_n890_), .ZN(new_n894_) );
  NAND2_X1 g0758 ( .A1(new_n892_), .A2(new_n894_), .ZN(new_n895_) );
  NAND2_X1 g0759 ( .A1(new_n756_), .A2(new_n730_), .ZN(new_n896_) );
  INV_X1 g0760 ( .A(new_n896_), .ZN(new_n897_) );
  NAND2_X1 g0761 ( .A1(new_n895_), .A2(new_n897_), .ZN(new_n898_) );
  INV_X1 g0762 ( .A(KEYINPUT53), .ZN(new_n899_) );
  NAND2_X1 g0763 ( .A1(new_n613_), .A2(new_n631_), .ZN(new_n900_) );
  NAND2_X1 g0764 ( .A1(new_n900_), .A2(new_n528_), .ZN(new_n901_) );
  NAND2_X1 g0765 ( .A1(new_n610_), .A2(new_n564_), .ZN(new_n902_) );
  NAND3_X1 g0766 ( .A1(new_n902_), .A2(new_n529_), .A3(new_n631_), .ZN(new_n903_) );
  NAND3_X1 g0767 ( .A1(new_n901_), .A2(new_n899_), .A3(new_n903_), .ZN(new_n904_) );
  NAND4_X1 g0768 ( .A1(new_n506_), .A2(new_n522_), .A3(new_n523_), .A4(new_n618_), .ZN(new_n905_) );
  NAND2_X1 g0769 ( .A1(new_n901_), .A2(new_n903_), .ZN(new_n906_) );
  NAND2_X1 g0770 ( .A1(new_n906_), .A2(KEYINPUT53), .ZN(new_n907_) );
  NAND3_X1 g0771 ( .A1(new_n907_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n908_) );
  NAND2_X1 g0772 ( .A1(new_n566_), .A2(new_n875_), .ZN(new_n909_) );
  NAND4_X1 g0773 ( .A1(new_n562_), .A2(new_n561_), .A3(new_n563_), .A4(new_n618_), .ZN(new_n910_) );
  NAND2_X1 g0774 ( .A1(new_n909_), .A2(new_n910_), .ZN(new_n911_) );
  NAND2_X1 g0775 ( .A1(new_n629_), .A2(new_n911_), .ZN(new_n912_) );
  NAND2_X1 g0776 ( .A1(new_n908_), .A2(new_n912_), .ZN(new_n913_) );
  INV_X1 g0777 ( .A(new_n913_), .ZN(new_n914_) );
  INV_X1 g0778 ( .A(new_n912_), .ZN(new_n915_) );
  NAND4_X1 g0779 ( .A1(new_n907_), .A2(new_n904_), .A3(new_n905_), .A4(new_n915_), .ZN(new_n916_) );
  NAND2_X1 g0780 ( .A1(new_n916_), .A2(new_n731_), .ZN(new_n917_) );
  NOR2_X1 g0781 ( .A1(new_n914_), .A2(new_n917_), .ZN(new_n918_) );
  NAND2_X1 g0782 ( .A1(new_n918_), .A2(new_n898_), .ZN(new_n919_) );
  NAND2_X1 g0783 ( .A1(new_n529_), .A2(new_n663_), .ZN(new_n920_) );
  NAND2_X1 g0784 ( .A1(new_n735_), .A2(G317), .ZN(new_n921_) );
  NAND2_X1 g0785 ( .A1(new_n701_), .A2(G294), .ZN(new_n922_) );
  NAND2_X1 g0786 ( .A1(new_n733_), .A2(G107), .ZN(new_n923_) );
  NAND2_X1 g0787 ( .A1(new_n690_), .A2(G283), .ZN(new_n924_) );
  NAND4_X1 g0788 ( .A1(new_n923_), .A2(new_n921_), .A3(new_n922_), .A4(new_n924_), .ZN(new_n925_) );
  INV_X1 g0789 ( .A(KEYINPUT54), .ZN(new_n926_) );
  NAND2_X1 g0790 ( .A1(new_n714_), .A2(G311), .ZN(new_n927_) );
  NAND2_X1 g0791 ( .A1(new_n927_), .A2(new_n926_), .ZN(new_n928_) );
  NAND2_X1 g0792 ( .A1(new_n716_), .A2(G116), .ZN(new_n929_) );
  NAND2_X1 g0793 ( .A1(new_n720_), .A2(G303), .ZN(new_n930_) );
  NOR2_X1 g0794 ( .A1(new_n927_), .A2(new_n926_), .ZN(new_n931_) );
  NOR2_X1 g0795 ( .A1(new_n711_), .A2(new_n493_), .ZN(new_n932_) );
  NOR2_X1 g0796 ( .A1(new_n931_), .A2(new_n932_), .ZN(new_n933_) );
  NAND4_X1 g0797 ( .A1(new_n933_), .A2(new_n928_), .A3(new_n929_), .A4(new_n930_), .ZN(new_n934_) );
  NOR3_X1 g0798 ( .A1(new_n925_), .A2(new_n738_), .A3(new_n934_), .ZN(new_n935_) );
  INV_X1 g0799 ( .A(new_n710_), .ZN(new_n936_) );
  NAND2_X1 g0800 ( .A1(new_n744_), .A2(G77), .ZN(new_n937_) );
  NOR2_X1 g0801 ( .A1(new_n702_), .A2(new_n256_), .ZN(new_n938_) );
  INV_X1 g0802 ( .A(G137), .ZN(new_n939_) );
  NOR2_X1 g0803 ( .A1(new_n694_), .A2(new_n939_), .ZN(new_n940_) );
  NOR2_X1 g0804 ( .A1(new_n938_), .A2(new_n940_), .ZN(new_n941_) );
  NOR2_X1 g0805 ( .A1(new_n717_), .A2(new_n261_), .ZN(new_n942_) );
  NAND2_X1 g0806 ( .A1(new_n714_), .A2(G143), .ZN(new_n943_) );
  NAND2_X1 g0807 ( .A1(new_n720_), .A2(G150), .ZN(new_n944_) );
  NAND2_X1 g0808 ( .A1(new_n944_), .A2(new_n943_), .ZN(new_n945_) );
  NOR2_X1 g0809 ( .A1(new_n691_), .A2(new_n139_), .ZN(new_n946_) );
  NOR2_X1 g0810 ( .A1(new_n699_), .A2(new_n359_), .ZN(new_n947_) );
  NOR4_X1 g0811 ( .A1(new_n947_), .A2(new_n945_), .A3(new_n942_), .A4(new_n946_), .ZN(new_n948_) );
  NAND4_X1 g0812 ( .A1(new_n948_), .A2(new_n936_), .A3(new_n937_), .A4(new_n941_), .ZN(new_n949_) );
  NAND2_X1 g0813 ( .A1(new_n672_), .A2(new_n206_), .ZN(new_n950_) );
  NAND2_X1 g0814 ( .A1(new_n653_), .A2(G87), .ZN(new_n951_) );
  NAND3_X1 g0815 ( .A1(new_n686_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_) );
  NAND3_X1 g0816 ( .A1(new_n949_), .A2(new_n732_), .A3(new_n952_), .ZN(new_n953_) );
  NOR2_X1 g0817 ( .A1(new_n953_), .A2(new_n935_), .ZN(new_n954_) );
  NAND2_X1 g0818 ( .A1(new_n920_), .A2(new_n954_), .ZN(new_n955_) );
  NAND2_X1 g0819 ( .A1(new_n919_), .A2(new_n955_), .ZN(new_n956_) );
  NAND2_X1 g0820 ( .A1(new_n956_), .A2(new_n874_), .ZN(new_n957_) );
  NAND3_X1 g0821 ( .A1(new_n919_), .A2(KEYINPUT55), .A3(new_n955_), .ZN(new_n958_) );
  NAND2_X1 g0822 ( .A1(new_n957_), .A2(new_n958_), .ZN(G387) );
  NAND3_X1 g0823 ( .A1(new_n896_), .A2(new_n731_), .A3(new_n890_), .ZN(new_n960_) );
  NAND2_X1 g0824 ( .A1(new_n623_), .A2(new_n663_), .ZN(new_n961_) );
  NAND2_X1 g0825 ( .A1(new_n208_), .A2(G45), .ZN(new_n962_) );
  INV_X1 g0826 ( .A(KEYINPUT23), .ZN(new_n963_) );
  NAND2_X1 g0827 ( .A1(G68), .A2(G77), .ZN(new_n964_) );
  NAND4_X1 g0828 ( .A1(new_n657_), .A2(new_n139_), .A3(G58), .A4(new_n964_), .ZN(new_n965_) );
  NAND2_X1 g0829 ( .A1(new_n965_), .A2(new_n292_), .ZN(new_n966_) );
  NAND2_X1 g0830 ( .A1(new_n966_), .A2(new_n963_), .ZN(new_n967_) );
  NAND3_X1 g0831 ( .A1(new_n965_), .A2(new_n292_), .A3(KEYINPUT23), .ZN(new_n968_) );
  NAND2_X1 g0832 ( .A1(new_n967_), .A2(new_n968_), .ZN(new_n969_) );
  NAND2_X1 g0833 ( .A1(new_n962_), .A2(new_n969_), .ZN(new_n970_) );
  NAND2_X1 g0834 ( .A1(new_n970_), .A2(new_n672_), .ZN(new_n971_) );
  NAND2_X1 g0835 ( .A1(new_n653_), .A2(new_n460_), .ZN(new_n972_) );
  INV_X1 g0836 ( .A(new_n657_), .ZN(new_n973_) );
  NAND2_X1 g0837 ( .A1(new_n973_), .A2(new_n661_), .ZN(new_n974_) );
  NAND3_X1 g0838 ( .A1(new_n971_), .A2(new_n972_), .A3(new_n974_), .ZN(new_n975_) );
  NAND2_X1 g0839 ( .A1(new_n975_), .A2(new_n686_), .ZN(new_n976_) );
  NAND2_X1 g0840 ( .A1(new_n744_), .A2(G116), .ZN(new_n977_) );
  NAND2_X1 g0841 ( .A1(new_n977_), .A2(KEYINPUT25), .ZN(new_n978_) );
  INV_X1 g0842 ( .A(KEYINPUT25), .ZN(new_n979_) );
  NAND3_X1 g0843 ( .A1(new_n744_), .A2(G116), .A3(new_n979_), .ZN(new_n980_) );
  NAND2_X1 g0844 ( .A1(new_n716_), .A2(G294), .ZN(new_n981_) );
  NAND2_X1 g0845 ( .A1(new_n714_), .A2(G322), .ZN(new_n982_) );
  NAND2_X1 g0846 ( .A1(new_n981_), .A2(new_n982_), .ZN(new_n983_) );
  NAND2_X1 g0847 ( .A1(new_n983_), .A2(KEYINPUT26), .ZN(new_n984_) );
  INV_X1 g0848 ( .A(KEYINPUT26), .ZN(new_n985_) );
  NAND3_X1 g0849 ( .A1(new_n981_), .A2(new_n985_), .A3(new_n982_), .ZN(new_n986_) );
  NAND4_X1 g0850 ( .A1(new_n978_), .A2(new_n984_), .A3(new_n980_), .A4(new_n986_), .ZN(new_n987_) );
  NAND2_X1 g0851 ( .A1(new_n701_), .A2(G311), .ZN(new_n988_) );
  NAND2_X1 g0852 ( .A1(new_n733_), .A2(G283), .ZN(new_n989_) );
  NAND2_X1 g0853 ( .A1(new_n735_), .A2(G326), .ZN(new_n990_) );
  NAND3_X1 g0854 ( .A1(new_n989_), .A2(new_n988_), .A3(new_n990_), .ZN(new_n991_) );
  INV_X1 g0855 ( .A(new_n738_), .ZN(new_n992_) );
  NAND2_X1 g0856 ( .A1(new_n690_), .A2(G303), .ZN(new_n993_) );
  NAND2_X1 g0857 ( .A1(new_n720_), .A2(G317), .ZN(new_n994_) );
  NAND3_X1 g0858 ( .A1(new_n992_), .A2(new_n993_), .A3(new_n994_), .ZN(new_n995_) );
  NOR3_X1 g0859 ( .A1(new_n995_), .A2(new_n991_), .A3(new_n987_), .ZN(new_n996_) );
  NAND2_X1 g0860 ( .A1(new_n735_), .A2(G150), .ZN(new_n997_) );
  NAND2_X1 g0861 ( .A1(new_n690_), .A2(G68), .ZN(new_n998_) );
  NAND2_X1 g0862 ( .A1(new_n733_), .A2(G87), .ZN(new_n999_) );
  NAND3_X1 g0863 ( .A1(new_n999_), .A2(new_n997_), .A3(new_n998_), .ZN(new_n1000_) );
  NOR2_X1 g0864 ( .A1(new_n717_), .A2(new_n140_), .ZN(new_n1001_) );
  INV_X1 g0865 ( .A(new_n1001_), .ZN(new_n1002_) );
  NAND2_X1 g0866 ( .A1(new_n714_), .A2(G159), .ZN(new_n1003_) );
  NAND2_X1 g0867 ( .A1(new_n720_), .A2(G50), .ZN(new_n1004_) );
  NOR2_X1 g0868 ( .A1(new_n702_), .A2(new_n261_), .ZN(new_n1005_) );
  NOR2_X1 g0869 ( .A1(new_n1005_), .A2(new_n932_), .ZN(new_n1006_) );
  NAND4_X1 g0870 ( .A1(new_n1006_), .A2(new_n1002_), .A3(new_n1003_), .A4(new_n1004_), .ZN(new_n1007_) );
  NOR3_X1 g0871 ( .A1(new_n1000_), .A2(new_n710_), .A3(new_n1007_), .ZN(new_n1008_) );
  NOR3_X1 g0872 ( .A1(new_n996_), .A2(new_n1008_), .A3(new_n731_), .ZN(new_n1009_) );
  NAND3_X1 g0873 ( .A1(new_n961_), .A2(new_n976_), .A3(new_n1009_), .ZN(new_n1010_) );
  NAND4_X1 g0874 ( .A1(new_n756_), .A2(new_n654_), .A3(new_n888_), .A4(new_n889_), .ZN(new_n1011_) );
  NAND2_X1 g0875 ( .A1(new_n1011_), .A2(new_n1010_), .ZN(new_n1012_) );
  INV_X1 g0876 ( .A(new_n1012_), .ZN(new_n1013_) );
  NAND2_X1 g0877 ( .A1(new_n1013_), .A2(new_n960_), .ZN(G393) );
  NAND2_X1 g0878 ( .A1(new_n756_), .A2(new_n890_), .ZN(new_n1015_) );
  NAND3_X1 g0879 ( .A1(new_n1015_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n1016_) );
  NAND3_X1 g0880 ( .A1(new_n895_), .A2(new_n654_), .A3(new_n1016_), .ZN(new_n1017_) );
  NAND3_X1 g0881 ( .A1(new_n896_), .A2(new_n882_), .A3(new_n731_), .ZN(new_n1018_) );
  NAND3_X1 g0882 ( .A1(new_n909_), .A2(new_n663_), .A3(new_n910_), .ZN(new_n1019_) );
  INV_X1 g0883 ( .A(KEYINPUT58), .ZN(new_n1020_) );
  INV_X1 g0884 ( .A(new_n720_), .ZN(new_n1021_) );
  NOR2_X1 g0885 ( .A1(new_n1021_), .A2(new_n808_), .ZN(new_n1022_) );
  NAND2_X1 g0886 ( .A1(new_n690_), .A2(G294), .ZN(new_n1023_) );
  NAND2_X1 g0887 ( .A1(new_n701_), .A2(G303), .ZN(new_n1024_) );
  NAND2_X1 g0888 ( .A1(new_n733_), .A2(G116), .ZN(new_n1025_) );
  NAND2_X1 g0889 ( .A1(new_n735_), .A2(G322), .ZN(new_n1026_) );
  NAND4_X1 g0890 ( .A1(new_n1025_), .A2(new_n1023_), .A3(new_n1024_), .A4(new_n1026_), .ZN(new_n1027_) );
  NOR4_X1 g0891 ( .A1(new_n1027_), .A2(new_n258_), .A3(new_n712_), .A4(new_n1022_), .ZN(new_n1028_) );
  NAND2_X1 g0892 ( .A1(new_n1028_), .A2(new_n1020_), .ZN(new_n1029_) );
  NAND2_X1 g0893 ( .A1(new_n716_), .A2(G283), .ZN(new_n1030_) );
  NAND2_X1 g0894 ( .A1(new_n714_), .A2(G317), .ZN(new_n1031_) );
  NAND2_X1 g0895 ( .A1(new_n1030_), .A2(new_n1031_), .ZN(new_n1032_) );
  NAND2_X1 g0896 ( .A1(new_n1032_), .A2(KEYINPUT59), .ZN(new_n1033_) );
  INV_X1 g0897 ( .A(KEYINPUT59), .ZN(new_n1034_) );
  NAND3_X1 g0898 ( .A1(new_n1030_), .A2(new_n1034_), .A3(new_n1031_), .ZN(new_n1035_) );
  NAND2_X1 g0899 ( .A1(new_n1033_), .A2(new_n1035_), .ZN(new_n1036_) );
  INV_X1 g0900 ( .A(new_n1028_), .ZN(new_n1037_) );
  NAND2_X1 g0901 ( .A1(new_n1037_), .A2(KEYINPUT58), .ZN(new_n1038_) );
  NAND3_X1 g0902 ( .A1(new_n1038_), .A2(new_n1029_), .A3(new_n1036_), .ZN(new_n1039_) );
  NAND2_X1 g0903 ( .A1(new_n714_), .A2(G150), .ZN(new_n1040_) );
  NAND2_X1 g0904 ( .A1(new_n1040_), .A2(KEYINPUT56), .ZN(new_n1041_) );
  INV_X1 g0905 ( .A(KEYINPUT56), .ZN(new_n1042_) );
  NAND3_X1 g0906 ( .A1(new_n714_), .A2(G150), .A3(new_n1042_), .ZN(new_n1043_) );
  NAND2_X1 g0907 ( .A1(new_n1041_), .A2(new_n1043_), .ZN(new_n1044_) );
  NAND2_X1 g0908 ( .A1(new_n716_), .A2(G68), .ZN(new_n1045_) );
  NAND2_X1 g0909 ( .A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1046_) );
  NAND2_X1 g0910 ( .A1(new_n1046_), .A2(KEYINPUT57), .ZN(new_n1047_) );
  INV_X1 g0911 ( .A(KEYINPUT57), .ZN(new_n1048_) );
  NAND3_X1 g0912 ( .A1(new_n1044_), .A2(new_n1048_), .A3(new_n1045_), .ZN(new_n1049_) );
  NAND2_X1 g0913 ( .A1(new_n1047_), .A2(new_n1049_), .ZN(new_n1050_) );
  NOR2_X1 g0914 ( .A1(new_n691_), .A2(new_n261_), .ZN(new_n1051_) );
  NOR2_X1 g0915 ( .A1(new_n1021_), .A2(new_n256_), .ZN(new_n1052_) );
  NAND2_X1 g0916 ( .A1(new_n735_), .A2(G143), .ZN(new_n1053_) );
  NAND2_X1 g0917 ( .A1(new_n701_), .A2(G50), .ZN(new_n1054_) );
  NAND2_X1 g0918 ( .A1(new_n733_), .A2(G77), .ZN(new_n1055_) );
  NAND3_X1 g0919 ( .A1(new_n1055_), .A2(new_n1053_), .A3(new_n1054_), .ZN(new_n1056_) );
  NOR4_X1 g0920 ( .A1(new_n1056_), .A2(G33), .A3(new_n1051_), .A4(new_n1052_), .ZN(new_n1057_) );
  NAND3_X1 g0921 ( .A1(new_n1057_), .A2(new_n805_), .A3(new_n1050_), .ZN(new_n1058_) );
  NAND2_X1 g0922 ( .A1(new_n1039_), .A2(new_n1058_), .ZN(new_n1059_) );
  NAND2_X1 g0923 ( .A1(new_n1059_), .A2(new_n709_), .ZN(new_n1060_) );
  NAND2_X1 g0924 ( .A1(new_n226_), .A2(new_n672_), .ZN(new_n1061_) );
  NAND2_X1 g0925 ( .A1(new_n653_), .A2(G97), .ZN(new_n1062_) );
  NAND3_X1 g0926 ( .A1(new_n1061_), .A2(new_n686_), .A3(new_n1062_), .ZN(new_n1063_) );
  NAND4_X1 g0927 ( .A1(new_n1019_), .A2(new_n732_), .A3(new_n1060_), .A4(new_n1063_), .ZN(new_n1064_) );
  NAND2_X1 g0928 ( .A1(new_n1018_), .A2(new_n1064_), .ZN(new_n1065_) );
  INV_X1 g0929 ( .A(new_n1065_), .ZN(new_n1066_) );
  NAND2_X1 g0930 ( .A1(new_n1017_), .A2(new_n1066_), .ZN(G390) );
  INV_X1 g0931 ( .A(KEYINPUT38), .ZN(new_n1068_) );
  NAND3_X1 g0932 ( .A1(new_n432_), .A2(new_n648_), .A3(G330), .ZN(new_n1069_) );
  NAND3_X1 g0933 ( .A1(new_n844_), .A2(new_n606_), .A3(new_n1069_), .ZN(new_n1070_) );
  NAND2_X1 g0934 ( .A1(new_n1070_), .A2(new_n1068_), .ZN(new_n1071_) );
  NAND4_X1 g0935 ( .A1(new_n844_), .A2(new_n1069_), .A3(new_n606_), .A4(KEYINPUT38), .ZN(new_n1072_) );
  NAND2_X1 g0936 ( .A1(new_n1071_), .A2(new_n1072_), .ZN(new_n1073_) );
  NAND2_X1 g0937 ( .A1(new_n833_), .A2(new_n631_), .ZN(new_n1074_) );
  NAND2_X1 g0938 ( .A1(new_n850_), .A2(new_n764_), .ZN(new_n1075_) );
  NAND2_X1 g0939 ( .A1(new_n1074_), .A2(new_n1075_), .ZN(new_n1076_) );
  NAND2_X1 g0940 ( .A1(new_n1076_), .A2(new_n829_), .ZN(new_n1077_) );
  NAND3_X1 g0941 ( .A1(new_n1074_), .A2(new_n828_), .A3(new_n1075_), .ZN(new_n1078_) );
  NAND2_X1 g0942 ( .A1(new_n1077_), .A2(new_n1078_), .ZN(new_n1079_) );
  INV_X1 g0943 ( .A(new_n1079_), .ZN(new_n1080_) );
  NAND2_X1 g0944 ( .A1(new_n842_), .A2(KEYINPUT40), .ZN(new_n1081_) );
  INV_X1 g0945 ( .A(KEYINPUT40), .ZN(new_n1082_) );
  NAND2_X1 g0946 ( .A1(new_n841_), .A2(new_n1082_), .ZN(new_n1083_) );
  NAND2_X1 g0947 ( .A1(new_n1081_), .A2(new_n1083_), .ZN(new_n1084_) );
  INV_X1 g0948 ( .A(new_n1084_), .ZN(new_n1085_) );
  INV_X1 g0949 ( .A(KEYINPUT39), .ZN(new_n1086_) );
  NAND3_X1 g0950 ( .A1(new_n648_), .A2(G330), .A3(new_n851_), .ZN(new_n1087_) );
  NAND2_X1 g0951 ( .A1(new_n1087_), .A2(new_n1086_), .ZN(new_n1088_) );
  NAND4_X1 g0952 ( .A1(new_n648_), .A2(new_n851_), .A3(G330), .A4(KEYINPUT39), .ZN(new_n1089_) );
  NAND2_X1 g0953 ( .A1(new_n1088_), .A2(new_n1089_), .ZN(new_n1090_) );
  NAND3_X1 g0954 ( .A1(new_n834_), .A2(new_n1090_), .A3(new_n835_), .ZN(new_n1091_) );
  NAND2_X1 g0955 ( .A1(new_n1091_), .A2(new_n1085_), .ZN(new_n1092_) );
  NAND4_X1 g0956 ( .A1(new_n834_), .A2(new_n1090_), .A3(new_n835_), .A4(new_n1084_), .ZN(new_n1093_) );
  NAND2_X1 g0957 ( .A1(new_n1092_), .A2(new_n1093_), .ZN(new_n1094_) );
  NAND3_X1 g0958 ( .A1(new_n1080_), .A2(new_n1094_), .A3(new_n1073_), .ZN(new_n1095_) );
  NAND3_X1 g0959 ( .A1(new_n1077_), .A2(new_n1073_), .A3(new_n1078_), .ZN(new_n1096_) );
  NAND3_X1 g0960 ( .A1(new_n1096_), .A2(new_n1092_), .A3(new_n1093_), .ZN(new_n1097_) );
  NAND3_X1 g0961 ( .A1(new_n1095_), .A2(new_n654_), .A3(new_n1097_), .ZN(new_n1098_) );
  INV_X1 g0962 ( .A(new_n730_), .ZN(new_n1099_) );
  NAND2_X1 g0963 ( .A1(new_n1094_), .A2(new_n1099_), .ZN(new_n1100_) );
  NAND2_X1 g0964 ( .A1(new_n841_), .A2(new_n661_), .ZN(new_n1101_) );
  NAND2_X1 g0965 ( .A1(new_n733_), .A2(G159), .ZN(new_n1102_) );
  NAND2_X1 g0966 ( .A1(new_n690_), .A2(G143), .ZN(new_n1103_) );
  NAND2_X1 g0967 ( .A1(new_n744_), .A2(G50), .ZN(new_n1104_) );
  NAND2_X1 g0968 ( .A1(new_n716_), .A2(G150), .ZN(new_n1105_) );
  NAND2_X1 g0969 ( .A1(new_n714_), .A2(G128), .ZN(new_n1106_) );
  NAND2_X1 g0970 ( .A1(new_n720_), .A2(G132), .ZN(new_n1107_) );
  NAND3_X1 g0971 ( .A1(new_n1107_), .A2(new_n1105_), .A3(new_n1106_), .ZN(new_n1108_) );
  NAND2_X1 g0972 ( .A1(new_n701_), .A2(G137), .ZN(new_n1109_) );
  NAND2_X1 g0973 ( .A1(new_n735_), .A2(G125), .ZN(new_n1110_) );
  NAND2_X1 g0974 ( .A1(new_n1110_), .A2(new_n1109_), .ZN(new_n1111_) );
  NOR3_X1 g0975 ( .A1(new_n710_), .A2(new_n1108_), .A3(new_n1111_), .ZN(new_n1112_) );
  NAND4_X1 g0976 ( .A1(new_n1112_), .A2(new_n1102_), .A3(new_n1103_), .A4(new_n1104_), .ZN(new_n1113_) );
  INV_X1 g0977 ( .A(new_n714_), .ZN(new_n1114_) );
  NOR2_X1 g0978 ( .A1(new_n1114_), .A2(new_n806_), .ZN(new_n1115_) );
  NOR2_X1 g0979 ( .A1(new_n718_), .A2(new_n1115_), .ZN(new_n1116_) );
  NAND2_X1 g0980 ( .A1(new_n701_), .A2(G107), .ZN(new_n1117_) );
  NAND4_X1 g0981 ( .A1(new_n1055_), .A2(new_n781_), .A3(new_n1116_), .A4(new_n1117_), .ZN(new_n1118_) );
  INV_X1 g0982 ( .A(KEYINPUT47), .ZN(new_n1119_) );
  NAND2_X1 g0983 ( .A1(new_n720_), .A2(G116), .ZN(new_n1120_) );
  NAND2_X1 g0984 ( .A1(new_n1120_), .A2(new_n1119_), .ZN(new_n1121_) );
  NAND3_X1 g0985 ( .A1(new_n720_), .A2(G116), .A3(KEYINPUT47), .ZN(new_n1122_) );
  NAND2_X1 g0986 ( .A1(new_n1121_), .A2(new_n1122_), .ZN(new_n1123_) );
  NAND2_X1 g0987 ( .A1(new_n992_), .A2(new_n1123_), .ZN(new_n1124_) );
  NAND2_X1 g0988 ( .A1(new_n735_), .A2(G294), .ZN(new_n1125_) );
  NAND2_X1 g0989 ( .A1(new_n690_), .A2(G97), .ZN(new_n1126_) );
  NAND2_X1 g0990 ( .A1(new_n1125_), .A2(new_n1126_), .ZN(new_n1127_) );
  NAND2_X1 g0991 ( .A1(new_n1127_), .A2(KEYINPUT48), .ZN(new_n1128_) );
  INV_X1 g0992 ( .A(KEYINPUT48), .ZN(new_n1129_) );
  NAND3_X1 g0993 ( .A1(new_n1125_), .A2(new_n1129_), .A3(new_n1126_), .ZN(new_n1130_) );
  NAND2_X1 g0994 ( .A1(new_n1128_), .A2(new_n1130_), .ZN(new_n1131_) );
  NOR3_X1 g0995 ( .A1(new_n1118_), .A2(new_n1124_), .A3(new_n1131_), .ZN(new_n1132_) );
  NAND2_X1 g0996 ( .A1(new_n813_), .A2(new_n261_), .ZN(new_n1133_) );
  INV_X1 g0997 ( .A(new_n1133_), .ZN(new_n1134_) );
  NOR3_X1 g0998 ( .A1(new_n1132_), .A2(new_n731_), .A3(new_n1134_), .ZN(new_n1135_) );
  NAND3_X1 g0999 ( .A1(new_n1101_), .A2(new_n1113_), .A3(new_n1135_), .ZN(new_n1136_) );
  NAND2_X1 g1000 ( .A1(new_n1100_), .A2(new_n1136_), .ZN(new_n1137_) );
  INV_X1 g1001 ( .A(new_n1137_), .ZN(new_n1138_) );
  NAND2_X1 g1002 ( .A1(new_n1138_), .A2(new_n1098_), .ZN(G378) );
  INV_X1 g1003 ( .A(KEYINPUT41), .ZN(new_n1140_) );
  NAND2_X1 g1004 ( .A1(new_n1080_), .A2(new_n1094_), .ZN(new_n1141_) );
  NAND2_X1 g1005 ( .A1(new_n1141_), .A2(new_n1140_), .ZN(new_n1142_) );
  NAND3_X1 g1006 ( .A1(new_n1080_), .A2(new_n1094_), .A3(KEYINPUT41), .ZN(new_n1143_) );
  NAND2_X1 g1007 ( .A1(new_n1142_), .A2(new_n1143_), .ZN(new_n1144_) );
  NAND2_X1 g1008 ( .A1(new_n1073_), .A2(new_n730_), .ZN(new_n1145_) );
  INV_X1 g1009 ( .A(new_n1145_), .ZN(new_n1146_) );
  NAND2_X1 g1010 ( .A1(new_n1144_), .A2(new_n1146_), .ZN(new_n1147_) );
  NAND2_X1 g1011 ( .A1(new_n854_), .A2(new_n850_), .ZN(new_n1148_) );
  NAND3_X1 g1012 ( .A1(new_n843_), .A2(new_n819_), .A3(new_n1148_), .ZN(new_n1149_) );
  NAND2_X1 g1013 ( .A1(new_n406_), .A2(new_n837_), .ZN(new_n1150_) );
  NAND2_X1 g1014 ( .A1(new_n430_), .A2(new_n1150_), .ZN(new_n1151_) );
  NAND4_X1 g1015 ( .A1(new_n406_), .A2(new_n420_), .A3(new_n421_), .A4(new_n837_), .ZN(new_n1152_) );
  NAND2_X1 g1016 ( .A1(new_n1151_), .A2(new_n1152_), .ZN(new_n1153_) );
  INV_X1 g1017 ( .A(new_n1153_), .ZN(new_n1154_) );
  NAND2_X1 g1018 ( .A1(new_n1149_), .A2(new_n1154_), .ZN(new_n1155_) );
  NAND4_X1 g1019 ( .A1(new_n843_), .A2(new_n819_), .A3(new_n1148_), .A4(new_n1153_), .ZN(new_n1156_) );
  NAND2_X1 g1020 ( .A1(new_n1155_), .A2(new_n1156_), .ZN(new_n1157_) );
  NAND2_X1 g1021 ( .A1(new_n1157_), .A2(new_n731_), .ZN(new_n1158_) );
  INV_X1 g1022 ( .A(new_n1158_), .ZN(new_n1159_) );
  NAND2_X1 g1023 ( .A1(new_n1147_), .A2(new_n1159_), .ZN(new_n1160_) );
  NAND2_X1 g1024 ( .A1(new_n1154_), .A2(new_n661_), .ZN(new_n1161_) );
  INV_X1 g1025 ( .A(KEYINPUT44), .ZN(new_n1162_) );
  NAND2_X1 g1026 ( .A1(new_n744_), .A2(G159), .ZN(new_n1163_) );
  NAND2_X1 g1027 ( .A1(new_n701_), .A2(G132), .ZN(new_n1164_) );
  NAND2_X1 g1028 ( .A1(new_n1163_), .A2(new_n1164_), .ZN(new_n1165_) );
  NAND2_X1 g1029 ( .A1(new_n1165_), .A2(new_n1162_), .ZN(new_n1166_) );
  NAND3_X1 g1030 ( .A1(new_n1163_), .A2(KEYINPUT44), .A3(new_n1164_), .ZN(new_n1167_) );
  NAND2_X1 g1031 ( .A1(new_n1166_), .A2(new_n1167_), .ZN(new_n1168_) );
  NAND2_X1 g1032 ( .A1(new_n716_), .A2(G143), .ZN(new_n1169_) );
  NAND2_X1 g1033 ( .A1(new_n714_), .A2(G125), .ZN(new_n1170_) );
  NAND2_X1 g1034 ( .A1(new_n720_), .A2(G128), .ZN(new_n1171_) );
  NAND3_X1 g1035 ( .A1(new_n1171_), .A2(new_n1169_), .A3(new_n1170_), .ZN(new_n1172_) );
  NAND2_X1 g1036 ( .A1(new_n733_), .A2(G150), .ZN(new_n1173_) );
  NAND2_X1 g1037 ( .A1(new_n735_), .A2(G124), .ZN(new_n1174_) );
  NAND2_X1 g1038 ( .A1(new_n1173_), .A2(new_n1174_), .ZN(new_n1175_) );
  NOR3_X1 g1039 ( .A1(new_n691_), .A2(new_n939_), .A3(KEYINPUT43), .ZN(new_n1176_) );
  INV_X1 g1040 ( .A(KEYINPUT43), .ZN(new_n1177_) );
  NOR2_X1 g1041 ( .A1(new_n691_), .A2(new_n939_), .ZN(new_n1178_) );
  NOR2_X1 g1042 ( .A1(new_n1178_), .A2(new_n1177_), .ZN(new_n1179_) );
  NOR4_X1 g1043 ( .A1(new_n1175_), .A2(new_n1179_), .A3(new_n1172_), .A4(new_n1176_), .ZN(new_n1180_) );
  NAND2_X1 g1044 ( .A1(new_n1180_), .A2(new_n1168_), .ZN(new_n1181_) );
  NAND2_X1 g1045 ( .A1(new_n1181_), .A2(new_n258_), .ZN(new_n1182_) );
  NOR2_X1 g1046 ( .A1(new_n691_), .A2(new_n218_), .ZN(new_n1183_) );
  NOR2_X1 g1047 ( .A1(new_n711_), .A2(new_n261_), .ZN(new_n1184_) );
  NOR2_X1 g1048 ( .A1(new_n1021_), .A2(new_n460_), .ZN(new_n1185_) );
  NOR2_X1 g1049 ( .A1(new_n1185_), .A2(KEYINPUT42), .ZN(new_n1186_) );
  INV_X1 g1050 ( .A(KEYINPUT42), .ZN(new_n1187_) );
  NOR3_X1 g1051 ( .A1(new_n1021_), .A2(new_n460_), .A3(new_n1187_), .ZN(new_n1188_) );
  NOR4_X1 g1052 ( .A1(new_n1186_), .A2(new_n1188_), .A3(new_n1183_), .A4(new_n1184_), .ZN(new_n1189_) );
  NOR2_X1 g1053 ( .A1(new_n1114_), .A2(new_n220_), .ZN(new_n1190_) );
  NOR3_X1 g1054 ( .A1(new_n947_), .A2(new_n1001_), .A3(new_n1190_), .ZN(new_n1191_) );
  NAND2_X1 g1055 ( .A1(new_n701_), .A2(G97), .ZN(new_n1192_) );
  NAND2_X1 g1056 ( .A1(new_n735_), .A2(G283), .ZN(new_n1193_) );
  NAND4_X1 g1057 ( .A1(new_n1189_), .A2(new_n1191_), .A3(new_n1192_), .A4(new_n1193_), .ZN(new_n1194_) );
  NAND2_X1 g1058 ( .A1(new_n1194_), .A2(G33), .ZN(new_n1195_) );
  NAND4_X1 g1059 ( .A1(new_n1182_), .A2(new_n1195_), .A3(new_n291_), .A4(new_n709_), .ZN(new_n1196_) );
  NAND2_X1 g1060 ( .A1(new_n709_), .A2(new_n291_), .ZN(new_n1197_) );
  NAND3_X1 g1061 ( .A1(new_n1197_), .A2(new_n139_), .A3(new_n662_), .ZN(new_n1198_) );
  NAND4_X1 g1062 ( .A1(new_n1161_), .A2(new_n732_), .A3(new_n1196_), .A4(new_n1198_), .ZN(new_n1199_) );
  NAND2_X1 g1063 ( .A1(new_n1160_), .A2(new_n1199_), .ZN(G375) );
  INV_X1 g1064 ( .A(KEYINPUT46), .ZN(new_n1201_) );
  INV_X1 g1065 ( .A(new_n1073_), .ZN(new_n1202_) );
  NAND2_X1 g1066 ( .A1(new_n1079_), .A2(new_n1202_), .ZN(new_n1203_) );
  NAND2_X1 g1067 ( .A1(new_n1203_), .A2(new_n1096_), .ZN(new_n1204_) );
  NAND2_X1 g1068 ( .A1(new_n1204_), .A2(new_n1201_), .ZN(new_n1205_) );
  NAND3_X1 g1069 ( .A1(new_n1203_), .A2(KEYINPUT46), .A3(new_n1096_), .ZN(new_n1206_) );
  NAND2_X1 g1070 ( .A1(new_n1205_), .A2(new_n1206_), .ZN(new_n1207_) );
  NAND2_X1 g1071 ( .A1(new_n1207_), .A2(new_n654_), .ZN(new_n1208_) );
  NAND2_X1 g1072 ( .A1(new_n1080_), .A2(new_n1099_), .ZN(new_n1209_) );
  NAND2_X1 g1073 ( .A1(new_n828_), .A2(new_n661_), .ZN(new_n1210_) );
  INV_X1 g1074 ( .A(KEYINPUT45), .ZN(new_n1211_) );
  NAND2_X1 g1075 ( .A1(new_n733_), .A2(G50), .ZN(new_n1212_) );
  NAND2_X1 g1076 ( .A1(new_n735_), .A2(G128), .ZN(new_n1213_) );
  NAND2_X1 g1077 ( .A1(new_n701_), .A2(G143), .ZN(new_n1214_) );
  NAND2_X1 g1078 ( .A1(new_n716_), .A2(G159), .ZN(new_n1215_) );
  NAND2_X1 g1079 ( .A1(new_n714_), .A2(G132), .ZN(new_n1216_) );
  NAND2_X1 g1080 ( .A1(new_n720_), .A2(G137), .ZN(new_n1217_) );
  NAND3_X1 g1081 ( .A1(new_n1217_), .A2(new_n1215_), .A3(new_n1216_), .ZN(new_n1218_) );
  INV_X1 g1082 ( .A(G150), .ZN(new_n1219_) );
  NOR2_X1 g1083 ( .A1(new_n691_), .A2(new_n1219_), .ZN(new_n1220_) );
  NOR4_X1 g1084 ( .A1(new_n710_), .A2(new_n1218_), .A3(new_n1184_), .A4(new_n1220_), .ZN(new_n1221_) );
  NAND4_X1 g1085 ( .A1(new_n1221_), .A2(new_n1212_), .A3(new_n1213_), .A4(new_n1214_), .ZN(new_n1222_) );
  NAND2_X1 g1086 ( .A1(new_n690_), .A2(G107), .ZN(new_n1223_) );
  NAND2_X1 g1087 ( .A1(new_n701_), .A2(G116), .ZN(new_n1224_) );
  NAND2_X1 g1088 ( .A1(new_n735_), .A2(G303), .ZN(new_n1225_) );
  NOR2_X1 g1089 ( .A1(new_n1021_), .A2(new_n806_), .ZN(new_n1226_) );
  NAND2_X1 g1090 ( .A1(new_n716_), .A2(G97), .ZN(new_n1227_) );
  NAND2_X1 g1091 ( .A1(new_n714_), .A2(G294), .ZN(new_n1228_) );
  NAND2_X1 g1092 ( .A1(new_n1227_), .A2(new_n1228_), .ZN(new_n1229_) );
  NAND2_X1 g1093 ( .A1(new_n999_), .A2(new_n937_), .ZN(new_n1230_) );
  NOR4_X1 g1094 ( .A1(new_n1230_), .A2(new_n738_), .A3(new_n1226_), .A4(new_n1229_), .ZN(new_n1231_) );
  NAND4_X1 g1095 ( .A1(new_n1231_), .A2(new_n1223_), .A3(new_n1224_), .A4(new_n1225_), .ZN(new_n1232_) );
  NAND2_X1 g1096 ( .A1(new_n813_), .A2(new_n359_), .ZN(new_n1233_) );
  NAND4_X1 g1097 ( .A1(new_n1232_), .A2(new_n1222_), .A3(new_n732_), .A4(new_n1233_), .ZN(new_n1234_) );
  INV_X1 g1098 ( .A(new_n1234_), .ZN(new_n1235_) );
  NAND2_X1 g1099 ( .A1(new_n1235_), .A2(new_n1211_), .ZN(new_n1236_) );
  NAND2_X1 g1100 ( .A1(new_n1234_), .A2(KEYINPUT45), .ZN(new_n1237_) );
  NAND2_X1 g1101 ( .A1(new_n1236_), .A2(new_n1237_), .ZN(new_n1238_) );
  NAND2_X1 g1102 ( .A1(new_n1210_), .A2(new_n1238_), .ZN(new_n1239_) );
  NAND2_X1 g1103 ( .A1(new_n1209_), .A2(new_n1239_), .ZN(new_n1240_) );
  INV_X1 g1104 ( .A(new_n1240_), .ZN(new_n1241_) );
  NAND2_X1 g1105 ( .A1(new_n1208_), .A2(new_n1241_), .ZN(G381) );
  INV_X1 g1106 ( .A(G378), .ZN(new_n1243_) );
  NAND3_X1 g1107 ( .A1(new_n1160_), .A2(new_n1243_), .A3(new_n1199_), .ZN(new_n1244_) );
  INV_X1 g1108 ( .A(new_n1244_), .ZN(new_n1245_) );
  INV_X1 g1109 ( .A(G396), .ZN(new_n1246_) );
  NAND3_X1 g1110 ( .A1(new_n1017_), .A2(new_n1246_), .A3(new_n1066_), .ZN(new_n1247_) );
  NAND4_X1 g1111 ( .A1(new_n1013_), .A2(new_n769_), .A3(new_n817_), .A4(new_n960_), .ZN(new_n1248_) );
  NOR4_X1 g1112 ( .A1(G387), .A2(G381), .A3(new_n1247_), .A4(new_n1248_), .ZN(new_n1249_) );
  NAND2_X1 g1113 ( .A1(new_n1249_), .A2(new_n1245_), .ZN(G407) );
  NAND2_X1 g1114 ( .A1(new_n1245_), .A2(new_n616_), .ZN(new_n1251_) );
  NAND3_X1 g1115 ( .A1(G407), .A2(new_n1251_), .A3(G213), .ZN(G409) );
  NAND2_X1 g1116 ( .A1(G390), .A2(G396), .ZN(new_n1253_) );
  NAND2_X1 g1117 ( .A1(new_n1253_), .A2(new_n1247_), .ZN(new_n1254_) );
  NAND2_X1 g1118 ( .A1(G381), .A2(new_n1254_), .ZN(new_n1255_) );
  NAND4_X1 g1119 ( .A1(new_n1208_), .A2(new_n1241_), .A3(new_n1247_), .A4(new_n1253_), .ZN(new_n1256_) );
  NAND2_X1 g1120 ( .A1(new_n1255_), .A2(new_n1256_), .ZN(new_n1257_) );
  NAND2_X1 g1121 ( .A1(G393), .A2(G384), .ZN(new_n1258_) );
  NAND2_X1 g1122 ( .A1(new_n1258_), .A2(new_n1248_), .ZN(new_n1259_) );
  NAND2_X1 g1123 ( .A1(G387), .A2(new_n1259_), .ZN(new_n1260_) );
  NAND4_X1 g1124 ( .A1(new_n957_), .A2(new_n958_), .A3(new_n1248_), .A4(new_n1258_), .ZN(new_n1261_) );
  NAND2_X1 g1125 ( .A1(new_n1260_), .A2(new_n1261_), .ZN(new_n1262_) );
  NAND2_X1 g1126 ( .A1(new_n1262_), .A2(new_n1257_), .ZN(new_n1263_) );
  NAND4_X1 g1127 ( .A1(new_n1260_), .A2(new_n1255_), .A3(new_n1256_), .A4(new_n1261_), .ZN(new_n1264_) );
  NAND2_X1 g1128 ( .A1(new_n1263_), .A2(new_n1264_), .ZN(new_n1265_) );
  NAND2_X1 g1129 ( .A1(new_n616_), .A2(G213), .ZN(new_n1266_) );
  NAND2_X1 g1130 ( .A1(G375), .A2(G378), .ZN(new_n1267_) );
  NAND3_X1 g1131 ( .A1(new_n1267_), .A2(new_n1244_), .A3(new_n1266_), .ZN(new_n1268_) );
  INV_X1 g1132 ( .A(KEYINPUT63), .ZN(new_n1269_) );
  NAND3_X1 g1133 ( .A1(new_n616_), .A2(G213), .A3(G2897), .ZN(new_n1270_) );
  NAND2_X1 g1134 ( .A1(new_n1270_), .A2(new_n1269_), .ZN(new_n1271_) );
  NAND4_X1 g1135 ( .A1(new_n616_), .A2(G213), .A3(G2897), .A4(KEYINPUT63), .ZN(new_n1272_) );
  NAND2_X1 g1136 ( .A1(new_n1271_), .A2(new_n1272_), .ZN(new_n1273_) );
  NAND3_X1 g1137 ( .A1(new_n1265_), .A2(new_n1268_), .A3(new_n1273_), .ZN(new_n1274_) );
  NAND2_X1 g1138 ( .A1(new_n1268_), .A2(new_n1273_), .ZN(new_n1275_) );
  NAND3_X1 g1139 ( .A1(new_n1275_), .A2(new_n1263_), .A3(new_n1264_), .ZN(new_n1276_) );
  NAND2_X1 g1140 ( .A1(new_n1274_), .A2(new_n1276_), .ZN(G405) );
  NAND2_X1 g1141 ( .A1(new_n1267_), .A2(new_n1244_), .ZN(new_n1278_) );
  NAND2_X1 g1142 ( .A1(new_n1265_), .A2(new_n1278_), .ZN(new_n1279_) );
  NAND4_X1 g1143 ( .A1(new_n1263_), .A2(new_n1244_), .A3(new_n1264_), .A4(new_n1267_), .ZN(new_n1280_) );
  NAND2_X1 g1144 ( .A1(new_n1279_), .A2(new_n1280_), .ZN(G402) );
endmodule


