module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n373_, new_n376_, new_n378_, new_n379_, new_n381_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n390_, new_n391_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n483_, new_n484_, new_n486_, new_n487_, new_n488_, new_n490_, new_n491_, new_n492_, new_n493_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n511_, new_n512_, new_n513_, new_n514_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_;
  XNOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 g001 ( .A(G132), .ZN(G219) );
  INV_X1 g002 ( .A(G82), .ZN(G220) );
  INV_X1 g003 ( .A(G96), .ZN(G221) );
  INV_X1 g004 ( .A(G69), .ZN(G235) );
  INV_X1 g005 ( .A(G120), .ZN(G236) );
  INV_X1 g006 ( .A(G57), .ZN(G237) );
  INV_X1 g007 ( .A(G108), .ZN(G238) );
  INV_X1 g008 ( .A(G2072), .ZN(new_n367_) );
  AND2_X1 g009 ( .A1(G2078), .A2(G2084), .ZN(new_n368_) );
  XNOR2_X1 g010 ( .A(new_n368_), .B(KEYINPUT20), .ZN(new_n369_) );
  AND2_X1 g011 ( .A1(new_n369_), .A2(G2090), .ZN(new_n370_) );
  XNOR2_X1 g012 ( .A(new_n370_), .B(KEYINPUT21), .ZN(new_n371_) );
  OR2_X1 g013 ( .A1(new_n371_), .A2(new_n367_), .ZN(G158) );
  AND3_X1 g014 ( .A1(G2), .A2(G15), .A3(G661), .ZN(new_n373_) );
  INV_X1 g015 ( .A(new_n373_), .ZN(G259) );
  AND2_X1 g016 ( .A1(G94), .A2(G452), .ZN(G173) );
  AND2_X1 g017 ( .A1(G7), .A2(G661), .ZN(new_n376_) );
  XOR2_X1 g018 ( .A(new_n376_), .B(KEYINPUT10), .Z(G223) );
  INV_X1 g019 ( .A(G567), .ZN(new_n378_) );
  OR2_X1 g020 ( .A1(G223), .A2(new_n378_), .ZN(new_n379_) );
  XOR2_X1 g021 ( .A(new_n379_), .B(KEYINPUT11), .Z(G234) );
  INV_X1 g022 ( .A(G2106), .ZN(new_n381_) );
  OR2_X1 g023 ( .A1(G223), .A2(new_n381_), .ZN(G217) );
  INV_X1 g024 ( .A(G218), .ZN(new_n383_) );
  AND2_X1 g025 ( .A1(G82), .A2(G132), .ZN(new_n384_) );
  XNOR2_X1 g026 ( .A(new_n384_), .B(KEYINPUT22), .ZN(new_n385_) );
  AND3_X1 g027 ( .A1(new_n385_), .A2(G96), .A3(new_n383_), .ZN(new_n386_) );
  AND4_X1 g028 ( .A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n387_) );
  AND2_X1 g029 ( .A1(new_n386_), .A2(new_n387_), .ZN(G325) );
  INV_X1 g030 ( .A(G325), .ZN(G261) );
  OR2_X1 g031 ( .A1(new_n386_), .A2(new_n381_), .ZN(new_n390_) );
  OR2_X1 g032 ( .A1(new_n387_), .A2(new_n378_), .ZN(new_n391_) );
  AND2_X1 g033 ( .A1(new_n390_), .A2(new_n391_), .ZN(G319) );
  INV_X1 g034 ( .A(G137), .ZN(new_n393_) );
  INV_X1 g035 ( .A(KEYINPUT17), .ZN(new_n394_) );
  OR2_X1 g036 ( .A1(G2104), .A2(G2105), .ZN(new_n395_) );
  XNOR2_X1 g037 ( .A(new_n395_), .B(new_n394_), .ZN(new_n396_) );
  OR2_X1 g038 ( .A1(new_n396_), .A2(new_n393_), .ZN(new_n397_) );
  INV_X1 g039 ( .A(G2105), .ZN(new_n398_) );
  AND3_X1 g040 ( .A1(new_n398_), .A2(G101), .A3(G2104), .ZN(new_n399_) );
  XNOR2_X1 g041 ( .A(new_n399_), .B(KEYINPUT23), .ZN(new_n400_) );
  INV_X1 g042 ( .A(G125), .ZN(new_n401_) );
  OR2_X1 g043 ( .A1(new_n401_), .A2(G2104), .ZN(new_n402_) );
  AND2_X1 g044 ( .A1(G113), .A2(G2104), .ZN(new_n403_) );
  INV_X1 g045 ( .A(new_n403_), .ZN(new_n404_) );
  AND2_X1 g046 ( .A1(new_n402_), .A2(new_n404_), .ZN(new_n405_) );
  OR2_X1 g047 ( .A1(new_n405_), .A2(new_n398_), .ZN(new_n406_) );
  AND3_X1 g048 ( .A1(new_n397_), .A2(new_n400_), .A3(new_n406_), .ZN(G160) );
  XNOR2_X1 g049 ( .A(new_n395_), .B(KEYINPUT17), .ZN(new_n408_) );
  AND2_X1 g050 ( .A1(new_n408_), .A2(G136), .ZN(new_n409_) );
  INV_X1 g051 ( .A(G2104), .ZN(new_n410_) );
  AND2_X1 g052 ( .A1(new_n410_), .A2(G2105), .ZN(new_n411_) );
  AND2_X1 g053 ( .A1(new_n411_), .A2(G124), .ZN(new_n412_) );
  XNOR2_X1 g054 ( .A(new_n412_), .B(KEYINPUT44), .ZN(new_n413_) );
  AND2_X1 g055 ( .A1(G2104), .A2(G2105), .ZN(new_n414_) );
  AND2_X1 g056 ( .A1(new_n414_), .A2(G112), .ZN(new_n415_) );
  AND2_X1 g057 ( .A1(new_n398_), .A2(G2104), .ZN(new_n416_) );
  AND2_X1 g058 ( .A1(new_n416_), .A2(G100), .ZN(new_n417_) );
  OR4_X1 g059 ( .A1(new_n413_), .A2(new_n409_), .A3(new_n415_), .A4(new_n417_), .ZN(new_n418_) );
  INV_X1 g060 ( .A(new_n418_), .ZN(G162) );
  AND2_X1 g061 ( .A1(new_n408_), .A2(G138), .ZN(new_n420_) );
  AND3_X1 g062 ( .A1(new_n398_), .A2(G102), .A3(G2104), .ZN(new_n421_) );
  AND3_X1 g063 ( .A1(new_n410_), .A2(G126), .A3(G2105), .ZN(new_n422_) );
  AND2_X1 g064 ( .A1(new_n414_), .A2(G114), .ZN(new_n423_) );
  OR3_X1 g065 ( .A1(new_n423_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n424_) );
  OR2_X1 g066 ( .A1(new_n420_), .A2(new_n424_), .ZN(new_n425_) );
  INV_X1 g067 ( .A(new_n425_), .ZN(G164) );
  INV_X1 g068 ( .A(G543), .ZN(new_n427_) );
  AND2_X1 g069 ( .A1(new_n427_), .A2(G651), .ZN(new_n428_) );
  XNOR2_X1 g070 ( .A(new_n428_), .B(KEYINPUT1), .ZN(new_n429_) );
  INV_X1 g071 ( .A(new_n429_), .ZN(new_n430_) );
  AND2_X1 g072 ( .A1(new_n430_), .A2(G62), .ZN(new_n431_) );
  INV_X1 g073 ( .A(G651), .ZN(new_n432_) );
  AND2_X1 g074 ( .A1(new_n427_), .A2(new_n432_), .ZN(new_n433_) );
  AND2_X1 g075 ( .A1(new_n433_), .A2(G88), .ZN(new_n434_) );
  XNOR2_X1 g076 ( .A(G543), .B(KEYINPUT0), .ZN(new_n435_) );
  AND2_X1 g077 ( .A1(new_n435_), .A2(G651), .ZN(new_n436_) );
  AND2_X1 g078 ( .A1(new_n436_), .A2(G75), .ZN(new_n437_) );
  AND2_X1 g079 ( .A1(new_n435_), .A2(new_n432_), .ZN(new_n438_) );
  AND2_X1 g080 ( .A1(new_n438_), .A2(G50), .ZN(new_n439_) );
  OR4_X1 g081 ( .A1(new_n431_), .A2(new_n434_), .A3(new_n437_), .A4(new_n439_), .ZN(G303) );
  INV_X1 g082 ( .A(G303), .ZN(G166) );
  AND2_X1 g083 ( .A1(new_n430_), .A2(G63), .ZN(new_n442_) );
  AND2_X1 g084 ( .A1(new_n438_), .A2(G51), .ZN(new_n443_) );
  OR2_X1 g085 ( .A1(new_n442_), .A2(new_n443_), .ZN(new_n444_) );
  XOR2_X1 g086 ( .A(new_n444_), .B(KEYINPUT6), .Z(new_n445_) );
  AND2_X1 g087 ( .A1(new_n433_), .A2(G89), .ZN(new_n446_) );
  XNOR2_X1 g088 ( .A(new_n446_), .B(KEYINPUT4), .ZN(new_n447_) );
  AND2_X1 g089 ( .A1(new_n436_), .A2(G76), .ZN(new_n448_) );
  OR2_X1 g090 ( .A1(new_n447_), .A2(new_n448_), .ZN(new_n449_) );
  XNOR2_X1 g091 ( .A(new_n449_), .B(KEYINPUT5), .ZN(new_n450_) );
  AND2_X1 g092 ( .A1(new_n445_), .A2(new_n450_), .ZN(new_n451_) );
  XNOR2_X1 g093 ( .A(new_n451_), .B(KEYINPUT7), .ZN(new_n452_) );
  INV_X1 g094 ( .A(new_n452_), .ZN(G168) );
  AND2_X1 g095 ( .A1(new_n436_), .A2(G77), .ZN(new_n454_) );
  AND2_X1 g096 ( .A1(new_n433_), .A2(G90), .ZN(new_n455_) );
  OR2_X1 g097 ( .A1(new_n454_), .A2(new_n455_), .ZN(new_n456_) );
  INV_X1 g098 ( .A(new_n456_), .ZN(new_n457_) );
  AND2_X1 g099 ( .A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n458_) );
  OR2_X1 g100 ( .A1(new_n457_), .A2(KEYINPUT9), .ZN(new_n459_) );
  INV_X1 g101 ( .A(new_n459_), .ZN(new_n460_) );
  AND2_X1 g102 ( .A1(new_n430_), .A2(G64), .ZN(new_n461_) );
  AND2_X1 g103 ( .A1(new_n438_), .A2(G52), .ZN(new_n462_) );
  OR4_X1 g104 ( .A1(new_n460_), .A2(new_n458_), .A3(new_n461_), .A4(new_n462_), .ZN(G301) );
  INV_X1 g105 ( .A(G301), .ZN(G171) );
  INV_X1 g106 ( .A(KEYINPUT14), .ZN(new_n465_) );
  AND2_X1 g107 ( .A1(new_n430_), .A2(G56), .ZN(new_n466_) );
  INV_X1 g108 ( .A(new_n466_), .ZN(new_n467_) );
  OR2_X1 g109 ( .A1(new_n467_), .A2(new_n465_), .ZN(new_n468_) );
  AND2_X1 g110 ( .A1(new_n438_), .A2(G43), .ZN(new_n469_) );
  INV_X1 g111 ( .A(new_n469_), .ZN(new_n470_) );
  OR2_X1 g112 ( .A1(new_n466_), .A2(KEYINPUT14), .ZN(new_n471_) );
  INV_X1 g113 ( .A(KEYINPUT13), .ZN(new_n472_) );
  INV_X1 g114 ( .A(KEYINPUT12), .ZN(new_n473_) );
  AND2_X1 g115 ( .A1(new_n433_), .A2(G81), .ZN(new_n474_) );
  XNOR2_X1 g116 ( .A(new_n474_), .B(new_n473_), .ZN(new_n475_) );
  AND3_X1 g117 ( .A1(new_n435_), .A2(G68), .A3(G651), .ZN(new_n476_) );
  INV_X1 g118 ( .A(new_n476_), .ZN(new_n477_) );
  AND2_X1 g119 ( .A1(new_n475_), .A2(new_n477_), .ZN(new_n478_) );
  XNOR2_X1 g120 ( .A(new_n478_), .B(new_n472_), .ZN(new_n479_) );
  AND4_X1 g121 ( .A1(new_n479_), .A2(new_n468_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n480_) );
  AND2_X1 g122 ( .A1(new_n480_), .A2(G860), .ZN(new_n481_) );
  INV_X1 g123 ( .A(new_n481_), .ZN(G153) );
  AND3_X1 g124 ( .A1(G319), .A2(G483), .A3(G661), .ZN(new_n483_) );
  AND2_X1 g125 ( .A1(new_n483_), .A2(G36), .ZN(new_n484_) );
  INV_X1 g126 ( .A(new_n484_), .ZN(G176) );
  AND2_X1 g127 ( .A1(G1), .A2(G3), .ZN(new_n486_) );
  INV_X1 g128 ( .A(new_n486_), .ZN(new_n487_) );
  AND2_X1 g129 ( .A1(new_n483_), .A2(new_n487_), .ZN(new_n488_) );
  INV_X1 g130 ( .A(new_n488_), .ZN(G188) );
  AND2_X1 g131 ( .A1(new_n436_), .A2(G78), .ZN(new_n490_) );
  AND2_X1 g132 ( .A1(new_n433_), .A2(G91), .ZN(new_n491_) );
  AND2_X1 g133 ( .A1(new_n430_), .A2(G65), .ZN(new_n492_) );
  AND2_X1 g134 ( .A1(new_n438_), .A2(G53), .ZN(new_n493_) );
  OR4_X1 g135 ( .A1(new_n492_), .A2(new_n490_), .A3(new_n493_), .A4(new_n491_), .ZN(G299) );
  XNOR2_X1 g136 ( .A(new_n452_), .B(KEYINPUT8), .ZN(G286) );
  AND2_X1 g137 ( .A1(new_n438_), .A2(G49), .ZN(new_n496_) );
  INV_X1 g138 ( .A(new_n496_), .ZN(new_n497_) );
  INV_X1 g139 ( .A(G87), .ZN(new_n498_) );
  OR2_X1 g140 ( .A1(new_n435_), .A2(new_n498_), .ZN(new_n499_) );
  AND2_X1 g141 ( .A1(G74), .A2(G651), .ZN(new_n500_) );
  INV_X1 g142 ( .A(new_n500_), .ZN(new_n501_) );
  AND3_X1 g143 ( .A1(new_n429_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_) );
  AND2_X1 g144 ( .A1(new_n502_), .A2(new_n497_), .ZN(new_n503_) );
  INV_X1 g145 ( .A(new_n503_), .ZN(G288) );
  AND2_X1 g146 ( .A1(new_n436_), .A2(G73), .ZN(new_n505_) );
  XNOR2_X1 g147 ( .A(new_n505_), .B(KEYINPUT2), .ZN(new_n506_) );
  AND2_X1 g148 ( .A1(new_n438_), .A2(G48), .ZN(new_n507_) );
  AND2_X1 g149 ( .A1(new_n430_), .A2(G61), .ZN(new_n508_) );
  AND2_X1 g150 ( .A1(new_n433_), .A2(G86), .ZN(new_n509_) );
  OR4_X1 g151 ( .A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .A4(new_n509_), .ZN(G305) );
  AND2_X1 g152 ( .A1(new_n436_), .A2(G72), .ZN(new_n511_) );
  AND2_X1 g153 ( .A1(new_n433_), .A2(G85), .ZN(new_n512_) );
  AND2_X1 g154 ( .A1(new_n430_), .A2(G60), .ZN(new_n513_) );
  AND2_X1 g155 ( .A1(new_n438_), .A2(G47), .ZN(new_n514_) );
  OR4_X1 g156 ( .A1(new_n513_), .A2(new_n511_), .A3(new_n514_), .A4(new_n512_), .ZN(G290) );
  INV_X1 g157 ( .A(G868), .ZN(new_n516_) );
  AND2_X1 g158 ( .A1(new_n436_), .A2(G79), .ZN(new_n517_) );
  INV_X1 g159 ( .A(new_n517_), .ZN(new_n518_) );
  INV_X1 g160 ( .A(G92), .ZN(new_n519_) );
  OR3_X1 g161 ( .A1(new_n519_), .A2(G543), .A3(G651), .ZN(new_n520_) );
  INV_X1 g162 ( .A(G66), .ZN(new_n521_) );
  OR2_X1 g163 ( .A1(new_n429_), .A2(new_n521_), .ZN(new_n522_) );
  AND2_X1 g164 ( .A1(new_n438_), .A2(G54), .ZN(new_n523_) );
  INV_X1 g165 ( .A(new_n523_), .ZN(new_n524_) );
  AND4_X1 g166 ( .A1(new_n518_), .A2(new_n524_), .A3(new_n522_), .A4(new_n520_), .ZN(new_n525_) );
  XOR2_X1 g167 ( .A(new_n525_), .B(KEYINPUT15), .Z(new_n526_) );
  INV_X1 g168 ( .A(new_n526_), .ZN(new_n527_) );
  AND2_X1 g169 ( .A1(new_n527_), .A2(new_n516_), .ZN(new_n528_) );
  AND2_X1 g170 ( .A1(G301), .A2(G868), .ZN(new_n529_) );
  OR2_X1 g171 ( .A1(new_n529_), .A2(new_n528_), .ZN(G284) );
  OR2_X1 g172 ( .A1(G286), .A2(new_n516_), .ZN(new_n531_) );
  OR2_X1 g173 ( .A1(G299), .A2(G868), .ZN(new_n532_) );
  AND2_X1 g174 ( .A1(new_n531_), .A2(new_n532_), .ZN(G297) );
  INV_X1 g175 ( .A(G559), .ZN(new_n534_) );
  OR2_X1 g176 ( .A1(new_n534_), .A2(G860), .ZN(new_n535_) );
  AND2_X1 g177 ( .A1(new_n526_), .A2(new_n535_), .ZN(new_n536_) );
  XOR2_X1 g178 ( .A(new_n536_), .B(KEYINPUT16), .Z(G148) );
  OR3_X1 g179 ( .A1(new_n527_), .A2(G559), .A3(new_n516_), .ZN(new_n538_) );
  AND2_X1 g180 ( .A1(new_n480_), .A2(new_n516_), .ZN(new_n539_) );
  INV_X1 g181 ( .A(new_n539_), .ZN(new_n540_) );
  AND2_X1 g182 ( .A1(new_n538_), .A2(new_n540_), .ZN(G282) );
  INV_X1 g183 ( .A(G2096), .ZN(new_n542_) );
  AND2_X1 g184 ( .A1(new_n408_), .A2(G135), .ZN(new_n543_) );
  AND2_X1 g185 ( .A1(new_n411_), .A2(G123), .ZN(new_n544_) );
  XNOR2_X1 g186 ( .A(new_n544_), .B(KEYINPUT18), .ZN(new_n545_) );
  AND2_X1 g187 ( .A1(new_n414_), .A2(G111), .ZN(new_n546_) );
  AND2_X1 g188 ( .A1(new_n416_), .A2(G99), .ZN(new_n547_) );
  OR4_X1 g189 ( .A1(new_n545_), .A2(new_n543_), .A3(new_n546_), .A4(new_n547_), .ZN(new_n548_) );
  INV_X1 g190 ( .A(new_n548_), .ZN(new_n549_) );
  AND2_X1 g191 ( .A1(new_n549_), .A2(new_n542_), .ZN(new_n550_) );
  AND2_X1 g192 ( .A1(new_n548_), .A2(G2096), .ZN(new_n551_) );
  OR3_X1 g193 ( .A1(new_n550_), .A2(G2100), .A3(new_n551_), .ZN(G156) );
  XNOR2_X1 g194 ( .A(G2430), .B(G2454), .ZN(new_n553_) );
  XNOR2_X1 g195 ( .A(G1341), .B(G1348), .ZN(new_n554_) );
  XOR2_X1 g196 ( .A(new_n553_), .B(new_n554_), .Z(new_n555_) );
  XNOR2_X1 g197 ( .A(G2435), .B(G2438), .ZN(new_n556_) );
  XNOR2_X1 g198 ( .A(new_n555_), .B(new_n556_), .ZN(new_n557_) );
  XOR2_X1 g199 ( .A(G2446), .B(G2451), .Z(new_n558_) );
  XNOR2_X1 g200 ( .A(G2427), .B(G2443), .ZN(new_n559_) );
  XOR2_X1 g201 ( .A(new_n558_), .B(new_n559_), .Z(new_n560_) );
  XNOR2_X1 g202 ( .A(new_n557_), .B(new_n560_), .ZN(new_n561_) );
  INV_X1 g203 ( .A(new_n561_), .ZN(new_n562_) );
  AND2_X1 g204 ( .A1(new_n562_), .A2(G14), .ZN(G401) );
  XNOR2_X1 g205 ( .A(G2090), .B(KEYINPUT42), .ZN(new_n564_) );
  XNOR2_X1 g206 ( .A(G2067), .B(G2072), .ZN(new_n565_) );
  XNOR2_X1 g207 ( .A(new_n564_), .B(new_n565_), .ZN(new_n566_) );
  XNOR2_X1 g208 ( .A(G2096), .B(G2100), .ZN(new_n567_) );
  XNOR2_X1 g209 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n568_) );
  XNOR2_X1 g210 ( .A(new_n567_), .B(new_n568_), .ZN(new_n569_) );
  XNOR2_X1 g211 ( .A(new_n566_), .B(new_n569_), .ZN(new_n570_) );
  XOR2_X1 g212 ( .A(G2078), .B(G2084), .Z(new_n571_) );
  XOR2_X1 g213 ( .A(new_n570_), .B(new_n571_), .Z(new_n572_) );
  INV_X1 g214 ( .A(new_n572_), .ZN(G227) );
  XOR2_X1 g215 ( .A(G1976), .B(G1981), .Z(new_n574_) );
  XNOR2_X1 g216 ( .A(G1956), .B(G1966), .ZN(new_n575_) );
  XNOR2_X1 g217 ( .A(new_n574_), .B(new_n575_), .ZN(new_n576_) );
  XNOR2_X1 g218 ( .A(new_n576_), .B(G2474), .ZN(new_n577_) );
  XNOR2_X1 g219 ( .A(G1991), .B(G1996), .ZN(new_n578_) );
  XNOR2_X1 g220 ( .A(new_n577_), .B(new_n578_), .ZN(new_n579_) );
  XNOR2_X1 g221 ( .A(G1971), .B(KEYINPUT41), .ZN(new_n580_) );
  XNOR2_X1 g222 ( .A(G1961), .B(G1986), .ZN(new_n581_) );
  XNOR2_X1 g223 ( .A(new_n580_), .B(new_n581_), .ZN(new_n582_) );
  XOR2_X1 g224 ( .A(new_n579_), .B(new_n582_), .Z(new_n583_) );
  INV_X1 g225 ( .A(new_n583_), .ZN(G229) );
  INV_X1 g226 ( .A(G29), .ZN(new_n585_) );
  INV_X1 g227 ( .A(KEYINPUT55), .ZN(new_n586_) );
  INV_X1 g228 ( .A(KEYINPUT52), .ZN(new_n587_) );
  INV_X1 g229 ( .A(G2090), .ZN(new_n588_) );
  AND2_X1 g230 ( .A1(G162), .A2(new_n588_), .ZN(new_n589_) );
  AND2_X1 g231 ( .A1(new_n418_), .A2(G2090), .ZN(new_n590_) );
  INV_X1 g232 ( .A(G1996), .ZN(new_n591_) );
  AND2_X1 g233 ( .A1(new_n408_), .A2(G141), .ZN(new_n592_) );
  AND2_X1 g234 ( .A1(new_n416_), .A2(G105), .ZN(new_n593_) );
  OR2_X1 g235 ( .A1(new_n593_), .A2(KEYINPUT38), .ZN(new_n594_) );
  INV_X1 g236 ( .A(new_n594_), .ZN(new_n595_) );
  AND2_X1 g237 ( .A1(new_n593_), .A2(KEYINPUT38), .ZN(new_n596_) );
  AND2_X1 g238 ( .A1(new_n411_), .A2(G129), .ZN(new_n597_) );
  AND2_X1 g239 ( .A1(new_n414_), .A2(G117), .ZN(new_n598_) );
  OR2_X1 g240 ( .A1(new_n597_), .A2(new_n598_), .ZN(new_n599_) );
  OR4_X1 g241 ( .A1(new_n595_), .A2(new_n592_), .A3(new_n596_), .A4(new_n599_), .ZN(new_n600_) );
  INV_X1 g242 ( .A(new_n600_), .ZN(new_n601_) );
  AND2_X1 g243 ( .A1(new_n601_), .A2(new_n591_), .ZN(new_n602_) );
  OR3_X1 g244 ( .A1(new_n589_), .A2(new_n602_), .A3(new_n590_), .ZN(new_n603_) );
  INV_X1 g245 ( .A(new_n603_), .ZN(new_n604_) );
  OR2_X1 g246 ( .A1(new_n604_), .A2(KEYINPUT51), .ZN(new_n605_) );
  INV_X1 g247 ( .A(KEYINPUT51), .ZN(new_n606_) );
  OR2_X1 g248 ( .A1(new_n603_), .A2(new_n606_), .ZN(new_n607_) );
  INV_X1 g249 ( .A(KEYINPUT50), .ZN(new_n608_) );
  AND2_X1 g250 ( .A1(new_n414_), .A2(G115), .ZN(new_n609_) );
  AND2_X1 g251 ( .A1(new_n411_), .A2(G127), .ZN(new_n610_) );
  OR2_X1 g252 ( .A1(new_n610_), .A2(new_n609_), .ZN(new_n611_) );
  XOR2_X1 g253 ( .A(new_n611_), .B(KEYINPUT47), .Z(new_n612_) );
  AND2_X1 g254 ( .A1(new_n416_), .A2(G103), .ZN(new_n613_) );
  AND2_X1 g255 ( .A1(new_n408_), .A2(G139), .ZN(new_n614_) );
  OR3_X1 g256 ( .A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_) );
  INV_X1 g257 ( .A(new_n615_), .ZN(new_n616_) );
  OR2_X1 g258 ( .A1(new_n616_), .A2(new_n367_), .ZN(new_n617_) );
  OR2_X1 g259 ( .A1(new_n615_), .A2(G2072), .ZN(new_n618_) );
  XOR2_X1 g260 ( .A(new_n425_), .B(G2078), .Z(new_n619_) );
  AND3_X1 g261 ( .A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_) );
  OR2_X1 g262 ( .A1(new_n620_), .A2(new_n608_), .ZN(new_n621_) );
  AND3_X1 g263 ( .A1(new_n621_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n622_) );
  INV_X1 g264 ( .A(KEYINPUT34), .ZN(new_n623_) );
  AND2_X1 g265 ( .A1(new_n408_), .A2(G140), .ZN(new_n624_) );
  AND2_X1 g266 ( .A1(new_n416_), .A2(G104), .ZN(new_n625_) );
  OR2_X1 g267 ( .A1(new_n624_), .A2(new_n625_), .ZN(new_n626_) );
  INV_X1 g268 ( .A(new_n626_), .ZN(new_n627_) );
  OR2_X1 g269 ( .A1(new_n627_), .A2(new_n623_), .ZN(new_n628_) );
  AND2_X1 g270 ( .A1(new_n414_), .A2(G116), .ZN(new_n629_) );
  AND2_X1 g271 ( .A1(new_n411_), .A2(G128), .ZN(new_n630_) );
  OR2_X1 g272 ( .A1(new_n630_), .A2(new_n629_), .ZN(new_n631_) );
  XNOR2_X1 g273 ( .A(new_n631_), .B(KEYINPUT35), .ZN(new_n632_) );
  OR2_X1 g274 ( .A1(new_n626_), .A2(KEYINPUT34), .ZN(new_n633_) );
  AND3_X1 g275 ( .A1(new_n628_), .A2(new_n633_), .A3(new_n632_), .ZN(new_n634_) );
  XNOR2_X1 g276 ( .A(new_n634_), .B(KEYINPUT36), .ZN(new_n635_) );
  INV_X1 g277 ( .A(new_n635_), .ZN(new_n636_) );
  XNOR2_X1 g278 ( .A(G2067), .B(KEYINPUT37), .ZN(new_n637_) );
  INV_X1 g279 ( .A(new_n637_), .ZN(new_n638_) );
  AND2_X1 g280 ( .A1(new_n636_), .A2(new_n638_), .ZN(new_n639_) );
  INV_X1 g281 ( .A(new_n639_), .ZN(new_n640_) );
  OR2_X1 g282 ( .A1(new_n636_), .A2(new_n638_), .ZN(new_n641_) );
  AND2_X1 g283 ( .A1(new_n620_), .A2(new_n608_), .ZN(new_n642_) );
  INV_X1 g284 ( .A(new_n642_), .ZN(new_n643_) );
  AND2_X1 g285 ( .A1(new_n600_), .A2(G1996), .ZN(new_n644_) );
  AND2_X1 g286 ( .A1(new_n408_), .A2(G131), .ZN(new_n645_) );
  AND2_X1 g287 ( .A1(new_n411_), .A2(G119), .ZN(new_n646_) );
  AND2_X1 g288 ( .A1(new_n416_), .A2(G95), .ZN(new_n647_) );
  AND2_X1 g289 ( .A1(new_n414_), .A2(G107), .ZN(new_n648_) );
  OR4_X1 g290 ( .A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .A4(new_n648_), .ZN(new_n649_) );
  AND2_X1 g291 ( .A1(new_n649_), .A2(G1991), .ZN(new_n650_) );
  OR2_X1 g292 ( .A1(new_n644_), .A2(new_n650_), .ZN(new_n651_) );
  INV_X1 g293 ( .A(new_n651_), .ZN(new_n652_) );
  XNOR2_X1 g294 ( .A(G160), .B(G2084), .ZN(new_n653_) );
  OR2_X1 g295 ( .A1(new_n649_), .A2(G1991), .ZN(new_n654_) );
  AND4_X1 g296 ( .A1(new_n652_), .A2(new_n548_), .A3(new_n653_), .A4(new_n654_), .ZN(new_n655_) );
  AND2_X1 g297 ( .A1(new_n643_), .A2(new_n655_), .ZN(new_n656_) );
  AND4_X1 g298 ( .A1(new_n656_), .A2(new_n622_), .A3(new_n640_), .A4(new_n641_), .ZN(new_n657_) );
  AND2_X1 g299 ( .A1(new_n657_), .A2(new_n587_), .ZN(new_n658_) );
  INV_X1 g300 ( .A(new_n658_), .ZN(new_n659_) );
  OR2_X1 g301 ( .A1(new_n657_), .A2(new_n587_), .ZN(new_n660_) );
  AND3_X1 g302 ( .A1(new_n659_), .A2(new_n586_), .A3(new_n660_), .ZN(new_n661_) );
  OR2_X1 g303 ( .A1(new_n661_), .A2(new_n585_), .ZN(new_n662_) );
  XNOR2_X1 g304 ( .A(new_n452_), .B(G1966), .ZN(new_n663_) );
  INV_X1 g305 ( .A(G1981), .ZN(new_n664_) );
  XNOR2_X1 g306 ( .A(G305), .B(new_n664_), .ZN(new_n665_) );
  INV_X1 g307 ( .A(new_n665_), .ZN(new_n666_) );
  OR2_X1 g308 ( .A1(new_n663_), .A2(new_n666_), .ZN(new_n667_) );
  XNOR2_X1 g309 ( .A(new_n667_), .B(KEYINPUT57), .ZN(new_n668_) );
  XNOR2_X1 g310 ( .A(new_n526_), .B(G1348), .ZN(new_n669_) );
  INV_X1 g311 ( .A(G1956), .ZN(new_n670_) );
  XNOR2_X1 g312 ( .A(G299), .B(new_n670_), .ZN(new_n671_) );
  AND2_X1 g313 ( .A1(G288), .A2(G1976), .ZN(new_n672_) );
  INV_X1 g314 ( .A(new_n672_), .ZN(new_n673_) );
  INV_X1 g315 ( .A(G1971), .ZN(new_n674_) );
  OR2_X1 g316 ( .A1(G166), .A2(new_n674_), .ZN(new_n675_) );
  AND2_X1 g317 ( .A1(new_n675_), .A2(new_n673_), .ZN(new_n676_) );
  OR2_X1 g318 ( .A1(G303), .A2(G1971), .ZN(new_n677_) );
  INV_X1 g319 ( .A(G1976), .ZN(new_n678_) );
  AND2_X1 g320 ( .A1(new_n503_), .A2(new_n678_), .ZN(new_n679_) );
  INV_X1 g321 ( .A(new_n679_), .ZN(new_n680_) );
  AND2_X1 g322 ( .A1(new_n677_), .A2(new_n680_), .ZN(new_n681_) );
  INV_X1 g323 ( .A(G1986), .ZN(new_n682_) );
  XNOR2_X1 g324 ( .A(G290), .B(new_n682_), .ZN(new_n683_) );
  AND4_X1 g325 ( .A1(new_n676_), .A2(new_n671_), .A3(new_n681_), .A4(new_n683_), .ZN(new_n684_) );
  XOR2_X1 g326 ( .A(G301), .B(G1961), .Z(new_n685_) );
  XNOR2_X1 g327 ( .A(new_n480_), .B(G1341), .ZN(new_n686_) );
  AND4_X1 g328 ( .A1(new_n685_), .A2(new_n669_), .A3(new_n684_), .A4(new_n686_), .ZN(new_n687_) );
  AND2_X1 g329 ( .A1(new_n668_), .A2(new_n687_), .ZN(new_n688_) );
  XOR2_X1 g330 ( .A(G16), .B(KEYINPUT56), .Z(new_n689_) );
  OR2_X1 g331 ( .A1(new_n688_), .A2(new_n689_), .ZN(new_n690_) );
  OR2_X1 g332 ( .A1(G26), .A2(G2067), .ZN(new_n691_) );
  AND2_X1 g333 ( .A1(new_n691_), .A2(G28), .ZN(new_n692_) );
  AND2_X1 g334 ( .A1(G33), .A2(G2072), .ZN(new_n693_) );
  INV_X1 g335 ( .A(new_n693_), .ZN(new_n694_) );
  AND2_X1 g336 ( .A1(G26), .A2(G2067), .ZN(new_n695_) );
  INV_X1 g337 ( .A(new_n695_), .ZN(new_n696_) );
  XOR2_X1 g338 ( .A(G32), .B(G1996), .Z(new_n697_) );
  AND4_X1 g339 ( .A1(new_n692_), .A2(new_n697_), .A3(new_n694_), .A4(new_n696_), .ZN(new_n698_) );
  XNOR2_X1 g340 ( .A(G2078), .B(KEYINPUT25), .ZN(new_n699_) );
  INV_X1 g341 ( .A(new_n699_), .ZN(new_n700_) );
  OR2_X1 g342 ( .A1(new_n700_), .A2(G27), .ZN(new_n701_) );
  INV_X1 g343 ( .A(G27), .ZN(new_n702_) );
  OR2_X1 g344 ( .A1(new_n699_), .A2(new_n702_), .ZN(new_n703_) );
  OR2_X1 g345 ( .A1(G25), .A2(G1991), .ZN(new_n704_) );
  OR2_X1 g346 ( .A1(G33), .A2(G2072), .ZN(new_n705_) );
  AND2_X1 g347 ( .A1(G25), .A2(G1991), .ZN(new_n706_) );
  INV_X1 g348 ( .A(new_n706_), .ZN(new_n707_) );
  AND3_X1 g349 ( .A1(new_n707_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n708_) );
  AND4_X1 g350 ( .A1(new_n698_), .A2(new_n701_), .A3(new_n703_), .A4(new_n708_), .ZN(new_n709_) );
  OR2_X1 g351 ( .A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n710_) );
  AND2_X1 g352 ( .A1(new_n709_), .A2(KEYINPUT53), .ZN(new_n711_) );
  INV_X1 g353 ( .A(new_n711_), .ZN(new_n712_) );
  XOR2_X1 g354 ( .A(G35), .B(G2090), .Z(new_n713_) );
  XOR2_X1 g355 ( .A(G2084), .B(KEYINPUT54), .Z(new_n714_) );
  XNOR2_X1 g356 ( .A(new_n714_), .B(G34), .ZN(new_n715_) );
  AND4_X1 g357 ( .A1(new_n712_), .A2(new_n710_), .A3(new_n713_), .A4(new_n715_), .ZN(new_n716_) );
  AND2_X1 g358 ( .A1(new_n716_), .A2(new_n586_), .ZN(new_n717_) );
  INV_X1 g359 ( .A(new_n717_), .ZN(new_n718_) );
  OR2_X1 g360 ( .A1(new_n716_), .A2(new_n586_), .ZN(new_n719_) );
  AND3_X1 g361 ( .A1(new_n718_), .A2(new_n585_), .A3(new_n719_), .ZN(new_n720_) );
  INV_X1 g362 ( .A(new_n720_), .ZN(new_n721_) );
  INV_X1 g363 ( .A(KEYINPUT61), .ZN(new_n722_) );
  XOR2_X1 g364 ( .A(G20), .B(G1956), .Z(new_n723_) );
  OR2_X1 g365 ( .A1(G19), .A2(G1341), .ZN(new_n724_) );
  OR2_X1 g366 ( .A1(G6), .A2(G1981), .ZN(new_n725_) );
  AND2_X1 g367 ( .A1(G19), .A2(G1341), .ZN(new_n726_) );
  INV_X1 g368 ( .A(new_n726_), .ZN(new_n727_) );
  AND2_X1 g369 ( .A1(G6), .A2(G1981), .ZN(new_n728_) );
  INV_X1 g370 ( .A(new_n728_), .ZN(new_n729_) );
  AND4_X1 g371 ( .A1(new_n727_), .A2(new_n729_), .A3(new_n724_), .A4(new_n725_), .ZN(new_n730_) );
  XNOR2_X1 g372 ( .A(G1348), .B(KEYINPUT59), .ZN(new_n731_) );
  XNOR2_X1 g373 ( .A(new_n731_), .B(G4), .ZN(new_n732_) );
  AND3_X1 g374 ( .A1(new_n732_), .A2(new_n723_), .A3(new_n730_), .ZN(new_n733_) );
  XOR2_X1 g375 ( .A(new_n733_), .B(KEYINPUT60), .Z(new_n734_) );
  INV_X1 g376 ( .A(new_n734_), .ZN(new_n735_) );
  INV_X1 g377 ( .A(KEYINPUT58), .ZN(new_n736_) );
  XNOR2_X1 g378 ( .A(G24), .B(G1986), .ZN(new_n737_) );
  INV_X1 g379 ( .A(new_n737_), .ZN(new_n738_) );
  AND2_X1 g380 ( .A1(G23), .A2(G1976), .ZN(new_n739_) );
  INV_X1 g381 ( .A(new_n739_), .ZN(new_n740_) );
  AND2_X1 g382 ( .A1(G22), .A2(G1971), .ZN(new_n741_) );
  INV_X1 g383 ( .A(new_n741_), .ZN(new_n742_) );
  OR2_X1 g384 ( .A1(G23), .A2(G1976), .ZN(new_n743_) );
  OR2_X1 g385 ( .A1(G22), .A2(G1971), .ZN(new_n744_) );
  AND2_X1 g386 ( .A1(new_n743_), .A2(new_n744_), .ZN(new_n745_) );
  AND4_X1 g387 ( .A1(new_n745_), .A2(new_n738_), .A3(new_n740_), .A4(new_n742_), .ZN(new_n746_) );
  OR2_X1 g388 ( .A1(new_n746_), .A2(new_n736_), .ZN(new_n747_) );
  AND2_X1 g389 ( .A1(new_n746_), .A2(new_n736_), .ZN(new_n748_) );
  INV_X1 g390 ( .A(new_n748_), .ZN(new_n749_) );
  XOR2_X1 g391 ( .A(G5), .B(G1961), .Z(new_n750_) );
  XOR2_X1 g392 ( .A(G21), .B(G1966), .Z(new_n751_) );
  AND4_X1 g393 ( .A1(new_n749_), .A2(new_n747_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n752_) );
  AND2_X1 g394 ( .A1(new_n735_), .A2(new_n752_), .ZN(new_n753_) );
  AND2_X1 g395 ( .A1(new_n753_), .A2(new_n722_), .ZN(new_n754_) );
  INV_X1 g396 ( .A(new_n753_), .ZN(new_n755_) );
  AND2_X1 g397 ( .A1(new_n755_), .A2(KEYINPUT61), .ZN(new_n756_) );
  OR3_X1 g398 ( .A1(new_n756_), .A2(new_n754_), .A3(G16), .ZN(new_n757_) );
  AND3_X1 g399 ( .A1(new_n757_), .A2(G11), .A3(new_n721_), .ZN(new_n758_) );
  AND3_X1 g400 ( .A1(new_n662_), .A2(new_n690_), .A3(new_n758_), .ZN(new_n759_) );
  XNOR2_X1 g401 ( .A(new_n759_), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 g402 ( .A(G311), .ZN(G150) );
  AND2_X1 g403 ( .A1(new_n526_), .A2(G559), .ZN(new_n762_) );
  AND2_X1 g404 ( .A1(new_n762_), .A2(new_n480_), .ZN(new_n763_) );
  INV_X1 g405 ( .A(new_n480_), .ZN(new_n764_) );
  INV_X1 g406 ( .A(new_n762_), .ZN(new_n765_) );
  AND2_X1 g407 ( .A1(new_n765_), .A2(new_n764_), .ZN(new_n766_) );
  OR3_X1 g408 ( .A1(new_n766_), .A2(new_n763_), .A3(G860), .ZN(new_n767_) );
  AND2_X1 g409 ( .A1(new_n436_), .A2(G80), .ZN(new_n768_) );
  AND2_X1 g410 ( .A1(new_n433_), .A2(G93), .ZN(new_n769_) );
  AND2_X1 g411 ( .A1(new_n430_), .A2(G67), .ZN(new_n770_) );
  AND2_X1 g412 ( .A1(new_n438_), .A2(G55), .ZN(new_n771_) );
  OR4_X1 g413 ( .A1(new_n770_), .A2(new_n768_), .A3(new_n771_), .A4(new_n769_), .ZN(new_n772_) );
  XNOR2_X1 g414 ( .A(new_n767_), .B(new_n772_), .ZN(G145) );
  INV_X1 g415 ( .A(G37), .ZN(new_n774_) );
  XNOR2_X1 g416 ( .A(new_n615_), .B(G160), .ZN(new_n775_) );
  XNOR2_X1 g417 ( .A(new_n635_), .B(new_n775_), .ZN(new_n776_) );
  AND2_X1 g418 ( .A1(new_n408_), .A2(G142), .ZN(new_n777_) );
  AND2_X1 g419 ( .A1(new_n416_), .A2(G106), .ZN(new_n778_) );
  OR2_X1 g420 ( .A1(new_n777_), .A2(new_n778_), .ZN(new_n779_) );
  INV_X1 g421 ( .A(new_n779_), .ZN(new_n780_) );
  AND2_X1 g422 ( .A1(new_n780_), .A2(KEYINPUT45), .ZN(new_n781_) );
  INV_X1 g423 ( .A(KEYINPUT45), .ZN(new_n782_) );
  AND2_X1 g424 ( .A1(new_n779_), .A2(new_n782_), .ZN(new_n783_) );
  AND2_X1 g425 ( .A1(new_n411_), .A2(G130), .ZN(new_n784_) );
  AND2_X1 g426 ( .A1(new_n414_), .A2(G118), .ZN(new_n785_) );
  OR4_X1 g427 ( .A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .A4(new_n785_), .ZN(new_n786_) );
  XNOR2_X1 g428 ( .A(new_n786_), .B(new_n601_), .ZN(new_n787_) );
  XNOR2_X1 g429 ( .A(new_n787_), .B(new_n418_), .ZN(new_n788_) );
  XNOR2_X1 g430 ( .A(new_n788_), .B(new_n776_), .ZN(new_n789_) );
  XNOR2_X1 g431 ( .A(new_n548_), .B(new_n649_), .ZN(new_n790_) );
  XNOR2_X1 g432 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(new_n791_) );
  XNOR2_X1 g433 ( .A(new_n790_), .B(new_n791_), .ZN(new_n792_) );
  XNOR2_X1 g434 ( .A(new_n792_), .B(new_n425_), .ZN(new_n793_) );
  AND2_X1 g435 ( .A1(new_n789_), .A2(new_n793_), .ZN(new_n794_) );
  INV_X1 g436 ( .A(new_n794_), .ZN(new_n795_) );
  OR2_X1 g437 ( .A1(new_n789_), .A2(new_n793_), .ZN(new_n796_) );
  AND3_X1 g438 ( .A1(new_n795_), .A2(new_n774_), .A3(new_n796_), .ZN(G395) );
  XNOR2_X1 g439 ( .A(new_n480_), .B(G290), .ZN(new_n798_) );
  XNOR2_X1 g440 ( .A(new_n798_), .B(G288), .ZN(new_n799_) );
  XNOR2_X1 g441 ( .A(G299), .B(KEYINPUT19), .ZN(new_n800_) );
  XNOR2_X1 g442 ( .A(new_n800_), .B(G305), .ZN(new_n801_) );
  XNOR2_X1 g443 ( .A(new_n799_), .B(new_n801_), .ZN(new_n802_) );
  XNOR2_X1 g444 ( .A(G303), .B(new_n772_), .ZN(new_n803_) );
  XNOR2_X1 g445 ( .A(new_n802_), .B(new_n803_), .ZN(new_n804_) );
  XNOR2_X1 g446 ( .A(new_n804_), .B(new_n765_), .ZN(new_n805_) );
  AND2_X1 g447 ( .A1(new_n805_), .A2(G868), .ZN(new_n806_) );
  AND2_X1 g448 ( .A1(new_n772_), .A2(new_n516_), .ZN(new_n807_) );
  OR2_X1 g449 ( .A1(new_n806_), .A2(new_n807_), .ZN(G295) );
  XNOR2_X1 g450 ( .A(G286), .B(new_n526_), .ZN(new_n809_) );
  XNOR2_X1 g451 ( .A(new_n804_), .B(new_n809_), .ZN(new_n810_) );
  AND2_X1 g452 ( .A1(new_n810_), .A2(G301), .ZN(new_n811_) );
  INV_X1 g453 ( .A(new_n811_), .ZN(new_n812_) );
  OR2_X1 g454 ( .A1(new_n810_), .A2(G301), .ZN(new_n813_) );
  AND3_X1 g455 ( .A1(new_n812_), .A2(new_n774_), .A3(new_n813_), .ZN(G397) );
  INV_X1 g456 ( .A(KEYINPUT40), .ZN(new_n815_) );
  INV_X1 g457 ( .A(KEYINPUT33), .ZN(new_n816_) );
  INV_X1 g458 ( .A(G1384), .ZN(new_n817_) );
  AND4_X1 g459 ( .A1(new_n397_), .A2(G40), .A3(new_n400_), .A4(new_n406_), .ZN(new_n818_) );
  AND3_X1 g460 ( .A1(new_n818_), .A2(new_n817_), .A3(new_n425_), .ZN(new_n819_) );
  AND2_X1 g461 ( .A1(new_n819_), .A2(G2067), .ZN(new_n820_) );
  INV_X1 g462 ( .A(new_n820_), .ZN(new_n821_) );
  INV_X1 g463 ( .A(G1348), .ZN(new_n822_) );
  OR2_X1 g464 ( .A1(new_n819_), .A2(new_n822_), .ZN(new_n823_) );
  AND2_X1 g465 ( .A1(new_n821_), .A2(new_n823_), .ZN(new_n824_) );
  INV_X1 g466 ( .A(KEYINPUT26), .ZN(new_n825_) );
  AND4_X1 g467 ( .A1(new_n818_), .A2(new_n817_), .A3(G1996), .A4(new_n425_), .ZN(new_n826_) );
  XNOR2_X1 g468 ( .A(new_n826_), .B(new_n825_), .ZN(new_n827_) );
  INV_X1 g469 ( .A(G1341), .ZN(new_n828_) );
  OR2_X1 g470 ( .A1(new_n819_), .A2(new_n828_), .ZN(new_n829_) );
  AND4_X1 g471 ( .A1(new_n827_), .A2(new_n480_), .A3(new_n526_), .A4(new_n829_), .ZN(new_n830_) );
  OR2_X1 g472 ( .A1(new_n830_), .A2(new_n824_), .ZN(new_n831_) );
  AND3_X1 g473 ( .A1(new_n827_), .A2(new_n480_), .A3(new_n829_), .ZN(new_n832_) );
  OR2_X1 g474 ( .A1(new_n832_), .A2(new_n526_), .ZN(new_n833_) );
  AND2_X1 g475 ( .A1(new_n831_), .A2(new_n833_), .ZN(new_n834_) );
  INV_X1 g476 ( .A(G299), .ZN(new_n835_) );
  INV_X1 g477 ( .A(KEYINPUT27), .ZN(new_n836_) );
  AND2_X1 g478 ( .A1(new_n425_), .A2(new_n817_), .ZN(new_n837_) );
  AND3_X1 g479 ( .A1(new_n837_), .A2(G2072), .A3(new_n818_), .ZN(new_n838_) );
  AND2_X1 g480 ( .A1(new_n838_), .A2(new_n836_), .ZN(new_n839_) );
  INV_X1 g481 ( .A(new_n839_), .ZN(new_n840_) );
  OR2_X1 g482 ( .A1(new_n819_), .A2(new_n670_), .ZN(new_n841_) );
  OR2_X1 g483 ( .A1(new_n838_), .A2(new_n836_), .ZN(new_n842_) );
  AND3_X1 g484 ( .A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_) );
  AND2_X1 g485 ( .A1(new_n843_), .A2(new_n835_), .ZN(new_n844_) );
  OR2_X1 g486 ( .A1(new_n834_), .A2(new_n844_), .ZN(new_n845_) );
  OR2_X1 g487 ( .A1(new_n843_), .A2(new_n835_), .ZN(new_n846_) );
  XNOR2_X1 g488 ( .A(new_n846_), .B(KEYINPUT28), .ZN(new_n847_) );
  AND2_X1 g489 ( .A1(new_n845_), .A2(new_n847_), .ZN(new_n848_) );
  XNOR2_X1 g490 ( .A(new_n848_), .B(KEYINPUT29), .ZN(new_n849_) );
  AND2_X1 g491 ( .A1(new_n819_), .A2(new_n699_), .ZN(new_n850_) );
  INV_X1 g492 ( .A(new_n850_), .ZN(new_n851_) );
  OR2_X1 g493 ( .A1(new_n819_), .A2(G1961), .ZN(new_n852_) );
  AND2_X1 g494 ( .A1(new_n851_), .A2(new_n852_), .ZN(new_n853_) );
  OR2_X1 g495 ( .A1(new_n853_), .A2(G301), .ZN(new_n854_) );
  AND2_X1 g496 ( .A1(new_n849_), .A2(new_n854_), .ZN(new_n855_) );
  INV_X1 g497 ( .A(G8), .ZN(new_n856_) );
  OR2_X1 g498 ( .A1(new_n819_), .A2(new_n856_), .ZN(new_n857_) );
  OR2_X1 g499 ( .A1(new_n857_), .A2(G1966), .ZN(new_n858_) );
  INV_X1 g500 ( .A(new_n858_), .ZN(new_n859_) );
  INV_X1 g501 ( .A(G2084), .ZN(new_n860_) );
  AND2_X1 g502 ( .A1(new_n819_), .A2(new_n860_), .ZN(new_n861_) );
  OR4_X1 g503 ( .A1(new_n859_), .A2(new_n856_), .A3(KEYINPUT30), .A4(new_n861_), .ZN(new_n862_) );
  INV_X1 g504 ( .A(KEYINPUT30), .ZN(new_n863_) );
  INV_X1 g505 ( .A(new_n861_), .ZN(new_n864_) );
  AND3_X1 g506 ( .A1(new_n858_), .A2(G8), .A3(new_n864_), .ZN(new_n865_) );
  OR2_X1 g507 ( .A1(new_n865_), .A2(new_n863_), .ZN(new_n866_) );
  AND3_X1 g508 ( .A1(new_n866_), .A2(new_n452_), .A3(new_n862_), .ZN(new_n867_) );
  AND2_X1 g509 ( .A1(new_n853_), .A2(G301), .ZN(new_n868_) );
  OR2_X1 g510 ( .A1(new_n867_), .A2(new_n868_), .ZN(new_n869_) );
  XOR2_X1 g511 ( .A(new_n869_), .B(KEYINPUT31), .Z(new_n870_) );
  OR2_X1 g512 ( .A1(new_n855_), .A2(new_n870_), .ZN(new_n871_) );
  AND2_X1 g513 ( .A1(new_n871_), .A2(G286), .ZN(new_n872_) );
  OR2_X1 g514 ( .A1(new_n857_), .A2(G1971), .ZN(new_n873_) );
  AND2_X1 g515 ( .A1(new_n819_), .A2(new_n588_), .ZN(new_n874_) );
  INV_X1 g516 ( .A(new_n874_), .ZN(new_n875_) );
  AND3_X1 g517 ( .A1(new_n873_), .A2(G303), .A3(new_n875_), .ZN(new_n876_) );
  OR2_X1 g518 ( .A1(new_n872_), .A2(new_n876_), .ZN(new_n877_) );
  AND2_X1 g519 ( .A1(new_n877_), .A2(G8), .ZN(new_n878_) );
  XNOR2_X1 g520 ( .A(new_n878_), .B(KEYINPUT32), .ZN(new_n879_) );
  OR2_X1 g521 ( .A1(new_n864_), .A2(new_n856_), .ZN(new_n880_) );
  AND3_X1 g522 ( .A1(new_n871_), .A2(new_n858_), .A3(new_n880_), .ZN(new_n881_) );
  OR2_X1 g523 ( .A1(new_n879_), .A2(new_n881_), .ZN(new_n882_) );
  AND2_X1 g524 ( .A1(new_n882_), .A2(new_n681_), .ZN(new_n883_) );
  OR2_X1 g525 ( .A1(new_n857_), .A2(new_n672_), .ZN(new_n884_) );
  OR2_X1 g526 ( .A1(new_n883_), .A2(new_n884_), .ZN(new_n885_) );
  AND2_X1 g527 ( .A1(new_n885_), .A2(new_n816_), .ZN(new_n886_) );
  INV_X1 g528 ( .A(new_n857_), .ZN(new_n887_) );
  AND3_X1 g529 ( .A1(new_n887_), .A2(KEYINPUT33), .A3(new_n679_), .ZN(new_n888_) );
  OR2_X1 g530 ( .A1(new_n666_), .A2(new_n888_), .ZN(new_n889_) );
  OR2_X1 g531 ( .A1(new_n886_), .A2(new_n889_), .ZN(new_n890_) );
  OR3_X1 g532 ( .A1(G303), .A2(new_n856_), .A3(G2090), .ZN(new_n891_) );
  AND2_X1 g533 ( .A1(new_n882_), .A2(new_n891_), .ZN(new_n892_) );
  OR2_X1 g534 ( .A1(new_n892_), .A2(new_n887_), .ZN(new_n893_) );
  INV_X1 g535 ( .A(KEYINPUT24), .ZN(new_n894_) );
  INV_X1 g536 ( .A(G305), .ZN(new_n895_) );
  AND2_X1 g537 ( .A1(new_n895_), .A2(new_n664_), .ZN(new_n896_) );
  AND2_X1 g538 ( .A1(new_n896_), .A2(new_n894_), .ZN(new_n897_) );
  INV_X1 g539 ( .A(new_n896_), .ZN(new_n898_) );
  AND2_X1 g540 ( .A1(new_n898_), .A2(KEYINPUT24), .ZN(new_n899_) );
  OR3_X1 g541 ( .A1(new_n899_), .A2(new_n857_), .A3(new_n897_), .ZN(new_n900_) );
  AND2_X1 g542 ( .A1(new_n893_), .A2(new_n900_), .ZN(new_n901_) );
  AND2_X1 g543 ( .A1(new_n890_), .A2(new_n901_), .ZN(new_n902_) );
  INV_X1 g544 ( .A(new_n837_), .ZN(new_n903_) );
  AND2_X1 g545 ( .A1(new_n903_), .A2(new_n818_), .ZN(new_n904_) );
  AND2_X1 g546 ( .A1(new_n639_), .A2(new_n904_), .ZN(new_n905_) );
  INV_X1 g547 ( .A(new_n683_), .ZN(new_n906_) );
  AND2_X1 g548 ( .A1(new_n906_), .A2(new_n904_), .ZN(new_n907_) );
  AND2_X1 g549 ( .A1(new_n651_), .A2(new_n904_), .ZN(new_n908_) );
  OR3_X1 g550 ( .A1(new_n905_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_) );
  OR2_X1 g551 ( .A1(new_n902_), .A2(new_n909_), .ZN(new_n910_) );
  INV_X1 g552 ( .A(new_n904_), .ZN(new_n911_) );
  INV_X1 g553 ( .A(new_n602_), .ZN(new_n912_) );
  OR2_X1 g554 ( .A1(G290), .A2(G1986), .ZN(new_n913_) );
  AND2_X1 g555 ( .A1(new_n913_), .A2(new_n654_), .ZN(new_n914_) );
  OR2_X1 g556 ( .A1(new_n908_), .A2(new_n914_), .ZN(new_n915_) );
  AND2_X1 g557 ( .A1(new_n915_), .A2(new_n912_), .ZN(new_n916_) );
  XOR2_X1 g558 ( .A(new_n916_), .B(KEYINPUT39), .Z(new_n917_) );
  OR2_X1 g559 ( .A1(new_n917_), .A2(new_n905_), .ZN(new_n918_) );
  AND2_X1 g560 ( .A1(new_n918_), .A2(new_n641_), .ZN(new_n919_) );
  OR2_X1 g561 ( .A1(new_n919_), .A2(new_n911_), .ZN(new_n920_) );
  AND2_X1 g562 ( .A1(new_n910_), .A2(new_n920_), .ZN(new_n921_) );
  XNOR2_X1 g563 ( .A(new_n921_), .B(new_n815_), .ZN(G329) );
  INV_X1 g564 ( .A(G401), .ZN(new_n924_) );
  AND2_X1 g565 ( .A1(new_n583_), .A2(new_n572_), .ZN(new_n925_) );
  AND2_X1 g566 ( .A1(new_n925_), .A2(KEYINPUT49), .ZN(new_n926_) );
  INV_X1 g567 ( .A(new_n926_), .ZN(new_n927_) );
  OR2_X1 g568 ( .A1(new_n925_), .A2(KEYINPUT49), .ZN(new_n928_) );
  AND4_X1 g569 ( .A1(new_n927_), .A2(G319), .A3(new_n924_), .A4(new_n928_), .ZN(new_n929_) );
  INV_X1 g570 ( .A(new_n929_), .ZN(new_n930_) );
  OR3_X1 g571 ( .A1(G397), .A2(G395), .A3(new_n930_), .ZN(G225) );
  INV_X1 g572 ( .A(G225), .ZN(G308) );
  assign   G231 = 1'b0;
  BUF_X1 g573 ( .A(G452), .Z(G350) );
  BUF_X1 g574 ( .A(G452), .Z(G335) );
  BUF_X1 g575 ( .A(G452), .Z(G409) );
  BUF_X1 g576 ( .A(G1083), .Z(G369) );
  BUF_X1 g577 ( .A(G1083), .Z(G367) );
  BUF_X1 g578 ( .A(G2066), .Z(G411) );
  BUF_X1 g579 ( .A(G2066), .Z(G337) );
  BUF_X1 g580 ( .A(G2066), .Z(G384) );
  BUF_X1 g581 ( .A(G452), .Z(G391) );
  OR2_X1 g582 ( .A1(new_n529_), .A2(new_n528_), .ZN(G321) );
  AND2_X1 g583 ( .A1(new_n531_), .A2(new_n532_), .ZN(G280) );
  AND2_X1 g584 ( .A1(new_n538_), .A2(new_n540_), .ZN(G323) );
  OR2_X1 g585 ( .A1(new_n806_), .A2(new_n807_), .ZN(G331) );
endmodule


