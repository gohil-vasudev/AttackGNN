module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n716_, new_n153_, new_n701_, new_n257_, new_n481_, new_n212_, new_n449_, new_n580_, new_n639_, new_n484_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n150_, new_n683_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n310_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n605_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n163_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n119_, N75 );
nand g001 ( new_n120_, N29, N42 );
nor g002 ( N388, new_n120_, new_n119_ );
not g003 ( new_n122_, N80 );
nand g004 ( new_n123_, N29, N36 );
nor g005 ( N389, new_n123_, new_n122_ );
not g006 ( new_n125_, N42 );
nor g007 ( N390, new_n123_, new_n125_ );
nand g008 ( new_n127_, N85, N86 );
not g009 ( N391, new_n127_ );
not g010 ( new_n129_, N17 );
nand g011 ( new_n130_, N1, N8 );
not g012 ( new_n131_, new_n130_ );
nand g013 ( new_n132_, new_n131_, N13 );
nor g014 ( N418, new_n132_, new_n129_ );
not g015 ( new_n134_, N390 );
nand g016 ( new_n135_, N1, N26 );
nand g017 ( new_n136_, N13, N17 );
nor g018 ( new_n137_, new_n135_, new_n136_ );
nand g019 ( N419, new_n134_, new_n137_ );
nand g020 ( new_n139_, N59, N75 );
not g021 ( new_n140_, new_n139_ );
nand g022 ( N420, new_n140_, N80 );
nand g023 ( new_n142_, N36, N59 );
not g024 ( new_n143_, new_n142_ );
nand g025 ( N421, new_n143_, N80 );
nand g026 ( N422, new_n143_, N42 );
not g027 ( new_n146_, N90 );
nor g028 ( new_n147_, N87, N88 );
nor g029 ( N423, new_n147_, new_n146_ );
nand g030 ( N446, new_n137_, N390 );
not g031 ( new_n150_, new_n135_ );
nand g032 ( new_n151_, new_n150_, N51 );
nor g033 ( new_n152_, new_n151_, keyIn_0_0 );
not g034 ( new_n153_, keyIn_0_0 );
not g035 ( new_n154_, N51 );
nor g036 ( new_n155_, new_n135_, new_n154_ );
nor g037 ( new_n156_, new_n155_, new_n153_ );
nor g038 ( N447, new_n152_, new_n156_ );
not g039 ( new_n158_, new_n132_ );
nand g040 ( new_n159_, new_n158_, N55 );
nand g041 ( new_n160_, N29, N68 );
nor g042 ( N448, new_n159_, new_n160_ );
nand g043 ( new_n162_, N59, N68 );
not g044 ( new_n163_, new_n162_ );
nand g045 ( new_n164_, new_n163_, N74 );
nor g046 ( N449, new_n159_, new_n164_ );
not g047 ( new_n166_, N89 );
nor g048 ( N450, new_n147_, new_n166_ );
not g049 ( new_n168_, N130 );
nand g050 ( new_n169_, N91, N96 );
not g051 ( new_n170_, new_n169_ );
nor g052 ( new_n171_, N91, N96 );
nor g053 ( new_n172_, new_n170_, new_n171_ );
not g054 ( new_n173_, new_n172_ );
nand g055 ( new_n174_, N101, N106 );
not g056 ( new_n175_, new_n174_ );
nor g057 ( new_n176_, N101, N106 );
nor g058 ( new_n177_, new_n175_, new_n176_ );
not g059 ( new_n178_, new_n177_ );
nor g060 ( new_n179_, new_n173_, new_n178_ );
nor g061 ( new_n180_, new_n172_, new_n177_ );
nor g062 ( new_n181_, new_n179_, new_n180_ );
not g063 ( new_n182_, new_n181_ );
nand g064 ( new_n183_, new_n182_, new_n168_ );
not g065 ( new_n184_, new_n183_ );
nor g066 ( new_n185_, new_n182_, new_n168_ );
nor g067 ( new_n186_, new_n184_, new_n185_ );
not g068 ( new_n187_, new_n186_ );
not g069 ( new_n188_, N135 );
nand g070 ( new_n189_, N111, N116 );
not g071 ( new_n190_, new_n189_ );
nor g072 ( new_n191_, N111, N116 );
nor g073 ( new_n192_, new_n190_, new_n191_ );
not g074 ( new_n193_, new_n192_ );
nand g075 ( new_n194_, N121, N126 );
not g076 ( new_n195_, new_n194_ );
nor g077 ( new_n196_, N121, N126 );
nor g078 ( new_n197_, new_n195_, new_n196_ );
not g079 ( new_n198_, new_n197_ );
nor g080 ( new_n199_, new_n193_, new_n198_ );
nor g081 ( new_n200_, new_n192_, new_n197_ );
nor g082 ( new_n201_, new_n199_, new_n200_ );
not g083 ( new_n202_, new_n201_ );
nand g084 ( new_n203_, new_n202_, new_n188_ );
not g085 ( new_n204_, new_n203_ );
nor g086 ( new_n205_, new_n202_, new_n188_ );
nor g087 ( new_n206_, new_n204_, new_n205_ );
not g088 ( new_n207_, new_n206_ );
nor g089 ( new_n208_, new_n187_, new_n207_ );
nor g090 ( new_n209_, new_n186_, new_n206_ );
nor g091 ( N767, new_n208_, new_n209_ );
nand g092 ( new_n211_, N159, N165 );
not g093 ( new_n212_, new_n211_ );
nor g094 ( new_n213_, N159, N165 );
nor g095 ( new_n214_, new_n212_, new_n213_ );
not g096 ( new_n215_, new_n214_ );
nand g097 ( new_n216_, N171, N177 );
not g098 ( new_n217_, new_n216_ );
nor g099 ( new_n218_, N171, N177 );
nor g100 ( new_n219_, new_n217_, new_n218_ );
not g101 ( new_n220_, new_n219_ );
nor g102 ( new_n221_, new_n215_, new_n220_ );
nor g103 ( new_n222_, new_n214_, new_n219_ );
nor g104 ( new_n223_, new_n221_, new_n222_ );
not g105 ( new_n224_, new_n223_ );
nand g106 ( new_n225_, new_n224_, new_n168_ );
not g107 ( new_n226_, new_n225_ );
nor g108 ( new_n227_, new_n224_, new_n168_ );
nor g109 ( new_n228_, new_n226_, new_n227_ );
not g110 ( new_n229_, new_n228_ );
not g111 ( new_n230_, N207 );
nand g112 ( new_n231_, N183, N189 );
not g113 ( new_n232_, new_n231_ );
nor g114 ( new_n233_, N183, N189 );
nor g115 ( new_n234_, new_n232_, new_n233_ );
not g116 ( new_n235_, new_n234_ );
nand g117 ( new_n236_, N195, N201 );
not g118 ( new_n237_, new_n236_ );
nor g119 ( new_n238_, N195, N201 );
nor g120 ( new_n239_, new_n237_, new_n238_ );
not g121 ( new_n240_, new_n239_ );
nor g122 ( new_n241_, new_n235_, new_n240_ );
nor g123 ( new_n242_, new_n234_, new_n239_ );
nor g124 ( new_n243_, new_n241_, new_n242_ );
not g125 ( new_n244_, new_n243_ );
nand g126 ( new_n245_, new_n244_, new_n230_ );
not g127 ( new_n246_, new_n245_ );
nor g128 ( new_n247_, new_n244_, new_n230_ );
nor g129 ( new_n248_, new_n246_, new_n247_ );
not g130 ( new_n249_, new_n248_ );
nor g131 ( new_n250_, new_n229_, new_n249_ );
nor g132 ( new_n251_, new_n228_, new_n248_ );
nor g133 ( N768, new_n250_, new_n251_ );
not g134 ( new_n253_, keyIn_0_9 );
nor g135 ( new_n254_, N447, keyIn_0_4 );
not g136 ( new_n255_, keyIn_0_4 );
nand g137 ( new_n256_, new_n155_, new_n153_ );
nand g138 ( new_n257_, new_n151_, keyIn_0_0 );
nand g139 ( new_n258_, new_n257_, new_n256_ );
nor g140 ( new_n259_, new_n258_, new_n255_ );
nor g141 ( new_n260_, new_n254_, new_n259_ );
nand g142 ( new_n261_, new_n260_, keyIn_0_7 );
not g143 ( new_n262_, keyIn_0_7 );
nand g144 ( new_n263_, new_n258_, new_n255_ );
nand g145 ( new_n264_, N447, keyIn_0_4 );
nand g146 ( new_n265_, new_n264_, new_n263_ );
nand g147 ( new_n266_, new_n265_, new_n262_ );
nand g148 ( new_n267_, new_n261_, new_n266_ );
not g149 ( new_n268_, keyIn_0_6 );
nand g150 ( new_n269_, N17, N42 );
nand g151 ( new_n270_, new_n269_, keyIn_0_3 );
not g152 ( new_n271_, new_n270_ );
nor g153 ( new_n272_, new_n269_, keyIn_0_3 );
nor g154 ( new_n273_, new_n271_, new_n272_ );
nor g155 ( new_n274_, N17, N42 );
nor g156 ( new_n275_, new_n274_, keyIn_0_2 );
nand g157 ( new_n276_, new_n274_, keyIn_0_2 );
not g158 ( new_n277_, new_n276_ );
nor g159 ( new_n278_, new_n277_, new_n275_ );
nand g160 ( new_n279_, new_n278_, new_n273_ );
nor g161 ( new_n280_, new_n279_, new_n268_ );
nand g162 ( new_n281_, new_n279_, new_n268_ );
nand g163 ( new_n282_, N59, N156 );
not g164 ( new_n283_, new_n282_ );
nand g165 ( new_n284_, new_n281_, new_n283_ );
nor g166 ( new_n285_, new_n284_, new_n280_ );
nand g167 ( new_n286_, new_n267_, new_n285_ );
nand g168 ( new_n287_, new_n286_, new_n253_ );
not g169 ( new_n288_, new_n287_ );
nor g170 ( new_n289_, new_n286_, new_n253_ );
nor g171 ( new_n290_, new_n288_, new_n289_ );
not g172 ( new_n291_, keyIn_0_1 );
nand g173 ( new_n292_, N17, N51 );
nor g174 ( new_n293_, new_n130_, new_n292_ );
nor g175 ( new_n294_, new_n293_, new_n291_ );
nand g176 ( new_n295_, new_n293_, new_n291_ );
not g177 ( new_n296_, new_n295_ );
nor g178 ( new_n297_, new_n296_, new_n294_ );
not g179 ( new_n298_, new_n297_ );
nand g180 ( new_n299_, new_n298_, keyIn_0_5 );
nor g181 ( new_n300_, new_n298_, keyIn_0_5 );
nor g182 ( new_n301_, new_n139_, new_n125_ );
nor g183 ( new_n302_, new_n300_, new_n301_ );
nand g184 ( new_n303_, new_n302_, new_n299_ );
nor g185 ( new_n304_, new_n303_, keyIn_0_8 );
nand g186 ( new_n305_, new_n303_, keyIn_0_8 );
not g187 ( new_n306_, new_n305_ );
nor g188 ( new_n307_, new_n306_, new_n304_ );
nor g189 ( new_n308_, new_n290_, new_n307_ );
nand g190 ( new_n309_, new_n308_, keyIn_0_10 );
not g191 ( new_n310_, keyIn_0_10 );
not g192 ( new_n311_, new_n289_ );
nand g193 ( new_n312_, new_n311_, new_n287_ );
not g194 ( new_n313_, new_n307_ );
nand g195 ( new_n314_, new_n312_, new_n313_ );
nand g196 ( new_n315_, new_n314_, new_n310_ );
nand g197 ( new_n316_, new_n309_, new_n315_ );
nand g198 ( new_n317_, new_n316_, N126 );
not g199 ( new_n318_, N153 );
not g200 ( new_n319_, N1 );
nand g201 ( new_n320_, new_n267_, new_n282_ );
nor g202 ( new_n321_, new_n320_, new_n129_ );
nor g203 ( new_n322_, new_n321_, new_n319_ );
nor g204 ( new_n323_, new_n322_, new_n318_ );
nand g205 ( new_n324_, N29, N75 );
nor g206 ( new_n325_, new_n324_, new_n122_ );
nand g207 ( new_n326_, new_n267_, new_n325_ );
not g208 ( new_n327_, new_n326_ );
not g209 ( new_n328_, N55 );
nor g210 ( new_n329_, new_n328_, N268 );
nand g211 ( new_n330_, new_n327_, new_n329_ );
not g212 ( new_n331_, new_n330_ );
nor g213 ( new_n332_, new_n323_, new_n331_ );
nand g214 ( new_n333_, new_n317_, new_n332_ );
nand g215 ( new_n334_, new_n333_, N201 );
not g216 ( new_n335_, new_n334_ );
nor g217 ( new_n336_, new_n333_, N201 );
nor g218 ( new_n337_, new_n335_, new_n336_ );
nand g219 ( new_n338_, new_n337_, N261 );
not g220 ( new_n339_, N219 );
nor g221 ( new_n340_, new_n337_, N261 );
nor g222 ( new_n341_, new_n340_, new_n339_ );
nand g223 ( new_n342_, new_n341_, new_n338_ );
not g224 ( new_n343_, N228 );
not g225 ( new_n344_, new_n337_ );
nor g226 ( new_n345_, new_n344_, new_n343_ );
nand g227 ( new_n346_, new_n335_, N237 );
nand g228 ( new_n347_, new_n333_, N246 );
not g229 ( new_n348_, N73 );
nand g230 ( new_n349_, N42, N72 );
nor g231 ( new_n350_, new_n349_, new_n348_ );
nand g232 ( new_n351_, new_n350_, new_n163_ );
nor g233 ( new_n352_, new_n159_, new_n351_ );
nand g234 ( new_n353_, new_n352_, N201 );
nand g235 ( new_n354_, N255, N267 );
nand g236 ( new_n355_, N121, N210 );
nand g237 ( new_n356_, new_n354_, new_n355_ );
not g238 ( new_n357_, new_n356_ );
nand g239 ( new_n358_, new_n353_, new_n357_ );
not g240 ( new_n359_, new_n358_ );
nand g241 ( new_n360_, new_n347_, new_n359_ );
not g242 ( new_n361_, new_n360_ );
nand g243 ( new_n362_, new_n346_, new_n361_ );
nor g244 ( new_n363_, new_n345_, new_n362_ );
nand g245 ( N850, new_n342_, new_n363_ );
not g246 ( new_n365_, keyIn_0_14 );
not g247 ( new_n366_, keyIn_0_13 );
not g248 ( new_n367_, keyIn_0_11 );
nand g249 ( new_n368_, new_n316_, N111 );
nor g250 ( new_n369_, new_n368_, new_n367_ );
nand g251 ( new_n370_, new_n368_, new_n367_ );
not g252 ( new_n371_, new_n322_ );
nand g253 ( new_n372_, new_n371_, N143 );
nand g254 ( new_n373_, new_n370_, new_n372_ );
nor g255 ( new_n374_, new_n373_, new_n369_ );
nand g256 ( new_n375_, new_n374_, keyIn_0_12 );
not g257 ( new_n376_, new_n375_ );
not g258 ( new_n377_, keyIn_0_12 );
not g259 ( new_n378_, new_n369_ );
not g260 ( new_n379_, new_n373_ );
nand g261 ( new_n380_, new_n379_, new_n378_ );
nand g262 ( new_n381_, new_n380_, new_n377_ );
nand g263 ( new_n382_, new_n381_, new_n330_ );
nor g264 ( new_n383_, new_n382_, new_n376_ );
nand g265 ( new_n384_, new_n383_, new_n366_ );
nor g266 ( new_n385_, new_n374_, keyIn_0_12 );
nor g267 ( new_n386_, new_n385_, new_n331_ );
nand g268 ( new_n387_, new_n386_, new_n375_ );
nand g269 ( new_n388_, new_n387_, keyIn_0_13 );
nand g270 ( new_n389_, new_n384_, new_n388_ );
nand g271 ( new_n390_, new_n389_, N183 );
nand g272 ( new_n391_, new_n390_, new_n365_ );
not g273 ( new_n392_, new_n390_ );
nand g274 ( new_n393_, new_n392_, keyIn_0_14 );
nand g275 ( new_n394_, new_n393_, new_n391_ );
nor g276 ( new_n395_, new_n389_, N183 );
nand g277 ( new_n396_, new_n395_, keyIn_0_15 );
not g278 ( new_n397_, keyIn_0_15 );
not g279 ( new_n398_, N183 );
nor g280 ( new_n399_, new_n387_, keyIn_0_13 );
nor g281 ( new_n400_, new_n383_, new_n366_ );
nor g282 ( new_n401_, new_n400_, new_n399_ );
nand g283 ( new_n402_, new_n401_, new_n398_ );
nand g284 ( new_n403_, new_n402_, new_n397_ );
nand g285 ( new_n404_, new_n403_, new_n396_ );
nor g286 ( new_n405_, new_n394_, new_n404_ );
not g287 ( new_n406_, new_n405_ );
nand g288 ( new_n407_, new_n316_, N121 );
not g289 ( new_n408_, N149 );
nor g290 ( new_n409_, new_n322_, new_n408_ );
nor g291 ( new_n410_, new_n409_, new_n331_ );
nand g292 ( new_n411_, new_n407_, new_n410_ );
nor g293 ( new_n412_, new_n411_, N195 );
not g294 ( new_n413_, new_n412_ );
nor g295 ( new_n414_, new_n413_, keyIn_0_16 );
not g296 ( new_n415_, new_n414_ );
nand g297 ( new_n416_, new_n413_, keyIn_0_16 );
nand g298 ( new_n417_, new_n415_, new_n416_ );
nand g299 ( new_n418_, new_n316_, N116 );
not g300 ( new_n419_, N146 );
nor g301 ( new_n420_, new_n322_, new_n419_ );
nor g302 ( new_n421_, new_n420_, new_n331_ );
nand g303 ( new_n422_, new_n418_, new_n421_ );
nor g304 ( new_n423_, new_n422_, N189 );
not g305 ( new_n424_, new_n423_ );
nand g306 ( new_n425_, new_n417_, new_n424_ );
not g307 ( new_n426_, N261 );
nor g308 ( new_n427_, new_n336_, new_n426_ );
not g309 ( new_n428_, new_n427_ );
nor g310 ( new_n429_, new_n425_, new_n428_ );
nor g311 ( new_n430_, new_n429_, keyIn_0_18 );
not g312 ( new_n431_, keyIn_0_18 );
not g313 ( new_n432_, new_n416_ );
nor g314 ( new_n433_, new_n432_, new_n414_ );
nor g315 ( new_n434_, new_n433_, new_n423_ );
nand g316 ( new_n435_, new_n434_, new_n427_ );
nor g317 ( new_n436_, new_n435_, new_n431_ );
nor g318 ( new_n437_, new_n436_, new_n430_ );
nand g319 ( new_n438_, new_n434_, new_n335_ );
nand g320 ( new_n439_, new_n411_, N195 );
nor g321 ( new_n440_, new_n423_, new_n439_ );
nand g322 ( new_n441_, new_n422_, N189 );
not g323 ( new_n442_, new_n441_ );
nor g324 ( new_n443_, new_n440_, new_n442_ );
nand g325 ( new_n444_, new_n438_, new_n443_ );
nor g326 ( new_n445_, new_n437_, new_n444_ );
nand g327 ( new_n446_, new_n406_, new_n445_ );
nor g328 ( new_n447_, new_n406_, new_n445_ );
nor g329 ( new_n448_, new_n447_, new_n339_ );
nand g330 ( new_n449_, new_n448_, new_n446_ );
not g331 ( new_n450_, N237 );
not g332 ( new_n451_, keyIn_0_17 );
not g333 ( new_n452_, new_n391_ );
nor g334 ( new_n453_, new_n390_, new_n365_ );
nor g335 ( new_n454_, new_n452_, new_n453_ );
nand g336 ( new_n455_, new_n454_, new_n451_ );
nand g337 ( new_n456_, new_n394_, keyIn_0_17 );
nand g338 ( new_n457_, new_n455_, new_n456_ );
not g339 ( new_n458_, new_n457_ );
nor g340 ( new_n459_, new_n458_, new_n450_ );
nand g341 ( new_n460_, new_n405_, N228 );
nand g342 ( new_n461_, new_n389_, N246 );
nand g343 ( new_n462_, new_n352_, N183 );
nand g344 ( new_n463_, N106, N210 );
nand g345 ( new_n464_, new_n462_, new_n463_ );
not g346 ( new_n465_, new_n464_ );
nand g347 ( new_n466_, new_n461_, new_n465_ );
not g348 ( new_n467_, new_n466_ );
nand g349 ( new_n468_, new_n460_, new_n467_ );
nor g350 ( new_n469_, new_n459_, new_n468_ );
nand g351 ( N863, new_n449_, new_n469_ );
nor g352 ( new_n471_, new_n427_, new_n335_ );
not g353 ( new_n472_, new_n471_ );
nand g354 ( new_n473_, new_n417_, new_n472_ );
nand g355 ( new_n474_, new_n473_, new_n439_ );
nor g356 ( new_n475_, new_n442_, new_n423_ );
nand g357 ( new_n476_, new_n474_, new_n475_ );
nor g358 ( new_n477_, new_n474_, new_n475_ );
nor g359 ( new_n478_, new_n477_, new_n339_ );
nand g360 ( new_n479_, new_n478_, new_n476_ );
not g361 ( new_n480_, new_n475_ );
nor g362 ( new_n481_, new_n480_, new_n343_ );
nand g363 ( new_n482_, new_n442_, N237 );
nand g364 ( new_n483_, new_n422_, N246 );
nand g365 ( new_n484_, new_n352_, N189 );
nand g366 ( new_n485_, N255, N259 );
nand g367 ( new_n486_, N111, N210 );
nand g368 ( new_n487_, new_n485_, new_n486_ );
not g369 ( new_n488_, new_n487_ );
nand g370 ( new_n489_, new_n484_, new_n488_ );
not g371 ( new_n490_, new_n489_ );
nand g372 ( new_n491_, new_n483_, new_n490_ );
not g373 ( new_n492_, new_n491_ );
nand g374 ( new_n493_, new_n482_, new_n492_ );
nor g375 ( new_n494_, new_n481_, new_n493_ );
nand g376 ( N864, new_n479_, new_n494_ );
nand g377 ( new_n496_, new_n417_, new_n439_ );
nand g378 ( new_n497_, new_n496_, new_n471_ );
nor g379 ( new_n498_, new_n496_, new_n471_ );
nor g380 ( new_n499_, new_n498_, new_n339_ );
nand g381 ( new_n500_, new_n499_, new_n497_ );
nor g382 ( new_n501_, new_n496_, new_n343_ );
not g383 ( new_n502_, new_n439_ );
nand g384 ( new_n503_, new_n502_, N237 );
nand g385 ( new_n504_, new_n411_, N246 );
nand g386 ( new_n505_, new_n352_, N195 );
nand g387 ( new_n506_, N255, N260 );
nand g388 ( new_n507_, N116, N210 );
nand g389 ( new_n508_, new_n506_, new_n507_ );
not g390 ( new_n509_, new_n508_ );
nand g391 ( new_n510_, new_n505_, new_n509_ );
not g392 ( new_n511_, new_n510_ );
nand g393 ( new_n512_, new_n504_, new_n511_ );
not g394 ( new_n513_, new_n512_ );
nand g395 ( new_n514_, new_n503_, new_n513_ );
nor g396 ( new_n515_, new_n501_, new_n514_ );
nand g397 ( N865, new_n500_, new_n515_ );
not g398 ( new_n517_, keyIn_0_21 );
nor g399 ( new_n518_, new_n457_, new_n517_ );
not g400 ( new_n519_, new_n518_ );
nand g401 ( new_n520_, new_n457_, new_n517_ );
not g402 ( new_n521_, keyIn_0_22 );
nor g403 ( new_n522_, new_n402_, new_n397_ );
nor g404 ( new_n523_, new_n395_, keyIn_0_15 );
nor g405 ( new_n524_, new_n522_, new_n523_ );
not g406 ( new_n525_, new_n437_ );
not g407 ( new_n526_, new_n444_ );
nand g408 ( new_n527_, new_n525_, new_n526_ );
nand g409 ( new_n528_, new_n524_, new_n527_ );
nand g410 ( new_n529_, new_n528_, new_n521_ );
nor g411 ( new_n530_, new_n404_, new_n445_ );
nand g412 ( new_n531_, new_n530_, keyIn_0_22 );
nand g413 ( new_n532_, new_n529_, new_n531_ );
nand g414 ( new_n533_, new_n520_, new_n532_ );
not g415 ( new_n534_, new_n533_ );
nand g416 ( new_n535_, new_n534_, new_n519_ );
nand g417 ( new_n536_, new_n535_, keyIn_0_23 );
not g418 ( new_n537_, keyIn_0_23 );
nor g419 ( new_n538_, new_n533_, new_n518_ );
nand g420 ( new_n539_, new_n538_, new_n537_ );
nand g421 ( new_n540_, new_n536_, new_n539_ );
nand g422 ( new_n541_, new_n316_, N106 );
not g423 ( new_n542_, new_n320_ );
nand g424 ( new_n543_, new_n542_, N55 );
nor g425 ( new_n544_, new_n543_, new_n318_ );
nor g426 ( new_n545_, new_n129_, N268 );
nand g427 ( new_n546_, new_n327_, new_n545_ );
nand g428 ( new_n547_, N138, N152 );
nand g429 ( new_n548_, new_n546_, new_n547_ );
nor g430 ( new_n549_, new_n544_, new_n548_ );
nand g431 ( new_n550_, new_n541_, new_n549_ );
nor g432 ( new_n551_, new_n550_, N177 );
not g433 ( new_n552_, new_n551_ );
nand g434 ( new_n553_, new_n540_, new_n552_ );
nand g435 ( new_n554_, new_n550_, N177 );
nand g436 ( new_n555_, new_n553_, new_n554_ );
nand g437 ( new_n556_, new_n316_, N101 );
nor g438 ( new_n557_, new_n543_, new_n408_ );
nand g439 ( new_n558_, N17, N138 );
nand g440 ( new_n559_, new_n546_, new_n558_ );
nor g441 ( new_n560_, new_n557_, new_n559_ );
nand g442 ( new_n561_, new_n556_, new_n560_ );
nor g443 ( new_n562_, new_n561_, N171 );
not g444 ( new_n563_, new_n562_ );
nand g445 ( new_n564_, new_n555_, new_n563_ );
nand g446 ( new_n565_, new_n561_, N171 );
nand g447 ( new_n566_, new_n564_, new_n565_ );
nand g448 ( new_n567_, new_n316_, N96 );
nor g449 ( new_n568_, new_n543_, new_n419_ );
nand g450 ( new_n569_, N51, N138 );
nand g451 ( new_n570_, new_n546_, new_n569_ );
nor g452 ( new_n571_, new_n568_, new_n570_ );
nand g453 ( new_n572_, new_n567_, new_n571_ );
nor g454 ( new_n573_, new_n572_, N165 );
not g455 ( new_n574_, new_n573_ );
nand g456 ( new_n575_, new_n566_, new_n574_ );
nand g457 ( new_n576_, new_n572_, N165 );
nand g458 ( new_n577_, new_n575_, new_n576_ );
nand g459 ( new_n578_, new_n316_, N91 );
not g460 ( new_n579_, N143 );
nor g461 ( new_n580_, new_n543_, new_n579_ );
nand g462 ( new_n581_, N8, N138 );
nand g463 ( new_n582_, new_n546_, new_n581_ );
nor g464 ( new_n583_, new_n580_, new_n582_ );
nand g465 ( new_n584_, new_n578_, new_n583_ );
nor g466 ( new_n585_, new_n584_, N159 );
not g467 ( new_n586_, new_n585_ );
nand g468 ( new_n587_, new_n577_, new_n586_ );
nand g469 ( new_n588_, new_n584_, N159 );
nand g470 ( N866, new_n587_, new_n588_ );
not g471 ( new_n590_, keyIn_0_29 );
not g472 ( new_n591_, new_n554_ );
nor g473 ( new_n592_, new_n591_, new_n551_ );
nand g474 ( new_n593_, new_n540_, new_n592_ );
nor g475 ( new_n594_, new_n593_, keyIn_0_25 );
nor g476 ( new_n595_, new_n540_, new_n592_ );
nand g477 ( new_n596_, new_n595_, keyIn_0_24 );
not g478 ( new_n597_, keyIn_0_24 );
nor g479 ( new_n598_, new_n538_, new_n537_ );
nor g480 ( new_n599_, new_n535_, keyIn_0_23 );
nor g481 ( new_n600_, new_n599_, new_n598_ );
not g482 ( new_n601_, new_n592_ );
nand g483 ( new_n602_, new_n600_, new_n601_ );
nand g484 ( new_n603_, new_n602_, new_n597_ );
nand g485 ( new_n604_, new_n603_, new_n596_ );
nor g486 ( new_n605_, new_n604_, new_n594_ );
nand g487 ( new_n606_, new_n593_, keyIn_0_25 );
nand g488 ( new_n607_, new_n605_, new_n606_ );
nand g489 ( new_n608_, new_n607_, keyIn_0_26 );
not g490 ( new_n609_, new_n594_ );
nor g491 ( new_n610_, new_n602_, new_n597_ );
nor g492 ( new_n611_, new_n595_, keyIn_0_24 );
nor g493 ( new_n612_, new_n610_, new_n611_ );
nand g494 ( new_n613_, new_n612_, new_n609_ );
not g495 ( new_n614_, keyIn_0_26 );
nand g496 ( new_n615_, new_n606_, new_n614_ );
nor g497 ( new_n616_, new_n613_, new_n615_ );
nor g498 ( new_n617_, new_n616_, new_n339_ );
nand g499 ( new_n618_, new_n617_, new_n608_ );
nor g500 ( new_n619_, new_n618_, keyIn_0_27 );
nand g501 ( new_n620_, new_n618_, keyIn_0_27 );
nand g502 ( new_n621_, N101, N210 );
nand g503 ( new_n622_, new_n620_, new_n621_ );
nor g504 ( new_n623_, new_n622_, new_n619_ );
nand g505 ( new_n624_, new_n623_, keyIn_0_28 );
not g506 ( new_n625_, new_n624_ );
not g507 ( new_n626_, keyIn_0_28 );
not g508 ( new_n627_, new_n619_ );
not g509 ( new_n628_, keyIn_0_27 );
not g510 ( new_n629_, new_n606_ );
nor g511 ( new_n630_, new_n613_, new_n629_ );
nor g512 ( new_n631_, new_n630_, new_n614_ );
not g513 ( new_n632_, new_n615_ );
nand g514 ( new_n633_, new_n605_, new_n632_ );
nand g515 ( new_n634_, new_n633_, N219 );
nor g516 ( new_n635_, new_n631_, new_n634_ );
nor g517 ( new_n636_, new_n635_, new_n628_ );
not g518 ( new_n637_, new_n621_ );
nor g519 ( new_n638_, new_n636_, new_n637_ );
nand g520 ( new_n639_, new_n638_, new_n627_ );
nand g521 ( new_n640_, new_n639_, new_n626_ );
nor g522 ( new_n641_, new_n601_, new_n343_ );
not g523 ( new_n642_, new_n641_ );
nor g524 ( new_n643_, new_n642_, keyIn_0_20 );
nand g525 ( new_n644_, new_n642_, keyIn_0_20 );
nor g526 ( new_n645_, new_n554_, new_n450_ );
nand g527 ( new_n646_, new_n550_, N246 );
nand g528 ( new_n647_, new_n352_, N177 );
nand g529 ( new_n648_, new_n646_, new_n647_ );
nor g530 ( new_n649_, new_n645_, new_n648_ );
nand g531 ( new_n650_, new_n644_, new_n649_ );
nor g532 ( new_n651_, new_n650_, new_n643_ );
nand g533 ( new_n652_, new_n640_, new_n651_ );
nor g534 ( new_n653_, new_n652_, new_n625_ );
nor g535 ( new_n654_, new_n653_, new_n590_ );
nor g536 ( new_n655_, new_n623_, keyIn_0_28 );
not g537 ( new_n656_, new_n651_ );
nor g538 ( new_n657_, new_n655_, new_n656_ );
nand g539 ( new_n658_, new_n657_, new_n624_ );
nor g540 ( new_n659_, new_n658_, keyIn_0_29 );
nor g541 ( new_n660_, new_n654_, new_n659_ );
nor g542 ( new_n661_, new_n660_, keyIn_0_30 );
not g543 ( new_n662_, keyIn_0_30 );
nand g544 ( new_n663_, new_n658_, keyIn_0_29 );
nand g545 ( new_n664_, new_n653_, new_n590_ );
nand g546 ( new_n665_, new_n664_, new_n663_ );
nor g547 ( new_n666_, new_n665_, new_n662_ );
nor g548 ( new_n667_, new_n661_, new_n666_ );
nor g549 ( new_n668_, new_n667_, keyIn_0_31 );
not g550 ( new_n669_, keyIn_0_31 );
nand g551 ( new_n670_, new_n665_, new_n662_ );
nand g552 ( new_n671_, new_n660_, keyIn_0_30 );
nand g553 ( new_n672_, new_n671_, new_n670_ );
nor g554 ( new_n673_, new_n672_, new_n669_ );
nor g555 ( N874, new_n668_, new_n673_ );
not g556 ( new_n675_, new_n588_ );
nor g557 ( new_n676_, new_n675_, new_n585_ );
nand g558 ( new_n677_, new_n577_, new_n676_ );
nor g559 ( new_n678_, new_n577_, new_n676_ );
nor g560 ( new_n679_, new_n678_, new_n339_ );
nand g561 ( new_n680_, new_n679_, new_n677_ );
not g562 ( new_n681_, new_n676_ );
nor g563 ( new_n682_, new_n681_, new_n343_ );
nand g564 ( new_n683_, new_n675_, N237 );
nand g565 ( new_n684_, new_n584_, N246 );
nand g566 ( new_n685_, new_n352_, N159 );
nand g567 ( new_n686_, N210, N268 );
nand g568 ( new_n687_, new_n685_, new_n686_ );
not g569 ( new_n688_, new_n687_ );
nand g570 ( new_n689_, new_n684_, new_n688_ );
not g571 ( new_n690_, new_n689_ );
nand g572 ( new_n691_, new_n683_, new_n690_ );
nor g573 ( new_n692_, new_n682_, new_n691_ );
nand g574 ( N878, new_n680_, new_n692_ );
not g575 ( new_n694_, new_n576_ );
nor g576 ( new_n695_, new_n694_, new_n573_ );
nand g577 ( new_n696_, new_n566_, new_n695_ );
nor g578 ( new_n697_, new_n566_, new_n695_ );
nor g579 ( new_n698_, new_n697_, new_n339_ );
nand g580 ( new_n699_, new_n698_, new_n696_ );
not g581 ( new_n700_, new_n695_ );
nor g582 ( new_n701_, new_n700_, new_n343_ );
nand g583 ( new_n702_, new_n694_, N237 );
nand g584 ( new_n703_, new_n572_, N246 );
nand g585 ( new_n704_, new_n352_, N165 );
nand g586 ( new_n705_, N91, N210 );
nand g587 ( new_n706_, new_n704_, new_n705_ );
not g588 ( new_n707_, new_n706_ );
nand g589 ( new_n708_, new_n703_, new_n707_ );
not g590 ( new_n709_, new_n708_ );
nand g591 ( new_n710_, new_n702_, new_n709_ );
nor g592 ( new_n711_, new_n701_, new_n710_ );
nand g593 ( N879, new_n699_, new_n711_ );
not g594 ( new_n713_, new_n565_ );
nor g595 ( new_n714_, new_n713_, new_n562_ );
nand g596 ( new_n715_, new_n555_, new_n714_ );
nor g597 ( new_n716_, new_n555_, new_n714_ );
nor g598 ( new_n717_, new_n716_, new_n339_ );
nand g599 ( new_n718_, new_n717_, new_n715_ );
not g600 ( new_n719_, keyIn_0_19 );
nor g601 ( new_n720_, new_n565_, new_n450_ );
not g602 ( new_n721_, new_n720_ );
nor g603 ( new_n722_, new_n721_, new_n719_ );
nor g604 ( new_n723_, new_n720_, keyIn_0_19 );
nor g605 ( new_n724_, new_n722_, new_n723_ );
nand g606 ( new_n725_, new_n714_, N228 );
nand g607 ( new_n726_, new_n561_, N246 );
nand g608 ( new_n727_, new_n352_, N171 );
nand g609 ( new_n728_, N96, N210 );
nand g610 ( new_n729_, new_n727_, new_n728_ );
not g611 ( new_n730_, new_n729_ );
nand g612 ( new_n731_, new_n726_, new_n730_ );
not g613 ( new_n732_, new_n731_ );
nand g614 ( new_n733_, new_n725_, new_n732_ );
nor g615 ( new_n734_, new_n724_, new_n733_ );
nand g616 ( N880, new_n718_, new_n734_ );
endmodule