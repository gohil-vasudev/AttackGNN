module top ( G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, keyinput0_G223gat, keyinput1_G223gat, keyinput2_G223gat, keyinput3_G223gat, keyinput0_G329gat, keyinput1_G329gat, keyinput2_G329gat, keyinput3_G329gat, keyinput0_G370gat, keyinput1_G370gat, keyinput2_G370gat, keyinput3_G370gat, keyinput0_G421gat, keyinput1_G421gat, keyinput2_G421gat, keyinput3_G421gat, keyinput0_G430gat, keyinput1_G430gat, keyinput2_G430gat, keyinput3_G430gat, keyinput0_G431gat, keyinput1_G431gat, keyinput2_G431gat, keyinput3_G431gat, keyinput0_G432gat, keyinput1_G432gat, keyinput2_G432gat, keyinput3_G432gat, G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat );
input G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat, G115gat, keyinput0_G223gat, keyinput1_G223gat, keyinput2_G223gat, keyinput3_G223gat, keyinput0_G329gat, keyinput1_G329gat, keyinput2_G329gat, keyinput3_G329gat, keyinput0_G370gat, keyinput1_G370gat, keyinput2_G370gat, keyinput3_G370gat, keyinput0_G421gat, keyinput1_G421gat, keyinput2_G421gat, keyinput3_G421gat, keyinput0_G430gat, keyinput1_G430gat, keyinput2_G430gat, keyinput3_G430gat, keyinput0_G431gat, keyinput1_G431gat, keyinput2_G431gat, keyinput3_G431gat, keyinput0_G432gat, keyinput1_G432gat, keyinput2_G432gat, keyinput3_G432gat;
output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
wire new_n1668_, new_n595_, new_n2051_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n1743_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1988_, new_n1433_, new_n2260_, new_n1517_, new_n1472_, new_n1785_, new_n439_, new_n1532_, new_n223_, new_n743_, new_n1962_, new_n1327_, new_n241_, new_n1535_, new_n2041_, new_n641_, new_n339_, new_n1849_, new_n389_, new_n514_, new_n2431_, new_n1351_, new_n636_, new_n691_, new_n1024_, new_n2291_, new_n911_, new_n679_, new_n937_, new_n1879_, new_n173_, new_n2054_, new_n728_, new_n1071_, new_n2114_, new_n1294_, new_n214_, new_n853_, new_n695_, new_n660_, new_n2038_, new_n1311_, new_n2424_, new_n552_, new_n342_, new_n1662_, new_n706_, new_n2132_, new_n2063_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n1769_, new_n317_, new_n2107_, new_n1188_, new_n2231_, new_n2264_, new_n2244_, new_n504_, new_n1414_, new_n234_, new_n873_, new_n1300_, new_n2135_, new_n1898_, new_n774_, new_n1777_, new_n2176_, new_n1620_, new_n1786_, new_n1946_, new_n1580_, new_n766_, new_n1973_, new_n2387_, new_n2421_, new_n1262_, new_n1212_, new_n2452_, new_n1332_, new_n1447_, new_n2293_, new_n685_, new_n326_, new_n2348_, new_n903_, new_n1595_, new_n822_, new_n1760_, new_n1018_, new_n1884_, new_n1864_, new_n1054_, new_n1288_, new_n385_, new_n1049_, new_n1330_, new_n2318_, new_n461_, new_n2171_, new_n2369_, new_n1323_, new_n297_, new_n150_, new_n1196_, new_n1366_, new_n137_, new_n2104_, new_n303_, new_n2334_, new_n2251_, new_n325_, new_n1285_, new_n1733_, new_n1842_, new_n1216_, new_n1632_, new_n1889_, new_n1987_, new_n629_, new_n2320_, new_n1214_, new_n883_, new_n1647_, new_n960_, new_n2433_, new_n1377_, new_n1522_, new_n549_, new_n2248_, new_n995_, new_n1035_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n2072_, new_n1678_, new_n568_, new_n1950_, new_n1936_, new_n423_, new_n496_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n85_, new_n912_, new_n1424_, new_n2350_, new_n680_, new_n981_, new_n2102_, new_n2337_, new_n1527_, new_n1275_, new_n1800_, new_n1198_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n2414_, new_n2397_, new_n194_, new_n2012_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n2184_, new_n142_, new_n2155_, new_n657_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n165_, new_n785_, new_n1501_, new_n477_, new_n664_, new_n280_, new_n1041_, new_n1989_, new_n426_, new_n1036_, new_n235_, new_n2142_, new_n1576_, new_n301_, new_n1718_, new_n169_, new_n1333_, new_n1132_, new_n395_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n1740_, new_n473_, new_n1624_, new_n1147_, new_n2217_, new_n1827_, new_n2401_, new_n1468_, new_n969_, new_n2332_, new_n1234_, new_n2343_, new_n1360_, new_n378_, new_n621_, new_n1637_, new_n244_, new_n943_, new_n1798_, new_n1321_, new_n1690_, new_n1209_, new_n1709_, new_n347_, new_n2084_, new_n2100_, new_n700_, new_n1419_, new_n921_, new_n396_, new_n1003_, new_n208_, new_n1671_, new_n1239_, new_n528_, new_n1667_, new_n2331_, new_n2213_, new_n2195_, new_n1218_, new_n1346_, new_n1201_, new_n1282_, new_n1630_, new_n2274_, new_n1349_, new_n2317_, new_n1547_, new_n1994_, new_n1437_, new_n2128_, new_n1598_, new_n1205_, new_n1966_, new_n1154_, new_n2411_, new_n295_, new_n1453_, new_n1850_, new_n2194_, new_n628_, new_n409_, new_n1090_, new_n1489_, new_n553_, new_n1061_, new_n2447_, new_n333_, new_n290_, new_n834_, new_n1991_, new_n1781_, new_n1738_, new_n1171_, new_n867_, new_n954_, new_n1591_, new_n1626_, new_n276_, new_n688_, new_n1704_, new_n410_, new_n1518_, new_n932_, new_n878_, new_n1981_, new_n509_, new_n1761_, new_n202_, new_n296_, new_n2187_, new_n1358_, new_n724_, new_n1070_, new_n1686_, new_n1416_, new_n156_, new_n261_, new_n672_, new_n1496_, new_n616_, new_n529_, new_n323_, new_n914_, new_n1875_, new_n362_, new_n1600_, new_n1631_, new_n2432_, new_n1771_, new_n460_, new_n1267_, new_n2237_, new_n1705_, new_n2090_, new_n1466_, new_n2370_, new_n1707_, new_n1716_, new_n1516_, new_n380_, new_n861_, new_n1564_, new_n1656_, new_n2149_, new_n1252_, new_n1993_, new_n2288_, new_n2371_, new_n352_, new_n1553_, new_n1593_, new_n944_, new_n1542_, new_n1064_, new_n1949_, new_n2280_, new_n2444_, new_n1480_, new_n1745_, new_n1860_, new_n2436_, new_n273_, new_n224_, new_n586_, new_n963_, new_n993_, new_n1357_, new_n102_, new_n143_, new_n1628_, new_n2441_, new_n403_, new_n868_, new_n1242_, new_n2190_, new_n149_, new_n1612_, new_n1343_, new_n936_, new_n1459_, new_n189_, new_n1438_, new_n106_, new_n1016_, new_n1904_, new_n1144_, new_n1465_, new_n182_, new_n666_, new_n1290_, new_n2065_, new_n2233_, new_n2277_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n1700_, new_n219_, new_n382_, new_n2232_, new_n239_, new_n718_, new_n1310_, new_n2239_, new_n88_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n2103_, new_n95_, new_n1635_, new_n1509_, new_n1559_, new_n2152_, new_n1789_, new_n2440_, new_n544_, new_n2172_, new_n1941_, new_n1324_, new_n1293_, new_n1336_, new_n345_, new_n2066_, new_n2427_, new_n499_, new_n131_, new_n533_, new_n2416_, new_n795_, new_n459_, new_n1441_, new_n1728_, new_n2363_, new_n2354_, new_n1510_, new_n1174_, new_n1655_, new_n80_, new_n613_, new_n1464_, new_n417_, new_n837_, new_n801_, new_n2039_, new_n2336_, new_n631_, new_n453_, new_n2430_, new_n1723_, new_n2126_, new_n519_, new_n148_, new_n2319_, new_n662_, new_n864_, new_n2322_, new_n440_, new_n2218_, new_n1826_, new_n2407_, new_n1765_, new_n974_, new_n1907_, new_n2118_, new_n1565_, new_n751_, new_n2289_, new_n2141_, new_n1038_, new_n372_, new_n1758_, new_n2211_, new_n852_, new_n1474_, new_n1328_, new_n1430_, new_n213_, new_n769_, new_n433_, new_n2096_, new_n1956_, new_n109_, new_n1450_, new_n992_, new_n1098_, new_n1729_, new_n2069_, new_n732_, new_n1832_, new_n689_, new_n933_, new_n1608_, new_n1492_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n1379_, new_n712_, new_n550_, new_n1068_, new_n269_, new_n2106_, new_n512_, new_n2375_, new_n2131_, new_n1673_, new_n1220_, new_n989_, new_n1741_, new_n1421_, new_n644_, new_n1856_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n2366_, new_n913_, new_n594_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n881_, new_n1268_, new_n2052_, new_n1381_, new_n1566_, new_n684_, new_n1274_, new_n1893_, new_n1665_, new_n1787_, new_n905_, new_n1539_, new_n1643_, new_n1958_, new_n962_, new_n2399_, new_n86_, new_n627_, new_n760_, new_n1391_, new_n1986_, new_n2408_, new_n1353_, new_n1033_, new_n2050_, new_n2180_, new_n2273_, new_n1153_, new_n320_, new_n984_, new_n1183_, new_n2133_, new_n2353_, new_n89_, new_n2376_, new_n1316_, new_n2391_, new_n1460_, new_n1878_, new_n1602_, new_n128_, new_n610_, new_n1369_, new_n159_, new_n1694_, new_n2226_, new_n1401_, new_n175_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n2446_, new_n171_, new_n1320_, new_n1861_, new_n434_, new_n200_, new_n2021_, new_n2279_, new_n581_, new_n329_, new_n2301_, new_n686_, new_n1567_, new_n168_, new_n1389_, new_n1400_, new_n757_, new_n793_, new_n406_, new_n1597_, new_n1089_, new_n1192_, new_n135_, new_n2347_, new_n405_, new_n2115_, new_n942_, new_n2382_, new_n614_, new_n895_, new_n976_, new_n1405_, new_n1249_, new_n1354_, new_n847_, new_n250_, new_n288_, new_n798_, new_n1926_, new_n1969_, new_n1948_, new_n753_, new_n2345_, new_n1361_, new_n941_, new_n2073_, new_n827_, new_n1356_, new_n1747_, new_n366_, new_n779_, new_n1025_, new_n365_, new_n1207_, new_n1799_, new_n601_, new_n1057_, new_n1644_, new_n1677_, new_n2266_, new_n812_, new_n266_, new_n542_, new_n548_, new_n1397_, new_n1313_, new_n1120_, new_n819_, new_n451_, new_n489_, new_n804_, new_n602_, new_n114_, new_n1060_, new_n1303_, new_n413_, new_n1906_, new_n1544_, new_n1382_, new_n1896_, new_n442_, new_n677_, new_n642_, new_n211_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n1814_, new_n735_, new_n2146_, new_n2202_, new_n1304_, new_n1537_, new_n1834_, new_n1108_, new_n2246_, new_n862_, new_n1606_, new_n532_, new_n2159_, new_n393_, new_n2110_, new_n1617_, new_n292_, new_n2258_, new_n215_, new_n1319_, new_n626_, new_n1473_, new_n959_, new_n990_, new_n1629_, new_n2426_, new_n1238_, new_n2062_, new_n133_, new_n2037_, new_n2250_, new_n1880_, new_n1162_, new_n1730_, new_n2018_, new_n212_, new_n2003_, new_n1278_, new_n902_, new_n2113_, new_n2144_, new_n2309_, new_n201_, new_n1996_, new_n414_, new_n2028_, new_n2364_, new_n2011_, new_n1482_, new_n554_, new_n2303_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n2094_, new_n2212_, new_n855_, new_n103_, new_n1037_, new_n2154_, new_n759_, new_n167_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n1858_, new_n478_, new_n1307_, new_n73_, new_n2339_, new_n1486_, new_n361_, new_n764_, new_n2349_, new_n2081_, new_n2007_, new_n1955_, new_n1683_, new_n510_, new_n966_, new_n351_, new_n1877_, new_n1292_, new_n2036_, new_n609_, new_n180_, new_n1759_, new_n961_, new_n530_, new_n890_, new_n1006_, new_n1836_, new_n1701_, new_n1905_, new_n811_, new_n1445_, new_n1902_, new_n956_, new_n486_, new_n970_, new_n1618_, new_n768_, new_n1691_, new_n773_, new_n1452_, new_n2121_, new_n1823_, new_n492_, new_n1200_, new_n650_, new_n750_, new_n254_, new_n355_, new_n432_, new_n925_, new_n2040_, new_n1940_, new_n778_, new_n2267_, new_n452_, new_n1483_, new_n2177_, new_n820_, new_n1386_, new_n508_, new_n1844_, new_n714_, new_n1748_, new_n116_, new_n1007_, new_n1613_, new_n882_, new_n2162_, new_n1557_, new_n1159_, new_n118_, new_n1584_, new_n1337_, new_n77_, new_n1348_, new_n1555_, new_n1636_, new_n1322_, new_n1751_, new_n1133_, new_n2164_, new_n1177_, new_n2197_, new_n646_, new_n538_, new_n1026_, new_n2019_, new_n541_, new_n1388_, new_n1550_, new_n2372_, new_n311_, new_n587_, new_n2010_, new_n2220_, new_n465_, new_n84_, new_n783_, new_n1380_, new_n2016_, new_n263_, new_n2080_, new_n1601_, new_n488_, new_n524_, new_n1725_, new_n1245_, new_n663_, new_n1499_, new_n2392_, new_n1791_, new_n2035_, new_n1908_, new_n1689_, new_n198_, new_n1857_, new_n1393_, new_n1335_, new_n1364_, new_n965_, new_n572_, new_n397_, new_n975_, new_n1199_, new_n399_, new_n1581_, new_n945_, new_n1882_, new_n1115_, new_n1846_, new_n1231_, new_n1055_, new_n2043_, new_n1431_, new_n923_, new_n1674_, new_n469_, new_n437_, new_n1633_, new_n2242_, new_n1607_, new_n2373_, new_n1924_, new_n2368_, new_n2188_, new_n457_, new_n1852_, new_n2170_, new_n1301_, new_n1999_, new_n1128_, new_n1002_, new_n1169_, new_n384_, new_n900_, new_n1722_, new_n1824_, new_n2316_, new_n1788_, new_n113_, new_n1648_, new_n2191_, new_n2418_, new_n775_, new_n454_, new_n1872_, new_n1124_, new_n1000_, new_n2225_, new_n1947_, new_n1273_, new_n1491_, new_n1554_, new_n176_, new_n1923_, new_n2013_, new_n291_, new_n309_, new_n1160_, new_n82_, new_n259_, new_n1536_, new_n2305_, new_n2381_, new_n227_, new_n2393_, new_n690_, new_n416_, new_n744_, new_n1175_, new_n2125_, new_n1136_, new_n1272_, new_n1287_, new_n1462_, new_n619_, new_n2410_, new_n1890_, new_n577_, new_n2179_, new_n376_, new_n1538_, new_n1579_, new_n2147_, new_n2310_, new_n2183_, new_n749_, new_n1091_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n2429_, new_n1776_, new_n1030_, new_n485_, new_n578_, new_n918_, new_n126_, new_n1586_, new_n1805_, new_n2380_, new_n2390_, new_n1572_, new_n665_, new_n800_, new_n1387_, new_n719_, new_n1178_, new_n270_, new_n570_, new_n893_, new_n520_, new_n1347_, new_n145_, new_n253_, new_n825_, new_n2312_, new_n1627_, new_n557_, new_n1642_, new_n1807_, new_n2281_, new_n1742_, new_n507_, new_n741_, new_n1699_, new_n1224_, new_n2008_, new_n748_, new_n2117_, new_n1137_, new_n1286_, new_n107_, new_n813_, new_n830_, new_n1107_, new_n730_, new_n1326_, new_n592_, new_n1820_, new_n231_, new_n1080_, new_n1279_, new_n522_, new_n588_, new_n916_, new_n199_, new_n675_, new_n1155_, new_n1186_, new_n1848_, new_n2448_, new_n225_, new_n2002_, new_n1863_, new_n1246_, new_n2119_, new_n387_, new_n112_, new_n2105_, new_n1951_, new_n121_, new_n949_, new_n2048_, new_n221_, new_n450_, new_n1394_, new_n2379_, new_n1179_, new_n298_, new_n184_, new_n1088_, new_n2394_, new_n2374_, new_n1756_, new_n2163_, new_n569_, new_n555_, new_n1139_, new_n1793_, new_n392_, new_n2404_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n147_, new_n692_, new_n502_, new_n1821_, new_n209_, new_n623_, new_n446_, new_n316_, new_n826_, new_n2079_, new_n1476_, new_n1854_, new_n332_, new_n972_, new_n1634_, new_n2285_, new_n2287_, new_n2413_, new_n2178_, new_n1916_, new_n2046_, new_n733_, new_n1983_, new_n122_, new_n1021_, new_n585_, new_n2076_, new_n2116_, new_n2189_, new_n1976_, new_n2307_, new_n242_, new_n503_, new_n2323_, new_n772_, new_n1244_, new_n307_, new_n1736_, new_n1181_, new_n1093_, new_n1451_, new_n2138_, new_n1097_, new_n1069_, new_n1164_, new_n1779_, new_n1869_, new_n2265_, new_n1891_, new_n1719_, new_n1830_, new_n1885_, new_n687_, new_n1029_, new_n1862_, new_n1654_, new_n1688_, new_n1963_, new_n217_, new_n788_, new_n1457_, new_n1204_, new_n1610_, new_n129_, new_n1112_, new_n1715_, new_n1156_, new_n1938_, new_n930_, new_n1475_, new_n1604_, new_n412_, new_n607_, new_n1731_, new_n645_, new_n1087_, new_n723_, new_n2326_, new_n2282_, new_n1933_, new_n1577_, new_n574_, new_n1548_, new_n1578_, new_n2204_, new_n2435_, new_n1661_, new_n1615_, new_n957_, new_n1047_, new_n75_, new_n787_, new_n336_, new_n2243_, new_n1399_, new_n1531_, new_n1927_, new_n294_, new_n1589_, new_n1792_, new_n1965_, new_n1173_, new_n704_, new_n2087_, new_n1809_, new_n2315_, new_n2443_, new_n1570_, new_n1811_, new_n2004_, new_n2130_, new_n1502_, new_n1778_, new_n2325_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n2186_, new_n1243_, new_n1077_, new_n2196_, new_n2067_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1506_, new_n1583_, new_n2085_, new_n228_, new_n1011_, new_n802_, new_n104_, new_n1236_, new_n1829_, new_n2150_, new_n947_, new_n1813_, new_n982_, new_n1449_, new_n1961_, new_n2346_, new_n279_, new_n455_, new_n1982_, new_n1569_, new_n120_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n1918_, new_n2222_, new_n1605_, new_n2097_, new_n1964_, new_n1314_, new_n2292_, new_n1359_, new_n1233_, new_n1839_, new_n2236_, new_n501_, new_n1157_, new_n2086_, new_n1575_, new_n1048_, new_n885_, new_n1808_, new_n283_, new_n390_, new_n1910_, new_n1922_, new_n566_, new_n186_, new_n386_, new_n767_, new_n401_, new_n2454_, new_n2173_, new_n556_, new_n1899_, new_n670_, new_n456_, new_n1125_, new_n1590_, new_n2095_, new_n246_, new_n1881_, new_n2127_, new_n667_, new_n367_, new_n2099_, new_n1237_, new_n2026_, new_n1837_, new_n1568_, new_n1479_, new_n2240_, new_n2321_, new_n894_, new_n2199_, new_n526_, new_n908_, new_n1886_, new_n2023_, new_n2192_, new_n678_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n2033_, new_n2045_, new_n2160_, new_n2328_, new_n2169_, new_n2283_, new_n1415_, new_n1390_, new_n721_, new_n742_, new_n892_, new_n1368_, new_n2384_, new_n472_, new_n1919_, new_n1985_, new_n1768_, new_n2111_, new_n1167_, new_n1530_, new_n2070_, new_n1490_, new_n2313_, new_n2278_, new_n792_, new_n953_, new_n257_, new_n2403_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n272_, new_n282_, new_n1059_, new_n634_, new_n192_, new_n1851_, new_n635_, new_n1774_, new_n110_, new_n2108_, new_n648_, new_n2450_, new_n164_, new_n1803_, new_n983_, new_n1406_, new_n1990_, new_n1082_, new_n2238_, new_n606_, new_n796_, new_n655_, new_n630_, new_n1717_, new_n1670_, new_n694_, new_n565_, new_n1979_, new_n1984_, new_n108_, new_n183_, new_n511_, new_n2359_, new_n1714_, new_n2034_, new_n2165_, new_n1640_, new_n1031_, new_n2405_, new_n1281_, new_n2129_, new_n1911_, new_n1005_, new_n999_, new_n321_, new_n1816_, new_n324_, new_n1713_, new_n491_, new_n676_, new_n2300_, new_n2112_, new_n271_, new_n674_, new_n274_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n1753_, new_n420_, new_n876_, new_n1894_, new_n1900_, new_n498_, new_n1217_, new_n2032_, new_n1463_, new_n429_, new_n2109_, new_n2122_, new_n1222_, new_n353_, new_n734_, new_n1062_, new_n506_, new_n872_, new_n1277_, new_n1428_, new_n1440_, new_n656_, new_n2311_, new_n394_, new_n935_, new_n1972_, new_n139_, new_n1150_, new_n1735_, new_n441_, new_n1752_, new_n600_, new_n1737_, new_n1930_, new_n1657_, new_n1797_, new_n1562_, new_n1939_, new_n1953_, new_n398_, new_n2434_, new_n383_, new_n207_, new_n267_, new_n2161_, new_n1395_, new_n1682_, new_n1795_, new_n1373_, new_n1229_, new_n1422_, new_n187_, new_n1523_, new_n1698_, new_n1679_, new_n334_, new_n331_, new_n835_, new_n1574_, new_n1614_, new_n2261_, new_n1423_, new_n1732_, new_n172_, new_n705_, new_n874_, new_n402_, new_n335_, new_n659_, new_n346_, new_n1954_, new_n1315_, new_n696_, new_n1868_, new_n1039_, new_n1507_, new_n1439_, new_n1658_, new_n1952_, new_n1365_, new_n952_, new_n1870_, new_n179_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1385_, new_n2185_, new_n559_, new_n762_, new_n2134_, new_n1193_, new_n1780_, new_n1187_, new_n1253_, new_n1546_, new_n1256_, new_n166_, new_n1513_, new_n162_, new_n1669_, new_n745_, new_n161_, new_n1114_, new_n1084_, new_n668_, new_n1573_, new_n2200_, new_n369_, new_n1693_, new_n1032_, new_n1545_, new_n901_, new_n1757_, new_n1255_, new_n2205_, new_n155_, new_n985_, new_n2074_, new_n1995_, new_n851_, new_n543_, new_n1943_, new_n1975_, new_n886_, new_n371_, new_n1712_, new_n2058_, new_n2075_, new_n2284_, new_n661_, new_n797_, new_n232_, new_n2145_, new_n76_, new_n1109_, new_n1269_, new_n1653_, new_n2453_, new_n884_, new_n938_, new_n1592_, new_n809_, new_n1142_, new_n1623_, new_n2439_, new_n604_, new_n1461_, new_n1104_, new_n1703_, new_n1511_, new_n571_, new_n1859_, new_n1504_, new_n758_, new_n1802_, new_n328_, new_n2168_, new_n2015_, new_n2327_, new_n130_, new_n2329_, new_n1794_, new_n268_, new_n2124_, new_n1299_, new_n1477_, new_n1079_, new_n144_, new_n2271_, new_n1804_, new_n931_, new_n575_, new_n1493_, new_n2438_, new_n2451_, new_n562_, new_n1929_, new_n2254_, new_n1638_, new_n1065_, new_n1118_, new_n177_, new_n1645_, new_n493_, new_n547_, new_n1934_, new_n264_, new_n379_, new_n1825_, new_n1481_, new_n1325_, new_n1625_, new_n1191_, new_n1931_, new_n824_, new_n2304_, new_n125_, new_n717_, new_n1455_, new_n475_, new_n2249_, new_n237_, new_n858_, new_n2306_, new_n1384_, new_n1434_, new_n411_, new_n673_, new_n1766_, new_n2025_, new_n2082_, new_n407_, new_n1897_, new_n81_, new_n1833_, new_n1692_, new_n1726_, new_n736_, new_n513_, new_n1903_, new_n558_, new_n313_, new_n1370_, new_n2093_, new_n2042_, new_n2415_, new_n1710_, new_n146_, new_n2047_, new_n2167_, new_n919_, new_n302_, new_n755_, new_n2017_, new_n1040_, new_n615_, new_n2298_, new_n722_, new_n856_, new_n415_, new_n537_, new_n2068_, new_n255_, new_n2437_, new_n1130_, new_n2064_, new_n2256_, new_n2360_, new_n1122_, new_n1185_, new_n1240_, new_n2031_, new_n354_, new_n968_, new_n2001_, new_n105_, new_n2419_, new_n2055_, new_n2215_, new_n1508_, new_n337_, new_n1195_, new_n658_, new_n591_, new_n1458_, new_n2091_, new_n163_, new_n1818_, new_n997_, new_n563_, new_n2209_, new_n910_, new_n1521_, new_n1334_, new_n2044_, new_n531_, new_n1675_, new_n2308_, new_n593_, new_n111_, new_n1543_, new_n252_, new_n1248_, new_n1812_, new_n2259_, new_n1978_, new_n2208_, new_n2206_, new_n1454_, new_n978_, new_n1308_, new_n408_, new_n470_, new_n134_, new_n1660_, new_n871_, new_n265_, new_n584_, new_n815_, new_n2223_, new_n1619_, new_n1425_, new_n1980_, new_n857_, new_n1828_, new_n2207_, new_n2272_, new_n1017_, new_n2203_, new_n2314_, new_n1853_, new_n101_, new_n2140_, new_n1471_, new_n1117_, new_n1594_, new_n836_, new_n1684_, new_n2148_, new_n2378_, new_n327_, new_n681_, new_n561_, new_n1427_, new_n2210_, new_n196_, new_n818_, new_n1815_, new_n1376_, new_n1876_, new_n2092_, new_n1534_, new_n640_, new_n2262_, new_n754_, new_n653_, new_n1659_, new_n377_, new_n1258_, new_n2247_, new_n375_, new_n1841_, new_n1724_, new_n1436_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n1339_, new_n1784_, new_n1970_, new_n780_, new_n245_, new_n643_, new_n1194_, new_n1338_, new_n91_, new_n1230_, new_n1027_, new_n348_, new_n2409_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1639_, new_n1165_, new_n1259_, new_n2297_, new_n1208_, new_n2299_, new_n185_, new_n2241_, new_n1942_, new_n373_, new_n1235_, new_n540_, new_n1149_, new_n1928_, new_n1066_, new_n422_, new_n1944_, new_n99_, new_n1664_, new_n249_, new_n284_, new_n119_, new_n293_, new_n934_, new_n1651_, new_n770_, new_n1225_, new_n521_, new_n2123_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n2333_, new_n2083_, new_n1616_, new_n1806_, new_n2352_, new_n958_, new_n699_, new_n236_, new_n74_, new_n955_, new_n1895_, new_n79_, new_n888_, new_n1505_, new_n1340_, new_n1180_, new_n817_, new_n720_, new_n1801_, new_n620_, new_n368_, new_n1410_, new_n738_, new_n2201_, new_n1363_, new_n2198_, new_n1317_, new_n2385_, new_n1232_, new_n859_, new_n197_, new_n1211_, new_n1412_, new_n1176_, new_n1374_, new_n2269_, new_n2417_, new_n842_, new_n1552_, new_n170_, new_n682_, new_n1075_, new_n1790_, new_n2030_, new_n1563_, new_n821_, new_n1937_, new_n669_, new_n220_, new_n1402_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n637_, new_n1603_, new_n1971_, new_n1342_, new_n424_, new_n2422_, new_n2182_, new_n1210_, new_n188_, new_n240_, new_n1843_, new_n1487_, new_n1646_, new_n123_, new_n127_, new_n1418_, new_n1871_, new_n761_, new_n2027_, new_n2428_, new_n2156_, new_n840_, new_n1283_, new_n1913_, new_n1873_, new_n898_, new_n1734_, new_n799_, new_n946_, new_n1764_, new_n344_, new_n287_, new_n1977_, new_n2362_, new_n2166_, new_n1901_, new_n1469_, new_n1749_, new_n1838_, new_n427_, new_n2449_, new_n1739_, new_n418_, new_n746_, new_n1221_, new_n1585_, new_n1587_, new_n1264_, new_n1680_, new_n152_, new_n2005_, new_n157_, new_n716_, new_n153_, new_n701_, new_n1676_, new_n1058_, new_n2365_, new_n364_, new_n832_, new_n1696_, new_n2193_, new_n1968_, new_n1101_, new_n1250_, new_n1681_, new_n315_, new_n124_, new_n1050_, new_n2455_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n2234_, new_n589_, new_n248_, new_n350_, new_n117_, new_n1083_, new_n2295_, new_n1297_, new_n2361_, new_n1959_, new_n1720_, new_n2330_, new_n2358_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n2151_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n1685_, new_n1721_, new_n1184_, new_n1960_, new_n1426_, new_n517_, new_n2077_, new_n1892_, new_n1992_, new_n318_, new_n622_, new_n1706_, new_n2006_, new_n702_, new_n2014_, new_n2230_, new_n833_, new_n1560_, new_n715_, new_n443_, new_n1086_, new_n158_, new_n763_, new_n1622_, new_n1138_, new_n466_, new_n262_, new_n1652_, new_n2356_, new_n2137_, new_n1847_, new_n2406_, new_n2057_, new_n218_, new_n1170_, new_n2276_, new_n845_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n2398_, new_n1540_, new_n1611_, new_n2143_, new_n205_, new_n1708_, new_n1533_, new_n141_, new_n1754_, new_n1750_, new_n1767_, new_n2235_, new_n887_, new_n926_, new_n2060_, new_n875_, new_n256_, new_n1226_, new_n1727_, new_n381_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n771_, new_n979_, new_n1819_, new_n1435_, new_n2342_, new_n1280_, new_n1241_, new_n1145_, new_n929_, new_n986_, new_n314_, new_n216_, new_n1782_, new_n917_, new_n2275_, new_n2071_, new_n1822_, new_n1887_, new_n210_, new_n447_, new_n2181_, new_n1967_, new_n140_, new_n790_, new_n1081_, new_n1247_, new_n1411_, new_n2000_, new_n739_, new_n2221_, new_n341_, new_n996_, new_n1318_, new_n2088_, new_n846_, new_n915_, new_n349_, new_n2294_, new_n848_, new_n277_, new_n1921_, new_n1772_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1711_, new_n1254_, new_n2216_, new_n438_, new_n1344_, new_n939_, new_n632_, new_n671_, new_n83_, new_n1514_, new_n2253_, new_n850_, new_n1202_, new_n436_, new_n1526_, new_n1446_, new_n2136_, new_n596_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1866_, new_n1383_, new_n948_, new_n1520_, new_n838_, new_n1609_, new_n2324_, new_n2377_, new_n1755_, new_n233_, new_n391_, new_n96_, new_n178_, new_n1085_, new_n2245_, new_n359_, new_n132_, new_n794_, new_n2098_, new_n1582_, new_n2056_, new_n2009_, new_n1702_, new_n1909_, new_n2153_, new_n1810_, new_n448_, new_n1932_, new_n1329_, new_n1161_, new_n2341_, new_n2383_, new_n2367_, new_n2395_, new_n92_, new_n1914_, new_n924_, new_n1867_, new_n97_, new_n1034_, new_n1957_, new_n1663_, new_n308_, new_n2214_, new_n633_, new_n784_, new_n2396_, new_n1396_, new_n258_, new_n860_, new_n306_, new_n494_, new_n2286_, new_n2219_, new_n1166_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n1920_, new_n1043_, new_n222_, new_n400_, new_n693_, new_n1485_, new_n505_, new_n471_, new_n967_, new_n374_, new_n1135_, new_n1289_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n2252_, new_n138_, new_n310_, new_n2389_, new_n2388_, new_n1331_, new_n1094_, new_n1621_, new_n839_, new_n2078_, new_n525_, new_n1695_, new_n2412_, new_n940_, new_n810_, new_n2400_, new_n808_, new_n2101_, new_n1284_, new_n907_, new_n897_, new_n1012_, new_n869_, new_n1775_, new_n1525_, new_n2120_, new_n598_, new_n2255_, new_n1935_, new_n1063_, new_n1001_, new_n1917_, new_n90_, new_n260_, new_n251_, new_n300_, new_n1503_, new_n806_, new_n2229_, new_n605_, new_n1074_, new_n2175_, new_n93_, new_n1551_, new_n2423_, new_n480_, new_n625_, new_n1141_, new_n1650_, new_n807_, new_n151_, new_n726_, new_n1763_, new_n1263_, new_n1123_, new_n2020_, new_n2402_, new_n583_, new_n617_, new_n78_, new_n1467_, new_n1762_, new_n1997_, new_n781_, new_n1014_, new_n428_, new_n1855_, new_n487_, new_n360_, new_n98_, new_n2139_, new_n2302_, new_n1915_, new_n1596_, new_n191_, new_n1261_, new_n2445_, new_n2022_, new_n1488_, new_n2024_, new_n2224_, new_n922_, new_n2029_, new_n87_, new_n476_, new_n987_, new_n1641_, new_n2420_, new_n243_, new_n154_, new_n1148_, new_n1146_, new_n174_, new_n468_, new_n977_, new_n2049_, new_n782_, new_n444_, new_n518_, new_n1845_, new_n2174_, new_n285_, new_n1888_, new_n203_, new_n2089_, new_n590_, new_n2357_, new_n789_, new_n515_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n1835_, new_n2338_, new_n2425_, new_n1076_, new_n1350_, new_n160_, new_n312_, new_n535_, new_n725_, new_n100_, new_n814_, new_n527_, new_n115_, new_n1378_, new_n1945_, new_n190_, new_n1478_, new_n597_, new_n1092_, new_n1783_, new_n1143_, new_n1072_, new_n1190_, new_n2442_, new_n651_, new_n1296_, new_n1883_, new_n1309_, new_n1796_, new_n1010_, new_n776_, new_n2053_, new_n370_, new_n1649_, new_n1515_, new_n1746_, new_n638_, new_n523_, new_n909_, new_n1840_, new_n2296_, new_n1571_, new_n2386_, new_n1773_, new_n2351_, new_n1470_, new_n711_, new_n1298_, new_n731_, new_n599_, new_n2257_, new_n1260_, new_n973_, new_n1529_, new_n1541_, new_n1096_, new_n2344_, new_n1599_, new_n756_, new_n823_, new_n1549_, new_n2228_, new_n1500_, new_n928_, new_n319_, new_n1008_, new_n2059_, new_n1687_, new_n338_, new_n707_, new_n740_, new_n1134_, new_n1291_, new_n247_, new_n539_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1817_, new_n1672_, new_n2061_, new_n1295_, new_n1432_, new_n2158_, new_n1189_, new_n2268_, new_n2355_, new_n1197_, new_n1912_, new_n1312_, new_n1874_, new_n2340_, new_n467_, new_n404_, new_n193_, new_n2270_, new_n1666_, new_n1744_, new_n358_, new_n877_, new_n1697_, new_n545_, new_n611_, new_n1998_, new_n289_, new_n72_, new_n425_, new_n896_, new_n1831_, new_n1925_, new_n1770_, new_n866_, new_n1556_, new_n994_, new_n1494_, new_n2335_, new_n2157_, new_n964_, new_n1078_, new_n2227_, new_n136_, new_n551_, new_n1408_, new_n618_, new_n1140_, new_n2263_, new_n2290_, new_n464_, new_n1498_, new_n94_, new_n204_, new_n181_, new_n1588_, new_n1974_, new_n573_, new_n765_, new_n1103_;

not g0000 ( new_n72_, keyinput3_G223gat );
not g0001 ( new_n73_, keyinput2_G223gat );
not g0002 ( new_n74_, G99gat );
not g0003 ( new_n75_, G108gat );
or g0004 ( new_n76_, G112gat, G115gat );
and g0005 ( new_n77_, new_n76_, G102gat );
or g0006 ( new_n78_, new_n77_, new_n75_ );
and g0007 ( new_n79_, new_n78_, G105gat );
not g0008 ( new_n80_, G105gat );
or g0009 ( new_n81_, new_n75_, G102gat );
and g0010 ( new_n82_, new_n81_, new_n80_ );
or g0011 ( new_n83_, new_n79_, new_n82_ );
and g0012 ( new_n84_, new_n83_, new_n74_ );
and g0013 ( new_n85_, G102gat, G112gat );
not g0014 ( new_n86_, new_n85_ );
and g0015 ( new_n87_, new_n86_, G108gat );
not g0016 ( new_n88_, new_n87_ );
and g0017 ( new_n89_, new_n88_, G99gat );
and g0018 ( new_n90_, new_n89_, new_n80_ );
or g0019 ( new_n91_, new_n84_, new_n90_ );
and g0020 ( new_n92_, new_n91_, G89gat );
not g0021 ( new_n93_, G89gat );
and g0022 ( new_n94_, G112gat, G115gat );
or g0023 ( new_n95_, new_n81_, new_n94_ );
and g0024 ( new_n96_, new_n95_, G105gat );
or g0025 ( new_n97_, new_n81_, G112gat );
and g0026 ( new_n98_, new_n97_, new_n80_ );
or g0027 ( new_n99_, new_n96_, new_n98_ );
and g0028 ( new_n100_, new_n99_, G99gat );
not g0029 ( new_n101_, new_n76_ );
not g0030 ( new_n102_, new_n81_ );
and g0031 ( new_n103_, new_n102_, new_n101_ );
not g0032 ( new_n104_, new_n103_ );
or g0033 ( new_n105_, new_n104_, new_n80_ );
and g0034 ( new_n106_, new_n105_, new_n74_ );
or g0035 ( new_n107_, new_n100_, new_n106_ );
and g0036 ( new_n108_, new_n107_, new_n93_ );
or g0037 ( new_n109_, new_n92_, new_n108_ );
and g0038 ( new_n110_, new_n85_, G115gat );
or g0039 ( new_n111_, new_n110_, new_n75_ );
and g0040 ( new_n112_, new_n111_, G105gat );
and g0041 ( new_n113_, G89gat, G99gat );
and g0042 ( new_n114_, new_n112_, new_n113_ );
or g0043 ( new_n115_, new_n109_, new_n114_ );
and g0044 ( new_n116_, new_n115_, keyinput0_G223gat );
not g0045 ( new_n117_, keyinput0_G223gat );
and g0046 ( new_n118_, new_n89_, new_n117_ );
or g0047 ( new_n119_, new_n116_, new_n118_ );
and g0048 ( new_n120_, new_n119_, keyinput1_G223gat );
not g0049 ( new_n121_, keyinput1_G223gat );
not g0050 ( new_n122_, G115gat );
and g0051 ( new_n123_, new_n102_, new_n122_ );
or g0052 ( new_n124_, new_n98_, new_n123_ );
and g0053 ( new_n125_, new_n124_, G99gat );
or g0054 ( new_n126_, new_n103_, new_n80_ );
and g0055 ( new_n127_, new_n126_, new_n74_ );
or g0056 ( new_n128_, new_n125_, new_n127_ );
and g0057 ( new_n129_, new_n128_, new_n117_ );
and g0058 ( new_n130_, new_n126_, keyinput0_G223gat );
or g0059 ( new_n131_, new_n129_, new_n130_ );
and g0060 ( new_n132_, new_n131_, new_n121_ );
or g0061 ( new_n133_, new_n120_, new_n132_ );
and g0062 ( new_n134_, new_n133_, new_n73_ );
and g0063 ( new_n135_, new_n87_, new_n122_ );
or g0064 ( new_n136_, new_n135_, new_n80_ );
or g0065 ( new_n137_, new_n81_, new_n122_ );
and g0066 ( new_n138_, new_n136_, new_n137_ );
and g0067 ( new_n139_, new_n138_, new_n74_ );
or g0068 ( new_n140_, new_n88_, new_n122_ );
and g0069 ( new_n141_, new_n140_, G99gat );
and g0070 ( new_n142_, new_n122_, G108gat );
or g0071 ( new_n143_, new_n142_, new_n80_ );
and g0072 ( new_n144_, new_n141_, new_n143_ );
or g0073 ( new_n145_, new_n139_, new_n144_ );
and g0074 ( new_n146_, new_n145_, new_n117_ );
and g0075 ( new_n147_, new_n138_, keyinput0_G223gat );
or g0076 ( new_n148_, new_n146_, new_n147_ );
and g0077 ( new_n149_, new_n148_, new_n121_ );
not g0078 ( new_n150_, new_n97_ );
or g0079 ( new_n151_, new_n150_, new_n74_ );
and g0080 ( new_n152_, new_n151_, new_n93_ );
and g0081 ( new_n153_, new_n81_, new_n74_ );
not g0082 ( new_n154_, G112gat );
and g0083 ( new_n155_, new_n154_, G108gat );
or g0084 ( new_n156_, new_n153_, new_n155_ );
and g0085 ( new_n157_, new_n156_, G89gat );
or g0086 ( new_n158_, new_n152_, new_n157_ );
and g0087 ( new_n159_, new_n158_, keyinput0_G223gat );
not g0088 ( new_n160_, G95gat );
or g0089 ( new_n161_, new_n113_, new_n160_ );
and g0090 ( new_n162_, new_n88_, new_n161_ );
and g0091 ( new_n163_, new_n162_, new_n117_ );
or g0092 ( new_n164_, new_n159_, new_n163_ );
and g0093 ( new_n165_, new_n164_, keyinput1_G223gat );
or g0094 ( new_n166_, new_n149_, new_n165_ );
and g0095 ( new_n167_, new_n166_, keyinput2_G223gat );
or g0096 ( new_n168_, new_n134_, new_n167_ );
and g0097 ( new_n169_, new_n168_, new_n72_ );
and g0098 ( new_n170_, new_n93_, G95gat );
not g0099 ( new_n171_, new_n170_ );
and g0100 ( new_n172_, new_n171_, new_n81_ );
not g0101 ( new_n173_, G76gat );
and g0102 ( new_n174_, new_n173_, G82gat );
not g0103 ( new_n175_, new_n174_ );
and g0104 ( new_n176_, new_n172_, new_n175_ );
not g0105 ( new_n177_, G63gat );
and g0106 ( new_n178_, new_n177_, G69gat );
not g0107 ( new_n179_, new_n178_ );
and g0108 ( new_n180_, new_n176_, new_n179_ );
not g0109 ( new_n181_, G50gat );
and g0110 ( new_n182_, new_n181_, G56gat );
not g0111 ( new_n183_, new_n182_ );
and g0112 ( new_n184_, new_n180_, new_n183_ );
not g0113 ( new_n185_, G37gat );
and g0114 ( new_n186_, new_n185_, G43gat );
not g0115 ( new_n187_, new_n186_ );
and g0116 ( new_n188_, new_n184_, new_n187_ );
not g0117 ( new_n189_, G24gat );
and g0118 ( new_n190_, new_n189_, G30gat );
not g0119 ( new_n191_, new_n190_ );
and g0120 ( new_n192_, new_n188_, new_n191_ );
not g0121 ( new_n193_, G11gat );
and g0122 ( new_n194_, new_n193_, G17gat );
not g0123 ( new_n195_, new_n194_ );
not g0124 ( new_n196_, G4gat );
or g0125 ( new_n197_, new_n196_, G1gat );
and g0126 ( new_n198_, new_n195_, new_n197_ );
and g0127 ( new_n199_, new_n192_, new_n198_ );
not g0128 ( new_n200_, new_n199_ );
and g0129 ( new_n201_, new_n200_, keyinput0_G223gat );
and g0130 ( new_n202_, new_n117_, G108gat );
or g0131 ( new_n203_, new_n201_, new_n202_ );
and g0132 ( new_n204_, new_n203_, keyinput1_G223gat );
or g0133 ( new_n205_, new_n142_, new_n117_ );
not g0134 ( new_n206_, new_n202_ );
and g0135 ( new_n207_, new_n206_, new_n121_ );
and g0136 ( new_n208_, new_n207_, new_n205_ );
or g0137 ( new_n209_, new_n204_, new_n208_ );
and g0138 ( new_n210_, new_n209_, keyinput2_G223gat );
not g0139 ( new_n211_, new_n112_ );
and g0140 ( new_n212_, new_n211_, new_n117_ );
and g0141 ( new_n213_, new_n111_, keyinput0_G223gat );
or g0142 ( new_n214_, new_n212_, new_n213_ );
and g0143 ( new_n215_, new_n214_, keyinput1_G223gat );
and g0144 ( new_n216_, new_n113_, G105gat );
or g0145 ( new_n217_, new_n216_, new_n160_ );
and g0146 ( new_n218_, new_n111_, new_n217_ );
and g0147 ( new_n219_, new_n218_, keyinput0_G223gat );
or g0148 ( new_n220_, new_n219_, new_n118_ );
and g0149 ( new_n221_, new_n220_, new_n121_ );
or g0150 ( new_n222_, new_n215_, new_n221_ );
and g0151 ( new_n223_, new_n222_, new_n73_ );
or g0152 ( new_n224_, new_n210_, new_n223_ );
and g0153 ( new_n225_, new_n224_, keyinput3_G223gat );
or g0154 ( G223gat, new_n169_, new_n225_ );
not g0155 ( new_n227_, G86gat );
and g0156 ( new_n228_, new_n170_, new_n74_ );
not g0157 ( new_n229_, new_n228_ );
and g0158 ( new_n230_, new_n229_, new_n97_ );
not g0159 ( new_n231_, new_n230_ );
or g0160 ( new_n232_, new_n231_, new_n172_ );
and g0161 ( new_n233_, new_n232_, new_n227_ );
and g0162 ( new_n234_, G99gat, G102gat );
not g0163 ( new_n235_, new_n234_ );
or g0164 ( new_n236_, new_n171_, new_n235_ );
and g0165 ( new_n237_, G89gat, G112gat );
not g0166 ( new_n238_, new_n237_ );
or g0167 ( new_n239_, new_n81_, new_n238_ );
and g0168 ( new_n240_, new_n236_, new_n239_ );
and g0169 ( new_n241_, new_n74_, G95gat );
or g0170 ( new_n242_, new_n155_, new_n241_ );
and g0171 ( new_n243_, new_n242_, G86gat );
and g0172 ( new_n244_, new_n240_, new_n243_ );
or g0173 ( new_n245_, new_n233_, new_n244_ );
and g0174 ( new_n246_, new_n245_, G76gat );
or g0175 ( new_n247_, new_n231_, new_n227_ );
and g0176 ( new_n248_, new_n247_, new_n173_ );
or g0177 ( new_n249_, new_n246_, new_n248_ );
and g0178 ( new_n250_, new_n249_, G82gat );
not g0179 ( new_n251_, G82gat );
and g0180 ( new_n252_, new_n242_, new_n251_ );
and g0181 ( new_n253_, new_n240_, new_n252_ );
or g0182 ( new_n254_, new_n250_, new_n253_ );
and g0183 ( new_n255_, new_n254_, G73gat );
not g0184 ( new_n256_, G73gat );
and g0185 ( new_n257_, new_n174_, new_n227_ );
not g0186 ( new_n258_, new_n257_ );
and g0187 ( new_n259_, new_n230_, new_n258_ );
not g0188 ( new_n260_, new_n259_ );
or g0189 ( new_n261_, new_n260_, new_n176_ );
and g0190 ( new_n262_, new_n261_, new_n256_ );
or g0191 ( new_n263_, new_n255_, new_n262_ );
and g0192 ( new_n264_, new_n263_, G63gat );
not g0193 ( new_n265_, G69gat );
or g0194 ( new_n266_, new_n260_, new_n256_ );
and g0195 ( new_n267_, new_n266_, new_n177_ );
or g0196 ( new_n268_, new_n267_, new_n265_ );
or g0197 ( new_n269_, new_n264_, new_n268_ );
or g0198 ( new_n270_, new_n254_, G69gat );
and g0199 ( new_n271_, new_n269_, new_n270_ );
not g0200 ( new_n272_, G56gat );
and g0201 ( new_n273_, G50gat, G60gat );
or g0202 ( new_n274_, new_n273_, new_n272_ );
not g0203 ( new_n275_, new_n274_ );
or g0204 ( new_n276_, new_n271_, new_n275_ );
and g0205 ( new_n277_, new_n267_, G69gat );
and g0206 ( new_n278_, new_n261_, new_n179_ );
or g0207 ( new_n279_, new_n277_, new_n278_ );
or g0208 ( new_n280_, new_n279_, new_n181_ );
not g0209 ( new_n281_, G60gat );
and g0210 ( new_n282_, new_n178_, new_n256_ );
not g0211 ( new_n283_, new_n282_ );
and g0212 ( new_n284_, new_n259_, new_n283_ );
not g0213 ( new_n285_, new_n284_ );
or g0214 ( new_n286_, new_n285_, new_n281_ );
and g0215 ( new_n287_, new_n280_, new_n286_ );
or g0216 ( new_n288_, new_n287_, new_n274_ );
and g0217 ( new_n289_, new_n276_, new_n288_ );
not g0218 ( new_n290_, G43gat );
and g0219 ( new_n291_, G37gat, G47gat );
or g0220 ( new_n292_, new_n291_, new_n290_ );
not g0221 ( new_n293_, new_n292_ );
or g0222 ( new_n294_, new_n289_, new_n293_ );
or g0223 ( new_n295_, new_n279_, new_n182_ );
or g0224 ( new_n296_, new_n286_, new_n183_ );
and g0225 ( new_n297_, new_n295_, new_n296_ );
or g0226 ( new_n298_, new_n297_, new_n185_ );
and g0227 ( new_n299_, new_n182_, new_n281_ );
not g0228 ( new_n300_, new_n299_ );
and g0229 ( new_n301_, new_n284_, new_n300_ );
and g0230 ( new_n302_, new_n301_, G47gat );
not g0231 ( new_n303_, new_n302_ );
and g0232 ( new_n304_, new_n298_, new_n303_ );
or g0233 ( new_n305_, new_n304_, new_n292_ );
and g0234 ( new_n306_, new_n294_, new_n305_ );
not g0235 ( new_n307_, G30gat );
and g0236 ( new_n308_, G24gat, G34gat );
or g0237 ( new_n309_, new_n308_, new_n307_ );
not g0238 ( new_n310_, new_n309_ );
or g0239 ( new_n311_, new_n306_, new_n310_ );
or g0240 ( new_n312_, new_n297_, new_n186_ );
and g0241 ( new_n313_, new_n302_, new_n186_ );
not g0242 ( new_n314_, new_n313_ );
and g0243 ( new_n315_, new_n312_, new_n314_ );
not g0244 ( new_n316_, G34gat );
and g0245 ( new_n317_, new_n316_, G24gat );
not g0246 ( new_n318_, new_n317_ );
or g0247 ( new_n319_, new_n315_, new_n318_ );
not g0248 ( new_n320_, G47gat );
and g0249 ( new_n321_, new_n186_, new_n320_ );
not g0250 ( new_n322_, new_n321_ );
and g0251 ( new_n323_, new_n301_, new_n322_ );
and g0252 ( new_n324_, new_n189_, G34gat );
and g0253 ( new_n325_, new_n323_, new_n324_ );
not g0254 ( new_n326_, new_n325_ );
and g0255 ( new_n327_, new_n319_, new_n326_ );
or g0256 ( new_n328_, new_n327_, new_n307_ );
and g0257 ( new_n329_, G1gat, G8gat );
or g0258 ( new_n330_, new_n329_, new_n196_ );
not g0259 ( new_n331_, G17gat );
and g0260 ( new_n332_, G11gat, G21gat );
or g0261 ( new_n333_, new_n332_, new_n331_ );
and g0262 ( new_n334_, new_n330_, new_n333_ );
and g0263 ( new_n335_, new_n328_, new_n334_ );
and g0264 ( new_n336_, new_n311_, new_n335_ );
not g0265 ( new_n337_, G21gat );
or g0266 ( new_n338_, new_n315_, new_n190_ );
and g0267 ( new_n339_, new_n325_, G30gat );
not g0268 ( new_n340_, new_n339_ );
and g0269 ( new_n341_, new_n338_, new_n340_ );
and g0270 ( new_n342_, new_n341_, new_n337_ );
and g0271 ( new_n343_, new_n190_, new_n316_ );
not g0272 ( new_n344_, new_n343_ );
and g0273 ( new_n345_, new_n323_, new_n344_ );
and g0274 ( new_n346_, new_n345_, G21gat );
not g0275 ( new_n347_, new_n346_ );
and g0276 ( new_n348_, new_n347_, new_n193_ );
or g0277 ( new_n349_, new_n342_, new_n348_ );
and g0278 ( new_n350_, new_n197_, G17gat );
and g0279 ( new_n351_, new_n349_, new_n350_ );
not g0280 ( new_n352_, G8gat );
and g0281 ( new_n353_, new_n352_, G1gat );
and g0282 ( new_n354_, new_n195_, new_n353_ );
and g0283 ( new_n355_, new_n341_, new_n354_ );
not g0284 ( new_n356_, G1gat );
or g0285 ( new_n357_, new_n195_, G21gat );
and g0286 ( new_n358_, new_n357_, G8gat );
and g0287 ( new_n359_, new_n345_, new_n358_ );
not g0288 ( new_n360_, new_n359_ );
and g0289 ( new_n361_, new_n360_, new_n356_ );
or g0290 ( new_n362_, new_n355_, new_n361_ );
and g0291 ( new_n363_, new_n362_, G4gat );
or g0292 ( new_n364_, new_n351_, new_n363_ );
or g0293 ( new_n365_, new_n336_, new_n364_ );
and g0294 ( new_n366_, new_n365_, keyinput3_G329gat );
not g0295 ( new_n367_, keyinput3_G329gat );
and g0296 ( new_n368_, new_n87_, new_n367_ );
or g0297 ( new_n369_, new_n366_, new_n368_ );
and g0298 ( new_n370_, new_n369_, keyinput2_G329gat );
not g0299 ( new_n371_, keyinput2_G329gat );
or g0300 ( new_n372_, new_n80_, G115gat );
and g0301 ( new_n373_, new_n372_, new_n74_ );
or g0302 ( new_n374_, new_n373_, G112gat );
or g0303 ( new_n375_, new_n372_, new_n74_ );
and g0304 ( new_n376_, new_n374_, new_n375_ );
and g0305 ( new_n377_, new_n376_, new_n367_ );
or g0306 ( new_n378_, new_n377_, new_n81_ );
and g0307 ( new_n379_, new_n378_, new_n371_ );
or g0308 ( new_n380_, new_n370_, new_n379_ );
and g0309 ( new_n381_, new_n380_, keyinput1_G329gat );
or g0310 ( new_n382_, new_n170_, new_n174_ );
or g0311 ( new_n383_, new_n178_, new_n185_ );
or g0312 ( new_n384_, new_n383_, new_n182_ );
or g0313 ( new_n385_, new_n384_, new_n382_ );
and g0314 ( new_n386_, new_n385_, new_n367_ );
or g0315 ( new_n387_, new_n386_, new_n371_ );
or g0316 ( new_n388_, new_n382_, new_n367_ );
and g0317 ( new_n389_, new_n387_, new_n388_ );
or g0318 ( new_n390_, new_n389_, new_n102_ );
not g0319 ( new_n391_, keyinput1_G329gat );
and g0320 ( new_n392_, new_n74_, new_n80_ );
not g0321 ( new_n393_, new_n392_ );
and g0322 ( new_n394_, new_n393_, G89gat );
and g0323 ( new_n395_, new_n78_, new_n394_ );
or g0324 ( new_n396_, keyinput2_G329gat, keyinput3_G329gat );
or g0325 ( new_n397_, new_n395_, new_n396_ );
and g0326 ( new_n398_, new_n397_, new_n391_ );
and g0327 ( new_n399_, new_n390_, new_n398_ );
or g0328 ( new_n400_, new_n381_, new_n399_ );
and g0329 ( new_n401_, new_n400_, keyinput0_G329gat );
not g0330 ( new_n402_, keyinput0_G329gat );
and g0331 ( new_n403_, new_n93_, G102gat );
or g0332 ( new_n404_, new_n376_, new_n403_ );
or g0333 ( new_n405_, new_n93_, G102gat );
and g0334 ( new_n406_, new_n404_, new_n405_ );
or g0335 ( new_n407_, new_n406_, new_n75_ );
and g0336 ( new_n408_, new_n407_, new_n367_ );
and g0337 ( new_n409_, new_n211_, keyinput3_G329gat );
or g0338 ( new_n410_, new_n408_, new_n409_ );
and g0339 ( new_n411_, new_n410_, new_n371_ );
and g0340 ( new_n412_, new_n135_, new_n367_ );
and g0341 ( new_n413_, new_n75_, keyinput3_G329gat );
or g0342 ( new_n414_, new_n412_, new_n413_ );
and g0343 ( new_n415_, new_n414_, keyinput2_G329gat );
or g0344 ( new_n416_, new_n411_, new_n415_ );
and g0345 ( new_n417_, new_n416_, keyinput1_G329gat );
and g0346 ( new_n418_, new_n81_, G89gat );
and g0347 ( new_n419_, new_n93_, new_n74_ );
or g0348 ( new_n420_, new_n150_, new_n419_ );
or g0349 ( new_n421_, new_n420_, new_n418_ );
and g0350 ( new_n422_, new_n421_, new_n367_ );
not g0351 ( new_n423_, new_n418_ );
and g0352 ( new_n424_, new_n423_, keyinput3_G329gat );
or g0353 ( new_n425_, new_n422_, new_n424_ );
and g0354 ( new_n426_, new_n425_, keyinput2_G329gat );
and g0355 ( new_n427_, new_n124_, new_n367_ );
and g0356 ( new_n428_, new_n218_, keyinput3_G329gat );
or g0357 ( new_n429_, new_n427_, new_n428_ );
and g0358 ( new_n430_, new_n429_, new_n371_ );
or g0359 ( new_n431_, new_n426_, new_n430_ );
and g0360 ( new_n432_, new_n431_, new_n391_ );
or g0361 ( new_n433_, new_n417_, new_n432_ );
and g0362 ( new_n434_, new_n433_, new_n402_ );
or g0363 ( G329gat, new_n401_, new_n434_ );
and g0364 ( new_n436_, new_n145_, G89gat );
and g0365 ( new_n437_, new_n128_, new_n93_ );
or g0366 ( new_n438_, new_n436_, new_n437_ );
and g0367 ( new_n439_, new_n438_, G95gat );
and g0368 ( new_n440_, new_n142_, new_n160_ );
or g0369 ( new_n441_, new_n439_, new_n440_ );
and g0370 ( new_n442_, new_n441_, G92gat );
not g0371 ( new_n443_, G92gat );
or g0372 ( new_n444_, new_n139_, new_n141_ );
and g0373 ( new_n445_, new_n444_, G89gat );
or g0374 ( new_n446_, new_n445_, new_n437_ );
and g0375 ( new_n447_, new_n446_, G95gat );
and g0376 ( new_n448_, new_n140_, new_n160_ );
or g0377 ( new_n449_, new_n447_, new_n448_ );
and g0378 ( new_n450_, new_n449_, new_n443_ );
or g0379 ( new_n451_, new_n442_, new_n450_ );
and g0380 ( new_n452_, new_n451_, G86gat );
and g0381 ( new_n453_, new_n135_, G99gat );
or g0382 ( new_n454_, new_n139_, new_n453_ );
and g0383 ( new_n455_, new_n454_, G89gat );
or g0384 ( new_n456_, new_n455_, new_n437_ );
and g0385 ( new_n457_, new_n456_, G95gat );
and g0386 ( new_n458_, new_n440_, new_n86_ );
or g0387 ( new_n459_, new_n457_, new_n458_ );
and g0388 ( new_n460_, new_n459_, G92gat );
or g0389 ( new_n461_, new_n128_, new_n171_ );
or g0390 ( new_n462_, new_n137_, new_n170_ );
and g0391 ( new_n463_, new_n461_, new_n462_ );
and g0392 ( new_n464_, new_n463_, new_n443_ );
or g0393 ( new_n465_, new_n460_, new_n464_ );
and g0394 ( new_n466_, new_n465_, new_n227_ );
or g0395 ( new_n467_, new_n452_, new_n466_ );
and g0396 ( new_n468_, new_n467_, G76gat );
or g0397 ( new_n469_, new_n123_, new_n170_ );
and g0398 ( new_n470_, new_n461_, new_n469_ );
and g0399 ( new_n471_, new_n470_, G92gat );
or g0400 ( new_n472_, new_n126_, new_n229_ );
or g0401 ( new_n473_, new_n97_, new_n122_ );
or g0402 ( new_n474_, new_n473_, new_n228_ );
and g0403 ( new_n475_, new_n472_, new_n474_ );
and g0404 ( new_n476_, new_n475_, new_n443_ );
or g0405 ( new_n477_, new_n471_, new_n476_ );
and g0406 ( new_n478_, new_n477_, G86gat );
and g0407 ( new_n479_, new_n392_, new_n170_ );
or g0408 ( new_n480_, new_n103_, new_n479_ );
or g0409 ( new_n481_, new_n480_, new_n443_ );
and g0410 ( new_n482_, new_n481_, new_n227_ );
or g0411 ( new_n483_, new_n478_, new_n482_ );
and g0412 ( new_n484_, new_n483_, new_n173_ );
or g0413 ( new_n485_, new_n468_, new_n484_ );
and g0414 ( new_n486_, new_n485_, G82gat );
and g0415 ( new_n487_, new_n441_, new_n251_ );
or g0416 ( new_n488_, new_n486_, new_n487_ );
and g0417 ( new_n489_, new_n488_, G79gat );
not g0418 ( new_n490_, G79gat );
and g0419 ( new_n491_, new_n449_, G86gat );
or g0420 ( new_n492_, new_n466_, new_n491_ );
and g0421 ( new_n493_, new_n492_, G76gat );
or g0422 ( new_n494_, new_n493_, new_n484_ );
and g0423 ( new_n495_, new_n494_, G82gat );
and g0424 ( new_n496_, new_n449_, new_n251_ );
or g0425 ( new_n497_, new_n495_, new_n496_ );
and g0426 ( new_n498_, new_n497_, new_n490_ );
or g0427 ( new_n499_, new_n489_, new_n498_ );
and g0428 ( new_n500_, new_n499_, G73gat );
and g0429 ( new_n501_, new_n459_, G86gat );
or g0430 ( new_n502_, new_n466_, new_n501_ );
and g0431 ( new_n503_, new_n502_, G76gat );
or g0432 ( new_n504_, new_n503_, new_n484_ );
and g0433 ( new_n505_, new_n504_, G82gat );
and g0434 ( new_n506_, new_n459_, new_n251_ );
or g0435 ( new_n507_, new_n505_, new_n506_ );
and g0436 ( new_n508_, new_n507_, G79gat );
and g0437 ( new_n509_, new_n484_, G82gat );
and g0438 ( new_n510_, new_n463_, new_n175_ );
or g0439 ( new_n511_, new_n509_, new_n510_ );
and g0440 ( new_n512_, new_n511_, new_n490_ );
or g0441 ( new_n513_, new_n508_, new_n512_ );
and g0442 ( new_n514_, new_n513_, new_n256_ );
or g0443 ( new_n515_, new_n500_, new_n514_ );
and g0444 ( new_n516_, new_n515_, G63gat );
and g0445 ( new_n517_, new_n470_, new_n175_ );
or g0446 ( new_n518_, new_n509_, new_n517_ );
and g0447 ( new_n519_, new_n518_, G79gat );
or g0448 ( new_n520_, new_n475_, new_n257_ );
or g0449 ( new_n521_, new_n481_, new_n258_ );
and g0450 ( new_n522_, new_n520_, new_n521_ );
and g0451 ( new_n523_, new_n522_, new_n490_ );
or g0452 ( new_n524_, new_n519_, new_n523_ );
and g0453 ( new_n525_, new_n524_, G73gat );
not g0454 ( new_n526_, new_n480_ );
and g0455 ( new_n527_, new_n227_, new_n443_ );
and g0456 ( new_n528_, new_n527_, new_n174_ );
not g0457 ( new_n529_, new_n528_ );
and g0458 ( new_n530_, new_n526_, new_n529_ );
not g0459 ( new_n531_, new_n530_ );
or g0460 ( new_n532_, new_n531_, new_n490_ );
and g0461 ( new_n533_, new_n532_, new_n256_ );
or g0462 ( new_n534_, new_n525_, new_n533_ );
and g0463 ( new_n535_, new_n534_, new_n177_ );
or g0464 ( new_n536_, new_n516_, new_n535_ );
and g0465 ( new_n537_, new_n536_, G69gat );
and g0466 ( new_n538_, new_n488_, new_n265_ );
or g0467 ( new_n539_, new_n537_, new_n538_ );
and g0468 ( new_n540_, new_n539_, G66gat );
not g0469 ( new_n541_, G66gat );
and g0470 ( new_n542_, new_n497_, G73gat );
or g0471 ( new_n543_, new_n514_, new_n542_ );
and g0472 ( new_n544_, new_n543_, G63gat );
or g0473 ( new_n545_, new_n544_, new_n535_ );
and g0474 ( new_n546_, new_n545_, G69gat );
and g0475 ( new_n547_, new_n497_, new_n265_ );
or g0476 ( new_n548_, new_n546_, new_n547_ );
and g0477 ( new_n549_, new_n548_, new_n541_ );
or g0478 ( new_n550_, new_n540_, new_n549_ );
and g0479 ( new_n551_, new_n550_, G60gat );
and g0480 ( new_n552_, new_n507_, G73gat );
or g0481 ( new_n553_, new_n514_, new_n552_ );
and g0482 ( new_n554_, new_n553_, G63gat );
or g0483 ( new_n555_, new_n554_, new_n535_ );
and g0484 ( new_n556_, new_n555_, G69gat );
and g0485 ( new_n557_, new_n507_, new_n265_ );
or g0486 ( new_n558_, new_n556_, new_n557_ );
and g0487 ( new_n559_, new_n558_, G66gat );
and g0488 ( new_n560_, new_n535_, G69gat );
and g0489 ( new_n561_, new_n511_, new_n179_ );
or g0490 ( new_n562_, new_n560_, new_n561_ );
and g0491 ( new_n563_, new_n562_, new_n541_ );
or g0492 ( new_n564_, new_n559_, new_n563_ );
and g0493 ( new_n565_, new_n564_, new_n281_ );
or g0494 ( new_n566_, new_n551_, new_n565_ );
and g0495 ( new_n567_, new_n566_, G50gat );
and g0496 ( new_n568_, new_n518_, new_n179_ );
or g0497 ( new_n569_, new_n560_, new_n568_ );
and g0498 ( new_n570_, new_n569_, G66gat );
or g0499 ( new_n571_, new_n522_, new_n282_ );
or g0500 ( new_n572_, new_n532_, new_n283_ );
and g0501 ( new_n573_, new_n571_, new_n572_ );
and g0502 ( new_n574_, new_n573_, new_n541_ );
or g0503 ( new_n575_, new_n570_, new_n574_ );
and g0504 ( new_n576_, new_n575_, G60gat );
and g0505 ( new_n577_, new_n256_, new_n490_ );
and g0506 ( new_n578_, new_n577_, new_n178_ );
or g0507 ( new_n579_, new_n531_, new_n578_ );
or g0508 ( new_n580_, new_n579_, new_n541_ );
and g0509 ( new_n581_, new_n580_, new_n281_ );
or g0510 ( new_n582_, new_n576_, new_n581_ );
and g0511 ( new_n583_, new_n582_, new_n181_ );
or g0512 ( new_n584_, new_n567_, new_n583_ );
and g0513 ( new_n585_, new_n584_, G56gat );
and g0514 ( new_n586_, new_n539_, new_n272_ );
or g0515 ( new_n587_, new_n585_, new_n586_ );
and g0516 ( new_n588_, new_n587_, G53gat );
not g0517 ( new_n589_, G53gat );
and g0518 ( new_n590_, new_n548_, G60gat );
or g0519 ( new_n591_, new_n565_, new_n590_ );
and g0520 ( new_n592_, new_n591_, G50gat );
or g0521 ( new_n593_, new_n592_, new_n583_ );
and g0522 ( new_n594_, new_n593_, G56gat );
and g0523 ( new_n595_, new_n548_, new_n272_ );
or g0524 ( new_n596_, new_n594_, new_n595_ );
and g0525 ( new_n597_, new_n596_, new_n589_ );
or g0526 ( new_n598_, new_n588_, new_n597_ );
and g0527 ( new_n599_, new_n598_, G47gat );
and g0528 ( new_n600_, new_n558_, G60gat );
or g0529 ( new_n601_, new_n565_, new_n600_ );
and g0530 ( new_n602_, new_n601_, G50gat );
or g0531 ( new_n603_, new_n602_, new_n583_ );
and g0532 ( new_n604_, new_n603_, G56gat );
and g0533 ( new_n605_, new_n558_, new_n272_ );
or g0534 ( new_n606_, new_n604_, new_n605_ );
and g0535 ( new_n607_, new_n606_, G53gat );
and g0536 ( new_n608_, new_n583_, G56gat );
and g0537 ( new_n609_, new_n562_, new_n183_ );
or g0538 ( new_n610_, new_n608_, new_n609_ );
and g0539 ( new_n611_, new_n610_, new_n589_ );
or g0540 ( new_n612_, new_n607_, new_n611_ );
and g0541 ( new_n613_, new_n612_, new_n320_ );
or g0542 ( new_n614_, new_n599_, new_n613_ );
and g0543 ( new_n615_, new_n614_, G37gat );
and g0544 ( new_n616_, new_n569_, new_n183_ );
or g0545 ( new_n617_, new_n608_, new_n616_ );
and g0546 ( new_n618_, new_n617_, G53gat );
or g0547 ( new_n619_, new_n573_, new_n299_ );
or g0548 ( new_n620_, new_n580_, new_n300_ );
and g0549 ( new_n621_, new_n619_, new_n620_ );
and g0550 ( new_n622_, new_n621_, new_n589_ );
or g0551 ( new_n623_, new_n618_, new_n622_ );
and g0552 ( new_n624_, new_n623_, G47gat );
not g0553 ( new_n625_, new_n579_ );
and g0554 ( new_n626_, new_n299_, new_n541_ );
not g0555 ( new_n627_, new_n626_ );
and g0556 ( new_n628_, new_n625_, new_n627_ );
and g0557 ( new_n629_, new_n628_, G53gat );
not g0558 ( new_n630_, new_n629_ );
and g0559 ( new_n631_, new_n630_, new_n320_ );
or g0560 ( new_n632_, new_n624_, new_n631_ );
and g0561 ( new_n633_, new_n632_, new_n185_ );
or g0562 ( new_n634_, new_n615_, new_n633_ );
and g0563 ( new_n635_, new_n634_, G43gat );
and g0564 ( new_n636_, new_n587_, new_n290_ );
or g0565 ( new_n637_, new_n635_, new_n636_ );
and g0566 ( new_n638_, new_n637_, G40gat );
not g0567 ( new_n639_, G40gat );
and g0568 ( new_n640_, new_n596_, G47gat );
or g0569 ( new_n641_, new_n613_, new_n640_ );
and g0570 ( new_n642_, new_n641_, G37gat );
or g0571 ( new_n643_, new_n642_, new_n633_ );
and g0572 ( new_n644_, new_n643_, G43gat );
and g0573 ( new_n645_, new_n596_, new_n290_ );
or g0574 ( new_n646_, new_n644_, new_n645_ );
and g0575 ( new_n647_, new_n646_, new_n639_ );
or g0576 ( new_n648_, new_n638_, new_n647_ );
and g0577 ( new_n649_, new_n648_, G34gat );
and g0578 ( new_n650_, new_n606_, G47gat );
or g0579 ( new_n651_, new_n613_, new_n650_ );
and g0580 ( new_n652_, new_n651_, G37gat );
or g0581 ( new_n653_, new_n652_, new_n633_ );
and g0582 ( new_n654_, new_n653_, G43gat );
and g0583 ( new_n655_, new_n606_, new_n290_ );
or g0584 ( new_n656_, new_n654_, new_n655_ );
and g0585 ( new_n657_, new_n656_, G40gat );
and g0586 ( new_n658_, new_n633_, G43gat );
and g0587 ( new_n659_, new_n610_, new_n187_ );
or g0588 ( new_n660_, new_n658_, new_n659_ );
and g0589 ( new_n661_, new_n660_, new_n639_ );
or g0590 ( new_n662_, new_n657_, new_n661_ );
and g0591 ( new_n663_, new_n662_, new_n316_ );
or g0592 ( new_n664_, new_n649_, new_n663_ );
and g0593 ( new_n665_, new_n664_, G24gat );
and g0594 ( new_n666_, new_n617_, new_n187_ );
or g0595 ( new_n667_, new_n658_, new_n666_ );
and g0596 ( new_n668_, new_n667_, G40gat );
or g0597 ( new_n669_, new_n621_, new_n321_ );
and g0598 ( new_n670_, new_n629_, new_n321_ );
not g0599 ( new_n671_, new_n670_ );
and g0600 ( new_n672_, new_n669_, new_n671_ );
and g0601 ( new_n673_, new_n672_, new_n639_ );
or g0602 ( new_n674_, new_n668_, new_n673_ );
and g0603 ( new_n675_, new_n674_, G34gat );
and g0604 ( new_n676_, new_n320_, new_n589_ );
and g0605 ( new_n677_, new_n676_, new_n186_ );
not g0606 ( new_n678_, new_n677_ );
and g0607 ( new_n679_, new_n628_, new_n678_ );
and g0608 ( new_n680_, new_n679_, G40gat );
not g0609 ( new_n681_, new_n680_ );
and g0610 ( new_n682_, new_n681_, new_n316_ );
or g0611 ( new_n683_, new_n675_, new_n682_ );
and g0612 ( new_n684_, new_n683_, new_n189_ );
or g0613 ( new_n685_, new_n665_, new_n684_ );
and g0614 ( new_n686_, new_n685_, G30gat );
and g0615 ( new_n687_, new_n637_, new_n307_ );
or g0616 ( new_n688_, new_n686_, new_n687_ );
and g0617 ( new_n689_, new_n688_, G27gat );
not g0618 ( new_n690_, G27gat );
and g0619 ( new_n691_, new_n646_, G34gat );
or g0620 ( new_n692_, new_n663_, new_n691_ );
and g0621 ( new_n693_, new_n692_, G24gat );
or g0622 ( new_n694_, new_n693_, new_n684_ );
and g0623 ( new_n695_, new_n694_, G30gat );
and g0624 ( new_n696_, new_n646_, new_n307_ );
or g0625 ( new_n697_, new_n695_, new_n696_ );
and g0626 ( new_n698_, new_n697_, new_n690_ );
or g0627 ( new_n699_, new_n689_, new_n698_ );
and g0628 ( new_n700_, new_n699_, G14gat );
not g0629 ( new_n701_, G14gat );
and g0630 ( new_n702_, new_n697_, new_n701_ );
or g0631 ( new_n703_, new_n700_, new_n702_ );
and g0632 ( new_n704_, new_n703_, G21gat );
and g0633 ( new_n705_, new_n656_, G34gat );
or g0634 ( new_n706_, new_n663_, new_n705_ );
and g0635 ( new_n707_, new_n706_, G24gat );
or g0636 ( new_n708_, new_n707_, new_n684_ );
and g0637 ( new_n709_, new_n708_, G30gat );
and g0638 ( new_n710_, new_n656_, new_n307_ );
or g0639 ( new_n711_, new_n709_, new_n710_ );
and g0640 ( new_n712_, new_n711_, G27gat );
and g0641 ( new_n713_, new_n684_, G30gat );
and g0642 ( new_n714_, new_n660_, new_n191_ );
or g0643 ( new_n715_, new_n713_, new_n714_ );
and g0644 ( new_n716_, new_n715_, new_n690_ );
or g0645 ( new_n717_, new_n712_, new_n716_ );
and g0646 ( new_n718_, new_n717_, new_n337_ );
or g0647 ( new_n719_, new_n704_, new_n718_ );
and g0648 ( new_n720_, new_n719_, G8gat );
and g0649 ( new_n721_, new_n717_, G14gat );
and g0650 ( new_n722_, new_n715_, new_n701_ );
or g0651 ( new_n723_, new_n721_, new_n722_ );
and g0652 ( new_n724_, new_n723_, new_n337_ );
and g0653 ( new_n725_, new_n711_, G14gat );
or g0654 ( new_n726_, new_n725_, new_n722_ );
and g0655 ( new_n727_, new_n726_, G21gat );
or g0656 ( new_n728_, new_n724_, new_n727_ );
and g0657 ( new_n729_, new_n728_, new_n352_ );
or g0658 ( new_n730_, new_n720_, new_n729_ );
and g0659 ( new_n731_, new_n730_, G11gat );
and g0660 ( new_n732_, new_n667_, new_n191_ );
or g0661 ( new_n733_, new_n713_, new_n732_ );
and g0662 ( new_n734_, new_n733_, G27gat );
or g0663 ( new_n735_, new_n672_, new_n343_ );
and g0664 ( new_n736_, new_n680_, new_n343_ );
not g0665 ( new_n737_, new_n736_ );
and g0666 ( new_n738_, new_n735_, new_n737_ );
and g0667 ( new_n739_, new_n738_, new_n690_ );
or g0668 ( new_n740_, new_n734_, new_n739_ );
and g0669 ( new_n741_, new_n740_, G21gat );
and g0670 ( new_n742_, new_n316_, new_n639_ );
and g0671 ( new_n743_, new_n742_, new_n190_ );
not g0672 ( new_n744_, new_n743_ );
and g0673 ( new_n745_, new_n679_, new_n744_ );
and g0674 ( new_n746_, new_n745_, G27gat );
not g0675 ( new_n747_, new_n746_ );
and g0676 ( new_n748_, new_n747_, new_n337_ );
or g0677 ( new_n749_, new_n741_, new_n748_ );
and g0678 ( new_n750_, new_n749_, new_n193_ );
or g0679 ( new_n751_, new_n731_, new_n750_ );
and g0680 ( new_n752_, new_n751_, G17gat );
and g0681 ( new_n753_, new_n688_, G14gat );
or g0682 ( new_n754_, new_n753_, new_n702_ );
and g0683 ( new_n755_, new_n754_, G8gat );
and g0684 ( new_n756_, new_n726_, new_n352_ );
or g0685 ( new_n757_, new_n755_, new_n756_ );
and g0686 ( new_n758_, new_n757_, new_n331_ );
or g0687 ( new_n759_, new_n752_, new_n758_ );
and g0688 ( new_n760_, new_n759_, G1gat );
and g0689 ( new_n761_, G21gat, G27gat );
or g0690 ( new_n762_, new_n195_, new_n761_ );
and g0691 ( new_n763_, G8gat, G14gat );
and g0692 ( new_n764_, new_n762_, new_n763_ );
and g0693 ( new_n765_, new_n733_, new_n764_ );
and g0694 ( new_n766_, new_n739_, G8gat );
or g0695 ( new_n767_, new_n766_, new_n748_ );
and g0696 ( new_n768_, new_n767_, new_n194_ );
and g0697 ( new_n769_, new_n357_, new_n701_ );
and g0698 ( new_n770_, new_n738_, new_n769_ );
and g0699 ( new_n771_, new_n745_, G14gat );
not g0700 ( new_n772_, new_n771_ );
and g0701 ( new_n773_, new_n772_, new_n352_ );
or g0702 ( new_n774_, new_n770_, new_n773_ );
or g0703 ( new_n775_, new_n768_, new_n774_ );
or g0704 ( new_n776_, new_n765_, new_n775_ );
and g0705 ( new_n777_, new_n776_, new_n356_ );
or g0706 ( new_n778_, new_n760_, new_n777_ );
and g0707 ( new_n779_, new_n778_, G4gat );
and g0708 ( new_n780_, new_n699_, G21gat );
or g0709 ( new_n781_, new_n780_, new_n718_ );
and g0710 ( new_n782_, new_n781_, G11gat );
or g0711 ( new_n783_, new_n782_, new_n750_ );
and g0712 ( new_n784_, new_n783_, G17gat );
and g0713 ( new_n785_, new_n688_, new_n331_ );
or g0714 ( new_n786_, new_n784_, new_n785_ );
and g0715 ( new_n787_, new_n786_, new_n196_ );
or g0716 ( new_n788_, new_n779_, new_n787_ );
and g0717 ( new_n789_, new_n788_, keyinput0_G370gat );
not g0718 ( new_n790_, keyinput0_G370gat );
and g0719 ( new_n791_, new_n75_, new_n790_ );
or g0720 ( new_n792_, new_n789_, new_n791_ );
and g0721 ( new_n793_, new_n792_, keyinput1_G370gat );
not g0722 ( new_n794_, keyinput1_G370gat );
and g0723 ( new_n795_, new_n423_, new_n790_ );
and g0724 ( new_n796_, new_n102_, keyinput0_G370gat );
or g0725 ( new_n797_, new_n795_, new_n796_ );
and g0726 ( new_n798_, new_n797_, new_n794_ );
or g0727 ( new_n799_, new_n793_, new_n798_ );
and g0728 ( new_n800_, new_n799_, keyinput2_G370gat );
not g0729 ( new_n801_, keyinput2_G370gat );
and g0730 ( new_n802_, new_n114_, new_n790_ );
not g0731 ( new_n803_, new_n176_ );
and g0732 ( new_n804_, new_n803_, keyinput0_G370gat );
or g0733 ( new_n805_, new_n802_, new_n804_ );
and g0734 ( new_n806_, new_n805_, new_n794_ );
and g0735 ( new_n807_, new_n112_, new_n790_ );
not g0736 ( new_n808_, new_n807_ );
not g0737 ( new_n809_, new_n796_ );
and g0738 ( new_n810_, new_n809_, keyinput1_G370gat );
and g0739 ( new_n811_, new_n808_, new_n810_ );
or g0740 ( new_n812_, new_n806_, new_n811_ );
and g0741 ( new_n813_, new_n812_, new_n801_ );
or g0742 ( new_n814_, new_n800_, new_n813_ );
and g0743 ( new_n815_, new_n814_, keyinput3_G370gat );
not g0744 ( new_n816_, keyinput3_G370gat );
and g0745 ( new_n817_, new_n158_, G95gat );
and g0746 ( new_n818_, new_n155_, new_n160_ );
or g0747 ( new_n819_, new_n817_, new_n818_ );
and g0748 ( new_n820_, new_n819_, new_n790_ );
not g0749 ( new_n821_, new_n184_ );
and g0750 ( new_n822_, new_n821_, keyinput0_G370gat );
or g0751 ( new_n823_, new_n820_, new_n822_ );
and g0752 ( new_n824_, new_n823_, new_n794_ );
and g0753 ( new_n825_, new_n87_, new_n790_ );
or g0754 ( new_n826_, new_n825_, new_n796_ );
and g0755 ( new_n827_, new_n826_, keyinput1_G370gat );
or g0756 ( new_n828_, new_n824_, new_n827_ );
and g0757 ( new_n829_, new_n828_, keyinput2_G370gat );
and g0758 ( new_n830_, new_n79_, keyinput0_G370gat );
and g0759 ( new_n831_, new_n97_, new_n790_ );
or g0760 ( new_n832_, new_n830_, new_n831_ );
and g0761 ( new_n833_, new_n832_, new_n794_ );
and g0762 ( new_n834_, new_n80_, new_n790_ );
or g0763 ( new_n835_, new_n104_, new_n834_ );
and g0764 ( new_n836_, new_n835_, keyinput1_G370gat );
or g0765 ( new_n837_, new_n833_, new_n836_ );
and g0766 ( new_n838_, new_n837_, new_n801_ );
or g0767 ( new_n839_, new_n829_, new_n838_ );
and g0768 ( new_n840_, new_n839_, new_n816_ );
or g0769 ( G370gat, new_n815_, new_n840_ );
and g0770 ( new_n842_, G63gat, G73gat );
or g0771 ( new_n843_, new_n842_, new_n265_ );
and g0772 ( new_n844_, G76gat, G86gat );
or g0773 ( new_n845_, new_n844_, new_n251_ );
and g0774 ( new_n846_, new_n843_, new_n845_ );
and g0775 ( new_n847_, new_n162_, new_n846_ );
and g0776 ( new_n848_, new_n274_, new_n292_ );
and g0777 ( new_n849_, new_n848_, new_n309_ );
and g0778 ( new_n850_, new_n847_, new_n849_ );
or g0779 ( new_n851_, new_n850_, G14gat );
and g0780 ( new_n852_, G73gat, G79gat );
and g0781 ( new_n853_, new_n852_, G63gat );
or g0782 ( new_n854_, new_n853_, new_n265_ );
and g0783 ( new_n855_, new_n844_, G92gat );
or g0784 ( new_n856_, new_n855_, new_n251_ );
and g0785 ( new_n857_, new_n854_, new_n856_ );
and g0786 ( new_n858_, new_n218_, new_n857_ );
and g0787 ( new_n859_, new_n291_, G53gat );
or g0788 ( new_n860_, new_n859_, new_n290_ );
and g0789 ( new_n861_, new_n273_, G66gat );
or g0790 ( new_n862_, new_n861_, new_n272_ );
and g0791 ( new_n863_, new_n308_, G40gat );
or g0792 ( new_n864_, new_n863_, new_n307_ );
and g0793 ( new_n865_, new_n862_, new_n864_ );
and g0794 ( new_n866_, new_n865_, new_n860_ );
and g0795 ( new_n867_, new_n858_, new_n866_ );
or g0796 ( new_n868_, new_n867_, new_n701_ );
and g0797 ( new_n869_, new_n868_, new_n851_ );
and g0798 ( new_n870_, new_n690_, G14gat );
not g0799 ( new_n871_, new_n870_ );
and g0800 ( new_n872_, new_n869_, new_n871_ );
or g0801 ( new_n873_, new_n872_, new_n352_ );
or g0802 ( new_n874_, new_n192_, G14gat );
and g0803 ( new_n875_, new_n78_, new_n160_ );
or g0804 ( new_n876_, new_n395_, new_n875_ );
not g0805 ( new_n877_, new_n527_ );
and g0806 ( new_n878_, new_n877_, G76gat );
or g0807 ( new_n879_, new_n878_, new_n251_ );
not g0808 ( new_n880_, new_n577_ );
and g0809 ( new_n881_, new_n880_, G63gat );
or g0810 ( new_n882_, new_n881_, new_n265_ );
and g0811 ( new_n883_, new_n879_, new_n882_ );
and g0812 ( new_n884_, new_n876_, new_n883_ );
or g0813 ( new_n885_, new_n742_, new_n189_ );
and g0814 ( new_n886_, new_n885_, G30gat );
not g0815 ( new_n887_, new_n886_ );
and g0816 ( new_n888_, new_n281_, new_n541_ );
not g0817 ( new_n889_, new_n888_ );
and g0818 ( new_n890_, new_n889_, G50gat );
or g0819 ( new_n891_, new_n890_, new_n272_ );
not g0820 ( new_n892_, new_n676_ );
and g0821 ( new_n893_, new_n892_, G37gat );
or g0822 ( new_n894_, new_n893_, new_n290_ );
and g0823 ( new_n895_, new_n891_, new_n894_ );
and g0824 ( new_n896_, new_n895_, new_n887_ );
and g0825 ( new_n897_, new_n884_, new_n896_ );
or g0826 ( new_n898_, new_n897_, new_n701_ );
and g0827 ( new_n899_, new_n874_, new_n898_ );
or g0828 ( new_n900_, new_n899_, G8gat );
and g0829 ( new_n901_, new_n900_, G21gat );
and g0830 ( new_n902_, new_n901_, new_n873_ );
not g0831 ( new_n903_, new_n902_ );
and g0832 ( new_n904_, new_n897_, G27gat );
or g0833 ( new_n905_, new_n904_, new_n701_ );
and g0834 ( new_n906_, new_n352_, new_n337_ );
and g0835 ( new_n907_, new_n874_, new_n906_ );
and g0836 ( new_n908_, new_n907_, new_n905_ );
not g0837 ( new_n909_, new_n908_ );
and g0838 ( new_n910_, new_n903_, new_n909_ );
and g0839 ( new_n911_, G11gat, G17gat );
not g0840 ( new_n912_, new_n911_ );
or g0841 ( new_n913_, new_n910_, new_n912_ );
not g0842 ( new_n914_, new_n900_ );
not g0843 ( new_n915_, new_n869_ );
and g0844 ( new_n916_, new_n915_, G8gat );
or g0845 ( new_n917_, new_n916_, G17gat );
or g0846 ( new_n918_, new_n914_, new_n917_ );
and g0847 ( new_n919_, new_n913_, new_n918_ );
or g0848 ( new_n920_, new_n919_, new_n356_ );
not g0849 ( new_n921_, new_n345_ );
and g0850 ( new_n922_, new_n921_, G8gat );
or g0851 ( new_n923_, new_n922_, G14gat );
and g0852 ( new_n924_, new_n745_, new_n352_ );
not g0853 ( new_n925_, new_n924_ );
and g0854 ( new_n926_, G99gat, G105gat );
or g0855 ( new_n927_, new_n171_, new_n926_ );
not g0856 ( new_n928_, new_n927_ );
and g0857 ( new_n929_, G47gat, G53gat );
or g0858 ( new_n930_, new_n187_, new_n929_ );
not g0859 ( new_n931_, new_n930_ );
or g0860 ( new_n932_, new_n928_, new_n931_ );
and g0861 ( new_n933_, G60gat, G66gat );
or g0862 ( new_n934_, new_n183_, new_n933_ );
not g0863 ( new_n935_, new_n934_ );
and g0864 ( new_n936_, G34gat, G40gat );
or g0865 ( new_n937_, new_n191_, new_n936_ );
not g0866 ( new_n938_, new_n937_ );
or g0867 ( new_n939_, new_n935_, new_n938_ );
or g0868 ( new_n940_, new_n932_, new_n939_ );
and g0869 ( new_n941_, G86gat, G92gat );
or g0870 ( new_n942_, new_n175_, new_n941_ );
or g0871 ( new_n943_, new_n179_, new_n852_ );
and g0872 ( new_n944_, new_n942_, new_n943_ );
not g0873 ( new_n945_, new_n944_ );
not g0874 ( new_n946_, new_n95_ );
not g0875 ( new_n947_, new_n763_ );
or g0876 ( new_n948_, new_n946_, new_n947_ );
or g0877 ( new_n949_, new_n945_, new_n948_ );
or g0878 ( new_n950_, new_n940_, new_n949_ );
and g0879 ( new_n951_, new_n925_, new_n950_ );
and g0880 ( new_n952_, new_n951_, new_n923_ );
or g0881 ( new_n953_, new_n337_, G8gat );
and g0882 ( new_n954_, new_n953_, new_n870_ );
and g0883 ( new_n955_, new_n337_, G8gat );
or g0884 ( new_n956_, new_n954_, new_n955_ );
and g0885 ( new_n957_, new_n956_, new_n194_ );
or g0886 ( new_n958_, new_n957_, G1gat );
or g0887 ( new_n959_, new_n952_, new_n958_ );
and g0888 ( new_n960_, new_n959_, G4gat );
and g0889 ( new_n961_, new_n920_, new_n960_ );
or g0890 ( new_n962_, G69gat, G82gat );
or g0891 ( new_n963_, G95gat, G108gat );
or g0892 ( new_n964_, new_n962_, new_n963_ );
or g0893 ( new_n965_, G17gat, G30gat );
or g0894 ( new_n966_, G43gat, G56gat );
or g0895 ( new_n967_, new_n965_, new_n966_ );
or g0896 ( new_n968_, new_n964_, new_n967_ );
and g0897 ( new_n969_, new_n968_, new_n196_ );
or g0898 ( new_n970_, new_n961_, new_n969_ );
and g0899 ( new_n971_, new_n970_, keyinput3_G421gat );
not g0900 ( new_n972_, keyinput3_G421gat );
and g0901 ( new_n973_, new_n158_, new_n972_ );
or g0902 ( new_n974_, new_n971_, new_n973_ );
and g0903 ( new_n975_, new_n974_, keyinput2_G421gat );
not g0904 ( new_n976_, keyinput2_G421gat );
and g0905 ( new_n977_, new_n115_, new_n972_ );
and g0906 ( new_n978_, new_n111_, keyinput3_G421gat );
or g0907 ( new_n979_, new_n977_, new_n978_ );
and g0908 ( new_n980_, new_n979_, new_n976_ );
or g0909 ( new_n981_, new_n975_, new_n980_ );
and g0910 ( new_n982_, new_n981_, keyinput1_G421gat );
not g0911 ( new_n983_, keyinput1_G421gat );
and g0912 ( new_n984_, new_n138_, new_n972_ );
and g0913 ( new_n985_, new_n142_, keyinput3_G421gat );
or g0914 ( new_n986_, new_n984_, new_n985_ );
and g0915 ( new_n987_, new_n986_, keyinput2_G421gat );
and g0916 ( new_n988_, new_n218_, keyinput3_G421gat );
and g0917 ( new_n989_, new_n126_, new_n972_ );
or g0918 ( new_n990_, new_n988_, new_n989_ );
and g0919 ( new_n991_, new_n990_, new_n976_ );
or g0920 ( new_n992_, new_n987_, new_n991_ );
and g0921 ( new_n993_, new_n992_, new_n983_ );
or g0922 ( new_n994_, new_n982_, new_n993_ );
and g0923 ( new_n995_, new_n994_, keyinput0_G421gat );
not g0924 ( new_n996_, keyinput0_G421gat );
and g0925 ( new_n997_, new_n145_, new_n972_ );
and g0926 ( new_n998_, new_n75_, keyinput3_G421gat );
or g0927 ( new_n999_, new_n997_, new_n998_ );
and g0928 ( new_n1000_, new_n999_, keyinput2_G421gat );
and g0929 ( new_n1001_, new_n128_, new_n972_ );
and g0930 ( new_n1002_, new_n89_, keyinput3_G421gat );
or g0931 ( new_n1003_, new_n1001_, new_n1002_ );
and g0932 ( new_n1004_, new_n1003_, new_n976_ );
or g0933 ( new_n1005_, new_n1000_, new_n1004_ );
and g0934 ( new_n1006_, new_n1005_, new_n983_ );
and g0935 ( new_n1007_, new_n211_, keyinput3_G421gat );
and g0936 ( new_n1008_, new_n89_, new_n972_ );
or g0937 ( new_n1009_, new_n1007_, new_n1008_ );
and g0938 ( new_n1010_, new_n1009_, new_n976_ );
or g0939 ( new_n1011_, new_n162_, keyinput3_G421gat );
not g0940 ( new_n1012_, new_n998_ );
and g0941 ( new_n1013_, new_n1012_, keyinput2_G421gat );
and g0942 ( new_n1014_, new_n1011_, new_n1013_ );
or g0943 ( new_n1015_, new_n1010_, new_n1014_ );
and g0944 ( new_n1016_, new_n1015_, keyinput1_G421gat );
or g0945 ( new_n1017_, new_n1006_, new_n1016_ );
and g0946 ( new_n1018_, new_n1017_, new_n996_ );
or g0947 ( G421gat, new_n995_, new_n1018_ );
or g0948 ( new_n1020_, new_n625_, new_n541_ );
and g0949 ( new_n1021_, new_n1020_, new_n281_ );
and g0950 ( new_n1022_, new_n284_, new_n541_ );
or g0951 ( new_n1023_, new_n1021_, new_n1022_ );
and g0952 ( new_n1024_, new_n927_, new_n95_ );
and g0953 ( new_n1025_, new_n944_, new_n1024_ );
and g0954 ( new_n1026_, new_n1025_, new_n933_ );
or g0955 ( new_n1027_, new_n1023_, new_n1026_ );
and g0956 ( new_n1028_, new_n1027_, new_n181_ );
and g0957 ( new_n1029_, new_n884_, G66gat );
and g0958 ( new_n1030_, new_n180_, new_n541_ );
or g0959 ( new_n1031_, new_n1029_, new_n1030_ );
and g0960 ( new_n1032_, new_n1031_, new_n281_ );
and g0961 ( new_n1033_, new_n858_, G66gat );
and g0962 ( new_n1034_, new_n847_, new_n541_ );
or g0963 ( new_n1035_, new_n1033_, new_n1034_ );
and g0964 ( new_n1036_, new_n1035_, G60gat );
or g0965 ( new_n1037_, new_n1032_, new_n1036_ );
and g0966 ( new_n1038_, new_n1037_, G50gat );
or g0967 ( new_n1039_, new_n1028_, new_n1038_ );
and g0968 ( new_n1040_, new_n1039_, G56gat );
and g0969 ( new_n1041_, new_n858_, new_n272_ );
or g0970 ( new_n1042_, new_n1040_, new_n1041_ );
and g0971 ( new_n1043_, new_n1042_, G53gat );
and g0972 ( new_n1044_, new_n847_, G60gat );
or g0973 ( new_n1045_, new_n1032_, new_n1044_ );
and g0974 ( new_n1046_, new_n1045_, G50gat );
or g0975 ( new_n1047_, new_n1028_, new_n1046_ );
and g0976 ( new_n1048_, new_n1047_, G56gat );
and g0977 ( new_n1049_, new_n847_, new_n272_ );
or g0978 ( new_n1050_, new_n1048_, new_n1049_ );
and g0979 ( new_n1051_, new_n1050_, new_n589_ );
or g0980 ( new_n1052_, new_n1043_, new_n1051_ );
and g0981 ( new_n1053_, new_n1052_, G47gat );
and g0982 ( new_n1054_, new_n884_, G60gat );
or g0983 ( new_n1055_, new_n1032_, new_n1054_ );
and g0984 ( new_n1056_, new_n1055_, G50gat );
or g0985 ( new_n1057_, new_n1028_, new_n1056_ );
and g0986 ( new_n1058_, new_n1057_, G56gat );
and g0987 ( new_n1059_, new_n884_, new_n272_ );
or g0988 ( new_n1060_, new_n1058_, new_n1059_ );
or g0989 ( new_n1061_, new_n1060_, new_n589_ );
and g0990 ( new_n1062_, new_n1028_, G56gat );
or g0991 ( new_n1063_, new_n1062_, new_n184_ );
or g0992 ( new_n1064_, new_n1063_, G53gat );
and g0993 ( new_n1065_, new_n1064_, new_n320_ );
and g0994 ( new_n1066_, new_n1061_, new_n1065_ );
or g0995 ( new_n1067_, new_n1053_, new_n1066_ );
and g0996 ( new_n1068_, new_n1067_, G37gat );
and g0997 ( new_n1069_, new_n1025_, new_n183_ );
or g0998 ( new_n1070_, new_n1062_, new_n1069_ );
and g0999 ( new_n1071_, new_n1070_, G53gat );
and g1000 ( new_n1072_, new_n1020_, new_n299_ );
or g1001 ( new_n1073_, new_n1072_, new_n301_ );
and g1002 ( new_n1074_, new_n1073_, new_n589_ );
or g1003 ( new_n1075_, new_n1071_, new_n1074_ );
and g1004 ( new_n1076_, new_n1075_, G47gat );
and g1005 ( new_n1077_, new_n627_, G53gat );
not g1006 ( new_n1078_, new_n1077_ );
or g1007 ( new_n1079_, new_n625_, new_n1078_ );
and g1008 ( new_n1080_, new_n1079_, new_n320_ );
or g1009 ( new_n1081_, new_n1076_, new_n1080_ );
and g1010 ( new_n1082_, new_n1081_, new_n185_ );
or g1011 ( new_n1083_, new_n1068_, new_n1082_ );
and g1012 ( new_n1084_, new_n1083_, G43gat );
and g1013 ( new_n1085_, new_n1042_, new_n290_ );
or g1014 ( new_n1086_, new_n1084_, new_n1085_ );
and g1015 ( new_n1087_, new_n1086_, G40gat );
and g1016 ( new_n1088_, new_n1050_, G47gat );
or g1017 ( new_n1089_, new_n1066_, new_n1088_ );
and g1018 ( new_n1090_, new_n1089_, G37gat );
or g1019 ( new_n1091_, new_n1090_, new_n1082_ );
and g1020 ( new_n1092_, new_n1091_, G43gat );
and g1021 ( new_n1093_, new_n1050_, new_n290_ );
or g1022 ( new_n1094_, new_n1092_, new_n1093_ );
and g1023 ( new_n1095_, new_n1094_, new_n639_ );
or g1024 ( new_n1096_, new_n1087_, new_n1095_ );
and g1025 ( new_n1097_, new_n1096_, G34gat );
and g1026 ( new_n1098_, new_n1060_, G47gat );
or g1027 ( new_n1099_, new_n1066_, new_n1098_ );
and g1028 ( new_n1100_, new_n1099_, G37gat );
or g1029 ( new_n1101_, new_n1100_, new_n1082_ );
and g1030 ( new_n1102_, new_n1101_, G43gat );
and g1031 ( new_n1103_, new_n1060_, new_n290_ );
or g1032 ( new_n1104_, new_n1102_, new_n1103_ );
or g1033 ( new_n1105_, new_n1104_, new_n639_ );
and g1034 ( new_n1106_, new_n1082_, G43gat );
and g1035 ( new_n1107_, new_n1063_, new_n187_ );
or g1036 ( new_n1108_, new_n1106_, new_n1107_ );
or g1037 ( new_n1109_, new_n1108_, G40gat );
and g1038 ( new_n1110_, new_n1109_, new_n316_ );
and g1039 ( new_n1111_, new_n1105_, new_n1110_ );
or g1040 ( new_n1112_, new_n1097_, new_n1111_ );
and g1041 ( new_n1113_, new_n1112_, G24gat );
and g1042 ( new_n1114_, new_n1070_, new_n187_ );
or g1043 ( new_n1115_, new_n1106_, new_n1114_ );
and g1044 ( new_n1116_, new_n1115_, G40gat );
or g1045 ( new_n1117_, new_n1073_, new_n321_ );
or g1046 ( new_n1118_, new_n1079_, new_n322_ );
and g1047 ( new_n1119_, new_n1117_, new_n1118_ );
and g1048 ( new_n1120_, new_n1119_, new_n639_ );
or g1049 ( new_n1121_, new_n1116_, new_n1120_ );
and g1050 ( new_n1122_, new_n1121_, G34gat );
and g1051 ( new_n1123_, new_n627_, new_n678_ );
not g1052 ( new_n1124_, new_n1123_ );
or g1053 ( new_n1125_, new_n1124_, new_n639_ );
or g1054 ( new_n1126_, new_n625_, new_n1125_ );
and g1055 ( new_n1127_, new_n1126_, new_n316_ );
or g1056 ( new_n1128_, new_n1122_, new_n1127_ );
and g1057 ( new_n1129_, new_n1128_, new_n189_ );
or g1058 ( new_n1130_, new_n1113_, new_n1129_ );
and g1059 ( new_n1131_, new_n1130_, G30gat );
and g1060 ( new_n1132_, new_n1086_, new_n307_ );
or g1061 ( new_n1133_, new_n1131_, new_n1132_ );
and g1062 ( new_n1134_, new_n1133_, G14gat );
and g1063 ( new_n1135_, new_n1034_, G60gat );
or g1064 ( new_n1136_, new_n1032_, new_n1135_ );
and g1065 ( new_n1137_, new_n1136_, G50gat );
or g1066 ( new_n1138_, new_n1028_, new_n1137_ );
and g1067 ( new_n1139_, new_n1138_, G56gat );
and g1068 ( new_n1140_, new_n1139_, G53gat );
or g1069 ( new_n1141_, new_n1051_, new_n1140_ );
and g1070 ( new_n1142_, new_n1141_, G47gat );
or g1071 ( new_n1143_, new_n1142_, new_n1066_ );
and g1072 ( new_n1144_, new_n1143_, G37gat );
or g1073 ( new_n1145_, new_n1144_, new_n1082_ );
and g1074 ( new_n1146_, new_n1145_, G43gat );
and g1075 ( new_n1147_, new_n1139_, new_n290_ );
or g1076 ( new_n1148_, new_n1146_, new_n1147_ );
and g1077 ( new_n1149_, new_n1148_, G40gat );
or g1078 ( new_n1150_, new_n1149_, new_n1095_ );
and g1079 ( new_n1151_, new_n1150_, G34gat );
or g1080 ( new_n1152_, new_n1151_, new_n1111_ );
and g1081 ( new_n1153_, new_n1152_, G24gat );
or g1082 ( new_n1154_, new_n1153_, new_n1129_ );
and g1083 ( new_n1155_, new_n1154_, G30gat );
and g1084 ( new_n1156_, new_n1148_, new_n307_ );
or g1085 ( new_n1157_, new_n1155_, new_n1156_ );
and g1086 ( new_n1158_, new_n1157_, new_n701_ );
or g1087 ( new_n1159_, new_n1134_, new_n1158_ );
and g1088 ( new_n1160_, new_n1159_, G27gat );
and g1089 ( new_n1161_, new_n1111_, G24gat );
or g1090 ( new_n1162_, new_n1129_, new_n1161_ );
and g1091 ( new_n1163_, new_n1162_, G30gat );
and g1092 ( new_n1164_, new_n1094_, new_n309_ );
or g1093 ( new_n1165_, new_n1163_, new_n1164_ );
and g1094 ( new_n1166_, new_n1165_, new_n690_ );
or g1095 ( new_n1167_, new_n1160_, new_n1166_ );
and g1096 ( new_n1168_, new_n1167_, G21gat );
and g1097 ( new_n1169_, new_n1104_, G34gat );
or g1098 ( new_n1170_, new_n1111_, new_n1169_ );
and g1099 ( new_n1171_, new_n1170_, G24gat );
or g1100 ( new_n1172_, new_n1171_, new_n1129_ );
and g1101 ( new_n1173_, new_n1172_, G30gat );
and g1102 ( new_n1174_, new_n1104_, new_n307_ );
or g1103 ( new_n1175_, new_n1173_, new_n1174_ );
and g1104 ( new_n1176_, new_n1175_, G27gat );
and g1105 ( new_n1177_, new_n1129_, G30gat );
and g1106 ( new_n1178_, new_n1108_, new_n191_ );
or g1107 ( new_n1179_, new_n1177_, new_n1178_ );
and g1108 ( new_n1180_, new_n1179_, new_n690_ );
or g1109 ( new_n1181_, new_n1176_, new_n1180_ );
and g1110 ( new_n1182_, new_n1181_, new_n337_ );
or g1111 ( new_n1183_, new_n1168_, new_n1182_ );
and g1112 ( new_n1184_, new_n1183_, G8gat );
and g1113 ( new_n1185_, new_n1175_, G14gat );
and g1114 ( new_n1186_, new_n317_, new_n639_ );
and g1115 ( new_n1187_, new_n1108_, new_n1186_ );
or g1116 ( new_n1188_, new_n1129_, new_n1187_ );
and g1117 ( new_n1189_, new_n1188_, G30gat );
and g1118 ( new_n1190_, new_n676_, G37gat );
and g1119 ( new_n1191_, new_n1063_, new_n1190_ );
or g1120 ( new_n1192_, new_n1082_, new_n1191_ );
and g1121 ( new_n1193_, new_n1192_, G43gat );
and g1122 ( new_n1194_, new_n281_, G50gat );
and g1123 ( new_n1195_, new_n1030_, new_n1194_ );
or g1124 ( new_n1196_, new_n1028_, new_n1195_ );
and g1125 ( new_n1197_, new_n894_, G56gat );
and g1126 ( new_n1198_, new_n1196_, new_n1197_ );
or g1127 ( new_n1199_, new_n1193_, new_n1198_ );
and g1128 ( new_n1200_, new_n1199_, new_n887_ );
or g1129 ( new_n1201_, new_n1189_, new_n1200_ );
and g1130 ( new_n1202_, new_n1201_, new_n701_ );
or g1131 ( new_n1203_, new_n1185_, new_n1202_ );
and g1132 ( new_n1204_, new_n1203_, G27gat );
or g1133 ( new_n1205_, new_n1204_, new_n1180_ );
and g1134 ( new_n1206_, new_n1205_, new_n337_ );
and g1135 ( new_n1207_, new_n1032_, G50gat );
or g1136 ( new_n1208_, new_n1028_, new_n1207_ );
and g1137 ( new_n1209_, new_n1208_, G56gat );
and g1138 ( new_n1210_, new_n1209_, G47gat );
or g1139 ( new_n1211_, new_n1066_, new_n1210_ );
and g1140 ( new_n1212_, new_n1211_, G37gat );
or g1141 ( new_n1213_, new_n1212_, new_n1082_ );
and g1142 ( new_n1214_, new_n1213_, G43gat );
and g1143 ( new_n1215_, new_n1209_, new_n290_ );
or g1144 ( new_n1216_, new_n1214_, new_n1215_ );
and g1145 ( new_n1217_, new_n1216_, G34gat );
or g1146 ( new_n1218_, new_n1111_, new_n1217_ );
and g1147 ( new_n1219_, new_n1218_, G24gat );
or g1148 ( new_n1220_, new_n1219_, new_n1129_ );
and g1149 ( new_n1221_, new_n1220_, G30gat );
and g1150 ( new_n1222_, new_n1216_, new_n307_ );
or g1151 ( new_n1223_, new_n1221_, new_n1222_ );
and g1152 ( new_n1224_, new_n1223_, G14gat );
or g1153 ( new_n1225_, new_n1224_, new_n1202_ );
and g1154 ( new_n1226_, new_n1225_, G21gat );
or g1155 ( new_n1227_, new_n1206_, new_n1226_ );
and g1156 ( new_n1228_, new_n1227_, new_n352_ );
or g1157 ( new_n1229_, new_n1184_, new_n1228_ );
and g1158 ( new_n1230_, new_n1229_, G11gat );
and g1159 ( new_n1231_, new_n1115_, new_n191_ );
or g1160 ( new_n1232_, new_n1177_, new_n1231_ );
and g1161 ( new_n1233_, new_n1232_, G27gat );
or g1162 ( new_n1234_, new_n1119_, new_n343_ );
or g1163 ( new_n1235_, new_n1126_, new_n344_ );
and g1164 ( new_n1236_, new_n1235_, new_n690_ );
and g1165 ( new_n1237_, new_n1234_, new_n1236_ );
or g1166 ( new_n1238_, new_n1233_, new_n1237_ );
or g1167 ( new_n1239_, new_n1238_, new_n337_ );
or g1168 ( new_n1240_, new_n743_, new_n690_ );
or g1169 ( new_n1241_, new_n1124_, new_n1240_ );
or g1170 ( new_n1242_, new_n625_, G21gat );
or g1171 ( new_n1243_, new_n1242_, new_n1241_ );
and g1172 ( new_n1244_, new_n1243_, new_n193_ );
and g1173 ( new_n1245_, new_n1239_, new_n1244_ );
or g1174 ( new_n1246_, new_n1230_, new_n1245_ );
and g1175 ( new_n1247_, new_n1246_, G17gat );
and g1176 ( new_n1248_, new_n1040_, new_n290_ );
or g1177 ( new_n1249_, new_n1084_, new_n1248_ );
and g1178 ( new_n1250_, new_n1249_, new_n307_ );
or g1179 ( new_n1251_, new_n1131_, new_n1250_ );
and g1180 ( new_n1252_, new_n1251_, G14gat );
or g1181 ( new_n1253_, new_n1252_, new_n1158_ );
and g1182 ( new_n1254_, new_n1253_, G8gat );
and g1183 ( new_n1255_, new_n1225_, new_n352_ );
or g1184 ( new_n1256_, new_n1254_, new_n1255_ );
and g1185 ( new_n1257_, new_n1256_, new_n331_ );
or g1186 ( new_n1258_, new_n1247_, new_n1257_ );
and g1187 ( new_n1259_, new_n1258_, G1gat );
and g1188 ( new_n1260_, new_n1238_, G14gat );
and g1189 ( new_n1261_, new_n1023_, new_n182_ );
and g1190 ( new_n1262_, new_n1261_, G53gat );
or g1191 ( new_n1263_, new_n1262_, new_n1074_ );
and g1192 ( new_n1264_, new_n1263_, G47gat );
or g1193 ( new_n1265_, new_n1264_, new_n1080_ );
and g1194 ( new_n1266_, new_n1265_, new_n186_ );
and g1195 ( new_n1267_, new_n1261_, new_n187_ );
or g1196 ( new_n1268_, new_n1266_, new_n1267_ );
and g1197 ( new_n1269_, new_n1268_, new_n937_ );
and g1198 ( new_n1270_, new_n1120_, G34gat );
or g1199 ( new_n1271_, new_n1270_, new_n1127_ );
and g1200 ( new_n1272_, new_n1271_, new_n190_ );
or g1201 ( new_n1273_, new_n1269_, new_n1272_ );
and g1202 ( new_n1274_, new_n1273_, G27gat );
or g1203 ( new_n1275_, new_n1274_, new_n1237_ );
and g1204 ( new_n1276_, new_n1275_, new_n701_ );
or g1205 ( new_n1277_, new_n1276_, new_n337_ );
or g1206 ( new_n1278_, new_n1260_, new_n1277_ );
and g1207 ( new_n1279_, new_n1278_, new_n1243_ );
or g1208 ( new_n1280_, new_n1279_, new_n352_ );
or g1209 ( new_n1281_, new_n1072_, new_n321_ );
and g1210 ( new_n1282_, new_n1281_, new_n1118_ );
or g1211 ( new_n1283_, new_n1282_, new_n343_ );
and g1212 ( new_n1284_, new_n1283_, new_n1235_ );
or g1213 ( new_n1285_, new_n1284_, new_n701_ );
and g1214 ( new_n1286_, new_n744_, new_n701_ );
not g1215 ( new_n1287_, new_n1286_ );
or g1216 ( new_n1288_, new_n1124_, new_n1287_ );
and g1217 ( new_n1289_, new_n1285_, new_n1288_ );
and g1218 ( new_n1290_, new_n1289_, G21gat );
and g1219 ( new_n1291_, new_n625_, G14gat );
or g1220 ( new_n1292_, new_n1291_, new_n1241_ );
and g1221 ( new_n1293_, new_n1292_, new_n337_ );
or g1222 ( new_n1294_, new_n1293_, G8gat );
or g1223 ( new_n1295_, new_n1290_, new_n1294_ );
and g1224 ( new_n1296_, new_n1280_, new_n1295_ );
or g1225 ( new_n1297_, new_n1296_, new_n195_ );
and g1226 ( new_n1298_, new_n1062_, new_n187_ );
or g1227 ( new_n1299_, new_n1106_, new_n1298_ );
and g1228 ( new_n1300_, new_n1299_, new_n191_ );
or g1229 ( new_n1301_, new_n1177_, new_n1300_ );
and g1230 ( new_n1302_, new_n1301_, G14gat );
and g1231 ( new_n1303_, new_n1273_, new_n701_ );
or g1232 ( new_n1304_, new_n1303_, new_n352_ );
or g1233 ( new_n1305_, new_n1302_, new_n1304_ );
or g1234 ( new_n1306_, new_n1289_, G8gat );
and g1235 ( new_n1307_, new_n1305_, new_n1306_ );
or g1236 ( new_n1308_, new_n1307_, new_n194_ );
and g1237 ( new_n1309_, new_n1308_, new_n356_ );
and g1238 ( new_n1310_, new_n1297_, new_n1309_ );
or g1239 ( new_n1311_, new_n1259_, new_n1310_ );
and g1240 ( new_n1312_, new_n1311_, G4gat );
and g1241 ( new_n1313_, new_n1133_, G27gat );
or g1242 ( new_n1314_, new_n1313_, new_n1166_ );
and g1243 ( new_n1315_, new_n1314_, G21gat );
or g1244 ( new_n1316_, new_n1315_, new_n1182_ );
and g1245 ( new_n1317_, new_n1316_, G11gat );
or g1246 ( new_n1318_, new_n1317_, new_n1245_ );
and g1247 ( new_n1319_, new_n1318_, G17gat );
and g1248 ( new_n1320_, new_n1251_, new_n331_ );
or g1249 ( new_n1321_, new_n1319_, new_n1320_ );
and g1250 ( new_n1322_, new_n1321_, new_n196_ );
or g1251 ( new_n1323_, new_n1312_, new_n1322_ );
and g1252 ( new_n1324_, new_n1323_, keyinput0_G430gat );
not g1253 ( new_n1325_, keyinput0_G430gat );
and g1254 ( new_n1326_, new_n75_, new_n1325_ );
or g1255 ( new_n1327_, new_n1324_, new_n1326_ );
and g1256 ( new_n1328_, new_n1327_, keyinput1_G430gat );
not g1257 ( new_n1329_, keyinput1_G430gat );
and g1258 ( new_n1330_, new_n423_, new_n1325_ );
and g1259 ( new_n1331_, new_n102_, keyinput0_G430gat );
or g1260 ( new_n1332_, new_n1330_, new_n1331_ );
and g1261 ( new_n1333_, new_n1332_, new_n1329_ );
or g1262 ( new_n1334_, new_n1328_, new_n1333_ );
and g1263 ( new_n1335_, new_n1334_, keyinput2_G430gat );
not g1264 ( new_n1336_, keyinput2_G430gat );
and g1265 ( new_n1337_, new_n114_, new_n1325_ );
and g1266 ( new_n1338_, new_n803_, keyinput0_G430gat );
or g1267 ( new_n1339_, new_n1337_, new_n1338_ );
and g1268 ( new_n1340_, new_n1339_, new_n1329_ );
and g1269 ( new_n1341_, new_n112_, new_n1325_ );
not g1270 ( new_n1342_, new_n1341_ );
not g1271 ( new_n1343_, new_n1331_ );
and g1272 ( new_n1344_, new_n1343_, keyinput1_G430gat );
and g1273 ( new_n1345_, new_n1342_, new_n1344_ );
or g1274 ( new_n1346_, new_n1340_, new_n1345_ );
and g1275 ( new_n1347_, new_n1346_, new_n1336_ );
or g1276 ( new_n1348_, new_n1335_, new_n1347_ );
and g1277 ( new_n1349_, new_n1348_, keyinput3_G430gat );
not g1278 ( new_n1350_, keyinput3_G430gat );
and g1279 ( new_n1351_, new_n819_, new_n1325_ );
and g1280 ( new_n1352_, new_n821_, keyinput0_G430gat );
or g1281 ( new_n1353_, new_n1351_, new_n1352_ );
and g1282 ( new_n1354_, new_n1353_, new_n1329_ );
and g1283 ( new_n1355_, new_n87_, new_n1325_ );
or g1284 ( new_n1356_, new_n1355_, new_n1331_ );
and g1285 ( new_n1357_, new_n1356_, keyinput1_G430gat );
or g1286 ( new_n1358_, new_n1354_, new_n1357_ );
and g1287 ( new_n1359_, new_n1358_, keyinput2_G430gat );
and g1288 ( new_n1360_, new_n79_, keyinput0_G430gat );
and g1289 ( new_n1361_, new_n97_, new_n1325_ );
or g1290 ( new_n1362_, new_n1360_, new_n1361_ );
and g1291 ( new_n1363_, new_n1362_, new_n1329_ );
and g1292 ( new_n1364_, new_n80_, new_n1325_ );
or g1293 ( new_n1365_, new_n104_, new_n1364_ );
and g1294 ( new_n1366_, new_n1365_, keyinput1_G430gat );
or g1295 ( new_n1367_, new_n1363_, new_n1366_ );
and g1296 ( new_n1368_, new_n1367_, new_n1336_ );
or g1297 ( new_n1369_, new_n1359_, new_n1368_ );
and g1298 ( new_n1370_, new_n1369_, new_n1350_ );
or g1299 ( G430gat, new_n1349_, new_n1370_ );
and g1300 ( new_n1372_, new_n876_, G92gat );
and g1301 ( new_n1373_, new_n172_, new_n443_ );
or g1302 ( new_n1374_, new_n1372_, new_n1373_ );
and g1303 ( new_n1375_, new_n1374_, new_n227_ );
and g1304 ( new_n1376_, new_n218_, G92gat );
and g1305 ( new_n1377_, new_n162_, new_n443_ );
or g1306 ( new_n1378_, new_n1376_, new_n1377_ );
and g1307 ( new_n1379_, new_n1378_, G86gat );
or g1308 ( new_n1380_, new_n1375_, new_n1379_ );
and g1309 ( new_n1381_, new_n1380_, G76gat );
and g1310 ( new_n1382_, new_n1024_, G92gat );
and g1311 ( new_n1383_, new_n230_, new_n443_ );
or g1312 ( new_n1384_, new_n1382_, new_n1383_ );
and g1313 ( new_n1385_, new_n1384_, G86gat );
or g1314 ( new_n1386_, new_n526_, new_n443_ );
and g1315 ( new_n1387_, new_n1386_, new_n227_ );
or g1316 ( new_n1388_, new_n1385_, new_n1387_ );
and g1317 ( new_n1389_, new_n1388_, new_n173_ );
or g1318 ( new_n1390_, new_n1381_, new_n1389_ );
and g1319 ( new_n1391_, new_n1390_, G82gat );
and g1320 ( new_n1392_, new_n218_, new_n251_ );
or g1321 ( new_n1393_, new_n1391_, new_n1392_ );
and g1322 ( new_n1394_, new_n1393_, G79gat );
and g1323 ( new_n1395_, new_n162_, G86gat );
or g1324 ( new_n1396_, new_n1375_, new_n1395_ );
and g1325 ( new_n1397_, new_n1396_, G76gat );
or g1326 ( new_n1398_, new_n1397_, new_n1389_ );
and g1327 ( new_n1399_, new_n1398_, G82gat );
and g1328 ( new_n1400_, new_n162_, new_n251_ );
or g1329 ( new_n1401_, new_n1399_, new_n1400_ );
and g1330 ( new_n1402_, new_n1401_, new_n490_ );
or g1331 ( new_n1403_, new_n1394_, new_n1402_ );
and g1332 ( new_n1404_, new_n1403_, G73gat );
and g1333 ( new_n1405_, new_n876_, G86gat );
or g1334 ( new_n1406_, new_n1375_, new_n1405_ );
and g1335 ( new_n1407_, new_n1406_, G76gat );
or g1336 ( new_n1408_, new_n1407_, new_n1389_ );
and g1337 ( new_n1409_, new_n1408_, G82gat );
and g1338 ( new_n1410_, new_n876_, new_n251_ );
or g1339 ( new_n1411_, new_n1409_, new_n1410_ );
or g1340 ( new_n1412_, new_n1411_, new_n490_ );
and g1341 ( new_n1413_, new_n1389_, G82gat );
or g1342 ( new_n1414_, new_n1413_, new_n176_ );
or g1343 ( new_n1415_, new_n1414_, G79gat );
and g1344 ( new_n1416_, new_n1415_, new_n256_ );
and g1345 ( new_n1417_, new_n1412_, new_n1416_ );
or g1346 ( new_n1418_, new_n1404_, new_n1417_ );
and g1347 ( new_n1419_, new_n1418_, G63gat );
and g1348 ( new_n1420_, new_n1024_, new_n175_ );
or g1349 ( new_n1421_, new_n1413_, new_n1420_ );
and g1350 ( new_n1422_, new_n1421_, G79gat );
and g1351 ( new_n1423_, new_n1387_, new_n174_ );
or g1352 ( new_n1424_, new_n1423_, new_n259_ );
and g1353 ( new_n1425_, new_n1424_, new_n490_ );
or g1354 ( new_n1426_, new_n1422_, new_n1425_ );
and g1355 ( new_n1427_, new_n1426_, G73gat );
or g1356 ( new_n1428_, new_n528_, new_n490_ );
or g1357 ( new_n1429_, new_n526_, new_n1428_ );
and g1358 ( new_n1430_, new_n1429_, new_n256_ );
or g1359 ( new_n1431_, new_n1427_, new_n1430_ );
and g1360 ( new_n1432_, new_n1431_, new_n177_ );
or g1361 ( new_n1433_, new_n1419_, new_n1432_ );
and g1362 ( new_n1434_, new_n1433_, G69gat );
and g1363 ( new_n1435_, new_n1393_, new_n265_ );
or g1364 ( new_n1436_, new_n1434_, new_n1435_ );
and g1365 ( new_n1437_, new_n1436_, G66gat );
and g1366 ( new_n1438_, new_n1375_, G76gat );
or g1367 ( new_n1439_, new_n1438_, new_n1389_ );
and g1368 ( new_n1440_, new_n1439_, G82gat );
and g1369 ( new_n1441_, new_n1440_, G73gat );
or g1370 ( new_n1442_, new_n1417_, new_n1441_ );
and g1371 ( new_n1443_, new_n1442_, G63gat );
or g1372 ( new_n1444_, new_n1443_, new_n1432_ );
and g1373 ( new_n1445_, new_n1444_, G69gat );
and g1374 ( new_n1446_, new_n1440_, new_n265_ );
or g1375 ( new_n1447_, new_n1445_, new_n1446_ );
and g1376 ( new_n1448_, new_n1447_, new_n541_ );
or g1377 ( new_n1449_, new_n1437_, new_n1448_ );
and g1378 ( new_n1450_, new_n1449_, G60gat );
and g1379 ( new_n1451_, new_n577_, G63gat );
and g1380 ( new_n1452_, new_n1414_, new_n1451_ );
or g1381 ( new_n1453_, new_n1432_, new_n1452_ );
and g1382 ( new_n1454_, new_n1453_, G69gat );
and g1383 ( new_n1455_, new_n227_, G76gat );
and g1384 ( new_n1456_, new_n1373_, new_n1455_ );
or g1385 ( new_n1457_, new_n1389_, new_n1456_ );
and g1386 ( new_n1458_, new_n882_, G82gat );
and g1387 ( new_n1459_, new_n1457_, new_n1458_ );
or g1388 ( new_n1460_, new_n1454_, new_n1459_ );
and g1389 ( new_n1461_, new_n1460_, G66gat );
and g1390 ( new_n1462_, new_n1432_, G69gat );
and g1391 ( new_n1463_, new_n1413_, new_n179_ );
or g1392 ( new_n1464_, new_n1462_, new_n1463_ );
and g1393 ( new_n1465_, new_n1464_, new_n541_ );
or g1394 ( new_n1466_, new_n1461_, new_n1465_ );
and g1395 ( new_n1467_, new_n1466_, new_n281_ );
or g1396 ( new_n1468_, new_n1450_, new_n1467_ );
and g1397 ( new_n1469_, new_n1468_, G50gat );
or g1398 ( new_n1470_, new_n1430_, new_n943_ );
or g1399 ( new_n1471_, new_n1425_, new_n1470_ );
not g1400 ( new_n1472_, new_n943_ );
or g1401 ( new_n1473_, new_n1387_, new_n1383_ );
and g1402 ( new_n1474_, new_n1473_, new_n174_ );
or g1403 ( new_n1475_, new_n1474_, new_n1472_ );
and g1404 ( new_n1476_, new_n1471_, new_n1475_ );
and g1405 ( new_n1477_, new_n1476_, G66gat );
and g1406 ( new_n1478_, new_n1423_, new_n283_ );
and g1407 ( new_n1479_, new_n1429_, new_n282_ );
or g1408 ( new_n1480_, new_n1478_, new_n1479_ );
and g1409 ( new_n1481_, new_n1480_, new_n541_ );
or g1410 ( new_n1482_, new_n1477_, new_n1481_ );
and g1411 ( new_n1483_, new_n1482_, G60gat );
or g1412 ( new_n1484_, new_n528_, new_n578_ );
and g1413 ( new_n1485_, new_n1484_, G66gat );
and g1414 ( new_n1486_, new_n1485_, new_n281_ );
or g1415 ( new_n1487_, new_n1483_, new_n1486_ );
and g1416 ( new_n1488_, new_n1487_, new_n181_ );
or g1417 ( new_n1489_, new_n1469_, new_n1488_ );
and g1418 ( new_n1490_, new_n1489_, G56gat );
and g1419 ( new_n1491_, new_n1436_, new_n272_ );
or g1420 ( new_n1492_, new_n1490_, new_n1491_ );
and g1421 ( new_n1493_, new_n1492_, G53gat );
and g1422 ( new_n1494_, new_n1447_, G60gat );
or g1423 ( new_n1495_, new_n1467_, new_n1494_ );
and g1424 ( new_n1496_, new_n1495_, G50gat );
or g1425 ( new_n1497_, new_n1496_, new_n1488_ );
and g1426 ( new_n1498_, new_n1497_, G56gat );
and g1427 ( new_n1499_, new_n1447_, new_n272_ );
or g1428 ( new_n1500_, new_n1498_, new_n1499_ );
and g1429 ( new_n1501_, new_n1500_, new_n589_ );
or g1430 ( new_n1502_, new_n1493_, new_n1501_ );
and g1431 ( new_n1503_, new_n1502_, G47gat );
and g1432 ( new_n1504_, new_n1465_, new_n281_ );
and g1433 ( new_n1505_, new_n1504_, G50gat );
or g1434 ( new_n1506_, new_n1505_, new_n1488_ );
and g1435 ( new_n1507_, new_n1506_, G56gat );
and g1436 ( new_n1508_, new_n1460_, new_n891_ );
or g1437 ( new_n1509_, new_n1507_, new_n1508_ );
and g1438 ( new_n1510_, new_n1509_, G53gat );
and g1439 ( new_n1511_, new_n1464_, new_n183_ );
and g1440 ( new_n1512_, new_n1488_, G56gat );
or g1441 ( new_n1513_, new_n1511_, new_n1512_ );
and g1442 ( new_n1514_, new_n1513_, new_n589_ );
or g1443 ( new_n1515_, new_n1510_, new_n1514_ );
and g1444 ( new_n1516_, new_n1515_, new_n320_ );
or g1445 ( new_n1517_, new_n1503_, new_n1516_ );
and g1446 ( new_n1518_, new_n1517_, G37gat );
and g1447 ( new_n1519_, new_n1476_, new_n183_ );
or g1448 ( new_n1520_, new_n1512_, new_n1519_ );
and g1449 ( new_n1521_, new_n1520_, G53gat );
and g1450 ( new_n1522_, new_n1480_, new_n300_ );
and g1451 ( new_n1523_, new_n1485_, new_n299_ );
or g1452 ( new_n1524_, new_n1522_, new_n1523_ );
and g1453 ( new_n1525_, new_n1524_, new_n589_ );
or g1454 ( new_n1526_, new_n1521_, new_n1525_ );
and g1455 ( new_n1527_, new_n1526_, G47gat );
and g1456 ( new_n1528_, new_n1484_, new_n320_ );
and g1457 ( new_n1529_, new_n1077_, new_n1528_ );
or g1458 ( new_n1530_, new_n1527_, new_n1529_ );
and g1459 ( new_n1531_, new_n1530_, new_n185_ );
or g1460 ( new_n1532_, new_n1518_, new_n1531_ );
and g1461 ( new_n1533_, new_n1532_, G43gat );
and g1462 ( new_n1534_, new_n1492_, new_n290_ );
or g1463 ( new_n1535_, new_n1533_, new_n1534_ );
and g1464 ( new_n1536_, new_n1535_, G40gat );
and g1465 ( new_n1537_, new_n1401_, G73gat );
or g1466 ( new_n1538_, new_n1417_, new_n1537_ );
and g1467 ( new_n1539_, new_n1538_, G63gat );
or g1468 ( new_n1540_, new_n1539_, new_n1432_ );
and g1469 ( new_n1541_, new_n1540_, G69gat );
and g1470 ( new_n1542_, new_n1401_, new_n265_ );
or g1471 ( new_n1543_, new_n1541_, new_n1542_ );
and g1472 ( new_n1544_, new_n1543_, G60gat );
or g1473 ( new_n1545_, new_n1467_, new_n1544_ );
and g1474 ( new_n1546_, new_n1545_, G50gat );
or g1475 ( new_n1547_, new_n1546_, new_n1488_ );
and g1476 ( new_n1548_, new_n1547_, G56gat );
and g1477 ( new_n1549_, new_n1543_, new_n272_ );
or g1478 ( new_n1550_, new_n1548_, new_n1549_ );
and g1479 ( new_n1551_, new_n1550_, G47gat );
or g1480 ( new_n1552_, new_n1551_, new_n1516_ );
and g1481 ( new_n1553_, new_n1552_, G37gat );
or g1482 ( new_n1554_, new_n1553_, new_n1531_ );
and g1483 ( new_n1555_, new_n1554_, G43gat );
and g1484 ( new_n1556_, new_n1550_, new_n290_ );
or g1485 ( new_n1557_, new_n1555_, new_n1556_ );
and g1486 ( new_n1558_, new_n1557_, new_n639_ );
or g1487 ( new_n1559_, new_n1536_, new_n1558_ );
and g1488 ( new_n1560_, new_n1559_, G34gat );
and g1489 ( new_n1561_, new_n1411_, G73gat );
or g1490 ( new_n1562_, new_n1417_, new_n1561_ );
and g1491 ( new_n1563_, new_n1562_, G63gat );
or g1492 ( new_n1564_, new_n1563_, new_n1432_ );
and g1493 ( new_n1565_, new_n1564_, G69gat );
and g1494 ( new_n1566_, new_n1411_, new_n265_ );
or g1495 ( new_n1567_, new_n1565_, new_n1566_ );
and g1496 ( new_n1568_, new_n1567_, new_n889_ );
or g1497 ( new_n1569_, new_n1568_, new_n1504_ );
and g1498 ( new_n1570_, new_n1569_, G50gat );
or g1499 ( new_n1571_, new_n1570_, new_n1488_ );
and g1500 ( new_n1572_, new_n1571_, G56gat );
and g1501 ( new_n1573_, new_n1567_, new_n272_ );
or g1502 ( new_n1574_, new_n1572_, new_n1573_ );
or g1503 ( new_n1575_, new_n1574_, new_n676_ );
or g1504 ( new_n1576_, new_n1513_, new_n892_ );
and g1505 ( new_n1577_, new_n1576_, G37gat );
and g1506 ( new_n1578_, new_n1575_, new_n1577_ );
or g1507 ( new_n1579_, new_n1578_, new_n1531_ );
and g1508 ( new_n1580_, new_n1579_, G43gat );
and g1509 ( new_n1581_, new_n1574_, new_n290_ );
or g1510 ( new_n1582_, new_n1580_, new_n1581_ );
and g1511 ( new_n1583_, new_n1582_, G40gat );
and g1512 ( new_n1584_, new_n1531_, G43gat );
and g1513 ( new_n1585_, new_n1414_, new_n179_ );
or g1514 ( new_n1586_, new_n1462_, new_n1585_ );
and g1515 ( new_n1587_, new_n1586_, new_n183_ );
or g1516 ( new_n1588_, new_n1587_, new_n1512_ );
and g1517 ( new_n1589_, new_n1588_, new_n187_ );
or g1518 ( new_n1590_, new_n1584_, new_n1589_ );
and g1519 ( new_n1591_, new_n1590_, new_n639_ );
or g1520 ( new_n1592_, new_n1583_, new_n1591_ );
and g1521 ( new_n1593_, new_n1592_, new_n316_ );
or g1522 ( new_n1594_, new_n1560_, new_n1593_ );
and g1523 ( new_n1595_, new_n1594_, G24gat );
and g1524 ( new_n1596_, new_n1481_, G60gat );
or g1525 ( new_n1597_, new_n1596_, new_n1486_ );
and g1526 ( new_n1598_, new_n1597_, new_n182_ );
or g1527 ( new_n1599_, new_n1421_, new_n1472_ );
and g1528 ( new_n1600_, new_n1471_, new_n934_ );
and g1529 ( new_n1601_, new_n1599_, new_n1600_ );
or g1530 ( new_n1602_, new_n1598_, new_n1601_ );
and g1531 ( new_n1603_, new_n1602_, new_n930_ );
and g1532 ( new_n1604_, new_n1525_, G47gat );
or g1533 ( new_n1605_, new_n1604_, new_n1529_ );
and g1534 ( new_n1606_, new_n1605_, new_n186_ );
or g1535 ( new_n1607_, new_n1603_, new_n1606_ );
and g1536 ( new_n1608_, new_n1607_, G40gat );
and g1537 ( new_n1609_, new_n1424_, new_n283_ );
or g1538 ( new_n1610_, new_n1609_, new_n1479_ );
and g1539 ( new_n1611_, new_n1610_, new_n300_ );
or g1540 ( new_n1612_, new_n1611_, new_n1523_ );
and g1541 ( new_n1613_, new_n1612_, new_n322_ );
and g1542 ( new_n1614_, new_n1529_, new_n186_ );
or g1543 ( new_n1615_, new_n1613_, new_n1614_ );
and g1544 ( new_n1616_, new_n1615_, new_n639_ );
or g1545 ( new_n1617_, new_n1608_, new_n1616_ );
and g1546 ( new_n1618_, new_n1617_, G34gat );
or g1547 ( new_n1619_, new_n526_, new_n1484_ );
and g1548 ( new_n1620_, new_n1619_, new_n1123_ );
or g1549 ( new_n1621_, new_n1620_, new_n639_ );
and g1550 ( new_n1622_, new_n1621_, new_n316_ );
or g1551 ( new_n1623_, new_n1618_, new_n1622_ );
and g1552 ( new_n1624_, new_n1623_, new_n189_ );
or g1553 ( new_n1625_, new_n1595_, new_n1624_ );
and g1554 ( new_n1626_, new_n1625_, G30gat );
and g1555 ( new_n1627_, new_n1535_, new_n307_ );
or g1556 ( new_n1628_, new_n1626_, new_n1627_ );
and g1557 ( new_n1629_, new_n1628_, G14gat );
and g1558 ( new_n1630_, new_n1402_, G73gat );
or g1559 ( new_n1631_, new_n1417_, new_n1630_ );
and g1560 ( new_n1632_, new_n1631_, G63gat );
or g1561 ( new_n1633_, new_n1632_, new_n1432_ );
and g1562 ( new_n1634_, new_n1633_, G69gat );
and g1563 ( new_n1635_, new_n1395_, new_n443_ );
or g1564 ( new_n1636_, new_n1375_, new_n1635_ );
and g1565 ( new_n1637_, new_n1636_, G76gat );
or g1566 ( new_n1638_, new_n1637_, new_n1389_ );
and g1567 ( new_n1639_, new_n854_, G82gat );
and g1568 ( new_n1640_, new_n1638_, new_n1639_ );
or g1569 ( new_n1641_, new_n1634_, new_n1640_ );
and g1570 ( new_n1642_, new_n1641_, G66gat );
or g1571 ( new_n1643_, new_n1642_, new_n1448_ );
and g1572 ( new_n1644_, new_n1643_, G60gat );
or g1573 ( new_n1645_, new_n1644_, new_n1467_ );
and g1574 ( new_n1646_, new_n1645_, G50gat );
or g1575 ( new_n1647_, new_n1646_, new_n1488_ );
and g1576 ( new_n1648_, new_n1647_, G56gat );
and g1577 ( new_n1649_, new_n1641_, new_n272_ );
or g1578 ( new_n1650_, new_n1648_, new_n1649_ );
and g1579 ( new_n1651_, new_n1650_, G53gat );
or g1580 ( new_n1652_, new_n1651_, new_n1501_ );
and g1581 ( new_n1653_, new_n1652_, G47gat );
or g1582 ( new_n1654_, new_n1653_, new_n1516_ );
and g1583 ( new_n1655_, new_n1654_, G37gat );
or g1584 ( new_n1656_, new_n1655_, new_n1531_ );
and g1585 ( new_n1657_, new_n1656_, G43gat );
and g1586 ( new_n1658_, new_n1650_, new_n290_ );
or g1587 ( new_n1659_, new_n1657_, new_n1658_ );
and g1588 ( new_n1660_, new_n1659_, G40gat );
or g1589 ( new_n1661_, new_n1660_, new_n1558_ );
and g1590 ( new_n1662_, new_n1661_, G34gat );
or g1591 ( new_n1663_, new_n1662_, new_n1593_ );
and g1592 ( new_n1664_, new_n1663_, G24gat );
or g1593 ( new_n1665_, new_n1664_, new_n1624_ );
and g1594 ( new_n1666_, new_n1665_, G30gat );
and g1595 ( new_n1667_, new_n1659_, new_n307_ );
or g1596 ( new_n1668_, new_n1666_, new_n1667_ );
and g1597 ( new_n1669_, new_n1668_, new_n701_ );
or g1598 ( new_n1670_, new_n1629_, new_n1669_ );
and g1599 ( new_n1671_, new_n1670_, G27gat );
and g1600 ( new_n1672_, new_n1592_, new_n317_ );
or g1601 ( new_n1673_, new_n1672_, new_n1624_ );
and g1602 ( new_n1674_, new_n1673_, G30gat );
and g1603 ( new_n1675_, new_n1557_, new_n309_ );
or g1604 ( new_n1676_, new_n1674_, new_n1675_ );
and g1605 ( new_n1677_, new_n1676_, new_n690_ );
or g1606 ( new_n1678_, new_n1671_, new_n1677_ );
and g1607 ( new_n1679_, new_n1678_, G21gat );
and g1608 ( new_n1680_, new_n1582_, G34gat );
or g1609 ( new_n1681_, new_n1593_, new_n1680_ );
and g1610 ( new_n1682_, new_n1681_, G24gat );
or g1611 ( new_n1683_, new_n1682_, new_n1624_ );
and g1612 ( new_n1684_, new_n1683_, G30gat );
and g1613 ( new_n1685_, new_n1582_, new_n307_ );
or g1614 ( new_n1686_, new_n1684_, new_n1685_ );
and g1615 ( new_n1687_, new_n1686_, G27gat );
and g1616 ( new_n1688_, new_n1590_, new_n191_ );
and g1617 ( new_n1689_, new_n1624_, G30gat );
or g1618 ( new_n1690_, new_n1688_, new_n1689_ );
and g1619 ( new_n1691_, new_n1690_, new_n690_ );
or g1620 ( new_n1692_, new_n1687_, new_n1691_ );
and g1621 ( new_n1693_, new_n1692_, new_n337_ );
or g1622 ( new_n1694_, new_n1679_, new_n1693_ );
and g1623 ( new_n1695_, new_n1694_, G8gat );
and g1624 ( new_n1696_, new_n1686_, G14gat );
and g1625 ( new_n1697_, new_n1591_, new_n317_ );
or g1626 ( new_n1698_, new_n1697_, new_n1624_ );
and g1627 ( new_n1699_, new_n1698_, G30gat );
and g1628 ( new_n1700_, new_n1513_, new_n1190_ );
or g1629 ( new_n1701_, new_n1531_, new_n1700_ );
and g1630 ( new_n1702_, new_n1701_, G43gat );
and g1631 ( new_n1703_, new_n1509_, new_n894_ );
or g1632 ( new_n1704_, new_n1702_, new_n1703_ );
and g1633 ( new_n1705_, new_n1704_, new_n887_ );
or g1634 ( new_n1706_, new_n1699_, new_n1705_ );
and g1635 ( new_n1707_, new_n1706_, new_n701_ );
or g1636 ( new_n1708_, new_n1696_, new_n1707_ );
and g1637 ( new_n1709_, new_n1708_, G27gat );
or g1638 ( new_n1710_, new_n1709_, new_n1691_ );
and g1639 ( new_n1711_, new_n1710_, new_n337_ );
and g1640 ( new_n1712_, new_n1516_, G37gat );
or g1641 ( new_n1713_, new_n1712_, new_n1531_ );
and g1642 ( new_n1714_, new_n1713_, G43gat );
and g1643 ( new_n1715_, new_n1500_, new_n292_ );
or g1644 ( new_n1716_, new_n1714_, new_n1715_ );
and g1645 ( new_n1717_, new_n1716_, new_n309_ );
or g1646 ( new_n1718_, new_n1674_, new_n1717_ );
and g1647 ( new_n1719_, new_n1718_, G14gat );
or g1648 ( new_n1720_, new_n1719_, new_n1707_ );
and g1649 ( new_n1721_, new_n1720_, G21gat );
or g1650 ( new_n1722_, new_n1711_, new_n1721_ );
and g1651 ( new_n1723_, new_n1722_, new_n352_ );
or g1652 ( new_n1724_, new_n1695_, new_n1723_ );
and g1653 ( new_n1725_, new_n1724_, G11gat );
and g1654 ( new_n1726_, new_n1607_, new_n191_ );
or g1655 ( new_n1727_, new_n1689_, new_n1726_ );
and g1656 ( new_n1728_, new_n1727_, G27gat );
or g1657 ( new_n1729_, new_n1615_, new_n343_ );
or g1658 ( new_n1730_, new_n1621_, new_n344_ );
and g1659 ( new_n1731_, new_n1730_, new_n690_ );
and g1660 ( new_n1732_, new_n1729_, new_n1731_ );
or g1661 ( new_n1733_, new_n1728_, new_n1732_ );
and g1662 ( new_n1734_, new_n1733_, G21gat );
or g1663 ( new_n1735_, new_n1620_, new_n1240_ );
and g1664 ( new_n1736_, new_n1735_, new_n337_ );
or g1665 ( new_n1737_, new_n1734_, new_n1736_ );
and g1666 ( new_n1738_, new_n1737_, new_n193_ );
or g1667 ( new_n1739_, new_n1725_, new_n1738_ );
and g1668 ( new_n1740_, new_n1739_, G17gat );
and g1669 ( new_n1741_, new_n1391_, new_n265_ );
or g1670 ( new_n1742_, new_n1434_, new_n1741_ );
and g1671 ( new_n1743_, new_n1742_, new_n272_ );
or g1672 ( new_n1744_, new_n1648_, new_n1743_ );
and g1673 ( new_n1745_, new_n1744_, new_n290_ );
or g1674 ( new_n1746_, new_n1657_, new_n1745_ );
and g1675 ( new_n1747_, new_n1746_, new_n307_ );
or g1676 ( new_n1748_, new_n1626_, new_n1747_ );
and g1677 ( new_n1749_, new_n1748_, G14gat );
or g1678 ( new_n1750_, new_n1749_, new_n1669_ );
and g1679 ( new_n1751_, new_n1750_, G8gat );
and g1680 ( new_n1752_, new_n1720_, new_n352_ );
or g1681 ( new_n1753_, new_n1751_, new_n1752_ );
and g1682 ( new_n1754_, new_n1753_, new_n331_ );
or g1683 ( new_n1755_, new_n1740_, new_n1754_ );
and g1684 ( new_n1756_, new_n1755_, G1gat );
and g1685 ( new_n1757_, new_n1520_, new_n930_ );
or g1686 ( new_n1758_, new_n1757_, new_n1606_ );
and g1687 ( new_n1759_, new_n1758_, G40gat );
or g1688 ( new_n1760_, new_n1759_, new_n1616_ );
and g1689 ( new_n1761_, new_n1760_, G34gat );
or g1690 ( new_n1762_, new_n1622_, new_n191_ );
or g1691 ( new_n1763_, new_n1761_, new_n1762_ );
or g1692 ( new_n1764_, new_n1758_, new_n190_ );
and g1693 ( new_n1765_, new_n1764_, new_n701_ );
and g1694 ( new_n1766_, new_n1763_, new_n1765_ );
and g1695 ( new_n1767_, new_n1727_, G14gat );
or g1696 ( new_n1768_, new_n1766_, new_n1767_ );
and g1697 ( new_n1769_, new_n1768_, G27gat );
or g1698 ( new_n1770_, new_n1769_, new_n1732_ );
and g1699 ( new_n1771_, new_n1770_, G21gat );
or g1700 ( new_n1772_, new_n1771_, new_n1736_ );
and g1701 ( new_n1773_, new_n1772_, G8gat );
and g1702 ( new_n1774_, new_n1524_, new_n322_ );
or g1703 ( new_n1775_, new_n1614_, new_n343_ );
or g1704 ( new_n1776_, new_n1774_, new_n1775_ );
and g1705 ( new_n1777_, new_n1730_, G14gat );
and g1706 ( new_n1778_, new_n1776_, new_n1777_ );
and g1707 ( new_n1779_, new_n1123_, new_n1484_ );
or g1708 ( new_n1780_, new_n1779_, new_n743_ );
and g1709 ( new_n1781_, new_n1780_, new_n701_ );
or g1710 ( new_n1782_, new_n1778_, new_n1781_ );
and g1711 ( new_n1783_, new_n1782_, G21gat );
or g1712 ( new_n1784_, new_n1780_, new_n690_ );
and g1713 ( new_n1785_, new_n1784_, new_n701_ );
and g1714 ( new_n1786_, new_n1735_, G14gat );
or g1715 ( new_n1787_, new_n1785_, new_n1786_ );
and g1716 ( new_n1788_, new_n1787_, new_n337_ );
or g1717 ( new_n1789_, new_n1783_, new_n1788_ );
and g1718 ( new_n1790_, new_n1789_, new_n352_ );
or g1719 ( new_n1791_, new_n1773_, new_n1790_ );
and g1720 ( new_n1792_, new_n1791_, new_n194_ );
and g1721 ( new_n1793_, new_n1513_, new_n187_ );
or g1722 ( new_n1794_, new_n1584_, new_n1793_ );
and g1723 ( new_n1795_, new_n1794_, new_n191_ );
or g1724 ( new_n1796_, new_n1795_, new_n1689_ );
and g1725 ( new_n1797_, new_n1796_, G14gat );
or g1726 ( new_n1798_, new_n1797_, new_n1766_ );
and g1727 ( new_n1799_, new_n1798_, G8gat );
and g1728 ( new_n1800_, new_n1782_, new_n352_ );
or g1729 ( new_n1801_, new_n1799_, new_n1800_ );
and g1730 ( new_n1802_, new_n1801_, new_n195_ );
or g1731 ( new_n1803_, new_n1792_, new_n1802_ );
and g1732 ( new_n1804_, new_n1803_, new_n356_ );
or g1733 ( new_n1805_, new_n1756_, new_n1804_ );
and g1734 ( new_n1806_, new_n1805_, G4gat );
and g1735 ( new_n1807_, new_n1628_, G27gat );
or g1736 ( new_n1808_, new_n1807_, new_n1677_ );
and g1737 ( new_n1809_, new_n1808_, G21gat );
or g1738 ( new_n1810_, new_n1809_, new_n1693_ );
and g1739 ( new_n1811_, new_n1810_, G11gat );
or g1740 ( new_n1812_, new_n1811_, new_n1738_ );
and g1741 ( new_n1813_, new_n1812_, G17gat );
and g1742 ( new_n1814_, new_n1748_, new_n331_ );
or g1743 ( new_n1815_, new_n1813_, new_n1814_ );
and g1744 ( new_n1816_, new_n1815_, new_n196_ );
or g1745 ( new_n1817_, new_n1806_, new_n1816_ );
and g1746 ( new_n1818_, new_n1817_, keyinput0_G431gat );
not g1747 ( new_n1819_, keyinput0_G431gat );
and g1748 ( new_n1820_, new_n75_, new_n1819_ );
or g1749 ( new_n1821_, new_n1818_, new_n1820_ );
and g1750 ( new_n1822_, new_n1821_, keyinput1_G431gat );
not g1751 ( new_n1823_, keyinput1_G431gat );
and g1752 ( new_n1824_, new_n423_, new_n1819_ );
and g1753 ( new_n1825_, new_n102_, keyinput0_G431gat );
or g1754 ( new_n1826_, new_n1824_, new_n1825_ );
and g1755 ( new_n1827_, new_n1826_, new_n1823_ );
or g1756 ( new_n1828_, new_n1822_, new_n1827_ );
and g1757 ( new_n1829_, new_n1828_, keyinput2_G431gat );
not g1758 ( new_n1830_, keyinput2_G431gat );
and g1759 ( new_n1831_, new_n114_, new_n1819_ );
and g1760 ( new_n1832_, new_n803_, keyinput0_G431gat );
or g1761 ( new_n1833_, new_n1831_, new_n1832_ );
and g1762 ( new_n1834_, new_n1833_, new_n1823_ );
and g1763 ( new_n1835_, new_n112_, new_n1819_ );
not g1764 ( new_n1836_, new_n1835_ );
not g1765 ( new_n1837_, new_n1825_ );
and g1766 ( new_n1838_, new_n1837_, keyinput1_G431gat );
and g1767 ( new_n1839_, new_n1836_, new_n1838_ );
or g1768 ( new_n1840_, new_n1834_, new_n1839_ );
and g1769 ( new_n1841_, new_n1840_, new_n1830_ );
or g1770 ( new_n1842_, new_n1829_, new_n1841_ );
and g1771 ( new_n1843_, new_n1842_, keyinput3_G431gat );
not g1772 ( new_n1844_, keyinput3_G431gat );
and g1773 ( new_n1845_, new_n819_, new_n1819_ );
and g1774 ( new_n1846_, new_n821_, keyinput0_G431gat );
or g1775 ( new_n1847_, new_n1845_, new_n1846_ );
and g1776 ( new_n1848_, new_n1847_, new_n1823_ );
and g1777 ( new_n1849_, new_n87_, new_n1819_ );
or g1778 ( new_n1850_, new_n1849_, new_n1825_ );
and g1779 ( new_n1851_, new_n1850_, keyinput1_G431gat );
or g1780 ( new_n1852_, new_n1848_, new_n1851_ );
and g1781 ( new_n1853_, new_n1852_, keyinput2_G431gat );
and g1782 ( new_n1854_, new_n79_, keyinput0_G431gat );
and g1783 ( new_n1855_, new_n97_, new_n1819_ );
or g1784 ( new_n1856_, new_n1854_, new_n1855_ );
and g1785 ( new_n1857_, new_n1856_, new_n1823_ );
and g1786 ( new_n1858_, new_n80_, new_n1819_ );
or g1787 ( new_n1859_, new_n104_, new_n1858_ );
and g1788 ( new_n1860_, new_n1859_, keyinput1_G431gat );
or g1789 ( new_n1861_, new_n1857_, new_n1860_ );
and g1790 ( new_n1862_, new_n1861_, new_n1830_ );
or g1791 ( new_n1863_, new_n1853_, new_n1862_ );
and g1792 ( new_n1864_, new_n1863_, new_n1844_ );
or g1793 ( G431gat, new_n1843_, new_n1864_ );
and g1794 ( new_n1866_, new_n84_, G89gat );
or g1795 ( new_n1867_, new_n108_, new_n1866_ );
and g1796 ( new_n1868_, new_n1867_, G95gat );
and g1797 ( new_n1869_, new_n1868_, new_n443_ );
and g1798 ( new_n1870_, G92gat, G95gat );
and g1799 ( new_n1871_, new_n109_, new_n1870_ );
or g1800 ( new_n1872_, new_n1869_, new_n1871_ );
and g1801 ( new_n1873_, new_n1872_, G86gat );
and g1802 ( new_n1874_, new_n418_, new_n392_ );
or g1803 ( new_n1875_, new_n108_, new_n1874_ );
and g1804 ( new_n1876_, new_n1875_, G95gat );
and g1805 ( new_n1877_, new_n1876_, G92gat );
and g1806 ( new_n1878_, new_n108_, G95gat );
and g1807 ( new_n1879_, new_n1878_, new_n443_ );
or g1808 ( new_n1880_, new_n1877_, new_n1879_ );
and g1809 ( new_n1881_, new_n1880_, new_n227_ );
or g1810 ( new_n1882_, new_n1873_, new_n1881_ );
and g1811 ( new_n1883_, new_n1882_, G76gat );
or g1812 ( new_n1884_, new_n106_, new_n98_ );
and g1813 ( new_n1885_, new_n1884_, new_n170_ );
and g1814 ( new_n1886_, new_n1885_, G92gat );
and g1815 ( new_n1887_, new_n106_, new_n170_ );
and g1816 ( new_n1888_, new_n1887_, new_n443_ );
or g1817 ( new_n1889_, new_n1886_, new_n1888_ );
and g1818 ( new_n1890_, new_n1889_, G86gat );
and g1819 ( new_n1891_, new_n479_, G92gat );
and g1820 ( new_n1892_, new_n1891_, new_n227_ );
or g1821 ( new_n1893_, new_n1890_, new_n1892_ );
and g1822 ( new_n1894_, new_n1893_, new_n173_ );
or g1823 ( new_n1895_, new_n1883_, new_n1894_ );
and g1824 ( new_n1896_, new_n1895_, G82gat );
and g1825 ( new_n1897_, new_n251_, G95gat );
and g1826 ( new_n1898_, new_n109_, new_n1897_ );
or g1827 ( new_n1899_, new_n1896_, new_n1898_ );
and g1828 ( new_n1900_, new_n1899_, G79gat );
or g1829 ( new_n1901_, new_n84_, new_n89_ );
and g1830 ( new_n1902_, new_n1901_, G89gat );
or g1831 ( new_n1903_, new_n1902_, new_n108_ );
and g1832 ( new_n1904_, new_n1903_, G95gat );
and g1833 ( new_n1905_, new_n88_, new_n160_ );
or g1834 ( new_n1906_, new_n1904_, new_n1905_ );
and g1835 ( new_n1907_, new_n1906_, G86gat );
or g1836 ( new_n1908_, new_n1881_, new_n1907_ );
and g1837 ( new_n1909_, new_n1908_, G76gat );
or g1838 ( new_n1910_, new_n1909_, new_n1894_ );
and g1839 ( new_n1911_, new_n1910_, G82gat );
and g1840 ( new_n1912_, new_n1906_, new_n251_ );
or g1841 ( new_n1913_, new_n1911_, new_n1912_ );
and g1842 ( new_n1914_, new_n1913_, new_n490_ );
or g1843 ( new_n1915_, new_n1900_, new_n1914_ );
and g1844 ( new_n1916_, new_n1915_, G73gat );
and g1845 ( new_n1917_, new_n78_, G99gat );
or g1846 ( new_n1918_, new_n84_, new_n1917_ );
and g1847 ( new_n1919_, new_n1918_, G89gat );
or g1848 ( new_n1920_, new_n1919_, new_n108_ );
and g1849 ( new_n1921_, new_n1920_, G95gat );
or g1850 ( new_n1922_, new_n1921_, new_n875_ );
or g1851 ( new_n1923_, new_n1922_, new_n527_ );
or g1852 ( new_n1924_, new_n1878_, new_n877_ );
and g1853 ( new_n1925_, new_n1924_, G76gat );
and g1854 ( new_n1926_, new_n1923_, new_n1925_ );
or g1855 ( new_n1927_, new_n1926_, new_n1894_ );
and g1856 ( new_n1928_, new_n1927_, G82gat );
and g1857 ( new_n1929_, new_n1922_, new_n251_ );
or g1858 ( new_n1930_, new_n1928_, new_n1929_ );
and g1859 ( new_n1931_, new_n1930_, G79gat );
and g1860 ( new_n1932_, new_n1894_, G82gat );
and g1861 ( new_n1933_, new_n1878_, new_n175_ );
or g1862 ( new_n1934_, new_n1932_, new_n1933_ );
or g1863 ( new_n1935_, new_n1934_, new_n176_ );
and g1864 ( new_n1936_, new_n1935_, new_n490_ );
or g1865 ( new_n1937_, new_n1931_, new_n1936_ );
and g1866 ( new_n1938_, new_n1937_, new_n256_ );
or g1867 ( new_n1939_, new_n1916_, new_n1938_ );
and g1868 ( new_n1940_, new_n1939_, G63gat );
and g1869 ( new_n1941_, new_n95_, new_n171_ );
or g1870 ( new_n1942_, new_n1878_, new_n1941_ );
and g1871 ( new_n1943_, new_n1942_, new_n942_ );
and g1872 ( new_n1944_, new_n1888_, G86gat );
or g1873 ( new_n1945_, new_n1944_, new_n1892_ );
and g1874 ( new_n1946_, new_n1945_, new_n174_ );
or g1875 ( new_n1947_, new_n1943_, new_n1946_ );
and g1876 ( new_n1948_, new_n1947_, G79gat );
and g1877 ( new_n1949_, new_n228_, new_n372_ );
or g1878 ( new_n1950_, new_n1949_, new_n97_ );
and g1879 ( new_n1951_, new_n1950_, new_n258_ );
or g1880 ( new_n1952_, new_n1951_, new_n1891_ );
and g1881 ( new_n1953_, new_n1952_, new_n490_ );
or g1882 ( new_n1954_, new_n1948_, new_n1953_ );
and g1883 ( new_n1955_, new_n1954_, G73gat );
or g1884 ( new_n1956_, new_n104_, new_n479_ );
and g1885 ( new_n1957_, new_n1956_, new_n529_ );
or g1886 ( new_n1958_, new_n1957_, new_n490_ );
and g1887 ( new_n1959_, new_n1958_, new_n256_ );
or g1888 ( new_n1960_, new_n1955_, new_n1959_ );
and g1889 ( new_n1961_, new_n1960_, new_n177_ );
or g1890 ( new_n1962_, new_n1940_, new_n1961_ );
and g1891 ( new_n1963_, new_n1962_, G69gat );
and g1892 ( new_n1964_, new_n1899_, new_n265_ );
or g1893 ( new_n1965_, new_n1963_, new_n1964_ );
and g1894 ( new_n1966_, new_n1965_, G66gat );
and g1895 ( new_n1967_, new_n1899_, G73gat );
or g1896 ( new_n1968_, new_n1938_, new_n1967_ );
and g1897 ( new_n1969_, new_n1968_, G63gat );
or g1898 ( new_n1970_, new_n1969_, new_n1961_ );
and g1899 ( new_n1971_, new_n1970_, G69gat );
or g1900 ( new_n1972_, new_n1971_, new_n1964_ );
and g1901 ( new_n1973_, new_n1972_, new_n541_ );
or g1902 ( new_n1974_, new_n1966_, new_n1973_ );
and g1903 ( new_n1975_, new_n1974_, G60gat );
and g1904 ( new_n1976_, new_n1868_, G86gat );
or g1905 ( new_n1977_, new_n1881_, new_n1976_ );
and g1906 ( new_n1978_, new_n1977_, G76gat );
or g1907 ( new_n1979_, new_n1978_, new_n1894_ );
and g1908 ( new_n1980_, new_n1979_, G82gat );
and g1909 ( new_n1981_, new_n1868_, new_n251_ );
or g1910 ( new_n1982_, new_n1980_, new_n1981_ );
and g1911 ( new_n1983_, new_n1982_, new_n882_ );
and g1912 ( new_n1984_, new_n1935_, new_n577_ );
and g1913 ( new_n1985_, G63gat, G69gat );
and g1914 ( new_n1986_, new_n1984_, new_n1985_ );
or g1915 ( new_n1987_, new_n1983_, new_n1986_ );
and g1916 ( new_n1988_, new_n1987_, G66gat );
and g1917 ( new_n1989_, new_n1961_, G69gat );
and g1918 ( new_n1990_, new_n1879_, new_n1455_ );
or g1919 ( new_n1991_, new_n1894_, new_n1990_ );
and g1920 ( new_n1992_, new_n1991_, G82gat );
and g1921 ( new_n1993_, new_n1876_, new_n879_ );
or g1922 ( new_n1994_, new_n1992_, new_n1993_ );
and g1923 ( new_n1995_, new_n1994_, new_n179_ );
and g1924 ( new_n1996_, new_n1995_, new_n541_ );
or g1925 ( new_n1997_, new_n1989_, new_n1996_ );
or g1926 ( new_n1998_, new_n1988_, new_n1997_ );
and g1927 ( new_n1999_, new_n1998_, new_n281_ );
or g1928 ( new_n2000_, new_n1975_, new_n1999_ );
and g1929 ( new_n2001_, new_n2000_, G50gat );
and g1930 ( new_n2002_, new_n1934_, new_n943_ );
or g1931 ( new_n2003_, new_n1959_, new_n1953_ );
and g1932 ( new_n2004_, new_n2003_, new_n178_ );
or g1933 ( new_n2005_, new_n2002_, new_n2004_ );
and g1934 ( new_n2006_, new_n2005_, G66gat );
and g1935 ( new_n2007_, new_n1885_, new_n942_ );
or g1936 ( new_n2008_, new_n1946_, new_n2007_ );
or g1937 ( new_n2009_, new_n2008_, new_n282_ );
or g1938 ( new_n2010_, new_n1958_, new_n283_ );
and g1939 ( new_n2011_, new_n2010_, new_n541_ );
and g1940 ( new_n2012_, new_n2009_, new_n2011_ );
or g1941 ( new_n2013_, new_n2006_, new_n2012_ );
and g1942 ( new_n2014_, new_n2013_, G60gat );
and g1943 ( new_n2015_, new_n1887_, new_n258_ );
and g1944 ( new_n2016_, new_n1891_, new_n257_ );
or g1945 ( new_n2017_, new_n2015_, new_n2016_ );
or g1946 ( new_n2018_, new_n2017_, new_n578_ );
and g1947 ( new_n2019_, new_n2018_, G66gat );
and g1948 ( new_n2020_, new_n529_, new_n479_ );
and g1949 ( new_n2021_, new_n2020_, new_n541_ );
or g1950 ( new_n2022_, new_n2019_, new_n2021_ );
and g1951 ( new_n2023_, new_n2022_, new_n281_ );
or g1952 ( new_n2024_, new_n2014_, new_n2023_ );
and g1953 ( new_n2025_, new_n2024_, new_n181_ );
or g1954 ( new_n2026_, new_n2001_, new_n2025_ );
and g1955 ( new_n2027_, new_n2026_, G56gat );
and g1956 ( new_n2028_, new_n1965_, new_n272_ );
or g1957 ( new_n2029_, new_n2027_, new_n2028_ );
and g1958 ( new_n2030_, new_n2029_, G53gat );
not g1959 ( new_n2031_, new_n1194_ );
or g1960 ( new_n2032_, new_n1998_, new_n2031_ );
or g1961 ( new_n2033_, new_n2024_, G50gat );
and g1962 ( new_n2034_, new_n2032_, new_n2033_ );
or g1963 ( new_n2035_, new_n2034_, new_n272_ );
and g1964 ( new_n2036_, new_n1913_, G73gat );
or g1965 ( new_n2037_, new_n1938_, new_n2036_ );
and g1966 ( new_n2038_, new_n2037_, G63gat );
or g1967 ( new_n2039_, new_n1961_, new_n265_ );
or g1968 ( new_n2040_, new_n2038_, new_n2039_ );
or g1969 ( new_n2041_, new_n1913_, G69gat );
and g1970 ( new_n2042_, new_n2040_, new_n2041_ );
or g1971 ( new_n2043_, new_n2042_, new_n275_ );
and g1972 ( new_n2044_, new_n2035_, new_n2043_ );
and g1973 ( new_n2045_, new_n2044_, new_n589_ );
or g1974 ( new_n2046_, new_n2030_, new_n2045_ );
and g1975 ( new_n2047_, new_n2046_, G47gat );
not g1976 ( new_n2048_, new_n891_ );
and g1977 ( new_n2049_, new_n1930_, G73gat );
or g1978 ( new_n2050_, new_n1938_, new_n2049_ );
and g1979 ( new_n2051_, new_n2050_, G63gat );
or g1980 ( new_n2052_, new_n2051_, new_n2039_ );
or g1981 ( new_n2053_, new_n1930_, G69gat );
and g1982 ( new_n2054_, new_n2052_, new_n2053_ );
or g1983 ( new_n2055_, new_n2054_, new_n2048_ );
or g1984 ( new_n2056_, new_n889_, new_n181_ );
or g1985 ( new_n2057_, new_n1995_, new_n2056_ );
or g1986 ( new_n2058_, new_n1989_, new_n2057_ );
and g1987 ( new_n2059_, new_n2033_, new_n2058_ );
or g1988 ( new_n2060_, new_n2059_, new_n272_ );
and g1989 ( new_n2061_, new_n2055_, new_n2060_ );
and g1990 ( new_n2062_, new_n2061_, G53gat );
and g1991 ( new_n2063_, new_n2025_, G56gat );
and g1992 ( new_n2064_, new_n1935_, new_n179_ );
or g1993 ( new_n2065_, new_n1989_, new_n2064_ );
and g1994 ( new_n2066_, new_n2065_, new_n183_ );
or g1995 ( new_n2067_, new_n2063_, new_n2066_ );
and g1996 ( new_n2068_, new_n2067_, new_n589_ );
or g1997 ( new_n2069_, new_n2062_, new_n2068_ );
and g1998 ( new_n2070_, new_n2069_, new_n320_ );
or g1999 ( new_n2071_, new_n2047_, new_n2070_ );
and g2000 ( new_n2072_, new_n2071_, G37gat );
and g2001 ( new_n2073_, new_n1947_, new_n179_ );
or g2002 ( new_n2074_, new_n1989_, new_n2073_ );
and g2003 ( new_n2075_, new_n2074_, G66gat );
or g2004 ( new_n2076_, new_n2075_, new_n2012_ );
and g2005 ( new_n2077_, new_n2076_, G60gat );
or g2006 ( new_n2078_, new_n2023_, new_n183_ );
or g2007 ( new_n2079_, new_n2077_, new_n2078_ );
or g2008 ( new_n2080_, new_n2074_, new_n182_ );
and g2009 ( new_n2081_, new_n2079_, new_n2080_ );
or g2010 ( new_n2082_, new_n2081_, new_n589_ );
and g2011 ( new_n2083_, new_n2023_, new_n182_ );
or g2012 ( new_n2084_, new_n1952_, new_n282_ );
and g2013 ( new_n2085_, new_n2010_, new_n300_ );
and g2014 ( new_n2086_, new_n2085_, new_n2084_ );
or g2015 ( new_n2087_, new_n2083_, new_n2086_ );
or g2016 ( new_n2088_, new_n2087_, G53gat );
and g2017 ( new_n2089_, new_n2082_, new_n2088_ );
or g2018 ( new_n2090_, new_n2089_, new_n320_ );
or g2019 ( new_n2091_, new_n1957_, new_n578_ );
or g2020 ( new_n2092_, new_n2020_, new_n627_ );
and g2021 ( new_n2093_, new_n2091_, new_n2092_ );
or g2022 ( new_n2094_, new_n2093_, new_n589_ );
or g2023 ( new_n2095_, new_n2094_, G47gat );
and g2024 ( new_n2096_, new_n2090_, new_n2095_ );
and g2025 ( new_n2097_, new_n2096_, new_n185_ );
or g2026 ( new_n2098_, new_n2072_, new_n2097_ );
and g2027 ( new_n2099_, new_n2098_, G43gat );
and g2028 ( new_n2100_, new_n2029_, new_n290_ );
or g2029 ( new_n2101_, new_n2099_, new_n2100_ );
and g2030 ( new_n2102_, new_n2101_, G40gat );
and g2031 ( new_n2103_, new_n1982_, G73gat );
or g2032 ( new_n2104_, new_n1938_, new_n2103_ );
and g2033 ( new_n2105_, new_n2104_, G63gat );
or g2034 ( new_n2106_, new_n2105_, new_n2039_ );
or g2035 ( new_n2107_, new_n1982_, G69gat );
and g2036 ( new_n2108_, new_n2106_, new_n2107_ );
or g2037 ( new_n2109_, new_n2108_, new_n275_ );
and g2038 ( new_n2110_, new_n2035_, new_n2109_ );
and g2039 ( new_n2111_, new_n2110_, G47gat );
or g2040 ( new_n2112_, new_n2070_, new_n2111_ );
and g2041 ( new_n2113_, new_n2112_, G37gat );
or g2042 ( new_n2114_, new_n2113_, new_n2097_ );
and g2043 ( new_n2115_, new_n2114_, G43gat );
and g2044 ( new_n2116_, new_n2110_, new_n290_ );
or g2045 ( new_n2117_, new_n2115_, new_n2116_ );
and g2046 ( new_n2118_, new_n2117_, new_n639_ );
or g2047 ( new_n2119_, new_n2102_, new_n2118_ );
and g2048 ( new_n2120_, new_n2119_, G34gat );
and g2049 ( new_n2121_, new_n2067_, G37gat );
or g2050 ( new_n2122_, new_n2121_, new_n894_ );
or g2051 ( new_n2123_, new_n2097_, new_n2122_ );
not g2052 ( new_n2124_, new_n894_ );
and g2053 ( new_n2125_, new_n1994_, new_n880_ );
or g2054 ( new_n2126_, new_n1984_, new_n2125_ );
and g2055 ( new_n2127_, new_n2126_, G63gat );
or g2056 ( new_n2128_, new_n2127_, new_n2039_ );
or g2057 ( new_n2129_, new_n1994_, G69gat );
and g2058 ( new_n2130_, new_n2128_, new_n2129_ );
or g2059 ( new_n2131_, new_n2130_, new_n2048_ );
and g2060 ( new_n2132_, new_n2060_, new_n2131_ );
or g2061 ( new_n2133_, new_n2132_, new_n2124_ );
and g2062 ( new_n2134_, new_n2123_, new_n2133_ );
and g2063 ( new_n2135_, new_n2134_, G40gat );
or g2064 ( new_n2136_, new_n2096_, new_n187_ );
or g2065 ( new_n2137_, new_n2063_, new_n186_ );
and g2066 ( new_n2138_, new_n1934_, new_n179_ );
or g2067 ( new_n2139_, new_n1989_, new_n2138_ );
and g2068 ( new_n2140_, new_n2139_, new_n183_ );
or g2069 ( new_n2141_, new_n2137_, new_n2140_ );
and g2070 ( new_n2142_, new_n2136_, new_n2141_ );
and g2071 ( new_n2143_, new_n2142_, new_n639_ );
or g2072 ( new_n2144_, new_n2135_, new_n2143_ );
and g2073 ( new_n2145_, new_n2144_, new_n316_ );
or g2074 ( new_n2146_, new_n2120_, new_n2145_ );
and g2075 ( new_n2147_, new_n2146_, G24gat );
and g2076 ( new_n2148_, new_n2008_, new_n943_ );
or g2077 ( new_n2149_, new_n2148_, new_n2004_ );
and g2078 ( new_n2150_, new_n2149_, G66gat );
or g2079 ( new_n2151_, new_n2150_, new_n2012_ );
and g2080 ( new_n2152_, new_n2151_, G60gat );
or g2081 ( new_n2153_, new_n2152_, new_n2023_ );
and g2082 ( new_n2154_, new_n2153_, new_n182_ );
and g2083 ( new_n2155_, new_n2149_, new_n183_ );
or g2084 ( new_n2156_, new_n2155_, new_n931_ );
or g2085 ( new_n2157_, new_n2154_, new_n2156_ );
or g2086 ( new_n2158_, new_n2088_, new_n320_ );
and g2087 ( new_n2159_, new_n2158_, new_n2095_ );
or g2088 ( new_n2160_, new_n2159_, new_n187_ );
and g2089 ( new_n2161_, new_n2157_, new_n2160_ );
and g2090 ( new_n2162_, new_n2161_, G40gat );
or g2091 ( new_n2163_, new_n2022_, new_n300_ );
or g2092 ( new_n2164_, new_n2017_, new_n282_ );
and g2093 ( new_n2165_, new_n2164_, new_n2010_ );
or g2094 ( new_n2166_, new_n2165_, new_n299_ );
and g2095 ( new_n2167_, new_n2166_, new_n322_ );
and g2096 ( new_n2168_, new_n2163_, new_n2167_ );
and g2097 ( new_n2169_, new_n2094_, new_n321_ );
or g2098 ( new_n2170_, new_n2168_, new_n2169_ );
and g2099 ( new_n2171_, new_n2170_, new_n639_ );
or g2100 ( new_n2172_, new_n2162_, new_n2171_ );
and g2101 ( new_n2173_, new_n2172_, G34gat );
and g2102 ( new_n2174_, new_n627_, new_n578_ );
or g2103 ( new_n2175_, new_n2020_, new_n677_ );
or g2104 ( new_n2176_, new_n2175_, new_n2174_ );
and g2105 ( new_n2177_, new_n2176_, G40gat );
and g2106 ( new_n2178_, new_n2177_, new_n316_ );
or g2107 ( new_n2179_, new_n2173_, new_n2178_ );
and g2108 ( new_n2180_, new_n2179_, new_n189_ );
or g2109 ( new_n2181_, new_n2147_, new_n2180_ );
and g2110 ( new_n2182_, new_n2181_, G30gat );
and g2111 ( new_n2183_, new_n2101_, new_n307_ );
or g2112 ( new_n2184_, new_n2182_, new_n2183_ );
and g2113 ( new_n2185_, new_n2184_, new_n701_ );
and g2114 ( new_n2186_, new_n115_, G95gat );
and g2115 ( new_n2187_, new_n111_, new_n160_ );
or g2116 ( new_n2188_, new_n2186_, new_n2187_ );
and g2117 ( new_n2189_, new_n2188_, G92gat );
or g2118 ( new_n2190_, new_n2189_, new_n1869_ );
and g2119 ( new_n2191_, new_n2190_, G86gat );
or g2120 ( new_n2192_, new_n2191_, new_n1881_ );
and g2121 ( new_n2193_, new_n2192_, G76gat );
or g2122 ( new_n2194_, new_n2193_, new_n1894_ );
and g2123 ( new_n2195_, new_n2194_, G82gat );
and g2124 ( new_n2196_, new_n2188_, new_n251_ );
or g2125 ( new_n2197_, new_n2195_, new_n2196_ );
and g2126 ( new_n2198_, new_n2197_, G79gat );
or g2127 ( new_n2199_, new_n2198_, new_n1914_ );
and g2128 ( new_n2200_, new_n2199_, G73gat );
or g2129 ( new_n2201_, new_n2200_, new_n1938_ );
and g2130 ( new_n2202_, new_n2201_, G63gat );
or g2131 ( new_n2203_, new_n2202_, new_n1961_ );
and g2132 ( new_n2204_, new_n2203_, G69gat );
and g2133 ( new_n2205_, new_n2197_, new_n265_ );
or g2134 ( new_n2206_, new_n2204_, new_n2205_ );
and g2135 ( new_n2207_, new_n2206_, G66gat );
or g2136 ( new_n2208_, new_n2207_, new_n1973_ );
and g2137 ( new_n2209_, new_n2208_, G60gat );
or g2138 ( new_n2210_, new_n2209_, new_n1999_ );
and g2139 ( new_n2211_, new_n2210_, G50gat );
or g2140 ( new_n2212_, new_n2211_, new_n2025_ );
and g2141 ( new_n2213_, new_n2212_, G56gat );
and g2142 ( new_n2214_, new_n2206_, new_n272_ );
or g2143 ( new_n2215_, new_n2213_, new_n2214_ );
and g2144 ( new_n2216_, new_n2215_, G53gat );
or g2145 ( new_n2217_, new_n2216_, new_n2045_ );
and g2146 ( new_n2218_, new_n2217_, G47gat );
or g2147 ( new_n2219_, new_n2218_, new_n2070_ );
and g2148 ( new_n2220_, new_n2219_, G37gat );
or g2149 ( new_n2221_, new_n2220_, new_n2097_ );
and g2150 ( new_n2222_, new_n2221_, G43gat );
and g2151 ( new_n2223_, new_n2215_, new_n290_ );
or g2152 ( new_n2224_, new_n2222_, new_n2223_ );
and g2153 ( new_n2225_, new_n2224_, new_n864_ );
and g2154 ( new_n2226_, new_n2118_, G34gat );
or g2155 ( new_n2227_, new_n2226_, new_n2145_ );
and g2156 ( new_n2228_, new_n2227_, G24gat );
or g2157 ( new_n2229_, new_n2228_, new_n2180_ );
and g2158 ( new_n2230_, new_n2229_, G30gat );
or g2159 ( new_n2231_, new_n2225_, new_n2230_ );
and g2160 ( new_n2232_, new_n2231_, G14gat );
or g2161 ( new_n2233_, new_n2185_, new_n2232_ );
and g2162 ( new_n2234_, new_n2233_, G27gat );
or g2163 ( new_n2235_, new_n2144_, new_n318_ );
or g2164 ( new_n2236_, new_n2179_, G24gat );
and g2165 ( new_n2237_, new_n2235_, new_n2236_ );
or g2166 ( new_n2238_, new_n2237_, new_n307_ );
and g2167 ( new_n2239_, new_n2070_, G37gat );
or g2168 ( new_n2240_, new_n2239_, new_n2097_ );
and g2169 ( new_n2241_, new_n2240_, G43gat );
and g2170 ( new_n2242_, new_n2044_, new_n292_ );
or g2171 ( new_n2243_, new_n2242_, new_n310_ );
or g2172 ( new_n2244_, new_n2241_, new_n2243_ );
and g2173 ( new_n2245_, new_n2244_, new_n690_ );
and g2174 ( new_n2246_, new_n2238_, new_n2245_ );
or g2175 ( new_n2247_, new_n2234_, new_n2246_ );
and g2176 ( new_n2248_, new_n2247_, G21gat );
not g2177 ( new_n2249_, new_n1186_ );
or g2178 ( new_n2250_, new_n2142_, new_n2249_ );
and g2179 ( new_n2251_, new_n2250_, new_n2236_ );
or g2180 ( new_n2252_, new_n2251_, new_n307_ );
and g2181 ( new_n2253_, new_n2121_, new_n676_ );
or g2182 ( new_n2254_, new_n2097_, new_n2253_ );
and g2183 ( new_n2255_, new_n2254_, G43gat );
and g2184 ( new_n2256_, new_n2061_, new_n894_ );
or g2185 ( new_n2257_, new_n2256_, new_n886_ );
or g2186 ( new_n2258_, new_n2255_, new_n2257_ );
and g2187 ( new_n2259_, new_n2258_, G27gat );
and g2188 ( new_n2260_, new_n2252_, new_n2259_ );
or g2189 ( new_n2261_, new_n2137_, new_n2066_ );
and g2190 ( new_n2262_, new_n2136_, new_n2261_ );
or g2191 ( new_n2263_, new_n2262_, new_n190_ );
or g2192 ( new_n2264_, new_n2236_, new_n307_ );
and g2193 ( new_n2265_, new_n2264_, new_n690_ );
and g2194 ( new_n2266_, new_n2263_, new_n2265_ );
or g2195 ( new_n2267_, new_n2260_, new_n2266_ );
and g2196 ( new_n2268_, new_n2267_, new_n337_ );
or g2197 ( new_n2269_, new_n2248_, new_n2268_ );
and g2198 ( new_n2270_, new_n2269_, G8gat );
and g2199 ( new_n2271_, new_n2144_, new_n317_ );
or g2200 ( new_n2272_, new_n2271_, new_n2180_ );
and g2201 ( new_n2273_, new_n2272_, G30gat );
and g2202 ( new_n2274_, new_n2117_, new_n309_ );
or g2203 ( new_n2275_, new_n2273_, new_n2274_ );
and g2204 ( new_n2276_, new_n2275_, G14gat );
and g2205 ( new_n2277_, new_n2143_, new_n317_ );
or g2206 ( new_n2278_, new_n2277_, new_n2180_ );
and g2207 ( new_n2279_, new_n2278_, G30gat );
and g2208 ( new_n2280_, new_n2134_, new_n887_ );
or g2209 ( new_n2281_, new_n2279_, new_n2280_ );
and g2210 ( new_n2282_, new_n2281_, new_n701_ );
or g2211 ( new_n2283_, new_n2276_, new_n2282_ );
and g2212 ( new_n2284_, new_n2283_, G21gat );
and g2213 ( new_n2285_, new_n2281_, G27gat );
or g2214 ( new_n2286_, new_n2285_, new_n2266_ );
and g2215 ( new_n2287_, new_n2286_, new_n701_ );
and g2216 ( new_n2288_, new_n2267_, G14gat );
or g2217 ( new_n2289_, new_n2287_, new_n2288_ );
and g2218 ( new_n2290_, new_n2289_, new_n337_ );
or g2219 ( new_n2291_, new_n2284_, new_n2290_ );
and g2220 ( new_n2292_, new_n2291_, new_n352_ );
or g2221 ( new_n2293_, new_n2270_, new_n2292_ );
and g2222 ( new_n2294_, new_n2293_, G11gat );
or g2223 ( new_n2295_, new_n2081_, new_n931_ );
and g2224 ( new_n2296_, new_n2160_, new_n937_ );
and g2225 ( new_n2297_, new_n2295_, new_n2296_ );
and g2226 ( new_n2298_, new_n2171_, G34gat );
or g2227 ( new_n2299_, new_n2298_, new_n2178_ );
and g2228 ( new_n2300_, new_n2299_, new_n190_ );
or g2229 ( new_n2301_, new_n2297_, new_n2300_ );
and g2230 ( new_n2302_, new_n2301_, G27gat );
and g2231 ( new_n2303_, new_n2087_, new_n322_ );
or g2232 ( new_n2304_, new_n2303_, new_n2169_ );
and g2233 ( new_n2305_, new_n2304_, new_n344_ );
and g2234 ( new_n2306_, new_n2177_, new_n343_ );
or g2235 ( new_n2307_, new_n2305_, new_n2306_ );
and g2236 ( new_n2308_, new_n2307_, new_n690_ );
or g2237 ( new_n2309_, new_n2302_, new_n2308_ );
and g2238 ( new_n2310_, new_n2309_, G21gat );
or g2239 ( new_n2311_, new_n2093_, new_n677_ );
and g2240 ( new_n2312_, new_n2311_, new_n744_ );
or g2241 ( new_n2313_, new_n2312_, new_n690_ );
and g2242 ( new_n2314_, new_n2313_, new_n337_ );
or g2243 ( new_n2315_, new_n2310_, new_n2314_ );
and g2244 ( new_n2316_, new_n2315_, new_n193_ );
or g2245 ( new_n2317_, new_n2294_, new_n2316_ );
and g2246 ( new_n2318_, new_n2317_, G17gat );
and g2247 ( new_n2319_, new_n2036_, new_n490_ );
or g2248 ( new_n2320_, new_n2319_, new_n1938_ );
and g2249 ( new_n2321_, new_n2320_, G63gat );
or g2250 ( new_n2322_, new_n2321_, new_n1961_ );
and g2251 ( new_n2323_, new_n2322_, G69gat );
and g2252 ( new_n2324_, new_n2186_, new_n251_ );
or g2253 ( new_n2325_, new_n1896_, new_n2324_ );
and g2254 ( new_n2326_, new_n2325_, new_n854_ );
or g2255 ( new_n2327_, new_n2323_, new_n2326_ );
and g2256 ( new_n2328_, new_n2327_, G66gat );
or g2257 ( new_n2329_, new_n2328_, new_n1973_ );
and g2258 ( new_n2330_, new_n2329_, G60gat );
or g2259 ( new_n2331_, new_n2330_, new_n1999_ );
and g2260 ( new_n2332_, new_n2331_, G50gat );
or g2261 ( new_n2333_, new_n2332_, new_n2025_ );
and g2262 ( new_n2334_, new_n2333_, G56gat );
and g2263 ( new_n2335_, new_n2325_, new_n265_ );
or g2264 ( new_n2336_, new_n2204_, new_n2335_ );
and g2265 ( new_n2337_, new_n2336_, new_n272_ );
or g2266 ( new_n2338_, new_n2334_, new_n2337_ );
and g2267 ( new_n2339_, new_n2338_, new_n290_ );
or g2268 ( new_n2340_, new_n2222_, new_n2339_ );
and g2269 ( new_n2341_, new_n2340_, new_n307_ );
or g2270 ( new_n2342_, new_n2182_, new_n2341_ );
and g2271 ( new_n2343_, new_n2342_, G14gat );
or g2272 ( new_n2344_, new_n2185_, new_n2343_ );
and g2273 ( new_n2345_, new_n2344_, G8gat );
and g2274 ( new_n2346_, new_n2283_, new_n352_ );
or g2275 ( new_n2347_, new_n2345_, new_n2346_ );
and g2276 ( new_n2348_, new_n2347_, new_n331_ );
or g2277 ( new_n2349_, new_n2318_, new_n2348_ );
and g2278 ( new_n2350_, new_n2349_, G1gat );
and g2279 ( new_n2351_, new_n2142_, new_n191_ );
and g2280 ( new_n2352_, new_n2180_, G30gat );
or g2281 ( new_n2353_, new_n2352_, new_n701_ );
or g2282 ( new_n2354_, new_n2351_, new_n2353_ );
and g2283 ( new_n2355_, new_n2161_, new_n937_ );
or g2284 ( new_n2356_, new_n2355_, new_n2300_ );
or g2285 ( new_n2357_, new_n2356_, G14gat );
and g2286 ( new_n2358_, new_n2354_, new_n2357_ );
or g2287 ( new_n2359_, new_n2358_, new_n352_ );
and g2288 ( new_n2360_, new_n2170_, new_n344_ );
or g2289 ( new_n2361_, new_n2360_, new_n2306_ );
and g2290 ( new_n2362_, new_n2361_, G14gat );
and g2291 ( new_n2363_, new_n2176_, new_n1286_ );
or g2292 ( new_n2364_, new_n2362_, new_n2363_ );
or g2293 ( new_n2365_, new_n2364_, G8gat );
and g2294 ( new_n2366_, new_n2359_, new_n2365_ );
or g2295 ( new_n2367_, new_n2366_, new_n194_ );
and g2296 ( new_n2368_, new_n2309_, G14gat );
and g2297 ( new_n2369_, new_n2356_, G27gat );
or g2298 ( new_n2370_, new_n2369_, new_n2308_ );
and g2299 ( new_n2371_, new_n2370_, new_n701_ );
or g2300 ( new_n2372_, new_n2368_, new_n2371_ );
and g2301 ( new_n2373_, new_n2372_, G21gat );
or g2302 ( new_n2374_, new_n2314_, new_n352_ );
or g2303 ( new_n2375_, new_n2373_, new_n2374_ );
and g2304 ( new_n2376_, new_n2364_, G21gat );
and g2305 ( new_n2377_, new_n2312_, G14gat );
or g2306 ( new_n2378_, new_n2363_, new_n690_ );
or g2307 ( new_n2379_, new_n2377_, new_n2378_ );
and g2308 ( new_n2380_, new_n2379_, new_n337_ );
or g2309 ( new_n2381_, new_n2380_, G8gat );
or g2310 ( new_n2382_, new_n2376_, new_n2381_ );
and g2311 ( new_n2383_, new_n2375_, new_n2382_ );
or g2312 ( new_n2384_, new_n2383_, new_n195_ );
and g2313 ( new_n2385_, new_n2384_, new_n356_ );
and g2314 ( new_n2386_, new_n2367_, new_n2385_ );
or g2315 ( new_n2387_, new_n2350_, new_n2386_ );
and g2316 ( new_n2388_, new_n2387_, G4gat );
and g2317 ( new_n2389_, new_n2231_, G27gat );
or g2318 ( new_n2390_, new_n2389_, new_n2246_ );
and g2319 ( new_n2391_, new_n2390_, G21gat );
or g2320 ( new_n2392_, new_n2391_, new_n2268_ );
and g2321 ( new_n2393_, new_n2392_, G11gat );
or g2322 ( new_n2394_, new_n2393_, new_n2316_ );
and g2323 ( new_n2395_, new_n2394_, G17gat );
and g2324 ( new_n2396_, new_n2342_, new_n331_ );
or g2325 ( new_n2397_, new_n2395_, new_n2396_ );
and g2326 ( new_n2398_, new_n2397_, new_n196_ );
or g2327 ( new_n2399_, new_n2388_, new_n2398_ );
and g2328 ( new_n2400_, new_n2399_, keyinput2_G432gat );
not g2329 ( new_n2401_, keyinput2_G432gat );
and g2330 ( new_n2402_, new_n111_, new_n2401_ );
or g2331 ( new_n2403_, new_n2400_, new_n2402_ );
and g2332 ( new_n2404_, new_n2403_, keyinput3_G432gat );
not g2333 ( new_n2405_, keyinput3_G432gat );
not g2334 ( new_n2406_, new_n188_ );
and g2335 ( new_n2407_, new_n2406_, new_n2401_ );
and g2336 ( new_n2408_, new_n218_, keyinput2_G432gat );
or g2337 ( new_n2409_, new_n2407_, new_n2408_ );
and g2338 ( new_n2410_, new_n2409_, new_n2405_ );
or g2339 ( new_n2411_, new_n2404_, new_n2410_ );
and g2340 ( new_n2412_, new_n2411_, keyinput1_G432gat );
not g2341 ( new_n2413_, keyinput1_G432gat );
and g2342 ( new_n2414_, new_n140_, new_n2401_ );
and g2343 ( new_n2415_, new_n102_, keyinput2_G432gat );
or g2344 ( new_n2416_, new_n2414_, new_n2415_ );
and g2345 ( new_n2417_, new_n2416_, keyinput3_G432gat );
and g2346 ( new_n2418_, new_n852_, new_n2401_ );
and g2347 ( new_n2419_, new_n856_, new_n2418_ );
and g2348 ( new_n2420_, new_n941_, keyinput2_G432gat );
or g2349 ( new_n2421_, new_n2419_, new_n2420_ );
and g2350 ( new_n2422_, new_n218_, new_n2405_ );
and g2351 ( new_n2423_, new_n2421_, new_n2422_ );
or g2352 ( new_n2424_, new_n2417_, new_n2423_ );
and g2353 ( new_n2425_, new_n2424_, new_n2413_ );
or g2354 ( new_n2426_, new_n2412_, new_n2425_ );
and g2355 ( new_n2427_, new_n2426_, keyinput0_G432gat );
not g2356 ( new_n2428_, keyinput0_G432gat );
and g2357 ( new_n2429_, new_n192_, G11gat );
not g2358 ( new_n2430_, new_n2429_ );
and g2359 ( new_n2431_, new_n2430_, new_n2401_ );
and g2360 ( new_n2432_, new_n184_, G37gat );
not g2361 ( new_n2433_, new_n2432_ );
and g2362 ( new_n2434_, new_n2433_, keyinput2_G432gat );
or g2363 ( new_n2435_, new_n2431_, new_n2434_ );
and g2364 ( new_n2436_, new_n2435_, new_n2405_ );
or g2365 ( new_n2437_, new_n177_, keyinput2_G432gat );
or g2366 ( new_n2438_, new_n803_, new_n2437_ );
and g2367 ( new_n2439_, new_n87_, keyinput2_G432gat );
not g2368 ( new_n2440_, new_n2439_ );
and g2369 ( new_n2441_, new_n2440_, keyinput3_G432gat );
and g2370 ( new_n2442_, new_n2438_, new_n2441_ );
or g2371 ( new_n2443_, new_n2436_, new_n2442_ );
and g2372 ( new_n2444_, new_n2443_, new_n2413_ );
and g2373 ( new_n2445_, new_n145_, new_n2401_ );
or g2374 ( new_n2446_, new_n2445_, new_n2439_ );
and g2375 ( new_n2447_, new_n2446_, new_n2405_ );
and g2376 ( new_n2448_, new_n112_, new_n2401_ );
and g2377 ( new_n2449_, G108gat, keyinput2_G432gat );
or g2378 ( new_n2450_, new_n2448_, new_n2449_ );
and g2379 ( new_n2451_, new_n2450_, keyinput3_G432gat );
or g2380 ( new_n2452_, new_n2447_, new_n2451_ );
and g2381 ( new_n2453_, new_n2452_, keyinput1_G432gat );
or g2382 ( new_n2454_, new_n2444_, new_n2453_ );
and g2383 ( new_n2455_, new_n2454_, new_n2428_ );
or g2384 ( G432gat, new_n2427_, new_n2455_ );
endmodule