module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n955_, new_n608_, new_n888_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n401_, new_n389_, new_n514_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n342_, new_n649_, new_n706_, new_n462_, new_n761_, new_n752_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n890_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n935_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n528_, new_n952_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n948_, new_n762_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n851_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n555_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n756_, new_n495_, new_n823_, new_n431_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n947_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n889_, new_n229_, new_n536_, new_n464_, new_n204_, new_n573_, new_n765_, new_n405_;

xor g000 ( new_n202_, N81, N85 );
xnor g001 ( new_n203_, new_n202_, keyIn_0_10 );
xnor g002 ( new_n204_, N89, N93 );
xnor g003 ( new_n205_, new_n204_, keyIn_0_11 );
xnor g004 ( new_n206_, new_n203_, new_n205_ );
xnor g005 ( new_n207_, new_n206_, keyIn_0_33 );
xnor g006 ( new_n208_, N65, N69 );
xnor g007 ( new_n209_, new_n208_, keyIn_0_8 );
xnor g008 ( new_n210_, N73, N77 );
xnor g009 ( new_n211_, new_n210_, keyIn_0_9 );
xnor g010 ( new_n212_, new_n209_, new_n211_ );
xnor g011 ( new_n213_, new_n212_, keyIn_0_32 );
xnor g012 ( new_n214_, new_n207_, new_n213_ );
or g013 ( new_n215_, new_n214_, keyIn_0_43 );
nand g014 ( new_n216_, new_n214_, keyIn_0_43 );
nand g015 ( new_n217_, N129, N137 );
nand g016 ( new_n218_, new_n215_, new_n216_, new_n217_ );
nand g017 ( new_n219_, new_n215_, new_n216_ );
not g018 ( new_n220_, new_n217_ );
nand g019 ( new_n221_, new_n219_, new_n220_ );
nand g020 ( new_n222_, new_n221_, new_n218_ );
nand g021 ( new_n223_, new_n222_, keyIn_0_47 );
not g022 ( new_n224_, keyIn_0_47 );
nand g023 ( new_n225_, new_n221_, new_n224_, new_n218_ );
xnor g024 ( new_n226_, N1, N17 );
xnor g025 ( new_n227_, N33, N49 );
xnor g026 ( new_n228_, new_n226_, new_n227_ );
nand g027 ( new_n229_, new_n223_, new_n225_, new_n228_ );
nand g028 ( new_n230_, new_n223_, new_n225_ );
not g029 ( new_n231_, new_n228_ );
nand g030 ( new_n232_, new_n230_, new_n231_ );
nand g031 ( new_n233_, new_n232_, keyIn_0_55, new_n229_ );
not g032 ( new_n234_, keyIn_0_55 );
nand g033 ( new_n235_, new_n232_, new_n229_ );
nand g034 ( new_n236_, new_n235_, new_n234_ );
nand g035 ( new_n237_, new_n236_, new_n233_ );
not g036 ( new_n238_, new_n237_ );
not g037 ( new_n239_, keyIn_0_56 );
xnor g038 ( new_n240_, N97, N101 );
xnor g039 ( new_n241_, new_n240_, keyIn_0_12 );
xnor g040 ( new_n242_, N105, N109 );
xnor g041 ( new_n243_, new_n242_, keyIn_0_13 );
xnor g042 ( new_n244_, new_n241_, new_n243_ );
xnor g043 ( new_n245_, new_n244_, keyIn_0_34 );
xnor g044 ( new_n246_, N121, N125 );
xnor g045 ( new_n247_, new_n246_, keyIn_0_15 );
xnor g046 ( new_n248_, N113, N117 );
xnor g047 ( new_n249_, new_n248_, keyIn_0_14 );
xnor g048 ( new_n250_, new_n247_, new_n249_ );
xnor g049 ( new_n251_, new_n250_, keyIn_0_35 );
xnor g050 ( new_n252_, new_n245_, new_n251_ );
nand g051 ( new_n253_, new_n252_, keyIn_0_44 );
not g052 ( new_n254_, keyIn_0_44 );
nand g053 ( new_n255_, new_n245_, new_n251_ );
or g054 ( new_n256_, new_n245_, new_n251_ );
nand g055 ( new_n257_, new_n256_, new_n254_, new_n255_ );
nand g056 ( new_n258_, N130, N137 );
nand g057 ( new_n259_, new_n253_, new_n257_, new_n258_ );
nand g058 ( new_n260_, new_n253_, new_n257_ );
nand g059 ( new_n261_, new_n260_, N130, N137 );
nand g060 ( new_n262_, new_n261_, new_n259_ );
nand g061 ( new_n263_, new_n262_, keyIn_0_48 );
not g062 ( new_n264_, keyIn_0_48 );
nand g063 ( new_n265_, new_n261_, new_n264_, new_n259_ );
xnor g064 ( new_n266_, N5, N21 );
xnor g065 ( new_n267_, N37, N53 );
xnor g066 ( new_n268_, new_n266_, new_n267_ );
nand g067 ( new_n269_, new_n263_, new_n265_, new_n268_ );
nand g068 ( new_n270_, new_n263_, new_n265_ );
not g069 ( new_n271_, new_n268_ );
nand g070 ( new_n272_, new_n270_, new_n271_ );
nand g071 ( new_n273_, new_n272_, new_n239_, new_n269_ );
nand g072 ( new_n274_, new_n272_, new_n269_ );
nand g073 ( new_n275_, new_n274_, keyIn_0_56 );
nand g074 ( new_n276_, new_n275_, new_n273_ );
not g075 ( new_n277_, keyIn_0_50 );
not g076 ( new_n278_, keyIn_0_46 );
nand g077 ( new_n279_, new_n207_, new_n251_ );
or g078 ( new_n280_, new_n207_, new_n251_ );
nand g079 ( new_n281_, new_n280_, new_n278_, new_n279_ );
nand g080 ( new_n282_, new_n280_, new_n279_ );
nand g081 ( new_n283_, new_n282_, keyIn_0_46 );
nand g082 ( new_n284_, new_n283_, new_n281_ );
nand g083 ( new_n285_, N132, N137 );
not g084 ( new_n286_, new_n285_ );
nand g085 ( new_n287_, new_n284_, new_n286_ );
nand g086 ( new_n288_, new_n283_, new_n281_, new_n285_ );
nand g087 ( new_n289_, new_n287_, new_n277_, new_n288_ );
nand g088 ( new_n290_, new_n287_, new_n288_ );
nand g089 ( new_n291_, new_n290_, keyIn_0_50 );
nand g090 ( new_n292_, new_n291_, new_n289_ );
xor g091 ( new_n293_, N13, N29 );
xnor g092 ( new_n294_, new_n293_, keyIn_0_23 );
xnor g093 ( new_n295_, N45, N61 );
xnor g094 ( new_n296_, new_n294_, new_n295_ );
not g095 ( new_n297_, new_n296_ );
nand g096 ( new_n298_, new_n292_, new_n297_ );
nand g097 ( new_n299_, new_n291_, new_n289_, new_n296_ );
nand g098 ( new_n300_, new_n298_, keyIn_0_58, new_n299_ );
not g099 ( new_n301_, keyIn_0_58 );
nand g100 ( new_n302_, new_n298_, new_n299_ );
nand g101 ( new_n303_, new_n302_, new_n301_ );
nand g102 ( new_n304_, new_n303_, new_n300_ );
not g103 ( new_n305_, keyIn_0_45 );
xnor g104 ( new_n306_, new_n213_, new_n245_ );
xnor g105 ( new_n307_, new_n306_, new_n305_ );
nand g106 ( new_n308_, N131, N137 );
xor g107 ( new_n309_, new_n308_, keyIn_0_16 );
not g108 ( new_n310_, new_n309_ );
nand g109 ( new_n311_, new_n307_, new_n310_ );
or g110 ( new_n312_, new_n306_, new_n305_ );
nand g111 ( new_n313_, new_n306_, new_n305_ );
nand g112 ( new_n314_, new_n312_, new_n313_, new_n309_ );
nand g113 ( new_n315_, new_n311_, new_n314_ );
nand g114 ( new_n316_, new_n315_, keyIn_0_49 );
not g115 ( new_n317_, keyIn_0_49 );
nand g116 ( new_n318_, new_n311_, new_n317_, new_n314_ );
xor g117 ( new_n319_, N41, N57 );
xnor g118 ( new_n320_, new_n319_, keyIn_0_22 );
xnor g119 ( new_n321_, N9, N25 );
xnor g120 ( new_n322_, new_n321_, keyIn_0_21 );
xnor g121 ( new_n323_, new_n320_, new_n322_ );
xor g122 ( new_n324_, new_n323_, keyIn_0_36 );
nand g123 ( new_n325_, new_n316_, new_n318_, new_n324_ );
nand g124 ( new_n326_, new_n316_, new_n318_ );
not g125 ( new_n327_, new_n324_ );
nand g126 ( new_n328_, new_n326_, new_n327_ );
nand g127 ( new_n329_, new_n328_, new_n325_ );
nand g128 ( new_n330_, new_n329_, keyIn_0_57 );
not g129 ( new_n331_, keyIn_0_57 );
nand g130 ( new_n332_, new_n328_, new_n331_, new_n325_ );
nand g131 ( new_n333_, new_n330_, new_n332_ );
nand g132 ( new_n334_, new_n333_, new_n276_, new_n304_ );
nand g133 ( new_n335_, new_n276_, new_n304_ );
and g134 ( new_n336_, new_n330_, new_n332_ );
nand g135 ( new_n337_, new_n335_, new_n336_ );
nand g136 ( new_n338_, new_n275_, new_n303_, new_n273_, new_n300_ );
nand g137 ( new_n339_, new_n337_, new_n237_, new_n334_, new_n338_ );
not g138 ( new_n340_, keyIn_0_63 );
nand g139 ( new_n341_, new_n330_, new_n340_, new_n332_ );
nand g140 ( new_n342_, new_n333_, keyIn_0_63 );
nand g141 ( new_n343_, new_n342_, new_n341_ );
and g142 ( new_n344_, new_n233_, new_n276_, new_n304_, new_n236_ );
nand g143 ( new_n345_, new_n343_, new_n344_ );
nand g144 ( new_n346_, new_n339_, new_n345_ );
not g145 ( new_n347_, keyIn_0_62 );
not g146 ( new_n348_, keyIn_0_42 );
not g147 ( new_n349_, N61 );
nand g148 ( new_n350_, new_n349_, N57 );
not g149 ( new_n351_, N57 );
nand g150 ( new_n352_, new_n351_, N61 );
nand g151 ( new_n353_, new_n350_, new_n352_ );
nand g152 ( new_n354_, new_n353_, keyIn_0_7 );
not g153 ( new_n355_, keyIn_0_7 );
nand g154 ( new_n356_, new_n350_, new_n352_, new_n355_ );
nand g155 ( new_n357_, new_n354_, new_n356_ );
not g156 ( new_n358_, keyIn_0_6 );
nand g157 ( new_n359_, N49, N53 );
or g158 ( new_n360_, N49, N53 );
nand g159 ( new_n361_, new_n360_, new_n359_ );
nand g160 ( new_n362_, new_n361_, new_n358_ );
nand g161 ( new_n363_, new_n360_, keyIn_0_6, new_n359_ );
nand g162 ( new_n364_, new_n362_, new_n363_ );
nand g163 ( new_n365_, new_n364_, new_n357_ );
nand g164 ( new_n366_, new_n362_, new_n354_, new_n356_, new_n363_ );
nand g165 ( new_n367_, new_n365_, keyIn_0_31, new_n366_ );
not g166 ( new_n368_, keyIn_0_31 );
nand g167 ( new_n369_, new_n365_, new_n366_ );
nand g168 ( new_n370_, new_n369_, new_n368_ );
not g169 ( new_n371_, keyIn_0_29 );
not g170 ( new_n372_, N21 );
nand g171 ( new_n373_, new_n372_, N17 );
not g172 ( new_n374_, N17 );
nand g173 ( new_n375_, new_n374_, N21 );
nand g174 ( new_n376_, new_n373_, new_n375_ );
nand g175 ( new_n377_, new_n376_, keyIn_0_2 );
not g176 ( new_n378_, keyIn_0_2 );
nand g177 ( new_n379_, new_n373_, new_n375_, new_n378_ );
nand g178 ( new_n380_, new_n377_, new_n379_ );
nand g179 ( new_n381_, N25, N29 );
or g180 ( new_n382_, N25, N29 );
nand g181 ( new_n383_, new_n382_, new_n381_ );
nand g182 ( new_n384_, new_n383_, keyIn_0_3 );
not g183 ( new_n385_, keyIn_0_3 );
nand g184 ( new_n386_, new_n382_, new_n385_, new_n381_ );
nand g185 ( new_n387_, new_n384_, new_n386_ );
nand g186 ( new_n388_, new_n387_, new_n380_ );
nand g187 ( new_n389_, new_n384_, new_n377_, new_n379_, new_n386_ );
nand g188 ( new_n390_, new_n388_, new_n371_, new_n389_ );
nand g189 ( new_n391_, new_n388_, new_n389_ );
nand g190 ( new_n392_, new_n391_, keyIn_0_29 );
nand g191 ( new_n393_, new_n370_, new_n392_, new_n367_, new_n390_ );
nand g192 ( new_n394_, new_n370_, new_n367_ );
nand g193 ( new_n395_, new_n392_, new_n390_ );
nand g194 ( new_n396_, new_n394_, new_n395_ );
nand g195 ( new_n397_, new_n396_, new_n348_, new_n393_ );
nand g196 ( new_n398_, new_n396_, new_n393_ );
nand g197 ( new_n399_, new_n398_, keyIn_0_42 );
nand g198 ( new_n400_, N136, N137 );
xnor g199 ( new_n401_, new_n400_, keyIn_0_20 );
nand g200 ( new_n402_, new_n399_, new_n397_, new_n401_ );
nand g201 ( new_n403_, new_n399_, new_n397_ );
not g202 ( new_n404_, new_n401_ );
nand g203 ( new_n405_, new_n403_, new_n404_ );
nand g204 ( new_n406_, new_n405_, new_n402_ );
nand g205 ( new_n407_, new_n406_, keyIn_0_54 );
not g206 ( new_n408_, keyIn_0_54 );
nand g207 ( new_n409_, new_n405_, new_n408_, new_n402_ );
xnor g208 ( new_n410_, N77, N93 );
xnor g209 ( new_n411_, N109, N125 );
xnor g210 ( new_n412_, new_n410_, new_n411_ );
nand g211 ( new_n413_, new_n407_, new_n409_, new_n412_ );
nand g212 ( new_n414_, new_n407_, new_n409_ );
not g213 ( new_n415_, new_n412_ );
nand g214 ( new_n416_, new_n414_, new_n415_ );
nand g215 ( new_n417_, new_n416_, new_n347_, new_n413_ );
nand g216 ( new_n418_, new_n416_, new_n413_ );
nand g217 ( new_n419_, new_n418_, keyIn_0_62 );
and g218 ( new_n420_, new_n419_, new_n417_ );
not g219 ( new_n421_, keyIn_0_61 );
not g220 ( new_n422_, keyIn_0_4 );
not g221 ( new_n423_, N33 );
not g222 ( new_n424_, N37 );
nand g223 ( new_n425_, new_n423_, new_n424_ );
nand g224 ( new_n426_, N33, N37 );
nand g225 ( new_n427_, new_n425_, new_n426_ );
nand g226 ( new_n428_, new_n427_, new_n422_ );
nand g227 ( new_n429_, new_n425_, keyIn_0_4, new_n426_ );
nand g228 ( new_n430_, new_n428_, new_n429_ );
not g229 ( new_n431_, keyIn_0_5 );
nand g230 ( new_n432_, N41, N45 );
not g231 ( new_n433_, N41 );
not g232 ( new_n434_, N45 );
nand g233 ( new_n435_, new_n433_, new_n434_ );
nand g234 ( new_n436_, new_n435_, new_n431_, new_n432_ );
xnor g235 ( new_n437_, N41, N45 );
nand g236 ( new_n438_, new_n437_, keyIn_0_5 );
nand g237 ( new_n439_, new_n438_, new_n436_ );
nand g238 ( new_n440_, new_n430_, new_n439_ );
nand g239 ( new_n441_, new_n428_, new_n438_, new_n429_, new_n436_ );
nand g240 ( new_n442_, new_n440_, keyIn_0_30, new_n441_ );
not g241 ( new_n443_, keyIn_0_30 );
nand g242 ( new_n444_, new_n440_, new_n441_ );
nand g243 ( new_n445_, new_n444_, new_n443_ );
nand g244 ( new_n446_, new_n445_, new_n442_ );
not g245 ( new_n447_, keyIn_0_0 );
nand g246 ( new_n448_, N1, N5 );
or g247 ( new_n449_, N1, N5 );
nand g248 ( new_n450_, new_n449_, new_n447_, new_n448_ );
nand g249 ( new_n451_, new_n449_, new_n448_ );
nand g250 ( new_n452_, new_n451_, keyIn_0_0 );
nand g251 ( new_n453_, new_n452_, new_n450_ );
not g252 ( new_n454_, keyIn_0_1 );
nand g253 ( new_n455_, N9, N13 );
or g254 ( new_n456_, N9, N13 );
nand g255 ( new_n457_, new_n456_, new_n454_, new_n455_ );
xnor g256 ( new_n458_, N9, N13 );
nand g257 ( new_n459_, new_n458_, keyIn_0_1 );
nand g258 ( new_n460_, new_n459_, new_n457_ );
nand g259 ( new_n461_, new_n453_, new_n460_ );
nand g260 ( new_n462_, new_n452_, new_n459_, new_n450_, new_n457_ );
nand g261 ( new_n463_, new_n461_, keyIn_0_28, new_n462_ );
not g262 ( new_n464_, keyIn_0_28 );
nand g263 ( new_n465_, new_n461_, new_n462_ );
nand g264 ( new_n466_, new_n465_, new_n464_ );
nand g265 ( new_n467_, new_n466_, new_n463_ );
nand g266 ( new_n468_, new_n446_, new_n467_ );
nand g267 ( new_n469_, new_n445_, new_n466_, new_n442_, new_n463_ );
nand g268 ( new_n470_, new_n468_, new_n469_ );
nand g269 ( new_n471_, new_n470_, keyIn_0_41 );
not g270 ( new_n472_, keyIn_0_41 );
nand g271 ( new_n473_, new_n468_, new_n472_, new_n469_ );
nand g272 ( new_n474_, new_n471_, new_n473_ );
nand g273 ( new_n475_, N135, N137 );
xor g274 ( new_n476_, new_n475_, keyIn_0_19 );
not g275 ( new_n477_, new_n476_ );
nand g276 ( new_n478_, new_n474_, new_n477_ );
nand g277 ( new_n479_, new_n471_, new_n473_, new_n476_ );
nand g278 ( new_n480_, new_n478_, new_n479_ );
nand g279 ( new_n481_, new_n480_, keyIn_0_53 );
not g280 ( new_n482_, keyIn_0_53 );
nand g281 ( new_n483_, new_n478_, new_n482_, new_n479_ );
nand g282 ( new_n484_, new_n481_, new_n483_ );
xor g283 ( new_n485_, N105, N121 );
xnor g284 ( new_n486_, new_n485_, keyIn_0_27 );
xnor g285 ( new_n487_, N73, N89 );
xnor g286 ( new_n488_, new_n487_, keyIn_0_26 );
xnor g287 ( new_n489_, new_n486_, new_n488_ );
xor g288 ( new_n490_, new_n489_, keyIn_0_38 );
not g289 ( new_n491_, new_n490_ );
nand g290 ( new_n492_, new_n484_, new_n491_ );
nand g291 ( new_n493_, new_n481_, new_n483_, new_n490_ );
nand g292 ( new_n494_, new_n492_, new_n493_ );
nand g293 ( new_n495_, new_n494_, new_n421_ );
nand g294 ( new_n496_, new_n492_, keyIn_0_61, new_n493_ );
nand g295 ( new_n497_, new_n495_, new_n496_ );
nor g296 ( new_n498_, new_n420_, new_n497_ );
not g297 ( new_n499_, keyIn_0_52 );
not g298 ( new_n500_, keyIn_0_40 );
nand g299 ( new_n501_, new_n394_, new_n446_ );
nand g300 ( new_n502_, new_n370_, new_n445_, new_n367_, new_n442_ );
nand g301 ( new_n503_, new_n501_, new_n500_, new_n502_ );
nand g302 ( new_n504_, new_n501_, new_n502_ );
nand g303 ( new_n505_, new_n504_, keyIn_0_40 );
nand g304 ( new_n506_, new_n505_, new_n503_ );
nand g305 ( new_n507_, N134, N137 );
xor g306 ( new_n508_, new_n507_, keyIn_0_18 );
not g307 ( new_n509_, new_n508_ );
nand g308 ( new_n510_, new_n506_, new_n509_ );
nand g309 ( new_n511_, new_n505_, new_n503_, new_n508_ );
nand g310 ( new_n512_, new_n510_, new_n499_, new_n511_ );
nand g311 ( new_n513_, new_n510_, new_n511_ );
nand g312 ( new_n514_, new_n513_, keyIn_0_52 );
nand g313 ( new_n515_, new_n514_, new_n512_ );
xor g314 ( new_n516_, N101, N117 );
xnor g315 ( new_n517_, new_n516_, keyIn_0_25 );
xnor g316 ( new_n518_, N69, N85 );
xnor g317 ( new_n519_, new_n518_, keyIn_0_24 );
xnor g318 ( new_n520_, new_n517_, new_n519_ );
xor g319 ( new_n521_, new_n520_, keyIn_0_37 );
not g320 ( new_n522_, new_n521_ );
nand g321 ( new_n523_, new_n515_, new_n522_ );
nand g322 ( new_n524_, new_n514_, new_n512_, new_n521_ );
nand g323 ( new_n525_, new_n523_, keyIn_0_60, new_n524_ );
not g324 ( new_n526_, keyIn_0_60 );
nand g325 ( new_n527_, new_n523_, new_n524_ );
nand g326 ( new_n528_, new_n527_, new_n526_ );
nand g327 ( new_n529_, new_n528_, new_n525_ );
nand g328 ( new_n530_, new_n395_, new_n467_ );
nand g329 ( new_n531_, new_n392_, new_n466_, new_n390_, new_n463_ );
nand g330 ( new_n532_, new_n530_, new_n531_ );
nand g331 ( new_n533_, new_n532_, keyIn_0_39 );
not g332 ( new_n534_, keyIn_0_39 );
nand g333 ( new_n535_, new_n530_, new_n534_, new_n531_ );
nand g334 ( new_n536_, new_n533_, new_n535_ );
nand g335 ( new_n537_, N133, N137 );
xnor g336 ( new_n538_, new_n537_, keyIn_0_17 );
not g337 ( new_n539_, new_n538_ );
nand g338 ( new_n540_, new_n536_, new_n539_ );
nand g339 ( new_n541_, new_n533_, new_n535_, new_n538_ );
nand g340 ( new_n542_, new_n540_, new_n541_ );
nand g341 ( new_n543_, new_n542_, keyIn_0_51 );
not g342 ( new_n544_, keyIn_0_51 );
nand g343 ( new_n545_, new_n540_, new_n544_, new_n541_ );
nand g344 ( new_n546_, new_n543_, new_n545_ );
xnor g345 ( new_n547_, N65, N81 );
xnor g346 ( new_n548_, N97, N113 );
xor g347 ( new_n549_, new_n547_, new_n548_ );
not g348 ( new_n550_, new_n549_ );
nand g349 ( new_n551_, new_n546_, new_n550_ );
nand g350 ( new_n552_, new_n543_, new_n545_, new_n549_ );
nand g351 ( new_n553_, new_n551_, keyIn_0_59, new_n552_ );
not g352 ( new_n554_, keyIn_0_59 );
nand g353 ( new_n555_, new_n551_, new_n552_ );
nand g354 ( new_n556_, new_n555_, new_n554_ );
nand g355 ( new_n557_, new_n556_, new_n553_ );
and g356 ( new_n558_, new_n529_, new_n557_ );
and g357 ( new_n559_, new_n346_, new_n498_, new_n558_ );
nand g358 ( new_n560_, new_n559_, new_n238_ );
xnor g359 ( N724, new_n560_, N1 );
not g360 ( new_n562_, new_n276_ );
nand g361 ( new_n563_, new_n559_, new_n562_ );
xnor g362 ( N725, new_n563_, N5 );
nand g363 ( new_n565_, new_n559_, new_n336_ );
xnor g364 ( N726, new_n565_, N9 );
not g365 ( new_n567_, new_n304_ );
nand g366 ( new_n568_, new_n559_, new_n567_ );
xnor g367 ( N727, new_n568_, N13 );
not g368 ( new_n570_, keyIn_0_105 );
nand g369 ( new_n571_, new_n419_, new_n417_ );
not g370 ( new_n572_, new_n497_ );
nor g371 ( new_n573_, new_n572_, new_n571_ );
nand g372 ( new_n574_, new_n346_, keyIn_0_76, new_n558_, new_n573_ );
not g373 ( new_n575_, keyIn_0_76 );
nand g374 ( new_n576_, new_n346_, new_n558_, new_n573_ );
nand g375 ( new_n577_, new_n576_, new_n575_ );
nand g376 ( new_n578_, new_n577_, new_n574_ );
nand g377 ( new_n579_, new_n578_, new_n238_ );
nand g378 ( new_n580_, new_n579_, keyIn_0_82 );
not g379 ( new_n581_, keyIn_0_82 );
nand g380 ( new_n582_, new_n578_, new_n581_, new_n238_ );
nand g381 ( new_n583_, new_n580_, new_n582_ );
nand g382 ( new_n584_, new_n583_, N17 );
nand g383 ( new_n585_, new_n580_, new_n374_, new_n582_ );
nand g384 ( new_n586_, new_n584_, new_n570_, new_n585_ );
nand g385 ( new_n587_, new_n584_, new_n585_ );
nand g386 ( new_n588_, new_n587_, keyIn_0_105 );
nand g387 ( N728, new_n588_, new_n586_ );
nand g388 ( new_n590_, new_n578_, new_n562_ );
nand g389 ( new_n591_, new_n590_, keyIn_0_83 );
not g390 ( new_n592_, keyIn_0_83 );
nand g391 ( new_n593_, new_n578_, new_n592_, new_n562_ );
nand g392 ( new_n594_, new_n591_, new_n593_ );
nand g393 ( new_n595_, new_n594_, N21 );
nand g394 ( new_n596_, new_n591_, new_n372_, new_n593_ );
nand g395 ( new_n597_, new_n595_, keyIn_0_106, new_n596_ );
not g396 ( new_n598_, keyIn_0_106 );
nand g397 ( new_n599_, new_n595_, new_n596_ );
nand g398 ( new_n600_, new_n599_, new_n598_ );
nand g399 ( N729, new_n600_, new_n597_ );
nand g400 ( new_n602_, new_n578_, new_n336_ );
xnor g401 ( N730, new_n602_, N25 );
not g402 ( new_n604_, keyIn_0_84 );
nand g403 ( new_n605_, new_n578_, new_n567_ );
nand g404 ( new_n606_, new_n605_, new_n604_ );
nand g405 ( new_n607_, new_n578_, keyIn_0_84, new_n567_ );
nand g406 ( new_n608_, new_n606_, new_n607_ );
nand g407 ( new_n609_, new_n608_, N29 );
not g408 ( new_n610_, N29 );
nand g409 ( new_n611_, new_n606_, new_n610_, new_n607_ );
nand g410 ( new_n612_, new_n609_, keyIn_0_107, new_n611_ );
not g411 ( new_n613_, keyIn_0_107 );
nand g412 ( new_n614_, new_n609_, new_n611_ );
nand g413 ( new_n615_, new_n614_, new_n613_ );
nand g414 ( N731, new_n615_, new_n612_ );
not g415 ( new_n617_, keyIn_0_108 );
nand g416 ( new_n618_, new_n528_, new_n556_, new_n525_, new_n553_ );
not g417 ( new_n619_, new_n618_ );
nand g418 ( new_n620_, new_n346_, keyIn_0_77, new_n498_, new_n619_ );
not g419 ( new_n621_, keyIn_0_77 );
nand g420 ( new_n622_, new_n346_, new_n498_, new_n619_ );
nand g421 ( new_n623_, new_n622_, new_n621_ );
nand g422 ( new_n624_, new_n623_, new_n620_ );
nand g423 ( new_n625_, new_n624_, new_n238_ );
nand g424 ( new_n626_, new_n625_, keyIn_0_85 );
not g425 ( new_n627_, keyIn_0_85 );
nand g426 ( new_n628_, new_n624_, new_n627_, new_n238_ );
nand g427 ( new_n629_, new_n626_, new_n628_ );
nand g428 ( new_n630_, new_n629_, N33 );
nand g429 ( new_n631_, new_n626_, new_n423_, new_n628_ );
nand g430 ( new_n632_, new_n630_, new_n617_, new_n631_ );
nand g431 ( new_n633_, new_n630_, new_n631_ );
nand g432 ( new_n634_, new_n633_, keyIn_0_108 );
nand g433 ( N732, new_n634_, new_n632_ );
not g434 ( new_n636_, keyIn_0_86 );
nand g435 ( new_n637_, new_n624_, new_n562_ );
nand g436 ( new_n638_, new_n637_, new_n636_ );
nand g437 ( new_n639_, new_n624_, keyIn_0_86, new_n562_ );
nand g438 ( new_n640_, new_n638_, new_n639_ );
nand g439 ( new_n641_, new_n640_, N37 );
nand g440 ( new_n642_, new_n638_, new_n424_, new_n639_ );
nand g441 ( new_n643_, new_n641_, keyIn_0_109, new_n642_ );
not g442 ( new_n644_, keyIn_0_109 );
nand g443 ( new_n645_, new_n641_, new_n642_ );
nand g444 ( new_n646_, new_n645_, new_n644_ );
nand g445 ( N733, new_n646_, new_n643_ );
not g446 ( new_n648_, keyIn_0_110 );
nand g447 ( new_n649_, new_n624_, new_n336_ );
nand g448 ( new_n650_, new_n649_, keyIn_0_87 );
not g449 ( new_n651_, keyIn_0_87 );
nand g450 ( new_n652_, new_n624_, new_n651_, new_n336_ );
nand g451 ( new_n653_, new_n650_, new_n652_ );
nand g452 ( new_n654_, new_n653_, N41 );
nand g453 ( new_n655_, new_n650_, new_n433_, new_n652_ );
nand g454 ( new_n656_, new_n654_, new_n648_, new_n655_ );
nand g455 ( new_n657_, new_n654_, new_n655_ );
nand g456 ( new_n658_, new_n657_, keyIn_0_110 );
nand g457 ( N734, new_n658_, new_n656_ );
not g458 ( new_n660_, keyIn_0_111 );
nand g459 ( new_n661_, new_n624_, new_n567_ );
nand g460 ( new_n662_, new_n661_, keyIn_0_88 );
not g461 ( new_n663_, keyIn_0_88 );
nand g462 ( new_n664_, new_n624_, new_n663_, new_n567_ );
nand g463 ( new_n665_, new_n662_, new_n664_ );
nand g464 ( new_n666_, new_n665_, N45 );
nand g465 ( new_n667_, new_n662_, new_n434_, new_n664_ );
nand g466 ( new_n668_, new_n666_, new_n660_, new_n667_ );
nand g467 ( new_n669_, new_n666_, new_n667_ );
nand g468 ( new_n670_, new_n669_, keyIn_0_111 );
nand g469 ( N735, new_n670_, new_n668_ );
and g470 ( new_n672_, new_n346_, new_n573_, new_n619_ );
nand g471 ( new_n673_, new_n672_, new_n238_ );
xnor g472 ( N736, new_n673_, N49 );
nand g473 ( new_n675_, new_n672_, new_n562_ );
xnor g474 ( N737, new_n675_, N53 );
nand g475 ( new_n677_, new_n672_, new_n336_ );
xnor g476 ( N738, new_n677_, N57 );
nand g477 ( new_n679_, new_n672_, new_n567_ );
xnor g478 ( N739, new_n679_, N61 );
not g479 ( new_n681_, keyIn_0_112 );
not g480 ( new_n682_, keyIn_0_89 );
not g481 ( new_n683_, keyIn_0_75 );
not g482 ( new_n684_, keyIn_0_74 );
not g483 ( new_n685_, keyIn_0_66 );
nand g484 ( new_n686_, new_n495_, new_n685_, new_n496_ );
nand g485 ( new_n687_, new_n497_, keyIn_0_66 );
nand g486 ( new_n688_, new_n687_, new_n686_ );
and g487 ( new_n689_, new_n571_, new_n529_, new_n557_ );
nand g488 ( new_n690_, new_n688_, new_n689_, new_n684_ );
nand g489 ( new_n691_, new_n688_, new_n689_ );
nand g490 ( new_n692_, new_n691_, keyIn_0_74 );
nand g491 ( new_n693_, new_n692_, new_n690_ );
and g492 ( new_n694_, new_n528_, new_n525_ );
nor g493 ( new_n695_, new_n694_, new_n557_ );
nand g494 ( new_n696_, new_n498_, new_n695_ );
nand g495 ( new_n697_, new_n696_, keyIn_0_72 );
not g496 ( new_n698_, keyIn_0_72 );
nand g497 ( new_n699_, new_n498_, new_n695_, new_n698_ );
nand g498 ( new_n700_, new_n697_, new_n699_ );
and g499 ( new_n701_, new_n693_, new_n700_ );
nand g500 ( new_n702_, new_n497_, keyIn_0_65 );
not g501 ( new_n703_, keyIn_0_65 );
nand g502 ( new_n704_, new_n495_, new_n703_, new_n496_ );
nand g503 ( new_n705_, new_n702_, new_n704_ );
nor g504 ( new_n706_, new_n618_, new_n420_ );
nand g505 ( new_n707_, new_n706_, new_n705_, keyIn_0_73 );
not g506 ( new_n708_, keyIn_0_73 );
nand g507 ( new_n709_, new_n706_, new_n705_ );
nand g508 ( new_n710_, new_n709_, new_n708_ );
nand g509 ( new_n711_, new_n710_, new_n707_ );
not g510 ( new_n712_, keyIn_0_71 );
nor g511 ( new_n713_, new_n694_, new_n571_, new_n557_ );
nand g512 ( new_n714_, new_n495_, keyIn_0_64, new_n496_ );
not g513 ( new_n715_, keyIn_0_64 );
nand g514 ( new_n716_, new_n497_, new_n715_ );
nand g515 ( new_n717_, new_n713_, new_n712_, new_n714_, new_n716_ );
nand g516 ( new_n718_, new_n695_, new_n420_, new_n714_, new_n716_ );
nand g517 ( new_n719_, new_n718_, keyIn_0_71 );
nand g518 ( new_n720_, new_n719_, new_n717_ );
and g519 ( new_n721_, new_n720_, new_n711_ );
nand g520 ( new_n722_, new_n721_, new_n701_, new_n683_ );
nand g521 ( new_n723_, new_n720_, new_n711_, new_n693_, new_n700_ );
nand g522 ( new_n724_, new_n723_, keyIn_0_75 );
xnor g523 ( new_n725_, new_n276_, keyIn_0_67 );
and g524 ( new_n726_, new_n238_, new_n725_, new_n304_, new_n336_ );
nand g525 ( new_n727_, new_n722_, new_n724_, new_n726_ );
nand g526 ( new_n728_, new_n727_, keyIn_0_78 );
not g527 ( new_n729_, keyIn_0_78 );
nand g528 ( new_n730_, new_n722_, new_n724_, new_n729_, new_n726_ );
nand g529 ( new_n731_, new_n728_, new_n682_, new_n557_, new_n730_ );
nand g530 ( new_n732_, new_n728_, new_n557_, new_n730_ );
nand g531 ( new_n733_, new_n732_, keyIn_0_89 );
nand g532 ( new_n734_, new_n733_, new_n731_ );
nand g533 ( new_n735_, new_n734_, N65 );
not g534 ( new_n736_, N65 );
nand g535 ( new_n737_, new_n733_, new_n736_, new_n731_ );
nand g536 ( new_n738_, new_n735_, new_n681_, new_n737_ );
nand g537 ( new_n739_, new_n735_, new_n737_ );
nand g538 ( new_n740_, new_n739_, keyIn_0_112 );
nand g539 ( N740, new_n740_, new_n738_ );
nand g540 ( new_n742_, new_n728_, keyIn_0_90, new_n694_, new_n730_ );
not g541 ( new_n743_, keyIn_0_90 );
nand g542 ( new_n744_, new_n728_, new_n694_, new_n730_ );
nand g543 ( new_n745_, new_n744_, new_n743_ );
nand g544 ( new_n746_, new_n745_, new_n742_ );
nand g545 ( new_n747_, new_n746_, N69 );
not g546 ( new_n748_, N69 );
nand g547 ( new_n749_, new_n745_, new_n748_, new_n742_ );
nand g548 ( new_n750_, new_n747_, keyIn_0_113, new_n749_ );
not g549 ( new_n751_, keyIn_0_113 );
nand g550 ( new_n752_, new_n747_, new_n749_ );
nand g551 ( new_n753_, new_n752_, new_n751_ );
nand g552 ( N741, new_n753_, new_n750_ );
nand g553 ( new_n755_, new_n728_, keyIn_0_91, new_n572_, new_n730_ );
not g554 ( new_n756_, keyIn_0_91 );
nand g555 ( new_n757_, new_n728_, new_n572_, new_n730_ );
nand g556 ( new_n758_, new_n757_, new_n756_ );
nand g557 ( new_n759_, new_n758_, new_n755_ );
nand g558 ( new_n760_, new_n759_, N73 );
not g559 ( new_n761_, N73 );
nand g560 ( new_n762_, new_n758_, new_n761_, new_n755_ );
nand g561 ( new_n763_, new_n760_, keyIn_0_114, new_n762_ );
not g562 ( new_n764_, keyIn_0_114 );
nand g563 ( new_n765_, new_n760_, new_n762_ );
nand g564 ( new_n766_, new_n765_, new_n764_ );
nand g565 ( N742, new_n766_, new_n763_ );
not g566 ( new_n768_, keyIn_0_115 );
nand g567 ( new_n769_, new_n728_, keyIn_0_92, new_n420_, new_n730_ );
not g568 ( new_n770_, keyIn_0_92 );
nand g569 ( new_n771_, new_n728_, new_n420_, new_n730_ );
nand g570 ( new_n772_, new_n771_, new_n770_ );
nand g571 ( new_n773_, new_n772_, new_n769_ );
nand g572 ( new_n774_, new_n773_, N77 );
not g573 ( new_n775_, N77 );
nand g574 ( new_n776_, new_n772_, new_n775_, new_n769_ );
nand g575 ( new_n777_, new_n774_, new_n768_, new_n776_ );
nand g576 ( new_n778_, new_n774_, new_n776_ );
nand g577 ( new_n779_, new_n778_, keyIn_0_115 );
nand g578 ( N743, new_n779_, new_n777_ );
xnor g579 ( new_n781_, new_n333_, keyIn_0_68 );
nor g580 ( new_n782_, new_n781_, new_n237_, new_n562_, new_n304_ );
nand g581 ( new_n783_, new_n722_, new_n724_, new_n782_, keyIn_0_79 );
not g582 ( new_n784_, keyIn_0_79 );
nand g583 ( new_n785_, new_n722_, new_n724_, new_n782_ );
nand g584 ( new_n786_, new_n785_, new_n784_ );
nand g585 ( new_n787_, new_n786_, keyIn_0_93, new_n557_, new_n783_ );
not g586 ( new_n788_, keyIn_0_93 );
nand g587 ( new_n789_, new_n786_, new_n557_, new_n783_ );
nand g588 ( new_n790_, new_n789_, new_n788_ );
nand g589 ( new_n791_, new_n790_, new_n787_ );
nand g590 ( new_n792_, new_n791_, N81 );
not g591 ( new_n793_, N81 );
nand g592 ( new_n794_, new_n790_, new_n793_, new_n787_ );
nand g593 ( new_n795_, new_n792_, keyIn_0_116, new_n794_ );
not g594 ( new_n796_, keyIn_0_116 );
nand g595 ( new_n797_, new_n792_, new_n794_ );
nand g596 ( new_n798_, new_n797_, new_n796_ );
nand g597 ( N744, new_n798_, new_n795_ );
not g598 ( new_n800_, keyIn_0_117 );
nand g599 ( new_n801_, new_n786_, keyIn_0_94, new_n694_, new_n783_ );
not g600 ( new_n802_, keyIn_0_94 );
nand g601 ( new_n803_, new_n786_, new_n694_, new_n783_ );
nand g602 ( new_n804_, new_n803_, new_n802_ );
nand g603 ( new_n805_, new_n804_, new_n801_ );
nand g604 ( new_n806_, new_n805_, N85 );
not g605 ( new_n807_, N85 );
nand g606 ( new_n808_, new_n804_, new_n807_, new_n801_ );
nand g607 ( new_n809_, new_n806_, new_n800_, new_n808_ );
nand g608 ( new_n810_, new_n806_, new_n808_ );
nand g609 ( new_n811_, new_n810_, keyIn_0_117 );
nand g610 ( N745, new_n811_, new_n809_ );
nand g611 ( new_n813_, new_n786_, keyIn_0_95, new_n572_, new_n783_ );
not g612 ( new_n814_, keyIn_0_95 );
nand g613 ( new_n815_, new_n786_, new_n572_, new_n783_ );
nand g614 ( new_n816_, new_n815_, new_n814_ );
nand g615 ( new_n817_, new_n816_, new_n813_ );
nand g616 ( new_n818_, new_n817_, N89 );
not g617 ( new_n819_, N89 );
nand g618 ( new_n820_, new_n816_, new_n819_, new_n813_ );
nand g619 ( new_n821_, new_n818_, keyIn_0_118, new_n820_ );
not g620 ( new_n822_, keyIn_0_118 );
nand g621 ( new_n823_, new_n818_, new_n820_ );
nand g622 ( new_n824_, new_n823_, new_n822_ );
nand g623 ( N746, new_n824_, new_n821_ );
nand g624 ( new_n826_, new_n786_, keyIn_0_96, new_n420_, new_n783_ );
not g625 ( new_n827_, keyIn_0_96 );
nand g626 ( new_n828_, new_n786_, new_n420_, new_n783_ );
nand g627 ( new_n829_, new_n828_, new_n827_ );
nand g628 ( new_n830_, new_n829_, new_n826_ );
nand g629 ( new_n831_, new_n830_, N93 );
not g630 ( new_n832_, N93 );
nand g631 ( new_n833_, new_n829_, new_n832_, new_n826_ );
nand g632 ( new_n834_, new_n831_, keyIn_0_119, new_n833_ );
not g633 ( new_n835_, keyIn_0_119 );
nand g634 ( new_n836_, new_n831_, new_n833_ );
nand g635 ( new_n837_, new_n836_, new_n835_ );
nand g636 ( N747, new_n837_, new_n834_ );
not g637 ( new_n839_, keyIn_0_97 );
not g638 ( new_n840_, keyIn_0_80 );
nor g639 ( new_n841_, new_n238_, new_n567_, new_n333_, new_n276_ );
nand g640 ( new_n842_, new_n722_, new_n724_, new_n840_, new_n841_ );
nand g641 ( new_n843_, new_n722_, new_n724_, new_n841_ );
nand g642 ( new_n844_, new_n843_, keyIn_0_80 );
nand g643 ( new_n845_, new_n844_, new_n839_, new_n557_, new_n842_ );
nand g644 ( new_n846_, new_n844_, new_n557_, new_n842_ );
nand g645 ( new_n847_, new_n846_, keyIn_0_97 );
nand g646 ( new_n848_, new_n847_, new_n845_ );
nand g647 ( new_n849_, new_n848_, N97 );
not g648 ( new_n850_, N97 );
nand g649 ( new_n851_, new_n847_, new_n850_, new_n845_ );
nand g650 ( new_n852_, new_n849_, keyIn_0_120, new_n851_ );
not g651 ( new_n853_, keyIn_0_120 );
nand g652 ( new_n854_, new_n849_, new_n851_ );
nand g653 ( new_n855_, new_n854_, new_n853_ );
nand g654 ( N748, new_n855_, new_n852_ );
not g655 ( new_n857_, keyIn_0_121 );
nand g656 ( new_n858_, new_n844_, keyIn_0_98, new_n694_, new_n842_ );
not g657 ( new_n859_, keyIn_0_98 );
nand g658 ( new_n860_, new_n844_, new_n694_, new_n842_ );
nand g659 ( new_n861_, new_n860_, new_n859_ );
nand g660 ( new_n862_, new_n861_, new_n858_ );
nand g661 ( new_n863_, new_n862_, N101 );
not g662 ( new_n864_, N101 );
nand g663 ( new_n865_, new_n861_, new_n864_, new_n858_ );
nand g664 ( new_n866_, new_n863_, new_n857_, new_n865_ );
nand g665 ( new_n867_, new_n863_, new_n865_ );
nand g666 ( new_n868_, new_n867_, keyIn_0_121 );
nand g667 ( N749, new_n868_, new_n866_ );
not g668 ( new_n870_, keyIn_0_122 );
not g669 ( new_n871_, keyIn_0_99 );
nand g670 ( new_n872_, new_n844_, new_n871_, new_n572_, new_n842_ );
nand g671 ( new_n873_, new_n844_, new_n572_, new_n842_ );
nand g672 ( new_n874_, new_n873_, keyIn_0_99 );
nand g673 ( new_n875_, new_n874_, new_n872_ );
nand g674 ( new_n876_, new_n875_, N105 );
not g675 ( new_n877_, N105 );
nand g676 ( new_n878_, new_n874_, new_n877_, new_n872_ );
nand g677 ( new_n879_, new_n876_, new_n870_, new_n878_ );
nand g678 ( new_n880_, new_n876_, new_n878_ );
nand g679 ( new_n881_, new_n880_, keyIn_0_122 );
nand g680 ( N750, new_n881_, new_n879_ );
not g681 ( new_n883_, keyIn_0_100 );
nand g682 ( new_n884_, new_n844_, new_n883_, new_n420_, new_n842_ );
nand g683 ( new_n885_, new_n844_, new_n420_, new_n842_ );
nand g684 ( new_n886_, new_n885_, keyIn_0_100 );
nand g685 ( new_n887_, new_n886_, new_n884_ );
nand g686 ( new_n888_, new_n887_, N109 );
not g687 ( new_n889_, N109 );
nand g688 ( new_n890_, new_n886_, new_n889_, new_n884_ );
nand g689 ( new_n891_, new_n888_, keyIn_0_123, new_n890_ );
not g690 ( new_n892_, keyIn_0_123 );
nand g691 ( new_n893_, new_n888_, new_n890_ );
nand g692 ( new_n894_, new_n893_, new_n892_ );
nand g693 ( N751, new_n894_, new_n891_ );
not g694 ( new_n896_, keyIn_0_124 );
not g695 ( new_n897_, keyIn_0_81 );
not g696 ( new_n898_, keyIn_0_69 );
nor g697 ( new_n899_, new_n237_, new_n898_ );
nor g698 ( new_n900_, new_n333_, keyIn_0_70 );
nand g699 ( new_n901_, new_n333_, keyIn_0_70 );
nand g700 ( new_n902_, new_n237_, new_n898_ );
nand g701 ( new_n903_, new_n902_, new_n901_ );
nor g702 ( new_n904_, new_n903_, new_n899_, new_n338_, new_n900_ );
nand g703 ( new_n905_, new_n722_, new_n724_, new_n897_, new_n904_ );
nand g704 ( new_n906_, new_n722_, new_n724_, new_n904_ );
nand g705 ( new_n907_, new_n906_, keyIn_0_81 );
nand g706 ( new_n908_, new_n907_, keyIn_0_101, new_n557_, new_n905_ );
not g707 ( new_n909_, keyIn_0_101 );
nand g708 ( new_n910_, new_n907_, new_n557_, new_n905_ );
nand g709 ( new_n911_, new_n910_, new_n909_ );
nand g710 ( new_n912_, new_n911_, new_n908_ );
nand g711 ( new_n913_, new_n912_, N113 );
not g712 ( new_n914_, N113 );
nand g713 ( new_n915_, new_n911_, new_n914_, new_n908_ );
nand g714 ( new_n916_, new_n913_, new_n896_, new_n915_ );
nand g715 ( new_n917_, new_n913_, new_n915_ );
nand g716 ( new_n918_, new_n917_, keyIn_0_124 );
nand g717 ( N752, new_n918_, new_n916_ );
nand g718 ( new_n920_, new_n907_, keyIn_0_102, new_n694_, new_n905_ );
not g719 ( new_n921_, keyIn_0_102 );
nand g720 ( new_n922_, new_n907_, new_n694_, new_n905_ );
nand g721 ( new_n923_, new_n922_, new_n921_ );
nand g722 ( new_n924_, new_n923_, new_n920_ );
nand g723 ( new_n925_, new_n924_, N117 );
not g724 ( new_n926_, N117 );
nand g725 ( new_n927_, new_n923_, new_n926_, new_n920_ );
nand g726 ( new_n928_, new_n925_, keyIn_0_125, new_n927_ );
not g727 ( new_n929_, keyIn_0_125 );
nand g728 ( new_n930_, new_n925_, new_n927_ );
nand g729 ( new_n931_, new_n930_, new_n929_ );
nand g730 ( N753, new_n931_, new_n928_ );
not g731 ( new_n933_, keyIn_0_126 );
not g732 ( new_n934_, keyIn_0_103 );
nand g733 ( new_n935_, new_n907_, new_n934_, new_n572_, new_n905_ );
nand g734 ( new_n936_, new_n907_, new_n572_, new_n905_ );
nand g735 ( new_n937_, new_n936_, keyIn_0_103 );
nand g736 ( new_n938_, new_n937_, new_n935_ );
nand g737 ( new_n939_, new_n938_, N121 );
not g738 ( new_n940_, N121 );
nand g739 ( new_n941_, new_n937_, new_n940_, new_n935_ );
nand g740 ( new_n942_, new_n939_, new_n933_, new_n941_ );
nand g741 ( new_n943_, new_n939_, new_n941_ );
nand g742 ( new_n944_, new_n943_, keyIn_0_126 );
nand g743 ( N754, new_n944_, new_n942_ );
nand g744 ( new_n946_, new_n907_, keyIn_0_104, new_n420_, new_n905_ );
not g745 ( new_n947_, keyIn_0_104 );
nand g746 ( new_n948_, new_n907_, new_n420_, new_n905_ );
nand g747 ( new_n949_, new_n948_, new_n947_ );
nand g748 ( new_n950_, new_n949_, new_n946_ );
nand g749 ( new_n951_, new_n950_, N125 );
not g750 ( new_n952_, N125 );
nand g751 ( new_n953_, new_n949_, new_n952_, new_n946_ );
nand g752 ( new_n954_, new_n951_, keyIn_0_127, new_n953_ );
not g753 ( new_n955_, keyIn_0_127 );
nand g754 ( new_n956_, new_n951_, new_n953_ );
nand g755 ( new_n957_, new_n956_, new_n955_ );
nand g756 ( N755, new_n957_, new_n954_ );
endmodule