module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n1233_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1517_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n706_, new_n649_, new_n1119_, new_n1213_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1447_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n1377_, new_n1522_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n1512_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1198_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n473_, new_n1147_, new_n1373_, new_n1422_, new_n1523_, new_n1468_, new_n969_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n621_, new_n1423_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1507_, new_n1439_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n762_, new_n1349_, new_n1193_, new_n1437_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1171_, new_n867_, new_n1032_, new_n901_, new_n276_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n1109_, new_n261_, new_n672_, new_n1496_, new_n1269_, new_n616_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1461_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n861_, new_n1252_, new_n352_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n1064_, new_n1065_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1325_, new_n993_, new_n1191_, new_n824_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n302_, new_n755_, new_n1040_, new_n1509_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1185_, new_n1240_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1334_, new_n531_, new_n593_, new_n974_, new_n252_, new_n1248_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1492_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n1421_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1534_, new_n684_, new_n640_, new_n1274_, new_n754_, new_n653_, new_n905_, new_n377_, new_n1258_, new_n1539_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n984_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n1340_, new_n798_, new_n1180_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n601_, new_n842_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n1264_, new_n215_, new_n1319_, new_n626_, new_n1473_, new_n990_, new_n716_, new_n701_, new_n1238_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n1203_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n906_, new_n361_, new_n764_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n216_, new_n1348_, new_n917_, new_n1322_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1202_, new_n436_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1329_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n1536_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n400_, new_n1175_, new_n1136_, new_n693_, new_n1287_, new_n1485_, new_n505_, new_n1462_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n520_, new_n1347_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1470_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1529_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n756_, new_n823_, new_n574_, new_n1500_, new_n928_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n1399_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1243_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n1449_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n1498_, new_n204_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_55 );
not g0001 ( new_n203_, keyIn_0_32 );
nand g0002 ( new_n204_, N65, N69 );
not g0003 ( new_n205_, new_n204_ );
nor g0004 ( new_n206_, N65, N69 );
nor g0005 ( new_n207_, new_n205_, new_n206_ );
nor g0006 ( new_n208_, new_n207_, keyIn_0_8 );
nand g0007 ( new_n209_, new_n207_, keyIn_0_8 );
not g0008 ( new_n210_, new_n209_ );
nor g0009 ( new_n211_, new_n210_, new_n208_ );
not g0010 ( new_n212_, new_n211_ );
not g0011 ( new_n213_, keyIn_0_9 );
nand g0012 ( new_n214_, N73, N77 );
not g0013 ( new_n215_, new_n214_ );
nor g0014 ( new_n216_, N73, N77 );
nor g0015 ( new_n217_, new_n215_, new_n216_ );
nor g0016 ( new_n218_, new_n217_, new_n213_ );
nand g0017 ( new_n219_, new_n217_, new_n213_ );
not g0018 ( new_n220_, new_n219_ );
nor g0019 ( new_n221_, new_n220_, new_n218_ );
not g0020 ( new_n222_, new_n221_ );
nand g0021 ( new_n223_, new_n212_, new_n222_ );
nor g0022 ( new_n224_, new_n212_, new_n222_ );
not g0023 ( new_n225_, new_n224_ );
nand g0024 ( new_n226_, new_n225_, new_n223_ );
nand g0025 ( new_n227_, new_n226_, new_n203_ );
not g0026 ( new_n228_, new_n227_ );
nor g0027 ( new_n229_, new_n226_, new_n203_ );
nor g0028 ( new_n230_, new_n228_, new_n229_ );
not g0029 ( new_n231_, new_n230_ );
not g0030 ( new_n232_, keyIn_0_33 );
not g0031 ( new_n233_, N81 );
nor g0032 ( new_n234_, new_n233_, N85 );
not g0033 ( new_n235_, N85 );
nor g0034 ( new_n236_, new_n235_, N81 );
nor g0035 ( new_n237_, new_n234_, new_n236_ );
not g0036 ( new_n238_, new_n237_ );
nand g0037 ( new_n239_, new_n238_, keyIn_0_10 );
not g0038 ( new_n240_, new_n239_ );
nor g0039 ( new_n241_, new_n238_, keyIn_0_10 );
nor g0040 ( new_n242_, new_n240_, new_n241_ );
not g0041 ( new_n243_, keyIn_0_11 );
nand g0042 ( new_n244_, N89, N93 );
not g0043 ( new_n245_, new_n244_ );
nor g0044 ( new_n246_, N89, N93 );
nor g0045 ( new_n247_, new_n245_, new_n246_ );
nor g0046 ( new_n248_, new_n247_, new_n243_ );
nand g0047 ( new_n249_, new_n247_, new_n243_ );
not g0048 ( new_n250_, new_n249_ );
nor g0049 ( new_n251_, new_n250_, new_n248_ );
nor g0050 ( new_n252_, new_n242_, new_n251_ );
nand g0051 ( new_n253_, new_n242_, new_n251_ );
not g0052 ( new_n254_, new_n253_ );
nor g0053 ( new_n255_, new_n254_, new_n252_ );
nor g0054 ( new_n256_, new_n255_, new_n232_ );
not g0055 ( new_n257_, new_n256_ );
nand g0056 ( new_n258_, new_n255_, new_n232_ );
nand g0057 ( new_n259_, new_n257_, new_n258_ );
nand g0058 ( new_n260_, new_n231_, new_n259_ );
not g0059 ( new_n261_, new_n260_ );
nor g0060 ( new_n262_, new_n231_, new_n259_ );
nor g0061 ( new_n263_, new_n261_, new_n262_ );
not g0062 ( new_n264_, new_n263_ );
nand g0063 ( new_n265_, new_n264_, keyIn_0_43 );
not g0064 ( new_n266_, keyIn_0_43 );
nand g0065 ( new_n267_, new_n263_, new_n266_ );
nand g0066 ( new_n268_, new_n265_, new_n267_ );
nand g0067 ( new_n269_, N129, N137 );
nand g0068 ( new_n270_, new_n268_, new_n269_ );
not g0069 ( new_n271_, new_n270_ );
nor g0070 ( new_n272_, new_n268_, new_n269_ );
nor g0071 ( new_n273_, new_n271_, new_n272_ );
not g0072 ( new_n274_, new_n273_ );
nand g0073 ( new_n275_, new_n274_, keyIn_0_47 );
not g0074 ( new_n276_, keyIn_0_47 );
nand g0075 ( new_n277_, new_n273_, new_n276_ );
nand g0076 ( new_n278_, new_n275_, new_n277_ );
not g0077 ( new_n279_, N1 );
nor g0078 ( new_n280_, new_n279_, N17 );
not g0079 ( new_n281_, N17 );
nor g0080 ( new_n282_, new_n281_, N1 );
nor g0081 ( new_n283_, new_n280_, new_n282_ );
nand g0082 ( new_n284_, N33, N49 );
not g0083 ( new_n285_, new_n284_ );
nor g0084 ( new_n286_, N33, N49 );
nor g0085 ( new_n287_, new_n285_, new_n286_ );
nor g0086 ( new_n288_, new_n283_, new_n287_ );
nand g0087 ( new_n289_, new_n283_, new_n287_ );
not g0088 ( new_n290_, new_n289_ );
nor g0089 ( new_n291_, new_n290_, new_n288_ );
not g0090 ( new_n292_, new_n291_ );
nand g0091 ( new_n293_, new_n278_, new_n292_ );
nor g0092 ( new_n294_, new_n278_, new_n292_ );
not g0093 ( new_n295_, new_n294_ );
nand g0094 ( new_n296_, new_n295_, new_n293_ );
nand g0095 ( new_n297_, new_n296_, new_n202_ );
not g0096 ( new_n298_, new_n293_ );
nor g0097 ( new_n299_, new_n298_, new_n294_ );
nand g0098 ( new_n300_, new_n299_, keyIn_0_55 );
nand g0099 ( new_n301_, new_n300_, new_n297_ );
not g0100 ( new_n302_, new_n301_ );
not g0101 ( new_n303_, keyIn_0_35 );
not g0102 ( new_n304_, keyIn_0_14 );
nand g0103 ( new_n305_, N113, N117 );
not g0104 ( new_n306_, new_n305_ );
nor g0105 ( new_n307_, N113, N117 );
nor g0106 ( new_n308_, new_n306_, new_n307_ );
nor g0107 ( new_n309_, new_n308_, new_n304_ );
nand g0108 ( new_n310_, new_n308_, new_n304_ );
not g0109 ( new_n311_, new_n310_ );
nor g0110 ( new_n312_, new_n311_, new_n309_ );
not g0111 ( new_n313_, new_n312_ );
not g0112 ( new_n314_, keyIn_0_15 );
nand g0113 ( new_n315_, N121, N125 );
not g0114 ( new_n316_, new_n315_ );
nor g0115 ( new_n317_, N121, N125 );
nor g0116 ( new_n318_, new_n316_, new_n317_ );
nor g0117 ( new_n319_, new_n318_, new_n314_ );
nand g0118 ( new_n320_, new_n318_, new_n314_ );
not g0119 ( new_n321_, new_n320_ );
nor g0120 ( new_n322_, new_n321_, new_n319_ );
not g0121 ( new_n323_, new_n322_ );
nand g0122 ( new_n324_, new_n313_, new_n323_ );
nor g0123 ( new_n325_, new_n313_, new_n323_ );
not g0124 ( new_n326_, new_n325_ );
nand g0125 ( new_n327_, new_n326_, new_n324_ );
nand g0126 ( new_n328_, new_n327_, new_n303_ );
not g0127 ( new_n329_, new_n328_ );
nor g0128 ( new_n330_, new_n327_, new_n303_ );
nor g0129 ( new_n331_, new_n329_, new_n330_ );
not g0130 ( new_n332_, new_n331_ );
nand g0131 ( new_n333_, new_n332_, new_n259_ );
not g0132 ( new_n334_, new_n333_ );
nor g0133 ( new_n335_, new_n332_, new_n259_ );
nor g0134 ( new_n336_, new_n334_, new_n335_ );
not g0135 ( new_n337_, new_n336_ );
nand g0136 ( new_n338_, new_n337_, keyIn_0_46 );
not g0137 ( new_n339_, keyIn_0_46 );
nand g0138 ( new_n340_, new_n336_, new_n339_ );
nand g0139 ( new_n341_, new_n338_, new_n340_ );
nand g0140 ( new_n342_, N132, N137 );
not g0141 ( new_n343_, new_n342_ );
nand g0142 ( new_n344_, new_n341_, new_n343_ );
not g0143 ( new_n345_, new_n344_ );
nor g0144 ( new_n346_, new_n341_, new_n343_ );
nor g0145 ( new_n347_, new_n345_, new_n346_ );
not g0146 ( new_n348_, new_n347_ );
nand g0147 ( new_n349_, new_n348_, keyIn_0_50 );
not g0148 ( new_n350_, keyIn_0_50 );
nand g0149 ( new_n351_, new_n347_, new_n350_ );
nand g0150 ( new_n352_, new_n349_, new_n351_ );
not g0151 ( new_n353_, keyIn_0_23 );
nand g0152 ( new_n354_, N13, N29 );
not g0153 ( new_n355_, new_n354_ );
nor g0154 ( new_n356_, N13, N29 );
nor g0155 ( new_n357_, new_n355_, new_n356_ );
nor g0156 ( new_n358_, new_n357_, new_n353_ );
nand g0157 ( new_n359_, new_n357_, new_n353_ );
not g0158 ( new_n360_, new_n359_ );
nor g0159 ( new_n361_, new_n360_, new_n358_ );
nand g0160 ( new_n362_, N45, N61 );
not g0161 ( new_n363_, new_n362_ );
nor g0162 ( new_n364_, N45, N61 );
nor g0163 ( new_n365_, new_n363_, new_n364_ );
nor g0164 ( new_n366_, new_n361_, new_n365_ );
nand g0165 ( new_n367_, new_n361_, new_n365_ );
not g0166 ( new_n368_, new_n367_ );
nor g0167 ( new_n369_, new_n368_, new_n366_ );
not g0168 ( new_n370_, new_n369_ );
nand g0169 ( new_n371_, new_n352_, new_n370_ );
nor g0170 ( new_n372_, new_n352_, new_n370_ );
not g0171 ( new_n373_, new_n372_ );
nand g0172 ( new_n374_, new_n373_, new_n371_ );
nand g0173 ( new_n375_, new_n374_, keyIn_0_58 );
not g0174 ( new_n376_, keyIn_0_58 );
not g0175 ( new_n377_, new_n371_ );
nor g0176 ( new_n378_, new_n377_, new_n372_ );
nand g0177 ( new_n379_, new_n378_, new_n376_ );
nand g0178 ( new_n380_, new_n379_, new_n375_ );
not g0179 ( new_n381_, new_n380_ );
not g0180 ( new_n382_, keyIn_0_56 );
nand g0181 ( new_n383_, N97, N101 );
not g0182 ( new_n384_, new_n383_ );
nor g0183 ( new_n385_, N97, N101 );
nor g0184 ( new_n386_, new_n384_, new_n385_ );
nor g0185 ( new_n387_, new_n386_, keyIn_0_12 );
nand g0186 ( new_n388_, new_n386_, keyIn_0_12 );
not g0187 ( new_n389_, new_n388_ );
nor g0188 ( new_n390_, new_n389_, new_n387_ );
not g0189 ( new_n391_, new_n390_ );
not g0190 ( new_n392_, keyIn_0_13 );
nand g0191 ( new_n393_, N105, N109 );
not g0192 ( new_n394_, new_n393_ );
nor g0193 ( new_n395_, N105, N109 );
nor g0194 ( new_n396_, new_n394_, new_n395_ );
nor g0195 ( new_n397_, new_n396_, new_n392_ );
nand g0196 ( new_n398_, new_n396_, new_n392_ );
not g0197 ( new_n399_, new_n398_ );
nor g0198 ( new_n400_, new_n399_, new_n397_ );
not g0199 ( new_n401_, new_n400_ );
nand g0200 ( new_n402_, new_n391_, new_n401_ );
not g0201 ( new_n403_, new_n402_ );
nor g0202 ( new_n404_, new_n391_, new_n401_ );
nor g0203 ( new_n405_, new_n403_, new_n404_ );
not g0204 ( new_n406_, new_n405_ );
nand g0205 ( new_n407_, new_n406_, keyIn_0_34 );
not g0206 ( new_n408_, keyIn_0_34 );
nand g0207 ( new_n409_, new_n405_, new_n408_ );
nand g0208 ( new_n410_, new_n407_, new_n409_ );
nand g0209 ( new_n411_, new_n331_, new_n410_ );
not g0210 ( new_n412_, new_n410_ );
nand g0211 ( new_n413_, new_n332_, new_n412_ );
nand g0212 ( new_n414_, new_n413_, new_n411_ );
nand g0213 ( new_n415_, new_n414_, keyIn_0_44 );
not g0214 ( new_n416_, new_n415_ );
nor g0215 ( new_n417_, new_n414_, keyIn_0_44 );
nor g0216 ( new_n418_, new_n416_, new_n417_ );
nand g0217 ( new_n419_, N130, N137 );
nor g0218 ( new_n420_, new_n418_, new_n419_ );
not g0219 ( new_n421_, new_n420_ );
nand g0220 ( new_n422_, new_n418_, new_n419_ );
nand g0221 ( new_n423_, new_n421_, new_n422_ );
nand g0222 ( new_n424_, new_n423_, keyIn_0_48 );
nor g0223 ( new_n425_, new_n423_, keyIn_0_48 );
not g0224 ( new_n426_, new_n425_ );
nand g0225 ( new_n427_, new_n426_, new_n424_ );
nand g0226 ( new_n428_, N5, N21 );
not g0227 ( new_n429_, new_n428_ );
nor g0228 ( new_n430_, N5, N21 );
nor g0229 ( new_n431_, new_n429_, new_n430_ );
nand g0230 ( new_n432_, N37, N53 );
not g0231 ( new_n433_, new_n432_ );
nor g0232 ( new_n434_, N37, N53 );
nor g0233 ( new_n435_, new_n433_, new_n434_ );
not g0234 ( new_n436_, new_n435_ );
nor g0235 ( new_n437_, new_n436_, new_n431_ );
nand g0236 ( new_n438_, new_n436_, new_n431_ );
not g0237 ( new_n439_, new_n438_ );
nor g0238 ( new_n440_, new_n439_, new_n437_ );
not g0239 ( new_n441_, new_n440_ );
nand g0240 ( new_n442_, new_n427_, new_n441_ );
not g0241 ( new_n443_, new_n424_ );
nor g0242 ( new_n444_, new_n443_, new_n425_ );
nand g0243 ( new_n445_, new_n444_, new_n440_ );
nand g0244 ( new_n446_, new_n445_, new_n442_ );
nand g0245 ( new_n447_, new_n446_, new_n382_ );
nor g0246 ( new_n448_, new_n446_, new_n382_ );
not g0247 ( new_n449_, new_n448_ );
nand g0248 ( new_n450_, new_n449_, new_n447_ );
not g0249 ( new_n451_, keyIn_0_49 );
nand g0250 ( new_n452_, new_n231_, new_n412_ );
nand g0251 ( new_n453_, new_n230_, new_n410_ );
nand g0252 ( new_n454_, new_n452_, new_n453_ );
nand g0253 ( new_n455_, new_n454_, keyIn_0_45 );
not g0254 ( new_n456_, new_n455_ );
nor g0255 ( new_n457_, new_n454_, keyIn_0_45 );
nor g0256 ( new_n458_, new_n456_, new_n457_ );
nand g0257 ( new_n459_, N131, N137 );
nand g0258 ( new_n460_, new_n459_, keyIn_0_16 );
not g0259 ( new_n461_, new_n460_ );
nor g0260 ( new_n462_, new_n459_, keyIn_0_16 );
nor g0261 ( new_n463_, new_n461_, new_n462_ );
nor g0262 ( new_n464_, new_n458_, new_n463_ );
nand g0263 ( new_n465_, new_n458_, new_n463_ );
not g0264 ( new_n466_, new_n465_ );
nor g0265 ( new_n467_, new_n466_, new_n464_ );
nor g0266 ( new_n468_, new_n467_, new_n451_ );
not g0267 ( new_n469_, new_n468_ );
nand g0268 ( new_n470_, new_n467_, new_n451_ );
nand g0269 ( new_n471_, new_n469_, new_n470_ );
not g0270 ( new_n472_, keyIn_0_36 );
not g0271 ( new_n473_, N41 );
nor g0272 ( new_n474_, new_n473_, N57 );
not g0273 ( new_n475_, N57 );
nor g0274 ( new_n476_, new_n475_, N41 );
nor g0275 ( new_n477_, new_n474_, new_n476_ );
not g0276 ( new_n478_, new_n477_ );
nand g0277 ( new_n479_, new_n478_, keyIn_0_22 );
not g0278 ( new_n480_, new_n479_ );
nor g0279 ( new_n481_, new_n478_, keyIn_0_22 );
nor g0280 ( new_n482_, new_n480_, new_n481_ );
not g0281 ( new_n483_, keyIn_0_21 );
nand g0282 ( new_n484_, N9, N25 );
not g0283 ( new_n485_, new_n484_ );
nor g0284 ( new_n486_, N9, N25 );
nor g0285 ( new_n487_, new_n485_, new_n486_ );
nor g0286 ( new_n488_, new_n487_, new_n483_ );
nand g0287 ( new_n489_, new_n487_, new_n483_ );
not g0288 ( new_n490_, new_n489_ );
nor g0289 ( new_n491_, new_n490_, new_n488_ );
nor g0290 ( new_n492_, new_n482_, new_n491_ );
nand g0291 ( new_n493_, new_n482_, new_n491_ );
not g0292 ( new_n494_, new_n493_ );
nor g0293 ( new_n495_, new_n494_, new_n492_ );
nor g0294 ( new_n496_, new_n495_, new_n472_ );
nand g0295 ( new_n497_, new_n495_, new_n472_ );
not g0296 ( new_n498_, new_n497_ );
nor g0297 ( new_n499_, new_n498_, new_n496_ );
not g0298 ( new_n500_, new_n499_ );
nand g0299 ( new_n501_, new_n471_, new_n500_ );
not g0300 ( new_n502_, new_n470_ );
nor g0301 ( new_n503_, new_n502_, new_n468_ );
nand g0302 ( new_n504_, new_n503_, new_n499_ );
nand g0303 ( new_n505_, new_n504_, new_n501_ );
nand g0304 ( new_n506_, new_n505_, keyIn_0_57 );
not g0305 ( new_n507_, new_n506_ );
nor g0306 ( new_n508_, new_n505_, keyIn_0_57 );
nor g0307 ( new_n509_, new_n507_, new_n508_ );
nand g0308 ( new_n510_, new_n509_, new_n450_ );
nor g0309 ( new_n511_, new_n381_, new_n510_ );
not g0310 ( new_n512_, new_n511_ );
not g0311 ( new_n513_, new_n447_ );
nor g0312 ( new_n514_, new_n513_, new_n448_ );
not g0313 ( new_n515_, new_n508_ );
nand g0314 ( new_n516_, new_n515_, new_n506_ );
nor g0315 ( new_n517_, new_n514_, new_n516_ );
nor g0316 ( new_n518_, new_n517_, new_n380_ );
nand g0317 ( new_n519_, new_n514_, new_n516_ );
nand g0318 ( new_n520_, new_n302_, new_n519_ );
nor g0319 ( new_n521_, new_n518_, new_n520_ );
nand g0320 ( new_n522_, new_n521_, new_n512_ );
nand g0321 ( new_n523_, new_n516_, keyIn_0_63 );
nand g0322 ( new_n524_, new_n523_, new_n380_ );
not g0323 ( new_n525_, new_n524_ );
nor g0324 ( new_n526_, new_n516_, keyIn_0_63 );
nand g0325 ( new_n527_, new_n301_, new_n450_ );
nor g0326 ( new_n528_, new_n527_, new_n526_ );
nand g0327 ( new_n529_, new_n528_, new_n525_ );
nand g0328 ( new_n530_, new_n522_, new_n529_ );
not g0329 ( new_n531_, keyIn_0_60 );
not g0330 ( new_n532_, keyIn_0_30 );
not g0331 ( new_n533_, N37 );
nand g0332 ( new_n534_, new_n533_, N33 );
not g0333 ( new_n535_, N33 );
nand g0334 ( new_n536_, new_n535_, N37 );
nand g0335 ( new_n537_, new_n534_, new_n536_ );
nand g0336 ( new_n538_, new_n537_, keyIn_0_4 );
nor g0337 ( new_n539_, new_n537_, keyIn_0_4 );
not g0338 ( new_n540_, new_n539_ );
nand g0339 ( new_n541_, new_n540_, new_n538_ );
not g0340 ( new_n542_, N45 );
nand g0341 ( new_n543_, new_n542_, N41 );
nand g0342 ( new_n544_, new_n473_, N45 );
nand g0343 ( new_n545_, new_n543_, new_n544_ );
nand g0344 ( new_n546_, new_n545_, keyIn_0_5 );
not g0345 ( new_n547_, keyIn_0_5 );
not g0346 ( new_n548_, new_n545_ );
nand g0347 ( new_n549_, new_n548_, new_n547_ );
nand g0348 ( new_n550_, new_n549_, new_n546_ );
nand g0349 ( new_n551_, new_n541_, new_n550_ );
not g0350 ( new_n552_, new_n538_ );
nor g0351 ( new_n553_, new_n552_, new_n539_ );
not g0352 ( new_n554_, new_n546_ );
nor g0353 ( new_n555_, new_n545_, keyIn_0_5 );
nor g0354 ( new_n556_, new_n554_, new_n555_ );
nand g0355 ( new_n557_, new_n553_, new_n556_ );
nand g0356 ( new_n558_, new_n557_, new_n551_ );
nand g0357 ( new_n559_, new_n558_, new_n532_ );
nor g0358 ( new_n560_, new_n553_, new_n556_ );
nor g0359 ( new_n561_, new_n541_, new_n550_ );
nor g0360 ( new_n562_, new_n560_, new_n561_ );
nand g0361 ( new_n563_, new_n562_, keyIn_0_30 );
nand g0362 ( new_n564_, new_n563_, new_n559_ );
not g0363 ( new_n565_, keyIn_0_31 );
not g0364 ( new_n566_, keyIn_0_6 );
not g0365 ( new_n567_, N53 );
nand g0366 ( new_n568_, new_n567_, N49 );
not g0367 ( new_n569_, N49 );
nand g0368 ( new_n570_, new_n569_, N53 );
nand g0369 ( new_n571_, new_n568_, new_n570_ );
nand g0370 ( new_n572_, new_n571_, new_n566_ );
not g0371 ( new_n573_, new_n571_ );
nand g0372 ( new_n574_, new_n573_, keyIn_0_6 );
nand g0373 ( new_n575_, new_n574_, new_n572_ );
not g0374 ( new_n576_, N61 );
nand g0375 ( new_n577_, new_n576_, N57 );
nand g0376 ( new_n578_, new_n475_, N61 );
nand g0377 ( new_n579_, new_n577_, new_n578_ );
nand g0378 ( new_n580_, new_n579_, keyIn_0_7 );
not g0379 ( new_n581_, keyIn_0_7 );
not g0380 ( new_n582_, new_n579_ );
nand g0381 ( new_n583_, new_n582_, new_n581_ );
nand g0382 ( new_n584_, new_n583_, new_n580_ );
nand g0383 ( new_n585_, new_n575_, new_n584_ );
not g0384 ( new_n586_, new_n572_ );
nor g0385 ( new_n587_, new_n571_, new_n566_ );
nor g0386 ( new_n588_, new_n586_, new_n587_ );
not g0387 ( new_n589_, new_n580_ );
nor g0388 ( new_n590_, new_n579_, keyIn_0_7 );
nor g0389 ( new_n591_, new_n589_, new_n590_ );
nand g0390 ( new_n592_, new_n588_, new_n591_ );
nand g0391 ( new_n593_, new_n592_, new_n585_ );
nand g0392 ( new_n594_, new_n593_, new_n565_ );
not g0393 ( new_n595_, new_n593_ );
nand g0394 ( new_n596_, new_n595_, keyIn_0_31 );
nand g0395 ( new_n597_, new_n596_, new_n594_ );
nand g0396 ( new_n598_, new_n597_, new_n564_ );
not g0397 ( new_n599_, new_n559_ );
nor g0398 ( new_n600_, new_n558_, new_n532_ );
nor g0399 ( new_n601_, new_n599_, new_n600_ );
not g0400 ( new_n602_, new_n594_ );
nor g0401 ( new_n603_, new_n593_, new_n565_ );
nor g0402 ( new_n604_, new_n602_, new_n603_ );
nand g0403 ( new_n605_, new_n601_, new_n604_ );
nand g0404 ( new_n606_, new_n605_, new_n598_ );
nand g0405 ( new_n607_, new_n606_, keyIn_0_40 );
not g0406 ( new_n608_, new_n607_ );
nor g0407 ( new_n609_, new_n606_, keyIn_0_40 );
nor g0408 ( new_n610_, new_n608_, new_n609_ );
not g0409 ( new_n611_, keyIn_0_18 );
nand g0410 ( new_n612_, N134, N137 );
nand g0411 ( new_n613_, new_n612_, new_n611_ );
not g0412 ( new_n614_, new_n613_ );
nor g0413 ( new_n615_, new_n612_, new_n611_ );
nor g0414 ( new_n616_, new_n614_, new_n615_ );
nor g0415 ( new_n617_, new_n610_, new_n616_ );
not g0416 ( new_n618_, keyIn_0_40 );
not g0417 ( new_n619_, new_n606_ );
nand g0418 ( new_n620_, new_n619_, new_n618_ );
nand g0419 ( new_n621_, new_n620_, new_n607_ );
not g0420 ( new_n622_, new_n616_ );
nor g0421 ( new_n623_, new_n621_, new_n622_ );
nor g0422 ( new_n624_, new_n617_, new_n623_ );
nor g0423 ( new_n625_, new_n624_, keyIn_0_52 );
not g0424 ( new_n626_, keyIn_0_52 );
nand g0425 ( new_n627_, new_n621_, new_n622_ );
nand g0426 ( new_n628_, new_n610_, new_n616_ );
nand g0427 ( new_n629_, new_n628_, new_n627_ );
nor g0428 ( new_n630_, new_n629_, new_n626_ );
nor g0429 ( new_n631_, new_n625_, new_n630_ );
not g0430 ( new_n632_, keyIn_0_37 );
not g0431 ( new_n633_, N69 );
nor g0432 ( new_n634_, new_n633_, N85 );
nor g0433 ( new_n635_, new_n235_, N69 );
nor g0434 ( new_n636_, new_n634_, new_n635_ );
not g0435 ( new_n637_, new_n636_ );
nand g0436 ( new_n638_, new_n637_, keyIn_0_24 );
not g0437 ( new_n639_, new_n638_ );
nor g0438 ( new_n640_, new_n637_, keyIn_0_24 );
nor g0439 ( new_n641_, new_n639_, new_n640_ );
not g0440 ( new_n642_, N101 );
nor g0441 ( new_n643_, new_n642_, N117 );
not g0442 ( new_n644_, N117 );
nor g0443 ( new_n645_, new_n644_, N101 );
nor g0444 ( new_n646_, new_n643_, new_n645_ );
not g0445 ( new_n647_, new_n646_ );
nand g0446 ( new_n648_, new_n647_, keyIn_0_25 );
not g0447 ( new_n649_, new_n648_ );
nor g0448 ( new_n650_, new_n647_, keyIn_0_25 );
nor g0449 ( new_n651_, new_n649_, new_n650_ );
nor g0450 ( new_n652_, new_n641_, new_n651_ );
nand g0451 ( new_n653_, new_n641_, new_n651_ );
not g0452 ( new_n654_, new_n653_ );
nor g0453 ( new_n655_, new_n654_, new_n652_ );
not g0454 ( new_n656_, new_n655_ );
nand g0455 ( new_n657_, new_n656_, new_n632_ );
not g0456 ( new_n658_, new_n657_ );
nor g0457 ( new_n659_, new_n656_, new_n632_ );
nor g0458 ( new_n660_, new_n658_, new_n659_ );
not g0459 ( new_n661_, new_n660_ );
nor g0460 ( new_n662_, new_n631_, new_n661_ );
nand g0461 ( new_n663_, new_n629_, new_n626_ );
nand g0462 ( new_n664_, new_n624_, keyIn_0_52 );
nand g0463 ( new_n665_, new_n664_, new_n663_ );
nor g0464 ( new_n666_, new_n665_, new_n660_ );
nor g0465 ( new_n667_, new_n662_, new_n666_ );
nor g0466 ( new_n668_, new_n667_, new_n531_ );
nand g0467 ( new_n669_, new_n665_, new_n660_ );
nand g0468 ( new_n670_, new_n631_, new_n661_ );
nand g0469 ( new_n671_, new_n670_, new_n669_ );
nor g0470 ( new_n672_, new_n671_, keyIn_0_60 );
nor g0471 ( new_n673_, new_n668_, new_n672_ );
not g0472 ( new_n674_, keyIn_0_59 );
not g0473 ( new_n675_, keyIn_0_51 );
not g0474 ( new_n676_, keyIn_0_39 );
nand g0475 ( new_n677_, N9, N13 );
not g0476 ( new_n678_, new_n677_ );
nor g0477 ( new_n679_, N9, N13 );
nor g0478 ( new_n680_, new_n678_, new_n679_ );
nand g0479 ( new_n681_, new_n680_, keyIn_0_1 );
not g0480 ( new_n682_, keyIn_0_1 );
not g0481 ( new_n683_, N9 );
not g0482 ( new_n684_, N13 );
nand g0483 ( new_n685_, new_n683_, new_n684_ );
nand g0484 ( new_n686_, new_n685_, new_n677_ );
nand g0485 ( new_n687_, new_n686_, new_n682_ );
nand g0486 ( new_n688_, new_n681_, new_n687_ );
not g0487 ( new_n689_, N5 );
nand g0488 ( new_n690_, new_n689_, N1 );
nand g0489 ( new_n691_, new_n279_, N5 );
nand g0490 ( new_n692_, new_n690_, new_n691_ );
nand g0491 ( new_n693_, new_n692_, keyIn_0_0 );
not g0492 ( new_n694_, new_n693_ );
nor g0493 ( new_n695_, new_n692_, keyIn_0_0 );
nor g0494 ( new_n696_, new_n694_, new_n695_ );
nand g0495 ( new_n697_, new_n696_, new_n688_ );
nor g0496 ( new_n698_, new_n686_, new_n682_ );
nor g0497 ( new_n699_, new_n680_, keyIn_0_1 );
nor g0498 ( new_n700_, new_n699_, new_n698_ );
not g0499 ( new_n701_, keyIn_0_0 );
nor g0500 ( new_n702_, new_n279_, N5 );
nor g0501 ( new_n703_, new_n689_, N1 );
nor g0502 ( new_n704_, new_n702_, new_n703_ );
nand g0503 ( new_n705_, new_n704_, new_n701_ );
nand g0504 ( new_n706_, new_n705_, new_n693_ );
nand g0505 ( new_n707_, new_n700_, new_n706_ );
nand g0506 ( new_n708_, new_n697_, new_n707_ );
nand g0507 ( new_n709_, new_n708_, keyIn_0_28 );
not g0508 ( new_n710_, keyIn_0_28 );
nor g0509 ( new_n711_, new_n700_, new_n706_ );
nor g0510 ( new_n712_, new_n696_, new_n688_ );
nor g0511 ( new_n713_, new_n712_, new_n711_ );
nand g0512 ( new_n714_, new_n713_, new_n710_ );
nand g0513 ( new_n715_, new_n714_, new_n709_ );
not g0514 ( new_n716_, keyIn_0_2 );
not g0515 ( new_n717_, N21 );
nand g0516 ( new_n718_, new_n717_, N17 );
nand g0517 ( new_n719_, new_n281_, N21 );
nand g0518 ( new_n720_, new_n718_, new_n719_ );
nand g0519 ( new_n721_, new_n720_, new_n716_ );
not g0520 ( new_n722_, new_n720_ );
nand g0521 ( new_n723_, new_n722_, keyIn_0_2 );
nand g0522 ( new_n724_, new_n723_, new_n721_ );
not g0523 ( new_n725_, N29 );
nand g0524 ( new_n726_, new_n725_, N25 );
not g0525 ( new_n727_, N25 );
nand g0526 ( new_n728_, new_n727_, N29 );
nand g0527 ( new_n729_, new_n726_, new_n728_ );
nor g0528 ( new_n730_, new_n729_, keyIn_0_3 );
nand g0529 ( new_n731_, new_n729_, keyIn_0_3 );
not g0530 ( new_n732_, new_n731_ );
nor g0531 ( new_n733_, new_n732_, new_n730_ );
nand g0532 ( new_n734_, new_n733_, new_n724_ );
not g0533 ( new_n735_, new_n721_ );
nor g0534 ( new_n736_, new_n720_, new_n716_ );
nor g0535 ( new_n737_, new_n735_, new_n736_ );
not g0536 ( new_n738_, keyIn_0_3 );
not g0537 ( new_n739_, new_n729_ );
nand g0538 ( new_n740_, new_n739_, new_n738_ );
nand g0539 ( new_n741_, new_n740_, new_n731_ );
nand g0540 ( new_n742_, new_n737_, new_n741_ );
nand g0541 ( new_n743_, new_n734_, new_n742_ );
nand g0542 ( new_n744_, new_n743_, keyIn_0_29 );
not g0543 ( new_n745_, keyIn_0_29 );
not g0544 ( new_n746_, new_n743_ );
nand g0545 ( new_n747_, new_n746_, new_n745_ );
nand g0546 ( new_n748_, new_n747_, new_n744_ );
nand g0547 ( new_n749_, new_n748_, new_n715_ );
nor g0548 ( new_n750_, new_n713_, new_n710_ );
nor g0549 ( new_n751_, new_n708_, keyIn_0_28 );
nor g0550 ( new_n752_, new_n750_, new_n751_ );
not g0551 ( new_n753_, new_n744_ );
nor g0552 ( new_n754_, new_n743_, keyIn_0_29 );
nor g0553 ( new_n755_, new_n753_, new_n754_ );
nand g0554 ( new_n756_, new_n755_, new_n752_ );
nand g0555 ( new_n757_, new_n756_, new_n749_ );
nand g0556 ( new_n758_, new_n757_, new_n676_ );
nor g0557 ( new_n759_, new_n755_, new_n752_ );
nor g0558 ( new_n760_, new_n748_, new_n715_ );
nor g0559 ( new_n761_, new_n759_, new_n760_ );
nand g0560 ( new_n762_, new_n761_, keyIn_0_39 );
nand g0561 ( new_n763_, new_n762_, new_n758_ );
nand g0562 ( new_n764_, N133, N137 );
nand g0563 ( new_n765_, new_n764_, keyIn_0_17 );
not g0564 ( new_n766_, new_n765_ );
nor g0565 ( new_n767_, new_n764_, keyIn_0_17 );
nor g0566 ( new_n768_, new_n766_, new_n767_ );
not g0567 ( new_n769_, new_n768_ );
nand g0568 ( new_n770_, new_n763_, new_n769_ );
not g0569 ( new_n771_, new_n758_ );
nor g0570 ( new_n772_, new_n757_, new_n676_ );
nor g0571 ( new_n773_, new_n771_, new_n772_ );
nand g0572 ( new_n774_, new_n773_, new_n768_ );
nand g0573 ( new_n775_, new_n774_, new_n770_ );
nand g0574 ( new_n776_, new_n775_, new_n675_ );
not g0575 ( new_n777_, new_n770_ );
nor g0576 ( new_n778_, new_n763_, new_n769_ );
nor g0577 ( new_n779_, new_n777_, new_n778_ );
nand g0578 ( new_n780_, new_n779_, keyIn_0_51 );
nand g0579 ( new_n781_, new_n780_, new_n776_ );
nand g0580 ( new_n782_, N65, N81 );
not g0581 ( new_n783_, new_n782_ );
nor g0582 ( new_n784_, N65, N81 );
nor g0583 ( new_n785_, new_n783_, new_n784_ );
nand g0584 ( new_n786_, N97, N113 );
not g0585 ( new_n787_, new_n786_ );
nor g0586 ( new_n788_, N97, N113 );
nor g0587 ( new_n789_, new_n787_, new_n788_ );
not g0588 ( new_n790_, new_n789_ );
nor g0589 ( new_n791_, new_n790_, new_n785_ );
nand g0590 ( new_n792_, new_n790_, new_n785_ );
not g0591 ( new_n793_, new_n792_ );
nor g0592 ( new_n794_, new_n793_, new_n791_ );
not g0593 ( new_n795_, new_n794_ );
nand g0594 ( new_n796_, new_n781_, new_n795_ );
nor g0595 ( new_n797_, new_n779_, keyIn_0_51 );
nor g0596 ( new_n798_, new_n775_, new_n675_ );
nor g0597 ( new_n799_, new_n797_, new_n798_ );
nand g0598 ( new_n800_, new_n799_, new_n794_ );
nand g0599 ( new_n801_, new_n800_, new_n796_ );
nand g0600 ( new_n802_, new_n801_, new_n674_ );
nor g0601 ( new_n803_, new_n799_, new_n794_ );
nor g0602 ( new_n804_, new_n781_, new_n795_ );
nor g0603 ( new_n805_, new_n803_, new_n804_ );
nand g0604 ( new_n806_, new_n805_, keyIn_0_59 );
nand g0605 ( new_n807_, new_n806_, new_n802_ );
nor g0606 ( new_n808_, new_n673_, new_n807_ );
nand g0607 ( new_n809_, new_n530_, new_n808_ );
not g0608 ( new_n810_, keyIn_0_61 );
not g0609 ( new_n811_, keyIn_0_41 );
nor g0610 ( new_n812_, new_n752_, new_n564_ );
nor g0611 ( new_n813_, new_n601_, new_n715_ );
nor g0612 ( new_n814_, new_n813_, new_n812_ );
nor g0613 ( new_n815_, new_n814_, new_n811_ );
nand g0614 ( new_n816_, new_n601_, new_n715_ );
nand g0615 ( new_n817_, new_n752_, new_n564_ );
nand g0616 ( new_n818_, new_n816_, new_n817_ );
nor g0617 ( new_n819_, new_n818_, keyIn_0_41 );
nor g0618 ( new_n820_, new_n815_, new_n819_ );
not g0619 ( new_n821_, keyIn_0_19 );
nand g0620 ( new_n822_, N135, N137 );
nand g0621 ( new_n823_, new_n822_, new_n821_ );
not g0622 ( new_n824_, new_n823_ );
nor g0623 ( new_n825_, new_n822_, new_n821_ );
nor g0624 ( new_n826_, new_n824_, new_n825_ );
nor g0625 ( new_n827_, new_n820_, new_n826_ );
nand g0626 ( new_n828_, new_n818_, keyIn_0_41 );
nand g0627 ( new_n829_, new_n814_, new_n811_ );
nand g0628 ( new_n830_, new_n829_, new_n828_ );
not g0629 ( new_n831_, new_n826_ );
nor g0630 ( new_n832_, new_n830_, new_n831_ );
nor g0631 ( new_n833_, new_n827_, new_n832_ );
nor g0632 ( new_n834_, new_n833_, keyIn_0_53 );
not g0633 ( new_n835_, keyIn_0_53 );
nand g0634 ( new_n836_, new_n830_, new_n831_ );
nand g0635 ( new_n837_, new_n820_, new_n826_ );
nand g0636 ( new_n838_, new_n837_, new_n836_ );
nor g0637 ( new_n839_, new_n838_, new_n835_ );
nor g0638 ( new_n840_, new_n834_, new_n839_ );
not g0639 ( new_n841_, keyIn_0_38 );
not g0640 ( new_n842_, keyIn_0_26 );
nand g0641 ( new_n843_, N73, N89 );
not g0642 ( new_n844_, new_n843_ );
nor g0643 ( new_n845_, N73, N89 );
nor g0644 ( new_n846_, new_n844_, new_n845_ );
nor g0645 ( new_n847_, new_n846_, new_n842_ );
nand g0646 ( new_n848_, new_n846_, new_n842_ );
not g0647 ( new_n849_, new_n848_ );
nor g0648 ( new_n850_, new_n849_, new_n847_ );
not g0649 ( new_n851_, new_n850_ );
not g0650 ( new_n852_, keyIn_0_27 );
nand g0651 ( new_n853_, N105, N121 );
not g0652 ( new_n854_, new_n853_ );
nor g0653 ( new_n855_, N105, N121 );
nor g0654 ( new_n856_, new_n854_, new_n855_ );
nor g0655 ( new_n857_, new_n856_, new_n852_ );
nand g0656 ( new_n858_, new_n856_, new_n852_ );
not g0657 ( new_n859_, new_n858_ );
nor g0658 ( new_n860_, new_n859_, new_n857_ );
not g0659 ( new_n861_, new_n860_ );
nand g0660 ( new_n862_, new_n851_, new_n861_ );
not g0661 ( new_n863_, new_n862_ );
nor g0662 ( new_n864_, new_n851_, new_n861_ );
nor g0663 ( new_n865_, new_n863_, new_n864_ );
nor g0664 ( new_n866_, new_n865_, new_n841_ );
nand g0665 ( new_n867_, new_n865_, new_n841_ );
not g0666 ( new_n868_, new_n867_ );
nor g0667 ( new_n869_, new_n868_, new_n866_ );
nor g0668 ( new_n870_, new_n840_, new_n869_ );
nand g0669 ( new_n871_, new_n838_, new_n835_ );
nand g0670 ( new_n872_, new_n833_, keyIn_0_53 );
nand g0671 ( new_n873_, new_n872_, new_n871_ );
not g0672 ( new_n874_, new_n869_ );
nor g0673 ( new_n875_, new_n873_, new_n874_ );
nor g0674 ( new_n876_, new_n870_, new_n875_ );
nor g0675 ( new_n877_, new_n876_, new_n810_ );
nand g0676 ( new_n878_, new_n873_, new_n874_ );
nand g0677 ( new_n879_, new_n840_, new_n869_ );
nand g0678 ( new_n880_, new_n879_, new_n878_ );
nor g0679 ( new_n881_, new_n880_, keyIn_0_61 );
nor g0680 ( new_n882_, new_n877_, new_n881_ );
not g0681 ( new_n883_, keyIn_0_62 );
not g0682 ( new_n884_, keyIn_0_54 );
nand g0683 ( new_n885_, new_n604_, new_n748_ );
nand g0684 ( new_n886_, new_n755_, new_n597_ );
nand g0685 ( new_n887_, new_n885_, new_n886_ );
nand g0686 ( new_n888_, new_n887_, keyIn_0_42 );
not g0687 ( new_n889_, new_n888_ );
nor g0688 ( new_n890_, new_n887_, keyIn_0_42 );
nor g0689 ( new_n891_, new_n889_, new_n890_ );
nand g0690 ( new_n892_, N136, N137 );
nand g0691 ( new_n893_, new_n892_, keyIn_0_20 );
not g0692 ( new_n894_, new_n893_ );
nor g0693 ( new_n895_, new_n892_, keyIn_0_20 );
nor g0694 ( new_n896_, new_n894_, new_n895_ );
not g0695 ( new_n897_, new_n896_ );
nor g0696 ( new_n898_, new_n891_, new_n897_ );
not g0697 ( new_n899_, keyIn_0_42 );
not g0698 ( new_n900_, new_n887_ );
nand g0699 ( new_n901_, new_n900_, new_n899_ );
nand g0700 ( new_n902_, new_n901_, new_n888_ );
nor g0701 ( new_n903_, new_n902_, new_n896_ );
nor g0702 ( new_n904_, new_n898_, new_n903_ );
nor g0703 ( new_n905_, new_n904_, new_n884_ );
nand g0704 ( new_n906_, new_n902_, new_n896_ );
nand g0705 ( new_n907_, new_n891_, new_n897_ );
nand g0706 ( new_n908_, new_n907_, new_n906_ );
nor g0707 ( new_n909_, new_n908_, keyIn_0_54 );
nor g0708 ( new_n910_, new_n905_, new_n909_ );
nand g0709 ( new_n911_, N77, N93 );
not g0710 ( new_n912_, new_n911_ );
nor g0711 ( new_n913_, N77, N93 );
nor g0712 ( new_n914_, new_n912_, new_n913_ );
nand g0713 ( new_n915_, N109, N125 );
not g0714 ( new_n916_, new_n915_ );
nor g0715 ( new_n917_, N109, N125 );
nor g0716 ( new_n918_, new_n916_, new_n917_ );
not g0717 ( new_n919_, new_n918_ );
nor g0718 ( new_n920_, new_n919_, new_n914_ );
nand g0719 ( new_n921_, new_n919_, new_n914_ );
not g0720 ( new_n922_, new_n921_ );
nor g0721 ( new_n923_, new_n922_, new_n920_ );
nor g0722 ( new_n924_, new_n910_, new_n923_ );
nand g0723 ( new_n925_, new_n908_, keyIn_0_54 );
nand g0724 ( new_n926_, new_n904_, new_n884_ );
nand g0725 ( new_n927_, new_n926_, new_n925_ );
not g0726 ( new_n928_, new_n923_ );
nor g0727 ( new_n929_, new_n927_, new_n928_ );
nor g0728 ( new_n930_, new_n924_, new_n929_ );
nor g0729 ( new_n931_, new_n930_, new_n883_ );
nand g0730 ( new_n932_, new_n927_, new_n928_ );
nand g0731 ( new_n933_, new_n910_, new_n923_ );
nand g0732 ( new_n934_, new_n933_, new_n932_ );
nor g0733 ( new_n935_, new_n934_, keyIn_0_62 );
nor g0734 ( new_n936_, new_n931_, new_n935_ );
nand g0735 ( new_n937_, new_n936_, new_n882_ );
nor g0736 ( new_n938_, new_n809_, new_n937_ );
not g0737 ( new_n939_, new_n938_ );
nor g0738 ( new_n940_, new_n939_, new_n302_ );
not g0739 ( new_n941_, new_n940_ );
nand g0740 ( new_n942_, new_n941_, N1 );
nand g0741 ( new_n943_, new_n940_, new_n279_ );
nand g0742 ( N724, new_n942_, new_n943_ );
nor g0743 ( new_n945_, new_n939_, new_n450_ );
not g0744 ( new_n946_, new_n945_ );
nand g0745 ( new_n947_, new_n946_, N5 );
nand g0746 ( new_n948_, new_n945_, new_n689_ );
nand g0747 ( N725, new_n947_, new_n948_ );
nor g0748 ( new_n950_, new_n939_, new_n509_ );
not g0749 ( new_n951_, new_n950_ );
nand g0750 ( new_n952_, new_n951_, N9 );
nand g0751 ( new_n953_, new_n950_, new_n683_ );
nand g0752 ( N726, new_n952_, new_n953_ );
nor g0753 ( new_n955_, new_n939_, new_n380_ );
not g0754 ( new_n956_, new_n955_ );
nand g0755 ( new_n957_, new_n956_, N13 );
nand g0756 ( new_n958_, new_n955_, new_n684_ );
nand g0757 ( N727, new_n957_, new_n958_ );
not g0758 ( new_n960_, keyIn_0_105 );
nand g0759 ( new_n961_, new_n381_, new_n510_ );
nor g0760 ( new_n962_, new_n509_, new_n450_ );
nor g0761 ( new_n963_, new_n962_, new_n301_ );
nand g0762 ( new_n964_, new_n963_, new_n961_ );
nor g0763 ( new_n965_, new_n964_, new_n511_ );
not g0764 ( new_n966_, new_n529_ );
nor g0765 ( new_n967_, new_n965_, new_n966_ );
nand g0766 ( new_n968_, new_n671_, keyIn_0_60 );
nand g0767 ( new_n969_, new_n667_, new_n531_ );
nand g0768 ( new_n970_, new_n969_, new_n968_ );
nor g0769 ( new_n971_, new_n805_, keyIn_0_59 );
nor g0770 ( new_n972_, new_n801_, new_n674_ );
nor g0771 ( new_n973_, new_n971_, new_n972_ );
nand g0772 ( new_n974_, new_n973_, new_n970_ );
nor g0773 ( new_n975_, new_n967_, new_n974_ );
nor g0774 ( new_n976_, new_n936_, new_n882_ );
nand g0775 ( new_n977_, new_n975_, new_n976_ );
nor g0776 ( new_n978_, new_n977_, keyIn_0_76 );
not g0777 ( new_n979_, new_n978_ );
not g0778 ( new_n980_, keyIn_0_76 );
not g0779 ( new_n981_, new_n976_ );
nor g0780 ( new_n982_, new_n809_, new_n981_ );
nor g0781 ( new_n983_, new_n982_, new_n980_ );
nor g0782 ( new_n984_, new_n983_, new_n302_ );
nand g0783 ( new_n985_, new_n984_, new_n979_ );
nand g0784 ( new_n986_, new_n985_, keyIn_0_82 );
not g0785 ( new_n987_, keyIn_0_82 );
nand g0786 ( new_n988_, new_n977_, keyIn_0_76 );
nand g0787 ( new_n989_, new_n988_, new_n301_ );
nor g0788 ( new_n990_, new_n989_, new_n978_ );
nand g0789 ( new_n991_, new_n990_, new_n987_ );
nand g0790 ( new_n992_, new_n986_, new_n991_ );
nand g0791 ( new_n993_, new_n992_, new_n281_ );
nor g0792 ( new_n994_, new_n992_, new_n281_ );
not g0793 ( new_n995_, new_n994_ );
nand g0794 ( new_n996_, new_n995_, new_n993_ );
nand g0795 ( new_n997_, new_n996_, new_n960_ );
not g0796 ( new_n998_, new_n993_ );
nor g0797 ( new_n999_, new_n998_, new_n994_ );
nand g0798 ( new_n1000_, new_n999_, keyIn_0_105 );
nand g0799 ( N728, new_n1000_, new_n997_ );
not g0800 ( new_n1002_, keyIn_0_83 );
nor g0801 ( new_n1003_, new_n983_, new_n450_ );
nand g0802 ( new_n1004_, new_n1003_, new_n979_ );
nand g0803 ( new_n1005_, new_n1004_, new_n1002_ );
nand g0804 ( new_n1006_, new_n988_, new_n514_ );
nor g0805 ( new_n1007_, new_n1006_, new_n978_ );
nand g0806 ( new_n1008_, new_n1007_, keyIn_0_83 );
nand g0807 ( new_n1009_, new_n1005_, new_n1008_ );
nand g0808 ( new_n1010_, new_n1009_, N21 );
nor g0809 ( new_n1011_, new_n1009_, N21 );
not g0810 ( new_n1012_, new_n1011_ );
nand g0811 ( new_n1013_, new_n1012_, new_n1010_ );
nand g0812 ( new_n1014_, new_n1013_, keyIn_0_106 );
not g0813 ( new_n1015_, keyIn_0_106 );
not g0814 ( new_n1016_, new_n1010_ );
nor g0815 ( new_n1017_, new_n1016_, new_n1011_ );
nand g0816 ( new_n1018_, new_n1017_, new_n1015_ );
nand g0817 ( N729, new_n1018_, new_n1014_ );
nor g0818 ( new_n1020_, new_n983_, new_n509_ );
nand g0819 ( new_n1021_, new_n1020_, new_n979_ );
nand g0820 ( new_n1022_, new_n1021_, N25 );
not g0821 ( new_n1023_, new_n1021_ );
nand g0822 ( new_n1024_, new_n1023_, new_n727_ );
nand g0823 ( N730, new_n1024_, new_n1022_ );
not g0824 ( new_n1026_, keyIn_0_84 );
nor g0825 ( new_n1027_, new_n983_, new_n380_ );
nand g0826 ( new_n1028_, new_n1027_, new_n979_ );
nand g0827 ( new_n1029_, new_n1028_, new_n1026_ );
nand g0828 ( new_n1030_, new_n988_, new_n381_ );
nor g0829 ( new_n1031_, new_n1030_, new_n978_ );
nand g0830 ( new_n1032_, new_n1031_, keyIn_0_84 );
nand g0831 ( new_n1033_, new_n1029_, new_n1032_ );
nand g0832 ( new_n1034_, new_n1033_, new_n725_ );
nor g0833 ( new_n1035_, new_n1033_, new_n725_ );
not g0834 ( new_n1036_, new_n1035_ );
nand g0835 ( new_n1037_, new_n1036_, new_n1034_ );
nand g0836 ( new_n1038_, new_n1037_, keyIn_0_107 );
not g0837 ( new_n1039_, keyIn_0_107 );
not g0838 ( new_n1040_, new_n1034_ );
nor g0839 ( new_n1041_, new_n1040_, new_n1035_ );
nand g0840 ( new_n1042_, new_n1041_, new_n1039_ );
nand g0841 ( N731, new_n1042_, new_n1038_ );
not g0842 ( new_n1044_, keyIn_0_108 );
nand g0843 ( new_n1045_, new_n673_, new_n807_ );
nor g0844 ( new_n1046_, new_n937_, new_n1045_ );
nand g0845 ( new_n1047_, new_n530_, new_n1046_ );
nor g0846 ( new_n1048_, new_n1047_, keyIn_0_77 );
nand g0847 ( new_n1049_, new_n1047_, keyIn_0_77 );
nand g0848 ( new_n1050_, new_n1049_, new_n301_ );
nor g0849 ( new_n1051_, new_n1050_, new_n1048_ );
nor g0850 ( new_n1052_, new_n1051_, keyIn_0_85 );
nand g0851 ( new_n1053_, new_n1051_, keyIn_0_85 );
not g0852 ( new_n1054_, new_n1053_ );
nor g0853 ( new_n1055_, new_n1054_, new_n1052_ );
nor g0854 ( new_n1056_, new_n1055_, new_n535_ );
not g0855 ( new_n1057_, new_n1056_ );
nand g0856 ( new_n1058_, new_n1055_, new_n535_ );
nand g0857 ( new_n1059_, new_n1057_, new_n1058_ );
nand g0858 ( new_n1060_, new_n1059_, new_n1044_ );
not g0859 ( new_n1061_, new_n1059_ );
nand g0860 ( new_n1062_, new_n1061_, keyIn_0_108 );
nand g0861 ( N732, new_n1062_, new_n1060_ );
not g0862 ( new_n1064_, keyIn_0_86 );
nand g0863 ( new_n1065_, new_n1049_, new_n514_ );
nor g0864 ( new_n1066_, new_n1065_, new_n1048_ );
nor g0865 ( new_n1067_, new_n1066_, new_n1064_ );
nand g0866 ( new_n1068_, new_n1066_, new_n1064_ );
not g0867 ( new_n1069_, new_n1068_ );
nor g0868 ( new_n1070_, new_n1069_, new_n1067_ );
nor g0869 ( new_n1071_, new_n1070_, new_n533_ );
not g0870 ( new_n1072_, new_n1071_ );
nand g0871 ( new_n1073_, new_n1070_, new_n533_ );
nand g0872 ( new_n1074_, new_n1072_, new_n1073_ );
nand g0873 ( new_n1075_, new_n1074_, keyIn_0_109 );
not g0874 ( new_n1076_, keyIn_0_109 );
not g0875 ( new_n1077_, new_n1074_ );
nand g0876 ( new_n1078_, new_n1077_, new_n1076_ );
nand g0877 ( N733, new_n1078_, new_n1075_ );
not g0878 ( new_n1080_, keyIn_0_110 );
not g0879 ( new_n1081_, keyIn_0_87 );
nand g0880 ( new_n1082_, new_n1049_, new_n516_ );
nor g0881 ( new_n1083_, new_n1082_, new_n1048_ );
nor g0882 ( new_n1084_, new_n1083_, new_n1081_ );
nand g0883 ( new_n1085_, new_n1083_, new_n1081_ );
not g0884 ( new_n1086_, new_n1085_ );
nor g0885 ( new_n1087_, new_n1086_, new_n1084_ );
nor g0886 ( new_n1088_, new_n1087_, N41 );
not g0887 ( new_n1089_, new_n1088_ );
nand g0888 ( new_n1090_, new_n1087_, N41 );
nand g0889 ( new_n1091_, new_n1089_, new_n1090_ );
nand g0890 ( new_n1092_, new_n1091_, new_n1080_ );
not g0891 ( new_n1093_, new_n1091_ );
nand g0892 ( new_n1094_, new_n1093_, keyIn_0_110 );
nand g0893 ( N734, new_n1094_, new_n1092_ );
not g0894 ( new_n1096_, keyIn_0_111 );
not g0895 ( new_n1097_, keyIn_0_88 );
nand g0896 ( new_n1098_, new_n1049_, new_n381_ );
nor g0897 ( new_n1099_, new_n1098_, new_n1048_ );
nor g0898 ( new_n1100_, new_n1099_, new_n1097_ );
nand g0899 ( new_n1101_, new_n1099_, new_n1097_ );
not g0900 ( new_n1102_, new_n1101_ );
nor g0901 ( new_n1103_, new_n1102_, new_n1100_ );
nor g0902 ( new_n1104_, new_n1103_, N45 );
not g0903 ( new_n1105_, new_n1104_ );
nand g0904 ( new_n1106_, new_n1103_, N45 );
nand g0905 ( new_n1107_, new_n1105_, new_n1106_ );
nand g0906 ( new_n1108_, new_n1107_, new_n1096_ );
not g0907 ( new_n1109_, new_n1107_ );
nand g0908 ( new_n1110_, new_n1109_, keyIn_0_111 );
nand g0909 ( N735, new_n1110_, new_n1108_ );
nor g0910 ( new_n1112_, new_n981_, new_n1045_ );
nand g0911 ( new_n1113_, new_n530_, new_n1112_ );
nor g0912 ( new_n1114_, new_n1113_, new_n302_ );
not g0913 ( new_n1115_, new_n1114_ );
nand g0914 ( new_n1116_, new_n1115_, N49 );
nand g0915 ( new_n1117_, new_n1114_, new_n569_ );
nand g0916 ( N736, new_n1116_, new_n1117_ );
nor g0917 ( new_n1119_, new_n1113_, new_n450_ );
not g0918 ( new_n1120_, new_n1119_ );
nand g0919 ( new_n1121_, new_n1120_, N53 );
nand g0920 ( new_n1122_, new_n1119_, new_n567_ );
nand g0921 ( N737, new_n1121_, new_n1122_ );
nor g0922 ( new_n1124_, new_n1113_, new_n509_ );
not g0923 ( new_n1125_, new_n1124_ );
nand g0924 ( new_n1126_, new_n1125_, N57 );
nand g0925 ( new_n1127_, new_n1124_, new_n475_ );
nand g0926 ( N738, new_n1126_, new_n1127_ );
nor g0927 ( new_n1129_, new_n1113_, new_n380_ );
not g0928 ( new_n1130_, new_n1129_ );
nand g0929 ( new_n1131_, new_n1130_, N61 );
nand g0930 ( new_n1132_, new_n1129_, new_n576_ );
nand g0931 ( N739, new_n1131_, new_n1132_ );
not g0932 ( new_n1134_, keyIn_0_112 );
not g0933 ( new_n1135_, N65 );
not g0934 ( new_n1136_, keyIn_0_75 );
nand g0935 ( new_n1137_, new_n880_, keyIn_0_61 );
nand g0936 ( new_n1138_, new_n876_, new_n810_ );
nand g0937 ( new_n1139_, new_n1138_, new_n1137_ );
nand g0938 ( new_n1140_, new_n1139_, keyIn_0_65 );
not g0939 ( new_n1141_, keyIn_0_65 );
nand g0940 ( new_n1142_, new_n882_, new_n1141_ );
nand g0941 ( new_n1143_, new_n1142_, new_n1140_ );
nand g0942 ( new_n1144_, new_n934_, keyIn_0_62 );
nand g0943 ( new_n1145_, new_n930_, new_n883_ );
nand g0944 ( new_n1146_, new_n1145_, new_n1144_ );
nor g0945 ( new_n1147_, new_n1045_, new_n1146_ );
nand g0946 ( new_n1148_, new_n1147_, new_n1143_ );
nor g0947 ( new_n1149_, new_n1148_, keyIn_0_73 );
nor g0948 ( new_n1150_, new_n1146_, new_n1139_ );
nand g0949 ( new_n1151_, new_n970_, new_n807_ );
not g0950 ( new_n1152_, new_n1151_ );
nand g0951 ( new_n1153_, new_n1152_, new_n1150_ );
nand g0952 ( new_n1154_, new_n1153_, keyIn_0_72 );
not g0953 ( new_n1155_, keyIn_0_72 );
nor g0954 ( new_n1156_, new_n937_, new_n1151_ );
nand g0955 ( new_n1157_, new_n1156_, new_n1155_ );
nand g0956 ( new_n1158_, new_n1154_, new_n1157_ );
nand g0957 ( new_n1159_, new_n1148_, keyIn_0_73 );
nand g0958 ( new_n1160_, new_n1158_, new_n1159_ );
nor g0959 ( new_n1161_, new_n1160_, new_n1149_ );
not g0960 ( new_n1162_, keyIn_0_71 );
nand g0961 ( new_n1163_, new_n882_, keyIn_0_64 );
nand g0962 ( new_n1164_, new_n1163_, new_n1146_ );
not g0963 ( new_n1165_, keyIn_0_64 );
nand g0964 ( new_n1166_, new_n1139_, new_n1165_ );
nand g0965 ( new_n1167_, new_n1152_, new_n1166_ );
nor g0966 ( new_n1168_, new_n1167_, new_n1164_ );
nor g0967 ( new_n1169_, new_n1168_, new_n1162_ );
nor g0968 ( new_n1170_, new_n1139_, new_n1165_ );
nor g0969 ( new_n1171_, new_n1170_, new_n936_ );
not g0970 ( new_n1172_, new_n1166_ );
nor g0971 ( new_n1173_, new_n1172_, new_n1151_ );
nand g0972 ( new_n1174_, new_n1173_, new_n1171_ );
nor g0973 ( new_n1175_, new_n1174_, keyIn_0_71 );
nor g0974 ( new_n1176_, new_n1169_, new_n1175_ );
nand g0975 ( new_n1177_, new_n1139_, keyIn_0_66 );
not g0976 ( new_n1178_, keyIn_0_66 );
nand g0977 ( new_n1179_, new_n882_, new_n1178_ );
nand g0978 ( new_n1180_, new_n1179_, new_n1177_ );
nor g0979 ( new_n1181_, new_n974_, new_n1146_ );
nand g0980 ( new_n1182_, new_n1181_, new_n1180_ );
nand g0981 ( new_n1183_, new_n1182_, keyIn_0_74 );
not g0982 ( new_n1184_, new_n1183_ );
nor g0983 ( new_n1185_, new_n1182_, keyIn_0_74 );
nor g0984 ( new_n1186_, new_n1184_, new_n1185_ );
nor g0985 ( new_n1187_, new_n1186_, new_n1176_ );
nand g0986 ( new_n1188_, new_n1187_, new_n1161_ );
nand g0987 ( new_n1189_, new_n1188_, new_n1136_ );
not g0988 ( new_n1190_, new_n1149_ );
not g0989 ( new_n1191_, new_n1160_ );
nand g0990 ( new_n1192_, new_n1191_, new_n1190_ );
nand g0991 ( new_n1193_, new_n1174_, keyIn_0_71 );
nand g0992 ( new_n1194_, new_n1168_, new_n1162_ );
nand g0993 ( new_n1195_, new_n1194_, new_n1193_ );
not g0994 ( new_n1196_, keyIn_0_74 );
not g0995 ( new_n1197_, new_n1182_ );
nand g0996 ( new_n1198_, new_n1197_, new_n1196_ );
nand g0997 ( new_n1199_, new_n1198_, new_n1183_ );
nand g0998 ( new_n1200_, new_n1199_, new_n1195_ );
nor g0999 ( new_n1201_, new_n1192_, new_n1200_ );
nand g1000 ( new_n1202_, new_n1201_, keyIn_0_75 );
nand g1001 ( new_n1203_, new_n1189_, new_n1202_ );
nand g1002 ( new_n1204_, new_n450_, keyIn_0_67 );
not g1003 ( new_n1205_, keyIn_0_67 );
nand g1004 ( new_n1206_, new_n514_, new_n1205_ );
nand g1005 ( new_n1207_, new_n1206_, new_n1204_ );
nand g1006 ( new_n1208_, new_n301_, new_n516_ );
nor g1007 ( new_n1209_, new_n1208_, new_n381_ );
nand g1008 ( new_n1210_, new_n1209_, new_n1207_ );
not g1009 ( new_n1211_, new_n1210_ );
nand g1010 ( new_n1212_, new_n1203_, new_n1211_ );
nand g1011 ( new_n1213_, new_n1212_, keyIn_0_78 );
nor g1012 ( new_n1214_, new_n1212_, keyIn_0_78 );
nor g1013 ( new_n1215_, new_n1214_, new_n807_ );
nand g1014 ( new_n1216_, new_n1215_, new_n1213_ );
nand g1015 ( new_n1217_, new_n1216_, keyIn_0_89 );
nor g1016 ( new_n1218_, new_n1216_, keyIn_0_89 );
not g1017 ( new_n1219_, new_n1218_ );
nand g1018 ( new_n1220_, new_n1219_, new_n1217_ );
nand g1019 ( new_n1221_, new_n1220_, new_n1135_ );
not g1020 ( new_n1222_, new_n1217_ );
nor g1021 ( new_n1223_, new_n1222_, new_n1218_ );
nand g1022 ( new_n1224_, new_n1223_, N65 );
nand g1023 ( new_n1225_, new_n1224_, new_n1221_ );
nand g1024 ( new_n1226_, new_n1225_, new_n1134_ );
not g1025 ( new_n1227_, new_n1225_ );
nand g1026 ( new_n1228_, new_n1227_, keyIn_0_112 );
nand g1027 ( N740, new_n1228_, new_n1226_ );
not g1028 ( new_n1230_, new_n1213_ );
not g1029 ( new_n1231_, keyIn_0_78 );
not g1030 ( new_n1232_, new_n1212_ );
nand g1031 ( new_n1233_, new_n1232_, new_n1231_ );
nand g1032 ( new_n1234_, new_n1233_, new_n673_ );
nor g1033 ( new_n1235_, new_n1234_, new_n1230_ );
nor g1034 ( new_n1236_, new_n1235_, keyIn_0_90 );
not g1035 ( new_n1237_, keyIn_0_90 );
nor g1036 ( new_n1238_, new_n1214_, new_n970_ );
nand g1037 ( new_n1239_, new_n1238_, new_n1213_ );
nor g1038 ( new_n1240_, new_n1239_, new_n1237_ );
nor g1039 ( new_n1241_, new_n1236_, new_n1240_ );
nor g1040 ( new_n1242_, new_n1241_, N69 );
nand g1041 ( new_n1243_, new_n1239_, new_n1237_ );
nand g1042 ( new_n1244_, new_n1235_, keyIn_0_90 );
nand g1043 ( new_n1245_, new_n1244_, new_n1243_ );
nor g1044 ( new_n1246_, new_n1245_, new_n633_ );
nor g1045 ( new_n1247_, new_n1242_, new_n1246_ );
nor g1046 ( new_n1248_, new_n1247_, keyIn_0_113 );
not g1047 ( new_n1249_, keyIn_0_113 );
nand g1048 ( new_n1250_, new_n1245_, new_n633_ );
nand g1049 ( new_n1251_, new_n1241_, N69 );
nand g1050 ( new_n1252_, new_n1251_, new_n1250_ );
nor g1051 ( new_n1253_, new_n1252_, new_n1249_ );
nor g1052 ( N741, new_n1248_, new_n1253_ );
not g1053 ( new_n1255_, N73 );
not g1054 ( new_n1256_, keyIn_0_91 );
nor g1055 ( new_n1257_, new_n1214_, new_n1139_ );
nand g1056 ( new_n1258_, new_n1257_, new_n1213_ );
nand g1057 ( new_n1259_, new_n1258_, new_n1256_ );
nor g1058 ( new_n1260_, new_n1258_, new_n1256_ );
not g1059 ( new_n1261_, new_n1260_ );
nand g1060 ( new_n1262_, new_n1261_, new_n1259_ );
nand g1061 ( new_n1263_, new_n1262_, new_n1255_ );
not g1062 ( new_n1264_, new_n1259_ );
nor g1063 ( new_n1265_, new_n1264_, new_n1260_ );
nand g1064 ( new_n1266_, new_n1265_, N73 );
nand g1065 ( new_n1267_, new_n1266_, new_n1263_ );
nand g1066 ( new_n1268_, new_n1267_, keyIn_0_114 );
not g1067 ( new_n1269_, keyIn_0_114 );
not g1068 ( new_n1270_, new_n1267_ );
nand g1069 ( new_n1271_, new_n1270_, new_n1269_ );
nand g1070 ( N742, new_n1271_, new_n1268_ );
not g1071 ( new_n1273_, N77 );
nor g1072 ( new_n1274_, new_n1214_, new_n936_ );
nand g1073 ( new_n1275_, new_n1274_, new_n1213_ );
nand g1074 ( new_n1276_, new_n1275_, keyIn_0_92 );
nor g1075 ( new_n1277_, new_n1275_, keyIn_0_92 );
not g1076 ( new_n1278_, new_n1277_ );
nand g1077 ( new_n1279_, new_n1278_, new_n1276_ );
nand g1078 ( new_n1280_, new_n1279_, new_n1273_ );
not g1079 ( new_n1281_, new_n1276_ );
nor g1080 ( new_n1282_, new_n1281_, new_n1277_ );
nand g1081 ( new_n1283_, new_n1282_, N77 );
nand g1082 ( new_n1284_, new_n1283_, new_n1280_ );
nand g1083 ( new_n1285_, new_n1284_, keyIn_0_115 );
not g1084 ( new_n1286_, keyIn_0_115 );
not g1085 ( new_n1287_, new_n1284_ );
nand g1086 ( new_n1288_, new_n1287_, new_n1286_ );
nand g1087 ( N743, new_n1288_, new_n1285_ );
not g1088 ( new_n1290_, keyIn_0_79 );
nand g1089 ( new_n1291_, new_n516_, keyIn_0_68 );
not g1090 ( new_n1292_, keyIn_0_68 );
nand g1091 ( new_n1293_, new_n509_, new_n1292_ );
nand g1092 ( new_n1294_, new_n1293_, new_n1291_ );
nor g1093 ( new_n1295_, new_n527_, new_n380_ );
nand g1094 ( new_n1296_, new_n1295_, new_n1294_ );
not g1095 ( new_n1297_, new_n1296_ );
nand g1096 ( new_n1298_, new_n1203_, new_n1297_ );
nor g1097 ( new_n1299_, new_n1298_, new_n1290_ );
nand g1098 ( new_n1300_, new_n1298_, new_n1290_ );
nand g1099 ( new_n1301_, new_n1300_, new_n973_ );
nor g1100 ( new_n1302_, new_n1301_, new_n1299_ );
nor g1101 ( new_n1303_, new_n1302_, keyIn_0_93 );
nand g1102 ( new_n1304_, new_n1302_, keyIn_0_93 );
not g1103 ( new_n1305_, new_n1304_ );
nor g1104 ( new_n1306_, new_n1305_, new_n1303_ );
nor g1105 ( new_n1307_, new_n1306_, N81 );
not g1106 ( new_n1308_, new_n1303_ );
nand g1107 ( new_n1309_, new_n1308_, new_n1304_ );
nor g1108 ( new_n1310_, new_n1309_, new_n233_ );
nor g1109 ( new_n1311_, new_n1307_, new_n1310_ );
nor g1110 ( new_n1312_, new_n1311_, keyIn_0_116 );
not g1111 ( new_n1313_, keyIn_0_116 );
nand g1112 ( new_n1314_, new_n1309_, new_n233_ );
nand g1113 ( new_n1315_, new_n1306_, N81 );
nand g1114 ( new_n1316_, new_n1315_, new_n1314_ );
nor g1115 ( new_n1317_, new_n1316_, new_n1313_ );
nor g1116 ( N744, new_n1312_, new_n1317_ );
not g1117 ( new_n1319_, keyIn_0_94 );
nand g1118 ( new_n1320_, new_n1300_, new_n673_ );
nor g1119 ( new_n1321_, new_n1320_, new_n1299_ );
nor g1120 ( new_n1322_, new_n1321_, new_n1319_ );
nand g1121 ( new_n1323_, new_n1321_, new_n1319_ );
not g1122 ( new_n1324_, new_n1323_ );
nor g1123 ( new_n1325_, new_n1324_, new_n1322_ );
nor g1124 ( new_n1326_, new_n1325_, N85 );
not g1125 ( new_n1327_, new_n1322_ );
nand g1126 ( new_n1328_, new_n1327_, new_n1323_ );
nor g1127 ( new_n1329_, new_n1328_, new_n235_ );
nor g1128 ( new_n1330_, new_n1326_, new_n1329_ );
nor g1129 ( new_n1331_, new_n1330_, keyIn_0_117 );
not g1130 ( new_n1332_, keyIn_0_117 );
nand g1131 ( new_n1333_, new_n1328_, new_n235_ );
nand g1132 ( new_n1334_, new_n1325_, N85 );
nand g1133 ( new_n1335_, new_n1334_, new_n1333_ );
nor g1134 ( new_n1336_, new_n1335_, new_n1332_ );
nor g1135 ( N745, new_n1331_, new_n1336_ );
not g1136 ( new_n1338_, N89 );
not g1137 ( new_n1339_, keyIn_0_95 );
nand g1138 ( new_n1340_, new_n1300_, new_n882_ );
nor g1139 ( new_n1341_, new_n1340_, new_n1299_ );
nor g1140 ( new_n1342_, new_n1341_, new_n1339_ );
nand g1141 ( new_n1343_, new_n1341_, new_n1339_ );
not g1142 ( new_n1344_, new_n1343_ );
nor g1143 ( new_n1345_, new_n1344_, new_n1342_ );
nor g1144 ( new_n1346_, new_n1345_, new_n1338_ );
not g1145 ( new_n1347_, new_n1342_ );
nand g1146 ( new_n1348_, new_n1347_, new_n1343_ );
nor g1147 ( new_n1349_, new_n1348_, N89 );
nor g1148 ( new_n1350_, new_n1346_, new_n1349_ );
nor g1149 ( new_n1351_, new_n1350_, keyIn_0_118 );
not g1150 ( new_n1352_, keyIn_0_118 );
nand g1151 ( new_n1353_, new_n1348_, N89 );
nand g1152 ( new_n1354_, new_n1345_, new_n1338_ );
nand g1153 ( new_n1355_, new_n1354_, new_n1353_ );
nor g1154 ( new_n1356_, new_n1355_, new_n1352_ );
nor g1155 ( N746, new_n1351_, new_n1356_ );
not g1156 ( new_n1358_, keyIn_0_96 );
nand g1157 ( new_n1359_, new_n1300_, new_n1146_ );
nor g1158 ( new_n1360_, new_n1359_, new_n1299_ );
nor g1159 ( new_n1361_, new_n1360_, new_n1358_ );
not g1160 ( new_n1362_, new_n1361_ );
nand g1161 ( new_n1363_, new_n1360_, new_n1358_ );
nand g1162 ( new_n1364_, new_n1362_, new_n1363_ );
nand g1163 ( new_n1365_, new_n1364_, N93 );
nor g1164 ( new_n1366_, new_n1364_, N93 );
not g1165 ( new_n1367_, new_n1366_ );
nand g1166 ( new_n1368_, new_n1367_, new_n1365_ );
nand g1167 ( new_n1369_, new_n1368_, keyIn_0_119 );
not g1168 ( new_n1370_, keyIn_0_119 );
not g1169 ( new_n1371_, new_n1365_ );
nor g1170 ( new_n1372_, new_n1371_, new_n1366_ );
nand g1171 ( new_n1373_, new_n1372_, new_n1370_ );
nand g1172 ( N747, new_n1373_, new_n1369_ );
nand g1173 ( new_n1375_, new_n302_, new_n380_ );
nor g1174 ( new_n1376_, new_n1375_, new_n519_ );
nand g1175 ( new_n1377_, new_n1203_, new_n1376_ );
nor g1176 ( new_n1378_, new_n1377_, keyIn_0_80 );
nand g1177 ( new_n1379_, new_n1377_, keyIn_0_80 );
nand g1178 ( new_n1380_, new_n1379_, new_n973_ );
nor g1179 ( new_n1381_, new_n1380_, new_n1378_ );
nor g1180 ( new_n1382_, new_n1381_, keyIn_0_97 );
not g1181 ( new_n1383_, new_n1382_ );
nand g1182 ( new_n1384_, new_n1381_, keyIn_0_97 );
nand g1183 ( new_n1385_, new_n1383_, new_n1384_ );
nand g1184 ( new_n1386_, new_n1385_, N97 );
nor g1185 ( new_n1387_, new_n1385_, N97 );
not g1186 ( new_n1388_, new_n1387_ );
nand g1187 ( new_n1389_, new_n1388_, new_n1386_ );
nand g1188 ( new_n1390_, new_n1389_, keyIn_0_120 );
not g1189 ( new_n1391_, keyIn_0_120 );
not g1190 ( new_n1392_, new_n1386_ );
nor g1191 ( new_n1393_, new_n1392_, new_n1387_ );
nand g1192 ( new_n1394_, new_n1393_, new_n1391_ );
nand g1193 ( N748, new_n1394_, new_n1390_ );
not g1194 ( new_n1396_, keyIn_0_98 );
nand g1195 ( new_n1397_, new_n1379_, new_n673_ );
nor g1196 ( new_n1398_, new_n1397_, new_n1378_ );
nor g1197 ( new_n1399_, new_n1398_, new_n1396_ );
nand g1198 ( new_n1400_, new_n1398_, new_n1396_ );
not g1199 ( new_n1401_, new_n1400_ );
nor g1200 ( new_n1402_, new_n1401_, new_n1399_ );
nor g1201 ( new_n1403_, new_n1402_, N101 );
not g1202 ( new_n1404_, new_n1399_ );
nand g1203 ( new_n1405_, new_n1404_, new_n1400_ );
nor g1204 ( new_n1406_, new_n1405_, new_n642_ );
nor g1205 ( new_n1407_, new_n1403_, new_n1406_ );
nor g1206 ( new_n1408_, new_n1407_, keyIn_0_121 );
not g1207 ( new_n1409_, keyIn_0_121 );
nand g1208 ( new_n1410_, new_n1405_, new_n642_ );
nand g1209 ( new_n1411_, new_n1402_, N101 );
nand g1210 ( new_n1412_, new_n1411_, new_n1410_ );
nor g1211 ( new_n1413_, new_n1412_, new_n1409_ );
nor g1212 ( N749, new_n1408_, new_n1413_ );
not g1213 ( new_n1415_, keyIn_0_122 );
not g1214 ( new_n1416_, N105 );
nand g1215 ( new_n1417_, new_n1379_, new_n882_ );
nor g1216 ( new_n1418_, new_n1417_, new_n1378_ );
nor g1217 ( new_n1419_, new_n1418_, keyIn_0_99 );
nand g1218 ( new_n1420_, new_n1418_, keyIn_0_99 );
not g1219 ( new_n1421_, new_n1420_ );
nor g1220 ( new_n1422_, new_n1421_, new_n1419_ );
nor g1221 ( new_n1423_, new_n1422_, new_n1416_ );
not g1222 ( new_n1424_, new_n1419_ );
nand g1223 ( new_n1425_, new_n1424_, new_n1420_ );
nor g1224 ( new_n1426_, new_n1425_, N105 );
nor g1225 ( new_n1427_, new_n1423_, new_n1426_ );
nor g1226 ( new_n1428_, new_n1427_, new_n1415_ );
nand g1227 ( new_n1429_, new_n1425_, N105 );
nand g1228 ( new_n1430_, new_n1422_, new_n1416_ );
nand g1229 ( new_n1431_, new_n1430_, new_n1429_ );
nor g1230 ( new_n1432_, new_n1431_, keyIn_0_122 );
nor g1231 ( N750, new_n1428_, new_n1432_ );
not g1232 ( new_n1434_, N109 );
nand g1233 ( new_n1435_, new_n1379_, new_n1146_ );
nor g1234 ( new_n1436_, new_n1435_, new_n1378_ );
nor g1235 ( new_n1437_, new_n1436_, keyIn_0_100 );
nand g1236 ( new_n1438_, new_n1436_, keyIn_0_100 );
not g1237 ( new_n1439_, new_n1438_ );
nor g1238 ( new_n1440_, new_n1439_, new_n1437_ );
nor g1239 ( new_n1441_, new_n1440_, new_n1434_ );
not g1240 ( new_n1442_, new_n1437_ );
nand g1241 ( new_n1443_, new_n1442_, new_n1438_ );
nor g1242 ( new_n1444_, new_n1443_, N109 );
nor g1243 ( new_n1445_, new_n1441_, new_n1444_ );
nor g1244 ( new_n1446_, new_n1445_, keyIn_0_123 );
not g1245 ( new_n1447_, keyIn_0_123 );
nand g1246 ( new_n1448_, new_n1443_, N109 );
nand g1247 ( new_n1449_, new_n1440_, new_n1434_ );
nand g1248 ( new_n1450_, new_n1449_, new_n1448_ );
nor g1249 ( new_n1451_, new_n1450_, new_n1447_ );
nor g1250 ( N751, new_n1446_, new_n1451_ );
not g1251 ( new_n1453_, keyIn_0_124 );
not g1252 ( new_n1454_, keyIn_0_69 );
nand g1253 ( new_n1455_, new_n302_, new_n1454_ );
nor g1254 ( new_n1456_, new_n380_, new_n450_ );
nand g1255 ( new_n1457_, new_n1455_, new_n1456_ );
nand g1256 ( new_n1458_, new_n509_, keyIn_0_70 );
nand g1257 ( new_n1459_, new_n301_, keyIn_0_69 );
not g1258 ( new_n1460_, keyIn_0_70 );
nand g1259 ( new_n1461_, new_n516_, new_n1460_ );
nand g1260 ( new_n1462_, new_n1459_, new_n1461_ );
not g1261 ( new_n1463_, new_n1462_ );
nand g1262 ( new_n1464_, new_n1463_, new_n1458_ );
nor g1263 ( new_n1465_, new_n1464_, new_n1457_ );
nand g1264 ( new_n1466_, new_n1203_, new_n1465_ );
nor g1265 ( new_n1467_, new_n1466_, keyIn_0_81 );
nand g1266 ( new_n1468_, new_n1466_, keyIn_0_81 );
nand g1267 ( new_n1469_, new_n1468_, new_n973_ );
nor g1268 ( new_n1470_, new_n1469_, new_n1467_ );
nor g1269 ( new_n1471_, new_n1470_, keyIn_0_101 );
nand g1270 ( new_n1472_, new_n1470_, keyIn_0_101 );
not g1271 ( new_n1473_, new_n1472_ );
nor g1272 ( new_n1474_, new_n1473_, new_n1471_ );
nor g1273 ( new_n1475_, new_n1474_, N113 );
not g1274 ( new_n1476_, N113 );
not g1275 ( new_n1477_, new_n1471_ );
nand g1276 ( new_n1478_, new_n1477_, new_n1472_ );
nor g1277 ( new_n1479_, new_n1478_, new_n1476_ );
nor g1278 ( new_n1480_, new_n1475_, new_n1479_ );
nor g1279 ( new_n1481_, new_n1480_, new_n1453_ );
nand g1280 ( new_n1482_, new_n1478_, new_n1476_ );
nand g1281 ( new_n1483_, new_n1474_, N113 );
nand g1282 ( new_n1484_, new_n1483_, new_n1482_ );
nor g1283 ( new_n1485_, new_n1484_, keyIn_0_124 );
nor g1284 ( N752, new_n1481_, new_n1485_ );
not g1285 ( new_n1487_, keyIn_0_102 );
nand g1286 ( new_n1488_, new_n1468_, new_n673_ );
nor g1287 ( new_n1489_, new_n1488_, new_n1467_ );
nor g1288 ( new_n1490_, new_n1489_, new_n1487_ );
not g1289 ( new_n1491_, new_n1490_ );
nand g1290 ( new_n1492_, new_n1489_, new_n1487_ );
nand g1291 ( new_n1493_, new_n1491_, new_n1492_ );
nand g1292 ( new_n1494_, new_n1493_, N117 );
nor g1293 ( new_n1495_, new_n1493_, N117 );
not g1294 ( new_n1496_, new_n1495_ );
nand g1295 ( new_n1497_, new_n1496_, new_n1494_ );
nand g1296 ( new_n1498_, new_n1497_, keyIn_0_125 );
not g1297 ( new_n1499_, keyIn_0_125 );
not g1298 ( new_n1500_, new_n1494_ );
nor g1299 ( new_n1501_, new_n1500_, new_n1495_ );
nand g1300 ( new_n1502_, new_n1501_, new_n1499_ );
nand g1301 ( N753, new_n1502_, new_n1498_ );
not g1302 ( new_n1504_, keyIn_0_126 );
not g1303 ( new_n1505_, N121 );
not g1304 ( new_n1506_, keyIn_0_103 );
nand g1305 ( new_n1507_, new_n1468_, new_n882_ );
nor g1306 ( new_n1508_, new_n1507_, new_n1467_ );
nor g1307 ( new_n1509_, new_n1508_, new_n1506_ );
not g1308 ( new_n1510_, new_n1509_ );
nand g1309 ( new_n1511_, new_n1508_, new_n1506_ );
nand g1310 ( new_n1512_, new_n1510_, new_n1511_ );
nand g1311 ( new_n1513_, new_n1512_, new_n1505_ );
nor g1312 ( new_n1514_, new_n1512_, new_n1505_ );
not g1313 ( new_n1515_, new_n1514_ );
nand g1314 ( new_n1516_, new_n1515_, new_n1513_ );
nand g1315 ( new_n1517_, new_n1516_, new_n1504_ );
not g1316 ( new_n1518_, new_n1513_ );
nor g1317 ( new_n1519_, new_n1518_, new_n1514_ );
nand g1318 ( new_n1520_, new_n1519_, keyIn_0_126 );
nand g1319 ( N754, new_n1520_, new_n1517_ );
not g1320 ( new_n1522_, N125 );
not g1321 ( new_n1523_, keyIn_0_104 );
nand g1322 ( new_n1524_, new_n1468_, new_n1146_ );
nor g1323 ( new_n1525_, new_n1524_, new_n1467_ );
nor g1324 ( new_n1526_, new_n1525_, new_n1523_ );
nand g1325 ( new_n1527_, new_n1525_, new_n1523_ );
not g1326 ( new_n1528_, new_n1527_ );
nor g1327 ( new_n1529_, new_n1528_, new_n1526_ );
nor g1328 ( new_n1530_, new_n1529_, new_n1522_ );
not g1329 ( new_n1531_, new_n1526_ );
nand g1330 ( new_n1532_, new_n1531_, new_n1527_ );
nor g1331 ( new_n1533_, new_n1532_, N125 );
nor g1332 ( new_n1534_, new_n1530_, new_n1533_ );
nor g1333 ( new_n1535_, new_n1534_, keyIn_0_127 );
not g1334 ( new_n1536_, keyIn_0_127 );
nand g1335 ( new_n1537_, new_n1532_, N125 );
nand g1336 ( new_n1538_, new_n1529_, new_n1522_ );
nand g1337 ( new_n1539_, new_n1538_, new_n1537_ );
nor g1338 ( new_n1540_, new_n1539_, new_n1536_ );
nor g1339 ( N755, new_n1535_, new_n1540_ );
endmodule