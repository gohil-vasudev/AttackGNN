module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n377_, new_n380_, new_n382_, new_n383_, new_n385_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n394_, new_n395_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n490_, new_n491_, new_n493_, new_n494_, new_n495_, new_n497_, new_n498_, new_n499_, new_n500_, new_n503_, new_n504_, new_n505_, new_n506_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n515_, new_n516_, new_n517_, new_n518_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n535_, new_n536_, new_n538_, new_n539_, new_n540_, new_n542_, new_n543_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_;
  XNOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 g001 ( .A(G132), .ZN(G219) );
  INV_X1 g002 ( .A(G82), .ZN(G220) );
  INV_X1 g003 ( .A(G96), .ZN(G221) );
  INV_X1 g004 ( .A(G69), .ZN(G235) );
  INV_X1 g005 ( .A(G120), .ZN(G236) );
  INV_X1 g006 ( .A(G57), .ZN(G237) );
  INV_X1 g007 ( .A(G108), .ZN(G238) );
  INV_X1 g008 ( .A(G2072), .ZN(new_n367_) );
  INV_X1 g009 ( .A(KEYINPUT21), .ZN(new_n368_) );
  INV_X1 g010 ( .A(G2090), .ZN(new_n369_) );
  AND2_X1 g011 ( .A1(G2078), .A2(G2084), .ZN(new_n370_) );
  XOR2_X1 g012 ( .A(new_n370_), .B(KEYINPUT20), .Z(new_n371_) );
  OR2_X1 g013 ( .A1(new_n371_), .A2(new_n369_), .ZN(new_n372_) );
  AND2_X1 g014 ( .A1(new_n372_), .A2(new_n368_), .ZN(new_n373_) );
  INV_X1 g015 ( .A(new_n372_), .ZN(new_n374_) );
  AND2_X1 g016 ( .A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n375_) );
  OR3_X1 g017 ( .A1(new_n375_), .A2(new_n367_), .A3(new_n373_), .ZN(G158) );
  AND3_X1 g018 ( .A1(G2), .A2(G15), .A3(G661), .ZN(new_n377_) );
  INV_X1 g019 ( .A(new_n377_), .ZN(G259) );
  AND2_X1 g020 ( .A1(G94), .A2(G452), .ZN(G173) );
  AND2_X1 g021 ( .A1(G7), .A2(G661), .ZN(new_n380_) );
  XOR2_X1 g022 ( .A(new_n380_), .B(KEYINPUT10), .Z(G223) );
  INV_X1 g023 ( .A(G567), .ZN(new_n382_) );
  OR2_X1 g024 ( .A1(G223), .A2(new_n382_), .ZN(new_n383_) );
  XOR2_X1 g025 ( .A(new_n383_), .B(KEYINPUT11), .Z(G234) );
  INV_X1 g026 ( .A(G2106), .ZN(new_n385_) );
  OR2_X1 g027 ( .A1(G223), .A2(new_n385_), .ZN(G217) );
  INV_X1 g028 ( .A(G218), .ZN(new_n387_) );
  AND2_X1 g029 ( .A1(G82), .A2(G132), .ZN(new_n388_) );
  XNOR2_X1 g030 ( .A(new_n388_), .B(KEYINPUT22), .ZN(new_n389_) );
  AND3_X1 g031 ( .A1(new_n389_), .A2(G96), .A3(new_n387_), .ZN(new_n390_) );
  AND4_X1 g032 ( .A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n391_) );
  AND2_X1 g033 ( .A1(new_n390_), .A2(new_n391_), .ZN(G325) );
  INV_X1 g034 ( .A(G325), .ZN(G261) );
  OR2_X1 g035 ( .A1(new_n390_), .A2(new_n385_), .ZN(new_n394_) );
  OR2_X1 g036 ( .A1(new_n391_), .A2(new_n382_), .ZN(new_n395_) );
  AND2_X1 g037 ( .A1(new_n394_), .A2(new_n395_), .ZN(G319) );
  INV_X1 g038 ( .A(G137), .ZN(new_n397_) );
  INV_X1 g039 ( .A(KEYINPUT17), .ZN(new_n398_) );
  OR2_X1 g040 ( .A1(G2104), .A2(G2105), .ZN(new_n399_) );
  XNOR2_X1 g041 ( .A(new_n399_), .B(new_n398_), .ZN(new_n400_) );
  OR2_X1 g042 ( .A1(new_n400_), .A2(new_n397_), .ZN(new_n401_) );
  INV_X1 g043 ( .A(G2105), .ZN(new_n402_) );
  AND3_X1 g044 ( .A1(new_n402_), .A2(G101), .A3(G2104), .ZN(new_n403_) );
  XNOR2_X1 g045 ( .A(new_n403_), .B(KEYINPUT23), .ZN(new_n404_) );
  INV_X1 g046 ( .A(G125), .ZN(new_n405_) );
  OR2_X1 g047 ( .A1(new_n402_), .A2(G2104), .ZN(new_n406_) );
  OR2_X1 g048 ( .A1(new_n406_), .A2(new_n405_), .ZN(new_n407_) );
  AND2_X1 g049 ( .A1(G2104), .A2(G2105), .ZN(new_n408_) );
  AND2_X1 g050 ( .A1(new_n408_), .A2(G113), .ZN(new_n409_) );
  INV_X1 g051 ( .A(new_n409_), .ZN(new_n410_) );
  AND2_X1 g052 ( .A1(new_n407_), .A2(new_n410_), .ZN(new_n411_) );
  AND3_X1 g053 ( .A1(new_n401_), .A2(new_n404_), .A3(new_n411_), .ZN(G160) );
  INV_X1 g054 ( .A(G136), .ZN(new_n413_) );
  OR2_X1 g055 ( .A1(new_n400_), .A2(new_n413_), .ZN(new_n414_) );
  INV_X1 g056 ( .A(new_n406_), .ZN(new_n415_) );
  AND2_X1 g057 ( .A1(new_n415_), .A2(G124), .ZN(new_n416_) );
  AND2_X1 g058 ( .A1(new_n416_), .A2(KEYINPUT44), .ZN(new_n417_) );
  INV_X1 g059 ( .A(new_n417_), .ZN(new_n418_) );
  OR2_X1 g060 ( .A1(new_n416_), .A2(KEYINPUT44), .ZN(new_n419_) );
  AND2_X1 g061 ( .A1(new_n408_), .A2(G112), .ZN(new_n420_) );
  INV_X1 g062 ( .A(new_n420_), .ZN(new_n421_) );
  INV_X1 g063 ( .A(G100), .ZN(new_n422_) );
  AND2_X1 g064 ( .A1(new_n402_), .A2(G2104), .ZN(new_n423_) );
  INV_X1 g065 ( .A(new_n423_), .ZN(new_n424_) );
  OR2_X1 g066 ( .A1(new_n424_), .A2(new_n422_), .ZN(new_n425_) );
  AND2_X1 g067 ( .A1(new_n425_), .A2(new_n421_), .ZN(new_n426_) );
  AND4_X1 g068 ( .A1(new_n418_), .A2(new_n414_), .A3(new_n419_), .A4(new_n426_), .ZN(G162) );
  XNOR2_X1 g069 ( .A(new_n399_), .B(KEYINPUT17), .ZN(new_n428_) );
  AND2_X1 g070 ( .A1(new_n428_), .A2(G138), .ZN(new_n429_) );
  AND2_X1 g071 ( .A1(new_n408_), .A2(G114), .ZN(new_n430_) );
  INV_X1 g072 ( .A(G2104), .ZN(new_n431_) );
  AND3_X1 g073 ( .A1(new_n431_), .A2(G126), .A3(G2105), .ZN(new_n432_) );
  AND3_X1 g074 ( .A1(new_n402_), .A2(G102), .A3(G2104), .ZN(new_n433_) );
  OR3_X1 g075 ( .A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_) );
  OR2_X1 g076 ( .A1(new_n429_), .A2(new_n434_), .ZN(new_n435_) );
  INV_X1 g077 ( .A(new_n435_), .ZN(G164) );
  INV_X1 g078 ( .A(G651), .ZN(new_n437_) );
  XNOR2_X1 g079 ( .A(G543), .B(KEYINPUT0), .ZN(new_n438_) );
  AND2_X1 g080 ( .A1(new_n438_), .A2(new_n437_), .ZN(new_n439_) );
  AND2_X1 g081 ( .A1(new_n439_), .A2(G50), .ZN(new_n440_) );
  INV_X1 g082 ( .A(G543), .ZN(new_n441_) );
  AND2_X1 g083 ( .A1(new_n441_), .A2(new_n437_), .ZN(new_n442_) );
  AND2_X1 g084 ( .A1(new_n442_), .A2(G88), .ZN(new_n443_) );
  AND2_X1 g085 ( .A1(new_n441_), .A2(G651), .ZN(new_n444_) );
  XNOR2_X1 g086 ( .A(new_n444_), .B(KEYINPUT1), .ZN(new_n445_) );
  INV_X1 g087 ( .A(new_n445_), .ZN(new_n446_) );
  AND2_X1 g088 ( .A1(new_n446_), .A2(G62), .ZN(new_n447_) );
  AND2_X1 g089 ( .A1(new_n438_), .A2(G651), .ZN(new_n448_) );
  AND2_X1 g090 ( .A1(new_n448_), .A2(G75), .ZN(new_n449_) );
  OR4_X1 g091 ( .A1(new_n447_), .A2(new_n440_), .A3(new_n449_), .A4(new_n443_), .ZN(G303) );
  INV_X1 g092 ( .A(G303), .ZN(G166) );
  AND2_X1 g093 ( .A1(new_n446_), .A2(G63), .ZN(new_n452_) );
  AND2_X1 g094 ( .A1(new_n439_), .A2(G51), .ZN(new_n453_) );
  OR2_X1 g095 ( .A1(new_n452_), .A2(new_n453_), .ZN(new_n454_) );
  XOR2_X1 g096 ( .A(new_n454_), .B(KEYINPUT6), .Z(new_n455_) );
  AND2_X1 g097 ( .A1(new_n442_), .A2(G89), .ZN(new_n456_) );
  XNOR2_X1 g098 ( .A(new_n456_), .B(KEYINPUT4), .ZN(new_n457_) );
  AND2_X1 g099 ( .A1(new_n448_), .A2(G76), .ZN(new_n458_) );
  OR2_X1 g100 ( .A1(new_n457_), .A2(new_n458_), .ZN(new_n459_) );
  XNOR2_X1 g101 ( .A(new_n459_), .B(KEYINPUT5), .ZN(new_n460_) );
  AND2_X1 g102 ( .A1(new_n455_), .A2(new_n460_), .ZN(new_n461_) );
  XOR2_X1 g103 ( .A(new_n461_), .B(KEYINPUT7), .Z(G168) );
  AND2_X1 g104 ( .A1(new_n448_), .A2(G77), .ZN(new_n463_) );
  AND2_X1 g105 ( .A1(new_n442_), .A2(G90), .ZN(new_n464_) );
  OR2_X1 g106 ( .A1(new_n463_), .A2(new_n464_), .ZN(new_n465_) );
  INV_X1 g107 ( .A(new_n465_), .ZN(new_n466_) );
  AND2_X1 g108 ( .A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n467_) );
  OR2_X1 g109 ( .A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n468_) );
  INV_X1 g110 ( .A(new_n468_), .ZN(new_n469_) );
  AND2_X1 g111 ( .A1(new_n446_), .A2(G64), .ZN(new_n470_) );
  AND2_X1 g112 ( .A1(new_n439_), .A2(G52), .ZN(new_n471_) );
  OR4_X1 g113 ( .A1(new_n469_), .A2(new_n467_), .A3(new_n470_), .A4(new_n471_), .ZN(G301) );
  INV_X1 g114 ( .A(G301), .ZN(G171) );
  INV_X1 g115 ( .A(G860), .ZN(new_n474_) );
  AND3_X1 g116 ( .A1(new_n441_), .A2(new_n437_), .A3(G81), .ZN(new_n475_) );
  XNOR2_X1 g117 ( .A(new_n475_), .B(KEYINPUT12), .ZN(new_n476_) );
  AND3_X1 g118 ( .A1(new_n438_), .A2(G68), .A3(G651), .ZN(new_n477_) );
  OR2_X1 g119 ( .A1(new_n476_), .A2(new_n477_), .ZN(new_n478_) );
  XNOR2_X1 g120 ( .A(new_n478_), .B(KEYINPUT13), .ZN(new_n479_) );
  AND2_X1 g121 ( .A1(new_n446_), .A2(G56), .ZN(new_n480_) );
  OR2_X1 g122 ( .A1(new_n480_), .A2(KEYINPUT14), .ZN(new_n481_) );
  AND2_X1 g123 ( .A1(new_n439_), .A2(G43), .ZN(new_n482_) );
  INV_X1 g124 ( .A(new_n482_), .ZN(new_n483_) );
  INV_X1 g125 ( .A(G56), .ZN(new_n484_) );
  INV_X1 g126 ( .A(KEYINPUT14), .ZN(new_n485_) );
  OR3_X1 g127 ( .A1(new_n445_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_) );
  AND4_X1 g128 ( .A1(new_n479_), .A2(new_n481_), .A3(new_n483_), .A4(new_n486_), .ZN(new_n487_) );
  INV_X1 g129 ( .A(new_n487_), .ZN(new_n488_) );
  OR2_X1 g130 ( .A1(new_n488_), .A2(new_n474_), .ZN(G153) );
  AND3_X1 g131 ( .A1(G319), .A2(G483), .A3(G661), .ZN(new_n490_) );
  AND2_X1 g132 ( .A1(new_n490_), .A2(G36), .ZN(new_n491_) );
  INV_X1 g133 ( .A(new_n491_), .ZN(G176) );
  AND2_X1 g134 ( .A1(G1), .A2(G3), .ZN(new_n493_) );
  INV_X1 g135 ( .A(new_n493_), .ZN(new_n494_) );
  AND2_X1 g136 ( .A1(new_n490_), .A2(new_n494_), .ZN(new_n495_) );
  INV_X1 g137 ( .A(new_n495_), .ZN(G188) );
  AND2_X1 g138 ( .A1(new_n448_), .A2(G78), .ZN(new_n497_) );
  AND2_X1 g139 ( .A1(new_n442_), .A2(G91), .ZN(new_n498_) );
  AND2_X1 g140 ( .A1(new_n446_), .A2(G65), .ZN(new_n499_) );
  AND2_X1 g141 ( .A1(new_n439_), .A2(G53), .ZN(new_n500_) );
  OR4_X1 g142 ( .A1(new_n499_), .A2(new_n497_), .A3(new_n498_), .A4(new_n500_), .ZN(G299) );
  XOR2_X1 g143 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 g144 ( .A1(new_n439_), .A2(G49), .ZN(new_n503_) );
  XOR2_X1 g145 ( .A(G543), .B(KEYINPUT0), .Z(new_n504_) );
  AND2_X1 g146 ( .A1(new_n504_), .A2(G87), .ZN(new_n505_) );
  AND2_X1 g147 ( .A1(G74), .A2(G651), .ZN(new_n506_) );
  OR4_X1 g148 ( .A1(new_n503_), .A2(new_n446_), .A3(new_n505_), .A4(new_n506_), .ZN(G288) );
  AND2_X1 g149 ( .A1(new_n439_), .A2(G48), .ZN(new_n508_) );
  AND2_X1 g150 ( .A1(new_n442_), .A2(G86), .ZN(new_n509_) );
  AND2_X1 g151 ( .A1(new_n446_), .A2(G61), .ZN(new_n510_) );
  AND2_X1 g152 ( .A1(new_n448_), .A2(G73), .ZN(new_n511_) );
  XOR2_X1 g153 ( .A(new_n511_), .B(KEYINPUT2), .Z(new_n512_) );
  INV_X1 g154 ( .A(new_n512_), .ZN(new_n513_) );
  OR4_X1 g155 ( .A1(new_n513_), .A2(new_n508_), .A3(new_n509_), .A4(new_n510_), .ZN(G305) );
  AND2_X1 g156 ( .A1(new_n448_), .A2(G72), .ZN(new_n515_) );
  AND2_X1 g157 ( .A1(new_n442_), .A2(G85), .ZN(new_n516_) );
  AND2_X1 g158 ( .A1(new_n446_), .A2(G60), .ZN(new_n517_) );
  AND2_X1 g159 ( .A1(new_n439_), .A2(G47), .ZN(new_n518_) );
  OR4_X1 g160 ( .A1(new_n517_), .A2(new_n515_), .A3(new_n518_), .A4(new_n516_), .ZN(G290) );
  INV_X1 g161 ( .A(G868), .ZN(new_n520_) );
  AND2_X1 g162 ( .A1(new_n439_), .A2(G54), .ZN(new_n521_) );
  INV_X1 g163 ( .A(new_n521_), .ZN(new_n522_) );
  INV_X1 g164 ( .A(G92), .ZN(new_n523_) );
  OR3_X1 g165 ( .A1(new_n523_), .A2(G543), .A3(G651), .ZN(new_n524_) );
  INV_X1 g166 ( .A(G66), .ZN(new_n525_) );
  OR2_X1 g167 ( .A1(new_n445_), .A2(new_n525_), .ZN(new_n526_) );
  AND2_X1 g168 ( .A1(new_n448_), .A2(G79), .ZN(new_n527_) );
  INV_X1 g169 ( .A(new_n527_), .ZN(new_n528_) );
  AND4_X1 g170 ( .A1(new_n522_), .A2(new_n528_), .A3(new_n526_), .A4(new_n524_), .ZN(new_n529_) );
  XOR2_X1 g171 ( .A(new_n529_), .B(KEYINPUT15), .Z(new_n530_) );
  INV_X1 g172 ( .A(new_n530_), .ZN(new_n531_) );
  AND2_X1 g173 ( .A1(new_n531_), .A2(new_n520_), .ZN(new_n532_) );
  AND2_X1 g174 ( .A1(G301), .A2(G868), .ZN(new_n533_) );
  OR2_X1 g175 ( .A1(new_n533_), .A2(new_n532_), .ZN(G284) );
  OR2_X1 g176 ( .A1(G286), .A2(new_n520_), .ZN(new_n535_) );
  OR2_X1 g177 ( .A1(G299), .A2(G868), .ZN(new_n536_) );
  AND2_X1 g178 ( .A1(new_n535_), .A2(new_n536_), .ZN(G297) );
  INV_X1 g179 ( .A(G559), .ZN(new_n538_) );
  OR2_X1 g180 ( .A1(new_n538_), .A2(G860), .ZN(new_n539_) );
  AND2_X1 g181 ( .A1(new_n530_), .A2(new_n539_), .ZN(new_n540_) );
  XOR2_X1 g182 ( .A(new_n540_), .B(KEYINPUT16), .Z(G148) );
  OR2_X1 g183 ( .A1(new_n488_), .A2(G868), .ZN(new_n542_) );
  OR3_X1 g184 ( .A1(new_n531_), .A2(G559), .A3(new_n520_), .ZN(new_n543_) );
  AND2_X1 g185 ( .A1(new_n543_), .A2(new_n542_), .ZN(G282) );
  INV_X1 g186 ( .A(G2100), .ZN(new_n545_) );
  INV_X1 g187 ( .A(G2096), .ZN(new_n546_) );
  INV_X1 g188 ( .A(G135), .ZN(new_n547_) );
  OR2_X1 g189 ( .A1(new_n400_), .A2(new_n547_), .ZN(new_n548_) );
  AND2_X1 g190 ( .A1(new_n415_), .A2(G123), .ZN(new_n549_) );
  AND2_X1 g191 ( .A1(new_n549_), .A2(KEYINPUT18), .ZN(new_n550_) );
  INV_X1 g192 ( .A(new_n550_), .ZN(new_n551_) );
  OR2_X1 g193 ( .A1(new_n549_), .A2(KEYINPUT18), .ZN(new_n552_) );
  AND2_X1 g194 ( .A1(new_n408_), .A2(G111), .ZN(new_n553_) );
  INV_X1 g195 ( .A(new_n553_), .ZN(new_n554_) );
  INV_X1 g196 ( .A(G99), .ZN(new_n555_) );
  OR2_X1 g197 ( .A1(new_n424_), .A2(new_n555_), .ZN(new_n556_) );
  AND4_X1 g198 ( .A1(new_n551_), .A2(new_n552_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n557_) );
  AND2_X1 g199 ( .A1(new_n557_), .A2(new_n548_), .ZN(new_n558_) );
  AND2_X1 g200 ( .A1(new_n558_), .A2(new_n546_), .ZN(new_n559_) );
  INV_X1 g201 ( .A(new_n559_), .ZN(new_n560_) );
  OR2_X1 g202 ( .A1(new_n558_), .A2(new_n546_), .ZN(new_n561_) );
  AND3_X1 g203 ( .A1(new_n560_), .A2(new_n545_), .A3(new_n561_), .ZN(new_n562_) );
  INV_X1 g204 ( .A(new_n562_), .ZN(G156) );
  XNOR2_X1 g205 ( .A(G2430), .B(G2454), .ZN(new_n564_) );
  XNOR2_X1 g206 ( .A(G1341), .B(G1348), .ZN(new_n565_) );
  XNOR2_X1 g207 ( .A(new_n564_), .B(new_n565_), .ZN(new_n566_) );
  XOR2_X1 g208 ( .A(G2435), .B(G2438), .Z(new_n567_) );
  XNOR2_X1 g209 ( .A(new_n566_), .B(new_n567_), .ZN(new_n568_) );
  XOR2_X1 g210 ( .A(G2446), .B(G2451), .Z(new_n569_) );
  XNOR2_X1 g211 ( .A(G2427), .B(G2443), .ZN(new_n570_) );
  XNOR2_X1 g212 ( .A(new_n569_), .B(new_n570_), .ZN(new_n571_) );
  INV_X1 g213 ( .A(new_n571_), .ZN(new_n572_) );
  AND2_X1 g214 ( .A1(new_n568_), .A2(new_n572_), .ZN(new_n573_) );
  INV_X1 g215 ( .A(new_n573_), .ZN(new_n574_) );
  OR2_X1 g216 ( .A1(new_n568_), .A2(new_n572_), .ZN(new_n575_) );
  AND3_X1 g217 ( .A1(new_n574_), .A2(new_n575_), .A3(G14), .ZN(G401) );
  XNOR2_X1 g218 ( .A(G2096), .B(G2100), .ZN(new_n577_) );
  XNOR2_X1 g219 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n578_) );
  XNOR2_X1 g220 ( .A(new_n577_), .B(new_n578_), .ZN(new_n579_) );
  XNOR2_X1 g221 ( .A(G2090), .B(KEYINPUT42), .ZN(new_n580_) );
  XNOR2_X1 g222 ( .A(G2067), .B(G2072), .ZN(new_n581_) );
  XNOR2_X1 g223 ( .A(new_n580_), .B(new_n581_), .ZN(new_n582_) );
  XNOR2_X1 g224 ( .A(new_n579_), .B(new_n582_), .ZN(new_n583_) );
  XOR2_X1 g225 ( .A(G2078), .B(G2084), .Z(new_n584_) );
  XNOR2_X1 g226 ( .A(new_n583_), .B(new_n584_), .ZN(G227) );
  XNOR2_X1 g227 ( .A(G1976), .B(G1981), .ZN(new_n586_) );
  XNOR2_X1 g228 ( .A(G1956), .B(G1966), .ZN(new_n587_) );
  XNOR2_X1 g229 ( .A(new_n586_), .B(new_n587_), .ZN(new_n588_) );
  XNOR2_X1 g230 ( .A(new_n588_), .B(G2474), .ZN(new_n589_) );
  XNOR2_X1 g231 ( .A(G1991), .B(G1996), .ZN(new_n590_) );
  XNOR2_X1 g232 ( .A(new_n589_), .B(new_n590_), .ZN(new_n591_) );
  XOR2_X1 g233 ( .A(G1971), .B(KEYINPUT41), .Z(new_n592_) );
  XNOR2_X1 g234 ( .A(G1961), .B(G1986), .ZN(new_n593_) );
  XOR2_X1 g235 ( .A(new_n592_), .B(new_n593_), .Z(new_n594_) );
  XNOR2_X1 g236 ( .A(new_n591_), .B(new_n594_), .ZN(new_n595_) );
  INV_X1 g237 ( .A(new_n595_), .ZN(G229) );
  INV_X1 g238 ( .A(G29), .ZN(new_n597_) );
  INV_X1 g239 ( .A(KEYINPUT55), .ZN(new_n598_) );
  INV_X1 g240 ( .A(KEYINPUT50), .ZN(new_n599_) );
  AND2_X1 g241 ( .A1(new_n415_), .A2(G127), .ZN(new_n600_) );
  AND2_X1 g242 ( .A1(new_n408_), .A2(G115), .ZN(new_n601_) );
  OR2_X1 g243 ( .A1(new_n600_), .A2(new_n601_), .ZN(new_n602_) );
  XOR2_X1 g244 ( .A(new_n602_), .B(KEYINPUT47), .Z(new_n603_) );
  AND2_X1 g245 ( .A1(new_n423_), .A2(G103), .ZN(new_n604_) );
  AND2_X1 g246 ( .A1(new_n428_), .A2(G139), .ZN(new_n605_) );
  OR3_X1 g247 ( .A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_) );
  OR2_X1 g248 ( .A1(new_n606_), .A2(G2072), .ZN(new_n607_) );
  XOR2_X1 g249 ( .A(new_n435_), .B(G2078), .Z(new_n608_) );
  INV_X1 g250 ( .A(new_n606_), .ZN(new_n609_) );
  OR2_X1 g251 ( .A1(new_n609_), .A2(new_n367_), .ZN(new_n610_) );
  AND3_X1 g252 ( .A1(new_n610_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n611_) );
  AND2_X1 g253 ( .A1(new_n611_), .A2(new_n599_), .ZN(new_n612_) );
  INV_X1 g254 ( .A(new_n612_), .ZN(new_n613_) );
  OR2_X1 g255 ( .A1(new_n611_), .A2(new_n599_), .ZN(new_n614_) );
  AND2_X1 g256 ( .A1(new_n428_), .A2(G131), .ZN(new_n615_) );
  AND2_X1 g257 ( .A1(new_n415_), .A2(G119), .ZN(new_n616_) );
  AND2_X1 g258 ( .A1(new_n408_), .A2(G107), .ZN(new_n617_) );
  AND2_X1 g259 ( .A1(new_n423_), .A2(G95), .ZN(new_n618_) );
  OR4_X1 g260 ( .A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .A4(new_n618_), .ZN(new_n619_) );
  AND2_X1 g261 ( .A1(new_n619_), .A2(G1991), .ZN(new_n620_) );
  INV_X1 g262 ( .A(G141), .ZN(new_n621_) );
  OR2_X1 g263 ( .A1(new_n400_), .A2(new_n621_), .ZN(new_n622_) );
  AND2_X1 g264 ( .A1(new_n423_), .A2(G105), .ZN(new_n623_) );
  AND2_X1 g265 ( .A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n624_) );
  INV_X1 g266 ( .A(new_n624_), .ZN(new_n625_) );
  OR2_X1 g267 ( .A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n626_) );
  AND2_X1 g268 ( .A1(new_n408_), .A2(G117), .ZN(new_n627_) );
  INV_X1 g269 ( .A(new_n627_), .ZN(new_n628_) );
  INV_X1 g270 ( .A(G129), .ZN(new_n629_) );
  OR2_X1 g271 ( .A1(new_n406_), .A2(new_n629_), .ZN(new_n630_) );
  AND4_X1 g272 ( .A1(new_n625_), .A2(new_n626_), .A3(new_n628_), .A4(new_n630_), .ZN(new_n631_) );
  AND2_X1 g273 ( .A1(new_n631_), .A2(new_n622_), .ZN(new_n632_) );
  INV_X1 g274 ( .A(new_n632_), .ZN(new_n633_) );
  AND2_X1 g275 ( .A1(new_n633_), .A2(G1996), .ZN(new_n634_) );
  OR2_X1 g276 ( .A1(new_n634_), .A2(new_n620_), .ZN(new_n635_) );
  INV_X1 g277 ( .A(new_n635_), .ZN(new_n636_) );
  INV_X1 g278 ( .A(G2084), .ZN(new_n637_) );
  OR2_X1 g279 ( .A1(G160), .A2(new_n637_), .ZN(new_n638_) );
  INV_X1 g280 ( .A(new_n558_), .ZN(new_n639_) );
  INV_X1 g281 ( .A(G160), .ZN(new_n640_) );
  OR2_X1 g282 ( .A1(new_n640_), .A2(G2084), .ZN(new_n641_) );
  OR2_X1 g283 ( .A1(new_n619_), .A2(G1991), .ZN(new_n642_) );
  AND3_X1 g284 ( .A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_) );
  AND3_X1 g285 ( .A1(new_n636_), .A2(new_n638_), .A3(new_n643_), .ZN(new_n644_) );
  AND2_X1 g286 ( .A1(new_n428_), .A2(G140), .ZN(new_n645_) );
  AND2_X1 g287 ( .A1(new_n423_), .A2(G104), .ZN(new_n646_) );
  OR2_X1 g288 ( .A1(new_n645_), .A2(new_n646_), .ZN(new_n647_) );
  OR2_X1 g289 ( .A1(new_n647_), .A2(KEYINPUT34), .ZN(new_n648_) );
  AND2_X1 g290 ( .A1(new_n415_), .A2(G128), .ZN(new_n649_) );
  AND2_X1 g291 ( .A1(new_n408_), .A2(G116), .ZN(new_n650_) );
  OR2_X1 g292 ( .A1(new_n649_), .A2(new_n650_), .ZN(new_n651_) );
  XNOR2_X1 g293 ( .A(new_n651_), .B(KEYINPUT35), .ZN(new_n652_) );
  INV_X1 g294 ( .A(KEYINPUT34), .ZN(new_n653_) );
  INV_X1 g295 ( .A(new_n647_), .ZN(new_n654_) );
  OR2_X1 g296 ( .A1(new_n654_), .A2(new_n653_), .ZN(new_n655_) );
  AND3_X1 g297 ( .A1(new_n655_), .A2(new_n648_), .A3(new_n652_), .ZN(new_n656_) );
  XNOR2_X1 g298 ( .A(new_n656_), .B(KEYINPUT36), .ZN(new_n657_) );
  XNOR2_X1 g299 ( .A(G2067), .B(KEYINPUT37), .ZN(new_n658_) );
  AND2_X1 g300 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n659_) );
  INV_X1 g301 ( .A(new_n659_), .ZN(new_n660_) );
  OR2_X1 g302 ( .A1(new_n657_), .A2(new_n658_), .ZN(new_n661_) );
  XNOR2_X1 g303 ( .A(G162), .B(new_n369_), .ZN(new_n662_) );
  INV_X1 g304 ( .A(G1996), .ZN(new_n663_) );
  AND2_X1 g305 ( .A1(new_n632_), .A2(new_n663_), .ZN(new_n664_) );
  OR2_X1 g306 ( .A1(new_n662_), .A2(new_n664_), .ZN(new_n665_) );
  XNOR2_X1 g307 ( .A(new_n665_), .B(KEYINPUT51), .ZN(new_n666_) );
  AND3_X1 g308 ( .A1(new_n660_), .A2(new_n661_), .A3(new_n666_), .ZN(new_n667_) );
  AND4_X1 g309 ( .A1(new_n667_), .A2(new_n613_), .A3(new_n614_), .A4(new_n644_), .ZN(new_n668_) );
  XNOR2_X1 g310 ( .A(new_n668_), .B(KEYINPUT52), .ZN(new_n669_) );
  AND2_X1 g311 ( .A1(new_n669_), .A2(new_n598_), .ZN(new_n670_) );
  OR2_X1 g312 ( .A1(new_n670_), .A2(new_n597_), .ZN(new_n671_) );
  XNOR2_X1 g313 ( .A(G168), .B(G1966), .ZN(new_n672_) );
  INV_X1 g314 ( .A(G1981), .ZN(new_n673_) );
  XNOR2_X1 g315 ( .A(G305), .B(new_n673_), .ZN(new_n674_) );
  AND2_X1 g316 ( .A1(new_n672_), .A2(new_n674_), .ZN(new_n675_) );
  XOR2_X1 g317 ( .A(new_n675_), .B(KEYINPUT57), .Z(new_n676_) );
  XNOR2_X1 g318 ( .A(new_n487_), .B(G1341), .ZN(new_n677_) );
  XNOR2_X1 g319 ( .A(new_n530_), .B(G1348), .ZN(new_n678_) );
  INV_X1 g320 ( .A(G1961), .ZN(new_n679_) );
  XNOR2_X1 g321 ( .A(G301), .B(new_n679_), .ZN(new_n680_) );
  INV_X1 g322 ( .A(G1976), .ZN(new_n681_) );
  INV_X1 g323 ( .A(G288), .ZN(new_n682_) );
  OR2_X1 g324 ( .A1(new_n682_), .A2(new_n681_), .ZN(new_n683_) );
  INV_X1 g325 ( .A(G1956), .ZN(new_n684_) );
  INV_X1 g326 ( .A(G299), .ZN(new_n685_) );
  OR2_X1 g327 ( .A1(new_n685_), .A2(new_n684_), .ZN(new_n686_) );
  AND2_X1 g328 ( .A1(new_n686_), .A2(new_n683_), .ZN(new_n687_) );
  OR2_X1 g329 ( .A1(G299), .A2(G1956), .ZN(new_n688_) );
  INV_X1 g330 ( .A(G1971), .ZN(new_n689_) );
  OR2_X1 g331 ( .A1(G166), .A2(new_n689_), .ZN(new_n690_) );
  AND2_X1 g332 ( .A1(new_n690_), .A2(new_n688_), .ZN(new_n691_) );
  AND2_X1 g333 ( .A1(G166), .A2(new_n689_), .ZN(new_n692_) );
  AND2_X1 g334 ( .A1(new_n682_), .A2(new_n681_), .ZN(new_n693_) );
  OR2_X1 g335 ( .A1(new_n692_), .A2(new_n693_), .ZN(new_n694_) );
  INV_X1 g336 ( .A(new_n694_), .ZN(new_n695_) );
  XOR2_X1 g337 ( .A(G290), .B(G1986), .Z(new_n696_) );
  AND4_X1 g338 ( .A1(new_n695_), .A2(new_n687_), .A3(new_n691_), .A4(new_n696_), .ZN(new_n697_) );
  AND4_X1 g339 ( .A1(new_n697_), .A2(new_n680_), .A3(new_n677_), .A4(new_n678_), .ZN(new_n698_) );
  AND2_X1 g340 ( .A1(new_n676_), .A2(new_n698_), .ZN(new_n699_) );
  XOR2_X1 g341 ( .A(G16), .B(KEYINPUT56), .Z(new_n700_) );
  OR2_X1 g342 ( .A1(new_n699_), .A2(new_n700_), .ZN(new_n701_) );
  XOR2_X1 g343 ( .A(G25), .B(G1991), .Z(new_n702_) );
  OR2_X1 g344 ( .A1(G33), .A2(G2072), .ZN(new_n703_) );
  AND2_X1 g345 ( .A1(new_n703_), .A2(G28), .ZN(new_n704_) );
  AND2_X1 g346 ( .A1(G32), .A2(G1996), .ZN(new_n705_) );
  INV_X1 g347 ( .A(new_n705_), .ZN(new_n706_) );
  AND2_X1 g348 ( .A1(G26), .A2(G2067), .ZN(new_n707_) );
  INV_X1 g349 ( .A(new_n707_), .ZN(new_n708_) );
  AND4_X1 g350 ( .A1(new_n704_), .A2(new_n702_), .A3(new_n706_), .A4(new_n708_), .ZN(new_n709_) );
  INV_X1 g351 ( .A(G27), .ZN(new_n710_) );
  XNOR2_X1 g352 ( .A(G2078), .B(KEYINPUT25), .ZN(new_n711_) );
  OR2_X1 g353 ( .A1(new_n711_), .A2(new_n710_), .ZN(new_n712_) );
  INV_X1 g354 ( .A(new_n711_), .ZN(new_n713_) );
  OR2_X1 g355 ( .A1(new_n713_), .A2(G27), .ZN(new_n714_) );
  OR2_X1 g356 ( .A1(G32), .A2(G1996), .ZN(new_n715_) );
  OR2_X1 g357 ( .A1(G26), .A2(G2067), .ZN(new_n716_) );
  AND2_X1 g358 ( .A1(G33), .A2(G2072), .ZN(new_n717_) );
  INV_X1 g359 ( .A(new_n717_), .ZN(new_n718_) );
  AND3_X1 g360 ( .A1(new_n718_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n719_) );
  AND4_X1 g361 ( .A1(new_n709_), .A2(new_n714_), .A3(new_n712_), .A4(new_n719_), .ZN(new_n720_) );
  OR2_X1 g362 ( .A1(new_n720_), .A2(KEYINPUT53), .ZN(new_n721_) );
  AND2_X1 g363 ( .A1(new_n720_), .A2(KEYINPUT53), .ZN(new_n722_) );
  INV_X1 g364 ( .A(new_n722_), .ZN(new_n723_) );
  XNOR2_X1 g365 ( .A(G2084), .B(KEYINPUT54), .ZN(new_n724_) );
  OR2_X1 g366 ( .A1(new_n724_), .A2(G34), .ZN(new_n725_) );
  XOR2_X1 g367 ( .A(G35), .B(G2090), .Z(new_n726_) );
  INV_X1 g368 ( .A(G34), .ZN(new_n727_) );
  INV_X1 g369 ( .A(new_n724_), .ZN(new_n728_) );
  OR2_X1 g370 ( .A1(new_n728_), .A2(new_n727_), .ZN(new_n729_) );
  AND3_X1 g371 ( .A1(new_n729_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n730_) );
  AND3_X1 g372 ( .A1(new_n723_), .A2(new_n721_), .A3(new_n730_), .ZN(new_n731_) );
  INV_X1 g373 ( .A(new_n731_), .ZN(new_n732_) );
  AND2_X1 g374 ( .A1(new_n732_), .A2(KEYINPUT55), .ZN(new_n733_) );
  AND2_X1 g375 ( .A1(new_n731_), .A2(new_n598_), .ZN(new_n734_) );
  OR3_X1 g376 ( .A1(new_n733_), .A2(G29), .A3(new_n734_), .ZN(new_n735_) );
  XNOR2_X1 g377 ( .A(G1348), .B(KEYINPUT59), .ZN(new_n736_) );
  XNOR2_X1 g378 ( .A(new_n736_), .B(G4), .ZN(new_n737_) );
  XOR2_X1 g379 ( .A(G6), .B(G1981), .Z(new_n738_) );
  XOR2_X1 g380 ( .A(G20), .B(G1956), .Z(new_n739_) );
  XOR2_X1 g381 ( .A(G19), .B(G1341), .Z(new_n740_) );
  AND4_X1 g382 ( .A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .A4(new_n740_), .ZN(new_n741_) );
  XOR2_X1 g383 ( .A(new_n741_), .B(KEYINPUT60), .Z(new_n742_) );
  INV_X1 g384 ( .A(KEYINPUT58), .ZN(new_n743_) );
  XNOR2_X1 g385 ( .A(G22), .B(G1971), .ZN(new_n744_) );
  INV_X1 g386 ( .A(new_n744_), .ZN(new_n745_) );
  XOR2_X1 g387 ( .A(G23), .B(G1976), .Z(new_n746_) );
  XOR2_X1 g388 ( .A(G24), .B(G1986), .Z(new_n747_) );
  AND3_X1 g389 ( .A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_) );
  AND2_X1 g390 ( .A1(new_n748_), .A2(new_n743_), .ZN(new_n749_) );
  OR2_X1 g391 ( .A1(new_n748_), .A2(new_n743_), .ZN(new_n750_) );
  INV_X1 g392 ( .A(new_n750_), .ZN(new_n751_) );
  XNOR2_X1 g393 ( .A(G5), .B(G1961), .ZN(new_n752_) );
  XNOR2_X1 g394 ( .A(G21), .B(G1966), .ZN(new_n753_) );
  OR4_X1 g395 ( .A1(new_n751_), .A2(new_n749_), .A3(new_n752_), .A4(new_n753_), .ZN(new_n754_) );
  OR2_X1 g396 ( .A1(new_n742_), .A2(new_n754_), .ZN(new_n755_) );
  AND2_X1 g397 ( .A1(new_n755_), .A2(KEYINPUT61), .ZN(new_n756_) );
  INV_X1 g398 ( .A(KEYINPUT61), .ZN(new_n757_) );
  INV_X1 g399 ( .A(new_n755_), .ZN(new_n758_) );
  AND2_X1 g400 ( .A1(new_n758_), .A2(new_n757_), .ZN(new_n759_) );
  OR3_X1 g401 ( .A1(new_n759_), .A2(G16), .A3(new_n756_), .ZN(new_n760_) );
  AND3_X1 g402 ( .A1(new_n760_), .A2(G11), .A3(new_n735_), .ZN(new_n761_) );
  AND3_X1 g403 ( .A1(new_n701_), .A2(new_n671_), .A3(new_n761_), .ZN(new_n762_) );
  XNOR2_X1 g404 ( .A(new_n762_), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 g405 ( .A(G311), .ZN(G150) );
  OR3_X1 g406 ( .A1(new_n531_), .A2(new_n488_), .A3(new_n538_), .ZN(new_n765_) );
  AND2_X1 g407 ( .A1(new_n530_), .A2(G559), .ZN(new_n766_) );
  OR2_X1 g408 ( .A1(new_n766_), .A2(new_n487_), .ZN(new_n767_) );
  AND3_X1 g409 ( .A1(new_n767_), .A2(new_n474_), .A3(new_n765_), .ZN(new_n768_) );
  AND2_X1 g410 ( .A1(new_n448_), .A2(G80), .ZN(new_n769_) );
  AND2_X1 g411 ( .A1(new_n442_), .A2(G93), .ZN(new_n770_) );
  AND2_X1 g412 ( .A1(new_n446_), .A2(G67), .ZN(new_n771_) );
  AND2_X1 g413 ( .A1(new_n439_), .A2(G55), .ZN(new_n772_) );
  OR4_X1 g414 ( .A1(new_n771_), .A2(new_n769_), .A3(new_n772_), .A4(new_n770_), .ZN(new_n773_) );
  XOR2_X1 g415 ( .A(new_n768_), .B(new_n773_), .Z(G145) );
  INV_X1 g416 ( .A(G37), .ZN(new_n775_) );
  XNOR2_X1 g417 ( .A(new_n606_), .B(G160), .ZN(new_n776_) );
  XNOR2_X1 g418 ( .A(new_n657_), .B(new_n776_), .ZN(new_n777_) );
  AND2_X1 g419 ( .A1(new_n428_), .A2(G142), .ZN(new_n778_) );
  AND2_X1 g420 ( .A1(new_n423_), .A2(G106), .ZN(new_n779_) );
  OR2_X1 g421 ( .A1(new_n778_), .A2(new_n779_), .ZN(new_n780_) );
  INV_X1 g422 ( .A(new_n780_), .ZN(new_n781_) );
  AND2_X1 g423 ( .A1(new_n781_), .A2(KEYINPUT45), .ZN(new_n782_) );
  INV_X1 g424 ( .A(KEYINPUT45), .ZN(new_n783_) );
  AND2_X1 g425 ( .A1(new_n780_), .A2(new_n783_), .ZN(new_n784_) );
  AND2_X1 g426 ( .A1(new_n408_), .A2(G118), .ZN(new_n785_) );
  AND2_X1 g427 ( .A1(new_n415_), .A2(G130), .ZN(new_n786_) );
  OR4_X1 g428 ( .A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .A4(new_n786_), .ZN(new_n787_) );
  XNOR2_X1 g429 ( .A(new_n787_), .B(new_n632_), .ZN(new_n788_) );
  XNOR2_X1 g430 ( .A(new_n788_), .B(G162), .ZN(new_n789_) );
  XNOR2_X1 g431 ( .A(new_n789_), .B(new_n777_), .ZN(new_n790_) );
  XNOR2_X1 g432 ( .A(new_n558_), .B(new_n619_), .ZN(new_n791_) );
  XNOR2_X1 g433 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(new_n792_) );
  XNOR2_X1 g434 ( .A(new_n791_), .B(new_n792_), .ZN(new_n793_) );
  XNOR2_X1 g435 ( .A(new_n793_), .B(G164), .ZN(new_n794_) );
  INV_X1 g436 ( .A(new_n794_), .ZN(new_n795_) );
  AND2_X1 g437 ( .A1(new_n790_), .A2(new_n795_), .ZN(new_n796_) );
  INV_X1 g438 ( .A(new_n796_), .ZN(new_n797_) );
  OR2_X1 g439 ( .A1(new_n790_), .A2(new_n795_), .ZN(new_n798_) );
  AND3_X1 g440 ( .A1(new_n797_), .A2(new_n775_), .A3(new_n798_), .ZN(G395) );
  XNOR2_X1 g441 ( .A(new_n487_), .B(G290), .ZN(new_n800_) );
  XNOR2_X1 g442 ( .A(new_n800_), .B(G288), .ZN(new_n801_) );
  XNOR2_X1 g443 ( .A(G299), .B(KEYINPUT19), .ZN(new_n802_) );
  XNOR2_X1 g444 ( .A(G305), .B(new_n802_), .ZN(new_n803_) );
  XNOR2_X1 g445 ( .A(new_n801_), .B(new_n803_), .ZN(new_n804_) );
  XOR2_X1 g446 ( .A(G303), .B(new_n773_), .Z(new_n805_) );
  XNOR2_X1 g447 ( .A(new_n804_), .B(new_n805_), .ZN(new_n806_) );
  XNOR2_X1 g448 ( .A(new_n806_), .B(new_n766_), .ZN(new_n807_) );
  AND2_X1 g449 ( .A1(new_n807_), .A2(G868), .ZN(new_n808_) );
  AND2_X1 g450 ( .A1(new_n773_), .A2(new_n520_), .ZN(new_n809_) );
  OR2_X1 g451 ( .A1(new_n808_), .A2(new_n809_), .ZN(G295) );
  XNOR2_X1 g452 ( .A(G286), .B(new_n530_), .ZN(new_n811_) );
  XNOR2_X1 g453 ( .A(new_n811_), .B(new_n806_), .ZN(new_n812_) );
  AND2_X1 g454 ( .A1(new_n812_), .A2(G171), .ZN(new_n813_) );
  INV_X1 g455 ( .A(new_n813_), .ZN(new_n814_) );
  OR2_X1 g456 ( .A1(new_n812_), .A2(G171), .ZN(new_n815_) );
  AND3_X1 g457 ( .A1(new_n814_), .A2(new_n775_), .A3(new_n815_), .ZN(G397) );
  INV_X1 g458 ( .A(KEYINPUT32), .ZN(new_n817_) );
  INV_X1 g459 ( .A(G1348), .ZN(new_n818_) );
  INV_X1 g460 ( .A(G1384), .ZN(new_n819_) );
  AND4_X1 g461 ( .A1(new_n401_), .A2(G40), .A3(new_n404_), .A4(new_n411_), .ZN(new_n820_) );
  AND3_X1 g462 ( .A1(new_n820_), .A2(new_n819_), .A3(new_n435_), .ZN(new_n821_) );
  OR2_X1 g463 ( .A1(new_n821_), .A2(new_n818_), .ZN(new_n822_) );
  AND2_X1 g464 ( .A1(new_n821_), .A2(G2067), .ZN(new_n823_) );
  INV_X1 g465 ( .A(new_n823_), .ZN(new_n824_) );
  AND2_X1 g466 ( .A1(new_n824_), .A2(new_n822_), .ZN(new_n825_) );
  INV_X1 g467 ( .A(KEYINPUT26), .ZN(new_n826_) );
  INV_X1 g468 ( .A(new_n821_), .ZN(new_n827_) );
  OR3_X1 g469 ( .A1(new_n827_), .A2(new_n663_), .A3(new_n826_), .ZN(new_n828_) );
  AND2_X1 g470 ( .A1(new_n435_), .A2(new_n819_), .ZN(new_n829_) );
  AND3_X1 g471 ( .A1(new_n829_), .A2(G1996), .A3(new_n820_), .ZN(new_n830_) );
  OR2_X1 g472 ( .A1(new_n830_), .A2(KEYINPUT26), .ZN(new_n831_) );
  INV_X1 g473 ( .A(G1341), .ZN(new_n832_) );
  OR2_X1 g474 ( .A1(new_n821_), .A2(new_n832_), .ZN(new_n833_) );
  AND2_X1 g475 ( .A1(new_n833_), .A2(new_n487_), .ZN(new_n834_) );
  AND4_X1 g476 ( .A1(new_n834_), .A2(new_n530_), .A3(new_n828_), .A4(new_n831_), .ZN(new_n835_) );
  OR2_X1 g477 ( .A1(new_n835_), .A2(new_n825_), .ZN(new_n836_) );
  AND3_X1 g478 ( .A1(new_n834_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n837_) );
  OR2_X1 g479 ( .A1(new_n837_), .A2(new_n530_), .ZN(new_n838_) );
  AND2_X1 g480 ( .A1(new_n836_), .A2(new_n838_), .ZN(new_n839_) );
  OR3_X1 g481 ( .A1(new_n827_), .A2(new_n367_), .A3(KEYINPUT27), .ZN(new_n840_) );
  OR2_X1 g482 ( .A1(new_n821_), .A2(new_n684_), .ZN(new_n841_) );
  INV_X1 g483 ( .A(KEYINPUT27), .ZN(new_n842_) );
  AND2_X1 g484 ( .A1(new_n821_), .A2(G2072), .ZN(new_n843_) );
  OR2_X1 g485 ( .A1(new_n843_), .A2(new_n842_), .ZN(new_n844_) );
  AND3_X1 g486 ( .A1(new_n844_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n845_) );
  AND2_X1 g487 ( .A1(new_n845_), .A2(new_n685_), .ZN(new_n846_) );
  OR2_X1 g488 ( .A1(new_n839_), .A2(new_n846_), .ZN(new_n847_) );
  OR2_X1 g489 ( .A1(new_n845_), .A2(new_n685_), .ZN(new_n848_) );
  XNOR2_X1 g490 ( .A(new_n848_), .B(KEYINPUT28), .ZN(new_n849_) );
  AND2_X1 g491 ( .A1(new_n847_), .A2(new_n849_), .ZN(new_n850_) );
  XNOR2_X1 g492 ( .A(new_n850_), .B(KEYINPUT29), .ZN(new_n851_) );
  AND2_X1 g493 ( .A1(new_n827_), .A2(new_n679_), .ZN(new_n852_) );
  AND2_X1 g494 ( .A1(new_n821_), .A2(new_n711_), .ZN(new_n853_) );
  OR2_X1 g495 ( .A1(new_n852_), .A2(new_n853_), .ZN(new_n854_) );
  AND2_X1 g496 ( .A1(G171), .A2(new_n854_), .ZN(new_n855_) );
  INV_X1 g497 ( .A(new_n855_), .ZN(new_n856_) );
  AND2_X1 g498 ( .A1(new_n851_), .A2(new_n856_), .ZN(new_n857_) );
  INV_X1 g499 ( .A(G168), .ZN(new_n858_) );
  INV_X1 g500 ( .A(G8), .ZN(new_n859_) );
  AND2_X1 g501 ( .A1(new_n827_), .A2(G8), .ZN(new_n860_) );
  INV_X1 g502 ( .A(new_n860_), .ZN(new_n861_) );
  OR2_X1 g503 ( .A1(new_n861_), .A2(G1966), .ZN(new_n862_) );
  INV_X1 g504 ( .A(new_n862_), .ZN(new_n863_) );
  AND2_X1 g505 ( .A1(new_n821_), .A2(new_n637_), .ZN(new_n864_) );
  OR4_X1 g506 ( .A1(new_n863_), .A2(new_n859_), .A3(KEYINPUT30), .A4(new_n864_), .ZN(new_n865_) );
  INV_X1 g507 ( .A(KEYINPUT30), .ZN(new_n866_) );
  INV_X1 g508 ( .A(new_n864_), .ZN(new_n867_) );
  AND3_X1 g509 ( .A1(new_n862_), .A2(G8), .A3(new_n867_), .ZN(new_n868_) );
  OR2_X1 g510 ( .A1(new_n868_), .A2(new_n866_), .ZN(new_n869_) );
  AND3_X1 g511 ( .A1(new_n869_), .A2(new_n858_), .A3(new_n865_), .ZN(new_n870_) );
  INV_X1 g512 ( .A(new_n854_), .ZN(new_n871_) );
  AND2_X1 g513 ( .A1(new_n871_), .A2(G301), .ZN(new_n872_) );
  OR2_X1 g514 ( .A1(new_n870_), .A2(new_n872_), .ZN(new_n873_) );
  XOR2_X1 g515 ( .A(new_n873_), .B(KEYINPUT31), .Z(new_n874_) );
  OR2_X1 g516 ( .A1(new_n857_), .A2(new_n874_), .ZN(new_n875_) );
  AND2_X1 g517 ( .A1(new_n875_), .A2(G286), .ZN(new_n876_) );
  OR2_X1 g518 ( .A1(new_n861_), .A2(G1971), .ZN(new_n877_) );
  AND2_X1 g519 ( .A1(new_n821_), .A2(new_n369_), .ZN(new_n878_) );
  INV_X1 g520 ( .A(new_n878_), .ZN(new_n879_) );
  AND3_X1 g521 ( .A1(new_n877_), .A2(G303), .A3(new_n879_), .ZN(new_n880_) );
  OR2_X1 g522 ( .A1(new_n876_), .A2(new_n880_), .ZN(new_n881_) );
  AND2_X1 g523 ( .A1(new_n881_), .A2(G8), .ZN(new_n882_) );
  XNOR2_X1 g524 ( .A(new_n882_), .B(new_n817_), .ZN(new_n883_) );
  INV_X1 g525 ( .A(new_n875_), .ZN(new_n884_) );
  AND2_X1 g526 ( .A1(new_n864_), .A2(G8), .ZN(new_n885_) );
  OR3_X1 g527 ( .A1(new_n884_), .A2(new_n863_), .A3(new_n885_), .ZN(new_n886_) );
  AND2_X1 g528 ( .A1(new_n883_), .A2(new_n886_), .ZN(new_n887_) );
  OR2_X1 g529 ( .A1(new_n887_), .A2(new_n694_), .ZN(new_n888_) );
  AND2_X1 g530 ( .A1(new_n860_), .A2(new_n683_), .ZN(new_n889_) );
  AND2_X1 g531 ( .A1(new_n888_), .A2(new_n889_), .ZN(new_n890_) );
  OR2_X1 g532 ( .A1(new_n890_), .A2(KEYINPUT33), .ZN(new_n891_) );
  INV_X1 g533 ( .A(KEYINPUT33), .ZN(new_n892_) );
  OR4_X1 g534 ( .A1(new_n861_), .A2(G1976), .A3(new_n892_), .A4(G288), .ZN(new_n893_) );
  AND2_X1 g535 ( .A1(new_n893_), .A2(new_n674_), .ZN(new_n894_) );
  AND2_X1 g536 ( .A1(new_n891_), .A2(new_n894_), .ZN(new_n895_) );
  AND3_X1 g537 ( .A1(G166), .A2(G8), .A3(new_n369_), .ZN(new_n896_) );
  OR2_X1 g538 ( .A1(new_n887_), .A2(new_n896_), .ZN(new_n897_) );
  AND2_X1 g539 ( .A1(new_n897_), .A2(new_n861_), .ZN(new_n898_) );
  INV_X1 g540 ( .A(KEYINPUT24), .ZN(new_n899_) );
  INV_X1 g541 ( .A(G305), .ZN(new_n900_) );
  AND2_X1 g542 ( .A1(new_n900_), .A2(new_n673_), .ZN(new_n901_) );
  OR2_X1 g543 ( .A1(new_n901_), .A2(new_n899_), .ZN(new_n902_) );
  AND2_X1 g544 ( .A1(new_n901_), .A2(new_n899_), .ZN(new_n903_) );
  INV_X1 g545 ( .A(new_n903_), .ZN(new_n904_) );
  AND3_X1 g546 ( .A1(new_n904_), .A2(new_n860_), .A3(new_n902_), .ZN(new_n905_) );
  OR2_X1 g547 ( .A1(new_n898_), .A2(new_n905_), .ZN(new_n906_) );
  OR2_X1 g548 ( .A1(new_n895_), .A2(new_n906_), .ZN(new_n907_) );
  INV_X1 g549 ( .A(new_n829_), .ZN(new_n908_) );
  AND2_X1 g550 ( .A1(new_n908_), .A2(new_n820_), .ZN(new_n909_) );
  INV_X1 g551 ( .A(new_n909_), .ZN(new_n910_) );
  OR2_X1 g552 ( .A1(new_n661_), .A2(new_n910_), .ZN(new_n911_) );
  AND2_X1 g553 ( .A1(new_n635_), .A2(new_n909_), .ZN(new_n912_) );
  INV_X1 g554 ( .A(new_n912_), .ZN(new_n913_) );
  OR2_X1 g555 ( .A1(new_n696_), .A2(new_n910_), .ZN(new_n914_) );
  AND3_X1 g556 ( .A1(new_n911_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_) );
  AND2_X1 g557 ( .A1(new_n907_), .A2(new_n915_), .ZN(new_n916_) );
  INV_X1 g558 ( .A(new_n664_), .ZN(new_n917_) );
  OR2_X1 g559 ( .A1(G290), .A2(G1986), .ZN(new_n918_) );
  AND2_X1 g560 ( .A1(new_n918_), .A2(new_n642_), .ZN(new_n919_) );
  OR2_X1 g561 ( .A1(new_n912_), .A2(new_n919_), .ZN(new_n920_) );
  AND2_X1 g562 ( .A1(new_n920_), .A2(new_n917_), .ZN(new_n921_) );
  INV_X1 g563 ( .A(new_n921_), .ZN(new_n922_) );
  OR2_X1 g564 ( .A1(new_n922_), .A2(KEYINPUT39), .ZN(new_n923_) );
  INV_X1 g565 ( .A(KEYINPUT39), .ZN(new_n924_) );
  OR2_X1 g566 ( .A1(new_n921_), .A2(new_n924_), .ZN(new_n925_) );
  AND3_X1 g567 ( .A1(new_n923_), .A2(new_n911_), .A3(new_n925_), .ZN(new_n926_) );
  OR2_X1 g568 ( .A1(new_n926_), .A2(new_n659_), .ZN(new_n927_) );
  AND2_X1 g569 ( .A1(new_n927_), .A2(new_n909_), .ZN(new_n928_) );
  OR2_X1 g570 ( .A1(new_n916_), .A2(new_n928_), .ZN(new_n929_) );
  XNOR2_X1 g571 ( .A(new_n929_), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 g572 ( .A(G401), .ZN(new_n932_) );
  OR2_X1 g573 ( .A1(G229), .A2(G227), .ZN(new_n933_) );
  INV_X1 g574 ( .A(new_n933_), .ZN(new_n934_) );
  AND2_X1 g575 ( .A1(new_n934_), .A2(KEYINPUT49), .ZN(new_n935_) );
  INV_X1 g576 ( .A(new_n935_), .ZN(new_n936_) );
  OR2_X1 g577 ( .A1(new_n934_), .A2(KEYINPUT49), .ZN(new_n937_) );
  AND4_X1 g578 ( .A1(new_n936_), .A2(G319), .A3(new_n932_), .A4(new_n937_), .ZN(new_n938_) );
  INV_X1 g579 ( .A(new_n938_), .ZN(new_n939_) );
  OR3_X1 g580 ( .A1(G397), .A2(G395), .A3(new_n939_), .ZN(G225) );
  INV_X1 g581 ( .A(G225), .ZN(G308) );
  assign   G231 = 1'b0;
  BUF_X1 g582 ( .A(G452), .Z(G350) );
  BUF_X1 g583 ( .A(G452), .Z(G335) );
  BUF_X1 g584 ( .A(G452), .Z(G409) );
  BUF_X1 g585 ( .A(G1083), .Z(G369) );
  BUF_X1 g586 ( .A(G1083), .Z(G367) );
  BUF_X1 g587 ( .A(G2066), .Z(G411) );
  BUF_X1 g588 ( .A(G2066), .Z(G337) );
  BUF_X1 g589 ( .A(G2066), .Z(G384) );
  BUF_X1 g590 ( .A(G452), .Z(G391) );
  OR2_X1 g591 ( .A1(new_n533_), .A2(new_n532_), .ZN(G321) );
  AND2_X1 g592 ( .A1(new_n535_), .A2(new_n536_), .ZN(G280) );
  AND2_X1 g593 ( .A1(new_n543_), .A2(new_n542_), .ZN(G323) );
  OR2_X1 g594 ( .A1(new_n808_), .A2(new_n809_), .ZN(G331) );
endmodule


