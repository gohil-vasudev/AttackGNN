module add_mul_mix_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, 
        c_9_, c_10_, c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, 
        d_4_, d_5_, d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, 
        d_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_, c_7_, c_8_, c_9_, c_10_,
         c_11_, c_12_, c_13_, c_14_, c_15_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_,
         d_6_, d_7_, d_8_, d_9_, d_10_, d_11_, d_12_, d_13_, d_14_, d_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995;

  OR2_X1 U2036 ( .A1(n2406), .A2(n2480), .ZN(n2609) );
  XNOR2_X2 U2037 ( .A(n3788), .B(n3789), .ZN(n2187) );
  XOR2_X2 U2038 ( .A(n2685), .B(n2686), .Z(n2406) );
  XNOR2_X2 U2039 ( .A(n3919), .B(n3920), .ZN(n3669) );
  XOR2_X2 U2040 ( .A(n2547), .B(n2598), .Z(n2050) );
  XNOR2_X1 U2041 ( .A(n2005), .B(n2006), .ZN(Result_9_) );
  OR2_X1 U2042 ( .A1(n2007), .A2(n2008), .ZN(n2005) );
  AND2_X1 U2043 ( .A1(n2009), .A2(n2010), .ZN(n2007) );
  XOR2_X1 U2044 ( .A(n2011), .B(n2012), .Z(Result_8_) );
  XOR2_X1 U2045 ( .A(n2013), .B(n2014), .Z(Result_7_) );
  AND2_X1 U2046 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
  OR2_X1 U2047 ( .A1(n2017), .A2(n2018), .ZN(n2016) );
  INV_X1 U2048 ( .A(n2019), .ZN(n2015) );
  XOR2_X1 U2049 ( .A(n2020), .B(n2021), .Z(Result_6_) );
  XOR2_X1 U2050 ( .A(n2022), .B(n2023), .Z(Result_5_) );
  AND2_X1 U2051 ( .A1(n2024), .A2(n2025), .ZN(n2023) );
  OR2_X1 U2052 ( .A1(n2026), .A2(n2027), .ZN(n2025) );
  INV_X1 U2053 ( .A(n2028), .ZN(n2024) );
  XOR2_X1 U2054 ( .A(n2029), .B(n2030), .Z(Result_4_) );
  XOR2_X1 U2055 ( .A(n2031), .B(n2032), .Z(Result_3_) );
  AND2_X1 U2056 ( .A1(n2033), .A2(n2034), .ZN(n2032) );
  OR2_X1 U2057 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  INV_X1 U2058 ( .A(n2037), .ZN(n2033) );
  AND2_X1 U2059 ( .A1(n2038), .A2(n2039), .ZN(Result_31_) );
  OR2_X1 U2060 ( .A1(n2040), .A2(n2041), .ZN(Result_30_) );
  AND2_X1 U2061 ( .A1(n2042), .A2(n2043), .ZN(n2041) );
  OR2_X1 U2062 ( .A1(n2044), .A2(n2045), .ZN(n2043) );
  AND2_X1 U2063 ( .A1(n2039), .A2(n2046), .ZN(n2044) );
  AND2_X1 U2064 ( .A1(n2038), .A2(n2047), .ZN(n2040) );
  OR2_X1 U2065 ( .A1(n2048), .A2(n2049), .ZN(n2047) );
  AND2_X1 U2066 ( .A1(n2050), .A2(n2051), .ZN(n2048) );
  XOR2_X1 U2067 ( .A(n2052), .B(n2053), .Z(Result_2_) );
  XNOR2_X1 U2068 ( .A(n2054), .B(n2055), .ZN(Result_29_) );
  XNOR2_X1 U2069 ( .A(n2056), .B(n2057), .ZN(n2054) );
  XNOR2_X1 U2070 ( .A(n2058), .B(n2059), .ZN(Result_28_) );
  XOR2_X1 U2071 ( .A(n2060), .B(n2061), .Z(n2059) );
  XNOR2_X1 U2072 ( .A(n2062), .B(n2063), .ZN(Result_27_) );
  XOR2_X1 U2073 ( .A(n2064), .B(n2065), .Z(n2063) );
  XNOR2_X1 U2074 ( .A(n2066), .B(n2067), .ZN(Result_26_) );
  XOR2_X1 U2075 ( .A(n2068), .B(n2069), .Z(n2067) );
  XNOR2_X1 U2076 ( .A(n2070), .B(n2071), .ZN(Result_25_) );
  XOR2_X1 U2077 ( .A(n2072), .B(n2073), .Z(n2071) );
  XNOR2_X1 U2078 ( .A(n2074), .B(n2075), .ZN(Result_24_) );
  XOR2_X1 U2079 ( .A(n2076), .B(n2077), .Z(n2075) );
  XOR2_X1 U2080 ( .A(n2078), .B(n2079), .Z(Result_23_) );
  XNOR2_X1 U2081 ( .A(n2080), .B(n2081), .ZN(n2078) );
  XOR2_X1 U2082 ( .A(n2082), .B(n2083), .Z(Result_22_) );
  XNOR2_X1 U2083 ( .A(n2084), .B(n2085), .ZN(n2082) );
  XOR2_X1 U2084 ( .A(n2086), .B(n2087), .Z(Result_21_) );
  XNOR2_X1 U2085 ( .A(n2088), .B(n2089), .ZN(n2086) );
  XOR2_X1 U2086 ( .A(n2090), .B(n2091), .Z(Result_20_) );
  XNOR2_X1 U2087 ( .A(n2092), .B(n2093), .ZN(n2090) );
  XOR2_X1 U2088 ( .A(n2094), .B(n2095), .Z(Result_1_) );
  AND2_X1 U2089 ( .A1(n2096), .A2(n2097), .ZN(n2095) );
  OR2_X1 U2090 ( .A1(n2098), .A2(n2099), .ZN(n2097) );
  AND2_X1 U2091 ( .A1(n2100), .A2(n2101), .ZN(n2098) );
  INV_X1 U2092 ( .A(n2102), .ZN(n2096) );
  XOR2_X1 U2093 ( .A(n2103), .B(n2104), .Z(Result_19_) );
  XNOR2_X1 U2094 ( .A(n2105), .B(n2106), .ZN(n2103) );
  XOR2_X1 U2095 ( .A(n2107), .B(n2108), .Z(Result_18_) );
  XNOR2_X1 U2096 ( .A(n2109), .B(n2110), .ZN(n2107) );
  XOR2_X1 U2097 ( .A(n2111), .B(n2112), .Z(Result_17_) );
  XNOR2_X1 U2098 ( .A(n2113), .B(n2114), .ZN(n2111) );
  XOR2_X1 U2099 ( .A(n2115), .B(n2116), .Z(Result_16_) );
  XNOR2_X1 U2100 ( .A(n2117), .B(n2118), .ZN(n2115) );
  XNOR2_X1 U2101 ( .A(n2119), .B(n2120), .ZN(Result_15_) );
  AND2_X1 U2102 ( .A1(n2121), .A2(n2122), .ZN(Result_14_) );
  INV_X1 U2103 ( .A(n2123), .ZN(n2122) );
  OR2_X1 U2104 ( .A1(n2124), .A2(n2125), .ZN(n2121) );
  AND2_X1 U2105 ( .A1(n2126), .A2(n2120), .ZN(n2124) );
  XOR2_X1 U2106 ( .A(n2127), .B(n2128), .Z(Result_13_) );
  OR2_X1 U2107 ( .A1(n2123), .A2(n2129), .ZN(n2127) );
  XNOR2_X1 U2108 ( .A(n2130), .B(n2131), .ZN(Result_12_) );
  OR2_X1 U2109 ( .A1(n2132), .A2(n2133), .ZN(n2130) );
  AND2_X1 U2110 ( .A1(n2134), .A2(n2135), .ZN(n2132) );
  OR2_X1 U2111 ( .A1(n2136), .A2(n2137), .ZN(n2135) );
  XNOR2_X1 U2112 ( .A(n2138), .B(n2139), .ZN(Result_11_) );
  OR2_X1 U2113 ( .A1(n2140), .A2(n2141), .ZN(n2138) );
  AND2_X1 U2114 ( .A1(n2142), .A2(n2143), .ZN(n2140) );
  OR2_X1 U2115 ( .A1(n2144), .A2(n2145), .ZN(n2143) );
  XNOR2_X1 U2116 ( .A(n2146), .B(n2147), .ZN(Result_10_) );
  OR2_X1 U2117 ( .A1(n2148), .A2(n2149), .ZN(n2146) );
  AND2_X1 U2118 ( .A1(n2150), .A2(n2151), .ZN(n2148) );
  OR2_X1 U2119 ( .A1(n2152), .A2(n2153), .ZN(n2151) );
  OR2_X1 U2120 ( .A1(n2154), .A2(n2155), .ZN(Result_0_) );
  OR2_X1 U2121 ( .A1(n2102), .A2(n2156), .ZN(n2155) );
  AND2_X1 U2122 ( .A1(n2094), .A2(n2099), .ZN(n2156) );
  AND2_X1 U2123 ( .A1(n2052), .A2(n2053), .ZN(n2094) );
  XNOR2_X1 U2124 ( .A(n2101), .B(n2157), .ZN(n2053) );
  OR2_X1 U2125 ( .A1(n2158), .A2(n2159), .ZN(n2052) );
  OR2_X1 U2126 ( .A1(n2160), .A2(n2037), .ZN(n2158) );
  AND2_X1 U2127 ( .A1(n2035), .A2(n2036), .ZN(n2037) );
  AND2_X1 U2128 ( .A1(n2161), .A2(n2162), .ZN(n2036) );
  INV_X1 U2129 ( .A(n2163), .ZN(n2161) );
  AND2_X1 U2130 ( .A1(n2031), .A2(n2035), .ZN(n2160) );
  INV_X1 U2131 ( .A(n2164), .ZN(n2035) );
  OR2_X1 U2132 ( .A1(n2165), .A2(n2159), .ZN(n2164) );
  INV_X1 U2133 ( .A(n2166), .ZN(n2159) );
  OR2_X1 U2134 ( .A1(n2167), .A2(n2168), .ZN(n2166) );
  AND2_X1 U2135 ( .A1(n2167), .A2(n2168), .ZN(n2165) );
  OR2_X1 U2136 ( .A1(n2169), .A2(n2170), .ZN(n2168) );
  AND2_X1 U2137 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
  AND2_X1 U2138 ( .A1(n2173), .A2(n2174), .ZN(n2169) );
  OR2_X1 U2139 ( .A1(n2172), .A2(n2171), .ZN(n2174) );
  XOR2_X1 U2140 ( .A(n2175), .B(n2176), .Z(n2167) );
  XOR2_X1 U2141 ( .A(n2177), .B(n2178), .Z(n2176) );
  AND2_X1 U2142 ( .A1(n2029), .A2(n2030), .ZN(n2031) );
  XNOR2_X1 U2143 ( .A(n2162), .B(n2163), .ZN(n2030) );
  OR2_X1 U2144 ( .A1(n2179), .A2(n2180), .ZN(n2163) );
  AND2_X1 U2145 ( .A1(n2181), .A2(n2182), .ZN(n2180) );
  AND2_X1 U2146 ( .A1(n2183), .A2(n2184), .ZN(n2179) );
  OR2_X1 U2147 ( .A1(n2182), .A2(n2181), .ZN(n2184) );
  XNOR2_X1 U2148 ( .A(n2173), .B(n2185), .ZN(n2162) );
  XOR2_X1 U2149 ( .A(n2172), .B(n2171), .Z(n2185) );
  OR2_X1 U2150 ( .A1(n2186), .A2(n2187), .ZN(n2171) );
  OR2_X1 U2151 ( .A1(n2188), .A2(n2189), .ZN(n2172) );
  AND2_X1 U2152 ( .A1(n2190), .A2(n2191), .ZN(n2189) );
  AND2_X1 U2153 ( .A1(n2192), .A2(n2193), .ZN(n2188) );
  OR2_X1 U2154 ( .A1(n2191), .A2(n2190), .ZN(n2193) );
  XOR2_X1 U2155 ( .A(n2194), .B(n2195), .Z(n2173) );
  XOR2_X1 U2156 ( .A(n2196), .B(n2197), .Z(n2195) );
  OR2_X1 U2157 ( .A1(n2198), .A2(n2199), .ZN(n2029) );
  OR2_X1 U2158 ( .A1(n2200), .A2(n2028), .ZN(n2198) );
  AND2_X1 U2159 ( .A1(n2026), .A2(n2027), .ZN(n2028) );
  AND2_X1 U2160 ( .A1(n2201), .A2(n2202), .ZN(n2027) );
  INV_X1 U2161 ( .A(n2203), .ZN(n2201) );
  AND2_X1 U2162 ( .A1(n2022), .A2(n2026), .ZN(n2200) );
  INV_X1 U2163 ( .A(n2204), .ZN(n2026) );
  OR2_X1 U2164 ( .A1(n2205), .A2(n2199), .ZN(n2204) );
  INV_X1 U2165 ( .A(n2206), .ZN(n2199) );
  OR2_X1 U2166 ( .A1(n2207), .A2(n2208), .ZN(n2206) );
  AND2_X1 U2167 ( .A1(n2207), .A2(n2208), .ZN(n2205) );
  OR2_X1 U2168 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
  AND2_X1 U2169 ( .A1(n2211), .A2(n2212), .ZN(n2210) );
  AND2_X1 U2170 ( .A1(n2213), .A2(n2214), .ZN(n2209) );
  OR2_X1 U2171 ( .A1(n2212), .A2(n2211), .ZN(n2214) );
  XOR2_X1 U2172 ( .A(n2183), .B(n2215), .Z(n2207) );
  XOR2_X1 U2173 ( .A(n2182), .B(n2181), .Z(n2215) );
  OR2_X1 U2174 ( .A1(n2216), .A2(n2187), .ZN(n2181) );
  OR2_X1 U2175 ( .A1(n2217), .A2(n2218), .ZN(n2182) );
  AND2_X1 U2176 ( .A1(n2219), .A2(n2220), .ZN(n2218) );
  AND2_X1 U2177 ( .A1(n2221), .A2(n2222), .ZN(n2217) );
  OR2_X1 U2178 ( .A1(n2220), .A2(n2219), .ZN(n2222) );
  XOR2_X1 U2179 ( .A(n2192), .B(n2223), .Z(n2183) );
  XOR2_X1 U2180 ( .A(n2191), .B(n2190), .Z(n2223) );
  OR2_X1 U2181 ( .A1(n2186), .A2(n2224), .ZN(n2190) );
  OR2_X1 U2182 ( .A1(n2225), .A2(n2226), .ZN(n2191) );
  AND2_X1 U2183 ( .A1(n2227), .A2(n2228), .ZN(n2226) );
  AND2_X1 U2184 ( .A1(n2229), .A2(n2230), .ZN(n2225) );
  OR2_X1 U2185 ( .A1(n2228), .A2(n2227), .ZN(n2230) );
  XOR2_X1 U2186 ( .A(n2231), .B(n2232), .Z(n2192) );
  XOR2_X1 U2187 ( .A(n2233), .B(n2234), .Z(n2232) );
  AND2_X1 U2188 ( .A1(n2020), .A2(n2021), .ZN(n2022) );
  XNOR2_X1 U2189 ( .A(n2202), .B(n2203), .ZN(n2021) );
  OR2_X1 U2190 ( .A1(n2235), .A2(n2236), .ZN(n2203) );
  AND2_X1 U2191 ( .A1(n2237), .A2(n2238), .ZN(n2236) );
  AND2_X1 U2192 ( .A1(n2239), .A2(n2240), .ZN(n2235) );
  OR2_X1 U2193 ( .A1(n2238), .A2(n2237), .ZN(n2240) );
  XNOR2_X1 U2194 ( .A(n2213), .B(n2241), .ZN(n2202) );
  XOR2_X1 U2195 ( .A(n2212), .B(n2211), .Z(n2241) );
  OR2_X1 U2196 ( .A1(n2242), .A2(n2187), .ZN(n2211) );
  OR2_X1 U2197 ( .A1(n2243), .A2(n2244), .ZN(n2212) );
  AND2_X1 U2198 ( .A1(n2245), .A2(n2246), .ZN(n2244) );
  AND2_X1 U2199 ( .A1(n2247), .A2(n2248), .ZN(n2243) );
  OR2_X1 U2200 ( .A1(n2246), .A2(n2245), .ZN(n2248) );
  XOR2_X1 U2201 ( .A(n2221), .B(n2249), .Z(n2213) );
  XOR2_X1 U2202 ( .A(n2220), .B(n2219), .Z(n2249) );
  OR2_X1 U2203 ( .A1(n2216), .A2(n2224), .ZN(n2219) );
  OR2_X1 U2204 ( .A1(n2250), .A2(n2251), .ZN(n2220) );
  AND2_X1 U2205 ( .A1(n2252), .A2(n2253), .ZN(n2251) );
  AND2_X1 U2206 ( .A1(n2254), .A2(n2255), .ZN(n2250) );
  OR2_X1 U2207 ( .A1(n2253), .A2(n2252), .ZN(n2255) );
  XOR2_X1 U2208 ( .A(n2229), .B(n2256), .Z(n2221) );
  XOR2_X1 U2209 ( .A(n2228), .B(n2227), .Z(n2256) );
  OR2_X1 U2210 ( .A1(n2186), .A2(n2257), .ZN(n2227) );
  OR2_X1 U2211 ( .A1(n2258), .A2(n2259), .ZN(n2228) );
  AND2_X1 U2212 ( .A1(n2260), .A2(n2261), .ZN(n2259) );
  AND2_X1 U2213 ( .A1(n2262), .A2(n2263), .ZN(n2258) );
  OR2_X1 U2214 ( .A1(n2261), .A2(n2260), .ZN(n2263) );
  XOR2_X1 U2215 ( .A(n2264), .B(n2265), .Z(n2229) );
  XOR2_X1 U2216 ( .A(n2266), .B(n2267), .Z(n2265) );
  OR2_X1 U2217 ( .A1(n2268), .A2(n2269), .ZN(n2020) );
  OR2_X1 U2218 ( .A1(n2270), .A2(n2019), .ZN(n2268) );
  AND2_X1 U2219 ( .A1(n2017), .A2(n2018), .ZN(n2019) );
  AND2_X1 U2220 ( .A1(n2271), .A2(n2272), .ZN(n2018) );
  INV_X1 U2221 ( .A(n2273), .ZN(n2271) );
  AND2_X1 U2222 ( .A1(n2013), .A2(n2017), .ZN(n2270) );
  INV_X1 U2223 ( .A(n2274), .ZN(n2017) );
  OR2_X1 U2224 ( .A1(n2275), .A2(n2269), .ZN(n2274) );
  INV_X1 U2225 ( .A(n2276), .ZN(n2269) );
  OR2_X1 U2226 ( .A1(n2277), .A2(n2278), .ZN(n2276) );
  AND2_X1 U2227 ( .A1(n2277), .A2(n2278), .ZN(n2275) );
  OR2_X1 U2228 ( .A1(n2279), .A2(n2280), .ZN(n2278) );
  AND2_X1 U2229 ( .A1(n2281), .A2(n2282), .ZN(n2280) );
  AND2_X1 U2230 ( .A1(n2283), .A2(n2284), .ZN(n2279) );
  OR2_X1 U2231 ( .A1(n2282), .A2(n2281), .ZN(n2284) );
  XOR2_X1 U2232 ( .A(n2239), .B(n2285), .Z(n2277) );
  XOR2_X1 U2233 ( .A(n2238), .B(n2237), .Z(n2285) );
  OR2_X1 U2234 ( .A1(n2286), .A2(n2187), .ZN(n2237) );
  OR2_X1 U2235 ( .A1(n2287), .A2(n2288), .ZN(n2238) );
  AND2_X1 U2236 ( .A1(n2289), .A2(n2290), .ZN(n2288) );
  AND2_X1 U2237 ( .A1(n2291), .A2(n2292), .ZN(n2287) );
  OR2_X1 U2238 ( .A1(n2290), .A2(n2289), .ZN(n2292) );
  XOR2_X1 U2239 ( .A(n2247), .B(n2293), .Z(n2239) );
  XOR2_X1 U2240 ( .A(n2246), .B(n2245), .Z(n2293) );
  OR2_X1 U2241 ( .A1(n2242), .A2(n2224), .ZN(n2245) );
  OR2_X1 U2242 ( .A1(n2294), .A2(n2295), .ZN(n2246) );
  AND2_X1 U2243 ( .A1(n2296), .A2(n2297), .ZN(n2295) );
  AND2_X1 U2244 ( .A1(n2298), .A2(n2299), .ZN(n2294) );
  OR2_X1 U2245 ( .A1(n2297), .A2(n2296), .ZN(n2299) );
  XOR2_X1 U2246 ( .A(n2254), .B(n2300), .Z(n2247) );
  XOR2_X1 U2247 ( .A(n2253), .B(n2252), .Z(n2300) );
  OR2_X1 U2248 ( .A1(n2216), .A2(n2257), .ZN(n2252) );
  OR2_X1 U2249 ( .A1(n2301), .A2(n2302), .ZN(n2253) );
  AND2_X1 U2250 ( .A1(n2303), .A2(n2304), .ZN(n2302) );
  AND2_X1 U2251 ( .A1(n2305), .A2(n2306), .ZN(n2301) );
  OR2_X1 U2252 ( .A1(n2304), .A2(n2303), .ZN(n2306) );
  XOR2_X1 U2253 ( .A(n2262), .B(n2307), .Z(n2254) );
  XOR2_X1 U2254 ( .A(n2261), .B(n2260), .Z(n2307) );
  OR2_X1 U2255 ( .A1(n2186), .A2(n2308), .ZN(n2260) );
  OR2_X1 U2256 ( .A1(n2309), .A2(n2310), .ZN(n2261) );
  AND2_X1 U2257 ( .A1(n2311), .A2(n2312), .ZN(n2310) );
  AND2_X1 U2258 ( .A1(n2313), .A2(n2314), .ZN(n2309) );
  OR2_X1 U2259 ( .A1(n2312), .A2(n2311), .ZN(n2314) );
  XOR2_X1 U2260 ( .A(n2315), .B(n2316), .Z(n2262) );
  XOR2_X1 U2261 ( .A(n2317), .B(n2318), .Z(n2316) );
  AND2_X1 U2262 ( .A1(n2011), .A2(n2012), .ZN(n2013) );
  XNOR2_X1 U2263 ( .A(n2272), .B(n2273), .ZN(n2012) );
  OR2_X1 U2264 ( .A1(n2319), .A2(n2320), .ZN(n2273) );
  AND2_X1 U2265 ( .A1(n2321), .A2(n2322), .ZN(n2320) );
  AND2_X1 U2266 ( .A1(n2323), .A2(n2324), .ZN(n2319) );
  OR2_X1 U2267 ( .A1(n2322), .A2(n2321), .ZN(n2324) );
  XNOR2_X1 U2268 ( .A(n2283), .B(n2325), .ZN(n2272) );
  XOR2_X1 U2269 ( .A(n2282), .B(n2281), .Z(n2325) );
  OR2_X1 U2270 ( .A1(n2326), .A2(n2187), .ZN(n2281) );
  OR2_X1 U2271 ( .A1(n2327), .A2(n2328), .ZN(n2282) );
  AND2_X1 U2272 ( .A1(n2329), .A2(n2330), .ZN(n2328) );
  AND2_X1 U2273 ( .A1(n2331), .A2(n2332), .ZN(n2327) );
  OR2_X1 U2274 ( .A1(n2330), .A2(n2329), .ZN(n2332) );
  XOR2_X1 U2275 ( .A(n2291), .B(n2333), .Z(n2283) );
  XOR2_X1 U2276 ( .A(n2290), .B(n2289), .Z(n2333) );
  OR2_X1 U2277 ( .A1(n2286), .A2(n2224), .ZN(n2289) );
  OR2_X1 U2278 ( .A1(n2334), .A2(n2335), .ZN(n2290) );
  AND2_X1 U2279 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  AND2_X1 U2280 ( .A1(n2338), .A2(n2339), .ZN(n2334) );
  OR2_X1 U2281 ( .A1(n2337), .A2(n2336), .ZN(n2339) );
  XOR2_X1 U2282 ( .A(n2298), .B(n2340), .Z(n2291) );
  XOR2_X1 U2283 ( .A(n2297), .B(n2296), .Z(n2340) );
  OR2_X1 U2284 ( .A1(n2242), .A2(n2257), .ZN(n2296) );
  OR2_X1 U2285 ( .A1(n2341), .A2(n2342), .ZN(n2297) );
  AND2_X1 U2286 ( .A1(n2343), .A2(n2344), .ZN(n2342) );
  AND2_X1 U2287 ( .A1(n2345), .A2(n2346), .ZN(n2341) );
  OR2_X1 U2288 ( .A1(n2344), .A2(n2343), .ZN(n2346) );
  XOR2_X1 U2289 ( .A(n2305), .B(n2347), .Z(n2298) );
  XOR2_X1 U2290 ( .A(n2304), .B(n2303), .Z(n2347) );
  OR2_X1 U2291 ( .A1(n2216), .A2(n2308), .ZN(n2303) );
  OR2_X1 U2292 ( .A1(n2348), .A2(n2349), .ZN(n2304) );
  AND2_X1 U2293 ( .A1(n2350), .A2(n2351), .ZN(n2349) );
  AND2_X1 U2294 ( .A1(n2352), .A2(n2353), .ZN(n2348) );
  OR2_X1 U2295 ( .A1(n2351), .A2(n2350), .ZN(n2353) );
  XOR2_X1 U2296 ( .A(n2313), .B(n2354), .Z(n2305) );
  XOR2_X1 U2297 ( .A(n2312), .B(n2311), .Z(n2354) );
  OR2_X1 U2298 ( .A1(n2186), .A2(n2355), .ZN(n2311) );
  OR2_X1 U2299 ( .A1(n2356), .A2(n2357), .ZN(n2312) );
  AND2_X1 U2300 ( .A1(n2358), .A2(n2359), .ZN(n2357) );
  AND2_X1 U2301 ( .A1(n2360), .A2(n2361), .ZN(n2356) );
  OR2_X1 U2302 ( .A1(n2359), .A2(n2358), .ZN(n2361) );
  XOR2_X1 U2303 ( .A(n2362), .B(n2363), .Z(n2313) );
  XOR2_X1 U2304 ( .A(n2364), .B(n2365), .Z(n2363) );
  OR2_X1 U2305 ( .A1(n2366), .A2(n2367), .ZN(n2011) );
  OR2_X1 U2306 ( .A1(n2368), .A2(n2008), .ZN(n2366) );
  AND2_X1 U2307 ( .A1(n2369), .A2(n2370), .ZN(n2008) );
  INV_X1 U2308 ( .A(n2009), .ZN(n2370) );
  OR2_X1 U2309 ( .A1(n2371), .A2(n2372), .ZN(n2009) );
  AND2_X1 U2310 ( .A1(n2369), .A2(n2006), .ZN(n2368) );
  OR2_X1 U2311 ( .A1(n2373), .A2(n2149), .ZN(n2006) );
  INV_X1 U2312 ( .A(n2374), .ZN(n2149) );
  OR2_X1 U2313 ( .A1(n2153), .A2(n2375), .ZN(n2374) );
  OR2_X1 U2314 ( .A1(n2152), .A2(n2150), .ZN(n2375) );
  INV_X1 U2315 ( .A(n2376), .ZN(n2150) );
  AND2_X1 U2316 ( .A1(n2376), .A2(n2147), .ZN(n2373) );
  OR2_X1 U2317 ( .A1(n2377), .A2(n2141), .ZN(n2147) );
  INV_X1 U2318 ( .A(n2378), .ZN(n2141) );
  OR2_X1 U2319 ( .A1(n2145), .A2(n2379), .ZN(n2378) );
  OR2_X1 U2320 ( .A1(n2144), .A2(n2142), .ZN(n2379) );
  INV_X1 U2321 ( .A(n2380), .ZN(n2142) );
  AND2_X1 U2322 ( .A1(n2380), .A2(n2139), .ZN(n2377) );
  OR2_X1 U2323 ( .A1(n2381), .A2(n2133), .ZN(n2139) );
  INV_X1 U2324 ( .A(n2382), .ZN(n2133) );
  OR2_X1 U2325 ( .A1(n2137), .A2(n2383), .ZN(n2382) );
  OR2_X1 U2326 ( .A1(n2136), .A2(n2134), .ZN(n2383) );
  INV_X1 U2327 ( .A(n2384), .ZN(n2134) );
  AND2_X1 U2328 ( .A1(n2384), .A2(n2131), .ZN(n2381) );
  OR2_X1 U2329 ( .A1(n2385), .A2(n2386), .ZN(n2131) );
  AND2_X1 U2330 ( .A1(n2129), .A2(n2128), .ZN(n2386) );
  INV_X1 U2331 ( .A(n2387), .ZN(n2129) );
  OR2_X1 U2332 ( .A1(n2388), .A2(n2389), .ZN(n2387) );
  AND2_X1 U2333 ( .A1(n2123), .A2(n2128), .ZN(n2385) );
  XOR2_X1 U2334 ( .A(n2137), .B(n2136), .Z(n2128) );
  XOR2_X1 U2335 ( .A(n2390), .B(n2391), .Z(n2136) );
  XOR2_X1 U2336 ( .A(n2392), .B(n2393), .Z(n2391) );
  OR2_X1 U2337 ( .A1(n2394), .A2(n2395), .ZN(n2137) );
  AND2_X1 U2338 ( .A1(n2396), .A2(n2397), .ZN(n2395) );
  AND2_X1 U2339 ( .A1(n2398), .A2(n2399), .ZN(n2394) );
  OR2_X1 U2340 ( .A1(n2397), .A2(n2396), .ZN(n2399) );
  AND2_X1 U2341 ( .A1(n2126), .A2(n2400), .ZN(n2123) );
  AND2_X1 U2342 ( .A1(n2120), .A2(n2125), .ZN(n2400) );
  XOR2_X1 U2343 ( .A(n2389), .B(n2388), .Z(n2125) );
  XNOR2_X1 U2344 ( .A(n2401), .B(n2398), .ZN(n2388) );
  XOR2_X1 U2345 ( .A(n2402), .B(n2403), .Z(n2398) );
  XOR2_X1 U2346 ( .A(n2404), .B(n2405), .Z(n2403) );
  XNOR2_X1 U2347 ( .A(n2397), .B(n2396), .ZN(n2401) );
  OR2_X1 U2348 ( .A1(n2406), .A2(n2187), .ZN(n2396) );
  OR2_X1 U2349 ( .A1(n2407), .A2(n2408), .ZN(n2397) );
  AND2_X1 U2350 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  AND2_X1 U2351 ( .A1(n2411), .A2(n2412), .ZN(n2407) );
  OR2_X1 U2352 ( .A1(n2410), .A2(n2409), .ZN(n2412) );
  OR2_X1 U2353 ( .A1(n2413), .A2(n2414), .ZN(n2389) );
  AND2_X1 U2354 ( .A1(n2415), .A2(n2416), .ZN(n2414) );
  AND2_X1 U2355 ( .A1(n2417), .A2(n2418), .ZN(n2413) );
  OR2_X1 U2356 ( .A1(n2415), .A2(n2416), .ZN(n2418) );
  XOR2_X1 U2357 ( .A(n2419), .B(n2417), .Z(n2120) );
  XNOR2_X1 U2358 ( .A(n2420), .B(n2411), .ZN(n2417) );
  XNOR2_X1 U2359 ( .A(n2421), .B(n2422), .ZN(n2411) );
  XNOR2_X1 U2360 ( .A(n2423), .B(n2424), .ZN(n2421) );
  XNOR2_X1 U2361 ( .A(n2410), .B(n2409), .ZN(n2420) );
  OR2_X1 U2362 ( .A1(n2224), .A2(n2406), .ZN(n2409) );
  OR2_X1 U2363 ( .A1(n2425), .A2(n2426), .ZN(n2410) );
  AND2_X1 U2364 ( .A1(n2427), .A2(n2428), .ZN(n2426) );
  AND2_X1 U2365 ( .A1(n2429), .A2(n2430), .ZN(n2425) );
  OR2_X1 U2366 ( .A1(n2428), .A2(n2427), .ZN(n2430) );
  XNOR2_X1 U2367 ( .A(n2416), .B(n2415), .ZN(n2419) );
  OR2_X1 U2368 ( .A1(n2050), .A2(n2187), .ZN(n2415) );
  OR2_X1 U2369 ( .A1(n2431), .A2(n2432), .ZN(n2416) );
  AND2_X1 U2370 ( .A1(n2433), .A2(n2434), .ZN(n2432) );
  AND2_X1 U2371 ( .A1(n2435), .A2(n2436), .ZN(n2431) );
  OR2_X1 U2372 ( .A1(n2434), .A2(n2433), .ZN(n2436) );
  INV_X1 U2373 ( .A(n2119), .ZN(n2126) );
  OR2_X1 U2374 ( .A1(n2437), .A2(n2438), .ZN(n2119) );
  AND2_X1 U2375 ( .A1(n2118), .A2(n2117), .ZN(n2438) );
  AND2_X1 U2376 ( .A1(n2116), .A2(n2439), .ZN(n2437) );
  OR2_X1 U2377 ( .A1(n2118), .A2(n2117), .ZN(n2439) );
  OR2_X1 U2378 ( .A1(n2440), .A2(n2441), .ZN(n2117) );
  AND2_X1 U2379 ( .A1(n2114), .A2(n2113), .ZN(n2441) );
  AND2_X1 U2380 ( .A1(n2112), .A2(n2442), .ZN(n2440) );
  OR2_X1 U2381 ( .A1(n2114), .A2(n2113), .ZN(n2442) );
  OR2_X1 U2382 ( .A1(n2443), .A2(n2444), .ZN(n2113) );
  AND2_X1 U2383 ( .A1(n2110), .A2(n2109), .ZN(n2444) );
  AND2_X1 U2384 ( .A1(n2108), .A2(n2445), .ZN(n2443) );
  OR2_X1 U2385 ( .A1(n2110), .A2(n2109), .ZN(n2445) );
  OR2_X1 U2386 ( .A1(n2446), .A2(n2447), .ZN(n2109) );
  AND2_X1 U2387 ( .A1(n2106), .A2(n2105), .ZN(n2447) );
  AND2_X1 U2388 ( .A1(n2104), .A2(n2448), .ZN(n2446) );
  OR2_X1 U2389 ( .A1(n2106), .A2(n2105), .ZN(n2448) );
  OR2_X1 U2390 ( .A1(n2449), .A2(n2450), .ZN(n2105) );
  AND2_X1 U2391 ( .A1(n2093), .A2(n2092), .ZN(n2450) );
  AND2_X1 U2392 ( .A1(n2091), .A2(n2451), .ZN(n2449) );
  OR2_X1 U2393 ( .A1(n2093), .A2(n2092), .ZN(n2451) );
  OR2_X1 U2394 ( .A1(n2452), .A2(n2453), .ZN(n2092) );
  AND2_X1 U2395 ( .A1(n2089), .A2(n2088), .ZN(n2453) );
  AND2_X1 U2396 ( .A1(n2087), .A2(n2454), .ZN(n2452) );
  OR2_X1 U2397 ( .A1(n2089), .A2(n2088), .ZN(n2454) );
  OR2_X1 U2398 ( .A1(n2455), .A2(n2456), .ZN(n2088) );
  AND2_X1 U2399 ( .A1(n2085), .A2(n2084), .ZN(n2456) );
  AND2_X1 U2400 ( .A1(n2083), .A2(n2457), .ZN(n2455) );
  OR2_X1 U2401 ( .A1(n2085), .A2(n2084), .ZN(n2457) );
  OR2_X1 U2402 ( .A1(n2458), .A2(n2459), .ZN(n2084) );
  AND2_X1 U2403 ( .A1(n2081), .A2(n2080), .ZN(n2459) );
  AND2_X1 U2404 ( .A1(n2079), .A2(n2460), .ZN(n2458) );
  OR2_X1 U2405 ( .A1(n2081), .A2(n2080), .ZN(n2460) );
  OR2_X1 U2406 ( .A1(n2461), .A2(n2462), .ZN(n2080) );
  AND2_X1 U2407 ( .A1(n2077), .A2(n2076), .ZN(n2462) );
  AND2_X1 U2408 ( .A1(n2074), .A2(n2463), .ZN(n2461) );
  OR2_X1 U2409 ( .A1(n2077), .A2(n2076), .ZN(n2463) );
  OR2_X1 U2410 ( .A1(n2464), .A2(n2465), .ZN(n2076) );
  AND2_X1 U2411 ( .A1(n2073), .A2(n2072), .ZN(n2465) );
  AND2_X1 U2412 ( .A1(n2070), .A2(n2466), .ZN(n2464) );
  OR2_X1 U2413 ( .A1(n2073), .A2(n2072), .ZN(n2466) );
  OR2_X1 U2414 ( .A1(n2467), .A2(n2468), .ZN(n2072) );
  AND2_X1 U2415 ( .A1(n2069), .A2(n2068), .ZN(n2468) );
  AND2_X1 U2416 ( .A1(n2066), .A2(n2469), .ZN(n2467) );
  OR2_X1 U2417 ( .A1(n2069), .A2(n2068), .ZN(n2469) );
  OR2_X1 U2418 ( .A1(n2470), .A2(n2471), .ZN(n2068) );
  AND2_X1 U2419 ( .A1(n2065), .A2(n2064), .ZN(n2471) );
  AND2_X1 U2420 ( .A1(n2062), .A2(n2472), .ZN(n2470) );
  OR2_X1 U2421 ( .A1(n2065), .A2(n2064), .ZN(n2472) );
  OR2_X1 U2422 ( .A1(n2473), .A2(n2474), .ZN(n2064) );
  AND2_X1 U2423 ( .A1(n2061), .A2(n2060), .ZN(n2474) );
  AND2_X1 U2424 ( .A1(n2058), .A2(n2475), .ZN(n2473) );
  OR2_X1 U2425 ( .A1(n2061), .A2(n2060), .ZN(n2475) );
  OR2_X1 U2426 ( .A1(n2476), .A2(n2477), .ZN(n2060) );
  AND2_X1 U2427 ( .A1(n2055), .A2(n2057), .ZN(n2477) );
  AND2_X1 U2428 ( .A1(n2478), .A2(n2479), .ZN(n2476) );
  OR2_X1 U2429 ( .A1(n2055), .A2(n2057), .ZN(n2479) );
  OR2_X1 U2430 ( .A1(n2480), .A2(n2046), .ZN(n2057) );
  OR2_X1 U2431 ( .A1(n2481), .A2(n2482), .ZN(n2055) );
  OR2_X1 U2432 ( .A1(n2050), .A2(n2046), .ZN(n2482) );
  INV_X1 U2433 ( .A(n2056), .ZN(n2478) );
  OR2_X1 U2434 ( .A1(n2483), .A2(n2484), .ZN(n2056) );
  AND2_X1 U2435 ( .A1(n2485), .A2(n2486), .ZN(n2484) );
  OR2_X1 U2436 ( .A1(n2487), .A2(n2045), .ZN(n2486) );
  AND2_X1 U2437 ( .A1(n2039), .A2(n2050), .ZN(n2487) );
  AND2_X1 U2438 ( .A1(n2042), .A2(n2488), .ZN(n2483) );
  OR2_X1 U2439 ( .A1(n2489), .A2(n2049), .ZN(n2488) );
  AND2_X1 U2440 ( .A1(n2406), .A2(n2051), .ZN(n2489) );
  INV_X1 U2441 ( .A(n2050), .ZN(n2042) );
  OR2_X1 U2442 ( .A1(n2490), .A2(n2046), .ZN(n2061) );
  XOR2_X1 U2443 ( .A(n2491), .B(n2492), .Z(n2058) );
  XNOR2_X1 U2444 ( .A(n2493), .B(n2494), .ZN(n2491) );
  OR2_X1 U2445 ( .A1(n2495), .A2(n2046), .ZN(n2065) );
  XNOR2_X1 U2446 ( .A(n2496), .B(n2497), .ZN(n2062) );
  XNOR2_X1 U2447 ( .A(n2498), .B(n2499), .ZN(n2496) );
  OR2_X1 U2448 ( .A1(n2500), .A2(n2046), .ZN(n2069) );
  XNOR2_X1 U2449 ( .A(n2501), .B(n2502), .ZN(n2066) );
  XNOR2_X1 U2450 ( .A(n2503), .B(n2504), .ZN(n2501) );
  OR2_X1 U2451 ( .A1(n2505), .A2(n2046), .ZN(n2073) );
  XNOR2_X1 U2452 ( .A(n2506), .B(n2507), .ZN(n2070) );
  XNOR2_X1 U2453 ( .A(n2508), .B(n2509), .ZN(n2506) );
  OR2_X1 U2454 ( .A1(n2510), .A2(n2046), .ZN(n2077) );
  XNOR2_X1 U2455 ( .A(n2511), .B(n2512), .ZN(n2074) );
  XNOR2_X1 U2456 ( .A(n2513), .B(n2514), .ZN(n2511) );
  OR2_X1 U2457 ( .A1(n2515), .A2(n2046), .ZN(n2081) );
  XNOR2_X1 U2458 ( .A(n2516), .B(n2517), .ZN(n2079) );
  XNOR2_X1 U2459 ( .A(n2518), .B(n2519), .ZN(n2516) );
  OR2_X1 U2460 ( .A1(n2520), .A2(n2046), .ZN(n2085) );
  XNOR2_X1 U2461 ( .A(n2521), .B(n2522), .ZN(n2083) );
  XNOR2_X1 U2462 ( .A(n2523), .B(n2524), .ZN(n2521) );
  OR2_X1 U2463 ( .A1(n2525), .A2(n2046), .ZN(n2089) );
  XNOR2_X1 U2464 ( .A(n2526), .B(n2527), .ZN(n2087) );
  XNOR2_X1 U2465 ( .A(n2528), .B(n2529), .ZN(n2526) );
  OR2_X1 U2466 ( .A1(n2355), .A2(n2046), .ZN(n2093) );
  XNOR2_X1 U2467 ( .A(n2530), .B(n2531), .ZN(n2091) );
  XNOR2_X1 U2468 ( .A(n2532), .B(n2533), .ZN(n2530) );
  OR2_X1 U2469 ( .A1(n2308), .A2(n2046), .ZN(n2106) );
  XNOR2_X1 U2470 ( .A(n2534), .B(n2535), .ZN(n2104) );
  XNOR2_X1 U2471 ( .A(n2536), .B(n2537), .ZN(n2534) );
  OR2_X1 U2472 ( .A1(n2257), .A2(n2046), .ZN(n2110) );
  XNOR2_X1 U2473 ( .A(n2538), .B(n2539), .ZN(n2108) );
  XNOR2_X1 U2474 ( .A(n2540), .B(n2541), .ZN(n2538) );
  OR2_X1 U2475 ( .A1(n2224), .A2(n2046), .ZN(n2114) );
  XNOR2_X1 U2476 ( .A(n2542), .B(n2543), .ZN(n2112) );
  XNOR2_X1 U2477 ( .A(n2544), .B(n2545), .ZN(n2542) );
  OR2_X1 U2478 ( .A1(n2046), .A2(n2187), .ZN(n2118) );
  INV_X1 U2479 ( .A(n2038), .ZN(n2046) );
  AND2_X1 U2480 ( .A1(n2546), .A2(n2547), .ZN(n2038) );
  OR2_X1 U2481 ( .A1(c_15_), .A2(d_15_), .ZN(n2546) );
  XNOR2_X1 U2482 ( .A(n2548), .B(n2435), .ZN(n2116) );
  XNOR2_X1 U2483 ( .A(n2549), .B(n2429), .ZN(n2435) );
  XNOR2_X1 U2484 ( .A(n2550), .B(n2551), .ZN(n2429) );
  XNOR2_X1 U2485 ( .A(n2552), .B(n2553), .ZN(n2550) );
  XNOR2_X1 U2486 ( .A(n2428), .B(n2427), .ZN(n2549) );
  OR2_X1 U2487 ( .A1(n2257), .A2(n2406), .ZN(n2427) );
  OR2_X1 U2488 ( .A1(n2554), .A2(n2555), .ZN(n2428) );
  AND2_X1 U2489 ( .A1(n2556), .A2(n2557), .ZN(n2555) );
  AND2_X1 U2490 ( .A1(n2558), .A2(n2559), .ZN(n2554) );
  OR2_X1 U2491 ( .A1(n2557), .A2(n2556), .ZN(n2559) );
  XNOR2_X1 U2492 ( .A(n2434), .B(n2433), .ZN(n2548) );
  OR2_X1 U2493 ( .A1(n2224), .A2(n2050), .ZN(n2433) );
  OR2_X1 U2494 ( .A1(n2560), .A2(n2561), .ZN(n2434) );
  AND2_X1 U2495 ( .A1(n2545), .A2(n2544), .ZN(n2561) );
  AND2_X1 U2496 ( .A1(n2543), .A2(n2562), .ZN(n2560) );
  OR2_X1 U2497 ( .A1(n2544), .A2(n2545), .ZN(n2562) );
  OR2_X1 U2498 ( .A1(n2257), .A2(n2050), .ZN(n2545) );
  OR2_X1 U2499 ( .A1(n2563), .A2(n2564), .ZN(n2544) );
  AND2_X1 U2500 ( .A1(n2541), .A2(n2540), .ZN(n2564) );
  AND2_X1 U2501 ( .A1(n2539), .A2(n2565), .ZN(n2563) );
  OR2_X1 U2502 ( .A1(n2540), .A2(n2541), .ZN(n2565) );
  OR2_X1 U2503 ( .A1(n2308), .A2(n2050), .ZN(n2541) );
  OR2_X1 U2504 ( .A1(n2566), .A2(n2567), .ZN(n2540) );
  AND2_X1 U2505 ( .A1(n2537), .A2(n2536), .ZN(n2567) );
  AND2_X1 U2506 ( .A1(n2535), .A2(n2568), .ZN(n2566) );
  OR2_X1 U2507 ( .A1(n2536), .A2(n2537), .ZN(n2568) );
  OR2_X1 U2508 ( .A1(n2355), .A2(n2050), .ZN(n2537) );
  OR2_X1 U2509 ( .A1(n2569), .A2(n2570), .ZN(n2536) );
  AND2_X1 U2510 ( .A1(n2533), .A2(n2532), .ZN(n2570) );
  AND2_X1 U2511 ( .A1(n2531), .A2(n2571), .ZN(n2569) );
  OR2_X1 U2512 ( .A1(n2532), .A2(n2533), .ZN(n2571) );
  OR2_X1 U2513 ( .A1(n2525), .A2(n2050), .ZN(n2533) );
  OR2_X1 U2514 ( .A1(n2572), .A2(n2573), .ZN(n2532) );
  AND2_X1 U2515 ( .A1(n2529), .A2(n2528), .ZN(n2573) );
  AND2_X1 U2516 ( .A1(n2527), .A2(n2574), .ZN(n2572) );
  OR2_X1 U2517 ( .A1(n2528), .A2(n2529), .ZN(n2574) );
  OR2_X1 U2518 ( .A1(n2520), .A2(n2050), .ZN(n2529) );
  OR2_X1 U2519 ( .A1(n2575), .A2(n2576), .ZN(n2528) );
  AND2_X1 U2520 ( .A1(n2524), .A2(n2523), .ZN(n2576) );
  AND2_X1 U2521 ( .A1(n2522), .A2(n2577), .ZN(n2575) );
  OR2_X1 U2522 ( .A1(n2523), .A2(n2524), .ZN(n2577) );
  OR2_X1 U2523 ( .A1(n2515), .A2(n2050), .ZN(n2524) );
  OR2_X1 U2524 ( .A1(n2578), .A2(n2579), .ZN(n2523) );
  AND2_X1 U2525 ( .A1(n2519), .A2(n2518), .ZN(n2579) );
  AND2_X1 U2526 ( .A1(n2517), .A2(n2580), .ZN(n2578) );
  OR2_X1 U2527 ( .A1(n2518), .A2(n2519), .ZN(n2580) );
  OR2_X1 U2528 ( .A1(n2510), .A2(n2050), .ZN(n2519) );
  OR2_X1 U2529 ( .A1(n2581), .A2(n2582), .ZN(n2518) );
  AND2_X1 U2530 ( .A1(n2514), .A2(n2513), .ZN(n2582) );
  AND2_X1 U2531 ( .A1(n2512), .A2(n2583), .ZN(n2581) );
  OR2_X1 U2532 ( .A1(n2513), .A2(n2514), .ZN(n2583) );
  OR2_X1 U2533 ( .A1(n2505), .A2(n2050), .ZN(n2514) );
  OR2_X1 U2534 ( .A1(n2584), .A2(n2585), .ZN(n2513) );
  AND2_X1 U2535 ( .A1(n2509), .A2(n2508), .ZN(n2585) );
  AND2_X1 U2536 ( .A1(n2507), .A2(n2586), .ZN(n2584) );
  OR2_X1 U2537 ( .A1(n2508), .A2(n2509), .ZN(n2586) );
  OR2_X1 U2538 ( .A1(n2500), .A2(n2050), .ZN(n2509) );
  OR2_X1 U2539 ( .A1(n2587), .A2(n2588), .ZN(n2508) );
  AND2_X1 U2540 ( .A1(n2504), .A2(n2503), .ZN(n2588) );
  AND2_X1 U2541 ( .A1(n2502), .A2(n2589), .ZN(n2587) );
  OR2_X1 U2542 ( .A1(n2503), .A2(n2504), .ZN(n2589) );
  OR2_X1 U2543 ( .A1(n2495), .A2(n2050), .ZN(n2504) );
  OR2_X1 U2544 ( .A1(n2590), .A2(n2591), .ZN(n2503) );
  AND2_X1 U2545 ( .A1(n2499), .A2(n2498), .ZN(n2591) );
  AND2_X1 U2546 ( .A1(n2497), .A2(n2592), .ZN(n2590) );
  OR2_X1 U2547 ( .A1(n2498), .A2(n2499), .ZN(n2592) );
  OR2_X1 U2548 ( .A1(n2490), .A2(n2050), .ZN(n2499) );
  OR2_X1 U2549 ( .A1(n2593), .A2(n2594), .ZN(n2498) );
  AND2_X1 U2550 ( .A1(n2492), .A2(n2494), .ZN(n2594) );
  AND2_X1 U2551 ( .A1(n2595), .A2(n2596), .ZN(n2593) );
  OR2_X1 U2552 ( .A1(n2494), .A2(n2492), .ZN(n2596) );
  OR2_X1 U2553 ( .A1(n2050), .A2(n2480), .ZN(n2492) );
  OR2_X1 U2554 ( .A1(n2481), .A2(n2597), .ZN(n2494) );
  OR2_X1 U2555 ( .A1(n2050), .A2(n2406), .ZN(n2597) );
  XOR2_X1 U2556 ( .A(d_14_), .B(c_14_), .Z(n2598) );
  INV_X1 U2557 ( .A(n2599), .ZN(n2547) );
  INV_X1 U2558 ( .A(n2493), .ZN(n2595) );
  OR2_X1 U2559 ( .A1(n2600), .A2(n2601), .ZN(n2493) );
  AND2_X1 U2560 ( .A1(n2602), .A2(n2603), .ZN(n2601) );
  OR2_X1 U2561 ( .A1(n2604), .A2(n2045), .ZN(n2603) );
  AND2_X1 U2562 ( .A1(n2039), .A2(n2406), .ZN(n2604) );
  AND2_X1 U2563 ( .A1(n2485), .A2(n2605), .ZN(n2600) );
  OR2_X1 U2564 ( .A1(n2606), .A2(n2049), .ZN(n2605) );
  AND2_X1 U2565 ( .A1(n2607), .A2(n2051), .ZN(n2606) );
  INV_X1 U2566 ( .A(n2406), .ZN(n2485) );
  XOR2_X1 U2567 ( .A(n2608), .B(n2609), .Z(n2497) );
  XNOR2_X1 U2568 ( .A(n2610), .B(n2611), .ZN(n2608) );
  XNOR2_X1 U2569 ( .A(n2612), .B(n2613), .ZN(n2502) );
  XNOR2_X1 U2570 ( .A(n2614), .B(n2615), .ZN(n2612) );
  XNOR2_X1 U2571 ( .A(n2616), .B(n2617), .ZN(n2507) );
  XNOR2_X1 U2572 ( .A(n2618), .B(n2619), .ZN(n2616) );
  XNOR2_X1 U2573 ( .A(n2620), .B(n2621), .ZN(n2512) );
  XNOR2_X1 U2574 ( .A(n2622), .B(n2623), .ZN(n2620) );
  XNOR2_X1 U2575 ( .A(n2624), .B(n2625), .ZN(n2517) );
  XNOR2_X1 U2576 ( .A(n2626), .B(n2627), .ZN(n2624) );
  XNOR2_X1 U2577 ( .A(n2628), .B(n2629), .ZN(n2522) );
  XNOR2_X1 U2578 ( .A(n2630), .B(n2631), .ZN(n2628) );
  XNOR2_X1 U2579 ( .A(n2632), .B(n2633), .ZN(n2527) );
  XNOR2_X1 U2580 ( .A(n2634), .B(n2635), .ZN(n2632) );
  XNOR2_X1 U2581 ( .A(n2636), .B(n2637), .ZN(n2531) );
  XNOR2_X1 U2582 ( .A(n2638), .B(n2639), .ZN(n2636) );
  XNOR2_X1 U2583 ( .A(n2640), .B(n2641), .ZN(n2535) );
  XNOR2_X1 U2584 ( .A(n2642), .B(n2643), .ZN(n2640) );
  XNOR2_X1 U2585 ( .A(n2644), .B(n2645), .ZN(n2539) );
  XNOR2_X1 U2586 ( .A(n2646), .B(n2647), .ZN(n2644) );
  XNOR2_X1 U2587 ( .A(n2648), .B(n2558), .ZN(n2543) );
  XNOR2_X1 U2588 ( .A(n2649), .B(n2650), .ZN(n2558) );
  XNOR2_X1 U2589 ( .A(n2651), .B(n2652), .ZN(n2649) );
  XNOR2_X1 U2590 ( .A(n2557), .B(n2556), .ZN(n2648) );
  OR2_X1 U2591 ( .A1(n2308), .A2(n2406), .ZN(n2556) );
  OR2_X1 U2592 ( .A1(n2653), .A2(n2654), .ZN(n2557) );
  AND2_X1 U2593 ( .A1(n2647), .A2(n2646), .ZN(n2654) );
  AND2_X1 U2594 ( .A1(n2645), .A2(n2655), .ZN(n2653) );
  OR2_X1 U2595 ( .A1(n2646), .A2(n2647), .ZN(n2655) );
  OR2_X1 U2596 ( .A1(n2355), .A2(n2406), .ZN(n2647) );
  OR2_X1 U2597 ( .A1(n2656), .A2(n2657), .ZN(n2646) );
  AND2_X1 U2598 ( .A1(n2643), .A2(n2642), .ZN(n2657) );
  AND2_X1 U2599 ( .A1(n2641), .A2(n2658), .ZN(n2656) );
  OR2_X1 U2600 ( .A1(n2642), .A2(n2643), .ZN(n2658) );
  OR2_X1 U2601 ( .A1(n2525), .A2(n2406), .ZN(n2643) );
  OR2_X1 U2602 ( .A1(n2659), .A2(n2660), .ZN(n2642) );
  AND2_X1 U2603 ( .A1(n2639), .A2(n2638), .ZN(n2660) );
  AND2_X1 U2604 ( .A1(n2637), .A2(n2661), .ZN(n2659) );
  OR2_X1 U2605 ( .A1(n2638), .A2(n2639), .ZN(n2661) );
  OR2_X1 U2606 ( .A1(n2520), .A2(n2406), .ZN(n2639) );
  OR2_X1 U2607 ( .A1(n2662), .A2(n2663), .ZN(n2638) );
  AND2_X1 U2608 ( .A1(n2635), .A2(n2634), .ZN(n2663) );
  AND2_X1 U2609 ( .A1(n2633), .A2(n2664), .ZN(n2662) );
  OR2_X1 U2610 ( .A1(n2634), .A2(n2635), .ZN(n2664) );
  OR2_X1 U2611 ( .A1(n2515), .A2(n2406), .ZN(n2635) );
  OR2_X1 U2612 ( .A1(n2665), .A2(n2666), .ZN(n2634) );
  AND2_X1 U2613 ( .A1(n2631), .A2(n2630), .ZN(n2666) );
  AND2_X1 U2614 ( .A1(n2629), .A2(n2667), .ZN(n2665) );
  OR2_X1 U2615 ( .A1(n2630), .A2(n2631), .ZN(n2667) );
  OR2_X1 U2616 ( .A1(n2510), .A2(n2406), .ZN(n2631) );
  OR2_X1 U2617 ( .A1(n2668), .A2(n2669), .ZN(n2630) );
  AND2_X1 U2618 ( .A1(n2627), .A2(n2626), .ZN(n2669) );
  AND2_X1 U2619 ( .A1(n2625), .A2(n2670), .ZN(n2668) );
  OR2_X1 U2620 ( .A1(n2626), .A2(n2627), .ZN(n2670) );
  OR2_X1 U2621 ( .A1(n2505), .A2(n2406), .ZN(n2627) );
  OR2_X1 U2622 ( .A1(n2671), .A2(n2672), .ZN(n2626) );
  AND2_X1 U2623 ( .A1(n2623), .A2(n2622), .ZN(n2672) );
  AND2_X1 U2624 ( .A1(n2621), .A2(n2673), .ZN(n2671) );
  OR2_X1 U2625 ( .A1(n2622), .A2(n2623), .ZN(n2673) );
  OR2_X1 U2626 ( .A1(n2500), .A2(n2406), .ZN(n2623) );
  OR2_X1 U2627 ( .A1(n2674), .A2(n2675), .ZN(n2622) );
  AND2_X1 U2628 ( .A1(n2619), .A2(n2618), .ZN(n2675) );
  AND2_X1 U2629 ( .A1(n2617), .A2(n2676), .ZN(n2674) );
  OR2_X1 U2630 ( .A1(n2618), .A2(n2619), .ZN(n2676) );
  OR2_X1 U2631 ( .A1(n2495), .A2(n2406), .ZN(n2619) );
  OR2_X1 U2632 ( .A1(n2677), .A2(n2678), .ZN(n2618) );
  AND2_X1 U2633 ( .A1(n2615), .A2(n2614), .ZN(n2678) );
  AND2_X1 U2634 ( .A1(n2613), .A2(n2679), .ZN(n2677) );
  OR2_X1 U2635 ( .A1(n2614), .A2(n2615), .ZN(n2679) );
  OR2_X1 U2636 ( .A1(n2490), .A2(n2406), .ZN(n2615) );
  OR2_X1 U2637 ( .A1(n2680), .A2(n2681), .ZN(n2614) );
  AND2_X1 U2638 ( .A1(n2609), .A2(n2611), .ZN(n2681) );
  AND2_X1 U2639 ( .A1(n2682), .A2(n2683), .ZN(n2680) );
  OR2_X1 U2640 ( .A1(n2611), .A2(n2609), .ZN(n2683) );
  OR2_X1 U2641 ( .A1(n2481), .A2(n2684), .ZN(n2611) );
  OR2_X1 U2642 ( .A1(n2607), .A2(n2406), .ZN(n2684) );
  XNOR2_X1 U2643 ( .A(n2687), .B(c_13_), .ZN(n2686) );
  INV_X1 U2644 ( .A(n2610), .ZN(n2682) );
  OR2_X1 U2645 ( .A1(n2688), .A2(n2689), .ZN(n2610) );
  AND2_X1 U2646 ( .A1(n2690), .A2(n2691), .ZN(n2689) );
  OR2_X1 U2647 ( .A1(n2692), .A2(n2045), .ZN(n2691) );
  AND2_X1 U2648 ( .A1(n2607), .A2(n2039), .ZN(n2692) );
  AND2_X1 U2649 ( .A1(n2602), .A2(n2693), .ZN(n2688) );
  OR2_X1 U2650 ( .A1(n2694), .A2(n2049), .ZN(n2693) );
  AND2_X1 U2651 ( .A1(n2695), .A2(n2051), .ZN(n2694) );
  XOR2_X1 U2652 ( .A(n2696), .B(n2697), .Z(n2613) );
  XNOR2_X1 U2653 ( .A(n2698), .B(n2699), .ZN(n2696) );
  XNOR2_X1 U2654 ( .A(n2700), .B(n2701), .ZN(n2617) );
  XNOR2_X1 U2655 ( .A(n2702), .B(n2703), .ZN(n2700) );
  XNOR2_X1 U2656 ( .A(n2704), .B(n2705), .ZN(n2621) );
  XNOR2_X1 U2657 ( .A(n2706), .B(n2707), .ZN(n2704) );
  XNOR2_X1 U2658 ( .A(n2708), .B(n2709), .ZN(n2625) );
  XNOR2_X1 U2659 ( .A(n2710), .B(n2711), .ZN(n2708) );
  XNOR2_X1 U2660 ( .A(n2712), .B(n2713), .ZN(n2629) );
  XNOR2_X1 U2661 ( .A(n2714), .B(n2715), .ZN(n2712) );
  XNOR2_X1 U2662 ( .A(n2716), .B(n2717), .ZN(n2633) );
  XNOR2_X1 U2663 ( .A(n2718), .B(n2719), .ZN(n2716) );
  XNOR2_X1 U2664 ( .A(n2720), .B(n2721), .ZN(n2637) );
  XNOR2_X1 U2665 ( .A(n2722), .B(n2723), .ZN(n2720) );
  XNOR2_X1 U2666 ( .A(n2724), .B(n2725), .ZN(n2641) );
  XNOR2_X1 U2667 ( .A(n2726), .B(n2727), .ZN(n2724) );
  XNOR2_X1 U2668 ( .A(n2728), .B(n2729), .ZN(n2645) );
  XNOR2_X1 U2669 ( .A(n2730), .B(n2731), .ZN(n2728) );
  XOR2_X1 U2670 ( .A(n2144), .B(n2145), .Z(n2384) );
  OR2_X1 U2671 ( .A1(n2732), .A2(n2733), .ZN(n2145) );
  AND2_X1 U2672 ( .A1(n2393), .A2(n2392), .ZN(n2733) );
  AND2_X1 U2673 ( .A1(n2390), .A2(n2734), .ZN(n2732) );
  OR2_X1 U2674 ( .A1(n2392), .A2(n2393), .ZN(n2734) );
  OR2_X1 U2675 ( .A1(n2607), .A2(n2187), .ZN(n2393) );
  OR2_X1 U2676 ( .A1(n2735), .A2(n2736), .ZN(n2392) );
  AND2_X1 U2677 ( .A1(n2405), .A2(n2404), .ZN(n2736) );
  AND2_X1 U2678 ( .A1(n2402), .A2(n2737), .ZN(n2735) );
  OR2_X1 U2679 ( .A1(n2404), .A2(n2405), .ZN(n2737) );
  OR2_X1 U2680 ( .A1(n2607), .A2(n2224), .ZN(n2405) );
  OR2_X1 U2681 ( .A1(n2738), .A2(n2739), .ZN(n2404) );
  AND2_X1 U2682 ( .A1(n2424), .A2(n2423), .ZN(n2739) );
  AND2_X1 U2683 ( .A1(n2422), .A2(n2740), .ZN(n2738) );
  OR2_X1 U2684 ( .A1(n2423), .A2(n2424), .ZN(n2740) );
  OR2_X1 U2685 ( .A1(n2607), .A2(n2257), .ZN(n2424) );
  OR2_X1 U2686 ( .A1(n2741), .A2(n2742), .ZN(n2423) );
  AND2_X1 U2687 ( .A1(n2553), .A2(n2552), .ZN(n2742) );
  AND2_X1 U2688 ( .A1(n2551), .A2(n2743), .ZN(n2741) );
  OR2_X1 U2689 ( .A1(n2552), .A2(n2553), .ZN(n2743) );
  OR2_X1 U2690 ( .A1(n2308), .A2(n2607), .ZN(n2553) );
  OR2_X1 U2691 ( .A1(n2744), .A2(n2745), .ZN(n2552) );
  AND2_X1 U2692 ( .A1(n2652), .A2(n2651), .ZN(n2745) );
  AND2_X1 U2693 ( .A1(n2650), .A2(n2746), .ZN(n2744) );
  OR2_X1 U2694 ( .A1(n2651), .A2(n2652), .ZN(n2746) );
  OR2_X1 U2695 ( .A1(n2355), .A2(n2607), .ZN(n2652) );
  OR2_X1 U2696 ( .A1(n2747), .A2(n2748), .ZN(n2651) );
  AND2_X1 U2697 ( .A1(n2731), .A2(n2730), .ZN(n2748) );
  AND2_X1 U2698 ( .A1(n2729), .A2(n2749), .ZN(n2747) );
  OR2_X1 U2699 ( .A1(n2730), .A2(n2731), .ZN(n2749) );
  OR2_X1 U2700 ( .A1(n2525), .A2(n2607), .ZN(n2731) );
  OR2_X1 U2701 ( .A1(n2750), .A2(n2751), .ZN(n2730) );
  AND2_X1 U2702 ( .A1(n2727), .A2(n2726), .ZN(n2751) );
  AND2_X1 U2703 ( .A1(n2725), .A2(n2752), .ZN(n2750) );
  OR2_X1 U2704 ( .A1(n2726), .A2(n2727), .ZN(n2752) );
  OR2_X1 U2705 ( .A1(n2520), .A2(n2607), .ZN(n2727) );
  OR2_X1 U2706 ( .A1(n2753), .A2(n2754), .ZN(n2726) );
  AND2_X1 U2707 ( .A1(n2723), .A2(n2722), .ZN(n2754) );
  AND2_X1 U2708 ( .A1(n2721), .A2(n2755), .ZN(n2753) );
  OR2_X1 U2709 ( .A1(n2722), .A2(n2723), .ZN(n2755) );
  OR2_X1 U2710 ( .A1(n2515), .A2(n2607), .ZN(n2723) );
  OR2_X1 U2711 ( .A1(n2756), .A2(n2757), .ZN(n2722) );
  AND2_X1 U2712 ( .A1(n2719), .A2(n2718), .ZN(n2757) );
  AND2_X1 U2713 ( .A1(n2717), .A2(n2758), .ZN(n2756) );
  OR2_X1 U2714 ( .A1(n2718), .A2(n2719), .ZN(n2758) );
  OR2_X1 U2715 ( .A1(n2510), .A2(n2607), .ZN(n2719) );
  OR2_X1 U2716 ( .A1(n2759), .A2(n2760), .ZN(n2718) );
  AND2_X1 U2717 ( .A1(n2715), .A2(n2714), .ZN(n2760) );
  AND2_X1 U2718 ( .A1(n2713), .A2(n2761), .ZN(n2759) );
  OR2_X1 U2719 ( .A1(n2714), .A2(n2715), .ZN(n2761) );
  OR2_X1 U2720 ( .A1(n2505), .A2(n2607), .ZN(n2715) );
  OR2_X1 U2721 ( .A1(n2762), .A2(n2763), .ZN(n2714) );
  AND2_X1 U2722 ( .A1(n2711), .A2(n2710), .ZN(n2763) );
  AND2_X1 U2723 ( .A1(n2709), .A2(n2764), .ZN(n2762) );
  OR2_X1 U2724 ( .A1(n2710), .A2(n2711), .ZN(n2764) );
  OR2_X1 U2725 ( .A1(n2500), .A2(n2607), .ZN(n2711) );
  OR2_X1 U2726 ( .A1(n2765), .A2(n2766), .ZN(n2710) );
  AND2_X1 U2727 ( .A1(n2707), .A2(n2706), .ZN(n2766) );
  AND2_X1 U2728 ( .A1(n2705), .A2(n2767), .ZN(n2765) );
  OR2_X1 U2729 ( .A1(n2706), .A2(n2707), .ZN(n2767) );
  OR2_X1 U2730 ( .A1(n2495), .A2(n2607), .ZN(n2707) );
  OR2_X1 U2731 ( .A1(n2768), .A2(n2769), .ZN(n2706) );
  AND2_X1 U2732 ( .A1(n2703), .A2(n2702), .ZN(n2769) );
  AND2_X1 U2733 ( .A1(n2701), .A2(n2770), .ZN(n2768) );
  OR2_X1 U2734 ( .A1(n2702), .A2(n2703), .ZN(n2770) );
  OR2_X1 U2735 ( .A1(n2490), .A2(n2607), .ZN(n2703) );
  OR2_X1 U2736 ( .A1(n2771), .A2(n2772), .ZN(n2702) );
  AND2_X1 U2737 ( .A1(n2697), .A2(n2699), .ZN(n2772) );
  AND2_X1 U2738 ( .A1(n2773), .A2(n2774), .ZN(n2771) );
  OR2_X1 U2739 ( .A1(n2699), .A2(n2697), .ZN(n2774) );
  OR2_X1 U2740 ( .A1(n2607), .A2(n2480), .ZN(n2697) );
  OR2_X1 U2741 ( .A1(n2481), .A2(n2775), .ZN(n2699) );
  OR2_X1 U2742 ( .A1(n2695), .A2(n2607), .ZN(n2775) );
  INV_X1 U2743 ( .A(n2602), .ZN(n2607) );
  XOR2_X1 U2744 ( .A(n2776), .B(n2777), .Z(n2602) );
  XNOR2_X1 U2745 ( .A(c_12_), .B(d_12_), .ZN(n2776) );
  INV_X1 U2746 ( .A(n2698), .ZN(n2773) );
  OR2_X1 U2747 ( .A1(n2778), .A2(n2779), .ZN(n2698) );
  AND2_X1 U2748 ( .A1(n2780), .A2(n2781), .ZN(n2779) );
  OR2_X1 U2749 ( .A1(n2782), .A2(n2045), .ZN(n2781) );
  AND2_X1 U2750 ( .A1(n2695), .A2(n2039), .ZN(n2782) );
  AND2_X1 U2751 ( .A1(n2690), .A2(n2783), .ZN(n2778) );
  OR2_X1 U2752 ( .A1(n2784), .A2(n2049), .ZN(n2783) );
  AND2_X1 U2753 ( .A1(n2785), .A2(n2051), .ZN(n2784) );
  XOR2_X1 U2754 ( .A(n2786), .B(n2787), .Z(n2701) );
  XNOR2_X1 U2755 ( .A(n2788), .B(n2789), .ZN(n2786) );
  XNOR2_X1 U2756 ( .A(n2790), .B(n2791), .ZN(n2705) );
  XNOR2_X1 U2757 ( .A(n2792), .B(n2793), .ZN(n2790) );
  XNOR2_X1 U2758 ( .A(n2794), .B(n2795), .ZN(n2709) );
  XNOR2_X1 U2759 ( .A(n2796), .B(n2797), .ZN(n2794) );
  XNOR2_X1 U2760 ( .A(n2798), .B(n2799), .ZN(n2713) );
  XNOR2_X1 U2761 ( .A(n2800), .B(n2801), .ZN(n2798) );
  XNOR2_X1 U2762 ( .A(n2802), .B(n2803), .ZN(n2717) );
  XNOR2_X1 U2763 ( .A(n2804), .B(n2805), .ZN(n2802) );
  XNOR2_X1 U2764 ( .A(n2806), .B(n2807), .ZN(n2721) );
  XNOR2_X1 U2765 ( .A(n2808), .B(n2809), .ZN(n2806) );
  XNOR2_X1 U2766 ( .A(n2810), .B(n2811), .ZN(n2725) );
  XNOR2_X1 U2767 ( .A(n2812), .B(n2813), .ZN(n2810) );
  XNOR2_X1 U2768 ( .A(n2814), .B(n2815), .ZN(n2729) );
  XNOR2_X1 U2769 ( .A(n2816), .B(n2817), .ZN(n2814) );
  XNOR2_X1 U2770 ( .A(n2818), .B(n2819), .ZN(n2650) );
  XNOR2_X1 U2771 ( .A(n2820), .B(n2821), .ZN(n2818) );
  XNOR2_X1 U2772 ( .A(n2822), .B(n2823), .ZN(n2551) );
  XNOR2_X1 U2773 ( .A(n2824), .B(n2825), .ZN(n2822) );
  XOR2_X1 U2774 ( .A(n2826), .B(n2827), .Z(n2422) );
  XOR2_X1 U2775 ( .A(n2828), .B(n2829), .Z(n2827) );
  XOR2_X1 U2776 ( .A(n2830), .B(n2831), .Z(n2402) );
  XOR2_X1 U2777 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR2_X1 U2778 ( .A(n2834), .B(n2835), .Z(n2390) );
  XOR2_X1 U2779 ( .A(n2836), .B(n2837), .Z(n2835) );
  XOR2_X1 U2780 ( .A(n2838), .B(n2839), .Z(n2144) );
  XOR2_X1 U2781 ( .A(n2840), .B(n2841), .Z(n2839) );
  XOR2_X1 U2782 ( .A(n2152), .B(n2153), .Z(n2380) );
  OR2_X1 U2783 ( .A1(n2842), .A2(n2843), .ZN(n2153) );
  AND2_X1 U2784 ( .A1(n2841), .A2(n2840), .ZN(n2843) );
  AND2_X1 U2785 ( .A1(n2838), .A2(n2844), .ZN(n2842) );
  OR2_X1 U2786 ( .A1(n2840), .A2(n2841), .ZN(n2844) );
  OR2_X1 U2787 ( .A1(n2695), .A2(n2187), .ZN(n2841) );
  OR2_X1 U2788 ( .A1(n2845), .A2(n2846), .ZN(n2840) );
  AND2_X1 U2789 ( .A1(n2837), .A2(n2836), .ZN(n2846) );
  AND2_X1 U2790 ( .A1(n2834), .A2(n2847), .ZN(n2845) );
  OR2_X1 U2791 ( .A1(n2836), .A2(n2837), .ZN(n2847) );
  OR2_X1 U2792 ( .A1(n2695), .A2(n2224), .ZN(n2837) );
  OR2_X1 U2793 ( .A1(n2848), .A2(n2849), .ZN(n2836) );
  AND2_X1 U2794 ( .A1(n2833), .A2(n2832), .ZN(n2849) );
  AND2_X1 U2795 ( .A1(n2830), .A2(n2850), .ZN(n2848) );
  OR2_X1 U2796 ( .A1(n2832), .A2(n2833), .ZN(n2850) );
  OR2_X1 U2797 ( .A1(n2695), .A2(n2257), .ZN(n2833) );
  OR2_X1 U2798 ( .A1(n2851), .A2(n2852), .ZN(n2832) );
  AND2_X1 U2799 ( .A1(n2829), .A2(n2828), .ZN(n2852) );
  AND2_X1 U2800 ( .A1(n2826), .A2(n2853), .ZN(n2851) );
  OR2_X1 U2801 ( .A1(n2828), .A2(n2829), .ZN(n2853) );
  OR2_X1 U2802 ( .A1(n2695), .A2(n2308), .ZN(n2829) );
  OR2_X1 U2803 ( .A1(n2854), .A2(n2855), .ZN(n2828) );
  AND2_X1 U2804 ( .A1(n2825), .A2(n2824), .ZN(n2855) );
  AND2_X1 U2805 ( .A1(n2823), .A2(n2856), .ZN(n2854) );
  OR2_X1 U2806 ( .A1(n2824), .A2(n2825), .ZN(n2856) );
  OR2_X1 U2807 ( .A1(n2355), .A2(n2695), .ZN(n2825) );
  OR2_X1 U2808 ( .A1(n2857), .A2(n2858), .ZN(n2824) );
  AND2_X1 U2809 ( .A1(n2821), .A2(n2820), .ZN(n2858) );
  AND2_X1 U2810 ( .A1(n2819), .A2(n2859), .ZN(n2857) );
  OR2_X1 U2811 ( .A1(n2820), .A2(n2821), .ZN(n2859) );
  OR2_X1 U2812 ( .A1(n2525), .A2(n2695), .ZN(n2821) );
  OR2_X1 U2813 ( .A1(n2860), .A2(n2861), .ZN(n2820) );
  AND2_X1 U2814 ( .A1(n2817), .A2(n2816), .ZN(n2861) );
  AND2_X1 U2815 ( .A1(n2815), .A2(n2862), .ZN(n2860) );
  OR2_X1 U2816 ( .A1(n2816), .A2(n2817), .ZN(n2862) );
  OR2_X1 U2817 ( .A1(n2520), .A2(n2695), .ZN(n2817) );
  OR2_X1 U2818 ( .A1(n2863), .A2(n2864), .ZN(n2816) );
  AND2_X1 U2819 ( .A1(n2813), .A2(n2812), .ZN(n2864) );
  AND2_X1 U2820 ( .A1(n2811), .A2(n2865), .ZN(n2863) );
  OR2_X1 U2821 ( .A1(n2812), .A2(n2813), .ZN(n2865) );
  OR2_X1 U2822 ( .A1(n2515), .A2(n2695), .ZN(n2813) );
  OR2_X1 U2823 ( .A1(n2866), .A2(n2867), .ZN(n2812) );
  AND2_X1 U2824 ( .A1(n2809), .A2(n2808), .ZN(n2867) );
  AND2_X1 U2825 ( .A1(n2807), .A2(n2868), .ZN(n2866) );
  OR2_X1 U2826 ( .A1(n2808), .A2(n2809), .ZN(n2868) );
  OR2_X1 U2827 ( .A1(n2510), .A2(n2695), .ZN(n2809) );
  OR2_X1 U2828 ( .A1(n2869), .A2(n2870), .ZN(n2808) );
  AND2_X1 U2829 ( .A1(n2805), .A2(n2804), .ZN(n2870) );
  AND2_X1 U2830 ( .A1(n2803), .A2(n2871), .ZN(n2869) );
  OR2_X1 U2831 ( .A1(n2804), .A2(n2805), .ZN(n2871) );
  OR2_X1 U2832 ( .A1(n2505), .A2(n2695), .ZN(n2805) );
  OR2_X1 U2833 ( .A1(n2872), .A2(n2873), .ZN(n2804) );
  AND2_X1 U2834 ( .A1(n2801), .A2(n2800), .ZN(n2873) );
  AND2_X1 U2835 ( .A1(n2799), .A2(n2874), .ZN(n2872) );
  OR2_X1 U2836 ( .A1(n2800), .A2(n2801), .ZN(n2874) );
  OR2_X1 U2837 ( .A1(n2500), .A2(n2695), .ZN(n2801) );
  OR2_X1 U2838 ( .A1(n2875), .A2(n2876), .ZN(n2800) );
  AND2_X1 U2839 ( .A1(n2797), .A2(n2796), .ZN(n2876) );
  AND2_X1 U2840 ( .A1(n2795), .A2(n2877), .ZN(n2875) );
  OR2_X1 U2841 ( .A1(n2796), .A2(n2797), .ZN(n2877) );
  OR2_X1 U2842 ( .A1(n2495), .A2(n2695), .ZN(n2797) );
  OR2_X1 U2843 ( .A1(n2878), .A2(n2879), .ZN(n2796) );
  AND2_X1 U2844 ( .A1(n2793), .A2(n2792), .ZN(n2879) );
  AND2_X1 U2845 ( .A1(n2791), .A2(n2880), .ZN(n2878) );
  OR2_X1 U2846 ( .A1(n2792), .A2(n2793), .ZN(n2880) );
  OR2_X1 U2847 ( .A1(n2490), .A2(n2695), .ZN(n2793) );
  OR2_X1 U2848 ( .A1(n2881), .A2(n2882), .ZN(n2792) );
  AND2_X1 U2849 ( .A1(n2787), .A2(n2789), .ZN(n2882) );
  AND2_X1 U2850 ( .A1(n2883), .A2(n2884), .ZN(n2881) );
  OR2_X1 U2851 ( .A1(n2789), .A2(n2787), .ZN(n2884) );
  OR2_X1 U2852 ( .A1(n2695), .A2(n2480), .ZN(n2787) );
  OR2_X1 U2853 ( .A1(n2481), .A2(n2885), .ZN(n2789) );
  OR2_X1 U2854 ( .A1(n2785), .A2(n2695), .ZN(n2885) );
  INV_X1 U2855 ( .A(n2690), .ZN(n2695) );
  XOR2_X1 U2856 ( .A(n2886), .B(n2887), .Z(n2690) );
  XNOR2_X1 U2857 ( .A(c_11_), .B(d_11_), .ZN(n2886) );
  INV_X1 U2858 ( .A(n2788), .ZN(n2883) );
  OR2_X1 U2859 ( .A1(n2888), .A2(n2889), .ZN(n2788) );
  AND2_X1 U2860 ( .A1(n2890), .A2(n2891), .ZN(n2889) );
  OR2_X1 U2861 ( .A1(n2892), .A2(n2045), .ZN(n2891) );
  AND2_X1 U2862 ( .A1(n2785), .A2(n2039), .ZN(n2892) );
  AND2_X1 U2863 ( .A1(n2780), .A2(n2893), .ZN(n2888) );
  OR2_X1 U2864 ( .A1(n2894), .A2(n2049), .ZN(n2893) );
  AND2_X1 U2865 ( .A1(n2895), .A2(n2051), .ZN(n2894) );
  XOR2_X1 U2866 ( .A(n2896), .B(n2897), .Z(n2791) );
  XNOR2_X1 U2867 ( .A(n2898), .B(n2899), .ZN(n2896) );
  XNOR2_X1 U2868 ( .A(n2900), .B(n2901), .ZN(n2795) );
  XNOR2_X1 U2869 ( .A(n2902), .B(n2903), .ZN(n2900) );
  XNOR2_X1 U2870 ( .A(n2904), .B(n2905), .ZN(n2799) );
  XNOR2_X1 U2871 ( .A(n2906), .B(n2907), .ZN(n2904) );
  XNOR2_X1 U2872 ( .A(n2908), .B(n2909), .ZN(n2803) );
  XNOR2_X1 U2873 ( .A(n2910), .B(n2911), .ZN(n2908) );
  XNOR2_X1 U2874 ( .A(n2912), .B(n2913), .ZN(n2807) );
  XNOR2_X1 U2875 ( .A(n2914), .B(n2915), .ZN(n2912) );
  XNOR2_X1 U2876 ( .A(n2916), .B(n2917), .ZN(n2811) );
  XNOR2_X1 U2877 ( .A(n2918), .B(n2919), .ZN(n2916) );
  XNOR2_X1 U2878 ( .A(n2920), .B(n2921), .ZN(n2815) );
  XNOR2_X1 U2879 ( .A(n2922), .B(n2923), .ZN(n2920) );
  XNOR2_X1 U2880 ( .A(n2924), .B(n2925), .ZN(n2819) );
  XNOR2_X1 U2881 ( .A(n2926), .B(n2927), .ZN(n2924) );
  XNOR2_X1 U2882 ( .A(n2928), .B(n2929), .ZN(n2823) );
  XNOR2_X1 U2883 ( .A(n2930), .B(n2931), .ZN(n2928) );
  XOR2_X1 U2884 ( .A(n2932), .B(n2933), .Z(n2826) );
  XOR2_X1 U2885 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR2_X1 U2886 ( .A(n2936), .B(n2937), .Z(n2830) );
  XOR2_X1 U2887 ( .A(n2938), .B(n2939), .Z(n2937) );
  XOR2_X1 U2888 ( .A(n2940), .B(n2941), .Z(n2834) );
  XOR2_X1 U2889 ( .A(n2942), .B(n2943), .Z(n2941) );
  XOR2_X1 U2890 ( .A(n2944), .B(n2945), .Z(n2838) );
  XOR2_X1 U2891 ( .A(n2946), .B(n2947), .Z(n2945) );
  XOR2_X1 U2892 ( .A(n2948), .B(n2949), .Z(n2152) );
  XOR2_X1 U2893 ( .A(n2950), .B(n2951), .Z(n2949) );
  XOR2_X1 U2894 ( .A(n2371), .B(n2372), .Z(n2376) );
  OR2_X1 U2895 ( .A1(n2952), .A2(n2953), .ZN(n2372) );
  AND2_X1 U2896 ( .A1(n2951), .A2(n2950), .ZN(n2953) );
  AND2_X1 U2897 ( .A1(n2948), .A2(n2954), .ZN(n2952) );
  OR2_X1 U2898 ( .A1(n2950), .A2(n2951), .ZN(n2954) );
  OR2_X1 U2899 ( .A1(n2785), .A2(n2187), .ZN(n2951) );
  OR2_X1 U2900 ( .A1(n2955), .A2(n2956), .ZN(n2950) );
  AND2_X1 U2901 ( .A1(n2947), .A2(n2946), .ZN(n2956) );
  AND2_X1 U2902 ( .A1(n2944), .A2(n2957), .ZN(n2955) );
  OR2_X1 U2903 ( .A1(n2946), .A2(n2947), .ZN(n2957) );
  OR2_X1 U2904 ( .A1(n2785), .A2(n2224), .ZN(n2947) );
  OR2_X1 U2905 ( .A1(n2958), .A2(n2959), .ZN(n2946) );
  AND2_X1 U2906 ( .A1(n2943), .A2(n2942), .ZN(n2959) );
  AND2_X1 U2907 ( .A1(n2940), .A2(n2960), .ZN(n2958) );
  OR2_X1 U2908 ( .A1(n2942), .A2(n2943), .ZN(n2960) );
  OR2_X1 U2909 ( .A1(n2785), .A2(n2257), .ZN(n2943) );
  OR2_X1 U2910 ( .A1(n2961), .A2(n2962), .ZN(n2942) );
  AND2_X1 U2911 ( .A1(n2936), .A2(n2939), .ZN(n2962) );
  AND2_X1 U2912 ( .A1(n2963), .A2(n2938), .ZN(n2961) );
  OR2_X1 U2913 ( .A1(n2964), .A2(n2965), .ZN(n2938) );
  AND2_X1 U2914 ( .A1(n2935), .A2(n2934), .ZN(n2965) );
  AND2_X1 U2915 ( .A1(n2932), .A2(n2966), .ZN(n2964) );
  OR2_X1 U2916 ( .A1(n2934), .A2(n2935), .ZN(n2966) );
  OR2_X1 U2917 ( .A1(n2785), .A2(n2355), .ZN(n2935) );
  OR2_X1 U2918 ( .A1(n2967), .A2(n2968), .ZN(n2934) );
  AND2_X1 U2919 ( .A1(n2929), .A2(n2930), .ZN(n2968) );
  AND2_X1 U2920 ( .A1(n2969), .A2(n2931), .ZN(n2967) );
  OR2_X1 U2921 ( .A1(n2970), .A2(n2971), .ZN(n2931) );
  AND2_X1 U2922 ( .A1(n2925), .A2(n2926), .ZN(n2971) );
  AND2_X1 U2923 ( .A1(n2972), .A2(n2927), .ZN(n2970) );
  OR2_X1 U2924 ( .A1(n2973), .A2(n2974), .ZN(n2927) );
  AND2_X1 U2925 ( .A1(n2921), .A2(n2922), .ZN(n2974) );
  AND2_X1 U2926 ( .A1(n2975), .A2(n2923), .ZN(n2973) );
  OR2_X1 U2927 ( .A1(n2976), .A2(n2977), .ZN(n2923) );
  AND2_X1 U2928 ( .A1(n2917), .A2(n2918), .ZN(n2977) );
  AND2_X1 U2929 ( .A1(n2978), .A2(n2919), .ZN(n2976) );
  OR2_X1 U2930 ( .A1(n2979), .A2(n2980), .ZN(n2919) );
  AND2_X1 U2931 ( .A1(n2913), .A2(n2914), .ZN(n2980) );
  AND2_X1 U2932 ( .A1(n2981), .A2(n2915), .ZN(n2979) );
  OR2_X1 U2933 ( .A1(n2982), .A2(n2983), .ZN(n2915) );
  AND2_X1 U2934 ( .A1(n2909), .A2(n2910), .ZN(n2983) );
  AND2_X1 U2935 ( .A1(n2984), .A2(n2911), .ZN(n2982) );
  OR2_X1 U2936 ( .A1(n2985), .A2(n2986), .ZN(n2911) );
  AND2_X1 U2937 ( .A1(n2905), .A2(n2906), .ZN(n2986) );
  AND2_X1 U2938 ( .A1(n2987), .A2(n2907), .ZN(n2985) );
  OR2_X1 U2939 ( .A1(n2988), .A2(n2989), .ZN(n2907) );
  AND2_X1 U2940 ( .A1(n2901), .A2(n2903), .ZN(n2989) );
  AND2_X1 U2941 ( .A1(n2990), .A2(n2902), .ZN(n2988) );
  OR2_X1 U2942 ( .A1(n2991), .A2(n2992), .ZN(n2902) );
  AND2_X1 U2943 ( .A1(n2897), .A2(n2899), .ZN(n2992) );
  AND2_X1 U2944 ( .A1(n2993), .A2(n2994), .ZN(n2991) );
  OR2_X1 U2945 ( .A1(n2899), .A2(n2897), .ZN(n2994) );
  OR2_X1 U2946 ( .A1(n2785), .A2(n2480), .ZN(n2897) );
  OR2_X1 U2947 ( .A1(n2481), .A2(n2995), .ZN(n2899) );
  OR2_X1 U2948 ( .A1(n2895), .A2(n2785), .ZN(n2995) );
  INV_X1 U2949 ( .A(n2898), .ZN(n2993) );
  OR2_X1 U2950 ( .A1(n2996), .A2(n2997), .ZN(n2898) );
  AND2_X1 U2951 ( .A1(n2998), .A2(n2999), .ZN(n2997) );
  OR2_X1 U2952 ( .A1(n3000), .A2(n2045), .ZN(n2999) );
  AND2_X1 U2953 ( .A1(n2895), .A2(n2039), .ZN(n3000) );
  AND2_X1 U2954 ( .A1(n2890), .A2(n3001), .ZN(n2996) );
  OR2_X1 U2955 ( .A1(n3002), .A2(n2049), .ZN(n3001) );
  AND2_X1 U2956 ( .A1(n3003), .A2(n2051), .ZN(n3002) );
  OR2_X1 U2957 ( .A1(n2903), .A2(n2901), .ZN(n2990) );
  XOR2_X1 U2958 ( .A(n3004), .B(n3005), .Z(n2901) );
  XNOR2_X1 U2959 ( .A(n3006), .B(n3007), .ZN(n3004) );
  OR2_X1 U2960 ( .A1(n2490), .A2(n2785), .ZN(n2903) );
  OR2_X1 U2961 ( .A1(n2906), .A2(n2905), .ZN(n2987) );
  XNOR2_X1 U2962 ( .A(n3008), .B(n3009), .ZN(n2905) );
  XNOR2_X1 U2963 ( .A(n3010), .B(n3011), .ZN(n3008) );
  OR2_X1 U2964 ( .A1(n2495), .A2(n2785), .ZN(n2906) );
  OR2_X1 U2965 ( .A1(n2910), .A2(n2909), .ZN(n2984) );
  XNOR2_X1 U2966 ( .A(n3012), .B(n3013), .ZN(n2909) );
  XNOR2_X1 U2967 ( .A(n3014), .B(n3015), .ZN(n3012) );
  OR2_X1 U2968 ( .A1(n2500), .A2(n2785), .ZN(n2910) );
  OR2_X1 U2969 ( .A1(n2914), .A2(n2913), .ZN(n2981) );
  XNOR2_X1 U2970 ( .A(n3016), .B(n3017), .ZN(n2913) );
  XNOR2_X1 U2971 ( .A(n3018), .B(n3019), .ZN(n3016) );
  OR2_X1 U2972 ( .A1(n2505), .A2(n2785), .ZN(n2914) );
  OR2_X1 U2973 ( .A1(n2918), .A2(n2917), .ZN(n2978) );
  XNOR2_X1 U2974 ( .A(n3020), .B(n3021), .ZN(n2917) );
  XNOR2_X1 U2975 ( .A(n3022), .B(n3023), .ZN(n3020) );
  OR2_X1 U2976 ( .A1(n2510), .A2(n2785), .ZN(n2918) );
  OR2_X1 U2977 ( .A1(n2922), .A2(n2921), .ZN(n2975) );
  XNOR2_X1 U2978 ( .A(n3024), .B(n3025), .ZN(n2921) );
  XNOR2_X1 U2979 ( .A(n3026), .B(n3027), .ZN(n3024) );
  OR2_X1 U2980 ( .A1(n2515), .A2(n2785), .ZN(n2922) );
  OR2_X1 U2981 ( .A1(n2926), .A2(n2925), .ZN(n2972) );
  XNOR2_X1 U2982 ( .A(n3028), .B(n3029), .ZN(n2925) );
  XNOR2_X1 U2983 ( .A(n3030), .B(n3031), .ZN(n3028) );
  OR2_X1 U2984 ( .A1(n2520), .A2(n2785), .ZN(n2926) );
  OR2_X1 U2985 ( .A1(n2930), .A2(n2929), .ZN(n2969) );
  XNOR2_X1 U2986 ( .A(n3032), .B(n3033), .ZN(n2929) );
  XNOR2_X1 U2987 ( .A(n3034), .B(n3035), .ZN(n3032) );
  OR2_X1 U2988 ( .A1(n2525), .A2(n2785), .ZN(n2930) );
  XOR2_X1 U2989 ( .A(n3036), .B(n3037), .Z(n2932) );
  XOR2_X1 U2990 ( .A(n3038), .B(n3039), .Z(n3037) );
  OR2_X1 U2991 ( .A1(n2939), .A2(n2936), .ZN(n2963) );
  XOR2_X1 U2992 ( .A(n3040), .B(n3041), .Z(n2936) );
  XOR2_X1 U2993 ( .A(n3042), .B(n3043), .Z(n3041) );
  OR2_X1 U2994 ( .A1(n2785), .A2(n2308), .ZN(n2939) );
  INV_X1 U2995 ( .A(n2780), .ZN(n2785) );
  XOR2_X1 U2996 ( .A(n3044), .B(n3045), .Z(n2780) );
  XNOR2_X1 U2997 ( .A(c_10_), .B(d_10_), .ZN(n3044) );
  XOR2_X1 U2998 ( .A(n3046), .B(n3047), .Z(n2940) );
  XOR2_X1 U2999 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR2_X1 U3000 ( .A(n3050), .B(n3051), .Z(n2944) );
  XOR2_X1 U3001 ( .A(n3052), .B(n3053), .Z(n3051) );
  XNOR2_X1 U3002 ( .A(n3054), .B(n3055), .ZN(n2948) );
  XNOR2_X1 U3003 ( .A(n3056), .B(n3057), .ZN(n3054) );
  XNOR2_X1 U3004 ( .A(n3058), .B(n3059), .ZN(n2371) );
  XNOR2_X1 U3005 ( .A(n3060), .B(n3061), .ZN(n3058) );
  INV_X1 U3006 ( .A(n2010), .ZN(n2369) );
  OR2_X1 U3007 ( .A1(n3062), .A2(n2367), .ZN(n2010) );
  INV_X1 U3008 ( .A(n3063), .ZN(n2367) );
  OR2_X1 U3009 ( .A1(n3064), .A2(n3065), .ZN(n3063) );
  AND2_X1 U3010 ( .A1(n3064), .A2(n3065), .ZN(n3062) );
  OR2_X1 U3011 ( .A1(n3066), .A2(n3067), .ZN(n3065) );
  AND2_X1 U3012 ( .A1(n3061), .A2(n3060), .ZN(n3067) );
  AND2_X1 U3013 ( .A1(n3059), .A2(n3068), .ZN(n3066) );
  OR2_X1 U3014 ( .A1(n3060), .A2(n3061), .ZN(n3068) );
  OR2_X1 U3015 ( .A1(n2895), .A2(n2187), .ZN(n3061) );
  OR2_X1 U3016 ( .A1(n3069), .A2(n3070), .ZN(n3060) );
  AND2_X1 U3017 ( .A1(n3057), .A2(n3056), .ZN(n3070) );
  AND2_X1 U3018 ( .A1(n3055), .A2(n3071), .ZN(n3069) );
  OR2_X1 U3019 ( .A1(n3056), .A2(n3057), .ZN(n3071) );
  OR2_X1 U3020 ( .A1(n2895), .A2(n2224), .ZN(n3057) );
  OR2_X1 U3021 ( .A1(n3072), .A2(n3073), .ZN(n3056) );
  AND2_X1 U3022 ( .A1(n3053), .A2(n3052), .ZN(n3073) );
  AND2_X1 U3023 ( .A1(n3050), .A2(n3074), .ZN(n3072) );
  OR2_X1 U3024 ( .A1(n3052), .A2(n3053), .ZN(n3074) );
  OR2_X1 U3025 ( .A1(n2895), .A2(n2257), .ZN(n3053) );
  OR2_X1 U3026 ( .A1(n3075), .A2(n3076), .ZN(n3052) );
  AND2_X1 U3027 ( .A1(n3049), .A2(n3048), .ZN(n3076) );
  AND2_X1 U3028 ( .A1(n3046), .A2(n3077), .ZN(n3075) );
  OR2_X1 U3029 ( .A1(n3048), .A2(n3049), .ZN(n3077) );
  OR2_X1 U3030 ( .A1(n2895), .A2(n2308), .ZN(n3049) );
  OR2_X1 U3031 ( .A1(n3078), .A2(n3079), .ZN(n3048) );
  AND2_X1 U3032 ( .A1(n3040), .A2(n3043), .ZN(n3079) );
  AND2_X1 U3033 ( .A1(n3080), .A2(n3042), .ZN(n3078) );
  OR2_X1 U3034 ( .A1(n3081), .A2(n3082), .ZN(n3042) );
  AND2_X1 U3035 ( .A1(n3039), .A2(n3038), .ZN(n3082) );
  AND2_X1 U3036 ( .A1(n3036), .A2(n3083), .ZN(n3081) );
  OR2_X1 U3037 ( .A1(n3038), .A2(n3039), .ZN(n3083) );
  OR2_X1 U3038 ( .A1(n2895), .A2(n2525), .ZN(n3039) );
  OR2_X1 U3039 ( .A1(n3084), .A2(n3085), .ZN(n3038) );
  AND2_X1 U3040 ( .A1(n3033), .A2(n3034), .ZN(n3085) );
  AND2_X1 U3041 ( .A1(n3086), .A2(n3035), .ZN(n3084) );
  OR2_X1 U3042 ( .A1(n3087), .A2(n3088), .ZN(n3035) );
  AND2_X1 U3043 ( .A1(n3029), .A2(n3030), .ZN(n3088) );
  AND2_X1 U3044 ( .A1(n3089), .A2(n3031), .ZN(n3087) );
  OR2_X1 U3045 ( .A1(n3090), .A2(n3091), .ZN(n3031) );
  AND2_X1 U3046 ( .A1(n3025), .A2(n3026), .ZN(n3091) );
  AND2_X1 U3047 ( .A1(n3092), .A2(n3027), .ZN(n3090) );
  OR2_X1 U3048 ( .A1(n3093), .A2(n3094), .ZN(n3027) );
  AND2_X1 U3049 ( .A1(n3021), .A2(n3022), .ZN(n3094) );
  AND2_X1 U3050 ( .A1(n3095), .A2(n3023), .ZN(n3093) );
  OR2_X1 U3051 ( .A1(n3096), .A2(n3097), .ZN(n3023) );
  AND2_X1 U3052 ( .A1(n3017), .A2(n3018), .ZN(n3097) );
  AND2_X1 U3053 ( .A1(n3098), .A2(n3019), .ZN(n3096) );
  OR2_X1 U3054 ( .A1(n3099), .A2(n3100), .ZN(n3019) );
  AND2_X1 U3055 ( .A1(n3013), .A2(n3014), .ZN(n3100) );
  AND2_X1 U3056 ( .A1(n3101), .A2(n3015), .ZN(n3099) );
  OR2_X1 U3057 ( .A1(n3102), .A2(n3103), .ZN(n3015) );
  AND2_X1 U3058 ( .A1(n3009), .A2(n3011), .ZN(n3103) );
  AND2_X1 U3059 ( .A1(n3104), .A2(n3010), .ZN(n3102) );
  OR2_X1 U3060 ( .A1(n3105), .A2(n3106), .ZN(n3010) );
  AND2_X1 U3061 ( .A1(n3005), .A2(n3007), .ZN(n3106) );
  AND2_X1 U3062 ( .A1(n3107), .A2(n3108), .ZN(n3105) );
  OR2_X1 U3063 ( .A1(n3007), .A2(n3005), .ZN(n3108) );
  OR2_X1 U3064 ( .A1(n2895), .A2(n2480), .ZN(n3005) );
  OR2_X1 U3065 ( .A1(n2481), .A2(n3109), .ZN(n3007) );
  OR2_X1 U3066 ( .A1(n3003), .A2(n2895), .ZN(n3109) );
  INV_X1 U3067 ( .A(n3006), .ZN(n3107) );
  OR2_X1 U3068 ( .A1(n3110), .A2(n3111), .ZN(n3006) );
  AND2_X1 U3069 ( .A1(n3112), .A2(n3113), .ZN(n3111) );
  OR2_X1 U3070 ( .A1(n3114), .A2(n2045), .ZN(n3113) );
  AND2_X1 U3071 ( .A1(n3003), .A2(n2039), .ZN(n3114) );
  AND2_X1 U3072 ( .A1(n2998), .A2(n3115), .ZN(n3110) );
  OR2_X1 U3073 ( .A1(n3116), .A2(n2049), .ZN(n3115) );
  AND2_X1 U3074 ( .A1(n2326), .A2(n2051), .ZN(n3116) );
  OR2_X1 U3075 ( .A1(n3011), .A2(n3009), .ZN(n3104) );
  XOR2_X1 U3076 ( .A(n3117), .B(n3118), .Z(n3009) );
  XNOR2_X1 U3077 ( .A(n3119), .B(n3120), .ZN(n3117) );
  OR2_X1 U3078 ( .A1(n2490), .A2(n2895), .ZN(n3011) );
  OR2_X1 U3079 ( .A1(n3014), .A2(n3013), .ZN(n3101) );
  XNOR2_X1 U3080 ( .A(n3121), .B(n3122), .ZN(n3013) );
  XNOR2_X1 U3081 ( .A(n3123), .B(n3124), .ZN(n3121) );
  OR2_X1 U3082 ( .A1(n2495), .A2(n2895), .ZN(n3014) );
  OR2_X1 U3083 ( .A1(n3018), .A2(n3017), .ZN(n3098) );
  XNOR2_X1 U3084 ( .A(n3125), .B(n3126), .ZN(n3017) );
  XNOR2_X1 U3085 ( .A(n3127), .B(n3128), .ZN(n3125) );
  OR2_X1 U3086 ( .A1(n2500), .A2(n2895), .ZN(n3018) );
  OR2_X1 U3087 ( .A1(n3022), .A2(n3021), .ZN(n3095) );
  XNOR2_X1 U3088 ( .A(n3129), .B(n3130), .ZN(n3021) );
  XNOR2_X1 U3089 ( .A(n3131), .B(n3132), .ZN(n3129) );
  OR2_X1 U3090 ( .A1(n2505), .A2(n2895), .ZN(n3022) );
  OR2_X1 U3091 ( .A1(n3026), .A2(n3025), .ZN(n3092) );
  XNOR2_X1 U3092 ( .A(n3133), .B(n3134), .ZN(n3025) );
  XNOR2_X1 U3093 ( .A(n3135), .B(n3136), .ZN(n3133) );
  OR2_X1 U3094 ( .A1(n2510), .A2(n2895), .ZN(n3026) );
  OR2_X1 U3095 ( .A1(n3030), .A2(n3029), .ZN(n3089) );
  XNOR2_X1 U3096 ( .A(n3137), .B(n3138), .ZN(n3029) );
  XNOR2_X1 U3097 ( .A(n3139), .B(n3140), .ZN(n3137) );
  OR2_X1 U3098 ( .A1(n2515), .A2(n2895), .ZN(n3030) );
  OR2_X1 U3099 ( .A1(n3034), .A2(n3033), .ZN(n3086) );
  XNOR2_X1 U3100 ( .A(n3141), .B(n3142), .ZN(n3033) );
  XNOR2_X1 U3101 ( .A(n3143), .B(n3144), .ZN(n3141) );
  OR2_X1 U3102 ( .A1(n2520), .A2(n2895), .ZN(n3034) );
  XOR2_X1 U3103 ( .A(n3145), .B(n3146), .Z(n3036) );
  XOR2_X1 U3104 ( .A(n3147), .B(n3148), .Z(n3146) );
  OR2_X1 U3105 ( .A1(n3043), .A2(n3040), .ZN(n3080) );
  XOR2_X1 U3106 ( .A(n3149), .B(n3150), .Z(n3040) );
  XOR2_X1 U3107 ( .A(n3151), .B(n3152), .Z(n3150) );
  OR2_X1 U3108 ( .A1(n2895), .A2(n2355), .ZN(n3043) );
  INV_X1 U3109 ( .A(n2890), .ZN(n2895) );
  XOR2_X1 U3110 ( .A(n3153), .B(n3154), .Z(n2890) );
  XNOR2_X1 U3111 ( .A(c_9_), .B(d_9_), .ZN(n3153) );
  XOR2_X1 U3112 ( .A(n3155), .B(n3156), .Z(n3046) );
  XOR2_X1 U3113 ( .A(n3157), .B(n3158), .Z(n3156) );
  XOR2_X1 U3114 ( .A(n3159), .B(n3160), .Z(n3050) );
  XOR2_X1 U3115 ( .A(n3161), .B(n3162), .Z(n3160) );
  XOR2_X1 U3116 ( .A(n3163), .B(n3164), .Z(n3055) );
  XOR2_X1 U3117 ( .A(n3165), .B(n3166), .Z(n3164) );
  XNOR2_X1 U3118 ( .A(n3167), .B(n3168), .ZN(n3059) );
  XNOR2_X1 U3119 ( .A(n3169), .B(n3170), .ZN(n3167) );
  XOR2_X1 U3120 ( .A(n2323), .B(n3171), .Z(n3064) );
  XOR2_X1 U3121 ( .A(n2322), .B(n2321), .Z(n3171) );
  OR2_X1 U3122 ( .A1(n3003), .A2(n2187), .ZN(n2321) );
  OR2_X1 U3123 ( .A1(n3172), .A2(n3173), .ZN(n2322) );
  AND2_X1 U3124 ( .A1(n3170), .A2(n3169), .ZN(n3173) );
  AND2_X1 U3125 ( .A1(n3168), .A2(n3174), .ZN(n3172) );
  OR2_X1 U3126 ( .A1(n3169), .A2(n3170), .ZN(n3174) );
  OR2_X1 U3127 ( .A1(n3003), .A2(n2224), .ZN(n3170) );
  OR2_X1 U3128 ( .A1(n3175), .A2(n3176), .ZN(n3169) );
  AND2_X1 U3129 ( .A1(n3166), .A2(n3165), .ZN(n3176) );
  AND2_X1 U3130 ( .A1(n3163), .A2(n3177), .ZN(n3175) );
  OR2_X1 U3131 ( .A1(n3165), .A2(n3166), .ZN(n3177) );
  OR2_X1 U3132 ( .A1(n3003), .A2(n2257), .ZN(n3166) );
  OR2_X1 U3133 ( .A1(n3178), .A2(n3179), .ZN(n3165) );
  AND2_X1 U3134 ( .A1(n3162), .A2(n3161), .ZN(n3179) );
  AND2_X1 U3135 ( .A1(n3159), .A2(n3180), .ZN(n3178) );
  OR2_X1 U3136 ( .A1(n3161), .A2(n3162), .ZN(n3180) );
  OR2_X1 U3137 ( .A1(n3003), .A2(n2308), .ZN(n3162) );
  OR2_X1 U3138 ( .A1(n3181), .A2(n3182), .ZN(n3161) );
  AND2_X1 U3139 ( .A1(n3158), .A2(n3157), .ZN(n3182) );
  AND2_X1 U3140 ( .A1(n3155), .A2(n3183), .ZN(n3181) );
  OR2_X1 U3141 ( .A1(n3157), .A2(n3158), .ZN(n3183) );
  OR2_X1 U3142 ( .A1(n3003), .A2(n2355), .ZN(n3158) );
  OR2_X1 U3143 ( .A1(n3184), .A2(n3185), .ZN(n3157) );
  AND2_X1 U3144 ( .A1(n3149), .A2(n3152), .ZN(n3185) );
  AND2_X1 U3145 ( .A1(n3186), .A2(n3151), .ZN(n3184) );
  OR2_X1 U3146 ( .A1(n3187), .A2(n3188), .ZN(n3151) );
  AND2_X1 U3147 ( .A1(n3148), .A2(n3147), .ZN(n3188) );
  AND2_X1 U3148 ( .A1(n3145), .A2(n3189), .ZN(n3187) );
  OR2_X1 U3149 ( .A1(n3147), .A2(n3148), .ZN(n3189) );
  OR2_X1 U3150 ( .A1(n3003), .A2(n2520), .ZN(n3148) );
  OR2_X1 U3151 ( .A1(n3190), .A2(n3191), .ZN(n3147) );
  AND2_X1 U3152 ( .A1(n3142), .A2(n3143), .ZN(n3191) );
  AND2_X1 U3153 ( .A1(n3192), .A2(n3144), .ZN(n3190) );
  OR2_X1 U3154 ( .A1(n3193), .A2(n3194), .ZN(n3144) );
  AND2_X1 U3155 ( .A1(n3138), .A2(n3139), .ZN(n3194) );
  AND2_X1 U3156 ( .A1(n3195), .A2(n3140), .ZN(n3193) );
  OR2_X1 U3157 ( .A1(n3196), .A2(n3197), .ZN(n3140) );
  AND2_X1 U3158 ( .A1(n3134), .A2(n3135), .ZN(n3197) );
  AND2_X1 U3159 ( .A1(n3198), .A2(n3136), .ZN(n3196) );
  OR2_X1 U3160 ( .A1(n3199), .A2(n3200), .ZN(n3136) );
  AND2_X1 U3161 ( .A1(n3130), .A2(n3131), .ZN(n3200) );
  AND2_X1 U3162 ( .A1(n3201), .A2(n3132), .ZN(n3199) );
  OR2_X1 U3163 ( .A1(n3202), .A2(n3203), .ZN(n3132) );
  AND2_X1 U3164 ( .A1(n3126), .A2(n3127), .ZN(n3203) );
  AND2_X1 U3165 ( .A1(n3204), .A2(n3128), .ZN(n3202) );
  OR2_X1 U3166 ( .A1(n3205), .A2(n3206), .ZN(n3128) );
  AND2_X1 U3167 ( .A1(n3122), .A2(n3124), .ZN(n3206) );
  AND2_X1 U3168 ( .A1(n3207), .A2(n3123), .ZN(n3205) );
  OR2_X1 U3169 ( .A1(n3208), .A2(n3209), .ZN(n3123) );
  AND2_X1 U3170 ( .A1(n3118), .A2(n3120), .ZN(n3209) );
  AND2_X1 U3171 ( .A1(n3210), .A2(n3211), .ZN(n3208) );
  OR2_X1 U3172 ( .A1(n3120), .A2(n3118), .ZN(n3211) );
  OR2_X1 U3173 ( .A1(n3003), .A2(n2480), .ZN(n3118) );
  OR2_X1 U3174 ( .A1(n2481), .A2(n3212), .ZN(n3120) );
  OR2_X1 U3175 ( .A1(n2326), .A2(n3003), .ZN(n3212) );
  INV_X1 U3176 ( .A(n3119), .ZN(n3210) );
  OR2_X1 U3177 ( .A1(n3213), .A2(n3214), .ZN(n3119) );
  AND2_X1 U3178 ( .A1(n3215), .A2(n3216), .ZN(n3214) );
  OR2_X1 U3179 ( .A1(n3217), .A2(n2045), .ZN(n3216) );
  AND2_X1 U3180 ( .A1(n2326), .A2(n2039), .ZN(n3217) );
  AND2_X1 U3181 ( .A1(n3112), .A2(n3218), .ZN(n3213) );
  OR2_X1 U3182 ( .A1(n3219), .A2(n2049), .ZN(n3218) );
  AND2_X1 U3183 ( .A1(n2286), .A2(n2051), .ZN(n3219) );
  OR2_X1 U3184 ( .A1(n3124), .A2(n3122), .ZN(n3207) );
  XOR2_X1 U3185 ( .A(n3220), .B(n3221), .Z(n3122) );
  XNOR2_X1 U3186 ( .A(n3222), .B(n3223), .ZN(n3220) );
  OR2_X1 U3187 ( .A1(n2490), .A2(n3003), .ZN(n3124) );
  OR2_X1 U3188 ( .A1(n3127), .A2(n3126), .ZN(n3204) );
  XNOR2_X1 U3189 ( .A(n3224), .B(n3225), .ZN(n3126) );
  XNOR2_X1 U3190 ( .A(n3226), .B(n3227), .ZN(n3224) );
  OR2_X1 U3191 ( .A1(n2495), .A2(n3003), .ZN(n3127) );
  OR2_X1 U3192 ( .A1(n3131), .A2(n3130), .ZN(n3201) );
  XNOR2_X1 U3193 ( .A(n3228), .B(n3229), .ZN(n3130) );
  XNOR2_X1 U3194 ( .A(n3230), .B(n3231), .ZN(n3228) );
  OR2_X1 U3195 ( .A1(n2500), .A2(n3003), .ZN(n3131) );
  OR2_X1 U3196 ( .A1(n3135), .A2(n3134), .ZN(n3198) );
  XNOR2_X1 U3197 ( .A(n3232), .B(n3233), .ZN(n3134) );
  XNOR2_X1 U3198 ( .A(n3234), .B(n3235), .ZN(n3232) );
  OR2_X1 U3199 ( .A1(n2505), .A2(n3003), .ZN(n3135) );
  OR2_X1 U3200 ( .A1(n3139), .A2(n3138), .ZN(n3195) );
  XNOR2_X1 U3201 ( .A(n3236), .B(n3237), .ZN(n3138) );
  XNOR2_X1 U3202 ( .A(n3238), .B(n3239), .ZN(n3236) );
  OR2_X1 U3203 ( .A1(n2510), .A2(n3003), .ZN(n3139) );
  OR2_X1 U3204 ( .A1(n3143), .A2(n3142), .ZN(n3192) );
  XNOR2_X1 U3205 ( .A(n3240), .B(n3241), .ZN(n3142) );
  XNOR2_X1 U3206 ( .A(n3242), .B(n3243), .ZN(n3240) );
  OR2_X1 U3207 ( .A1(n2515), .A2(n3003), .ZN(n3143) );
  XOR2_X1 U3208 ( .A(n3244), .B(n3245), .Z(n3145) );
  XOR2_X1 U3209 ( .A(n3246), .B(n3247), .Z(n3245) );
  OR2_X1 U3210 ( .A1(n3152), .A2(n3149), .ZN(n3186) );
  XOR2_X1 U3211 ( .A(n3248), .B(n3249), .Z(n3149) );
  XOR2_X1 U3212 ( .A(n3250), .B(n3251), .Z(n3249) );
  OR2_X1 U3213 ( .A1(n3003), .A2(n2525), .ZN(n3152) );
  INV_X1 U3214 ( .A(n2998), .ZN(n3003) );
  XOR2_X1 U3215 ( .A(n3252), .B(n3253), .Z(n2998) );
  XNOR2_X1 U3216 ( .A(c_8_), .B(d_8_), .ZN(n3252) );
  XOR2_X1 U3217 ( .A(n3254), .B(n3255), .Z(n3155) );
  XOR2_X1 U3218 ( .A(n3256), .B(n3257), .Z(n3255) );
  XOR2_X1 U3219 ( .A(n3258), .B(n3259), .Z(n3159) );
  XOR2_X1 U3220 ( .A(n3260), .B(n3261), .Z(n3259) );
  XNOR2_X1 U3221 ( .A(n3262), .B(n3263), .ZN(n3163) );
  XNOR2_X1 U3222 ( .A(n3264), .B(n3265), .ZN(n3262) );
  XOR2_X1 U3223 ( .A(n3266), .B(n3267), .Z(n3168) );
  XOR2_X1 U3224 ( .A(n3268), .B(n3269), .Z(n3267) );
  XOR2_X1 U3225 ( .A(n2331), .B(n3270), .Z(n2323) );
  XOR2_X1 U3226 ( .A(n2330), .B(n2329), .Z(n3270) );
  OR2_X1 U3227 ( .A1(n2326), .A2(n2224), .ZN(n2329) );
  OR2_X1 U3228 ( .A1(n3271), .A2(n3272), .ZN(n2330) );
  AND2_X1 U3229 ( .A1(n3269), .A2(n3268), .ZN(n3272) );
  AND2_X1 U3230 ( .A1(n3266), .A2(n3273), .ZN(n3271) );
  OR2_X1 U3231 ( .A1(n3268), .A2(n3269), .ZN(n3273) );
  OR2_X1 U3232 ( .A1(n2326), .A2(n2257), .ZN(n3269) );
  OR2_X1 U3233 ( .A1(n3274), .A2(n3275), .ZN(n3268) );
  AND2_X1 U3234 ( .A1(n3265), .A2(n3264), .ZN(n3275) );
  AND2_X1 U3235 ( .A1(n3263), .A2(n3276), .ZN(n3274) );
  OR2_X1 U3236 ( .A1(n3264), .A2(n3265), .ZN(n3276) );
  OR2_X1 U3237 ( .A1(n2326), .A2(n2308), .ZN(n3265) );
  OR2_X1 U3238 ( .A1(n3277), .A2(n3278), .ZN(n3264) );
  AND2_X1 U3239 ( .A1(n3261), .A2(n3260), .ZN(n3278) );
  AND2_X1 U3240 ( .A1(n3258), .A2(n3279), .ZN(n3277) );
  OR2_X1 U3241 ( .A1(n3260), .A2(n3261), .ZN(n3279) );
  OR2_X1 U3242 ( .A1(n2326), .A2(n2355), .ZN(n3261) );
  OR2_X1 U3243 ( .A1(n3280), .A2(n3281), .ZN(n3260) );
  AND2_X1 U3244 ( .A1(n3257), .A2(n3256), .ZN(n3281) );
  AND2_X1 U3245 ( .A1(n3254), .A2(n3282), .ZN(n3280) );
  OR2_X1 U3246 ( .A1(n3256), .A2(n3257), .ZN(n3282) );
  OR2_X1 U3247 ( .A1(n2326), .A2(n2525), .ZN(n3257) );
  OR2_X1 U3248 ( .A1(n3283), .A2(n3284), .ZN(n3256) );
  AND2_X1 U3249 ( .A1(n3248), .A2(n3251), .ZN(n3284) );
  AND2_X1 U3250 ( .A1(n3285), .A2(n3250), .ZN(n3283) );
  OR2_X1 U3251 ( .A1(n3286), .A2(n3287), .ZN(n3250) );
  AND2_X1 U3252 ( .A1(n3247), .A2(n3246), .ZN(n3287) );
  AND2_X1 U3253 ( .A1(n3244), .A2(n3288), .ZN(n3286) );
  OR2_X1 U3254 ( .A1(n3246), .A2(n3247), .ZN(n3288) );
  OR2_X1 U3255 ( .A1(n2326), .A2(n2515), .ZN(n3247) );
  OR2_X1 U3256 ( .A1(n3289), .A2(n3290), .ZN(n3246) );
  AND2_X1 U3257 ( .A1(n3241), .A2(n3242), .ZN(n3290) );
  AND2_X1 U3258 ( .A1(n3291), .A2(n3243), .ZN(n3289) );
  OR2_X1 U3259 ( .A1(n3292), .A2(n3293), .ZN(n3243) );
  AND2_X1 U3260 ( .A1(n3237), .A2(n3238), .ZN(n3293) );
  AND2_X1 U3261 ( .A1(n3294), .A2(n3239), .ZN(n3292) );
  OR2_X1 U3262 ( .A1(n3295), .A2(n3296), .ZN(n3239) );
  AND2_X1 U3263 ( .A1(n3233), .A2(n3234), .ZN(n3296) );
  AND2_X1 U3264 ( .A1(n3297), .A2(n3235), .ZN(n3295) );
  OR2_X1 U3265 ( .A1(n3298), .A2(n3299), .ZN(n3235) );
  AND2_X1 U3266 ( .A1(n3229), .A2(n3230), .ZN(n3299) );
  AND2_X1 U3267 ( .A1(n3300), .A2(n3231), .ZN(n3298) );
  OR2_X1 U3268 ( .A1(n3301), .A2(n3302), .ZN(n3231) );
  AND2_X1 U3269 ( .A1(n3225), .A2(n3227), .ZN(n3302) );
  AND2_X1 U3270 ( .A1(n3303), .A2(n3226), .ZN(n3301) );
  OR2_X1 U3271 ( .A1(n3304), .A2(n3305), .ZN(n3226) );
  AND2_X1 U3272 ( .A1(n3221), .A2(n3223), .ZN(n3305) );
  AND2_X1 U3273 ( .A1(n3306), .A2(n3307), .ZN(n3304) );
  OR2_X1 U3274 ( .A1(n3223), .A2(n3221), .ZN(n3307) );
  OR2_X1 U3275 ( .A1(n2326), .A2(n2480), .ZN(n3221) );
  OR2_X1 U3276 ( .A1(n2481), .A2(n3308), .ZN(n3223) );
  OR2_X1 U3277 ( .A1(n2286), .A2(n2326), .ZN(n3308) );
  INV_X1 U3278 ( .A(n3222), .ZN(n3306) );
  OR2_X1 U3279 ( .A1(n3309), .A2(n3310), .ZN(n3222) );
  AND2_X1 U3280 ( .A1(n3311), .A2(n3312), .ZN(n3310) );
  OR2_X1 U3281 ( .A1(n3313), .A2(n2045), .ZN(n3312) );
  AND2_X1 U3282 ( .A1(n2286), .A2(n2039), .ZN(n3313) );
  AND2_X1 U3283 ( .A1(n3215), .A2(n3314), .ZN(n3309) );
  OR2_X1 U3284 ( .A1(n3315), .A2(n2049), .ZN(n3314) );
  AND2_X1 U3285 ( .A1(n2242), .A2(n2051), .ZN(n3315) );
  OR2_X1 U3286 ( .A1(n3227), .A2(n3225), .ZN(n3303) );
  XOR2_X1 U3287 ( .A(n3316), .B(n3317), .Z(n3225) );
  XNOR2_X1 U3288 ( .A(n3318), .B(n3319), .ZN(n3316) );
  OR2_X1 U3289 ( .A1(n2490), .A2(n2326), .ZN(n3227) );
  OR2_X1 U3290 ( .A1(n3230), .A2(n3229), .ZN(n3300) );
  XNOR2_X1 U3291 ( .A(n3320), .B(n3321), .ZN(n3229) );
  XNOR2_X1 U3292 ( .A(n3322), .B(n3323), .ZN(n3320) );
  OR2_X1 U3293 ( .A1(n2495), .A2(n2326), .ZN(n3230) );
  OR2_X1 U3294 ( .A1(n3234), .A2(n3233), .ZN(n3297) );
  XNOR2_X1 U3295 ( .A(n3324), .B(n3325), .ZN(n3233) );
  XNOR2_X1 U3296 ( .A(n3326), .B(n3327), .ZN(n3324) );
  OR2_X1 U3297 ( .A1(n2500), .A2(n2326), .ZN(n3234) );
  OR2_X1 U3298 ( .A1(n3238), .A2(n3237), .ZN(n3294) );
  XNOR2_X1 U3299 ( .A(n3328), .B(n3329), .ZN(n3237) );
  XNOR2_X1 U3300 ( .A(n3330), .B(n3331), .ZN(n3328) );
  OR2_X1 U3301 ( .A1(n2505), .A2(n2326), .ZN(n3238) );
  OR2_X1 U3302 ( .A1(n3242), .A2(n3241), .ZN(n3291) );
  XNOR2_X1 U3303 ( .A(n3332), .B(n3333), .ZN(n3241) );
  XNOR2_X1 U3304 ( .A(n3334), .B(n3335), .ZN(n3332) );
  OR2_X1 U3305 ( .A1(n2510), .A2(n2326), .ZN(n3242) );
  XOR2_X1 U3306 ( .A(n3336), .B(n3337), .Z(n3244) );
  XOR2_X1 U3307 ( .A(n3338), .B(n3339), .Z(n3337) );
  OR2_X1 U3308 ( .A1(n3251), .A2(n3248), .ZN(n3285) );
  XOR2_X1 U3309 ( .A(n3340), .B(n3341), .Z(n3248) );
  XOR2_X1 U3310 ( .A(n3342), .B(n3343), .Z(n3341) );
  OR2_X1 U3311 ( .A1(n2326), .A2(n2520), .ZN(n3251) );
  INV_X1 U3312 ( .A(n3112), .ZN(n2326) );
  XOR2_X1 U3313 ( .A(n3344), .B(n3345), .Z(n3112) );
  XNOR2_X1 U3314 ( .A(c_7_), .B(d_7_), .ZN(n3344) );
  XOR2_X1 U3315 ( .A(n3346), .B(n3347), .Z(n3254) );
  XOR2_X1 U3316 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR2_X1 U3317 ( .A(n3350), .B(n3351), .Z(n3258) );
  XOR2_X1 U3318 ( .A(n3352), .B(n3353), .Z(n3351) );
  XOR2_X1 U3319 ( .A(n3354), .B(n3355), .Z(n3263) );
  XOR2_X1 U3320 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR2_X1 U3321 ( .A(n3358), .B(n3359), .Z(n3266) );
  XOR2_X1 U3322 ( .A(n3360), .B(n3361), .Z(n3359) );
  XOR2_X1 U3323 ( .A(n2338), .B(n3362), .Z(n2331) );
  XOR2_X1 U3324 ( .A(n2337), .B(n2336), .Z(n3362) );
  OR2_X1 U3325 ( .A1(n2286), .A2(n2257), .ZN(n2336) );
  OR2_X1 U3326 ( .A1(n3363), .A2(n3364), .ZN(n2337) );
  AND2_X1 U3327 ( .A1(n3361), .A2(n3360), .ZN(n3364) );
  AND2_X1 U3328 ( .A1(n3358), .A2(n3365), .ZN(n3363) );
  OR2_X1 U3329 ( .A1(n3360), .A2(n3361), .ZN(n3365) );
  OR2_X1 U3330 ( .A1(n2286), .A2(n2308), .ZN(n3361) );
  OR2_X1 U3331 ( .A1(n3366), .A2(n3367), .ZN(n3360) );
  AND2_X1 U3332 ( .A1(n3357), .A2(n3356), .ZN(n3367) );
  AND2_X1 U3333 ( .A1(n3354), .A2(n3368), .ZN(n3366) );
  OR2_X1 U3334 ( .A1(n3356), .A2(n3357), .ZN(n3368) );
  OR2_X1 U3335 ( .A1(n2286), .A2(n2355), .ZN(n3357) );
  OR2_X1 U3336 ( .A1(n3369), .A2(n3370), .ZN(n3356) );
  AND2_X1 U3337 ( .A1(n3353), .A2(n3352), .ZN(n3370) );
  AND2_X1 U3338 ( .A1(n3350), .A2(n3371), .ZN(n3369) );
  OR2_X1 U3339 ( .A1(n3352), .A2(n3353), .ZN(n3371) );
  OR2_X1 U3340 ( .A1(n2286), .A2(n2525), .ZN(n3353) );
  OR2_X1 U3341 ( .A1(n3372), .A2(n3373), .ZN(n3352) );
  AND2_X1 U3342 ( .A1(n3349), .A2(n3348), .ZN(n3373) );
  AND2_X1 U3343 ( .A1(n3346), .A2(n3374), .ZN(n3372) );
  OR2_X1 U3344 ( .A1(n3348), .A2(n3349), .ZN(n3374) );
  OR2_X1 U3345 ( .A1(n2286), .A2(n2520), .ZN(n3349) );
  OR2_X1 U3346 ( .A1(n3375), .A2(n3376), .ZN(n3348) );
  AND2_X1 U3347 ( .A1(n3340), .A2(n3343), .ZN(n3376) );
  AND2_X1 U3348 ( .A1(n3377), .A2(n3342), .ZN(n3375) );
  OR2_X1 U3349 ( .A1(n3378), .A2(n3379), .ZN(n3342) );
  AND2_X1 U3350 ( .A1(n3339), .A2(n3338), .ZN(n3379) );
  AND2_X1 U3351 ( .A1(n3336), .A2(n3380), .ZN(n3378) );
  OR2_X1 U3352 ( .A1(n3338), .A2(n3339), .ZN(n3380) );
  OR2_X1 U3353 ( .A1(n2286), .A2(n2510), .ZN(n3339) );
  OR2_X1 U3354 ( .A1(n3381), .A2(n3382), .ZN(n3338) );
  AND2_X1 U3355 ( .A1(n3333), .A2(n3334), .ZN(n3382) );
  AND2_X1 U3356 ( .A1(n3383), .A2(n3335), .ZN(n3381) );
  OR2_X1 U3357 ( .A1(n3384), .A2(n3385), .ZN(n3335) );
  AND2_X1 U3358 ( .A1(n3329), .A2(n3330), .ZN(n3385) );
  AND2_X1 U3359 ( .A1(n3386), .A2(n3331), .ZN(n3384) );
  OR2_X1 U3360 ( .A1(n3387), .A2(n3388), .ZN(n3331) );
  AND2_X1 U3361 ( .A1(n3325), .A2(n3326), .ZN(n3388) );
  AND2_X1 U3362 ( .A1(n3389), .A2(n3327), .ZN(n3387) );
  OR2_X1 U3363 ( .A1(n3390), .A2(n3391), .ZN(n3327) );
  AND2_X1 U3364 ( .A1(n3321), .A2(n3323), .ZN(n3391) );
  AND2_X1 U3365 ( .A1(n3392), .A2(n3322), .ZN(n3390) );
  OR2_X1 U3366 ( .A1(n3393), .A2(n3394), .ZN(n3322) );
  AND2_X1 U3367 ( .A1(n3317), .A2(n3319), .ZN(n3394) );
  AND2_X1 U3368 ( .A1(n3395), .A2(n3396), .ZN(n3393) );
  OR2_X1 U3369 ( .A1(n3319), .A2(n3317), .ZN(n3396) );
  OR2_X1 U3370 ( .A1(n2286), .A2(n2480), .ZN(n3317) );
  OR2_X1 U3371 ( .A1(n2481), .A2(n3397), .ZN(n3319) );
  OR2_X1 U3372 ( .A1(n2242), .A2(n2286), .ZN(n3397) );
  INV_X1 U3373 ( .A(n3318), .ZN(n3395) );
  OR2_X1 U3374 ( .A1(n3398), .A2(n3399), .ZN(n3318) );
  AND2_X1 U3375 ( .A1(n3400), .A2(n3401), .ZN(n3399) );
  OR2_X1 U3376 ( .A1(n3402), .A2(n2045), .ZN(n3401) );
  AND2_X1 U3377 ( .A1(n2242), .A2(n2039), .ZN(n3402) );
  AND2_X1 U3378 ( .A1(n3311), .A2(n3403), .ZN(n3398) );
  OR2_X1 U3379 ( .A1(n3404), .A2(n2049), .ZN(n3403) );
  AND2_X1 U3380 ( .A1(n2216), .A2(n2051), .ZN(n3404) );
  OR2_X1 U3381 ( .A1(n3323), .A2(n3321), .ZN(n3392) );
  XOR2_X1 U3382 ( .A(n3405), .B(n3406), .Z(n3321) );
  XNOR2_X1 U3383 ( .A(n3407), .B(n3408), .ZN(n3405) );
  OR2_X1 U3384 ( .A1(n2490), .A2(n2286), .ZN(n3323) );
  OR2_X1 U3385 ( .A1(n3326), .A2(n3325), .ZN(n3389) );
  XNOR2_X1 U3386 ( .A(n3409), .B(n3410), .ZN(n3325) );
  XNOR2_X1 U3387 ( .A(n3411), .B(n3412), .ZN(n3409) );
  OR2_X1 U3388 ( .A1(n2495), .A2(n2286), .ZN(n3326) );
  OR2_X1 U3389 ( .A1(n3330), .A2(n3329), .ZN(n3386) );
  XNOR2_X1 U3390 ( .A(n3413), .B(n3414), .ZN(n3329) );
  XNOR2_X1 U3391 ( .A(n3415), .B(n3416), .ZN(n3413) );
  OR2_X1 U3392 ( .A1(n2500), .A2(n2286), .ZN(n3330) );
  OR2_X1 U3393 ( .A1(n3334), .A2(n3333), .ZN(n3383) );
  XNOR2_X1 U3394 ( .A(n3417), .B(n3418), .ZN(n3333) );
  XNOR2_X1 U3395 ( .A(n3419), .B(n3420), .ZN(n3417) );
  OR2_X1 U3396 ( .A1(n2505), .A2(n2286), .ZN(n3334) );
  XOR2_X1 U3397 ( .A(n3421), .B(n3422), .Z(n3336) );
  XOR2_X1 U3398 ( .A(n3423), .B(n3424), .Z(n3422) );
  OR2_X1 U3399 ( .A1(n3343), .A2(n3340), .ZN(n3377) );
  XOR2_X1 U3400 ( .A(n3425), .B(n3426), .Z(n3340) );
  XOR2_X1 U3401 ( .A(n3427), .B(n3428), .Z(n3426) );
  OR2_X1 U3402 ( .A1(n2286), .A2(n2515), .ZN(n3343) );
  INV_X1 U3403 ( .A(n3215), .ZN(n2286) );
  XOR2_X1 U3404 ( .A(n3429), .B(n3430), .Z(n3215) );
  XNOR2_X1 U3405 ( .A(c_6_), .B(d_6_), .ZN(n3429) );
  XOR2_X1 U3406 ( .A(n3431), .B(n3432), .Z(n3346) );
  XOR2_X1 U3407 ( .A(n3433), .B(n3434), .Z(n3432) );
  XOR2_X1 U3408 ( .A(n3435), .B(n3436), .Z(n3350) );
  XOR2_X1 U3409 ( .A(n3437), .B(n3438), .Z(n3436) );
  XOR2_X1 U3410 ( .A(n3439), .B(n3440), .Z(n3354) );
  XOR2_X1 U3411 ( .A(n3441), .B(n3442), .Z(n3440) );
  XOR2_X1 U3412 ( .A(n3443), .B(n3444), .Z(n3358) );
  XOR2_X1 U3413 ( .A(n3445), .B(n3446), .Z(n3444) );
  XOR2_X1 U3414 ( .A(n2345), .B(n3447), .Z(n2338) );
  XOR2_X1 U3415 ( .A(n2344), .B(n2343), .Z(n3447) );
  OR2_X1 U3416 ( .A1(n2242), .A2(n2308), .ZN(n2343) );
  OR2_X1 U3417 ( .A1(n3448), .A2(n3449), .ZN(n2344) );
  AND2_X1 U3418 ( .A1(n3446), .A2(n3445), .ZN(n3449) );
  AND2_X1 U3419 ( .A1(n3443), .A2(n3450), .ZN(n3448) );
  OR2_X1 U3420 ( .A1(n3445), .A2(n3446), .ZN(n3450) );
  OR2_X1 U3421 ( .A1(n2242), .A2(n2355), .ZN(n3446) );
  OR2_X1 U3422 ( .A1(n3451), .A2(n3452), .ZN(n3445) );
  AND2_X1 U3423 ( .A1(n3442), .A2(n3441), .ZN(n3452) );
  AND2_X1 U3424 ( .A1(n3439), .A2(n3453), .ZN(n3451) );
  OR2_X1 U3425 ( .A1(n3441), .A2(n3442), .ZN(n3453) );
  OR2_X1 U3426 ( .A1(n2242), .A2(n2525), .ZN(n3442) );
  OR2_X1 U3427 ( .A1(n3454), .A2(n3455), .ZN(n3441) );
  AND2_X1 U3428 ( .A1(n3438), .A2(n3437), .ZN(n3455) );
  AND2_X1 U3429 ( .A1(n3435), .A2(n3456), .ZN(n3454) );
  OR2_X1 U3430 ( .A1(n3437), .A2(n3438), .ZN(n3456) );
  OR2_X1 U3431 ( .A1(n2242), .A2(n2520), .ZN(n3438) );
  OR2_X1 U3432 ( .A1(n3457), .A2(n3458), .ZN(n3437) );
  AND2_X1 U3433 ( .A1(n3434), .A2(n3433), .ZN(n3458) );
  AND2_X1 U3434 ( .A1(n3431), .A2(n3459), .ZN(n3457) );
  OR2_X1 U3435 ( .A1(n3433), .A2(n3434), .ZN(n3459) );
  OR2_X1 U3436 ( .A1(n2242), .A2(n2515), .ZN(n3434) );
  OR2_X1 U3437 ( .A1(n3460), .A2(n3461), .ZN(n3433) );
  AND2_X1 U3438 ( .A1(n3425), .A2(n3428), .ZN(n3461) );
  AND2_X1 U3439 ( .A1(n3462), .A2(n3427), .ZN(n3460) );
  OR2_X1 U3440 ( .A1(n3463), .A2(n3464), .ZN(n3427) );
  AND2_X1 U3441 ( .A1(n3424), .A2(n3423), .ZN(n3464) );
  AND2_X1 U3442 ( .A1(n3421), .A2(n3465), .ZN(n3463) );
  OR2_X1 U3443 ( .A1(n3423), .A2(n3424), .ZN(n3465) );
  OR2_X1 U3444 ( .A1(n2242), .A2(n2505), .ZN(n3424) );
  OR2_X1 U3445 ( .A1(n3466), .A2(n3467), .ZN(n3423) );
  AND2_X1 U3446 ( .A1(n3418), .A2(n3419), .ZN(n3467) );
  AND2_X1 U3447 ( .A1(n3468), .A2(n3420), .ZN(n3466) );
  OR2_X1 U3448 ( .A1(n3469), .A2(n3470), .ZN(n3420) );
  AND2_X1 U3449 ( .A1(n3414), .A2(n3415), .ZN(n3470) );
  AND2_X1 U3450 ( .A1(n3471), .A2(n3416), .ZN(n3469) );
  OR2_X1 U3451 ( .A1(n3472), .A2(n3473), .ZN(n3416) );
  AND2_X1 U3452 ( .A1(n3410), .A2(n3412), .ZN(n3473) );
  AND2_X1 U3453 ( .A1(n3474), .A2(n3411), .ZN(n3472) );
  OR2_X1 U3454 ( .A1(n3475), .A2(n3476), .ZN(n3411) );
  AND2_X1 U3455 ( .A1(n3406), .A2(n3408), .ZN(n3476) );
  AND2_X1 U3456 ( .A1(n3477), .A2(n3478), .ZN(n3475) );
  OR2_X1 U3457 ( .A1(n3408), .A2(n3406), .ZN(n3478) );
  OR2_X1 U3458 ( .A1(n2242), .A2(n2480), .ZN(n3406) );
  OR2_X1 U3459 ( .A1(n2481), .A2(n3479), .ZN(n3408) );
  OR2_X1 U3460 ( .A1(n2216), .A2(n2242), .ZN(n3479) );
  INV_X1 U3461 ( .A(n3407), .ZN(n3477) );
  OR2_X1 U3462 ( .A1(n3480), .A2(n3481), .ZN(n3407) );
  AND2_X1 U3463 ( .A1(n3482), .A2(n3483), .ZN(n3481) );
  OR2_X1 U3464 ( .A1(n3484), .A2(n2045), .ZN(n3483) );
  AND2_X1 U3465 ( .A1(n2216), .A2(n2039), .ZN(n3484) );
  AND2_X1 U3466 ( .A1(n3400), .A2(n3485), .ZN(n3480) );
  OR2_X1 U3467 ( .A1(n3486), .A2(n2049), .ZN(n3485) );
  AND2_X1 U3468 ( .A1(n2186), .A2(n2051), .ZN(n3486) );
  OR2_X1 U3469 ( .A1(n3412), .A2(n3410), .ZN(n3474) );
  XOR2_X1 U3470 ( .A(n3487), .B(n3488), .Z(n3410) );
  XNOR2_X1 U3471 ( .A(n3489), .B(n3490), .ZN(n3487) );
  OR2_X1 U3472 ( .A1(n2490), .A2(n2242), .ZN(n3412) );
  OR2_X1 U3473 ( .A1(n3415), .A2(n3414), .ZN(n3471) );
  XNOR2_X1 U3474 ( .A(n3491), .B(n3492), .ZN(n3414) );
  XNOR2_X1 U3475 ( .A(n3493), .B(n3494), .ZN(n3491) );
  OR2_X1 U3476 ( .A1(n2495), .A2(n2242), .ZN(n3415) );
  OR2_X1 U3477 ( .A1(n3419), .A2(n3418), .ZN(n3468) );
  XNOR2_X1 U3478 ( .A(n3495), .B(n3496), .ZN(n3418) );
  XNOR2_X1 U3479 ( .A(n3497), .B(n3498), .ZN(n3495) );
  OR2_X1 U3480 ( .A1(n2500), .A2(n2242), .ZN(n3419) );
  XOR2_X1 U3481 ( .A(n3499), .B(n3500), .Z(n3421) );
  XOR2_X1 U3482 ( .A(n3501), .B(n3502), .Z(n3500) );
  OR2_X1 U3483 ( .A1(n3428), .A2(n3425), .ZN(n3462) );
  XOR2_X1 U3484 ( .A(n3503), .B(n3504), .Z(n3425) );
  XOR2_X1 U3485 ( .A(n3505), .B(n3506), .Z(n3504) );
  OR2_X1 U3486 ( .A1(n2242), .A2(n2510), .ZN(n3428) );
  INV_X1 U3487 ( .A(n3311), .ZN(n2242) );
  XOR2_X1 U3488 ( .A(n3507), .B(n3508), .Z(n3311) );
  XNOR2_X1 U3489 ( .A(c_5_), .B(d_5_), .ZN(n3507) );
  XOR2_X1 U3490 ( .A(n3509), .B(n3510), .Z(n3431) );
  XOR2_X1 U3491 ( .A(n3511), .B(n3512), .Z(n3510) );
  XOR2_X1 U3492 ( .A(n3513), .B(n3514), .Z(n3435) );
  XOR2_X1 U3493 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR2_X1 U3494 ( .A(n3517), .B(n3518), .Z(n3439) );
  XOR2_X1 U3495 ( .A(n3519), .B(n3520), .Z(n3518) );
  XOR2_X1 U3496 ( .A(n3521), .B(n3522), .Z(n3443) );
  XOR2_X1 U3497 ( .A(n3523), .B(n3524), .Z(n3522) );
  XOR2_X1 U3498 ( .A(n2352), .B(n3525), .Z(n2345) );
  XOR2_X1 U3499 ( .A(n2351), .B(n2350), .Z(n3525) );
  OR2_X1 U3500 ( .A1(n2216), .A2(n2355), .ZN(n2350) );
  OR2_X1 U3501 ( .A1(n3526), .A2(n3527), .ZN(n2351) );
  AND2_X1 U3502 ( .A1(n3524), .A2(n3523), .ZN(n3527) );
  AND2_X1 U3503 ( .A1(n3521), .A2(n3528), .ZN(n3526) );
  OR2_X1 U3504 ( .A1(n3523), .A2(n3524), .ZN(n3528) );
  OR2_X1 U3505 ( .A1(n2216), .A2(n2525), .ZN(n3524) );
  OR2_X1 U3506 ( .A1(n3529), .A2(n3530), .ZN(n3523) );
  AND2_X1 U3507 ( .A1(n3520), .A2(n3519), .ZN(n3530) );
  AND2_X1 U3508 ( .A1(n3517), .A2(n3531), .ZN(n3529) );
  OR2_X1 U3509 ( .A1(n3519), .A2(n3520), .ZN(n3531) );
  OR2_X1 U3510 ( .A1(n2216), .A2(n2520), .ZN(n3520) );
  OR2_X1 U3511 ( .A1(n3532), .A2(n3533), .ZN(n3519) );
  AND2_X1 U3512 ( .A1(n3516), .A2(n3515), .ZN(n3533) );
  AND2_X1 U3513 ( .A1(n3513), .A2(n3534), .ZN(n3532) );
  OR2_X1 U3514 ( .A1(n3515), .A2(n3516), .ZN(n3534) );
  OR2_X1 U3515 ( .A1(n2216), .A2(n2515), .ZN(n3516) );
  OR2_X1 U3516 ( .A1(n3535), .A2(n3536), .ZN(n3515) );
  AND2_X1 U3517 ( .A1(n3512), .A2(n3511), .ZN(n3536) );
  AND2_X1 U3518 ( .A1(n3509), .A2(n3537), .ZN(n3535) );
  OR2_X1 U3519 ( .A1(n3511), .A2(n3512), .ZN(n3537) );
  OR2_X1 U3520 ( .A1(n2216), .A2(n2510), .ZN(n3512) );
  OR2_X1 U3521 ( .A1(n3538), .A2(n3539), .ZN(n3511) );
  AND2_X1 U3522 ( .A1(n3503), .A2(n3506), .ZN(n3539) );
  AND2_X1 U3523 ( .A1(n3540), .A2(n3505), .ZN(n3538) );
  OR2_X1 U3524 ( .A1(n3541), .A2(n3542), .ZN(n3505) );
  AND2_X1 U3525 ( .A1(n3502), .A2(n3501), .ZN(n3542) );
  AND2_X1 U3526 ( .A1(n3499), .A2(n3543), .ZN(n3541) );
  OR2_X1 U3527 ( .A1(n3501), .A2(n3502), .ZN(n3543) );
  OR2_X1 U3528 ( .A1(n2216), .A2(n2500), .ZN(n3502) );
  OR2_X1 U3529 ( .A1(n3544), .A2(n3545), .ZN(n3501) );
  AND2_X1 U3530 ( .A1(n3496), .A2(n3497), .ZN(n3545) );
  AND2_X1 U3531 ( .A1(n3546), .A2(n3498), .ZN(n3544) );
  OR2_X1 U3532 ( .A1(n3547), .A2(n3548), .ZN(n3498) );
  AND2_X1 U3533 ( .A1(n3492), .A2(n3494), .ZN(n3548) );
  AND2_X1 U3534 ( .A1(n3549), .A2(n3493), .ZN(n3547) );
  OR2_X1 U3535 ( .A1(n3550), .A2(n3551), .ZN(n3493) );
  AND2_X1 U3536 ( .A1(n3488), .A2(n3490), .ZN(n3551) );
  AND2_X1 U3537 ( .A1(n3552), .A2(n3553), .ZN(n3550) );
  OR2_X1 U3538 ( .A1(n3490), .A2(n3488), .ZN(n3553) );
  OR2_X1 U3539 ( .A1(n2216), .A2(n2480), .ZN(n3488) );
  OR2_X1 U3540 ( .A1(n2481), .A2(n3554), .ZN(n3490) );
  OR2_X1 U3541 ( .A1(n2186), .A2(n2216), .ZN(n3554) );
  INV_X1 U3542 ( .A(n3489), .ZN(n3552) );
  OR2_X1 U3543 ( .A1(n3555), .A2(n3556), .ZN(n3489) );
  AND2_X1 U3544 ( .A1(n3557), .A2(n3558), .ZN(n3556) );
  OR2_X1 U3545 ( .A1(n3559), .A2(n2045), .ZN(n3558) );
  AND2_X1 U3546 ( .A1(n2186), .A2(n2039), .ZN(n3559) );
  AND2_X1 U3547 ( .A1(n3482), .A2(n3560), .ZN(n3555) );
  OR2_X1 U3548 ( .A1(n3561), .A2(n2049), .ZN(n3560) );
  AND2_X1 U3549 ( .A1(n3562), .A2(n2051), .ZN(n3561) );
  OR2_X1 U3550 ( .A1(n3494), .A2(n3492), .ZN(n3549) );
  XOR2_X1 U3551 ( .A(n3563), .B(n3564), .Z(n3492) );
  XNOR2_X1 U3552 ( .A(n3565), .B(n3566), .ZN(n3563) );
  OR2_X1 U3553 ( .A1(n2490), .A2(n2216), .ZN(n3494) );
  OR2_X1 U3554 ( .A1(n3497), .A2(n3496), .ZN(n3546) );
  XOR2_X1 U3555 ( .A(n3567), .B(n3568), .Z(n3496) );
  XOR2_X1 U3556 ( .A(n3569), .B(n3570), .Z(n3568) );
  OR2_X1 U3557 ( .A1(n2495), .A2(n2216), .ZN(n3497) );
  XOR2_X1 U3558 ( .A(n3571), .B(n3572), .Z(n3499) );
  XOR2_X1 U3559 ( .A(n3573), .B(n3574), .Z(n3572) );
  OR2_X1 U3560 ( .A1(n3506), .A2(n3503), .ZN(n3540) );
  XOR2_X1 U3561 ( .A(n3575), .B(n3576), .Z(n3503) );
  XOR2_X1 U3562 ( .A(n3577), .B(n3578), .Z(n3576) );
  OR2_X1 U3563 ( .A1(n2216), .A2(n2505), .ZN(n3506) );
  INV_X1 U3564 ( .A(n3400), .ZN(n2216) );
  XOR2_X1 U3565 ( .A(n3579), .B(n3580), .Z(n3400) );
  XNOR2_X1 U3566 ( .A(c_4_), .B(d_4_), .ZN(n3579) );
  XOR2_X1 U3567 ( .A(n3581), .B(n3582), .Z(n3509) );
  XOR2_X1 U3568 ( .A(n3583), .B(n3584), .Z(n3582) );
  XOR2_X1 U3569 ( .A(n3585), .B(n3586), .Z(n3513) );
  XOR2_X1 U3570 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR2_X1 U3571 ( .A(n3589), .B(n3590), .Z(n3517) );
  XOR2_X1 U3572 ( .A(n3591), .B(n3592), .Z(n3590) );
  XOR2_X1 U3573 ( .A(n3593), .B(n3594), .Z(n3521) );
  XOR2_X1 U3574 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR2_X1 U3575 ( .A(n2360), .B(n3597), .Z(n2352) );
  XOR2_X1 U3576 ( .A(n2359), .B(n2358), .Z(n3597) );
  OR2_X1 U3577 ( .A1(n2186), .A2(n2525), .ZN(n2358) );
  OR2_X1 U3578 ( .A1(n3598), .A2(n3599), .ZN(n2359) );
  AND2_X1 U3579 ( .A1(n3596), .A2(n3595), .ZN(n3599) );
  AND2_X1 U3580 ( .A1(n3593), .A2(n3600), .ZN(n3598) );
  OR2_X1 U3581 ( .A1(n3595), .A2(n3596), .ZN(n3600) );
  OR2_X1 U3582 ( .A1(n2186), .A2(n2520), .ZN(n3596) );
  OR2_X1 U3583 ( .A1(n3601), .A2(n3602), .ZN(n3595) );
  AND2_X1 U3584 ( .A1(n3592), .A2(n3591), .ZN(n3602) );
  AND2_X1 U3585 ( .A1(n3589), .A2(n3603), .ZN(n3601) );
  OR2_X1 U3586 ( .A1(n3591), .A2(n3592), .ZN(n3603) );
  OR2_X1 U3587 ( .A1(n2186), .A2(n2515), .ZN(n3592) );
  OR2_X1 U3588 ( .A1(n3604), .A2(n3605), .ZN(n3591) );
  AND2_X1 U3589 ( .A1(n3588), .A2(n3587), .ZN(n3605) );
  AND2_X1 U3590 ( .A1(n3585), .A2(n3606), .ZN(n3604) );
  OR2_X1 U3591 ( .A1(n3587), .A2(n3588), .ZN(n3606) );
  OR2_X1 U3592 ( .A1(n2186), .A2(n2510), .ZN(n3588) );
  OR2_X1 U3593 ( .A1(n3607), .A2(n3608), .ZN(n3587) );
  AND2_X1 U3594 ( .A1(n3584), .A2(n3583), .ZN(n3608) );
  AND2_X1 U3595 ( .A1(n3581), .A2(n3609), .ZN(n3607) );
  OR2_X1 U3596 ( .A1(n3583), .A2(n3584), .ZN(n3609) );
  OR2_X1 U3597 ( .A1(n2186), .A2(n2505), .ZN(n3584) );
  OR2_X1 U3598 ( .A1(n3610), .A2(n3611), .ZN(n3583) );
  AND2_X1 U3599 ( .A1(n3575), .A2(n3578), .ZN(n3611) );
  AND2_X1 U3600 ( .A1(n3612), .A2(n3577), .ZN(n3610) );
  OR2_X1 U3601 ( .A1(n3613), .A2(n3614), .ZN(n3577) );
  AND2_X1 U3602 ( .A1(n3574), .A2(n3573), .ZN(n3614) );
  AND2_X1 U3603 ( .A1(n3571), .A2(n3615), .ZN(n3613) );
  OR2_X1 U3604 ( .A1(n3573), .A2(n3574), .ZN(n3615) );
  OR2_X1 U3605 ( .A1(n2186), .A2(n2495), .ZN(n3574) );
  OR2_X1 U3606 ( .A1(n3616), .A2(n3617), .ZN(n3573) );
  AND2_X1 U3607 ( .A1(n3567), .A2(n3570), .ZN(n3617) );
  AND2_X1 U3608 ( .A1(n3618), .A2(n3569), .ZN(n3616) );
  OR2_X1 U3609 ( .A1(n3619), .A2(n3620), .ZN(n3569) );
  AND2_X1 U3610 ( .A1(n3564), .A2(n3566), .ZN(n3620) );
  AND2_X1 U3611 ( .A1(n3621), .A2(n3622), .ZN(n3619) );
  OR2_X1 U3612 ( .A1(n3566), .A2(n3564), .ZN(n3622) );
  OR2_X1 U3613 ( .A1(n2186), .A2(n2480), .ZN(n3564) );
  OR2_X1 U3614 ( .A1(n2481), .A2(n3623), .ZN(n3566) );
  OR2_X1 U3615 ( .A1(n3562), .A2(n2186), .ZN(n3623) );
  INV_X1 U3616 ( .A(n3565), .ZN(n3621) );
  OR2_X1 U3617 ( .A1(n3624), .A2(n3625), .ZN(n3565) );
  AND2_X1 U3618 ( .A1(n3626), .A2(n3627), .ZN(n3625) );
  OR2_X1 U3619 ( .A1(n3628), .A2(n2045), .ZN(n3627) );
  AND2_X1 U3620 ( .A1(n3562), .A2(n2039), .ZN(n3628) );
  AND2_X1 U3621 ( .A1(n3557), .A2(n3629), .ZN(n3624) );
  OR2_X1 U3622 ( .A1(n3630), .A2(n2049), .ZN(n3629) );
  AND2_X1 U3623 ( .A1(n3631), .A2(n2051), .ZN(n3630) );
  OR2_X1 U3624 ( .A1(n3570), .A2(n3567), .ZN(n3618) );
  XOR2_X1 U3625 ( .A(n3632), .B(n3633), .Z(n3567) );
  XNOR2_X1 U3626 ( .A(n3634), .B(n3635), .ZN(n3632) );
  OR2_X1 U3627 ( .A1(n2490), .A2(n2186), .ZN(n3570) );
  XNOR2_X1 U3628 ( .A(n3636), .B(n3637), .ZN(n3571) );
  XNOR2_X1 U3629 ( .A(n3638), .B(n3639), .ZN(n3636) );
  OR2_X1 U3630 ( .A1(n3578), .A2(n3575), .ZN(n3612) );
  XOR2_X1 U3631 ( .A(n3640), .B(n3641), .Z(n3575) );
  XOR2_X1 U3632 ( .A(n3642), .B(n3643), .Z(n3641) );
  OR2_X1 U3633 ( .A1(n2186), .A2(n2500), .ZN(n3578) );
  INV_X1 U3634 ( .A(n3482), .ZN(n2186) );
  XOR2_X1 U3635 ( .A(n3644), .B(n3645), .Z(n3482) );
  XNOR2_X1 U3636 ( .A(c_3_), .B(d_3_), .ZN(n3644) );
  XOR2_X1 U3637 ( .A(n3646), .B(n3647), .Z(n3581) );
  XOR2_X1 U3638 ( .A(n3648), .B(n3649), .Z(n3647) );
  XOR2_X1 U3639 ( .A(n3650), .B(n3651), .Z(n3585) );
  XOR2_X1 U3640 ( .A(n3652), .B(n3653), .Z(n3651) );
  XOR2_X1 U3641 ( .A(n3654), .B(n3655), .Z(n3589) );
  XOR2_X1 U3642 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR2_X1 U3643 ( .A(n3658), .B(n3659), .Z(n3593) );
  XOR2_X1 U3644 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR2_X1 U3645 ( .A(n3662), .B(n3663), .Z(n2360) );
  XOR2_X1 U3646 ( .A(n3664), .B(n3665), .Z(n3663) );
  AND2_X1 U3647 ( .A1(n2100), .A2(n3666), .ZN(n2102) );
  AND2_X1 U3648 ( .A1(n2101), .A2(n2099), .ZN(n3666) );
  XOR2_X1 U3649 ( .A(n3667), .B(n3668), .Z(n2099) );
  OR2_X1 U3650 ( .A1(n2187), .A2(n3669), .ZN(n3667) );
  XNOR2_X1 U3651 ( .A(n3670), .B(n3671), .ZN(n2101) );
  XOR2_X1 U3652 ( .A(n3672), .B(n3673), .Z(n3671) );
  INV_X1 U3653 ( .A(n2157), .ZN(n2100) );
  OR2_X1 U3654 ( .A1(n3674), .A2(n3675), .ZN(n2157) );
  AND2_X1 U3655 ( .A1(n2178), .A2(n2177), .ZN(n3675) );
  AND2_X1 U3656 ( .A1(n2175), .A2(n3676), .ZN(n3674) );
  OR2_X1 U3657 ( .A1(n2177), .A2(n2178), .ZN(n3676) );
  OR2_X1 U3658 ( .A1(n3562), .A2(n2187), .ZN(n2178) );
  OR2_X1 U3659 ( .A1(n3677), .A2(n3678), .ZN(n2177) );
  AND2_X1 U3660 ( .A1(n2197), .A2(n2196), .ZN(n3678) );
  AND2_X1 U3661 ( .A1(n2194), .A2(n3679), .ZN(n3677) );
  OR2_X1 U3662 ( .A1(n2196), .A2(n2197), .ZN(n3679) );
  OR2_X1 U3663 ( .A1(n3562), .A2(n2224), .ZN(n2197) );
  OR2_X1 U3664 ( .A1(n3680), .A2(n3681), .ZN(n2196) );
  AND2_X1 U3665 ( .A1(n2234), .A2(n2233), .ZN(n3681) );
  AND2_X1 U3666 ( .A1(n2231), .A2(n3682), .ZN(n3680) );
  OR2_X1 U3667 ( .A1(n2233), .A2(n2234), .ZN(n3682) );
  OR2_X1 U3668 ( .A1(n3562), .A2(n2257), .ZN(n2234) );
  OR2_X1 U3669 ( .A1(n3683), .A2(n3684), .ZN(n2233) );
  AND2_X1 U3670 ( .A1(n2267), .A2(n2266), .ZN(n3684) );
  AND2_X1 U3671 ( .A1(n2264), .A2(n3685), .ZN(n3683) );
  OR2_X1 U3672 ( .A1(n2266), .A2(n2267), .ZN(n3685) );
  OR2_X1 U3673 ( .A1(n3562), .A2(n2308), .ZN(n2267) );
  OR2_X1 U3674 ( .A1(n3686), .A2(n3687), .ZN(n2266) );
  AND2_X1 U3675 ( .A1(n2318), .A2(n2317), .ZN(n3687) );
  AND2_X1 U3676 ( .A1(n2315), .A2(n3688), .ZN(n3686) );
  OR2_X1 U3677 ( .A1(n2317), .A2(n2318), .ZN(n3688) );
  OR2_X1 U3678 ( .A1(n3562), .A2(n2355), .ZN(n2318) );
  OR2_X1 U3679 ( .A1(n3689), .A2(n3690), .ZN(n2317) );
  AND2_X1 U3680 ( .A1(n2365), .A2(n2364), .ZN(n3690) );
  AND2_X1 U3681 ( .A1(n2362), .A2(n3691), .ZN(n3689) );
  OR2_X1 U3682 ( .A1(n2364), .A2(n2365), .ZN(n3691) );
  OR2_X1 U3683 ( .A1(n3562), .A2(n2525), .ZN(n2365) );
  OR2_X1 U3684 ( .A1(n3692), .A2(n3693), .ZN(n2364) );
  AND2_X1 U3685 ( .A1(n3665), .A2(n3664), .ZN(n3693) );
  AND2_X1 U3686 ( .A1(n3662), .A2(n3694), .ZN(n3692) );
  OR2_X1 U3687 ( .A1(n3664), .A2(n3665), .ZN(n3694) );
  OR2_X1 U3688 ( .A1(n3562), .A2(n2520), .ZN(n3665) );
  OR2_X1 U3689 ( .A1(n3695), .A2(n3696), .ZN(n3664) );
  AND2_X1 U3690 ( .A1(n3661), .A2(n3660), .ZN(n3696) );
  AND2_X1 U3691 ( .A1(n3658), .A2(n3697), .ZN(n3695) );
  OR2_X1 U3692 ( .A1(n3660), .A2(n3661), .ZN(n3697) );
  OR2_X1 U3693 ( .A1(n3562), .A2(n2515), .ZN(n3661) );
  OR2_X1 U3694 ( .A1(n3698), .A2(n3699), .ZN(n3660) );
  AND2_X1 U3695 ( .A1(n3657), .A2(n3656), .ZN(n3699) );
  AND2_X1 U3696 ( .A1(n3654), .A2(n3700), .ZN(n3698) );
  OR2_X1 U3697 ( .A1(n3656), .A2(n3657), .ZN(n3700) );
  OR2_X1 U3698 ( .A1(n3562), .A2(n2510), .ZN(n3657) );
  OR2_X1 U3699 ( .A1(n3701), .A2(n3702), .ZN(n3656) );
  AND2_X1 U3700 ( .A1(n3653), .A2(n3652), .ZN(n3702) );
  AND2_X1 U3701 ( .A1(n3650), .A2(n3703), .ZN(n3701) );
  OR2_X1 U3702 ( .A1(n3652), .A2(n3653), .ZN(n3703) );
  OR2_X1 U3703 ( .A1(n3562), .A2(n2505), .ZN(n3653) );
  OR2_X1 U3704 ( .A1(n3704), .A2(n3705), .ZN(n3652) );
  AND2_X1 U3705 ( .A1(n3649), .A2(n3648), .ZN(n3705) );
  AND2_X1 U3706 ( .A1(n3646), .A2(n3706), .ZN(n3704) );
  OR2_X1 U3707 ( .A1(n3648), .A2(n3649), .ZN(n3706) );
  OR2_X1 U3708 ( .A1(n3562), .A2(n2500), .ZN(n3649) );
  OR2_X1 U3709 ( .A1(n3707), .A2(n3708), .ZN(n3648) );
  AND2_X1 U3710 ( .A1(n3640), .A2(n3643), .ZN(n3708) );
  AND2_X1 U3711 ( .A1(n3709), .A2(n3642), .ZN(n3707) );
  OR2_X1 U3712 ( .A1(n3710), .A2(n3711), .ZN(n3642) );
  AND2_X1 U3713 ( .A1(n3639), .A2(n3638), .ZN(n3711) );
  AND2_X1 U3714 ( .A1(n3637), .A2(n3712), .ZN(n3710) );
  OR2_X1 U3715 ( .A1(n3638), .A2(n3639), .ZN(n3712) );
  OR2_X1 U3716 ( .A1(n3562), .A2(n2490), .ZN(n3639) );
  OR2_X1 U3717 ( .A1(n3713), .A2(n3714), .ZN(n3638) );
  AND2_X1 U3718 ( .A1(n3633), .A2(n3635), .ZN(n3714) );
  AND2_X1 U3719 ( .A1(n3715), .A2(n3716), .ZN(n3713) );
  OR2_X1 U3720 ( .A1(n3635), .A2(n3633), .ZN(n3716) );
  OR2_X1 U3721 ( .A1(n3562), .A2(n2480), .ZN(n3633) );
  OR2_X1 U3722 ( .A1(n2481), .A2(n3717), .ZN(n3635) );
  OR2_X1 U3723 ( .A1(n3631), .A2(n3562), .ZN(n3717) );
  INV_X1 U3724 ( .A(n3634), .ZN(n3715) );
  OR2_X1 U3725 ( .A1(n3718), .A2(n3719), .ZN(n3634) );
  AND2_X1 U3726 ( .A1(n3720), .A2(n3721), .ZN(n3719) );
  OR2_X1 U3727 ( .A1(n3722), .A2(n2045), .ZN(n3721) );
  AND2_X1 U3728 ( .A1(n2039), .A2(n3723), .ZN(n2045) );
  AND2_X1 U3729 ( .A1(n3631), .A2(n2039), .ZN(n3722) );
  INV_X1 U3730 ( .A(n3669), .ZN(n3720) );
  AND2_X1 U3731 ( .A1(n3626), .A2(n3724), .ZN(n3718) );
  OR2_X1 U3732 ( .A1(n3725), .A2(n2049), .ZN(n3724) );
  AND2_X1 U3733 ( .A1(n3726), .A2(n2051), .ZN(n2049) );
  AND2_X1 U3734 ( .A1(n3669), .A2(n2051), .ZN(n3725) );
  INV_X1 U3735 ( .A(n3723), .ZN(n2051) );
  XNOR2_X1 U3736 ( .A(n3727), .B(n3728), .ZN(n3637) );
  OR2_X1 U3737 ( .A1(n3729), .A2(n3730), .ZN(n3727) );
  INV_X1 U3738 ( .A(n3731), .ZN(n3730) );
  AND2_X1 U3739 ( .A1(n3732), .A2(n3733), .ZN(n3729) );
  OR2_X1 U3740 ( .A1(n3643), .A2(n3640), .ZN(n3709) );
  XNOR2_X1 U3741 ( .A(n3734), .B(n3735), .ZN(n3640) );
  XNOR2_X1 U3742 ( .A(n3736), .B(n3737), .ZN(n3735) );
  OR2_X1 U3743 ( .A1(n3562), .A2(n2495), .ZN(n3643) );
  INV_X1 U3744 ( .A(n3557), .ZN(n3562) );
  XOR2_X1 U3745 ( .A(n3738), .B(n3739), .Z(n3557) );
  XNOR2_X1 U3746 ( .A(c_2_), .B(d_2_), .ZN(n3738) );
  XNOR2_X1 U3747 ( .A(n3740), .B(n3741), .ZN(n3646) );
  XNOR2_X1 U3748 ( .A(n3742), .B(n3743), .ZN(n3740) );
  XNOR2_X1 U3749 ( .A(n3744), .B(n3745), .ZN(n3650) );
  XNOR2_X1 U3750 ( .A(n3746), .B(n3747), .ZN(n3744) );
  XNOR2_X1 U3751 ( .A(n3748), .B(n3749), .ZN(n3654) );
  XNOR2_X1 U3752 ( .A(n3750), .B(n3751), .ZN(n3748) );
  XOR2_X1 U3753 ( .A(n3752), .B(n3753), .Z(n3658) );
  XOR2_X1 U3754 ( .A(n3754), .B(n3755), .Z(n3753) );
  XOR2_X1 U3755 ( .A(n3756), .B(n3757), .Z(n3662) );
  XOR2_X1 U3756 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR2_X1 U3757 ( .A(n3760), .B(n3761), .Z(n2362) );
  XOR2_X1 U3758 ( .A(n3762), .B(n3763), .Z(n3761) );
  XOR2_X1 U3759 ( .A(n3764), .B(n3765), .Z(n2315) );
  XOR2_X1 U3760 ( .A(n3766), .B(n3767), .Z(n3765) );
  XOR2_X1 U3761 ( .A(n3768), .B(n3769), .Z(n2264) );
  XOR2_X1 U3762 ( .A(n3770), .B(n3771), .Z(n3769) );
  XOR2_X1 U3763 ( .A(n3772), .B(n3773), .Z(n2231) );
  XOR2_X1 U3764 ( .A(n3774), .B(n3775), .Z(n3773) );
  XOR2_X1 U3765 ( .A(n3776), .B(n3777), .Z(n2194) );
  XOR2_X1 U3766 ( .A(n3778), .B(n3779), .Z(n3777) );
  XOR2_X1 U3767 ( .A(n3780), .B(n3781), .Z(n2175) );
  XOR2_X1 U3768 ( .A(n3782), .B(n3783), .Z(n3781) );
  INV_X1 U3769 ( .A(n3784), .ZN(n2154) );
  OR2_X1 U3770 ( .A1(n3668), .A2(n2187), .ZN(n3784) );
  OR2_X1 U3771 ( .A1(n3785), .A2(n3786), .ZN(n3668) );
  AND2_X1 U3772 ( .A1(n3670), .A2(n3672), .ZN(n3786) );
  AND2_X1 U3773 ( .A1(n3787), .A2(n3673), .ZN(n3785) );
  OR2_X1 U3774 ( .A1(n2224), .A2(n3669), .ZN(n3673) );
  OR2_X1 U3775 ( .A1(n3672), .A2(n3670), .ZN(n3787) );
  OR2_X1 U3776 ( .A1(n3631), .A2(n2187), .ZN(n3670) );
  XOR2_X1 U3777 ( .A(b_0_), .B(a_0_), .Z(n3789) );
  OR2_X1 U3778 ( .A1(n3790), .A2(n3791), .ZN(n3788) );
  AND2_X1 U3779 ( .A1(n3792), .A2(a_1_), .ZN(n3791) );
  AND2_X1 U3780 ( .A1(b_1_), .A2(n3793), .ZN(n3790) );
  OR2_X1 U3781 ( .A1(n3792), .A2(a_1_), .ZN(n3793) );
  INV_X1 U3782 ( .A(n3794), .ZN(n3792) );
  OR2_X1 U3783 ( .A1(n3795), .A2(n3796), .ZN(n3672) );
  AND2_X1 U3784 ( .A1(n3780), .A2(n3782), .ZN(n3796) );
  AND2_X1 U3785 ( .A1(n3797), .A2(n3783), .ZN(n3795) );
  OR2_X1 U3786 ( .A1(n3631), .A2(n2224), .ZN(n3783) );
  XNOR2_X1 U3787 ( .A(n3798), .B(n3794), .ZN(n2224) );
  OR2_X1 U3788 ( .A1(n3799), .A2(n3800), .ZN(n3794) );
  AND2_X1 U3789 ( .A1(n3801), .A2(n3802), .ZN(n3800) );
  AND2_X1 U3790 ( .A1(n3803), .A2(n3804), .ZN(n3799) );
  INV_X1 U3791 ( .A(b_2_), .ZN(n3804) );
  OR2_X1 U3792 ( .A1(n3802), .A2(n3801), .ZN(n3803) );
  INV_X1 U3793 ( .A(a_2_), .ZN(n3802) );
  XNOR2_X1 U3794 ( .A(a_1_), .B(b_1_), .ZN(n3798) );
  OR2_X1 U3795 ( .A1(n3782), .A2(n3780), .ZN(n3797) );
  OR2_X1 U3796 ( .A1(n2257), .A2(n3669), .ZN(n3780) );
  OR2_X1 U3797 ( .A1(n3805), .A2(n3806), .ZN(n3782) );
  AND2_X1 U3798 ( .A1(n3776), .A2(n3778), .ZN(n3806) );
  AND2_X1 U3799 ( .A1(n3807), .A2(n3779), .ZN(n3805) );
  OR2_X1 U3800 ( .A1(n2308), .A2(n3669), .ZN(n3779) );
  OR2_X1 U3801 ( .A1(n3778), .A2(n3776), .ZN(n3807) );
  OR2_X1 U3802 ( .A1(n3631), .A2(n2257), .ZN(n3776) );
  XNOR2_X1 U3803 ( .A(n3808), .B(n3801), .ZN(n2257) );
  OR2_X1 U3804 ( .A1(n3809), .A2(n3810), .ZN(n3801) );
  AND2_X1 U3805 ( .A1(n3811), .A2(n3812), .ZN(n3810) );
  AND2_X1 U3806 ( .A1(n3813), .A2(n3814), .ZN(n3809) );
  INV_X1 U3807 ( .A(b_3_), .ZN(n3814) );
  OR2_X1 U3808 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  INV_X1 U3809 ( .A(a_3_), .ZN(n3812) );
  XNOR2_X1 U3810 ( .A(a_2_), .B(b_2_), .ZN(n3808) );
  OR2_X1 U3811 ( .A1(n3815), .A2(n3816), .ZN(n3778) );
  AND2_X1 U3812 ( .A1(n3772), .A2(n3774), .ZN(n3816) );
  AND2_X1 U3813 ( .A1(n3817), .A2(n3775), .ZN(n3815) );
  OR2_X1 U3814 ( .A1(n2355), .A2(n3669), .ZN(n3775) );
  OR2_X1 U3815 ( .A1(n3774), .A2(n3772), .ZN(n3817) );
  OR2_X1 U3816 ( .A1(n3631), .A2(n2308), .ZN(n3772) );
  XNOR2_X1 U3817 ( .A(n3818), .B(n3811), .ZN(n2308) );
  OR2_X1 U3818 ( .A1(n3819), .A2(n3820), .ZN(n3811) );
  AND2_X1 U3819 ( .A1(n3821), .A2(n3822), .ZN(n3820) );
  AND2_X1 U3820 ( .A1(n3823), .A2(n3824), .ZN(n3819) );
  INV_X1 U3821 ( .A(b_4_), .ZN(n3824) );
  OR2_X1 U3822 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  INV_X1 U3823 ( .A(a_4_), .ZN(n3822) );
  XNOR2_X1 U3824 ( .A(a_3_), .B(b_3_), .ZN(n3818) );
  OR2_X1 U3825 ( .A1(n3825), .A2(n3826), .ZN(n3774) );
  AND2_X1 U3826 ( .A1(n3768), .A2(n3770), .ZN(n3826) );
  AND2_X1 U3827 ( .A1(n3827), .A2(n3771), .ZN(n3825) );
  OR2_X1 U3828 ( .A1(n2525), .A2(n3669), .ZN(n3771) );
  OR2_X1 U3829 ( .A1(n3770), .A2(n3768), .ZN(n3827) );
  OR2_X1 U3830 ( .A1(n3631), .A2(n2355), .ZN(n3768) );
  XNOR2_X1 U3831 ( .A(n3828), .B(n3821), .ZN(n2355) );
  OR2_X1 U3832 ( .A1(n3829), .A2(n3830), .ZN(n3821) );
  AND2_X1 U3833 ( .A1(n3831), .A2(n3832), .ZN(n3830) );
  AND2_X1 U3834 ( .A1(n3833), .A2(n3834), .ZN(n3829) );
  INV_X1 U3835 ( .A(b_5_), .ZN(n3834) );
  OR2_X1 U3836 ( .A1(n3832), .A2(n3831), .ZN(n3833) );
  INV_X1 U3837 ( .A(a_5_), .ZN(n3832) );
  XNOR2_X1 U3838 ( .A(a_4_), .B(b_4_), .ZN(n3828) );
  OR2_X1 U3839 ( .A1(n3835), .A2(n3836), .ZN(n3770) );
  AND2_X1 U3840 ( .A1(n3764), .A2(n3766), .ZN(n3836) );
  AND2_X1 U3841 ( .A1(n3837), .A2(n3767), .ZN(n3835) );
  OR2_X1 U3842 ( .A1(n2520), .A2(n3669), .ZN(n3767) );
  OR2_X1 U3843 ( .A1(n3766), .A2(n3764), .ZN(n3837) );
  OR2_X1 U3844 ( .A1(n3631), .A2(n2525), .ZN(n3764) );
  XNOR2_X1 U3845 ( .A(n3838), .B(n3831), .ZN(n2525) );
  OR2_X1 U3846 ( .A1(n3839), .A2(n3840), .ZN(n3831) );
  AND2_X1 U3847 ( .A1(n3841), .A2(n3842), .ZN(n3840) );
  AND2_X1 U3848 ( .A1(n3843), .A2(n3844), .ZN(n3839) );
  INV_X1 U3849 ( .A(b_6_), .ZN(n3844) );
  OR2_X1 U3850 ( .A1(n3842), .A2(n3841), .ZN(n3843) );
  INV_X1 U3851 ( .A(a_6_), .ZN(n3842) );
  XNOR2_X1 U3852 ( .A(a_5_), .B(b_5_), .ZN(n3838) );
  OR2_X1 U3853 ( .A1(n3845), .A2(n3846), .ZN(n3766) );
  AND2_X1 U3854 ( .A1(n3760), .A2(n3762), .ZN(n3846) );
  AND2_X1 U3855 ( .A1(n3847), .A2(n3763), .ZN(n3845) );
  OR2_X1 U3856 ( .A1(n2515), .A2(n3669), .ZN(n3763) );
  OR2_X1 U3857 ( .A1(n3762), .A2(n3760), .ZN(n3847) );
  OR2_X1 U3858 ( .A1(n3631), .A2(n2520), .ZN(n3760) );
  XNOR2_X1 U3859 ( .A(n3848), .B(n3841), .ZN(n2520) );
  OR2_X1 U3860 ( .A1(n3849), .A2(n3850), .ZN(n3841) );
  AND2_X1 U3861 ( .A1(n3851), .A2(n3852), .ZN(n3850) );
  AND2_X1 U3862 ( .A1(n3853), .A2(n3854), .ZN(n3849) );
  INV_X1 U3863 ( .A(b_7_), .ZN(n3854) );
  OR2_X1 U3864 ( .A1(n3852), .A2(n3851), .ZN(n3853) );
  INV_X1 U3865 ( .A(a_7_), .ZN(n3852) );
  XNOR2_X1 U3866 ( .A(a_6_), .B(b_6_), .ZN(n3848) );
  OR2_X1 U3867 ( .A1(n3855), .A2(n3856), .ZN(n3762) );
  AND2_X1 U3868 ( .A1(n3756), .A2(n3758), .ZN(n3856) );
  AND2_X1 U3869 ( .A1(n3857), .A2(n3759), .ZN(n3855) );
  OR2_X1 U3870 ( .A1(n2510), .A2(n3669), .ZN(n3759) );
  OR2_X1 U3871 ( .A1(n3758), .A2(n3756), .ZN(n3857) );
  OR2_X1 U3872 ( .A1(n3631), .A2(n2515), .ZN(n3756) );
  XNOR2_X1 U3873 ( .A(n3858), .B(n3851), .ZN(n2515) );
  OR2_X1 U3874 ( .A1(n3859), .A2(n3860), .ZN(n3851) );
  AND2_X1 U3875 ( .A1(n3861), .A2(n3862), .ZN(n3860) );
  AND2_X1 U3876 ( .A1(n3863), .A2(n3864), .ZN(n3859) );
  INV_X1 U3877 ( .A(b_8_), .ZN(n3864) );
  OR2_X1 U3878 ( .A1(n3862), .A2(n3861), .ZN(n3863) );
  INV_X1 U3879 ( .A(a_8_), .ZN(n3862) );
  XNOR2_X1 U3880 ( .A(a_7_), .B(b_7_), .ZN(n3858) );
  OR2_X1 U3881 ( .A1(n3865), .A2(n3866), .ZN(n3758) );
  AND2_X1 U3882 ( .A1(n3752), .A2(n3754), .ZN(n3866) );
  AND2_X1 U3883 ( .A1(n3867), .A2(n3755), .ZN(n3865) );
  OR2_X1 U3884 ( .A1(n2505), .A2(n3669), .ZN(n3755) );
  OR2_X1 U3885 ( .A1(n3754), .A2(n3752), .ZN(n3867) );
  OR2_X1 U3886 ( .A1(n3631), .A2(n2510), .ZN(n3752) );
  XNOR2_X1 U3887 ( .A(n3868), .B(n3861), .ZN(n2510) );
  OR2_X1 U3888 ( .A1(n3869), .A2(n3870), .ZN(n3861) );
  AND2_X1 U3889 ( .A1(n3871), .A2(n3872), .ZN(n3870) );
  AND2_X1 U3890 ( .A1(n3873), .A2(n3874), .ZN(n3869) );
  INV_X1 U3891 ( .A(b_9_), .ZN(n3874) );
  OR2_X1 U3892 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  INV_X1 U3893 ( .A(a_9_), .ZN(n3872) );
  XNOR2_X1 U3894 ( .A(a_8_), .B(b_8_), .ZN(n3868) );
  OR2_X1 U3895 ( .A1(n3875), .A2(n3876), .ZN(n3754) );
  AND2_X1 U3896 ( .A1(n3749), .A2(n3751), .ZN(n3876) );
  AND2_X1 U3897 ( .A1(n3877), .A2(n3750), .ZN(n3875) );
  OR2_X1 U3898 ( .A1(n2500), .A2(n3669), .ZN(n3750) );
  OR2_X1 U3899 ( .A1(n3751), .A2(n3749), .ZN(n3877) );
  OR2_X1 U3900 ( .A1(n3631), .A2(n2505), .ZN(n3749) );
  XNOR2_X1 U3901 ( .A(n3878), .B(n3871), .ZN(n2505) );
  OR2_X1 U3902 ( .A1(n3879), .A2(n3880), .ZN(n3871) );
  AND2_X1 U3903 ( .A1(n3881), .A2(n3882), .ZN(n3880) );
  AND2_X1 U3904 ( .A1(n3883), .A2(n3884), .ZN(n3879) );
  INV_X1 U3905 ( .A(b_10_), .ZN(n3884) );
  OR2_X1 U3906 ( .A1(n3882), .A2(n3881), .ZN(n3883) );
  INV_X1 U3907 ( .A(a_10_), .ZN(n3882) );
  XNOR2_X1 U3908 ( .A(a_9_), .B(b_9_), .ZN(n3878) );
  OR2_X1 U3909 ( .A1(n3885), .A2(n3886), .ZN(n3751) );
  AND2_X1 U3910 ( .A1(n3745), .A2(n3747), .ZN(n3886) );
  AND2_X1 U3911 ( .A1(n3887), .A2(n3746), .ZN(n3885) );
  OR2_X1 U3912 ( .A1(n2495), .A2(n3669), .ZN(n3746) );
  OR2_X1 U3913 ( .A1(n3747), .A2(n3745), .ZN(n3887) );
  OR2_X1 U3914 ( .A1(n3631), .A2(n2500), .ZN(n3745) );
  XNOR2_X1 U3915 ( .A(n3888), .B(n3881), .ZN(n2500) );
  OR2_X1 U3916 ( .A1(n3889), .A2(n3890), .ZN(n3881) );
  AND2_X1 U3917 ( .A1(n3891), .A2(n3892), .ZN(n3890) );
  AND2_X1 U3918 ( .A1(n3893), .A2(n3894), .ZN(n3889) );
  INV_X1 U3919 ( .A(b_11_), .ZN(n3894) );
  OR2_X1 U3920 ( .A1(n3892), .A2(n3891), .ZN(n3893) );
  INV_X1 U3921 ( .A(a_11_), .ZN(n3892) );
  XNOR2_X1 U3922 ( .A(a_10_), .B(b_10_), .ZN(n3888) );
  OR2_X1 U3923 ( .A1(n3895), .A2(n3896), .ZN(n3747) );
  AND2_X1 U3924 ( .A1(n3741), .A2(n3743), .ZN(n3896) );
  AND2_X1 U3925 ( .A1(n3897), .A2(n3742), .ZN(n3895) );
  OR2_X1 U3926 ( .A1(n2490), .A2(n3669), .ZN(n3742) );
  OR2_X1 U3927 ( .A1(n3743), .A2(n3741), .ZN(n3897) );
  OR2_X1 U3928 ( .A1(n3631), .A2(n2495), .ZN(n3741) );
  XNOR2_X1 U3929 ( .A(n3898), .B(n3891), .ZN(n2495) );
  OR2_X1 U3930 ( .A1(n3899), .A2(n3900), .ZN(n3891) );
  AND2_X1 U3931 ( .A1(n3901), .A2(n3902), .ZN(n3900) );
  AND2_X1 U3932 ( .A1(n3903), .A2(n3904), .ZN(n3899) );
  INV_X1 U3933 ( .A(b_12_), .ZN(n3904) );
  OR2_X1 U3934 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  INV_X1 U3935 ( .A(a_12_), .ZN(n3902) );
  XNOR2_X1 U3936 ( .A(a_11_), .B(b_11_), .ZN(n3898) );
  OR2_X1 U3937 ( .A1(n3905), .A2(n3906), .ZN(n3743) );
  AND2_X1 U3938 ( .A1(n3734), .A2(n3737), .ZN(n3906) );
  AND2_X1 U3939 ( .A1(n3736), .A2(n3907), .ZN(n3905) );
  OR2_X1 U3940 ( .A1(n3737), .A2(n3734), .ZN(n3907) );
  OR2_X1 U3941 ( .A1(n3631), .A2(n2490), .ZN(n3734) );
  XNOR2_X1 U3942 ( .A(n3908), .B(n3901), .ZN(n2490) );
  OR2_X1 U3943 ( .A1(n3909), .A2(n3910), .ZN(n3901) );
  AND2_X1 U3944 ( .A1(n3911), .A2(n3912), .ZN(n3910) );
  AND2_X1 U3945 ( .A1(n3913), .A2(n3914), .ZN(n3909) );
  OR2_X1 U3946 ( .A1(n3911), .A2(n3912), .ZN(n3913) );
  INV_X1 U3947 ( .A(a_13_), .ZN(n3912) );
  INV_X1 U3948 ( .A(n3915), .ZN(n3911) );
  XNOR2_X1 U3949 ( .A(a_12_), .B(b_12_), .ZN(n3908) );
  OR2_X1 U3950 ( .A1(n2480), .A2(n3669), .ZN(n3737) );
  AND2_X1 U3951 ( .A1(n3731), .A2(n3728), .ZN(n3736) );
  OR2_X1 U3952 ( .A1(n3669), .A2(n3916), .ZN(n3728) );
  OR2_X1 U3953 ( .A1(n3631), .A2(n2481), .ZN(n3916) );
  OR2_X1 U3954 ( .A1(n3723), .A2(n3726), .ZN(n2481) );
  INV_X1 U3955 ( .A(n2039), .ZN(n3726) );
  AND2_X1 U3956 ( .A1(n3917), .A2(n3918), .ZN(n2039) );
  OR2_X1 U3957 ( .A1(b_15_), .A2(a_15_), .ZN(n3918) );
  OR2_X1 U3958 ( .A1(n3733), .A2(n3732), .ZN(n3731) );
  OR2_X1 U3959 ( .A1(n3723), .A2(n3669), .ZN(n3732) );
  XOR2_X1 U3960 ( .A(d_0_), .B(c_0_), .Z(n3920) );
  OR2_X1 U3961 ( .A1(n3921), .A2(n3922), .ZN(n3919) );
  AND2_X1 U3962 ( .A1(n3923), .A2(c_1_), .ZN(n3922) );
  AND2_X1 U3963 ( .A1(d_1_), .A2(n3924), .ZN(n3921) );
  OR2_X1 U3964 ( .A1(n3923), .A2(c_1_), .ZN(n3924) );
  INV_X1 U3965 ( .A(n3925), .ZN(n3923) );
  XOR2_X1 U3966 ( .A(n3917), .B(n3926), .Z(n3723) );
  XOR2_X1 U3967 ( .A(b_14_), .B(a_14_), .Z(n3926) );
  INV_X1 U3968 ( .A(n3927), .ZN(n3917) );
  OR2_X1 U3969 ( .A1(n3631), .A2(n2480), .ZN(n3733) );
  XNOR2_X1 U3970 ( .A(n3915), .B(n3928), .ZN(n2480) );
  XNOR2_X1 U3971 ( .A(n3914), .B(a_13_), .ZN(n3928) );
  INV_X1 U3972 ( .A(b_13_), .ZN(n3914) );
  OR2_X1 U3973 ( .A1(n3929), .A2(n3930), .ZN(n3915) );
  AND2_X1 U3974 ( .A1(n3927), .A2(a_14_), .ZN(n3930) );
  AND2_X1 U3975 ( .A1(b_14_), .A2(n3931), .ZN(n3929) );
  OR2_X1 U3976 ( .A1(n3927), .A2(a_14_), .ZN(n3931) );
  AND2_X1 U3977 ( .A1(a_15_), .A2(b_15_), .ZN(n3927) );
  INV_X1 U3978 ( .A(n3626), .ZN(n3631) );
  XOR2_X1 U3979 ( .A(n3932), .B(n3925), .Z(n3626) );
  OR2_X1 U3980 ( .A1(n3933), .A2(n3934), .ZN(n3925) );
  AND2_X1 U3981 ( .A1(n3739), .A2(n3935), .ZN(n3934) );
  AND2_X1 U3982 ( .A1(n3936), .A2(n3937), .ZN(n3933) );
  INV_X1 U3983 ( .A(d_2_), .ZN(n3937) );
  OR2_X1 U3984 ( .A1(n3935), .A2(n3739), .ZN(n3936) );
  OR2_X1 U3985 ( .A1(n3938), .A2(n3939), .ZN(n3739) );
  AND2_X1 U3986 ( .A1(n3645), .A2(n3940), .ZN(n3939) );
  AND2_X1 U3987 ( .A1(n3941), .A2(n3942), .ZN(n3938) );
  INV_X1 U3988 ( .A(d_3_), .ZN(n3942) );
  OR2_X1 U3989 ( .A1(n3940), .A2(n3645), .ZN(n3941) );
  OR2_X1 U3990 ( .A1(n3943), .A2(n3944), .ZN(n3645) );
  AND2_X1 U3991 ( .A1(n3580), .A2(n3945), .ZN(n3944) );
  AND2_X1 U3992 ( .A1(n3946), .A2(n3947), .ZN(n3943) );
  INV_X1 U3993 ( .A(d_4_), .ZN(n3947) );
  OR2_X1 U3994 ( .A1(n3945), .A2(n3580), .ZN(n3946) );
  OR2_X1 U3995 ( .A1(n3948), .A2(n3949), .ZN(n3580) );
  AND2_X1 U3996 ( .A1(n3508), .A2(n3950), .ZN(n3949) );
  AND2_X1 U3997 ( .A1(n3951), .A2(n3952), .ZN(n3948) );
  INV_X1 U3998 ( .A(d_5_), .ZN(n3952) );
  OR2_X1 U3999 ( .A1(n3950), .A2(n3508), .ZN(n3951) );
  OR2_X1 U4000 ( .A1(n3953), .A2(n3954), .ZN(n3508) );
  AND2_X1 U4001 ( .A1(n3430), .A2(n3955), .ZN(n3954) );
  AND2_X1 U4002 ( .A1(n3956), .A2(n3957), .ZN(n3953) );
  INV_X1 U4003 ( .A(d_6_), .ZN(n3957) );
  OR2_X1 U4004 ( .A1(n3955), .A2(n3430), .ZN(n3956) );
  OR2_X1 U4005 ( .A1(n3958), .A2(n3959), .ZN(n3430) );
  AND2_X1 U4006 ( .A1(n3345), .A2(n3960), .ZN(n3959) );
  AND2_X1 U4007 ( .A1(n3961), .A2(n3962), .ZN(n3958) );
  INV_X1 U4008 ( .A(d_7_), .ZN(n3962) );
  OR2_X1 U4009 ( .A1(n3960), .A2(n3345), .ZN(n3961) );
  OR2_X1 U4010 ( .A1(n3963), .A2(n3964), .ZN(n3345) );
  AND2_X1 U4011 ( .A1(n3253), .A2(n3965), .ZN(n3964) );
  AND2_X1 U4012 ( .A1(n3966), .A2(n3967), .ZN(n3963) );
  INV_X1 U4013 ( .A(d_8_), .ZN(n3967) );
  OR2_X1 U4014 ( .A1(n3965), .A2(n3253), .ZN(n3966) );
  OR2_X1 U4015 ( .A1(n3968), .A2(n3969), .ZN(n3253) );
  AND2_X1 U4016 ( .A1(n3154), .A2(n3970), .ZN(n3969) );
  AND2_X1 U4017 ( .A1(n3971), .A2(n3972), .ZN(n3968) );
  INV_X1 U4018 ( .A(d_9_), .ZN(n3972) );
  OR2_X1 U4019 ( .A1(n3970), .A2(n3154), .ZN(n3971) );
  OR2_X1 U4020 ( .A1(n3973), .A2(n3974), .ZN(n3154) );
  AND2_X1 U4021 ( .A1(n3045), .A2(n3975), .ZN(n3974) );
  AND2_X1 U4022 ( .A1(n3976), .A2(n3977), .ZN(n3973) );
  INV_X1 U4023 ( .A(d_10_), .ZN(n3977) );
  OR2_X1 U4024 ( .A1(n3975), .A2(n3045), .ZN(n3976) );
  OR2_X1 U4025 ( .A1(n3978), .A2(n3979), .ZN(n3045) );
  AND2_X1 U4026 ( .A1(n2887), .A2(n3980), .ZN(n3979) );
  AND2_X1 U4027 ( .A1(n3981), .A2(n3982), .ZN(n3978) );
  INV_X1 U4028 ( .A(d_11_), .ZN(n3982) );
  OR2_X1 U4029 ( .A1(n3980), .A2(n2887), .ZN(n3981) );
  OR2_X1 U4030 ( .A1(n3983), .A2(n3984), .ZN(n2887) );
  AND2_X1 U4031 ( .A1(n2777), .A2(n3985), .ZN(n3984) );
  AND2_X1 U4032 ( .A1(n3986), .A2(n3987), .ZN(n3983) );
  INV_X1 U4033 ( .A(d_12_), .ZN(n3987) );
  OR2_X1 U4034 ( .A1(n3985), .A2(n2777), .ZN(n3986) );
  OR2_X1 U4035 ( .A1(n3988), .A2(n3989), .ZN(n2777) );
  AND2_X1 U4036 ( .A1(n2685), .A2(n3990), .ZN(n3989) );
  AND2_X1 U4037 ( .A1(n3991), .A2(n2687), .ZN(n3988) );
  INV_X1 U4038 ( .A(d_13_), .ZN(n2687) );
  OR2_X1 U4039 ( .A1(n2685), .A2(n3990), .ZN(n3991) );
  INV_X1 U4040 ( .A(c_13_), .ZN(n3990) );
  INV_X1 U4041 ( .A(n3992), .ZN(n2685) );
  OR2_X1 U4042 ( .A1(n3993), .A2(n3994), .ZN(n3992) );
  AND2_X1 U4043 ( .A1(c_14_), .A2(n2599), .ZN(n3994) );
  AND2_X1 U4044 ( .A1(d_14_), .A2(n3995), .ZN(n3993) );
  OR2_X1 U4045 ( .A1(n2599), .A2(c_14_), .ZN(n3995) );
  AND2_X1 U4046 ( .A1(c_15_), .A2(d_15_), .ZN(n2599) );
  INV_X1 U4047 ( .A(c_12_), .ZN(n3985) );
  INV_X1 U4048 ( .A(c_11_), .ZN(n3980) );
  INV_X1 U4049 ( .A(c_10_), .ZN(n3975) );
  INV_X1 U4050 ( .A(c_9_), .ZN(n3970) );
  INV_X1 U4051 ( .A(c_8_), .ZN(n3965) );
  INV_X1 U4052 ( .A(c_7_), .ZN(n3960) );
  INV_X1 U4053 ( .A(c_6_), .ZN(n3955) );
  INV_X1 U4054 ( .A(c_5_), .ZN(n3950) );
  INV_X1 U4055 ( .A(c_4_), .ZN(n3945) );
  INV_X1 U4056 ( .A(c_3_), .ZN(n3940) );
  INV_X1 U4057 ( .A(c_2_), .ZN(n3935) );
  XNOR2_X1 U4058 ( .A(c_1_), .B(d_1_), .ZN(n3932) );
endmodule

