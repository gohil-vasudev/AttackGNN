module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n543_, new_n113_, new_n924_, new_n886_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n914_, new_n938_, new_n259_, new_n362_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n126_, new_n810_, new_n940_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n904_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_2 );
not g001 ( new_n107_, N37 );
and g002 ( new_n108_, new_n107_, N33 );
not g003 ( new_n109_, N33 );
and g004 ( new_n110_, new_n109_, N37 );
or g005 ( new_n111_, new_n108_, new_n110_ );
not g006 ( new_n112_, N41 );
or g007 ( new_n113_, new_n112_, N45 );
not g008 ( new_n114_, N45 );
or g009 ( new_n115_, new_n114_, N41 );
and g010 ( new_n116_, new_n113_, new_n115_ );
and g011 ( new_n117_, new_n111_, new_n116_ );
or g012 ( new_n118_, new_n109_, N37 );
or g013 ( new_n119_, new_n107_, N33 );
and g014 ( new_n120_, new_n118_, new_n119_ );
and g015 ( new_n121_, new_n114_, N41 );
and g016 ( new_n122_, new_n112_, N45 );
or g017 ( new_n123_, new_n121_, new_n122_ );
and g018 ( new_n124_, new_n123_, new_n120_ );
or g019 ( new_n125_, new_n117_, new_n124_ );
and g020 ( new_n126_, new_n125_, new_n106_ );
or g021 ( new_n127_, new_n123_, new_n120_ );
or g022 ( new_n128_, new_n111_, new_n116_ );
and g023 ( new_n129_, new_n127_, new_n128_ );
and g024 ( new_n130_, new_n129_, keyIn_0_2 );
or g025 ( new_n131_, new_n126_, new_n130_ );
not g026 ( new_n132_, keyIn_0_0 );
not g027 ( new_n133_, N5 );
and g028 ( new_n134_, new_n133_, N1 );
not g029 ( new_n135_, N1 );
and g030 ( new_n136_, new_n135_, N5 );
or g031 ( new_n137_, new_n134_, new_n136_ );
not g032 ( new_n138_, N9 );
or g033 ( new_n139_, new_n138_, N13 );
not g034 ( new_n140_, N13 );
or g035 ( new_n141_, new_n140_, N9 );
and g036 ( new_n142_, new_n139_, new_n141_ );
and g037 ( new_n143_, new_n137_, new_n142_ );
or g038 ( new_n144_, new_n135_, N5 );
or g039 ( new_n145_, new_n133_, N1 );
and g040 ( new_n146_, new_n144_, new_n145_ );
and g041 ( new_n147_, new_n140_, N9 );
and g042 ( new_n148_, new_n138_, N13 );
or g043 ( new_n149_, new_n147_, new_n148_ );
and g044 ( new_n150_, new_n149_, new_n146_ );
or g045 ( new_n151_, new_n143_, new_n150_ );
or g046 ( new_n152_, new_n151_, new_n132_ );
or g047 ( new_n153_, new_n149_, new_n146_ );
or g048 ( new_n154_, new_n137_, new_n142_ );
and g049 ( new_n155_, new_n153_, new_n154_ );
or g050 ( new_n156_, new_n155_, keyIn_0_0 );
and g051 ( new_n157_, new_n152_, new_n156_ );
and g052 ( new_n158_, new_n131_, new_n157_ );
or g053 ( new_n159_, new_n129_, keyIn_0_2 );
or g054 ( new_n160_, new_n125_, new_n106_ );
and g055 ( new_n161_, new_n160_, new_n159_ );
and g056 ( new_n162_, new_n155_, keyIn_0_0 );
and g057 ( new_n163_, new_n151_, new_n132_ );
or g058 ( new_n164_, new_n163_, new_n162_ );
and g059 ( new_n165_, new_n164_, new_n161_ );
or g060 ( new_n166_, new_n158_, new_n165_ );
and g061 ( new_n167_, new_n166_, keyIn_0_18 );
not g062 ( new_n168_, new_n167_ );
or g063 ( new_n169_, new_n166_, keyIn_0_18 );
and g064 ( new_n170_, new_n168_, new_n169_ );
and g065 ( new_n171_, N135, N137 );
not g066 ( new_n172_, new_n171_ );
and g067 ( new_n173_, new_n170_, new_n172_ );
or g068 ( new_n174_, new_n170_, new_n172_ );
not g069 ( new_n175_, new_n174_ );
or g070 ( new_n176_, new_n175_, new_n173_ );
and g071 ( new_n177_, new_n176_, keyIn_0_30 );
not g072 ( new_n178_, keyIn_0_30 );
not g073 ( new_n179_, new_n173_ );
and g074 ( new_n180_, new_n179_, new_n174_ );
and g075 ( new_n181_, new_n180_, new_n178_ );
or g076 ( new_n182_, new_n177_, new_n181_ );
not g077 ( new_n183_, keyIn_0_14 );
not g078 ( new_n184_, N89 );
and g079 ( new_n185_, new_n184_, N73 );
not g080 ( new_n186_, N73 );
and g081 ( new_n187_, new_n186_, N89 );
or g082 ( new_n188_, new_n185_, new_n187_ );
not g083 ( new_n189_, N121 );
and g084 ( new_n190_, new_n189_, N105 );
not g085 ( new_n191_, N105 );
and g086 ( new_n192_, new_n191_, N121 );
or g087 ( new_n193_, new_n190_, new_n192_ );
not g088 ( new_n194_, new_n193_ );
and g089 ( new_n195_, new_n194_, new_n188_ );
not g090 ( new_n196_, new_n195_ );
or g091 ( new_n197_, new_n194_, new_n188_ );
and g092 ( new_n198_, new_n196_, new_n197_ );
not g093 ( new_n199_, new_n198_ );
and g094 ( new_n200_, new_n199_, new_n183_ );
and g095 ( new_n201_, new_n198_, keyIn_0_14 );
or g096 ( new_n202_, new_n200_, new_n201_ );
and g097 ( new_n203_, new_n182_, new_n202_ );
or g098 ( new_n204_, new_n180_, new_n178_ );
not g099 ( new_n205_, new_n181_ );
and g100 ( new_n206_, new_n205_, new_n204_ );
not g101 ( new_n207_, new_n202_ );
and g102 ( new_n208_, new_n206_, new_n207_ );
or g103 ( new_n209_, new_n208_, new_n203_ );
not g104 ( new_n210_, keyIn_0_15 );
not g105 ( new_n211_, N93 );
and g106 ( new_n212_, new_n211_, N77 );
not g107 ( new_n213_, N77 );
and g108 ( new_n214_, new_n213_, N93 );
or g109 ( new_n215_, new_n212_, new_n214_ );
not g110 ( new_n216_, N125 );
and g111 ( new_n217_, new_n216_, N109 );
not g112 ( new_n218_, N109 );
and g113 ( new_n219_, new_n218_, N125 );
or g114 ( new_n220_, new_n217_, new_n219_ );
not g115 ( new_n221_, new_n220_ );
and g116 ( new_n222_, new_n221_, new_n215_ );
not g117 ( new_n223_, new_n222_ );
or g118 ( new_n224_, new_n221_, new_n215_ );
and g119 ( new_n225_, new_n223_, new_n224_ );
not g120 ( new_n226_, new_n225_ );
and g121 ( new_n227_, new_n226_, new_n210_ );
and g122 ( new_n228_, new_n225_, keyIn_0_15 );
or g123 ( new_n229_, new_n227_, new_n228_ );
not g124 ( new_n230_, new_n229_ );
not g125 ( new_n231_, N53 );
and g126 ( new_n232_, new_n231_, N49 );
not g127 ( new_n233_, N49 );
and g128 ( new_n234_, new_n233_, N53 );
or g129 ( new_n235_, new_n232_, new_n234_ );
not g130 ( new_n236_, N57 );
or g131 ( new_n237_, new_n236_, N61 );
not g132 ( new_n238_, N61 );
or g133 ( new_n239_, new_n238_, N57 );
and g134 ( new_n240_, new_n237_, new_n239_ );
and g135 ( new_n241_, new_n235_, new_n240_ );
or g136 ( new_n242_, new_n233_, N53 );
or g137 ( new_n243_, new_n231_, N49 );
and g138 ( new_n244_, new_n242_, new_n243_ );
and g139 ( new_n245_, new_n238_, N57 );
and g140 ( new_n246_, new_n236_, N61 );
or g141 ( new_n247_, new_n245_, new_n246_ );
and g142 ( new_n248_, new_n247_, new_n244_ );
or g143 ( new_n249_, new_n241_, new_n248_ );
or g144 ( new_n250_, new_n249_, keyIn_0_3 );
not g145 ( new_n251_, keyIn_0_3 );
or g146 ( new_n252_, new_n247_, new_n244_ );
or g147 ( new_n253_, new_n235_, new_n240_ );
and g148 ( new_n254_, new_n252_, new_n253_ );
or g149 ( new_n255_, new_n254_, new_n251_ );
and g150 ( new_n256_, new_n250_, new_n255_ );
not g151 ( new_n257_, keyIn_0_1 );
not g152 ( new_n258_, N21 );
and g153 ( new_n259_, new_n258_, N17 );
not g154 ( new_n260_, N17 );
and g155 ( new_n261_, new_n260_, N21 );
or g156 ( new_n262_, new_n259_, new_n261_ );
not g157 ( new_n263_, N25 );
or g158 ( new_n264_, new_n263_, N29 );
not g159 ( new_n265_, N29 );
or g160 ( new_n266_, new_n265_, N25 );
and g161 ( new_n267_, new_n264_, new_n266_ );
and g162 ( new_n268_, new_n262_, new_n267_ );
or g163 ( new_n269_, new_n260_, N21 );
or g164 ( new_n270_, new_n258_, N17 );
and g165 ( new_n271_, new_n269_, new_n270_ );
and g166 ( new_n272_, new_n265_, N25 );
and g167 ( new_n273_, new_n263_, N29 );
or g168 ( new_n274_, new_n272_, new_n273_ );
and g169 ( new_n275_, new_n274_, new_n271_ );
or g170 ( new_n276_, new_n268_, new_n275_ );
and g171 ( new_n277_, new_n276_, new_n257_ );
or g172 ( new_n278_, new_n274_, new_n271_ );
or g173 ( new_n279_, new_n262_, new_n267_ );
and g174 ( new_n280_, new_n278_, new_n279_ );
and g175 ( new_n281_, new_n280_, keyIn_0_1 );
or g176 ( new_n282_, new_n277_, new_n281_ );
and g177 ( new_n283_, new_n282_, new_n256_ );
and g178 ( new_n284_, new_n254_, new_n251_ );
and g179 ( new_n285_, new_n249_, keyIn_0_3 );
or g180 ( new_n286_, new_n285_, new_n284_ );
or g181 ( new_n287_, new_n280_, keyIn_0_1 );
or g182 ( new_n288_, new_n276_, new_n257_ );
and g183 ( new_n289_, new_n288_, new_n287_ );
and g184 ( new_n290_, new_n286_, new_n289_ );
or g185 ( new_n291_, new_n283_, new_n290_ );
and g186 ( new_n292_, new_n291_, keyIn_0_19 );
not g187 ( new_n293_, new_n292_ );
or g188 ( new_n294_, new_n291_, keyIn_0_19 );
and g189 ( new_n295_, new_n293_, new_n294_ );
and g190 ( new_n296_, N136, N137 );
or g191 ( new_n297_, new_n295_, new_n296_ );
and g192 ( new_n298_, new_n295_, new_n296_ );
not g193 ( new_n299_, new_n298_ );
and g194 ( new_n300_, new_n299_, new_n297_ );
not g195 ( new_n301_, new_n300_ );
and g196 ( new_n302_, new_n301_, keyIn_0_31 );
not g197 ( new_n303_, keyIn_0_31 );
and g198 ( new_n304_, new_n300_, new_n303_ );
or g199 ( new_n305_, new_n302_, new_n304_ );
or g200 ( new_n306_, new_n305_, new_n230_ );
or g201 ( new_n307_, new_n300_, new_n303_ );
not g202 ( new_n308_, new_n304_ );
and g203 ( new_n309_, new_n308_, new_n307_ );
or g204 ( new_n310_, new_n309_, new_n229_ );
and g205 ( new_n311_, new_n306_, new_n310_ );
and g206 ( new_n312_, new_n311_, new_n209_ );
not g207 ( new_n313_, keyIn_0_29 );
not g208 ( new_n314_, keyIn_0_17 );
or g209 ( new_n315_, new_n161_, new_n256_ );
or g210 ( new_n316_, new_n131_, new_n286_ );
and g211 ( new_n317_, new_n316_, new_n315_ );
or g212 ( new_n318_, new_n317_, new_n314_ );
and g213 ( new_n319_, new_n131_, new_n286_ );
and g214 ( new_n320_, new_n161_, new_n256_ );
or g215 ( new_n321_, new_n319_, new_n320_ );
or g216 ( new_n322_, new_n321_, keyIn_0_17 );
and g217 ( new_n323_, new_n318_, new_n322_ );
and g218 ( new_n324_, N134, N137 );
or g219 ( new_n325_, new_n323_, new_n324_ );
and g220 ( new_n326_, new_n321_, keyIn_0_17 );
and g221 ( new_n327_, new_n317_, new_n314_ );
or g222 ( new_n328_, new_n327_, new_n326_ );
not g223 ( new_n329_, new_n324_ );
or g224 ( new_n330_, new_n328_, new_n329_ );
and g225 ( new_n331_, new_n330_, new_n325_ );
or g226 ( new_n332_, new_n331_, new_n313_ );
and g227 ( new_n333_, new_n328_, new_n329_ );
and g228 ( new_n334_, new_n323_, new_n324_ );
or g229 ( new_n335_, new_n333_, new_n334_ );
or g230 ( new_n336_, new_n335_, keyIn_0_29 );
and g231 ( new_n337_, new_n336_, new_n332_ );
not g232 ( new_n338_, N85 );
and g233 ( new_n339_, new_n338_, N69 );
not g234 ( new_n340_, N69 );
and g235 ( new_n341_, new_n340_, N85 );
or g236 ( new_n342_, new_n339_, new_n341_ );
not g237 ( new_n343_, N117 );
and g238 ( new_n344_, new_n343_, N101 );
not g239 ( new_n345_, N101 );
and g240 ( new_n346_, new_n345_, N117 );
or g241 ( new_n347_, new_n344_, new_n346_ );
not g242 ( new_n348_, new_n347_ );
and g243 ( new_n349_, new_n348_, new_n342_ );
not g244 ( new_n350_, new_n349_ );
or g245 ( new_n351_, new_n348_, new_n342_ );
and g246 ( new_n352_, new_n350_, new_n351_ );
not g247 ( new_n353_, new_n352_ );
and g248 ( new_n354_, new_n353_, keyIn_0_13 );
not g249 ( new_n355_, new_n354_ );
or g250 ( new_n356_, new_n353_, keyIn_0_13 );
and g251 ( new_n357_, new_n355_, new_n356_ );
or g252 ( new_n358_, new_n337_, new_n357_ );
and g253 ( new_n359_, new_n335_, keyIn_0_29 );
and g254 ( new_n360_, new_n331_, new_n313_ );
or g255 ( new_n361_, new_n359_, new_n360_ );
not g256 ( new_n362_, new_n357_ );
or g257 ( new_n363_, new_n361_, new_n362_ );
and g258 ( new_n364_, new_n363_, new_n358_ );
not g259 ( new_n365_, keyIn_0_16 );
and g260 ( new_n366_, new_n164_, new_n282_ );
and g261 ( new_n367_, new_n157_, new_n289_ );
or g262 ( new_n368_, new_n366_, new_n367_ );
and g263 ( new_n369_, new_n368_, new_n365_ );
or g264 ( new_n370_, new_n157_, new_n289_ );
or g265 ( new_n371_, new_n164_, new_n282_ );
and g266 ( new_n372_, new_n371_, new_n370_ );
and g267 ( new_n373_, new_n372_, keyIn_0_16 );
or g268 ( new_n374_, new_n373_, new_n369_ );
and g269 ( new_n375_, N133, N137 );
and g270 ( new_n376_, new_n374_, new_n375_ );
or g271 ( new_n377_, new_n372_, keyIn_0_16 );
or g272 ( new_n378_, new_n368_, new_n365_ );
and g273 ( new_n379_, new_n377_, new_n378_ );
not g274 ( new_n380_, new_n375_ );
and g275 ( new_n381_, new_n379_, new_n380_ );
or g276 ( new_n382_, new_n376_, new_n381_ );
and g277 ( new_n383_, new_n382_, keyIn_0_28 );
not g278 ( new_n384_, keyIn_0_28 );
or g279 ( new_n385_, new_n379_, new_n380_ );
or g280 ( new_n386_, new_n374_, new_n375_ );
and g281 ( new_n387_, new_n386_, new_n385_ );
and g282 ( new_n388_, new_n387_, new_n384_ );
or g283 ( new_n389_, new_n383_, new_n388_ );
not g284 ( new_n390_, N81 );
and g285 ( new_n391_, new_n390_, N65 );
not g286 ( new_n392_, N65 );
and g287 ( new_n393_, new_n392_, N81 );
or g288 ( new_n394_, new_n391_, new_n393_ );
not g289 ( new_n395_, N113 );
and g290 ( new_n396_, new_n395_, N97 );
not g291 ( new_n397_, N97 );
and g292 ( new_n398_, new_n397_, N113 );
or g293 ( new_n399_, new_n396_, new_n398_ );
not g294 ( new_n400_, new_n399_ );
and g295 ( new_n401_, new_n400_, new_n394_ );
not g296 ( new_n402_, new_n401_ );
or g297 ( new_n403_, new_n400_, new_n394_ );
and g298 ( new_n404_, new_n402_, new_n403_ );
not g299 ( new_n405_, new_n404_ );
and g300 ( new_n406_, new_n405_, keyIn_0_12 );
not g301 ( new_n407_, new_n406_ );
or g302 ( new_n408_, new_n405_, keyIn_0_12 );
and g303 ( new_n409_, new_n407_, new_n408_ );
and g304 ( new_n410_, new_n389_, new_n409_ );
or g305 ( new_n411_, new_n387_, new_n384_ );
or g306 ( new_n412_, new_n382_, keyIn_0_28 );
and g307 ( new_n413_, new_n412_, new_n411_ );
not g308 ( new_n414_, new_n409_ );
and g309 ( new_n415_, new_n413_, new_n414_ );
or g310 ( new_n416_, new_n410_, new_n415_ );
and g311 ( new_n417_, new_n416_, new_n364_ );
and g312 ( new_n418_, new_n312_, new_n417_ );
not g313 ( new_n419_, new_n418_ );
not g314 ( new_n420_, keyIn_0_24 );
not g315 ( new_n421_, keyIn_0_20 );
not g316 ( new_n422_, keyIn_0_4 );
and g317 ( new_n423_, new_n340_, N65 );
and g318 ( new_n424_, new_n392_, N69 );
or g319 ( new_n425_, new_n423_, new_n424_ );
or g320 ( new_n426_, new_n186_, N77 );
or g321 ( new_n427_, new_n213_, N73 );
and g322 ( new_n428_, new_n426_, new_n427_ );
and g323 ( new_n429_, new_n425_, new_n428_ );
or g324 ( new_n430_, new_n392_, N69 );
or g325 ( new_n431_, new_n340_, N65 );
and g326 ( new_n432_, new_n430_, new_n431_ );
and g327 ( new_n433_, new_n213_, N73 );
and g328 ( new_n434_, new_n186_, N77 );
or g329 ( new_n435_, new_n433_, new_n434_ );
and g330 ( new_n436_, new_n435_, new_n432_ );
or g331 ( new_n437_, new_n429_, new_n436_ );
and g332 ( new_n438_, new_n437_, new_n422_ );
or g333 ( new_n439_, new_n435_, new_n432_ );
or g334 ( new_n440_, new_n425_, new_n428_ );
and g335 ( new_n441_, new_n439_, new_n440_ );
and g336 ( new_n442_, new_n441_, keyIn_0_4 );
or g337 ( new_n443_, new_n438_, new_n442_ );
not g338 ( new_n444_, keyIn_0_5 );
or g339 ( new_n445_, new_n390_, N85 );
or g340 ( new_n446_, new_n338_, N81 );
and g341 ( new_n447_, new_n445_, new_n446_ );
and g342 ( new_n448_, new_n211_, N89 );
and g343 ( new_n449_, new_n184_, N93 );
or g344 ( new_n450_, new_n448_, new_n449_ );
or g345 ( new_n451_, new_n450_, new_n447_ );
and g346 ( new_n452_, new_n338_, N81 );
and g347 ( new_n453_, new_n390_, N85 );
or g348 ( new_n454_, new_n452_, new_n453_ );
or g349 ( new_n455_, new_n184_, N93 );
or g350 ( new_n456_, new_n211_, N89 );
and g351 ( new_n457_, new_n455_, new_n456_ );
or g352 ( new_n458_, new_n454_, new_n457_ );
and g353 ( new_n459_, new_n451_, new_n458_ );
or g354 ( new_n460_, new_n459_, new_n444_ );
and g355 ( new_n461_, new_n454_, new_n457_ );
and g356 ( new_n462_, new_n450_, new_n447_ );
or g357 ( new_n463_, new_n461_, new_n462_ );
or g358 ( new_n464_, new_n463_, keyIn_0_5 );
and g359 ( new_n465_, new_n464_, new_n460_ );
and g360 ( new_n466_, new_n443_, new_n465_ );
or g361 ( new_n467_, new_n441_, keyIn_0_4 );
or g362 ( new_n468_, new_n437_, new_n422_ );
and g363 ( new_n469_, new_n468_, new_n467_ );
and g364 ( new_n470_, new_n463_, keyIn_0_5 );
and g365 ( new_n471_, new_n459_, new_n444_ );
or g366 ( new_n472_, new_n470_, new_n471_ );
and g367 ( new_n473_, new_n472_, new_n469_ );
or g368 ( new_n474_, new_n466_, new_n473_ );
and g369 ( new_n475_, new_n474_, new_n421_ );
or g370 ( new_n476_, new_n472_, new_n469_ );
or g371 ( new_n477_, new_n443_, new_n465_ );
and g372 ( new_n478_, new_n476_, new_n477_ );
and g373 ( new_n479_, new_n478_, keyIn_0_20 );
or g374 ( new_n480_, new_n475_, new_n479_ );
and g375 ( new_n481_, N129, N137 );
or g376 ( new_n482_, new_n480_, new_n481_ );
or g377 ( new_n483_, new_n478_, keyIn_0_20 );
or g378 ( new_n484_, new_n474_, new_n421_ );
and g379 ( new_n485_, new_n484_, new_n483_ );
not g380 ( new_n486_, new_n481_ );
or g381 ( new_n487_, new_n485_, new_n486_ );
and g382 ( new_n488_, new_n482_, new_n487_ );
or g383 ( new_n489_, new_n488_, new_n420_ );
and g384 ( new_n490_, new_n485_, new_n486_ );
and g385 ( new_n491_, new_n480_, new_n481_ );
or g386 ( new_n492_, new_n491_, new_n490_ );
or g387 ( new_n493_, new_n492_, keyIn_0_24 );
and g388 ( new_n494_, new_n493_, new_n489_ );
not g389 ( new_n495_, keyIn_0_8 );
and g390 ( new_n496_, new_n260_, N1 );
and g391 ( new_n497_, new_n135_, N17 );
or g392 ( new_n498_, new_n496_, new_n497_ );
and g393 ( new_n499_, new_n233_, N33 );
and g394 ( new_n500_, new_n109_, N49 );
or g395 ( new_n501_, new_n499_, new_n500_ );
not g396 ( new_n502_, new_n501_ );
and g397 ( new_n503_, new_n502_, new_n498_ );
not g398 ( new_n504_, new_n503_ );
or g399 ( new_n505_, new_n502_, new_n498_ );
and g400 ( new_n506_, new_n504_, new_n505_ );
not g401 ( new_n507_, new_n506_ );
and g402 ( new_n508_, new_n507_, new_n495_ );
and g403 ( new_n509_, new_n506_, keyIn_0_8 );
or g404 ( new_n510_, new_n508_, new_n509_ );
not g405 ( new_n511_, new_n510_ );
or g406 ( new_n512_, new_n494_, new_n511_ );
and g407 ( new_n513_, new_n492_, keyIn_0_24 );
and g408 ( new_n514_, new_n488_, new_n420_ );
or g409 ( new_n515_, new_n513_, new_n514_ );
or g410 ( new_n516_, new_n515_, new_n510_ );
and g411 ( new_n517_, new_n516_, new_n512_ );
not g412 ( new_n518_, keyIn_0_22 );
and g413 ( new_n519_, new_n345_, N97 );
and g414 ( new_n520_, new_n397_, N101 );
or g415 ( new_n521_, new_n519_, new_n520_ );
or g416 ( new_n522_, new_n191_, N109 );
or g417 ( new_n523_, new_n218_, N105 );
and g418 ( new_n524_, new_n522_, new_n523_ );
and g419 ( new_n525_, new_n521_, new_n524_ );
or g420 ( new_n526_, new_n397_, N101 );
or g421 ( new_n527_, new_n345_, N97 );
and g422 ( new_n528_, new_n526_, new_n527_ );
and g423 ( new_n529_, new_n218_, N105 );
and g424 ( new_n530_, new_n191_, N109 );
or g425 ( new_n531_, new_n529_, new_n530_ );
and g426 ( new_n532_, new_n531_, new_n528_ );
or g427 ( new_n533_, new_n525_, new_n532_ );
and g428 ( new_n534_, new_n533_, keyIn_0_6 );
not g429 ( new_n535_, keyIn_0_6 );
or g430 ( new_n536_, new_n531_, new_n528_ );
or g431 ( new_n537_, new_n521_, new_n524_ );
and g432 ( new_n538_, new_n536_, new_n537_ );
and g433 ( new_n539_, new_n538_, new_n535_ );
or g434 ( new_n540_, new_n534_, new_n539_ );
and g435 ( new_n541_, new_n443_, new_n540_ );
or g436 ( new_n542_, new_n538_, new_n535_ );
or g437 ( new_n543_, new_n533_, keyIn_0_6 );
and g438 ( new_n544_, new_n543_, new_n542_ );
and g439 ( new_n545_, new_n469_, new_n544_ );
or g440 ( new_n546_, new_n541_, new_n545_ );
and g441 ( new_n547_, new_n546_, new_n518_ );
not g442 ( new_n548_, new_n547_ );
or g443 ( new_n549_, new_n546_, new_n518_ );
and g444 ( new_n550_, new_n548_, new_n549_ );
and g445 ( new_n551_, N131, N137 );
not g446 ( new_n552_, new_n551_ );
or g447 ( new_n553_, new_n550_, new_n552_ );
and g448 ( new_n554_, new_n550_, new_n552_ );
not g449 ( new_n555_, new_n554_ );
and g450 ( new_n556_, new_n555_, new_n553_ );
not g451 ( new_n557_, new_n556_ );
and g452 ( new_n558_, new_n557_, keyIn_0_26 );
not g453 ( new_n559_, keyIn_0_26 );
and g454 ( new_n560_, new_n556_, new_n559_ );
or g455 ( new_n561_, new_n558_, new_n560_ );
not g456 ( new_n562_, keyIn_0_10 );
and g457 ( new_n563_, new_n263_, N9 );
and g458 ( new_n564_, new_n138_, N25 );
or g459 ( new_n565_, new_n563_, new_n564_ );
and g460 ( new_n566_, new_n236_, N41 );
and g461 ( new_n567_, new_n112_, N57 );
or g462 ( new_n568_, new_n566_, new_n567_ );
not g463 ( new_n569_, new_n568_ );
and g464 ( new_n570_, new_n569_, new_n565_ );
not g465 ( new_n571_, new_n570_ );
or g466 ( new_n572_, new_n569_, new_n565_ );
and g467 ( new_n573_, new_n571_, new_n572_ );
not g468 ( new_n574_, new_n573_ );
and g469 ( new_n575_, new_n574_, new_n562_ );
and g470 ( new_n576_, new_n573_, keyIn_0_10 );
or g471 ( new_n577_, new_n575_, new_n576_ );
not g472 ( new_n578_, new_n577_ );
and g473 ( new_n579_, new_n561_, new_n578_ );
or g474 ( new_n580_, new_n556_, new_n559_ );
not g475 ( new_n581_, new_n560_ );
and g476 ( new_n582_, new_n581_, new_n580_ );
and g477 ( new_n583_, new_n582_, new_n577_ );
or g478 ( new_n584_, new_n579_, new_n583_ );
and g479 ( new_n585_, new_n515_, new_n510_ );
and g480 ( new_n586_, new_n494_, new_n511_ );
or g481 ( new_n587_, new_n585_, new_n586_ );
not g482 ( new_n588_, keyIn_0_21 );
or g483 ( new_n589_, new_n395_, N117 );
or g484 ( new_n590_, new_n343_, N113 );
and g485 ( new_n591_, new_n589_, new_n590_ );
and g486 ( new_n592_, new_n216_, N121 );
and g487 ( new_n593_, new_n189_, N125 );
or g488 ( new_n594_, new_n592_, new_n593_ );
or g489 ( new_n595_, new_n594_, new_n591_ );
and g490 ( new_n596_, new_n343_, N113 );
and g491 ( new_n597_, new_n395_, N117 );
or g492 ( new_n598_, new_n596_, new_n597_ );
or g493 ( new_n599_, new_n189_, N125 );
or g494 ( new_n600_, new_n216_, N121 );
and g495 ( new_n601_, new_n599_, new_n600_ );
or g496 ( new_n602_, new_n598_, new_n601_ );
and g497 ( new_n603_, new_n595_, new_n602_ );
or g498 ( new_n604_, new_n603_, keyIn_0_7 );
not g499 ( new_n605_, keyIn_0_7 );
and g500 ( new_n606_, new_n598_, new_n601_ );
and g501 ( new_n607_, new_n594_, new_n591_ );
or g502 ( new_n608_, new_n606_, new_n607_ );
or g503 ( new_n609_, new_n608_, new_n605_ );
and g504 ( new_n610_, new_n609_, new_n604_ );
or g505 ( new_n611_, new_n544_, new_n610_ );
and g506 ( new_n612_, new_n608_, new_n605_ );
and g507 ( new_n613_, new_n603_, keyIn_0_7 );
or g508 ( new_n614_, new_n612_, new_n613_ );
or g509 ( new_n615_, new_n540_, new_n614_ );
and g510 ( new_n616_, new_n615_, new_n611_ );
or g511 ( new_n617_, new_n616_, new_n588_ );
and g512 ( new_n618_, new_n540_, new_n614_ );
and g513 ( new_n619_, new_n544_, new_n610_ );
or g514 ( new_n620_, new_n618_, new_n619_ );
or g515 ( new_n621_, new_n620_, keyIn_0_21 );
and g516 ( new_n622_, new_n617_, new_n621_ );
and g517 ( new_n623_, N130, N137 );
or g518 ( new_n624_, new_n622_, new_n623_ );
and g519 ( new_n625_, new_n620_, keyIn_0_21 );
and g520 ( new_n626_, new_n616_, new_n588_ );
or g521 ( new_n627_, new_n626_, new_n625_ );
not g522 ( new_n628_, new_n623_ );
or g523 ( new_n629_, new_n627_, new_n628_ );
and g524 ( new_n630_, new_n629_, new_n624_ );
or g525 ( new_n631_, new_n630_, keyIn_0_25 );
not g526 ( new_n632_, keyIn_0_25 );
and g527 ( new_n633_, new_n627_, new_n628_ );
and g528 ( new_n634_, new_n622_, new_n623_ );
or g529 ( new_n635_, new_n633_, new_n634_ );
or g530 ( new_n636_, new_n635_, new_n632_ );
and g531 ( new_n637_, new_n636_, new_n631_ );
and g532 ( new_n638_, new_n258_, N5 );
and g533 ( new_n639_, new_n133_, N21 );
or g534 ( new_n640_, new_n638_, new_n639_ );
and g535 ( new_n641_, new_n231_, N37 );
and g536 ( new_n642_, new_n107_, N53 );
or g537 ( new_n643_, new_n641_, new_n642_ );
not g538 ( new_n644_, new_n643_ );
and g539 ( new_n645_, new_n644_, new_n640_ );
not g540 ( new_n646_, new_n645_ );
or g541 ( new_n647_, new_n644_, new_n640_ );
and g542 ( new_n648_, new_n646_, new_n647_ );
not g543 ( new_n649_, new_n648_ );
and g544 ( new_n650_, new_n649_, keyIn_0_9 );
not g545 ( new_n651_, new_n650_ );
or g546 ( new_n652_, new_n649_, keyIn_0_9 );
and g547 ( new_n653_, new_n651_, new_n652_ );
or g548 ( new_n654_, new_n637_, new_n653_ );
and g549 ( new_n655_, new_n635_, new_n632_ );
and g550 ( new_n656_, new_n630_, keyIn_0_25 );
or g551 ( new_n657_, new_n655_, new_n656_ );
not g552 ( new_n658_, new_n653_ );
or g553 ( new_n659_, new_n657_, new_n658_ );
and g554 ( new_n660_, new_n659_, new_n654_ );
or g555 ( new_n661_, new_n587_, new_n660_ );
or g556 ( new_n662_, new_n661_, new_n584_ );
and g557 ( new_n663_, new_n657_, new_n658_ );
and g558 ( new_n664_, new_n637_, new_n653_ );
or g559 ( new_n665_, new_n663_, new_n664_ );
or g560 ( new_n666_, new_n665_, new_n517_ );
or g561 ( new_n667_, new_n666_, new_n584_ );
and g562 ( new_n668_, new_n662_, new_n667_ );
not g563 ( new_n669_, keyIn_0_27 );
and g564 ( new_n670_, new_n614_, new_n465_ );
and g565 ( new_n671_, new_n472_, new_n610_ );
or g566 ( new_n672_, new_n670_, new_n671_ );
and g567 ( new_n673_, new_n672_, keyIn_0_23 );
not g568 ( new_n674_, new_n673_ );
or g569 ( new_n675_, new_n672_, keyIn_0_23 );
and g570 ( new_n676_, new_n674_, new_n675_ );
and g571 ( new_n677_, N132, N137 );
or g572 ( new_n678_, new_n676_, new_n677_ );
and g573 ( new_n679_, new_n676_, new_n677_ );
not g574 ( new_n680_, new_n679_ );
and g575 ( new_n681_, new_n680_, new_n678_ );
not g576 ( new_n682_, new_n681_ );
and g577 ( new_n683_, new_n682_, new_n669_ );
and g578 ( new_n684_, new_n681_, keyIn_0_27 );
or g579 ( new_n685_, new_n683_, new_n684_ );
and g580 ( new_n686_, new_n265_, N13 );
and g581 ( new_n687_, new_n140_, N29 );
or g582 ( new_n688_, new_n686_, new_n687_ );
and g583 ( new_n689_, new_n238_, N45 );
and g584 ( new_n690_, new_n114_, N61 );
or g585 ( new_n691_, new_n689_, new_n690_ );
not g586 ( new_n692_, new_n691_ );
and g587 ( new_n693_, new_n692_, new_n688_ );
not g588 ( new_n694_, new_n693_ );
or g589 ( new_n695_, new_n692_, new_n688_ );
and g590 ( new_n696_, new_n694_, new_n695_ );
not g591 ( new_n697_, new_n696_ );
and g592 ( new_n698_, new_n697_, keyIn_0_11 );
not g593 ( new_n699_, new_n698_ );
or g594 ( new_n700_, new_n697_, keyIn_0_11 );
and g595 ( new_n701_, new_n699_, new_n700_ );
and g596 ( new_n702_, new_n685_, new_n701_ );
or g597 ( new_n703_, new_n681_, keyIn_0_27 );
not g598 ( new_n704_, new_n684_ );
and g599 ( new_n705_, new_n704_, new_n703_ );
not g600 ( new_n706_, new_n701_ );
and g601 ( new_n707_, new_n705_, new_n706_ );
or g602 ( new_n708_, new_n702_, new_n707_ );
or g603 ( new_n709_, new_n668_, new_n708_ );
or g604 ( new_n710_, new_n705_, new_n706_ );
or g605 ( new_n711_, new_n685_, new_n701_ );
and g606 ( new_n712_, new_n711_, new_n710_ );
or g607 ( new_n713_, new_n712_, new_n584_ );
or g608 ( new_n714_, new_n582_, new_n577_ );
or g609 ( new_n715_, new_n561_, new_n578_ );
and g610 ( new_n716_, new_n715_, new_n714_ );
or g611 ( new_n717_, new_n708_, new_n716_ );
and g612 ( new_n718_, new_n713_, new_n717_ );
and g613 ( new_n719_, new_n517_, new_n660_ );
not g614 ( new_n720_, new_n719_ );
or g615 ( new_n721_, new_n718_, new_n720_ );
and g616 ( new_n722_, new_n709_, new_n721_ );
or g617 ( new_n723_, new_n722_, new_n517_ );
or g618 ( new_n724_, new_n723_, new_n419_ );
and g619 ( new_n725_, new_n724_, N1 );
and g620 ( new_n726_, new_n665_, new_n517_ );
and g621 ( new_n727_, new_n726_, new_n716_ );
and g622 ( new_n728_, new_n587_, new_n660_ );
and g623 ( new_n729_, new_n728_, new_n716_ );
or g624 ( new_n730_, new_n727_, new_n729_ );
and g625 ( new_n731_, new_n730_, new_n712_ );
and g626 ( new_n732_, new_n708_, new_n716_ );
and g627 ( new_n733_, new_n712_, new_n584_ );
or g628 ( new_n734_, new_n733_, new_n732_ );
and g629 ( new_n735_, new_n734_, new_n719_ );
or g630 ( new_n736_, new_n731_, new_n735_ );
and g631 ( new_n737_, new_n736_, new_n587_ );
and g632 ( new_n738_, new_n737_, new_n418_ );
and g633 ( new_n739_, new_n738_, new_n135_ );
or g634 ( N724, new_n725_, new_n739_ );
or g635 ( new_n741_, new_n722_, new_n660_ );
or g636 ( new_n742_, new_n741_, new_n419_ );
and g637 ( new_n743_, new_n742_, N5 );
and g638 ( new_n744_, new_n736_, new_n665_ );
and g639 ( new_n745_, new_n744_, new_n418_ );
and g640 ( new_n746_, new_n745_, new_n133_ );
or g641 ( N725, new_n743_, new_n746_ );
or g642 ( new_n748_, new_n722_, new_n716_ );
or g643 ( new_n749_, new_n748_, new_n419_ );
and g644 ( new_n750_, new_n749_, N9 );
and g645 ( new_n751_, new_n736_, new_n584_ );
and g646 ( new_n752_, new_n751_, new_n418_ );
and g647 ( new_n753_, new_n752_, new_n138_ );
or g648 ( N726, new_n750_, new_n753_ );
or g649 ( new_n755_, new_n722_, new_n712_ );
or g650 ( new_n756_, new_n755_, new_n419_ );
and g651 ( new_n757_, new_n756_, N13 );
and g652 ( new_n758_, new_n736_, new_n708_ );
and g653 ( new_n759_, new_n758_, new_n418_ );
and g654 ( new_n760_, new_n759_, new_n140_ );
or g655 ( N727, new_n757_, new_n760_ );
and g656 ( new_n762_, new_n309_, new_n229_ );
and g657 ( new_n763_, new_n305_, new_n230_ );
or g658 ( new_n764_, new_n763_, new_n762_ );
or g659 ( new_n765_, new_n206_, new_n207_ );
or g660 ( new_n766_, new_n182_, new_n202_ );
and g661 ( new_n767_, new_n765_, new_n766_ );
and g662 ( new_n768_, new_n417_, new_n767_ );
and g663 ( new_n769_, new_n768_, new_n764_ );
not g664 ( new_n770_, new_n769_ );
or g665 ( new_n771_, new_n723_, new_n770_ );
and g666 ( new_n772_, new_n771_, N17 );
and g667 ( new_n773_, new_n737_, new_n769_ );
and g668 ( new_n774_, new_n773_, new_n260_ );
or g669 ( N728, new_n772_, new_n774_ );
or g670 ( new_n776_, new_n741_, new_n770_ );
and g671 ( new_n777_, new_n776_, N21 );
and g672 ( new_n778_, new_n744_, new_n769_ );
and g673 ( new_n779_, new_n778_, new_n258_ );
or g674 ( N729, new_n777_, new_n779_ );
or g675 ( new_n781_, new_n748_, new_n770_ );
and g676 ( new_n782_, new_n781_, N25 );
and g677 ( new_n783_, new_n751_, new_n769_ );
and g678 ( new_n784_, new_n783_, new_n263_ );
or g679 ( N730, new_n782_, new_n784_ );
or g680 ( new_n786_, new_n755_, new_n770_ );
and g681 ( new_n787_, new_n786_, N29 );
and g682 ( new_n788_, new_n758_, new_n769_ );
and g683 ( new_n789_, new_n788_, new_n265_ );
or g684 ( N731, new_n787_, new_n789_ );
and g685 ( new_n791_, new_n361_, new_n362_ );
and g686 ( new_n792_, new_n337_, new_n357_ );
or g687 ( new_n793_, new_n791_, new_n792_ );
or g688 ( new_n794_, new_n413_, new_n414_ );
or g689 ( new_n795_, new_n389_, new_n409_ );
and g690 ( new_n796_, new_n795_, new_n794_ );
and g691 ( new_n797_, new_n793_, new_n796_ );
and g692 ( new_n798_, new_n312_, new_n797_ );
not g693 ( new_n799_, new_n798_ );
or g694 ( new_n800_, new_n723_, new_n799_ );
and g695 ( new_n801_, new_n800_, N33 );
and g696 ( new_n802_, new_n737_, new_n798_ );
and g697 ( new_n803_, new_n802_, new_n109_ );
or g698 ( N732, new_n801_, new_n803_ );
or g699 ( new_n805_, new_n741_, new_n799_ );
and g700 ( new_n806_, new_n805_, N37 );
and g701 ( new_n807_, new_n744_, new_n798_ );
and g702 ( new_n808_, new_n807_, new_n107_ );
or g703 ( N733, new_n806_, new_n808_ );
or g704 ( new_n810_, new_n748_, new_n799_ );
and g705 ( new_n811_, new_n810_, N41 );
and g706 ( new_n812_, new_n751_, new_n798_ );
and g707 ( new_n813_, new_n812_, new_n112_ );
or g708 ( N734, new_n811_, new_n813_ );
or g709 ( new_n815_, new_n755_, new_n799_ );
and g710 ( new_n816_, new_n815_, N45 );
and g711 ( new_n817_, new_n758_, new_n798_ );
and g712 ( new_n818_, new_n817_, new_n114_ );
or g713 ( N735, new_n816_, new_n818_ );
and g714 ( new_n820_, new_n797_, new_n767_ );
and g715 ( new_n821_, new_n820_, new_n764_ );
not g716 ( new_n822_, new_n821_ );
or g717 ( new_n823_, new_n723_, new_n822_ );
and g718 ( new_n824_, new_n823_, N49 );
and g719 ( new_n825_, new_n737_, new_n821_ );
and g720 ( new_n826_, new_n825_, new_n233_ );
or g721 ( N736, new_n824_, new_n826_ );
or g722 ( new_n828_, new_n741_, new_n822_ );
and g723 ( new_n829_, new_n828_, N53 );
and g724 ( new_n830_, new_n744_, new_n821_ );
and g725 ( new_n831_, new_n830_, new_n231_ );
or g726 ( N737, new_n829_, new_n831_ );
or g727 ( new_n833_, new_n748_, new_n822_ );
and g728 ( new_n834_, new_n833_, N57 );
and g729 ( new_n835_, new_n751_, new_n821_ );
and g730 ( new_n836_, new_n835_, new_n236_ );
or g731 ( N738, new_n834_, new_n836_ );
or g732 ( new_n838_, new_n755_, new_n822_ );
and g733 ( new_n839_, new_n838_, N61 );
and g734 ( new_n840_, new_n758_, new_n821_ );
and g735 ( new_n841_, new_n840_, new_n238_ );
or g736 ( N739, new_n839_, new_n841_ );
or g737 ( new_n843_, new_n793_, new_n796_ );
or g738 ( new_n844_, new_n843_, new_n209_ );
or g739 ( new_n845_, new_n416_, new_n364_ );
or g740 ( new_n846_, new_n845_, new_n209_ );
and g741 ( new_n847_, new_n844_, new_n846_ );
or g742 ( new_n848_, new_n847_, new_n764_ );
or g743 ( new_n849_, new_n764_, new_n767_ );
or g744 ( new_n850_, new_n311_, new_n209_ );
and g745 ( new_n851_, new_n849_, new_n850_ );
and g746 ( new_n852_, new_n364_, new_n796_ );
not g747 ( new_n853_, new_n852_ );
or g748 ( new_n854_, new_n851_, new_n853_ );
and g749 ( new_n855_, new_n848_, new_n854_ );
or g750 ( new_n856_, new_n855_, new_n796_ );
and g751 ( new_n857_, new_n733_, new_n728_ );
not g752 ( new_n858_, new_n857_ );
or g753 ( new_n859_, new_n856_, new_n858_ );
and g754 ( new_n860_, new_n859_, N65 );
or g755 ( new_n861_, new_n768_, new_n820_ );
and g756 ( new_n862_, new_n861_, new_n311_ );
and g757 ( new_n863_, new_n764_, new_n767_ );
or g758 ( new_n864_, new_n863_, new_n312_ );
and g759 ( new_n865_, new_n864_, new_n852_ );
or g760 ( new_n866_, new_n862_, new_n865_ );
and g761 ( new_n867_, new_n866_, new_n416_ );
and g762 ( new_n868_, new_n867_, new_n857_ );
and g763 ( new_n869_, new_n868_, new_n392_ );
or g764 ( N740, new_n860_, new_n869_ );
or g765 ( new_n871_, new_n855_, new_n364_ );
or g766 ( new_n872_, new_n871_, new_n858_ );
and g767 ( new_n873_, new_n872_, N69 );
and g768 ( new_n874_, new_n866_, new_n793_ );
and g769 ( new_n875_, new_n874_, new_n857_ );
and g770 ( new_n876_, new_n875_, new_n340_ );
or g771 ( N741, new_n873_, new_n876_ );
or g772 ( new_n878_, new_n855_, new_n767_ );
or g773 ( new_n879_, new_n878_, new_n858_ );
and g774 ( new_n880_, new_n879_, N73 );
and g775 ( new_n881_, new_n866_, new_n209_ );
and g776 ( new_n882_, new_n881_, new_n857_ );
and g777 ( new_n883_, new_n882_, new_n186_ );
or g778 ( N742, new_n880_, new_n883_ );
or g779 ( new_n885_, new_n855_, new_n311_ );
or g780 ( new_n886_, new_n885_, new_n858_ );
and g781 ( new_n887_, new_n886_, N77 );
and g782 ( new_n888_, new_n866_, new_n764_ );
and g783 ( new_n889_, new_n888_, new_n857_ );
and g784 ( new_n890_, new_n889_, new_n213_ );
or g785 ( N743, new_n887_, new_n890_ );
and g786 ( new_n892_, new_n729_, new_n708_ );
not g787 ( new_n893_, new_n892_ );
or g788 ( new_n894_, new_n856_, new_n893_ );
and g789 ( new_n895_, new_n894_, N81 );
and g790 ( new_n896_, new_n867_, new_n892_ );
and g791 ( new_n897_, new_n896_, new_n390_ );
or g792 ( N744, new_n895_, new_n897_ );
or g793 ( new_n899_, new_n871_, new_n893_ );
and g794 ( new_n900_, new_n899_, N85 );
and g795 ( new_n901_, new_n874_, new_n892_ );
and g796 ( new_n902_, new_n901_, new_n338_ );
or g797 ( N745, new_n900_, new_n902_ );
or g798 ( new_n904_, new_n878_, new_n893_ );
and g799 ( new_n905_, new_n904_, N89 );
and g800 ( new_n906_, new_n881_, new_n892_ );
and g801 ( new_n907_, new_n906_, new_n184_ );
or g802 ( N746, new_n905_, new_n907_ );
or g803 ( new_n909_, new_n885_, new_n893_ );
and g804 ( new_n910_, new_n909_, N93 );
and g805 ( new_n911_, new_n888_, new_n892_ );
and g806 ( new_n912_, new_n911_, new_n211_ );
or g807 ( N747, new_n910_, new_n912_ );
and g808 ( new_n914_, new_n733_, new_n726_ );
not g809 ( new_n915_, new_n914_ );
or g810 ( new_n916_, new_n856_, new_n915_ );
and g811 ( new_n917_, new_n916_, N97 );
and g812 ( new_n918_, new_n867_, new_n914_ );
and g813 ( new_n919_, new_n918_, new_n397_ );
or g814 ( N748, new_n917_, new_n919_ );
or g815 ( new_n921_, new_n871_, new_n915_ );
and g816 ( new_n922_, new_n921_, N101 );
and g817 ( new_n923_, new_n874_, new_n914_ );
and g818 ( new_n924_, new_n923_, new_n345_ );
or g819 ( N749, new_n922_, new_n924_ );
or g820 ( new_n926_, new_n878_, new_n915_ );
and g821 ( new_n927_, new_n926_, N105 );
and g822 ( new_n928_, new_n881_, new_n914_ );
and g823 ( new_n929_, new_n928_, new_n191_ );
or g824 ( N750, new_n927_, new_n929_ );
or g825 ( new_n931_, new_n885_, new_n915_ );
and g826 ( new_n932_, new_n931_, N109 );
and g827 ( new_n933_, new_n888_, new_n914_ );
and g828 ( new_n934_, new_n933_, new_n218_ );
or g829 ( N751, new_n932_, new_n934_ );
and g830 ( new_n936_, new_n727_, new_n708_ );
not g831 ( new_n937_, new_n936_ );
or g832 ( new_n938_, new_n856_, new_n937_ );
and g833 ( new_n939_, new_n938_, N113 );
and g834 ( new_n940_, new_n867_, new_n936_ );
and g835 ( new_n941_, new_n940_, new_n395_ );
or g836 ( N752, new_n939_, new_n941_ );
or g837 ( new_n943_, new_n871_, new_n937_ );
and g838 ( new_n944_, new_n943_, N117 );
and g839 ( new_n945_, new_n874_, new_n936_ );
and g840 ( new_n946_, new_n945_, new_n343_ );
or g841 ( N753, new_n944_, new_n946_ );
or g842 ( new_n948_, new_n878_, new_n937_ );
and g843 ( new_n949_, new_n948_, N121 );
and g844 ( new_n950_, new_n881_, new_n936_ );
and g845 ( new_n951_, new_n950_, new_n189_ );
or g846 ( N754, new_n949_, new_n951_ );
or g847 ( new_n953_, new_n885_, new_n937_ );
and g848 ( new_n954_, new_n953_, N125 );
and g849 ( new_n955_, new_n888_, new_n936_ );
and g850 ( new_n956_, new_n955_, new_n216_ );
or g851 ( N755, new_n954_, new_n956_ );
endmodule