module add_mul_comp_sub_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, 
        a_17_, a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, 
        a_27_, a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, 
        b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, 
        b_16_, b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, 
        b_26_, b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, 
        Result_32_, Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, 
        Result_38_, Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, 
        Result_44_, Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, 
        Result_50_, Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, 
        Result_56_, Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, 
        Result_62_, Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   Result_9_, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_31_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_28_ = Result_9_;
  assign Result_26_ = Result_9_;
  assign Result_24_ = Result_9_;
  assign Result_22_ = Result_9_;
  assign Result_20_ = Result_9_;
  assign Result_19_ = Result_9_;
  assign Result_17_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_16_ = Result_9_;
  assign Result_18_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_21_ = Result_9_;
  assign Result_23_ = Result_9_;
  assign Result_25_ = Result_9_;
  assign Result_27_ = Result_9_;
  assign Result_29_ = Result_9_;
  assign Result_30_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  OR2_X2 U749 ( .A1(n1241), .A2(n1242), .ZN(Result_9_) );
  INV_X1 U750 ( .A(n716), .ZN(Result_63_) );
  AND2_X1 U751 ( .A1(n717), .A2(n718), .ZN(n716) );
  OR2_X1 U752 ( .A1(n719), .A2(n720), .ZN(Result_62_) );
  AND2_X1 U753 ( .A1(n721), .A2(n722), .ZN(n720) );
  OR2_X1 U754 ( .A1(n723), .A2(n724), .ZN(n722) );
  AND2_X1 U755 ( .A1(Result_9_), .A2(n717), .ZN(n724) );
  INV_X1 U756 ( .A(n725), .ZN(n717) );
  INV_X1 U757 ( .A(n726), .ZN(n723) );
  OR2_X1 U758 ( .A1(n727), .A2(n728), .ZN(n726) );
  AND2_X1 U759 ( .A1(n729), .A2(n730), .ZN(n719) );
  OR2_X1 U760 ( .A1(n731), .A2(n732), .ZN(n730) );
  AND2_X1 U761 ( .A1(n725), .A2(Result_9_), .ZN(n732) );
  AND2_X1 U762 ( .A1(n728), .A2(n733), .ZN(n731) );
  AND2_X1 U763 ( .A1(a_31_), .A2(b_31_), .ZN(n728) );
  INV_X1 U764 ( .A(n721), .ZN(n729) );
  OR2_X1 U765 ( .A1(n734), .A2(n735), .ZN(n721) );
  INV_X1 U766 ( .A(n736), .ZN(n735) );
  OR2_X1 U767 ( .A1(n737), .A2(n738), .ZN(Result_61_) );
  AND2_X1 U768 ( .A1(n739), .A2(Result_9_), .ZN(n738) );
  OR2_X1 U769 ( .A1(n740), .A2(n741), .ZN(n739) );
  INV_X1 U770 ( .A(n742), .ZN(n741) );
  OR2_X1 U771 ( .A1(n743), .A2(n744), .ZN(n742) );
  AND2_X1 U772 ( .A1(n744), .A2(n743), .ZN(n740) );
  AND2_X1 U773 ( .A1(n733), .A2(n745), .ZN(n737) );
  OR2_X1 U774 ( .A1(n746), .A2(n747), .ZN(n745) );
  INV_X1 U775 ( .A(n748), .ZN(n747) );
  OR2_X1 U776 ( .A1(n749), .A2(n744), .ZN(n748) );
  AND2_X1 U777 ( .A1(n744), .A2(n749), .ZN(n746) );
  AND2_X1 U778 ( .A1(n750), .A2(n751), .ZN(n744) );
  OR2_X1 U779 ( .A1(n752), .A2(b_29_), .ZN(n751) );
  OR2_X1 U780 ( .A1(n753), .A2(n754), .ZN(Result_60_) );
  AND2_X1 U781 ( .A1(n755), .A2(Result_9_), .ZN(n754) );
  OR2_X1 U782 ( .A1(n756), .A2(n757), .ZN(n755) );
  INV_X1 U783 ( .A(n758), .ZN(n757) );
  OR2_X1 U784 ( .A1(n759), .A2(n760), .ZN(n758) );
  AND2_X1 U785 ( .A1(n760), .A2(n759), .ZN(n756) );
  AND2_X1 U786 ( .A1(n761), .A2(n733), .ZN(n753) );
  AND2_X1 U787 ( .A1(n762), .A2(n763), .ZN(n761) );
  INV_X1 U788 ( .A(n764), .ZN(n763) );
  AND2_X1 U789 ( .A1(n765), .A2(n760), .ZN(n764) );
  OR2_X1 U790 ( .A1(n760), .A2(n765), .ZN(n762) );
  AND2_X1 U791 ( .A1(n766), .A2(n767), .ZN(n760) );
  OR2_X1 U792 ( .A1(n768), .A2(b_28_), .ZN(n767) );
  OR2_X1 U793 ( .A1(n769), .A2(n770), .ZN(Result_59_) );
  AND2_X1 U794 ( .A1(n771), .A2(Result_9_), .ZN(n770) );
  OR2_X1 U795 ( .A1(n772), .A2(n773), .ZN(n771) );
  INV_X1 U796 ( .A(n774), .ZN(n773) );
  OR2_X1 U797 ( .A1(n775), .A2(n776), .ZN(n774) );
  AND2_X1 U798 ( .A1(n776), .A2(n775), .ZN(n772) );
  AND2_X1 U799 ( .A1(n777), .A2(n733), .ZN(n769) );
  AND2_X1 U800 ( .A1(n778), .A2(n779), .ZN(n777) );
  INV_X1 U801 ( .A(n780), .ZN(n779) );
  AND2_X1 U802 ( .A1(n781), .A2(n776), .ZN(n780) );
  OR2_X1 U803 ( .A1(n776), .A2(n781), .ZN(n778) );
  AND2_X1 U804 ( .A1(n782), .A2(n783), .ZN(n776) );
  OR2_X1 U805 ( .A1(n784), .A2(b_27_), .ZN(n783) );
  OR2_X1 U806 ( .A1(n785), .A2(n786), .ZN(Result_58_) );
  AND2_X1 U807 ( .A1(n787), .A2(Result_9_), .ZN(n786) );
  OR2_X1 U808 ( .A1(n788), .A2(n789), .ZN(n787) );
  INV_X1 U809 ( .A(n790), .ZN(n789) );
  OR2_X1 U810 ( .A1(n791), .A2(n792), .ZN(n790) );
  AND2_X1 U811 ( .A1(n792), .A2(n791), .ZN(n788) );
  AND2_X1 U812 ( .A1(n793), .A2(n733), .ZN(n785) );
  AND2_X1 U813 ( .A1(n794), .A2(n795), .ZN(n793) );
  INV_X1 U814 ( .A(n796), .ZN(n795) );
  AND2_X1 U815 ( .A1(n797), .A2(n792), .ZN(n796) );
  OR2_X1 U816 ( .A1(n792), .A2(n797), .ZN(n794) );
  AND2_X1 U817 ( .A1(n798), .A2(n799), .ZN(n792) );
  OR2_X1 U818 ( .A1(n800), .A2(b_26_), .ZN(n799) );
  OR2_X1 U819 ( .A1(n801), .A2(n802), .ZN(Result_57_) );
  AND2_X1 U820 ( .A1(n803), .A2(Result_9_), .ZN(n802) );
  OR2_X1 U821 ( .A1(n804), .A2(n805), .ZN(n803) );
  INV_X1 U822 ( .A(n806), .ZN(n805) );
  OR2_X1 U823 ( .A1(n807), .A2(n808), .ZN(n806) );
  AND2_X1 U824 ( .A1(n808), .A2(n807), .ZN(n804) );
  AND2_X1 U825 ( .A1(n809), .A2(n733), .ZN(n801) );
  AND2_X1 U826 ( .A1(n810), .A2(n811), .ZN(n809) );
  INV_X1 U827 ( .A(n812), .ZN(n811) );
  AND2_X1 U828 ( .A1(n813), .A2(n808), .ZN(n812) );
  OR2_X1 U829 ( .A1(n808), .A2(n813), .ZN(n810) );
  AND2_X1 U830 ( .A1(n814), .A2(n815), .ZN(n808) );
  OR2_X1 U831 ( .A1(n816), .A2(b_25_), .ZN(n815) );
  OR2_X1 U832 ( .A1(n817), .A2(n818), .ZN(Result_56_) );
  AND2_X1 U833 ( .A1(n819), .A2(Result_9_), .ZN(n818) );
  OR2_X1 U834 ( .A1(n820), .A2(n821), .ZN(n819) );
  INV_X1 U835 ( .A(n822), .ZN(n821) );
  OR2_X1 U836 ( .A1(n823), .A2(n824), .ZN(n822) );
  AND2_X1 U837 ( .A1(n824), .A2(n823), .ZN(n820) );
  AND2_X1 U838 ( .A1(n825), .A2(n733), .ZN(n817) );
  AND2_X1 U839 ( .A1(n826), .A2(n827), .ZN(n825) );
  INV_X1 U840 ( .A(n828), .ZN(n827) );
  AND2_X1 U841 ( .A1(n829), .A2(n824), .ZN(n828) );
  OR2_X1 U842 ( .A1(n824), .A2(n829), .ZN(n826) );
  AND2_X1 U843 ( .A1(n830), .A2(n831), .ZN(n824) );
  OR2_X1 U844 ( .A1(n832), .A2(b_24_), .ZN(n831) );
  OR2_X1 U845 ( .A1(n833), .A2(n834), .ZN(Result_55_) );
  AND2_X1 U846 ( .A1(n835), .A2(Result_9_), .ZN(n834) );
  OR2_X1 U847 ( .A1(n836), .A2(n837), .ZN(n835) );
  INV_X1 U848 ( .A(n838), .ZN(n837) );
  OR2_X1 U849 ( .A1(n839), .A2(n840), .ZN(n838) );
  AND2_X1 U850 ( .A1(n840), .A2(n839), .ZN(n836) );
  AND2_X1 U851 ( .A1(n841), .A2(n733), .ZN(n833) );
  AND2_X1 U852 ( .A1(n842), .A2(n843), .ZN(n841) );
  INV_X1 U853 ( .A(n844), .ZN(n843) );
  AND2_X1 U854 ( .A1(n845), .A2(n840), .ZN(n844) );
  OR2_X1 U855 ( .A1(n840), .A2(n845), .ZN(n842) );
  AND2_X1 U856 ( .A1(n846), .A2(n847), .ZN(n840) );
  OR2_X1 U857 ( .A1(n848), .A2(b_23_), .ZN(n847) );
  OR2_X1 U858 ( .A1(n849), .A2(n850), .ZN(Result_54_) );
  AND2_X1 U859 ( .A1(n851), .A2(Result_9_), .ZN(n850) );
  OR2_X1 U860 ( .A1(n852), .A2(n853), .ZN(n851) );
  INV_X1 U861 ( .A(n854), .ZN(n853) );
  OR2_X1 U862 ( .A1(n855), .A2(n856), .ZN(n854) );
  AND2_X1 U863 ( .A1(n856), .A2(n855), .ZN(n852) );
  AND2_X1 U864 ( .A1(n857), .A2(n733), .ZN(n849) );
  AND2_X1 U865 ( .A1(n858), .A2(n859), .ZN(n857) );
  INV_X1 U866 ( .A(n860), .ZN(n859) );
  AND2_X1 U867 ( .A1(n861), .A2(n856), .ZN(n860) );
  OR2_X1 U868 ( .A1(n856), .A2(n861), .ZN(n858) );
  AND2_X1 U869 ( .A1(n862), .A2(n863), .ZN(n856) );
  OR2_X1 U870 ( .A1(n864), .A2(b_22_), .ZN(n863) );
  OR2_X1 U871 ( .A1(n865), .A2(n866), .ZN(Result_53_) );
  AND2_X1 U872 ( .A1(n867), .A2(Result_9_), .ZN(n866) );
  OR2_X1 U873 ( .A1(n868), .A2(n869), .ZN(n867) );
  INV_X1 U874 ( .A(n870), .ZN(n869) );
  OR2_X1 U875 ( .A1(n871), .A2(n872), .ZN(n870) );
  AND2_X1 U876 ( .A1(n872), .A2(n871), .ZN(n868) );
  AND2_X1 U877 ( .A1(n873), .A2(n733), .ZN(n865) );
  AND2_X1 U878 ( .A1(n874), .A2(n875), .ZN(n873) );
  INV_X1 U879 ( .A(n876), .ZN(n875) );
  AND2_X1 U880 ( .A1(n877), .A2(n872), .ZN(n876) );
  OR2_X1 U881 ( .A1(n872), .A2(n877), .ZN(n874) );
  AND2_X1 U882 ( .A1(n878), .A2(n879), .ZN(n872) );
  OR2_X1 U883 ( .A1(n880), .A2(b_21_), .ZN(n879) );
  OR2_X1 U884 ( .A1(n881), .A2(n882), .ZN(Result_52_) );
  AND2_X1 U885 ( .A1(n883), .A2(Result_9_), .ZN(n882) );
  OR2_X1 U886 ( .A1(n884), .A2(n885), .ZN(n883) );
  INV_X1 U887 ( .A(n886), .ZN(n885) );
  OR2_X1 U888 ( .A1(n887), .A2(n888), .ZN(n886) );
  AND2_X1 U889 ( .A1(n888), .A2(n887), .ZN(n884) );
  AND2_X1 U890 ( .A1(n889), .A2(n733), .ZN(n881) );
  AND2_X1 U891 ( .A1(n890), .A2(n891), .ZN(n889) );
  INV_X1 U892 ( .A(n892), .ZN(n891) );
  AND2_X1 U893 ( .A1(n893), .A2(n888), .ZN(n892) );
  OR2_X1 U894 ( .A1(n888), .A2(n893), .ZN(n890) );
  AND2_X1 U895 ( .A1(n894), .A2(n895), .ZN(n888) );
  OR2_X1 U896 ( .A1(n896), .A2(b_20_), .ZN(n895) );
  OR2_X1 U897 ( .A1(n897), .A2(n898), .ZN(Result_51_) );
  AND2_X1 U898 ( .A1(n899), .A2(Result_9_), .ZN(n898) );
  OR2_X1 U899 ( .A1(n900), .A2(n901), .ZN(n899) );
  INV_X1 U900 ( .A(n902), .ZN(n901) );
  OR2_X1 U901 ( .A1(n903), .A2(n904), .ZN(n902) );
  AND2_X1 U902 ( .A1(n904), .A2(n903), .ZN(n900) );
  AND2_X1 U903 ( .A1(n905), .A2(n733), .ZN(n897) );
  AND2_X1 U904 ( .A1(n906), .A2(n907), .ZN(n905) );
  INV_X1 U905 ( .A(n908), .ZN(n907) );
  AND2_X1 U906 ( .A1(n909), .A2(n904), .ZN(n908) );
  OR2_X1 U907 ( .A1(n904), .A2(n909), .ZN(n906) );
  AND2_X1 U908 ( .A1(n910), .A2(n911), .ZN(n904) );
  OR2_X1 U909 ( .A1(n912), .A2(b_19_), .ZN(n911) );
  OR2_X1 U910 ( .A1(n913), .A2(n914), .ZN(Result_50_) );
  AND2_X1 U911 ( .A1(n915), .A2(Result_9_), .ZN(n914) );
  OR2_X1 U912 ( .A1(n916), .A2(n917), .ZN(n915) );
  INV_X1 U913 ( .A(n918), .ZN(n917) );
  OR2_X1 U914 ( .A1(n919), .A2(n920), .ZN(n918) );
  AND2_X1 U915 ( .A1(n920), .A2(n919), .ZN(n916) );
  AND2_X1 U916 ( .A1(n921), .A2(n733), .ZN(n913) );
  AND2_X1 U917 ( .A1(n922), .A2(n923), .ZN(n921) );
  INV_X1 U918 ( .A(n924), .ZN(n923) );
  AND2_X1 U919 ( .A1(n925), .A2(n920), .ZN(n924) );
  OR2_X1 U920 ( .A1(n920), .A2(n925), .ZN(n922) );
  AND2_X1 U921 ( .A1(n926), .A2(n927), .ZN(n920) );
  OR2_X1 U922 ( .A1(n928), .A2(b_18_), .ZN(n927) );
  OR2_X1 U923 ( .A1(n929), .A2(n930), .ZN(Result_49_) );
  AND2_X1 U924 ( .A1(n931), .A2(Result_9_), .ZN(n930) );
  OR2_X1 U925 ( .A1(n932), .A2(n933), .ZN(n931) );
  INV_X1 U926 ( .A(n934), .ZN(n933) );
  OR2_X1 U927 ( .A1(n935), .A2(n936), .ZN(n934) );
  AND2_X1 U928 ( .A1(n936), .A2(n935), .ZN(n932) );
  AND2_X1 U929 ( .A1(n937), .A2(n733), .ZN(n929) );
  AND2_X1 U930 ( .A1(n938), .A2(n939), .ZN(n937) );
  INV_X1 U931 ( .A(n940), .ZN(n939) );
  AND2_X1 U932 ( .A1(n941), .A2(n936), .ZN(n940) );
  OR2_X1 U933 ( .A1(n936), .A2(n941), .ZN(n938) );
  AND2_X1 U934 ( .A1(n942), .A2(n943), .ZN(n936) );
  OR2_X1 U935 ( .A1(n944), .A2(b_17_), .ZN(n943) );
  OR2_X1 U936 ( .A1(n945), .A2(n946), .ZN(Result_48_) );
  AND2_X1 U937 ( .A1(n947), .A2(Result_9_), .ZN(n946) );
  OR2_X1 U938 ( .A1(n948), .A2(n949), .ZN(n947) );
  INV_X1 U939 ( .A(n950), .ZN(n949) );
  OR2_X1 U940 ( .A1(n951), .A2(n952), .ZN(n950) );
  AND2_X1 U941 ( .A1(n952), .A2(n951), .ZN(n948) );
  AND2_X1 U942 ( .A1(n953), .A2(n733), .ZN(n945) );
  AND2_X1 U943 ( .A1(n954), .A2(n955), .ZN(n953) );
  INV_X1 U944 ( .A(n956), .ZN(n955) );
  AND2_X1 U945 ( .A1(n957), .A2(n952), .ZN(n956) );
  OR2_X1 U946 ( .A1(n952), .A2(n957), .ZN(n954) );
  AND2_X1 U947 ( .A1(n958), .A2(n959), .ZN(n952) );
  OR2_X1 U948 ( .A1(n960), .A2(b_16_), .ZN(n959) );
  OR2_X1 U949 ( .A1(n961), .A2(n962), .ZN(Result_47_) );
  AND2_X1 U950 ( .A1(n963), .A2(Result_9_), .ZN(n962) );
  OR2_X1 U951 ( .A1(n964), .A2(n965), .ZN(n963) );
  INV_X1 U952 ( .A(n966), .ZN(n965) );
  OR2_X1 U953 ( .A1(n967), .A2(n968), .ZN(n966) );
  AND2_X1 U954 ( .A1(n968), .A2(n967), .ZN(n964) );
  AND2_X1 U955 ( .A1(n969), .A2(n733), .ZN(n961) );
  AND2_X1 U956 ( .A1(n970), .A2(n971), .ZN(n969) );
  INV_X1 U957 ( .A(n972), .ZN(n971) );
  AND2_X1 U958 ( .A1(n973), .A2(n968), .ZN(n972) );
  OR2_X1 U959 ( .A1(n968), .A2(n973), .ZN(n970) );
  AND2_X1 U960 ( .A1(n974), .A2(n975), .ZN(n968) );
  OR2_X1 U961 ( .A1(n976), .A2(b_15_), .ZN(n975) );
  OR2_X1 U962 ( .A1(n977), .A2(n978), .ZN(Result_46_) );
  AND2_X1 U963 ( .A1(n979), .A2(Result_9_), .ZN(n978) );
  OR2_X1 U964 ( .A1(n980), .A2(n981), .ZN(n979) );
  INV_X1 U965 ( .A(n982), .ZN(n981) );
  OR2_X1 U966 ( .A1(n983), .A2(n984), .ZN(n982) );
  AND2_X1 U967 ( .A1(n984), .A2(n983), .ZN(n980) );
  AND2_X1 U968 ( .A1(n985), .A2(n733), .ZN(n977) );
  AND2_X1 U969 ( .A1(n986), .A2(n987), .ZN(n985) );
  INV_X1 U970 ( .A(n988), .ZN(n987) );
  AND2_X1 U971 ( .A1(n989), .A2(n984), .ZN(n988) );
  OR2_X1 U972 ( .A1(n984), .A2(n989), .ZN(n986) );
  AND2_X1 U973 ( .A1(n990), .A2(n991), .ZN(n984) );
  OR2_X1 U974 ( .A1(n992), .A2(b_14_), .ZN(n991) );
  OR2_X1 U975 ( .A1(n993), .A2(n994), .ZN(Result_45_) );
  AND2_X1 U976 ( .A1(n995), .A2(Result_9_), .ZN(n994) );
  OR2_X1 U977 ( .A1(n996), .A2(n997), .ZN(n995) );
  INV_X1 U978 ( .A(n998), .ZN(n997) );
  OR2_X1 U979 ( .A1(n999), .A2(n1000), .ZN(n998) );
  AND2_X1 U980 ( .A1(n1000), .A2(n999), .ZN(n996) );
  AND2_X1 U981 ( .A1(n1001), .A2(n733), .ZN(n993) );
  AND2_X1 U982 ( .A1(n1002), .A2(n1003), .ZN(n1001) );
  INV_X1 U983 ( .A(n1004), .ZN(n1003) );
  AND2_X1 U984 ( .A1(n1005), .A2(n1000), .ZN(n1004) );
  OR2_X1 U985 ( .A1(n1000), .A2(n1005), .ZN(n1002) );
  AND2_X1 U986 ( .A1(n1006), .A2(n1007), .ZN(n1000) );
  OR2_X1 U987 ( .A1(n1008), .A2(b_13_), .ZN(n1007) );
  OR2_X1 U988 ( .A1(n1009), .A2(n1010), .ZN(Result_44_) );
  AND2_X1 U989 ( .A1(n1011), .A2(Result_9_), .ZN(n1010) );
  OR2_X1 U990 ( .A1(n1012), .A2(n1013), .ZN(n1011) );
  INV_X1 U991 ( .A(n1014), .ZN(n1013) );
  OR2_X1 U992 ( .A1(n1015), .A2(n1016), .ZN(n1014) );
  AND2_X1 U993 ( .A1(n1016), .A2(n1015), .ZN(n1012) );
  AND2_X1 U994 ( .A1(n1017), .A2(n733), .ZN(n1009) );
  AND2_X1 U995 ( .A1(n1018), .A2(n1019), .ZN(n1017) );
  INV_X1 U996 ( .A(n1020), .ZN(n1019) );
  AND2_X1 U997 ( .A1(n1021), .A2(n1016), .ZN(n1020) );
  OR2_X1 U998 ( .A1(n1016), .A2(n1021), .ZN(n1018) );
  AND2_X1 U999 ( .A1(n1022), .A2(n1023), .ZN(n1016) );
  OR2_X1 U1000 ( .A1(n1024), .A2(b_12_), .ZN(n1023) );
  OR2_X1 U1001 ( .A1(n1025), .A2(n1026), .ZN(Result_43_) );
  AND2_X1 U1002 ( .A1(n1027), .A2(Result_9_), .ZN(n1026) );
  OR2_X1 U1003 ( .A1(n1028), .A2(n1029), .ZN(n1027) );
  INV_X1 U1004 ( .A(n1030), .ZN(n1029) );
  OR2_X1 U1005 ( .A1(n1031), .A2(n1032), .ZN(n1030) );
  AND2_X1 U1006 ( .A1(n1032), .A2(n1031), .ZN(n1028) );
  AND2_X1 U1007 ( .A1(n1033), .A2(n733), .ZN(n1025) );
  AND2_X1 U1008 ( .A1(n1034), .A2(n1035), .ZN(n1033) );
  INV_X1 U1009 ( .A(n1036), .ZN(n1035) );
  AND2_X1 U1010 ( .A1(n1037), .A2(n1032), .ZN(n1036) );
  OR2_X1 U1011 ( .A1(n1032), .A2(n1037), .ZN(n1034) );
  AND2_X1 U1012 ( .A1(n1038), .A2(n1039), .ZN(n1032) );
  OR2_X1 U1013 ( .A1(n1040), .A2(b_11_), .ZN(n1039) );
  OR2_X1 U1014 ( .A1(n1041), .A2(n1042), .ZN(Result_42_) );
  AND2_X1 U1015 ( .A1(n1043), .A2(Result_9_), .ZN(n1042) );
  OR2_X1 U1016 ( .A1(n1044), .A2(n1045), .ZN(n1043) );
  INV_X1 U1017 ( .A(n1046), .ZN(n1045) );
  OR2_X1 U1018 ( .A1(n1047), .A2(n1048), .ZN(n1046) );
  AND2_X1 U1019 ( .A1(n1048), .A2(n1047), .ZN(n1044) );
  AND2_X1 U1020 ( .A1(n1049), .A2(n733), .ZN(n1041) );
  AND2_X1 U1021 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
  INV_X1 U1022 ( .A(n1052), .ZN(n1051) );
  AND2_X1 U1023 ( .A1(n1053), .A2(n1048), .ZN(n1052) );
  OR2_X1 U1024 ( .A1(n1048), .A2(n1053), .ZN(n1050) );
  AND2_X1 U1025 ( .A1(n1054), .A2(n1055), .ZN(n1048) );
  OR2_X1 U1026 ( .A1(n1056), .A2(b_10_), .ZN(n1055) );
  OR2_X1 U1027 ( .A1(n1057), .A2(n1058), .ZN(Result_41_) );
  AND2_X1 U1028 ( .A1(n1059), .A2(Result_9_), .ZN(n1058) );
  OR2_X1 U1029 ( .A1(n1060), .A2(n1061), .ZN(n1059) );
  INV_X1 U1030 ( .A(n1062), .ZN(n1061) );
  OR2_X1 U1031 ( .A1(n1063), .A2(n1064), .ZN(n1062) );
  AND2_X1 U1032 ( .A1(n1064), .A2(n1063), .ZN(n1060) );
  AND2_X1 U1033 ( .A1(n1065), .A2(n733), .ZN(n1057) );
  AND2_X1 U1034 ( .A1(n1066), .A2(n1067), .ZN(n1065) );
  INV_X1 U1035 ( .A(n1068), .ZN(n1067) );
  AND2_X1 U1036 ( .A1(n1069), .A2(n1064), .ZN(n1068) );
  OR2_X1 U1037 ( .A1(n1064), .A2(n1069), .ZN(n1066) );
  AND2_X1 U1038 ( .A1(n1070), .A2(n1071), .ZN(n1064) );
  OR2_X1 U1039 ( .A1(n1072), .A2(b_9_), .ZN(n1071) );
  OR2_X1 U1040 ( .A1(n1073), .A2(n1074), .ZN(Result_40_) );
  AND2_X1 U1041 ( .A1(n1075), .A2(Result_9_), .ZN(n1074) );
  OR2_X1 U1042 ( .A1(n1076), .A2(n1077), .ZN(n1075) );
  INV_X1 U1043 ( .A(n1078), .ZN(n1077) );
  OR2_X1 U1044 ( .A1(n1079), .A2(n1080), .ZN(n1078) );
  AND2_X1 U1045 ( .A1(n1080), .A2(n1079), .ZN(n1076) );
  AND2_X1 U1046 ( .A1(n1081), .A2(n733), .ZN(n1073) );
  AND2_X1 U1047 ( .A1(n1082), .A2(n1083), .ZN(n1081) );
  INV_X1 U1048 ( .A(n1084), .ZN(n1083) );
  AND2_X1 U1049 ( .A1(n1085), .A2(n1080), .ZN(n1084) );
  OR2_X1 U1050 ( .A1(n1080), .A2(n1085), .ZN(n1082) );
  AND2_X1 U1051 ( .A1(n1086), .A2(n1087), .ZN(n1080) );
  OR2_X1 U1052 ( .A1(n1088), .A2(b_8_), .ZN(n1087) );
  OR2_X1 U1053 ( .A1(n1089), .A2(n1090), .ZN(Result_39_) );
  AND2_X1 U1054 ( .A1(n1091), .A2(Result_9_), .ZN(n1090) );
  OR2_X1 U1055 ( .A1(n1092), .A2(n1093), .ZN(n1091) );
  INV_X1 U1056 ( .A(n1094), .ZN(n1093) );
  OR2_X1 U1057 ( .A1(n1095), .A2(n1096), .ZN(n1094) );
  AND2_X1 U1058 ( .A1(n1096), .A2(n1095), .ZN(n1092) );
  AND2_X1 U1059 ( .A1(n1097), .A2(n733), .ZN(n1089) );
  AND2_X1 U1060 ( .A1(n1098), .A2(n1099), .ZN(n1097) );
  INV_X1 U1061 ( .A(n1100), .ZN(n1099) );
  AND2_X1 U1062 ( .A1(n1101), .A2(n1096), .ZN(n1100) );
  OR2_X1 U1063 ( .A1(n1096), .A2(n1101), .ZN(n1098) );
  AND2_X1 U1064 ( .A1(n1102), .A2(n1103), .ZN(n1096) );
  OR2_X1 U1065 ( .A1(n1104), .A2(b_7_), .ZN(n1103) );
  OR2_X1 U1066 ( .A1(n1105), .A2(n1106), .ZN(Result_38_) );
  AND2_X1 U1067 ( .A1(n1107), .A2(Result_9_), .ZN(n1106) );
  OR2_X1 U1068 ( .A1(n1108), .A2(n1109), .ZN(n1107) );
  INV_X1 U1069 ( .A(n1110), .ZN(n1109) );
  OR2_X1 U1070 ( .A1(n1111), .A2(n1112), .ZN(n1110) );
  AND2_X1 U1071 ( .A1(n1112), .A2(n1111), .ZN(n1108) );
  AND2_X1 U1072 ( .A1(n1113), .A2(n733), .ZN(n1105) );
  AND2_X1 U1073 ( .A1(n1114), .A2(n1115), .ZN(n1113) );
  INV_X1 U1074 ( .A(n1116), .ZN(n1115) );
  AND2_X1 U1075 ( .A1(n1117), .A2(n1112), .ZN(n1116) );
  OR2_X1 U1076 ( .A1(n1112), .A2(n1117), .ZN(n1114) );
  AND2_X1 U1077 ( .A1(n1118), .A2(n1119), .ZN(n1112) );
  OR2_X1 U1078 ( .A1(n1120), .A2(b_6_), .ZN(n1119) );
  OR2_X1 U1079 ( .A1(n1121), .A2(n1122), .ZN(Result_37_) );
  AND2_X1 U1080 ( .A1(n1123), .A2(Result_9_), .ZN(n1122) );
  OR2_X1 U1081 ( .A1(n1124), .A2(n1125), .ZN(n1123) );
  INV_X1 U1082 ( .A(n1126), .ZN(n1125) );
  OR2_X1 U1083 ( .A1(n1127), .A2(n1128), .ZN(n1126) );
  AND2_X1 U1084 ( .A1(n1128), .A2(n1127), .ZN(n1124) );
  AND2_X1 U1085 ( .A1(n1129), .A2(n733), .ZN(n1121) );
  AND2_X1 U1086 ( .A1(n1130), .A2(n1131), .ZN(n1129) );
  INV_X1 U1087 ( .A(n1132), .ZN(n1131) );
  AND2_X1 U1088 ( .A1(n1133), .A2(n1128), .ZN(n1132) );
  OR2_X1 U1089 ( .A1(n1128), .A2(n1133), .ZN(n1130) );
  AND2_X1 U1090 ( .A1(n1134), .A2(n1135), .ZN(n1128) );
  OR2_X1 U1091 ( .A1(n1136), .A2(b_5_), .ZN(n1135) );
  OR2_X1 U1092 ( .A1(n1137), .A2(n1138), .ZN(Result_36_) );
  AND2_X1 U1093 ( .A1(n1139), .A2(Result_9_), .ZN(n1138) );
  OR2_X1 U1094 ( .A1(n1140), .A2(n1141), .ZN(n1139) );
  INV_X1 U1095 ( .A(n1142), .ZN(n1141) );
  OR2_X1 U1096 ( .A1(n1143), .A2(n1144), .ZN(n1142) );
  AND2_X1 U1097 ( .A1(n1144), .A2(n1143), .ZN(n1140) );
  AND2_X1 U1098 ( .A1(n1145), .A2(n733), .ZN(n1137) );
  AND2_X1 U1099 ( .A1(n1146), .A2(n1147), .ZN(n1145) );
  INV_X1 U1100 ( .A(n1148), .ZN(n1147) );
  AND2_X1 U1101 ( .A1(n1149), .A2(n1144), .ZN(n1148) );
  OR2_X1 U1102 ( .A1(n1144), .A2(n1149), .ZN(n1146) );
  AND2_X1 U1103 ( .A1(n1150), .A2(n1151), .ZN(n1144) );
  OR2_X1 U1104 ( .A1(n1152), .A2(b_4_), .ZN(n1151) );
  OR2_X1 U1105 ( .A1(n1153), .A2(n1154), .ZN(Result_35_) );
  AND2_X1 U1106 ( .A1(n1155), .A2(Result_9_), .ZN(n1154) );
  OR2_X1 U1107 ( .A1(n1156), .A2(n1157), .ZN(n1155) );
  INV_X1 U1108 ( .A(n1158), .ZN(n1157) );
  OR2_X1 U1109 ( .A1(n1159), .A2(n1160), .ZN(n1158) );
  AND2_X1 U1110 ( .A1(n1160), .A2(n1159), .ZN(n1156) );
  AND2_X1 U1111 ( .A1(n1161), .A2(n733), .ZN(n1153) );
  AND2_X1 U1112 ( .A1(n1162), .A2(n1163), .ZN(n1161) );
  INV_X1 U1113 ( .A(n1164), .ZN(n1163) );
  AND2_X1 U1114 ( .A1(n1165), .A2(n1160), .ZN(n1164) );
  OR2_X1 U1115 ( .A1(n1160), .A2(n1165), .ZN(n1162) );
  AND2_X1 U1116 ( .A1(n1166), .A2(n1167), .ZN(n1160) );
  OR2_X1 U1117 ( .A1(n1168), .A2(b_3_), .ZN(n1167) );
  OR2_X1 U1118 ( .A1(n1169), .A2(n1170), .ZN(Result_34_) );
  AND2_X1 U1119 ( .A1(n1171), .A2(Result_9_), .ZN(n1170) );
  OR2_X1 U1120 ( .A1(n1172), .A2(n1173), .ZN(n1171) );
  INV_X1 U1121 ( .A(n1174), .ZN(n1173) );
  OR2_X1 U1122 ( .A1(n1175), .A2(n1176), .ZN(n1174) );
  AND2_X1 U1123 ( .A1(n1176), .A2(n1175), .ZN(n1172) );
  AND2_X1 U1124 ( .A1(n1177), .A2(n733), .ZN(n1169) );
  AND2_X1 U1125 ( .A1(n1178), .A2(n1179), .ZN(n1177) );
  INV_X1 U1126 ( .A(n1180), .ZN(n1179) );
  AND2_X1 U1127 ( .A1(n1181), .A2(n1176), .ZN(n1180) );
  OR2_X1 U1128 ( .A1(n1176), .A2(n1181), .ZN(n1178) );
  AND2_X1 U1129 ( .A1(n1182), .A2(n1183), .ZN(n1176) );
  OR2_X1 U1130 ( .A1(n1184), .A2(b_2_), .ZN(n1183) );
  OR2_X1 U1131 ( .A1(n1185), .A2(n1186), .ZN(Result_33_) );
  AND2_X1 U1132 ( .A1(n1187), .A2(Result_9_), .ZN(n1186) );
  OR2_X1 U1133 ( .A1(n1188), .A2(n1189), .ZN(n1187) );
  INV_X1 U1134 ( .A(n1190), .ZN(n1189) );
  OR2_X1 U1135 ( .A1(n1191), .A2(n1192), .ZN(n1190) );
  AND2_X1 U1136 ( .A1(n1192), .A2(n1191), .ZN(n1188) );
  AND2_X1 U1137 ( .A1(n1193), .A2(n733), .ZN(n1185) );
  AND2_X1 U1138 ( .A1(n1194), .A2(n1195), .ZN(n1193) );
  INV_X1 U1139 ( .A(n1196), .ZN(n1195) );
  AND2_X1 U1140 ( .A1(n1197), .A2(n1192), .ZN(n1196) );
  OR2_X1 U1141 ( .A1(n1192), .A2(n1197), .ZN(n1194) );
  AND2_X1 U1142 ( .A1(n1198), .A2(n1199), .ZN(n1192) );
  OR2_X1 U1143 ( .A1(n1200), .A2(b_1_), .ZN(n1199) );
  OR2_X1 U1144 ( .A1(n1201), .A2(n1202), .ZN(Result_32_) );
  AND2_X1 U1145 ( .A1(n1203), .A2(Result_9_), .ZN(n1202) );
  OR2_X1 U1146 ( .A1(n1204), .A2(n1205), .ZN(n1203) );
  INV_X1 U1147 ( .A(n1206), .ZN(n1204) );
  AND2_X1 U1148 ( .A1(n1207), .A2(n733), .ZN(n1201) );
  INV_X1 U1149 ( .A(n727), .ZN(n733) );
  OR2_X1 U1150 ( .A1(Result_9_), .A2(n1208), .ZN(n727) );
  AND2_X1 U1151 ( .A1(n1209), .A2(n1210), .ZN(n1208) );
  AND2_X1 U1152 ( .A1(n1211), .A2(n1212), .ZN(n1210) );
  AND2_X1 U1153 ( .A1(n1213), .A2(n1214), .ZN(n1212) );
  AND2_X1 U1154 ( .A1(n1215), .A2(n1216), .ZN(n1214) );
  AND2_X1 U1155 ( .A1(n736), .A2(n1217), .ZN(n1216) );
  AND2_X1 U1156 ( .A1(n766), .A2(n750), .ZN(n1215) );
  AND2_X1 U1157 ( .A1(n1218), .A2(n1219), .ZN(n1213) );
  AND2_X1 U1158 ( .A1(n798), .A2(n782), .ZN(n1219) );
  AND2_X1 U1159 ( .A1(n830), .A2(n814), .ZN(n1218) );
  AND2_X1 U1160 ( .A1(n1220), .A2(n1221), .ZN(n1211) );
  AND2_X1 U1161 ( .A1(n1222), .A2(n1223), .ZN(n1221) );
  AND2_X1 U1162 ( .A1(n862), .A2(n846), .ZN(n1223) );
  AND2_X1 U1163 ( .A1(n894), .A2(n878), .ZN(n1222) );
  AND2_X1 U1164 ( .A1(n1224), .A2(n1225), .ZN(n1220) );
  AND2_X1 U1165 ( .A1(n926), .A2(n910), .ZN(n1225) );
  AND2_X1 U1166 ( .A1(n958), .A2(n942), .ZN(n1224) );
  AND2_X1 U1167 ( .A1(n1226), .A2(n1227), .ZN(n1209) );
  AND2_X1 U1168 ( .A1(n1228), .A2(n1229), .ZN(n1227) );
  AND2_X1 U1169 ( .A1(n1230), .A2(n1231), .ZN(n1229) );
  AND2_X1 U1170 ( .A1(n990), .A2(n974), .ZN(n1231) );
  AND2_X1 U1171 ( .A1(n1022), .A2(n1006), .ZN(n1230) );
  AND2_X1 U1172 ( .A1(n1232), .A2(n1233), .ZN(n1228) );
  AND2_X1 U1173 ( .A1(n1054), .A2(n1038), .ZN(n1233) );
  AND2_X1 U1174 ( .A1(n1086), .A2(n1070), .ZN(n1232) );
  AND2_X1 U1175 ( .A1(n1234), .A2(n1235), .ZN(n1226) );
  AND2_X1 U1176 ( .A1(n1236), .A2(n1237), .ZN(n1235) );
  AND2_X1 U1177 ( .A1(n1118), .A2(n1102), .ZN(n1237) );
  AND2_X1 U1178 ( .A1(n1150), .A2(n1134), .ZN(n1236) );
  AND2_X1 U1179 ( .A1(n1238), .A2(n1239), .ZN(n1234) );
  AND2_X1 U1180 ( .A1(n1182), .A2(n1166), .ZN(n1239) );
  AND2_X1 U1181 ( .A1(n718), .A2(n1198), .ZN(n1238) );
  OR2_X1 U1182 ( .A1(a_31_), .A2(n1240), .ZN(n718) );
  AND2_X1 U1183 ( .A1(n1206), .A2(n1217), .ZN(n1241) );
  OR2_X1 U1184 ( .A1(n1243), .A2(n1244), .ZN(n1206) );
  AND2_X1 U1185 ( .A1(a_1_), .A2(n1245), .ZN(n1244) );
  AND2_X1 U1186 ( .A1(n1198), .A2(n1191), .ZN(n1243) );
  OR2_X1 U1187 ( .A1(n1246), .A2(n1247), .ZN(n1191) );
  AND2_X1 U1188 ( .A1(a_2_), .A2(n1248), .ZN(n1247) );
  AND2_X1 U1189 ( .A1(n1182), .A2(n1175), .ZN(n1246) );
  OR2_X1 U1190 ( .A1(n1249), .A2(n1250), .ZN(n1175) );
  AND2_X1 U1191 ( .A1(a_3_), .A2(n1251), .ZN(n1250) );
  AND2_X1 U1192 ( .A1(n1166), .A2(n1159), .ZN(n1249) );
  OR2_X1 U1193 ( .A1(n1252), .A2(n1253), .ZN(n1159) );
  AND2_X1 U1194 ( .A1(a_4_), .A2(n1254), .ZN(n1253) );
  AND2_X1 U1195 ( .A1(n1150), .A2(n1143), .ZN(n1252) );
  OR2_X1 U1196 ( .A1(n1255), .A2(n1256), .ZN(n1143) );
  AND2_X1 U1197 ( .A1(a_5_), .A2(n1257), .ZN(n1256) );
  AND2_X1 U1198 ( .A1(n1134), .A2(n1127), .ZN(n1255) );
  OR2_X1 U1199 ( .A1(n1258), .A2(n1259), .ZN(n1127) );
  AND2_X1 U1200 ( .A1(a_6_), .A2(n1260), .ZN(n1259) );
  AND2_X1 U1201 ( .A1(n1118), .A2(n1111), .ZN(n1258) );
  OR2_X1 U1202 ( .A1(n1261), .A2(n1262), .ZN(n1111) );
  AND2_X1 U1203 ( .A1(a_7_), .A2(n1263), .ZN(n1262) );
  AND2_X1 U1204 ( .A1(n1102), .A2(n1095), .ZN(n1261) );
  OR2_X1 U1205 ( .A1(n1264), .A2(n1265), .ZN(n1095) );
  AND2_X1 U1206 ( .A1(a_8_), .A2(n1266), .ZN(n1265) );
  AND2_X1 U1207 ( .A1(n1086), .A2(n1079), .ZN(n1264) );
  OR2_X1 U1208 ( .A1(n1267), .A2(n1268), .ZN(n1079) );
  AND2_X1 U1209 ( .A1(a_9_), .A2(n1269), .ZN(n1268) );
  AND2_X1 U1210 ( .A1(n1070), .A2(n1063), .ZN(n1267) );
  OR2_X1 U1211 ( .A1(n1270), .A2(n1271), .ZN(n1063) );
  AND2_X1 U1212 ( .A1(a_10_), .A2(n1272), .ZN(n1271) );
  AND2_X1 U1213 ( .A1(n1054), .A2(n1047), .ZN(n1270) );
  OR2_X1 U1214 ( .A1(n1273), .A2(n1274), .ZN(n1047) );
  AND2_X1 U1215 ( .A1(a_11_), .A2(n1275), .ZN(n1274) );
  AND2_X1 U1216 ( .A1(n1038), .A2(n1031), .ZN(n1273) );
  OR2_X1 U1217 ( .A1(n1276), .A2(n1277), .ZN(n1031) );
  AND2_X1 U1218 ( .A1(a_12_), .A2(n1278), .ZN(n1277) );
  AND2_X1 U1219 ( .A1(n1022), .A2(n1015), .ZN(n1276) );
  OR2_X1 U1220 ( .A1(n1279), .A2(n1280), .ZN(n1015) );
  AND2_X1 U1221 ( .A1(a_13_), .A2(n1281), .ZN(n1280) );
  AND2_X1 U1222 ( .A1(n1006), .A2(n999), .ZN(n1279) );
  OR2_X1 U1223 ( .A1(n1282), .A2(n1283), .ZN(n999) );
  AND2_X1 U1224 ( .A1(a_14_), .A2(n1284), .ZN(n1283) );
  AND2_X1 U1225 ( .A1(n990), .A2(n983), .ZN(n1282) );
  OR2_X1 U1226 ( .A1(n1285), .A2(n1286), .ZN(n983) );
  AND2_X1 U1227 ( .A1(a_15_), .A2(n1287), .ZN(n1286) );
  AND2_X1 U1228 ( .A1(n974), .A2(n967), .ZN(n1285) );
  OR2_X1 U1229 ( .A1(n1288), .A2(n1289), .ZN(n967) );
  AND2_X1 U1230 ( .A1(a_16_), .A2(n1290), .ZN(n1289) );
  AND2_X1 U1231 ( .A1(n958), .A2(n951), .ZN(n1288) );
  OR2_X1 U1232 ( .A1(n1291), .A2(n1292), .ZN(n951) );
  AND2_X1 U1233 ( .A1(a_17_), .A2(n1293), .ZN(n1292) );
  AND2_X1 U1234 ( .A1(n942), .A2(n935), .ZN(n1291) );
  OR2_X1 U1235 ( .A1(n1294), .A2(n1295), .ZN(n935) );
  AND2_X1 U1236 ( .A1(a_18_), .A2(n1296), .ZN(n1295) );
  AND2_X1 U1237 ( .A1(n926), .A2(n919), .ZN(n1294) );
  OR2_X1 U1238 ( .A1(n1297), .A2(n1298), .ZN(n919) );
  AND2_X1 U1239 ( .A1(a_19_), .A2(n1299), .ZN(n1298) );
  AND2_X1 U1240 ( .A1(n910), .A2(n903), .ZN(n1297) );
  OR2_X1 U1241 ( .A1(n1300), .A2(n1301), .ZN(n903) );
  AND2_X1 U1242 ( .A1(a_20_), .A2(n1302), .ZN(n1301) );
  AND2_X1 U1243 ( .A1(n894), .A2(n887), .ZN(n1300) );
  OR2_X1 U1244 ( .A1(n1303), .A2(n1304), .ZN(n887) );
  AND2_X1 U1245 ( .A1(a_21_), .A2(n1305), .ZN(n1304) );
  AND2_X1 U1246 ( .A1(n878), .A2(n871), .ZN(n1303) );
  OR2_X1 U1247 ( .A1(n1306), .A2(n1307), .ZN(n871) );
  AND2_X1 U1248 ( .A1(a_22_), .A2(n1308), .ZN(n1307) );
  AND2_X1 U1249 ( .A1(n862), .A2(n855), .ZN(n1306) );
  OR2_X1 U1250 ( .A1(n1309), .A2(n1310), .ZN(n855) );
  AND2_X1 U1251 ( .A1(a_23_), .A2(n1311), .ZN(n1310) );
  AND2_X1 U1252 ( .A1(n846), .A2(n839), .ZN(n1309) );
  OR2_X1 U1253 ( .A1(n1312), .A2(n1313), .ZN(n839) );
  AND2_X1 U1254 ( .A1(a_24_), .A2(n1314), .ZN(n1313) );
  AND2_X1 U1255 ( .A1(n830), .A2(n823), .ZN(n1312) );
  OR2_X1 U1256 ( .A1(n1315), .A2(n1316), .ZN(n823) );
  AND2_X1 U1257 ( .A1(a_25_), .A2(n1317), .ZN(n1316) );
  AND2_X1 U1258 ( .A1(n814), .A2(n807), .ZN(n1315) );
  OR2_X1 U1259 ( .A1(n1318), .A2(n1319), .ZN(n807) );
  AND2_X1 U1260 ( .A1(a_26_), .A2(n1320), .ZN(n1319) );
  AND2_X1 U1261 ( .A1(n798), .A2(n791), .ZN(n1318) );
  OR2_X1 U1262 ( .A1(n1321), .A2(n1322), .ZN(n791) );
  AND2_X1 U1263 ( .A1(a_27_), .A2(n1323), .ZN(n1322) );
  AND2_X1 U1264 ( .A1(n782), .A2(n775), .ZN(n1321) );
  OR2_X1 U1265 ( .A1(n1324), .A2(n1325), .ZN(n775) );
  AND2_X1 U1266 ( .A1(a_28_), .A2(n1326), .ZN(n1325) );
  AND2_X1 U1267 ( .A1(n766), .A2(n759), .ZN(n1324) );
  OR2_X1 U1268 ( .A1(n1327), .A2(n1328), .ZN(n759) );
  AND2_X1 U1269 ( .A1(a_29_), .A2(n1329), .ZN(n1328) );
  AND2_X1 U1270 ( .A1(n750), .A2(n743), .ZN(n1327) );
  OR2_X1 U1271 ( .A1(n1330), .A2(n734), .ZN(n743) );
  AND2_X1 U1272 ( .A1(n1331), .A2(a_30_), .ZN(n734) );
  AND2_X1 U1273 ( .A1(n725), .A2(n736), .ZN(n1330) );
  OR2_X1 U1274 ( .A1(a_30_), .A2(n1331), .ZN(n736) );
  INV_X1 U1275 ( .A(b_30_), .ZN(n1331) );
  AND2_X1 U1276 ( .A1(n1240), .A2(a_31_), .ZN(n725) );
  INV_X1 U1277 ( .A(b_31_), .ZN(n1240) );
  OR2_X1 U1278 ( .A1(a_29_), .A2(n1329), .ZN(n750) );
  OR2_X1 U1279 ( .A1(a_28_), .A2(n1326), .ZN(n766) );
  OR2_X1 U1280 ( .A1(a_27_), .A2(n1323), .ZN(n782) );
  OR2_X1 U1281 ( .A1(a_26_), .A2(n1320), .ZN(n798) );
  OR2_X1 U1282 ( .A1(a_25_), .A2(n1317), .ZN(n814) );
  OR2_X1 U1283 ( .A1(a_24_), .A2(n1314), .ZN(n830) );
  OR2_X1 U1284 ( .A1(a_23_), .A2(n1311), .ZN(n846) );
  OR2_X1 U1285 ( .A1(a_22_), .A2(n1308), .ZN(n862) );
  OR2_X1 U1286 ( .A1(a_21_), .A2(n1305), .ZN(n878) );
  OR2_X1 U1287 ( .A1(a_20_), .A2(n1302), .ZN(n894) );
  OR2_X1 U1288 ( .A1(a_19_), .A2(n1299), .ZN(n910) );
  OR2_X1 U1289 ( .A1(a_18_), .A2(n1296), .ZN(n926) );
  OR2_X1 U1290 ( .A1(a_17_), .A2(n1293), .ZN(n942) );
  OR2_X1 U1291 ( .A1(a_16_), .A2(n1290), .ZN(n958) );
  OR2_X1 U1292 ( .A1(a_15_), .A2(n1287), .ZN(n974) );
  OR2_X1 U1293 ( .A1(a_14_), .A2(n1284), .ZN(n990) );
  OR2_X1 U1294 ( .A1(a_13_), .A2(n1281), .ZN(n1006) );
  OR2_X1 U1295 ( .A1(a_12_), .A2(n1278), .ZN(n1022) );
  OR2_X1 U1296 ( .A1(a_11_), .A2(n1275), .ZN(n1038) );
  OR2_X1 U1297 ( .A1(a_10_), .A2(n1272), .ZN(n1054) );
  OR2_X1 U1298 ( .A1(a_9_), .A2(n1269), .ZN(n1070) );
  OR2_X1 U1299 ( .A1(a_8_), .A2(n1266), .ZN(n1086) );
  OR2_X1 U1300 ( .A1(a_7_), .A2(n1263), .ZN(n1102) );
  OR2_X1 U1301 ( .A1(a_6_), .A2(n1260), .ZN(n1118) );
  OR2_X1 U1302 ( .A1(a_5_), .A2(n1257), .ZN(n1134) );
  OR2_X1 U1303 ( .A1(a_4_), .A2(n1254), .ZN(n1150) );
  OR2_X1 U1304 ( .A1(a_3_), .A2(n1251), .ZN(n1166) );
  OR2_X1 U1305 ( .A1(a_2_), .A2(n1248), .ZN(n1182) );
  OR2_X1 U1306 ( .A1(a_1_), .A2(n1245), .ZN(n1198) );
  AND2_X1 U1307 ( .A1(n1332), .A2(n1333), .ZN(n1207) );
  INV_X1 U1308 ( .A(n1334), .ZN(n1333) );
  AND2_X1 U1309 ( .A1(n1335), .A2(n1205), .ZN(n1334) );
  OR2_X1 U1310 ( .A1(n1205), .A2(n1335), .ZN(n1332) );
  OR2_X1 U1311 ( .A1(n1336), .A2(n1337), .ZN(n1335) );
  AND2_X1 U1312 ( .A1(n1197), .A2(n1200), .ZN(n1337) );
  AND2_X1 U1313 ( .A1(n1338), .A2(n1245), .ZN(n1336) );
  INV_X1 U1314 ( .A(b_1_), .ZN(n1245) );
  OR2_X1 U1315 ( .A1(n1200), .A2(n1197), .ZN(n1338) );
  OR2_X1 U1316 ( .A1(n1339), .A2(n1340), .ZN(n1197) );
  AND2_X1 U1317 ( .A1(n1181), .A2(n1184), .ZN(n1340) );
  AND2_X1 U1318 ( .A1(n1341), .A2(n1248), .ZN(n1339) );
  INV_X1 U1319 ( .A(b_2_), .ZN(n1248) );
  OR2_X1 U1320 ( .A1(n1184), .A2(n1181), .ZN(n1341) );
  OR2_X1 U1321 ( .A1(n1342), .A2(n1343), .ZN(n1181) );
  AND2_X1 U1322 ( .A1(n1165), .A2(n1168), .ZN(n1343) );
  AND2_X1 U1323 ( .A1(n1344), .A2(n1251), .ZN(n1342) );
  INV_X1 U1324 ( .A(b_3_), .ZN(n1251) );
  OR2_X1 U1325 ( .A1(n1168), .A2(n1165), .ZN(n1344) );
  OR2_X1 U1326 ( .A1(n1345), .A2(n1346), .ZN(n1165) );
  AND2_X1 U1327 ( .A1(n1149), .A2(n1152), .ZN(n1346) );
  AND2_X1 U1328 ( .A1(n1347), .A2(n1254), .ZN(n1345) );
  INV_X1 U1329 ( .A(b_4_), .ZN(n1254) );
  OR2_X1 U1330 ( .A1(n1152), .A2(n1149), .ZN(n1347) );
  OR2_X1 U1331 ( .A1(n1348), .A2(n1349), .ZN(n1149) );
  AND2_X1 U1332 ( .A1(n1133), .A2(n1136), .ZN(n1349) );
  AND2_X1 U1333 ( .A1(n1350), .A2(n1257), .ZN(n1348) );
  INV_X1 U1334 ( .A(b_5_), .ZN(n1257) );
  OR2_X1 U1335 ( .A1(n1136), .A2(n1133), .ZN(n1350) );
  OR2_X1 U1336 ( .A1(n1351), .A2(n1352), .ZN(n1133) );
  AND2_X1 U1337 ( .A1(n1117), .A2(n1120), .ZN(n1352) );
  AND2_X1 U1338 ( .A1(n1353), .A2(n1260), .ZN(n1351) );
  INV_X1 U1339 ( .A(b_6_), .ZN(n1260) );
  OR2_X1 U1340 ( .A1(n1120), .A2(n1117), .ZN(n1353) );
  OR2_X1 U1341 ( .A1(n1354), .A2(n1355), .ZN(n1117) );
  AND2_X1 U1342 ( .A1(n1101), .A2(n1104), .ZN(n1355) );
  AND2_X1 U1343 ( .A1(n1356), .A2(n1263), .ZN(n1354) );
  INV_X1 U1344 ( .A(b_7_), .ZN(n1263) );
  OR2_X1 U1345 ( .A1(n1104), .A2(n1101), .ZN(n1356) );
  OR2_X1 U1346 ( .A1(n1357), .A2(n1358), .ZN(n1101) );
  AND2_X1 U1347 ( .A1(n1085), .A2(n1088), .ZN(n1358) );
  AND2_X1 U1348 ( .A1(n1359), .A2(n1266), .ZN(n1357) );
  INV_X1 U1349 ( .A(b_8_), .ZN(n1266) );
  OR2_X1 U1350 ( .A1(n1088), .A2(n1085), .ZN(n1359) );
  OR2_X1 U1351 ( .A1(n1360), .A2(n1361), .ZN(n1085) );
  AND2_X1 U1352 ( .A1(n1069), .A2(n1072), .ZN(n1361) );
  AND2_X1 U1353 ( .A1(n1362), .A2(n1269), .ZN(n1360) );
  INV_X1 U1354 ( .A(b_9_), .ZN(n1269) );
  OR2_X1 U1355 ( .A1(n1072), .A2(n1069), .ZN(n1362) );
  OR2_X1 U1356 ( .A1(n1363), .A2(n1364), .ZN(n1069) );
  AND2_X1 U1357 ( .A1(n1053), .A2(n1056), .ZN(n1364) );
  AND2_X1 U1358 ( .A1(n1365), .A2(n1272), .ZN(n1363) );
  INV_X1 U1359 ( .A(b_10_), .ZN(n1272) );
  OR2_X1 U1360 ( .A1(n1056), .A2(n1053), .ZN(n1365) );
  OR2_X1 U1361 ( .A1(n1366), .A2(n1367), .ZN(n1053) );
  AND2_X1 U1362 ( .A1(n1037), .A2(n1040), .ZN(n1367) );
  AND2_X1 U1363 ( .A1(n1368), .A2(n1275), .ZN(n1366) );
  INV_X1 U1364 ( .A(b_11_), .ZN(n1275) );
  OR2_X1 U1365 ( .A1(n1040), .A2(n1037), .ZN(n1368) );
  OR2_X1 U1366 ( .A1(n1369), .A2(n1370), .ZN(n1037) );
  AND2_X1 U1367 ( .A1(n1021), .A2(n1024), .ZN(n1370) );
  AND2_X1 U1368 ( .A1(n1371), .A2(n1278), .ZN(n1369) );
  INV_X1 U1369 ( .A(b_12_), .ZN(n1278) );
  OR2_X1 U1370 ( .A1(n1024), .A2(n1021), .ZN(n1371) );
  OR2_X1 U1371 ( .A1(n1372), .A2(n1373), .ZN(n1021) );
  AND2_X1 U1372 ( .A1(n1005), .A2(n1008), .ZN(n1373) );
  AND2_X1 U1373 ( .A1(n1374), .A2(n1281), .ZN(n1372) );
  INV_X1 U1374 ( .A(b_13_), .ZN(n1281) );
  OR2_X1 U1375 ( .A1(n1008), .A2(n1005), .ZN(n1374) );
  OR2_X1 U1376 ( .A1(n1375), .A2(n1376), .ZN(n1005) );
  AND2_X1 U1377 ( .A1(n989), .A2(n992), .ZN(n1376) );
  AND2_X1 U1378 ( .A1(n1377), .A2(n1284), .ZN(n1375) );
  INV_X1 U1379 ( .A(b_14_), .ZN(n1284) );
  OR2_X1 U1380 ( .A1(n992), .A2(n989), .ZN(n1377) );
  OR2_X1 U1381 ( .A1(n1378), .A2(n1379), .ZN(n989) );
  AND2_X1 U1382 ( .A1(n973), .A2(n976), .ZN(n1379) );
  AND2_X1 U1383 ( .A1(n1380), .A2(n1287), .ZN(n1378) );
  INV_X1 U1384 ( .A(b_15_), .ZN(n1287) );
  OR2_X1 U1385 ( .A1(n976), .A2(n973), .ZN(n1380) );
  OR2_X1 U1386 ( .A1(n1381), .A2(n1382), .ZN(n973) );
  AND2_X1 U1387 ( .A1(n957), .A2(n960), .ZN(n1382) );
  AND2_X1 U1388 ( .A1(n1383), .A2(n1290), .ZN(n1381) );
  INV_X1 U1389 ( .A(b_16_), .ZN(n1290) );
  OR2_X1 U1390 ( .A1(n960), .A2(n957), .ZN(n1383) );
  OR2_X1 U1391 ( .A1(n1384), .A2(n1385), .ZN(n957) );
  AND2_X1 U1392 ( .A1(n941), .A2(n944), .ZN(n1385) );
  AND2_X1 U1393 ( .A1(n1386), .A2(n1293), .ZN(n1384) );
  INV_X1 U1394 ( .A(b_17_), .ZN(n1293) );
  OR2_X1 U1395 ( .A1(n944), .A2(n941), .ZN(n1386) );
  OR2_X1 U1396 ( .A1(n1387), .A2(n1388), .ZN(n941) );
  AND2_X1 U1397 ( .A1(n925), .A2(n928), .ZN(n1388) );
  AND2_X1 U1398 ( .A1(n1389), .A2(n1296), .ZN(n1387) );
  INV_X1 U1399 ( .A(b_18_), .ZN(n1296) );
  OR2_X1 U1400 ( .A1(n928), .A2(n925), .ZN(n1389) );
  OR2_X1 U1401 ( .A1(n1390), .A2(n1391), .ZN(n925) );
  AND2_X1 U1402 ( .A1(n909), .A2(n912), .ZN(n1391) );
  AND2_X1 U1403 ( .A1(n1392), .A2(n1299), .ZN(n1390) );
  INV_X1 U1404 ( .A(b_19_), .ZN(n1299) );
  OR2_X1 U1405 ( .A1(n912), .A2(n909), .ZN(n1392) );
  OR2_X1 U1406 ( .A1(n1393), .A2(n1394), .ZN(n909) );
  AND2_X1 U1407 ( .A1(n893), .A2(n896), .ZN(n1394) );
  AND2_X1 U1408 ( .A1(n1395), .A2(n1302), .ZN(n1393) );
  INV_X1 U1409 ( .A(b_20_), .ZN(n1302) );
  OR2_X1 U1410 ( .A1(n896), .A2(n893), .ZN(n1395) );
  OR2_X1 U1411 ( .A1(n1396), .A2(n1397), .ZN(n893) );
  AND2_X1 U1412 ( .A1(n877), .A2(n880), .ZN(n1397) );
  AND2_X1 U1413 ( .A1(n1398), .A2(n1305), .ZN(n1396) );
  INV_X1 U1414 ( .A(b_21_), .ZN(n1305) );
  OR2_X1 U1415 ( .A1(n880), .A2(n877), .ZN(n1398) );
  OR2_X1 U1416 ( .A1(n1399), .A2(n1400), .ZN(n877) );
  AND2_X1 U1417 ( .A1(n861), .A2(n864), .ZN(n1400) );
  AND2_X1 U1418 ( .A1(n1401), .A2(n1308), .ZN(n1399) );
  INV_X1 U1419 ( .A(b_22_), .ZN(n1308) );
  OR2_X1 U1420 ( .A1(n864), .A2(n861), .ZN(n1401) );
  OR2_X1 U1421 ( .A1(n1402), .A2(n1403), .ZN(n861) );
  AND2_X1 U1422 ( .A1(n845), .A2(n848), .ZN(n1403) );
  AND2_X1 U1423 ( .A1(n1404), .A2(n1311), .ZN(n1402) );
  INV_X1 U1424 ( .A(b_23_), .ZN(n1311) );
  OR2_X1 U1425 ( .A1(n848), .A2(n845), .ZN(n1404) );
  OR2_X1 U1426 ( .A1(n1405), .A2(n1406), .ZN(n845) );
  AND2_X1 U1427 ( .A1(n829), .A2(n832), .ZN(n1406) );
  AND2_X1 U1428 ( .A1(n1407), .A2(n1314), .ZN(n1405) );
  INV_X1 U1429 ( .A(b_24_), .ZN(n1314) );
  OR2_X1 U1430 ( .A1(n832), .A2(n829), .ZN(n1407) );
  OR2_X1 U1431 ( .A1(n1408), .A2(n1409), .ZN(n829) );
  AND2_X1 U1432 ( .A1(n813), .A2(n816), .ZN(n1409) );
  AND2_X1 U1433 ( .A1(n1410), .A2(n1317), .ZN(n1408) );
  INV_X1 U1434 ( .A(b_25_), .ZN(n1317) );
  OR2_X1 U1435 ( .A1(n816), .A2(n813), .ZN(n1410) );
  OR2_X1 U1436 ( .A1(n1411), .A2(n1412), .ZN(n813) );
  AND2_X1 U1437 ( .A1(n797), .A2(n800), .ZN(n1412) );
  AND2_X1 U1438 ( .A1(n1413), .A2(n1320), .ZN(n1411) );
  INV_X1 U1439 ( .A(b_26_), .ZN(n1320) );
  OR2_X1 U1440 ( .A1(n800), .A2(n797), .ZN(n1413) );
  OR2_X1 U1441 ( .A1(n1414), .A2(n1415), .ZN(n797) );
  AND2_X1 U1442 ( .A1(n781), .A2(n784), .ZN(n1415) );
  AND2_X1 U1443 ( .A1(n1416), .A2(n1323), .ZN(n1414) );
  INV_X1 U1444 ( .A(b_27_), .ZN(n1323) );
  OR2_X1 U1445 ( .A1(n784), .A2(n781), .ZN(n1416) );
  OR2_X1 U1446 ( .A1(n1417), .A2(n1418), .ZN(n781) );
  AND2_X1 U1447 ( .A1(n765), .A2(n768), .ZN(n1418) );
  AND2_X1 U1448 ( .A1(n1419), .A2(n1326), .ZN(n1417) );
  INV_X1 U1449 ( .A(b_28_), .ZN(n1326) );
  OR2_X1 U1450 ( .A1(n768), .A2(n765), .ZN(n1419) );
  OR2_X1 U1451 ( .A1(n1420), .A2(n1421), .ZN(n765) );
  AND2_X1 U1452 ( .A1(n1422), .A2(n752), .ZN(n1421) );
  AND2_X1 U1453 ( .A1(n1423), .A2(n1329), .ZN(n1420) );
  INV_X1 U1454 ( .A(b_29_), .ZN(n1329) );
  OR2_X1 U1455 ( .A1(n1422), .A2(n752), .ZN(n1423) );
  INV_X1 U1456 ( .A(a_29_), .ZN(n752) );
  INV_X1 U1457 ( .A(n749), .ZN(n1422) );
  OR2_X1 U1458 ( .A1(n1424), .A2(n1425), .ZN(n749) );
  AND2_X1 U1459 ( .A1(a_30_), .A2(b_30_), .ZN(n1425) );
  AND2_X1 U1460 ( .A1(n1426), .A2(b_31_), .ZN(n1424) );
  AND2_X1 U1461 ( .A1(a_31_), .A2(n1427), .ZN(n1426) );
  OR2_X1 U1462 ( .A1(a_30_), .A2(b_30_), .ZN(n1427) );
  INV_X1 U1463 ( .A(a_28_), .ZN(n768) );
  INV_X1 U1464 ( .A(a_27_), .ZN(n784) );
  INV_X1 U1465 ( .A(a_26_), .ZN(n800) );
  INV_X1 U1466 ( .A(a_25_), .ZN(n816) );
  INV_X1 U1467 ( .A(a_24_), .ZN(n832) );
  INV_X1 U1468 ( .A(a_23_), .ZN(n848) );
  INV_X1 U1469 ( .A(a_22_), .ZN(n864) );
  INV_X1 U1470 ( .A(a_21_), .ZN(n880) );
  INV_X1 U1471 ( .A(a_20_), .ZN(n896) );
  INV_X1 U1472 ( .A(a_19_), .ZN(n912) );
  INV_X1 U1473 ( .A(a_18_), .ZN(n928) );
  INV_X1 U1474 ( .A(a_17_), .ZN(n944) );
  INV_X1 U1475 ( .A(a_16_), .ZN(n960) );
  INV_X1 U1476 ( .A(a_15_), .ZN(n976) );
  INV_X1 U1477 ( .A(a_14_), .ZN(n992) );
  INV_X1 U1478 ( .A(a_13_), .ZN(n1008) );
  INV_X1 U1479 ( .A(a_12_), .ZN(n1024) );
  INV_X1 U1480 ( .A(a_11_), .ZN(n1040) );
  INV_X1 U1481 ( .A(a_10_), .ZN(n1056) );
  INV_X1 U1482 ( .A(a_9_), .ZN(n1072) );
  INV_X1 U1483 ( .A(a_8_), .ZN(n1088) );
  INV_X1 U1484 ( .A(a_7_), .ZN(n1104) );
  INV_X1 U1485 ( .A(a_6_), .ZN(n1120) );
  INV_X1 U1486 ( .A(a_5_), .ZN(n1136) );
  INV_X1 U1487 ( .A(a_4_), .ZN(n1152) );
  INV_X1 U1488 ( .A(a_3_), .ZN(n1168) );
  INV_X1 U1489 ( .A(a_2_), .ZN(n1184) );
  INV_X1 U1490 ( .A(a_1_), .ZN(n1200) );
  AND2_X1 U1491 ( .A1(n1217), .A2(n1428), .ZN(n1205) );
  INV_X1 U1492 ( .A(n1242), .ZN(n1428) );
  AND2_X1 U1493 ( .A1(a_0_), .A2(n1429), .ZN(n1242) );
  OR2_X1 U1494 ( .A1(a_0_), .A2(n1429), .ZN(n1217) );
  INV_X1 U1495 ( .A(b_0_), .ZN(n1429) );
endmodule

