module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g10722, g10664, g1289, g8943, g1882, n1663,
         g255, g312, g11257, g452, g7032, g123, g6830, g207, g8920, g713,
         g4340, g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695, g11372,
         g461, n1594, g8260, g940, g11391, g976, g8432, g709, n1719, g6088,
         g1092, g6478, g1574, g1864, g11320, g369, g6500, g1580, g5392, g1736,
         g10663, n1637, g10782, n3065, g6216, g1424, g1737, g10858, g1672,
         g5914, g1077, g7590, g1231, g6656, g4, g6728, g5126, g1104, n1658,
         g7290, g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064, g8019,
         g6545, g1543, g256, g315, g6533, g1534, g8820, g622, n1713, g8941,
         g1927, g10859, g1660, g6922, g278, g8772, g1436, g8433, g718, g6526,
         g10793, g554, g11333, g496, n1689, g11392, g981, g794, g829, g6093,
         g1095, g8889, g704, g7302, g1265, g6525, g1786, g8429, g682, g7292,
         g1296, g6621, g7134, n3062, g260, g327, g6333, g1389, n1603, g6826,
         g1371, g1955, g1956, g10860, g1675, g11483, g354, g6392, g113, g7626,
         g639, n1692, g10866, g1684, g8193, g1639, g6983, g1791, n1702, g6839,
         g248, g4076, g1707, g4293, g1759, g11482, g351, g6507, g1604, g6096,
         g1098, g8250, g932, g8282, g1896, g8435, g736, g6924, g1019, g6819,
         n3061, g746, g745, g6244, g1419, n1602, g6627, g32, n1865, g6071,
         g1086, g8046, g1486, g10707, g1730, g6198, g1504, g8051, g1470, g8024,
         g822, g10862, g1678, g8050, g174, g7133, g1766, g7930, g1801, g6832,
         g186, g11308, g959, g6918, g8769, g1407, g6909, g1868, g4940, g5404,
         g1718, n1611, g11265, g396, g6930, g1015, g10726, n1650, g4891, n3059,
         n1874, g6224, g1415, g7586, g1227, g10770, g1721, n3058, n3057, g6934,
         g284, g11256, g426, g6824, g219, g1360, n3056, g6126, g806, g8767,
         g1428, g6546, g1564, g4238, g1741, g6823, g225, g6928, g281, g11602,
         g1308, g9721, g611, n1609, g4890, n3055, n1586, g1217, g6524, g1589,
         g8045, g1466, g6469, g1571, g6471, g1861, g6821, n3054, g11514, g1448,
         g1133, n1706, g11610, g1333, g7843, g153, g11310, g962, g5536, g11331,
         g486, n1621, g11380, g471, n1606, g6838, g1397, g8288, g1950, g755,
         g756, n3053, g10855, g1101, g549, g10898, g105, g10865, g1669, g6822,
         g6528, g1531, g6180, g1458, g10718, g572, g6912, g1011, g10719, n3051,
         g6234, g1411, g6099, g1074, g11259, g444, g8039, g1474, g6059, g1080,
         g5396, g1713, n1610, g262, g333, g6906, g269, g11266, g401, g11294,
         g1857, n1682, g5421, g9, g8649, g664, g11312, g965, g6840, g1400,
         g254, g309, g7202, g814, g6834, g231, g10795, g557, g875, g869, g6831,
         g1383, g8060, g158, g4893, g627, g7244, g1023, g6026, g259, n3050,
         g11608, g1327, g654, g6911, g293, g11640, g1346, g8777, g1633, g4274,
         g1753, g1508, n1707, g7297, g1240, g11326, g538, g11269, g416, g11325,
         g542, g10864, g1681, g11290, g374, g10798, g563, g8284, g1914, g11328,
         g530, g10800, g575, g8944, g1936, n1694, g7183, g4465, g1356, g1317,
         g11484, g357, g11263, g386, g6501, g1601, g6757, g166, g11334, g501,
         n1690, g6042, g8384, g1840, g6653, g257, g318, g5849, n3048, g6929,
         g302, g11488, g342, g7299, g1250, g4330, g1163, g1958, n3047, g7257,
         g1032, g8775, g1432, g5770, g1453, n1628, g11486, g363, g261, g330,
         g4338, g1157, g4500, n3046, g10721, n3045, g8147, g928, g6038, g11337,
         g516, n1620, g6045, g7191, g826, g861, g8774, g1627, g7293, g1292,
         g6907, g290, g4903, n3044, n1873, g6123, g6506, g1583, g11376, g466,
         n1646, g6542, g1561, g6551, g1546, g6901, g287, g10797, g560, g8505,
         g617, n1645, n1631, g11647, g336, g11340, g456, n1641, g253, g305,
         n1681, g11625, g345, g636, g8, g6502, N599, g6049, g8945, g1945,
         n1697, g4231, g1738, g8040, g1478, n3042, g6155, g1690, n1653, g8043,
         g1482, g5173, g1110, n1677, g6916, g296, g10861, g1663, g8431, g700,
         g4309, g1762, g11485, g360, g6334, g192, g10767, g1657, g8923, g722,
         n1693, g7189, g10799, g566, g6747, n3041, g6080, g1089, g3381, g5910,
         g1071, g11393, g986, g11349, g971, g6439, g143, g9266, g1814, n1608,
         g1212, g8940, g1918, g9269, g1822, n1643, g6820, g237, g8042, g1462,
         g6759, g178, g11487, g366, g802, g837, g9124, g599, n1644, g11293,
         g1854, g11298, g944, g8287, g1941, g8047, g170, g6205, g1520, g8885,
         g686, n1676, g11305, g953, n3040, g2478, g1765, g10711, g1733, g7303,
         g5194, g1610, g7541, g1796, n1626, g11607, g1324, g6541, g1540, g6827,
         n3038, g11332, g491, n1691, g4902, n3037, g6828, g213, g6516, g1781,
         n1659, g8938, g1900, n1675, g7298, g1245, n3036, g6672, n3035, g8048,
         g148, g798, g833, g8285, g1923, g8254, g936, g11604, g1314, g849,
         g11636, g1336, g6910, g272, g8173, g1806, g8245, n1716, g8281, g1887,
         g10724, n3034, g11314, g968, g4905, n3033, g4484, g1137, g8937, g1891,
         n1657, g7300, g1255, g6002, n1588, g874, g9110, g591, n1607, g8926,
         g731, n1696, g8631, g7632, g1218, g9150, g605, n1593, g6531, g6786,
         g182, g11303, g950, g1129, n1705, g857, g11258, g448, g9272, g1828,
         n1605, g10773, g1727, g6470, g1592, g5083, g1703, g8286, g1932, g8773,
         g1624, g6054, g11260, g440, g11338, g476, n1599, g5918, g119, n1613,
         g8922, g668, n1662, g8049, g139, g4342, g1149, n1685, g10720, n3031,
         g6755, n3030, g6897, g263, g7709, g818, g4255, g1747, g5543, n1622,
         g6915, g275, g6513, g1524, g6480, g1577, g6733, g810, g11264, g391,
         g8973, g658, n1615, g6833, g1386, g5996, n1587, g1125, n1708, g5755,
         g201, n1619, g7295, g1280, n1862, g6068, g1083, g7137, g650, n1709,
         g8779, g1636, g853, g11270, g421, g5529, g11306, g956, g11291, g378,
         g4283, g1756, g841, g6894, g1027, g6902, g1003, g8765, g1403, g4498,
         g1145, g5148, g1107, n1614, g7581, g1223, g11267, g406, g10936, g1811,
         n1699, g10784, n3029, g10765, g1654, g6332, g197, n1678, g6479, g1595,
         g6537, g1537, g8434, g727, g6908, g6243, n1717, g11324, g481, n1680,
         n1647, g11609, g1330, g845, g8244, g8194, g1512, n3027, DFF_436_n1,
         g8052, g1490, g4325, g1166, g11481, g348, n3026, g7301, g1260, g6035,
         g8059, g131, n3025, g6015, g258, g11330, g521, n1698, g11605, g1318,
         g8921, g1872, n1616, g8883, g677, n1656, n3024, g6523, g1549, g11300,
         g947, g9555, g1834, n1655, g6481, g1598, g1121, g11606, g1321, g11335,
         g506, n1600, g10791, g546, g8939, g1909, g6529, g1552, g10776, g1687,
         g6514, g1586, g324, g1141, n1660, g11639, g1341, g4089, g1710, g10785,
         n3023, g6179, n3022, g8053, g135, g11329, g525, n1695, g6515, g1607,
         g321, g7204, g11443, g1275, g11603, g8770, g1615, g11292, g382, g6331,
         n3020, g6900, g266, g7294, g1284, n1864, g6829, n3019, g8428, g673,
         n3018, g8054, g162, g11268, g411, g11262, g431, n1876, g8283, g1905,
         g6193, g1515, n1627, g8776, g1630, g7143, g6898, g991, g7291, g1300,
         g11478, g339, g6000, g4264, g1750, g8768, g1440, g10863, g1666, g6522,
         g1528, g11641, g1351, n1721, g10780, n3017, g8044, g127, n1704,
         g11579, g1618, g7296, g1235, g6923, g299, g11261, g435, n1878, g6638,
         g6534, g1555, g6895, g995, g8771, g1621, g4506, n3016, g643, n1612,
         g8055, g1494, g6468, g1567, g8430, g691, g11327, g534, g6508, g1776,
         n1715, g10717, g569, g4334, g1160, n1585, g6679, g1, g11336, g511,
         n1679, g10771, g1724, g5445, g12, g8559, g1878, g7219, g5390, n1654,
         n1512, n1574, n1486, n1485, n1544, n1545, n1548, n1530, n1420, n1855,
         n1566, n1567, n1479, n1858, n1480, n1478, n1137, n1195, n1404, n1229,
         n1227, n1450, n916, n822, n809, n958, n918, n1159, n812, n1056, n817,
         n837, n804, n1380, n926, n1385, n1391, n1564, n1231, n1226, n1232,
         n1260, n1132, n1107, n1154, n1093, n1214, n931, n962, n1147, n1193,
         n1153, n1125, n1099, n917, n806, n808, n1097, n1123, n1151, n1090,
         n1161, n967, n921, n898, n1055, n938, n1150, n1096, n1098, n1213,
         n1152, n836, Tg1_OUT1, Tg1_OUT2, Tg1_OUT3, Tg1_OUT4, Tg1_OUT5,
         Tg1_OUT6, Tg1_OUT7, Tg1_OUT8, Tg2_OUT1, Tg2_OUT2, Tg2_OUT3, Tg2_OUT4,
         Tg2_OUT5, Tg2_OUT6, Tg2_OUT7, Tg2_OUT8, test_se_NOT, Trigger_select,
         n1, n7, n12, n40, n42, n45, n46, n57, n68, n84, n86, n106, n112, n113,
         n114, n118, n119, n124, n155, n167, n192, n227, n257, n274, n319,
         n324, n363, n369, n371, n395, n435, n443, n491, n493, n505, n507,
         n510, n517, n2199, n2200, n2201, n2279, n2322, n2323, n2326, n2329,
         n2330, n2331, n2333, n2334, n2335, n2336, n2337, n2343, n2344, n2345,
         n2347, n2348, n2352, n2353, n2354, n2355, n2356, n2358, n2360, n2362,
         n2363, n2364, n2365, n2366, n2367, n2369, n2373, n2374, n2375, n2376,
         n2378, n2380, n2383, n2391, n2392, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2431, n2432,
         n2433, n2434, n2435, n2436, n2439, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2468, n2469, n2471,
         n2472, n2473, n2474, n2476, n2477, n2478, n2482, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3021, n3028, n3032, n3039, n3043, n3049,
         n3052, n3060, n3063, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, U1586_n1, U1754_n1, U1798_n1, U1839_n1, U1843_n1, U1877_n1,
         U1908_n1, U1909_n1, U1987_n1, U2031_n1, U2035_n1, U2418_n1, U2468_n1,
         U2478_n1, U2488_n1, U2533_n1, U2534_n1, U2639_n1, U2641_n1, U2654_n1,
         U2658_n1, U2683_n1, U2699_n1, U2846_n1, U2847_n1, U2848_n1, U2859_n1,
         U2860_n1, U2861_n1, U2867_n1, U2879_n1, U2881_n1, U2882_n1, U2883_n1,
         U2884_n1, U2885_n1, U2886_n1, U2887_n1, U2888_n1, U2889_n1, U2890_n1,
         U2891_n1, U2892_n1, U2893_n1, U2894_n1, U2895_n1, U2896_n1, U2897_n1,
         U2898_n1, U2899_n1, U2900_n1, U2901_n1, U2902_n1, U3090_n1, U3092_n1,
         U3094_n1, U3096_n1, U3098_n1, U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(n1), .SI(test_si1), .SE(n2590), .CLK(n2630), .Q(
        g1289), .QN(n2391) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n2512), .CLK(n2669), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n2512), .CLK(n2669), .Q(g312), 
        .QN(n2367) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n2557), .CLK(n2646), .Q(g452) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n2508), .CLK(n2671), .Q(g123)
         );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n2565), .CLK(n2642), .Q(g207), 
        .QN(n2458) );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n2582), .CLK(n2634), .Q(g713), 
        .QN(n2445) );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n2582), .CLK(n2634), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n2522), .CLK(n2664), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n2519), .CLK(n2665), .Q(
        g1558) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n2567), .CLK(n2641), .Q(
        g695), .QN(n2419) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n2567), .CLK(n2641), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n2559), .CLK(n2645), .Q(g940) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n2577), .CLK(n2636), .Q(
        g976) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n2577), .CLK(n2636), .Q(g709), .QN(n1719) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n2562), .CLK(n2643), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n2538), .CLK(n2656), .Q(
        g1574) );
  SDFFX1 DFF_18_Q_reg ( .D(n68), .SI(g1574), .SE(n2509), .CLK(n2670), .Q(g1864), .QN(n2416) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n2548), .CLK(n2651), .Q(
        g369), .QN(n2489) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n2561), .CLK(n2644), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n2561), .CLK(n2644), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(n2561), .CLK(n2644), .Q(
        n1637) );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(n2561), .CLK(n2644), .Q(
        n3065), .QN(n4321) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n2561), .CLK(n2644), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n2561), .CLK(n2644), .Q(
        g1737), .QN(n2398) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n2544), .CLK(n2653), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n2569), .CLK(n2640), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n2590), .CLK(n2630), .Q(
        g1231), .QN(n2462) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n2586), .CLK(n2632), .Q(g4)
         );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(n2531), .CLK(n2659), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n2523), .CLK(n2663), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n2522), .CLK(n2663), .Q(
        g1304), .QN(n2337) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n2516), .CLK(n2667), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n2579), .CLK(n2635), .Q(
        g1499), .QN(n2365) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n2573), .CLK(n2638), .Q(
        g1444), .QN(n2405) );
  SDFFX1 DFF_37_Q_reg ( .D(n2490), .SI(g1444), .SE(n2573), .CLK(n2638), .Q(
        n3064) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n2521), .CLK(n2664), .Q(
        g4180), .QN(n2466) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n2519), .CLK(n2665), .Q(
        g1543) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n2510), .CLK(n2670), .Q(g315), .QN(n2378) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n2567), .CLK(n2641), .Q(
        g1534) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n2567), .CLK(n2641), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n2585), .CLK(n2632), .Q(
        g1927), .QN(n2444) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n2543), .CLK(n2653), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n2547), .CLK(n2651), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n2547), .CLK(n2651), .Q(
        g1436), .QN(n2402) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n2576), .CLK(n2636), .Q(
        g718), .QN(n2279) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n2550), .CLK(n2649), .Q(
        g8985) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n2543), .CLK(n2653), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n2541), .CLK(n2654), .Q(
        g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n2505), .CLK(n2672), .Q(
        g981) );
  SDFFX1 DFF_53_Q_reg ( .D(n2494), .SI(g981), .SE(n2580), .CLK(n2634), .Q(
        g3007) );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n2580), .CLK(n2634), .Q(
        test_so1), .QN(n2503) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n2551), .CLK(n2649), .Q(
        g829) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n2508), .CLK(n2670), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n2575), .CLK(n2637), .Q(
        g704), .QN(n2418) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n2575), .CLK(n2637), .Q(
        g1265), .QN(n2333) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n2530), .CLK(n2660), .Q(
        g1786), .QN(n2439) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n2530), .CLK(n2660), .Q(
        g682) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n2566), .CLK(n2642), .Q(
        g1296), .QN(n2335) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n2565), .CLK(n2642), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n2550), .CLK(n2649), .Q(
        g8977) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n2583), .CLK(n2633), .Q(
        n3062), .QN(n4311) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n2509), .CLK(n2670), .Q(g327), .QN(n2360) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n2588), .CLK(n2630), .Q(
        g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n2586), .CLK(n2631), .Q(
        g1371) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n2577), .CLK(n2636), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n2543), .CLK(n2653), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n2560), .CLK(n2645), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n2560), .CLK(n2645), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n2539), .CLK(n2655), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n2568), .CLK(n2641), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n2568), .CLK(n2641), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n2529), .CLK(n2660), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n2529), .CLK(n2660), .Q(
        g248) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n2529), .CLK(n2660), .Q(
        g1707), .QN(n2397) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n2527), .CLK(n2661), .Q(
        g1759) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n2567), .CLK(n2641), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n2566), .CLK(n2641), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n2566), .CLK(n2641), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n2539), .CLK(n2655), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n2539), .CLK(n2655), .Q(
        g932) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n2509), .CLK(n2670), .Q(
        g1896) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n2576), .CLK(n2636), .Q(
        g736) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n2539), .CLK(n2655), .Q(
        g1019), .QN(n2323) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n2539), .CLK(n2655), .Q(
        n3061) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n2538), .CLK(n2655), .Q(g745), .QN(n2464) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n2538), .CLK(n2655), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n2538), .CLK(n2655), .Q(
        g8979) );
  SDFFX1 DFF_92_Q_reg ( .D(n2491), .SI(g8979), .SE(n2581), .CLK(n2634), .Q(g32), .QN(n2199) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n2581), .CLK(n2634), .Q(n1865), .QN(n4317) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n2506), .CLK(n2672), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n2564), .CLK(n2642), .Q(
        g1486) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n2553), .CLK(n2648), .Q(
        g1730) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n2552), .CLK(n2648), .Q(
        g1504) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n2573), .CLK(n2638), .Q(
        g1470), .QN(n2413) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n2516), .CLK(n2666), .Q(
        g822), .QN(n2428) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n2515), .CLK(n2667), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n2507), .CLK(n2671), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n2547), .CLK(n2651), .Q(
        g174) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n2563), .CLK(n2643), .Q(
        g1766), .QN(n2461) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n2529), .CLK(n2660), .Q(
        g1801), .QN(n2427) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n2529), .CLK(n2660), .Q(
        g186) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n2517), .CLK(n2666), .Q(
        g959) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n2508), .CLK(n2671), .Q(
        test_so2) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n2570), .CLK(n2639), 
        .Q(g1407) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n2570), .CLK(n2640), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n2570), .CLK(n2640), .Q(
        g4173), .QN(n2451) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n2553), .CLK(n2648), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n2558), .CLK(n2646), .Q(
        g396) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n2574), .CLK(n2637), .Q(
        g1015), .QN(n2322) );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(n2574), .CLK(n2638), .Q(
        n1650) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n2574), .CLK(n2638), .Q(
        n3059), .QN(n1874) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n2524), .CLK(n2662), .Q(
        g1415) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n2589), .CLK(n2630), .Q(
        g1227), .QN(n2448) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n2589), .CLK(n2630), .Q(
        g1721) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n2506), .CLK(n2671), .Q(
        n3058) );
  SDFFX1 DFF_122_Q_reg ( .D(n2499), .SI(n3058), .SE(n2506), .CLK(n2671), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(n2506), .CLK(n2672), .Q(
        g284) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n2578), .CLK(n2636), .Q(
        g426) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n2577), .CLK(n2636), .Q(
        g219), .QN(n2460) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n2523), .CLK(n2663), .Q(
        n3056) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n2523), .CLK(n2663), .Q(
        g806), .QN(n2432) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n2570), .CLK(n2639), .Q(
        g1428), .QN(n2404) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n2570), .CLK(n2639), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n2578), .CLK(n2635), .Q(
        g1564) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n2553), .CLK(n2648), .Q(
        g1741) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n2586), .CLK(n2631), .Q(
        g225), .QN(n2457) );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(n2537), .CLK(n2656), .Q(
        g281) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n2537), .CLK(n2656), .Q(
        g1308) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n2567), .CLK(n2641), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n2533), .CLK(n2658), .Q(
        n3055) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n2533), .CLK(n2658), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n2505), .CLK(n2672), .Q(
        g1589) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n2573), .CLK(n2638), .Q(
        g1466) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n2513), .CLK(n2668), .Q(
        g1571) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n2525), .CLK(n2662), .Q(
        g1861), .QN(n2417) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n2525), .CLK(n2662), .Q(
        n3054) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n2578), .CLK(n2635), .Q(
        g1448), .QN(n2473) );
  SDFFX1 DFF_145_Q_reg ( .D(n192), .SI(g1448), .SE(n2578), .CLK(n2636), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n2575), .CLK(n2637), .Q(
        g1333) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n2575), .CLK(n2637), .Q(
        g153), .QN(n2362) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n2514), .CLK(n2668), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(n2569), .CLK(n2640), .Q(
        g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n2569), .CLK(n2640), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n2569), .CLK(n2640), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n2545), .CLK(n2652), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n2545), .CLK(n2652), .Q(
        g1397) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n2545), .CLK(n2652), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n2555), .CLK(n2647), .Q(
        g1950) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n2552), .CLK(n2649), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(n167), .SI(g756), .SE(n2574), .CLK(n2638), .Q(
        n3053) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n2543), .CLK(n2653), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n2587), .CLK(n2631), .Q(
        g105), .QN(n2482) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n2587), .CLK(n2631), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n2587), .CLK(n2631), .Q(
        test_so3) );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(n2579), .CLK(n2635), 
        .Q(g1531) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n2578), .CLK(n2635), .Q(
        g1458) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n2553), .CLK(n2648), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n2562), .CLK(n2644), .Q(
        g1011), .QN(n2354) );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(n2562), .CLK(n2644), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n2562), .CLK(n2644), .Q(
        g1411) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n2574), .CLK(n2637), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n2556), .CLK(n2646), .Q(
        g444) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n2586), .CLK(n2632), .Q(
        g1474), .QN(n2412) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n2564), .CLK(n2643), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n2563), .CLK(n2643), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n2515), .CLK(n2667), .Q(
        g333), .QN(n2369) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n2515), .CLK(n2667), .Q(
        g269) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n2557), .CLK(n2646), .Q(
        g401) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n2589), .CLK(n2630), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n2588), .CLK(n2631), .Q(g9) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n2576), .CLK(n2637), .Q(g664), 
        .QN(n2429) );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n2516), .CLK(n2666), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n2516), .CLK(n2667), .Q(
        g1400) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n2518), .CLK(n2665), .Q(
        g309), .QN(n2201) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n2518), .CLK(n2665), .Q(
        g814), .QN(n2431) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n2525), .CLK(n2662), .Q(
        g231), .QN(n2459) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n2546), .CLK(n2651), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n2546), .CLK(n2651), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n2528), .CLK(n2661), .Q(
        g869) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n2528), .CLK(n2661), .Q(
        g1383) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n2508), .CLK(n2671), .Q(
        g158), .QN(n2348) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n2583), .CLK(n2633), .Q(
        g627) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n2559), .CLK(n2645), .Q(
        g1023) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n2559), .CLK(n2645), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n2559), .CLK(n2645), .Q(
        n3050), .QN(n4318) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n2526), .CLK(n2662), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(n119), .SI(g1327), .SE(n2583), .CLK(n2633), .Q(
        g654), .QN(n2450) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n2542), .CLK(n2653), .Q(
        g293) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n2542), .CLK(n2654), .Q(
        g1346) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n2513), .CLK(n2668), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n2513), .CLK(n2668), .Q(
        g1753) );
  SDFFX1 DFF_201_Q_reg ( .D(n2496), .SI(g1753), .SE(n2512), .CLK(n2668), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n2534), .CLK(n2657), .Q(
        g1240), .QN(n2375) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n2534), .CLK(n2657), .Q(
        g538), .QN(n2409) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n2557), .CLK(n2646), .Q(
        g416) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n2536), .CLK(n2656), .Q(
        g542), .QN(n2410) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n2536), .CLK(n2656), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n2548), .CLK(n2651), .Q(
        g374), .QN(n2434) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n2548), .CLK(n2651), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n2555), .CLK(n2647), .Q(
        g1914), .QN(n2326) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n2522), .CLK(n2664), .Q(
        g530), .QN(n2407) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n2521), .CLK(n2664), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n2580), .CLK(n2635), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n2579), .CLK(n2635), .Q(
        g8978) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n2579), .CLK(n2635), .Q(
        test_so4) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n2558), .CLK(n2645), 
        .Q(g1317), .QN(n2478) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n2558), .CLK(n2645), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n2558), .CLK(n2646), .Q(
        g386) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n2510), .CLK(n2669), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n2510), .CLK(n2669), .Q(
        g166) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n2541), .CLK(n2654), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n2516), .CLK(n2667), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n2554), .CLK(n2647), .Q(
        g1840), .QN(n2442) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n2550), .CLK(n2650), .Q(
        g8983) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n2546), .CLK(n2652), .Q(
        g318), .QN(n2358) );
  SDFFX1 DFF_226_Q_reg ( .D(n227), .SI(g318), .SE(n2558), .CLK(n2645), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n2551), .CLK(n2649), .Q(
        g794), .QN(n2443) );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(n2551), .CLK(n2649), .Q(
        n3048) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n2575), .CLK(n2637), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n2574), .CLK(n2637), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n2533), .CLK(n2658), .Q(
        g1250), .QN(n2355) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n2533), .CLK(n2658), .Q(
        g1163), .QN(n2424) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n2506), .CLK(n2672), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n2569), .CLK(n2640), .Q(
        g1032), .QN(n2477) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n2568), .CLK(n2640), .Q(
        g1432), .QN(n2474) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n2579), .CLK(n2635), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n2545), .CLK(n2652), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n2544), .CLK(n2652), .Q(g330), .QN(n2200) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n2544), .CLK(n2652), .Q(
        g1157), .QN(n2422) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n2544), .CLK(n2652), .Q(
        n3046), .QN(n4323) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(n2544), .CLK(n2653), .Q(
        n3045) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n2544), .CLK(n2653), .Q(
        g928) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n2537), .CLK(n2656), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n2537), .CLK(n2656), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n2521), .CLK(n2664), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n2521), .CLK(n2664), .Q(
        g4178), .QN(n2446) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n2515), .CLK(n2667), .Q(
        g861) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n2515), .CLK(n2667), .Q(
        g1627) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n2565), .CLK(n2642), .Q(
        g1292), .QN(n2334) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n2532), .CLK(n2659), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n2532), .CLK(n2659), .Q(
        n3044), .QN(n1873) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n2531), .CLK(n2659), .Q(
        g4176), .QN(n2447) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n2560), .CLK(n2644), .Q(
        g1583) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n2560), .CLK(n2644), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n2560), .CLK(n2644), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n2584), .CLK(n2633), .Q(
        g1546) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n2536), .CLK(n2657), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n2536), .CLK(n2657), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n2536), .CLK(n2657), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n2497), .SI(g617), .SE(n2535), .CLK(n2657), .Q(
        n1631) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n2571), .CLK(n2639), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n2545), .CLK(n2652), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n2528), .CLK(n2660), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n2569), .CLK(n2640), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n2581), .CLK(n2634), .Q(g8)
         );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n2553), .CLK(n2648), .Q(
        test_so5), .QN(n2504) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n2519), .CLK(n2665), .Q(
        g2648) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n2518), .CLK(n2665), .Q(
        g255) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n2585), .CLK(n2632), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n2584), .CLK(n2632), .Q(
        g1738) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n2584), .CLK(n2632), .Q(
        g1478), .QN(n2401) );
  SDFFX1 DFF_275_Q_reg ( .D(n507), .SI(g1478), .SE(n2584), .CLK(n2632), .Q(
        n3042) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n2529), .CLK(n2660), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n2519), .CLK(n2665), .Q(
        g1482) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n2519), .CLK(n2665), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n2509), .CLK(n2670), .Q(
        g296) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n2508), .CLK(n2670), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n2508), .CLK(n2670), .Q(
        g700), .QN(n2366) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n2563), .CLK(n2643), .Q(
        g1762) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n2562), .CLK(n2643), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n2562), .CLK(n2643), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n2584), .CLK(n2633), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n2584), .CLK(n2633), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n2549), .CLK(n2650), .Q(
        g8980) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n2514), .CLK(n2667), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n2587), .CLK(n2631), .Q(
        n3041) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n2587), .CLK(n2631), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n2559), .CLK(n2645), .Q(
        g2986), .QN(n2476) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n2559), .CLK(n2645), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n2581), .CLK(n2634), .Q(
        g986) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n2577), .CLK(n2636), .Q(
        g971) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n2577), .CLK(n2636), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n2575), .CLK(n2637), .Q(
        g143), .QN(n2363) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n2580), .CLK(n2635), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n2533), .CLK(n2658), .Q(
        g1212), .QN(n2465) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n2506), .CLK(n2671), .Q(
        g1918), .QN(n2420) );
  SDFFX1 DFF_301_Q_reg ( .D(n106), .SI(g1918), .SE(n2580), .CLK(n2634), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n2580), .CLK(n2635), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n2538), .CLK(n2656), .Q(
        g237) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n2551), .CLK(n2649), .Q(g746), .QN(n2463) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n2520), .CLK(n2664), .Q(
        g1462), .QN(n2400) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n2520), .CLK(n2664), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n2540), .CLK(n2654), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n2540), .CLK(n2654), .Q(g837) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n2540), .CLK(n2655), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n2589), .CLK(n2630), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n2589), .CLK(n2630), .Q(
        g944) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n2555), .CLK(n2647), .Q(
        g1941) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n2525), .CLK(n2662), .Q(
        g170) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n2525), .CLK(n2662), .Q(
        g1520) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n2513), .CLK(n2668), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n2513), .CLK(n2668), .Q(
        g953) );
  SDFFX1 DFF_318_Q_reg ( .D(n112), .SI(g953), .SE(n2563), .CLK(n2643), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(n2563), .CLK(n2643), .Q(
        n3040) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n2563), .CLK(n2643), .Q(
        g1765), .QN(n2469) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n2552), .CLK(n2648), .Q(
        g1733) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n2552), .CLK(n2648), .Q(
        test_so6), .QN(n2502) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n2553), .CLK(n2648), 
        .Q(g1610), .QN(n2468) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n2526), .CLK(n2661), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n2526), .CLK(n2661), .Q(
        g1324) );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(n2526), .CLK(n2661), .Q(
        g1540) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n2526), .CLK(n2662), .Q(
        n3038), .QN(n4315) );
  SDFFX1 DFF_328_Q_reg ( .D(n2498), .SI(n3038), .SE(n2541), .CLK(n2654), .Q(
        g3069) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n2541), .CLK(n2654), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n2530), .CLK(n2659), .Q(
        n3037) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n2530), .CLK(n2659), .Q(
        g213) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n2530), .CLK(n2659), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n2510), .CLK(n2670), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n2534), .CLK(n2658), .Q(
        g1245), .QN(n2352) );
  SDFFX1 DFF_335_Q_reg ( .D(n7), .SI(g1245), .SE(n2534), .CLK(n2658), .Q(n3036) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(n2534), .CLK(n2658), .Q(
        n3035) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n2527), .CLK(n2661), .Q(
        g148), .QN(n2364) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n2527), .CLK(n2661), .Q(g833) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n2555), .CLK(n2647), .Q(
        g1923) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n2555), .CLK(n2647), .Q(
        g936) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n2522), .CLK(n2664), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n2518), .CLK(n2666), .Q(
        g849) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n2518), .CLK(n2666), .Q(
        g1336), .QN(n2383) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n2517), .CLK(n2666), .Q(
        g272) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n2517), .CLK(n2666), .Q(
        g1806), .QN(n2426) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n2515), .CLK(n2667), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n2512), .CLK(n2668), .Q(
        g1887) );
  SDFFX1 DFF_350_Q_reg ( .D(g10724), .SI(g1887), .SE(n2512), .CLK(n2668), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n2512), .CLK(n2669), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n2531), .CLK(n2659), .Q(
        n3033), .QN(n4313) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(n2531), .CLK(n2659), .Q(
        g1137) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n2585), .CLK(n2632), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n2533), .CLK(n2658), .Q(
        g1255), .QN(n2330) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n2546), .CLK(n2652), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n2546), .CLK(n2652), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n2583), .CLK(n2633), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n2581), .CLK(n2634), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n2581), .CLK(n2634), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n2589), .CLK(n2630), .Q(
        g1218), .QN(n2472) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n2540), .CLK(n2655), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n2540), .CLK(n2655), .Q(
        g8986) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n2520), .CLK(n2664), .Q(
        g182), .QN(n2471) );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(n2520), .CLK(n2665), .Q(
        g950) );
  SDFFX1 DFF_366_Q_reg ( .D(n363), .SI(g950), .SE(n2520), .CLK(n2665), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n2516), .CLK(n2666), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n2556), .CLK(n2646), .Q(
        g448) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n2554), .CLK(n2647), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n2554), .CLK(n2648), .Q(
        g1727) );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(n2554), .CLK(n2648), .Q(
        g1592) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n2554), .CLK(n2648), .Q(
        g1703), .QN(n2406) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n2555), .CLK(n2647), .Q(
        g1932), .QN(n2329) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n2520), .CLK(n2665), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n2571), .CLK(n2639), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n2590), .CLK(n2630), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n2556), .CLK(n2646), .Q(
        g440) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n2537), .CLK(n2656), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n2537), .CLK(n2656), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n2576), .CLK(n2637), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n2543), .CLK(n2653), .Q(
        g139), .QN(n2344) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n2543), .CLK(n2653), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(n2542), .CLK(n2653), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n2531), .CLK(n2659), .Q(
        n3030) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n2519), .CLK(n2665), .Q(
        g263) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n2517), .CLK(n2666), .Q(
        g818), .QN(n2395) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n2514), .CLK(n2667), .Q(
        g1747) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n2549), .CLK(n2650), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n2507), .CLK(n2671), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n2507), .CLK(n2671), .Q(
        g1524) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n2507), .CLK(n2671), .Q(
        g1577) );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(n2549), .CLK(n2650), .Q(
        g810), .QN(n2396) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n2558), .CLK(n2646), .Q(
        g391) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n2583), .CLK(n2633), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n2528), .CLK(n2660), .Q(
        g1386) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n2528), .CLK(n2660), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n2528), .CLK(n2661), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(n395), .SI(g875), .SE(n2527), .CLK(n2661), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n2588), .CLK(n2631), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n2505), .CLK(n2672), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n2566), .CLK(n2641), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n2539), .CLK(n2655), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n2573), .CLK(n2638), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n2514), .CLK(n2667), .Q(
        g853) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n2557), .CLK(n2646), .Q(
        g421) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n2570), .CLK(n2640), .Q(
        g4174), .QN(n2452) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n2548), .CLK(n2650), .Q(
        g956) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n2548), .CLK(n2650), .Q(
        g378), .QN(n2433) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n2526), .CLK(n2662), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n2525), .CLK(n2662), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n2523), .CLK(n2663), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n2571), .CLK(n2639), .Q(
        g1027), .QN(n2392) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n2571), .CLK(n2639), .Q(
        g1003), .QN(n2376) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n2571), .CLK(n2639), .Q(
        g1403) );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(n2571), .CLK(n2639), .Q(
        g1145) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n2522), .CLK(n2663), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n2522), .CLK(n2663), .Q(
        g1223), .QN(n2449) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n2557), .CLK(n2646), .Q(
        g406) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n2505), .CLK(n2672), .Q(
        g1811), .QN(n1699) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(n2505), .CLK(n2672), .Q(
        n3029), .QN(n4320) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n2588), .CLK(n2630), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(n2588), .CLK(n2630), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n2568), .CLK(n2640), .Q(
        g1595) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n2568), .CLK(n2640), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n2576), .CLK(n2636), .Q(
        g727) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n2587), .CLK(n2631), .Q(
        test_so8) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n2551), .CLK(n2649), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n2551), .CLK(n2649), .Q(
        g481), .QN(n1680) );
  SDFFX1 DFF_431_Q_reg ( .D(n319), .SI(g481), .SE(n2550), .CLK(n2649), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n2527), .CLK(n2661), .Q(
        g1330) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n2549), .CLK(n2650), .Q(
        g845) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n2521), .CLK(n2664), .Q(
        g4181), .QN(n2441) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n2521), .CLK(n2664), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n2560), .CLK(n2645), .Q(
        n3027), .QN(DFF_436_n1) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n2564), .CLK(n2642), .Q(
        g1490), .QN(n2399) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n2564), .CLK(n2643), .Q(
        g1166), .QN(n2425) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n2564), .CLK(n2643), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n2545), .CLK(n2652), .Q(
        n3026) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n2532), .CLK(n2658), .Q(
        g1260), .QN(n2331) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n2532), .CLK(n2658), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n2532), .CLK(n2658), .Q(
        g131), .QN(n2343) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n2532), .CLK(n2659), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n2535), .CLK(n2657), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n2509), .CLK(n2670), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n2509), .CLK(n2670), .Q(
        g1318) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n2585), .CLK(n2632), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n2582), .CLK(n2633), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n2582), .CLK(n2633), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n2493), .SI(g2608), .SE(n2582), .CLK(n2633), .Q(
        n3024) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n2582), .CLK(n2634), .Q(
        g1549) );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(n2527), .CLK(n2661), .Q(
        g947) );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(n2554), .CLK(n2647), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n2547), .CLK(n2651), .Q(
        g1598) );
  SDFFX1 DFF_457_Q_reg ( .D(n435), .SI(g1598), .SE(n2547), .CLK(n2651), .Q(
        g1121) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n2530), .CLK(n2660), .Q(
        g1321) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n2541), .CLK(n2654), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n2541), .CLK(n2654), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n2552), .CLK(n2649), .Q(
        g1909), .QN(n2421) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n2552), .CLK(n2649), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n2572), .CLK(n2638), .Q(
        g1552) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n2572), .CLK(n2638), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n2572), .CLK(n2638), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(n2572), .CLK(n2639), .Q(
        g1586) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n2572), .CLK(n2639), .Q(
        g324), .QN(n2356) );
  SDFFX1 DFF_468_Q_reg ( .D(n443), .SI(g324), .SE(n2572), .CLK(n2639), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n2518), .CLK(n2666), .Q(
        g1341) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n2517), .CLK(n2666), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(n2517), .CLK(n2666), .Q(
        n3023), .QN(n4319) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(n2588), .CLK(n2631), .Q(
        n3022), .QN(n4312) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n2542), .CLK(n2653), .Q(
        g135), .QN(n2345) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n2514), .CLK(n2668), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n2514), .CLK(n2668), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n2513), .CLK(n2668), .Q(
        g1607) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n2535), .CLK(n2657), .Q(
        g321), .QN(n2380) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n2535), .CLK(n2657), .Q(
        g8982) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n2535), .CLK(n2657), .Q(
        g1275), .QN(n2373) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n2535), .CLK(n2657), .Q(
        test_so9) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n2546), .CLK(n2651), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n2548), .CLK(n2650), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(n2507), .CLK(n2671), .Q(
        n3020) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n2507), .CLK(n2671), .Q(
        g266) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n2565), .CLK(n2642), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n2565), .CLK(n2642), .Q(
        n3019), .QN(n4314) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n2576), .CLK(n2637), .Q(
        g673) );
  SDFFX1 DFF_489_Q_reg ( .D(n274), .SI(g673), .SE(n2531), .CLK(n2659), .Q(
        n3018) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n2547), .CLK(n2651), .Q(
        g162), .QN(n2347) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n2557), .CLK(n2646), .Q(
        g411) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n2556), .CLK(n2647), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n2556), .CLK(n2647), .Q(
        g1905), .QN(n2436) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n2538), .CLK(n2656), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n2586), .CLK(n2631), .Q(
        g1630) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n2549), .CLK(n2650), .Q(
        g8976) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n2566), .CLK(n2642), .Q(
        g991) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n2566), .CLK(n2642), .Q(
        g1300), .QN(n2336) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n2511), .CLK(n2669), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n2511), .CLK(n2669), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n2511), .CLK(n2669), .Q(
        g1750) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n2511), .CLK(n2669), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n2511), .CLK(n2669), .Q(
        g1440), .QN(n2403) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n2511), .CLK(n2669), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(n2510), .CLK(n2669), .Q(
        g1528) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n2542), .CLK(n2654), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(n2542), .CLK(n2654), .Q(
        n3017), .QN(n4322) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n2536), .CLK(n2656), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n2579), .CLK(n2635), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n2534), .CLK(n2657), .Q(
        g1235), .QN(n2353) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n2510), .CLK(n2670), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n2556), .CLK(n2647), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n2550), .CLK(n2650), .Q(
        g8981) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(n2550), .CLK(n2650), .Q(
        g1555) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n2505), .CLK(n2672), .Q(
        g995), .QN(n2374) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n2565), .CLK(n2642), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n2564), .CLK(n2642), .Q(
        n3016), .QN(n4316) );
  SDFFX1 DFF_518_Q_reg ( .D(n118), .SI(n3016), .SE(n2583), .CLK(n2633), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n2568), .CLK(n2641), .Q(
        g1494), .QN(n2411) );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(n2524), .CLK(n2662), .Q(
        g1567) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n2524), .CLK(n2662), .Q(
        g691), .QN(n2435) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n2524), .CLK(n2663), .Q(
        g534), .QN(n2408) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n2524), .CLK(n2663), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n2524), .CLK(n2663), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n2523), .CLK(n2663), .Q(
        g1160), .QN(n2423) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n2523), .CLK(n2663), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n2578), .CLK(n2636), .Q(g1) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n2540), .CLK(n2654), .Q(g511), .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n2586), .CLK(n2632), .Q(
        g1724) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n2585), .CLK(n2632), .Q(
        g12) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n2585), .CLK(n2632), .Q(
        g1878) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n2549), .CLK(n2650), .Q(
        test_so10) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n2573), .CLK(n2638), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(g6179), .IN2(n2493), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n42), .IN2(n1132), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n1226), .IN2(n1858), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(n112), .IN2(n898), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n12), .IN2(n57), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n40), .IN2(n40), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n124), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n938), .IN2(n2492), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n2492), .IN2(n2492), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n2492), .IN2(n2492), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n2492), .IN2(n2492), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n113), .IN2(n84), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n86), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n257), .IN2(n155), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n2590), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n371), .S(Trigger_select), .Q(
        g4207) );
  NBUFFX2 U2511 ( .INP(n2681), .Z(n2631) );
  NBUFFX2 U2512 ( .INP(n2681), .Z(n2632) );
  NBUFFX2 U2513 ( .INP(n2681), .Z(n2630) );
  NBUFFX2 U2514 ( .INP(n2677), .Z(n2650) );
  NBUFFX2 U2515 ( .INP(n2676), .Z(n2657) );
  NBUFFX2 U2516 ( .INP(n2678), .Z(n2647) );
  NBUFFX2 U2517 ( .INP(n2677), .Z(n2652) );
  NBUFFX2 U2518 ( .INP(n2673), .Z(n2668) );
  NBUFFX2 U2519 ( .INP(n2675), .Z(n2658) );
  NBUFFX2 U2520 ( .INP(n2675), .Z(n2662) );
  NBUFFX2 U2521 ( .INP(n2679), .Z(n2639) );
  NBUFFX2 U2522 ( .INP(n2674), .Z(n2666) );
  NBUFFX2 U2523 ( .INP(n2677), .Z(n2648) );
  NBUFFX2 U2524 ( .INP(n2675), .Z(n2661) );
  NBUFFX2 U2525 ( .INP(n2676), .Z(n2655) );
  NBUFFX2 U2526 ( .INP(n2680), .Z(n2633) );
  NBUFFX2 U2527 ( .INP(n2675), .Z(n2660) );
  NBUFFX2 U2528 ( .INP(n2680), .Z(n2637) );
  NBUFFX2 U2529 ( .INP(n2676), .Z(n2654) );
  NBUFFX2 U2530 ( .INP(n2677), .Z(n2649) );
  NBUFFX2 U2531 ( .INP(n2679), .Z(n2638) );
  NBUFFX2 U2532 ( .INP(n2680), .Z(n2635) );
  NBUFFX2 U2535 ( .INP(n2674), .Z(n2667) );
  NBUFFX2 U2536 ( .INP(n2674), .Z(n2663) );
  NBUFFX2 U2537 ( .INP(n2675), .Z(n2659) );
  NBUFFX2 U2538 ( .INP(n2679), .Z(n2640) );
  NBUFFX2 U2539 ( .INP(n2676), .Z(n2653) );
  NBUFFX2 U2540 ( .INP(n2678), .Z(n2644) );
  NBUFFX2 U2541 ( .INP(n2677), .Z(n2651) );
  NBUFFX2 U2542 ( .INP(n2673), .Z(n2670) );
  NBUFFX2 U2543 ( .INP(n2676), .Z(n2656) );
  NBUFFX2 U2544 ( .INP(n2678), .Z(n2643) );
  NBUFFX2 U2545 ( .INP(n2680), .Z(n2636) );
  NBUFFX2 U2546 ( .INP(n2678), .Z(n2645) );
  NBUFFX2 U2547 ( .INP(n2679), .Z(n2641) );
  NBUFFX2 U2548 ( .INP(n2674), .Z(n2665) );
  NBUFFX2 U2549 ( .INP(n2674), .Z(n2664) );
  NBUFFX2 U2550 ( .INP(n2680), .Z(n2634) );
  NBUFFX2 U2551 ( .INP(n2679), .Z(n2642) );
  NBUFFX2 U2552 ( .INP(n2673), .Z(n2671) );
  NBUFFX2 U2553 ( .INP(n2678), .Z(n2646) );
  NBUFFX2 U2554 ( .INP(n2673), .Z(n2669) );
  NBUFFX2 U2555 ( .INP(n2673), .Z(n2672) );
  NBUFFX2 U2556 ( .INP(n2619), .Z(n2505) );
  NBUFFX2 U2557 ( .INP(n2619), .Z(n2506) );
  NBUFFX2 U2558 ( .INP(n2618), .Z(n2507) );
  NBUFFX2 U2559 ( .INP(n2618), .Z(n2508) );
  NBUFFX2 U2560 ( .INP(n2618), .Z(n2509) );
  NBUFFX2 U2561 ( .INP(n2617), .Z(n2510) );
  NBUFFX2 U2562 ( .INP(n2617), .Z(n2511) );
  NBUFFX2 U2563 ( .INP(n2617), .Z(n2512) );
  NBUFFX2 U2564 ( .INP(n2616), .Z(n2513) );
  NBUFFX2 U2565 ( .INP(n2616), .Z(n2514) );
  NBUFFX2 U2566 ( .INP(n2616), .Z(n2515) );
  NBUFFX2 U2567 ( .INP(n2615), .Z(n2516) );
  NBUFFX2 U2568 ( .INP(n2615), .Z(n2517) );
  NBUFFX2 U2569 ( .INP(n2615), .Z(n2518) );
  NBUFFX2 U2570 ( .INP(n2614), .Z(n2519) );
  NBUFFX2 U2571 ( .INP(n2614), .Z(n2520) );
  NBUFFX2 U2572 ( .INP(n2614), .Z(n2521) );
  NBUFFX2 U2573 ( .INP(n2613), .Z(n2522) );
  NBUFFX2 U2574 ( .INP(n2613), .Z(n2523) );
  NBUFFX2 U2575 ( .INP(n2613), .Z(n2524) );
  NBUFFX2 U2576 ( .INP(n2612), .Z(n2525) );
  NBUFFX2 U2577 ( .INP(n2612), .Z(n2526) );
  NBUFFX2 U2578 ( .INP(n2612), .Z(n2527) );
  NBUFFX2 U2579 ( .INP(n2611), .Z(n2528) );
  NBUFFX2 U2580 ( .INP(n2611), .Z(n2529) );
  NBUFFX2 U2581 ( .INP(n2611), .Z(n2530) );
  NBUFFX2 U2582 ( .INP(n2610), .Z(n2531) );
  NBUFFX2 U2583 ( .INP(n2610), .Z(n2532) );
  NBUFFX2 U2584 ( .INP(n2610), .Z(n2533) );
  NBUFFX2 U2585 ( .INP(n2609), .Z(n2534) );
  NBUFFX2 U2586 ( .INP(n2609), .Z(n2535) );
  NBUFFX2 U2587 ( .INP(n2609), .Z(n2536) );
  NBUFFX2 U2588 ( .INP(n2608), .Z(n2537) );
  NBUFFX2 U2589 ( .INP(n2608), .Z(n2538) );
  NBUFFX2 U2590 ( .INP(n2608), .Z(n2539) );
  NBUFFX2 U2591 ( .INP(n2607), .Z(n2540) );
  NBUFFX2 U2592 ( .INP(n2607), .Z(n2541) );
  NBUFFX2 U2593 ( .INP(n2607), .Z(n2542) );
  NBUFFX2 U2594 ( .INP(n2606), .Z(n2543) );
  NBUFFX2 U2595 ( .INP(n2606), .Z(n2544) );
  NBUFFX2 U2596 ( .INP(n2606), .Z(n2545) );
  NBUFFX2 U2597 ( .INP(n2605), .Z(n2546) );
  NBUFFX2 U2598 ( .INP(n2605), .Z(n2547) );
  NBUFFX2 U2599 ( .INP(n2605), .Z(n2548) );
  NBUFFX2 U2600 ( .INP(n2604), .Z(n2549) );
  NBUFFX2 U2601 ( .INP(n2604), .Z(n2550) );
  NBUFFX2 U2602 ( .INP(n2604), .Z(n2551) );
  NBUFFX2 U2603 ( .INP(n2603), .Z(n2552) );
  NBUFFX2 U2604 ( .INP(n2603), .Z(n2553) );
  NBUFFX2 U2605 ( .INP(n2603), .Z(n2554) );
  NBUFFX2 U2606 ( .INP(n2602), .Z(n2555) );
  NBUFFX2 U2607 ( .INP(n2602), .Z(n2556) );
  NBUFFX2 U2608 ( .INP(n2602), .Z(n2557) );
  NBUFFX2 U2609 ( .INP(n2601), .Z(n2558) );
  NBUFFX2 U2610 ( .INP(n2601), .Z(n2559) );
  NBUFFX2 U2611 ( .INP(n2601), .Z(n2560) );
  NBUFFX2 U2612 ( .INP(n2600), .Z(n2561) );
  NBUFFX2 U2613 ( .INP(n2600), .Z(n2562) );
  NBUFFX2 U2614 ( .INP(n2600), .Z(n2563) );
  NBUFFX2 U2615 ( .INP(n2599), .Z(n2564) );
  NBUFFX2 U2616 ( .INP(n2599), .Z(n2565) );
  NBUFFX2 U2617 ( .INP(n2599), .Z(n2566) );
  NBUFFX2 U2618 ( .INP(n2598), .Z(n2567) );
  NBUFFX2 U2619 ( .INP(n2598), .Z(n2568) );
  NBUFFX2 U2620 ( .INP(n2598), .Z(n2569) );
  NBUFFX2 U2621 ( .INP(n2597), .Z(n2570) );
  NBUFFX2 U2622 ( .INP(n2597), .Z(n2571) );
  NBUFFX2 U2623 ( .INP(n2597), .Z(n2572) );
  NBUFFX2 U2624 ( .INP(n2596), .Z(n2573) );
  NBUFFX2 U2625 ( .INP(n2596), .Z(n2574) );
  NBUFFX2 U2626 ( .INP(n2596), .Z(n2575) );
  NBUFFX2 U2627 ( .INP(n2595), .Z(n2576) );
  NBUFFX2 U2628 ( .INP(n2595), .Z(n2577) );
  NBUFFX2 U2629 ( .INP(n2595), .Z(n2578) );
  NBUFFX2 U2630 ( .INP(n2594), .Z(n2579) );
  NBUFFX2 U2631 ( .INP(n2594), .Z(n2580) );
  NBUFFX2 U2632 ( .INP(n2594), .Z(n2581) );
  NBUFFX2 U2633 ( .INP(n2593), .Z(n2582) );
  NBUFFX2 U2634 ( .INP(n2593), .Z(n2583) );
  NBUFFX2 U2635 ( .INP(n2593), .Z(n2584) );
  NBUFFX2 U2636 ( .INP(n2592), .Z(n2585) );
  NBUFFX2 U2637 ( .INP(n2592), .Z(n2586) );
  NBUFFX2 U2638 ( .INP(n2592), .Z(n2587) );
  NBUFFX2 U2640 ( .INP(n2591), .Z(n2588) );
  NBUFFX2 U2642 ( .INP(n2591), .Z(n2589) );
  NBUFFX2 U2643 ( .INP(n2591), .Z(n2590) );
  NBUFFX2 U2644 ( .INP(n2629), .Z(n2591) );
  NBUFFX2 U2645 ( .INP(n2629), .Z(n2592) );
  NBUFFX2 U2646 ( .INP(n2628), .Z(n2593) );
  NBUFFX2 U2647 ( .INP(n2628), .Z(n2594) );
  NBUFFX2 U2648 ( .INP(n2628), .Z(n2595) );
  NBUFFX2 U2649 ( .INP(n2627), .Z(n2596) );
  NBUFFX2 U2650 ( .INP(n2627), .Z(n2597) );
  NBUFFX2 U2651 ( .INP(n2627), .Z(n2598) );
  NBUFFX2 U2652 ( .INP(n2626), .Z(n2599) );
  NBUFFX2 U2653 ( .INP(n2626), .Z(n2600) );
  NBUFFX2 U2655 ( .INP(n2626), .Z(n2601) );
  NBUFFX2 U2656 ( .INP(n2625), .Z(n2602) );
  NBUFFX2 U2657 ( .INP(n2625), .Z(n2603) );
  NBUFFX2 U2659 ( .INP(n2625), .Z(n2604) );
  NBUFFX2 U2660 ( .INP(n2624), .Z(n2605) );
  NBUFFX2 U2661 ( .INP(n2624), .Z(n2606) );
  NBUFFX2 U2662 ( .INP(n2624), .Z(n2607) );
  NBUFFX2 U2663 ( .INP(n2623), .Z(n2608) );
  NBUFFX2 U2664 ( .INP(n2623), .Z(n2609) );
  NBUFFX2 U2665 ( .INP(n2623), .Z(n2610) );
  NBUFFX2 U2666 ( .INP(n2622), .Z(n2611) );
  NBUFFX2 U2667 ( .INP(n2622), .Z(n2612) );
  NBUFFX2 U2668 ( .INP(n2622), .Z(n2613) );
  NBUFFX2 U2669 ( .INP(n2621), .Z(n2614) );
  NBUFFX2 U2670 ( .INP(n2621), .Z(n2615) );
  NBUFFX2 U2671 ( .INP(n2621), .Z(n2616) );
  NBUFFX2 U2672 ( .INP(n2620), .Z(n2617) );
  NBUFFX2 U2673 ( .INP(n2620), .Z(n2618) );
  NBUFFX2 U2674 ( .INP(n2620), .Z(n2619) );
  NBUFFX2 U2675 ( .INP(test_se), .Z(n2620) );
  NBUFFX2 U2676 ( .INP(n2625), .Z(n2621) );
  NBUFFX2 U2677 ( .INP(n2602), .Z(n2622) );
  NBUFFX2 U2678 ( .INP(n2603), .Z(n2623) );
  NBUFFX2 U2679 ( .INP(n2604), .Z(n2624) );
  NBUFFX2 U2680 ( .INP(test_se), .Z(n2625) );
  NBUFFX2 U2681 ( .INP(test_se), .Z(n2626) );
  NBUFFX2 U2682 ( .INP(n2619), .Z(n2627) );
  NBUFFX2 U2684 ( .INP(test_se), .Z(n2628) );
  NBUFFX2 U2685 ( .INP(n2620), .Z(n2629) );
  NBUFFX2 U2686 ( .INP(n2684), .Z(n2673) );
  NBUFFX2 U2687 ( .INP(n2684), .Z(n2674) );
  NBUFFX2 U2688 ( .INP(n2684), .Z(n2675) );
  NBUFFX2 U2689 ( .INP(n2683), .Z(n2676) );
  NBUFFX2 U2690 ( .INP(n2683), .Z(n2677) );
  NBUFFX2 U2691 ( .INP(n2683), .Z(n2678) );
  NBUFFX2 U2692 ( .INP(n2682), .Z(n2679) );
  NBUFFX2 U2693 ( .INP(n2682), .Z(n2680) );
  NBUFFX2 U2694 ( .INP(n2682), .Z(n2681) );
  NBUFFX2 U2695 ( .INP(CK), .Z(n2682) );
  NBUFFX2 U2696 ( .INP(CK), .Z(n2683) );
  NBUFFX2 U2697 ( .INP(CK), .Z(n2684) );
  OR2X1 U2700 ( .IN1(n2685), .IN2(n2686), .Q(n962) );
  AND2X1 U2701 ( .IN1(n2687), .IN2(n1696), .Q(n2686) );
  INVX0 U2702 ( .INP(n2688), .ZN(n2685) );
  OR2X1 U2703 ( .IN1(n57), .IN2(n1696), .Q(n2688) );
  OR2X1 U2704 ( .IN1(n2689), .IN2(n2690), .Q(n917) );
  AND2X1 U2705 ( .IN1(n2691), .IN2(n1697), .Q(n2690) );
  INVX0 U2706 ( .INP(n2692), .ZN(n2689) );
  OR2X1 U2707 ( .IN1(n12), .IN2(n1697), .Q(n2692) );
  INVX0 U2708 ( .INP(n2693), .ZN(n68) );
  OR2X1 U2709 ( .IN1(n2694), .IN2(n2695), .Q(n2693) );
  AND2X1 U2710 ( .IN1(n2696), .IN2(n2697), .Q(n2695) );
  OR2X1 U2711 ( .IN1(n2698), .IN2(n2416), .Q(n2696) );
  AND2X1 U2712 ( .IN1(n3033), .IN2(n2417), .Q(n2698) );
  INVX0 U2713 ( .INP(n2699), .ZN(n57) );
  INVX0 U2714 ( .INP(n2700), .ZN(n517) );
  INVX0 U2715 ( .INP(n2701), .ZN(n510) );
  INVX0 U2716 ( .INP(n2702), .ZN(n491) );
  INVX0 U2717 ( .INP(n2703), .ZN(n45) );
  AND2X1 U2718 ( .IN1(g109), .IN2(g1141), .Q(n443) );
  AND2X1 U2719 ( .IN1(g109), .IN2(g1121), .Q(n435) );
  INVX0 U2720 ( .INP(n2704), .ZN(n395) );
  OR2X1 U2721 ( .IN1(n505), .IN2(n1708), .Q(n2704) );
  INVX0 U2722 ( .INP(n2705), .ZN(n363) );
  OR2X1 U2723 ( .IN1(n505), .IN2(n1705), .Q(n2705) );
  AND2X1 U2724 ( .IN1(n804), .IN2(n2706), .Q(n324) );
  INVX0 U2725 ( .INP(n2707), .ZN(n319) );
  OR2X1 U2726 ( .IN1(n2708), .IN2(n2463), .Q(n2707) );
  AND2X1 U2727 ( .IN1(n2709), .IN2(n2710), .Q(n2708) );
  OR2X1 U2728 ( .IN1(g750), .IN2(n1647), .Q(n2709) );
  INVX0 U2729 ( .INP(n2711), .ZN(n274) );
  AND2X1 U2730 ( .IN1(n2712), .IN2(g986), .Q(n2494) );
  INVX0 U2731 ( .INP(n2713), .ZN(n227) );
  INVX0 U2732 ( .INP(n2714), .ZN(n192) );
  OR2X1 U2733 ( .IN1(n505), .IN2(n1706), .Q(n2714) );
  INVX0 U2734 ( .INP(n2715), .ZN(n167) );
  OR4X1 U2735 ( .IN1(n2716), .IN2(n2717), .IN3(g42), .IN4(n2718), .Q(n1588) );
  OR3X1 U2736 ( .IN1(n2718), .IN2(n2717), .IN3(n2719), .Q(n1587) );
  OR2X1 U2737 ( .IN1(n2719), .IN2(n2720), .Q(n1586) );
  OR3X1 U2738 ( .IN1(g42), .IN2(n2716), .IN3(n2720), .Q(n1585) );
  OR3X1 U2739 ( .IN1(g46), .IN2(n2721), .IN3(n2722), .Q(n2720) );
  OR2X1 U2740 ( .IN1(n2451), .IN2(n2452), .Q(n1214) );
  INVX0 U2741 ( .INP(n2723), .ZN(n12) );
  INVX0 U2742 ( .INP(n2724), .ZN(n119) );
  AND2X1 U2743 ( .IN1(n2725), .IN2(n2726), .Q(n2724) );
  OR2X1 U2744 ( .IN1(n2727), .IN2(n2450), .Q(n2725) );
  AND2X1 U2745 ( .IN1(n2728), .IN2(n1709), .Q(n2727) );
  INVX0 U2746 ( .INP(n2729), .ZN(n118) );
  AND3X1 U2747 ( .IN1(n2730), .IN2(n2731), .IN3(n2726), .Q(n2729) );
  OR2X1 U2748 ( .IN1(g627), .IN2(n1612), .Q(n2731) );
  OR2X1 U2749 ( .IN1(n2447), .IN2(n2732), .Q(n1153) );
  OR2X1 U2750 ( .IN1(n2432), .IN2(n2733), .Q(n1151) );
  INVX0 U2751 ( .INP(n2734), .ZN(n114) );
  INVX0 U2752 ( .INP(n2735), .ZN(n112) );
  OR4X1 U2753 ( .IN1(n2736), .IN2(n1626), .IN3(n2737), .IN4(n2738), .Q(n2735)
         );
  INVX0 U2754 ( .INP(n2739), .ZN(n2738) );
  AND4X1 U2755 ( .IN1(g1690), .IN2(g1707), .IN3(g1806), .IN4(g1801), .Q(n2739)
         );
  OR2X1 U2756 ( .IN1(g1781), .IN2(n2740), .Q(n2737) );
  OR2X1 U2757 ( .IN1(n2446), .IN2(n2741), .Q(n1099) );
  OR2X1 U2758 ( .IN1(n2431), .IN2(n2742), .Q(n1097) );
  AND3X1 U2759 ( .IN1(n2743), .IN2(n2744), .IN3(n2745), .Q(n106) );
  INVX0 U2760 ( .INP(n1098), .ZN(n2744) );
  INVX0 U2761 ( .INP(n2746), .ZN(n1) );
  AND2X1 U2762 ( .IN1(n2391), .IN2(n2465), .Q(n2746) );
  AND2X1 U2763 ( .IN1(g18), .IN2(n2747), .Q(g9721) );
  XOR2X1 U2764 ( .IN1(n1609), .IN2(n2748), .Q(n2747) );
  AND2X1 U2765 ( .IN1(n2749), .IN2(n2750), .Q(n2748) );
  OR2X1 U2766 ( .IN1(n2751), .IN2(n2752), .Q(n2749) );
  AND2X1 U2767 ( .IN1(n1645), .IN2(n2753), .Q(n2751) );
  OR2X1 U2768 ( .IN1(n804), .IN2(n2754), .Q(n2753) );
  AND3X1 U2769 ( .IN1(n2755), .IN2(n2756), .IN3(g18), .Q(g9555) );
  OR2X1 U2770 ( .IN1(n806), .IN2(g1834), .Q(n2756) );
  INVX0 U2771 ( .INP(n2757), .ZN(n2755) );
  AND3X1 U2772 ( .IN1(n808), .IN2(n926), .IN3(g1834), .Q(n2757) );
  OR2X1 U2773 ( .IN1(n2758), .IN2(g1840), .Q(n808) );
  AND2X1 U2774 ( .IN1(n809), .IN2(n2759), .Q(n2758) );
  OR3X1 U2775 ( .IN1(g31), .IN2(g30), .IN3(n2721), .Q(g9451) );
  AND3X1 U2776 ( .IN1(n2760), .IN2(n2761), .IN3(g18), .Q(g9272) );
  OR2X1 U2777 ( .IN1(n1605), .IN2(n2762), .Q(n2761) );
  INVX0 U2778 ( .INP(n2763), .ZN(n2760) );
  AND3X1 U2779 ( .IN1(n2764), .IN2(n2762), .IN3(n1605), .Q(n2763) );
  OR2X1 U2780 ( .IN1(n2765), .IN2(n2759), .Q(n2762) );
  AND3X1 U2781 ( .IN1(n2766), .IN2(n2767), .IN3(n2768), .Q(n2765) );
  OR2X1 U2782 ( .IN1(n1643), .IN2(n817), .Q(n2768) );
  AND2X1 U2783 ( .IN1(g18), .IN2(n2769), .Q(g9269) );
  XOR2X1 U2784 ( .IN1(n1643), .IN2(n2770), .Q(n2769) );
  AND2X1 U2785 ( .IN1(n2771), .IN2(n2772), .Q(n2770) );
  OR2X1 U2786 ( .IN1(n2759), .IN2(n2773), .Q(n2772) );
  AND2X1 U2787 ( .IN1(n2767), .IN2(n822), .Q(n2773) );
  AND2X1 U2788 ( .IN1(g18), .IN2(n2774), .Q(g9266) );
  XOR2X1 U2789 ( .IN1(n1608), .IN2(n2775), .Q(n2774) );
  AND2X1 U2790 ( .IN1(n2776), .IN2(n2771), .Q(n2775) );
  OR3X1 U2791 ( .IN1(n817), .IN2(g1822), .IN3(n2759), .Q(n2771) );
  OR2X1 U2792 ( .IN1(n2777), .IN2(n2759), .Q(n2776) );
  INVX0 U2793 ( .INP(n812), .ZN(n2759) );
  AND2X1 U2794 ( .IN1(n2778), .IN2(n2779), .Q(n2777) );
  AND3X1 U2795 ( .IN1(n2780), .IN2(n2781), .IN3(g18), .Q(g9150) );
  OR2X1 U2796 ( .IN1(n1593), .IN2(n2782), .Q(n2781) );
  INVX0 U2797 ( .INP(n2783), .ZN(n2782) );
  OR3X1 U2798 ( .IN1(n2784), .IN2(n2783), .IN3(g605), .Q(n2780) );
  OR2X1 U2799 ( .IN1(n2785), .IN2(n2786), .Q(n2783) );
  AND2X1 U2800 ( .IN1(n804), .IN2(n2787), .Q(n2786) );
  OR3X1 U2801 ( .IN1(n2788), .IN2(n2789), .IN3(n2790), .Q(n2787) );
  AND2X1 U2802 ( .IN1(n2791), .IN2(g599), .Q(n2790) );
  AND2X1 U2803 ( .IN1(g18), .IN2(n2792), .Q(g9124) );
  XOR2X1 U2804 ( .IN1(n836), .IN2(n1644), .Q(n2792) );
  AND2X1 U2805 ( .IN1(g18), .IN2(n2793), .Q(g9110) );
  XOR2X1 U2806 ( .IN1(n1607), .IN2(n2794), .Q(n2793) );
  AND3X1 U2807 ( .IN1(n2795), .IN2(n837), .IN3(n2796), .Q(n2794) );
  OR2X1 U2808 ( .IN1(n2797), .IN2(n2798), .Q(n2796) );
  OR3X1 U2809 ( .IN1(g599), .IN2(n2799), .IN3(n2798), .Q(n837) );
  OR2X1 U2810 ( .IN1(n2800), .IN2(n2801), .Q(g8973) );
  AND2X1 U2811 ( .IN1(n2802), .IN2(n2803), .Q(n2800) );
  XOR2X1 U2812 ( .IN1(n2804), .IN2(n1615), .Q(n2802) );
  OR2X1 U2813 ( .IN1(n2805), .IN2(n2806), .Q(n2804) );
  AND2X1 U2814 ( .IN1(n2429), .IN2(n2807), .Q(n2805) );
  OR2X1 U2815 ( .IN1(n2808), .IN2(n2809), .Q(g8945) );
  AND2X1 U2816 ( .IN1(n2810), .IN2(n2811), .Q(n2808) );
  XNOR2X1 U2817 ( .IN1(n1697), .IN2(n2812), .Q(n2811) );
  OR2X1 U2818 ( .IN1(n2813), .IN2(n2814), .Q(n2812) );
  AND2X1 U2819 ( .IN1(n2815), .IN2(g1950), .Q(n2814) );
  AND2X1 U2820 ( .IN1(n2816), .IN2(n2817), .Q(n2813) );
  OR2X1 U2821 ( .IN1(n2691), .IN2(n2723), .Q(n2817) );
  AND3X1 U2822 ( .IN1(g1936), .IN2(n2818), .IN3(n921), .Q(n2723) );
  AND3X1 U2823 ( .IN1(n2819), .IN2(n2820), .IN3(n1694), .Q(n2691) );
  OR2X1 U2824 ( .IN1(n2821), .IN2(n2809), .Q(g8944) );
  AND2X1 U2825 ( .IN1(n2810), .IN2(n2822), .Q(n2821) );
  XOR2X1 U2826 ( .IN1(g1936), .IN2(n2823), .Q(n2822) );
  OR2X1 U2827 ( .IN1(n2824), .IN2(n2825), .Q(n2823) );
  AND2X1 U2828 ( .IN1(n2815), .IN2(g1941), .Q(n2825) );
  AND2X1 U2829 ( .IN1(n2816), .IN2(n2826), .Q(n2824) );
  OR2X1 U2830 ( .IN1(n2827), .IN2(n2828), .Q(n2826) );
  AND2X1 U2831 ( .IN1(n2820), .IN2(n2819), .Q(n2828) );
  AND4X1 U2832 ( .IN1(n2829), .IN2(n1675), .IN3(n2420), .IN4(n2830), .Q(n2819)
         );
  AND2X1 U2833 ( .IN1(n2421), .IN2(n2444), .Q(n2830) );
  AND2X1 U2834 ( .IN1(n921), .IN2(n2818), .Q(n2827) );
  AND4X1 U2835 ( .IN1(g1900), .IN2(n2831), .IN3(g1909), .IN4(g1918), .Q(n2818)
         );
  OR2X1 U2836 ( .IN1(n2832), .IN2(n2809), .Q(g8943) );
  AND2X1 U2837 ( .IN1(n2833), .IN2(n2810), .Q(n2832) );
  XNOR2X1 U2838 ( .IN1(n1663), .IN2(n2834), .Q(n2833) );
  AND3X1 U2839 ( .IN1(n2835), .IN2(n2836), .IN3(n2837), .Q(n2834) );
  OR2X1 U2840 ( .IN1(n2838), .IN2(g1887), .Q(n2836) );
  OR2X1 U2841 ( .IN1(n2815), .IN2(n2839), .Q(n2835) );
  XNOR2X1 U2842 ( .IN1(n2820), .IN2(n1616), .Q(n2839) );
  OR2X1 U2843 ( .IN1(n2840), .IN2(n2809), .Q(g8941) );
  AND2X1 U2844 ( .IN1(n2841), .IN2(n2810), .Q(n2840) );
  XOR2X1 U2845 ( .IN1(n2842), .IN2(n2444), .Q(n2841) );
  OR2X1 U2849 ( .IN1(n2843), .IN2(n2844), .Q(n2842) );
  AND3X1 U2850 ( .IN1(n2845), .IN2(n2846), .IN3(n2847), .Q(n2843) );
  OR2X1 U2851 ( .IN1(n2838), .IN2(n2329), .Q(n2847) );
  OR4X1 U2852 ( .IN1(n2420), .IN2(n1675), .IN3(n2848), .IN4(n2421), .Q(n2846)
         );
  OR4X1 U2853 ( .IN1(g1900), .IN2(g1918), .IN3(n2849), .IN4(g1909), .Q(n2845)
         );
  OR2X1 U2854 ( .IN1(n2850), .IN2(n2809), .Q(g8940) );
  AND2X1 U2855 ( .IN1(n2851), .IN2(n2810), .Q(n2850) );
  XOR2X1 U2856 ( .IN1(g1918), .IN2(n2852), .Q(n2851) );
  AND2X1 U2857 ( .IN1(n2853), .IN2(n2837), .Q(n2852) );
  OR3X1 U2858 ( .IN1(n2854), .IN2(n2855), .IN3(n2856), .Q(n2853) );
  AND2X1 U2862 ( .IN1(n2815), .IN2(g1923), .Q(n2856) );
  AND3X1 U2863 ( .IN1(n2857), .IN2(n1675), .IN3(n2421), .Q(n2855) );
  AND3X1 U2864 ( .IN1(n2858), .IN2(g1900), .IN3(g1909), .Q(n2854) );
  INVX0 U2865 ( .INP(n2848), .ZN(n2858) );
  OR2X1 U2866 ( .IN1(n2859), .IN2(n2809), .Q(g8939) );
  AND2X1 U2868 ( .IN1(n2860), .IN2(n2810), .Q(n2859) );
  XOR2X1 U2869 ( .IN1(n2861), .IN2(n2421), .Q(n2860) );
  OR2X1 U2870 ( .IN1(n2862), .IN2(n2844), .Q(n2861) );
  AND3X1 U2871 ( .IN1(n2863), .IN2(n2864), .IN3(n2865), .Q(n2862) );
  OR2X1 U2872 ( .IN1(n2838), .IN2(n2326), .Q(n2865) );
  OR2X1 U2873 ( .IN1(n1675), .IN2(n2848), .Q(n2864) );
  OR2X1 U2874 ( .IN1(g1900), .IN2(n2849), .Q(n2863) );
  OR2X1 U2875 ( .IN1(n2866), .IN2(n2809), .Q(g8938) );
  AND2X1 U2876 ( .IN1(n2867), .IN2(n2810), .Q(n2866) );
  XOR2X1 U2877 ( .IN1(n2868), .IN2(n1675), .Q(n2867) );
  OR2X1 U2878 ( .IN1(n2869), .IN2(n2844), .Q(n2868) );
  AND3X1 U2880 ( .IN1(n2848), .IN2(n2849), .IN3(n2870), .Q(n2869) );
  OR2X1 U2903 ( .IN1(n2838), .IN2(n2436), .Q(n2870) );
  INVX0 U2904 ( .INP(n2857), .ZN(n2849) );
  AND3X1 U2905 ( .IN1(n2829), .IN2(n2820), .IN3(n2838), .Q(n2857) );
  AND3X1 U2906 ( .IN1(n1616), .IN2(n1657), .IN3(n1663), .Q(n2829) );
  OR3X1 U2907 ( .IN1(n1657), .IN2(n2871), .IN3(n2815), .Q(n2848) );
  OR2X1 U2908 ( .IN1(n2872), .IN2(n2809), .Q(g8937) );
  AND2X1 U2909 ( .IN1(n2810), .IN2(n2873), .Q(n2872) );
  XNOR2X1 U2910 ( .IN1(n1657), .IN2(n2874), .Q(n2873) );
  OR2X1 U2911 ( .IN1(n2875), .IN2(n2876), .Q(n2874) );
  AND2X1 U2912 ( .IN1(n2815), .IN2(g1896), .Q(n2876) );
  AND2X1 U2913 ( .IN1(n2816), .IN2(n2877), .Q(n2875) );
  OR2X1 U2914 ( .IN1(n2878), .IN2(n2831), .Q(n2877) );
  INVX0 U2915 ( .INP(n2871), .ZN(n2831) );
  OR3X1 U2916 ( .IN1(n1663), .IN2(n1616), .IN3(n2820), .Q(n2871) );
  AND3X1 U2917 ( .IN1(n1663), .IN2(n1616), .IN3(n2820), .Q(n2878) );
  AND3X1 U2918 ( .IN1(n2767), .IN2(n2766), .IN3(n2879), .Q(n2820) );
  OR2X1 U2919 ( .IN1(g1828), .IN2(n2778), .Q(n2766) );
  AND2X1 U2920 ( .IN1(n2837), .IN2(n2838), .Q(n2816) );
  OR2X1 U2921 ( .IN1(n2880), .IN2(n2801), .Q(g8926) );
  AND2X1 U2922 ( .IN1(n2803), .IN2(n2881), .Q(n2880) );
  XNOR2X1 U2923 ( .IN1(n1696), .IN2(n898), .Q(n2881) );
  OR2X1 U2924 ( .IN1(n2882), .IN2(n2883), .Q(n898) );
  AND2X1 U2925 ( .IN1(n2807), .IN2(g736), .Q(n2883) );
  AND2X1 U2926 ( .IN1(n2884), .IN2(n2885), .Q(n2882) );
  OR2X1 U2927 ( .IN1(n2687), .IN2(n2699), .Q(n2885) );
  AND3X1 U2928 ( .IN1(g722), .IN2(n2886), .IN3(n967), .Q(n2699) );
  AND3X1 U2929 ( .IN1(n2887), .IN2(n2888), .IN3(n1693), .Q(n2687) );
  OR2X1 U2930 ( .IN1(n2889), .IN2(n2801), .Q(g8923) );
  AND2X1 U2931 ( .IN1(n2803), .IN2(n2890), .Q(n2889) );
  XOR2X1 U2932 ( .IN1(g722), .IN2(n2891), .Q(n2890) );
  OR2X1 U2933 ( .IN1(n2892), .IN2(n2893), .Q(n2891) );
  AND2X1 U2934 ( .IN1(n2807), .IN2(g727), .Q(n2893) );
  AND2X1 U2935 ( .IN1(n2884), .IN2(n2894), .Q(n2892) );
  OR2X1 U2936 ( .IN1(n2895), .IN2(n2896), .Q(n2894) );
  AND2X1 U2937 ( .IN1(n2888), .IN2(n2887), .Q(n2896) );
  AND4X1 U2938 ( .IN1(n2897), .IN2(n1676), .IN3(n2418), .IN4(n2898), .Q(n2887)
         );
  AND2X1 U2939 ( .IN1(n2419), .IN2(n2445), .Q(n2898) );
  AND2X1 U2940 ( .IN1(n967), .IN2(n2886), .Q(n2895) );
  AND4X1 U2941 ( .IN1(g686), .IN2(n2899), .IN3(g695), .IN4(g704), .Q(n2886) );
  OR2X1 U2942 ( .IN1(n2900), .IN2(n2801), .Q(g8922) );
  AND2X1 U2943 ( .IN1(n2901), .IN2(n2803), .Q(n2900) );
  XNOR2X1 U2944 ( .IN1(n1662), .IN2(n2902), .Q(n2901) );
  AND3X1 U2945 ( .IN1(n2903), .IN2(n2904), .IN3(n2905), .Q(n2902) );
  OR2X1 U2946 ( .IN1(n2906), .IN2(g673), .Q(n2904) );
  OR2X1 U2947 ( .IN1(n2807), .IN2(n2907), .Q(n2903) );
  XOR2X1 U2948 ( .IN1(n2908), .IN2(n1615), .Q(n2907) );
  OR2X1 U2949 ( .IN1(n2909), .IN2(n2809), .Q(g8921) );
  AND4X1 U2950 ( .IN1(n2910), .IN2(n916), .IN3(n2764), .IN4(n2767), .Q(n2809)
         );
  AND2X1 U2951 ( .IN1(n2911), .IN2(n2810), .Q(n2909) );
  INVX0 U2952 ( .INP(n2910), .ZN(n2810) );
  OR2X1 U2953 ( .IN1(n812), .IN2(n2912), .Q(n2910) );
  XNOR2X1 U2954 ( .IN1(n1616), .IN2(n2913), .Q(n2911) );
  AND2X1 U2955 ( .IN1(n2837), .IN2(n2914), .Q(n2913) );
  OR2X1 U2956 ( .IN1(n2838), .IN2(g1878), .Q(n2914) );
  INVX0 U2957 ( .INP(n2844), .ZN(n2837) );
  AND2X1 U2958 ( .IN1(n918), .IN2(n2838), .Q(n2844) );
  INVX0 U2959 ( .INP(n2815), .ZN(n2838) );
  OR2X1 U2960 ( .IN1(n2915), .IN2(n257), .Q(n2815) );
  AND2X1 U2961 ( .IN1(n926), .IN2(g1840), .Q(n2915) );
  OR2X1 U2962 ( .IN1(n493), .IN2(n2916), .Q(n918) );
  AND2X1 U2963 ( .IN1(n2917), .IN2(n2779), .Q(n2916) );
  INVX0 U2964 ( .INP(n809), .ZN(n2779) );
  AND3X1 U2965 ( .IN1(g1834), .IN2(g1814), .IN3(n2442), .Q(n809) );
  OR2X1 U2966 ( .IN1(n2918), .IN2(n1682), .Q(n2917) );
  AND2X1 U2967 ( .IN1(n1643), .IN2(n1605), .Q(n2918) );
  OR2X1 U2968 ( .IN1(n2919), .IN2(n2801), .Q(g8920) );
  AND2X1 U2969 ( .IN1(n2920), .IN2(n2803), .Q(n2919) );
  XOR2X1 U2970 ( .IN1(n2445), .IN2(n931), .Q(n2920) );
  OR2X1 U2971 ( .IN1(n2921), .IN2(n2806), .Q(n931) );
  AND3X1 U2972 ( .IN1(n2922), .IN2(n2923), .IN3(n2924), .Q(n2921) );
  OR2X1 U2973 ( .IN1(n2906), .IN2(n2279), .Q(n2924) );
  OR4X1 U2974 ( .IN1(n2418), .IN2(n1676), .IN3(n2925), .IN4(n2419), .Q(n2923)
         );
  OR4X1 U2975 ( .IN1(g686), .IN2(g704), .IN3(n2926), .IN4(g695), .Q(n2922) );
  OR2X1 U2976 ( .IN1(n2927), .IN2(n2801), .Q(g8889) );
  AND2X1 U2977 ( .IN1(n2928), .IN2(n2803), .Q(n2927) );
  XOR2X1 U2978 ( .IN1(g704), .IN2(n938), .Q(n2928) );
  INVX0 U2979 ( .INP(n2929), .ZN(n938) );
  OR2X1 U2980 ( .IN1(n2806), .IN2(n2930), .Q(n2929) );
  AND3X1 U2981 ( .IN1(n2931), .IN2(n2932), .IN3(n2933), .Q(n2930) );
  OR2X1 U2982 ( .IN1(n1719), .IN2(n2906), .Q(n2933) );
  OR3X1 U2983 ( .IN1(n1676), .IN2(n2925), .IN3(n2419), .Q(n2932) );
  OR3X1 U2984 ( .IN1(g686), .IN2(n2926), .IN3(g695), .Q(n2931) );
  OR2X1 U2985 ( .IN1(n2934), .IN2(n2801), .Q(g8887) );
  AND2X1 U2986 ( .IN1(n2935), .IN2(n2803), .Q(n2934) );
  XOR2X1 U2987 ( .IN1(n2936), .IN2(n2419), .Q(n2935) );
  OR2X1 U2988 ( .IN1(n2937), .IN2(n2806), .Q(n2936) );
  AND3X1 U2989 ( .IN1(n2938), .IN2(n2939), .IN3(n2940), .Q(n2937) );
  OR2X1 U2990 ( .IN1(n2906), .IN2(n2366), .Q(n2940) );
  OR2X1 U2991 ( .IN1(n1676), .IN2(n2925), .Q(n2939) );
  OR2X1 U2992 ( .IN1(g686), .IN2(n2926), .Q(n2938) );
  OR2X1 U2993 ( .IN1(n2941), .IN2(n2801), .Q(g8885) );
  AND2X1 U2994 ( .IN1(n2942), .IN2(n2803), .Q(n2941) );
  XOR2X1 U2995 ( .IN1(n2943), .IN2(n1676), .Q(n2942) );
  OR2X1 U2996 ( .IN1(n2944), .IN2(n2806), .Q(n2943) );
  AND3X1 U2997 ( .IN1(n2925), .IN2(n2926), .IN3(n2945), .Q(n2944) );
  OR2X1 U2998 ( .IN1(n2906), .IN2(n2435), .Q(n2945) );
  INVX0 U2999 ( .INP(n2946), .ZN(n2926) );
  AND3X1 U3000 ( .IN1(n2897), .IN2(n2888), .IN3(n2906), .Q(n2946) );
  AND3X1 U3001 ( .IN1(n1615), .IN2(n1656), .IN3(n1662), .Q(n2897) );
  OR3X1 U3002 ( .IN1(n1656), .IN2(n2947), .IN3(n2807), .Q(n2925) );
  OR2X1 U3003 ( .IN1(n2948), .IN2(n2801), .Q(g8883) );
  INVX0 U3004 ( .INP(n2949), .ZN(n2801) );
  OR4X1 U3005 ( .IN1(n2950), .IN2(n2706), .IN3(n2784), .IN4(n2803), .Q(n2949)
         );
  AND2X1 U3006 ( .IN1(n2803), .IN2(n2951), .Q(n2948) );
  XNOR2X1 U3007 ( .IN1(n1656), .IN2(n2952), .Q(n2951) );
  OR2X1 U3008 ( .IN1(n2953), .IN2(n2954), .Q(n2952) );
  AND2X1 U3009 ( .IN1(n2807), .IN2(g682), .Q(n2954) );
  AND2X1 U3010 ( .IN1(n2884), .IN2(n2955), .Q(n2953) );
  OR2X1 U3011 ( .IN1(n2956), .IN2(n2899), .Q(n2955) );
  INVX0 U3012 ( .INP(n2947), .ZN(n2899) );
  OR3X1 U3013 ( .IN1(n1662), .IN2(n1615), .IN3(n2888), .Q(n2947) );
  AND3X1 U3014 ( .IN1(n1662), .IN2(n1615), .IN3(n2888), .Q(n2956) );
  INVX0 U3015 ( .INP(n2908), .ZN(n2888) );
  OR3X1 U3016 ( .IN1(n2788), .IN2(n2789), .IN3(n2957), .Q(n2908) );
  AND2X1 U3017 ( .IN1(n2958), .IN2(n1593), .Q(n2789) );
  AND2X1 U3018 ( .IN1(n2905), .IN2(n2906), .Q(n2884) );
  INVX0 U3019 ( .INP(n2806), .ZN(n2905) );
  AND2X1 U3020 ( .IN1(n958), .IN2(n2906), .Q(n2806) );
  INVX0 U3021 ( .INP(n2807), .ZN(n2906) );
  OR2X1 U3022 ( .IN1(n2959), .IN2(n2960), .Q(n2807) );
  AND2X1 U3023 ( .IN1(n2961), .IN2(g617), .Q(n2960) );
  OR2X1 U3024 ( .IN1(n2962), .IN2(n2752), .Q(n958) );
  AND2X1 U3025 ( .IN1(n2963), .IN2(n2754), .Q(n2962) );
  OR2X1 U3026 ( .IN1(n2964), .IN2(n1692), .Q(n2963) );
  AND2X1 U3027 ( .IN1(n1593), .IN2(n1644), .Q(n2964) );
  AND2X1 U3028 ( .IN1(n2798), .IN2(n2965), .Q(n2803) );
  AND2X1 U3029 ( .IN1(n2966), .IN2(n2965), .Q(g8820) );
  OR2X1 U3030 ( .IN1(n2967), .IN2(n2785), .Q(n2966) );
  INVX0 U3031 ( .INP(n2750), .ZN(n2785) );
  OR2X1 U3032 ( .IN1(n2795), .IN2(g622), .Q(n2750) );
  AND2X1 U3033 ( .IN1(n2795), .IN2(g622), .Q(n2967) );
  OR2X1 U3034 ( .IN1(n2798), .IN2(n2754), .Q(n2795) );
  INVX0 U3035 ( .INP(n2950), .ZN(n2754) );
  AND3X1 U3036 ( .IN1(g611), .IN2(g591), .IN3(n1645), .Q(n2950) );
  INVX0 U3037 ( .INP(n804), .ZN(n2798) );
  OR2X1 U3038 ( .IN1(n2968), .IN2(n2969), .Q(g8779) );
  AND2X1 U3039 ( .IN1(n2970), .IN2(n2971), .Q(n2969) );
  AND2X1 U3040 ( .IN1(n371), .IN2(g1636), .Q(n2968) );
  OR2X1 U3041 ( .IN1(n2972), .IN2(n2973), .Q(g8777) );
  AND2X1 U3042 ( .IN1(n2974), .IN2(n2971), .Q(n2973) );
  AND2X1 U3043 ( .IN1(n371), .IN2(g1633), .Q(n2972) );
  OR2X1 U3044 ( .IN1(n2975), .IN2(n2976), .Q(g8776) );
  AND2X1 U3045 ( .IN1(n2977), .IN2(n2971), .Q(n2976) );
  AND2X1 U3046 ( .IN1(n371), .IN2(g1630), .Q(n2975) );
  AND2X1 U3047 ( .IN1(n2978), .IN2(g109), .Q(g8775) );
  XNOR2X1 U3048 ( .IN1(n2402), .IN2(n2979), .Q(n2978) );
  OR2X1 U3049 ( .IN1(n2980), .IN2(n2981), .Q(g8774) );
  AND2X1 U3050 ( .IN1(n2979), .IN2(n2971), .Q(n2981) );
  OR2X1 U3051 ( .IN1(n2982), .IN2(n2983), .Q(n2979) );
  AND2X1 U3052 ( .IN1(n2984), .IN2(n2985), .Q(n2982) );
  XNOR2X1 U3053 ( .IN1(n1706), .IN2(n2986), .Q(n2984) );
  AND3X1 U3054 ( .IN1(n1654), .IN2(g1107), .IN3(n2987), .Q(n2986) );
  AND2X1 U3055 ( .IN1(n371), .IN2(g1627), .Q(n2980) );
  OR2X1 U3056 ( .IN1(n2988), .IN2(n2989), .Q(g8773) );
  AND2X1 U3057 ( .IN1(n2990), .IN2(n2971), .Q(n2989) );
  AND2X1 U3058 ( .IN1(n371), .IN2(g1624), .Q(n2988) );
  AND2X1 U3059 ( .IN1(n2991), .IN2(g109), .Q(g8772) );
  XNOR2X1 U3060 ( .IN1(n2403), .IN2(n2977), .Q(n2991) );
  OR2X1 U3061 ( .IN1(n2992), .IN2(n2993), .Q(n2977) );
  AND2X1 U3062 ( .IN1(n2994), .IN2(n2985), .Q(n2992) );
  XOR2X1 U3063 ( .IN1(g1137), .IN2(n2995), .Q(n2994) );
  AND3X1 U3064 ( .IN1(g1107), .IN2(g1101), .IN3(n2987), .Q(n2995) );
  OR2X1 U3065 ( .IN1(n2996), .IN2(n2997), .Q(g8771) );
  AND2X1 U3066 ( .IN1(n2998), .IN2(n2971), .Q(n2997) );
  AND2X1 U3067 ( .IN1(n371), .IN2(g1621), .Q(n2996) );
  OR2X1 U3068 ( .IN1(n2999), .IN2(n3000), .Q(g8770) );
  AND2X1 U3069 ( .IN1(n3001), .IN2(n2971), .Q(n3000) );
  AND2X1 U3070 ( .IN1(n371), .IN2(g1615), .Q(n2999) );
  AND2X1 U3071 ( .IN1(n3002), .IN2(g109), .Q(g8769) );
  XNOR2X1 U3072 ( .IN1(n2404), .IN2(n3001), .Q(n3002) );
  OR2X1 U3073 ( .IN1(n3003), .IN2(n3004), .Q(n3001) );
  AND2X1 U3074 ( .IN1(n3005), .IN2(n2985), .Q(n3003) );
  XOR2X1 U3075 ( .IN1(n3006), .IN2(g1121), .Q(n3005) );
  AND2X1 U3076 ( .IN1(n3007), .IN2(n2987), .Q(n3006) );
  AND2X1 U3077 ( .IN1(n3008), .IN2(g109), .Q(g8768) );
  XNOR2X1 U3078 ( .IN1(n2405), .IN2(n2974), .Q(n3008) );
  OR2X1 U3079 ( .IN1(n3009), .IN2(n3010), .Q(n2974) );
  AND2X1 U3080 ( .IN1(n3011), .IN2(n2985), .Q(n3009) );
  XOR2X1 U3081 ( .IN1(n3012), .IN2(g1141), .Q(n3011) );
  AND2X1 U3082 ( .IN1(n3013), .IN2(n1654), .Q(n3012) );
  AND2X1 U3083 ( .IN1(n3014), .IN2(g109), .Q(g8767) );
  XOR2X1 U3084 ( .IN1(g1403), .IN2(n2998), .Q(n3014) );
  OR2X1 U3085 ( .IN1(n3015), .IN2(n3021), .Q(n2998) );
  AND2X1 U3086 ( .IN1(n3028), .IN2(n2985), .Q(n3015) );
  XNOR2X1 U3087 ( .IN1(n1708), .IN2(n3032), .Q(n3028) );
  AND2X1 U3088 ( .IN1(n3039), .IN2(n1654), .Q(n3032) );
  AND2X1 U3089 ( .IN1(n3043), .IN2(g109), .Q(g8766) );
  XNOR2X1 U3091 ( .IN1(n2473), .IN2(n2970), .Q(n3043) );
  OR2X1 U3093 ( .IN1(n3049), .IN2(n3052), .Q(n2970) );
  AND2X1 U3095 ( .IN1(n3060), .IN2(n2985), .Q(n3049) );
  XOR2X1 U3097 ( .IN1(g1145), .IN2(n3063), .Q(n3060) );
  AND2X1 U3099 ( .IN1(n3013), .IN2(g1101), .Q(n3063) );
  AND3X1 U3100 ( .IN1(g1110), .IN2(n1614), .IN3(n1658), .Q(n3013) );
  AND2X1 U3101 ( .IN1(n3066), .IN2(g109), .Q(g8765) );
  XNOR2X1 U3102 ( .IN1(n2474), .IN2(n2990), .Q(n3066) );
  OR2X1 U3103 ( .IN1(n3067), .IN2(n3068), .Q(n2990) );
  AND2X1 U3104 ( .IN1(n3069), .IN2(n2985), .Q(n3067) );
  XNOR2X1 U3105 ( .IN1(n1705), .IN2(n3070), .Q(n3069) );
  AND2X1 U3106 ( .IN1(n3039), .IN2(g1101), .Q(n3070) );
  AND3X1 U3107 ( .IN1(g1107), .IN2(n1658), .IN3(n1677), .Q(n3039) );
  OR3X1 U3108 ( .IN1(n2784), .IN2(n3071), .IN3(n3072), .Q(g8649) );
  AND2X1 U3109 ( .IN1(n124), .IN2(g664), .Q(n3072) );
  OR2X1 U3110 ( .IN1(n3073), .IN2(n3074), .Q(g8631) );
  AND2X1 U3111 ( .IN1(n2784), .IN2(n3075), .Q(n3074) );
  OR3X1 U3112 ( .IN1(n1716), .IN2(n3076), .IN3(n3077), .Q(n3075) );
  AND2X1 U3113 ( .IN1(n3078), .IN2(n3079), .Q(n3077) );
  OR2X1 U3114 ( .IN1(n1622), .IN2(n2432), .Q(n3078) );
  AND2X1 U3115 ( .IN1(n3080), .IN2(n3081), .Q(n3076) );
  OR2X1 U3116 ( .IN1(n2396), .IN2(n2431), .Q(n3081) );
  OR2X1 U3117 ( .IN1(n2395), .IN2(n2428), .Q(n3080) );
  AND2X1 U3118 ( .IN1(n3082), .IN2(n2965), .Q(n3073) );
  OR2X1 U3119 ( .IN1(n3083), .IN2(n3084), .Q(n3082) );
  AND2X1 U3120 ( .IN1(n2788), .IN2(n1713), .Q(n3084) );
  AND2X1 U3121 ( .IN1(n3085), .IN2(g636), .Q(n3083) );
  OR3X1 U3122 ( .IN1(n3086), .IN2(n2715), .IN3(n3087), .Q(n3085) );
  XOR2X1 U3123 ( .IN1(n3088), .IN2(n3089), .Q(n3087) );
  AND2X1 U3125 ( .IN1(g255), .IN2(g622), .Q(n3089) );
  OR2X1 U3126 ( .IN1(n3090), .IN2(n3091), .Q(n3088) );
  AND3X1 U3127 ( .IN1(n1609), .IN2(n2799), .IN3(n1692), .Q(n3091) );
  AND2X1 U3128 ( .IN1(n2797), .IN2(g639), .Q(n3090) );
  OR2X1 U3129 ( .IN1(n2497), .IN2(n1874), .Q(n2715) );
  AND3X1 U3130 ( .IN1(n1609), .IN2(n3092), .IN3(n3093), .Q(n3086) );
  AND3X1 U3131 ( .IN1(n3094), .IN2(n2797), .IN3(n2799), .Q(n3093) );
  INVX0 U3132 ( .INP(n3095), .ZN(n3094) );
  OR2X1 U3133 ( .IN1(n3096), .IN2(n3097), .Q(g8566) );
  AND2X1 U3134 ( .IN1(g1690), .IN2(g1687), .Q(n3097) );
  AND2X1 U3135 ( .IN1(n1653), .IN2(g1669), .Q(n3096) );
  OR2X1 U3136 ( .IN1(n3098), .IN2(n3099), .Q(g8565) );
  AND2X1 U3137 ( .IN1(g1690), .IN2(g1684), .Q(n3099) );
  AND2X1 U3138 ( .IN1(n1653), .IN2(g1666), .Q(n3098) );
  OR2X1 U3139 ( .IN1(n3100), .IN2(n3101), .Q(g8564) );
  AND2X1 U3140 ( .IN1(g1690), .IN2(g1681), .Q(n3101) );
  AND2X1 U3141 ( .IN1(n1653), .IN2(g1663), .Q(n3100) );
  OR2X1 U3142 ( .IN1(n3102), .IN2(n3103), .Q(g8563) );
  AND2X1 U3143 ( .IN1(g1690), .IN2(g1678), .Q(n3103) );
  AND2X1 U3144 ( .IN1(n1653), .IN2(g1660), .Q(n3102) );
  OR2X1 U3145 ( .IN1(n3104), .IN2(n3105), .Q(g8562) );
  AND2X1 U3146 ( .IN1(g1690), .IN2(g1675), .Q(n3105) );
  AND2X1 U3147 ( .IN1(n1653), .IN2(g1657), .Q(n3104) );
  OR2X1 U3148 ( .IN1(n3106), .IN2(n3107), .Q(g8561) );
  AND2X1 U3149 ( .IN1(g1690), .IN2(g1672), .Q(n3107) );
  AND2X1 U3150 ( .IN1(n1653), .IN2(g1654), .Q(n3106) );
  OR3X1 U3151 ( .IN1(n3108), .IN2(n3109), .IN3(n2912), .Q(g8559) );
  AND2X1 U3152 ( .IN1(n3110), .IN2(g1878), .Q(n3109) );
  AND2X1 U3153 ( .IN1(g18), .IN2(n3111), .Q(g8505) );
  XOR2X1 U3154 ( .IN1(g617), .IN2(n3112), .Q(n3111) );
  OR2X1 U3155 ( .IN1(n2959), .IN2(n3071), .Q(n3112) );
  AND2X1 U3156 ( .IN1(g736), .IN2(n3113), .Q(n3071) );
  AND2X1 U3157 ( .IN1(n2961), .IN2(n3095), .Q(n2959) );
  AND4X1 U3158 ( .IN1(n2957), .IN2(n1609), .IN3(n1593), .IN4(n1645), .Q(n3095)
         );
  AND2X1 U3159 ( .IN1(g591), .IN2(n1644), .Q(n2957) );
  OR2X1 U3160 ( .IN1(n3114), .IN2(n3115), .Q(g8435) );
  AND2X1 U3161 ( .IN1(n3113), .IN2(g727), .Q(n3115) );
  AND2X1 U3162 ( .IN1(n3116), .IN2(g736), .Q(n3114) );
  OR2X1 U3163 ( .IN1(n3117), .IN2(n3118), .Q(g8434) );
  AND2X1 U3164 ( .IN1(n3113), .IN2(g718), .Q(n3118) );
  AND2X1 U3165 ( .IN1(n3116), .IN2(g727), .Q(n3117) );
  OR2X1 U3166 ( .IN1(n3119), .IN2(n3120), .Q(g8433) );
  AND2X1 U3167 ( .IN1(n3113), .IN2(g709), .Q(n3120) );
  AND2X1 U3168 ( .IN1(n3116), .IN2(g718), .Q(n3119) );
  OR2X1 U3169 ( .IN1(n3121), .IN2(n3122), .Q(g8432) );
  AND2X1 U3170 ( .IN1(n3113), .IN2(g700), .Q(n3122) );
  AND2X1 U3172 ( .IN1(n3116), .IN2(g709), .Q(n3121) );
  OR2X1 U3173 ( .IN1(n3123), .IN2(n3124), .Q(g8431) );
  AND2X1 U3174 ( .IN1(n3113), .IN2(g691), .Q(n3124) );
  AND2X1 U3175 ( .IN1(n3116), .IN2(g700), .Q(n3123) );
  OR2X1 U3176 ( .IN1(n3125), .IN2(n3126), .Q(g8430) );
  AND2X1 U3177 ( .IN1(n3113), .IN2(g682), .Q(n3126) );
  AND2X1 U3178 ( .IN1(n3116), .IN2(g691), .Q(n3125) );
  OR2X1 U3179 ( .IN1(n3127), .IN2(n3128), .Q(g8429) );
  AND2X1 U3180 ( .IN1(n3113), .IN2(g673), .Q(n3128) );
  AND2X1 U3181 ( .IN1(n3116), .IN2(g682), .Q(n3127) );
  OR2X1 U3182 ( .IN1(n3129), .IN2(n3130), .Q(g8428) );
  AND2X1 U3183 ( .IN1(n3113), .IN2(g664), .Q(n3130) );
  AND2X1 U3184 ( .IN1(n3116), .IN2(g673), .Q(n3129) );
  AND2X1 U3185 ( .IN1(n2965), .IN2(n124), .Q(n3116) );
  INVX0 U3186 ( .INP(n3113), .ZN(n124) );
  AND3X1 U3187 ( .IN1(g617), .IN2(n2961), .IN3(n1609), .Q(n3113) );
  AND2X1 U3188 ( .IN1(g18), .IN2(n3131), .Q(g8384) );
  XOR2X1 U3189 ( .IN1(g1840), .IN2(n3132), .Q(n3131) );
  OR2X1 U3190 ( .IN1(n3108), .IN2(n257), .Q(n3132) );
  INVX0 U3191 ( .INP(n3133), .ZN(n257) );
  OR2X1 U3192 ( .IN1(n493), .IN2(n3134), .Q(n3133) );
  INVX0 U3193 ( .INP(n926), .ZN(n493) );
  AND2X1 U3194 ( .IN1(n3135), .IN2(g1950), .Q(n3108) );
  OR2X1 U3195 ( .IN1(g82), .IN2(g8986), .Q(g8352) );
  OR2X1 U3196 ( .IN1(g82), .IN2(g8985), .Q(g8349) );
  OR2X1 U3197 ( .IN1(g82), .IN2(g8976), .Q(g8347) );
  OR2X1 U3198 ( .IN1(g82), .IN2(test_so10), .Q(g8340) );
  OR2X1 U3199 ( .IN1(g82), .IN2(g8983), .Q(g8335) );
  OR2X1 U3200 ( .IN1(g82), .IN2(g8982), .Q(g8331) );
  OR2X1 U3201 ( .IN1(g82), .IN2(g8981), .Q(g8328) );
  OR2X1 U3202 ( .IN1(g82), .IN2(g8980), .Q(g8323) );
  OR2X1 U3203 ( .IN1(g82), .IN2(g8979), .Q(g8318) );
  OR2X1 U3204 ( .IN1(g82), .IN2(g8978), .Q(g8316) );
  OR2X1 U3205 ( .IN1(g82), .IN2(g8977), .Q(g8313) );
  OR2X1 U3206 ( .IN1(n3136), .IN2(n3137), .Q(g8288) );
  AND2X1 U3207 ( .IN1(n3135), .IN2(g1941), .Q(n3137) );
  AND2X1 U3208 ( .IN1(n3138), .IN2(g1950), .Q(n3136) );
  OR2X1 U3209 ( .IN1(n3139), .IN2(n3140), .Q(g8287) );
  AND2X1 U3210 ( .IN1(n3135), .IN2(g1932), .Q(n3140) );
  AND2X1 U3211 ( .IN1(n3138), .IN2(g1941), .Q(n3139) );
  OR2X1 U3212 ( .IN1(n3141), .IN2(n3142), .Q(g8286) );
  AND2X1 U3213 ( .IN1(n3135), .IN2(g1923), .Q(n3142) );
  AND2X1 U3214 ( .IN1(n3138), .IN2(g1932), .Q(n3141) );
  OR2X1 U3215 ( .IN1(n3143), .IN2(n3144), .Q(g8285) );
  AND2X1 U3216 ( .IN1(n3135), .IN2(g1914), .Q(n3144) );
  AND2X1 U3217 ( .IN1(n3138), .IN2(g1923), .Q(n3143) );
  OR2X1 U3218 ( .IN1(n3145), .IN2(n3146), .Q(g8284) );
  AND2X1 U3219 ( .IN1(n3135), .IN2(g1905), .Q(n3146) );
  AND2X1 U3220 ( .IN1(n3138), .IN2(g1914), .Q(n3145) );
  OR2X1 U3221 ( .IN1(n3147), .IN2(n3148), .Q(g8283) );
  AND2X1 U3222 ( .IN1(n3135), .IN2(g1896), .Q(n3148) );
  AND2X1 U3223 ( .IN1(n3138), .IN2(g1905), .Q(n3147) );
  OR2X1 U3224 ( .IN1(n3149), .IN2(n3150), .Q(g8282) );
  AND2X1 U3225 ( .IN1(n3135), .IN2(g1887), .Q(n3150) );
  AND2X1 U3226 ( .IN1(n3138), .IN2(g1896), .Q(n3149) );
  OR2X1 U3227 ( .IN1(n3151), .IN2(n3152), .Q(g8281) );
  AND2X1 U3228 ( .IN1(n3135), .IN2(g1878), .Q(n3152) );
  AND2X1 U3229 ( .IN1(n3138), .IN2(g1887), .Q(n3151) );
  AND2X1 U3230 ( .IN1(n2764), .IN2(n3110), .Q(n3138) );
  INVX0 U3231 ( .INP(n3135), .ZN(n3110) );
  AND3X1 U3232 ( .IN1(g1840), .IN2(n926), .IN3(n1655), .Q(n3135) );
  AND2X1 U3233 ( .IN1(n3153), .IN2(g940), .Q(g8260) );
  AND2X1 U3234 ( .IN1(n3153), .IN2(g936), .Q(g8254) );
  AND2X1 U3235 ( .IN1(n3153), .IN2(g932), .Q(g8250) );
  AND2X1 U3236 ( .IN1(n3154), .IN2(n3155), .Q(g8245) );
  XOR2X1 U3237 ( .IN1(n3156), .IN2(n1716), .Q(n3154) );
  OR2X1 U3238 ( .IN1(n2428), .IN2(n3157), .Q(n3156) );
  AND3X1 U3239 ( .IN1(n3158), .IN2(n3159), .IN3(n2745), .Q(g8244) );
  INVX0 U3240 ( .INP(n3160), .ZN(n3158) );
  AND2X1 U3241 ( .IN1(n3161), .IN2(n2441), .Q(n3160) );
  OR2X1 U3242 ( .IN1(n2743), .IN2(n2466), .Q(n3161) );
  OR2X1 U3243 ( .IN1(n3162), .IN2(n3163), .Q(g8194) );
  AND2X1 U3244 ( .IN1(n3164), .IN2(n2971), .Q(n3163) );
  XNOR2X1 U3245 ( .IN1(n4316), .IN2(n3165), .Q(n3164) );
  AND3X1 U3246 ( .IN1(g1104), .IN2(g1110), .IN3(n3166), .Q(n3165) );
  AND2X1 U3247 ( .IN1(n371), .IN2(g1512), .Q(n3162) );
  OR2X1 U3248 ( .IN1(n3167), .IN2(n3168), .Q(g8193) );
  AND2X1 U3249 ( .IN1(n3169), .IN2(n2971), .Q(n3168) );
  XOR2X1 U3250 ( .IN1(test_so4), .IN2(n3170), .Q(n3169) );
  AND2X1 U3251 ( .IN1(n3166), .IN2(n2987), .Q(n3170) );
  AND2X1 U3252 ( .IN1(g1104), .IN2(n1677), .Q(n2987) );
  AND2X1 U3253 ( .IN1(n1614), .IN2(n1654), .Q(n3166) );
  AND2X1 U3254 ( .IN1(n371), .IN2(g1639), .Q(n3167) );
  AND2X1 U3255 ( .IN1(n1610), .IN2(n3171), .Q(g8173) );
  OR2X1 U3256 ( .IN1(n3172), .IN2(n3173), .Q(n3171) );
  AND2X1 U3257 ( .IN1(n3174), .IN2(g1806), .Q(n3173) );
  OR2X1 U3258 ( .IN1(n369), .IN2(n1055), .Q(n3174) );
  AND3X1 U3259 ( .IN1(n1055), .IN2(g1801), .IN3(n1056), .Q(n3172) );
  OR3X1 U3260 ( .IN1(n2427), .IN2(n2426), .IN3(n2734), .Q(n1055) );
  OR2X1 U3261 ( .IN1(n1626), .IN2(n3175), .Q(n2734) );
  AND2X1 U3262 ( .IN1(n3153), .IN2(g928), .Q(g8147) );
  INVX0 U3263 ( .INP(n3176), .ZN(n3153) );
  OR2X1 U3264 ( .IN1(n505), .IN2(n3177), .Q(n3176) );
  AND3X1 U3265 ( .IN1(n3178), .IN2(DFF_436_n1), .IN3(n3179), .Q(n3177) );
  AND2X1 U3266 ( .IN1(n3180), .IN2(g109), .Q(g8060) );
  XNOR2X1 U3267 ( .IN1(n2347), .IN2(g6002), .Q(n3180) );
  AND2X1 U3268 ( .IN1(n3181), .IN2(g109), .Q(g8059) );
  XNOR2X1 U3269 ( .IN1(n2345), .IN2(g6042), .Q(n3181) );
  AND2X1 U3270 ( .IN1(n3182), .IN2(g109), .Q(g8055) );
  XNOR2X1 U3271 ( .IN1(n2399), .IN2(n3183), .Q(n3182) );
  AND2X1 U3272 ( .IN1(n3184), .IN2(g109), .Q(g8054) );
  XOR2X1 U3273 ( .IN1(g174), .IN2(g6015), .Q(n3184) );
  AND2X1 U3274 ( .IN1(n3185), .IN2(g109), .Q(g8053) );
  XNOR2X1 U3275 ( .IN1(n2344), .IN2(g6045), .Q(n3185) );
  AND2X1 U3276 ( .IN1(n3186), .IN2(g109), .Q(g8052) );
  XOR2X1 U3277 ( .IN1(g1486), .IN2(n3187), .Q(n3186) );
  AND2X1 U3278 ( .IN1(n3188), .IN2(g109), .Q(g8051) );
  XOR2X1 U3279 ( .IN1(g1466), .IN2(n3189), .Q(n3188) );
  AND2X1 U3280 ( .IN1(n3190), .IN2(g109), .Q(g8050) );
  XOR2X1 U3281 ( .IN1(g170), .IN2(g6026), .Q(n3190) );
  AND2X1 U3282 ( .IN1(n3191), .IN2(g109), .Q(g8049) );
  XOR2X1 U3283 ( .IN1(g166), .IN2(g6049), .Q(n3191) );
  AND2X1 U3284 ( .IN1(n3192), .IN2(g109), .Q(g8048) );
  XNOR2X1 U3285 ( .IN1(n2362), .IN2(g5996), .Q(n3192) );
  AND2X1 U3286 ( .IN1(n3193), .IN2(g109), .Q(g8047) );
  XNOR2X1 U3287 ( .IN1(n1704), .IN2(g6035), .Q(n3193) );
  AND2X1 U3288 ( .IN1(n3194), .IN2(g109), .Q(g8046) );
  XOR2X1 U3289 ( .IN1(g1482), .IN2(n3195), .Q(n3194) );
  AND2X1 U3290 ( .IN1(n3196), .IN2(g109), .Q(g8045) );
  XNOR2X1 U3291 ( .IN1(n2400), .IN2(n3197), .Q(n3196) );
  AND2X1 U3292 ( .IN1(n3198), .IN2(g109), .Q(g8044) );
  XNOR2X1 U3293 ( .IN1(n2343), .IN2(g6038), .Q(n3198) );
  AND2X1 U3294 ( .IN1(n3199), .IN2(g109), .Q(g8043) );
  XNOR2X1 U3295 ( .IN1(n2401), .IN2(n3200), .Q(n3199) );
  AND2X1 U3296 ( .IN1(n3201), .IN2(g109), .Q(g8042) );
  XOR2X1 U3297 ( .IN1(g1458), .IN2(n3202), .Q(n3201) );
  AND2X1 U3298 ( .IN1(n3203), .IN2(g109), .Q(g8041) );
  XNOR2X1 U3299 ( .IN1(n2411), .IN2(n3204), .Q(n3203) );
  AND2X1 U3300 ( .IN1(n3205), .IN2(g109), .Q(g8040) );
  XNOR2X1 U3301 ( .IN1(n2412), .IN2(n3206), .Q(n3205) );
  AND2X1 U3302 ( .IN1(n3207), .IN2(g109), .Q(g8039) );
  XNOR2X1 U3303 ( .IN1(n2413), .IN2(n3208), .Q(n3207) );
  AND2X1 U3304 ( .IN1(n3209), .IN2(n3155), .Q(g8024) );
  XOR2X1 U3305 ( .IN1(n3157), .IN2(n2428), .Q(n3209) );
  AND2X1 U3306 ( .IN1(n3210), .IN2(n2745), .Q(g8019) );
  XOR2X1 U3307 ( .IN1(n2466), .IN2(n2743), .Q(n3210) );
  AND2X1 U3308 ( .IN1(n3211), .IN2(n1610), .Q(g7930) );
  XOR2X1 U3309 ( .IN1(n1056), .IN2(g1801), .Q(n3211) );
  AND2X1 U3310 ( .IN1(n3212), .IN2(g109), .Q(g7843) );
  XNOR2X1 U3311 ( .IN1(n2348), .IN2(g6000), .Q(n3212) );
  AND3X1 U3312 ( .IN1(n3157), .IN2(n3213), .IN3(n3155), .Q(g7709) );
  INVX0 U3313 ( .INP(n1096), .ZN(n3213) );
  INVX0 U3314 ( .INP(n1090), .ZN(n3157) );
  AND3X1 U3315 ( .IN1(n3214), .IN2(n3215), .IN3(n3216), .Q(g7632) );
  INVX0 U3316 ( .INP(n3217), .ZN(n3215) );
  OR2X1 U3317 ( .IN1(n3218), .IN2(g1218), .Q(n3214) );
  OR3X1 U3318 ( .IN1(n3219), .IN2(n3220), .IN3(n2784), .Q(g7626) );
  AND3X1 U3319 ( .IN1(n2961), .IN2(n3221), .IN3(n1692), .Q(n3220) );
  OR3X1 U3320 ( .IN1(n2958), .IN2(n2791), .IN3(n2706), .Q(n3221) );
  OR2X1 U3321 ( .IN1(n2788), .IN2(n3222), .Q(n2706) );
  INVX0 U3322 ( .INP(n3092), .ZN(n3222) );
  OR2X1 U3323 ( .IN1(n1644), .IN2(g605), .Q(n3092) );
  AND3X1 U3324 ( .IN1(g605), .IN2(n1607), .IN3(n1644), .Q(n2788) );
  INVX0 U3325 ( .INP(n2799), .ZN(n2791) );
  OR2X1 U3326 ( .IN1(n1593), .IN2(n1607), .Q(n2799) );
  INVX0 U3327 ( .INP(n2797), .ZN(n2958) );
  OR2X1 U3328 ( .IN1(n1644), .IN2(g591), .Q(n2797) );
  AND2X1 U3329 ( .IN1(n2752), .IN2(g639), .Q(n3219) );
  AND2X1 U3330 ( .IN1(n3216), .IN2(n3223), .Q(g7590) );
  INVX0 U3331 ( .INP(n3224), .ZN(n3223) );
  AND2X1 U3332 ( .IN1(n3225), .IN2(n2462), .Q(n3224) );
  AND2X1 U3333 ( .IN1(n3216), .IN2(n3226), .Q(g7586) );
  OR2X1 U3334 ( .IN1(n3227), .IN2(n1107), .Q(n3226) );
  AND3X1 U3335 ( .IN1(g1223), .IN2(n3228), .IN3(n3217), .Q(n1107) );
  AND2X1 U3336 ( .IN1(n3225), .IN2(g1227), .Q(n3227) );
  OR3X1 U3337 ( .IN1(n3229), .IN2(n3228), .IN3(n3230), .Q(n3225) );
  AND2X1 U3338 ( .IN1(n3231), .IN2(n3216), .Q(g7581) );
  XNOR2X1 U3339 ( .IN1(n3217), .IN2(n2449), .Q(n3231) );
  AND3X1 U3340 ( .IN1(g1218), .IN2(n3232), .IN3(n3218), .Q(n3217) );
  AND3X1 U3341 ( .IN1(n3233), .IN2(n3234), .IN3(n1610), .Q(g7541) );
  OR2X1 U3342 ( .IN1(n1626), .IN2(n3235), .Q(n3234) );
  INVX0 U3343 ( .INP(n1056), .ZN(n3235) );
  OR2X1 U3344 ( .IN1(n113), .IN2(g1796), .Q(n3233) );
  INVX0 U3345 ( .INP(n3236), .ZN(n113) );
  OR2X1 U3346 ( .IN1(n3237), .IN2(n3238), .Q(g7303) );
  AND2X1 U3347 ( .IN1(n3218), .IN2(g1265), .Q(n3238) );
  AND2X1 U3348 ( .IN1(n3239), .IN2(test_so6), .Q(n3237) );
  OR2X1 U3349 ( .IN1(n3240), .IN2(n3241), .Q(g7302) );
  AND2X1 U3350 ( .IN1(n3218), .IN2(g1260), .Q(n3241) );
  AND2X1 U3351 ( .IN1(n3239), .IN2(g1265), .Q(n3240) );
  OR2X1 U3352 ( .IN1(n3242), .IN2(n3243), .Q(g7301) );
  AND2X1 U3353 ( .IN1(n3218), .IN2(g1255), .Q(n3243) );
  AND2X1 U3354 ( .IN1(n3239), .IN2(g1260), .Q(n3242) );
  OR2X1 U3355 ( .IN1(n3244), .IN2(n3245), .Q(g7300) );
  AND2X1 U3356 ( .IN1(n3218), .IN2(g1250), .Q(n3245) );
  AND2X1 U3357 ( .IN1(n3239), .IN2(g1255), .Q(n3244) );
  OR2X1 U3358 ( .IN1(n3246), .IN2(n3247), .Q(g7299) );
  AND2X1 U3359 ( .IN1(n3218), .IN2(g1245), .Q(n3247) );
  AND2X1 U3360 ( .IN1(n3239), .IN2(g1250), .Q(n3246) );
  OR2X1 U3361 ( .IN1(n3248), .IN2(n3249), .Q(g7298) );
  AND2X1 U3362 ( .IN1(n3218), .IN2(g1240), .Q(n3249) );
  AND2X1 U3363 ( .IN1(n3239), .IN2(g1245), .Q(n3248) );
  OR2X1 U3364 ( .IN1(n3250), .IN2(n3251), .Q(g7297) );
  AND2X1 U3365 ( .IN1(n3218), .IN2(g1235), .Q(n3251) );
  AND2X1 U3366 ( .IN1(n3239), .IN2(g1240), .Q(n3250) );
  OR2X1 U3367 ( .IN1(n3252), .IN2(n3253), .Q(g7296) );
  AND2X1 U3368 ( .IN1(n3218), .IN2(g1275), .Q(n3253) );
  AND2X1 U3369 ( .IN1(n3239), .IN2(g1235), .Q(n3252) );
  OR2X1 U3370 ( .IN1(n3254), .IN2(n3255), .Q(g7295) );
  AND2X1 U3371 ( .IN1(n3218), .IN2(g1284), .Q(n3255) );
  AND2X1 U3372 ( .IN1(n3239), .IN2(g1280), .Q(n3254) );
  OR2X1 U3373 ( .IN1(n3256), .IN2(n3257), .Q(g7294) );
  AND2X1 U3374 ( .IN1(n3218), .IN2(g1292), .Q(n3257) );
  AND2X1 U3375 ( .IN1(n3239), .IN2(g1284), .Q(n3256) );
  OR2X1 U3376 ( .IN1(n3258), .IN2(n3259), .Q(g7293) );
  AND2X1 U3377 ( .IN1(n3218), .IN2(g1296), .Q(n3259) );
  AND2X1 U3378 ( .IN1(n3239), .IN2(g1292), .Q(n3258) );
  OR2X1 U3379 ( .IN1(n3260), .IN2(n3261), .Q(g7292) );
  AND2X1 U3380 ( .IN1(n3218), .IN2(g1300), .Q(n3261) );
  AND2X1 U3381 ( .IN1(n3239), .IN2(g1296), .Q(n3260) );
  OR2X1 U3382 ( .IN1(n3262), .IN2(n3263), .Q(g7291) );
  AND2X1 U3383 ( .IN1(n3218), .IN2(g1304), .Q(n3263) );
  AND2X1 U3384 ( .IN1(n3239), .IN2(g1300), .Q(n3262) );
  OR2X1 U3385 ( .IN1(n3264), .IN2(n3265), .Q(g7290) );
  AND2X1 U3386 ( .IN1(n3218), .IN2(test_so6), .Q(n3265) );
  AND2X1 U3387 ( .IN1(n3239), .IN2(g1304), .Q(n3264) );
  OR2X1 U3388 ( .IN1(n3266), .IN2(n3267), .Q(g7257) );
  AND2X1 U3389 ( .IN1(n371), .IN2(g1032), .Q(n3267) );
  AND2X1 U3390 ( .IN1(n2971), .IN2(g1077), .Q(n3266) );
  OR2X1 U3391 ( .IN1(n3268), .IN2(n3269), .Q(g7244) );
  AND2X1 U3392 ( .IN1(n371), .IN2(g1023), .Q(n3269) );
  AND2X1 U3393 ( .IN1(n2971), .IN2(g1071), .Q(n3268) );
  OR2X1 U3394 ( .IN1(n3270), .IN2(test_so10), .Q(g7219) );
  OR2X1 U3395 ( .IN1(n3270), .IN2(g8982), .Q(g7204) );
  AND2X1 U3396 ( .IN1(n3271), .IN2(n3155), .Q(g7202) );
  XOR2X1 U3397 ( .IN1(n2742), .IN2(n2431), .Q(n3271) );
  AND2X1 U3398 ( .IN1(n3272), .IN2(n2745), .Q(g7191) );
  XOR2X1 U3399 ( .IN1(n2741), .IN2(n2446), .Q(n3272) );
  OR2X1 U3400 ( .IN1(n3270), .IN2(g8980), .Q(g7189) );
  OR2X1 U3401 ( .IN1(n3270), .IN2(g8978), .Q(g7183) );
  OR2X1 U3402 ( .IN1(n3270), .IN2(g8976), .Q(g7143) );
  AND2X1 U3403 ( .IN1(n3273), .IN2(n2726), .Q(g7137) );
  XNOR2X1 U3404 ( .IN1(n2728), .IN2(n1709), .Q(n3273) );
  AND2X1 U3405 ( .IN1(n2726), .IN2(n3274), .Q(g7134) );
  OR2X1 U3406 ( .IN1(n3275), .IN2(n2728), .Q(n3274) );
  AND2X1 U3407 ( .IN1(n2730), .IN2(n3062), .Q(n3275) );
  INVX0 U3408 ( .INP(n3276), .ZN(n2730) );
  AND2X1 U3409 ( .IN1(n2965), .IN2(n2752), .Q(n2726) );
  INVX0 U3410 ( .INP(n2961), .ZN(n2752) );
  AND3X1 U3411 ( .IN1(n2728), .IN2(n1709), .IN3(n2450), .Q(n2961) );
  AND2X1 U3412 ( .IN1(n3276), .IN2(n4311), .Q(n2728) );
  AND2X1 U3413 ( .IN1(g627), .IN2(n1612), .Q(n3276) );
  OR2X1 U3414 ( .IN1(n3277), .IN2(g1713), .Q(g7133) );
  AND2X1 U3415 ( .IN1(n3278), .IN2(n3279), .Q(n3277) );
  OR2X1 U3416 ( .IN1(n2500), .IN2(g1766), .Q(n3278) );
  OR2X1 U3417 ( .IN1(n3280), .IN2(n1132), .Q(g7032) );
  AND4X1 U3418 ( .IN1(n3281), .IN2(n3282), .IN3(n3283), .IN4(n3284), .Q(n1132)
         );
  AND4X1 U3419 ( .IN1(g174), .IN2(g170), .IN3(g166), .IN4(g182), .Q(n3284) );
  AND4X1 U3420 ( .IN1(n1704), .IN2(n1613), .IN3(g6786), .IN4(n1137), .Q(n3283)
         );
  AND4X1 U3421 ( .IN1(n2347), .IN2(n2345), .IN3(n2344), .IN4(n2343), .Q(n3282)
         );
  AND4X1 U3422 ( .IN1(n2364), .IN2(n2363), .IN3(n2362), .IN4(n2348), .Q(n3281)
         );
  AND2X1 U3423 ( .IN1(g109), .IN2(g123), .Q(n3280) );
  AND2X1 U3424 ( .IN1(n1610), .IN2(n3285), .Q(g6983) );
  OR2X1 U3425 ( .IN1(n3286), .IN2(n3287), .Q(n3285) );
  AND2X1 U3426 ( .IN1(n3236), .IN2(g1791), .Q(n3287) );
  OR2X1 U3427 ( .IN1(n369), .IN2(n3175), .Q(n3236) );
  AND3X1 U3428 ( .IN1(n3175), .IN2(g1786), .IN3(n155), .Q(n3286) );
  OR3X1 U3429 ( .IN1(n1659), .IN2(n2736), .IN3(n2740), .Q(n3175) );
  OR2X1 U3430 ( .IN1(n3288), .IN2(n3289), .Q(g6934) );
  AND2X1 U3431 ( .IN1(n3290), .IN2(g170), .Q(n3289) );
  AND2X1 U3432 ( .IN1(n3291), .IN2(g284), .Q(n3288) );
  OR2X1 U3433 ( .IN1(n3292), .IN2(n3293), .Q(g6930) );
  AND2X1 U3434 ( .IN1(n371), .IN2(g1015), .Q(n3293) );
  AND2X1 U3435 ( .IN1(n2971), .IN2(g1074), .Q(n3292) );
  OR2X1 U3436 ( .IN1(n3294), .IN2(n3295), .Q(g6929) );
  AND2X1 U3437 ( .IN1(n3290), .IN2(g143), .Q(n3295) );
  AND2X1 U3438 ( .IN1(n3291), .IN2(g302), .Q(n3294) );
  OR2X1 U3439 ( .IN1(n3296), .IN2(n3297), .Q(g6928) );
  AND2X1 U3440 ( .IN1(n3290), .IN2(g174), .Q(n3297) );
  AND2X1 U3441 ( .IN1(n3291), .IN2(g281), .Q(n3296) );
  OR2X1 U3442 ( .IN1(n3298), .IN2(n3299), .Q(g6924) );
  AND2X1 U3443 ( .IN1(n371), .IN2(g1019), .Q(n3299) );
  AND2X1 U3444 ( .IN1(n2971), .IN2(g1098), .Q(n3298) );
  OR2X1 U3445 ( .IN1(n3300), .IN2(n3301), .Q(g6923) );
  AND2X1 U3446 ( .IN1(n3290), .IN2(g166), .Q(n3301) );
  AND2X1 U3447 ( .IN1(n3291), .IN2(g299), .Q(n3300) );
  OR2X1 U3448 ( .IN1(n3302), .IN2(n3303), .Q(g6922) );
  AND2X1 U3449 ( .IN1(n3290), .IN2(g162), .Q(n3303) );
  AND2X1 U3450 ( .IN1(n3291), .IN2(g278), .Q(n3302) );
  OR2X1 U3451 ( .IN1(n3304), .IN2(n3305), .Q(g6918) );
  AND2X1 U3452 ( .IN1(test_so2), .IN2(n371), .Q(n3305) );
  AND2X1 U3453 ( .IN1(n2971), .IN2(g1095), .Q(n3304) );
  OR2X1 U3454 ( .IN1(n3306), .IN2(n3307), .Q(g6916) );
  AND2X1 U3455 ( .IN1(n3290), .IN2(g139), .Q(n3307) );
  AND2X1 U3456 ( .IN1(n3291), .IN2(g296), .Q(n3306) );
  OR2X1 U3457 ( .IN1(n3308), .IN2(n3309), .Q(g6915) );
  AND2X1 U3458 ( .IN1(n3290), .IN2(g158), .Q(n3309) );
  AND2X1 U3459 ( .IN1(n3291), .IN2(g275), .Q(n3308) );
  OR2X1 U3460 ( .IN1(n3310), .IN2(n3311), .Q(g6912) );
  AND2X1 U3461 ( .IN1(n371), .IN2(g1011), .Q(n3311) );
  AND2X1 U3462 ( .IN1(n2971), .IN2(g1092), .Q(n3310) );
  OR2X1 U3463 ( .IN1(n3312), .IN2(n3313), .Q(g6911) );
  AND2X1 U3464 ( .IN1(n3290), .IN2(g135), .Q(n3313) );
  AND2X1 U3465 ( .IN1(n3291), .IN2(g293), .Q(n3312) );
  OR2X1 U3466 ( .IN1(n3314), .IN2(n3315), .Q(g6910) );
  AND2X1 U3467 ( .IN1(n3290), .IN2(g153), .Q(n3315) );
  AND2X1 U3468 ( .IN1(n3291), .IN2(g272), .Q(n3314) );
  OR2X1 U3469 ( .IN1(n3316), .IN2(n2694), .Q(g6909) );
  AND2X1 U3470 ( .IN1(n2697), .IN2(g1868), .Q(n3316) );
  INVX0 U3471 ( .INP(n1147), .ZN(n2697) );
  AND3X1 U3472 ( .IN1(n3033), .IN2(n2417), .IN3(n2416), .Q(n1147) );
  OR2X1 U3473 ( .IN1(n3317), .IN2(n3318), .Q(g6908) );
  AND2X1 U3474 ( .IN1(test_so8), .IN2(n371), .Q(n3318) );
  AND2X1 U3475 ( .IN1(n2971), .IN2(g1089), .Q(n3317) );
  OR2X1 U3476 ( .IN1(n3319), .IN2(n3320), .Q(g6907) );
  AND2X1 U3477 ( .IN1(n3290), .IN2(g131), .Q(n3320) );
  AND2X1 U3478 ( .IN1(n3291), .IN2(g290), .Q(n3319) );
  OR2X1 U3479 ( .IN1(n3321), .IN2(n3322), .Q(g6906) );
  AND2X1 U3480 ( .IN1(n3290), .IN2(g148), .Q(n3322) );
  AND2X1 U3481 ( .IN1(n3291), .IN2(g269), .Q(n3321) );
  OR2X1 U3482 ( .IN1(n3323), .IN2(n3324), .Q(g6902) );
  AND2X1 U3483 ( .IN1(n371), .IN2(g1003), .Q(n3324) );
  AND2X1 U3484 ( .IN1(n2971), .IN2(g1086), .Q(n3323) );
  OR2X1 U3485 ( .IN1(n3325), .IN2(n3326), .Q(g6901) );
  AND2X1 U3486 ( .IN1(n3290), .IN2(g127), .Q(n3326) );
  AND2X1 U3487 ( .IN1(n3291), .IN2(g287), .Q(n3325) );
  OR2X1 U3488 ( .IN1(n3327), .IN2(n3328), .Q(g6900) );
  AND2X1 U3489 ( .IN1(n3290), .IN2(g178), .Q(n3328) );
  AND2X1 U3490 ( .IN1(n3291), .IN2(g266), .Q(n3327) );
  OR2X1 U3491 ( .IN1(n3329), .IN2(n3330), .Q(g6898) );
  AND2X1 U3492 ( .IN1(n371), .IN2(g991), .Q(n3330) );
  AND2X1 U3493 ( .IN1(n2971), .IN2(g1083), .Q(n3329) );
  OR2X1 U3494 ( .IN1(n3331), .IN2(n3332), .Q(g6897) );
  AND2X1 U3495 ( .IN1(n3290), .IN2(g182), .Q(n3332) );
  AND2X1 U3496 ( .IN1(n3291), .IN2(g263), .Q(n3331) );
  INVX0 U3497 ( .INP(n3290), .ZN(n3291) );
  OR2X1 U3498 ( .IN1(n505), .IN2(n3333), .Q(n3290) );
  AND2X1 U3499 ( .IN1(n1613), .IN2(n1137), .Q(n3333) );
  INVX0 U3500 ( .INP(n3334), .ZN(n1137) );
  OR2X1 U3501 ( .IN1(n4312), .IN2(n2985), .Q(n3334) );
  OR2X1 U3502 ( .IN1(n3335), .IN2(n3336), .Q(g6895) );
  AND2X1 U3503 ( .IN1(n371), .IN2(g995), .Q(n3336) );
  AND2X1 U3504 ( .IN1(n2971), .IN2(g1080), .Q(n3335) );
  OR2X1 U3505 ( .IN1(n3337), .IN2(n3338), .Q(g6894) );
  AND2X1 U3506 ( .IN1(n371), .IN2(g1027), .Q(n3338) );
  AND2X1 U3507 ( .IN1(test_so7), .IN2(n2971), .Q(n3337) );
  AND2X1 U3508 ( .IN1(n3339), .IN2(n3340), .Q(g6842) );
  AND2X1 U3509 ( .IN1(g109), .IN2(g1400), .Q(g6841) );
  AND2X1 U3510 ( .IN1(g109), .IN2(g248), .Q(g6840) );
  AND2X1 U3511 ( .IN1(g109), .IN2(g1397), .Q(g6839) );
  AND2X1 U3512 ( .IN1(g109), .IN2(n3054), .Q(g6834) );
  AND2X1 U3513 ( .IN1(g109), .IN2(n3019), .Q(g6830) );
  AND2X1 U3514 ( .IN1(g109), .IN2(n3038), .Q(g6828) );
  AND2X1 U3515 ( .IN1(g109), .IN2(n3061), .Q(g6820) );
  OR2X1 U3516 ( .IN1(n2499), .IN2(n3033), .Q(g6755) );
  AND3X1 U3517 ( .IN1(n3341), .IN2(g109), .IN3(n4312), .Q(g6747) );
  OR2X1 U3518 ( .IN1(n3041), .IN2(n3024), .Q(n3341) );
  AND3X1 U3519 ( .IN1(n2742), .IN2(n3342), .IN3(n3155), .Q(g6733) );
  INVX0 U3520 ( .INP(n1150), .ZN(n3342) );
  INVX0 U3521 ( .INP(n1123), .ZN(n2742) );
  AND3X1 U3522 ( .IN1(n2741), .IN2(n3343), .IN3(n2745), .Q(g6728) );
  INVX0 U3523 ( .INP(n1152), .ZN(n3343) );
  INVX0 U3524 ( .INP(n1125), .ZN(n2741) );
  OR2X1 U3525 ( .IN1(n3344), .IN2(n3345), .Q(g6679) );
  AND2X1 U3526 ( .IN1(g109), .IN2(g1), .Q(n3345) );
  AND2X1 U3527 ( .IN1(n1154), .IN2(n86), .Q(n3344) );
  INVX0 U3528 ( .INP(n3346), .ZN(n86) );
  OR2X1 U3529 ( .IN1(n3347), .IN2(n3348), .Q(n3346) );
  OR4X1 U3530 ( .IN1(g1411), .IN2(g1403), .IN3(g1415), .IN4(g1407), .Q(n3348)
         );
  OR4X1 U3531 ( .IN1(n2403), .IN2(n2402), .IN3(n2405), .IN4(n2404), .Q(n3347)
         );
  AND4X1 U3532 ( .IN1(g1419), .IN2(n1159), .IN3(g6234), .IN4(n3349), .Q(n1154)
         );
  AND4X1 U3533 ( .IN1(g1520), .IN2(g1515), .IN3(g1432), .IN4(g1448), .Q(n3349)
         );
  OR2X1 U3534 ( .IN1(n2497), .IN2(g627), .Q(g6672) );
  OR2X1 U3535 ( .IN1(n3350), .IN2(n3351), .Q(g6656) );
  AND2X1 U3536 ( .IN1(g109), .IN2(g4), .Q(n3351) );
  AND2X1 U3537 ( .IN1(n1161), .IN2(n84), .Q(n3350) );
  INVX0 U3538 ( .INP(n3352), .ZN(n84) );
  OR2X1 U3539 ( .IN1(n3353), .IN2(n3354), .Q(n3352) );
  OR4X1 U3540 ( .IN1(g1482), .IN2(g1499), .IN3(g1486), .IN4(g1466), .Q(n3354)
         );
  OR4X1 U3541 ( .IN1(n2399), .IN2(g1458), .IN3(n2401), .IN4(n2400), .Q(n3353)
         );
  AND4X1 U3542 ( .IN1(g1453), .IN2(n2496), .IN3(n1159), .IN4(n3355), .Q(n1161)
         );
  AND4X1 U3543 ( .IN1(g1494), .IN2(g1508), .IN3(g1470), .IN4(g1474), .Q(n3355)
         );
  AND2X1 U3544 ( .IN1(g1504), .IN2(g109), .Q(n2496) );
  AND2X1 U3545 ( .IN1(n2710), .IN2(g8983), .Q(g6653) );
  AND2X1 U3546 ( .IN1(n2710), .IN2(g8981), .Q(g6638) );
  AND2X1 U3547 ( .IN1(n2710), .IN2(g8979), .Q(g6627) );
  AND2X1 U3548 ( .IN1(n2710), .IN2(g8977), .Q(g6621) );
  OR2X1 U3549 ( .IN1(n3356), .IN2(n3357), .Q(g6551) );
  AND2X1 U3550 ( .IN1(n3358), .IN2(g1478), .Q(n3357) );
  AND2X1 U3551 ( .IN1(n3359), .IN2(g1546), .Q(n3356) );
  OR2X1 U3552 ( .IN1(n3360), .IN2(n3361), .Q(g6546) );
  AND2X1 U3553 ( .IN1(n3358), .IN2(g1453), .Q(n3361) );
  AND2X1 U3554 ( .IN1(n3359), .IN2(g1564), .Q(n3360) );
  OR2X1 U3555 ( .IN1(n3362), .IN2(n3363), .Q(g6545) );
  AND2X1 U3556 ( .IN1(n3358), .IN2(g1482), .Q(n3363) );
  AND2X1 U3557 ( .IN1(n3359), .IN2(g1543), .Q(n3362) );
  OR2X1 U3558 ( .IN1(n3364), .IN2(n3365), .Q(g6542) );
  AND2X1 U3559 ( .IN1(n3358), .IN2(g1458), .Q(n3365) );
  AND2X1 U3560 ( .IN1(n3359), .IN2(g1561), .Q(n3364) );
  OR2X1 U3561 ( .IN1(n3366), .IN2(n3367), .Q(g6541) );
  AND2X1 U3562 ( .IN1(n3358), .IN2(g1486), .Q(n3367) );
  AND2X1 U3563 ( .IN1(n3359), .IN2(g1540), .Q(n3366) );
  OR2X1 U3564 ( .IN1(n3368), .IN2(n3369), .Q(g6538) );
  AND2X1 U3565 ( .IN1(n3358), .IN2(g1462), .Q(n3369) );
  AND2X1 U3566 ( .IN1(n3359), .IN2(g1558), .Q(n3368) );
  OR2X1 U3567 ( .IN1(n3370), .IN2(n3371), .Q(g6537) );
  AND2X1 U3568 ( .IN1(n3358), .IN2(g1490), .Q(n3371) );
  AND2X1 U3569 ( .IN1(n3359), .IN2(g1537), .Q(n3370) );
  OR2X1 U3570 ( .IN1(n3372), .IN2(n3373), .Q(g6534) );
  AND2X1 U3571 ( .IN1(n3358), .IN2(g1466), .Q(n3373) );
  AND2X1 U3572 ( .IN1(n3359), .IN2(g1555), .Q(n3372) );
  OR2X1 U3573 ( .IN1(n3374), .IN2(n3375), .Q(g6533) );
  AND2X1 U3574 ( .IN1(n3358), .IN2(g1494), .Q(n3375) );
  AND2X1 U3575 ( .IN1(n3359), .IN2(g1534), .Q(n3374) );
  AND2X1 U3576 ( .IN1(n2710), .IN2(g8986), .Q(g6531) );
  OR2X1 U3577 ( .IN1(n3376), .IN2(n3377), .Q(g6529) );
  AND2X1 U3578 ( .IN1(n3358), .IN2(g1470), .Q(n3377) );
  AND2X1 U3579 ( .IN1(n3359), .IN2(g1552), .Q(n3376) );
  OR2X1 U3580 ( .IN1(n3378), .IN2(n3379), .Q(g6528) );
  AND2X1 U3581 ( .IN1(n3358), .IN2(g1499), .Q(n3379) );
  AND2X1 U3582 ( .IN1(n3359), .IN2(g1531), .Q(n3378) );
  AND2X1 U3583 ( .IN1(n2710), .IN2(g8985), .Q(g6526) );
  AND2X1 U3584 ( .IN1(n3380), .IN2(n1610), .Q(g6525) );
  XOR2X1 U3585 ( .IN1(g1786), .IN2(n155), .Q(n3380) );
  INVX0 U3586 ( .INP(n3381), .ZN(n155) );
  OR2X1 U3587 ( .IN1(n3382), .IN2(n3383), .Q(g6524) );
  AND2X1 U3588 ( .IN1(n3358), .IN2(g1428), .Q(n3383) );
  AND2X1 U3589 ( .IN1(n3359), .IN2(g1589), .Q(n3382) );
  OR2X1 U3590 ( .IN1(n3384), .IN2(n3385), .Q(g6523) );
  AND2X1 U3591 ( .IN1(n3358), .IN2(g1474), .Q(n3385) );
  AND2X1 U3592 ( .IN1(n3359), .IN2(g1549), .Q(n3384) );
  OR2X1 U3593 ( .IN1(n3386), .IN2(n3387), .Q(g6522) );
  AND2X1 U3594 ( .IN1(n3358), .IN2(g1504), .Q(n3387) );
  AND2X1 U3595 ( .IN1(n3359), .IN2(g1528), .Q(n3386) );
  AND3X1 U3596 ( .IN1(n3388), .IN2(n3381), .IN3(n1610), .Q(g6516) );
  OR2X1 U3597 ( .IN1(n1659), .IN2(n3389), .Q(n3381) );
  OR2X1 U3598 ( .IN1(n3390), .IN2(g1781), .Q(n3388) );
  INVX0 U3599 ( .INP(n3389), .ZN(n3390) );
  OR2X1 U3600 ( .IN1(n3391), .IN2(n3392), .Q(g6515) );
  AND2X1 U3601 ( .IN1(n3358), .IN2(g1448), .Q(n3392) );
  AND2X1 U3602 ( .IN1(n3359), .IN2(g1607), .Q(n3391) );
  OR2X1 U3603 ( .IN1(n3393), .IN2(n3394), .Q(g6514) );
  AND2X1 U3604 ( .IN1(n3358), .IN2(g1407), .Q(n3394) );
  AND2X1 U3605 ( .IN1(n3359), .IN2(g1586), .Q(n3393) );
  OR2X1 U3606 ( .IN1(n3395), .IN2(n3396), .Q(g6513) );
  AND2X1 U3607 ( .IN1(n3358), .IN2(g1508), .Q(n3396) );
  AND2X1 U3608 ( .IN1(n3359), .IN2(g1524), .Q(n3395) );
  AND2X1 U3609 ( .IN1(n1610), .IN2(n3397), .Q(g6508) );
  OR2X1 U3610 ( .IN1(n3398), .IN2(n3399), .Q(n3397) );
  AND2X1 U3611 ( .IN1(n3389), .IN2(g1776), .Q(n3399) );
  OR2X1 U3612 ( .IN1(n369), .IN2(n2736), .Q(n3389) );
  AND3X1 U3613 ( .IN1(test_so5), .IN2(n2736), .IN3(n3400), .Q(n3398) );
  OR2X1 U3614 ( .IN1(n1715), .IN2(n3401), .Q(n2736) );
  OR2X1 U3615 ( .IN1(n3402), .IN2(n3403), .Q(g6507) );
  AND2X1 U3616 ( .IN1(n3358), .IN2(g1444), .Q(n3403) );
  AND2X1 U3617 ( .IN1(n3359), .IN2(g1604), .Q(n3402) );
  OR2X1 U3618 ( .IN1(n3404), .IN2(n3405), .Q(g6506) );
  AND2X1 U3619 ( .IN1(n3358), .IN2(g1424), .Q(n3405) );
  AND2X1 U3620 ( .IN1(n3359), .IN2(g1583), .Q(n3404) );
  AND2X1 U3621 ( .IN1(n1610), .IN2(n3406), .Q(g6502) );
  XOR2X1 U3622 ( .IN1(test_so5), .IN2(n3400), .Q(n3406) );
  INVX0 U3623 ( .INP(n3279), .ZN(n3400) );
  OR2X1 U3624 ( .IN1(n2461), .IN2(n369), .Q(n3279) );
  OR2X1 U3625 ( .IN1(n3407), .IN2(n3408), .Q(g6501) );
  AND2X1 U3626 ( .IN1(n3358), .IN2(g1440), .Q(n3408) );
  AND2X1 U3627 ( .IN1(n3359), .IN2(g1601), .Q(n3407) );
  OR2X1 U3628 ( .IN1(n3409), .IN2(n3410), .Q(g6500) );
  AND2X1 U3629 ( .IN1(n3358), .IN2(g1411), .Q(n3410) );
  AND2X1 U3630 ( .IN1(n3359), .IN2(g1580), .Q(n3409) );
  OR2X1 U3631 ( .IN1(n3411), .IN2(n3412), .Q(g6481) );
  AND2X1 U3632 ( .IN1(n3358), .IN2(g1436), .Q(n3412) );
  AND2X1 U3633 ( .IN1(n3359), .IN2(g1598), .Q(n3411) );
  OR2X1 U3634 ( .IN1(n3413), .IN2(n3414), .Q(g6480) );
  AND2X1 U3635 ( .IN1(n3358), .IN2(g1419), .Q(n3414) );
  AND2X1 U3636 ( .IN1(n3359), .IN2(g1577), .Q(n3413) );
  OR2X1 U3637 ( .IN1(n3415), .IN2(n3416), .Q(g6479) );
  AND2X1 U3638 ( .IN1(n3358), .IN2(g1432), .Q(n3416) );
  AND2X1 U3639 ( .IN1(n3359), .IN2(g1595), .Q(n3415) );
  OR2X1 U3640 ( .IN1(n3417), .IN2(n3418), .Q(g6478) );
  AND2X1 U3641 ( .IN1(n3358), .IN2(g1515), .Q(n3418) );
  AND2X1 U3642 ( .IN1(n3359), .IN2(g1574), .Q(n3417) );
  AND2X1 U3643 ( .IN1(n3419), .IN2(n3420), .Q(g6471) );
  XOR2X1 U3644 ( .IN1(n4313), .IN2(n2417), .Q(n3420) );
  OR2X1 U3645 ( .IN1(n3421), .IN2(n3422), .Q(g6470) );
  AND2X1 U3646 ( .IN1(n3358), .IN2(g1403), .Q(n3422) );
  AND2X1 U3647 ( .IN1(n3359), .IN2(g1592), .Q(n3421) );
  OR2X1 U3648 ( .IN1(n3423), .IN2(n3424), .Q(g6469) );
  AND2X1 U3649 ( .IN1(n3358), .IN2(g1520), .Q(n3424) );
  AND2X1 U3650 ( .IN1(n3359), .IN2(g1571), .Q(n3423) );
  OR2X1 U3651 ( .IN1(n3425), .IN2(n3426), .Q(g6468) );
  AND2X1 U3652 ( .IN1(n3358), .IN2(g1415), .Q(n3426) );
  AND2X1 U3653 ( .IN1(n3359), .IN2(g1567), .Q(n3425) );
  INVX0 U3654 ( .INP(n3358), .ZN(n3359) );
  OR2X1 U3655 ( .IN1(n1159), .IN2(n505), .Q(n3358) );
  AND2X1 U3656 ( .IN1(n3427), .IN2(g109), .Q(g6439) );
  XNOR3X1 U3657 ( .IN1(g143), .IN2(n2362), .IN3(n3428), .Q(n3427) );
  XOR2X1 U3658 ( .IN1(n2471), .IN2(n2364), .Q(n3428) );
  AND2X1 U3659 ( .IN1(n3429), .IN2(n3179), .Q(g6392) );
  OR2X1 U3660 ( .IN1(n505), .IN2(n3178), .Q(n3429) );
  INVX0 U3661 ( .INP(g881), .ZN(n3178) );
  AND2X1 U3662 ( .IN1(g109), .IN2(g197), .Q(g6333) );
  AND2X1 U3663 ( .IN1(g109), .IN2(n3020), .Q(g6332) );
  OR2X1 U3664 ( .IN1(n3430), .IN2(n3431), .Q(g6243) );
  XOR2X1 U3665 ( .IN1(n2443), .IN2(n1717), .Q(n3431) );
  AND2X1 U3666 ( .IN1(g109), .IN2(g1520), .Q(g6224) );
  AND2X1 U3667 ( .IN1(g109), .IN2(g1515), .Q(g6205) );
  AND2X1 U3668 ( .IN1(n2493), .IN2(n3041), .Q(g6179) );
  AND2X1 U3669 ( .IN1(n3432), .IN2(g6331), .Q(n2493) );
  AND2X1 U3670 ( .IN1(g201), .IN2(g109), .Q(g6331) );
  OR2X1 U3671 ( .IN1(n3433), .IN2(n3434), .Q(g6155) );
  AND3X1 U3672 ( .IN1(g1700), .IN2(g1707), .IN3(n1653), .Q(n3434) );
  AND2X1 U3673 ( .IN1(g4076), .IN2(g1690), .Q(n3433) );
  AND2X1 U3674 ( .IN1(n3435), .IN2(n3155), .Q(g6126) );
  INVX0 U3675 ( .INP(n3430), .ZN(n3155) );
  XOR2X1 U3676 ( .IN1(n2733), .IN2(n2432), .Q(n3435) );
  AND2X1 U3677 ( .IN1(n3436), .IN2(n2745), .Q(g6123) );
  XOR2X1 U3678 ( .IN1(n2732), .IN2(n2447), .Q(n3436) );
  OR2X1 U3679 ( .IN1(n3437), .IN2(n3438), .Q(g6099) );
  AND2X1 U3680 ( .IN1(n3439), .IN2(g1074), .Q(n3438) );
  AND2X1 U3681 ( .IN1(n3440), .IN2(g342), .Q(n3437) );
  OR2X1 U3682 ( .IN1(n3441), .IN2(n3442), .Q(g6096) );
  AND2X1 U3683 ( .IN1(n3439), .IN2(g1098), .Q(n3442) );
  AND2X1 U3684 ( .IN1(n3440), .IN2(g366), .Q(n3441) );
  OR2X1 U3685 ( .IN1(n3443), .IN2(n3444), .Q(g6093) );
  AND2X1 U3686 ( .IN1(n3439), .IN2(g1095), .Q(n3444) );
  AND2X1 U3687 ( .IN1(n3440), .IN2(g363), .Q(n3443) );
  OR2X1 U3688 ( .IN1(n3445), .IN2(n3446), .Q(g6088) );
  AND2X1 U3689 ( .IN1(n3439), .IN2(g1092), .Q(n3446) );
  AND2X1 U3690 ( .IN1(n3440), .IN2(g360), .Q(n3445) );
  OR2X1 U3691 ( .IN1(n3447), .IN2(n3448), .Q(g6080) );
  AND2X1 U3692 ( .IN1(n3439), .IN2(g1089), .Q(n3448) );
  AND2X1 U3693 ( .IN1(n3440), .IN2(g357), .Q(n3447) );
  OR2X1 U3694 ( .IN1(n3449), .IN2(n3450), .Q(g6071) );
  AND2X1 U3695 ( .IN1(n3439), .IN2(g1086), .Q(n3450) );
  AND2X1 U3696 ( .IN1(n3440), .IN2(g354), .Q(n3449) );
  OR2X1 U3697 ( .IN1(n3451), .IN2(n3452), .Q(g6068) );
  AND2X1 U3698 ( .IN1(n3439), .IN2(g1083), .Q(n3452) );
  AND2X1 U3699 ( .IN1(n3440), .IN2(g351), .Q(n3451) );
  OR2X1 U3700 ( .IN1(n3453), .IN2(n3454), .Q(g6059) );
  AND2X1 U3701 ( .IN1(n3439), .IN2(g1080), .Q(n3454) );
  AND2X1 U3702 ( .IN1(n3440), .IN2(g348), .Q(n3453) );
  OR2X1 U3703 ( .IN1(n3455), .IN2(n3456), .Q(g6054) );
  AND2X1 U3704 ( .IN1(test_so7), .IN2(n3439), .Q(n3456) );
  AND2X1 U3705 ( .IN1(n3440), .IN2(g336), .Q(n3455) );
  OR2X1 U3706 ( .IN1(n3457), .IN2(n3458), .Q(g6049) );
  AND2X1 U3707 ( .IN1(n2985), .IN2(g549), .Q(n3458) );
  OR2X1 U3708 ( .IN1(n3459), .IN2(n3460), .Q(g6045) );
  AND2X1 U3709 ( .IN1(n2985), .IN2(g575), .Q(n3460) );
  OR2X1 U3710 ( .IN1(n3461), .IN2(n3462), .Q(g6042) );
  AND2X1 U3711 ( .IN1(n2985), .IN2(g572), .Q(n3462) );
  OR2X1 U3712 ( .IN1(n3463), .IN2(n3052), .Q(g6038) );
  AND2X1 U3713 ( .IN1(n2985), .IN2(g569), .Q(n3463) );
  OR2X1 U3714 ( .IN1(n3464), .IN2(n3010), .Q(g6035) );
  AND2X1 U3715 ( .IN1(n2985), .IN2(g566), .Q(n3464) );
  OR2X1 U3716 ( .IN1(n3465), .IN2(n2993), .Q(g6026) );
  AND2X1 U3717 ( .IN1(n2985), .IN2(g563), .Q(n3465) );
  OR2X1 U3718 ( .IN1(n3466), .IN2(n2983), .Q(g6015) );
  AND2X1 U3719 ( .IN1(n2985), .IN2(g560), .Q(n3466) );
  OR2X1 U3720 ( .IN1(n3467), .IN2(n3068), .Q(g6002) );
  AND2X1 U3721 ( .IN1(n2985), .IN2(g557), .Q(n3467) );
  OR2X1 U3722 ( .IN1(n3468), .IN2(n3021), .Q(g6000) );
  AND2X1 U3723 ( .IN1(n2985), .IN2(g554), .Q(n3468) );
  OR2X1 U3724 ( .IN1(n3469), .IN2(n3004), .Q(g5996) );
  AND2X1 U3725 ( .IN1(n2985), .IN2(g546), .Q(n3469) );
  OR2X1 U3726 ( .IN1(n3470), .IN2(n1195), .Q(g5918) );
  AND2X1 U3727 ( .IN1(g109), .IN2(g119), .Q(n3470) );
  OR2X1 U3728 ( .IN1(n3471), .IN2(n3472), .Q(g5914) );
  AND2X1 U3729 ( .IN1(n3439), .IN2(g1077), .Q(n3472) );
  AND2X1 U3730 ( .IN1(n3440), .IN2(g345), .Q(n3471) );
  OR2X1 U3731 ( .IN1(n3473), .IN2(n3474), .Q(g5910) );
  AND2X1 U3732 ( .IN1(n3439), .IN2(g1071), .Q(n3474) );
  AND2X1 U3733 ( .IN1(n3440), .IN2(g339), .Q(n3473) );
  OR2X1 U3734 ( .IN1(n3475), .IN2(n3476), .Q(g5770) );
  AND2X1 U3735 ( .IN1(g6180), .IN2(n3477), .Q(n3476) );
  INVX0 U3736 ( .INP(n3478), .ZN(n3477) );
  AND2X1 U3737 ( .IN1(g1453), .IN2(g109), .Q(g6180) );
  AND3X1 U3738 ( .IN1(n1628), .IN2(g109), .IN3(n3478), .Q(n3475) );
  XOR3X1 U3739 ( .IN1(g1494), .IN2(n2365), .IN3(n1707), .Q(n3478) );
  OR2X1 U3740 ( .IN1(n3479), .IN2(n3480), .Q(g5755) );
  AND2X1 U3741 ( .IN1(g6334), .IN2(n3481), .Q(n3480) );
  AND2X1 U3742 ( .IN1(g1389), .IN2(g109), .Q(g6334) );
  AND3X1 U3743 ( .IN1(n1603), .IN2(g109), .IN3(n3482), .Q(n3479) );
  INVX0 U3744 ( .INP(n3481), .ZN(n3482) );
  XNOR3X1 U3745 ( .IN1(n1678), .IN2(n1619), .IN3(n3483), .Q(n3481) );
  OR2X1 U3746 ( .IN1(n42), .IN2(g1386), .Q(n3483) );
  AND2X1 U3747 ( .IN1(n3432), .IN2(n1619), .Q(n42) );
  INVX0 U3748 ( .INP(n3484), .ZN(n3432) );
  OR4X1 U3749 ( .IN1(n3485), .IN2(n3486), .IN3(n3487), .IN4(n3488), .Q(n3484)
         );
  OR4X1 U3750 ( .IN1(g213), .IN2(g237), .IN3(g186), .IN4(n3489), .Q(n3488) );
  OR3X1 U3751 ( .IN1(g243), .IN2(g1386), .IN3(g192), .Q(n3489) );
  OR4X1 U3752 ( .IN1(test_so3), .IN2(g248), .IN3(g1389), .IN4(n3490), .Q(n3487) );
  OR3X1 U3753 ( .IN1(g1400), .IN2(g197), .IN3(g1397), .Q(n3490) );
  OR4X1 U3754 ( .IN1(g1371), .IN2(n3020), .IN3(n3061), .IN4(n3491), .Q(n3486)
         );
  OR2X1 U3755 ( .IN1(g1383), .IN2(n3054), .Q(n3491) );
  INVX0 U3756 ( .INP(n3492), .ZN(n3485) );
  AND4X1 U3757 ( .IN1(n2460), .IN2(n4315), .IN3(n4314), .IN4(n3493), .Q(n3492)
         );
  AND3X1 U3758 ( .IN1(n2457), .IN2(n2458), .IN3(n2459), .Q(n3493) );
  AND3X1 U3759 ( .IN1(g743), .IN2(g109), .IN3(g744), .Q(g5659) );
  AND3X1 U3760 ( .IN1(g741), .IN2(g109), .IN3(g742), .Q(g5658) );
  AND2X1 U3761 ( .IN1(n3494), .IN2(n2733), .Q(g5543) );
  OR2X1 U3762 ( .IN1(n1622), .IN2(n3079), .Q(n2733) );
  OR2X1 U3763 ( .IN1(n1717), .IN2(n2443), .Q(n3079) );
  INVX0 U3764 ( .INP(n3495), .ZN(n3494) );
  AND2X1 U3765 ( .IN1(n3496), .IN2(n3497), .Q(n3495) );
  OR2X1 U3766 ( .IN1(g5849), .IN2(n1717), .Q(n3497) );
  OR2X1 U3767 ( .IN1(n2443), .IN2(n3430), .Q(g5849) );
  OR2X1 U3768 ( .IN1(n3430), .IN2(n1622), .Q(n3496) );
  OR3X1 U3769 ( .IN1(n2464), .IN2(n2463), .IN3(n505), .Q(n3430) );
  AND3X1 U3770 ( .IN1(n2732), .IN2(n3498), .IN3(n2745), .Q(g5536) );
  INVX0 U3771 ( .INP(n1213), .ZN(n3498) );
  INVX0 U3772 ( .INP(n1193), .ZN(n2732) );
  OR2X1 U3773 ( .IN1(n3499), .IN2(n3500), .Q(g5529) );
  AND3X1 U3774 ( .IN1(n2745), .IN2(g4173), .IN3(n2452), .Q(n3500) );
  AND2X1 U3775 ( .IN1(g4940), .IN2(g4174), .Q(n3499) );
  OR2X1 U3776 ( .IN1(n3501), .IN2(n1195), .Q(g5445) );
  AND2X1 U3777 ( .IN1(g109), .IN2(g12), .Q(n3501) );
  OR2X1 U3778 ( .IN1(n3502), .IN2(n1195), .Q(g5421) );
  AND2X1 U3779 ( .IN1(g109), .IN2(g9), .Q(n3502) );
  OR2X1 U3780 ( .IN1(n3503), .IN2(n3504), .Q(g5404) );
  AND2X1 U3781 ( .IN1(n371), .IN2(g1718), .Q(n3504) );
  AND2X1 U3782 ( .IN1(n2971), .IN2(g1713), .Q(n3503) );
  OR2X1 U3783 ( .IN1(n3505), .IN2(n3506), .Q(g5396) );
  AND2X1 U3784 ( .IN1(n371), .IN2(g1713), .Q(n3506) );
  AND2X1 U3785 ( .IN1(n2971), .IN2(g1710), .Q(n3505) );
  AND2X1 U3786 ( .IN1(n3507), .IN2(g1101), .Q(g5390) );
  AND2X1 U3787 ( .IN1(n3507), .IN2(g1110), .Q(g5173) );
  AND2X1 U3788 ( .IN1(n3507), .IN2(g1107), .Q(g5148) );
  AND2X1 U3789 ( .IN1(n3507), .IN2(g1104), .Q(g5126) );
  INVX0 U3790 ( .INP(n3508), .ZN(n3507) );
  OR2X1 U3791 ( .IN1(n505), .IN2(n3056), .Q(n3508) );
  AND3X1 U3792 ( .IN1(n371), .IN2(n3339), .IN3(n3509), .Q(g5083) );
  INVX0 U3793 ( .INP(g4089), .ZN(n3339) );
  AND2X1 U3794 ( .IN1(n2745), .IN2(n2451), .Q(g4940) );
  AND2X1 U3795 ( .IN1(n2503), .IN2(g109), .Q(n2745) );
  AND2X1 U3796 ( .IN1(n3510), .IN2(n3018), .Q(g4905) );
  AND2X1 U3797 ( .IN1(n3510), .IN2(n3037), .Q(g4903) );
  AND2X1 U3798 ( .IN1(n3510), .IN2(n3030), .Q(g4902) );
  INVX0 U3799 ( .INP(n2499), .ZN(n3510) );
  AND2X1 U3800 ( .IN1(n3511), .IN2(n3053), .Q(g4893) );
  AND2X1 U3801 ( .IN1(n3511), .IN2(n3055), .Q(g4891) );
  AND2X1 U3802 ( .IN1(n3511), .IN2(n3035), .Q(g4890) );
  INVX0 U3803 ( .INP(n2497), .ZN(n3511) );
  OR2X1 U3804 ( .IN1(n3512), .IN2(n2784), .Q(n2497) );
  INVX0 U3805 ( .INP(n2965), .ZN(n2784) );
  OR4X1 U3806 ( .IN1(g605), .IN2(g611), .IN3(g591), .IN4(g599), .Q(n2965) );
  AND2X1 U3807 ( .IN1(n1607), .IN2(g611), .Q(n3512) );
  AND2X1 U3808 ( .IN1(g109), .IN2(n3016), .Q(g4506) );
  AND2X1 U3809 ( .IN1(n371), .IN2(n3046), .Q(g4500) );
  AND2X1 U3810 ( .IN1(g109), .IN2(g1145), .Q(g4498) );
  AND2X1 U3811 ( .IN1(g109), .IN2(g1137), .Q(g4484) );
  AND2X1 U3812 ( .IN1(test_so4), .IN2(g109), .Q(g4465) );
  AND2X1 U3813 ( .IN1(g109), .IN2(g1149), .Q(g4342) );
  AND2X1 U3814 ( .IN1(g109), .IN2(g1153), .Q(g4340) );
  OR2X1 U3815 ( .IN1(n3513), .IN2(n3514), .Q(g4309) );
  AND2X1 U3816 ( .IN1(n3515), .IN2(g1762), .Q(n3514) );
  AND2X1 U3817 ( .IN1(n3516), .IN2(g1806), .Q(n3513) );
  OR2X1 U3818 ( .IN1(n3517), .IN2(n3518), .Q(g4293) );
  AND2X1 U3819 ( .IN1(n3515), .IN2(g1759), .Q(n3518) );
  AND2X1 U3820 ( .IN1(n3516), .IN2(g1801), .Q(n3517) );
  OR2X1 U3821 ( .IN1(n3519), .IN2(n3520), .Q(g4283) );
  AND2X1 U3822 ( .IN1(n3515), .IN2(g1756), .Q(n3520) );
  AND2X1 U3823 ( .IN1(n3516), .IN2(g1796), .Q(n3519) );
  OR2X1 U3824 ( .IN1(n3521), .IN2(n3522), .Q(g4274) );
  AND2X1 U3825 ( .IN1(n3515), .IN2(g1753), .Q(n3522) );
  AND2X1 U3826 ( .IN1(n3516), .IN2(g1791), .Q(n3521) );
  OR2X1 U3827 ( .IN1(n3523), .IN2(n3524), .Q(g4264) );
  AND2X1 U3828 ( .IN1(n3515), .IN2(g1750), .Q(n3524) );
  AND2X1 U3829 ( .IN1(n3516), .IN2(g1786), .Q(n3523) );
  OR2X1 U3830 ( .IN1(n3525), .IN2(n3526), .Q(g4255) );
  AND2X1 U3831 ( .IN1(n3515), .IN2(g1747), .Q(n3526) );
  AND2X1 U3832 ( .IN1(n3516), .IN2(g1781), .Q(n3525) );
  OR2X1 U3833 ( .IN1(n3527), .IN2(n3528), .Q(g4239) );
  AND2X1 U3834 ( .IN1(n3515), .IN2(g1744), .Q(n3528) );
  AND2X1 U3835 ( .IN1(n3516), .IN2(g1776), .Q(n3527) );
  OR2X1 U3836 ( .IN1(n3529), .IN2(n3530), .Q(g4238) );
  AND2X1 U3837 ( .IN1(n3515), .IN2(g1741), .Q(n3530) );
  AND2X1 U3838 ( .IN1(n3516), .IN2(test_so5), .Q(n3529) );
  OR2X1 U3839 ( .IN1(n3531), .IN2(n3532), .Q(g4231) );
  AND2X1 U3840 ( .IN1(n3515), .IN2(g1738), .Q(n3532) );
  AND2X1 U3841 ( .IN1(n3516), .IN2(g1766), .Q(n3531) );
  OR2X1 U3842 ( .IN1(n507), .IN2(n3042), .Q(g4089) );
  INVX0 U3843 ( .INP(g1700), .ZN(n507) );
  AND2X1 U3844 ( .IN1(g1700), .IN2(n2397), .Q(g4076) );
  AND4X1 U3845 ( .IN1(g932), .IN2(g928), .IN3(g936), .IN4(g940), .Q(g3381) );
  INVX0 U3846 ( .INP(g23), .ZN(g3327) );
  AND2X1 U3847 ( .IN1(n2468), .IN2(n2398), .Q(g2478) );
  OR2X1 U3848 ( .IN1(n3533), .IN2(n3534), .Q(g11647) );
  AND2X1 U3849 ( .IN1(n3270), .IN2(n3535), .Q(n3534) );
  OR2X1 U3850 ( .IN1(n3536), .IN2(n3537), .Q(n3535) );
  AND2X1 U3851 ( .IN1(n3538), .IN2(n3539), .Q(n3537) );
  AND2X1 U3852 ( .IN1(n3540), .IN2(n3541), .Q(n3536) );
  INVX0 U3853 ( .INP(n3538), .ZN(n3541) );
  AND2X1 U3854 ( .IN1(n2710), .IN2(g336), .Q(n3533) );
  AND2X1 U3855 ( .IN1(n3542), .IN2(n3543), .Q(g11641) );
  INVX0 U3856 ( .INP(n3544), .ZN(n3542) );
  AND2X1 U3857 ( .IN1(n3545), .IN2(n3546), .Q(n3544) );
  OR2X1 U3858 ( .IN1(n1226), .IN2(n1721), .Q(n3546) );
  AND2X1 U3859 ( .IN1(n7), .IN2(n2498), .Q(n1226) );
  INVX0 U3860 ( .INP(n1227), .ZN(n7) );
  OR2X1 U3861 ( .IN1(n3547), .IN2(n2498), .Q(n3545) );
  AND2X1 U3862 ( .IN1(g1351), .IN2(n1229), .Q(n2498) );
  AND2X1 U3863 ( .IN1(n3548), .IN2(n3543), .Q(g11640) );
  OR2X1 U3864 ( .IN1(n3549), .IN2(n3550), .Q(n3548) );
  AND2X1 U3865 ( .IN1(n1232), .IN2(n1231), .Q(n3550) );
  AND2X1 U3866 ( .IN1(n3547), .IN2(g1346), .Q(n3549) );
  OR2X1 U3867 ( .IN1(n1227), .IN2(n3551), .Q(n3547) );
  INVX0 U3868 ( .INP(n1229), .ZN(n3551) );
  AND3X1 U3869 ( .IN1(g1336), .IN2(g1346), .IN3(g1341), .Q(n1229) );
  AND2X1 U3870 ( .IN1(n3552), .IN2(n3543), .Q(g11639) );
  XOR2X1 U3871 ( .IN1(n1231), .IN2(g1341), .Q(n3552) );
  AND2X1 U3872 ( .IN1(n3553), .IN2(n3543), .Q(g11636) );
  OR2X1 U3873 ( .IN1(n3216), .IN2(n2713), .Q(n3543) );
  AND2X1 U3874 ( .IN1(g109), .IN2(n3554), .Q(n2713) );
  OR2X1 U3875 ( .IN1(n3036), .IN2(n3555), .Q(n3554) );
  AND2X1 U3876 ( .IN1(g3069), .IN2(n4318), .Q(n3555) );
  AND2X1 U3877 ( .IN1(g109), .IN2(n2465), .Q(n3216) );
  XOR2X1 U3878 ( .IN1(n1227), .IN2(n2383), .Q(n3553) );
  OR2X1 U3879 ( .IN1(n3556), .IN2(n3557), .Q(g11625) );
  AND2X1 U3880 ( .IN1(n3270), .IN2(n3558), .Q(n3557) );
  XOR2X1 U3881 ( .IN1(n3540), .IN2(n3539), .Q(n3558) );
  AND2X1 U3882 ( .IN1(n3559), .IN2(n3560), .Q(n3539) );
  OR2X1 U3883 ( .IN1(n3561), .IN2(n2492), .Q(n3560) );
  XNOR2X1 U3884 ( .IN1(n3562), .IN2(n3563), .Q(n3561) );
  AND2X1 U3885 ( .IN1(n1594), .IN2(n3564), .Q(n3563) );
  OR2X1 U3886 ( .IN1(n40), .IN2(n1681), .Q(n3559) );
  XOR3X1 U3887 ( .IN1(n3565), .IN2(n3566), .IN3(n3567), .Q(n3540) );
  XOR3X1 U3888 ( .IN1(n3568), .IN2(n3569), .IN3(n3570), .Q(n3567) );
  XOR2X1 U3889 ( .IN1(n3571), .IN2(n3572), .Q(n3570) );
  XOR3X1 U3890 ( .IN1(n3573), .IN2(n3574), .IN3(n3575), .Q(n3565) );
  XOR2X1 U3891 ( .IN1(n3576), .IN2(n3577), .Q(n3575) );
  AND2X1 U3892 ( .IN1(n2710), .IN2(g345), .Q(n3556) );
  OR2X1 U3893 ( .IN1(n3578), .IN2(n3579), .Q(g11610) );
  AND2X1 U3894 ( .IN1(n3580), .IN2(g1333), .Q(n3579) );
  AND2X1 U3895 ( .IN1(n3581), .IN2(g1806), .Q(n3578) );
  OR2X1 U3896 ( .IN1(n3582), .IN2(n3583), .Q(g11609) );
  AND2X1 U3897 ( .IN1(n3580), .IN2(g1330), .Q(n3583) );
  AND2X1 U3898 ( .IN1(n3581), .IN2(g1801), .Q(n3582) );
  OR2X1 U3899 ( .IN1(n3584), .IN2(n3585), .Q(g11608) );
  AND2X1 U3900 ( .IN1(n3580), .IN2(g1327), .Q(n3585) );
  AND2X1 U3901 ( .IN1(n3581), .IN2(g1796), .Q(n3584) );
  OR2X1 U3902 ( .IN1(n3586), .IN2(n3587), .Q(g11607) );
  AND2X1 U3903 ( .IN1(n3580), .IN2(g1324), .Q(n3587) );
  AND2X1 U3904 ( .IN1(n3581), .IN2(g1791), .Q(n3586) );
  OR2X1 U3905 ( .IN1(n3588), .IN2(n3589), .Q(g11606) );
  AND2X1 U3906 ( .IN1(n3580), .IN2(g1321), .Q(n3589) );
  AND2X1 U3907 ( .IN1(n3581), .IN2(g1786), .Q(n3588) );
  OR2X1 U3908 ( .IN1(n3590), .IN2(n3591), .Q(g11605) );
  AND2X1 U3909 ( .IN1(n3580), .IN2(g1318), .Q(n3591) );
  AND2X1 U3910 ( .IN1(n3581), .IN2(g1781), .Q(n3590) );
  OR2X1 U3911 ( .IN1(n3592), .IN2(n3593), .Q(g11604) );
  AND2X1 U3912 ( .IN1(n3580), .IN2(g1314), .Q(n3593) );
  AND2X1 U3913 ( .IN1(n3581), .IN2(g1776), .Q(n3592) );
  OR2X1 U3914 ( .IN1(n3594), .IN2(n3595), .Q(g11603) );
  AND2X1 U3915 ( .IN1(n3581), .IN2(test_so5), .Q(n3595) );
  AND2X1 U3916 ( .IN1(test_so9), .IN2(n3580), .Q(n3594) );
  OR2X1 U3917 ( .IN1(n3596), .IN2(n3597), .Q(g11602) );
  AND2X1 U3918 ( .IN1(n3580), .IN2(g1308), .Q(n3597) );
  AND2X1 U3919 ( .IN1(n3581), .IN2(g1766), .Q(n3596) );
  INVX0 U3920 ( .INP(n3580), .ZN(n3581) );
  OR2X1 U3921 ( .IN1(n2478), .IN2(n1227), .Q(n3580) );
  OR3X1 U3922 ( .IN1(n3598), .IN2(n3232), .IN3(n3230), .Q(n1227) );
  AND4X1 U3923 ( .IN1(n3599), .IN2(n3600), .IN3(n3601), .IN4(n3602), .Q(n3598)
         );
  AND3X1 U3924 ( .IN1(n3603), .IN2(n3604), .IN3(n3605), .Q(n3602) );
  AND3X1 U3925 ( .IN1(n3606), .IN2(n3607), .IN3(n3608), .Q(n3605) );
  XOR2X1 U3926 ( .IN1(n2323), .IN2(g1260), .Q(n3608) );
  XOR2X1 U3927 ( .IN1(n2322), .IN2(g1265), .Q(n3607) );
  XOR2X1 U3928 ( .IN1(n2374), .IN2(g1275), .Q(n3606) );
  XOR2X1 U3929 ( .IN1(n2376), .IN2(g1240), .Q(n3604) );
  XOR2X1 U3930 ( .IN1(g991), .IN2(n2353), .Q(n3603) );
  AND3X1 U3931 ( .IN1(n3609), .IN2(n3610), .IN3(n3611), .Q(n3601) );
  XOR2X1 U3932 ( .IN1(test_so2), .IN2(n2330), .Q(n3611) );
  XOR2X1 U3933 ( .IN1(n2502), .IN2(g1023), .Q(n3610) );
  XNOR2X1 U3934 ( .IN1(n3612), .IN2(n3613), .Q(n3609) );
  XOR2X1 U3935 ( .IN1(test_so8), .IN2(n2352), .Q(n3600) );
  XOR2X1 U3936 ( .IN1(n2354), .IN2(g1250), .Q(n3599) );
  OR2X1 U3937 ( .IN1(n3614), .IN2(n3615), .Q(g11579) );
  AND2X1 U3938 ( .IN1(n3616), .IN2(n2971), .Q(n3615) );
  XNOR2X1 U3939 ( .IN1(n2468), .IN2(n3617), .Q(n3616) );
  OR2X1 U3940 ( .IN1(n3618), .IN2(n3619), .Q(n3617) );
  AND2X1 U3941 ( .IN1(n1260), .IN2(n3620), .Q(n3619) );
  INVX0 U3942 ( .INP(n3621), .ZN(n3620) );
  AND2X1 U3943 ( .IN1(n3621), .IN2(n3622), .Q(n3618) );
  OR2X1 U3944 ( .IN1(n46), .IN2(n2703), .Q(n3622) );
  AND4X1 U3945 ( .IN1(n1658), .IN2(n1677), .IN3(n3623), .IN4(n3007), .Q(n2703)
         );
  INVX0 U3946 ( .INP(n3624), .ZN(n46) );
  OR2X1 U3947 ( .IN1(n3625), .IN2(n3623), .Q(n3624) );
  OR2X1 U3948 ( .IN1(n3626), .IN2(n3627), .Q(n3623) );
  AND2X1 U3949 ( .IN1(n1685), .IN2(n3628), .Q(n3627) );
  OR2X1 U3950 ( .IN1(n3629), .IN2(g1153), .Q(n3628) );
  AND4X1 U3951 ( .IN1(n3630), .IN2(n3631), .IN3(n3632), .IN4(n3633), .Q(n3629)
         );
  INVX0 U3952 ( .INP(n3634), .ZN(n3633) );
  OR4X1 U3953 ( .IN1(g1121), .IN2(g1145), .IN3(g1137), .IN4(test_so4), .Q(
        n3634) );
  AND3X1 U3954 ( .IN1(n1705), .IN2(n1660), .IN3(n1706), .Q(n3632) );
  AND3X1 U3955 ( .IN1(n2422), .IN2(n1708), .IN3(n2423), .Q(n3631) );
  AND3X1 U3956 ( .IN1(n2425), .IN2(n2424), .IN3(n4316), .Q(n3630) );
  AND2X1 U3957 ( .IN1(n1686), .IN2(g1149), .Q(n3626) );
  AND3X1 U3958 ( .IN1(n1658), .IN2(n3007), .IN3(n1677), .Q(n3625) );
  AND2X1 U3959 ( .IN1(g1101), .IN2(n1614), .Q(n3007) );
  AND2X1 U3960 ( .IN1(n371), .IN2(g1618), .Q(n3614) );
  OR2X1 U3961 ( .IN1(n3635), .IN2(n3636), .Q(g11514) );
  AND2X1 U3962 ( .IN1(g6193), .IN2(n3637), .Q(n3636) );
  INVX0 U3963 ( .INP(n3638), .ZN(n3637) );
  AND2X1 U3964 ( .IN1(g1419), .IN2(g109), .Q(g6193) );
  AND3X1 U3965 ( .IN1(n1602), .IN2(g109), .IN3(n3638), .Q(n3635) );
  XNOR3X1 U3966 ( .IN1(n1627), .IN2(n3639), .IN3(n3621), .Q(n3638) );
  OR2X1 U3967 ( .IN1(n3640), .IN2(n3641), .Q(n3621) );
  AND2X1 U3968 ( .IN1(n3642), .IN2(n2985), .Q(n3641) );
  OR2X1 U3969 ( .IN1(n3643), .IN2(n3644), .Q(n3642) );
  INVX0 U3970 ( .INP(n3645), .ZN(n3644) );
  OR2X1 U3971 ( .IN1(n3646), .IN2(n3647), .Q(n3645) );
  AND2X1 U3972 ( .IN1(n3648), .IN2(n3649), .Q(n3646) );
  AND2X1 U3973 ( .IN1(n3647), .IN2(n1699), .Q(n3643) );
  AND4X1 U3974 ( .IN1(n4320), .IN2(n4319), .IN3(n4322), .IN4(n4321), .Q(n3647)
         );
  AND2X1 U3975 ( .IN1(g18), .IN2(g201), .Q(n3640) );
  XOR2X1 U3976 ( .IN1(g1448), .IN2(g1415), .Q(n3639) );
  OR2X1 U3977 ( .IN1(n3650), .IN2(n3651), .Q(g11488) );
  INVX0 U3978 ( .INP(n3652), .ZN(n3651) );
  OR2X1 U3979 ( .IN1(n2710), .IN2(n3577), .Q(n3652) );
  AND2X1 U3980 ( .IN1(n3653), .IN2(n3654), .Q(n3577) );
  OR2X1 U3981 ( .IN1(n3655), .IN2(n2492), .Q(n3654) );
  XOR2X1 U3982 ( .IN1(n3656), .IN2(g516), .Q(n3655) );
  OR4X1 U3983 ( .IN1(g466), .IN2(g461), .IN3(n1641), .IN4(n1606), .Q(n3656) );
  OR2X1 U3984 ( .IN1(n40), .IN2(n2201), .Q(n3653) );
  AND2X1 U3985 ( .IN1(n2710), .IN2(g342), .Q(n3650) );
  OR2X1 U3986 ( .IN1(n3657), .IN2(n3658), .Q(g11487) );
  AND2X1 U3987 ( .IN1(n3270), .IN2(n3574), .Q(n3658) );
  OR2X1 U3988 ( .IN1(n3659), .IN2(n3660), .Q(n3574) );
  AND2X1 U3989 ( .IN1(n3661), .IN2(n40), .Q(n3660) );
  XOR2X1 U3990 ( .IN1(g511), .IN2(n3662), .Q(n3661) );
  AND2X1 U3991 ( .IN1(n3663), .IN2(n1594), .Q(n3662) );
  AND2X1 U3992 ( .IN1(n2492), .IN2(g333), .Q(n3659) );
  AND2X1 U3993 ( .IN1(n2710), .IN2(g366), .Q(n3657) );
  OR2X1 U3994 ( .IN1(n3664), .IN2(n3665), .Q(g11486) );
  AND2X1 U3995 ( .IN1(n3270), .IN2(n3576), .Q(n3665) );
  OR2X1 U3996 ( .IN1(n3666), .IN2(n3667), .Q(n3576) );
  AND2X1 U3997 ( .IN1(n3668), .IN2(n40), .Q(n3667) );
  XOR2X1 U3998 ( .IN1(n3669), .IN2(n1600), .Q(n3668) );
  OR2X1 U3999 ( .IN1(g471), .IN2(n3670), .Q(n3669) );
  AND2X1 U4000 ( .IN1(n2492), .IN2(g330), .Q(n3666) );
  AND2X1 U4001 ( .IN1(n2710), .IN2(g363), .Q(n3664) );
  OR2X1 U4002 ( .IN1(n3671), .IN2(n3672), .Q(g11485) );
  INVX0 U4003 ( .INP(n3673), .ZN(n3672) );
  OR2X1 U4004 ( .IN1(n2710), .IN2(n3573), .Q(n3673) );
  AND2X1 U4005 ( .IN1(n3674), .IN2(n3675), .Q(n3573) );
  OR2X1 U4006 ( .IN1(n3676), .IN2(n2492), .Q(n3675) );
  XOR2X1 U4007 ( .IN1(n3677), .IN2(g501), .Q(n3676) );
  OR2X1 U4008 ( .IN1(n1646), .IN2(n3678), .Q(n3677) );
  OR2X1 U4009 ( .IN1(n40), .IN2(n2360), .Q(n3674) );
  AND2X1 U4010 ( .IN1(n2710), .IN2(g360), .Q(n3671) );
  OR2X1 U4011 ( .IN1(n3679), .IN2(n3680), .Q(g11484) );
  AND2X1 U4012 ( .IN1(n3270), .IN2(n3571), .Q(n3680) );
  OR2X1 U4013 ( .IN1(n3681), .IN2(n3682), .Q(n3571) );
  AND2X1 U4014 ( .IN1(n3683), .IN2(n40), .Q(n3682) );
  XOR2X1 U4015 ( .IN1(g496), .IN2(n3684), .Q(n3683) );
  AND2X1 U4016 ( .IN1(n3685), .IN2(g456), .Q(n3684) );
  AND2X1 U4017 ( .IN1(n2492), .IN2(g324), .Q(n3681) );
  AND2X1 U4018 ( .IN1(n2710), .IN2(g357), .Q(n3679) );
  OR2X1 U4019 ( .IN1(n3686), .IN2(n3687), .Q(g11483) );
  INVX0 U4020 ( .INP(n3688), .ZN(n3687) );
  OR2X1 U4021 ( .IN1(n2710), .IN2(n3572), .Q(n3688) );
  AND2X1 U4022 ( .IN1(n3689), .IN2(n3690), .Q(n3572) );
  OR2X1 U4023 ( .IN1(n3691), .IN2(n2492), .Q(n3690) );
  XOR2X1 U4024 ( .IN1(n1691), .IN2(n3692), .Q(n3691) );
  AND2X1 U4025 ( .IN1(n3685), .IN2(n1641), .Q(n3692) );
  AND3X1 U4026 ( .IN1(g466), .IN2(n1606), .IN3(n1594), .Q(n3685) );
  OR2X1 U4027 ( .IN1(n40), .IN2(n2380), .Q(n3689) );
  AND2X1 U4028 ( .IN1(n2710), .IN2(g354), .Q(n3686) );
  OR2X1 U4029 ( .IN1(n3693), .IN2(n3694), .Q(g11482) );
  INVX0 U4030 ( .INP(n3695), .ZN(n3694) );
  OR2X1 U4031 ( .IN1(n2710), .IN2(n3566), .Q(n3695) );
  AND2X1 U4032 ( .IN1(n3696), .IN2(n3697), .Q(n3566) );
  OR2X1 U4033 ( .IN1(n3698), .IN2(n2492), .Q(n3697) );
  XOR2X1 U4034 ( .IN1(n1621), .IN2(n3699), .Q(n3698) );
  AND2X1 U4035 ( .IN1(n3564), .IN2(g461), .Q(n3699) );
  AND3X1 U4036 ( .IN1(g456), .IN2(n1606), .IN3(n1646), .Q(n3564) );
  OR2X1 U4037 ( .IN1(n40), .IN2(n2358), .Q(n3696) );
  AND2X1 U4038 ( .IN1(n2710), .IN2(g351), .Q(n3693) );
  OR2X1 U4039 ( .IN1(n3700), .IN2(n3701), .Q(g11481) );
  AND2X1 U4040 ( .IN1(n3270), .IN2(n3568), .Q(n3701) );
  OR2X1 U4041 ( .IN1(n3702), .IN2(n3703), .Q(n3568) );
  AND2X1 U4042 ( .IN1(n3704), .IN2(n40), .Q(n3703) );
  XOR2X1 U4043 ( .IN1(n3705), .IN2(n1680), .Q(n3704) );
  OR2X1 U4044 ( .IN1(g466), .IN2(n3678), .Q(n3705) );
  OR3X1 U4045 ( .IN1(n1594), .IN2(g471), .IN3(g456), .Q(n3678) );
  AND2X1 U4046 ( .IN1(n2492), .IN2(g315), .Q(n3702) );
  AND2X1 U4047 ( .IN1(n2710), .IN2(g348), .Q(n3700) );
  OR2X1 U4048 ( .IN1(n3706), .IN2(n3707), .Q(g11478) );
  AND2X1 U4049 ( .IN1(n3270), .IN2(n3569), .Q(n3707) );
  OR2X1 U4050 ( .IN1(n3708), .IN2(n3709), .Q(n3569) );
  AND2X1 U4051 ( .IN1(n3710), .IN2(n40), .Q(n3709) );
  XOR2X1 U4052 ( .IN1(g476), .IN2(n3711), .Q(n3710) );
  AND2X1 U4053 ( .IN1(n3663), .IN2(g461), .Q(n3711) );
  AND3X1 U4054 ( .IN1(g471), .IN2(n1646), .IN3(n1641), .Q(n3663) );
  AND2X1 U4055 ( .IN1(n2492), .IN2(g312), .Q(n3708) );
  AND2X1 U4056 ( .IN1(n2710), .IN2(g339), .Q(n3706) );
  INVX0 U4057 ( .INP(n3270), .ZN(n2710) );
  AND2X1 U4058 ( .IN1(g750), .IN2(n1647), .Q(n3270) );
  OR2X1 U4059 ( .IN1(n3712), .IN2(n3713), .Q(g11443) );
  AND2X1 U4060 ( .IN1(n3239), .IN2(g1275), .Q(n3713) );
  AND2X1 U4061 ( .IN1(g109), .IN2(n3230), .Q(n3239) );
  AND2X1 U4062 ( .IN1(n3218), .IN2(n3612), .Q(n3712) );
  OR2X1 U4063 ( .IN1(n3714), .IN2(n3715), .Q(n3612) );
  AND2X1 U4064 ( .IN1(n3716), .IN2(n3229), .Q(n3715) );
  INVX0 U4065 ( .INP(n3232), .ZN(n3229) );
  OR2X1 U4066 ( .IN1(n3717), .IN2(n3718), .Q(n3716) );
  AND2X1 U4067 ( .IN1(n1862), .IN2(n3719), .Q(n3718) );
  OR2X1 U4068 ( .IN1(n3720), .IN2(g1284), .Q(n3719) );
  AND4X1 U4069 ( .IN1(n3721), .IN2(n3722), .IN3(n3723), .IN4(n3724), .Q(n3720)
         );
  AND4X1 U4070 ( .IN1(n2333), .IN2(n2331), .IN3(n2330), .IN4(n2502), .Q(n3724)
         );
  AND3X1 U4071 ( .IN1(n2335), .IN2(n2334), .IN3(n2336), .Q(n3723) );
  AND3X1 U4072 ( .IN1(n2352), .IN2(n2337), .IN3(n2353), .Q(n3722) );
  AND3X1 U4073 ( .IN1(n2373), .IN2(n2355), .IN3(n2375), .Q(n3721) );
  AND2X1 U4074 ( .IN1(n1864), .IN2(g1280), .Q(n3717) );
  AND2X1 U4075 ( .IN1(n3613), .IN2(n3232), .Q(n3714) );
  OR2X1 U4076 ( .IN1(n2462), .IN2(n3228), .Q(n3232) );
  OR3X1 U4077 ( .IN1(n2472), .IN2(n2449), .IN3(n2448), .Q(n3228) );
  XNOR2X1 U4078 ( .IN1(n3725), .IN2(g1027), .Q(n3613) );
  OR2X1 U4079 ( .IN1(n3538), .IN2(n2477), .Q(n3725) );
  INVX0 U4080 ( .INP(n3230), .ZN(n3218) );
  OR3X1 U4081 ( .IN1(n2391), .IN2(n371), .IN3(g1713), .Q(n3230) );
  AND2X1 U4082 ( .IN1(n3726), .IN2(n3727), .Q(g11393) );
  XOR2X1 U4083 ( .IN1(g986), .IN2(n3728), .Q(n3726) );
  AND2X1 U4084 ( .IN1(n3729), .IN2(n3727), .Q(g11392) );
  OR2X1 U4085 ( .IN1(n3730), .IN2(n3731), .Q(n3729) );
  AND2X1 U4086 ( .IN1(n3732), .IN2(g981), .Q(n3731) );
  INVX0 U4087 ( .INP(n3728), .ZN(n3732) );
  AND2X1 U4088 ( .IN1(n2712), .IN2(n2490), .Q(n3728) );
  AND3X1 U4089 ( .IN1(n3733), .IN2(g976), .IN3(n3734), .Q(n3730) );
  INVX0 U4090 ( .INP(n2712), .ZN(n3733) );
  AND3X1 U4091 ( .IN1(g976), .IN2(g971), .IN3(g981), .Q(n2712) );
  AND2X1 U4092 ( .IN1(n3735), .IN2(n3727), .Q(g11391) );
  XOR2X1 U4093 ( .IN1(g976), .IN2(n3734), .Q(n3735) );
  AND2X1 U4094 ( .IN1(n3736), .IN2(n3737), .Q(g11380) );
  OR2X1 U4095 ( .IN1(n3738), .IN2(g471), .Q(n3737) );
  AND2X1 U4096 ( .IN1(n3739), .IN2(n3740), .Q(n3738) );
  AND2X1 U4097 ( .IN1(n3736), .IN2(n3741), .Q(g11376) );
  OR2X1 U4098 ( .IN1(n3742), .IN2(n3743), .Q(n3741) );
  AND2X1 U4099 ( .IN1(n3744), .IN2(g466), .Q(n3743) );
  OR2X1 U4100 ( .IN1(n3670), .IN2(n3745), .Q(n3744) );
  AND3X1 U4101 ( .IN1(n3670), .IN2(g461), .IN3(n3746), .Q(n3742) );
  INVX0 U4102 ( .INP(n3740), .ZN(n3670) );
  AND2X1 U4103 ( .IN1(n3747), .IN2(n3736), .Q(g11372) );
  XOR2X1 U4104 ( .IN1(g461), .IN2(n3746), .Q(n3747) );
  INVX0 U4105 ( .INP(n3748), .ZN(n3746) );
  AND3X1 U4106 ( .IN1(n3727), .IN2(n3749), .IN3(n3750), .Q(g11349) );
  OR2X1 U4107 ( .IN1(n2490), .IN2(g971), .Q(n3750) );
  INVX0 U4108 ( .INP(n3734), .ZN(n3749) );
  AND2X1 U4109 ( .IN1(g971), .IN2(n2490), .Q(n3734) );
  AND3X1 U4110 ( .IN1(n40), .IN2(n3751), .IN3(n1420), .Q(n2490) );
  INVX0 U4111 ( .INP(n3752), .ZN(n3751) );
  AND4X1 U4112 ( .IN1(n3753), .IN2(n3754), .IN3(n3755), .IN4(n3756), .Q(n3752)
         );
  AND3X1 U4113 ( .IN1(n3757), .IN2(n3758), .IN3(n3759), .Q(n3756) );
  AND3X1 U4114 ( .IN1(n3760), .IN2(n3761), .IN3(n3762), .Q(n3759) );
  XOR2X1 U4115 ( .IN1(n2367), .IN2(g421), .Q(n3762) );
  XOR2X1 U4116 ( .IN1(n2369), .IN2(g411), .Q(n3761) );
  XOR2X1 U4117 ( .IN1(n2360), .IN2(g401), .Q(n3760) );
  XOR2X1 U4118 ( .IN1(n2378), .IN2(g426), .Q(n3758) );
  XOR2X1 U4119 ( .IN1(n2380), .IN2(g391), .Q(n3757) );
  AND3X1 U4120 ( .IN1(n3763), .IN2(n3764), .IN3(n3765), .Q(n3755) );
  XOR2X1 U4121 ( .IN1(n2200), .IN2(g406), .Q(n3765) );
  XOR2X1 U4122 ( .IN1(n2201), .IN2(g416), .Q(n3764) );
  XOR2X1 U4123 ( .IN1(n1681), .IN2(n3766), .Q(n3763) );
  XOR2X1 U4124 ( .IN1(n2356), .IN2(g396), .Q(n3754) );
  XOR2X1 U4125 ( .IN1(n2358), .IN2(g386), .Q(n3753) );
  OR2X1 U4126 ( .IN1(n3767), .IN2(n2495), .Q(n3727) );
  AND2X1 U4127 ( .IN1(g109), .IN2(n3768), .Q(n2495) );
  OR2X1 U4128 ( .IN1(n3064), .IN2(n3769), .Q(n3768) );
  AND2X1 U4129 ( .IN1(g3007), .IN2(n4317), .Q(n3769) );
  AND3X1 U4130 ( .IN1(n3770), .IN2(n3748), .IN3(n3736), .Q(g11340) );
  INVX0 U4131 ( .INP(n3771), .ZN(n3736) );
  OR2X1 U4132 ( .IN1(n505), .IN2(n3026), .Q(n3771) );
  OR2X1 U4133 ( .IN1(n1641), .IN2(n3745), .Q(n3748) );
  OR2X1 U4134 ( .IN1(n3739), .IN2(g456), .Q(n3770) );
  INVX0 U4135 ( .INP(n3745), .ZN(n3739) );
  OR2X1 U4136 ( .IN1(n3772), .IN2(n2492), .Q(n3745) );
  AND2X1 U4137 ( .IN1(n3740), .IN2(g471), .Q(n3772) );
  AND3X1 U4138 ( .IN1(g466), .IN2(g456), .IN3(g461), .Q(n3740) );
  OR2X1 U4139 ( .IN1(n3773), .IN2(n3774), .Q(g11338) );
  AND2X1 U4140 ( .IN1(n40), .IN2(g516), .Q(n3774) );
  AND2X1 U4141 ( .IN1(n2492), .IN2(g476), .Q(n3773) );
  OR2X1 U4142 ( .IN1(n3775), .IN2(n3776), .Q(g11337) );
  AND2X1 U4143 ( .IN1(n40), .IN2(g511), .Q(n3776) );
  AND2X1 U4144 ( .IN1(n2492), .IN2(g516), .Q(n3775) );
  OR2X1 U4145 ( .IN1(n3777), .IN2(n3778), .Q(g11336) );
  AND2X1 U4146 ( .IN1(n40), .IN2(g506), .Q(n3778) );
  AND2X1 U4147 ( .IN1(n2492), .IN2(g511), .Q(n3777) );
  OR2X1 U4148 ( .IN1(n3779), .IN2(n3780), .Q(g11335) );
  AND2X1 U4149 ( .IN1(n40), .IN2(g501), .Q(n3780) );
  AND2X1 U4150 ( .IN1(n2492), .IN2(g506), .Q(n3779) );
  OR2X1 U4151 ( .IN1(n3781), .IN2(n3782), .Q(g11334) );
  AND2X1 U4152 ( .IN1(n40), .IN2(g496), .Q(n3782) );
  AND2X1 U4153 ( .IN1(n2492), .IN2(g501), .Q(n3781) );
  OR2X1 U4154 ( .IN1(n3783), .IN2(n3784), .Q(g11333) );
  AND2X1 U4155 ( .IN1(n40), .IN2(g491), .Q(n3784) );
  AND2X1 U4156 ( .IN1(n2492), .IN2(g496), .Q(n3783) );
  OR2X1 U4157 ( .IN1(n3785), .IN2(n3786), .Q(g11332) );
  AND2X1 U4158 ( .IN1(n40), .IN2(g486), .Q(n3786) );
  AND2X1 U4159 ( .IN1(n2492), .IN2(g491), .Q(n3785) );
  OR2X1 U4160 ( .IN1(n3787), .IN2(n3788), .Q(g11331) );
  AND2X1 U4161 ( .IN1(n40), .IN2(g481), .Q(n3788) );
  AND2X1 U4162 ( .IN1(n2492), .IN2(g486), .Q(n3787) );
  OR2X1 U4163 ( .IN1(n3789), .IN2(n3790), .Q(g11330) );
  AND2X1 U4164 ( .IN1(n40), .IN2(g525), .Q(n3790) );
  AND2X1 U4165 ( .IN1(n2492), .IN2(g521), .Q(n3789) );
  OR2X1 U4166 ( .IN1(n3791), .IN2(n3792), .Q(g11329) );
  AND2X1 U4167 ( .IN1(n40), .IN2(g530), .Q(n3792) );
  AND2X1 U4168 ( .IN1(n2492), .IN2(g525), .Q(n3791) );
  OR2X1 U4169 ( .IN1(n3793), .IN2(n3794), .Q(g11328) );
  AND2X1 U4170 ( .IN1(n40), .IN2(g534), .Q(n3794) );
  AND2X1 U4171 ( .IN1(n2492), .IN2(g530), .Q(n3793) );
  OR2X1 U4172 ( .IN1(n3795), .IN2(n3796), .Q(g11327) );
  AND2X1 U4173 ( .IN1(n40), .IN2(g538), .Q(n3796) );
  AND2X1 U4174 ( .IN1(n2492), .IN2(g534), .Q(n3795) );
  OR2X1 U4175 ( .IN1(n3797), .IN2(n3798), .Q(g11326) );
  AND2X1 U4176 ( .IN1(n40), .IN2(g542), .Q(n3798) );
  AND2X1 U4177 ( .IN1(n2492), .IN2(g538), .Q(n3797) );
  OR2X1 U4178 ( .IN1(n3799), .IN2(n3800), .Q(g11325) );
  AND2X1 U4179 ( .IN1(n40), .IN2(g476), .Q(n3800) );
  AND2X1 U4180 ( .IN1(n2492), .IN2(g542), .Q(n3799) );
  OR2X1 U4181 ( .IN1(n3801), .IN2(n3802), .Q(g11324) );
  AND2X1 U4182 ( .IN1(n3562), .IN2(n40), .Q(n3802) );
  OR2X1 U4183 ( .IN1(n3803), .IN2(n3804), .Q(n3562) );
  AND2X1 U4184 ( .IN1(n1698), .IN2(n3805), .Q(n3804) );
  OR2X1 U4185 ( .IN1(n3806), .IN2(g525), .Q(n3805) );
  AND4X1 U4186 ( .IN1(n3807), .IN2(n3808), .IN3(n3809), .IN4(n3810), .Q(n3806)
         );
  AND4X1 U4187 ( .IN1(n1621), .IN2(n1620), .IN3(n1600), .IN4(n1599), .Q(n3810)
         );
  AND3X1 U4188 ( .IN1(n1680), .IN2(n1679), .IN3(n1689), .Q(n3809) );
  AND3X1 U4189 ( .IN1(n1691), .IN2(n1690), .IN3(n2407), .Q(n3808) );
  AND3X1 U4190 ( .IN1(n2409), .IN2(n2408), .IN3(n2410), .Q(n3807) );
  AND2X1 U4191 ( .IN1(n1695), .IN2(g521), .Q(n3803) );
  AND2X1 U4192 ( .IN1(n2492), .IN2(g481), .Q(n3801) );
  AND3X1 U4193 ( .IN1(n3811), .IN2(n3812), .IN3(n3767), .Q(g11320) );
  INVX0 U4194 ( .INP(n3813), .ZN(n3812) );
  OR2X1 U4195 ( .IN1(n3814), .IN2(g369), .Q(n3811) );
  OR2X1 U4196 ( .IN1(n3815), .IN2(n3816), .Q(g11314) );
  AND2X1 U4197 ( .IN1(n3817), .IN2(g968), .Q(n3816) );
  AND2X1 U4198 ( .IN1(n1855), .IN2(g861), .Q(n3815) );
  OR2X1 U4199 ( .IN1(n3818), .IN2(n3819), .Q(g11312) );
  AND2X1 U4200 ( .IN1(g965), .IN2(n3817), .Q(n3819) );
  AND2X1 U4201 ( .IN1(n1855), .IN2(g857), .Q(n3818) );
  OR2X1 U4202 ( .IN1(n3820), .IN2(n3821), .Q(g11310) );
  AND2X1 U4203 ( .IN1(g962), .IN2(n3817), .Q(n3821) );
  AND2X1 U4204 ( .IN1(n1855), .IN2(g853), .Q(n3820) );
  OR2X1 U4205 ( .IN1(n3822), .IN2(n3823), .Q(g11308) );
  AND2X1 U4206 ( .IN1(n3817), .IN2(g959), .Q(n3823) );
  AND2X1 U4207 ( .IN1(n1855), .IN2(g849), .Q(n3822) );
  OR2X1 U4208 ( .IN1(n3824), .IN2(n3825), .Q(g11306) );
  AND2X1 U4209 ( .IN1(n3817), .IN2(g956), .Q(n3825) );
  AND2X1 U4210 ( .IN1(n1855), .IN2(g845), .Q(n3824) );
  OR2X1 U4211 ( .IN1(n3826), .IN2(n3827), .Q(g11305) );
  AND2X1 U4212 ( .IN1(n3817), .IN2(g953), .Q(n3827) );
  AND2X1 U4213 ( .IN1(n1855), .IN2(g841), .Q(n3826) );
  OR2X1 U4214 ( .IN1(n3828), .IN2(n3829), .Q(g11303) );
  AND2X1 U4215 ( .IN1(n3817), .IN2(g950), .Q(n3829) );
  AND2X1 U4216 ( .IN1(n1855), .IN2(g837), .Q(n3828) );
  OR2X1 U4217 ( .IN1(n3830), .IN2(n3831), .Q(g11300) );
  AND2X1 U4218 ( .IN1(n3817), .IN2(g947), .Q(n3831) );
  AND2X1 U4219 ( .IN1(n1855), .IN2(g833), .Q(n3830) );
  OR2X1 U4220 ( .IN1(n3832), .IN2(n3833), .Q(g11298) );
  AND2X1 U4221 ( .IN1(n1855), .IN2(g829), .Q(n3833) );
  AND2X1 U4222 ( .IN1(n3817), .IN2(g944), .Q(n3832) );
  INVX0 U4223 ( .INP(n1855), .ZN(n3817) );
  OR3X1 U4224 ( .IN1(n3834), .IN2(n3835), .IN3(n3836), .Q(g11294) );
  AND2X1 U4225 ( .IN1(n2912), .IN2(n3837), .Q(n3836) );
  OR3X1 U4226 ( .IN1(n3838), .IN2(n3839), .IN3(n3840), .Q(n3837) );
  AND3X1 U4227 ( .IN1(n3841), .IN2(g1690), .IN3(n3842), .Q(n3840) );
  OR2X1 U4228 ( .IN1(n3843), .IN2(n3844), .Q(n3842) );
  OR2X1 U4229 ( .IN1(n3845), .IN2(n3846), .Q(n3841) );
  AND3X1 U4230 ( .IN1(n3847), .IN2(n3848), .IN3(g1690), .Q(n3839) );
  OR2X1 U4231 ( .IN1(n3849), .IN2(n3850), .Q(n3848) );
  OR2X1 U4232 ( .IN1(n3851), .IN2(n3648), .Q(n3847) );
  AND2X1 U4233 ( .IN1(n1653), .IN2(n3852), .Q(n3838) );
  OR2X1 U4234 ( .IN1(n3853), .IN2(n3854), .Q(n3852) );
  AND2X1 U4235 ( .IN1(n3855), .IN2(n3401), .Q(n3854) );
  OR2X1 U4236 ( .IN1(n2461), .IN2(n2504), .Q(n3401) );
  OR2X1 U4237 ( .IN1(n1659), .IN2(n1715), .Q(n3855) );
  AND2X1 U4238 ( .IN1(n3856), .IN2(n2740), .Q(n3853) );
  OR2X1 U4239 ( .IN1(n1702), .IN2(n2439), .Q(n2740) );
  OR2X1 U4240 ( .IN1(n1626), .IN2(n2427), .Q(n3856) );
  AND3X1 U4241 ( .IN1(n926), .IN2(n3857), .IN3(n1682), .Q(n3835) );
  INVX0 U4242 ( .INP(n3858), .ZN(n3857) );
  AND4X1 U4243 ( .IN1(n822), .IN2(n817), .IN3(n2767), .IN4(n2778), .Q(n3858)
         );
  INVX0 U4244 ( .INP(n3859), .ZN(n2767) );
  OR2X1 U4245 ( .IN1(n1605), .IN2(n1608), .Q(n817) );
  AND2X1 U4246 ( .IN1(n3419), .IN2(g1857), .Q(n3834) );
  INVX0 U4247 ( .INP(n2694), .ZN(n3419) );
  OR2X1 U4248 ( .IN1(n926), .IN2(n2912), .Q(n2694) );
  OR2X1 U4249 ( .IN1(n3860), .IN2(n3861), .Q(g11293) );
  AND2X1 U4250 ( .IN1(n3862), .IN2(n2912), .Q(n3861) );
  OR2X1 U4251 ( .IN1(n3863), .IN2(n3864), .Q(n3862) );
  AND2X1 U4252 ( .IN1(n1653), .IN2(n2426), .Q(n3864) );
  AND2X1 U4253 ( .IN1(n3846), .IN2(g1690), .Q(n3863) );
  AND2X1 U4254 ( .IN1(n3865), .IN2(n2764), .Q(n3860) );
  OR2X1 U4255 ( .IN1(n3866), .IN2(n3859), .Q(n3865) );
  AND3X1 U4256 ( .IN1(g1828), .IN2(n1643), .IN3(n1608), .Q(n3859) );
  AND2X1 U4257 ( .IN1(n3867), .IN2(g1854), .Q(n3866) );
  OR4X1 U4258 ( .IN1(n3868), .IN2(n2711), .IN3(n3869), .IN4(n3870), .Q(n3867)
         );
  AND2X1 U4259 ( .IN1(n1682), .IN2(n3871), .Q(n3870) );
  XOR2X1 U4260 ( .IN1(n1380), .IN2(n3872), .Q(n3871) );
  AND2X1 U4261 ( .IN1(n3873), .IN2(g1857), .Q(n3869) );
  XOR2X1 U4262 ( .IN1(n2778), .IN2(n3872), .Q(n3873) );
  OR2X1 U4263 ( .IN1(n2499), .IN2(n1873), .Q(n2711) );
  OR2X1 U4264 ( .IN1(n3874), .IN2(n2912), .Q(n2499) );
  INVX0 U4265 ( .INP(n2764), .ZN(n2912) );
  OR4X1 U4266 ( .IN1(g1814), .IN2(g1834), .IN3(g1828), .IN4(g1822), .Q(n2764)
         );
  AND2X1 U4267 ( .IN1(n1608), .IN2(g1834), .Q(n3874) );
  AND4X1 U4268 ( .IN1(n1380), .IN2(n3134), .IN3(n822), .IN4(n2778), .Q(n3868)
         );
  OR2X1 U4269 ( .IN1(n1643), .IN2(g1814), .Q(n2778) );
  OR2X1 U4270 ( .IN1(n1643), .IN2(g1828), .Q(n822) );
  OR4X1 U4271 ( .IN1(g1834), .IN2(n2879), .IN3(g1840), .IN4(g1828), .Q(n3134)
         );
  OR2X1 U4272 ( .IN1(n1608), .IN2(g1822), .Q(n2879) );
  AND2X1 U4273 ( .IN1(n3767), .IN2(n3875), .Q(g11292) );
  OR2X1 U4274 ( .IN1(n3876), .IN2(g382), .Q(n3875) );
  AND2X1 U4275 ( .IN1(n3767), .IN2(n3877), .Q(g11291) );
  OR2X1 U4276 ( .IN1(n3878), .IN2(n3879), .Q(n3877) );
  INVX0 U4277 ( .INP(n3880), .ZN(n3879) );
  OR2X1 U4278 ( .IN1(n3876), .IN2(n2433), .Q(n3880) );
  AND2X1 U4279 ( .IN1(n3881), .IN2(n3814), .Q(n3876) );
  INVX0 U4280 ( .INP(n1385), .ZN(n3881) );
  AND3X1 U4281 ( .IN1(n1385), .IN2(g374), .IN3(n3813), .Q(n3878) );
  OR3X1 U4282 ( .IN1(n2489), .IN2(n2434), .IN3(n2433), .Q(n1385) );
  AND2X1 U4283 ( .IN1(n3882), .IN2(n3767), .Q(g11290) );
  INVX0 U4284 ( .INP(n3883), .ZN(n3767) );
  OR2X1 U4285 ( .IN1(n505), .IN2(g869), .Q(n3883) );
  XOR2X1 U4286 ( .IN1(g374), .IN2(n3813), .Q(n3882) );
  AND2X1 U4287 ( .IN1(g369), .IN2(n3814), .Q(n3813) );
  AND2X1 U4288 ( .IN1(n40), .IN2(n3884), .Q(n3814) );
  OR2X1 U4289 ( .IN1(n3885), .IN2(n3886), .Q(g11270) );
  AND2X1 U4290 ( .IN1(n40), .IN2(g416), .Q(n3886) );
  AND2X1 U4291 ( .IN1(n2492), .IN2(g421), .Q(n3885) );
  OR2X1 U4292 ( .IN1(n3887), .IN2(n3888), .Q(g11269) );
  AND2X1 U4293 ( .IN1(n40), .IN2(g411), .Q(n3888) );
  AND2X1 U4294 ( .IN1(n2492), .IN2(g416), .Q(n3887) );
  OR2X1 U4295 ( .IN1(n3889), .IN2(n3890), .Q(g11268) );
  AND2X1 U4296 ( .IN1(n40), .IN2(g406), .Q(n3890) );
  AND2X1 U4297 ( .IN1(n2492), .IN2(g411), .Q(n3889) );
  OR2X1 U4298 ( .IN1(n3891), .IN2(n3892), .Q(g11267) );
  AND2X1 U4299 ( .IN1(n40), .IN2(g401), .Q(n3892) );
  AND2X1 U4300 ( .IN1(n2492), .IN2(g406), .Q(n3891) );
  OR2X1 U4301 ( .IN1(n3893), .IN2(n3894), .Q(g11266) );
  AND2X1 U4302 ( .IN1(n40), .IN2(g396), .Q(n3894) );
  AND2X1 U4303 ( .IN1(n2492), .IN2(g401), .Q(n3893) );
  OR2X1 U4304 ( .IN1(n3895), .IN2(n3896), .Q(g11265) );
  AND2X1 U4305 ( .IN1(n40), .IN2(g391), .Q(n3896) );
  AND2X1 U4306 ( .IN1(n2492), .IN2(g396), .Q(n3895) );
  OR2X1 U4307 ( .IN1(n3897), .IN2(n3898), .Q(g11264) );
  AND2X1 U4308 ( .IN1(n40), .IN2(g386), .Q(n3898) );
  AND2X1 U4309 ( .IN1(n2492), .IN2(g391), .Q(n3897) );
  OR2X1 U4310 ( .IN1(n3899), .IN2(n3900), .Q(g11263) );
  AND2X1 U4311 ( .IN1(n40), .IN2(g426), .Q(n3900) );
  AND2X1 U4312 ( .IN1(n2492), .IN2(g386), .Q(n3899) );
  OR2X1 U4313 ( .IN1(n3901), .IN2(n3902), .Q(g11262) );
  AND2X1 U4314 ( .IN1(n40), .IN2(g435), .Q(n3902) );
  AND2X1 U4315 ( .IN1(n2492), .IN2(g431), .Q(n3901) );
  OR2X1 U4316 ( .IN1(n3903), .IN2(n3904), .Q(g11261) );
  AND2X1 U4317 ( .IN1(n40), .IN2(g440), .Q(n3904) );
  AND2X1 U4318 ( .IN1(n2492), .IN2(g435), .Q(n3903) );
  OR2X1 U4319 ( .IN1(n3905), .IN2(n3906), .Q(g11260) );
  AND2X1 U4320 ( .IN1(n40), .IN2(g444), .Q(n3906) );
  AND2X1 U4321 ( .IN1(n2492), .IN2(g440), .Q(n3905) );
  OR2X1 U4322 ( .IN1(n3907), .IN2(n3908), .Q(g11259) );
  AND2X1 U4323 ( .IN1(n40), .IN2(g448), .Q(n3908) );
  AND2X1 U4324 ( .IN1(n2492), .IN2(g444), .Q(n3907) );
  OR2X1 U4325 ( .IN1(n3909), .IN2(n3910), .Q(g11258) );
  AND2X1 U4326 ( .IN1(n40), .IN2(g452), .Q(n3910) );
  AND2X1 U4327 ( .IN1(n2492), .IN2(g448), .Q(n3909) );
  OR2X1 U4328 ( .IN1(n3911), .IN2(n3912), .Q(g11257) );
  AND2X1 U4329 ( .IN1(n40), .IN2(g421), .Q(n3912) );
  AND2X1 U4330 ( .IN1(n2492), .IN2(g452), .Q(n3911) );
  OR2X1 U4331 ( .IN1(n3913), .IN2(n3914), .Q(g11256) );
  AND2X1 U4332 ( .IN1(n3766), .IN2(n40), .Q(n3914) );
  INVX0 U4333 ( .INP(n3915), .ZN(n3766) );
  OR2X1 U4334 ( .IN1(n3916), .IN2(n3917), .Q(n3915) );
  AND2X1 U4335 ( .IN1(n3918), .IN2(n1420), .Q(n3917) );
  OR2X1 U4336 ( .IN1(n3919), .IN2(n3920), .Q(n3918) );
  AND3X1 U4337 ( .IN1(n1876), .IN2(n3921), .IN3(n1878), .Q(n3920) );
  OR2X1 U4338 ( .IN1(n3922), .IN2(n3923), .Q(n3921) );
  OR4X1 U4339 ( .IN1(g411), .IN2(g426), .IN3(g391), .IN4(n3924), .Q(n3923) );
  OR3X1 U4340 ( .IN1(g386), .IN2(g401), .IN3(g421), .Q(n3924) );
  OR4X1 U4341 ( .IN1(g448), .IN2(g452), .IN3(g396), .IN4(n3925), .Q(n3922) );
  OR4X1 U4342 ( .IN1(g440), .IN2(g444), .IN3(g416), .IN4(g406), .Q(n3925) );
  AND2X1 U4343 ( .IN1(g431), .IN2(g435), .Q(n3919) );
  AND2X1 U4344 ( .IN1(n1681), .IN2(n3884), .Q(n3916) );
  INVX0 U4345 ( .INP(n1420), .ZN(n3884) );
  AND2X1 U4346 ( .IN1(n2492), .IN2(g426), .Q(n3913) );
  INVX0 U4347 ( .INP(n40), .ZN(n2492) );
  OR4X1 U4348 ( .IN1(g845), .IN2(g857), .IN3(n3926), .IN4(n3927), .Q(n40) );
  OR4X1 U4349 ( .IN1(g841), .IN2(g833), .IN3(g837), .IN4(n3928), .Q(n3927) );
  OR2X1 U4350 ( .IN1(g861), .IN2(g853), .Q(n3928) );
  OR3X1 U4351 ( .IN1(n3929), .IN2(g829), .IN3(g849), .Q(n3926) );
  AND3X1 U4352 ( .IN1(n3930), .IN2(n3931), .IN3(n3932), .Q(n3929) );
  OR2X1 U4353 ( .IN1(n505), .IN2(n3933), .Q(n3932) );
  AND2X1 U4354 ( .IN1(n3934), .IN2(n3935), .Q(n3933) );
  AND2X1 U4355 ( .IN1(g10628), .IN2(n3936), .Q(g11206) );
  XOR2X1 U4356 ( .IN1(n3936), .IN2(n2491), .Q(g11163) );
  INVX0 U4357 ( .INP(n3937), .ZN(n3936) );
  OR2X1 U4358 ( .IN1(n3938), .IN2(n3939), .Q(n3937) );
  AND2X1 U4359 ( .IN1(g5392), .IN2(g10663), .Q(n3939) );
  AND2X1 U4360 ( .IN1(g109), .IN2(n3516), .Q(g5392) );
  INVX0 U4361 ( .INP(n3515), .ZN(n3516) );
  OR2X1 U4362 ( .IN1(n2468), .IN2(n2469), .Q(n3515) );
  AND2X1 U4363 ( .IN1(n3940), .IN2(g109), .Q(n3938) );
  OR4X1 U4364 ( .IN1(n3941), .IN2(n3942), .IN3(n3943), .IN4(n3944), .Q(n3940)
         );
  AND2X1 U4365 ( .IN1(n3945), .IN2(n3036), .Q(n3944) );
  AND3X1 U4366 ( .IN1(g10724), .IN2(g3069), .IN3(n4318), .Q(n3943) );
  AND2X1 U4367 ( .IN1(n2482), .IN2(g10726), .Q(n3942) );
  AND2X1 U4368 ( .IN1(g10664), .IN2(g2648), .Q(n3941) );
  OR2X1 U4369 ( .IN1(n3946), .IN2(n3947), .Q(g10936) );
  AND2X1 U4370 ( .IN1(n1391), .IN2(n2500), .Q(n3947) );
  INVX0 U4371 ( .INP(n3948), .ZN(n1391) );
  AND4X1 U4372 ( .IN1(n3935), .IN2(n3945), .IN3(n3844), .IN4(n3649), .Q(n3948)
         );
  AND3X1 U4373 ( .IN1(n3851), .IN2(n3845), .IN3(n3846), .Q(n3935) );
  AND2X1 U4374 ( .IN1(n369), .IN2(g1811), .Q(n3946) );
  OR2X1 U4375 ( .IN1(n3949), .IN2(n3950), .Q(g10898) );
  AND2X1 U4376 ( .IN1(n3951), .IN2(n2971), .Q(n3950) );
  OR2X1 U4377 ( .IN1(n3538), .IN2(n3952), .Q(n3951) );
  XNOR3X1 U4378 ( .IN1(test_so8), .IN2(g1019), .IN3(n3953), .Q(n3952) );
  XOR3X1 U4379 ( .IN1(n3954), .IN2(n3955), .IN3(n3956), .Q(n3953) );
  XNOR3X1 U4380 ( .IN1(g1003), .IN2(n2374), .IN3(n3957), .Q(n3956) );
  XOR2X1 U4381 ( .IN1(test_so2), .IN2(n2392), .Q(n3957) );
  XOR2X1 U4382 ( .IN1(g1023), .IN2(g991), .Q(n3955) );
  XNOR2X1 U4383 ( .IN1(g1011), .IN2(n2322), .Q(n3954) );
  AND2X1 U4384 ( .IN1(n3849), .IN2(n3649), .Q(n3538) );
  OR3X1 U4385 ( .IN1(g46), .IN2(n2717), .IN3(n2719), .Q(n3649) );
  OR2X1 U4386 ( .IN1(n3958), .IN2(n2716), .Q(n2719) );
  OR4X1 U4387 ( .IN1(g44), .IN2(g43), .IN3(g48), .IN4(g45), .Q(n2716) );
  OR2X1 U4388 ( .IN1(g47), .IN2(n2721), .Q(n2717) );
  AND2X1 U4389 ( .IN1(n371), .IN2(g105), .Q(n3949) );
  OR2X1 U4390 ( .IN1(n3959), .IN2(n3960), .Q(g10866) );
  AND2X1 U4391 ( .IN1(n371), .IN2(g1684), .Q(n3959) );
  OR2X1 U4392 ( .IN1(n3961), .IN2(n3962), .Q(g10865) );
  AND3X1 U4393 ( .IN1(n1404), .IN2(n3963), .IN3(n3440), .Q(n3962) );
  OR2X1 U4394 ( .IN1(n505), .IN2(g10722), .Q(n3963) );
  AND2X1 U4395 ( .IN1(n3439), .IN2(g1669), .Q(n3961) );
  OR2X1 U4396 ( .IN1(n3964), .IN2(n3965), .Q(g10864) );
  AND2X1 U4397 ( .IN1(n371), .IN2(g1681), .Q(n3964) );
  OR2X1 U4398 ( .IN1(n3966), .IN2(n3967), .Q(g10863) );
  AND3X1 U4399 ( .IN1(n3968), .IN2(n3969), .IN3(n3440), .Q(n3967) );
  OR2X1 U4400 ( .IN1(n3970), .IN2(g1718), .Q(n3968) );
  AND2X1 U4401 ( .IN1(n3439), .IN2(g1666), .Q(n3966) );
  OR2X1 U4402 ( .IN1(n3971), .IN2(n3972), .Q(g10862) );
  AND2X1 U4403 ( .IN1(n371), .IN2(g1678), .Q(n3971) );
  OR2X1 U4404 ( .IN1(n3973), .IN2(n3974), .Q(g10861) );
  AND2X1 U4405 ( .IN1(n3975), .IN2(n3440), .Q(n3974) );
  AND2X1 U4406 ( .IN1(n3439), .IN2(g1663), .Q(n3973) );
  OR2X1 U4407 ( .IN1(n3976), .IN2(n3977), .Q(g10860) );
  AND2X1 U4408 ( .IN1(n371), .IN2(g1675), .Q(n3976) );
  OR2X1 U4409 ( .IN1(n3978), .IN2(n3979), .Q(g10859) );
  AND2X1 U4410 ( .IN1(n3980), .IN2(n3440), .Q(n3979) );
  AND2X1 U4411 ( .IN1(n3439), .IN2(g1660), .Q(n3978) );
  OR2X1 U4412 ( .IN1(n3981), .IN2(n3982), .Q(g10858) );
  AND2X1 U4413 ( .IN1(n371), .IN2(g1672), .Q(n3981) );
  OR2X1 U4414 ( .IN1(n3983), .IN2(n3984), .Q(g10855) );
  AND2X1 U4415 ( .IN1(n3975), .IN2(n2971), .Q(n3984) );
  OR2X1 U4416 ( .IN1(n3985), .IN2(n3986), .Q(n3975) );
  AND2X1 U4417 ( .IN1(n3202), .IN2(n3987), .Q(n3986) );
  OR2X1 U4418 ( .IN1(n3457), .IN2(n3988), .Q(n3202) );
  AND2X1 U4419 ( .IN1(n2985), .IN2(g1512), .Q(n3988) );
  AND2X1 U4420 ( .IN1(g18), .IN2(g192), .Q(n3457) );
  AND2X1 U4421 ( .IN1(n3989), .IN2(n3969), .Q(n3985) );
  OR2X1 U4422 ( .IN1(n3990), .IN2(g1718), .Q(n3989) );
  AND2X1 U4423 ( .IN1(g10720), .IN2(g109), .Q(n3990) );
  AND2X1 U4424 ( .IN1(n371), .IN2(g549), .Q(n3983) );
  OR2X1 U4425 ( .IN1(n2491), .IN2(n2701), .Q(g10801) );
  XOR3X1 U4426 ( .IN1(n1858), .IN2(n3991), .IN3(n3992), .Q(n2491) );
  XOR3X1 U4427 ( .IN1(n3993), .IN2(n3851), .IN3(n3994), .Q(n3992) );
  OR3X1 U4428 ( .IN1(n3995), .IN2(n3996), .IN3(n3934), .Q(n3994) );
  AND3X1 U4429 ( .IN1(n3648), .IN2(n3850), .IN3(n3849), .Q(n3934) );
  AND3X1 U4430 ( .IN1(g10664), .IN2(g10726), .IN3(n3849), .Q(n3996) );
  INVX0 U4431 ( .INP(g10663), .ZN(n3849) );
  AND2X1 U4432 ( .IN1(n3997), .IN2(g10663), .Q(n3995) );
  XOR2X1 U4433 ( .IN1(n3648), .IN2(n3850), .Q(n3997) );
  INVX0 U4434 ( .INP(g10664), .ZN(n3850) );
  INVX0 U4435 ( .INP(g10724), .ZN(n3851) );
  AND2X1 U4436 ( .IN1(n2199), .IN2(n3998), .Q(n3993) );
  XOR2X1 U4437 ( .IN1(n3845), .IN2(n3846), .Q(n3991) );
  INVX0 U4438 ( .INP(g10720), .ZN(n3845) );
  XNOR2X1 U4439 ( .IN1(n3843), .IN2(n3844), .Q(n1858) );
  OR2X1 U4440 ( .IN1(n3999), .IN2(n4000), .Q(g10800) );
  AND2X1 U4441 ( .IN1(n3980), .IN2(n2971), .Q(n4000) );
  OR2X1 U4442 ( .IN1(n4001), .IN2(n4002), .Q(n3980) );
  AND2X1 U4443 ( .IN1(n3197), .IN2(n3987), .Q(n4002) );
  OR2X1 U4444 ( .IN1(n3459), .IN2(n4003), .Q(n3197) );
  AND2X1 U4445 ( .IN1(n2985), .IN2(g1636), .Q(n4003) );
  AND2X1 U4446 ( .IN1(g18), .IN2(g248), .Q(n3459) );
  AND2X1 U4447 ( .IN1(n4004), .IN2(n3969), .Q(n4001) );
  OR2X1 U4448 ( .IN1(g10719), .IN2(n4005), .Q(n4004) );
  AND2X1 U4449 ( .IN1(n371), .IN2(g575), .Q(n3999) );
  OR2X1 U4450 ( .IN1(n4006), .IN2(n4007), .Q(g10799) );
  AND2X1 U4451 ( .IN1(n371), .IN2(g566), .Q(n4006) );
  OR2X1 U4452 ( .IN1(n4008), .IN2(n3960), .Q(g10798) );
  AND2X1 U4453 ( .IN1(n4009), .IN2(n2971), .Q(n3960) );
  OR2X1 U4454 ( .IN1(n4010), .IN2(n4011), .Q(n4009) );
  AND2X1 U4455 ( .IN1(n1404), .IN2(n3872), .Q(n4011) );
  AND2X1 U4456 ( .IN1(n3987), .IN2(n3200), .Q(n4010) );
  OR2X1 U4457 ( .IN1(n4012), .IN2(n2993), .Q(n3200) );
  INVX0 U4458 ( .INP(n4013), .ZN(n2993) );
  OR2X1 U4459 ( .IN1(n2457), .IN2(n2985), .Q(n4013) );
  AND2X1 U4460 ( .IN1(n2985), .IN2(g1624), .Q(n4012) );
  AND2X1 U4461 ( .IN1(n371), .IN2(g563), .Q(n4008) );
  OR2X1 U4462 ( .IN1(n4014), .IN2(n3965), .Q(g10797) );
  AND2X1 U4463 ( .IN1(n4015), .IN2(n2971), .Q(n3965) );
  OR2X1 U4464 ( .IN1(n4016), .IN2(n4017), .Q(n4015) );
  AND2X1 U4465 ( .IN1(n1404), .IN2(n3945), .Q(n4017) );
  AND2X1 U4466 ( .IN1(n3987), .IN2(n3195), .Q(n4016) );
  OR2X1 U4467 ( .IN1(n4018), .IN2(n2983), .Q(n3195) );
  INVX0 U4468 ( .INP(n4019), .ZN(n2983) );
  OR2X1 U4469 ( .IN1(n2460), .IN2(n2985), .Q(n4019) );
  AND2X1 U4470 ( .IN1(n2985), .IN2(g1621), .Q(n4018) );
  AND2X1 U4471 ( .IN1(n371), .IN2(g560), .Q(n4014) );
  OR2X1 U4472 ( .IN1(n4020), .IN2(n3972), .Q(g10795) );
  AND2X1 U4473 ( .IN1(n4021), .IN2(n2971), .Q(n3972) );
  OR2X1 U4474 ( .IN1(n4022), .IN2(n4023), .Q(n4021) );
  AND2X1 U4475 ( .IN1(n1404), .IN2(n3970), .Q(n4023) );
  AND2X1 U4476 ( .IN1(n3987), .IN2(n3187), .Q(n4022) );
  OR2X1 U4477 ( .IN1(n4024), .IN2(n3068), .Q(n3187) );
  AND2X1 U4478 ( .IN1(g213), .IN2(g18), .Q(n3068) );
  AND2X1 U4479 ( .IN1(n2985), .IN2(g1615), .Q(n4024) );
  AND2X1 U4480 ( .IN1(n371), .IN2(g557), .Q(n4020) );
  OR2X1 U4481 ( .IN1(n4025), .IN2(n3977), .Q(g10793) );
  AND3X1 U4482 ( .IN1(n4026), .IN2(n4027), .IN3(n2971), .Q(n3977) );
  OR2X1 U4483 ( .IN1(n3183), .IN2(n3969), .Q(n4027) );
  OR2X1 U4484 ( .IN1(n4028), .IN2(n3021), .Q(n3183) );
  INVX0 U4485 ( .INP(n4029), .ZN(n3021) );
  OR2X1 U4486 ( .IN1(n2458), .IN2(n2985), .Q(n4029) );
  AND2X1 U4487 ( .IN1(n2985), .IN2(g1639), .Q(n4028) );
  OR3X1 U4488 ( .IN1(n4005), .IN2(g10720), .IN3(n3987), .Q(n4026) );
  OR2X1 U4489 ( .IN1(n505), .IN2(g1718), .Q(n4005) );
  AND2X1 U4490 ( .IN1(n371), .IN2(g554), .Q(n4025) );
  OR2X1 U4491 ( .IN1(n4030), .IN2(n3982), .Q(g10791) );
  INVX0 U4492 ( .INP(n4031), .ZN(n3982) );
  OR2X1 U4493 ( .IN1(n371), .IN2(n4032), .Q(n4031) );
  AND2X1 U4494 ( .IN1(n4033), .IN2(n4034), .Q(n4032) );
  OR3X1 U4495 ( .IN1(n505), .IN2(n3846), .IN3(n4035), .Q(n4034) );
  INVX0 U4496 ( .INP(g10719), .ZN(n3846) );
  OR2X1 U4497 ( .IN1(n4036), .IN2(n3969), .Q(n4033) );
  INVX0 U4498 ( .INP(n3204), .ZN(n4036) );
  OR2X1 U4499 ( .IN1(n4037), .IN2(n3004), .Q(n3204) );
  AND2X1 U4500 ( .IN1(g186), .IN2(g18), .Q(n3004) );
  AND2X1 U4501 ( .IN1(n2985), .IN2(g1618), .Q(n4037) );
  AND2X1 U4502 ( .IN1(n371), .IN2(g546), .Q(n4030) );
  AND2X1 U4503 ( .IN1(n369), .IN2(n3023), .Q(g10785) );
  AND2X1 U4504 ( .IN1(n369), .IN2(n3029), .Q(g10784) );
  AND2X1 U4505 ( .IN1(n369), .IN2(n3065), .Q(g10782) );
  AND2X1 U4506 ( .IN1(n369), .IN2(n3017), .Q(g10780) );
  INVX0 U4507 ( .INP(n2500), .ZN(n369) );
  AND2X1 U4508 ( .IN1(n2406), .IN2(g1696), .Q(n2500) );
  OR2X1 U4509 ( .IN1(n4038), .IN2(n4007), .Q(g10776) );
  INVX0 U4510 ( .INP(n4039), .ZN(n4007) );
  OR2X1 U4511 ( .IN1(n371), .IN2(n4040), .Q(n4039) );
  AND3X1 U4512 ( .IN1(n4041), .IN2(n4042), .IN3(n4043), .Q(n4040) );
  OR2X1 U4513 ( .IN1(n3648), .IN2(n4035), .Q(n4043) );
  INVX0 U4514 ( .INP(g10726), .ZN(n3648) );
  INVX0 U4515 ( .INP(n1450), .ZN(n4042) );
  OR2X1 U4516 ( .IN1(n4044), .IN2(n3969), .Q(n4041) );
  INVX0 U4517 ( .INP(n3206), .ZN(n4044) );
  OR2X1 U4518 ( .IN1(n4045), .IN2(n3010), .Q(n3206) );
  INVX0 U4519 ( .INP(n4046), .ZN(n3010) );
  OR2X1 U4520 ( .IN1(n2459), .IN2(n2985), .Q(n4046) );
  AND2X1 U4521 ( .IN1(n2985), .IN2(g1627), .Q(n4045) );
  AND2X1 U4522 ( .IN1(n371), .IN2(g1687), .Q(n4038) );
  OR2X1 U4523 ( .IN1(n4047), .IN2(n4048), .Q(g10773) );
  AND2X1 U4524 ( .IN1(n3509), .IN2(g1727), .Q(n4048) );
  AND2X1 U4525 ( .IN1(n4049), .IN2(n3970), .Q(n4047) );
  INVX0 U4526 ( .INP(n3930), .ZN(n3970) );
  OR2X1 U4527 ( .IN1(n4050), .IN2(n4051), .Q(g10771) );
  AND3X1 U4528 ( .IN1(g109), .IN2(g10720), .IN3(n4049), .Q(n4051) );
  AND2X1 U4529 ( .IN1(n3509), .IN2(g1724), .Q(n4050) );
  OR2X1 U4530 ( .IN1(n4052), .IN2(n4053), .Q(g10770) );
  AND3X1 U4531 ( .IN1(g109), .IN2(g10719), .IN3(n4049), .Q(n4053) );
  AND2X1 U4532 ( .IN1(n3509), .IN2(g1721), .Q(n4052) );
  OR2X1 U4533 ( .IN1(n4054), .IN2(n4055), .Q(g10767) );
  AND2X1 U4534 ( .IN1(n4056), .IN2(n3440), .Q(n4055) );
  AND2X1 U4535 ( .IN1(n3439), .IN2(g1657), .Q(n4054) );
  OR2X1 U4536 ( .IN1(n4057), .IN2(n4058), .Q(g10765) );
  AND2X1 U4537 ( .IN1(n3440), .IN2(n4059), .Q(n4058) );
  INVX0 U4538 ( .INP(n3439), .ZN(n3440) );
  AND2X1 U4539 ( .IN1(n3439), .IN2(g1654), .Q(n4057) );
  OR2X1 U4540 ( .IN1(g1696), .IN2(n2406), .Q(n3439) );
  OR2X1 U4541 ( .IN1(n4060), .IN2(n4061), .Q(g10718) );
  AND2X1 U4542 ( .IN1(n4056), .IN2(n2971), .Q(n4061) );
  OR2X1 U4543 ( .IN1(n4062), .IN2(n4063), .Q(n4056) );
  AND2X1 U4544 ( .IN1(n3189), .IN2(n3987), .Q(n4063) );
  OR2X1 U4545 ( .IN1(n3461), .IN2(n4064), .Q(n3189) );
  AND2X1 U4546 ( .IN1(n2985), .IN2(g1633), .Q(n4064) );
  AND2X1 U4547 ( .IN1(g18), .IN2(g243), .Q(n3461) );
  AND2X1 U4548 ( .IN1(n4065), .IN2(n3969), .Q(n4062) );
  INVX0 U4549 ( .INP(n3987), .ZN(n3969) );
  OR2X1 U4550 ( .IN1(n4066), .IN2(g1718), .Q(n4065) );
  AND2X1 U4551 ( .IN1(g10664), .IN2(g109), .Q(n4066) );
  AND2X1 U4552 ( .IN1(n371), .IN2(g572), .Q(n4060) );
  OR2X1 U4553 ( .IN1(n4067), .IN2(n4068), .Q(g10717) );
  AND2X1 U4554 ( .IN1(n4059), .IN2(n2971), .Q(n4068) );
  OR3X1 U4555 ( .IN1(n1450), .IN2(n4069), .IN3(n4070), .Q(n4059) );
  AND2X1 U4556 ( .IN1(n1404), .IN2(g10663), .Q(n4070) );
  INVX0 U4557 ( .INP(n4035), .ZN(n1404) );
  OR2X1 U4558 ( .IN1(n3987), .IN2(g1718), .Q(n4035) );
  AND2X1 U4559 ( .IN1(n3987), .IN2(n3208), .Q(n4069) );
  OR2X1 U4560 ( .IN1(n4071), .IN2(n3052), .Q(n3208) );
  AND2X1 U4561 ( .IN1(g237), .IN2(g18), .Q(n3052) );
  AND2X1 U4562 ( .IN1(n2985), .IN2(g1630), .Q(n4071) );
  INVX0 U4563 ( .INP(g18), .ZN(n2985) );
  AND2X1 U4564 ( .IN1(n1611), .IN2(n4323), .Q(n3987) );
  AND2X1 U4565 ( .IN1(n371), .IN2(g569), .Q(n4067) );
  INVX0 U4566 ( .INP(n2971), .ZN(n371) );
  AND2X1 U4567 ( .IN1(n3340), .IN2(n2406), .Q(n2971) );
  OR2X1 U4568 ( .IN1(n4072), .IN2(n4073), .Q(g10711) );
  AND2X1 U4569 ( .IN1(n4049), .IN2(n3872), .Q(n4073) );
  OR2X1 U4570 ( .IN1(n505), .IN2(g10724), .Q(n3872) );
  AND2X1 U4571 ( .IN1(n3509), .IN2(g1733), .Q(n4072) );
  OR2X1 U4572 ( .IN1(n4074), .IN2(n4075), .Q(g10707) );
  AND2X1 U4573 ( .IN1(n3509), .IN2(g1730), .Q(n4075) );
  AND2X1 U4574 ( .IN1(n4049), .IN2(n3945), .Q(n4074) );
  INVX0 U4575 ( .INP(n3509), .ZN(n4049) );
  OR2X1 U4576 ( .IN1(n2406), .IN2(n3340), .Q(n3509) );
  INVX0 U4577 ( .INP(g1696), .ZN(n3340) );
  OR4X1 U4578 ( .IN1(n4076), .IN2(n4077), .IN3(n4078), .IN4(n4079), .Q(g10664)
         );
  OR4X1 U4579 ( .IN1(n4080), .IN2(n4081), .IN3(n4082), .IN4(n4083), .Q(n4079)
         );
  OR2X1 U4580 ( .IN1(n4084), .IN2(n4085), .Q(n4083) );
  AND2X1 U4581 ( .IN1(n4086), .IN2(g1741), .Q(n4085) );
  AND2X1 U4582 ( .IN1(n1486), .IN2(g1546), .Q(n4084) );
  AND2X1 U4583 ( .IN1(test_so9), .IN2(n4087), .Q(n4082) );
  AND2X1 U4584 ( .IN1(g1191), .IN2(n4088), .Q(n4081) );
  INVX0 U4585 ( .INP(n4089), .ZN(n4080) );
  OR4X1 U4586 ( .IN1(n4090), .IN2(n4091), .IN3(n4092), .IN4(n4088), .Q(n4089)
         );
  OR2X1 U4587 ( .IN1(n4087), .IN2(n4086), .Q(n4092) );
  INVX0 U4588 ( .INP(n1478), .ZN(n4090) );
  OR3X1 U4589 ( .IN1(n4093), .IN2(n4094), .IN3(n4095), .Q(n4078) );
  AND2X1 U4590 ( .IN1(n4096), .IN2(g284), .Q(n4095) );
  AND2X1 U4591 ( .IN1(n4097), .IN2(g947), .Q(n4094) );
  AND2X1 U4592 ( .IN1(g919), .IN2(n4098), .Q(n4093) );
  AND2X1 U4593 ( .IN1(n1485), .IN2(g1589), .Q(n4077) );
  AND2X1 U4594 ( .IN1(n3998), .IN2(n3040), .Q(n4076) );
  AND2X1 U4595 ( .IN1(n4099), .IN2(n4100), .Q(g10628) );
  OR2X1 U4596 ( .IN1(n3930), .IN2(n3179), .Q(n4100) );
  OR3X1 U4597 ( .IN1(n2476), .IN2(n505), .IN3(n3058), .Q(n3179) );
  OR2X1 U4598 ( .IN1(n505), .IN2(n3844), .Q(n3930) );
  INVX0 U4599 ( .INP(g10721), .ZN(n3844) );
  OR2X1 U4600 ( .IN1(n4101), .IN2(n505), .Q(n4099) );
  INVX0 U4601 ( .INP(n4102), .ZN(n4101) );
  OR4X1 U4602 ( .IN1(n4103), .IN2(n4104), .IN3(n4105), .IN4(n4106), .Q(n4102)
         );
  AND2X1 U4603 ( .IN1(n3064), .IN2(n3945), .Q(n4106) );
  INVX0 U4604 ( .INP(n3931), .ZN(n3945) );
  OR2X1 U4605 ( .IN1(n505), .IN2(n3843), .Q(n3931) );
  INVX0 U4606 ( .INP(g10722), .ZN(n3843) );
  OR4X1 U4607 ( .IN1(n4107), .IN2(n4108), .IN3(n4109), .IN4(n4110), .Q(g10722)
         );
  OR4X1 U4608 ( .IN1(n4111), .IN2(n4112), .IN3(n4113), .IN4(n4114), .Q(n4110)
         );
  OR2X1 U4609 ( .IN1(n4115), .IN2(n4116), .Q(n4114) );
  AND2X1 U4610 ( .IN1(n4097), .IN2(g986), .Q(n4116) );
  AND2X1 U4611 ( .IN1(g907), .IN2(n4098), .Q(n4115) );
  AND2X1 U4612 ( .IN1(n4087), .IN2(g1351), .Q(n4113) );
  AND2X1 U4613 ( .IN1(g1179), .IN2(n4088), .Q(n4112) );
  AND2X1 U4614 ( .IN1(n4117), .IN2(g1324), .Q(n4111) );
  OR4X1 U4615 ( .IN1(n4118), .IN2(n4119), .IN3(n4120), .IN4(n4121), .Q(n4109)
         );
  OR3X1 U4616 ( .IN1(n4122), .IN2(n4123), .IN3(n4124), .Q(n4121) );
  AND2X1 U4617 ( .IN1(n4125), .IN2(g8), .Q(n4124) );
  AND2X1 U4618 ( .IN1(n4126), .IN2(n1631), .Q(n4123) );
  AND2X1 U4619 ( .IN1(n2700), .IN2(g959), .Q(n4122) );
  AND2X1 U4620 ( .IN1(n4127), .IN2(g940), .Q(n4120) );
  AND2X1 U4621 ( .IN1(g895), .IN2(n4128), .Q(n4119) );
  OR4X1 U4622 ( .IN1(n4129), .IN2(n4130), .IN3(n4131), .IN4(n4132), .Q(n4108)
         );
  OR2X1 U4623 ( .IN1(n4133), .IN2(n4134), .Q(n4132) );
  AND2X1 U4624 ( .IN1(n1486), .IN2(g1534), .Q(n4134) );
  AND2X1 U4625 ( .IN1(n1485), .IN2(g1577), .Q(n4133) );
  AND2X1 U4626 ( .IN1(n1479), .IN2(g1558), .Q(n4131) );
  AND2X1 U4627 ( .IN1(n1512), .IN2(g1203), .Q(n4130) );
  AND2X1 U4628 ( .IN1(n1480), .IN2(g1601), .Q(n4129) );
  OR4X1 U4629 ( .IN1(n4135), .IN2(n4136), .IN3(n4137), .IN4(n4138), .Q(n4107)
         );
  OR2X1 U4630 ( .IN1(n4139), .IN2(n4140), .Q(n4138) );
  AND2X1 U4631 ( .IN1(n3998), .IN2(n3048), .Q(n4140) );
  AND2X1 U4632 ( .IN1(n4086), .IN2(g1730), .Q(n4139) );
  AND2X1 U4633 ( .IN1(n4141), .IN2(g296), .Q(n4137) );
  AND2X1 U4634 ( .IN1(n4096), .IN2(g272), .Q(n4136) );
  AND2X1 U4635 ( .IN1(n4142), .IN2(g1753), .Q(n4135) );
  INVX0 U4636 ( .INP(g109), .ZN(n505) );
  AND3X1 U4637 ( .IN1(g10724), .IN2(g3007), .IN3(n4317), .Q(n4105) );
  AND2X1 U4638 ( .IN1(g881), .IN2(g10720), .Q(n4104) );
  AND2X1 U4639 ( .IN1(g877), .IN2(g10719), .Q(n4103) );
  OR2X1 U4640 ( .IN1(g10726), .IN2(n2701), .Q(g10465) );
  OR4X1 U4641 ( .IN1(n4143), .IN2(n4144), .IN3(n4145), .IN4(n4146), .Q(g10726)
         );
  OR4X1 U4642 ( .IN1(n4147), .IN2(n4148), .IN3(n4149), .IN4(n4150), .Q(n4146)
         );
  OR3X1 U4643 ( .IN1(n4151), .IN2(n4152), .IN3(n4153), .Q(n4150) );
  AND2X1 U4644 ( .IN1(n1486), .IN2(g1540), .Q(n4153) );
  AND2X1 U4645 ( .IN1(n1485), .IN2(g1583), .Q(n4152) );
  AND2X1 U4646 ( .IN1(n1479), .IN2(g1564), .Q(n4151) );
  AND2X1 U4647 ( .IN1(n1480), .IN2(g1607), .Q(n4149) );
  AND2X1 U4648 ( .IN1(n3998), .IN2(n1650), .Q(n4148) );
  AND2X1 U4649 ( .IN1(n4141), .IN2(g302), .Q(n4147) );
  OR4X1 U4650 ( .IN1(n4154), .IN2(n4155), .IN3(n4156), .IN4(n4157), .Q(n4145)
         );
  AND2X1 U4651 ( .IN1(n2700), .IN2(g965), .Q(n4157) );
  AND2X1 U4652 ( .IN1(n1478), .IN2(n4158), .Q(n4156) );
  AND2X1 U4653 ( .IN1(n4117), .IN2(g1330), .Q(n4155) );
  AND2X1 U4654 ( .IN1(g913), .IN2(n4098), .Q(n4154) );
  OR2X1 U4655 ( .IN1(n4159), .IN2(n4160), .Q(n4144) );
  AND2X1 U4656 ( .IN1(n4142), .IN2(g1759), .Q(n4160) );
  AND2X1 U4657 ( .IN1(g1185), .IN2(n4088), .Q(n4159) );
  AND2X1 U4658 ( .IN1(n4096), .IN2(g278), .Q(n4143) );
  OR2X1 U4659 ( .IN1(g10724), .IN2(n2701), .Q(g10463) );
  OR4X1 U4660 ( .IN1(n4161), .IN2(n4162), .IN3(n4163), .IN4(n4164), .Q(g10724)
         );
  OR4X1 U4661 ( .IN1(n4165), .IN2(n4166), .IN3(n4167), .IN4(n4168), .Q(n4164)
         );
  AND2X1 U4662 ( .IN1(n4142), .IN2(g1756), .Q(n4168) );
  AND2X1 U4663 ( .IN1(g1182), .IN2(n4088), .Q(n4167) );
  AND2X1 U4664 ( .IN1(n4141), .IN2(g299), .Q(n4166) );
  AND2X1 U4665 ( .IN1(n4096), .IN2(g275), .Q(n4165) );
  OR4X1 U4666 ( .IN1(n4169), .IN2(n4170), .IN3(n4171), .IN4(n4172), .Q(n4163)
         );
  AND2X1 U4667 ( .IN1(n4125), .IN2(n3025), .Q(n4172) );
  AND2X1 U4668 ( .IN1(n2700), .IN2(g962), .Q(n4171) );
  AND2X1 U4669 ( .IN1(n4117), .IN2(g1327), .Q(n4170) );
  AND2X1 U4670 ( .IN1(g910), .IN2(n4098), .Q(n4169) );
  OR4X1 U4671 ( .IN1(n4173), .IN2(n4174), .IN3(n4175), .IN4(n4176), .Q(n4162)
         );
  INVX0 U4672 ( .INP(n4177), .ZN(n4176) );
  OR2X1 U4673 ( .IN1(n4178), .IN2(n4126), .Q(n4177) );
  AND2X1 U4674 ( .IN1(n4126), .IN2(n3057), .Q(n4175) );
  AND2X1 U4675 ( .IN1(n1486), .IN2(g1537), .Q(n4174) );
  AND2X1 U4676 ( .IN1(n1485), .IN2(g1580), .Q(n4173) );
  OR4X1 U4677 ( .IN1(n4179), .IN2(n4180), .IN3(n4181), .IN4(n4182), .Q(n4161)
         );
  AND2X1 U4678 ( .IN1(n3998), .IN2(n3034), .Q(n4182) );
  AND2X1 U4679 ( .IN1(n4086), .IN2(g1733), .Q(n4181) );
  AND2X1 U4680 ( .IN1(n1479), .IN2(g1561), .Q(n4180) );
  AND2X1 U4681 ( .IN1(n1480), .IN2(g1604), .Q(n4179) );
  OR2X1 U4682 ( .IN1(g10721), .IN2(n2701), .Q(g10459) );
  OR4X1 U4683 ( .IN1(n4183), .IN2(n4184), .IN3(n4185), .IN4(n4186), .Q(g10721)
         );
  OR4X1 U4684 ( .IN1(n4187), .IN2(n4188), .IN3(n4189), .IN4(n4190), .Q(n4186)
         );
  OR2X1 U4685 ( .IN1(n4191), .IN2(n4192), .Q(n4190) );
  AND2X1 U4686 ( .IN1(n4097), .IN2(g981), .Q(n4192) );
  AND2X1 U4687 ( .IN1(g904), .IN2(n4098), .Q(n4191) );
  AND2X1 U4688 ( .IN1(n4087), .IN2(g1346), .Q(n4189) );
  AND2X1 U4689 ( .IN1(g1176), .IN2(n4088), .Q(n4188) );
  AND2X1 U4690 ( .IN1(n4117), .IN2(g1321), .Q(n4187) );
  OR4X1 U4691 ( .IN1(n4118), .IN2(n4193), .IN3(n4194), .IN4(n4195), .Q(n4185)
         );
  OR3X1 U4692 ( .IN1(n4196), .IN2(n4197), .IN3(n4198), .Q(n4195) );
  AND2X1 U4693 ( .IN1(n4125), .IN2(g1), .Q(n4198) );
  AND2X1 U4694 ( .IN1(n4126), .IN2(g9), .Q(n4197) );
  AND2X1 U4695 ( .IN1(n2700), .IN2(g956), .Q(n4196) );
  AND2X1 U4696 ( .IN1(n4127), .IN2(g936), .Q(n4194) );
  AND2X1 U4697 ( .IN1(g892), .IN2(n4128), .Q(n4193) );
  OR4X1 U4698 ( .IN1(n4199), .IN2(n4200), .IN3(n4201), .IN4(n4202), .Q(n4184)
         );
  OR2X1 U4699 ( .IN1(n4203), .IN2(n4204), .Q(n4202) );
  AND2X1 U4700 ( .IN1(n1486), .IN2(g1531), .Q(n4204) );
  AND2X1 U4701 ( .IN1(n1485), .IN2(g1574), .Q(n4203) );
  AND2X1 U4702 ( .IN1(n1479), .IN2(g1555), .Q(n4201) );
  AND2X1 U4703 ( .IN1(g1200), .IN2(n1512), .Q(n4200) );
  AND2X1 U4704 ( .IN1(n1480), .IN2(g1598), .Q(n4199) );
  OR4X1 U4705 ( .IN1(n4205), .IN2(n4206), .IN3(n4207), .IN4(n4208), .Q(n4183)
         );
  OR2X1 U4706 ( .IN1(n4209), .IN2(n4210), .Q(n4208) );
  AND2X1 U4707 ( .IN1(n3998), .IN2(n3045), .Q(n4210) );
  AND2X1 U4708 ( .IN1(n4086), .IN2(g1727), .Q(n4209) );
  AND2X1 U4709 ( .IN1(n4141), .IN2(g293), .Q(n4207) );
  AND2X1 U4710 ( .IN1(n4096), .IN2(g269), .Q(n4206) );
  AND2X1 U4711 ( .IN1(n4142), .IN2(g1750), .Q(n4205) );
  OR2X1 U4712 ( .IN1(g10720), .IN2(n2701), .Q(g10457) );
  OR4X1 U4713 ( .IN1(n4211), .IN2(n4212), .IN3(n4213), .IN4(n4214), .Q(g10720)
         );
  OR4X1 U4714 ( .IN1(n4215), .IN2(n4216), .IN3(n4217), .IN4(n4218), .Q(n4214)
         );
  OR2X1 U4715 ( .IN1(n4219), .IN2(n4220), .Q(n4218) );
  AND2X1 U4716 ( .IN1(n4097), .IN2(g976), .Q(n4220) );
  AND2X1 U4717 ( .IN1(g901), .IN2(n4098), .Q(n4219) );
  AND2X1 U4718 ( .IN1(n4087), .IN2(g1341), .Q(n4217) );
  AND2X1 U4719 ( .IN1(g1173), .IN2(n4088), .Q(n4216) );
  AND2X1 U4720 ( .IN1(n4117), .IN2(g1318), .Q(n4215) );
  OR4X1 U4721 ( .IN1(n4118), .IN2(n4221), .IN3(n4222), .IN4(n4223), .Q(n4213)
         );
  OR3X1 U4722 ( .IN1(n4224), .IN2(n4225), .IN3(n4226), .Q(n4223) );
  AND2X1 U4723 ( .IN1(n4125), .IN2(g4), .Q(n4226) );
  AND2X1 U4724 ( .IN1(n4126), .IN2(g12), .Q(n4225) );
  AND2X1 U4725 ( .IN1(n2700), .IN2(g953), .Q(n4224) );
  AND2X1 U4726 ( .IN1(n4127), .IN2(g932), .Q(n4222) );
  AND2X1 U4727 ( .IN1(g889), .IN2(n4128), .Q(n4221) );
  OR4X1 U4728 ( .IN1(n4227), .IN2(n4228), .IN3(n4229), .IN4(n4230), .Q(n4212)
         );
  OR2X1 U4729 ( .IN1(n4231), .IN2(n4232), .Q(n4230) );
  AND2X1 U4730 ( .IN1(n1530), .IN2(g925), .Q(n4232) );
  AND2X1 U4731 ( .IN1(g1197), .IN2(n1512), .Q(n4231) );
  AND2X1 U4732 ( .IN1(n1479), .IN2(g1552), .Q(n4229) );
  AND2X1 U4733 ( .IN1(n1486), .IN2(g1528), .Q(n4228) );
  AND2X1 U4734 ( .IN1(n1485), .IN2(g1571), .Q(n4227) );
  OR4X1 U4735 ( .IN1(n4233), .IN2(n4234), .IN3(n4235), .IN4(n4236), .Q(n4211)
         );
  OR3X1 U4736 ( .IN1(n4237), .IN2(n4238), .IN3(n4239), .Q(n4236) );
  AND2X1 U4737 ( .IN1(n1480), .IN2(g1595), .Q(n4239) );
  AND2X1 U4738 ( .IN1(n3998), .IN2(n3031), .Q(n4238) );
  AND2X1 U4739 ( .IN1(n4086), .IN2(g1724), .Q(n4237) );
  AND2X1 U4740 ( .IN1(n4141), .IN2(g290), .Q(n4235) );
  AND2X1 U4741 ( .IN1(n4096), .IN2(g266), .Q(n4234) );
  AND2X1 U4742 ( .IN1(n4142), .IN2(g1747), .Q(n4233) );
  OR2X1 U4743 ( .IN1(g10719), .IN2(n2701), .Q(g10455) );
  OR4X1 U4744 ( .IN1(n4240), .IN2(n4241), .IN3(n4242), .IN4(n4243), .Q(g10719)
         );
  OR4X1 U4745 ( .IN1(n4244), .IN2(n4245), .IN3(n4246), .IN4(n4247), .Q(n4243)
         );
  OR3X1 U4746 ( .IN1(n4248), .IN2(n4249), .IN3(n4250), .Q(n4247) );
  AND2X1 U4747 ( .IN1(g1170), .IN2(n4088), .Q(n4250) );
  AND2X1 U4748 ( .IN1(n4117), .IN2(g1314), .Q(n4249) );
  AND2X1 U4749 ( .IN1(n4087), .IN2(g1336), .Q(n4248) );
  AND2X1 U4750 ( .IN1(n4097), .IN2(g971), .Q(n4246) );
  AND2X1 U4751 ( .IN1(g898), .IN2(n4098), .Q(n4245) );
  AND2X1 U4752 ( .IN1(n4125), .IN2(g123), .Q(n4244) );
  OR4X1 U4753 ( .IN1(n2501), .IN2(n4118), .IN3(n4251), .IN4(n4252), .Q(n4242)
         );
  OR3X1 U4754 ( .IN1(n4253), .IN2(n4254), .IN3(n4255), .Q(n4252) );
  AND2X1 U4755 ( .IN1(n4126), .IN2(g119), .Q(n4255) );
  AND2X1 U4756 ( .IN1(n2700), .IN2(g950), .Q(n4254) );
  AND2X1 U4757 ( .IN1(n4127), .IN2(g928), .Q(n4253) );
  AND2X1 U4758 ( .IN1(g886), .IN2(n4128), .Q(n4251) );
  INVX0 U4759 ( .INP(n4256), .ZN(n4118) );
  OR4X1 U4760 ( .IN1(n4126), .IN2(n4178), .IN3(n1512), .IN4(n4087), .Q(n4256)
         );
  OR4X1 U4761 ( .IN1(n4257), .IN2(n2702), .IN3(n2501), .IN4(n4125), .Q(n4178)
         );
  AND2X1 U4762 ( .IN1(g42), .IN2(n4258), .Q(n4125) );
  OR2X1 U4763 ( .IN1(n4259), .IN2(n4260), .Q(n2702) );
  OR4X1 U4764 ( .IN1(n4261), .IN2(n3998), .IN3(n4127), .IN4(n4128), .Q(n4260)
         );
  AND4X1 U4765 ( .IN1(n1574), .IN2(n4262), .IN3(g43), .IN4(g42), .Q(n4128) );
  AND4X1 U4766 ( .IN1(n1574), .IN2(g45), .IN3(g42), .IN4(n4263), .Q(n4127) );
  AND2X1 U4767 ( .IN1(n4264), .IN2(g44), .Q(n4263) );
  OR4X1 U4768 ( .IN1(n4098), .IN2(n2700), .IN3(n1530), .IN4(n4097), .Q(n4259)
         );
  AND2X1 U4769 ( .IN1(n1574), .IN2(n4265), .Q(n2700) );
  AND2X1 U4770 ( .IN1(n3958), .IN2(n4258), .Q(n4126) );
  AND4X1 U4771 ( .IN1(g43), .IN2(n1548), .IN3(n4266), .IN4(n4267), .Q(n4258)
         );
  OR4X1 U4772 ( .IN1(n4268), .IN2(n4269), .IN3(n4270), .IN4(n4271), .Q(n4241)
         );
  OR2X1 U4773 ( .IN1(n4272), .IN2(n4273), .Q(n4271) );
  AND2X1 U4774 ( .IN1(g922), .IN2(n1530), .Q(n4273) );
  AND2X1 U4775 ( .IN1(g1194), .IN2(n1512), .Q(n4272) );
  AND2X1 U4776 ( .IN1(n1479), .IN2(g1549), .Q(n4270) );
  AND2X1 U4777 ( .IN1(n1486), .IN2(g1524), .Q(n4269) );
  AND2X1 U4778 ( .IN1(n1485), .IN2(g1567), .Q(n4268) );
  OR4X1 U4779 ( .IN1(n4274), .IN2(n4275), .IN3(n4276), .IN4(n4277), .Q(n4240)
         );
  OR3X1 U4780 ( .IN1(n4278), .IN2(n4279), .IN3(n4280), .Q(n4277) );
  AND2X1 U4781 ( .IN1(n1480), .IN2(g1592), .Q(n4280) );
  AND2X1 U4782 ( .IN1(n3998), .IN2(n3051), .Q(n4279) );
  AND2X1 U4783 ( .IN1(n4086), .IN2(g1721), .Q(n4278) );
  AND2X1 U4784 ( .IN1(n4141), .IN2(g287), .Q(n4276) );
  AND2X1 U4785 ( .IN1(n4096), .IN2(g263), .Q(n4275) );
  AND2X1 U4786 ( .IN1(n4142), .IN2(g1744), .Q(n4274) );
  OR2X1 U4787 ( .IN1(g10663), .IN2(n2701), .Q(g10377) );
  OR2X1 U4788 ( .IN1(g30), .IN2(n3998), .Q(n2701) );
  OR4X1 U4789 ( .IN1(n4281), .IN2(n4282), .IN3(n4283), .IN4(n4284), .Q(g10663)
         );
  OR4X1 U4790 ( .IN1(n4285), .IN2(n4286), .IN3(n4287), .IN4(n4288), .Q(n4284)
         );
  OR4X1 U4791 ( .IN1(n4289), .IN2(n4290), .IN3(n1564), .IN4(n2501), .Q(n4288)
         );
  AND4X1 U4792 ( .IN1(g46), .IN2(g47), .IN3(n4291), .IN4(n4292), .Q(n2501) );
  INVX0 U4793 ( .INP(n1545), .ZN(n4291) );
  OR4X1 U4794 ( .IN1(n4264), .IN2(n4267), .IN3(g45), .IN4(g42), .Q(n1545) );
  AND2X1 U4795 ( .IN1(n4097), .IN2(g944), .Q(n4290) );
  AND2X1 U4796 ( .IN1(n1574), .IN2(n4293), .Q(n4097) );
  AND2X1 U4797 ( .IN1(g916), .IN2(n4098), .Q(n4289) );
  AND2X1 U4798 ( .IN1(n4294), .IN2(n1574), .Q(n4098) );
  AND3X1 U4799 ( .IN1(n2722), .IN2(n4292), .IN3(g46), .Q(n1574) );
  AND2X1 U4800 ( .IN1(n4142), .IN2(g1762), .Q(n4287) );
  AND2X1 U4801 ( .IN1(g1188), .IN2(n4088), .Q(n4286) );
  AND2X1 U4802 ( .IN1(n4117), .IN2(g1333), .Q(n4285) );
  OR4X1 U4803 ( .IN1(n4295), .IN2(n4296), .IN3(n4297), .IN4(n4298), .Q(n4283)
         );
  AND3X1 U4804 ( .IN1(n1478), .IN2(n4158), .IN3(n4299), .Q(n4298) );
  INVX0 U4805 ( .INP(n4087), .ZN(n4299) );
  INVX0 U4806 ( .INP(n4257), .ZN(n4158) );
  OR4X1 U4807 ( .IN1(n4117), .IN2(n4091), .IN3(n4088), .IN4(n4300), .Q(n4257)
         );
  OR2X1 U4808 ( .IN1(n4086), .IN2(n4142), .Q(n4300) );
  AND2X1 U4809 ( .IN1(n3958), .IN2(n4301), .Q(n4142) );
  AND2X1 U4810 ( .IN1(n4294), .IN2(n1544), .Q(n4088) );
  OR2X1 U4811 ( .IN1(n1567), .IN2(n1566), .Q(n4091) );
  OR2X1 U4812 ( .IN1(n4302), .IN2(n1479), .Q(n1566) );
  AND2X1 U4813 ( .IN1(n1548), .IN2(n4294), .Q(n4302) );
  AND4X1 U4814 ( .IN1(g44), .IN2(g42), .IN3(n4266), .IN4(g43), .Q(n4294) );
  OR2X1 U4815 ( .IN1(n4303), .IN2(n1480), .Q(n1567) );
  AND2X1 U4816 ( .IN1(n4265), .IN2(n1548), .Q(n1480) );
  AND2X1 U4817 ( .IN1(n1548), .IN2(n4293), .Q(n4303) );
  AND2X1 U4818 ( .IN1(n4265), .IN2(n1544), .Q(n4117) );
  AND3X1 U4819 ( .IN1(n4264), .IN2(n3958), .IN3(n4262), .Q(n4265) );
  AND2X1 U4820 ( .IN1(n4087), .IN2(g1308), .Q(n4297) );
  AND2X1 U4821 ( .IN1(n4293), .IN2(n1544), .Q(n4087) );
  AND3X1 U4822 ( .IN1(n4264), .IN2(g42), .IN3(n4262), .Q(n4293) );
  AND2X1 U4823 ( .IN1(n4267), .IN2(g45), .Q(n4262) );
  INVX0 U4824 ( .INP(g44), .ZN(n4267) );
  AND2X1 U4825 ( .IN1(n1486), .IN2(g1543), .Q(n4296) );
  AND2X1 U4826 ( .IN1(n1485), .IN2(g1586), .Q(n4295) );
  OR2X1 U4827 ( .IN1(n4304), .IN2(n4305), .Q(n4282) );
  AND2X1 U4828 ( .IN1(n4086), .IN2(g1738), .Q(n4305) );
  AND2X1 U4829 ( .IN1(g42), .IN2(n4301), .Q(n4086) );
  AND4X1 U4830 ( .IN1(g45), .IN2(n1544), .IN3(g43), .IN4(g44), .Q(n4301) );
  AND3X1 U4831 ( .IN1(n2718), .IN2(n4292), .IN3(g47), .Q(n1544) );
  AND2X1 U4832 ( .IN1(n4096), .IN2(g281), .Q(n4304) );
  AND2X1 U4833 ( .IN1(n4306), .IN2(n4261), .Q(n4096) );
  INVX0 U4834 ( .INP(n4141), .ZN(n4306) );
  AND2X1 U4835 ( .IN1(n3958), .IN2(n4261), .Q(n4141) );
  AND4X1 U4836 ( .IN1(g44), .IN2(n1548), .IN3(n4266), .IN4(n4264), .Q(n4261)
         );
  INVX0 U4837 ( .INP(g43), .ZN(n4264) );
  INVX0 U4838 ( .INP(g45), .ZN(n4266) );
  AND3X1 U4839 ( .IN1(n2722), .IN2(n2718), .IN3(n4292), .Q(n1548) );
  AND2X1 U4840 ( .IN1(n4307), .IN2(g48), .Q(n4292) );
  INVX0 U4841 ( .INP(n2721), .ZN(n4307) );
  AND2X1 U4842 ( .IN1(n4308), .IN2(n4309), .Q(n2721) );
  OR3X1 U4843 ( .IN1(g41), .IN2(g48), .IN3(g30), .Q(n4309) );
  OR2X1 U4844 ( .IN1(n3998), .IN2(g41), .Q(n4308) );
  INVX0 U4845 ( .INP(g46), .ZN(n2718) );
  INVX0 U4846 ( .INP(g47), .ZN(n2722) );
  INVX0 U4847 ( .INP(g42), .ZN(n3958) );
  AND2X1 U4848 ( .IN1(n3998), .IN2(n1637), .Q(n4281) );
  OR2X1 U4849 ( .IN1(g31), .IN2(n4310), .Q(n3998) );
  INVX0 U4850 ( .INP(g48), .ZN(n4310) );
  XOR2X1 U4851 ( .IN1(n2503), .IN2(n3159), .Q(N599) );
  OR3X1 U4852 ( .IN1(n2466), .IN2(n2441), .IN3(n2743), .Q(n3159) );
  INVX0 U4853 ( .INP(n1093), .ZN(n2743) );
  OR2X1 U1550_U1 ( .IN1(g10722), .IN2(n510), .Q(g10461) );
  OR2X1 U1551_U1 ( .IN1(g10664), .IN2(n510), .Q(g10379) );
  INVX0 U1586_U2 ( .INP(n2495), .ZN(U1586_n1) );
  AND2X1 U1586_U1 ( .IN1(n2490), .IN2(U1586_n1), .Q(n1855) );
  INVX0 U1754_U2 ( .INP(n1545), .ZN(U1754_n1) );
  AND2X1 U1754_U1 ( .IN1(n1548), .IN2(U1754_n1), .Q(n1479) );
  INVX0 U1798_U2 ( .INP(n1480), .ZN(U1798_n1) );
  AND2X1 U1798_U1 ( .IN1(n1567), .IN2(U1798_n1), .Q(n1485) );
  INVX0 U1839_U2 ( .INP(n1479), .ZN(U1839_n1) );
  AND2X1 U1839_U1 ( .IN1(n1566), .IN2(U1839_n1), .Q(n1486) );
  INVX0 U1843_U2 ( .INP(n2501), .ZN(U1843_n1) );
  AND2X1 U1843_U1 ( .IN1(n491), .IN2(U1843_n1), .Q(n1478) );
  INVX0 U1877_U2 ( .INP(n505), .ZN(U1877_n1) );
  AND2X1 U1877_U1 ( .IN1(n1137), .IN2(U1877_n1), .Q(n1195) );
  INVX0 U1908_U2 ( .INP(n1545), .ZN(U1908_n1) );
  AND2X1 U1908_U1 ( .IN1(n1544), .IN2(U1908_n1), .Q(n1512) );
  INVX0 U1909_U2 ( .INP(n1545), .ZN(U1909_n1) );
  AND2X1 U1909_U1 ( .IN1(n1574), .IN2(U1909_n1), .Q(n1530) );
  INVX0 U1987_U2 ( .INP(n809), .ZN(U1987_n1) );
  AND2X1 U1987_U1 ( .IN1(n822), .IN2(U1987_n1), .Q(n916) );
  INVX0 U2031_U2 ( .INP(n369), .ZN(U2031_n1) );
  AND2X1 U2031_U1 ( .IN1(n114), .IN2(U2031_n1), .Q(n1056) );
  INVX0 U2035_U2 ( .INP(g109), .ZN(U2035_n1) );
  AND2X1 U2035_U1 ( .IN1(n1404), .IN2(U2035_n1), .Q(n1450) );
  INVX0 U2418_U2 ( .INP(n517), .ZN(U2418_n1) );
  AND2X1 U2418_U1 ( .IN1(g968), .IN2(U2418_n1), .Q(n1564) );
  INVX0 U2468_U2 ( .INP(n1227), .ZN(U2468_n1) );
  AND2X1 U2468_U1 ( .IN1(g1336), .IN2(U2468_n1), .Q(n1231) );
  INVX0 U2478_U2 ( .INP(n1229), .ZN(U2478_n1) );
  AND2X1 U2478_U1 ( .IN1(g1341), .IN2(U2478_n1), .Q(n1232) );
  INVX0 U2488_U2 ( .INP(n46), .ZN(U2488_n1) );
  AND2X1 U2488_U1 ( .IN1(n45), .IN2(U2488_n1), .Q(n1260) );
  INVX0 U2533_U2 ( .INP(n505), .ZN(U2533_n1) );
  AND2X1 U2533_U1 ( .IN1(g178), .IN2(U2533_n1), .Q(g6786) );
  INVX0 U2534_U2 ( .INP(n505), .ZN(U2534_n1) );
  AND2X1 U2534_U1 ( .IN1(g1424), .IN2(U2534_n1), .Q(g6234) );
  INVX0 U2639_U2 ( .INP(n958), .ZN(U2639_n1) );
  AND2X1 U2639_U1 ( .IN1(n962), .IN2(U2639_n1), .Q(n804) );
  INVX0 U2641_U2 ( .INP(g1868), .ZN(U2641_n1) );
  AND2X1 U2641_U1 ( .IN1(n1147), .IN2(U2641_n1), .Q(n926) );
  INVX0 U2654_U2 ( .INP(g750), .ZN(U2654_n1) );
  AND2X1 U2654_U1 ( .IN1(g746), .IN2(U2654_n1), .Q(g4171) );
  INVX0 U2658_U2 ( .INP(n918), .ZN(U2658_n1) );
  AND2X1 U2658_U1 ( .IN1(n917), .IN2(U2658_n1), .Q(n812) );
  INVX0 U2683_U2 ( .INP(n1385), .ZN(U2683_n1) );
  AND2X1 U2683_U1 ( .IN1(g382), .IN2(U2683_n1), .Q(n1420) );
  INVX0 U2699_U2 ( .INP(n493), .ZN(U2699_n1) );
  AND2X1 U2699_U1 ( .IN1(n808), .IN2(U2699_n1), .Q(n806) );
  INVX0 U2846_U2 ( .INP(n1214), .ZN(U2846_n1) );
  AND2X1 U2846_U1 ( .IN1(g4175), .IN2(U2846_n1), .Q(n1193) );
  INVX0 U2847_U2 ( .INP(n1153), .ZN(U2847_n1) );
  AND2X1 U2847_U1 ( .IN1(g4177), .IN2(U2847_n1), .Q(n1125) );
  INVX0 U2848_U2 ( .INP(n1099), .ZN(U2848_n1) );
  AND2X1 U2848_U1 ( .IN1(g4179), .IN2(U2848_n1), .Q(n1093) );
  INVX0 U2859_U2 ( .INP(g12), .ZN(U2859_n1) );
  AND2X1 U2859_U1 ( .IN1(n1137), .IN2(U2859_n1), .Q(n1159) );
  INVX0 U2860_U2 ( .INP(n1151), .ZN(U2860_n1) );
  AND2X1 U2860_U1 ( .IN1(g810), .IN2(U2860_n1), .Q(n1123) );
  INVX0 U2861_U2 ( .INP(n1097), .ZN(U2861_n1) );
  AND2X1 U2861_U1 ( .IN1(g818), .IN2(U2861_n1), .Q(n1090) );
  INVX0 U2867_U2 ( .INP(g1834), .ZN(U2867_n1) );
  AND2X1 U2867_U1 ( .IN1(n817), .IN2(U2867_n1), .Q(n1380) );
  INVX0 U2879_U2 ( .INP(n1656), .ZN(U2879_n1) );
  AND2X1 U2879_U1 ( .IN1(g713), .IN2(U2879_n1), .Q(n967) );
  INVX0 U2881_U2 ( .INP(n1657), .ZN(U2881_n1) );
  AND2X1 U2881_U1 ( .IN1(g1927), .IN2(U2881_n1), .Q(n921) );
  INVX0 U2882_U2 ( .INP(n505), .ZN(U2882_n1) );
  AND2X1 U2882_U1 ( .IN1(g1160), .IN2(U2882_n1), .Q(g4334) );
  INVX0 U2883_U2 ( .INP(n505), .ZN(U2883_n1) );
  AND2X1 U2883_U1 ( .IN1(g1166), .IN2(U2883_n1), .Q(g4325) );
  INVX0 U2884_U2 ( .INP(n505), .ZN(U2884_n1) );
  AND2X1 U2884_U1 ( .IN1(g148), .IN2(U2884_n1), .Q(g6759) );
  INVX0 U2885_U2 ( .INP(n505), .ZN(U2885_n1) );
  AND2X1 U2885_U1 ( .IN1(g1157), .IN2(U2885_n1), .Q(g4338) );
  INVX0 U2886_U2 ( .INP(n505), .ZN(U2886_n1) );
  AND2X1 U2886_U1 ( .IN1(g1163), .IN2(U2886_n1), .Q(g4330) );
  INVX0 U2887_U2 ( .INP(n505), .ZN(U2887_n1) );
  AND2X1 U2887_U1 ( .IN1(g237), .IN2(U2887_n1), .Q(g6821) );
  INVX0 U2888_U2 ( .INP(n505), .ZN(U2888_n1) );
  AND2X1 U2888_U1 ( .IN1(g1499), .IN2(U2888_n1), .Q(g6198) );
  INVX0 U2889_U2 ( .INP(n505), .ZN(U2889_n1) );
  AND2X1 U2889_U1 ( .IN1(g1411), .IN2(U2889_n1), .Q(g6244) );
  INVX0 U2890_U2 ( .INP(n505), .ZN(U2890_n1) );
  AND2X1 U2890_U1 ( .IN1(g225), .IN2(U2890_n1), .Q(g6826) );
  INVX0 U2891_U2 ( .INP(n505), .ZN(U2891_n1) );
  AND2X1 U2891_U1 ( .IN1(g1407), .IN2(U2891_n1), .Q(g6216) );
  INVX0 U2892_U2 ( .INP(n505), .ZN(U2892_n1) );
  AND2X1 U2892_U1 ( .IN1(g213), .IN2(U2892_n1), .Q(g6829) );
  INVX0 U2893_U2 ( .INP(n505), .ZN(U2893_n1) );
  AND2X1 U2893_U1 ( .IN1(g186), .IN2(U2893_n1), .Q(g6833) );
  INVX0 U2894_U2 ( .INP(n505), .ZN(U2894_n1) );
  AND2X1 U2894_U1 ( .IN1(g219), .IN2(U2894_n1), .Q(g6827) );
  INVX0 U2895_U2 ( .INP(n505), .ZN(U2895_n1) );
  AND2X1 U2895_U1 ( .IN1(g143), .IN2(U2895_n1), .Q(g6757) );
  INVX0 U2896_U2 ( .INP(n505), .ZN(U2896_n1) );
  AND2X1 U2896_U1 ( .IN1(g207), .IN2(U2896_n1), .Q(g6831) );
  INVX0 U2897_U2 ( .INP(n505), .ZN(U2897_n1) );
  AND2X1 U2897_U1 ( .IN1(g231), .IN2(U2897_n1), .Q(g6822) );
  INVX0 U2898_U2 ( .INP(n505), .ZN(U2898_n1) );
  AND2X1 U2898_U1 ( .IN1(g192), .IN2(U2898_n1), .Q(g6838) );
  INVX0 U2899_U2 ( .INP(n505), .ZN(U2899_n1) );
  AND2X1 U2899_U1 ( .IN1(test_so3), .IN2(U2899_n1), .Q(g6823) );
  INVX0 U2900_U2 ( .INP(n505), .ZN(U2900_n1) );
  AND2X1 U2900_U1 ( .IN1(g1371), .IN2(U2900_n1), .Q(g6824) );
  INVX0 U2901_U2 ( .INP(n505), .ZN(U2901_n1) );
  AND2X1 U2901_U1 ( .IN1(g1383), .IN2(U2901_n1), .Q(g6832) );
  INVX0 U2902_U2 ( .INP(n505), .ZN(U2902_n1) );
  AND2X1 U2902_U1 ( .IN1(g243), .IN2(U2902_n1), .Q(g6819) );
  INVX0 U3090_U2 ( .INP(g810), .ZN(U3090_n1) );
  AND2X1 U3090_U1 ( .IN1(n1151), .IN2(U3090_n1), .Q(n1150) );
  INVX0 U3092_U2 ( .INP(g818), .ZN(U3092_n1) );
  AND2X1 U3092_U1 ( .IN1(n1097), .IN2(U3092_n1), .Q(n1096) );
  INVX0 U3094_U2 ( .INP(g4179), .ZN(U3094_n1) );
  AND2X1 U3094_U1 ( .IN1(n1099), .IN2(U3094_n1), .Q(n1098) );
  INVX0 U3096_U2 ( .INP(g4175), .ZN(U3096_n1) );
  AND2X1 U3096_U1 ( .IN1(n1214), .IN2(U3096_n1), .Q(n1213) );
  INVX0 U3098_U2 ( .INP(g4177), .ZN(U3098_n1) );
  AND2X1 U3098_U1 ( .IN1(n1153), .IN2(U3098_n1), .Q(n1152) );
  INVX0 U3124_U2 ( .INP(n324), .ZN(U3124_n1) );
  AND2X1 U3124_U1 ( .IN1(n837), .IN2(U3124_n1), .Q(n836) );
  INVX0 U3171_U2 ( .INP(n2500), .ZN(U3171_n1) );
  AND2X1 U3171_U1 ( .IN1(g1610), .IN2(U3171_n1), .Q(g5194) );
endmodule

