module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n236_, new_n238_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n246_, new_n170_, new_n266_, new_n173_, new_n220_, new_n419_, new_n214_, new_n424_, new_n114_, new_n188_, new_n240_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n344_, new_n287_, new_n427_, new_n234_, new_n393_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n124_, new_n164_, new_n230_, new_n281_, new_n430_, new_n248_, new_n117_, new_n167_, new_n385_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n324_, new_n158_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n381_, new_n388_, new_n194_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n216_, new_n280_, new_n426_, new_n235_, new_n301_, new_n169_, new_n395_, new_n383_, new_n210_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n263_, new_n334_, new_n331_, new_n378_, new_n349_, new_n244_, new_n172_, new_n277_, new_n286_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n161_, new_n333_, new_n290_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n227_, new_n416_, new_n222_, new_n328_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n107_, new_n182_, new_n407_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n199_, new_n146_, new_n302_, new_n191_, new_n225_, new_n387_, new_n112_, new_n121_, new_n221_, new_n243_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n174_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n203_, new_n316_, new_n417_, new_n332_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n193_, new_n128_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n175_, new_n226_, new_n185_, new_n171_, new_n434_, new_n200_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n120_, new_n406_, new_n229_, new_n204_, new_n181_, new_n135_, new_n405_;

xnor g000 ( new_n106_, N65, N69 );
xnor g001 ( new_n107_, N73, N77 );
xnor g002 ( new_n108_, new_n106_, new_n107_ );
xnor g003 ( new_n109_, N81, N85 );
xnor g004 ( new_n110_, N89, N93 );
xnor g005 ( new_n111_, new_n109_, new_n110_ );
nand g006 ( new_n112_, new_n108_, new_n111_ );
not g007 ( new_n113_, new_n108_ );
not g008 ( new_n114_, new_n111_ );
nand g009 ( new_n115_, new_n113_, new_n114_ );
nand g010 ( new_n116_, new_n115_, new_n112_ );
nand g011 ( new_n117_, N129, N137 );
nand g012 ( new_n118_, new_n116_, new_n117_ );
nand g013 ( new_n119_, new_n115_, N129, N137, new_n112_ );
nand g014 ( new_n120_, new_n118_, new_n119_ );
xor g015 ( new_n121_, N1, N17 );
xnor g016 ( new_n122_, N33, N49 );
xnor g017 ( new_n123_, new_n121_, new_n122_ );
xor g018 ( new_n124_, new_n123_, keyIn_0_9 );
not g019 ( new_n125_, new_n124_ );
nand g020 ( new_n126_, new_n120_, new_n125_ );
nand g021 ( new_n127_, new_n118_, new_n124_, new_n119_ );
nand g022 ( new_n128_, new_n126_, new_n127_ );
xnor g023 ( new_n129_, N105, N109 );
xnor g024 ( new_n130_, new_n129_, keyIn_0_3 );
xor g025 ( new_n131_, N97, N101 );
nand g026 ( new_n132_, new_n130_, new_n131_ );
or g027 ( new_n133_, new_n130_, new_n131_ );
nand g028 ( new_n134_, new_n133_, new_n132_ );
nand g029 ( new_n135_, new_n134_, new_n108_ );
nand g030 ( new_n136_, new_n133_, new_n113_, new_n132_ );
nand g031 ( new_n137_, new_n135_, new_n136_ );
nand g032 ( new_n138_, N131, N137 );
nand g033 ( new_n139_, new_n137_, new_n138_ );
nand g034 ( new_n140_, new_n135_, N131, N137, new_n136_ );
nand g035 ( new_n141_, new_n139_, new_n140_ );
xnor g036 ( new_n142_, N41, N57 );
xnor g037 ( new_n143_, new_n142_, keyIn_0_6 );
xor g038 ( new_n144_, N9, N25 );
xnor g039 ( new_n145_, new_n143_, new_n144_ );
not g040 ( new_n146_, new_n145_ );
nand g041 ( new_n147_, new_n141_, new_n146_ );
nand g042 ( new_n148_, new_n139_, new_n140_, new_n145_ );
and g043 ( new_n149_, new_n147_, new_n148_ );
xnor g044 ( new_n150_, N113, N117 );
xnor g045 ( new_n151_, new_n150_, keyIn_0_4 );
xor g046 ( new_n152_, N121, N125 );
nand g047 ( new_n153_, new_n151_, new_n152_ );
or g048 ( new_n154_, new_n151_, new_n152_ );
nand g049 ( new_n155_, new_n154_, new_n153_ );
nand g050 ( new_n156_, new_n155_, new_n114_ );
nand g051 ( new_n157_, new_n154_, new_n111_, new_n153_ );
nand g052 ( new_n158_, new_n156_, new_n157_ );
nand g053 ( new_n159_, N132, N137 );
nand g054 ( new_n160_, new_n158_, new_n159_ );
nand g055 ( new_n161_, new_n156_, new_n157_, N132, N137 );
nand g056 ( new_n162_, new_n160_, new_n161_ );
xnor g057 ( new_n163_, N13, N29 );
xnor g058 ( new_n164_, N45, N61 );
xor g059 ( new_n165_, new_n163_, new_n164_ );
not g060 ( new_n166_, new_n165_ );
nand g061 ( new_n167_, new_n162_, new_n166_ );
nand g062 ( new_n168_, new_n160_, new_n161_, new_n165_ );
nand g063 ( new_n169_, new_n167_, new_n168_ );
nand g064 ( new_n170_, new_n134_, new_n155_ );
nand g065 ( new_n171_, new_n133_, new_n154_, new_n132_, new_n153_ );
nand g066 ( new_n172_, new_n170_, new_n171_ );
nand g067 ( new_n173_, N130, N137 );
nand g068 ( new_n174_, new_n172_, new_n173_ );
nand g069 ( new_n175_, new_n170_, N130, N137, new_n171_ );
nand g070 ( new_n176_, new_n174_, new_n175_ );
xor g071 ( new_n177_, N5, N21 );
xnor g072 ( new_n178_, N37, N53 );
xnor g073 ( new_n179_, new_n177_, new_n178_ );
xnor g074 ( new_n180_, new_n176_, new_n179_ );
not g075 ( new_n181_, keyIn_0_11 );
nand g076 ( new_n182_, new_n128_, new_n181_ );
nand g077 ( new_n183_, new_n126_, keyIn_0_11, new_n127_ );
nand g078 ( new_n184_, new_n182_, new_n183_ );
nand g079 ( new_n185_, new_n180_, new_n149_, new_n184_, new_n169_ );
nand g080 ( new_n186_, new_n185_, keyIn_0_19 );
not g081 ( new_n187_, keyIn_0_19 );
nand g082 ( new_n188_, new_n147_, new_n148_ );
and g083 ( new_n189_, new_n167_, new_n168_ );
nor g084 ( new_n190_, new_n189_, new_n188_ );
nand g085 ( new_n191_, new_n190_, new_n187_, new_n180_, new_n184_ );
nand g086 ( new_n192_, new_n191_, new_n186_ );
or g087 ( new_n193_, new_n180_, keyIn_0_13 );
nand g088 ( new_n194_, new_n180_, keyIn_0_13 );
not g089 ( new_n195_, new_n128_ );
nor g090 ( new_n196_, new_n169_, new_n195_ );
nand g091 ( new_n197_, new_n193_, new_n194_, new_n149_, new_n196_ );
not g092 ( new_n198_, new_n180_ );
nand g093 ( new_n199_, new_n198_, keyIn_0_12, new_n188_ );
nand g094 ( new_n200_, new_n188_, keyIn_0_12 );
nand g095 ( new_n201_, new_n200_, new_n180_ );
nor g096 ( new_n202_, new_n169_, new_n128_ );
nand g097 ( new_n203_, new_n199_, new_n201_, new_n202_ );
nand g098 ( new_n204_, new_n192_, new_n197_, new_n203_ );
xnor g099 ( new_n205_, N69, N85 );
xnor g100 ( new_n206_, N101, N117 );
xor g101 ( new_n207_, new_n205_, new_n206_ );
not g102 ( new_n208_, new_n207_ );
nand g103 ( new_n209_, N134, N137 );
not g104 ( new_n210_, keyIn_0_1 );
nand g105 ( new_n211_, N33, N37 );
or g106 ( new_n212_, N33, N37 );
nand g107 ( new_n213_, new_n212_, new_n210_, new_n211_ );
nand g108 ( new_n214_, new_n212_, new_n211_ );
nand g109 ( new_n215_, new_n214_, keyIn_0_1 );
nand g110 ( new_n216_, new_n215_, new_n213_ );
not g111 ( new_n217_, keyIn_0_2 );
nand g112 ( new_n218_, N41, N45 );
or g113 ( new_n219_, N41, N45 );
nand g114 ( new_n220_, new_n219_, new_n217_, new_n218_ );
xnor g115 ( new_n221_, N41, N45 );
nand g116 ( new_n222_, new_n221_, keyIn_0_2 );
nand g117 ( new_n223_, new_n222_, new_n220_ );
nand g118 ( new_n224_, new_n216_, new_n223_ );
nand g119 ( new_n225_, new_n215_, new_n222_, new_n213_, new_n220_ );
nand g120 ( new_n226_, new_n224_, keyIn_0_8, new_n225_ );
not g121 ( new_n227_, keyIn_0_8 );
nand g122 ( new_n228_, new_n224_, new_n225_ );
nand g123 ( new_n229_, new_n228_, new_n227_ );
xnor g124 ( new_n230_, N49, N53 );
xnor g125 ( new_n231_, N57, N61 );
xnor g126 ( new_n232_, new_n230_, new_n231_ );
nand g127 ( new_n233_, new_n229_, new_n226_, new_n232_ );
nand g128 ( new_n234_, new_n229_, new_n226_ );
not g129 ( new_n235_, new_n232_ );
nand g130 ( new_n236_, new_n234_, new_n235_ );
nand g131 ( new_n237_, new_n236_, new_n233_ );
nand g132 ( new_n238_, new_n237_, new_n209_ );
nand g133 ( new_n239_, new_n236_, N134, N137, new_n233_ );
nand g134 ( new_n240_, new_n238_, new_n239_ );
nand g135 ( new_n241_, new_n240_, new_n208_ );
nand g136 ( new_n242_, new_n238_, new_n207_, new_n239_ );
nand g137 ( new_n243_, new_n241_, new_n242_ );
not g138 ( new_n244_, new_n243_ );
nand g139 ( new_n245_, new_n244_, keyIn_0_14 );
nand g140 ( new_n246_, N17, N21 );
or g141 ( new_n247_, N17, N21 );
nand g142 ( new_n248_, new_n247_, keyIn_0_0, new_n246_ );
not g143 ( new_n249_, keyIn_0_0 );
xnor g144 ( new_n250_, N17, N21 );
nand g145 ( new_n251_, new_n250_, new_n249_ );
xor g146 ( new_n252_, N25, N29 );
not g147 ( new_n253_, new_n252_ );
nand g148 ( new_n254_, new_n253_, new_n248_, new_n251_ );
nand g149 ( new_n255_, new_n251_, new_n248_ );
nand g150 ( new_n256_, new_n255_, new_n252_ );
nand g151 ( new_n257_, new_n256_, new_n254_ );
xnor g152 ( new_n258_, N1, N5 );
xnor g153 ( new_n259_, N9, N13 );
xnor g154 ( new_n260_, new_n258_, new_n259_ );
xnor g155 ( new_n261_, new_n257_, new_n260_ );
nand g156 ( new_n262_, N133, N137 );
xnor g157 ( new_n263_, new_n261_, new_n262_ );
xnor g158 ( new_n264_, N65, N81 );
xnor g159 ( new_n265_, N97, N113 );
xnor g160 ( new_n266_, new_n264_, new_n265_ );
xnor g161 ( new_n267_, new_n263_, new_n266_ );
not g162 ( new_n268_, new_n267_ );
xnor g163 ( new_n269_, N105, N121 );
xnor g164 ( new_n270_, new_n269_, keyIn_0_7 );
xor g165 ( new_n271_, N73, N89 );
xnor g166 ( new_n272_, new_n270_, new_n271_ );
not g167 ( new_n273_, new_n272_ );
nand g168 ( new_n274_, N135, N137 );
xnor g169 ( new_n275_, new_n274_, keyIn_0_5 );
not g170 ( new_n276_, new_n275_ );
nand g171 ( new_n277_, new_n229_, new_n226_, new_n260_ );
not g172 ( new_n278_, new_n260_ );
nand g173 ( new_n279_, new_n234_, new_n278_ );
nand g174 ( new_n280_, new_n279_, new_n277_ );
nand g175 ( new_n281_, new_n280_, new_n276_ );
nand g176 ( new_n282_, new_n279_, new_n275_, new_n277_ );
nand g177 ( new_n283_, new_n281_, new_n282_ );
nand g178 ( new_n284_, new_n283_, new_n273_ );
nand g179 ( new_n285_, new_n281_, new_n272_, new_n282_ );
and g180 ( new_n286_, new_n284_, new_n285_ );
nand g181 ( new_n287_, new_n245_, new_n268_, new_n286_ );
nor g182 ( new_n288_, new_n244_, keyIn_0_14 );
not g183 ( new_n289_, keyIn_0_10 );
nand g184 ( new_n290_, N136, N137 );
nand g185 ( new_n291_, new_n257_, new_n232_ );
nand g186 ( new_n292_, new_n235_, new_n254_, new_n256_ );
nand g187 ( new_n293_, new_n291_, new_n292_ );
nand g188 ( new_n294_, new_n293_, new_n290_ );
nand g189 ( new_n295_, new_n291_, new_n292_, N136, N137 );
nand g190 ( new_n296_, new_n294_, new_n289_, new_n295_ );
nand g191 ( new_n297_, new_n294_, new_n295_ );
nand g192 ( new_n298_, new_n297_, keyIn_0_10 );
nand g193 ( new_n299_, new_n298_, new_n296_ );
xnor g194 ( new_n300_, N77, N93 );
xnor g195 ( new_n301_, N109, N125 );
xor g196 ( new_n302_, new_n300_, new_n301_ );
not g197 ( new_n303_, new_n302_ );
nand g198 ( new_n304_, new_n299_, new_n303_ );
nand g199 ( new_n305_, new_n298_, new_n296_, new_n302_ );
nand g200 ( new_n306_, new_n304_, new_n305_ );
xnor g201 ( new_n307_, new_n306_, keyIn_0_15 );
nor g202 ( new_n308_, new_n287_, new_n307_, new_n288_ );
nand g203 ( new_n309_, new_n204_, new_n308_ );
nand g204 ( new_n310_, new_n309_, keyIn_0_24 );
not g205 ( new_n311_, keyIn_0_24 );
nand g206 ( new_n312_, new_n204_, new_n308_, new_n311_ );
nand g207 ( new_n313_, new_n310_, new_n312_ );
nand g208 ( new_n314_, new_n313_, new_n128_ );
xnor g209 ( N724, new_n314_, N1 );
nand g210 ( new_n316_, new_n313_, new_n198_ );
xnor g211 ( N725, new_n316_, N5 );
nand g212 ( new_n318_, new_n313_, new_n188_ );
nand g213 ( new_n319_, new_n318_, N9 );
not g214 ( new_n320_, N9 );
nand g215 ( new_n321_, new_n313_, new_n320_, new_n188_ );
nand g216 ( new_n322_, new_n319_, new_n321_ );
nand g217 ( new_n323_, new_n322_, keyIn_0_30 );
not g218 ( new_n324_, keyIn_0_30 );
nand g219 ( new_n325_, new_n319_, new_n324_, new_n321_ );
nand g220 ( N726, new_n323_, new_n325_ );
nand g221 ( new_n327_, new_n313_, new_n169_ );
nand g222 ( new_n328_, new_n327_, N13 );
not g223 ( new_n329_, N13 );
nand g224 ( new_n330_, new_n313_, new_n329_, new_n169_ );
nand g225 ( new_n331_, new_n328_, new_n330_ );
nand g226 ( new_n332_, new_n331_, keyIn_0_31 );
not g227 ( new_n333_, keyIn_0_31 );
nand g228 ( new_n334_, new_n328_, new_n333_, new_n330_ );
nand g229 ( N727, new_n332_, new_n334_ );
nor g230 ( new_n336_, new_n244_, new_n267_ );
nand g231 ( new_n337_, new_n284_, new_n285_ );
and g232 ( new_n338_, new_n337_, new_n306_ );
and g233 ( new_n339_, new_n204_, new_n336_, new_n338_ );
nand g234 ( new_n340_, new_n339_, new_n128_ );
xnor g235 ( N728, new_n340_, N17 );
nand g236 ( new_n342_, new_n339_, new_n198_ );
xnor g237 ( N729, new_n342_, N21 );
not g238 ( new_n344_, keyIn_0_25 );
nand g239 ( new_n345_, new_n339_, new_n188_ );
xnor g240 ( new_n346_, new_n345_, new_n344_ );
xnor g241 ( N730, new_n346_, N25 );
nand g242 ( new_n348_, new_n339_, new_n169_ );
xnor g243 ( new_n349_, new_n348_, keyIn_0_26 );
xnor g244 ( N731, new_n349_, N29 );
nor g245 ( new_n351_, new_n243_, new_n306_ );
xnor g246 ( new_n352_, new_n267_, keyIn_0_16 );
nand g247 ( new_n353_, new_n204_, new_n286_, new_n351_, new_n352_ );
not g248 ( new_n354_, new_n353_ );
nand g249 ( new_n355_, new_n354_, new_n128_ );
xnor g250 ( N732, new_n355_, N33 );
nand g251 ( new_n357_, new_n354_, new_n198_ );
xnor g252 ( N733, new_n357_, N37 );
nand g253 ( new_n359_, new_n354_, new_n188_ );
xnor g254 ( N734, new_n359_, N41 );
nand g255 ( new_n361_, new_n354_, new_n169_ );
xnor g256 ( N735, new_n361_, N45 );
xor g257 ( new_n363_, new_n267_, keyIn_0_17 );
nand g258 ( new_n364_, new_n204_, new_n244_, new_n338_, new_n363_ );
not g259 ( new_n365_, new_n364_ );
nand g260 ( new_n366_, new_n365_, new_n128_ );
xnor g261 ( N736, new_n366_, N49 );
nand g262 ( new_n368_, new_n365_, new_n198_ );
xnor g263 ( N737, new_n368_, N53 );
nand g264 ( new_n370_, new_n365_, new_n188_ );
xnor g265 ( N738, new_n370_, N57 );
nand g266 ( new_n372_, new_n365_, new_n169_ );
xnor g267 ( N739, new_n372_, N61 );
nand g268 ( new_n374_, new_n243_, new_n337_, new_n306_, new_n267_ );
nand g269 ( new_n375_, new_n374_, keyIn_0_20 );
not g270 ( new_n376_, keyIn_0_20 );
and g271 ( new_n377_, new_n243_, new_n267_ );
nand g272 ( new_n378_, new_n338_, new_n377_, new_n376_ );
nand g273 ( new_n379_, new_n378_, new_n375_ );
and g274 ( new_n380_, new_n304_, new_n305_ );
xnor g275 ( new_n381_, new_n337_, keyIn_0_18 );
nand g276 ( new_n382_, new_n381_, new_n380_, new_n336_ );
nand g277 ( new_n383_, new_n244_, new_n380_, new_n267_, new_n337_ );
nand g278 ( new_n384_, new_n383_, keyIn_0_22 );
not g279 ( new_n385_, keyIn_0_22 );
nand g280 ( new_n386_, new_n351_, new_n385_, new_n267_, new_n337_ );
nand g281 ( new_n387_, new_n384_, new_n386_ );
nand g282 ( new_n388_, new_n286_, new_n380_, new_n243_, new_n267_ );
nand g283 ( new_n389_, new_n388_, keyIn_0_21 );
not g284 ( new_n390_, keyIn_0_21 );
nor g285 ( new_n391_, new_n337_, new_n306_ );
nand g286 ( new_n392_, new_n377_, new_n390_, new_n391_ );
nand g287 ( new_n393_, new_n389_, new_n392_ );
nand g288 ( new_n394_, new_n387_, new_n393_, new_n379_, new_n382_ );
xnor g289 ( new_n395_, new_n394_, keyIn_0_23 );
and g290 ( new_n396_, new_n196_, new_n188_, new_n180_ );
nand g291 ( new_n397_, new_n395_, new_n268_, new_n396_ );
xnor g292 ( N740, new_n397_, N65 );
nand g293 ( new_n399_, new_n395_, new_n244_, new_n396_ );
xnor g294 ( N741, new_n399_, N69 );
nand g295 ( new_n401_, new_n395_, new_n286_, new_n396_ );
xnor g296 ( N742, new_n401_, N73 );
nand g297 ( new_n403_, new_n395_, new_n306_, new_n396_ );
xnor g298 ( N743, new_n403_, N77 );
not g299 ( new_n405_, new_n190_ );
nor g300 ( new_n406_, new_n405_, new_n195_, new_n198_ );
nand g301 ( new_n407_, new_n395_, new_n268_, new_n406_ );
xnor g302 ( N744, new_n407_, N81 );
nand g303 ( new_n409_, new_n395_, new_n244_, new_n406_ );
xnor g304 ( new_n410_, keyIn_0_27, N85 );
xnor g305 ( N745, new_n409_, new_n410_ );
nand g306 ( new_n412_, new_n395_, new_n286_, new_n406_ );
xnor g307 ( N746, new_n412_, N89 );
nand g308 ( new_n414_, new_n395_, new_n306_, new_n406_ );
xnor g309 ( N747, new_n414_, N93 );
nor g310 ( new_n416_, new_n180_, new_n149_, new_n128_, new_n169_ );
nand g311 ( new_n417_, new_n395_, new_n268_, new_n416_ );
xnor g312 ( N748, new_n417_, N97 );
nand g313 ( new_n419_, new_n395_, new_n244_, new_n416_ );
xnor g314 ( N749, new_n419_, N101 );
nand g315 ( new_n421_, new_n395_, new_n286_, new_n416_ );
xnor g316 ( N750, new_n421_, N105 );
nand g317 ( new_n423_, new_n395_, new_n306_, new_n416_ );
xor g318 ( new_n424_, keyIn_0_28, N109 );
xnor g319 ( N751, new_n423_, new_n424_ );
nor g320 ( new_n426_, new_n405_, new_n128_, new_n180_ );
nand g321 ( new_n427_, new_n395_, new_n268_, new_n426_ );
xnor g322 ( N752, new_n427_, N113 );
not g323 ( new_n429_, N117 );
not g324 ( new_n430_, keyIn_0_29 );
and g325 ( new_n431_, new_n379_, new_n382_ );
nand g326 ( new_n432_, new_n431_, keyIn_0_23, new_n387_, new_n393_ );
not g327 ( new_n433_, keyIn_0_23 );
nand g328 ( new_n434_, new_n394_, new_n433_ );
nand g329 ( new_n435_, new_n432_, new_n434_, new_n244_, new_n426_ );
nand g330 ( new_n436_, new_n435_, new_n430_ );
nand g331 ( new_n437_, new_n395_, keyIn_0_29, new_n244_, new_n426_ );
nand g332 ( new_n438_, new_n437_, new_n436_ );
nand g333 ( new_n439_, new_n438_, new_n429_ );
nand g334 ( new_n440_, new_n437_, N117, new_n436_ );
nand g335 ( N753, new_n439_, new_n440_ );
nand g336 ( new_n442_, new_n395_, new_n286_, new_n426_ );
xnor g337 ( N754, new_n442_, N121 );
nand g338 ( new_n444_, new_n395_, new_n306_, new_n426_ );
xnor g339 ( N755, new_n444_, N125 );
endmodule