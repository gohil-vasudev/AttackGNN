module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n155_, new_n384_, new_n410_, new_n445_, new_n236_, new_n238_, new_n92_, new_n79_, new_n250_, new_n113_, new_n288_, new_n371_, new_n97_, new_n454_, new_n421_, new_n202_, new_n296_, new_n308_, new_n368_, new_n232_, new_n258_, new_n76_, new_n439_, new_n176_, new_n283_, new_n223_, new_n390_, new_n156_, new_n306_, new_n366_, new_n291_, new_n261_, new_n241_, new_n309_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n82_, new_n401_, new_n389_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n456_, new_n170_, new_n246_, new_n400_, new_n328_, new_n460_, new_n266_, new_n367_, new_n173_, new_n220_, new_n130_, new_n419_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n214_, new_n451_, new_n424_, new_n138_, new_n310_, new_n144_, new_n275_, new_n114_, new_n188_, new_n240_, new_n413_, new_n352_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n126_, new_n462_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n317_, new_n102_, new_n344_, new_n143_, new_n287_, new_n125_, new_n145_, new_n253_, new_n403_, new_n90_, new_n237_, new_n427_, new_n234_, new_n149_, new_n472_, new_n393_, new_n260_, new_n418_, new_n251_, new_n189_, new_n300_, new_n292_, new_n106_, new_n411_, new_n215_, new_n152_, new_n157_, new_n107_, new_n93_, new_n182_, new_n153_, new_n407_, new_n81_, new_n133_, new_n257_, new_n212_, new_n151_, new_n364_, new_n219_, new_n231_, new_n313_, new_n78_, new_n239_, new_n382_, new_n272_, new_n282_, new_n201_, new_n428_, new_n192_, new_n414_, new_n199_, new_n146_, new_n88_, new_n360_, new_n98_, new_n110_, new_n315_, new_n302_, new_n191_, new_n124_, new_n326_, new_n95_, new_n225_, new_n164_, new_n230_, new_n281_, new_n430_, new_n87_, new_n387_, new_n103_, new_n112_, new_n248_, new_n350_, new_n117_, new_n121_, new_n415_, new_n167_, new_n221_, new_n385_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n297_, new_n361_, new_n468_, new_n150_, new_n354_, new_n392_, new_n444_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n105_, new_n340_, new_n147_, new_n285_, new_n80_, new_n351_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n325_, new_n417_, new_n180_, new_n332_, new_n318_, new_n453_, new_n163_, new_n148_, new_n321_, new_n440_, new_n443_, new_n324_, new_n122_, new_n111_, new_n158_, new_n252_, new_n466_, new_n262_, new_n160_, new_n312_, new_n271_, new_n274_, new_n372_, new_n100_, new_n242_, new_n218_, new_n115_, new_n307_, new_n190_, new_n305_, new_n420_, new_n408_, new_n470_, new_n423_, new_n205_, new_n213_, new_n134_, new_n141_, new_n433_, new_n435_, new_n206_, new_n109_, new_n254_, new_n429_, new_n355_, new_n353_, new_n85_, new_n432_, new_n265_, new_n370_, new_n256_, new_n452_, new_n278_, new_n304_, new_n381_, new_n388_, new_n217_, new_n101_, new_n269_, new_n194_, new_n394_, new_n116_, new_n299_, new_n129_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n412_, new_n165_, new_n441_, new_n327_, new_n216_, new_n431_, new_n77_, new_n196_, new_n280_, new_n319_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n338_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n187_, new_n311_, new_n86_, new_n465_, new_n84_, new_n195_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n357_, new_n320_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n89_, new_n467_, new_n286_, new_n404_, new_n335_, new_n193_, new_n91_, new_n346_, new_n396_, new_n198_, new_n438_, new_n128_, new_n358_, new_n208_, new_n348_, new_n159_, new_n83_, new_n322_, new_n228_, new_n289_, new_n179_, new_n425_, new_n436_, new_n175_, new_n226_, new_n397_, new_n104_, new_n185_, new_n399_, new_n373_, new_n171_, new_n434_, new_n200_, new_n422_, new_n99_, new_n329_, new_n249_, new_n233_, new_n284_, new_n469_, new_n119_, new_n293_, new_n391_, new_n96_, new_n178_, new_n437_, new_n168_, new_n279_, new_n455_, new_n295_, new_n359_, new_n132_, new_n120_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n406_, new_n356_, new_n333_, new_n229_, new_n290_, new_n464_, new_n94_, new_n204_, new_n369_, new_n181_, new_n135_, new_n448_, new_n276_, new_n405_;

not g000 ( new_n76_, keyIn_0_6 );
not g001 ( new_n77_, N17 );
and g002 ( new_n78_, keyIn_0_0, N11 );
not g003 ( new_n79_, new_n78_ );
or g004 ( new_n80_, keyIn_0_0, N11 );
and g005 ( new_n81_, new_n79_, new_n80_ );
or g006 ( new_n82_, new_n81_, new_n77_ );
and g007 ( new_n83_, new_n82_, keyIn_0_3 );
not g008 ( new_n84_, keyIn_0_3 );
not g009 ( new_n85_, new_n81_ );
and g010 ( new_n86_, new_n85_, new_n84_, N17 );
or g011 ( new_n87_, new_n83_, new_n86_ );
not g012 ( new_n88_, N1 );
and g013 ( new_n89_, new_n88_, N4 );
not g014 ( new_n90_, new_n89_ );
not g015 ( new_n91_, N76 );
and g016 ( new_n92_, new_n91_, N82 );
not g017 ( new_n93_, new_n92_ );
and g018 ( new_n94_, new_n90_, new_n93_ );
not g019 ( new_n95_, N50 );
and g020 ( new_n96_, new_n95_, N56 );
not g021 ( new_n97_, new_n96_ );
not g022 ( new_n98_, N102 );
and g023 ( new_n99_, new_n98_, N108 );
not g024 ( new_n100_, new_n99_ );
not g025 ( new_n101_, N30 );
or g026 ( new_n102_, new_n101_, N24 );
not g027 ( new_n103_, N43 );
or g028 ( new_n104_, new_n103_, N37 );
and g029 ( new_n105_, new_n102_, new_n104_ );
and g030 ( new_n106_, new_n94_, new_n105_, new_n97_, new_n100_ );
not g031 ( new_n107_, N69 );
and g032 ( new_n108_, keyIn_0_1, N63 );
not g033 ( new_n109_, new_n108_ );
or g034 ( new_n110_, keyIn_0_1, N63 );
and g035 ( new_n111_, new_n109_, new_n110_ );
or g036 ( new_n112_, new_n111_, new_n107_ );
and g037 ( new_n113_, new_n112_, keyIn_0_4 );
not g038 ( new_n114_, keyIn_0_4 );
not g039 ( new_n115_, new_n111_ );
and g040 ( new_n116_, new_n115_, new_n114_, N69 );
or g041 ( new_n117_, new_n113_, new_n116_ );
not g042 ( new_n118_, keyIn_0_5 );
not g043 ( new_n119_, N95 );
not g044 ( new_n120_, keyIn_0_2 );
and g045 ( new_n121_, new_n120_, N89 );
not g046 ( new_n122_, N89 );
and g047 ( new_n123_, new_n122_, keyIn_0_2 );
or g048 ( new_n124_, new_n121_, new_n123_, new_n119_ );
and g049 ( new_n125_, new_n124_, new_n118_ );
not g050 ( new_n126_, new_n121_ );
not g051 ( new_n127_, new_n123_ );
and g052 ( new_n128_, new_n126_, new_n127_, keyIn_0_5, N95 );
or g053 ( new_n129_, new_n125_, new_n128_ );
and g054 ( new_n130_, new_n87_, new_n117_, new_n106_, new_n129_ );
not g055 ( new_n131_, new_n130_ );
and g056 ( new_n132_, new_n131_, new_n76_ );
and g057 ( new_n133_, new_n87_, new_n106_ );
and g058 ( new_n134_, new_n117_, new_n129_ );
and g059 ( new_n135_, new_n133_, new_n134_, keyIn_0_6 );
or g060 ( N223, new_n132_, new_n135_ );
not g061 ( new_n137_, new_n129_ );
or g062 ( new_n138_, new_n130_, keyIn_0_6 );
not g063 ( new_n139_, new_n135_ );
and g064 ( new_n140_, new_n139_, new_n138_ );
or g065 ( new_n141_, new_n140_, keyIn_0_7 );
not g066 ( new_n142_, keyIn_0_7 );
or g067 ( new_n143_, new_n132_, new_n142_, new_n135_ );
and g068 ( new_n144_, new_n141_, new_n143_ );
or g069 ( new_n145_, new_n144_, new_n137_ );
and g070 ( new_n146_, N223, new_n142_ );
not g071 ( new_n147_, new_n143_ );
or g072 ( new_n148_, new_n146_, new_n147_, new_n129_ );
and g073 ( new_n149_, new_n145_, new_n148_ );
or g074 ( new_n150_, new_n149_, keyIn_0_10 );
not g075 ( new_n151_, keyIn_0_10 );
or g076 ( new_n152_, new_n146_, new_n147_ );
and g077 ( new_n153_, new_n152_, new_n129_ );
not g078 ( new_n154_, new_n148_ );
or g079 ( new_n155_, new_n153_, new_n154_, new_n151_ );
and g080 ( new_n156_, new_n150_, new_n155_ );
or g081 ( new_n157_, new_n156_, new_n119_, N99 );
and g082 ( new_n158_, new_n157_, keyIn_0_12 );
not g083 ( new_n159_, keyIn_0_12 );
not g084 ( new_n160_, N99 );
or g085 ( new_n161_, new_n153_, new_n154_ );
and g086 ( new_n162_, new_n161_, new_n151_ );
not g087 ( new_n163_, new_n155_ );
or g088 ( new_n164_, new_n162_, new_n163_ );
and g089 ( new_n165_, new_n164_, new_n159_, N95, new_n160_ );
or g090 ( new_n166_, new_n158_, new_n165_ );
not g091 ( new_n167_, keyIn_0_11 );
or g092 ( new_n168_, new_n144_, new_n89_ );
or g093 ( new_n169_, new_n146_, new_n147_, new_n90_ );
and g094 ( new_n170_, new_n168_, new_n169_ );
or g095 ( new_n171_, new_n170_, keyIn_0_8 );
not g096 ( new_n172_, keyIn_0_8 );
and g097 ( new_n173_, new_n152_, new_n90_ );
not g098 ( new_n174_, new_n169_ );
or g099 ( new_n175_, new_n173_, new_n174_, new_n172_ );
and g100 ( new_n176_, new_n171_, new_n175_ );
not g101 ( new_n177_, N4 );
or g102 ( new_n178_, new_n177_, N8 );
or g103 ( new_n179_, new_n176_, new_n178_ );
and g104 ( new_n180_, new_n179_, new_n167_ );
not g105 ( new_n181_, N8 );
or g106 ( new_n182_, new_n173_, new_n174_ );
and g107 ( new_n183_, new_n182_, new_n172_ );
not g108 ( new_n184_, new_n175_ );
or g109 ( new_n185_, new_n183_, new_n184_ );
and g110 ( new_n186_, new_n185_, keyIn_0_11, N4, new_n181_ );
or g111 ( new_n187_, new_n180_, new_n186_ );
not g112 ( new_n188_, N21 );
not g113 ( new_n189_, keyIn_0_9 );
not g114 ( new_n190_, new_n87_ );
or g115 ( new_n191_, new_n144_, new_n190_ );
not g116 ( new_n192_, new_n191_ );
and g117 ( new_n193_, new_n144_, new_n190_ );
or g118 ( new_n194_, new_n192_, new_n193_, new_n189_ );
not g119 ( new_n195_, new_n193_ );
and g120 ( new_n196_, new_n195_, new_n191_ );
or g121 ( new_n197_, new_n196_, keyIn_0_9 );
and g122 ( new_n198_, new_n197_, N17, new_n194_ );
and g123 ( new_n199_, new_n198_, new_n188_ );
not g124 ( new_n200_, new_n199_ );
not g125 ( new_n201_, N56 );
or g126 ( new_n202_, new_n152_, new_n97_ );
or g127 ( new_n203_, new_n144_, new_n96_ );
and g128 ( new_n204_, new_n202_, new_n203_ );
or g129 ( new_n205_, new_n204_, new_n201_ );
or g130 ( new_n206_, new_n205_, N60 );
not g131 ( new_n207_, N108 );
or g132 ( new_n208_, new_n152_, new_n100_ );
or g133 ( new_n209_, new_n144_, new_n99_ );
and g134 ( new_n210_, new_n208_, new_n209_ );
or g135 ( new_n211_, new_n210_, new_n207_ );
or g136 ( new_n212_, new_n211_, N112 );
and g137 ( new_n213_, new_n206_, new_n212_ );
not g138 ( new_n214_, N82 );
or g139 ( new_n215_, new_n152_, new_n93_ );
or g140 ( new_n216_, new_n144_, new_n92_ );
and g141 ( new_n217_, new_n215_, new_n216_ );
or g142 ( new_n218_, new_n217_, new_n214_ );
or g143 ( new_n219_, new_n218_, N86 );
or g144 ( new_n220_, new_n152_, new_n104_ );
not g145 ( new_n221_, new_n104_ );
or g146 ( new_n222_, new_n144_, new_n221_ );
and g147 ( new_n223_, new_n220_, new_n222_ );
or g148 ( new_n224_, new_n223_, new_n103_ );
or g149 ( new_n225_, new_n224_, N47 );
or g150 ( new_n226_, new_n152_, new_n117_ );
not g151 ( new_n227_, new_n117_ );
or g152 ( new_n228_, new_n144_, new_n227_ );
and g153 ( new_n229_, new_n226_, new_n228_ );
or g154 ( new_n230_, new_n229_, new_n107_ );
or g155 ( new_n231_, new_n230_, N73 );
or g156 ( new_n232_, new_n152_, new_n102_ );
not g157 ( new_n233_, new_n102_ );
or g158 ( new_n234_, new_n144_, new_n233_ );
and g159 ( new_n235_, new_n232_, new_n234_ );
or g160 ( new_n236_, new_n235_, new_n101_ );
or g161 ( new_n237_, new_n236_, N34 );
and g162 ( new_n238_, new_n219_, new_n225_, new_n231_, new_n237_ );
and g163 ( new_n239_, new_n200_, new_n238_, new_n213_ );
and g164 ( new_n240_, new_n166_, new_n187_, new_n239_ );
or g165 ( new_n241_, new_n240_, keyIn_0_13 );
and g166 ( new_n242_, new_n166_, keyIn_0_13, new_n187_, new_n239_ );
not g167 ( new_n243_, new_n242_ );
and g168 ( new_n244_, new_n241_, new_n243_ );
not g169 ( N329, new_n244_ );
not g170 ( new_n246_, keyIn_0_18 );
not g171 ( new_n247_, keyIn_0_16 );
not g172 ( new_n248_, new_n180_ );
not g173 ( new_n249_, new_n186_ );
and g174 ( new_n250_, new_n248_, new_n249_ );
not g175 ( new_n251_, keyIn_0_15 );
or g176 ( new_n252_, new_n244_, new_n251_ );
and g177 ( new_n253_, new_n241_, new_n251_, new_n243_ );
not g178 ( new_n254_, new_n253_ );
and g179 ( new_n255_, new_n252_, new_n254_ );
or g180 ( new_n256_, new_n255_, new_n250_ );
and g181 ( new_n257_, new_n252_, new_n250_, new_n254_ );
not g182 ( new_n258_, new_n257_ );
and g183 ( new_n259_, new_n256_, new_n247_, new_n258_ );
not g184 ( new_n260_, new_n259_ );
or g185 ( new_n261_, new_n176_, new_n177_, N14 );
not g186 ( new_n262_, new_n261_ );
and g187 ( new_n263_, new_n262_, keyIn_0_14 );
not g188 ( new_n264_, keyIn_0_14 );
and g189 ( new_n265_, new_n261_, new_n264_ );
or g190 ( new_n266_, new_n263_, new_n265_ );
and g191 ( new_n267_, new_n256_, new_n258_ );
or g192 ( new_n268_, new_n267_, new_n247_ );
and g193 ( new_n269_, new_n268_, new_n260_, new_n266_ );
not g194 ( new_n270_, new_n269_ );
and g195 ( new_n271_, new_n270_, new_n246_ );
and g196 ( new_n272_, new_n269_, keyIn_0_18 );
or g197 ( new_n273_, new_n271_, new_n272_ );
not g198 ( new_n274_, keyIn_0_19 );
not g199 ( new_n275_, new_n206_ );
or g200 ( new_n276_, new_n255_, new_n275_ );
and g201 ( new_n277_, new_n252_, new_n275_, new_n254_ );
not g202 ( new_n278_, new_n277_ );
and g203 ( new_n279_, new_n276_, new_n278_ );
or g204 ( new_n280_, new_n279_, keyIn_0_17 );
and g205 ( new_n281_, new_n276_, keyIn_0_17, new_n278_ );
not g206 ( new_n282_, new_n281_ );
and g207 ( new_n283_, new_n280_, new_n282_ );
or g208 ( new_n284_, new_n205_, N66 );
or g209 ( new_n285_, new_n283_, new_n284_ );
and g210 ( new_n286_, new_n285_, new_n274_ );
not g211 ( new_n287_, N66 );
not g212 ( new_n288_, new_n205_ );
not g213 ( new_n289_, new_n283_ );
and g214 ( new_n290_, new_n289_, keyIn_0_19, new_n287_, new_n288_ );
or g215 ( new_n291_, new_n286_, new_n290_ );
not g216 ( new_n292_, new_n225_ );
and g217 ( new_n293_, new_n255_, new_n292_ );
not g218 ( new_n294_, new_n293_ );
or g219 ( new_n295_, new_n255_, new_n292_ );
and g220 ( new_n296_, new_n294_, new_n295_ );
or g221 ( new_n297_, new_n296_, N53, new_n224_ );
not g222 ( new_n298_, new_n212_ );
or g223 ( new_n299_, new_n255_, new_n298_ );
and g224 ( new_n300_, new_n255_, new_n298_ );
not g225 ( new_n301_, new_n300_ );
and g226 ( new_n302_, new_n301_, new_n299_ );
or g227 ( new_n303_, new_n302_, N115, new_n211_ );
not g228 ( new_n304_, new_n231_ );
and g229 ( new_n305_, new_n255_, new_n304_ );
not g230 ( new_n306_, new_n305_ );
or g231 ( new_n307_, new_n255_, new_n304_ );
and g232 ( new_n308_, new_n306_, new_n307_ );
or g233 ( new_n309_, new_n308_, N79, new_n230_ );
and g234 ( new_n310_, new_n297_, new_n303_, new_n309_ );
and g235 ( new_n311_, new_n255_, new_n199_ );
not g236 ( new_n312_, new_n311_ );
or g237 ( new_n313_, new_n255_, new_n199_ );
and g238 ( new_n314_, new_n312_, new_n313_ );
not g239 ( new_n315_, N27 );
and g240 ( new_n316_, new_n198_, new_n315_ );
not g241 ( new_n317_, new_n316_ );
or g242 ( new_n318_, new_n314_, new_n317_ );
not g243 ( new_n319_, new_n237_ );
and g244 ( new_n320_, new_n255_, new_n319_ );
not g245 ( new_n321_, new_n320_ );
or g246 ( new_n322_, new_n255_, new_n319_ );
and g247 ( new_n323_, new_n321_, new_n322_ );
or g248 ( new_n324_, new_n323_, N40, new_n236_ );
and g249 ( new_n325_, new_n324_, new_n318_ );
not g250 ( new_n326_, new_n219_ );
or g251 ( new_n327_, new_n255_, new_n326_ );
and g252 ( new_n328_, new_n255_, new_n326_ );
not g253 ( new_n329_, new_n328_ );
and g254 ( new_n330_, new_n329_, new_n327_ );
or g255 ( new_n331_, new_n330_, N92, new_n218_ );
and g256 ( new_n332_, new_n164_, N95, new_n160_ );
or g257 ( new_n333_, new_n332_, new_n159_ );
not g258 ( new_n334_, new_n165_ );
and g259 ( new_n335_, new_n333_, new_n334_ );
and g260 ( new_n336_, new_n255_, new_n335_ );
not g261 ( new_n337_, new_n336_ );
or g262 ( new_n338_, new_n255_, new_n335_ );
and g263 ( new_n339_, new_n337_, new_n338_ );
or g264 ( new_n340_, new_n339_, new_n119_, N105, new_n156_ );
and g265 ( new_n341_, new_n310_, new_n325_, new_n331_, new_n340_ );
and g266 ( new_n342_, new_n291_, keyIn_0_20, new_n273_, new_n341_ );
not g267 ( new_n343_, new_n342_ );
and g268 ( new_n344_, new_n291_, new_n273_, new_n341_ );
or g269 ( new_n345_, new_n344_, keyIn_0_20 );
and g270 ( new_n346_, new_n345_, new_n343_ );
not g271 ( N370, new_n346_ );
or g272 ( new_n348_, new_n346_, keyIn_0_21 );
and g273 ( new_n349_, new_n345_, keyIn_0_21, new_n343_ );
not g274 ( new_n350_, new_n349_ );
and g275 ( new_n351_, new_n348_, new_n350_ );
not g276 ( new_n352_, new_n351_ );
and g277 ( new_n353_, new_n352_, keyIn_0_22, N40 );
not g278 ( new_n354_, keyIn_0_22 );
not g279 ( new_n355_, N40 );
or g280 ( new_n356_, new_n351_, new_n355_ );
and g281 ( new_n357_, new_n356_, new_n354_ );
and g282 ( new_n358_, N329, N34 );
and g283 ( new_n359_, N223, N24 );
or g284 ( new_n360_, new_n358_, new_n101_, new_n359_ );
or g285 ( new_n361_, new_n357_, new_n353_, new_n360_ );
and g286 ( new_n362_, new_n361_, keyIn_0_24 );
not g287 ( new_n363_, keyIn_0_24 );
not g288 ( new_n364_, new_n353_ );
not g289 ( new_n365_, new_n357_ );
not g290 ( new_n366_, new_n360_ );
and g291 ( new_n367_, new_n365_, new_n363_, new_n364_, new_n366_ );
or g292 ( new_n368_, new_n362_, new_n367_ );
and g293 ( new_n369_, new_n352_, N27 );
and g294 ( new_n370_, N329, N21 );
and g295 ( new_n371_, N223, N11 );
or g296 ( new_n372_, new_n369_, new_n77_, new_n370_, new_n371_ );
and g297 ( new_n373_, new_n368_, new_n372_ );
and g298 ( new_n374_, new_n352_, N66 );
and g299 ( new_n375_, N329, N60 );
and g300 ( new_n376_, N223, N50 );
or g301 ( new_n377_, new_n374_, new_n201_, new_n375_, new_n376_ );
and g302 ( new_n378_, new_n373_, new_n377_ );
not g303 ( new_n379_, keyIn_0_25 );
and g304 ( new_n380_, new_n352_, keyIn_0_23, N53 );
not g305 ( new_n381_, keyIn_0_23 );
not g306 ( new_n382_, N53 );
or g307 ( new_n383_, new_n351_, new_n382_ );
and g308 ( new_n384_, new_n383_, new_n381_ );
and g309 ( new_n385_, N329, N47 );
and g310 ( new_n386_, N223, N37 );
or g311 ( new_n387_, new_n385_, new_n103_, new_n386_ );
or g312 ( new_n388_, new_n384_, new_n380_, new_n387_ );
and g313 ( new_n389_, new_n388_, new_n379_ );
not g314 ( new_n390_, new_n380_ );
not g315 ( new_n391_, new_n384_ );
not g316 ( new_n392_, new_n387_ );
and g317 ( new_n393_, new_n391_, keyIn_0_25, new_n390_, new_n392_ );
or g318 ( new_n394_, new_n389_, new_n393_ );
and g319 ( new_n395_, new_n352_, N79 );
not g320 ( new_n396_, new_n395_ );
and g321 ( new_n397_, N329, N73 );
not g322 ( new_n398_, new_n397_ );
and g323 ( new_n399_, N223, N63 );
not g324 ( new_n400_, new_n399_ );
and g325 ( new_n401_, new_n396_, N69, new_n398_, new_n400_ );
not g326 ( new_n402_, new_n401_ );
and g327 ( new_n403_, new_n352_, N115 );
and g328 ( new_n404_, N329, N112 );
and g329 ( new_n405_, N223, N102 );
or g330 ( new_n406_, new_n403_, new_n207_, new_n404_, new_n405_ );
not g331 ( new_n407_, N105 );
or g332 ( new_n408_, new_n351_, new_n407_ );
and g333 ( new_n409_, N329, N99 );
not g334 ( new_n410_, new_n409_ );
and g335 ( new_n411_, N223, N89 );
not g336 ( new_n412_, new_n411_ );
and g337 ( new_n413_, new_n408_, N95, new_n410_, new_n412_ );
not g338 ( new_n414_, new_n413_ );
and g339 ( new_n415_, new_n352_, N92 );
and g340 ( new_n416_, N329, N86 );
and g341 ( new_n417_, N223, N76 );
or g342 ( new_n418_, new_n415_, new_n214_, new_n416_, new_n417_ );
and g343 ( new_n419_, new_n402_, new_n406_, new_n414_, new_n418_ );
and g344 ( new_n420_, new_n378_, new_n394_, new_n419_ );
not g345 ( new_n421_, new_n420_ );
and g346 ( new_n422_, new_n352_, N14 );
and g347 ( new_n423_, N329, N8 );
and g348 ( new_n424_, N223, N1 );
or g349 ( new_n425_, new_n422_, new_n177_, new_n423_, new_n424_ );
and g350 ( N421, new_n421_, new_n425_ );
not g351 ( new_n427_, keyIn_0_30 );
not g352 ( new_n428_, new_n378_ );
not g353 ( new_n429_, keyIn_0_26 );
not g354 ( new_n430_, new_n389_ );
not g355 ( new_n431_, new_n393_ );
and g356 ( new_n432_, new_n430_, new_n429_, new_n431_ );
and g357 ( new_n433_, new_n394_, keyIn_0_26 );
or g358 ( new_n434_, new_n433_, new_n432_ );
and g359 ( new_n435_, new_n434_, new_n368_ );
not g360 ( new_n436_, new_n435_ );
and g361 ( new_n437_, new_n436_, keyIn_0_27 );
not g362 ( new_n438_, keyIn_0_27 );
and g363 ( new_n439_, new_n435_, new_n438_ );
or g364 ( new_n440_, new_n437_, new_n428_, new_n439_ );
and g365 ( new_n441_, new_n440_, new_n427_ );
or g366 ( new_n442_, new_n435_, new_n438_ );
not g367 ( new_n443_, new_n368_ );
not g368 ( new_n444_, new_n432_ );
not g369 ( new_n445_, new_n433_ );
and g370 ( new_n446_, new_n445_, new_n444_ );
or g371 ( new_n447_, new_n446_, keyIn_0_27, new_n443_ );
and g372 ( new_n448_, new_n442_, keyIn_0_30, new_n378_, new_n447_ );
or g373 ( N430, new_n441_, new_n448_ );
not g374 ( new_n450_, new_n373_ );
not g375 ( new_n451_, keyIn_0_28 );
and g376 ( new_n452_, new_n401_, new_n377_ );
and g377 ( new_n453_, new_n368_, new_n394_, new_n452_ );
not g378 ( new_n454_, new_n453_ );
and g379 ( new_n455_, new_n454_, new_n451_ );
and g380 ( new_n456_, new_n453_, keyIn_0_28 );
or g381 ( new_n457_, new_n455_, new_n456_ );
not g382 ( new_n458_, new_n457_ );
not g383 ( new_n459_, new_n418_ );
and g384 ( new_n460_, new_n394_, new_n377_, new_n459_ );
or g385 ( N431, new_n458_, new_n450_, new_n460_ );
not g386 ( new_n462_, keyIn_0_29 );
and g387 ( new_n463_, new_n418_, new_n413_ );
and g388 ( new_n464_, new_n368_, new_n394_, new_n463_ );
and g389 ( new_n465_, new_n464_, new_n462_ );
not g390 ( new_n466_, new_n465_ );
or g391 ( new_n467_, new_n464_, new_n462_ );
and g392 ( new_n468_, new_n466_, new_n372_, new_n467_ );
and g393 ( new_n469_, new_n442_, new_n447_, new_n457_, new_n468_ );
not g394 ( new_n470_, new_n469_ );
and g395 ( new_n471_, new_n470_, keyIn_0_31 );
not g396 ( new_n472_, keyIn_0_31 );
and g397 ( new_n473_, new_n469_, new_n472_ );
or g398 ( N432, new_n471_, new_n473_ );
endmodule