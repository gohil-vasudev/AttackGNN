module add_mul_comp_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, 
        a_7_, a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, 
        b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, 
        b_13_, b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   Result_9_, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593;
  assign Result_8_ = Result_9_;
  assign Result_6_ = Result_9_;
  assign Result_4_ = Result_9_;
  assign Result_2_ = Result_9_;
  assign Result_15_ = Result_9_;
  assign Result_13_ = Result_9_;
  assign Result_11_ = Result_9_;
  assign Result_0_ = Result_9_;
  assign Result_10_ = Result_9_;
  assign Result_12_ = Result_9_;
  assign Result_14_ = Result_9_;
  assign Result_1_ = Result_9_;
  assign Result_3_ = Result_9_;
  assign Result_5_ = Result_9_;
  assign Result_7_ = Result_9_;

  NOR2_X1 U329 ( .A1(n312), .A2(n313), .ZN(Result_9_) );
  NOR2_X1 U330 ( .A1(n314), .A2(n315), .ZN(n313) );
  INV_X1 U331 ( .A(n316), .ZN(n315) );
  XNOR2_X1 U332 ( .A(n317), .B(a_15_), .ZN(Result_31_) );
  NAND2_X1 U333 ( .A1(n318), .A2(n319), .ZN(Result_30_) );
  NAND2_X1 U334 ( .A1(n320), .A2(n321), .ZN(n319) );
  AND2_X1 U335 ( .A1(n322), .A2(n323), .ZN(n321) );
  NOR2_X1 U336 ( .A1(n324), .A2(n325), .ZN(n320) );
  NAND2_X1 U337 ( .A1(n326), .A2(n327), .ZN(n325) );
  NAND2_X1 U338 ( .A1(b_15_), .A2(n328), .ZN(n327) );
  NAND2_X1 U339 ( .A1(n329), .A2(n317), .ZN(n326) );
  NAND2_X1 U340 ( .A1(n330), .A2(n331), .ZN(n318) );
  XNOR2_X1 U341 ( .A(n332), .B(a_14_), .ZN(n331) );
  NOR2_X1 U342 ( .A1(n333), .A2(n334), .ZN(n330) );
  NOR2_X1 U343 ( .A1(n335), .A2(n336), .ZN(n334) );
  NOR2_X1 U344 ( .A1(n324), .A2(n337), .ZN(n333) );
  NAND2_X1 U345 ( .A1(n328), .A2(n317), .ZN(n337) );
  INV_X1 U346 ( .A(a_15_), .ZN(n324) );
  NAND2_X1 U347 ( .A1(n338), .A2(n339), .ZN(Result_29_) );
  NAND2_X1 U348 ( .A1(n340), .A2(n341), .ZN(n339) );
  XOR2_X1 U349 ( .A(n342), .B(n343), .Z(n341) );
  NAND2_X1 U350 ( .A1(n344), .A2(n335), .ZN(n338) );
  XNOR2_X1 U351 ( .A(n345), .B(n342), .ZN(n344) );
  NAND2_X1 U352 ( .A1(n346), .A2(n347), .ZN(n342) );
  NAND2_X1 U353 ( .A1(n348), .A2(n349), .ZN(Result_28_) );
  NAND2_X1 U354 ( .A1(n340), .A2(n350), .ZN(n349) );
  XNOR2_X1 U355 ( .A(n351), .B(n352), .ZN(n350) );
  NAND2_X1 U356 ( .A1(n353), .A2(n335), .ZN(n348) );
  XOR2_X1 U357 ( .A(n354), .B(n351), .Z(n353) );
  AND2_X1 U358 ( .A1(n355), .A2(n356), .ZN(n351) );
  NAND2_X1 U359 ( .A1(n357), .A2(n358), .ZN(Result_27_) );
  NAND2_X1 U360 ( .A1(n340), .A2(n359), .ZN(n358) );
  XOR2_X1 U361 ( .A(n360), .B(n361), .Z(n359) );
  NAND2_X1 U362 ( .A1(n362), .A2(n335), .ZN(n357) );
  XNOR2_X1 U363 ( .A(n363), .B(n360), .ZN(n362) );
  NAND2_X1 U364 ( .A1(n364), .A2(n365), .ZN(n360) );
  NAND2_X1 U365 ( .A1(n366), .A2(n367), .ZN(Result_26_) );
  NAND2_X1 U366 ( .A1(n340), .A2(n368), .ZN(n367) );
  XNOR2_X1 U367 ( .A(n369), .B(n370), .ZN(n368) );
  NAND2_X1 U368 ( .A1(n371), .A2(n335), .ZN(n366) );
  XOR2_X1 U369 ( .A(n372), .B(n369), .Z(n371) );
  AND2_X1 U370 ( .A1(n373), .A2(n374), .ZN(n369) );
  NAND2_X1 U371 ( .A1(n375), .A2(n376), .ZN(Result_25_) );
  NAND2_X1 U372 ( .A1(n340), .A2(n377), .ZN(n376) );
  XOR2_X1 U373 ( .A(n378), .B(n379), .Z(n377) );
  NAND2_X1 U374 ( .A1(n380), .A2(n335), .ZN(n375) );
  XNOR2_X1 U375 ( .A(n381), .B(n378), .ZN(n380) );
  NAND2_X1 U376 ( .A1(n382), .A2(n383), .ZN(n378) );
  NAND2_X1 U377 ( .A1(n384), .A2(n385), .ZN(Result_24_) );
  NAND2_X1 U378 ( .A1(n340), .A2(n386), .ZN(n385) );
  XNOR2_X1 U379 ( .A(n387), .B(n388), .ZN(n386) );
  NAND2_X1 U380 ( .A1(n389), .A2(n335), .ZN(n384) );
  XOR2_X1 U381 ( .A(n390), .B(n387), .Z(n389) );
  AND2_X1 U382 ( .A1(n391), .A2(n392), .ZN(n387) );
  NAND2_X1 U383 ( .A1(n393), .A2(n394), .ZN(Result_23_) );
  NAND2_X1 U384 ( .A1(n340), .A2(n395), .ZN(n394) );
  XOR2_X1 U385 ( .A(n396), .B(n397), .Z(n395) );
  NAND2_X1 U386 ( .A1(n398), .A2(n335), .ZN(n393) );
  XNOR2_X1 U387 ( .A(n399), .B(n396), .ZN(n398) );
  NAND2_X1 U388 ( .A1(n400), .A2(n401), .ZN(n396) );
  NAND2_X1 U389 ( .A1(n402), .A2(n403), .ZN(Result_22_) );
  NAND2_X1 U390 ( .A1(n340), .A2(n404), .ZN(n403) );
  XNOR2_X1 U391 ( .A(n405), .B(n406), .ZN(n404) );
  NAND2_X1 U392 ( .A1(n407), .A2(n335), .ZN(n402) );
  XOR2_X1 U393 ( .A(n408), .B(n405), .Z(n407) );
  AND2_X1 U394 ( .A1(n409), .A2(n410), .ZN(n405) );
  NAND2_X1 U395 ( .A1(n411), .A2(n412), .ZN(Result_21_) );
  NAND2_X1 U396 ( .A1(n340), .A2(n413), .ZN(n412) );
  XOR2_X1 U397 ( .A(n414), .B(n415), .Z(n413) );
  NAND2_X1 U398 ( .A1(n416), .A2(n335), .ZN(n411) );
  XNOR2_X1 U399 ( .A(n417), .B(n414), .ZN(n416) );
  NAND2_X1 U400 ( .A1(n418), .A2(n419), .ZN(n414) );
  NAND2_X1 U401 ( .A1(n420), .A2(n421), .ZN(Result_20_) );
  NAND2_X1 U402 ( .A1(n340), .A2(n422), .ZN(n421) );
  XNOR2_X1 U403 ( .A(n423), .B(n424), .ZN(n422) );
  NAND2_X1 U404 ( .A1(n425), .A2(n335), .ZN(n420) );
  XOR2_X1 U405 ( .A(n426), .B(n423), .Z(n425) );
  AND2_X1 U406 ( .A1(n427), .A2(n428), .ZN(n423) );
  NAND2_X1 U407 ( .A1(n429), .A2(n430), .ZN(Result_19_) );
  NAND2_X1 U408 ( .A1(n340), .A2(n431), .ZN(n430) );
  XOR2_X1 U409 ( .A(n432), .B(n433), .Z(n431) );
  NAND2_X1 U410 ( .A1(n434), .A2(n335), .ZN(n429) );
  XNOR2_X1 U411 ( .A(n435), .B(n432), .ZN(n434) );
  NAND2_X1 U412 ( .A1(n436), .A2(n437), .ZN(n432) );
  NAND2_X1 U413 ( .A1(n438), .A2(n439), .ZN(Result_18_) );
  NAND2_X1 U414 ( .A1(n340), .A2(n440), .ZN(n439) );
  XNOR2_X1 U415 ( .A(n441), .B(n442), .ZN(n440) );
  NAND2_X1 U416 ( .A1(n443), .A2(n335), .ZN(n438) );
  XOR2_X1 U417 ( .A(n444), .B(n441), .Z(n443) );
  AND2_X1 U418 ( .A1(n445), .A2(n446), .ZN(n441) );
  NAND2_X1 U419 ( .A1(n447), .A2(n448), .ZN(Result_17_) );
  NAND2_X1 U420 ( .A1(n340), .A2(n449), .ZN(n448) );
  XNOR2_X1 U421 ( .A(n450), .B(n451), .ZN(n449) );
  NAND2_X1 U422 ( .A1(n452), .A2(n335), .ZN(n447) );
  XNOR2_X1 U423 ( .A(n453), .B(n454), .ZN(n452) );
  INV_X1 U424 ( .A(n450), .ZN(n454) );
  NOR2_X1 U425 ( .A1(n455), .A2(n456), .ZN(n450) );
  INV_X1 U426 ( .A(n457), .ZN(n456) );
  NAND2_X1 U427 ( .A1(n458), .A2(n459), .ZN(Result_16_) );
  NAND2_X1 U428 ( .A1(n340), .A2(n460), .ZN(n459) );
  XNOR2_X1 U429 ( .A(n461), .B(n462), .ZN(n460) );
  NOR2_X1 U430 ( .A1(n463), .A2(n464), .ZN(n462) );
  AND2_X1 U431 ( .A1(n451), .A2(a_1_), .ZN(n464) );
  NOR2_X1 U432 ( .A1(n465), .A2(n466), .ZN(n463) );
  NOR2_X1 U433 ( .A1(a_1_), .A2(n451), .ZN(n465) );
  NAND2_X1 U434 ( .A1(n467), .A2(n468), .ZN(n451) );
  NAND2_X1 U435 ( .A1(b_2_), .A2(n469), .ZN(n468) );
  OR2_X1 U436 ( .A1(n442), .A2(a_2_), .ZN(n469) );
  NAND2_X1 U437 ( .A1(a_2_), .A2(n442), .ZN(n467) );
  NAND2_X1 U438 ( .A1(n470), .A2(n471), .ZN(n442) );
  NAND2_X1 U439 ( .A1(b_3_), .A2(n472), .ZN(n471) );
  OR2_X1 U440 ( .A1(n433), .A2(a_3_), .ZN(n472) );
  NAND2_X1 U441 ( .A1(a_3_), .A2(n433), .ZN(n470) );
  NAND2_X1 U442 ( .A1(n473), .A2(n474), .ZN(n433) );
  NAND2_X1 U443 ( .A1(b_4_), .A2(n475), .ZN(n474) );
  OR2_X1 U444 ( .A1(n424), .A2(a_4_), .ZN(n475) );
  NAND2_X1 U445 ( .A1(a_4_), .A2(n424), .ZN(n473) );
  NAND2_X1 U446 ( .A1(n476), .A2(n477), .ZN(n424) );
  NAND2_X1 U447 ( .A1(b_5_), .A2(n478), .ZN(n477) );
  OR2_X1 U448 ( .A1(n415), .A2(a_5_), .ZN(n478) );
  NAND2_X1 U449 ( .A1(a_5_), .A2(n415), .ZN(n476) );
  NAND2_X1 U450 ( .A1(n479), .A2(n480), .ZN(n415) );
  NAND2_X1 U451 ( .A1(b_6_), .A2(n481), .ZN(n480) );
  OR2_X1 U452 ( .A1(n406), .A2(a_6_), .ZN(n481) );
  NAND2_X1 U453 ( .A1(a_6_), .A2(n406), .ZN(n479) );
  NAND2_X1 U454 ( .A1(n482), .A2(n483), .ZN(n406) );
  NAND2_X1 U455 ( .A1(b_7_), .A2(n484), .ZN(n483) );
  OR2_X1 U456 ( .A1(n397), .A2(a_7_), .ZN(n484) );
  NAND2_X1 U457 ( .A1(a_7_), .A2(n397), .ZN(n482) );
  NAND2_X1 U458 ( .A1(n485), .A2(n486), .ZN(n397) );
  NAND2_X1 U459 ( .A1(b_8_), .A2(n487), .ZN(n486) );
  OR2_X1 U460 ( .A1(n388), .A2(a_8_), .ZN(n487) );
  NAND2_X1 U461 ( .A1(a_8_), .A2(n388), .ZN(n485) );
  NAND2_X1 U462 ( .A1(n488), .A2(n489), .ZN(n388) );
  NAND2_X1 U463 ( .A1(b_9_), .A2(n490), .ZN(n489) );
  OR2_X1 U464 ( .A1(n379), .A2(a_9_), .ZN(n490) );
  NAND2_X1 U465 ( .A1(a_9_), .A2(n379), .ZN(n488) );
  NAND2_X1 U466 ( .A1(n491), .A2(n492), .ZN(n379) );
  NAND2_X1 U467 ( .A1(b_10_), .A2(n493), .ZN(n492) );
  OR2_X1 U468 ( .A1(n370), .A2(a_10_), .ZN(n493) );
  NAND2_X1 U469 ( .A1(a_10_), .A2(n370), .ZN(n491) );
  NAND2_X1 U470 ( .A1(n494), .A2(n495), .ZN(n370) );
  NAND2_X1 U471 ( .A1(b_11_), .A2(n496), .ZN(n495) );
  OR2_X1 U472 ( .A1(n361), .A2(a_11_), .ZN(n496) );
  NAND2_X1 U473 ( .A1(a_11_), .A2(n361), .ZN(n494) );
  NAND2_X1 U474 ( .A1(n497), .A2(n498), .ZN(n361) );
  NAND2_X1 U475 ( .A1(b_12_), .A2(n499), .ZN(n498) );
  OR2_X1 U476 ( .A1(n352), .A2(a_12_), .ZN(n499) );
  NAND2_X1 U477 ( .A1(a_12_), .A2(n352), .ZN(n497) );
  NAND2_X1 U478 ( .A1(n500), .A2(n501), .ZN(n352) );
  NAND2_X1 U479 ( .A1(b_13_), .A2(n502), .ZN(n501) );
  OR2_X1 U480 ( .A1(n343), .A2(a_13_), .ZN(n502) );
  NAND2_X1 U481 ( .A1(a_13_), .A2(n343), .ZN(n500) );
  NAND2_X1 U482 ( .A1(n503), .A2(n504), .ZN(n343) );
  NAND2_X1 U483 ( .A1(b_14_), .A2(n505), .ZN(n504) );
  NAND2_X1 U484 ( .A1(n506), .A2(n336), .ZN(n505) );
  OR2_X1 U485 ( .A1(n336), .A2(n506), .ZN(n503) );
  INV_X1 U486 ( .A(a_14_), .ZN(n506) );
  NAND2_X1 U487 ( .A1(b_15_), .A2(a_15_), .ZN(n336) );
  INV_X1 U488 ( .A(n328), .ZN(n340) );
  NAND2_X1 U489 ( .A1(n329), .A2(n507), .ZN(n328) );
  NAND2_X1 U490 ( .A1(n508), .A2(n509), .ZN(n507) );
  NOR2_X1 U491 ( .A1(n510), .A2(n511), .ZN(n509) );
  NAND2_X1 U492 ( .A1(n512), .A2(n513), .ZN(n511) );
  NOR2_X1 U493 ( .A1(n514), .A2(n515), .ZN(n513) );
  NOR2_X1 U494 ( .A1(n516), .A2(n517), .ZN(n512) );
  NAND2_X1 U495 ( .A1(n518), .A2(n519), .ZN(n510) );
  NOR2_X1 U496 ( .A1(n455), .A2(n520), .ZN(n519) );
  NOR2_X1 U497 ( .A1(n521), .A2(n312), .ZN(n518) );
  NOR2_X1 U498 ( .A1(n522), .A2(n523), .ZN(n508) );
  NAND2_X1 U499 ( .A1(n524), .A2(n525), .ZN(n523) );
  NOR2_X1 U500 ( .A1(n526), .A2(n527), .ZN(n525) );
  NOR2_X1 U501 ( .A1(n528), .A2(n529), .ZN(n524) );
  NOR2_X1 U502 ( .A1(a_15_), .A2(n317), .ZN(n529) );
  NAND2_X1 U503 ( .A1(n530), .A2(n531), .ZN(n522) );
  NOR2_X1 U504 ( .A1(n532), .A2(n533), .ZN(n531) );
  NOR2_X1 U505 ( .A1(n534), .A2(n535), .ZN(n530) );
  INV_X1 U506 ( .A(n335), .ZN(n329) );
  NAND2_X1 U507 ( .A1(n536), .A2(n335), .ZN(n458) );
  NAND2_X1 U508 ( .A1(n316), .A2(n537), .ZN(n335) );
  NAND2_X1 U509 ( .A1(n538), .A2(n539), .ZN(n537) );
  NAND2_X1 U510 ( .A1(n457), .A2(n540), .ZN(n538) );
  NAND2_X1 U511 ( .A1(n541), .A2(n542), .ZN(n540) );
  NAND2_X1 U512 ( .A1(n543), .A2(n437), .ZN(n542) );
  NOR2_X1 U513 ( .A1(n544), .A2(n545), .ZN(n543) );
  AND2_X1 U514 ( .A1(n546), .A2(a_2_), .ZN(n545) );
  NOR2_X1 U515 ( .A1(n547), .A2(n548), .ZN(n544) );
  NAND2_X1 U516 ( .A1(n427), .A2(n436), .ZN(n548) );
  NOR2_X1 U517 ( .A1(n549), .A2(n550), .ZN(n547) );
  NAND2_X1 U518 ( .A1(n428), .A2(n551), .ZN(n550) );
  NAND2_X1 U519 ( .A1(n552), .A2(n553), .ZN(n551) );
  NAND2_X1 U520 ( .A1(n554), .A2(n401), .ZN(n553) );
  NOR2_X1 U521 ( .A1(n555), .A2(n556), .ZN(n554) );
  AND2_X1 U522 ( .A1(n557), .A2(a_6_), .ZN(n556) );
  NOR2_X1 U523 ( .A1(n558), .A2(n559), .ZN(n555) );
  NAND2_X1 U524 ( .A1(n391), .A2(n400), .ZN(n559) );
  NOR2_X1 U525 ( .A1(n560), .A2(n561), .ZN(n558) );
  NAND2_X1 U526 ( .A1(n392), .A2(n562), .ZN(n561) );
  NAND2_X1 U527 ( .A1(n563), .A2(n564), .ZN(n562) );
  NAND2_X1 U528 ( .A1(n565), .A2(n365), .ZN(n564) );
  NOR2_X1 U529 ( .A1(n566), .A2(n567), .ZN(n565) );
  AND2_X1 U530 ( .A1(n568), .A2(a_10_), .ZN(n567) );
  NOR2_X1 U531 ( .A1(n527), .A2(n363), .ZN(n566) );
  NOR2_X1 U532 ( .A1(n535), .A2(n526), .ZN(n563) );
  AND2_X1 U533 ( .A1(n569), .A2(a_9_), .ZN(n560) );
  NOR2_X1 U534 ( .A1(n517), .A2(n532), .ZN(n552) );
  AND2_X1 U535 ( .A1(n570), .A2(a_5_), .ZN(n549) );
  NOR2_X1 U536 ( .A1(n455), .A2(n514), .ZN(n541) );
  NAND2_X1 U537 ( .A1(n314), .A2(n461), .ZN(n536) );
  NAND2_X1 U538 ( .A1(n539), .A2(n316), .ZN(n461) );
  NAND2_X1 U539 ( .A1(a_0_), .A2(n571), .ZN(n316) );
  INV_X1 U540 ( .A(n312), .ZN(n539) );
  NOR2_X1 U541 ( .A1(n571), .A2(a_0_), .ZN(n312) );
  INV_X1 U542 ( .A(b_0_), .ZN(n571) );
  NOR2_X1 U543 ( .A1(n455), .A2(n572), .ZN(n314) );
  AND2_X1 U544 ( .A1(n453), .A2(n457), .ZN(n572) );
  NAND2_X1 U545 ( .A1(a_1_), .A2(n466), .ZN(n457) );
  NAND2_X1 U546 ( .A1(n445), .A2(n573), .ZN(n453) );
  NAND2_X1 U547 ( .A1(n446), .A2(n444), .ZN(n573) );
  NAND2_X1 U548 ( .A1(n436), .A2(n574), .ZN(n444) );
  NAND2_X1 U549 ( .A1(n437), .A2(n435), .ZN(n574) );
  NAND2_X1 U550 ( .A1(n427), .A2(n575), .ZN(n435) );
  NAND2_X1 U551 ( .A1(n428), .A2(n426), .ZN(n575) );
  NAND2_X1 U552 ( .A1(n418), .A2(n576), .ZN(n426) );
  NAND2_X1 U553 ( .A1(n419), .A2(n417), .ZN(n576) );
  NAND2_X1 U554 ( .A1(n409), .A2(n577), .ZN(n417) );
  NAND2_X1 U555 ( .A1(n410), .A2(n408), .ZN(n577) );
  NAND2_X1 U556 ( .A1(n400), .A2(n578), .ZN(n408) );
  NAND2_X1 U557 ( .A1(n401), .A2(n399), .ZN(n578) );
  NAND2_X1 U558 ( .A1(n391), .A2(n579), .ZN(n399) );
  NAND2_X1 U559 ( .A1(n392), .A2(n390), .ZN(n579) );
  NAND2_X1 U560 ( .A1(n382), .A2(n580), .ZN(n390) );
  NAND2_X1 U561 ( .A1(n383), .A2(n381), .ZN(n580) );
  NAND2_X1 U562 ( .A1(n373), .A2(n581), .ZN(n381) );
  NAND2_X1 U563 ( .A1(n374), .A2(n372), .ZN(n581) );
  NAND2_X1 U564 ( .A1(n364), .A2(n582), .ZN(n372) );
  NAND2_X1 U565 ( .A1(n365), .A2(n363), .ZN(n582) );
  NAND2_X1 U566 ( .A1(n355), .A2(n583), .ZN(n363) );
  NAND2_X1 U567 ( .A1(n356), .A2(n354), .ZN(n583) );
  NAND2_X1 U568 ( .A1(n346), .A2(n584), .ZN(n354) );
  NAND2_X1 U569 ( .A1(n347), .A2(n345), .ZN(n584) );
  NAND2_X1 U570 ( .A1(n322), .A2(n585), .ZN(n345) );
  NAND2_X1 U571 ( .A1(n586), .A2(n323), .ZN(n585) );
  NAND2_X1 U572 ( .A1(a_14_), .A2(n332), .ZN(n323) );
  NAND2_X1 U573 ( .A1(a_15_), .A2(n317), .ZN(n586) );
  INV_X1 U574 ( .A(b_15_), .ZN(n317) );
  INV_X1 U575 ( .A(n520), .ZN(n322) );
  NOR2_X1 U576 ( .A1(n332), .A2(a_14_), .ZN(n520) );
  INV_X1 U577 ( .A(b_14_), .ZN(n332) );
  NAND2_X1 U578 ( .A1(a_13_), .A2(n587), .ZN(n347) );
  INV_X1 U579 ( .A(n521), .ZN(n346) );
  NOR2_X1 U580 ( .A1(n587), .A2(a_13_), .ZN(n521) );
  INV_X1 U581 ( .A(b_13_), .ZN(n587) );
  NAND2_X1 U582 ( .A1(a_12_), .A2(n588), .ZN(n356) );
  INV_X1 U583 ( .A(n528), .ZN(n355) );
  NOR2_X1 U584 ( .A1(n588), .A2(a_12_), .ZN(n528) );
  INV_X1 U585 ( .A(b_12_), .ZN(n588) );
  NAND2_X1 U586 ( .A1(a_11_), .A2(n589), .ZN(n365) );
  INV_X1 U587 ( .A(n527), .ZN(n364) );
  NOR2_X1 U588 ( .A1(n589), .A2(a_11_), .ZN(n527) );
  INV_X1 U589 ( .A(b_11_), .ZN(n589) );
  NAND2_X1 U590 ( .A1(a_10_), .A2(n568), .ZN(n374) );
  INV_X1 U591 ( .A(n526), .ZN(n373) );
  NOR2_X1 U592 ( .A1(n568), .A2(a_10_), .ZN(n526) );
  INV_X1 U593 ( .A(b_10_), .ZN(n568) );
  NAND2_X1 U594 ( .A1(a_9_), .A2(n569), .ZN(n383) );
  INV_X1 U595 ( .A(n535), .ZN(n382) );
  NOR2_X1 U596 ( .A1(n569), .A2(a_9_), .ZN(n535) );
  INV_X1 U597 ( .A(b_9_), .ZN(n569) );
  NAND2_X1 U598 ( .A1(a_8_), .A2(n590), .ZN(n392) );
  INV_X1 U599 ( .A(n534), .ZN(n391) );
  NOR2_X1 U600 ( .A1(n590), .A2(a_8_), .ZN(n534) );
  INV_X1 U601 ( .A(b_8_), .ZN(n590) );
  NAND2_X1 U602 ( .A1(a_7_), .A2(n591), .ZN(n401) );
  INV_X1 U603 ( .A(n533), .ZN(n400) );
  NOR2_X1 U604 ( .A1(n591), .A2(a_7_), .ZN(n533) );
  INV_X1 U605 ( .A(b_7_), .ZN(n591) );
  NAND2_X1 U606 ( .A1(a_6_), .A2(n557), .ZN(n410) );
  INV_X1 U607 ( .A(n532), .ZN(n409) );
  NOR2_X1 U608 ( .A1(n557), .A2(a_6_), .ZN(n532) );
  INV_X1 U609 ( .A(b_6_), .ZN(n557) );
  NAND2_X1 U610 ( .A1(a_5_), .A2(n570), .ZN(n419) );
  INV_X1 U611 ( .A(n517), .ZN(n418) );
  NOR2_X1 U612 ( .A1(n570), .A2(a_5_), .ZN(n517) );
  INV_X1 U613 ( .A(b_5_), .ZN(n570) );
  NAND2_X1 U614 ( .A1(a_4_), .A2(n592), .ZN(n428) );
  INV_X1 U615 ( .A(n516), .ZN(n427) );
  NOR2_X1 U616 ( .A1(n592), .A2(a_4_), .ZN(n516) );
  INV_X1 U617 ( .A(b_4_), .ZN(n592) );
  NAND2_X1 U618 ( .A1(a_3_), .A2(n593), .ZN(n437) );
  INV_X1 U619 ( .A(n515), .ZN(n436) );
  NOR2_X1 U620 ( .A1(n593), .A2(a_3_), .ZN(n515) );
  INV_X1 U621 ( .A(b_3_), .ZN(n593) );
  NAND2_X1 U622 ( .A1(a_2_), .A2(n546), .ZN(n446) );
  INV_X1 U623 ( .A(n514), .ZN(n445) );
  NOR2_X1 U624 ( .A1(n546), .A2(a_2_), .ZN(n514) );
  INV_X1 U625 ( .A(b_2_), .ZN(n546) );
  NOR2_X1 U626 ( .A1(n466), .A2(a_1_), .ZN(n455) );
  INV_X1 U627 ( .A(b_1_), .ZN(n466) );
endmodule

