module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n153_, new_n701_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n878_, new_n543_, new_n113_, new_n886_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n789_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n881_, new_n319_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, N93 );
and g001 ( new_n107_, new_n106_, N89 );
not g002 ( new_n108_, N89 );
and g003 ( new_n109_, new_n108_, N93 );
or g004 ( new_n110_, new_n107_, new_n109_ );
not g005 ( new_n111_, new_n110_ );
not g006 ( new_n112_, N85 );
and g007 ( new_n113_, new_n112_, N81 );
not g008 ( new_n114_, N81 );
and g009 ( new_n115_, new_n114_, N85 );
or g010 ( new_n116_, new_n113_, new_n115_ );
and g011 ( new_n117_, new_n111_, new_n116_ );
not g012 ( new_n118_, new_n116_ );
and g013 ( new_n119_, new_n118_, new_n110_ );
or g014 ( new_n120_, new_n117_, new_n119_ );
not g015 ( new_n121_, new_n120_ );
not g016 ( new_n122_, N77 );
and g017 ( new_n123_, new_n122_, N73 );
not g018 ( new_n124_, N73 );
and g019 ( new_n125_, new_n124_, N77 );
or g020 ( new_n126_, new_n123_, new_n125_ );
not g021 ( new_n127_, new_n126_ );
not g022 ( new_n128_, N69 );
and g023 ( new_n129_, new_n128_, N65 );
not g024 ( new_n130_, N65 );
and g025 ( new_n131_, new_n130_, N69 );
or g026 ( new_n132_, new_n129_, new_n131_ );
and g027 ( new_n133_, new_n127_, new_n132_ );
not g028 ( new_n134_, new_n132_ );
and g029 ( new_n135_, new_n134_, new_n126_ );
or g030 ( new_n136_, new_n133_, new_n135_ );
and g031 ( new_n137_, new_n121_, new_n136_ );
not g032 ( new_n138_, new_n136_ );
and g033 ( new_n139_, new_n138_, new_n120_ );
or g034 ( new_n140_, new_n137_, new_n139_ );
not g035 ( new_n141_, new_n140_ );
and g036 ( new_n142_, N129, N137 );
and g037 ( new_n143_, new_n141_, new_n142_ );
not g038 ( new_n144_, new_n143_ );
or g039 ( new_n145_, new_n141_, new_n142_ );
and g040 ( new_n146_, new_n144_, new_n145_ );
not g041 ( new_n147_, N49 );
and g042 ( new_n148_, new_n147_, N33 );
not g043 ( new_n149_, N33 );
and g044 ( new_n150_, new_n149_, N49 );
or g045 ( new_n151_, new_n148_, new_n150_ );
not g046 ( new_n152_, new_n151_ );
not g047 ( new_n153_, N17 );
and g048 ( new_n154_, new_n153_, N1 );
not g049 ( new_n155_, N1 );
and g050 ( new_n156_, new_n155_, N17 );
or g051 ( new_n157_, new_n154_, new_n156_ );
and g052 ( new_n158_, new_n152_, new_n157_ );
not g053 ( new_n159_, new_n158_ );
or g054 ( new_n160_, new_n152_, new_n157_ );
and g055 ( new_n161_, new_n159_, new_n160_ );
and g056 ( new_n162_, new_n161_, keyIn_0_9 );
not g057 ( new_n163_, new_n162_ );
or g058 ( new_n164_, new_n161_, keyIn_0_9 );
and g059 ( new_n165_, new_n163_, new_n164_ );
or g060 ( new_n166_, new_n146_, new_n165_ );
not g061 ( new_n167_, new_n166_ );
and g062 ( new_n168_, new_n146_, new_n165_ );
or g063 ( new_n169_, new_n167_, new_n168_ );
not g064 ( new_n170_, N117 );
and g065 ( new_n171_, new_n170_, N113 );
not g066 ( new_n172_, N113 );
and g067 ( new_n173_, new_n172_, N117 );
or g068 ( new_n174_, new_n171_, new_n173_ );
and g069 ( new_n175_, new_n174_, keyIn_0_4 );
not g070 ( new_n176_, new_n175_ );
or g071 ( new_n177_, new_n174_, keyIn_0_4 );
and g072 ( new_n178_, new_n176_, new_n177_ );
not g073 ( new_n179_, N125 );
and g074 ( new_n180_, new_n179_, N121 );
not g075 ( new_n181_, N121 );
and g076 ( new_n182_, new_n181_, N125 );
or g077 ( new_n183_, new_n180_, new_n182_ );
not g078 ( new_n184_, new_n183_ );
and g079 ( new_n185_, new_n178_, new_n184_ );
not g080 ( new_n186_, new_n185_ );
or g081 ( new_n187_, new_n178_, new_n184_ );
and g082 ( new_n188_, new_n186_, new_n187_ );
not g083 ( new_n189_, new_n188_ );
not g084 ( new_n190_, N109 );
and g085 ( new_n191_, new_n190_, N105 );
not g086 ( new_n192_, N105 );
and g087 ( new_n193_, new_n192_, N109 );
or g088 ( new_n194_, new_n191_, new_n193_ );
and g089 ( new_n195_, new_n194_, keyIn_0_3 );
not g090 ( new_n196_, new_n195_ );
or g091 ( new_n197_, new_n194_, keyIn_0_3 );
and g092 ( new_n198_, new_n196_, new_n197_ );
not g093 ( new_n199_, N101 );
and g094 ( new_n200_, new_n199_, N97 );
not g095 ( new_n201_, N97 );
and g096 ( new_n202_, new_n201_, N101 );
or g097 ( new_n203_, new_n200_, new_n202_ );
and g098 ( new_n204_, new_n198_, new_n203_ );
not g099 ( new_n205_, new_n204_ );
or g100 ( new_n206_, new_n198_, new_n203_ );
and g101 ( new_n207_, new_n205_, new_n206_ );
and g102 ( new_n208_, new_n189_, new_n207_ );
not g103 ( new_n209_, new_n207_ );
and g104 ( new_n210_, new_n209_, new_n188_ );
or g105 ( new_n211_, new_n208_, new_n210_ );
not g106 ( new_n212_, new_n211_ );
and g107 ( new_n213_, N130, N137 );
and g108 ( new_n214_, new_n212_, new_n213_ );
not g109 ( new_n215_, new_n214_ );
or g110 ( new_n216_, new_n212_, new_n213_ );
and g111 ( new_n217_, new_n215_, new_n216_ );
not g112 ( new_n218_, new_n217_ );
not g113 ( new_n219_, N53 );
and g114 ( new_n220_, new_n219_, N37 );
not g115 ( new_n221_, N37 );
and g116 ( new_n222_, new_n221_, N53 );
or g117 ( new_n223_, new_n220_, new_n222_ );
not g118 ( new_n224_, new_n223_ );
not g119 ( new_n225_, N21 );
and g120 ( new_n226_, new_n225_, N5 );
not g121 ( new_n227_, N5 );
and g122 ( new_n228_, new_n227_, N21 );
or g123 ( new_n229_, new_n226_, new_n228_ );
and g124 ( new_n230_, new_n224_, new_n229_ );
not g125 ( new_n231_, new_n230_ );
or g126 ( new_n232_, new_n224_, new_n229_ );
and g127 ( new_n233_, new_n231_, new_n232_ );
and g128 ( new_n234_, new_n218_, new_n233_ );
not g129 ( new_n235_, new_n233_ );
and g130 ( new_n236_, new_n217_, new_n235_ );
or g131 ( new_n237_, new_n234_, new_n236_ );
and g132 ( new_n238_, new_n209_, new_n138_ );
and g133 ( new_n239_, new_n207_, new_n136_ );
or g134 ( new_n240_, new_n238_, new_n239_ );
not g135 ( new_n241_, new_n240_ );
and g136 ( new_n242_, N131, N137 );
and g137 ( new_n243_, new_n241_, new_n242_ );
not g138 ( new_n244_, new_n243_ );
or g139 ( new_n245_, new_n241_, new_n242_ );
and g140 ( new_n246_, new_n244_, new_n245_ );
not g141 ( new_n247_, N57 );
and g142 ( new_n248_, new_n247_, N41 );
not g143 ( new_n249_, N41 );
and g144 ( new_n250_, new_n249_, N57 );
or g145 ( new_n251_, new_n248_, new_n250_ );
not g146 ( new_n252_, new_n251_ );
and g147 ( new_n253_, new_n252_, keyIn_0_6 );
not g148 ( new_n254_, new_n253_ );
or g149 ( new_n255_, new_n252_, keyIn_0_6 );
and g150 ( new_n256_, new_n254_, new_n255_ );
not g151 ( new_n257_, new_n256_ );
not g152 ( new_n258_, N25 );
and g153 ( new_n259_, new_n258_, N9 );
not g154 ( new_n260_, N9 );
and g155 ( new_n261_, new_n260_, N25 );
or g156 ( new_n262_, new_n259_, new_n261_ );
and g157 ( new_n263_, new_n257_, new_n262_ );
not g158 ( new_n264_, new_n263_ );
or g159 ( new_n265_, new_n257_, new_n262_ );
and g160 ( new_n266_, new_n264_, new_n265_ );
not g161 ( new_n267_, new_n266_ );
or g162 ( new_n268_, new_n246_, new_n267_ );
not g163 ( new_n269_, new_n268_ );
and g164 ( new_n270_, new_n246_, new_n267_ );
or g165 ( new_n271_, new_n269_, new_n270_ );
and g166 ( new_n272_, new_n271_, keyIn_0_12 );
and g167 ( new_n273_, new_n272_, new_n237_ );
not g168 ( new_n274_, new_n273_ );
or g169 ( new_n275_, new_n272_, new_n237_ );
not g170 ( new_n276_, new_n168_ );
and g171 ( new_n277_, new_n276_, new_n166_ );
and g172 ( new_n278_, new_n189_, new_n121_ );
and g173 ( new_n279_, new_n188_, new_n120_ );
or g174 ( new_n280_, new_n278_, new_n279_ );
not g175 ( new_n281_, new_n280_ );
and g176 ( new_n282_, N132, N137 );
and g177 ( new_n283_, new_n281_, new_n282_ );
not g178 ( new_n284_, new_n283_ );
or g179 ( new_n285_, new_n281_, new_n282_ );
and g180 ( new_n286_, new_n284_, new_n285_ );
not g181 ( new_n287_, N61 );
and g182 ( new_n288_, new_n287_, N45 );
not g183 ( new_n289_, N45 );
and g184 ( new_n290_, new_n289_, N61 );
or g185 ( new_n291_, new_n288_, new_n290_ );
not g186 ( new_n292_, new_n291_ );
not g187 ( new_n293_, N29 );
and g188 ( new_n294_, new_n293_, N13 );
not g189 ( new_n295_, N13 );
and g190 ( new_n296_, new_n295_, N29 );
or g191 ( new_n297_, new_n294_, new_n296_ );
and g192 ( new_n298_, new_n292_, new_n297_ );
not g193 ( new_n299_, new_n298_ );
or g194 ( new_n300_, new_n292_, new_n297_ );
and g195 ( new_n301_, new_n299_, new_n300_ );
not g196 ( new_n302_, new_n301_ );
and g197 ( new_n303_, new_n286_, new_n302_ );
not g198 ( new_n304_, new_n303_ );
or g199 ( new_n305_, new_n286_, new_n302_ );
and g200 ( new_n306_, new_n304_, new_n305_ );
and g201 ( new_n307_, new_n306_, new_n277_ );
and g202 ( new_n308_, new_n275_, new_n307_ );
and g203 ( new_n309_, new_n308_, new_n274_ );
or g204 ( new_n310_, new_n271_, new_n306_ );
and g205 ( new_n311_, new_n169_, keyIn_0_11 );
not g206 ( new_n312_, keyIn_0_11 );
and g207 ( new_n313_, new_n277_, new_n312_ );
or g208 ( new_n314_, new_n311_, new_n313_ );
or g209 ( new_n315_, new_n237_, new_n314_ );
or g210 ( new_n316_, new_n315_, new_n310_ );
or g211 ( new_n317_, new_n316_, keyIn_0_19 );
not g212 ( new_n318_, keyIn_0_19 );
not g213 ( new_n319_, new_n270_ );
and g214 ( new_n320_, new_n319_, new_n268_ );
not g215 ( new_n321_, new_n305_ );
or g216 ( new_n322_, new_n321_, new_n303_ );
and g217 ( new_n323_, new_n322_, new_n320_ );
or g218 ( new_n324_, new_n217_, new_n235_ );
not g219 ( new_n325_, new_n236_ );
and g220 ( new_n326_, new_n325_, new_n324_ );
or g221 ( new_n327_, new_n277_, new_n312_ );
not g222 ( new_n328_, new_n313_ );
and g223 ( new_n329_, new_n328_, new_n327_ );
and g224 ( new_n330_, new_n329_, new_n326_ );
and g225 ( new_n331_, new_n330_, new_n323_ );
or g226 ( new_n332_, new_n331_, new_n318_ );
and g227 ( new_n333_, new_n317_, new_n332_ );
and g228 ( new_n334_, new_n237_, keyIn_0_13 );
not g229 ( new_n335_, new_n334_ );
or g230 ( new_n336_, new_n237_, keyIn_0_13 );
and g231 ( new_n337_, new_n335_, new_n336_ );
not g232 ( new_n338_, new_n337_ );
and g233 ( new_n339_, new_n320_, new_n169_ );
and g234 ( new_n340_, new_n339_, new_n306_ );
and g235 ( new_n341_, new_n338_, new_n340_ );
or g236 ( new_n342_, new_n333_, new_n341_ );
or g237 ( new_n343_, new_n342_, new_n309_ );
not g238 ( new_n344_, keyIn_0_10 );
and g239 ( new_n345_, new_n287_, N57 );
and g240 ( new_n346_, new_n247_, N61 );
or g241 ( new_n347_, new_n345_, new_n346_ );
not g242 ( new_n348_, new_n347_ );
and g243 ( new_n349_, new_n219_, N49 );
and g244 ( new_n350_, new_n147_, N53 );
or g245 ( new_n351_, new_n349_, new_n350_ );
and g246 ( new_n352_, new_n348_, new_n351_ );
not g247 ( new_n353_, new_n352_ );
or g248 ( new_n354_, new_n348_, new_n351_ );
and g249 ( new_n355_, new_n353_, new_n354_ );
and g250 ( new_n356_, new_n225_, N17 );
and g251 ( new_n357_, new_n153_, N21 );
or g252 ( new_n358_, new_n356_, new_n357_ );
and g253 ( new_n359_, new_n358_, keyIn_0_0 );
not g254 ( new_n360_, keyIn_0_0 );
or g255 ( new_n361_, new_n153_, N21 );
or g256 ( new_n362_, new_n225_, N17 );
and g257 ( new_n363_, new_n361_, new_n362_ );
and g258 ( new_n364_, new_n363_, new_n360_ );
or g259 ( new_n365_, new_n359_, new_n364_ );
and g260 ( new_n366_, new_n293_, N25 );
and g261 ( new_n367_, new_n258_, N29 );
or g262 ( new_n368_, new_n366_, new_n367_ );
not g263 ( new_n369_, new_n368_ );
and g264 ( new_n370_, new_n365_, new_n369_ );
or g265 ( new_n371_, new_n363_, new_n360_ );
or g266 ( new_n372_, new_n358_, keyIn_0_0 );
and g267 ( new_n373_, new_n372_, new_n371_ );
and g268 ( new_n374_, new_n373_, new_n368_ );
or g269 ( new_n375_, new_n370_, new_n374_ );
and g270 ( new_n376_, new_n375_, new_n355_ );
not g271 ( new_n377_, new_n355_ );
or g272 ( new_n378_, new_n373_, new_n368_ );
or g273 ( new_n379_, new_n365_, new_n369_ );
and g274 ( new_n380_, new_n379_, new_n378_ );
and g275 ( new_n381_, new_n380_, new_n377_ );
or g276 ( new_n382_, new_n376_, new_n381_ );
and g277 ( new_n383_, N136, N137 );
not g278 ( new_n384_, new_n383_ );
and g279 ( new_n385_, new_n382_, new_n384_ );
or g280 ( new_n386_, new_n380_, new_n377_ );
or g281 ( new_n387_, new_n375_, new_n355_ );
and g282 ( new_n388_, new_n387_, new_n386_ );
and g283 ( new_n389_, new_n388_, new_n383_ );
or g284 ( new_n390_, new_n385_, new_n389_ );
and g285 ( new_n391_, new_n390_, new_n344_ );
or g286 ( new_n392_, new_n388_, new_n383_ );
or g287 ( new_n393_, new_n382_, new_n384_ );
and g288 ( new_n394_, new_n393_, new_n392_ );
and g289 ( new_n395_, new_n394_, keyIn_0_10 );
or g290 ( new_n396_, new_n391_, new_n395_ );
and g291 ( new_n397_, new_n179_, N109 );
and g292 ( new_n398_, new_n190_, N125 );
or g293 ( new_n399_, new_n397_, new_n398_ );
not g294 ( new_n400_, new_n399_ );
and g295 ( new_n401_, new_n106_, N77 );
and g296 ( new_n402_, new_n122_, N93 );
or g297 ( new_n403_, new_n401_, new_n402_ );
and g298 ( new_n404_, new_n400_, new_n403_ );
not g299 ( new_n405_, new_n404_ );
or g300 ( new_n406_, new_n400_, new_n403_ );
and g301 ( new_n407_, new_n405_, new_n406_ );
or g302 ( new_n408_, new_n396_, new_n407_ );
or g303 ( new_n409_, new_n394_, keyIn_0_10 );
or g304 ( new_n410_, new_n390_, new_n344_ );
and g305 ( new_n411_, new_n410_, new_n409_ );
not g306 ( new_n412_, new_n407_ );
or g307 ( new_n413_, new_n411_, new_n412_ );
and g308 ( new_n414_, new_n408_, new_n413_ );
and g309 ( new_n415_, new_n414_, keyIn_0_15 );
not g310 ( new_n416_, new_n415_ );
or g311 ( new_n417_, new_n414_, keyIn_0_15 );
and g312 ( new_n418_, new_n416_, new_n417_ );
not g313 ( new_n419_, new_n418_ );
not g314 ( new_n420_, keyIn_0_14 );
not g315 ( new_n421_, keyIn_0_8 );
not g316 ( new_n422_, keyIn_0_1 );
or g317 ( new_n423_, new_n149_, N37 );
or g318 ( new_n424_, new_n221_, N33 );
and g319 ( new_n425_, new_n423_, new_n424_ );
or g320 ( new_n426_, new_n425_, new_n422_ );
and g321 ( new_n427_, new_n221_, N33 );
and g322 ( new_n428_, new_n149_, N37 );
or g323 ( new_n429_, new_n427_, new_n428_ );
or g324 ( new_n430_, new_n429_, keyIn_0_1 );
and g325 ( new_n431_, new_n430_, new_n426_ );
not g326 ( new_n432_, keyIn_0_2 );
or g327 ( new_n433_, new_n249_, N45 );
or g328 ( new_n434_, new_n289_, N41 );
and g329 ( new_n435_, new_n433_, new_n434_ );
and g330 ( new_n436_, new_n435_, new_n432_ );
and g331 ( new_n437_, new_n289_, N41 );
and g332 ( new_n438_, new_n249_, N45 );
or g333 ( new_n439_, new_n437_, new_n438_ );
and g334 ( new_n440_, new_n439_, keyIn_0_2 );
or g335 ( new_n441_, new_n440_, new_n436_ );
and g336 ( new_n442_, new_n441_, new_n431_ );
and g337 ( new_n443_, new_n429_, keyIn_0_1 );
and g338 ( new_n444_, new_n425_, new_n422_ );
or g339 ( new_n445_, new_n443_, new_n444_ );
or g340 ( new_n446_, new_n439_, keyIn_0_2 );
or g341 ( new_n447_, new_n435_, new_n432_ );
and g342 ( new_n448_, new_n446_, new_n447_ );
and g343 ( new_n449_, new_n445_, new_n448_ );
or g344 ( new_n450_, new_n442_, new_n449_ );
or g345 ( new_n451_, new_n450_, new_n421_ );
or g346 ( new_n452_, new_n445_, new_n448_ );
or g347 ( new_n453_, new_n441_, new_n431_ );
and g348 ( new_n454_, new_n452_, new_n453_ );
or g349 ( new_n455_, new_n454_, keyIn_0_8 );
and g350 ( new_n456_, new_n451_, new_n455_ );
or g351 ( new_n457_, new_n456_, new_n355_ );
and g352 ( new_n458_, new_n454_, keyIn_0_8 );
and g353 ( new_n459_, new_n450_, new_n421_ );
or g354 ( new_n460_, new_n458_, new_n459_ );
or g355 ( new_n461_, new_n460_, new_n377_ );
and g356 ( new_n462_, new_n461_, new_n457_ );
and g357 ( new_n463_, N134, N137 );
or g358 ( new_n464_, new_n462_, new_n463_ );
and g359 ( new_n465_, new_n460_, new_n377_ );
and g360 ( new_n466_, new_n456_, new_n355_ );
or g361 ( new_n467_, new_n465_, new_n466_ );
not g362 ( new_n468_, new_n463_ );
or g363 ( new_n469_, new_n467_, new_n468_ );
and g364 ( new_n470_, new_n469_, new_n464_ );
and g365 ( new_n471_, new_n170_, N101 );
and g366 ( new_n472_, new_n199_, N117 );
or g367 ( new_n473_, new_n471_, new_n472_ );
not g368 ( new_n474_, new_n473_ );
and g369 ( new_n475_, new_n112_, N69 );
and g370 ( new_n476_, new_n128_, N85 );
or g371 ( new_n477_, new_n475_, new_n476_ );
and g372 ( new_n478_, new_n474_, new_n477_ );
not g373 ( new_n479_, new_n478_ );
or g374 ( new_n480_, new_n474_, new_n477_ );
and g375 ( new_n481_, new_n479_, new_n480_ );
not g376 ( new_n482_, new_n481_ );
or g377 ( new_n483_, new_n470_, new_n482_ );
and g378 ( new_n484_, new_n467_, new_n468_ );
and g379 ( new_n485_, new_n462_, new_n463_ );
or g380 ( new_n486_, new_n484_, new_n485_ );
or g381 ( new_n487_, new_n486_, new_n481_ );
and g382 ( new_n488_, new_n487_, new_n483_ );
and g383 ( new_n489_, new_n488_, new_n420_ );
not g384 ( new_n490_, new_n489_ );
and g385 ( new_n491_, new_n486_, new_n481_ );
and g386 ( new_n492_, new_n470_, new_n482_ );
or g387 ( new_n493_, new_n491_, new_n492_ );
and g388 ( new_n494_, new_n493_, keyIn_0_14 );
not g389 ( new_n495_, new_n494_ );
and g390 ( new_n496_, new_n295_, N9 );
and g391 ( new_n497_, new_n260_, N13 );
or g392 ( new_n498_, new_n496_, new_n497_ );
not g393 ( new_n499_, new_n498_ );
and g394 ( new_n500_, new_n227_, N1 );
and g395 ( new_n501_, new_n155_, N5 );
or g396 ( new_n502_, new_n500_, new_n501_ );
and g397 ( new_n503_, new_n499_, new_n502_ );
not g398 ( new_n504_, new_n503_ );
or g399 ( new_n505_, new_n499_, new_n502_ );
and g400 ( new_n506_, new_n504_, new_n505_ );
not g401 ( new_n507_, new_n506_ );
and g402 ( new_n508_, new_n460_, new_n507_ );
and g403 ( new_n509_, new_n456_, new_n506_ );
or g404 ( new_n510_, new_n508_, new_n509_ );
and g405 ( new_n511_, N135, N137 );
and g406 ( new_n512_, new_n511_, keyIn_0_5 );
not g407 ( new_n513_, new_n512_ );
or g408 ( new_n514_, new_n511_, keyIn_0_5 );
and g409 ( new_n515_, new_n513_, new_n514_ );
not g410 ( new_n516_, new_n515_ );
and g411 ( new_n517_, new_n510_, new_n516_ );
or g412 ( new_n518_, new_n456_, new_n506_ );
or g413 ( new_n519_, new_n460_, new_n507_ );
and g414 ( new_n520_, new_n519_, new_n518_ );
and g415 ( new_n521_, new_n520_, new_n515_ );
or g416 ( new_n522_, new_n517_, new_n521_ );
and g417 ( new_n523_, new_n181_, N105 );
and g418 ( new_n524_, new_n192_, N121 );
or g419 ( new_n525_, new_n523_, new_n524_ );
not g420 ( new_n526_, new_n525_ );
and g421 ( new_n527_, new_n526_, keyIn_0_7 );
not g422 ( new_n528_, new_n527_ );
or g423 ( new_n529_, new_n526_, keyIn_0_7 );
and g424 ( new_n530_, new_n528_, new_n529_ );
not g425 ( new_n531_, new_n530_ );
and g426 ( new_n532_, new_n108_, N73 );
and g427 ( new_n533_, new_n124_, N89 );
or g428 ( new_n534_, new_n532_, new_n533_ );
and g429 ( new_n535_, new_n531_, new_n534_ );
not g430 ( new_n536_, new_n535_ );
or g431 ( new_n537_, new_n531_, new_n534_ );
and g432 ( new_n538_, new_n536_, new_n537_ );
and g433 ( new_n539_, new_n522_, new_n538_ );
or g434 ( new_n540_, new_n520_, new_n515_ );
or g435 ( new_n541_, new_n510_, new_n516_ );
and g436 ( new_n542_, new_n541_, new_n540_ );
not g437 ( new_n543_, new_n538_ );
and g438 ( new_n544_, new_n542_, new_n543_ );
or g439 ( new_n545_, new_n539_, new_n544_ );
and g440 ( new_n546_, new_n375_, new_n506_ );
and g441 ( new_n547_, new_n380_, new_n507_ );
or g442 ( new_n548_, new_n546_, new_n547_ );
and g443 ( new_n549_, N133, N137 );
not g444 ( new_n550_, new_n549_ );
and g445 ( new_n551_, new_n548_, new_n550_ );
not g446 ( new_n552_, new_n551_ );
or g447 ( new_n553_, new_n548_, new_n550_ );
and g448 ( new_n554_, new_n552_, new_n553_ );
not g449 ( new_n555_, new_n554_ );
and g450 ( new_n556_, new_n172_, N97 );
and g451 ( new_n557_, new_n201_, N113 );
or g452 ( new_n558_, new_n556_, new_n557_ );
not g453 ( new_n559_, new_n558_ );
and g454 ( new_n560_, new_n114_, N65 );
and g455 ( new_n561_, new_n130_, N81 );
or g456 ( new_n562_, new_n560_, new_n561_ );
and g457 ( new_n563_, new_n559_, new_n562_ );
not g458 ( new_n564_, new_n563_ );
or g459 ( new_n565_, new_n559_, new_n562_ );
and g460 ( new_n566_, new_n564_, new_n565_ );
and g461 ( new_n567_, new_n555_, new_n566_ );
not g462 ( new_n568_, new_n566_ );
and g463 ( new_n569_, new_n554_, new_n568_ );
or g464 ( new_n570_, new_n567_, new_n569_ );
and g465 ( new_n571_, new_n545_, new_n570_ );
and g466 ( new_n572_, new_n495_, new_n571_ );
and g467 ( new_n573_, new_n572_, new_n490_ );
and g468 ( new_n574_, new_n573_, new_n419_ );
and g469 ( new_n575_, new_n343_, new_n574_ );
or g470 ( new_n576_, new_n575_, keyIn_0_24 );
not g471 ( new_n577_, keyIn_0_24 );
not g472 ( new_n578_, new_n309_ );
and g473 ( new_n579_, new_n331_, new_n318_ );
and g474 ( new_n580_, new_n316_, keyIn_0_19 );
or g475 ( new_n581_, new_n580_, new_n579_ );
not g476 ( new_n582_, new_n341_ );
and g477 ( new_n583_, new_n581_, new_n582_ );
and g478 ( new_n584_, new_n583_, new_n578_ );
not g479 ( new_n585_, new_n574_ );
or g480 ( new_n586_, new_n584_, new_n585_ );
or g481 ( new_n587_, new_n586_, new_n577_ );
and g482 ( new_n588_, new_n576_, new_n587_ );
and g483 ( new_n589_, new_n588_, new_n169_ );
not g484 ( new_n590_, new_n589_ );
and g485 ( new_n591_, new_n590_, N1 );
and g486 ( new_n592_, new_n589_, new_n155_ );
or g487 ( N724, new_n591_, new_n592_ );
and g488 ( new_n594_, new_n588_, new_n237_ );
not g489 ( new_n595_, new_n594_ );
and g490 ( new_n596_, new_n595_, N5 );
and g491 ( new_n597_, new_n594_, new_n227_ );
or g492 ( N725, new_n596_, new_n597_ );
not g493 ( new_n599_, keyIn_0_30 );
and g494 ( new_n600_, new_n586_, new_n577_ );
and g495 ( new_n601_, new_n575_, keyIn_0_24 );
or g496 ( new_n602_, new_n601_, new_n600_ );
or g497 ( new_n603_, new_n602_, new_n320_ );
and g498 ( new_n604_, new_n603_, N9 );
and g499 ( new_n605_, new_n588_, new_n271_ );
and g500 ( new_n606_, new_n605_, new_n260_ );
or g501 ( new_n607_, new_n604_, new_n606_ );
or g502 ( new_n608_, new_n607_, new_n599_ );
or g503 ( new_n609_, new_n605_, new_n260_ );
or g504 ( new_n610_, new_n603_, N9 );
and g505 ( new_n611_, new_n610_, new_n609_ );
or g506 ( new_n612_, new_n611_, keyIn_0_30 );
and g507 ( N726, new_n608_, new_n612_ );
or g508 ( new_n614_, new_n602_, new_n306_ );
and g509 ( new_n615_, new_n614_, N13 );
and g510 ( new_n616_, new_n588_, new_n322_ );
and g511 ( new_n617_, new_n616_, new_n295_ );
or g512 ( new_n618_, new_n615_, new_n617_ );
and g513 ( new_n619_, new_n618_, keyIn_0_31 );
not g514 ( new_n620_, keyIn_0_31 );
or g515 ( new_n621_, new_n616_, new_n295_ );
or g516 ( new_n622_, new_n614_, N13 );
and g517 ( new_n623_, new_n622_, new_n621_ );
and g518 ( new_n624_, new_n623_, new_n620_ );
or g519 ( N727, new_n619_, new_n624_ );
and g520 ( new_n626_, new_n488_, new_n570_ );
and g521 ( new_n627_, new_n411_, new_n412_ );
and g522 ( new_n628_, new_n396_, new_n407_ );
or g523 ( new_n629_, new_n628_, new_n627_ );
or g524 ( new_n630_, new_n542_, new_n543_ );
or g525 ( new_n631_, new_n522_, new_n538_ );
and g526 ( new_n632_, new_n631_, new_n630_ );
and g527 ( new_n633_, new_n632_, new_n629_ );
and g528 ( new_n634_, new_n626_, new_n633_ );
and g529 ( new_n635_, new_n343_, new_n634_ );
and g530 ( new_n636_, new_n635_, new_n169_ );
not g531 ( new_n637_, new_n636_ );
and g532 ( new_n638_, new_n637_, N17 );
and g533 ( new_n639_, new_n636_, new_n153_ );
or g534 ( N728, new_n638_, new_n639_ );
and g535 ( new_n641_, new_n635_, new_n237_ );
not g536 ( new_n642_, new_n641_ );
and g537 ( new_n643_, new_n642_, N21 );
and g538 ( new_n644_, new_n641_, new_n225_ );
or g539 ( N729, new_n643_, new_n644_ );
and g540 ( new_n646_, new_n635_, new_n271_ );
and g541 ( new_n647_, new_n646_, keyIn_0_25 );
not g542 ( new_n648_, new_n647_ );
or g543 ( new_n649_, new_n646_, keyIn_0_25 );
and g544 ( new_n650_, new_n648_, new_n649_ );
not g545 ( new_n651_, new_n650_ );
and g546 ( new_n652_, new_n651_, N25 );
and g547 ( new_n653_, new_n650_, new_n258_ );
or g548 ( N730, new_n652_, new_n653_ );
and g549 ( new_n655_, new_n635_, new_n322_ );
not g550 ( new_n656_, new_n655_ );
and g551 ( new_n657_, new_n656_, keyIn_0_26 );
not g552 ( new_n658_, new_n657_ );
or g553 ( new_n659_, new_n656_, keyIn_0_26 );
and g554 ( new_n660_, new_n658_, new_n659_ );
not g555 ( new_n661_, new_n660_ );
and g556 ( new_n662_, new_n661_, N29 );
and g557 ( new_n663_, new_n660_, new_n293_ );
or g558 ( N731, new_n662_, new_n663_ );
or g559 ( new_n665_, new_n632_, new_n629_ );
not g560 ( new_n666_, new_n570_ );
and g561 ( new_n667_, new_n666_, keyIn_0_16 );
not g562 ( new_n668_, new_n667_ );
or g563 ( new_n669_, new_n666_, keyIn_0_16 );
and g564 ( new_n670_, new_n668_, new_n669_ );
or g565 ( new_n671_, new_n670_, new_n488_ );
or g566 ( new_n672_, new_n671_, new_n665_ );
or g567 ( new_n673_, new_n584_, new_n672_ );
not g568 ( new_n674_, new_n673_ );
and g569 ( new_n675_, new_n674_, new_n169_ );
not g570 ( new_n676_, new_n675_ );
and g571 ( new_n677_, new_n676_, N33 );
and g572 ( new_n678_, new_n675_, new_n149_ );
or g573 ( N732, new_n677_, new_n678_ );
and g574 ( new_n680_, new_n674_, new_n237_ );
not g575 ( new_n681_, new_n680_ );
and g576 ( new_n682_, new_n681_, N37 );
and g577 ( new_n683_, new_n680_, new_n221_ );
or g578 ( N733, new_n682_, new_n683_ );
and g579 ( new_n685_, new_n674_, new_n271_ );
not g580 ( new_n686_, new_n685_ );
and g581 ( new_n687_, new_n686_, N41 );
and g582 ( new_n688_, new_n685_, new_n249_ );
or g583 ( N734, new_n687_, new_n688_ );
and g584 ( new_n690_, new_n674_, new_n322_ );
not g585 ( new_n691_, new_n690_ );
and g586 ( new_n692_, new_n691_, N45 );
and g587 ( new_n693_, new_n690_, new_n289_ );
or g588 ( N735, new_n692_, new_n693_ );
and g589 ( new_n695_, new_n666_, keyIn_0_17 );
not g590 ( new_n696_, new_n695_ );
or g591 ( new_n697_, new_n666_, keyIn_0_17 );
and g592 ( new_n698_, new_n696_, new_n697_ );
and g593 ( new_n699_, new_n698_, new_n493_ );
and g594 ( new_n700_, new_n699_, new_n633_ );
and g595 ( new_n701_, new_n343_, new_n700_ );
and g596 ( new_n702_, new_n701_, new_n169_ );
not g597 ( new_n703_, new_n702_ );
and g598 ( new_n704_, new_n703_, N49 );
and g599 ( new_n705_, new_n702_, new_n147_ );
or g600 ( N736, new_n704_, new_n705_ );
and g601 ( new_n707_, new_n701_, new_n237_ );
not g602 ( new_n708_, new_n707_ );
and g603 ( new_n709_, new_n708_, N53 );
and g604 ( new_n710_, new_n707_, new_n219_ );
or g605 ( N737, new_n709_, new_n710_ );
and g606 ( new_n712_, new_n701_, new_n271_ );
not g607 ( new_n713_, new_n712_ );
and g608 ( new_n714_, new_n713_, N57 );
and g609 ( new_n715_, new_n712_, new_n247_ );
or g610 ( N738, new_n714_, new_n715_ );
and g611 ( new_n717_, new_n701_, new_n322_ );
not g612 ( new_n718_, new_n717_ );
and g613 ( new_n719_, new_n718_, N61 );
and g614 ( new_n720_, new_n717_, new_n287_ );
or g615 ( N739, new_n719_, new_n720_ );
or g616 ( new_n722_, new_n545_, new_n414_ );
or g617 ( new_n723_, new_n493_, new_n570_ );
or g618 ( new_n724_, new_n722_, new_n723_ );
and g619 ( new_n725_, new_n724_, keyIn_0_20 );
not g620 ( new_n726_, keyIn_0_20 );
and g621 ( new_n727_, new_n488_, new_n666_ );
and g622 ( new_n728_, new_n633_, new_n727_ );
and g623 ( new_n729_, new_n728_, new_n726_ );
or g624 ( new_n730_, new_n725_, new_n729_ );
and g625 ( new_n731_, new_n626_, new_n414_ );
and g626 ( new_n732_, new_n545_, keyIn_0_18 );
not g627 ( new_n733_, new_n732_ );
or g628 ( new_n734_, new_n545_, keyIn_0_18 );
and g629 ( new_n735_, new_n733_, new_n734_ );
and g630 ( new_n736_, new_n735_, new_n731_ );
not g631 ( new_n737_, new_n736_ );
and g632 ( new_n738_, new_n730_, new_n737_ );
or g633 ( new_n739_, new_n665_, new_n723_ );
and g634 ( new_n740_, new_n739_, keyIn_0_21 );
not g635 ( new_n741_, keyIn_0_21 );
and g636 ( new_n742_, new_n545_, new_n414_ );
and g637 ( new_n743_, new_n742_, new_n727_ );
and g638 ( new_n744_, new_n743_, new_n741_ );
or g639 ( new_n745_, new_n740_, new_n744_ );
or g640 ( new_n746_, new_n488_, new_n570_ );
or g641 ( new_n747_, new_n545_, new_n629_ );
or g642 ( new_n748_, new_n747_, new_n746_ );
and g643 ( new_n749_, new_n748_, keyIn_0_22 );
not g644 ( new_n750_, keyIn_0_22 );
and g645 ( new_n751_, new_n493_, new_n666_ );
and g646 ( new_n752_, new_n632_, new_n414_ );
and g647 ( new_n753_, new_n751_, new_n752_ );
and g648 ( new_n754_, new_n753_, new_n750_ );
or g649 ( new_n755_, new_n749_, new_n754_ );
and g650 ( new_n756_, new_n745_, new_n755_ );
and g651 ( new_n757_, new_n738_, new_n756_ );
and g652 ( new_n758_, new_n757_, keyIn_0_23 );
not g653 ( new_n759_, new_n758_ );
or g654 ( new_n760_, new_n757_, keyIn_0_23 );
and g655 ( new_n761_, new_n759_, new_n760_ );
and g656 ( new_n762_, new_n271_, new_n306_ );
and g657 ( new_n763_, new_n326_, new_n169_ );
and g658 ( new_n764_, new_n762_, new_n763_ );
and g659 ( new_n765_, new_n761_, new_n764_ );
and g660 ( new_n766_, new_n765_, new_n570_ );
not g661 ( new_n767_, new_n766_ );
and g662 ( new_n768_, new_n767_, N65 );
and g663 ( new_n769_, new_n766_, new_n130_ );
or g664 ( N740, new_n768_, new_n769_ );
and g665 ( new_n771_, new_n765_, new_n493_ );
not g666 ( new_n772_, new_n771_ );
and g667 ( new_n773_, new_n772_, N69 );
and g668 ( new_n774_, new_n771_, new_n128_ );
or g669 ( N741, new_n773_, new_n774_ );
and g670 ( new_n776_, new_n765_, new_n545_ );
not g671 ( new_n777_, new_n776_ );
and g672 ( new_n778_, new_n777_, N73 );
and g673 ( new_n779_, new_n776_, new_n124_ );
or g674 ( N742, new_n778_, new_n779_ );
and g675 ( new_n781_, new_n765_, new_n629_ );
not g676 ( new_n782_, new_n781_ );
and g677 ( new_n783_, new_n782_, N77 );
and g678 ( new_n784_, new_n781_, new_n122_ );
or g679 ( N743, new_n783_, new_n784_ );
and g680 ( new_n786_, new_n323_, new_n763_ );
and g681 ( new_n787_, new_n761_, new_n786_ );
and g682 ( new_n788_, new_n787_, new_n570_ );
not g683 ( new_n789_, new_n788_ );
and g684 ( new_n790_, new_n789_, N81 );
and g685 ( new_n791_, new_n788_, new_n114_ );
or g686 ( N744, new_n790_, new_n791_ );
not g687 ( new_n793_, keyIn_0_27 );
not g688 ( new_n794_, keyIn_0_23 );
or g689 ( new_n795_, new_n728_, new_n726_ );
or g690 ( new_n796_, new_n724_, keyIn_0_20 );
and g691 ( new_n797_, new_n796_, new_n795_ );
or g692 ( new_n798_, new_n797_, new_n736_ );
or g693 ( new_n799_, new_n743_, new_n741_ );
not g694 ( new_n800_, new_n744_ );
and g695 ( new_n801_, new_n800_, new_n799_ );
or g696 ( new_n802_, new_n753_, new_n750_ );
or g697 ( new_n803_, new_n748_, keyIn_0_22 );
and g698 ( new_n804_, new_n803_, new_n802_ );
or g699 ( new_n805_, new_n801_, new_n804_ );
or g700 ( new_n806_, new_n805_, new_n798_ );
and g701 ( new_n807_, new_n806_, new_n794_ );
or g702 ( new_n808_, new_n807_, new_n758_ );
not g703 ( new_n809_, new_n786_ );
or g704 ( new_n810_, new_n808_, new_n809_ );
or g705 ( new_n811_, new_n810_, new_n488_ );
or g706 ( new_n812_, new_n811_, new_n793_ );
and g707 ( new_n813_, new_n787_, new_n493_ );
or g708 ( new_n814_, new_n813_, keyIn_0_27 );
and g709 ( new_n815_, new_n812_, new_n814_ );
and g710 ( new_n816_, new_n815_, N85 );
and g711 ( new_n817_, new_n813_, keyIn_0_27 );
and g712 ( new_n818_, new_n811_, new_n793_ );
or g713 ( new_n819_, new_n818_, new_n817_ );
and g714 ( new_n820_, new_n819_, new_n112_ );
or g715 ( N745, new_n816_, new_n820_ );
and g716 ( new_n822_, new_n787_, new_n545_ );
not g717 ( new_n823_, new_n822_ );
and g718 ( new_n824_, new_n823_, N89 );
and g719 ( new_n825_, new_n822_, new_n108_ );
or g720 ( N746, new_n824_, new_n825_ );
and g721 ( new_n827_, new_n787_, new_n629_ );
not g722 ( new_n828_, new_n827_ );
and g723 ( new_n829_, new_n828_, N93 );
and g724 ( new_n830_, new_n827_, new_n106_ );
or g725 ( N747, new_n829_, new_n830_ );
and g726 ( new_n832_, new_n237_, new_n277_ );
and g727 ( new_n833_, new_n832_, new_n762_ );
and g728 ( new_n834_, new_n761_, new_n833_ );
and g729 ( new_n835_, new_n834_, new_n570_ );
not g730 ( new_n836_, new_n835_ );
and g731 ( new_n837_, new_n836_, N97 );
and g732 ( new_n838_, new_n835_, new_n201_ );
or g733 ( N748, new_n837_, new_n838_ );
and g734 ( new_n840_, new_n834_, new_n493_ );
not g735 ( new_n841_, new_n840_ );
and g736 ( new_n842_, new_n841_, N101 );
and g737 ( new_n843_, new_n840_, new_n199_ );
or g738 ( N749, new_n842_, new_n843_ );
and g739 ( new_n845_, new_n834_, new_n545_ );
not g740 ( new_n846_, new_n845_ );
and g741 ( new_n847_, new_n846_, N105 );
and g742 ( new_n848_, new_n845_, new_n192_ );
or g743 ( N750, new_n847_, new_n848_ );
not g744 ( new_n850_, new_n833_ );
or g745 ( new_n851_, new_n808_, new_n850_ );
or g746 ( new_n852_, new_n851_, new_n414_ );
or g747 ( new_n853_, new_n852_, keyIn_0_28 );
not g748 ( new_n854_, keyIn_0_28 );
and g749 ( new_n855_, new_n834_, new_n629_ );
or g750 ( new_n856_, new_n855_, new_n854_ );
and g751 ( new_n857_, new_n853_, new_n856_ );
and g752 ( new_n858_, new_n857_, N109 );
and g753 ( new_n859_, new_n855_, new_n854_ );
and g754 ( new_n860_, new_n852_, keyIn_0_28 );
or g755 ( new_n861_, new_n860_, new_n859_ );
and g756 ( new_n862_, new_n861_, new_n190_ );
or g757 ( N751, new_n858_, new_n862_ );
and g758 ( new_n864_, new_n832_, new_n323_ );
and g759 ( new_n865_, new_n761_, new_n864_ );
and g760 ( new_n866_, new_n865_, new_n570_ );
not g761 ( new_n867_, new_n866_ );
and g762 ( new_n868_, new_n867_, N113 );
and g763 ( new_n869_, new_n866_, new_n172_ );
or g764 ( N752, new_n868_, new_n869_ );
not g765 ( new_n871_, new_n864_ );
or g766 ( new_n872_, new_n808_, new_n871_ );
or g767 ( new_n873_, new_n872_, new_n488_ );
and g768 ( new_n874_, new_n873_, keyIn_0_29 );
not g769 ( new_n875_, keyIn_0_29 );
and g770 ( new_n876_, new_n865_, new_n493_ );
and g771 ( new_n877_, new_n876_, new_n875_ );
or g772 ( new_n878_, new_n874_, new_n877_ );
and g773 ( new_n879_, new_n878_, N117 );
or g774 ( new_n880_, new_n876_, new_n875_ );
or g775 ( new_n881_, new_n873_, keyIn_0_29 );
and g776 ( new_n882_, new_n881_, new_n880_ );
and g777 ( new_n883_, new_n882_, new_n170_ );
or g778 ( N753, new_n879_, new_n883_ );
and g779 ( new_n885_, new_n865_, new_n545_ );
not g780 ( new_n886_, new_n885_ );
and g781 ( new_n887_, new_n886_, N121 );
and g782 ( new_n888_, new_n885_, new_n181_ );
or g783 ( N754, new_n887_, new_n888_ );
and g784 ( new_n890_, new_n865_, new_n629_ );
not g785 ( new_n891_, new_n890_ );
and g786 ( new_n892_, new_n891_, N125 );
and g787 ( new_n893_, new_n890_, new_n179_ );
or g788 ( N755, new_n892_, new_n893_ );
endmodule