module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n888_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n777_, new_n720_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n641_, new_n339_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n630_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n961_, new_n890_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n498_, new_n496_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n302_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n837_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n852_, new_n307_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n226_, new_n802_, new_n697_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n947_, new_n994_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n618_, new_n521_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n202_, keyIn_0_60 );
not g001 ( new_n203_, N93 );
nand g002 ( new_n204_, new_n203_, N89 );
not g003 ( new_n205_, N89 );
nand g004 ( new_n206_, new_n205_, N93 );
nand g005 ( new_n207_, new_n204_, new_n206_ );
nand g006 ( new_n208_, new_n207_, keyIn_0_10 );
not g007 ( new_n209_, keyIn_0_10 );
xnor g008 ( new_n210_, N89, N93 );
nand g009 ( new_n211_, new_n210_, new_n209_ );
nand g010 ( new_n212_, new_n208_, new_n211_ );
not g011 ( new_n213_, keyIn_0_11 );
xnor g012 ( new_n214_, N81, N85 );
xnor g013 ( new_n215_, new_n214_, new_n213_ );
nand g014 ( new_n216_, new_n215_, new_n212_ );
xnor g015 ( new_n217_, new_n210_, keyIn_0_10 );
xnor g016 ( new_n218_, new_n214_, keyIn_0_11 );
nand g017 ( new_n219_, new_n217_, new_n218_ );
nand g018 ( new_n220_, new_n219_, new_n216_ );
xnor g019 ( new_n221_, new_n220_, keyIn_0_45 );
not g020 ( new_n222_, keyIn_0_44 );
xnor g021 ( new_n223_, N73, N77 );
xnor g022 ( new_n224_, new_n223_, keyIn_0_9 );
xnor g023 ( new_n225_, N65, N69 );
xnor g024 ( new_n226_, new_n225_, keyIn_0_8 );
nand g025 ( new_n227_, new_n224_, new_n226_ );
not g026 ( new_n228_, keyIn_0_9 );
xnor g027 ( new_n229_, new_n223_, new_n228_ );
not g028 ( new_n230_, keyIn_0_8 );
xnor g029 ( new_n231_, new_n225_, new_n230_ );
nand g030 ( new_n232_, new_n229_, new_n231_ );
nand g031 ( new_n233_, new_n227_, new_n232_ );
xnor g032 ( new_n234_, new_n233_, new_n222_ );
nand g033 ( new_n235_, new_n234_, new_n221_ );
xnor g034 ( new_n236_, new_n218_, new_n212_ );
nand g035 ( new_n237_, new_n236_, keyIn_0_45 );
not g036 ( new_n238_, keyIn_0_45 );
nand g037 ( new_n239_, new_n220_, new_n238_ );
nand g038 ( new_n240_, new_n237_, new_n239_ );
xnor g039 ( new_n241_, new_n233_, keyIn_0_44 );
nand g040 ( new_n242_, new_n241_, new_n240_ );
nand g041 ( new_n243_, new_n235_, new_n242_ );
nand g042 ( new_n244_, new_n243_, new_n202_ );
xnor g043 ( new_n245_, new_n234_, new_n240_ );
nand g044 ( new_n246_, new_n245_, keyIn_0_60 );
nand g045 ( new_n247_, new_n246_, new_n244_ );
nand g046 ( new_n248_, N129, N137 );
xor g047 ( new_n249_, new_n248_, keyIn_0_16 );
nand g048 ( new_n250_, new_n247_, new_n249_ );
xnor g049 ( new_n251_, new_n243_, keyIn_0_60 );
not g050 ( new_n252_, new_n249_ );
nand g051 ( new_n253_, new_n251_, new_n252_ );
nand g052 ( new_n254_, new_n253_, new_n250_ );
nand g053 ( new_n255_, new_n254_, keyIn_0_64 );
not g054 ( new_n256_, keyIn_0_64 );
xnor g055 ( new_n257_, new_n247_, new_n252_ );
nand g056 ( new_n258_, new_n257_, new_n256_ );
nand g057 ( new_n259_, new_n258_, new_n255_ );
xor g058 ( new_n260_, N33, N49 );
xnor g059 ( new_n261_, new_n260_, keyIn_0_25 );
xnor g060 ( new_n262_, N1, N17 );
xnor g061 ( new_n263_, new_n262_, keyIn_0_24 );
xnor g062 ( new_n264_, new_n261_, new_n263_ );
xnor g063 ( new_n265_, new_n264_, keyIn_0_48 );
not g064 ( new_n266_, new_n265_ );
nand g065 ( new_n267_, new_n259_, new_n266_ );
xnor g066 ( new_n268_, new_n254_, new_n256_ );
nand g067 ( new_n269_, new_n268_, new_n265_ );
nand g068 ( new_n270_, new_n269_, new_n267_ );
xnor g069 ( new_n271_, new_n270_, keyIn_0_72 );
not g070 ( new_n272_, keyIn_0_106 );
nor g071 ( new_n273_, new_n271_, keyIn_0_86 );
not g072 ( new_n274_, keyIn_0_87 );
not g073 ( new_n275_, keyIn_0_74 );
not g074 ( new_n276_, keyIn_0_46 );
xnor g075 ( new_n277_, N97, N101 );
xnor g076 ( new_n278_, new_n277_, keyIn_0_12 );
xnor g077 ( new_n279_, N105, N109 );
nand g078 ( new_n280_, new_n279_, keyIn_0_13 );
not g079 ( new_n281_, keyIn_0_13 );
xor g080 ( new_n282_, N105, N109 );
nand g081 ( new_n283_, new_n282_, new_n281_ );
nand g082 ( new_n284_, new_n283_, new_n280_ );
xnor g083 ( new_n285_, new_n278_, new_n284_ );
nand g084 ( new_n286_, new_n285_, new_n276_ );
not g085 ( new_n287_, keyIn_0_12 );
xnor g086 ( new_n288_, new_n277_, new_n287_ );
nand g087 ( new_n289_, new_n288_, new_n284_ );
xnor g088 ( new_n290_, new_n279_, new_n281_ );
nand g089 ( new_n291_, new_n278_, new_n290_ );
nand g090 ( new_n292_, new_n291_, new_n289_ );
nand g091 ( new_n293_, new_n292_, keyIn_0_46 );
nand g092 ( new_n294_, new_n286_, new_n293_ );
xnor g093 ( new_n295_, new_n241_, new_n294_ );
nand g094 ( new_n296_, new_n295_, keyIn_0_62 );
not g095 ( new_n297_, keyIn_0_62 );
xnor g096 ( new_n298_, new_n292_, new_n276_ );
nand g097 ( new_n299_, new_n241_, new_n298_ );
nand g098 ( new_n300_, new_n234_, new_n294_ );
nand g099 ( new_n301_, new_n299_, new_n300_ );
nand g100 ( new_n302_, new_n301_, new_n297_ );
nand g101 ( new_n303_, new_n296_, new_n302_ );
nand g102 ( new_n304_, N131, N137 );
xnor g103 ( new_n305_, new_n304_, keyIn_0_18 );
nand g104 ( new_n306_, new_n303_, new_n305_ );
xnor g105 ( new_n307_, new_n301_, keyIn_0_62 );
not g106 ( new_n308_, new_n305_ );
nand g107 ( new_n309_, new_n307_, new_n308_ );
nand g108 ( new_n310_, new_n309_, new_n306_ );
nand g109 ( new_n311_, new_n310_, keyIn_0_66 );
not g110 ( new_n312_, keyIn_0_66 );
xnor g111 ( new_n313_, new_n303_, new_n308_ );
nand g112 ( new_n314_, new_n313_, new_n312_ );
nand g113 ( new_n315_, new_n314_, new_n311_ );
xor g114 ( new_n316_, N9, N25 );
xnor g115 ( new_n317_, new_n316_, keyIn_0_28 );
xor g116 ( new_n318_, N41, N57 );
xnor g117 ( new_n319_, new_n318_, keyIn_0_29 );
xnor g118 ( new_n320_, new_n317_, new_n319_ );
xor g119 ( new_n321_, new_n320_, keyIn_0_50 );
not g120 ( new_n322_, new_n321_ );
xnor g121 ( new_n323_, new_n315_, new_n322_ );
nand g122 ( new_n324_, new_n323_, new_n275_ );
nand g123 ( new_n325_, new_n315_, new_n321_ );
xnor g124 ( new_n326_, new_n310_, new_n312_ );
nand g125 ( new_n327_, new_n326_, new_n322_ );
nand g126 ( new_n328_, new_n327_, new_n325_ );
nand g127 ( new_n329_, new_n328_, keyIn_0_74 );
nand g128 ( new_n330_, new_n324_, new_n329_ );
nand g129 ( new_n331_, new_n330_, new_n274_ );
nand g130 ( new_n332_, new_n271_, keyIn_0_86 );
nand g131 ( new_n333_, new_n332_, new_n331_ );
nor g132 ( new_n334_, new_n333_, new_n273_ );
not g133 ( new_n335_, keyIn_0_67 );
xnor g134 ( new_n336_, N121, N125 );
xnor g135 ( new_n337_, new_n336_, keyIn_0_15 );
xnor g136 ( new_n338_, N113, N117 );
nand g137 ( new_n339_, new_n338_, keyIn_0_14 );
not g138 ( new_n340_, keyIn_0_14 );
xor g139 ( new_n341_, N113, N117 );
nand g140 ( new_n342_, new_n341_, new_n340_ );
nand g141 ( new_n343_, new_n342_, new_n339_ );
nand g142 ( new_n344_, new_n337_, new_n343_ );
not g143 ( new_n345_, keyIn_0_15 );
xnor g144 ( new_n346_, new_n336_, new_n345_ );
xnor g145 ( new_n347_, new_n338_, new_n340_ );
nand g146 ( new_n348_, new_n346_, new_n347_ );
nand g147 ( new_n349_, new_n348_, new_n344_ );
nand g148 ( new_n350_, new_n349_, keyIn_0_47 );
not g149 ( new_n351_, keyIn_0_47 );
xnor g150 ( new_n352_, new_n346_, new_n343_ );
nand g151 ( new_n353_, new_n352_, new_n351_ );
nand g152 ( new_n354_, new_n353_, new_n350_ );
nand g153 ( new_n355_, new_n354_, new_n221_ );
xnor g154 ( new_n356_, new_n349_, new_n351_ );
nand g155 ( new_n357_, new_n356_, new_n240_ );
nand g156 ( new_n358_, new_n355_, new_n357_ );
nand g157 ( new_n359_, new_n358_, keyIn_0_63 );
not g158 ( new_n360_, keyIn_0_63 );
xnor g159 ( new_n361_, new_n354_, new_n240_ );
nand g160 ( new_n362_, new_n361_, new_n360_ );
nand g161 ( new_n363_, new_n362_, new_n359_ );
nand g162 ( new_n364_, N132, N137 );
xnor g163 ( new_n365_, new_n364_, keyIn_0_19 );
not g164 ( new_n366_, new_n365_ );
nand g165 ( new_n367_, new_n363_, new_n366_ );
xnor g166 ( new_n368_, new_n358_, new_n360_ );
nand g167 ( new_n369_, new_n368_, new_n365_ );
nand g168 ( new_n370_, new_n369_, new_n367_ );
nand g169 ( new_n371_, new_n370_, new_n335_ );
xnor g170 ( new_n372_, new_n363_, new_n365_ );
nand g171 ( new_n373_, new_n372_, keyIn_0_67 );
nand g172 ( new_n374_, new_n373_, new_n371_ );
xor g173 ( new_n375_, N13, N29 );
xnor g174 ( new_n376_, new_n375_, keyIn_0_30 );
xnor g175 ( new_n377_, N45, N61 );
xnor g176 ( new_n378_, new_n377_, keyIn_0_31 );
xnor g177 ( new_n379_, new_n376_, new_n378_ );
xor g178 ( new_n380_, new_n379_, keyIn_0_51 );
not g179 ( new_n381_, new_n380_ );
nand g180 ( new_n382_, new_n374_, new_n381_ );
xnor g181 ( new_n383_, new_n370_, keyIn_0_67 );
nand g182 ( new_n384_, new_n383_, new_n380_ );
nand g183 ( new_n385_, new_n384_, new_n382_ );
nand g184 ( new_n386_, new_n385_, keyIn_0_75 );
not g185 ( new_n387_, keyIn_0_75 );
xnor g186 ( new_n388_, new_n374_, new_n380_ );
nand g187 ( new_n389_, new_n388_, new_n387_ );
nand g188 ( new_n390_, new_n389_, new_n386_ );
nand g189 ( new_n391_, new_n390_, keyIn_0_88 );
not g190 ( new_n392_, keyIn_0_61 );
nand g191 ( new_n393_, new_n298_, new_n354_ );
nand g192 ( new_n394_, new_n356_, new_n294_ );
nand g193 ( new_n395_, new_n393_, new_n394_ );
nand g194 ( new_n396_, new_n395_, new_n392_ );
xnor g195 ( new_n397_, new_n294_, new_n354_ );
nand g196 ( new_n398_, new_n397_, keyIn_0_61 );
nand g197 ( new_n399_, new_n398_, new_n396_ );
nand g198 ( new_n400_, N130, N137 );
xnor g199 ( new_n401_, new_n400_, keyIn_0_17 );
not g200 ( new_n402_, new_n401_ );
nand g201 ( new_n403_, new_n399_, new_n402_ );
xnor g202 ( new_n404_, new_n395_, keyIn_0_61 );
nand g203 ( new_n405_, new_n404_, new_n401_ );
nand g204 ( new_n406_, new_n405_, new_n403_ );
nand g205 ( new_n407_, new_n406_, keyIn_0_65 );
not g206 ( new_n408_, keyIn_0_65 );
xnor g207 ( new_n409_, new_n399_, new_n401_ );
nand g208 ( new_n410_, new_n409_, new_n408_ );
nand g209 ( new_n411_, new_n410_, new_n407_ );
xor g210 ( new_n412_, N5, N21 );
xnor g211 ( new_n413_, new_n412_, keyIn_0_26 );
xnor g212 ( new_n414_, N37, N53 );
xnor g213 ( new_n415_, new_n414_, keyIn_0_27 );
xnor g214 ( new_n416_, new_n413_, new_n415_ );
xor g215 ( new_n417_, new_n416_, keyIn_0_49 );
nand g216 ( new_n418_, new_n411_, new_n417_ );
xnor g217 ( new_n419_, new_n406_, new_n408_ );
not g218 ( new_n420_, new_n417_ );
nand g219 ( new_n421_, new_n419_, new_n420_ );
nand g220 ( new_n422_, new_n421_, new_n418_ );
nand g221 ( new_n423_, new_n422_, keyIn_0_73 );
not g222 ( new_n424_, keyIn_0_73 );
xnor g223 ( new_n425_, new_n411_, new_n420_ );
nand g224 ( new_n426_, new_n425_, new_n424_ );
nand g225 ( new_n427_, new_n426_, new_n423_ );
nand g226 ( new_n428_, new_n391_, new_n427_ );
xnor g227 ( new_n429_, new_n328_, new_n275_ );
nand g228 ( new_n430_, new_n429_, keyIn_0_87 );
not g229 ( new_n431_, keyIn_0_88 );
xnor g230 ( new_n432_, new_n385_, new_n387_ );
nand g231 ( new_n433_, new_n432_, new_n431_ );
nand g232 ( new_n434_, new_n430_, new_n433_ );
nor g233 ( new_n435_, new_n434_, new_n428_ );
nand g234 ( new_n436_, new_n334_, new_n435_ );
xnor g235 ( new_n437_, new_n436_, new_n272_ );
not g236 ( new_n438_, keyIn_0_105 );
xnor g237 ( new_n439_, new_n422_, new_n424_ );
nor g238 ( new_n440_, new_n439_, keyIn_0_84 );
not g239 ( new_n441_, new_n440_ );
not g240 ( new_n442_, keyIn_0_84 );
nor g241 ( new_n443_, new_n427_, new_n442_ );
nor g242 ( new_n444_, new_n443_, new_n429_ );
nand g243 ( new_n445_, new_n444_, new_n441_ );
not g244 ( new_n446_, keyIn_0_85 );
nand g245 ( new_n447_, new_n432_, new_n446_ );
nand g246 ( new_n448_, new_n390_, keyIn_0_85 );
nand g247 ( new_n449_, new_n447_, new_n448_ );
nand g248 ( new_n450_, new_n271_, keyIn_0_83 );
not g249 ( new_n451_, keyIn_0_83 );
xnor g250 ( new_n452_, new_n259_, new_n265_ );
nand g251 ( new_n453_, new_n452_, keyIn_0_72 );
not g252 ( new_n454_, keyIn_0_72 );
nand g253 ( new_n455_, new_n270_, new_n454_ );
nand g254 ( new_n456_, new_n453_, new_n455_ );
nand g255 ( new_n457_, new_n456_, new_n451_ );
nand g256 ( new_n458_, new_n450_, new_n457_ );
nand g257 ( new_n459_, new_n458_, new_n449_ );
nor g258 ( new_n460_, new_n445_, new_n459_ );
xnor g259 ( new_n461_, new_n460_, new_n438_ );
nor g260 ( new_n462_, new_n461_, new_n437_ );
not g261 ( new_n463_, keyIn_0_107 );
not g262 ( new_n464_, keyIn_0_91 );
nor g263 ( new_n465_, new_n390_, new_n464_ );
not g264 ( new_n466_, keyIn_0_90 );
nand g265 ( new_n467_, new_n330_, new_n466_ );
not g266 ( new_n468_, keyIn_0_89 );
nand g267 ( new_n469_, new_n439_, new_n468_ );
nand g268 ( new_n470_, new_n469_, new_n467_ );
nor g269 ( new_n471_, new_n470_, new_n465_ );
nand g270 ( new_n472_, new_n427_, keyIn_0_89 );
nand g271 ( new_n473_, new_n472_, new_n271_ );
nand g272 ( new_n474_, new_n390_, new_n464_ );
nand g273 ( new_n475_, new_n429_, keyIn_0_90 );
nand g274 ( new_n476_, new_n475_, new_n474_ );
nor g275 ( new_n477_, new_n476_, new_n473_ );
nand g276 ( new_n478_, new_n477_, new_n471_ );
xnor g277 ( new_n479_, new_n478_, new_n463_ );
not g278 ( new_n480_, keyIn_0_104 );
nor g279 ( new_n481_, new_n429_, keyIn_0_82 );
not g280 ( new_n482_, new_n481_ );
not g281 ( new_n483_, keyIn_0_82 );
nor g282 ( new_n484_, new_n330_, new_n483_ );
nor g283 ( new_n485_, new_n484_, new_n390_ );
nand g284 ( new_n486_, new_n485_, new_n482_ );
not g285 ( new_n487_, keyIn_0_80 );
nand g286 ( new_n488_, new_n271_, new_n487_ );
nand g287 ( new_n489_, new_n456_, keyIn_0_80 );
nand g288 ( new_n490_, new_n488_, new_n489_ );
nand g289 ( new_n491_, new_n439_, keyIn_0_81 );
not g290 ( new_n492_, keyIn_0_81 );
nand g291 ( new_n493_, new_n427_, new_n492_ );
nand g292 ( new_n494_, new_n491_, new_n493_ );
nand g293 ( new_n495_, new_n494_, new_n490_ );
nor g294 ( new_n496_, new_n486_, new_n495_ );
xnor g295 ( new_n497_, new_n496_, new_n480_ );
nor g296 ( new_n498_, new_n497_, new_n479_ );
nand g297 ( new_n499_, new_n462_, new_n498_ );
nand g298 ( new_n500_, new_n499_, keyIn_0_112 );
not g299 ( new_n501_, keyIn_0_112 );
xnor g300 ( new_n502_, new_n436_, keyIn_0_106 );
nand g301 ( new_n503_, new_n460_, keyIn_0_105 );
nand g302 ( new_n504_, new_n439_, keyIn_0_84 );
nand g303 ( new_n505_, new_n504_, new_n330_ );
nor g304 ( new_n506_, new_n505_, new_n440_ );
not g305 ( new_n507_, new_n459_ );
nand g306 ( new_n508_, new_n507_, new_n506_ );
nand g307 ( new_n509_, new_n508_, new_n438_ );
nand g308 ( new_n510_, new_n509_, new_n503_ );
nand g309 ( new_n511_, new_n502_, new_n510_ );
xnor g310 ( new_n512_, new_n478_, keyIn_0_107 );
nand g311 ( new_n513_, new_n496_, keyIn_0_104 );
nand g312 ( new_n514_, new_n429_, keyIn_0_82 );
nand g313 ( new_n515_, new_n514_, new_n432_ );
nor g314 ( new_n516_, new_n515_, new_n481_ );
not g315 ( new_n517_, new_n495_ );
nand g316 ( new_n518_, new_n517_, new_n516_ );
nand g317 ( new_n519_, new_n518_, new_n480_ );
nand g318 ( new_n520_, new_n519_, new_n513_ );
nand g319 ( new_n521_, new_n512_, new_n520_ );
nor g320 ( new_n522_, new_n521_, new_n511_ );
nand g321 ( new_n523_, new_n522_, new_n501_ );
nand g322 ( new_n524_, new_n500_, new_n523_ );
not g323 ( new_n525_, new_n524_ );
not g324 ( new_n526_, keyIn_0_78 );
not g325 ( new_n527_, keyIn_0_4 );
xnor g326 ( new_n528_, N33, N37 );
xnor g327 ( new_n529_, new_n528_, new_n527_ );
not g328 ( new_n530_, keyIn_0_5 );
xnor g329 ( new_n531_, N41, N45 );
xnor g330 ( new_n532_, new_n531_, new_n530_ );
nand g331 ( new_n533_, new_n529_, new_n532_ );
xnor g332 ( new_n534_, new_n528_, keyIn_0_4 );
xnor g333 ( new_n535_, new_n531_, keyIn_0_5 );
nand g334 ( new_n536_, new_n534_, new_n535_ );
nand g335 ( new_n537_, new_n533_, new_n536_ );
xnor g336 ( new_n538_, new_n537_, keyIn_0_42 );
not g337 ( new_n539_, keyIn_0_40 );
not g338 ( new_n540_, keyIn_0_1 );
xnor g339 ( new_n541_, N9, N13 );
xnor g340 ( new_n542_, new_n541_, new_n540_ );
not g341 ( new_n543_, keyIn_0_0 );
xnor g342 ( new_n544_, N1, N5 );
nand g343 ( new_n545_, new_n544_, new_n543_ );
nor g344 ( new_n546_, N1, N5 );
nand g345 ( new_n547_, N1, N5 );
not g346 ( new_n548_, new_n547_ );
nor g347 ( new_n549_, new_n548_, new_n546_ );
nand g348 ( new_n550_, new_n549_, keyIn_0_0 );
nand g349 ( new_n551_, new_n550_, new_n545_ );
xnor g350 ( new_n552_, new_n542_, new_n551_ );
nand g351 ( new_n553_, new_n552_, new_n539_ );
xnor g352 ( new_n554_, new_n541_, keyIn_0_1 );
nand g353 ( new_n555_, new_n554_, new_n551_ );
xnor g354 ( new_n556_, new_n544_, keyIn_0_0 );
nand g355 ( new_n557_, new_n542_, new_n556_ );
nand g356 ( new_n558_, new_n557_, new_n555_ );
nand g357 ( new_n559_, new_n558_, keyIn_0_40 );
nand g358 ( new_n560_, new_n553_, new_n559_ );
xnor g359 ( new_n561_, new_n538_, new_n560_ );
nand g360 ( new_n562_, new_n561_, keyIn_0_58 );
not g361 ( new_n563_, keyIn_0_58 );
xnor g362 ( new_n564_, new_n558_, new_n539_ );
nand g363 ( new_n565_, new_n538_, new_n564_ );
not g364 ( new_n566_, keyIn_0_42 );
xnor g365 ( new_n567_, new_n537_, new_n566_ );
nand g366 ( new_n568_, new_n567_, new_n560_ );
nand g367 ( new_n569_, new_n565_, new_n568_ );
nand g368 ( new_n570_, new_n569_, new_n563_ );
nand g369 ( new_n571_, new_n562_, new_n570_ );
nand g370 ( new_n572_, N135, N137 );
xnor g371 ( new_n573_, new_n572_, keyIn_0_22 );
not g372 ( new_n574_, new_n573_ );
nand g373 ( new_n575_, new_n571_, new_n574_ );
xnor g374 ( new_n576_, new_n569_, keyIn_0_58 );
nand g375 ( new_n577_, new_n576_, new_n573_ );
nand g376 ( new_n578_, new_n577_, new_n575_ );
nand g377 ( new_n579_, new_n578_, keyIn_0_70 );
not g378 ( new_n580_, keyIn_0_70 );
xnor g379 ( new_n581_, new_n571_, new_n573_ );
nand g380 ( new_n582_, new_n581_, new_n580_ );
nand g381 ( new_n583_, new_n582_, new_n579_ );
xor g382 ( new_n584_, N73, N89 );
xnor g383 ( new_n585_, new_n584_, keyIn_0_36 );
xor g384 ( new_n586_, N105, N121 );
xnor g385 ( new_n587_, new_n586_, keyIn_0_37 );
xnor g386 ( new_n588_, new_n585_, new_n587_ );
xnor g387 ( new_n589_, new_n588_, keyIn_0_54 );
not g388 ( new_n590_, new_n589_ );
nand g389 ( new_n591_, new_n583_, new_n590_ );
xnor g390 ( new_n592_, new_n578_, new_n580_ );
nand g391 ( new_n593_, new_n592_, new_n589_ );
nand g392 ( new_n594_, new_n593_, new_n591_ );
xnor g393 ( new_n595_, new_n594_, new_n526_ );
not g394 ( new_n596_, keyIn_0_79 );
not g395 ( new_n597_, keyIn_0_41 );
xnor g396 ( new_n598_, N17, N21 );
xnor g397 ( new_n599_, new_n598_, keyIn_0_2 );
not g398 ( new_n600_, keyIn_0_3 );
xnor g399 ( new_n601_, N25, N29 );
nand g400 ( new_n602_, new_n601_, new_n600_ );
nor g401 ( new_n603_, N25, N29 );
nand g402 ( new_n604_, N25, N29 );
not g403 ( new_n605_, new_n604_ );
nor g404 ( new_n606_, new_n605_, new_n603_ );
nand g405 ( new_n607_, new_n606_, keyIn_0_3 );
nand g406 ( new_n608_, new_n607_, new_n602_ );
nand g407 ( new_n609_, new_n599_, new_n608_ );
not g408 ( new_n610_, keyIn_0_2 );
xnor g409 ( new_n611_, new_n598_, new_n610_ );
xnor g410 ( new_n612_, new_n601_, keyIn_0_3 );
nand g411 ( new_n613_, new_n611_, new_n612_ );
nand g412 ( new_n614_, new_n613_, new_n609_ );
nand g413 ( new_n615_, new_n614_, new_n597_ );
xnor g414 ( new_n616_, new_n611_, new_n608_ );
nand g415 ( new_n617_, new_n616_, keyIn_0_41 );
nand g416 ( new_n618_, new_n617_, new_n615_ );
not g417 ( new_n619_, keyIn_0_6 );
xnor g418 ( new_n620_, N49, N53 );
xnor g419 ( new_n621_, new_n620_, new_n619_ );
not g420 ( new_n622_, keyIn_0_7 );
xnor g421 ( new_n623_, N57, N61 );
nand g422 ( new_n624_, new_n623_, new_n622_ );
nor g423 ( new_n625_, N57, N61 );
nand g424 ( new_n626_, N57, N61 );
not g425 ( new_n627_, new_n626_ );
nor g426 ( new_n628_, new_n627_, new_n625_ );
nand g427 ( new_n629_, new_n628_, keyIn_0_7 );
nand g428 ( new_n630_, new_n629_, new_n624_ );
nand g429 ( new_n631_, new_n621_, new_n630_ );
xnor g430 ( new_n632_, new_n620_, keyIn_0_6 );
xnor g431 ( new_n633_, new_n623_, keyIn_0_7 );
nand g432 ( new_n634_, new_n632_, new_n633_ );
nand g433 ( new_n635_, new_n634_, new_n631_ );
nand g434 ( new_n636_, new_n635_, keyIn_0_43 );
not g435 ( new_n637_, keyIn_0_43 );
xnor g436 ( new_n638_, new_n632_, new_n630_ );
nand g437 ( new_n639_, new_n638_, new_n637_ );
nand g438 ( new_n640_, new_n639_, new_n636_ );
nand g439 ( new_n641_, new_n618_, new_n640_ );
xnor g440 ( new_n642_, new_n614_, keyIn_0_41 );
xnor g441 ( new_n643_, new_n635_, new_n637_ );
nand g442 ( new_n644_, new_n642_, new_n643_ );
nand g443 ( new_n645_, new_n644_, new_n641_ );
nand g444 ( new_n646_, new_n645_, keyIn_0_59 );
not g445 ( new_n647_, keyIn_0_59 );
xnor g446 ( new_n648_, new_n642_, new_n640_ );
nand g447 ( new_n649_, new_n648_, new_n647_ );
nand g448 ( new_n650_, new_n649_, new_n646_ );
nand g449 ( new_n651_, N136, N137 );
xor g450 ( new_n652_, new_n651_, keyIn_0_23 );
not g451 ( new_n653_, new_n652_ );
nand g452 ( new_n654_, new_n650_, new_n653_ );
xnor g453 ( new_n655_, new_n645_, new_n647_ );
nand g454 ( new_n656_, new_n655_, new_n652_ );
nand g455 ( new_n657_, new_n656_, new_n654_ );
nand g456 ( new_n658_, new_n657_, keyIn_0_71 );
not g457 ( new_n659_, keyIn_0_71 );
xnor g458 ( new_n660_, new_n650_, new_n652_ );
nand g459 ( new_n661_, new_n660_, new_n659_ );
nand g460 ( new_n662_, new_n661_, new_n658_ );
xor g461 ( new_n663_, N77, N93 );
xnor g462 ( new_n664_, new_n663_, keyIn_0_38 );
xnor g463 ( new_n665_, N109, N125 );
xnor g464 ( new_n666_, new_n665_, keyIn_0_39 );
xnor g465 ( new_n667_, new_n664_, new_n666_ );
xor g466 ( new_n668_, new_n667_, keyIn_0_55 );
not g467 ( new_n669_, new_n668_ );
xnor g468 ( new_n670_, new_n662_, new_n669_ );
nand g469 ( new_n671_, new_n670_, new_n596_ );
nand g470 ( new_n672_, new_n662_, new_n668_ );
xnor g471 ( new_n673_, new_n657_, new_n659_ );
nand g472 ( new_n674_, new_n673_, new_n669_ );
nand g473 ( new_n675_, new_n674_, new_n672_ );
nand g474 ( new_n676_, new_n675_, keyIn_0_79 );
nand g475 ( new_n677_, new_n671_, new_n676_ );
nor g476 ( new_n678_, new_n595_, new_n677_ );
not g477 ( new_n679_, keyIn_0_77 );
xnor g478 ( new_n680_, new_n538_, new_n640_ );
nand g479 ( new_n681_, new_n680_, keyIn_0_57 );
not g480 ( new_n682_, keyIn_0_57 );
nand g481 ( new_n683_, new_n538_, new_n643_ );
nand g482 ( new_n684_, new_n567_, new_n640_ );
nand g483 ( new_n685_, new_n683_, new_n684_ );
nand g484 ( new_n686_, new_n685_, new_n682_ );
nand g485 ( new_n687_, new_n681_, new_n686_ );
nand g486 ( new_n688_, N134, N137 );
xor g487 ( new_n689_, new_n688_, keyIn_0_21 );
nand g488 ( new_n690_, new_n687_, new_n689_ );
xnor g489 ( new_n691_, new_n685_, keyIn_0_57 );
not g490 ( new_n692_, new_n689_ );
nand g491 ( new_n693_, new_n691_, new_n692_ );
nand g492 ( new_n694_, new_n693_, new_n690_ );
nand g493 ( new_n695_, new_n694_, keyIn_0_69 );
not g494 ( new_n696_, keyIn_0_69 );
xnor g495 ( new_n697_, new_n687_, new_n692_ );
nand g496 ( new_n698_, new_n697_, new_n696_ );
nand g497 ( new_n699_, new_n698_, new_n695_ );
xnor g498 ( new_n700_, N69, N85 );
xnor g499 ( new_n701_, new_n700_, keyIn_0_34 );
xnor g500 ( new_n702_, N101, N117 );
xnor g501 ( new_n703_, new_n702_, keyIn_0_35 );
xnor g502 ( new_n704_, new_n701_, new_n703_ );
xor g503 ( new_n705_, new_n704_, keyIn_0_53 );
not g504 ( new_n706_, new_n705_ );
nand g505 ( new_n707_, new_n699_, new_n706_ );
xnor g506 ( new_n708_, new_n694_, new_n696_ );
nand g507 ( new_n709_, new_n708_, new_n705_ );
nand g508 ( new_n710_, new_n709_, new_n707_ );
xnor g509 ( new_n711_, new_n710_, new_n679_ );
not g510 ( new_n712_, keyIn_0_76 );
nand g511 ( new_n713_, new_n564_, new_n618_ );
nand g512 ( new_n714_, new_n642_, new_n560_ );
nand g513 ( new_n715_, new_n713_, new_n714_ );
nand g514 ( new_n716_, new_n715_, keyIn_0_56 );
not g515 ( new_n717_, keyIn_0_56 );
xnor g516 ( new_n718_, new_n560_, new_n618_ );
nand g517 ( new_n719_, new_n718_, new_n717_ );
nand g518 ( new_n720_, new_n719_, new_n716_ );
nand g519 ( new_n721_, N133, N137 );
xnor g520 ( new_n722_, new_n721_, keyIn_0_20 );
nand g521 ( new_n723_, new_n720_, new_n722_ );
xnor g522 ( new_n724_, new_n715_, new_n717_ );
not g523 ( new_n725_, new_n722_ );
nand g524 ( new_n726_, new_n724_, new_n725_ );
nand g525 ( new_n727_, new_n726_, new_n723_ );
nand g526 ( new_n728_, new_n727_, keyIn_0_68 );
not g527 ( new_n729_, keyIn_0_68 );
xnor g528 ( new_n730_, new_n720_, new_n725_ );
nand g529 ( new_n731_, new_n730_, new_n729_ );
nand g530 ( new_n732_, new_n731_, new_n728_ );
xor g531 ( new_n733_, N65, N81 );
xnor g532 ( new_n734_, new_n733_, keyIn_0_32 );
xor g533 ( new_n735_, N97, N113 );
xnor g534 ( new_n736_, new_n735_, keyIn_0_33 );
xnor g535 ( new_n737_, new_n734_, new_n736_ );
xor g536 ( new_n738_, new_n737_, keyIn_0_52 );
not g537 ( new_n739_, new_n738_ );
xnor g538 ( new_n740_, new_n732_, new_n739_ );
nand g539 ( new_n741_, new_n740_, new_n712_ );
nand g540 ( new_n742_, new_n732_, new_n738_ );
xnor g541 ( new_n743_, new_n727_, new_n729_ );
nand g542 ( new_n744_, new_n743_, new_n739_ );
nand g543 ( new_n745_, new_n744_, new_n742_ );
nand g544 ( new_n746_, new_n745_, keyIn_0_76 );
nand g545 ( new_n747_, new_n741_, new_n746_ );
nor g546 ( new_n748_, new_n711_, new_n747_ );
nand g547 ( new_n749_, new_n678_, new_n748_ );
nor g548 ( new_n750_, new_n525_, new_n749_ );
xor g549 ( new_n751_, new_n750_, keyIn_0_114 );
nand g550 ( new_n752_, new_n751_, new_n271_ );
xnor g551 ( N724, new_n752_, N1 );
nand g552 ( new_n754_, new_n751_, new_n427_ );
xnor g553 ( N725, new_n754_, N5 );
nand g554 ( new_n756_, new_n751_, new_n330_ );
xnor g555 ( N726, new_n756_, N9 );
nand g556 ( new_n758_, new_n751_, new_n432_ );
xnor g557 ( N727, new_n758_, N13 );
nand g558 ( new_n760_, new_n594_, keyIn_0_78 );
xnor g559 ( new_n761_, new_n583_, new_n589_ );
nand g560 ( new_n762_, new_n761_, new_n526_ );
nand g561 ( new_n763_, new_n762_, new_n760_ );
xnor g562 ( new_n764_, new_n675_, new_n596_ );
nor g563 ( new_n765_, new_n764_, new_n763_ );
nand g564 ( new_n766_, new_n765_, new_n748_ );
nor g565 ( new_n767_, new_n525_, new_n766_ );
xnor g566 ( new_n768_, new_n767_, keyIn_0_115 );
nand g567 ( new_n769_, new_n768_, new_n271_ );
xnor g568 ( N728, new_n769_, N17 );
nand g569 ( new_n771_, new_n768_, new_n427_ );
xnor g570 ( N729, new_n771_, N21 );
nand g571 ( new_n773_, new_n768_, new_n330_ );
xnor g572 ( N730, new_n773_, N25 );
nand g573 ( new_n775_, new_n768_, new_n432_ );
xnor g574 ( N731, new_n775_, N29 );
nand g575 ( new_n777_, new_n710_, keyIn_0_77 );
xnor g576 ( new_n778_, new_n699_, new_n705_ );
nand g577 ( new_n779_, new_n778_, new_n679_ );
nand g578 ( new_n780_, new_n779_, new_n777_ );
xnor g579 ( new_n781_, new_n745_, new_n712_ );
nor g580 ( new_n782_, new_n781_, new_n780_ );
nand g581 ( new_n783_, new_n782_, new_n678_ );
nor g582 ( new_n784_, new_n525_, new_n783_ );
xnor g583 ( new_n785_, new_n784_, keyIn_0_116 );
nand g584 ( new_n786_, new_n785_, new_n271_ );
xnor g585 ( N732, new_n786_, N33 );
nand g586 ( new_n788_, new_n785_, new_n427_ );
xnor g587 ( N733, new_n788_, N37 );
nand g588 ( new_n790_, new_n785_, new_n330_ );
xnor g589 ( N734, new_n790_, N41 );
nand g590 ( new_n792_, new_n785_, new_n432_ );
xnor g591 ( N735, new_n792_, N45 );
not g592 ( new_n794_, keyIn_0_117 );
not g593 ( new_n795_, new_n765_ );
not g594 ( new_n796_, new_n782_ );
nor g595 ( new_n797_, new_n795_, new_n796_ );
nand g596 ( new_n798_, new_n524_, new_n797_ );
xnor g597 ( new_n799_, new_n798_, new_n794_ );
nand g598 ( new_n800_, new_n799_, new_n271_ );
xnor g599 ( N736, new_n800_, N49 );
nand g600 ( new_n802_, new_n799_, new_n427_ );
xnor g601 ( N737, new_n802_, N53 );
nand g602 ( new_n804_, new_n799_, new_n330_ );
xnor g603 ( N738, new_n804_, N57 );
not g604 ( new_n806_, N61 );
nand g605 ( new_n807_, new_n799_, new_n432_ );
nand g606 ( new_n808_, new_n807_, keyIn_0_122 );
not g607 ( new_n809_, keyIn_0_122 );
xnor g608 ( new_n810_, new_n798_, keyIn_0_117 );
nor g609 ( new_n811_, new_n810_, new_n390_ );
nand g610 ( new_n812_, new_n811_, new_n809_ );
nand g611 ( new_n813_, new_n812_, new_n808_ );
nand g612 ( new_n814_, new_n813_, new_n806_ );
xnor g613 ( new_n815_, new_n807_, new_n809_ );
nand g614 ( new_n816_, new_n815_, N61 );
nand g615 ( N739, new_n816_, new_n814_ );
not g616 ( new_n818_, N65 );
not g617 ( new_n819_, keyIn_0_123 );
not g618 ( new_n820_, keyIn_0_113 );
not g619 ( new_n821_, keyIn_0_111 );
not g620 ( new_n822_, keyIn_0_103 );
nor g621 ( new_n823_, new_n764_, new_n822_ );
not g622 ( new_n824_, new_n823_ );
xnor g623 ( new_n825_, new_n780_, keyIn_0_101 );
nand g624 ( new_n826_, new_n825_, new_n824_ );
nand g625 ( new_n827_, new_n763_, keyIn_0_102 );
not g626 ( new_n828_, keyIn_0_102 );
nand g627 ( new_n829_, new_n595_, new_n828_ );
nand g628 ( new_n830_, new_n829_, new_n827_ );
nor g629 ( new_n831_, new_n677_, keyIn_0_103 );
nor g630 ( new_n832_, new_n831_, new_n747_ );
nand g631 ( new_n833_, new_n832_, new_n830_ );
nor g632 ( new_n834_, new_n826_, new_n833_ );
nor g633 ( new_n835_, new_n834_, new_n821_ );
not g634 ( new_n836_, keyIn_0_109 );
not g635 ( new_n837_, keyIn_0_97 );
nor g636 ( new_n838_, new_n764_, new_n837_ );
nand g637 ( new_n839_, new_n764_, new_n837_ );
nand g638 ( new_n840_, new_n839_, new_n763_ );
nor g639 ( new_n841_, new_n840_, new_n838_ );
not g640 ( new_n842_, keyIn_0_95 );
nand g641 ( new_n843_, new_n781_, new_n842_ );
nand g642 ( new_n844_, new_n747_, keyIn_0_95 );
nand g643 ( new_n845_, new_n843_, new_n844_ );
not g644 ( new_n846_, keyIn_0_96 );
nand g645 ( new_n847_, new_n711_, new_n846_ );
nand g646 ( new_n848_, new_n780_, keyIn_0_96 );
nand g647 ( new_n849_, new_n847_, new_n848_ );
nand g648 ( new_n850_, new_n849_, new_n845_ );
not g649 ( new_n851_, new_n850_ );
nand g650 ( new_n852_, new_n851_, new_n841_ );
nor g651 ( new_n853_, new_n852_, new_n836_ );
nor g652 ( new_n854_, new_n853_, new_n835_ );
not g653 ( new_n855_, new_n838_ );
nor g654 ( new_n856_, new_n677_, keyIn_0_97 );
nor g655 ( new_n857_, new_n856_, new_n595_ );
nand g656 ( new_n858_, new_n857_, new_n855_ );
nor g657 ( new_n859_, new_n858_, new_n850_ );
nor g658 ( new_n860_, new_n859_, keyIn_0_109 );
nand g659 ( new_n861_, new_n711_, keyIn_0_101 );
not g660 ( new_n862_, keyIn_0_101 );
nand g661 ( new_n863_, new_n780_, new_n862_ );
nand g662 ( new_n864_, new_n861_, new_n863_ );
nor g663 ( new_n865_, new_n864_, new_n823_ );
xnor g664 ( new_n866_, new_n763_, new_n828_ );
nand g665 ( new_n867_, new_n764_, new_n822_ );
nand g666 ( new_n868_, new_n867_, new_n781_ );
nor g667 ( new_n869_, new_n866_, new_n868_ );
nand g668 ( new_n870_, new_n869_, new_n865_ );
nor g669 ( new_n871_, new_n870_, keyIn_0_111 );
nor g670 ( new_n872_, new_n871_, new_n860_ );
nand g671 ( new_n873_, new_n854_, new_n872_ );
not g672 ( new_n874_, keyIn_0_99 );
nor g673 ( new_n875_, new_n763_, new_n874_ );
not g674 ( new_n876_, keyIn_0_100 );
nand g675 ( new_n877_, new_n764_, new_n876_ );
nand g676 ( new_n878_, new_n763_, new_n874_ );
nand g677 ( new_n879_, new_n877_, new_n878_ );
nor g678 ( new_n880_, new_n879_, new_n875_ );
not g679 ( new_n881_, keyIn_0_98 );
xnor g680 ( new_n882_, new_n747_, new_n881_ );
nand g681 ( new_n883_, new_n677_, keyIn_0_100 );
nand g682 ( new_n884_, new_n883_, new_n711_ );
nor g683 ( new_n885_, new_n882_, new_n884_ );
nand g684 ( new_n886_, new_n885_, new_n880_ );
nand g685 ( new_n887_, new_n886_, keyIn_0_110 );
not g686 ( new_n888_, keyIn_0_110 );
not g687 ( new_n889_, new_n875_ );
nor g688 ( new_n890_, new_n677_, keyIn_0_100 );
nor g689 ( new_n891_, new_n595_, keyIn_0_99 );
nor g690 ( new_n892_, new_n891_, new_n890_ );
nand g691 ( new_n893_, new_n892_, new_n889_ );
xnor g692 ( new_n894_, new_n747_, keyIn_0_98 );
not g693 ( new_n895_, new_n884_ );
nand g694 ( new_n896_, new_n895_, new_n894_ );
nor g695 ( new_n897_, new_n896_, new_n893_ );
nand g696 ( new_n898_, new_n897_, new_n888_ );
nand g697 ( new_n899_, new_n898_, new_n887_ );
not g698 ( new_n900_, keyIn_0_93 );
nor g699 ( new_n901_, new_n711_, new_n900_ );
not g700 ( new_n902_, keyIn_0_92 );
nand g701 ( new_n903_, new_n781_, new_n902_ );
nand g702 ( new_n904_, new_n747_, keyIn_0_92 );
nand g703 ( new_n905_, new_n903_, new_n904_ );
nor g704 ( new_n906_, new_n905_, new_n901_ );
not g705 ( new_n907_, keyIn_0_94 );
nand g706 ( new_n908_, new_n595_, new_n907_ );
nand g707 ( new_n909_, new_n908_, new_n677_ );
nand g708 ( new_n910_, new_n711_, new_n900_ );
nand g709 ( new_n911_, new_n763_, keyIn_0_94 );
nand g710 ( new_n912_, new_n910_, new_n911_ );
nor g711 ( new_n913_, new_n909_, new_n912_ );
nand g712 ( new_n914_, new_n913_, new_n906_ );
xnor g713 ( new_n915_, new_n914_, keyIn_0_108 );
nand g714 ( new_n916_, new_n915_, new_n899_ );
nor g715 ( new_n917_, new_n873_, new_n916_ );
nand g716 ( new_n918_, new_n917_, new_n820_ );
nand g717 ( new_n919_, new_n870_, keyIn_0_111 );
nand g718 ( new_n920_, new_n859_, keyIn_0_109 );
nand g719 ( new_n921_, new_n919_, new_n920_ );
nand g720 ( new_n922_, new_n852_, new_n836_ );
nand g721 ( new_n923_, new_n834_, new_n821_ );
nand g722 ( new_n924_, new_n922_, new_n923_ );
nor g723 ( new_n925_, new_n924_, new_n921_ );
xnor g724 ( new_n926_, new_n886_, new_n888_ );
not g725 ( new_n927_, keyIn_0_108 );
xnor g726 ( new_n928_, new_n914_, new_n927_ );
nor g727 ( new_n929_, new_n926_, new_n928_ );
nand g728 ( new_n930_, new_n929_, new_n925_ );
nand g729 ( new_n931_, new_n930_, keyIn_0_113 );
nand g730 ( new_n932_, new_n918_, new_n931_ );
nor g731 ( new_n933_, new_n429_, new_n432_ );
not g732 ( new_n934_, new_n933_ );
nand g733 ( new_n935_, new_n439_, new_n271_ );
nor g734 ( new_n936_, new_n934_, new_n935_ );
nand g735 ( new_n937_, new_n932_, new_n936_ );
xnor g736 ( new_n938_, new_n937_, keyIn_0_118 );
nand g737 ( new_n939_, new_n938_, new_n781_ );
nand g738 ( new_n940_, new_n939_, new_n819_ );
not g739 ( new_n941_, keyIn_0_118 );
xnor g740 ( new_n942_, new_n937_, new_n941_ );
nor g741 ( new_n943_, new_n942_, new_n747_ );
nand g742 ( new_n944_, new_n943_, keyIn_0_123 );
nand g743 ( new_n945_, new_n944_, new_n940_ );
nand g744 ( new_n946_, new_n945_, new_n818_ );
xnor g745 ( new_n947_, new_n939_, keyIn_0_123 );
nand g746 ( new_n948_, new_n947_, N65 );
nand g747 ( N740, new_n948_, new_n946_ );
not g748 ( new_n950_, N69 );
not g749 ( new_n951_, keyIn_0_124 );
nand g750 ( new_n952_, new_n938_, new_n711_ );
nand g751 ( new_n953_, new_n952_, new_n951_ );
nor g752 ( new_n954_, new_n942_, new_n780_ );
nand g753 ( new_n955_, new_n954_, keyIn_0_124 );
nand g754 ( new_n956_, new_n955_, new_n953_ );
nand g755 ( new_n957_, new_n956_, new_n950_ );
xnor g756 ( new_n958_, new_n952_, keyIn_0_124 );
nand g757 ( new_n959_, new_n958_, N69 );
nand g758 ( N741, new_n959_, new_n957_ );
not g759 ( new_n961_, N73 );
nand g760 ( new_n962_, new_n938_, new_n763_ );
nand g761 ( new_n963_, new_n962_, keyIn_0_125 );
not g762 ( new_n964_, keyIn_0_125 );
nor g763 ( new_n965_, new_n942_, new_n595_ );
nand g764 ( new_n966_, new_n965_, new_n964_ );
nand g765 ( new_n967_, new_n966_, new_n963_ );
nand g766 ( new_n968_, new_n967_, new_n961_ );
xnor g767 ( new_n969_, new_n962_, new_n964_ );
nand g768 ( new_n970_, new_n969_, N73 );
nand g769 ( N742, new_n970_, new_n968_ );
not g770 ( new_n972_, N77 );
not g771 ( new_n973_, keyIn_0_126 );
nand g772 ( new_n974_, new_n938_, new_n677_ );
nand g773 ( new_n975_, new_n974_, new_n973_ );
nor g774 ( new_n976_, new_n942_, new_n764_ );
nand g775 ( new_n977_, new_n976_, keyIn_0_126 );
nand g776 ( new_n978_, new_n977_, new_n975_ );
nand g777 ( new_n979_, new_n978_, new_n972_ );
xnor g778 ( new_n980_, new_n974_, keyIn_0_126 );
nand g779 ( new_n981_, new_n980_, N77 );
nand g780 ( N743, new_n981_, new_n979_ );
not g781 ( new_n983_, N81 );
not g782 ( new_n984_, keyIn_0_127 );
nor g783 ( new_n985_, new_n330_, new_n390_ );
not g784 ( new_n986_, new_n985_ );
nor g785 ( new_n987_, new_n986_, new_n935_ );
nand g786 ( new_n988_, new_n932_, new_n987_ );
xnor g787 ( new_n989_, new_n988_, keyIn_0_119 );
nand g788 ( new_n990_, new_n989_, new_n781_ );
nand g789 ( new_n991_, new_n990_, new_n984_ );
not g790 ( new_n992_, keyIn_0_119 );
xnor g791 ( new_n993_, new_n988_, new_n992_ );
nor g792 ( new_n994_, new_n993_, new_n747_ );
nand g793 ( new_n995_, new_n994_, keyIn_0_127 );
nand g794 ( new_n996_, new_n995_, new_n991_ );
nand g795 ( new_n997_, new_n996_, new_n983_ );
xnor g796 ( new_n998_, new_n990_, keyIn_0_127 );
nand g797 ( new_n999_, new_n998_, N81 );
nand g798 ( N744, new_n999_, new_n997_ );
nand g799 ( new_n1001_, new_n989_, new_n711_ );
xnor g800 ( N745, new_n1001_, N85 );
nand g801 ( new_n1003_, new_n989_, new_n763_ );
xnor g802 ( N746, new_n1003_, N89 );
nand g803 ( new_n1005_, new_n989_, new_n677_ );
xnor g804 ( N747, new_n1005_, N93 );
not g805 ( new_n1007_, new_n932_ );
nor g806 ( new_n1008_, new_n439_, new_n271_ );
nand g807 ( new_n1009_, new_n1008_, new_n933_ );
nor g808 ( new_n1010_, new_n1007_, new_n1009_ );
xnor g809 ( new_n1011_, new_n1010_, keyIn_0_120 );
nand g810 ( new_n1012_, new_n1011_, new_n781_ );
xnor g811 ( N748, new_n1012_, N97 );
nand g812 ( new_n1014_, new_n1011_, new_n711_ );
xnor g813 ( N749, new_n1014_, N101 );
nand g814 ( new_n1016_, new_n1011_, new_n763_ );
xnor g815 ( N750, new_n1016_, N105 );
nand g816 ( new_n1018_, new_n1011_, new_n677_ );
xnor g817 ( N751, new_n1018_, N109 );
nand g818 ( new_n1020_, new_n1008_, new_n985_ );
nor g819 ( new_n1021_, new_n1007_, new_n1020_ );
xor g820 ( new_n1022_, new_n1021_, keyIn_0_121 );
nand g821 ( new_n1023_, new_n1022_, new_n781_ );
xnor g822 ( N752, new_n1023_, N113 );
nand g823 ( new_n1025_, new_n1022_, new_n711_ );
xnor g824 ( N753, new_n1025_, N117 );
nand g825 ( new_n1027_, new_n1022_, new_n763_ );
xnor g826 ( N754, new_n1027_, N121 );
nand g827 ( new_n1029_, new_n1022_, new_n677_ );
xnor g828 ( N755, new_n1029_, N125 );
endmodule