module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n114_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n317_, new_n287_, new_n234_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n449_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n248_, new_n350_, new_n117_, new_n167_, new_n385_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n158_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n194_, new_n116_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n399_, new_n233_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n460_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n107_, new_n182_, new_n407_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n444_, new_n392_, new_n147_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n404_, new_n193_, new_n128_, new_n348_, new_n159_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n200_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n229_, new_n204_, new_n181_, new_n135_, new_n405_;

xor g000 ( new_n106_, N89, N93 );
xnor g001 ( new_n107_, N81, N85 );
xnor g002 ( new_n108_, new_n106_, new_n107_ );
xor g003 ( new_n109_, N65, N69 );
xnor g004 ( new_n110_, N73, N77 );
xnor g005 ( new_n111_, new_n109_, new_n110_ );
xor g006 ( new_n112_, new_n108_, new_n111_ );
nand g007 ( new_n113_, N129, N137 );
xnor g008 ( new_n114_, new_n112_, new_n113_ );
xor g009 ( new_n115_, N33, N49 );
xnor g010 ( new_n116_, N1, N17 );
xnor g011 ( new_n117_, new_n115_, new_n116_ );
xnor g012 ( new_n118_, new_n117_, keyIn_0_9 );
xnor g013 ( new_n119_, new_n114_, new_n118_ );
not g014 ( new_n120_, new_n119_ );
xnor g015 ( new_n121_, N113, N117 );
xnor g016 ( new_n122_, new_n121_, keyIn_0_4 );
xnor g017 ( new_n123_, N121, N125 );
xnor g018 ( new_n124_, new_n122_, new_n123_ );
xnor g019 ( new_n125_, N105, N109 );
xnor g020 ( new_n126_, new_n125_, keyIn_0_3 );
xor g021 ( new_n127_, N97, N101 );
xnor g022 ( new_n128_, new_n126_, new_n127_ );
xor g023 ( new_n129_, new_n124_, new_n128_ );
nand g024 ( new_n130_, N130, N137 );
xnor g025 ( new_n131_, new_n129_, new_n130_ );
xor g026 ( new_n132_, N37, N53 );
xnor g027 ( new_n133_, N5, N21 );
xnor g028 ( new_n134_, new_n132_, new_n133_ );
xor g029 ( new_n135_, new_n131_, new_n134_ );
not g030 ( new_n136_, new_n135_ );
xnor g031 ( new_n137_, new_n128_, new_n111_ );
nand g032 ( new_n138_, N131, N137 );
xor g033 ( new_n139_, new_n137_, new_n138_ );
xnor g034 ( new_n140_, N41, N57 );
xnor g035 ( new_n141_, new_n140_, keyIn_0_6 );
xor g036 ( new_n142_, N9, N25 );
xnor g037 ( new_n143_, new_n141_, new_n142_ );
xor g038 ( new_n144_, new_n139_, new_n143_ );
nand g039 ( new_n145_, new_n144_, keyIn_0_12 );
nor g040 ( new_n146_, new_n145_, new_n136_ );
nand g041 ( new_n147_, new_n145_, new_n136_ );
xnor g042 ( new_n148_, new_n124_, new_n108_ );
nand g043 ( new_n149_, N132, N137 );
xor g044 ( new_n150_, new_n148_, new_n149_ );
xor g045 ( new_n151_, N45, N61 );
xnor g046 ( new_n152_, N13, N29 );
xnor g047 ( new_n153_, new_n151_, new_n152_ );
xnor g048 ( new_n154_, new_n150_, new_n153_ );
not g049 ( new_n155_, new_n154_ );
nor g050 ( new_n156_, new_n155_, new_n120_ );
nand g051 ( new_n157_, new_n147_, new_n156_ );
nor g052 ( new_n158_, new_n157_, new_n146_ );
not g053 ( new_n159_, new_n158_ );
nor g054 ( new_n160_, new_n144_, new_n154_ );
xor g055 ( new_n161_, new_n119_, keyIn_0_11 );
nor g056 ( new_n162_, new_n161_, new_n135_ );
nand g057 ( new_n163_, new_n162_, new_n160_ );
xor g058 ( new_n164_, new_n163_, keyIn_0_19 );
xor g059 ( new_n165_, new_n135_, keyIn_0_13 );
nor g060 ( new_n166_, new_n144_, new_n119_ );
nand g061 ( new_n167_, new_n166_, new_n154_ );
nor g062 ( new_n168_, new_n165_, new_n167_ );
nor g063 ( new_n169_, new_n164_, new_n168_ );
nand g064 ( new_n170_, new_n169_, new_n159_ );
xnor g065 ( new_n171_, N57, N61 );
xnor g066 ( new_n172_, N49, N53 );
xnor g067 ( new_n173_, new_n171_, new_n172_ );
not g068 ( new_n174_, new_n173_ );
not g069 ( new_n175_, keyIn_0_8 );
not g070 ( new_n176_, N45 );
nand g071 ( new_n177_, new_n176_, N41 );
not g072 ( new_n178_, N41 );
nand g073 ( new_n179_, new_n178_, N45 );
nand g074 ( new_n180_, new_n177_, new_n179_ );
nand g075 ( new_n181_, new_n180_, keyIn_0_2 );
not g076 ( new_n182_, keyIn_0_2 );
xnor g077 ( new_n183_, N41, N45 );
nand g078 ( new_n184_, new_n183_, new_n182_ );
nand g079 ( new_n185_, new_n181_, new_n184_ );
not g080 ( new_n186_, keyIn_0_1 );
xnor g081 ( new_n187_, N33, N37 );
nand g082 ( new_n188_, new_n187_, new_n186_ );
not g083 ( new_n189_, N37 );
nand g084 ( new_n190_, new_n189_, N33 );
not g085 ( new_n191_, N33 );
nand g086 ( new_n192_, new_n191_, N37 );
nand g087 ( new_n193_, new_n190_, new_n192_ );
nand g088 ( new_n194_, new_n193_, keyIn_0_1 );
and g089 ( new_n195_, new_n194_, new_n188_ );
nand g090 ( new_n196_, new_n195_, new_n185_ );
xnor g091 ( new_n197_, new_n183_, keyIn_0_2 );
nand g092 ( new_n198_, new_n194_, new_n188_ );
nand g093 ( new_n199_, new_n197_, new_n198_ );
nand g094 ( new_n200_, new_n196_, new_n199_ );
nand g095 ( new_n201_, new_n200_, new_n175_ );
xnor g096 ( new_n202_, new_n185_, new_n198_ );
nand g097 ( new_n203_, new_n202_, keyIn_0_8 );
nand g098 ( new_n204_, new_n203_, new_n201_ );
nand g099 ( new_n205_, new_n204_, new_n174_ );
xnor g100 ( new_n206_, new_n200_, keyIn_0_8 );
nand g101 ( new_n207_, new_n206_, new_n173_ );
nand g102 ( new_n208_, new_n207_, new_n205_ );
nand g103 ( new_n209_, N134, N137 );
nand g104 ( new_n210_, new_n208_, new_n209_ );
xnor g105 ( new_n211_, new_n204_, new_n173_ );
not g106 ( new_n212_, new_n209_ );
nand g107 ( new_n213_, new_n211_, new_n212_ );
nand g108 ( new_n214_, new_n213_, new_n210_ );
xnor g109 ( new_n215_, N101, N117 );
xnor g110 ( new_n216_, N69, N85 );
xnor g111 ( new_n217_, new_n215_, new_n216_ );
xnor g112 ( new_n218_, new_n214_, new_n217_ );
nand g113 ( new_n219_, new_n218_, keyIn_0_14 );
nor g114 ( new_n220_, new_n218_, keyIn_0_14 );
xnor g115 ( new_n221_, N17, N21 );
xnor g116 ( new_n222_, new_n221_, keyIn_0_0 );
xnor g117 ( new_n223_, N25, N29 );
not g118 ( new_n224_, new_n223_ );
nand g119 ( new_n225_, new_n222_, new_n224_ );
not g120 ( new_n226_, N21 );
nand g121 ( new_n227_, new_n226_, N17 );
not g122 ( new_n228_, N17 );
nand g123 ( new_n229_, new_n228_, N21 );
nand g124 ( new_n230_, new_n227_, new_n229_ );
nand g125 ( new_n231_, new_n230_, keyIn_0_0 );
not g126 ( new_n232_, keyIn_0_0 );
nand g127 ( new_n233_, new_n221_, new_n232_ );
nand g128 ( new_n234_, new_n231_, new_n233_ );
nand g129 ( new_n235_, new_n234_, new_n223_ );
nand g130 ( new_n236_, new_n225_, new_n235_ );
xor g131 ( new_n237_, N9, N13 );
xnor g132 ( new_n238_, N1, N5 );
xnor g133 ( new_n239_, new_n237_, new_n238_ );
not g134 ( new_n240_, new_n239_ );
xnor g135 ( new_n241_, new_n236_, new_n240_ );
nand g136 ( new_n242_, N133, N137 );
xnor g137 ( new_n243_, new_n241_, new_n242_ );
xor g138 ( new_n244_, N97, N113 );
xnor g139 ( new_n245_, N65, N81 );
xnor g140 ( new_n246_, new_n244_, new_n245_ );
xnor g141 ( new_n247_, new_n243_, new_n246_ );
nor g142 ( new_n248_, new_n220_, new_n247_ );
nand g143 ( new_n249_, new_n248_, new_n219_ );
xnor g144 ( new_n250_, new_n234_, new_n224_ );
nand g145 ( new_n251_, new_n250_, new_n174_ );
nand g146 ( new_n252_, new_n236_, new_n173_ );
nand g147 ( new_n253_, new_n251_, new_n252_ );
nand g148 ( new_n254_, N136, N137 );
not g149 ( new_n255_, new_n254_ );
xnor g150 ( new_n256_, new_n253_, new_n255_ );
nand g151 ( new_n257_, new_n256_, keyIn_0_10 );
not g152 ( new_n258_, keyIn_0_10 );
xnor g153 ( new_n259_, new_n236_, new_n174_ );
nand g154 ( new_n260_, new_n259_, new_n255_ );
nand g155 ( new_n261_, new_n253_, new_n254_ );
nand g156 ( new_n262_, new_n260_, new_n261_ );
nand g157 ( new_n263_, new_n262_, new_n258_ );
nand g158 ( new_n264_, new_n257_, new_n263_ );
xnor g159 ( new_n265_, N109, N125 );
xnor g160 ( new_n266_, N77, N93 );
xnor g161 ( new_n267_, new_n265_, new_n266_ );
not g162 ( new_n268_, new_n267_ );
xnor g163 ( new_n269_, new_n264_, new_n268_ );
xnor g164 ( new_n270_, new_n269_, keyIn_0_15 );
nand g165 ( new_n271_, new_n204_, new_n239_ );
nand g166 ( new_n272_, new_n206_, new_n240_ );
nand g167 ( new_n273_, new_n272_, new_n271_ );
nand g168 ( new_n274_, new_n273_, keyIn_0_5 );
not g169 ( new_n275_, keyIn_0_5 );
xnor g170 ( new_n276_, new_n204_, new_n240_ );
nand g171 ( new_n277_, new_n276_, new_n275_ );
nand g172 ( new_n278_, new_n277_, new_n274_ );
nand g173 ( new_n279_, N135, N137 );
not g174 ( new_n280_, new_n279_ );
xnor g175 ( new_n281_, new_n278_, new_n280_ );
xnor g176 ( new_n282_, N105, N121 );
xnor g177 ( new_n283_, new_n282_, keyIn_0_7 );
xnor g178 ( new_n284_, N73, N89 );
xnor g179 ( new_n285_, new_n283_, new_n284_ );
nand g180 ( new_n286_, new_n281_, new_n285_ );
nand g181 ( new_n287_, new_n278_, new_n279_ );
xnor g182 ( new_n288_, new_n273_, new_n275_ );
nand g183 ( new_n289_, new_n288_, new_n280_ );
nand g184 ( new_n290_, new_n289_, new_n287_ );
not g185 ( new_n291_, new_n285_ );
nand g186 ( new_n292_, new_n290_, new_n291_ );
nand g187 ( new_n293_, new_n286_, new_n292_ );
nand g188 ( new_n294_, new_n270_, new_n293_ );
nor g189 ( new_n295_, new_n249_, new_n294_ );
nand g190 ( new_n296_, new_n170_, new_n295_ );
xnor g191 ( new_n297_, new_n296_, keyIn_0_24 );
nand g192 ( new_n298_, new_n297_, new_n120_ );
xnor g193 ( N724, new_n298_, N1 );
nand g194 ( new_n300_, new_n297_, new_n135_ );
xnor g195 ( N725, new_n300_, N5 );
nand g196 ( new_n302_, new_n297_, new_n144_ );
xnor g197 ( new_n303_, new_n302_, N9 );
xnor g198 ( N726, new_n303_, keyIn_0_30 );
not g199 ( new_n305_, N13 );
and g200 ( new_n306_, new_n297_, new_n155_ );
xnor g201 ( new_n307_, new_n306_, new_n305_ );
nand g202 ( new_n308_, new_n307_, keyIn_0_31 );
not g203 ( new_n309_, keyIn_0_31 );
xnor g204 ( new_n310_, new_n306_, N13 );
nand g205 ( new_n311_, new_n310_, new_n309_ );
nand g206 ( N727, new_n308_, new_n311_ );
nor g207 ( new_n313_, new_n293_, new_n269_ );
and g208 ( new_n314_, new_n170_, new_n313_ );
not g209 ( new_n315_, new_n217_ );
xnor g210 ( new_n316_, new_n214_, new_n315_ );
not g211 ( new_n317_, new_n247_ );
nand g212 ( new_n318_, new_n316_, new_n317_ );
not g213 ( new_n319_, new_n318_ );
nand g214 ( new_n320_, new_n314_, new_n319_ );
nor g215 ( new_n321_, new_n320_, new_n119_ );
xnor g216 ( N728, new_n321_, new_n228_ );
nor g217 ( new_n323_, new_n320_, new_n136_ );
xnor g218 ( N729, new_n323_, new_n226_ );
not g219 ( new_n325_, new_n144_ );
nor g220 ( new_n326_, new_n320_, new_n325_ );
xnor g221 ( new_n327_, new_n326_, keyIn_0_25 );
xnor g222 ( N730, new_n327_, N25 );
nor g223 ( new_n329_, new_n320_, new_n154_ );
xnor g224 ( new_n330_, new_n329_, keyIn_0_26 );
xor g225 ( N731, new_n330_, N29 );
xnor g226 ( new_n332_, new_n290_, new_n285_ );
xnor g227 ( new_n333_, new_n247_, keyIn_0_16 );
xnor g228 ( new_n334_, new_n264_, new_n267_ );
nor g229 ( new_n335_, new_n316_, new_n334_ );
nand g230 ( new_n336_, new_n335_, new_n333_ );
nor g231 ( new_n337_, new_n332_, new_n336_ );
nand g232 ( new_n338_, new_n170_, new_n337_ );
nor g233 ( new_n339_, new_n338_, new_n119_ );
xnor g234 ( N732, new_n339_, new_n191_ );
nor g235 ( new_n341_, new_n338_, new_n136_ );
xnor g236 ( N733, new_n341_, new_n189_ );
nor g237 ( new_n343_, new_n338_, new_n325_ );
xnor g238 ( N734, new_n343_, new_n178_ );
nor g239 ( new_n345_, new_n338_, new_n154_ );
xnor g240 ( N735, new_n345_, new_n176_ );
not g241 ( new_n347_, new_n314_ );
xor g242 ( new_n348_, new_n247_, keyIn_0_17 );
nand g243 ( new_n349_, new_n348_, new_n218_ );
nor g244 ( new_n350_, new_n347_, new_n349_ );
nand g245 ( new_n351_, new_n350_, new_n120_ );
xnor g246 ( N736, new_n351_, N49 );
nand g247 ( new_n353_, new_n350_, new_n135_ );
xnor g248 ( N737, new_n353_, N53 );
nand g249 ( new_n355_, new_n350_, new_n144_ );
xnor g250 ( N738, new_n355_, N57 );
nand g251 ( new_n357_, new_n350_, new_n155_ );
xnor g252 ( N739, new_n357_, N61 );
nor g253 ( new_n359_, new_n218_, new_n317_ );
nand g254 ( new_n360_, new_n313_, new_n359_ );
xnor g255 ( new_n361_, new_n360_, keyIn_0_20 );
and g256 ( new_n362_, new_n359_, new_n269_ );
nand g257 ( new_n363_, new_n362_, new_n293_ );
xor g258 ( new_n364_, new_n363_, keyIn_0_21 );
nand g259 ( new_n365_, new_n218_, new_n269_ );
nor g260 ( new_n366_, new_n365_, new_n317_ );
nand g261 ( new_n367_, new_n332_, new_n366_ );
nand g262 ( new_n368_, new_n367_, keyIn_0_22 );
not g263 ( new_n369_, keyIn_0_22 );
nand g264 ( new_n370_, new_n335_, new_n247_ );
nor g265 ( new_n371_, new_n370_, new_n293_ );
nand g266 ( new_n372_, new_n371_, new_n369_ );
nand g267 ( new_n373_, new_n372_, new_n368_ );
or g268 ( new_n374_, new_n293_, keyIn_0_18 );
nand g269 ( new_n375_, new_n293_, keyIn_0_18 );
nor g270 ( new_n376_, new_n318_, new_n334_ );
and g271 ( new_n377_, new_n375_, new_n376_ );
nand g272 ( new_n378_, new_n377_, new_n374_ );
nand g273 ( new_n379_, new_n378_, new_n373_ );
nor g274 ( new_n380_, new_n364_, new_n379_ );
nand g275 ( new_n381_, new_n380_, new_n361_ );
xnor g276 ( new_n382_, new_n381_, keyIn_0_23 );
nand g277 ( new_n383_, new_n382_, new_n317_ );
nor g278 ( new_n384_, new_n325_, new_n155_ );
nor g279 ( new_n385_, new_n135_, new_n119_ );
nand g280 ( new_n386_, new_n384_, new_n385_ );
nor g281 ( new_n387_, new_n383_, new_n386_ );
xor g282 ( N740, new_n387_, N65 );
nand g283 ( new_n389_, new_n382_, new_n218_ );
nor g284 ( new_n390_, new_n389_, new_n386_ );
xor g285 ( N741, new_n390_, N69 );
nand g286 ( new_n392_, new_n382_, new_n293_ );
nor g287 ( new_n393_, new_n392_, new_n386_ );
xor g288 ( N742, new_n393_, N73 );
nand g289 ( new_n395_, new_n382_, new_n334_ );
nor g290 ( new_n396_, new_n395_, new_n386_ );
xor g291 ( N743, new_n396_, N77 );
nand g292 ( new_n398_, new_n385_, new_n160_ );
nor g293 ( new_n399_, new_n383_, new_n398_ );
xor g294 ( N744, new_n399_, N81 );
not g295 ( new_n401_, N85 );
not g296 ( new_n402_, keyIn_0_27 );
not g297 ( new_n403_, new_n361_ );
xnor g298 ( new_n404_, new_n363_, keyIn_0_21 );
and g299 ( new_n405_, new_n378_, new_n373_ );
nand g300 ( new_n406_, new_n405_, new_n404_ );
nor g301 ( new_n407_, new_n406_, new_n403_ );
nand g302 ( new_n408_, new_n407_, keyIn_0_23 );
not g303 ( new_n409_, keyIn_0_23 );
nand g304 ( new_n410_, new_n381_, new_n409_ );
nand g305 ( new_n411_, new_n408_, new_n410_ );
nor g306 ( new_n412_, new_n411_, new_n316_ );
not g307 ( new_n413_, new_n398_ );
nand g308 ( new_n414_, new_n412_, new_n413_ );
nand g309 ( new_n415_, new_n414_, new_n402_ );
nor g310 ( new_n416_, new_n389_, new_n398_ );
nand g311 ( new_n417_, new_n416_, keyIn_0_27 );
nand g312 ( new_n418_, new_n417_, new_n415_ );
nand g313 ( new_n419_, new_n418_, new_n401_ );
xnor g314 ( new_n420_, new_n414_, keyIn_0_27 );
nand g315 ( new_n421_, new_n420_, N85 );
nand g316 ( N745, new_n421_, new_n419_ );
nor g317 ( new_n423_, new_n392_, new_n398_ );
xor g318 ( N746, new_n423_, N89 );
nor g319 ( new_n425_, new_n411_, new_n269_ );
nand g320 ( new_n426_, new_n425_, new_n413_ );
xnor g321 ( N747, new_n426_, N93 );
nor g322 ( new_n428_, new_n136_, new_n120_ );
nand g323 ( new_n429_, new_n428_, new_n384_ );
nor g324 ( new_n430_, new_n383_, new_n429_ );
xor g325 ( N748, new_n430_, N97 );
not g326 ( new_n432_, new_n429_ );
nand g327 ( new_n433_, new_n412_, new_n432_ );
xnor g328 ( N749, new_n433_, N101 );
nor g329 ( new_n435_, new_n392_, new_n429_ );
xor g330 ( N750, new_n435_, N105 );
not g331 ( new_n437_, N109 );
nand g332 ( new_n438_, new_n425_, new_n432_ );
nand g333 ( new_n439_, new_n438_, keyIn_0_28 );
not g334 ( new_n440_, keyIn_0_28 );
nor g335 ( new_n441_, new_n395_, new_n429_ );
nand g336 ( new_n442_, new_n441_, new_n440_ );
nand g337 ( new_n443_, new_n442_, new_n439_ );
nand g338 ( new_n444_, new_n443_, new_n437_ );
xnor g339 ( new_n445_, new_n438_, new_n440_ );
nand g340 ( new_n446_, new_n445_, N109 );
nand g341 ( N751, new_n446_, new_n444_ );
nand g342 ( new_n448_, new_n428_, new_n160_ );
nor g343 ( new_n449_, new_n383_, new_n448_ );
xor g344 ( N752, new_n449_, N113 );
not g345 ( new_n451_, new_n448_ );
nand g346 ( new_n452_, new_n412_, new_n451_ );
nand g347 ( new_n453_, new_n452_, keyIn_0_29 );
not g348 ( new_n454_, keyIn_0_29 );
nor g349 ( new_n455_, new_n389_, new_n448_ );
nand g350 ( new_n456_, new_n455_, new_n454_ );
nand g351 ( new_n457_, new_n456_, new_n453_ );
nand g352 ( new_n458_, new_n457_, N117 );
not g353 ( new_n459_, N117 );
xnor g354 ( new_n460_, new_n452_, new_n454_ );
nand g355 ( new_n461_, new_n460_, new_n459_ );
nand g356 ( N753, new_n461_, new_n458_ );
nor g357 ( new_n463_, new_n392_, new_n448_ );
xor g358 ( N754, new_n463_, N121 );
nand g359 ( new_n465_, new_n425_, new_n451_ );
xnor g360 ( N755, new_n465_, N125 );
endmodule