module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n720_, new_n620_, new_n368_, new_n738_, new_n439_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n679_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n735_, new_n500_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n716_, new_n153_, new_n701_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n321_, new_n715_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n562_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n480_, new_n625_, new_n730_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n687_, new_n370_, new_n689_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n757_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n108_, keyIn_0_36 );
not g001 ( new_n109_, N30 );
and g002 ( new_n110_, keyIn_0_4, N24 );
not g003 ( new_n111_, new_n110_ );
or g004 ( new_n112_, keyIn_0_4, N24 );
and g005 ( new_n113_, new_n111_, new_n112_ );
or g006 ( new_n114_, new_n113_, new_n109_ );
or g007 ( new_n115_, new_n114_, keyIn_0_21 );
and g008 ( new_n116_, new_n114_, keyIn_0_21 );
not g009 ( new_n117_, new_n116_ );
and g010 ( new_n118_, new_n117_, new_n115_ );
not g011 ( new_n119_, new_n118_ );
not g012 ( new_n120_, keyIn_0_26 );
not g013 ( new_n121_, N95 );
and g014 ( new_n122_, keyIn_0_14, N89 );
not g015 ( new_n123_, new_n122_ );
or g016 ( new_n124_, keyIn_0_14, N89 );
and g017 ( new_n125_, new_n123_, new_n124_ );
or g018 ( new_n126_, new_n125_, new_n121_ );
not g019 ( new_n127_, new_n126_ );
and g020 ( new_n128_, new_n127_, new_n120_ );
and g021 ( new_n129_, new_n126_, keyIn_0_26 );
or g022 ( new_n130_, new_n128_, new_n129_ );
not g023 ( new_n131_, N56 );
not g024 ( new_n132_, N50 );
and g025 ( new_n133_, new_n132_, keyIn_0_8 );
not g026 ( new_n134_, new_n133_ );
or g027 ( new_n135_, new_n132_, keyIn_0_8 );
and g028 ( new_n136_, new_n134_, new_n135_ );
or g029 ( new_n137_, new_n136_, new_n131_ );
not g030 ( new_n138_, new_n137_ );
and g031 ( new_n139_, new_n138_, keyIn_0_23 );
not g032 ( new_n140_, keyIn_0_23 );
and g033 ( new_n141_, new_n137_, new_n140_ );
or g034 ( new_n142_, new_n139_, new_n141_ );
and g035 ( new_n143_, new_n142_, new_n130_ );
and g036 ( new_n144_, new_n143_, new_n119_ );
or g037 ( new_n145_, keyIn_0_2, N11 );
not g038 ( new_n146_, N17 );
and g039 ( new_n147_, keyIn_0_2, N11 );
or g040 ( new_n148_, new_n147_, new_n146_ );
not g041 ( new_n149_, new_n148_ );
and g042 ( new_n150_, new_n149_, new_n145_ );
not g043 ( new_n151_, new_n150_ );
and g044 ( new_n152_, new_n151_, keyIn_0_20 );
or g045 ( new_n153_, new_n151_, keyIn_0_20 );
not g046 ( new_n154_, new_n153_ );
or g047 ( new_n155_, new_n154_, new_n152_ );
not g048 ( new_n156_, N69 );
and g049 ( new_n157_, keyIn_0_10, N63 );
not g050 ( new_n158_, new_n157_ );
or g051 ( new_n159_, keyIn_0_10, N63 );
and g052 ( new_n160_, new_n158_, new_n159_ );
or g053 ( new_n161_, new_n160_, new_n156_ );
not g054 ( new_n162_, new_n161_ );
and g055 ( new_n163_, new_n162_, keyIn_0_24 );
not g056 ( new_n164_, keyIn_0_24 );
and g057 ( new_n165_, new_n161_, new_n164_ );
or g058 ( new_n166_, new_n163_, new_n165_ );
and g059 ( new_n167_, new_n155_, new_n166_ );
not g060 ( new_n168_, keyIn_0_22 );
and g061 ( new_n169_, keyIn_0_6, N37 );
not g062 ( new_n170_, keyIn_0_6 );
not g063 ( new_n171_, N37 );
and g064 ( new_n172_, new_n170_, new_n171_ );
or g065 ( new_n173_, new_n172_, new_n169_ );
and g066 ( new_n174_, new_n173_, N43 );
and g067 ( new_n175_, new_n174_, new_n168_ );
not g068 ( new_n176_, N43 );
not g069 ( new_n177_, new_n169_ );
or g070 ( new_n178_, keyIn_0_6, N37 );
and g071 ( new_n179_, new_n177_, new_n178_ );
or g072 ( new_n180_, new_n179_, new_n176_ );
and g073 ( new_n181_, new_n180_, keyIn_0_22 );
or g074 ( new_n182_, new_n175_, new_n181_ );
or g075 ( new_n183_, keyIn_0_0, N1 );
not g076 ( new_n184_, new_n183_ );
not g077 ( new_n185_, N4 );
and g078 ( new_n186_, keyIn_0_0, N1 );
or g079 ( new_n187_, new_n186_, new_n185_ );
or g080 ( new_n188_, new_n187_, new_n184_ );
and g081 ( new_n189_, new_n188_, keyIn_0_18 );
not g082 ( new_n190_, keyIn_0_18 );
not g083 ( new_n191_, new_n186_ );
and g084 ( new_n192_, new_n191_, N4 );
and g085 ( new_n193_, new_n192_, new_n183_ );
and g086 ( new_n194_, new_n193_, new_n190_ );
or g087 ( new_n195_, new_n194_, new_n189_ );
and g088 ( new_n196_, new_n182_, new_n195_ );
not g089 ( new_n197_, keyIn_0_27 );
and g090 ( new_n198_, keyIn_0_16, N102 );
not g091 ( new_n199_, new_n198_ );
or g092 ( new_n200_, keyIn_0_16, N102 );
and g093 ( new_n201_, new_n200_, N108 );
and g094 ( new_n202_, new_n201_, new_n199_ );
and g095 ( new_n203_, new_n202_, new_n197_ );
not g096 ( new_n204_, new_n202_ );
and g097 ( new_n205_, new_n204_, keyIn_0_27 );
or g098 ( new_n206_, new_n205_, new_n203_ );
not g099 ( new_n207_, keyIn_0_25 );
and g100 ( new_n208_, keyIn_0_12, N76 );
not g101 ( new_n209_, keyIn_0_12 );
not g102 ( new_n210_, N76 );
and g103 ( new_n211_, new_n209_, new_n210_ );
or g104 ( new_n212_, new_n211_, new_n208_ );
and g105 ( new_n213_, new_n212_, N82 );
and g106 ( new_n214_, new_n213_, new_n207_ );
not g107 ( new_n215_, N82 );
not g108 ( new_n216_, new_n208_ );
or g109 ( new_n217_, keyIn_0_12, N76 );
and g110 ( new_n218_, new_n216_, new_n217_ );
or g111 ( new_n219_, new_n218_, new_n215_ );
and g112 ( new_n220_, new_n219_, keyIn_0_25 );
or g113 ( new_n221_, new_n214_, new_n220_ );
and g114 ( new_n222_, new_n221_, new_n206_ );
and g115 ( new_n223_, new_n196_, new_n222_ );
and g116 ( new_n224_, new_n223_, new_n167_ );
and g117 ( new_n225_, new_n224_, new_n144_ );
and g118 ( new_n226_, new_n225_, new_n108_ );
not g119 ( new_n227_, new_n130_ );
or g120 ( new_n228_, new_n137_, new_n140_ );
not g121 ( new_n229_, new_n141_ );
and g122 ( new_n230_, new_n229_, new_n228_ );
or g123 ( new_n231_, new_n227_, new_n230_ );
or g124 ( new_n232_, new_n231_, new_n118_ );
not g125 ( new_n233_, new_n152_ );
and g126 ( new_n234_, new_n233_, new_n153_ );
not g127 ( new_n235_, new_n166_ );
or g128 ( new_n236_, new_n235_, new_n234_ );
or g129 ( new_n237_, new_n180_, keyIn_0_22 );
or g130 ( new_n238_, new_n174_, new_n168_ );
and g131 ( new_n239_, new_n237_, new_n238_ );
or g132 ( new_n240_, new_n193_, new_n190_ );
or g133 ( new_n241_, new_n188_, keyIn_0_18 );
and g134 ( new_n242_, new_n240_, new_n241_ );
or g135 ( new_n243_, new_n239_, new_n242_ );
not g136 ( new_n244_, new_n203_ );
or g137 ( new_n245_, new_n202_, new_n197_ );
and g138 ( new_n246_, new_n244_, new_n245_ );
or g139 ( new_n247_, new_n219_, keyIn_0_25 );
or g140 ( new_n248_, new_n213_, new_n207_ );
and g141 ( new_n249_, new_n247_, new_n248_ );
or g142 ( new_n250_, new_n249_, new_n246_ );
or g143 ( new_n251_, new_n250_, new_n243_ );
or g144 ( new_n252_, new_n251_, new_n236_ );
or g145 ( new_n253_, new_n252_, new_n232_ );
and g146 ( new_n254_, new_n253_, keyIn_0_36 );
or g147 ( N223, new_n254_, new_n226_ );
not g148 ( new_n256_, keyIn_0_37 );
and g149 ( new_n257_, N223, new_n256_ );
not g150 ( new_n258_, new_n226_ );
or g151 ( new_n259_, new_n225_, new_n108_ );
and g152 ( new_n260_, new_n258_, new_n259_ );
and g153 ( new_n261_, new_n260_, keyIn_0_37 );
or g154 ( new_n262_, new_n257_, new_n261_ );
and g155 ( new_n263_, new_n262_, new_n155_ );
or g156 ( new_n264_, new_n260_, keyIn_0_37 );
or g157 ( new_n265_, N223, new_n256_ );
and g158 ( new_n266_, new_n265_, new_n264_ );
and g159 ( new_n267_, new_n266_, new_n234_ );
or g160 ( new_n268_, new_n263_, new_n267_ );
and g161 ( new_n269_, new_n268_, keyIn_0_39 );
not g162 ( new_n270_, new_n269_ );
or g163 ( new_n271_, new_n268_, keyIn_0_39 );
and g164 ( new_n272_, new_n270_, new_n271_ );
not g165 ( new_n273_, N21 );
and g166 ( new_n274_, keyIn_0_3, N17 );
not g167 ( new_n275_, new_n274_ );
or g168 ( new_n276_, keyIn_0_3, N17 );
and g169 ( new_n277_, new_n275_, new_n276_ );
and g170 ( new_n278_, new_n277_, new_n273_ );
not g171 ( new_n279_, new_n278_ );
and g172 ( new_n280_, new_n279_, keyIn_0_28 );
not g173 ( new_n281_, new_n280_ );
or g174 ( new_n282_, new_n279_, keyIn_0_28 );
and g175 ( new_n283_, new_n281_, new_n282_ );
and g176 ( new_n284_, new_n272_, new_n283_ );
not g177 ( new_n285_, new_n284_ );
and g178 ( new_n286_, new_n285_, keyIn_0_48 );
not g179 ( new_n287_, keyIn_0_48 );
and g180 ( new_n288_, new_n284_, new_n287_ );
or g181 ( new_n289_, new_n286_, new_n288_ );
not g182 ( new_n290_, keyIn_0_42 );
and g183 ( new_n291_, new_n262_, new_n142_ );
and g184 ( new_n292_, new_n266_, new_n230_ );
or g185 ( new_n293_, new_n291_, new_n292_ );
and g186 ( new_n294_, new_n293_, new_n290_ );
not g187 ( new_n295_, new_n294_ );
or g188 ( new_n296_, new_n293_, new_n290_ );
and g189 ( new_n297_, new_n295_, new_n296_ );
not g190 ( new_n298_, N60 );
and g191 ( new_n299_, keyIn_0_9, N56 );
not g192 ( new_n300_, new_n299_ );
or g193 ( new_n301_, keyIn_0_9, N56 );
and g194 ( new_n302_, new_n300_, new_n301_ );
and g195 ( new_n303_, new_n302_, new_n298_ );
not g196 ( new_n304_, new_n303_ );
and g197 ( new_n305_, new_n304_, keyIn_0_31 );
not g198 ( new_n306_, new_n305_ );
or g199 ( new_n307_, new_n304_, keyIn_0_31 );
and g200 ( new_n308_, new_n306_, new_n307_ );
or g201 ( new_n309_, new_n297_, new_n308_ );
not g202 ( new_n310_, new_n309_ );
and g203 ( new_n311_, new_n310_, keyIn_0_51 );
not g204 ( new_n312_, keyIn_0_51 );
and g205 ( new_n313_, new_n309_, new_n312_ );
or g206 ( new_n314_, new_n311_, new_n313_ );
and g207 ( new_n315_, new_n262_, new_n221_ );
and g208 ( new_n316_, new_n266_, new_n249_ );
or g209 ( new_n317_, new_n315_, new_n316_ );
and g210 ( new_n318_, new_n317_, keyIn_0_44 );
not g211 ( new_n319_, new_n318_ );
or g212 ( new_n320_, new_n317_, keyIn_0_44 );
and g213 ( new_n321_, new_n319_, new_n320_ );
or g214 ( new_n322_, keyIn_0_13, N82 );
not g215 ( new_n323_, N86 );
and g216 ( new_n324_, keyIn_0_13, N82 );
not g217 ( new_n325_, new_n324_ );
and g218 ( new_n326_, new_n325_, new_n323_ );
and g219 ( new_n327_, new_n326_, new_n322_ );
and g220 ( new_n328_, new_n327_, keyIn_0_33 );
not g221 ( new_n329_, new_n328_ );
or g222 ( new_n330_, new_n327_, keyIn_0_33 );
and g223 ( new_n331_, new_n329_, new_n330_ );
or g224 ( new_n332_, new_n321_, new_n331_ );
not g225 ( new_n333_, new_n332_ );
and g226 ( new_n334_, new_n333_, keyIn_0_53 );
not g227 ( new_n335_, keyIn_0_53 );
and g228 ( new_n336_, new_n332_, new_n335_ );
or g229 ( new_n337_, new_n334_, new_n336_ );
and g230 ( new_n338_, new_n314_, new_n337_ );
and g231 ( new_n339_, new_n338_, new_n289_ );
not g232 ( new_n340_, keyIn_0_50 );
not g233 ( new_n341_, keyIn_0_41 );
and g234 ( new_n342_, new_n262_, new_n182_ );
and g235 ( new_n343_, new_n266_, new_n239_ );
or g236 ( new_n344_, new_n342_, new_n343_ );
and g237 ( new_n345_, new_n344_, new_n341_ );
not g238 ( new_n346_, new_n345_ );
or g239 ( new_n347_, new_n344_, new_n341_ );
and g240 ( new_n348_, new_n346_, new_n347_ );
not g241 ( new_n349_, N47 );
and g242 ( new_n350_, keyIn_0_7, N43 );
not g243 ( new_n351_, new_n350_ );
or g244 ( new_n352_, keyIn_0_7, N43 );
and g245 ( new_n353_, new_n351_, new_n352_ );
not g246 ( new_n354_, new_n353_ );
and g247 ( new_n355_, new_n354_, new_n349_ );
not g248 ( new_n356_, new_n355_ );
and g249 ( new_n357_, new_n356_, keyIn_0_30 );
not g250 ( new_n358_, new_n357_ );
or g251 ( new_n359_, new_n356_, keyIn_0_30 );
and g252 ( new_n360_, new_n358_, new_n359_ );
or g253 ( new_n361_, new_n348_, new_n360_ );
not g254 ( new_n362_, new_n361_ );
and g255 ( new_n363_, new_n362_, new_n340_ );
and g256 ( new_n364_, new_n361_, keyIn_0_50 );
or g257 ( new_n365_, new_n363_, new_n364_ );
not g258 ( new_n366_, keyIn_0_54 );
and g259 ( new_n367_, new_n262_, new_n130_ );
and g260 ( new_n368_, new_n266_, new_n227_ );
or g261 ( new_n369_, new_n367_, new_n368_ );
and g262 ( new_n370_, new_n369_, keyIn_0_45 );
not g263 ( new_n371_, new_n370_ );
or g264 ( new_n372_, new_n369_, keyIn_0_45 );
and g265 ( new_n373_, new_n371_, new_n372_ );
not g266 ( new_n374_, N99 );
and g267 ( new_n375_, keyIn_0_15, N95 );
not g268 ( new_n376_, new_n375_ );
or g269 ( new_n377_, keyIn_0_15, N95 );
and g270 ( new_n378_, new_n376_, new_n377_ );
not g271 ( new_n379_, new_n378_ );
and g272 ( new_n380_, new_n379_, new_n374_ );
and g273 ( new_n381_, new_n380_, keyIn_0_34 );
not g274 ( new_n382_, new_n381_ );
or g275 ( new_n383_, new_n380_, keyIn_0_34 );
and g276 ( new_n384_, new_n382_, new_n383_ );
or g277 ( new_n385_, new_n373_, new_n384_ );
not g278 ( new_n386_, new_n385_ );
and g279 ( new_n387_, new_n386_, new_n366_ );
and g280 ( new_n388_, new_n385_, keyIn_0_54 );
or g281 ( new_n389_, new_n387_, new_n388_ );
and g282 ( new_n390_, new_n365_, new_n389_ );
and g283 ( new_n391_, new_n262_, new_n206_ );
and g284 ( new_n392_, new_n266_, new_n246_ );
or g285 ( new_n393_, new_n391_, new_n392_ );
and g286 ( new_n394_, new_n393_, keyIn_0_46 );
not g287 ( new_n395_, keyIn_0_46 );
or g288 ( new_n396_, new_n266_, new_n246_ );
or g289 ( new_n397_, new_n262_, new_n206_ );
and g290 ( new_n398_, new_n397_, new_n396_ );
and g291 ( new_n399_, new_n398_, new_n395_ );
or g292 ( new_n400_, new_n394_, new_n399_ );
not g293 ( new_n401_, keyIn_0_35 );
not g294 ( new_n402_, N112 );
and g295 ( new_n403_, keyIn_0_17, N108 );
not g296 ( new_n404_, new_n403_ );
or g297 ( new_n405_, keyIn_0_17, N108 );
and g298 ( new_n406_, new_n404_, new_n405_ );
not g299 ( new_n407_, new_n406_ );
and g300 ( new_n408_, new_n407_, new_n402_ );
and g301 ( new_n409_, new_n408_, new_n401_ );
not g302 ( new_n410_, new_n409_ );
or g303 ( new_n411_, new_n408_, new_n401_ );
and g304 ( new_n412_, new_n410_, new_n411_ );
not g305 ( new_n413_, new_n412_ );
and g306 ( new_n414_, new_n400_, new_n413_ );
and g307 ( new_n415_, new_n414_, keyIn_0_55 );
not g308 ( new_n416_, keyIn_0_55 );
or g309 ( new_n417_, new_n398_, new_n395_ );
or g310 ( new_n418_, new_n393_, keyIn_0_46 );
and g311 ( new_n419_, new_n418_, new_n417_ );
or g312 ( new_n420_, new_n419_, new_n412_ );
and g313 ( new_n421_, new_n420_, new_n416_ );
or g314 ( new_n422_, new_n421_, new_n415_ );
not g315 ( new_n423_, keyIn_0_47 );
and g316 ( new_n424_, new_n262_, new_n195_ );
and g317 ( new_n425_, new_n266_, new_n242_ );
or g318 ( new_n426_, new_n424_, new_n425_ );
and g319 ( new_n427_, new_n426_, keyIn_0_38 );
not g320 ( new_n428_, keyIn_0_38 );
or g321 ( new_n429_, new_n266_, new_n242_ );
or g322 ( new_n430_, new_n262_, new_n195_ );
and g323 ( new_n431_, new_n430_, new_n429_ );
and g324 ( new_n432_, new_n431_, new_n428_ );
or g325 ( new_n433_, new_n427_, new_n432_ );
not g326 ( new_n434_, keyIn_0_19 );
and g327 ( new_n435_, new_n185_, keyIn_0_1 );
not g328 ( new_n436_, new_n435_ );
or g329 ( new_n437_, new_n185_, keyIn_0_1 );
and g330 ( new_n438_, new_n436_, new_n437_ );
not g331 ( new_n439_, new_n438_ );
or g332 ( new_n440_, new_n439_, N8 );
and g333 ( new_n441_, new_n440_, new_n434_ );
not g334 ( new_n442_, new_n441_ );
or g335 ( new_n443_, new_n440_, new_n434_ );
and g336 ( new_n444_, new_n442_, new_n443_ );
not g337 ( new_n445_, new_n444_ );
and g338 ( new_n446_, new_n433_, new_n445_ );
and g339 ( new_n447_, new_n446_, new_n423_ );
or g340 ( new_n448_, new_n431_, new_n428_ );
or g341 ( new_n449_, new_n426_, keyIn_0_38 );
and g342 ( new_n450_, new_n449_, new_n448_ );
or g343 ( new_n451_, new_n450_, new_n444_ );
and g344 ( new_n452_, new_n451_, keyIn_0_47 );
or g345 ( new_n453_, new_n452_, new_n447_ );
and g346 ( new_n454_, new_n422_, new_n453_ );
not g347 ( new_n455_, keyIn_0_52 );
not g348 ( new_n456_, keyIn_0_43 );
and g349 ( new_n457_, new_n262_, new_n166_ );
and g350 ( new_n458_, new_n266_, new_n235_ );
or g351 ( new_n459_, new_n457_, new_n458_ );
and g352 ( new_n460_, new_n459_, new_n456_ );
or g353 ( new_n461_, new_n266_, new_n235_ );
or g354 ( new_n462_, new_n262_, new_n166_ );
and g355 ( new_n463_, new_n462_, new_n461_ );
and g356 ( new_n464_, new_n463_, keyIn_0_43 );
or g357 ( new_n465_, new_n460_, new_n464_ );
not g358 ( new_n466_, keyIn_0_32 );
not g359 ( new_n467_, N73 );
and g360 ( new_n468_, keyIn_0_11, N69 );
not g361 ( new_n469_, new_n468_ );
or g362 ( new_n470_, keyIn_0_11, N69 );
and g363 ( new_n471_, new_n469_, new_n470_ );
and g364 ( new_n472_, new_n471_, new_n467_ );
not g365 ( new_n473_, new_n472_ );
and g366 ( new_n474_, new_n473_, new_n466_ );
and g367 ( new_n475_, new_n472_, keyIn_0_32 );
or g368 ( new_n476_, new_n474_, new_n475_ );
and g369 ( new_n477_, new_n465_, new_n476_ );
and g370 ( new_n478_, new_n477_, new_n455_ );
or g371 ( new_n479_, new_n463_, keyIn_0_43 );
or g372 ( new_n480_, new_n459_, new_n456_ );
and g373 ( new_n481_, new_n480_, new_n479_ );
not g374 ( new_n482_, new_n476_ );
or g375 ( new_n483_, new_n481_, new_n482_ );
and g376 ( new_n484_, new_n483_, keyIn_0_52 );
or g377 ( new_n485_, new_n484_, new_n478_ );
not g378 ( new_n486_, keyIn_0_40 );
and g379 ( new_n487_, new_n262_, new_n119_ );
and g380 ( new_n488_, new_n266_, new_n118_ );
or g381 ( new_n489_, new_n487_, new_n488_ );
and g382 ( new_n490_, new_n489_, new_n486_ );
or g383 ( new_n491_, new_n266_, new_n118_ );
or g384 ( new_n492_, new_n262_, new_n119_ );
and g385 ( new_n493_, new_n492_, new_n491_ );
and g386 ( new_n494_, new_n493_, keyIn_0_40 );
or g387 ( new_n495_, new_n490_, new_n494_ );
not g388 ( new_n496_, N34 );
and g389 ( new_n497_, keyIn_0_5, N30 );
not g390 ( new_n498_, new_n497_ );
or g391 ( new_n499_, keyIn_0_5, N30 );
and g392 ( new_n500_, new_n498_, new_n499_ );
and g393 ( new_n501_, new_n500_, new_n496_ );
not g394 ( new_n502_, new_n501_ );
and g395 ( new_n503_, new_n502_, keyIn_0_29 );
not g396 ( new_n504_, new_n503_ );
or g397 ( new_n505_, new_n502_, keyIn_0_29 );
and g398 ( new_n506_, new_n504_, new_n505_ );
not g399 ( new_n507_, new_n506_ );
and g400 ( new_n508_, new_n495_, new_n507_ );
and g401 ( new_n509_, new_n508_, keyIn_0_49 );
not g402 ( new_n510_, keyIn_0_49 );
or g403 ( new_n511_, new_n493_, keyIn_0_40 );
or g404 ( new_n512_, new_n489_, new_n486_ );
and g405 ( new_n513_, new_n512_, new_n511_ );
or g406 ( new_n514_, new_n513_, new_n506_ );
and g407 ( new_n515_, new_n514_, new_n510_ );
or g408 ( new_n516_, new_n515_, new_n509_ );
and g409 ( new_n517_, new_n485_, new_n516_ );
and g410 ( new_n518_, new_n454_, new_n517_ );
and g411 ( new_n519_, new_n518_, new_n390_ );
and g412 ( new_n520_, new_n519_, new_n339_ );
and g413 ( new_n521_, new_n520_, keyIn_0_60 );
not g414 ( new_n522_, keyIn_0_60 );
not g415 ( new_n523_, new_n520_ );
and g416 ( new_n524_, new_n523_, new_n522_ );
or g417 ( N329, new_n524_, new_n521_ );
not g418 ( new_n526_, new_n422_ );
not g419 ( new_n527_, keyIn_0_61 );
not g420 ( new_n528_, new_n521_ );
or g421 ( new_n529_, new_n520_, keyIn_0_60 );
and g422 ( new_n530_, new_n528_, new_n529_ );
or g423 ( new_n531_, new_n530_, new_n527_ );
and g424 ( new_n532_, new_n530_, new_n527_ );
not g425 ( new_n533_, new_n532_ );
and g426 ( new_n534_, new_n533_, new_n531_ );
and g427 ( new_n535_, new_n534_, new_n526_ );
and g428 ( new_n536_, N329, keyIn_0_61 );
or g429 ( new_n537_, new_n536_, new_n532_ );
and g430 ( new_n538_, new_n537_, new_n422_ );
not g431 ( new_n539_, keyIn_0_59 );
not g432 ( new_n540_, N115 );
and g433 ( new_n541_, new_n407_, new_n540_ );
and g434 ( new_n542_, new_n400_, new_n541_ );
and g435 ( new_n543_, new_n542_, new_n539_ );
not g436 ( new_n544_, new_n543_ );
or g437 ( new_n545_, new_n542_, new_n539_ );
and g438 ( new_n546_, new_n544_, new_n545_ );
not g439 ( new_n547_, new_n546_ );
or g440 ( new_n548_, new_n538_, new_n547_ );
or g441 ( new_n549_, new_n548_, new_n535_ );
not g442 ( new_n550_, new_n516_ );
and g443 ( new_n551_, new_n534_, new_n550_ );
not g444 ( new_n552_, new_n551_ );
and g445 ( new_n553_, new_n537_, new_n516_ );
not g446 ( new_n554_, new_n553_ );
not g447 ( new_n555_, N40 );
and g448 ( new_n556_, new_n500_, new_n555_ );
and g449 ( new_n557_, new_n495_, new_n556_ );
and g450 ( new_n558_, new_n554_, new_n557_ );
and g451 ( new_n559_, new_n558_, new_n552_ );
not g452 ( new_n560_, new_n389_ );
and g453 ( new_n561_, new_n534_, new_n560_ );
not g454 ( new_n562_, new_n561_ );
and g455 ( new_n563_, new_n537_, new_n389_ );
not g456 ( new_n564_, new_n563_ );
not g457 ( new_n565_, new_n373_ );
not g458 ( new_n566_, N105 );
and g459 ( new_n567_, new_n379_, new_n566_ );
and g460 ( new_n568_, new_n565_, new_n567_ );
and g461 ( new_n569_, new_n568_, keyIn_0_58 );
not g462 ( new_n570_, new_n569_ );
or g463 ( new_n571_, new_n568_, keyIn_0_58 );
and g464 ( new_n572_, new_n570_, new_n571_ );
and g465 ( new_n573_, new_n564_, new_n572_ );
and g466 ( new_n574_, new_n573_, new_n562_ );
or g467 ( new_n575_, new_n559_, new_n574_ );
not g468 ( new_n576_, new_n575_ );
and g469 ( new_n577_, new_n576_, new_n549_ );
not g470 ( new_n578_, new_n337_ );
and g471 ( new_n579_, new_n534_, new_n578_ );
not g472 ( new_n580_, new_n579_ );
and g473 ( new_n581_, new_n537_, new_n337_ );
not g474 ( new_n582_, new_n581_ );
not g475 ( new_n583_, keyIn_0_57 );
not g476 ( new_n584_, new_n321_ );
not g477 ( new_n585_, N92 );
and g478 ( new_n586_, new_n325_, new_n585_ );
and g479 ( new_n587_, new_n586_, new_n322_ );
and g480 ( new_n588_, new_n584_, new_n587_ );
and g481 ( new_n589_, new_n588_, new_n583_ );
not g482 ( new_n590_, new_n589_ );
or g483 ( new_n591_, new_n588_, new_n583_ );
and g484 ( new_n592_, new_n590_, new_n591_ );
and g485 ( new_n593_, new_n582_, new_n592_ );
and g486 ( new_n594_, new_n593_, new_n580_ );
not g487 ( new_n595_, new_n365_ );
and g488 ( new_n596_, new_n534_, new_n595_ );
not g489 ( new_n597_, new_n596_ );
and g490 ( new_n598_, new_n537_, new_n365_ );
not g491 ( new_n599_, new_n598_ );
not g492 ( new_n600_, new_n348_ );
not g493 ( new_n601_, N53 );
and g494 ( new_n602_, new_n354_, new_n601_ );
and g495 ( new_n603_, new_n600_, new_n602_ );
and g496 ( new_n604_, new_n599_, new_n603_ );
and g497 ( new_n605_, new_n604_, new_n597_ );
or g498 ( new_n606_, new_n594_, new_n605_ );
not g499 ( new_n607_, new_n606_ );
not g500 ( new_n608_, new_n314_ );
and g501 ( new_n609_, new_n534_, new_n608_ );
and g502 ( new_n610_, new_n537_, new_n314_ );
not g503 ( new_n611_, new_n297_ );
not g504 ( new_n612_, N66 );
and g505 ( new_n613_, new_n302_, new_n612_ );
and g506 ( new_n614_, new_n611_, new_n613_ );
not g507 ( new_n615_, new_n614_ );
or g508 ( new_n616_, new_n610_, new_n615_ );
or g509 ( new_n617_, new_n616_, new_n609_ );
not g510 ( new_n618_, new_n485_ );
and g511 ( new_n619_, new_n534_, new_n618_ );
and g512 ( new_n620_, new_n537_, new_n485_ );
not g513 ( new_n621_, keyIn_0_56 );
not g514 ( new_n622_, N79 );
and g515 ( new_n623_, new_n471_, new_n622_ );
and g516 ( new_n624_, new_n465_, new_n623_ );
and g517 ( new_n625_, new_n624_, new_n621_ );
not g518 ( new_n626_, new_n625_ );
or g519 ( new_n627_, new_n624_, new_n621_ );
and g520 ( new_n628_, new_n626_, new_n627_ );
not g521 ( new_n629_, new_n628_ );
or g522 ( new_n630_, new_n620_, new_n629_ );
or g523 ( new_n631_, new_n630_, new_n619_ );
and g524 ( new_n632_, new_n617_, new_n631_ );
not g525 ( new_n633_, new_n453_ );
and g526 ( new_n634_, new_n534_, new_n633_ );
and g527 ( new_n635_, new_n537_, new_n453_ );
or g528 ( new_n636_, new_n439_, N14 );
or g529 ( new_n637_, new_n450_, new_n636_ );
or g530 ( new_n638_, new_n635_, new_n637_ );
or g531 ( new_n639_, new_n638_, new_n634_ );
not g532 ( new_n640_, new_n289_ );
and g533 ( new_n641_, new_n534_, new_n640_ );
and g534 ( new_n642_, new_n537_, new_n289_ );
not g535 ( new_n643_, N27 );
and g536 ( new_n644_, new_n277_, new_n643_ );
and g537 ( new_n645_, new_n272_, new_n644_ );
not g538 ( new_n646_, new_n645_ );
or g539 ( new_n647_, new_n642_, new_n646_ );
or g540 ( new_n648_, new_n647_, new_n641_ );
and g541 ( new_n649_, new_n639_, new_n648_ );
and g542 ( new_n650_, new_n632_, new_n649_ );
and g543 ( new_n651_, new_n650_, new_n607_ );
and g544 ( new_n652_, new_n651_, new_n577_ );
and g545 ( new_n653_, new_n652_, keyIn_0_62 );
or g546 ( new_n654_, new_n652_, keyIn_0_62 );
not g547 ( new_n655_, new_n654_ );
or g548 ( N370, new_n655_, new_n653_ );
not g549 ( new_n657_, keyIn_0_63 );
not g550 ( new_n658_, new_n653_ );
and g551 ( new_n659_, new_n658_, new_n654_ );
or g552 ( new_n660_, new_n659_, new_n643_ );
and g553 ( new_n661_, N329, N21 );
and g554 ( new_n662_, N223, N11 );
or g555 ( new_n663_, new_n662_, new_n146_ );
or g556 ( new_n664_, new_n661_, new_n663_ );
not g557 ( new_n665_, new_n664_ );
and g558 ( new_n666_, new_n660_, new_n665_ );
not g559 ( new_n667_, new_n666_ );
or g560 ( new_n668_, new_n659_, new_n555_ );
and g561 ( new_n669_, N329, N34 );
and g562 ( new_n670_, N223, N24 );
or g563 ( new_n671_, new_n670_, new_n109_ );
or g564 ( new_n672_, new_n669_, new_n671_ );
not g565 ( new_n673_, new_n672_ );
and g566 ( new_n674_, new_n668_, new_n673_ );
not g567 ( new_n675_, new_n674_ );
and g568 ( new_n676_, new_n667_, new_n675_ );
or g569 ( new_n677_, new_n659_, new_n601_ );
and g570 ( new_n678_, N329, N47 );
and g571 ( new_n679_, N223, N37 );
or g572 ( new_n680_, new_n679_, new_n176_ );
or g573 ( new_n681_, new_n678_, new_n680_ );
not g574 ( new_n682_, new_n681_ );
and g575 ( new_n683_, new_n677_, new_n682_ );
not g576 ( new_n684_, new_n683_ );
and g577 ( new_n685_, N370, N66 );
and g578 ( new_n686_, N329, N60 );
and g579 ( new_n687_, N223, N50 );
or g580 ( new_n688_, new_n687_, new_n131_ );
or g581 ( new_n689_, new_n686_, new_n688_ );
or g582 ( new_n690_, new_n685_, new_n689_ );
and g583 ( new_n691_, new_n684_, new_n690_ );
and g584 ( new_n692_, new_n676_, new_n691_ );
or g585 ( new_n693_, new_n659_, new_n566_ );
and g586 ( new_n694_, N329, N99 );
and g587 ( new_n695_, N223, N89 );
or g588 ( new_n696_, new_n695_, new_n121_ );
or g589 ( new_n697_, new_n694_, new_n696_ );
not g590 ( new_n698_, new_n697_ );
and g591 ( new_n699_, new_n693_, new_n698_ );
not g592 ( new_n700_, new_n699_ );
and g593 ( new_n701_, N370, N115 );
and g594 ( new_n702_, N329, N112 );
not g595 ( new_n703_, new_n702_ );
and g596 ( new_n704_, N223, N102 );
not g597 ( new_n705_, new_n704_ );
and g598 ( new_n706_, new_n705_, N108 );
and g599 ( new_n707_, new_n703_, new_n706_ );
not g600 ( new_n708_, new_n707_ );
or g601 ( new_n709_, new_n701_, new_n708_ );
and g602 ( new_n710_, new_n700_, new_n709_ );
and g603 ( new_n711_, N370, N79 );
and g604 ( new_n712_, N329, N73 );
and g605 ( new_n713_, N223, N63 );
or g606 ( new_n714_, new_n713_, new_n156_ );
or g607 ( new_n715_, new_n712_, new_n714_ );
or g608 ( new_n716_, new_n711_, new_n715_ );
and g609 ( new_n717_, N370, N92 );
and g610 ( new_n718_, N329, N86 );
and g611 ( new_n719_, N223, N76 );
or g612 ( new_n720_, new_n719_, new_n215_ );
or g613 ( new_n721_, new_n718_, new_n720_ );
or g614 ( new_n722_, new_n717_, new_n721_ );
and g615 ( new_n723_, new_n716_, new_n722_ );
and g616 ( new_n724_, new_n710_, new_n723_ );
and g617 ( new_n725_, new_n692_, new_n724_ );
and g618 ( new_n726_, new_n725_, new_n657_ );
or g619 ( new_n727_, new_n666_, new_n674_ );
or g620 ( new_n728_, new_n659_, new_n612_ );
not g621 ( new_n729_, new_n689_ );
and g622 ( new_n730_, new_n728_, new_n729_ );
or g623 ( new_n731_, new_n683_, new_n730_ );
or g624 ( N430, new_n727_, new_n731_ );
or g625 ( new_n733_, new_n659_, new_n540_ );
and g626 ( new_n734_, new_n733_, new_n707_ );
or g627 ( new_n735_, new_n699_, new_n734_ );
or g628 ( new_n736_, new_n659_, new_n622_ );
not g629 ( new_n737_, new_n715_ );
and g630 ( new_n738_, new_n736_, new_n737_ );
or g631 ( new_n739_, new_n659_, new_n585_ );
not g632 ( new_n740_, new_n721_ );
and g633 ( new_n741_, new_n739_, new_n740_ );
or g634 ( new_n742_, new_n738_, new_n741_ );
or g635 ( new_n743_, new_n735_, new_n742_ );
or g636 ( new_n744_, N430, new_n743_ );
and g637 ( new_n745_, new_n744_, keyIn_0_63 );
or g638 ( new_n746_, new_n745_, new_n726_ );
and g639 ( new_n747_, N370, N14 );
and g640 ( new_n748_, N329, N8 );
and g641 ( new_n749_, N223, N1 );
or g642 ( new_n750_, new_n749_, new_n185_ );
or g643 ( new_n751_, new_n748_, new_n750_ );
or g644 ( new_n752_, new_n747_, new_n751_ );
and g645 ( N421, new_n746_, new_n752_ );
and g646 ( new_n754_, new_n742_, new_n690_ );
and g647 ( new_n755_, new_n754_, new_n684_ );
or g648 ( N431, new_n755_, new_n727_ );
and g649 ( new_n757_, new_n722_, new_n699_ );
and g650 ( new_n758_, new_n690_, new_n738_ );
or g651 ( new_n759_, new_n758_, new_n683_ );
or g652 ( new_n760_, new_n759_, new_n757_ );
and g653 ( new_n761_, new_n760_, new_n675_ );
or g654 ( N432, new_n761_, new_n666_ );
endmodule