module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n214_, new_n451_, new_n114_, new_n188_, new_n240_, new_n211_, new_n123_, new_n127_, new_n342_, new_n317_, new_n344_, new_n287_, new_n427_, new_n234_, new_n472_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n212_, new_n364_, new_n449_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n248_, new_n350_, new_n117_, new_n167_, new_n385_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n388_, new_n194_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n165_, new_n441_, new_n216_, new_n280_, new_n235_, new_n398_, new_n301_, new_n169_, new_n383_, new_n343_, new_n210_, new_n458_, new_n207_, new_n267_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n126_, new_n177_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n145_, new_n253_, new_n403_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n107_, new_n182_, new_n151_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n112_, new_n121_, new_n221_, new_n243_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n174_, new_n354_, new_n392_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n203_, new_n316_, new_n332_, new_n163_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n115_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n327_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n128_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n434_, new_n200_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n120_, new_n406_, new_n356_, new_n229_, new_n204_, new_n181_, new_n135_, new_n405_;

not g000 ( new_n106_, N1 );
xor g001 ( new_n107_, N33, N49 );
xnor g002 ( new_n108_, N1, N17 );
xor g003 ( new_n109_, new_n107_, new_n108_ );
not g004 ( new_n110_, new_n109_ );
xor g005 ( new_n111_, N73, N77 );
xnor g006 ( new_n112_, N65, N69 );
xnor g007 ( new_n113_, new_n111_, new_n112_ );
xor g008 ( new_n114_, N81, N85 );
xnor g009 ( new_n115_, N89, N93 );
xnor g010 ( new_n116_, new_n114_, new_n115_ );
xnor g011 ( new_n117_, new_n113_, new_n116_ );
nand g012 ( new_n118_, N129, N137 );
xnor g013 ( new_n119_, new_n117_, new_n118_ );
xnor g014 ( new_n120_, new_n119_, new_n110_ );
not g015 ( new_n121_, keyIn_0_15 );
not g016 ( new_n122_, keyIn_0_13 );
not g017 ( new_n123_, keyIn_0_11 );
not g018 ( new_n124_, keyIn_0_9 );
not g019 ( new_n125_, N53 );
nand g020 ( new_n126_, new_n125_, N49 );
not g021 ( new_n127_, N49 );
nand g022 ( new_n128_, new_n127_, N53 );
nand g023 ( new_n129_, new_n126_, new_n128_ );
nand g024 ( new_n130_, new_n129_, keyIn_0_4 );
not g025 ( new_n131_, keyIn_0_4 );
nand g026 ( new_n132_, new_n126_, new_n128_, new_n131_ );
nand g027 ( new_n133_, new_n130_, new_n132_ );
not g028 ( new_n134_, keyIn_0_5 );
not g029 ( new_n135_, N61 );
nand g030 ( new_n136_, new_n135_, N57 );
not g031 ( new_n137_, N57 );
nand g032 ( new_n138_, new_n137_, N61 );
nand g033 ( new_n139_, new_n136_, new_n138_ );
nand g034 ( new_n140_, new_n139_, new_n134_ );
nand g035 ( new_n141_, new_n136_, new_n138_, keyIn_0_5 );
nand g036 ( new_n142_, new_n140_, new_n141_ );
nand g037 ( new_n143_, new_n133_, new_n142_ );
nand g038 ( new_n144_, new_n130_, new_n140_, new_n132_, new_n141_ );
nand g039 ( new_n145_, new_n143_, new_n144_ );
nand g040 ( new_n146_, new_n145_, keyIn_0_8 );
not g041 ( new_n147_, keyIn_0_8 );
nand g042 ( new_n148_, new_n143_, new_n147_, new_n144_ );
nand g043 ( new_n149_, new_n146_, new_n148_ );
not g044 ( new_n150_, keyIn_0_2 );
not g045 ( new_n151_, N37 );
nand g046 ( new_n152_, new_n151_, N33 );
not g047 ( new_n153_, N33 );
nand g048 ( new_n154_, new_n153_, N37 );
nand g049 ( new_n155_, new_n152_, new_n154_ );
nand g050 ( new_n156_, new_n155_, new_n150_ );
nand g051 ( new_n157_, new_n152_, new_n154_, keyIn_0_2 );
nand g052 ( new_n158_, new_n156_, new_n157_ );
not g053 ( new_n159_, keyIn_0_3 );
not g054 ( new_n160_, N45 );
nand g055 ( new_n161_, new_n160_, N41 );
not g056 ( new_n162_, N41 );
nand g057 ( new_n163_, new_n162_, N45 );
nand g058 ( new_n164_, new_n161_, new_n163_ );
nand g059 ( new_n165_, new_n164_, new_n159_ );
nand g060 ( new_n166_, new_n161_, new_n163_, keyIn_0_3 );
nand g061 ( new_n167_, new_n165_, new_n166_ );
nand g062 ( new_n168_, new_n158_, new_n167_ );
nand g063 ( new_n169_, new_n156_, new_n165_, new_n157_, new_n166_ );
nand g064 ( new_n170_, new_n168_, new_n169_ );
nand g065 ( new_n171_, new_n170_, keyIn_0_7 );
not g066 ( new_n172_, keyIn_0_7 );
nand g067 ( new_n173_, new_n168_, new_n172_, new_n169_ );
nand g068 ( new_n174_, new_n149_, new_n171_, new_n173_ );
nand g069 ( new_n175_, new_n171_, new_n173_ );
nand g070 ( new_n176_, new_n175_, new_n146_, new_n148_ );
nand g071 ( new_n177_, new_n174_, new_n176_ );
nand g072 ( new_n178_, new_n177_, new_n124_ );
nand g073 ( new_n179_, new_n174_, new_n176_, keyIn_0_9 );
nand g074 ( new_n180_, new_n178_, new_n179_ );
nand g075 ( new_n181_, N134, N137 );
nand g076 ( new_n182_, new_n180_, new_n181_ );
nand g077 ( new_n183_, new_n178_, N134, N137, new_n179_ );
nand g078 ( new_n184_, new_n182_, new_n183_ );
nand g079 ( new_n185_, new_n184_, new_n123_ );
nand g080 ( new_n186_, new_n182_, keyIn_0_11, new_n183_ );
nand g081 ( new_n187_, new_n185_, new_n186_ );
xor g082 ( new_n188_, N101, N117 );
xnor g083 ( new_n189_, N69, N85 );
xor g084 ( new_n190_, new_n188_, new_n189_ );
nand g085 ( new_n191_, new_n187_, new_n190_ );
not g086 ( new_n192_, new_n190_ );
nand g087 ( new_n193_, new_n185_, new_n186_, new_n192_ );
nand g088 ( new_n194_, new_n191_, new_n193_ );
nand g089 ( new_n195_, new_n194_, new_n122_ );
nand g090 ( new_n196_, new_n191_, keyIn_0_13, new_n193_ );
nand g091 ( new_n197_, new_n195_, new_n196_ );
nand g092 ( new_n198_, new_n197_, new_n121_ );
nand g093 ( new_n199_, new_n195_, keyIn_0_15, new_n196_ );
nand g094 ( new_n200_, new_n198_, new_n199_ );
not g095 ( new_n201_, keyIn_0_6 );
not g096 ( new_n202_, keyIn_0_0 );
not g097 ( new_n203_, N5 );
nand g098 ( new_n204_, new_n203_, N1 );
nand g099 ( new_n205_, new_n106_, N5 );
nand g100 ( new_n206_, new_n204_, new_n205_ );
nand g101 ( new_n207_, new_n206_, new_n202_ );
nand g102 ( new_n208_, new_n204_, new_n205_, keyIn_0_0 );
nand g103 ( new_n209_, new_n207_, new_n208_ );
not g104 ( new_n210_, N13 );
nand g105 ( new_n211_, new_n210_, N9 );
not g106 ( new_n212_, N9 );
nand g107 ( new_n213_, new_n212_, N13 );
nand g108 ( new_n214_, new_n211_, new_n213_ );
nand g109 ( new_n215_, new_n214_, keyIn_0_1 );
not g110 ( new_n216_, keyIn_0_1 );
nand g111 ( new_n217_, new_n211_, new_n213_, new_n216_ );
nand g112 ( new_n218_, new_n215_, new_n217_ );
nand g113 ( new_n219_, new_n209_, new_n218_ );
nand g114 ( new_n220_, new_n207_, new_n215_, new_n208_, new_n217_ );
nand g115 ( new_n221_, new_n219_, new_n220_ );
nand g116 ( new_n222_, new_n221_, new_n201_ );
nand g117 ( new_n223_, new_n219_, keyIn_0_6, new_n220_ );
nand g118 ( new_n224_, new_n222_, new_n223_ );
xnor g119 ( new_n225_, N25, N29 );
xnor g120 ( new_n226_, N17, N21 );
xnor g121 ( new_n227_, new_n225_, new_n226_ );
xor g122 ( new_n228_, new_n224_, new_n227_ );
nand g123 ( new_n229_, N133, N137 );
xnor g124 ( new_n230_, new_n228_, new_n229_ );
xnor g125 ( new_n231_, N97, N113 );
xnor g126 ( new_n232_, N65, N81 );
xnor g127 ( new_n233_, new_n231_, new_n232_ );
xnor g128 ( new_n234_, new_n230_, new_n233_ );
not g129 ( new_n235_, keyIn_0_17 );
xnor g130 ( new_n236_, new_n119_, new_n109_ );
xor g131 ( new_n237_, N121, N125 );
xnor g132 ( new_n238_, N113, N117 );
xnor g133 ( new_n239_, new_n237_, new_n238_ );
xor g134 ( new_n240_, N105, N109 );
xnor g135 ( new_n241_, N97, N101 );
xnor g136 ( new_n242_, new_n240_, new_n241_ );
xnor g137 ( new_n243_, new_n239_, new_n242_ );
nand g138 ( new_n244_, N130, N137 );
not g139 ( new_n245_, new_n244_ );
xnor g140 ( new_n246_, new_n243_, new_n245_ );
xor g141 ( new_n247_, N37, N53 );
xnor g142 ( new_n248_, N5, N21 );
xor g143 ( new_n249_, new_n247_, new_n248_ );
xnor g144 ( new_n250_, new_n246_, new_n249_ );
xnor g145 ( new_n251_, new_n113_, new_n242_ );
and g146 ( new_n252_, N131, N137 );
xnor g147 ( new_n253_, new_n251_, new_n252_ );
xor g148 ( new_n254_, N41, N57 );
xnor g149 ( new_n255_, N9, N25 );
xor g150 ( new_n256_, new_n254_, new_n255_ );
not g151 ( new_n257_, new_n256_ );
xnor g152 ( new_n258_, new_n253_, new_n257_ );
nand g153 ( new_n259_, new_n236_, new_n250_, new_n258_ );
not g154 ( new_n260_, new_n249_ );
xnor g155 ( new_n261_, new_n246_, new_n260_ );
nand g156 ( new_n262_, new_n120_, new_n258_, new_n261_ );
nand g157 ( new_n263_, new_n259_, new_n262_ );
xor g158 ( new_n264_, new_n116_, new_n239_ );
nand g159 ( new_n265_, N132, N137 );
xnor g160 ( new_n266_, new_n264_, new_n265_ );
xor g161 ( new_n267_, N45, N61 );
xnor g162 ( new_n268_, N13, N29 );
xor g163 ( new_n269_, new_n267_, new_n268_ );
nand g164 ( new_n270_, new_n266_, new_n269_ );
or g165 ( new_n271_, new_n264_, new_n265_ );
nand g166 ( new_n272_, new_n264_, new_n265_ );
not g167 ( new_n273_, new_n269_ );
nand g168 ( new_n274_, new_n271_, new_n272_, new_n273_ );
and g169 ( new_n275_, new_n270_, new_n274_ );
nand g170 ( new_n276_, new_n263_, new_n275_ );
nand g171 ( new_n277_, new_n270_, new_n274_ );
nand g172 ( new_n278_, new_n258_, new_n277_ );
xnor g173 ( new_n279_, new_n253_, new_n256_ );
nand g174 ( new_n280_, new_n275_, new_n279_ );
nand g175 ( new_n281_, new_n280_, new_n278_ );
nor g176 ( new_n282_, new_n120_, new_n250_ );
nand g177 ( new_n283_, new_n281_, new_n282_ );
nand g178 ( new_n284_, new_n276_, new_n283_ );
nand g179 ( new_n285_, new_n284_, new_n235_ );
nand g180 ( new_n286_, new_n276_, new_n283_, keyIn_0_17 );
and g181 ( new_n287_, new_n285_, new_n234_, new_n286_ );
not g182 ( new_n288_, keyIn_0_12 );
not g183 ( new_n289_, keyIn_0_10 );
nand g184 ( new_n290_, new_n224_, new_n171_, new_n173_ );
nand g185 ( new_n291_, new_n175_, new_n222_, new_n223_ );
nand g186 ( new_n292_, new_n290_, new_n291_ );
nand g187 ( new_n293_, new_n292_, new_n289_ );
nand g188 ( new_n294_, new_n290_, new_n291_, keyIn_0_10 );
nand g189 ( new_n295_, new_n293_, new_n294_ );
nand g190 ( new_n296_, N135, N137 );
not g191 ( new_n297_, new_n296_ );
nand g192 ( new_n298_, new_n295_, new_n297_ );
nand g193 ( new_n299_, new_n293_, new_n294_, new_n296_ );
nand g194 ( new_n300_, new_n298_, new_n299_ );
nand g195 ( new_n301_, new_n300_, new_n288_ );
nand g196 ( new_n302_, new_n298_, keyIn_0_12, new_n299_ );
nand g197 ( new_n303_, new_n301_, new_n302_ );
xor g198 ( new_n304_, N105, N121 );
xnor g199 ( new_n305_, N73, N89 );
xor g200 ( new_n306_, new_n304_, new_n305_ );
nand g201 ( new_n307_, new_n303_, new_n306_ );
not g202 ( new_n308_, new_n306_ );
nand g203 ( new_n309_, new_n301_, new_n302_, new_n308_ );
nand g204 ( new_n310_, new_n307_, new_n309_ );
nand g205 ( new_n311_, new_n310_, keyIn_0_14 );
not g206 ( new_n312_, keyIn_0_14 );
nand g207 ( new_n313_, new_n307_, new_n312_, new_n309_ );
nand g208 ( new_n314_, new_n311_, new_n313_ );
xor g209 ( new_n315_, new_n149_, new_n227_ );
nand g210 ( new_n316_, N136, N137 );
xnor g211 ( new_n317_, new_n315_, new_n316_ );
xor g212 ( new_n318_, N109, N125 );
xnor g213 ( new_n319_, N77, N93 );
xnor g214 ( new_n320_, new_n318_, new_n319_ );
xnor g215 ( new_n321_, new_n317_, new_n320_ );
and g216 ( new_n322_, new_n314_, new_n287_, new_n321_ );
nand g217 ( new_n323_, new_n200_, new_n322_ );
nand g218 ( new_n324_, new_n323_, keyIn_0_18 );
not g219 ( new_n325_, keyIn_0_18 );
nand g220 ( new_n326_, new_n200_, new_n322_, new_n325_ );
nand g221 ( new_n327_, new_n324_, new_n326_ );
nand g222 ( new_n328_, new_n327_, new_n120_ );
nand g223 ( new_n329_, new_n328_, keyIn_0_20 );
not g224 ( new_n330_, keyIn_0_20 );
nand g225 ( new_n331_, new_n327_, new_n330_, new_n120_ );
nand g226 ( new_n332_, new_n329_, new_n331_ );
nand g227 ( new_n333_, new_n332_, new_n106_ );
nand g228 ( new_n334_, new_n329_, N1, new_n331_ );
nand g229 ( new_n335_, new_n333_, new_n334_ );
nand g230 ( new_n336_, new_n335_, keyIn_0_26 );
not g231 ( new_n337_, keyIn_0_26 );
nand g232 ( new_n338_, new_n333_, new_n337_, new_n334_ );
and g233 ( N724, new_n336_, new_n338_ );
nand g234 ( new_n340_, new_n327_, new_n250_ );
nand g235 ( new_n341_, new_n340_, keyIn_0_21 );
not g236 ( new_n342_, keyIn_0_21 );
nand g237 ( new_n343_, new_n327_, new_n342_, new_n250_ );
nand g238 ( new_n344_, new_n341_, new_n343_ );
nand g239 ( new_n345_, new_n344_, N5 );
nand g240 ( new_n346_, new_n341_, new_n203_, new_n343_ );
nand g241 ( new_n347_, new_n345_, new_n346_ );
nand g242 ( new_n348_, new_n347_, keyIn_0_27 );
not g243 ( new_n349_, keyIn_0_27 );
nand g244 ( new_n350_, new_n345_, new_n349_, new_n346_ );
and g245 ( N725, new_n348_, new_n350_ );
not g246 ( new_n352_, keyIn_0_28 );
nand g247 ( new_n353_, new_n327_, new_n279_ );
nand g248 ( new_n354_, new_n353_, keyIn_0_22 );
not g249 ( new_n355_, keyIn_0_22 );
nand g250 ( new_n356_, new_n327_, new_n355_, new_n279_ );
nand g251 ( new_n357_, new_n354_, new_n356_ );
nand g252 ( new_n358_, new_n357_, new_n212_ );
nand g253 ( new_n359_, new_n354_, N9, new_n356_ );
nand g254 ( new_n360_, new_n358_, new_n359_ );
nand g255 ( new_n361_, new_n360_, new_n352_ );
nand g256 ( new_n362_, new_n358_, keyIn_0_28, new_n359_ );
and g257 ( N726, new_n361_, new_n362_ );
nand g258 ( new_n364_, new_n327_, new_n277_ );
nand g259 ( new_n365_, new_n364_, keyIn_0_23 );
not g260 ( new_n366_, keyIn_0_23 );
nand g261 ( new_n367_, new_n327_, new_n366_, new_n277_ );
nand g262 ( new_n368_, new_n365_, new_n367_ );
nand g263 ( new_n369_, new_n368_, new_n210_ );
nand g264 ( new_n370_, new_n365_, N13, new_n367_ );
nand g265 ( new_n371_, new_n369_, new_n370_ );
nand g266 ( new_n372_, new_n371_, keyIn_0_29 );
not g267 ( new_n373_, keyIn_0_29 );
nand g268 ( new_n374_, new_n369_, new_n373_, new_n370_ );
and g269 ( N727, new_n372_, new_n374_ );
nor g270 ( new_n376_, new_n314_, new_n321_ );
nand g271 ( new_n377_, new_n376_, new_n197_, new_n287_ );
or g272 ( new_n378_, new_n377_, keyIn_0_19 );
nand g273 ( new_n379_, new_n377_, keyIn_0_19 );
nand g274 ( new_n380_, new_n378_, new_n120_, new_n379_ );
xnor g275 ( N728, new_n380_, N17 );
not g276 ( new_n382_, keyIn_0_30 );
not g277 ( new_n383_, N21 );
not g278 ( new_n384_, keyIn_0_24 );
nand g279 ( new_n385_, new_n378_, new_n250_, new_n379_ );
xnor g280 ( new_n386_, new_n385_, new_n384_ );
nand g281 ( new_n387_, new_n386_, new_n383_ );
xnor g282 ( new_n388_, new_n385_, keyIn_0_24 );
nand g283 ( new_n389_, new_n388_, N21 );
nand g284 ( new_n390_, new_n387_, new_n389_ );
nand g285 ( new_n391_, new_n390_, new_n382_ );
nand g286 ( new_n392_, new_n387_, new_n389_, keyIn_0_30 );
nand g287 ( N729, new_n391_, new_n392_ );
nand g288 ( new_n394_, new_n378_, new_n279_, new_n379_ );
xnor g289 ( N730, new_n394_, N25 );
not g290 ( new_n396_, keyIn_0_25 );
nand g291 ( new_n397_, new_n378_, new_n277_, new_n379_ );
xnor g292 ( new_n398_, new_n397_, new_n396_ );
nand g293 ( new_n399_, new_n398_, N29 );
not g294 ( new_n400_, N29 );
xnor g295 ( new_n401_, new_n397_, keyIn_0_25 );
nand g296 ( new_n402_, new_n401_, new_n400_ );
nand g297 ( new_n403_, new_n399_, new_n402_ );
nand g298 ( new_n404_, new_n403_, keyIn_0_31 );
not g299 ( new_n405_, keyIn_0_31 );
nand g300 ( new_n406_, new_n399_, new_n402_, new_n405_ );
nand g301 ( N731, new_n404_, new_n406_ );
and g302 ( new_n408_, new_n314_, new_n321_ );
nor g303 ( new_n409_, new_n197_, new_n234_ );
and g304 ( new_n410_, new_n409_, new_n285_, new_n286_ );
nand g305 ( new_n411_, new_n410_, new_n408_ );
nor g306 ( new_n412_, new_n411_, new_n236_ );
xnor g307 ( N732, new_n412_, new_n153_ );
nor g308 ( new_n414_, new_n411_, new_n261_ );
xnor g309 ( N733, new_n414_, new_n151_ );
nor g310 ( new_n416_, new_n411_, new_n258_ );
xnor g311 ( N734, new_n416_, new_n162_ );
nor g312 ( new_n418_, new_n411_, new_n275_ );
xnor g313 ( N735, new_n418_, new_n160_ );
nand g314 ( new_n420_, new_n410_, new_n376_ );
nor g315 ( new_n421_, new_n420_, new_n236_ );
xnor g316 ( N736, new_n421_, new_n127_ );
nor g317 ( new_n423_, new_n420_, new_n261_ );
xnor g318 ( N737, new_n423_, new_n125_ );
nor g319 ( new_n425_, new_n420_, new_n258_ );
xnor g320 ( N738, new_n425_, new_n137_ );
nor g321 ( new_n427_, new_n420_, new_n275_ );
xnor g322 ( N739, new_n427_, new_n135_ );
nor g323 ( new_n429_, new_n280_, new_n236_, new_n250_ );
nand g324 ( new_n430_, new_n409_, new_n311_, new_n313_ );
or g325 ( new_n431_, new_n314_, keyIn_0_16 );
nand g326 ( new_n432_, new_n314_, keyIn_0_16 );
and g327 ( new_n433_, new_n197_, new_n234_ );
nand g328 ( new_n434_, new_n431_, new_n433_, new_n432_ );
nand g329 ( new_n435_, new_n434_, new_n430_ );
nand g330 ( new_n436_, new_n435_, new_n321_ );
not g331 ( new_n437_, new_n197_ );
nor g332 ( new_n438_, new_n408_, new_n376_ );
or g333 ( new_n439_, new_n438_, new_n437_, new_n234_ );
nand g334 ( new_n440_, new_n439_, new_n436_ );
nand g335 ( new_n441_, new_n440_, new_n234_, new_n429_ );
xnor g336 ( N740, new_n441_, N65 );
nand g337 ( new_n443_, new_n440_, new_n437_, new_n429_ );
xnor g338 ( N741, new_n443_, N69 );
nand g339 ( new_n445_, new_n440_, new_n314_, new_n429_ );
xnor g340 ( N742, new_n445_, N73 );
nor g341 ( new_n448_, new_n437_, new_n314_, new_n234_, new_n321_ );
nand g342 ( new_n449_, new_n448_, new_n429_ );
xnor g343 ( N743, new_n449_, N77 );
nor g344 ( new_n451_, new_n262_, new_n275_ );
nand g345 ( new_n452_, new_n440_, new_n234_, new_n451_ );
xnor g346 ( N744, new_n452_, N81 );
nand g347 ( new_n454_, new_n440_, new_n437_, new_n451_ );
xnor g348 ( N745, new_n454_, N85 );
nand g349 ( new_n456_, new_n440_, new_n314_, new_n451_ );
xnor g350 ( N746, new_n456_, N89 );
nand g351 ( new_n458_, new_n448_, new_n451_ );
xnor g352 ( N747, new_n458_, N93 );
nor g353 ( new_n460_, new_n280_, new_n120_, new_n261_ );
nand g354 ( new_n461_, new_n440_, new_n234_, new_n460_ );
xnor g355 ( N748, new_n461_, N97 );
nand g356 ( new_n463_, new_n440_, new_n437_, new_n460_ );
xnor g357 ( N749, new_n463_, N101 );
nand g358 ( new_n465_, new_n440_, new_n314_, new_n460_ );
xnor g359 ( N750, new_n465_, N105 );
nand g360 ( new_n467_, new_n448_, new_n460_ );
xnor g361 ( N751, new_n467_, N109 );
nor g362 ( new_n469_, new_n259_, new_n275_ );
nand g363 ( new_n470_, new_n440_, new_n234_, new_n469_ );
xnor g364 ( N752, new_n470_, N113 );
nand g365 ( new_n472_, new_n440_, new_n437_, new_n469_ );
xnor g366 ( N753, new_n472_, N117 );
nand g367 ( new_n474_, new_n440_, new_n314_, new_n469_ );
xnor g368 ( N754, new_n474_, N121 );
nand g369 ( new_n476_, new_n448_, new_n469_ );
xnor g370 ( N755, new_n476_, N125 );
endmodule