module add_mul_sub_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        operation_0_, operation_1_, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, operation_0_,
         operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521;

  OR2_X1 U264 ( .A1(n256), .A2(n257), .ZN(Result_7_) );
  AND2_X1 U265 ( .A1(n258), .A2(n259), .ZN(n257) );
  OR2_X1 U266 ( .A1(n260), .A2(n261), .ZN(n258) );
  AND2_X1 U267 ( .A1(n262), .A2(n263), .ZN(n256) );
  OR2_X1 U268 ( .A1(n264), .A2(n265), .ZN(Result_6_) );
  OR2_X1 U269 ( .A1(n266), .A2(n267), .ZN(n265) );
  AND2_X1 U270 ( .A1(n268), .A2(n269), .ZN(n267) );
  OR2_X1 U271 ( .A1(n270), .A2(n271), .ZN(n268) );
  AND2_X1 U272 ( .A1(a_2_), .A2(n272), .ZN(n271) );
  OR2_X1 U273 ( .A1(n273), .A2(n274), .ZN(n272) );
  AND2_X1 U274 ( .A1(n262), .A2(b_3_), .ZN(n273) );
  AND2_X1 U275 ( .A1(n275), .A2(n276), .ZN(n270) );
  AND2_X1 U276 ( .A1(b_2_), .A2(n277), .ZN(n266) );
  OR2_X1 U277 ( .A1(n278), .A2(n279), .ZN(n277) );
  OR2_X1 U278 ( .A1(n280), .A2(n281), .ZN(n279) );
  AND2_X1 U279 ( .A1(n282), .A2(n276), .ZN(n281) );
  OR2_X1 U280 ( .A1(n283), .A2(n274), .ZN(n282) );
  OR2_X1 U281 ( .A1(n284), .A2(n285), .ZN(n274) );
  OR2_X1 U282 ( .A1(n286), .A2(n287), .ZN(n285) );
  AND2_X1 U283 ( .A1(n288), .A2(n289), .ZN(n287) );
  AND2_X1 U284 ( .A1(n290), .A2(n291), .ZN(n286) );
  AND2_X1 U285 ( .A1(n292), .A2(n293), .ZN(n284) );
  AND2_X1 U286 ( .A1(n262), .A2(a_3_), .ZN(n283) );
  AND2_X1 U287 ( .A1(a_2_), .A2(n275), .ZN(n280) );
  OR2_X1 U288 ( .A1(n294), .A2(n295), .ZN(n275) );
  OR2_X1 U289 ( .A1(n296), .A2(n297), .ZN(n295) );
  AND2_X1 U290 ( .A1(n260), .A2(n288), .ZN(n297) );
  AND2_X1 U291 ( .A1(n290), .A2(n263), .ZN(n296) );
  AND2_X1 U292 ( .A1(n292), .A2(n261), .ZN(n294) );
  AND2_X1 U293 ( .A1(n260), .A2(n262), .ZN(n278) );
  AND2_X1 U294 ( .A1(n298), .A2(a_2_), .ZN(n264) );
  AND2_X1 U295 ( .A1(n261), .A2(n262), .ZN(n298) );
  OR2_X1 U296 ( .A1(n299), .A2(n300), .ZN(Result_5_) );
  OR2_X1 U297 ( .A1(n301), .A2(n302), .ZN(n300) );
  AND2_X1 U298 ( .A1(n303), .A2(n304), .ZN(n302) );
  OR2_X1 U299 ( .A1(n305), .A2(n306), .ZN(n304) );
  OR2_X1 U300 ( .A1(n307), .A2(n308), .ZN(n306) );
  AND2_X1 U301 ( .A1(n288), .A2(n309), .ZN(n308) );
  AND2_X1 U302 ( .A1(n290), .A2(n310), .ZN(n307) );
  AND2_X1 U303 ( .A1(n292), .A2(n311), .ZN(n305) );
  INV_X1 U304 ( .A(n312), .ZN(n303) );
  AND2_X1 U305 ( .A1(n312), .A2(n313), .ZN(n301) );
  OR2_X1 U306 ( .A1(n314), .A2(n315), .ZN(n313) );
  OR2_X1 U307 ( .A1(n316), .A2(n317), .ZN(n315) );
  AND2_X1 U308 ( .A1(n318), .A2(n288), .ZN(n317) );
  INV_X1 U309 ( .A(n309), .ZN(n318) );
  AND2_X1 U310 ( .A1(n319), .A2(n290), .ZN(n316) );
  INV_X1 U311 ( .A(n310), .ZN(n319) );
  AND2_X1 U312 ( .A1(n320), .A2(n292), .ZN(n314) );
  INV_X1 U313 ( .A(n311), .ZN(n320) );
  OR2_X1 U314 ( .A1(n321), .A2(n322), .ZN(n312) );
  AND2_X1 U315 ( .A1(a_1_), .A2(n323), .ZN(n322) );
  AND2_X1 U316 ( .A1(b_1_), .A2(n324), .ZN(n321) );
  AND2_X1 U317 ( .A1(n262), .A2(n325), .ZN(n299) );
  OR2_X1 U318 ( .A1(n326), .A2(n327), .ZN(n325) );
  AND2_X1 U319 ( .A1(n328), .A2(n329), .ZN(n327) );
  INV_X1 U320 ( .A(n330), .ZN(n326) );
  OR2_X1 U321 ( .A1(n329), .A2(n328), .ZN(n330) );
  OR2_X1 U322 ( .A1(n331), .A2(n332), .ZN(n328) );
  AND2_X1 U323 ( .A1(n333), .A2(n334), .ZN(n332) );
  AND2_X1 U324 ( .A1(n335), .A2(n336), .ZN(n331) );
  OR2_X1 U325 ( .A1(n337), .A2(n338), .ZN(Result_4_) );
  OR2_X1 U326 ( .A1(n339), .A2(n340), .ZN(n338) );
  AND2_X1 U327 ( .A1(n341), .A2(n342), .ZN(n340) );
  OR2_X1 U328 ( .A1(n343), .A2(n344), .ZN(n341) );
  OR2_X1 U329 ( .A1(n345), .A2(n346), .ZN(n344) );
  AND2_X1 U330 ( .A1(n347), .A2(n288), .ZN(n346) );
  INV_X1 U331 ( .A(n348), .ZN(n347) );
  AND2_X1 U332 ( .A1(n349), .A2(n290), .ZN(n345) );
  INV_X1 U333 ( .A(n350), .ZN(n349) );
  AND2_X1 U334 ( .A1(n351), .A2(n292), .ZN(n343) );
  INV_X1 U335 ( .A(n352), .ZN(n351) );
  AND2_X1 U336 ( .A1(n353), .A2(n354), .ZN(n339) );
  OR2_X1 U337 ( .A1(n355), .A2(n356), .ZN(n354) );
  OR2_X1 U338 ( .A1(n357), .A2(n358), .ZN(n356) );
  AND2_X1 U339 ( .A1(n288), .A2(n348), .ZN(n358) );
  AND2_X1 U340 ( .A1(n290), .A2(n350), .ZN(n357) );
  OR2_X1 U341 ( .A1(n359), .A2(n360), .ZN(n350) );
  AND2_X1 U342 ( .A1(a_1_), .A2(n310), .ZN(n360) );
  AND2_X1 U343 ( .A1(b_1_), .A2(n361), .ZN(n359) );
  OR2_X1 U344 ( .A1(a_1_), .A2(n310), .ZN(n361) );
  OR2_X1 U345 ( .A1(n362), .A2(n363), .ZN(n310) );
  AND2_X1 U346 ( .A1(n263), .A2(n364), .ZN(n362) );
  OR2_X1 U347 ( .A1(a_2_), .A2(b_2_), .ZN(n364) );
  AND2_X1 U348 ( .A1(n365), .A2(n366), .ZN(n290) );
  AND2_X1 U349 ( .A1(n292), .A2(n352), .ZN(n355) );
  INV_X1 U350 ( .A(n342), .ZN(n353) );
  OR2_X1 U351 ( .A1(n367), .A2(n368), .ZN(n342) );
  AND2_X1 U352 ( .A1(n369), .A2(n262), .ZN(n337) );
  AND2_X1 U353 ( .A1(n370), .A2(n371), .ZN(n369) );
  INV_X1 U354 ( .A(n372), .ZN(n371) );
  AND2_X1 U355 ( .A1(n373), .A2(n374), .ZN(n372) );
  OR2_X1 U356 ( .A1(n374), .A2(n373), .ZN(n370) );
  AND2_X1 U357 ( .A1(n375), .A2(n376), .ZN(n373) );
  OR2_X1 U358 ( .A1(n377), .A2(n378), .ZN(n376) );
  INV_X1 U359 ( .A(n379), .ZN(n378) );
  OR2_X1 U360 ( .A1(n379), .A2(n380), .ZN(n375) );
  INV_X1 U361 ( .A(n377), .ZN(n380) );
  OR2_X1 U362 ( .A1(n381), .A2(n382), .ZN(Result_3_) );
  AND2_X1 U363 ( .A1(n383), .A2(n262), .ZN(n381) );
  AND2_X1 U364 ( .A1(n384), .A2(n385), .ZN(n383) );
  OR2_X1 U365 ( .A1(n386), .A2(n387), .ZN(n384) );
  OR2_X1 U366 ( .A1(n388), .A2(n382), .ZN(Result_2_) );
  AND2_X1 U367 ( .A1(n389), .A2(n262), .ZN(n388) );
  AND2_X1 U368 ( .A1(n390), .A2(n391), .ZN(n389) );
  OR2_X1 U369 ( .A1(n392), .A2(n393), .ZN(n390) );
  AND2_X1 U370 ( .A1(n394), .A2(n395), .ZN(n393) );
  OR2_X1 U371 ( .A1(n396), .A2(n397), .ZN(n394) );
  AND2_X1 U372 ( .A1(n386), .A2(n387), .ZN(n392) );
  INV_X1 U373 ( .A(n398), .ZN(n387) );
  INV_X1 U374 ( .A(n399), .ZN(n386) );
  OR2_X1 U375 ( .A1(n400), .A2(n382), .ZN(Result_1_) );
  AND2_X1 U376 ( .A1(n262), .A2(n401), .ZN(n400) );
  OR2_X1 U377 ( .A1(n402), .A2(n403), .ZN(n401) );
  AND2_X1 U378 ( .A1(n404), .A2(n391), .ZN(n403) );
  AND2_X1 U379 ( .A1(n405), .A2(n406), .ZN(n402) );
  OR2_X1 U380 ( .A1(n407), .A2(n382), .ZN(Result_0_) );
  OR2_X1 U381 ( .A1(n408), .A2(n409), .ZN(n382) );
  AND2_X1 U382 ( .A1(n292), .A2(n410), .ZN(n409) );
  OR2_X1 U383 ( .A1(n411), .A2(n367), .ZN(n410) );
  INV_X1 U384 ( .A(n412), .ZN(n367) );
  AND2_X1 U385 ( .A1(n352), .A2(n413), .ZN(n411) );
  OR2_X1 U386 ( .A1(n414), .A2(n415), .ZN(n352) );
  AND2_X1 U387 ( .A1(n311), .A2(n324), .ZN(n415) );
  AND2_X1 U388 ( .A1(b_1_), .A2(n416), .ZN(n414) );
  OR2_X1 U389 ( .A1(n324), .A2(n311), .ZN(n416) );
  OR2_X1 U390 ( .A1(n417), .A2(n418), .ZN(n311) );
  AND2_X1 U391 ( .A1(n261), .A2(n276), .ZN(n418) );
  AND2_X1 U392 ( .A1(b_2_), .A2(n419), .ZN(n417) );
  OR2_X1 U393 ( .A1(n261), .A2(n276), .ZN(n419) );
  INV_X1 U394 ( .A(n293), .ZN(n261) );
  OR2_X1 U395 ( .A1(a_3_), .A2(n420), .ZN(n293) );
  AND2_X1 U396 ( .A1(n366), .A2(operation_1_), .ZN(n292) );
  AND2_X1 U397 ( .A1(n421), .A2(n288), .ZN(n408) );
  AND2_X1 U398 ( .A1(n365), .A2(operation_0_), .ZN(n288) );
  AND2_X1 U399 ( .A1(n422), .A2(n412), .ZN(n421) );
  OR2_X1 U400 ( .A1(a_0_), .A2(n423), .ZN(n412) );
  OR2_X1 U401 ( .A1(n368), .A2(n348), .ZN(n422) );
  OR2_X1 U402 ( .A1(n424), .A2(n425), .ZN(n348) );
  AND2_X1 U403 ( .A1(a_1_), .A2(n309), .ZN(n425) );
  AND2_X1 U404 ( .A1(n426), .A2(n323), .ZN(n424) );
  OR2_X1 U405 ( .A1(a_1_), .A2(n309), .ZN(n426) );
  OR2_X1 U406 ( .A1(n427), .A2(n428), .ZN(n309) );
  AND2_X1 U407 ( .A1(n260), .A2(a_2_), .ZN(n428) );
  AND2_X1 U408 ( .A1(n429), .A2(n269), .ZN(n427) );
  OR2_X1 U409 ( .A1(n260), .A2(a_2_), .ZN(n429) );
  INV_X1 U410 ( .A(n289), .ZN(n260) );
  OR2_X1 U411 ( .A1(b_3_), .A2(n430), .ZN(n289) );
  INV_X1 U412 ( .A(n413), .ZN(n368) );
  OR2_X1 U413 ( .A1(b_0_), .A2(n431), .ZN(n413) );
  AND2_X1 U414 ( .A1(n262), .A2(n432), .ZN(n407) );
  OR2_X1 U415 ( .A1(n433), .A2(n434), .ZN(n432) );
  OR2_X1 U416 ( .A1(n435), .A2(n436), .ZN(n434) );
  AND2_X1 U417 ( .A1(n404), .A2(n405), .ZN(n436) );
  INV_X1 U418 ( .A(n391), .ZN(n405) );
  OR2_X1 U419 ( .A1(n437), .A2(n385), .ZN(n391) );
  OR2_X1 U420 ( .A1(n399), .A2(n398), .ZN(n385) );
  OR2_X1 U421 ( .A1(n438), .A2(n439), .ZN(n398) );
  INV_X1 U422 ( .A(n440), .ZN(n439) );
  OR2_X1 U423 ( .A1(n441), .A2(n442), .ZN(n440) );
  AND2_X1 U424 ( .A1(n442), .A2(n441), .ZN(n438) );
  AND2_X1 U425 ( .A1(n443), .A2(n444), .ZN(n441) );
  OR2_X1 U426 ( .A1(n445), .A2(n446), .ZN(n444) );
  INV_X1 U427 ( .A(n447), .ZN(n446) );
  OR2_X1 U428 ( .A1(n447), .A2(n448), .ZN(n443) );
  INV_X1 U429 ( .A(n445), .ZN(n448) );
  OR2_X1 U430 ( .A1(n449), .A2(n450), .ZN(n399) );
  AND2_X1 U431 ( .A1(n377), .A2(n379), .ZN(n450) );
  AND2_X1 U432 ( .A1(n374), .A2(n451), .ZN(n449) );
  OR2_X1 U433 ( .A1(n379), .A2(n377), .ZN(n451) );
  OR2_X1 U434 ( .A1(n420), .A2(n431), .ZN(n377) );
  OR2_X1 U435 ( .A1(n452), .A2(n453), .ZN(n379) );
  AND2_X1 U436 ( .A1(n336), .A2(n334), .ZN(n453) );
  AND2_X1 U437 ( .A1(n329), .A2(n454), .ZN(n452) );
  OR2_X1 U438 ( .A1(n334), .A2(n336), .ZN(n454) );
  INV_X1 U439 ( .A(n333), .ZN(n336) );
  AND2_X1 U440 ( .A1(b_3_), .A2(a_1_), .ZN(n333) );
  INV_X1 U441 ( .A(n335), .ZN(n334) );
  AND2_X1 U442 ( .A1(n263), .A2(n363), .ZN(n335) );
  INV_X1 U443 ( .A(n291), .ZN(n263) );
  OR2_X1 U444 ( .A1(n430), .A2(n420), .ZN(n291) );
  INV_X1 U445 ( .A(b_3_), .ZN(n420) );
  AND2_X1 U446 ( .A1(n455), .A2(n456), .ZN(n329) );
  OR2_X1 U447 ( .A1(n457), .A2(n363), .ZN(n456) );
  INV_X1 U448 ( .A(n458), .ZN(n363) );
  OR2_X1 U449 ( .A1(n458), .A2(n459), .ZN(n455) );
  OR2_X1 U450 ( .A1(n460), .A2(n461), .ZN(n374) );
  AND2_X1 U451 ( .A1(n462), .A2(n463), .ZN(n461) );
  INV_X1 U452 ( .A(n464), .ZN(n460) );
  OR2_X1 U453 ( .A1(n462), .A2(n463), .ZN(n464) );
  OR2_X1 U454 ( .A1(n465), .A2(n466), .ZN(n462) );
  INV_X1 U455 ( .A(n467), .ZN(n466) );
  OR2_X1 U456 ( .A1(n468), .A2(n469), .ZN(n467) );
  AND2_X1 U457 ( .A1(n469), .A2(n468), .ZN(n465) );
  OR2_X1 U458 ( .A1(n470), .A2(n471), .ZN(n437) );
  AND2_X1 U459 ( .A1(n472), .A2(n473), .ZN(n471) );
  AND2_X1 U460 ( .A1(n397), .A2(n396), .ZN(n470) );
  INV_X1 U461 ( .A(n473), .ZN(n396) );
  INV_X1 U462 ( .A(n472), .ZN(n397) );
  INV_X1 U463 ( .A(n406), .ZN(n404) );
  OR2_X1 U464 ( .A1(n474), .A2(n435), .ZN(n406) );
  AND2_X1 U465 ( .A1(n475), .A2(n395), .ZN(n474) );
  INV_X1 U466 ( .A(n476), .ZN(n435) );
  OR2_X1 U467 ( .A1(n475), .A2(n395), .ZN(n476) );
  OR2_X1 U468 ( .A1(n473), .A2(n472), .ZN(n395) );
  OR2_X1 U469 ( .A1(n477), .A2(n478), .ZN(n472) );
  AND2_X1 U470 ( .A1(n479), .A2(n480), .ZN(n478) );
  INV_X1 U471 ( .A(n481), .ZN(n477) );
  OR2_X1 U472 ( .A1(n479), .A2(n480), .ZN(n481) );
  OR2_X1 U473 ( .A1(n482), .A2(n483), .ZN(n479) );
  AND2_X1 U474 ( .A1(n484), .A2(n485), .ZN(n483) );
  AND2_X1 U475 ( .A1(n486), .A2(n487), .ZN(n482) );
  OR2_X1 U476 ( .A1(n488), .A2(n489), .ZN(n473) );
  AND2_X1 U477 ( .A1(n445), .A2(n447), .ZN(n489) );
  AND2_X1 U478 ( .A1(n442), .A2(n490), .ZN(n488) );
  OR2_X1 U479 ( .A1(n447), .A2(n445), .ZN(n490) );
  OR2_X1 U480 ( .A1(n491), .A2(n492), .ZN(n445) );
  AND2_X1 U481 ( .A1(n463), .A2(n468), .ZN(n492) );
  AND2_X1 U482 ( .A1(n469), .A2(n493), .ZN(n491) );
  OR2_X1 U483 ( .A1(n468), .A2(n463), .ZN(n493) );
  OR2_X1 U484 ( .A1(n269), .A2(n324), .ZN(n463) );
  OR2_X1 U485 ( .A1(n458), .A2(n457), .ZN(n468) );
  INV_X1 U486 ( .A(n459), .ZN(n457) );
  OR2_X1 U487 ( .A1(n276), .A2(n269), .ZN(n458) );
  INV_X1 U488 ( .A(n494), .ZN(n469) );
  OR2_X1 U489 ( .A1(n495), .A2(n496), .ZN(n494) );
  AND2_X1 U490 ( .A1(n497), .A2(b_1_), .ZN(n496) );
  AND2_X1 U491 ( .A1(a_2_), .A2(n498), .ZN(n497) );
  OR2_X1 U492 ( .A1(n430), .A2(n423), .ZN(n498) );
  INV_X1 U493 ( .A(a_3_), .ZN(n430) );
  AND2_X1 U494 ( .A1(n499), .A2(b_0_), .ZN(n495) );
  AND2_X1 U495 ( .A1(a_3_), .A2(n500), .ZN(n499) );
  OR2_X1 U496 ( .A1(n276), .A2(n323), .ZN(n500) );
  OR2_X1 U497 ( .A1(n269), .A2(n431), .ZN(n447) );
  INV_X1 U498 ( .A(b_2_), .ZN(n269) );
  OR2_X1 U499 ( .A1(n501), .A2(n502), .ZN(n442) );
  INV_X1 U500 ( .A(n503), .ZN(n502) );
  OR2_X1 U501 ( .A1(n504), .A2(n505), .ZN(n503) );
  AND2_X1 U502 ( .A1(n505), .A2(n504), .ZN(n501) );
  OR2_X1 U503 ( .A1(n506), .A2(n507), .ZN(n504) );
  AND2_X1 U504 ( .A1(n508), .A2(b_0_), .ZN(n507) );
  AND2_X1 U505 ( .A1(a_2_), .A2(n509), .ZN(n508) );
  OR2_X1 U506 ( .A1(n323), .A2(n324), .ZN(n509) );
  AND2_X1 U507 ( .A1(n510), .A2(a_1_), .ZN(n506) );
  AND2_X1 U508 ( .A1(b_1_), .A2(n511), .ZN(n510) );
  OR2_X1 U509 ( .A1(n276), .A2(n423), .ZN(n511) );
  INV_X1 U510 ( .A(a_2_), .ZN(n276) );
  OR2_X1 U511 ( .A1(n433), .A2(n512), .ZN(n475) );
  AND2_X1 U512 ( .A1(n513), .A2(n514), .ZN(n512) );
  OR2_X1 U513 ( .A1(n423), .A2(n431), .ZN(n513) );
  AND2_X1 U514 ( .A1(n515), .A2(a_0_), .ZN(n433) );
  INV_X1 U515 ( .A(n514), .ZN(n515) );
  OR2_X1 U516 ( .A1(n516), .A2(n517), .ZN(n514) );
  AND2_X1 U517 ( .A1(n480), .A2(n485), .ZN(n517) );
  AND2_X1 U518 ( .A1(n484), .A2(n518), .ZN(n516) );
  OR2_X1 U519 ( .A1(n485), .A2(n480), .ZN(n518) );
  OR2_X1 U520 ( .A1(n323), .A2(n431), .ZN(n480) );
  INV_X1 U521 ( .A(a_0_), .ZN(n431) );
  INV_X1 U522 ( .A(b_1_), .ZN(n323) );
  INV_X1 U523 ( .A(n487), .ZN(n484) );
  OR2_X1 U524 ( .A1(n519), .A2(n505), .ZN(n487) );
  AND2_X1 U525 ( .A1(b_0_), .A2(n520), .ZN(n505) );
  AND2_X1 U526 ( .A1(a_2_), .A2(n459), .ZN(n520) );
  AND2_X1 U527 ( .A1(a_3_), .A2(b_1_), .ZN(n459) );
  AND2_X1 U528 ( .A1(n521), .A2(n486), .ZN(n519) );
  INV_X1 U529 ( .A(n485), .ZN(n486) );
  OR2_X1 U530 ( .A1(n324), .A2(n423), .ZN(n485) );
  INV_X1 U531 ( .A(b_0_), .ZN(n423) );
  INV_X1 U532 ( .A(a_1_), .ZN(n324) );
  AND2_X1 U533 ( .A1(b_1_), .A2(a_2_), .ZN(n521) );
  INV_X1 U534 ( .A(n259), .ZN(n262) );
  OR2_X1 U535 ( .A1(n366), .A2(n365), .ZN(n259) );
  INV_X1 U536 ( .A(operation_1_), .ZN(n365) );
  INV_X1 U537 ( .A(operation_0_), .ZN(n366) );
endmodule

