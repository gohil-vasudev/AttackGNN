module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n300_, new_n302_, new_n303_, new_n305_, new_n306_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n321_, new_n323_, new_n324_, new_n326_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n336_, new_n338_, new_n340_, new_n341_, new_n343_, new_n344_, new_n346_, new_n348_, new_n350_, new_n351_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n388_, new_n389_, new_n391_, new_n392_, new_n394_, new_n395_, new_n397_, new_n398_, new_n400_, new_n401_, new_n402_, new_n404_, new_n406_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_, new_n423_, new_n425_, new_n427_, new_n428_, new_n430_, new_n431_, new_n432_, new_n433_, new_n435_, new_n436_, new_n438_, new_n440_, new_n441_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XOR2_X1 g004 ( .A(G57GAT), .B(KEYINPUT1), .Z(new_n142_) );
  AND2_X1 g005 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n142_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(new_n144_), .B(new_n141_), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(G120GAT), .B(G127GAT), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n148_), .B(new_n138_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n145_), .B(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .ZN(new_n151_) );
  XNOR2_X1 g014 ( .A(new_n150_), .B(new_n151_), .ZN(new_n152_) );
  XNOR2_X1 g015 ( .A(G85GAT), .B(G162GAT), .ZN(new_n153_) );
  XNOR2_X1 g016 ( .A(new_n152_), .B(new_n153_), .ZN(new_n154_) );
  XNOR2_X1 g017 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(new_n155_) );
  XNOR2_X1 g018 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n156_) );
  XNOR2_X1 g019 ( .A(new_n155_), .B(new_n156_), .ZN(new_n157_) );
  XOR2_X1 g020 ( .A(new_n154_), .B(new_n157_), .Z(new_n158_) );
  INV_X1 g021 ( .A(new_n158_), .ZN(new_n159_) );
  INV_X1 g022 ( .A(G197GAT), .ZN(new_n160_) );
  XNOR2_X1 g023 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(G211GAT), .B(G218GAT), .ZN(new_n162_) );
  XNOR2_X1 g025 ( .A(new_n161_), .B(new_n162_), .ZN(new_n163_) );
  XNOR2_X1 g026 ( .A(new_n163_), .B(new_n160_), .ZN(new_n164_) );
  XNOR2_X1 g027 ( .A(new_n164_), .B(new_n141_), .ZN(new_n165_) );
  XOR2_X1 g028 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n166_) );
  XNOR2_X1 g029 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n167_) );
  XNOR2_X1 g030 ( .A(new_n166_), .B(new_n167_), .ZN(new_n168_) );
  XNOR2_X1 g031 ( .A(G78GAT), .B(G106GAT), .ZN(new_n169_) );
  AND2_X1 g032 ( .A1(new_n169_), .A2(G148GAT), .ZN(new_n170_) );
  INV_X1 g033 ( .A(G148GAT), .ZN(new_n171_) );
  AND2_X1 g034 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n172_) );
  INV_X1 g035 ( .A(new_n172_), .ZN(new_n173_) );
  OR2_X1 g036 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n174_) );
  AND3_X1 g037 ( .A1(new_n173_), .A2(new_n171_), .A3(new_n174_), .ZN(new_n175_) );
  OR2_X1 g038 ( .A1(new_n170_), .A2(new_n175_), .ZN(new_n176_) );
  XNOR2_X1 g039 ( .A(new_n176_), .B(new_n168_), .ZN(new_n177_) );
  XNOR2_X1 g040 ( .A(new_n165_), .B(new_n177_), .ZN(new_n178_) );
  XNOR2_X1 g041 ( .A(G50GAT), .B(G162GAT), .ZN(new_n179_) );
  XNOR2_X1 g042 ( .A(new_n178_), .B(new_n179_), .ZN(new_n180_) );
  AND2_X1 g043 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n181_) );
  XOR2_X1 g044 ( .A(new_n180_), .B(new_n181_), .Z(new_n182_) );
  XOR2_X1 g045 ( .A(new_n148_), .B(G15GAT), .Z(new_n183_) );
  AND2_X1 g046 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n184_) );
  XOR2_X1 g047 ( .A(new_n183_), .B(new_n184_), .Z(new_n185_) );
  XNOR2_X1 g048 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n186_) );
  XNOR2_X1 g049 ( .A(G176GAT), .B(G183GAT), .ZN(new_n187_) );
  XNOR2_X1 g050 ( .A(new_n186_), .B(new_n187_), .ZN(new_n188_) );
  XNOR2_X1 g051 ( .A(new_n185_), .B(new_n188_), .ZN(new_n189_) );
  XNOR2_X1 g052 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n190_) );
  XNOR2_X1 g053 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n191_) );
  XNOR2_X1 g054 ( .A(new_n190_), .B(new_n191_), .ZN(new_n192_) );
  XOR2_X1 g055 ( .A(G134GAT), .B(G190GAT), .Z(new_n193_) );
  XNOR2_X1 g056 ( .A(G43GAT), .B(G99GAT), .ZN(new_n194_) );
  XNOR2_X1 g057 ( .A(new_n193_), .B(new_n194_), .ZN(new_n195_) );
  XNOR2_X1 g058 ( .A(new_n195_), .B(new_n192_), .ZN(new_n196_) );
  XNOR2_X1 g059 ( .A(new_n189_), .B(new_n196_), .ZN(new_n197_) );
  AND2_X1 g060 ( .A1(new_n182_), .A2(new_n197_), .ZN(new_n198_) );
  XNOR2_X1 g061 ( .A(new_n198_), .B(KEYINPUT26), .ZN(new_n199_) );
  XOR2_X1 g062 ( .A(G36GAT), .B(G190GAT), .Z(new_n200_) );
  INV_X1 g063 ( .A(new_n200_), .ZN(new_n201_) );
  XNOR2_X1 g064 ( .A(new_n164_), .B(new_n201_), .ZN(new_n202_) );
  XNOR2_X1 g065 ( .A(G64GAT), .B(G176GAT), .ZN(new_n203_) );
  XNOR2_X1 g066 ( .A(new_n203_), .B(G92GAT), .ZN(new_n204_) );
  AND2_X1 g067 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n205_) );
  XNOR2_X1 g068 ( .A(new_n204_), .B(new_n205_), .ZN(new_n206_) );
  XNOR2_X1 g069 ( .A(G8GAT), .B(G183GAT), .ZN(new_n207_) );
  XNOR2_X1 g070 ( .A(new_n206_), .B(new_n207_), .ZN(new_n208_) );
  XNOR2_X1 g071 ( .A(new_n202_), .B(new_n208_), .ZN(new_n209_) );
  XOR2_X1 g072 ( .A(new_n209_), .B(new_n192_), .Z(new_n210_) );
  XOR2_X1 g073 ( .A(new_n210_), .B(KEYINPUT27), .Z(new_n211_) );
  AND2_X1 g074 ( .A1(new_n199_), .A2(new_n211_), .ZN(new_n212_) );
  INV_X1 g075 ( .A(new_n197_), .ZN(new_n213_) );
  INV_X1 g076 ( .A(new_n210_), .ZN(new_n214_) );
  AND2_X1 g077 ( .A1(new_n213_), .A2(new_n214_), .ZN(new_n215_) );
  OR2_X1 g078 ( .A1(new_n215_), .A2(new_n182_), .ZN(new_n216_) );
  XNOR2_X1 g079 ( .A(new_n216_), .B(KEYINPUT25), .ZN(new_n217_) );
  OR2_X1 g080 ( .A1(new_n212_), .A2(new_n217_), .ZN(new_n218_) );
  AND2_X1 g081 ( .A1(new_n218_), .A2(new_n159_), .ZN(new_n219_) );
  XOR2_X1 g082 ( .A(new_n182_), .B(KEYINPUT28), .Z(new_n220_) );
  AND2_X1 g083 ( .A1(new_n211_), .A2(new_n158_), .ZN(new_n221_) );
  AND3_X1 g084 ( .A1(new_n220_), .A2(new_n221_), .A3(new_n197_), .ZN(new_n222_) );
  OR2_X1 g085 ( .A1(new_n219_), .A2(new_n222_), .ZN(new_n223_) );
  INV_X1 g086 ( .A(KEYINPUT7), .ZN(new_n224_) );
  AND2_X1 g087 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n225_) );
  INV_X1 g088 ( .A(new_n225_), .ZN(new_n226_) );
  OR2_X1 g089 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n227_) );
  AND3_X1 g090 ( .A1(new_n226_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_) );
  XNOR2_X1 g091 ( .A(G43GAT), .B(KEYINPUT8), .ZN(new_n229_) );
  AND2_X1 g092 ( .A1(new_n229_), .A2(KEYINPUT7), .ZN(new_n230_) );
  OR2_X1 g093 ( .A1(new_n230_), .A2(new_n228_), .ZN(new_n231_) );
  XNOR2_X1 g094 ( .A(G85GAT), .B(G99GAT), .ZN(new_n232_) );
  AND2_X1 g095 ( .A1(new_n232_), .A2(G92GAT), .ZN(new_n233_) );
  INV_X1 g096 ( .A(G92GAT), .ZN(new_n234_) );
  OR2_X1 g097 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n235_) );
  AND2_X1 g098 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n236_) );
  INV_X1 g099 ( .A(new_n236_), .ZN(new_n237_) );
  AND3_X1 g100 ( .A1(new_n237_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n238_) );
  OR2_X1 g101 ( .A1(new_n233_), .A2(new_n238_), .ZN(new_n239_) );
  XNOR2_X1 g102 ( .A(new_n231_), .B(new_n239_), .ZN(new_n240_) );
  XOR2_X1 g103 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(new_n241_) );
  AND2_X1 g104 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n242_) );
  XNOR2_X1 g105 ( .A(new_n241_), .B(new_n242_), .ZN(new_n243_) );
  XNOR2_X1 g106 ( .A(new_n243_), .B(KEYINPUT9), .ZN(new_n244_) );
  XNOR2_X1 g107 ( .A(new_n240_), .B(new_n244_), .ZN(new_n245_) );
  XOR2_X1 g108 ( .A(G106GAT), .B(G218GAT), .Z(new_n246_) );
  XNOR2_X1 g109 ( .A(new_n246_), .B(new_n151_), .ZN(new_n247_) );
  XNOR2_X1 g110 ( .A(new_n245_), .B(new_n247_), .ZN(new_n248_) );
  XOR2_X1 g111 ( .A(new_n248_), .B(new_n179_), .Z(new_n249_) );
  XNOR2_X1 g112 ( .A(new_n249_), .B(new_n200_), .ZN(new_n250_) );
  XNOR2_X1 g113 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n251_) );
  XNOR2_X1 g114 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n252_) );
  XNOR2_X1 g115 ( .A(new_n251_), .B(new_n252_), .ZN(new_n253_) );
  XNOR2_X1 g116 ( .A(G78GAT), .B(G155GAT), .ZN(new_n254_) );
  XNOR2_X1 g117 ( .A(G127GAT), .B(G211GAT), .ZN(new_n255_) );
  XNOR2_X1 g118 ( .A(new_n254_), .B(new_n255_), .ZN(new_n256_) );
  XNOR2_X1 g119 ( .A(new_n253_), .B(new_n256_), .ZN(new_n257_) );
  XNOR2_X1 g120 ( .A(G57GAT), .B(G71GAT), .ZN(new_n258_) );
  XOR2_X1 g121 ( .A(new_n258_), .B(KEYINPUT13), .Z(new_n259_) );
  XNOR2_X1 g122 ( .A(G15GAT), .B(G22GAT), .ZN(new_n260_) );
  XNOR2_X1 g123 ( .A(new_n260_), .B(new_n138_), .ZN(new_n261_) );
  XNOR2_X1 g124 ( .A(new_n259_), .B(new_n261_), .ZN(new_n262_) );
  XNOR2_X1 g125 ( .A(new_n262_), .B(new_n257_), .ZN(new_n263_) );
  XNOR2_X1 g126 ( .A(new_n263_), .B(new_n207_), .ZN(new_n264_) );
  AND2_X1 g127 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n265_) );
  XNOR2_X1 g128 ( .A(new_n264_), .B(new_n265_), .ZN(new_n266_) );
  AND2_X1 g129 ( .A1(new_n250_), .A2(new_n266_), .ZN(new_n267_) );
  XNOR2_X1 g130 ( .A(new_n267_), .B(KEYINPUT16), .ZN(new_n268_) );
  AND2_X1 g131 ( .A1(new_n223_), .A2(new_n268_), .ZN(new_n269_) );
  INV_X1 g132 ( .A(new_n259_), .ZN(new_n270_) );
  XNOR2_X1 g133 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n271_) );
  AND2_X1 g134 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n272_) );
  XNOR2_X1 g135 ( .A(new_n271_), .B(new_n272_), .ZN(new_n273_) );
  XNOR2_X1 g136 ( .A(new_n273_), .B(KEYINPUT32), .ZN(new_n274_) );
  XNOR2_X1 g137 ( .A(new_n176_), .B(new_n239_), .ZN(new_n275_) );
  XNOR2_X1 g138 ( .A(new_n275_), .B(new_n274_), .ZN(new_n276_) );
  XNOR2_X1 g139 ( .A(new_n276_), .B(new_n203_), .ZN(new_n277_) );
  XOR2_X1 g140 ( .A(G120GAT), .B(G204GAT), .Z(new_n278_) );
  XNOR2_X1 g141 ( .A(new_n277_), .B(new_n278_), .ZN(new_n279_) );
  XNOR2_X1 g142 ( .A(new_n279_), .B(new_n270_), .ZN(new_n280_) );
  INV_X1 g143 ( .A(new_n280_), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n282_) );
  XNOR2_X1 g145 ( .A(G8GAT), .B(G169GAT), .ZN(new_n283_) );
  XNOR2_X1 g146 ( .A(new_n282_), .B(new_n283_), .ZN(new_n284_) );
  XNOR2_X1 g147 ( .A(G113GAT), .B(G197GAT), .ZN(new_n285_) );
  XNOR2_X1 g148 ( .A(G29GAT), .B(G141GAT), .ZN(new_n286_) );
  XNOR2_X1 g149 ( .A(new_n285_), .B(new_n286_), .ZN(new_n287_) );
  XNOR2_X1 g150 ( .A(new_n284_), .B(new_n287_), .ZN(new_n288_) );
  XNOR2_X1 g151 ( .A(new_n231_), .B(new_n261_), .ZN(new_n289_) );
  XOR2_X1 g152 ( .A(new_n289_), .B(new_n288_), .Z(new_n290_) );
  XOR2_X1 g153 ( .A(G36GAT), .B(G50GAT), .Z(new_n291_) );
  AND2_X1 g154 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n292_) );
  XNOR2_X1 g155 ( .A(new_n291_), .B(new_n292_), .ZN(new_n293_) );
  XOR2_X1 g156 ( .A(new_n290_), .B(new_n293_), .Z(new_n294_) );
  AND2_X1 g157 ( .A1(new_n281_), .A2(new_n294_), .ZN(new_n295_) );
  AND2_X1 g158 ( .A1(new_n269_), .A2(new_n295_), .ZN(new_n296_) );
  AND2_X1 g159 ( .A1(new_n296_), .A2(new_n158_), .ZN(new_n297_) );
  XNOR2_X1 g160 ( .A(new_n297_), .B(KEYINPUT34), .ZN(new_n298_) );
  XNOR2_X1 g161 ( .A(new_n298_), .B(new_n138_), .ZN(G1324GAT) );
  AND2_X1 g162 ( .A1(new_n296_), .A2(new_n214_), .ZN(new_n300_) );
  XOR2_X1 g163 ( .A(new_n300_), .B(G8GAT), .Z(G1325GAT) );
  AND2_X1 g164 ( .A1(new_n296_), .A2(new_n213_), .ZN(new_n302_) );
  XNOR2_X1 g165 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n303_) );
  XNOR2_X1 g166 ( .A(new_n302_), .B(new_n303_), .ZN(G1326GAT) );
  INV_X1 g167 ( .A(new_n220_), .ZN(new_n305_) );
  AND2_X1 g168 ( .A1(new_n296_), .A2(new_n305_), .ZN(new_n306_) );
  XOR2_X1 g169 ( .A(new_n306_), .B(G22GAT), .Z(G1327GAT) );
  INV_X1 g170 ( .A(new_n266_), .ZN(new_n308_) );
  OR2_X1 g171 ( .A1(new_n250_), .A2(KEYINPUT36), .ZN(new_n309_) );
  INV_X1 g172 ( .A(KEYINPUT36), .ZN(new_n310_) );
  XNOR2_X1 g173 ( .A(new_n249_), .B(new_n201_), .ZN(new_n311_) );
  OR2_X1 g174 ( .A1(new_n311_), .A2(new_n310_), .ZN(new_n312_) );
  AND2_X1 g175 ( .A1(new_n309_), .A2(new_n312_), .ZN(new_n313_) );
  AND3_X1 g176 ( .A1(new_n223_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_) );
  XOR2_X1 g177 ( .A(new_n314_), .B(KEYINPUT37), .Z(new_n315_) );
  AND2_X1 g178 ( .A1(new_n315_), .A2(new_n295_), .ZN(new_n316_) );
  XNOR2_X1 g179 ( .A(new_n316_), .B(KEYINPUT38), .ZN(new_n317_) );
  AND2_X1 g180 ( .A1(new_n317_), .A2(new_n158_), .ZN(new_n318_) );
  XNOR2_X1 g181 ( .A(G29GAT), .B(KEYINPUT39), .ZN(new_n319_) );
  XNOR2_X1 g182 ( .A(new_n318_), .B(new_n319_), .ZN(G1328GAT) );
  AND2_X1 g183 ( .A1(new_n317_), .A2(new_n214_), .ZN(new_n321_) );
  XOR2_X1 g184 ( .A(new_n321_), .B(G36GAT), .Z(G1329GAT) );
  AND2_X1 g185 ( .A1(new_n317_), .A2(new_n213_), .ZN(new_n323_) );
  XNOR2_X1 g186 ( .A(new_n323_), .B(KEYINPUT40), .ZN(new_n324_) );
  XOR2_X1 g187 ( .A(new_n324_), .B(G43GAT), .Z(G1330GAT) );
  AND2_X1 g188 ( .A1(new_n317_), .A2(new_n305_), .ZN(new_n326_) );
  XOR2_X1 g189 ( .A(new_n326_), .B(G50GAT), .Z(G1331GAT) );
  INV_X1 g190 ( .A(new_n294_), .ZN(new_n328_) );
  XNOR2_X1 g191 ( .A(new_n280_), .B(KEYINPUT41), .ZN(new_n329_) );
  INV_X1 g192 ( .A(new_n329_), .ZN(new_n330_) );
  AND2_X1 g193 ( .A1(new_n330_), .A2(new_n328_), .ZN(new_n331_) );
  AND2_X1 g194 ( .A1(new_n269_), .A2(new_n331_), .ZN(new_n332_) );
  AND2_X1 g195 ( .A1(new_n332_), .A2(new_n158_), .ZN(new_n333_) );
  XOR2_X1 g196 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n334_) );
  XNOR2_X1 g197 ( .A(new_n333_), .B(new_n334_), .ZN(G1332GAT) );
  AND2_X1 g198 ( .A1(new_n332_), .A2(new_n214_), .ZN(new_n336_) );
  XOR2_X1 g199 ( .A(new_n336_), .B(G64GAT), .Z(G1333GAT) );
  AND2_X1 g200 ( .A1(new_n332_), .A2(new_n213_), .ZN(new_n338_) );
  XOR2_X1 g201 ( .A(new_n338_), .B(G71GAT), .Z(G1334GAT) );
  AND2_X1 g202 ( .A1(new_n332_), .A2(new_n305_), .ZN(new_n340_) );
  XNOR2_X1 g203 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n341_) );
  XNOR2_X1 g204 ( .A(new_n340_), .B(new_n341_), .ZN(G1335GAT) );
  AND2_X1 g205 ( .A1(new_n315_), .A2(new_n331_), .ZN(new_n343_) );
  AND2_X1 g206 ( .A1(new_n343_), .A2(new_n158_), .ZN(new_n344_) );
  XOR2_X1 g207 ( .A(new_n344_), .B(G85GAT), .Z(G1336GAT) );
  AND2_X1 g208 ( .A1(new_n343_), .A2(new_n214_), .ZN(new_n346_) );
  XNOR2_X1 g209 ( .A(new_n346_), .B(new_n234_), .ZN(G1337GAT) );
  AND2_X1 g210 ( .A1(new_n343_), .A2(new_n213_), .ZN(new_n348_) );
  XOR2_X1 g211 ( .A(new_n348_), .B(G99GAT), .Z(G1338GAT) );
  AND2_X1 g212 ( .A1(new_n343_), .A2(new_n305_), .ZN(new_n350_) );
  XNOR2_X1 g213 ( .A(new_n350_), .B(KEYINPUT44), .ZN(new_n351_) );
  XOR2_X1 g214 ( .A(new_n351_), .B(G106GAT), .Z(G1339GAT) );
  INV_X1 g215 ( .A(KEYINPUT46), .ZN(new_n353_) );
  OR3_X1 g216 ( .A1(new_n329_), .A2(new_n353_), .A3(new_n328_), .ZN(new_n354_) );
  INV_X1 g217 ( .A(new_n354_), .ZN(new_n355_) );
  INV_X1 g218 ( .A(KEYINPUT41), .ZN(new_n356_) );
  AND2_X1 g219 ( .A1(new_n279_), .A2(new_n259_), .ZN(new_n357_) );
  OR2_X1 g220 ( .A1(new_n277_), .A2(new_n278_), .ZN(new_n358_) );
  INV_X1 g221 ( .A(new_n203_), .ZN(new_n359_) );
  XNOR2_X1 g222 ( .A(new_n276_), .B(new_n359_), .ZN(new_n360_) );
  INV_X1 g223 ( .A(new_n278_), .ZN(new_n361_) );
  OR2_X1 g224 ( .A1(new_n360_), .A2(new_n361_), .ZN(new_n362_) );
  AND3_X1 g225 ( .A1(new_n358_), .A2(new_n362_), .A3(new_n270_), .ZN(new_n363_) );
  OR3_X1 g226 ( .A1(new_n357_), .A2(new_n356_), .A3(new_n363_), .ZN(new_n364_) );
  OR2_X1 g227 ( .A1(new_n280_), .A2(KEYINPUT41), .ZN(new_n365_) );
  AND3_X1 g228 ( .A1(new_n365_), .A2(new_n294_), .A3(new_n364_), .ZN(new_n366_) );
  OR2_X1 g229 ( .A1(new_n366_), .A2(KEYINPUT46), .ZN(new_n367_) );
  INV_X1 g230 ( .A(new_n367_), .ZN(new_n368_) );
  AND2_X1 g231 ( .A1(new_n250_), .A2(new_n308_), .ZN(new_n369_) );
  INV_X1 g232 ( .A(new_n369_), .ZN(new_n370_) );
  OR4_X1 g233 ( .A1(new_n368_), .A2(new_n355_), .A3(KEYINPUT47), .A4(new_n370_), .ZN(new_n371_) );
  INV_X1 g234 ( .A(KEYINPUT47), .ZN(new_n372_) );
  AND3_X1 g235 ( .A1(new_n367_), .A2(new_n354_), .A3(new_n369_), .ZN(new_n373_) );
  OR2_X1 g236 ( .A1(new_n373_), .A2(new_n372_), .ZN(new_n374_) );
  INV_X1 g237 ( .A(KEYINPUT45), .ZN(new_n375_) );
  AND3_X1 g238 ( .A1(new_n309_), .A2(new_n312_), .A3(new_n266_), .ZN(new_n376_) );
  XNOR2_X1 g239 ( .A(new_n376_), .B(new_n375_), .ZN(new_n377_) );
  OR2_X1 g240 ( .A1(new_n280_), .A2(new_n294_), .ZN(new_n378_) );
  OR2_X1 g241 ( .A1(new_n377_), .A2(new_n378_), .ZN(new_n379_) );
  AND4_X1 g242 ( .A1(new_n374_), .A2(new_n371_), .A3(new_n379_), .A4(KEYINPUT48), .ZN(new_n380_) );
  INV_X1 g243 ( .A(new_n380_), .ZN(new_n381_) );
  AND3_X1 g244 ( .A1(new_n374_), .A2(new_n371_), .A3(new_n379_), .ZN(new_n382_) );
  OR2_X1 g245 ( .A1(new_n382_), .A2(KEYINPUT48), .ZN(new_n383_) );
  AND3_X1 g246 ( .A1(new_n383_), .A2(new_n221_), .A3(new_n381_), .ZN(new_n384_) );
  AND3_X1 g247 ( .A1(new_n384_), .A2(new_n213_), .A3(new_n220_), .ZN(new_n385_) );
  AND2_X1 g248 ( .A1(new_n385_), .A2(new_n294_), .ZN(new_n386_) );
  XOR2_X1 g249 ( .A(new_n386_), .B(G113GAT), .Z(G1340GAT) );
  AND2_X1 g250 ( .A1(new_n385_), .A2(new_n330_), .ZN(new_n388_) );
  XNOR2_X1 g251 ( .A(G120GAT), .B(KEYINPUT49), .ZN(new_n389_) );
  XNOR2_X1 g252 ( .A(new_n388_), .B(new_n389_), .ZN(G1341GAT) );
  AND2_X1 g253 ( .A1(new_n385_), .A2(new_n266_), .ZN(new_n391_) );
  XNOR2_X1 g254 ( .A(new_n391_), .B(KEYINPUT50), .ZN(new_n392_) );
  XOR2_X1 g255 ( .A(new_n392_), .B(G127GAT), .Z(G1342GAT) );
  AND2_X1 g256 ( .A1(new_n385_), .A2(new_n311_), .ZN(new_n394_) );
  XNOR2_X1 g257 ( .A(G134GAT), .B(KEYINPUT51), .ZN(new_n395_) );
  XNOR2_X1 g258 ( .A(new_n394_), .B(new_n395_), .ZN(G1343GAT) );
  AND2_X1 g259 ( .A1(new_n384_), .A2(new_n199_), .ZN(new_n397_) );
  AND2_X1 g260 ( .A1(new_n397_), .A2(new_n294_), .ZN(new_n398_) );
  XOR2_X1 g261 ( .A(new_n398_), .B(G141GAT), .Z(G1344GAT) );
  AND2_X1 g262 ( .A1(new_n397_), .A2(new_n330_), .ZN(new_n400_) );
  XOR2_X1 g263 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(new_n401_) );
  XNOR2_X1 g264 ( .A(new_n400_), .B(new_n401_), .ZN(new_n402_) );
  XNOR2_X1 g265 ( .A(new_n402_), .B(new_n171_), .ZN(G1345GAT) );
  AND2_X1 g266 ( .A1(new_n397_), .A2(new_n266_), .ZN(new_n404_) );
  XOR2_X1 g267 ( .A(new_n404_), .B(G155GAT), .Z(G1346GAT) );
  AND2_X1 g268 ( .A1(new_n397_), .A2(new_n311_), .ZN(new_n406_) );
  XOR2_X1 g269 ( .A(new_n406_), .B(G162GAT), .Z(G1347GAT) );
  INV_X1 g270 ( .A(KEYINPUT55), .ZN(new_n408_) );
  INV_X1 g271 ( .A(new_n182_), .ZN(new_n409_) );
  INV_X1 g272 ( .A(KEYINPUT54), .ZN(new_n410_) );
  AND4_X1 g273 ( .A1(new_n383_), .A2(new_n410_), .A3(new_n214_), .A4(new_n381_), .ZN(new_n411_) );
  INV_X1 g274 ( .A(new_n411_), .ZN(new_n412_) );
  AND3_X1 g275 ( .A1(new_n383_), .A2(new_n214_), .A3(new_n381_), .ZN(new_n413_) );
  OR2_X1 g276 ( .A1(new_n413_), .A2(new_n410_), .ZN(new_n414_) );
  AND4_X1 g277 ( .A1(new_n414_), .A2(new_n159_), .A3(new_n409_), .A4(new_n412_), .ZN(new_n415_) );
  XNOR2_X1 g278 ( .A(new_n415_), .B(new_n408_), .ZN(new_n416_) );
  AND2_X1 g279 ( .A1(new_n416_), .A2(new_n213_), .ZN(new_n417_) );
  AND2_X1 g280 ( .A1(new_n417_), .A2(new_n294_), .ZN(new_n418_) );
  XOR2_X1 g281 ( .A(new_n418_), .B(G169GAT), .Z(G1348GAT) );
  INV_X1 g282 ( .A(G176GAT), .ZN(new_n420_) );
  AND3_X1 g283 ( .A1(new_n416_), .A2(new_n213_), .A3(new_n330_), .ZN(new_n421_) );
  XOR2_X1 g284 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(new_n422_) );
  XNOR2_X1 g285 ( .A(new_n421_), .B(new_n422_), .ZN(new_n423_) );
  XNOR2_X1 g286 ( .A(new_n423_), .B(new_n420_), .ZN(G1349GAT) );
  AND2_X1 g287 ( .A1(new_n417_), .A2(new_n266_), .ZN(new_n425_) );
  XOR2_X1 g288 ( .A(new_n425_), .B(G183GAT), .Z(G1350GAT) );
  AND2_X1 g289 ( .A1(new_n417_), .A2(new_n311_), .ZN(new_n427_) );
  XOR2_X1 g290 ( .A(G190GAT), .B(KEYINPUT58), .Z(new_n428_) );
  XNOR2_X1 g291 ( .A(new_n427_), .B(new_n428_), .ZN(G1351GAT) );
  AND4_X1 g292 ( .A1(new_n414_), .A2(new_n159_), .A3(new_n199_), .A4(new_n412_), .ZN(new_n430_) );
  AND2_X1 g293 ( .A1(new_n430_), .A2(new_n294_), .ZN(new_n431_) );
  XOR2_X1 g294 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(new_n432_) );
  XNOR2_X1 g295 ( .A(new_n431_), .B(new_n432_), .ZN(new_n433_) );
  XNOR2_X1 g296 ( .A(new_n433_), .B(new_n160_), .ZN(G1352GAT) );
  AND2_X1 g297 ( .A1(new_n430_), .A2(new_n280_), .ZN(new_n435_) );
  XNOR2_X1 g298 ( .A(G204GAT), .B(KEYINPUT61), .ZN(new_n436_) );
  XNOR2_X1 g299 ( .A(new_n435_), .B(new_n436_), .ZN(G1353GAT) );
  AND2_X1 g300 ( .A1(new_n430_), .A2(new_n266_), .ZN(new_n438_) );
  XOR2_X1 g301 ( .A(new_n438_), .B(G211GAT), .Z(G1354GAT) );
  AND2_X1 g302 ( .A1(new_n430_), .A2(new_n313_), .ZN(new_n440_) );
  XNOR2_X1 g303 ( .A(new_n440_), .B(KEYINPUT62), .ZN(new_n441_) );
  XOR2_X1 g304 ( .A(new_n441_), .B(G218GAT), .Z(G1355GAT) );
endmodule


