module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917;

  AND2_X1 U1994 ( .A1(n1962), .A2(n1963), .ZN(Result_9_) );
  XOR2_X1 U1995 ( .A(n1964), .B(n1965), .Z(n1962) );
  AND2_X1 U1996 ( .A1(n1966), .A2(n1967), .ZN(n1965) );
  OR2_X1 U1997 ( .A1(n1968), .A2(n1969), .ZN(n1967) );
  AND2_X1 U1998 ( .A1(n1970), .A2(n1971), .ZN(n1969) );
  INV_X1 U1999 ( .A(n1972), .ZN(n1966) );
  AND2_X1 U2000 ( .A1(n1973), .A2(n1963), .ZN(Result_8_) );
  XOR2_X1 U2001 ( .A(n1974), .B(n1975), .Z(n1973) );
  AND2_X1 U2002 ( .A1(n1963), .A2(n1976), .ZN(Result_7_) );
  XOR2_X1 U2003 ( .A(n1977), .B(n1978), .Z(n1976) );
  AND2_X1 U2004 ( .A1(n1979), .A2(n1980), .ZN(n1978) );
  OR2_X1 U2005 ( .A1(n1981), .A2(n1982), .ZN(n1980) );
  AND2_X1 U2006 ( .A1(n1983), .A2(n1984), .ZN(n1982) );
  INV_X1 U2007 ( .A(n1985), .ZN(n1979) );
  AND2_X1 U2008 ( .A1(n1986), .A2(n1963), .ZN(Result_6_) );
  XOR2_X1 U2009 ( .A(n1987), .B(n1988), .Z(n1986) );
  AND2_X1 U2010 ( .A1(n1963), .A2(n1989), .ZN(Result_5_) );
  XOR2_X1 U2011 ( .A(n1990), .B(n1991), .Z(n1989) );
  AND2_X1 U2012 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
  OR2_X1 U2013 ( .A1(n1994), .A2(n1995), .ZN(n1993) );
  AND2_X1 U2014 ( .A1(n1996), .A2(n1997), .ZN(n1995) );
  INV_X1 U2015 ( .A(n1998), .ZN(n1992) );
  AND2_X1 U2016 ( .A1(n1999), .A2(n1963), .ZN(Result_4_) );
  XOR2_X1 U2017 ( .A(n2000), .B(n2001), .Z(n1999) );
  AND2_X1 U2018 ( .A1(n1963), .A2(n2002), .ZN(Result_3_) );
  XOR2_X1 U2019 ( .A(n2003), .B(n2004), .Z(n2002) );
  AND2_X1 U2020 ( .A1(n2005), .A2(n2006), .ZN(n2004) );
  OR2_X1 U2021 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
  AND2_X1 U2022 ( .A1(n2009), .A2(n2010), .ZN(n2008) );
  INV_X1 U2023 ( .A(n2011), .ZN(n2005) );
  OR2_X1 U2024 ( .A1(n2012), .A2(n2013), .ZN(Result_31_) );
  AND2_X1 U2025 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  AND2_X1 U2026 ( .A1(n2016), .A2(b_15_), .ZN(n2012) );
  XNOR2_X1 U2027 ( .A(n2017), .B(n2015), .ZN(n2016) );
  OR2_X1 U2028 ( .A1(n2018), .A2(n2019), .ZN(Result_30_) );
  AND2_X1 U2029 ( .A1(n2020), .A2(n2015), .ZN(n2019) );
  XOR2_X1 U2030 ( .A(n2021), .B(n2022), .Z(n2020) );
  XNOR2_X1 U2031 ( .A(n2023), .B(a_14_), .ZN(n2022) );
  AND2_X1 U2032 ( .A1(b_15_), .A2(a_15_), .ZN(n2021) );
  AND2_X1 U2033 ( .A1(n1963), .A2(n2024), .ZN(n2018) );
  OR2_X1 U2034 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
  AND2_X1 U2035 ( .A1(b_15_), .A2(n2027), .ZN(n2026) );
  OR2_X1 U2036 ( .A1(n2028), .A2(n2029), .ZN(n2027) );
  AND2_X1 U2037 ( .A1(a_14_), .A2(n2023), .ZN(n2028) );
  AND2_X1 U2038 ( .A1(b_14_), .A2(n2030), .ZN(n2025) );
  OR2_X1 U2039 ( .A1(n2014), .A2(n2031), .ZN(n2030) );
  AND2_X1 U2040 ( .A1(n2032), .A2(n1963), .ZN(Result_2_) );
  XOR2_X1 U2041 ( .A(n2033), .B(n2034), .Z(n2032) );
  OR2_X1 U2042 ( .A1(n2035), .A2(n2036), .ZN(Result_29_) );
  AND2_X1 U2043 ( .A1(n2037), .A2(n1963), .ZN(n2036) );
  XOR2_X1 U2044 ( .A(n2038), .B(n2039), .Z(n2037) );
  XNOR2_X1 U2045 ( .A(n2040), .B(n2041), .ZN(n2039) );
  AND2_X1 U2046 ( .A1(n2042), .A2(n2015), .ZN(n2035) );
  INV_X1 U2047 ( .A(n2043), .ZN(n2042) );
  AND3_X1 U2048 ( .A1(n2044), .A2(n2045), .A3(n2046), .ZN(n2043) );
  OR2_X1 U2049 ( .A1(n2047), .A2(b_13_), .ZN(n2046) );
  XNOR2_X1 U2050 ( .A(n2048), .B(a_13_), .ZN(n2047) );
  OR2_X1 U2051 ( .A1(n2049), .A2(n2048), .ZN(n2045) );
  OR2_X1 U2052 ( .A1(n2050), .A2(n2051), .ZN(n2044) );
  OR2_X1 U2053 ( .A1(n2052), .A2(n2053), .ZN(Result_28_) );
  AND2_X1 U2054 ( .A1(n2054), .A2(n1963), .ZN(n2053) );
  XOR2_X1 U2055 ( .A(n2055), .B(n2056), .Z(n2054) );
  XNOR2_X1 U2056 ( .A(n2057), .B(n2058), .ZN(n2055) );
  AND2_X1 U2057 ( .A1(n2059), .A2(n2015), .ZN(n2052) );
  XOR2_X1 U2058 ( .A(n2060), .B(n2061), .Z(n2059) );
  OR2_X1 U2059 ( .A1(n2062), .A2(n2063), .ZN(n2061) );
  OR2_X1 U2060 ( .A1(n2064), .A2(n2065), .ZN(Result_27_) );
  AND2_X1 U2061 ( .A1(n2066), .A2(n1963), .ZN(n2065) );
  XOR2_X1 U2062 ( .A(n2067), .B(n2068), .Z(n2066) );
  XNOR2_X1 U2063 ( .A(n2069), .B(n2070), .ZN(n2067) );
  AND2_X1 U2064 ( .A1(n2071), .A2(n2015), .ZN(n2064) );
  INV_X1 U2065 ( .A(n2072), .ZN(n2071) );
  AND3_X1 U2066 ( .A1(n2073), .A2(n2074), .A3(n2075), .ZN(n2072) );
  OR2_X1 U2067 ( .A1(n2076), .A2(b_11_), .ZN(n2075) );
  XNOR2_X1 U2068 ( .A(a_11_), .B(n2077), .ZN(n2076) );
  OR2_X1 U2069 ( .A1(n2078), .A2(n2079), .ZN(n2074) );
  OR2_X1 U2070 ( .A1(n2080), .A2(n2077), .ZN(n2073) );
  INV_X1 U2071 ( .A(n2078), .ZN(n2077) );
  OR2_X1 U2072 ( .A1(n2081), .A2(n2082), .ZN(Result_26_) );
  AND2_X1 U2073 ( .A1(n2083), .A2(n1963), .ZN(n2082) );
  XOR2_X1 U2074 ( .A(n2084), .B(n2085), .Z(n2083) );
  XNOR2_X1 U2075 ( .A(n2086), .B(n2087), .ZN(n2084) );
  AND2_X1 U2076 ( .A1(n2088), .A2(n2015), .ZN(n2081) );
  XOR2_X1 U2077 ( .A(n2089), .B(n2090), .Z(n2088) );
  OR2_X1 U2078 ( .A1(n2091), .A2(n2092), .ZN(n2090) );
  OR2_X1 U2079 ( .A1(n2093), .A2(n2094), .ZN(Result_25_) );
  AND2_X1 U2080 ( .A1(n2095), .A2(n1963), .ZN(n2094) );
  XNOR2_X1 U2081 ( .A(n2096), .B(n2097), .ZN(n2095) );
  XOR2_X1 U2082 ( .A(n2098), .B(n2099), .Z(n2097) );
  AND2_X1 U2083 ( .A1(n2100), .A2(n2015), .ZN(n2093) );
  XOR2_X1 U2084 ( .A(n2101), .B(n2102), .Z(n2100) );
  AND2_X1 U2085 ( .A1(n2103), .A2(n2104), .ZN(n2102) );
  INV_X1 U2086 ( .A(n2105), .ZN(n2104) );
  OR2_X1 U2087 ( .A1(n2106), .A2(n2107), .ZN(Result_24_) );
  AND2_X1 U2088 ( .A1(n2108), .A2(n1963), .ZN(n2107) );
  XNOR2_X1 U2089 ( .A(n2109), .B(n2110), .ZN(n2108) );
  XOR2_X1 U2090 ( .A(n2111), .B(n2112), .Z(n2110) );
  AND2_X1 U2091 ( .A1(n2113), .A2(n2015), .ZN(n2106) );
  XOR2_X1 U2092 ( .A(n2114), .B(n2115), .Z(n2113) );
  OR2_X1 U2093 ( .A1(n2116), .A2(n2117), .ZN(n2115) );
  OR2_X1 U2094 ( .A1(n2118), .A2(n2119), .ZN(Result_23_) );
  AND2_X1 U2095 ( .A1(n2120), .A2(n1963), .ZN(n2119) );
  XNOR2_X1 U2096 ( .A(n2121), .B(n2122), .ZN(n2120) );
  XOR2_X1 U2097 ( .A(n2123), .B(n2124), .Z(n2122) );
  AND2_X1 U2098 ( .A1(n2125), .A2(n2015), .ZN(n2118) );
  XOR2_X1 U2099 ( .A(n2126), .B(n2127), .Z(n2125) );
  AND2_X1 U2100 ( .A1(n2128), .A2(n2129), .ZN(n2127) );
  INV_X1 U2101 ( .A(n2130), .ZN(n2129) );
  OR2_X1 U2102 ( .A1(n2131), .A2(n2132), .ZN(Result_22_) );
  AND2_X1 U2103 ( .A1(n2133), .A2(n1963), .ZN(n2132) );
  XNOR2_X1 U2104 ( .A(n2134), .B(n2135), .ZN(n2133) );
  XOR2_X1 U2105 ( .A(n2136), .B(n2137), .Z(n2135) );
  AND2_X1 U2106 ( .A1(n2138), .A2(n2015), .ZN(n2131) );
  XOR2_X1 U2107 ( .A(n2139), .B(n2140), .Z(n2138) );
  OR2_X1 U2108 ( .A1(n2141), .A2(n2142), .ZN(n2140) );
  OR2_X1 U2109 ( .A1(n2143), .A2(n2144), .ZN(Result_21_) );
  AND2_X1 U2110 ( .A1(n2145), .A2(n1963), .ZN(n2144) );
  XNOR2_X1 U2111 ( .A(n2146), .B(n2147), .ZN(n2145) );
  XOR2_X1 U2112 ( .A(n2148), .B(n2149), .Z(n2147) );
  AND2_X1 U2113 ( .A1(n2150), .A2(n2015), .ZN(n2143) );
  XOR2_X1 U2114 ( .A(n2151), .B(n2152), .Z(n2150) );
  AND2_X1 U2115 ( .A1(n2153), .A2(n2154), .ZN(n2152) );
  INV_X1 U2116 ( .A(n2155), .ZN(n2154) );
  OR2_X1 U2117 ( .A1(n2156), .A2(n2157), .ZN(Result_20_) );
  AND2_X1 U2118 ( .A1(n2158), .A2(n1963), .ZN(n2157) );
  XNOR2_X1 U2119 ( .A(n2159), .B(n2160), .ZN(n2158) );
  XOR2_X1 U2120 ( .A(n2161), .B(n2162), .Z(n2160) );
  AND2_X1 U2121 ( .A1(n2163), .A2(n2015), .ZN(n2156) );
  XOR2_X1 U2122 ( .A(n2164), .B(n2165), .Z(n2163) );
  OR2_X1 U2123 ( .A1(n2166), .A2(n2167), .ZN(n2165) );
  AND2_X1 U2124 ( .A1(n1963), .A2(n2168), .ZN(Result_1_) );
  XOR2_X1 U2125 ( .A(n2169), .B(n2170), .Z(n2168) );
  AND2_X1 U2126 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
  OR2_X1 U2127 ( .A1(n2173), .A2(n2174), .ZN(n2172) );
  AND2_X1 U2128 ( .A1(n2175), .A2(n2176), .ZN(n2174) );
  INV_X1 U2129 ( .A(n2177), .ZN(n2171) );
  OR2_X1 U2130 ( .A1(n2178), .A2(n2179), .ZN(Result_19_) );
  AND2_X1 U2131 ( .A1(n2180), .A2(n1963), .ZN(n2179) );
  XNOR2_X1 U2132 ( .A(n2181), .B(n2182), .ZN(n2180) );
  XOR2_X1 U2133 ( .A(n2183), .B(n2184), .Z(n2182) );
  AND2_X1 U2134 ( .A1(n2185), .A2(n2015), .ZN(n2178) );
  XOR2_X1 U2135 ( .A(n2186), .B(n2187), .Z(n2185) );
  AND2_X1 U2136 ( .A1(n2188), .A2(n2189), .ZN(n2187) );
  INV_X1 U2137 ( .A(n2190), .ZN(n2189) );
  OR2_X1 U2138 ( .A1(n2191), .A2(n2192), .ZN(Result_18_) );
  AND2_X1 U2139 ( .A1(n2193), .A2(n1963), .ZN(n2192) );
  XNOR2_X1 U2140 ( .A(n2194), .B(n2195), .ZN(n2193) );
  XOR2_X1 U2141 ( .A(n2196), .B(n2197), .Z(n2195) );
  AND2_X1 U2142 ( .A1(n2198), .A2(n2015), .ZN(n2191) );
  XOR2_X1 U2143 ( .A(n2199), .B(n2200), .Z(n2198) );
  OR2_X1 U2144 ( .A1(n2201), .A2(n2202), .ZN(n2200) );
  OR2_X1 U2145 ( .A1(n2203), .A2(n2204), .ZN(Result_17_) );
  AND2_X1 U2146 ( .A1(n2205), .A2(n1963), .ZN(n2204) );
  XNOR2_X1 U2147 ( .A(n2206), .B(n2207), .ZN(n2205) );
  XOR2_X1 U2148 ( .A(n2208), .B(n2209), .Z(n2207) );
  AND2_X1 U2149 ( .A1(n2210), .A2(n2015), .ZN(n2203) );
  XOR2_X1 U2150 ( .A(n2211), .B(n2212), .Z(n2210) );
  AND2_X1 U2151 ( .A1(n2213), .A2(n2214), .ZN(n2212) );
  OR2_X1 U2152 ( .A1(n2215), .A2(n2216), .ZN(Result_16_) );
  AND2_X1 U2153 ( .A1(n2217), .A2(n1963), .ZN(n2216) );
  XNOR2_X1 U2154 ( .A(n2218), .B(n2219), .ZN(n2217) );
  XOR2_X1 U2155 ( .A(n2220), .B(n2221), .Z(n2219) );
  AND2_X1 U2156 ( .A1(n2222), .A2(n2015), .ZN(n2215) );
  XOR2_X1 U2157 ( .A(n2223), .B(n2224), .Z(n2222) );
  OR2_X1 U2158 ( .A1(a_0_), .A2(n2225), .ZN(n2224) );
  OR2_X1 U2159 ( .A1(n2226), .A2(n2227), .ZN(n2223) );
  AND2_X1 U2160 ( .A1(n2228), .A2(n2229), .ZN(n2227) );
  AND2_X1 U2161 ( .A1(n2211), .A2(n2230), .ZN(n2226) );
  OR2_X1 U2162 ( .A1(n2231), .A2(n2201), .ZN(n2211) );
  AND2_X1 U2163 ( .A1(n2232), .A2(n2233), .ZN(n2201) );
  AND2_X1 U2164 ( .A1(n2199), .A2(n2234), .ZN(n2231) );
  OR2_X1 U2165 ( .A1(n2235), .A2(n2236), .ZN(n2199) );
  AND2_X1 U2166 ( .A1(n2237), .A2(n2238), .ZN(n2236) );
  AND2_X1 U2167 ( .A1(n2186), .A2(n2239), .ZN(n2235) );
  OR2_X1 U2168 ( .A1(n2240), .A2(n2166), .ZN(n2186) );
  AND2_X1 U2169 ( .A1(n2241), .A2(n2242), .ZN(n2166) );
  AND2_X1 U2170 ( .A1(n2164), .A2(n2243), .ZN(n2240) );
  OR2_X1 U2171 ( .A1(n2244), .A2(n2245), .ZN(n2164) );
  AND2_X1 U2172 ( .A1(n2246), .A2(n2247), .ZN(n2245) );
  AND2_X1 U2173 ( .A1(n2151), .A2(n2248), .ZN(n2244) );
  OR2_X1 U2174 ( .A1(n2249), .A2(n2141), .ZN(n2151) );
  AND2_X1 U2175 ( .A1(n2250), .A2(n2251), .ZN(n2141) );
  AND2_X1 U2176 ( .A1(n2139), .A2(n2252), .ZN(n2249) );
  OR2_X1 U2177 ( .A1(n2253), .A2(n2254), .ZN(n2139) );
  AND2_X1 U2178 ( .A1(n2255), .A2(n2256), .ZN(n2254) );
  AND2_X1 U2179 ( .A1(n2126), .A2(n2257), .ZN(n2253) );
  OR2_X1 U2180 ( .A1(n2258), .A2(n2116), .ZN(n2126) );
  AND2_X1 U2181 ( .A1(n2259), .A2(n2260), .ZN(n2116) );
  AND2_X1 U2182 ( .A1(n2114), .A2(n2261), .ZN(n2258) );
  OR2_X1 U2183 ( .A1(n2262), .A2(n2263), .ZN(n2114) );
  AND2_X1 U2184 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  AND2_X1 U2185 ( .A1(n2101), .A2(n2266), .ZN(n2262) );
  OR2_X1 U2186 ( .A1(n2267), .A2(n2092), .ZN(n2101) );
  AND2_X1 U2187 ( .A1(n2268), .A2(n2269), .ZN(n2092) );
  AND2_X1 U2188 ( .A1(n2089), .A2(n2270), .ZN(n2267) );
  OR2_X1 U2189 ( .A1(n2271), .A2(n2272), .ZN(n2089) );
  AND2_X1 U2190 ( .A1(n2273), .A2(n2274), .ZN(n2272) );
  AND2_X1 U2191 ( .A1(n2078), .A2(n2079), .ZN(n2271) );
  OR2_X1 U2192 ( .A1(n2275), .A2(n2063), .ZN(n2078) );
  AND2_X1 U2193 ( .A1(n2276), .A2(n2277), .ZN(n2063) );
  AND2_X1 U2194 ( .A1(n2060), .A2(n2278), .ZN(n2275) );
  OR2_X1 U2195 ( .A1(n2279), .A2(n2280), .ZN(n2060) );
  AND2_X1 U2196 ( .A1(n2281), .A2(n2282), .ZN(n2280) );
  AND2_X1 U2197 ( .A1(n2051), .A2(n2050), .ZN(n2279) );
  INV_X1 U2198 ( .A(n2048), .ZN(n2051) );
  OR3_X1 U2199 ( .A1(n2283), .A2(n2284), .A3(n2285), .ZN(n2048) );
  AND2_X1 U2200 ( .A1(n2286), .A2(a_15_), .ZN(n2285) );
  INV_X1 U2201 ( .A(n2287), .ZN(n2286) );
  AND2_X1 U2202 ( .A1(n2288), .A2(b_15_), .ZN(n2284) );
  AND2_X1 U2203 ( .A1(n1963), .A2(n2289), .ZN(Result_15_) );
  XNOR2_X1 U2204 ( .A(n2290), .B(n2291), .ZN(n2289) );
  AND3_X1 U2205 ( .A1(n2292), .A2(n2293), .A3(n1963), .ZN(Result_14_) );
  OR2_X1 U2206 ( .A1(n2294), .A2(n2295), .ZN(n2292) );
  AND2_X1 U2207 ( .A1(n2296), .A2(n2291), .ZN(n2294) );
  AND2_X1 U2208 ( .A1(n1963), .A2(n2297), .ZN(Result_13_) );
  XNOR2_X1 U2209 ( .A(n2298), .B(n2299), .ZN(n2297) );
  OR2_X1 U2210 ( .A1(n2300), .A2(n2301), .ZN(n2299) );
  INV_X1 U2211 ( .A(n2302), .ZN(n2301) );
  AND2_X1 U2212 ( .A1(n2303), .A2(n2304), .ZN(n2300) );
  OR2_X1 U2213 ( .A1(n2305), .A2(n2306), .ZN(n2303) );
  AND2_X1 U2214 ( .A1(n2307), .A2(n1963), .ZN(Result_12_) );
  XNOR2_X1 U2215 ( .A(n2308), .B(n2309), .ZN(n2307) );
  AND2_X1 U2216 ( .A1(n2310), .A2(n2311), .ZN(n2309) );
  OR2_X1 U2217 ( .A1(n2312), .A2(n2313), .ZN(n2311) );
  INV_X1 U2218 ( .A(n2314), .ZN(n2310) );
  AND2_X1 U2219 ( .A1(n2315), .A2(n1963), .ZN(Result_11_) );
  XOR2_X1 U2220 ( .A(n2316), .B(n2317), .Z(n2315) );
  AND2_X1 U2221 ( .A1(n2318), .A2(n2319), .ZN(n2317) );
  OR2_X1 U2222 ( .A1(n2320), .A2(n2321), .ZN(n2319) );
  AND2_X1 U2223 ( .A1(n2322), .A2(n2323), .ZN(n2320) );
  INV_X1 U2224 ( .A(n2324), .ZN(n2318) );
  AND2_X1 U2225 ( .A1(n2325), .A2(n1963), .ZN(Result_10_) );
  XOR2_X1 U2226 ( .A(n2326), .B(n2327), .Z(n2325) );
  AND2_X1 U2227 ( .A1(n2328), .A2(n2329), .ZN(n2327) );
  OR2_X1 U2228 ( .A1(n2330), .A2(n2331), .ZN(n2329) );
  AND2_X1 U2229 ( .A1(n2332), .A2(n2333), .ZN(n2330) );
  INV_X1 U2230 ( .A(n2334), .ZN(n2328) );
  AND2_X1 U2231 ( .A1(n1963), .A2(n2335), .ZN(Result_0_) );
  OR3_X1 U2232 ( .A1(n2177), .A2(n2336), .A3(n2337), .ZN(n2335) );
  AND2_X1 U2233 ( .A1(n2169), .A2(n2173), .ZN(n2337) );
  AND2_X1 U2234 ( .A1(n2033), .A2(n2034), .ZN(n2169) );
  XOR2_X1 U2235 ( .A(n2176), .B(n2175), .Z(n2034) );
  OR2_X1 U2236 ( .A1(n2338), .A2(n2339), .ZN(n2033) );
  OR2_X1 U2237 ( .A1(n2340), .A2(n2011), .ZN(n2338) );
  AND3_X1 U2238 ( .A1(n2010), .A2(n2009), .A3(n2007), .ZN(n2011) );
  INV_X1 U2239 ( .A(n2341), .ZN(n2009) );
  AND2_X1 U2240 ( .A1(n2003), .A2(n2007), .ZN(n2340) );
  INV_X1 U2241 ( .A(n2342), .ZN(n2007) );
  OR2_X1 U2242 ( .A1(n2343), .A2(n2339), .ZN(n2342) );
  INV_X1 U2243 ( .A(n2344), .ZN(n2339) );
  OR2_X1 U2244 ( .A1(n2345), .A2(n2346), .ZN(n2344) );
  AND2_X1 U2245 ( .A1(n2345), .A2(n2346), .ZN(n2343) );
  OR2_X1 U2246 ( .A1(n2347), .A2(n2348), .ZN(n2346) );
  AND2_X1 U2247 ( .A1(n2349), .A2(n2350), .ZN(n2348) );
  AND2_X1 U2248 ( .A1(n2351), .A2(n2352), .ZN(n2347) );
  OR2_X1 U2249 ( .A1(n2350), .A2(n2349), .ZN(n2352) );
  XNOR2_X1 U2250 ( .A(n2353), .B(n2354), .ZN(n2345) );
  XOR2_X1 U2251 ( .A(n2355), .B(n2356), .Z(n2354) );
  AND2_X1 U2252 ( .A1(n2000), .A2(n2001), .ZN(n2003) );
  XNOR2_X1 U2253 ( .A(n2010), .B(n2341), .ZN(n2001) );
  OR2_X1 U2254 ( .A1(n2357), .A2(n2358), .ZN(n2341) );
  AND2_X1 U2255 ( .A1(n2359), .A2(n2360), .ZN(n2358) );
  AND2_X1 U2256 ( .A1(n2361), .A2(n2362), .ZN(n2357) );
  OR2_X1 U2257 ( .A1(n2360), .A2(n2359), .ZN(n2362) );
  XNOR2_X1 U2258 ( .A(n2351), .B(n2363), .ZN(n2010) );
  XOR2_X1 U2259 ( .A(n2350), .B(n2349), .Z(n2363) );
  OR2_X1 U2260 ( .A1(n2238), .A2(n2364), .ZN(n2349) );
  OR2_X1 U2261 ( .A1(n2365), .A2(n2366), .ZN(n2350) );
  AND2_X1 U2262 ( .A1(n2367), .A2(n2368), .ZN(n2366) );
  AND2_X1 U2263 ( .A1(n2369), .A2(n2370), .ZN(n2365) );
  OR2_X1 U2264 ( .A1(n2368), .A2(n2367), .ZN(n2370) );
  XOR2_X1 U2265 ( .A(n2371), .B(n2372), .Z(n2351) );
  XOR2_X1 U2266 ( .A(n2373), .B(n2374), .Z(n2372) );
  OR2_X1 U2267 ( .A1(n2375), .A2(n2376), .ZN(n2000) );
  OR2_X1 U2268 ( .A1(n2377), .A2(n1998), .ZN(n2375) );
  AND3_X1 U2269 ( .A1(n1997), .A2(n1996), .A3(n1994), .ZN(n1998) );
  INV_X1 U2270 ( .A(n2378), .ZN(n1996) );
  AND2_X1 U2271 ( .A1(n1990), .A2(n1994), .ZN(n2377) );
  INV_X1 U2272 ( .A(n2379), .ZN(n1994) );
  OR2_X1 U2273 ( .A1(n2380), .A2(n2376), .ZN(n2379) );
  INV_X1 U2274 ( .A(n2381), .ZN(n2376) );
  OR2_X1 U2275 ( .A1(n2382), .A2(n2383), .ZN(n2381) );
  AND2_X1 U2276 ( .A1(n2382), .A2(n2383), .ZN(n2380) );
  OR2_X1 U2277 ( .A1(n2384), .A2(n2385), .ZN(n2383) );
  AND2_X1 U2278 ( .A1(n2386), .A2(n2387), .ZN(n2385) );
  AND2_X1 U2279 ( .A1(n2388), .A2(n2389), .ZN(n2384) );
  OR2_X1 U2280 ( .A1(n2387), .A2(n2386), .ZN(n2389) );
  XOR2_X1 U2281 ( .A(n2361), .B(n2390), .Z(n2382) );
  XOR2_X1 U2282 ( .A(n2360), .B(n2359), .Z(n2390) );
  OR2_X1 U2283 ( .A1(n2242), .A2(n2364), .ZN(n2359) );
  OR2_X1 U2284 ( .A1(n2391), .A2(n2392), .ZN(n2360) );
  AND2_X1 U2285 ( .A1(n2393), .A2(n2394), .ZN(n2392) );
  AND2_X1 U2286 ( .A1(n2395), .A2(n2396), .ZN(n2391) );
  OR2_X1 U2287 ( .A1(n2394), .A2(n2393), .ZN(n2396) );
  XOR2_X1 U2288 ( .A(n2369), .B(n2397), .Z(n2361) );
  XOR2_X1 U2289 ( .A(n2368), .B(n2367), .Z(n2397) );
  OR2_X1 U2290 ( .A1(n2238), .A2(n2228), .ZN(n2367) );
  OR2_X1 U2291 ( .A1(n2398), .A2(n2399), .ZN(n2368) );
  AND2_X1 U2292 ( .A1(n2400), .A2(n2401), .ZN(n2399) );
  AND2_X1 U2293 ( .A1(n2402), .A2(n2403), .ZN(n2398) );
  OR2_X1 U2294 ( .A1(n2401), .A2(n2400), .ZN(n2403) );
  XNOR2_X1 U2295 ( .A(n2404), .B(n2405), .ZN(n2369) );
  XNOR2_X1 U2296 ( .A(n2234), .B(n2406), .ZN(n2404) );
  AND2_X1 U2297 ( .A1(n1987), .A2(n1988), .ZN(n1990) );
  XNOR2_X1 U2298 ( .A(n1997), .B(n2378), .ZN(n1988) );
  OR2_X1 U2299 ( .A1(n2407), .A2(n2408), .ZN(n2378) );
  AND2_X1 U2300 ( .A1(n2409), .A2(n2410), .ZN(n2408) );
  AND2_X1 U2301 ( .A1(n2411), .A2(n2412), .ZN(n2407) );
  OR2_X1 U2302 ( .A1(n2410), .A2(n2409), .ZN(n2412) );
  XNOR2_X1 U2303 ( .A(n2388), .B(n2413), .ZN(n1997) );
  XOR2_X1 U2304 ( .A(n2387), .B(n2386), .Z(n2413) );
  OR2_X1 U2305 ( .A1(n2247), .A2(n2364), .ZN(n2386) );
  OR2_X1 U2306 ( .A1(n2414), .A2(n2415), .ZN(n2387) );
  AND2_X1 U2307 ( .A1(n2416), .A2(n2417), .ZN(n2415) );
  AND2_X1 U2308 ( .A1(n2418), .A2(n2419), .ZN(n2414) );
  OR2_X1 U2309 ( .A1(n2417), .A2(n2416), .ZN(n2419) );
  XOR2_X1 U2310 ( .A(n2395), .B(n2420), .Z(n2388) );
  XOR2_X1 U2311 ( .A(n2394), .B(n2393), .Z(n2420) );
  OR2_X1 U2312 ( .A1(n2242), .A2(n2228), .ZN(n2393) );
  OR2_X1 U2313 ( .A1(n2421), .A2(n2422), .ZN(n2394) );
  AND2_X1 U2314 ( .A1(n2423), .A2(n2424), .ZN(n2422) );
  AND2_X1 U2315 ( .A1(n2425), .A2(n2426), .ZN(n2421) );
  OR2_X1 U2316 ( .A1(n2424), .A2(n2423), .ZN(n2426) );
  XOR2_X1 U2317 ( .A(n2402), .B(n2427), .Z(n2395) );
  XOR2_X1 U2318 ( .A(n2401), .B(n2400), .Z(n2427) );
  OR2_X1 U2319 ( .A1(n2238), .A2(n2232), .ZN(n2400) );
  OR2_X1 U2320 ( .A1(n2428), .A2(n2429), .ZN(n2401) );
  AND2_X1 U2321 ( .A1(n2239), .A2(n2430), .ZN(n2429) );
  AND2_X1 U2322 ( .A1(n2431), .A2(n2432), .ZN(n2428) );
  OR2_X1 U2323 ( .A1(n2430), .A2(n2239), .ZN(n2432) );
  XOR2_X1 U2324 ( .A(n2433), .B(n2434), .Z(n2402) );
  XOR2_X1 U2325 ( .A(n2435), .B(n2436), .Z(n2434) );
  OR2_X1 U2326 ( .A1(n2437), .A2(n2438), .ZN(n1987) );
  OR2_X1 U2327 ( .A1(n2439), .A2(n1985), .ZN(n2437) );
  AND3_X1 U2328 ( .A1(n1984), .A2(n1983), .A3(n1981), .ZN(n1985) );
  INV_X1 U2329 ( .A(n2440), .ZN(n1983) );
  AND2_X1 U2330 ( .A1(n1977), .A2(n1981), .ZN(n2439) );
  INV_X1 U2331 ( .A(n2441), .ZN(n1981) );
  OR2_X1 U2332 ( .A1(n2442), .A2(n2438), .ZN(n2441) );
  INV_X1 U2333 ( .A(n2443), .ZN(n2438) );
  OR2_X1 U2334 ( .A1(n2444), .A2(n2445), .ZN(n2443) );
  AND2_X1 U2335 ( .A1(n2444), .A2(n2445), .ZN(n2442) );
  OR2_X1 U2336 ( .A1(n2446), .A2(n2447), .ZN(n2445) );
  AND2_X1 U2337 ( .A1(n2448), .A2(n2449), .ZN(n2447) );
  AND2_X1 U2338 ( .A1(n2450), .A2(n2451), .ZN(n2446) );
  OR2_X1 U2339 ( .A1(n2449), .A2(n2448), .ZN(n2451) );
  XOR2_X1 U2340 ( .A(n2411), .B(n2452), .Z(n2444) );
  XOR2_X1 U2341 ( .A(n2410), .B(n2409), .Z(n2452) );
  OR2_X1 U2342 ( .A1(n2251), .A2(n2364), .ZN(n2409) );
  OR2_X1 U2343 ( .A1(n2453), .A2(n2454), .ZN(n2410) );
  AND2_X1 U2344 ( .A1(n2455), .A2(n2456), .ZN(n2454) );
  AND2_X1 U2345 ( .A1(n2457), .A2(n2458), .ZN(n2453) );
  OR2_X1 U2346 ( .A1(n2456), .A2(n2455), .ZN(n2458) );
  XOR2_X1 U2347 ( .A(n2418), .B(n2459), .Z(n2411) );
  XOR2_X1 U2348 ( .A(n2417), .B(n2416), .Z(n2459) );
  OR2_X1 U2349 ( .A1(n2247), .A2(n2228), .ZN(n2416) );
  OR2_X1 U2350 ( .A1(n2460), .A2(n2461), .ZN(n2417) );
  AND2_X1 U2351 ( .A1(n2462), .A2(n2463), .ZN(n2461) );
  AND2_X1 U2352 ( .A1(n2464), .A2(n2465), .ZN(n2460) );
  OR2_X1 U2353 ( .A1(n2463), .A2(n2462), .ZN(n2465) );
  XOR2_X1 U2354 ( .A(n2425), .B(n2466), .Z(n2418) );
  XOR2_X1 U2355 ( .A(n2424), .B(n2423), .Z(n2466) );
  OR2_X1 U2356 ( .A1(n2242), .A2(n2232), .ZN(n2423) );
  OR2_X1 U2357 ( .A1(n2467), .A2(n2468), .ZN(n2424) );
  AND2_X1 U2358 ( .A1(n2469), .A2(n2470), .ZN(n2468) );
  AND2_X1 U2359 ( .A1(n2471), .A2(n2472), .ZN(n2467) );
  OR2_X1 U2360 ( .A1(n2470), .A2(n2469), .ZN(n2472) );
  XOR2_X1 U2361 ( .A(n2431), .B(n2473), .Z(n2425) );
  XOR2_X1 U2362 ( .A(n2430), .B(n2239), .Z(n2473) );
  OR2_X1 U2363 ( .A1(n2237), .A2(n2238), .ZN(n2239) );
  OR2_X1 U2364 ( .A1(n2474), .A2(n2475), .ZN(n2430) );
  AND2_X1 U2365 ( .A1(n2476), .A2(n2477), .ZN(n2475) );
  AND2_X1 U2366 ( .A1(n2478), .A2(n2479), .ZN(n2474) );
  OR2_X1 U2367 ( .A1(n2477), .A2(n2476), .ZN(n2479) );
  XOR2_X1 U2368 ( .A(n2480), .B(n2481), .Z(n2431) );
  XOR2_X1 U2369 ( .A(n2482), .B(n2483), .Z(n2481) );
  AND2_X1 U2370 ( .A1(n1974), .A2(n1975), .ZN(n1977) );
  XNOR2_X1 U2371 ( .A(n1984), .B(n2440), .ZN(n1975) );
  OR2_X1 U2372 ( .A1(n2484), .A2(n2485), .ZN(n2440) );
  AND2_X1 U2373 ( .A1(n2486), .A2(n2487), .ZN(n2485) );
  AND2_X1 U2374 ( .A1(n2488), .A2(n2489), .ZN(n2484) );
  OR2_X1 U2375 ( .A1(n2487), .A2(n2486), .ZN(n2489) );
  XNOR2_X1 U2376 ( .A(n2450), .B(n2490), .ZN(n1984) );
  XOR2_X1 U2377 ( .A(n2449), .B(n2448), .Z(n2490) );
  OR2_X1 U2378 ( .A1(n2256), .A2(n2364), .ZN(n2448) );
  OR2_X1 U2379 ( .A1(n2491), .A2(n2492), .ZN(n2449) );
  AND2_X1 U2380 ( .A1(n2493), .A2(n2494), .ZN(n2492) );
  AND2_X1 U2381 ( .A1(n2495), .A2(n2496), .ZN(n2491) );
  OR2_X1 U2382 ( .A1(n2494), .A2(n2493), .ZN(n2496) );
  XOR2_X1 U2383 ( .A(n2457), .B(n2497), .Z(n2450) );
  XOR2_X1 U2384 ( .A(n2456), .B(n2455), .Z(n2497) );
  OR2_X1 U2385 ( .A1(n2251), .A2(n2228), .ZN(n2455) );
  OR2_X1 U2386 ( .A1(n2498), .A2(n2499), .ZN(n2456) );
  AND2_X1 U2387 ( .A1(n2500), .A2(n2501), .ZN(n2499) );
  AND2_X1 U2388 ( .A1(n2502), .A2(n2503), .ZN(n2498) );
  OR2_X1 U2389 ( .A1(n2501), .A2(n2500), .ZN(n2503) );
  XOR2_X1 U2390 ( .A(n2464), .B(n2504), .Z(n2457) );
  XOR2_X1 U2391 ( .A(n2463), .B(n2462), .Z(n2504) );
  OR2_X1 U2392 ( .A1(n2247), .A2(n2232), .ZN(n2462) );
  OR2_X1 U2393 ( .A1(n2505), .A2(n2506), .ZN(n2463) );
  AND2_X1 U2394 ( .A1(n2507), .A2(n2508), .ZN(n2506) );
  AND2_X1 U2395 ( .A1(n2509), .A2(n2510), .ZN(n2505) );
  OR2_X1 U2396 ( .A1(n2508), .A2(n2507), .ZN(n2510) );
  XOR2_X1 U2397 ( .A(n2471), .B(n2511), .Z(n2464) );
  XOR2_X1 U2398 ( .A(n2470), .B(n2469), .Z(n2511) );
  OR2_X1 U2399 ( .A1(n2237), .A2(n2242), .ZN(n2469) );
  OR2_X1 U2400 ( .A1(n2512), .A2(n2513), .ZN(n2470) );
  AND2_X1 U2401 ( .A1(n2514), .A2(n2243), .ZN(n2513) );
  AND2_X1 U2402 ( .A1(n2515), .A2(n2516), .ZN(n2512) );
  OR2_X1 U2403 ( .A1(n2243), .A2(n2514), .ZN(n2516) );
  XOR2_X1 U2404 ( .A(n2478), .B(n2517), .Z(n2471) );
  XOR2_X1 U2405 ( .A(n2477), .B(n2476), .Z(n2517) );
  OR2_X1 U2406 ( .A1(n2238), .A2(n2241), .ZN(n2476) );
  OR2_X1 U2407 ( .A1(n2518), .A2(n2519), .ZN(n2477) );
  AND2_X1 U2408 ( .A1(n2520), .A2(n2521), .ZN(n2519) );
  AND2_X1 U2409 ( .A1(n2522), .A2(n2523), .ZN(n2518) );
  OR2_X1 U2410 ( .A1(n2521), .A2(n2520), .ZN(n2523) );
  XOR2_X1 U2411 ( .A(n2524), .B(n2525), .Z(n2478) );
  XOR2_X1 U2412 ( .A(n2526), .B(n2527), .Z(n2525) );
  OR2_X1 U2413 ( .A1(n2528), .A2(n2529), .ZN(n1974) );
  OR2_X1 U2414 ( .A1(n2530), .A2(n1972), .ZN(n2528) );
  AND3_X1 U2415 ( .A1(n1971), .A2(n1970), .A3(n1968), .ZN(n1972) );
  INV_X1 U2416 ( .A(n2531), .ZN(n1970) );
  AND2_X1 U2417 ( .A1(n1968), .A2(n1964), .ZN(n2530) );
  OR2_X1 U2418 ( .A1(n2532), .A2(n2334), .ZN(n1964) );
  AND3_X1 U2419 ( .A1(n2333), .A2(n2331), .A3(n2332), .ZN(n2334) );
  INV_X1 U2420 ( .A(n2533), .ZN(n2332) );
  AND2_X1 U2421 ( .A1(n2331), .A2(n2326), .ZN(n2532) );
  OR2_X1 U2422 ( .A1(n2534), .A2(n2324), .ZN(n2326) );
  AND3_X1 U2423 ( .A1(n2323), .A2(n2321), .A3(n2322), .ZN(n2324) );
  INV_X1 U2424 ( .A(n2535), .ZN(n2322) );
  AND2_X1 U2425 ( .A1(n2321), .A2(n2316), .ZN(n2534) );
  OR2_X1 U2426 ( .A1(n2536), .A2(n2314), .ZN(n2316) );
  AND2_X1 U2427 ( .A1(n2313), .A2(n2312), .ZN(n2314) );
  AND2_X1 U2428 ( .A1(n2313), .A2(n2537), .ZN(n2536) );
  INV_X1 U2429 ( .A(n2308), .ZN(n2537) );
  AND2_X1 U2430 ( .A1(n2538), .A2(n2302), .ZN(n2308) );
  OR3_X1 U2431 ( .A1(n2306), .A2(n2305), .A3(n2304), .ZN(n2302) );
  OR2_X1 U2432 ( .A1(n2293), .A2(n2304), .ZN(n2538) );
  OR2_X1 U2433 ( .A1(n2539), .A2(n2312), .ZN(n2304) );
  INV_X1 U2434 ( .A(n2540), .ZN(n2312) );
  OR2_X1 U2435 ( .A1(n2541), .A2(n2542), .ZN(n2540) );
  AND2_X1 U2436 ( .A1(n2541), .A2(n2542), .ZN(n2539) );
  OR2_X1 U2437 ( .A1(n2543), .A2(n2544), .ZN(n2542) );
  AND2_X1 U2438 ( .A1(n2545), .A2(n2546), .ZN(n2544) );
  AND2_X1 U2439 ( .A1(n2547), .A2(n2548), .ZN(n2543) );
  OR2_X1 U2440 ( .A1(n2546), .A2(n2545), .ZN(n2548) );
  XOR2_X1 U2441 ( .A(n2549), .B(n2550), .Z(n2541) );
  XOR2_X1 U2442 ( .A(n2551), .B(n2552), .Z(n2550) );
  INV_X1 U2443 ( .A(n2298), .ZN(n2293) );
  AND3_X1 U2444 ( .A1(n2291), .A2(n2295), .A3(n2296), .ZN(n2298) );
  INV_X1 U2445 ( .A(n2290), .ZN(n2296) );
  OR2_X1 U2446 ( .A1(n2553), .A2(n2554), .ZN(n2290) );
  AND2_X1 U2447 ( .A1(n2221), .A2(n2220), .ZN(n2554) );
  AND2_X1 U2448 ( .A1(n2218), .A2(n2555), .ZN(n2553) );
  OR2_X1 U2449 ( .A1(n2221), .A2(n2220), .ZN(n2555) );
  OR2_X1 U2450 ( .A1(n2556), .A2(n2557), .ZN(n2220) );
  AND2_X1 U2451 ( .A1(n2209), .A2(n2208), .ZN(n2557) );
  AND2_X1 U2452 ( .A1(n2206), .A2(n2558), .ZN(n2556) );
  OR2_X1 U2453 ( .A1(n2209), .A2(n2208), .ZN(n2558) );
  OR2_X1 U2454 ( .A1(n2559), .A2(n2560), .ZN(n2208) );
  AND2_X1 U2455 ( .A1(n2197), .A2(n2196), .ZN(n2560) );
  AND2_X1 U2456 ( .A1(n2194), .A2(n2561), .ZN(n2559) );
  OR2_X1 U2457 ( .A1(n2197), .A2(n2196), .ZN(n2561) );
  OR2_X1 U2458 ( .A1(n2562), .A2(n2563), .ZN(n2196) );
  AND2_X1 U2459 ( .A1(n2184), .A2(n2183), .ZN(n2563) );
  AND2_X1 U2460 ( .A1(n2181), .A2(n2564), .ZN(n2562) );
  OR2_X1 U2461 ( .A1(n2184), .A2(n2183), .ZN(n2564) );
  OR2_X1 U2462 ( .A1(n2565), .A2(n2566), .ZN(n2183) );
  AND2_X1 U2463 ( .A1(n2162), .A2(n2161), .ZN(n2566) );
  AND2_X1 U2464 ( .A1(n2159), .A2(n2567), .ZN(n2565) );
  OR2_X1 U2465 ( .A1(n2162), .A2(n2161), .ZN(n2567) );
  OR2_X1 U2466 ( .A1(n2568), .A2(n2569), .ZN(n2161) );
  AND2_X1 U2467 ( .A1(n2149), .A2(n2148), .ZN(n2569) );
  AND2_X1 U2468 ( .A1(n2146), .A2(n2570), .ZN(n2568) );
  OR2_X1 U2469 ( .A1(n2149), .A2(n2148), .ZN(n2570) );
  OR2_X1 U2470 ( .A1(n2571), .A2(n2572), .ZN(n2148) );
  AND2_X1 U2471 ( .A1(n2137), .A2(n2136), .ZN(n2572) );
  AND2_X1 U2472 ( .A1(n2134), .A2(n2573), .ZN(n2571) );
  OR2_X1 U2473 ( .A1(n2137), .A2(n2136), .ZN(n2573) );
  OR2_X1 U2474 ( .A1(n2574), .A2(n2575), .ZN(n2136) );
  AND2_X1 U2475 ( .A1(n2124), .A2(n2123), .ZN(n2575) );
  AND2_X1 U2476 ( .A1(n2121), .A2(n2576), .ZN(n2574) );
  OR2_X1 U2477 ( .A1(n2124), .A2(n2123), .ZN(n2576) );
  OR2_X1 U2478 ( .A1(n2577), .A2(n2578), .ZN(n2123) );
  AND2_X1 U2479 ( .A1(n2112), .A2(n2111), .ZN(n2578) );
  AND2_X1 U2480 ( .A1(n2109), .A2(n2579), .ZN(n2577) );
  OR2_X1 U2481 ( .A1(n2112), .A2(n2111), .ZN(n2579) );
  OR2_X1 U2482 ( .A1(n2580), .A2(n2581), .ZN(n2111) );
  AND2_X1 U2483 ( .A1(n2099), .A2(n2098), .ZN(n2581) );
  AND2_X1 U2484 ( .A1(n2096), .A2(n2582), .ZN(n2580) );
  OR2_X1 U2485 ( .A1(n2099), .A2(n2098), .ZN(n2582) );
  OR2_X1 U2486 ( .A1(n2583), .A2(n2584), .ZN(n2098) );
  AND2_X1 U2487 ( .A1(n2087), .A2(n2086), .ZN(n2584) );
  AND2_X1 U2488 ( .A1(n2085), .A2(n2585), .ZN(n2583) );
  OR2_X1 U2489 ( .A1(n2087), .A2(n2086), .ZN(n2585) );
  OR2_X1 U2490 ( .A1(n2586), .A2(n2587), .ZN(n2086) );
  AND2_X1 U2491 ( .A1(n2070), .A2(n2069), .ZN(n2587) );
  AND2_X1 U2492 ( .A1(n2068), .A2(n2588), .ZN(n2586) );
  OR2_X1 U2493 ( .A1(n2070), .A2(n2069), .ZN(n2588) );
  OR2_X1 U2494 ( .A1(n2589), .A2(n2590), .ZN(n2069) );
  AND2_X1 U2495 ( .A1(n2058), .A2(n2057), .ZN(n2590) );
  AND2_X1 U2496 ( .A1(n2056), .A2(n2591), .ZN(n2589) );
  OR2_X1 U2497 ( .A1(n2058), .A2(n2057), .ZN(n2591) );
  OR2_X1 U2498 ( .A1(n2592), .A2(n2593), .ZN(n2057) );
  AND2_X1 U2499 ( .A1(n2038), .A2(n2041), .ZN(n2593) );
  AND2_X1 U2500 ( .A1(n2040), .A2(n2594), .ZN(n2592) );
  OR2_X1 U2501 ( .A1(n2038), .A2(n2041), .ZN(n2594) );
  OR2_X1 U2502 ( .A1(n2595), .A2(n2281), .ZN(n2041) );
  OR2_X1 U2503 ( .A1(n2287), .A2(n2596), .ZN(n2038) );
  INV_X1 U2504 ( .A(n2597), .ZN(n2040) );
  OR3_X1 U2505 ( .A1(n2598), .A2(n2599), .A3(n2600), .ZN(n2597) );
  AND2_X1 U2506 ( .A1(n2029), .A2(b_14_), .ZN(n2600) );
  AND2_X1 U2507 ( .A1(b_13_), .A2(n2601), .ZN(n2599) );
  OR2_X1 U2508 ( .A1(n2602), .A2(n2031), .ZN(n2601) );
  AND2_X1 U2509 ( .A1(a_15_), .A2(n2023), .ZN(n2602) );
  AND2_X1 U2510 ( .A1(n2283), .A2(n2282), .ZN(n2598) );
  AND2_X1 U2511 ( .A1(a_14_), .A2(b_14_), .ZN(n2283) );
  OR2_X1 U2512 ( .A1(n2595), .A2(n2276), .ZN(n2058) );
  XNOR2_X1 U2513 ( .A(n2603), .B(n2604), .ZN(n2056) );
  XNOR2_X1 U2514 ( .A(n2605), .B(n2606), .ZN(n2604) );
  OR2_X1 U2515 ( .A1(n2595), .A2(n2273), .ZN(n2070) );
  XOR2_X1 U2516 ( .A(n2607), .B(n2608), .Z(n2068) );
  XOR2_X1 U2517 ( .A(n2609), .B(n2610), .Z(n2608) );
  OR2_X1 U2518 ( .A1(n2595), .A2(n2268), .ZN(n2087) );
  XOR2_X1 U2519 ( .A(n2611), .B(n2612), .Z(n2085) );
  XOR2_X1 U2520 ( .A(n2613), .B(n2614), .Z(n2612) );
  OR2_X1 U2521 ( .A1(n2264), .A2(n2595), .ZN(n2099) );
  XOR2_X1 U2522 ( .A(n2615), .B(n2616), .Z(n2096) );
  XOR2_X1 U2523 ( .A(n2617), .B(n2618), .Z(n2616) );
  OR2_X1 U2524 ( .A1(n2595), .A2(n2259), .ZN(n2112) );
  XOR2_X1 U2525 ( .A(n2619), .B(n2620), .Z(n2109) );
  XOR2_X1 U2526 ( .A(n2621), .B(n2622), .Z(n2620) );
  OR2_X1 U2527 ( .A1(n2255), .A2(n2595), .ZN(n2124) );
  XOR2_X1 U2528 ( .A(n2623), .B(n2624), .Z(n2121) );
  XOR2_X1 U2529 ( .A(n2625), .B(n2626), .Z(n2624) );
  OR2_X1 U2530 ( .A1(n2595), .A2(n2250), .ZN(n2137) );
  XOR2_X1 U2531 ( .A(n2627), .B(n2628), .Z(n2134) );
  XOR2_X1 U2532 ( .A(n2629), .B(n2630), .Z(n2628) );
  OR2_X1 U2533 ( .A1(n2246), .A2(n2595), .ZN(n2149) );
  XOR2_X1 U2534 ( .A(n2631), .B(n2632), .Z(n2146) );
  XOR2_X1 U2535 ( .A(n2633), .B(n2634), .Z(n2632) );
  OR2_X1 U2536 ( .A1(n2595), .A2(n2241), .ZN(n2162) );
  XOR2_X1 U2537 ( .A(n2635), .B(n2636), .Z(n2159) );
  XOR2_X1 U2538 ( .A(n2637), .B(n2638), .Z(n2636) );
  OR2_X1 U2539 ( .A1(n2237), .A2(n2595), .ZN(n2184) );
  XOR2_X1 U2540 ( .A(n2639), .B(n2640), .Z(n2181) );
  XOR2_X1 U2541 ( .A(n2641), .B(n2642), .Z(n2640) );
  OR2_X1 U2542 ( .A1(n2595), .A2(n2232), .ZN(n2197) );
  XOR2_X1 U2543 ( .A(n2643), .B(n2644), .Z(n2194) );
  XOR2_X1 U2544 ( .A(n2645), .B(n2646), .Z(n2644) );
  OR2_X1 U2545 ( .A1(n2595), .A2(n2228), .ZN(n2209) );
  XOR2_X1 U2546 ( .A(n2647), .B(n2648), .Z(n2206) );
  XOR2_X1 U2547 ( .A(n2649), .B(n2650), .Z(n2648) );
  OR2_X1 U2548 ( .A1(n2595), .A2(n2364), .ZN(n2221) );
  XOR2_X1 U2549 ( .A(n2651), .B(n2652), .Z(n2218) );
  XOR2_X1 U2550 ( .A(n2653), .B(n2654), .Z(n2652) );
  XOR2_X1 U2551 ( .A(n2305), .B(n2306), .Z(n2295) );
  OR2_X1 U2552 ( .A1(n2655), .A2(n2656), .ZN(n2306) );
  AND2_X1 U2553 ( .A1(n2657), .A2(n2658), .ZN(n2656) );
  AND2_X1 U2554 ( .A1(n2659), .A2(n2660), .ZN(n2655) );
  OR2_X1 U2555 ( .A1(n2657), .A2(n2658), .ZN(n2660) );
  XOR2_X1 U2556 ( .A(n2547), .B(n2661), .Z(n2305) );
  XOR2_X1 U2557 ( .A(n2546), .B(n2545), .Z(n2661) );
  OR2_X1 U2558 ( .A1(n2282), .A2(n2364), .ZN(n2545) );
  OR2_X1 U2559 ( .A1(n2662), .A2(n2663), .ZN(n2546) );
  AND2_X1 U2560 ( .A1(n2664), .A2(n2665), .ZN(n2663) );
  AND2_X1 U2561 ( .A1(n2666), .A2(n2667), .ZN(n2662) );
  OR2_X1 U2562 ( .A1(n2665), .A2(n2664), .ZN(n2667) );
  XOR2_X1 U2563 ( .A(n2668), .B(n2669), .Z(n2547) );
  XOR2_X1 U2564 ( .A(n2670), .B(n2671), .Z(n2669) );
  XNOR2_X1 U2565 ( .A(n2659), .B(n2672), .ZN(n2291) );
  XOR2_X1 U2566 ( .A(n2658), .B(n2657), .Z(n2672) );
  OR2_X1 U2567 ( .A1(n2023), .A2(n2364), .ZN(n2657) );
  OR2_X1 U2568 ( .A1(n2673), .A2(n2674), .ZN(n2658) );
  AND2_X1 U2569 ( .A1(n2654), .A2(n2653), .ZN(n2674) );
  AND2_X1 U2570 ( .A1(n2651), .A2(n2675), .ZN(n2673) );
  OR2_X1 U2571 ( .A1(n2653), .A2(n2654), .ZN(n2675) );
  OR2_X1 U2572 ( .A1(n2023), .A2(n2228), .ZN(n2654) );
  OR2_X1 U2573 ( .A1(n2676), .A2(n2677), .ZN(n2653) );
  AND2_X1 U2574 ( .A1(n2650), .A2(n2649), .ZN(n2677) );
  AND2_X1 U2575 ( .A1(n2647), .A2(n2678), .ZN(n2676) );
  OR2_X1 U2576 ( .A1(n2649), .A2(n2650), .ZN(n2678) );
  OR2_X1 U2577 ( .A1(n2023), .A2(n2232), .ZN(n2650) );
  OR2_X1 U2578 ( .A1(n2679), .A2(n2680), .ZN(n2649) );
  AND2_X1 U2579 ( .A1(n2646), .A2(n2645), .ZN(n2680) );
  AND2_X1 U2580 ( .A1(n2643), .A2(n2681), .ZN(n2679) );
  OR2_X1 U2581 ( .A1(n2645), .A2(n2646), .ZN(n2681) );
  OR2_X1 U2582 ( .A1(n2237), .A2(n2023), .ZN(n2646) );
  OR2_X1 U2583 ( .A1(n2682), .A2(n2683), .ZN(n2645) );
  AND2_X1 U2584 ( .A1(n2642), .A2(n2641), .ZN(n2683) );
  AND2_X1 U2585 ( .A1(n2639), .A2(n2684), .ZN(n2682) );
  OR2_X1 U2586 ( .A1(n2641), .A2(n2642), .ZN(n2684) );
  OR2_X1 U2587 ( .A1(n2023), .A2(n2241), .ZN(n2642) );
  OR2_X1 U2588 ( .A1(n2685), .A2(n2686), .ZN(n2641) );
  AND2_X1 U2589 ( .A1(n2638), .A2(n2637), .ZN(n2686) );
  AND2_X1 U2590 ( .A1(n2635), .A2(n2687), .ZN(n2685) );
  OR2_X1 U2591 ( .A1(n2637), .A2(n2638), .ZN(n2687) );
  OR2_X1 U2592 ( .A1(n2246), .A2(n2023), .ZN(n2638) );
  OR2_X1 U2593 ( .A1(n2688), .A2(n2689), .ZN(n2637) );
  AND2_X1 U2594 ( .A1(n2634), .A2(n2633), .ZN(n2689) );
  AND2_X1 U2595 ( .A1(n2631), .A2(n2690), .ZN(n2688) );
  OR2_X1 U2596 ( .A1(n2633), .A2(n2634), .ZN(n2690) );
  OR2_X1 U2597 ( .A1(n2023), .A2(n2250), .ZN(n2634) );
  OR2_X1 U2598 ( .A1(n2691), .A2(n2692), .ZN(n2633) );
  AND2_X1 U2599 ( .A1(n2630), .A2(n2629), .ZN(n2692) );
  AND2_X1 U2600 ( .A1(n2627), .A2(n2693), .ZN(n2691) );
  OR2_X1 U2601 ( .A1(n2629), .A2(n2630), .ZN(n2693) );
  OR2_X1 U2602 ( .A1(n2255), .A2(n2023), .ZN(n2630) );
  OR2_X1 U2603 ( .A1(n2694), .A2(n2695), .ZN(n2629) );
  AND2_X1 U2604 ( .A1(n2626), .A2(n2625), .ZN(n2695) );
  AND2_X1 U2605 ( .A1(n2623), .A2(n2696), .ZN(n2694) );
  OR2_X1 U2606 ( .A1(n2625), .A2(n2626), .ZN(n2696) );
  OR2_X1 U2607 ( .A1(n2023), .A2(n2259), .ZN(n2626) );
  OR2_X1 U2608 ( .A1(n2697), .A2(n2698), .ZN(n2625) );
  AND2_X1 U2609 ( .A1(n2622), .A2(n2621), .ZN(n2698) );
  AND2_X1 U2610 ( .A1(n2619), .A2(n2699), .ZN(n2697) );
  OR2_X1 U2611 ( .A1(n2621), .A2(n2622), .ZN(n2699) );
  OR2_X1 U2612 ( .A1(n2264), .A2(n2023), .ZN(n2622) );
  OR2_X1 U2613 ( .A1(n2700), .A2(n2701), .ZN(n2621) );
  AND2_X1 U2614 ( .A1(n2618), .A2(n2617), .ZN(n2701) );
  AND2_X1 U2615 ( .A1(n2615), .A2(n2702), .ZN(n2700) );
  OR2_X1 U2616 ( .A1(n2617), .A2(n2618), .ZN(n2702) );
  OR2_X1 U2617 ( .A1(n2023), .A2(n2268), .ZN(n2618) );
  OR2_X1 U2618 ( .A1(n2703), .A2(n2704), .ZN(n2617) );
  AND2_X1 U2619 ( .A1(n2614), .A2(n2613), .ZN(n2704) );
  AND2_X1 U2620 ( .A1(n2611), .A2(n2705), .ZN(n2703) );
  OR2_X1 U2621 ( .A1(n2613), .A2(n2614), .ZN(n2705) );
  OR2_X1 U2622 ( .A1(n2023), .A2(n2273), .ZN(n2614) );
  OR2_X1 U2623 ( .A1(n2706), .A2(n2707), .ZN(n2613) );
  AND2_X1 U2624 ( .A1(n2610), .A2(n2609), .ZN(n2707) );
  AND2_X1 U2625 ( .A1(n2607), .A2(n2708), .ZN(n2706) );
  OR2_X1 U2626 ( .A1(n2609), .A2(n2610), .ZN(n2708) );
  OR2_X1 U2627 ( .A1(n2023), .A2(n2276), .ZN(n2610) );
  OR2_X1 U2628 ( .A1(n2709), .A2(n2710), .ZN(n2609) );
  AND2_X1 U2629 ( .A1(n2603), .A2(n2606), .ZN(n2710) );
  AND2_X1 U2630 ( .A1(n2605), .A2(n2711), .ZN(n2709) );
  OR2_X1 U2631 ( .A1(n2606), .A2(n2603), .ZN(n2711) );
  OR2_X1 U2632 ( .A1(n2023), .A2(n2281), .ZN(n2603) );
  OR3_X1 U2633 ( .A1(n2023), .A2(n2282), .A3(n2596), .ZN(n2606) );
  INV_X1 U2634 ( .A(n2712), .ZN(n2605) );
  OR2_X1 U2635 ( .A1(n2713), .A2(n2714), .ZN(n2712) );
  AND2_X1 U2636 ( .A1(b_13_), .A2(n2715), .ZN(n2714) );
  OR2_X1 U2637 ( .A1(n2716), .A2(n2029), .ZN(n2715) );
  AND2_X1 U2638 ( .A1(a_14_), .A2(n2277), .ZN(n2716) );
  AND2_X1 U2639 ( .A1(b_12_), .A2(n2717), .ZN(n2713) );
  OR2_X1 U2640 ( .A1(n2718), .A2(n2031), .ZN(n2717) );
  AND2_X1 U2641 ( .A1(a_15_), .A2(n2282), .ZN(n2718) );
  XNOR2_X1 U2642 ( .A(n2050), .B(n2719), .ZN(n2607) );
  XNOR2_X1 U2643 ( .A(n2720), .B(n2721), .ZN(n2719) );
  XOR2_X1 U2644 ( .A(n2722), .B(n2723), .Z(n2611) );
  XOR2_X1 U2645 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR2_X1 U2646 ( .A(n2726), .B(n2727), .Z(n2615) );
  XOR2_X1 U2647 ( .A(n2728), .B(n2729), .Z(n2727) );
  XOR2_X1 U2648 ( .A(n2730), .B(n2731), .Z(n2619) );
  XOR2_X1 U2649 ( .A(n2732), .B(n2733), .Z(n2731) );
  XOR2_X1 U2650 ( .A(n2734), .B(n2735), .Z(n2623) );
  XOR2_X1 U2651 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR2_X1 U2652 ( .A(n2738), .B(n2739), .Z(n2627) );
  XOR2_X1 U2653 ( .A(n2740), .B(n2741), .Z(n2739) );
  XOR2_X1 U2654 ( .A(n2742), .B(n2743), .Z(n2631) );
  XOR2_X1 U2655 ( .A(n2744), .B(n2745), .Z(n2743) );
  XOR2_X1 U2656 ( .A(n2746), .B(n2747), .Z(n2635) );
  XOR2_X1 U2657 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR2_X1 U2658 ( .A(n2750), .B(n2751), .Z(n2639) );
  XOR2_X1 U2659 ( .A(n2752), .B(n2753), .Z(n2751) );
  XOR2_X1 U2660 ( .A(n2754), .B(n2755), .Z(n2643) );
  XOR2_X1 U2661 ( .A(n2756), .B(n2757), .Z(n2755) );
  XOR2_X1 U2662 ( .A(n2758), .B(n2759), .Z(n2647) );
  XOR2_X1 U2663 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR2_X1 U2664 ( .A(n2762), .B(n2763), .Z(n2651) );
  XOR2_X1 U2665 ( .A(n2764), .B(n2765), .Z(n2763) );
  XOR2_X1 U2666 ( .A(n2666), .B(n2766), .Z(n2659) );
  XOR2_X1 U2667 ( .A(n2665), .B(n2664), .Z(n2766) );
  OR2_X1 U2668 ( .A1(n2282), .A2(n2228), .ZN(n2664) );
  OR2_X1 U2669 ( .A1(n2767), .A2(n2768), .ZN(n2665) );
  AND2_X1 U2670 ( .A1(n2765), .A2(n2764), .ZN(n2768) );
  AND2_X1 U2671 ( .A1(n2762), .A2(n2769), .ZN(n2767) );
  OR2_X1 U2672 ( .A1(n2764), .A2(n2765), .ZN(n2769) );
  OR2_X1 U2673 ( .A1(n2282), .A2(n2232), .ZN(n2765) );
  OR2_X1 U2674 ( .A1(n2770), .A2(n2771), .ZN(n2764) );
  AND2_X1 U2675 ( .A1(n2761), .A2(n2760), .ZN(n2771) );
  AND2_X1 U2676 ( .A1(n2758), .A2(n2772), .ZN(n2770) );
  OR2_X1 U2677 ( .A1(n2760), .A2(n2761), .ZN(n2772) );
  OR2_X1 U2678 ( .A1(n2237), .A2(n2282), .ZN(n2761) );
  OR2_X1 U2679 ( .A1(n2773), .A2(n2774), .ZN(n2760) );
  AND2_X1 U2680 ( .A1(n2757), .A2(n2756), .ZN(n2774) );
  AND2_X1 U2681 ( .A1(n2754), .A2(n2775), .ZN(n2773) );
  OR2_X1 U2682 ( .A1(n2756), .A2(n2757), .ZN(n2775) );
  OR2_X1 U2683 ( .A1(n2282), .A2(n2241), .ZN(n2757) );
  OR2_X1 U2684 ( .A1(n2776), .A2(n2777), .ZN(n2756) );
  AND2_X1 U2685 ( .A1(n2753), .A2(n2752), .ZN(n2777) );
  AND2_X1 U2686 ( .A1(n2750), .A2(n2778), .ZN(n2776) );
  OR2_X1 U2687 ( .A1(n2752), .A2(n2753), .ZN(n2778) );
  OR2_X1 U2688 ( .A1(n2246), .A2(n2282), .ZN(n2753) );
  OR2_X1 U2689 ( .A1(n2779), .A2(n2780), .ZN(n2752) );
  AND2_X1 U2690 ( .A1(n2749), .A2(n2748), .ZN(n2780) );
  AND2_X1 U2691 ( .A1(n2746), .A2(n2781), .ZN(n2779) );
  OR2_X1 U2692 ( .A1(n2748), .A2(n2749), .ZN(n2781) );
  OR2_X1 U2693 ( .A1(n2282), .A2(n2250), .ZN(n2749) );
  OR2_X1 U2694 ( .A1(n2782), .A2(n2783), .ZN(n2748) );
  AND2_X1 U2695 ( .A1(n2745), .A2(n2744), .ZN(n2783) );
  AND2_X1 U2696 ( .A1(n2742), .A2(n2784), .ZN(n2782) );
  OR2_X1 U2697 ( .A1(n2744), .A2(n2745), .ZN(n2784) );
  OR2_X1 U2698 ( .A1(n2255), .A2(n2282), .ZN(n2745) );
  OR2_X1 U2699 ( .A1(n2785), .A2(n2786), .ZN(n2744) );
  AND2_X1 U2700 ( .A1(n2741), .A2(n2740), .ZN(n2786) );
  AND2_X1 U2701 ( .A1(n2738), .A2(n2787), .ZN(n2785) );
  OR2_X1 U2702 ( .A1(n2740), .A2(n2741), .ZN(n2787) );
  OR2_X1 U2703 ( .A1(n2282), .A2(n2259), .ZN(n2741) );
  OR2_X1 U2704 ( .A1(n2788), .A2(n2789), .ZN(n2740) );
  AND2_X1 U2705 ( .A1(n2737), .A2(n2736), .ZN(n2789) );
  AND2_X1 U2706 ( .A1(n2734), .A2(n2790), .ZN(n2788) );
  OR2_X1 U2707 ( .A1(n2736), .A2(n2737), .ZN(n2790) );
  OR2_X1 U2708 ( .A1(n2264), .A2(n2282), .ZN(n2737) );
  OR2_X1 U2709 ( .A1(n2791), .A2(n2792), .ZN(n2736) );
  AND2_X1 U2710 ( .A1(n2733), .A2(n2732), .ZN(n2792) );
  AND2_X1 U2711 ( .A1(n2730), .A2(n2793), .ZN(n2791) );
  OR2_X1 U2712 ( .A1(n2732), .A2(n2733), .ZN(n2793) );
  OR2_X1 U2713 ( .A1(n2282), .A2(n2268), .ZN(n2733) );
  OR2_X1 U2714 ( .A1(n2794), .A2(n2795), .ZN(n2732) );
  AND2_X1 U2715 ( .A1(n2729), .A2(n2728), .ZN(n2795) );
  AND2_X1 U2716 ( .A1(n2726), .A2(n2796), .ZN(n2794) );
  OR2_X1 U2717 ( .A1(n2728), .A2(n2729), .ZN(n2796) );
  OR2_X1 U2718 ( .A1(n2282), .A2(n2273), .ZN(n2729) );
  OR2_X1 U2719 ( .A1(n2797), .A2(n2798), .ZN(n2728) );
  AND2_X1 U2720 ( .A1(n2725), .A2(n2724), .ZN(n2798) );
  AND2_X1 U2721 ( .A1(n2722), .A2(n2799), .ZN(n2797) );
  OR2_X1 U2722 ( .A1(n2724), .A2(n2725), .ZN(n2799) );
  OR2_X1 U2723 ( .A1(n2282), .A2(n2276), .ZN(n2725) );
  OR2_X1 U2724 ( .A1(n2800), .A2(n2801), .ZN(n2724) );
  AND2_X1 U2725 ( .A1(n2050), .A2(n2721), .ZN(n2801) );
  AND2_X1 U2726 ( .A1(n2720), .A2(n2802), .ZN(n2800) );
  OR2_X1 U2727 ( .A1(n2721), .A2(n2050), .ZN(n2802) );
  OR2_X1 U2728 ( .A1(n2282), .A2(n2281), .ZN(n2050) );
  OR3_X1 U2729 ( .A1(n2282), .A2(n2277), .A3(n2596), .ZN(n2721) );
  INV_X1 U2730 ( .A(n2803), .ZN(n2720) );
  OR2_X1 U2731 ( .A1(n2804), .A2(n2805), .ZN(n2803) );
  AND2_X1 U2732 ( .A1(b_12_), .A2(n2806), .ZN(n2805) );
  OR2_X1 U2733 ( .A1(n2807), .A2(n2029), .ZN(n2806) );
  AND2_X1 U2734 ( .A1(a_14_), .A2(n2274), .ZN(n2807) );
  AND2_X1 U2735 ( .A1(b_11_), .A2(n2808), .ZN(n2804) );
  OR2_X1 U2736 ( .A1(n2809), .A2(n2031), .ZN(n2808) );
  AND2_X1 U2737 ( .A1(a_15_), .A2(n2277), .ZN(n2809) );
  XNOR2_X1 U2738 ( .A(n2810), .B(n2811), .ZN(n2722) );
  XNOR2_X1 U2739 ( .A(n2812), .B(n2813), .ZN(n2811) );
  XOR2_X1 U2740 ( .A(n2814), .B(n2815), .Z(n2726) );
  XNOR2_X1 U2741 ( .A(n2816), .B(n2062), .ZN(n2815) );
  XOR2_X1 U2742 ( .A(n2817), .B(n2818), .Z(n2730) );
  XOR2_X1 U2743 ( .A(n2819), .B(n2820), .Z(n2818) );
  XOR2_X1 U2744 ( .A(n2821), .B(n2822), .Z(n2734) );
  XOR2_X1 U2745 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR2_X1 U2746 ( .A(n2825), .B(n2826), .Z(n2738) );
  XOR2_X1 U2747 ( .A(n2827), .B(n2828), .Z(n2826) );
  XOR2_X1 U2748 ( .A(n2829), .B(n2830), .Z(n2742) );
  XOR2_X1 U2749 ( .A(n2831), .B(n2832), .Z(n2830) );
  XOR2_X1 U2750 ( .A(n2833), .B(n2834), .Z(n2746) );
  XOR2_X1 U2751 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR2_X1 U2752 ( .A(n2837), .B(n2838), .Z(n2750) );
  XOR2_X1 U2753 ( .A(n2839), .B(n2840), .Z(n2838) );
  XOR2_X1 U2754 ( .A(n2841), .B(n2842), .Z(n2754) );
  XOR2_X1 U2755 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR2_X1 U2756 ( .A(n2845), .B(n2846), .Z(n2758) );
  XOR2_X1 U2757 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR2_X1 U2758 ( .A(n2849), .B(n2850), .Z(n2762) );
  XOR2_X1 U2759 ( .A(n2851), .B(n2852), .Z(n2850) );
  XOR2_X1 U2760 ( .A(n2853), .B(n2854), .Z(n2666) );
  XOR2_X1 U2761 ( .A(n2855), .B(n2856), .Z(n2854) );
  XNOR2_X1 U2762 ( .A(n2323), .B(n2535), .ZN(n2313) );
  OR2_X1 U2763 ( .A1(n2857), .A2(n2858), .ZN(n2535) );
  AND2_X1 U2764 ( .A1(n2552), .A2(n2551), .ZN(n2858) );
  AND2_X1 U2765 ( .A1(n2549), .A2(n2859), .ZN(n2857) );
  OR2_X1 U2766 ( .A1(n2551), .A2(n2552), .ZN(n2859) );
  OR2_X1 U2767 ( .A1(n2277), .A2(n2364), .ZN(n2552) );
  OR2_X1 U2768 ( .A1(n2860), .A2(n2861), .ZN(n2551) );
  AND2_X1 U2769 ( .A1(n2671), .A2(n2670), .ZN(n2861) );
  AND2_X1 U2770 ( .A1(n2668), .A2(n2862), .ZN(n2860) );
  OR2_X1 U2771 ( .A1(n2670), .A2(n2671), .ZN(n2862) );
  OR2_X1 U2772 ( .A1(n2277), .A2(n2228), .ZN(n2671) );
  OR2_X1 U2773 ( .A1(n2863), .A2(n2864), .ZN(n2670) );
  AND2_X1 U2774 ( .A1(n2856), .A2(n2855), .ZN(n2864) );
  AND2_X1 U2775 ( .A1(n2853), .A2(n2865), .ZN(n2863) );
  OR2_X1 U2776 ( .A1(n2855), .A2(n2856), .ZN(n2865) );
  OR2_X1 U2777 ( .A1(n2277), .A2(n2232), .ZN(n2856) );
  OR2_X1 U2778 ( .A1(n2866), .A2(n2867), .ZN(n2855) );
  AND2_X1 U2779 ( .A1(n2852), .A2(n2851), .ZN(n2867) );
  AND2_X1 U2780 ( .A1(n2849), .A2(n2868), .ZN(n2866) );
  OR2_X1 U2781 ( .A1(n2851), .A2(n2852), .ZN(n2868) );
  OR2_X1 U2782 ( .A1(n2237), .A2(n2277), .ZN(n2852) );
  OR2_X1 U2783 ( .A1(n2869), .A2(n2870), .ZN(n2851) );
  AND2_X1 U2784 ( .A1(n2848), .A2(n2847), .ZN(n2870) );
  AND2_X1 U2785 ( .A1(n2845), .A2(n2871), .ZN(n2869) );
  OR2_X1 U2786 ( .A1(n2847), .A2(n2848), .ZN(n2871) );
  OR2_X1 U2787 ( .A1(n2277), .A2(n2241), .ZN(n2848) );
  OR2_X1 U2788 ( .A1(n2872), .A2(n2873), .ZN(n2847) );
  AND2_X1 U2789 ( .A1(n2844), .A2(n2843), .ZN(n2873) );
  AND2_X1 U2790 ( .A1(n2841), .A2(n2874), .ZN(n2872) );
  OR2_X1 U2791 ( .A1(n2843), .A2(n2844), .ZN(n2874) );
  OR2_X1 U2792 ( .A1(n2246), .A2(n2277), .ZN(n2844) );
  OR2_X1 U2793 ( .A1(n2875), .A2(n2876), .ZN(n2843) );
  AND2_X1 U2794 ( .A1(n2840), .A2(n2839), .ZN(n2876) );
  AND2_X1 U2795 ( .A1(n2837), .A2(n2877), .ZN(n2875) );
  OR2_X1 U2796 ( .A1(n2839), .A2(n2840), .ZN(n2877) );
  OR2_X1 U2797 ( .A1(n2277), .A2(n2250), .ZN(n2840) );
  OR2_X1 U2798 ( .A1(n2878), .A2(n2879), .ZN(n2839) );
  AND2_X1 U2799 ( .A1(n2836), .A2(n2835), .ZN(n2879) );
  AND2_X1 U2800 ( .A1(n2833), .A2(n2880), .ZN(n2878) );
  OR2_X1 U2801 ( .A1(n2835), .A2(n2836), .ZN(n2880) );
  OR2_X1 U2802 ( .A1(n2255), .A2(n2277), .ZN(n2836) );
  OR2_X1 U2803 ( .A1(n2881), .A2(n2882), .ZN(n2835) );
  AND2_X1 U2804 ( .A1(n2832), .A2(n2831), .ZN(n2882) );
  AND2_X1 U2805 ( .A1(n2829), .A2(n2883), .ZN(n2881) );
  OR2_X1 U2806 ( .A1(n2831), .A2(n2832), .ZN(n2883) );
  OR2_X1 U2807 ( .A1(n2277), .A2(n2259), .ZN(n2832) );
  OR2_X1 U2808 ( .A1(n2884), .A2(n2885), .ZN(n2831) );
  AND2_X1 U2809 ( .A1(n2828), .A2(n2827), .ZN(n2885) );
  AND2_X1 U2810 ( .A1(n2825), .A2(n2886), .ZN(n2884) );
  OR2_X1 U2811 ( .A1(n2827), .A2(n2828), .ZN(n2886) );
  OR2_X1 U2812 ( .A1(n2264), .A2(n2277), .ZN(n2828) );
  OR2_X1 U2813 ( .A1(n2887), .A2(n2888), .ZN(n2827) );
  AND2_X1 U2814 ( .A1(n2824), .A2(n2823), .ZN(n2888) );
  AND2_X1 U2815 ( .A1(n2821), .A2(n2889), .ZN(n2887) );
  OR2_X1 U2816 ( .A1(n2823), .A2(n2824), .ZN(n2889) );
  OR2_X1 U2817 ( .A1(n2277), .A2(n2268), .ZN(n2824) );
  OR2_X1 U2818 ( .A1(n2890), .A2(n2891), .ZN(n2823) );
  AND2_X1 U2819 ( .A1(n2820), .A2(n2819), .ZN(n2891) );
  AND2_X1 U2820 ( .A1(n2817), .A2(n2892), .ZN(n2890) );
  OR2_X1 U2821 ( .A1(n2819), .A2(n2820), .ZN(n2892) );
  OR2_X1 U2822 ( .A1(n2277), .A2(n2273), .ZN(n2820) );
  OR2_X1 U2823 ( .A1(n2893), .A2(n2894), .ZN(n2819) );
  AND2_X1 U2824 ( .A1(n2278), .A2(n2816), .ZN(n2894) );
  AND2_X1 U2825 ( .A1(n2814), .A2(n2895), .ZN(n2893) );
  OR2_X1 U2826 ( .A1(n2816), .A2(n2278), .ZN(n2895) );
  INV_X1 U2827 ( .A(n2062), .ZN(n2278) );
  AND2_X1 U2828 ( .A1(a_12_), .A2(b_12_), .ZN(n2062) );
  OR2_X1 U2829 ( .A1(n2896), .A2(n2897), .ZN(n2816) );
  AND2_X1 U2830 ( .A1(n2810), .A2(n2813), .ZN(n2897) );
  AND2_X1 U2831 ( .A1(n2812), .A2(n2898), .ZN(n2896) );
  OR2_X1 U2832 ( .A1(n2813), .A2(n2810), .ZN(n2898) );
  OR2_X1 U2833 ( .A1(n2281), .A2(n2277), .ZN(n2810) );
  OR3_X1 U2834 ( .A1(n2277), .A2(n2274), .A3(n2596), .ZN(n2813) );
  INV_X1 U2835 ( .A(n2899), .ZN(n2812) );
  OR2_X1 U2836 ( .A1(n2900), .A2(n2901), .ZN(n2899) );
  AND2_X1 U2837 ( .A1(b_11_), .A2(n2902), .ZN(n2901) );
  OR2_X1 U2838 ( .A1(n2903), .A2(n2029), .ZN(n2902) );
  AND2_X1 U2839 ( .A1(a_14_), .A2(n2269), .ZN(n2903) );
  AND2_X1 U2840 ( .A1(b_10_), .A2(n2904), .ZN(n2900) );
  OR2_X1 U2841 ( .A1(n2905), .A2(n2031), .ZN(n2904) );
  AND2_X1 U2842 ( .A1(a_15_), .A2(n2274), .ZN(n2905) );
  XNOR2_X1 U2843 ( .A(n2906), .B(n2907), .ZN(n2814) );
  XNOR2_X1 U2844 ( .A(n2908), .B(n2909), .ZN(n2907) );
  XOR2_X1 U2845 ( .A(n2910), .B(n2911), .Z(n2817) );
  XOR2_X1 U2846 ( .A(n2912), .B(n2913), .Z(n2911) );
  XOR2_X1 U2847 ( .A(n2914), .B(n2915), .Z(n2821) );
  XOR2_X1 U2848 ( .A(n2916), .B(n2079), .Z(n2915) );
  XOR2_X1 U2849 ( .A(n2917), .B(n2918), .Z(n2825) );
  XOR2_X1 U2850 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR2_X1 U2851 ( .A(n2921), .B(n2922), .Z(n2829) );
  XOR2_X1 U2852 ( .A(n2923), .B(n2924), .Z(n2922) );
  XOR2_X1 U2853 ( .A(n2925), .B(n2926), .Z(n2833) );
  XOR2_X1 U2854 ( .A(n2927), .B(n2928), .Z(n2926) );
  XOR2_X1 U2855 ( .A(n2929), .B(n2930), .Z(n2837) );
  XOR2_X1 U2856 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR2_X1 U2857 ( .A(n2933), .B(n2934), .Z(n2841) );
  XOR2_X1 U2858 ( .A(n2935), .B(n2936), .Z(n2934) );
  XOR2_X1 U2859 ( .A(n2937), .B(n2938), .Z(n2845) );
  XOR2_X1 U2860 ( .A(n2939), .B(n2940), .Z(n2938) );
  XOR2_X1 U2861 ( .A(n2941), .B(n2942), .Z(n2849) );
  XOR2_X1 U2862 ( .A(n2943), .B(n2944), .Z(n2942) );
  XOR2_X1 U2863 ( .A(n2945), .B(n2946), .Z(n2853) );
  XOR2_X1 U2864 ( .A(n2947), .B(n2948), .Z(n2946) );
  XOR2_X1 U2865 ( .A(n2949), .B(n2950), .Z(n2668) );
  XOR2_X1 U2866 ( .A(n2951), .B(n2952), .Z(n2950) );
  XOR2_X1 U2867 ( .A(n2953), .B(n2954), .Z(n2549) );
  XOR2_X1 U2868 ( .A(n2955), .B(n2956), .Z(n2954) );
  XNOR2_X1 U2869 ( .A(n2957), .B(n2958), .ZN(n2323) );
  XOR2_X1 U2870 ( .A(n2959), .B(n2960), .Z(n2958) );
  XNOR2_X1 U2871 ( .A(n2333), .B(n2533), .ZN(n2321) );
  OR2_X1 U2872 ( .A1(n2961), .A2(n2962), .ZN(n2533) );
  AND2_X1 U2873 ( .A1(n2960), .A2(n2959), .ZN(n2962) );
  AND2_X1 U2874 ( .A1(n2957), .A2(n2963), .ZN(n2961) );
  OR2_X1 U2875 ( .A1(n2959), .A2(n2960), .ZN(n2963) );
  OR2_X1 U2876 ( .A1(n2274), .A2(n2364), .ZN(n2960) );
  OR2_X1 U2877 ( .A1(n2964), .A2(n2965), .ZN(n2959) );
  AND2_X1 U2878 ( .A1(n2956), .A2(n2955), .ZN(n2965) );
  AND2_X1 U2879 ( .A1(n2953), .A2(n2966), .ZN(n2964) );
  OR2_X1 U2880 ( .A1(n2955), .A2(n2956), .ZN(n2966) );
  OR2_X1 U2881 ( .A1(n2274), .A2(n2228), .ZN(n2956) );
  OR2_X1 U2882 ( .A1(n2967), .A2(n2968), .ZN(n2955) );
  AND2_X1 U2883 ( .A1(n2952), .A2(n2951), .ZN(n2968) );
  AND2_X1 U2884 ( .A1(n2949), .A2(n2969), .ZN(n2967) );
  OR2_X1 U2885 ( .A1(n2951), .A2(n2952), .ZN(n2969) );
  OR2_X1 U2886 ( .A1(n2274), .A2(n2232), .ZN(n2952) );
  OR2_X1 U2887 ( .A1(n2970), .A2(n2971), .ZN(n2951) );
  AND2_X1 U2888 ( .A1(n2948), .A2(n2947), .ZN(n2971) );
  AND2_X1 U2889 ( .A1(n2945), .A2(n2972), .ZN(n2970) );
  OR2_X1 U2890 ( .A1(n2947), .A2(n2948), .ZN(n2972) );
  OR2_X1 U2891 ( .A1(n2237), .A2(n2274), .ZN(n2948) );
  OR2_X1 U2892 ( .A1(n2973), .A2(n2974), .ZN(n2947) );
  AND2_X1 U2893 ( .A1(n2944), .A2(n2943), .ZN(n2974) );
  AND2_X1 U2894 ( .A1(n2941), .A2(n2975), .ZN(n2973) );
  OR2_X1 U2895 ( .A1(n2943), .A2(n2944), .ZN(n2975) );
  OR2_X1 U2896 ( .A1(n2274), .A2(n2241), .ZN(n2944) );
  OR2_X1 U2897 ( .A1(n2976), .A2(n2977), .ZN(n2943) );
  AND2_X1 U2898 ( .A1(n2940), .A2(n2939), .ZN(n2977) );
  AND2_X1 U2899 ( .A1(n2937), .A2(n2978), .ZN(n2976) );
  OR2_X1 U2900 ( .A1(n2939), .A2(n2940), .ZN(n2978) );
  OR2_X1 U2901 ( .A1(n2246), .A2(n2274), .ZN(n2940) );
  OR2_X1 U2902 ( .A1(n2979), .A2(n2980), .ZN(n2939) );
  AND2_X1 U2903 ( .A1(n2936), .A2(n2935), .ZN(n2980) );
  AND2_X1 U2904 ( .A1(n2933), .A2(n2981), .ZN(n2979) );
  OR2_X1 U2905 ( .A1(n2935), .A2(n2936), .ZN(n2981) );
  OR2_X1 U2906 ( .A1(n2274), .A2(n2250), .ZN(n2936) );
  OR2_X1 U2907 ( .A1(n2982), .A2(n2983), .ZN(n2935) );
  AND2_X1 U2908 ( .A1(n2932), .A2(n2931), .ZN(n2983) );
  AND2_X1 U2909 ( .A1(n2929), .A2(n2984), .ZN(n2982) );
  OR2_X1 U2910 ( .A1(n2931), .A2(n2932), .ZN(n2984) );
  OR2_X1 U2911 ( .A1(n2255), .A2(n2274), .ZN(n2932) );
  OR2_X1 U2912 ( .A1(n2985), .A2(n2986), .ZN(n2931) );
  AND2_X1 U2913 ( .A1(n2928), .A2(n2927), .ZN(n2986) );
  AND2_X1 U2914 ( .A1(n2925), .A2(n2987), .ZN(n2985) );
  OR2_X1 U2915 ( .A1(n2927), .A2(n2928), .ZN(n2987) );
  OR2_X1 U2916 ( .A1(n2274), .A2(n2259), .ZN(n2928) );
  OR2_X1 U2917 ( .A1(n2988), .A2(n2989), .ZN(n2927) );
  AND2_X1 U2918 ( .A1(n2924), .A2(n2923), .ZN(n2989) );
  AND2_X1 U2919 ( .A1(n2921), .A2(n2990), .ZN(n2988) );
  OR2_X1 U2920 ( .A1(n2923), .A2(n2924), .ZN(n2990) );
  OR2_X1 U2921 ( .A1(n2264), .A2(n2274), .ZN(n2924) );
  OR2_X1 U2922 ( .A1(n2991), .A2(n2992), .ZN(n2923) );
  AND2_X1 U2923 ( .A1(n2920), .A2(n2919), .ZN(n2992) );
  AND2_X1 U2924 ( .A1(n2917), .A2(n2993), .ZN(n2991) );
  OR2_X1 U2925 ( .A1(n2919), .A2(n2920), .ZN(n2993) );
  OR2_X1 U2926 ( .A1(n2274), .A2(n2268), .ZN(n2920) );
  OR2_X1 U2927 ( .A1(n2994), .A2(n2995), .ZN(n2919) );
  AND2_X1 U2928 ( .A1(n2079), .A2(n2916), .ZN(n2995) );
  AND2_X1 U2929 ( .A1(n2914), .A2(n2996), .ZN(n2994) );
  OR2_X1 U2930 ( .A1(n2916), .A2(n2079), .ZN(n2996) );
  OR2_X1 U2931 ( .A1(n2274), .A2(n2273), .ZN(n2079) );
  OR2_X1 U2932 ( .A1(n2997), .A2(n2998), .ZN(n2916) );
  AND2_X1 U2933 ( .A1(n2913), .A2(n2912), .ZN(n2998) );
  AND2_X1 U2934 ( .A1(n2910), .A2(n2999), .ZN(n2997) );
  OR2_X1 U2935 ( .A1(n2912), .A2(n2913), .ZN(n2999) );
  OR2_X1 U2936 ( .A1(n2276), .A2(n2274), .ZN(n2913) );
  OR2_X1 U2937 ( .A1(n3000), .A2(n3001), .ZN(n2912) );
  AND2_X1 U2938 ( .A1(n2906), .A2(n2909), .ZN(n3001) );
  AND2_X1 U2939 ( .A1(n2908), .A2(n3002), .ZN(n3000) );
  OR2_X1 U2940 ( .A1(n2909), .A2(n2906), .ZN(n3002) );
  OR2_X1 U2941 ( .A1(n2281), .A2(n2274), .ZN(n2906) );
  OR3_X1 U2942 ( .A1(n2274), .A2(n2269), .A3(n2596), .ZN(n2909) );
  INV_X1 U2943 ( .A(n3003), .ZN(n2908) );
  OR2_X1 U2944 ( .A1(n3004), .A2(n3005), .ZN(n3003) );
  AND2_X1 U2945 ( .A1(b_9_), .A2(n3006), .ZN(n3005) );
  OR2_X1 U2946 ( .A1(n3007), .A2(n2031), .ZN(n3006) );
  AND2_X1 U2947 ( .A1(a_15_), .A2(n2269), .ZN(n3007) );
  AND2_X1 U2948 ( .A1(b_10_), .A2(n3008), .ZN(n3004) );
  OR2_X1 U2949 ( .A1(n3009), .A2(n2029), .ZN(n3008) );
  AND2_X1 U2950 ( .A1(a_14_), .A2(n2265), .ZN(n3009) );
  XNOR2_X1 U2951 ( .A(n3010), .B(n3011), .ZN(n2910) );
  XNOR2_X1 U2952 ( .A(n3012), .B(n3013), .ZN(n3011) );
  XOR2_X1 U2953 ( .A(n3014), .B(n3015), .Z(n2914) );
  XOR2_X1 U2954 ( .A(n3016), .B(n3017), .Z(n3015) );
  XOR2_X1 U2955 ( .A(n3018), .B(n3019), .Z(n2917) );
  XOR2_X1 U2956 ( .A(n3020), .B(n3021), .Z(n3019) );
  XOR2_X1 U2957 ( .A(n3022), .B(n3023), .Z(n2921) );
  XNOR2_X1 U2958 ( .A(n3024), .B(n2091), .ZN(n3023) );
  XOR2_X1 U2959 ( .A(n3025), .B(n3026), .Z(n2925) );
  XOR2_X1 U2960 ( .A(n3027), .B(n3028), .Z(n3026) );
  XOR2_X1 U2961 ( .A(n3029), .B(n3030), .Z(n2929) );
  XOR2_X1 U2962 ( .A(n3031), .B(n3032), .Z(n3030) );
  XOR2_X1 U2963 ( .A(n3033), .B(n3034), .Z(n2933) );
  XOR2_X1 U2964 ( .A(n3035), .B(n3036), .Z(n3034) );
  XOR2_X1 U2965 ( .A(n3037), .B(n3038), .Z(n2937) );
  XOR2_X1 U2966 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR2_X1 U2967 ( .A(n3041), .B(n3042), .Z(n2941) );
  XOR2_X1 U2968 ( .A(n3043), .B(n3044), .Z(n3042) );
  XOR2_X1 U2969 ( .A(n3045), .B(n3046), .Z(n2945) );
  XOR2_X1 U2970 ( .A(n3047), .B(n3048), .Z(n3046) );
  XOR2_X1 U2971 ( .A(n3049), .B(n3050), .Z(n2949) );
  XOR2_X1 U2972 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR2_X1 U2973 ( .A(n3053), .B(n3054), .Z(n2953) );
  XOR2_X1 U2974 ( .A(n3055), .B(n3056), .Z(n3054) );
  XOR2_X1 U2975 ( .A(n3057), .B(n3058), .Z(n2957) );
  XOR2_X1 U2976 ( .A(n3059), .B(n3060), .Z(n3058) );
  XNOR2_X1 U2977 ( .A(n3061), .B(n3062), .ZN(n2333) );
  XOR2_X1 U2978 ( .A(n3063), .B(n3064), .Z(n3062) );
  XNOR2_X1 U2979 ( .A(n1971), .B(n2531), .ZN(n2331) );
  OR2_X1 U2980 ( .A1(n3065), .A2(n3066), .ZN(n2531) );
  AND2_X1 U2981 ( .A1(n3064), .A2(n3063), .ZN(n3066) );
  AND2_X1 U2982 ( .A1(n3061), .A2(n3067), .ZN(n3065) );
  OR2_X1 U2983 ( .A1(n3063), .A2(n3064), .ZN(n3067) );
  OR2_X1 U2984 ( .A1(n2269), .A2(n2364), .ZN(n3064) );
  OR2_X1 U2985 ( .A1(n3068), .A2(n3069), .ZN(n3063) );
  AND2_X1 U2986 ( .A1(n3060), .A2(n3059), .ZN(n3069) );
  AND2_X1 U2987 ( .A1(n3057), .A2(n3070), .ZN(n3068) );
  OR2_X1 U2988 ( .A1(n3059), .A2(n3060), .ZN(n3070) );
  OR2_X1 U2989 ( .A1(n2269), .A2(n2228), .ZN(n3060) );
  OR2_X1 U2990 ( .A1(n3071), .A2(n3072), .ZN(n3059) );
  AND2_X1 U2991 ( .A1(n3056), .A2(n3055), .ZN(n3072) );
  AND2_X1 U2992 ( .A1(n3053), .A2(n3073), .ZN(n3071) );
  OR2_X1 U2993 ( .A1(n3055), .A2(n3056), .ZN(n3073) );
  OR2_X1 U2994 ( .A1(n2269), .A2(n2232), .ZN(n3056) );
  OR2_X1 U2995 ( .A1(n3074), .A2(n3075), .ZN(n3055) );
  AND2_X1 U2996 ( .A1(n3049), .A2(n3052), .ZN(n3075) );
  AND2_X1 U2997 ( .A1(n3076), .A2(n3051), .ZN(n3074) );
  OR2_X1 U2998 ( .A1(n3077), .A2(n3078), .ZN(n3051) );
  AND2_X1 U2999 ( .A1(n3048), .A2(n3047), .ZN(n3078) );
  AND2_X1 U3000 ( .A1(n3045), .A2(n3079), .ZN(n3077) );
  OR2_X1 U3001 ( .A1(n3047), .A2(n3048), .ZN(n3079) );
  OR2_X1 U3002 ( .A1(n2269), .A2(n2241), .ZN(n3048) );
  OR2_X1 U3003 ( .A1(n3080), .A2(n3081), .ZN(n3047) );
  AND2_X1 U3004 ( .A1(n3041), .A2(n3044), .ZN(n3081) );
  AND2_X1 U3005 ( .A1(n3082), .A2(n3043), .ZN(n3080) );
  OR2_X1 U3006 ( .A1(n3083), .A2(n3084), .ZN(n3043) );
  AND2_X1 U3007 ( .A1(n3037), .A2(n3040), .ZN(n3084) );
  AND2_X1 U3008 ( .A1(n3085), .A2(n3039), .ZN(n3083) );
  OR2_X1 U3009 ( .A1(n3086), .A2(n3087), .ZN(n3039) );
  AND2_X1 U3010 ( .A1(n3033), .A2(n3036), .ZN(n3087) );
  AND2_X1 U3011 ( .A1(n3088), .A2(n3035), .ZN(n3086) );
  OR2_X1 U3012 ( .A1(n3089), .A2(n3090), .ZN(n3035) );
  AND2_X1 U3013 ( .A1(n3029), .A2(n3032), .ZN(n3090) );
  AND2_X1 U3014 ( .A1(n3091), .A2(n3031), .ZN(n3089) );
  OR2_X1 U3015 ( .A1(n3092), .A2(n3093), .ZN(n3031) );
  AND2_X1 U3016 ( .A1(n3025), .A2(n3028), .ZN(n3093) );
  AND2_X1 U3017 ( .A1(n3094), .A2(n3027), .ZN(n3092) );
  OR2_X1 U3018 ( .A1(n3095), .A2(n3096), .ZN(n3027) );
  AND2_X1 U3019 ( .A1(n3022), .A2(n2270), .ZN(n3096) );
  AND2_X1 U3020 ( .A1(n3097), .A2(n3024), .ZN(n3095) );
  OR2_X1 U3021 ( .A1(n3098), .A2(n3099), .ZN(n3024) );
  AND2_X1 U3022 ( .A1(n3018), .A2(n3021), .ZN(n3099) );
  AND2_X1 U3023 ( .A1(n3100), .A2(n3020), .ZN(n3098) );
  OR2_X1 U3024 ( .A1(n3101), .A2(n3102), .ZN(n3020) );
  AND2_X1 U3025 ( .A1(n3014), .A2(n3017), .ZN(n3102) );
  AND2_X1 U3026 ( .A1(n3103), .A2(n3016), .ZN(n3101) );
  OR2_X1 U3027 ( .A1(n3104), .A2(n3105), .ZN(n3016) );
  AND2_X1 U3028 ( .A1(n3010), .A2(n3013), .ZN(n3105) );
  AND2_X1 U3029 ( .A1(n3012), .A2(n3106), .ZN(n3104) );
  OR2_X1 U3030 ( .A1(n3013), .A2(n3010), .ZN(n3106) );
  OR2_X1 U3031 ( .A1(n2281), .A2(n2269), .ZN(n3010) );
  OR3_X1 U3032 ( .A1(n2265), .A2(n2269), .A3(n2596), .ZN(n3013) );
  INV_X1 U3033 ( .A(n3107), .ZN(n3012) );
  OR2_X1 U3034 ( .A1(n3108), .A2(n3109), .ZN(n3107) );
  AND2_X1 U3035 ( .A1(b_9_), .A2(n3110), .ZN(n3109) );
  OR2_X1 U3036 ( .A1(n3111), .A2(n2029), .ZN(n3110) );
  AND2_X1 U3037 ( .A1(a_14_), .A2(n2260), .ZN(n3111) );
  AND2_X1 U3038 ( .A1(b_8_), .A2(n3112), .ZN(n3108) );
  OR2_X1 U3039 ( .A1(n3113), .A2(n2031), .ZN(n3112) );
  AND2_X1 U3040 ( .A1(a_15_), .A2(n2265), .ZN(n3113) );
  OR2_X1 U3041 ( .A1(n3017), .A2(n3014), .ZN(n3103) );
  XNOR2_X1 U3042 ( .A(n3114), .B(n3115), .ZN(n3014) );
  XNOR2_X1 U3043 ( .A(n3116), .B(n3117), .ZN(n3115) );
  OR2_X1 U3044 ( .A1(n2276), .A2(n2269), .ZN(n3017) );
  OR2_X1 U3045 ( .A1(n3021), .A2(n3018), .ZN(n3100) );
  XOR2_X1 U3046 ( .A(n3118), .B(n3119), .Z(n3018) );
  XOR2_X1 U3047 ( .A(n3120), .B(n3121), .Z(n3119) );
  OR2_X1 U3048 ( .A1(n2273), .A2(n2269), .ZN(n3021) );
  OR2_X1 U3049 ( .A1(n2270), .A2(n3022), .ZN(n3097) );
  XOR2_X1 U3050 ( .A(n3122), .B(n3123), .Z(n3022) );
  XOR2_X1 U3051 ( .A(n3124), .B(n3125), .Z(n3123) );
  INV_X1 U3052 ( .A(n2091), .ZN(n2270) );
  AND2_X1 U3053 ( .A1(a_10_), .A2(b_10_), .ZN(n2091) );
  OR2_X1 U3054 ( .A1(n3028), .A2(n3025), .ZN(n3094) );
  XOR2_X1 U3055 ( .A(n3126), .B(n3127), .Z(n3025) );
  XOR2_X1 U3056 ( .A(n3128), .B(n3129), .Z(n3127) );
  OR2_X1 U3057 ( .A1(n2264), .A2(n2269), .ZN(n3028) );
  OR2_X1 U3058 ( .A1(n3032), .A2(n3029), .ZN(n3091) );
  XOR2_X1 U3059 ( .A(n3130), .B(n3131), .Z(n3029) );
  XOR2_X1 U3060 ( .A(n3132), .B(n2266), .Z(n3131) );
  OR2_X1 U3061 ( .A1(n2269), .A2(n2259), .ZN(n3032) );
  OR2_X1 U3062 ( .A1(n3036), .A2(n3033), .ZN(n3088) );
  XOR2_X1 U3063 ( .A(n3133), .B(n3134), .Z(n3033) );
  XOR2_X1 U3064 ( .A(n3135), .B(n3136), .Z(n3134) );
  OR2_X1 U3065 ( .A1(n2255), .A2(n2269), .ZN(n3036) );
  OR2_X1 U3066 ( .A1(n3040), .A2(n3037), .ZN(n3085) );
  XOR2_X1 U3067 ( .A(n3137), .B(n3138), .Z(n3037) );
  XOR2_X1 U3068 ( .A(n3139), .B(n3140), .Z(n3138) );
  OR2_X1 U3069 ( .A1(n2269), .A2(n2250), .ZN(n3040) );
  OR2_X1 U3070 ( .A1(n3044), .A2(n3041), .ZN(n3082) );
  XOR2_X1 U3071 ( .A(n3141), .B(n3142), .Z(n3041) );
  XOR2_X1 U3072 ( .A(n3143), .B(n3144), .Z(n3142) );
  OR2_X1 U3073 ( .A1(n2246), .A2(n2269), .ZN(n3044) );
  XOR2_X1 U3074 ( .A(n3145), .B(n3146), .Z(n3045) );
  XOR2_X1 U3075 ( .A(n3147), .B(n3148), .Z(n3146) );
  OR2_X1 U3076 ( .A1(n3052), .A2(n3049), .ZN(n3076) );
  XOR2_X1 U3077 ( .A(n3149), .B(n3150), .Z(n3049) );
  XOR2_X1 U3078 ( .A(n3151), .B(n3152), .Z(n3150) );
  OR2_X1 U3079 ( .A1(n2237), .A2(n2269), .ZN(n3052) );
  XOR2_X1 U3080 ( .A(n3153), .B(n3154), .Z(n3053) );
  XOR2_X1 U3081 ( .A(n3155), .B(n3156), .Z(n3154) );
  XOR2_X1 U3082 ( .A(n3157), .B(n3158), .Z(n3057) );
  XOR2_X1 U3083 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR2_X1 U3084 ( .A(n3161), .B(n3162), .Z(n3061) );
  XOR2_X1 U3085 ( .A(n3163), .B(n3164), .Z(n3162) );
  XNOR2_X1 U3086 ( .A(n3165), .B(n3166), .ZN(n1971) );
  XOR2_X1 U3087 ( .A(n3167), .B(n3168), .Z(n3166) );
  INV_X1 U3088 ( .A(n3169), .ZN(n1968) );
  OR2_X1 U3089 ( .A1(n3170), .A2(n2529), .ZN(n3169) );
  INV_X1 U3090 ( .A(n3171), .ZN(n2529) );
  OR2_X1 U3091 ( .A1(n3172), .A2(n3173), .ZN(n3171) );
  AND2_X1 U3092 ( .A1(n3172), .A2(n3173), .ZN(n3170) );
  OR2_X1 U3093 ( .A1(n3174), .A2(n3175), .ZN(n3173) );
  AND2_X1 U3094 ( .A1(n3168), .A2(n3167), .ZN(n3175) );
  AND2_X1 U3095 ( .A1(n3165), .A2(n3176), .ZN(n3174) );
  OR2_X1 U3096 ( .A1(n3167), .A2(n3168), .ZN(n3176) );
  OR2_X1 U3097 ( .A1(n2265), .A2(n2364), .ZN(n3168) );
  OR2_X1 U3098 ( .A1(n3177), .A2(n3178), .ZN(n3167) );
  AND2_X1 U3099 ( .A1(n3164), .A2(n3163), .ZN(n3178) );
  AND2_X1 U3100 ( .A1(n3161), .A2(n3179), .ZN(n3177) );
  OR2_X1 U3101 ( .A1(n3163), .A2(n3164), .ZN(n3179) );
  OR2_X1 U3102 ( .A1(n2265), .A2(n2228), .ZN(n3164) );
  OR2_X1 U3103 ( .A1(n3180), .A2(n3181), .ZN(n3163) );
  AND2_X1 U3104 ( .A1(n3160), .A2(n3159), .ZN(n3181) );
  AND2_X1 U3105 ( .A1(n3157), .A2(n3182), .ZN(n3180) );
  OR2_X1 U3106 ( .A1(n3159), .A2(n3160), .ZN(n3182) );
  OR2_X1 U3107 ( .A1(n2265), .A2(n2232), .ZN(n3160) );
  OR2_X1 U3108 ( .A1(n3183), .A2(n3184), .ZN(n3159) );
  AND2_X1 U3109 ( .A1(n3156), .A2(n3155), .ZN(n3184) );
  AND2_X1 U3110 ( .A1(n3153), .A2(n3185), .ZN(n3183) );
  OR2_X1 U3111 ( .A1(n3155), .A2(n3156), .ZN(n3185) );
  OR2_X1 U3112 ( .A1(n2237), .A2(n2265), .ZN(n3156) );
  OR2_X1 U3113 ( .A1(n3186), .A2(n3187), .ZN(n3155) );
  AND2_X1 U3114 ( .A1(n3149), .A2(n3152), .ZN(n3187) );
  AND2_X1 U3115 ( .A1(n3188), .A2(n3151), .ZN(n3186) );
  OR2_X1 U3116 ( .A1(n3189), .A2(n3190), .ZN(n3151) );
  AND2_X1 U3117 ( .A1(n3148), .A2(n3147), .ZN(n3190) );
  AND2_X1 U3118 ( .A1(n3145), .A2(n3191), .ZN(n3189) );
  OR2_X1 U3119 ( .A1(n3147), .A2(n3148), .ZN(n3191) );
  OR2_X1 U3120 ( .A1(n2246), .A2(n2265), .ZN(n3148) );
  OR2_X1 U3121 ( .A1(n3192), .A2(n3193), .ZN(n3147) );
  AND2_X1 U3122 ( .A1(n3141), .A2(n3144), .ZN(n3193) );
  AND2_X1 U3123 ( .A1(n3194), .A2(n3143), .ZN(n3192) );
  OR2_X1 U3124 ( .A1(n3195), .A2(n3196), .ZN(n3143) );
  AND2_X1 U3125 ( .A1(n3137), .A2(n3140), .ZN(n3196) );
  AND2_X1 U3126 ( .A1(n3197), .A2(n3139), .ZN(n3195) );
  OR2_X1 U3127 ( .A1(n3198), .A2(n3199), .ZN(n3139) );
  AND2_X1 U3128 ( .A1(n3133), .A2(n3136), .ZN(n3199) );
  AND2_X1 U3129 ( .A1(n3200), .A2(n3135), .ZN(n3198) );
  OR2_X1 U3130 ( .A1(n3201), .A2(n3202), .ZN(n3135) );
  AND2_X1 U3131 ( .A1(n3130), .A2(n2266), .ZN(n3202) );
  AND2_X1 U3132 ( .A1(n3203), .A2(n3132), .ZN(n3201) );
  OR2_X1 U3133 ( .A1(n3204), .A2(n3205), .ZN(n3132) );
  AND2_X1 U3134 ( .A1(n3126), .A2(n3129), .ZN(n3205) );
  AND2_X1 U3135 ( .A1(n3206), .A2(n3128), .ZN(n3204) );
  OR2_X1 U3136 ( .A1(n3207), .A2(n3208), .ZN(n3128) );
  AND2_X1 U3137 ( .A1(n3122), .A2(n3125), .ZN(n3208) );
  AND2_X1 U3138 ( .A1(n3209), .A2(n3124), .ZN(n3207) );
  OR2_X1 U3139 ( .A1(n3210), .A2(n3211), .ZN(n3124) );
  AND2_X1 U3140 ( .A1(n3118), .A2(n3121), .ZN(n3211) );
  AND2_X1 U3141 ( .A1(n3212), .A2(n3120), .ZN(n3210) );
  OR2_X1 U3142 ( .A1(n3213), .A2(n3214), .ZN(n3120) );
  AND2_X1 U3143 ( .A1(n3114), .A2(n3117), .ZN(n3214) );
  AND2_X1 U3144 ( .A1(n3116), .A2(n3215), .ZN(n3213) );
  OR2_X1 U3145 ( .A1(n3117), .A2(n3114), .ZN(n3215) );
  OR2_X1 U3146 ( .A1(n2281), .A2(n2265), .ZN(n3114) );
  OR3_X1 U3147 ( .A1(n2260), .A2(n2265), .A3(n2596), .ZN(n3117) );
  INV_X1 U3148 ( .A(n3216), .ZN(n3116) );
  OR2_X1 U3149 ( .A1(n3217), .A2(n3218), .ZN(n3216) );
  AND2_X1 U3150 ( .A1(b_8_), .A2(n3219), .ZN(n3218) );
  OR2_X1 U3151 ( .A1(n3220), .A2(n2029), .ZN(n3219) );
  AND2_X1 U3152 ( .A1(a_14_), .A2(n2256), .ZN(n3220) );
  AND2_X1 U3153 ( .A1(b_7_), .A2(n3221), .ZN(n3217) );
  OR2_X1 U3154 ( .A1(n3222), .A2(n2031), .ZN(n3221) );
  AND2_X1 U3155 ( .A1(a_15_), .A2(n2260), .ZN(n3222) );
  OR2_X1 U3156 ( .A1(n3121), .A2(n3118), .ZN(n3212) );
  XNOR2_X1 U3157 ( .A(n3223), .B(n3224), .ZN(n3118) );
  XNOR2_X1 U3158 ( .A(n3225), .B(n3226), .ZN(n3224) );
  OR2_X1 U3159 ( .A1(n2276), .A2(n2265), .ZN(n3121) );
  OR2_X1 U3160 ( .A1(n3125), .A2(n3122), .ZN(n3209) );
  XOR2_X1 U3161 ( .A(n3227), .B(n3228), .Z(n3122) );
  XOR2_X1 U3162 ( .A(n3229), .B(n3230), .Z(n3228) );
  OR2_X1 U3163 ( .A1(n2273), .A2(n2265), .ZN(n3125) );
  OR2_X1 U3164 ( .A1(n3129), .A2(n3126), .ZN(n3206) );
  XOR2_X1 U3165 ( .A(n3231), .B(n3232), .Z(n3126) );
  XOR2_X1 U3166 ( .A(n3233), .B(n3234), .Z(n3232) );
  OR2_X1 U3167 ( .A1(n2268), .A2(n2265), .ZN(n3129) );
  OR2_X1 U3168 ( .A1(n2266), .A2(n3130), .ZN(n3203) );
  XOR2_X1 U3169 ( .A(n3235), .B(n3236), .Z(n3130) );
  XOR2_X1 U3170 ( .A(n3237), .B(n3238), .Z(n3236) );
  OR2_X1 U3171 ( .A1(n2264), .A2(n2265), .ZN(n2266) );
  OR2_X1 U3172 ( .A1(n3136), .A2(n3133), .ZN(n3200) );
  XOR2_X1 U3173 ( .A(n3239), .B(n3240), .Z(n3133) );
  XOR2_X1 U3174 ( .A(n3241), .B(n3242), .Z(n3240) );
  OR2_X1 U3175 ( .A1(n2265), .A2(n2259), .ZN(n3136) );
  OR2_X1 U3176 ( .A1(n3140), .A2(n3137), .ZN(n3197) );
  XNOR2_X1 U3177 ( .A(n3243), .B(n3244), .ZN(n3137) );
  XNOR2_X1 U3178 ( .A(n2261), .B(n3245), .ZN(n3243) );
  OR2_X1 U3179 ( .A1(n2255), .A2(n2265), .ZN(n3140) );
  OR2_X1 U3180 ( .A1(n3144), .A2(n3141), .ZN(n3194) );
  XOR2_X1 U3181 ( .A(n3246), .B(n3247), .Z(n3141) );
  XOR2_X1 U3182 ( .A(n3248), .B(n3249), .Z(n3247) );
  OR2_X1 U3183 ( .A1(n2265), .A2(n2250), .ZN(n3144) );
  XOR2_X1 U3184 ( .A(n3250), .B(n3251), .Z(n3145) );
  XOR2_X1 U3185 ( .A(n3252), .B(n3253), .Z(n3251) );
  OR2_X1 U3186 ( .A1(n3152), .A2(n3149), .ZN(n3188) );
  XOR2_X1 U3187 ( .A(n3254), .B(n3255), .Z(n3149) );
  XOR2_X1 U3188 ( .A(n3256), .B(n3257), .Z(n3255) );
  OR2_X1 U3189 ( .A1(n2265), .A2(n2241), .ZN(n3152) );
  XOR2_X1 U3190 ( .A(n3258), .B(n3259), .Z(n3153) );
  XOR2_X1 U3191 ( .A(n3260), .B(n3261), .Z(n3259) );
  XOR2_X1 U3192 ( .A(n3262), .B(n3263), .Z(n3157) );
  XOR2_X1 U3193 ( .A(n3264), .B(n3265), .Z(n3263) );
  XOR2_X1 U3194 ( .A(n3266), .B(n3267), .Z(n3161) );
  XOR2_X1 U3195 ( .A(n3268), .B(n3269), .Z(n3267) );
  XOR2_X1 U3196 ( .A(n3270), .B(n3271), .Z(n3165) );
  XOR2_X1 U3197 ( .A(n3272), .B(n3273), .Z(n3271) );
  XOR2_X1 U3198 ( .A(n2488), .B(n3274), .Z(n3172) );
  XOR2_X1 U3199 ( .A(n2487), .B(n2486), .Z(n3274) );
  OR2_X1 U3200 ( .A1(n2260), .A2(n2364), .ZN(n2486) );
  OR2_X1 U3201 ( .A1(n3275), .A2(n3276), .ZN(n2487) );
  AND2_X1 U3202 ( .A1(n3273), .A2(n3272), .ZN(n3276) );
  AND2_X1 U3203 ( .A1(n3270), .A2(n3277), .ZN(n3275) );
  OR2_X1 U3204 ( .A1(n3272), .A2(n3273), .ZN(n3277) );
  OR2_X1 U3205 ( .A1(n2260), .A2(n2228), .ZN(n3273) );
  OR2_X1 U3206 ( .A1(n3278), .A2(n3279), .ZN(n3272) );
  AND2_X1 U3207 ( .A1(n3269), .A2(n3268), .ZN(n3279) );
  AND2_X1 U3208 ( .A1(n3266), .A2(n3280), .ZN(n3278) );
  OR2_X1 U3209 ( .A1(n3268), .A2(n3269), .ZN(n3280) );
  OR2_X1 U3210 ( .A1(n2260), .A2(n2232), .ZN(n3269) );
  OR2_X1 U3211 ( .A1(n3281), .A2(n3282), .ZN(n3268) );
  AND2_X1 U3212 ( .A1(n3265), .A2(n3264), .ZN(n3282) );
  AND2_X1 U3213 ( .A1(n3262), .A2(n3283), .ZN(n3281) );
  OR2_X1 U3214 ( .A1(n3264), .A2(n3265), .ZN(n3283) );
  OR2_X1 U3215 ( .A1(n2237), .A2(n2260), .ZN(n3265) );
  OR2_X1 U3216 ( .A1(n3284), .A2(n3285), .ZN(n3264) );
  AND2_X1 U3217 ( .A1(n3261), .A2(n3260), .ZN(n3285) );
  AND2_X1 U3218 ( .A1(n3258), .A2(n3286), .ZN(n3284) );
  OR2_X1 U3219 ( .A1(n3260), .A2(n3261), .ZN(n3286) );
  OR2_X1 U3220 ( .A1(n2260), .A2(n2241), .ZN(n3261) );
  OR2_X1 U3221 ( .A1(n3287), .A2(n3288), .ZN(n3260) );
  AND2_X1 U3222 ( .A1(n3254), .A2(n3257), .ZN(n3288) );
  AND2_X1 U3223 ( .A1(n3289), .A2(n3256), .ZN(n3287) );
  OR2_X1 U3224 ( .A1(n3290), .A2(n3291), .ZN(n3256) );
  AND2_X1 U3225 ( .A1(n3253), .A2(n3252), .ZN(n3291) );
  AND2_X1 U3226 ( .A1(n3250), .A2(n3292), .ZN(n3290) );
  OR2_X1 U3227 ( .A1(n3252), .A2(n3253), .ZN(n3292) );
  OR2_X1 U3228 ( .A1(n2260), .A2(n2250), .ZN(n3253) );
  OR2_X1 U3229 ( .A1(n3293), .A2(n3294), .ZN(n3252) );
  AND2_X1 U3230 ( .A1(n3246), .A2(n3249), .ZN(n3294) );
  AND2_X1 U3231 ( .A1(n3295), .A2(n3248), .ZN(n3293) );
  OR2_X1 U3232 ( .A1(n3296), .A2(n3297), .ZN(n3248) );
  AND2_X1 U3233 ( .A1(n3244), .A2(n2261), .ZN(n3297) );
  AND2_X1 U3234 ( .A1(n3298), .A2(n3245), .ZN(n3296) );
  OR2_X1 U3235 ( .A1(n3299), .A2(n3300), .ZN(n3245) );
  AND2_X1 U3236 ( .A1(n3239), .A2(n3242), .ZN(n3300) );
  AND2_X1 U3237 ( .A1(n3301), .A2(n3241), .ZN(n3299) );
  OR2_X1 U3238 ( .A1(n3302), .A2(n3303), .ZN(n3241) );
  AND2_X1 U3239 ( .A1(n3235), .A2(n3238), .ZN(n3303) );
  AND2_X1 U3240 ( .A1(n3304), .A2(n3237), .ZN(n3302) );
  OR2_X1 U3241 ( .A1(n3305), .A2(n3306), .ZN(n3237) );
  AND2_X1 U3242 ( .A1(n3231), .A2(n3234), .ZN(n3306) );
  AND2_X1 U3243 ( .A1(n3307), .A2(n3233), .ZN(n3305) );
  OR2_X1 U3244 ( .A1(n3308), .A2(n3309), .ZN(n3233) );
  AND2_X1 U3245 ( .A1(n3227), .A2(n3230), .ZN(n3309) );
  AND2_X1 U3246 ( .A1(n3310), .A2(n3229), .ZN(n3308) );
  OR2_X1 U3247 ( .A1(n3311), .A2(n3312), .ZN(n3229) );
  AND2_X1 U3248 ( .A1(n3223), .A2(n3226), .ZN(n3312) );
  AND2_X1 U3249 ( .A1(n3225), .A2(n3313), .ZN(n3311) );
  OR2_X1 U3250 ( .A1(n3226), .A2(n3223), .ZN(n3313) );
  OR2_X1 U3251 ( .A1(n2260), .A2(n2281), .ZN(n3223) );
  OR3_X1 U3252 ( .A1(n2256), .A2(n2260), .A3(n2596), .ZN(n3226) );
  INV_X1 U3253 ( .A(n3314), .ZN(n3225) );
  OR2_X1 U3254 ( .A1(n3315), .A2(n3316), .ZN(n3314) );
  AND2_X1 U3255 ( .A1(b_7_), .A2(n3317), .ZN(n3316) );
  OR2_X1 U3256 ( .A1(n3318), .A2(n2029), .ZN(n3317) );
  AND2_X1 U3257 ( .A1(a_14_), .A2(n2251), .ZN(n3318) );
  AND2_X1 U3258 ( .A1(b_6_), .A2(n3319), .ZN(n3315) );
  OR2_X1 U3259 ( .A1(n3320), .A2(n2031), .ZN(n3319) );
  AND2_X1 U3260 ( .A1(a_15_), .A2(n2256), .ZN(n3320) );
  OR2_X1 U3261 ( .A1(n3230), .A2(n3227), .ZN(n3310) );
  XNOR2_X1 U3262 ( .A(n3321), .B(n3322), .ZN(n3227) );
  XNOR2_X1 U3263 ( .A(n3323), .B(n3324), .ZN(n3322) );
  OR2_X1 U3264 ( .A1(n2260), .A2(n2276), .ZN(n3230) );
  OR2_X1 U3265 ( .A1(n3234), .A2(n3231), .ZN(n3307) );
  XOR2_X1 U3266 ( .A(n3325), .B(n3326), .Z(n3231) );
  XOR2_X1 U3267 ( .A(n3327), .B(n3328), .Z(n3326) );
  OR2_X1 U3268 ( .A1(n2260), .A2(n2273), .ZN(n3234) );
  OR2_X1 U3269 ( .A1(n3238), .A2(n3235), .ZN(n3304) );
  XOR2_X1 U3270 ( .A(n3329), .B(n3330), .Z(n3235) );
  XOR2_X1 U3271 ( .A(n3331), .B(n3332), .Z(n3330) );
  OR2_X1 U3272 ( .A1(n2260), .A2(n2268), .ZN(n3238) );
  OR2_X1 U3273 ( .A1(n3242), .A2(n3239), .ZN(n3301) );
  XOR2_X1 U3274 ( .A(n3333), .B(n3334), .Z(n3239) );
  XOR2_X1 U3275 ( .A(n3335), .B(n3336), .Z(n3334) );
  OR2_X1 U3276 ( .A1(n2260), .A2(n2264), .ZN(n3242) );
  OR2_X1 U3277 ( .A1(n2261), .A2(n3244), .ZN(n3298) );
  XOR2_X1 U3278 ( .A(n3337), .B(n3338), .Z(n3244) );
  XOR2_X1 U3279 ( .A(n3339), .B(n3340), .Z(n3338) );
  INV_X1 U3280 ( .A(n2117), .ZN(n2261) );
  AND2_X1 U3281 ( .A1(b_8_), .A2(a_8_), .ZN(n2117) );
  OR2_X1 U3282 ( .A1(n3249), .A2(n3246), .ZN(n3295) );
  XOR2_X1 U3283 ( .A(n3341), .B(n3342), .Z(n3246) );
  XOR2_X1 U3284 ( .A(n3343), .B(n3344), .Z(n3342) );
  OR2_X1 U3285 ( .A1(n2255), .A2(n2260), .ZN(n3249) );
  XOR2_X1 U3286 ( .A(n3345), .B(n3346), .Z(n3250) );
  XOR2_X1 U3287 ( .A(n3347), .B(n2257), .Z(n3346) );
  OR2_X1 U3288 ( .A1(n3257), .A2(n3254), .ZN(n3289) );
  XOR2_X1 U3289 ( .A(n3348), .B(n3349), .Z(n3254) );
  XOR2_X1 U3290 ( .A(n3350), .B(n3351), .Z(n3349) );
  OR2_X1 U3291 ( .A1(n2246), .A2(n2260), .ZN(n3257) );
  XOR2_X1 U3292 ( .A(n3352), .B(n3353), .Z(n3258) );
  XOR2_X1 U3293 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR2_X1 U3294 ( .A(n3356), .B(n3357), .Z(n3262) );
  XOR2_X1 U3295 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR2_X1 U3296 ( .A(n3360), .B(n3361), .Z(n3266) );
  XOR2_X1 U3297 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR2_X1 U3298 ( .A(n3364), .B(n3365), .Z(n3270) );
  XOR2_X1 U3299 ( .A(n3366), .B(n3367), .Z(n3365) );
  XOR2_X1 U3300 ( .A(n2495), .B(n3368), .Z(n2488) );
  XOR2_X1 U3301 ( .A(n2494), .B(n2493), .Z(n3368) );
  OR2_X1 U3302 ( .A1(n2256), .A2(n2228), .ZN(n2493) );
  OR2_X1 U3303 ( .A1(n3369), .A2(n3370), .ZN(n2494) );
  AND2_X1 U3304 ( .A1(n3367), .A2(n3366), .ZN(n3370) );
  AND2_X1 U3305 ( .A1(n3364), .A2(n3371), .ZN(n3369) );
  OR2_X1 U3306 ( .A1(n3366), .A2(n3367), .ZN(n3371) );
  OR2_X1 U3307 ( .A1(n2256), .A2(n2232), .ZN(n3367) );
  OR2_X1 U3308 ( .A1(n3372), .A2(n3373), .ZN(n3366) );
  AND2_X1 U3309 ( .A1(n3363), .A2(n3362), .ZN(n3373) );
  AND2_X1 U3310 ( .A1(n3360), .A2(n3374), .ZN(n3372) );
  OR2_X1 U3311 ( .A1(n3362), .A2(n3363), .ZN(n3374) );
  OR2_X1 U3312 ( .A1(n2237), .A2(n2256), .ZN(n3363) );
  OR2_X1 U3313 ( .A1(n3375), .A2(n3376), .ZN(n3362) );
  AND2_X1 U3314 ( .A1(n3359), .A2(n3358), .ZN(n3376) );
  AND2_X1 U3315 ( .A1(n3356), .A2(n3377), .ZN(n3375) );
  OR2_X1 U3316 ( .A1(n3358), .A2(n3359), .ZN(n3377) );
  OR2_X1 U3317 ( .A1(n2256), .A2(n2241), .ZN(n3359) );
  OR2_X1 U3318 ( .A1(n3378), .A2(n3379), .ZN(n3358) );
  AND2_X1 U3319 ( .A1(n3355), .A2(n3354), .ZN(n3379) );
  AND2_X1 U3320 ( .A1(n3352), .A2(n3380), .ZN(n3378) );
  OR2_X1 U3321 ( .A1(n3354), .A2(n3355), .ZN(n3380) );
  OR2_X1 U3322 ( .A1(n2246), .A2(n2256), .ZN(n3355) );
  OR2_X1 U3323 ( .A1(n3381), .A2(n3382), .ZN(n3354) );
  AND2_X1 U3324 ( .A1(n3348), .A2(n3351), .ZN(n3382) );
  AND2_X1 U3325 ( .A1(n3383), .A2(n3350), .ZN(n3381) );
  OR2_X1 U3326 ( .A1(n3384), .A2(n3385), .ZN(n3350) );
  AND2_X1 U3327 ( .A1(n2257), .A2(n3347), .ZN(n3385) );
  AND2_X1 U3328 ( .A1(n3345), .A2(n3386), .ZN(n3384) );
  OR2_X1 U3329 ( .A1(n3347), .A2(n2257), .ZN(n3386) );
  OR2_X1 U3330 ( .A1(n2255), .A2(n2256), .ZN(n2257) );
  OR2_X1 U3331 ( .A1(n3387), .A2(n3388), .ZN(n3347) );
  AND2_X1 U3332 ( .A1(n3341), .A2(n3344), .ZN(n3388) );
  AND2_X1 U3333 ( .A1(n3389), .A2(n3343), .ZN(n3387) );
  OR2_X1 U3334 ( .A1(n3390), .A2(n3391), .ZN(n3343) );
  AND2_X1 U3335 ( .A1(n3337), .A2(n3340), .ZN(n3391) );
  AND2_X1 U3336 ( .A1(n3392), .A2(n3339), .ZN(n3390) );
  OR2_X1 U3337 ( .A1(n3393), .A2(n3394), .ZN(n3339) );
  AND2_X1 U3338 ( .A1(n3333), .A2(n3336), .ZN(n3394) );
  AND2_X1 U3339 ( .A1(n3395), .A2(n3335), .ZN(n3393) );
  OR2_X1 U3340 ( .A1(n3396), .A2(n3397), .ZN(n3335) );
  AND2_X1 U3341 ( .A1(n3329), .A2(n3332), .ZN(n3397) );
  AND2_X1 U3342 ( .A1(n3398), .A2(n3331), .ZN(n3396) );
  OR2_X1 U3343 ( .A1(n3399), .A2(n3400), .ZN(n3331) );
  AND2_X1 U3344 ( .A1(n3325), .A2(n3328), .ZN(n3400) );
  AND2_X1 U3345 ( .A1(n3401), .A2(n3327), .ZN(n3399) );
  OR2_X1 U3346 ( .A1(n3402), .A2(n3403), .ZN(n3327) );
  AND2_X1 U3347 ( .A1(n3321), .A2(n3324), .ZN(n3403) );
  AND2_X1 U3348 ( .A1(n3323), .A2(n3404), .ZN(n3402) );
  OR2_X1 U3349 ( .A1(n3324), .A2(n3321), .ZN(n3404) );
  OR2_X1 U3350 ( .A1(n2256), .A2(n2281), .ZN(n3321) );
  OR3_X1 U3351 ( .A1(n2256), .A2(n2251), .A3(n2596), .ZN(n3324) );
  INV_X1 U3352 ( .A(n3405), .ZN(n3323) );
  OR2_X1 U3353 ( .A1(n3406), .A2(n3407), .ZN(n3405) );
  AND2_X1 U3354 ( .A1(b_6_), .A2(n3408), .ZN(n3407) );
  OR2_X1 U3355 ( .A1(n3409), .A2(n2029), .ZN(n3408) );
  AND2_X1 U3356 ( .A1(a_14_), .A2(n2247), .ZN(n3409) );
  AND2_X1 U3357 ( .A1(b_5_), .A2(n3410), .ZN(n3406) );
  OR2_X1 U3358 ( .A1(n3411), .A2(n2031), .ZN(n3410) );
  AND2_X1 U3359 ( .A1(a_15_), .A2(n2251), .ZN(n3411) );
  OR2_X1 U3360 ( .A1(n3328), .A2(n3325), .ZN(n3401) );
  XNOR2_X1 U3361 ( .A(n3412), .B(n3413), .ZN(n3325) );
  XNOR2_X1 U3362 ( .A(n3414), .B(n3415), .ZN(n3413) );
  OR2_X1 U3363 ( .A1(n2256), .A2(n2276), .ZN(n3328) );
  OR2_X1 U3364 ( .A1(n3332), .A2(n3329), .ZN(n3398) );
  XOR2_X1 U3365 ( .A(n3416), .B(n3417), .Z(n3329) );
  XOR2_X1 U3366 ( .A(n3418), .B(n3419), .Z(n3417) );
  OR2_X1 U3367 ( .A1(n2256), .A2(n2273), .ZN(n3332) );
  OR2_X1 U3368 ( .A1(n3336), .A2(n3333), .ZN(n3395) );
  XOR2_X1 U3369 ( .A(n3420), .B(n3421), .Z(n3333) );
  XOR2_X1 U3370 ( .A(n3422), .B(n3423), .Z(n3421) );
  OR2_X1 U3371 ( .A1(n2256), .A2(n2268), .ZN(n3336) );
  OR2_X1 U3372 ( .A1(n3340), .A2(n3337), .ZN(n3392) );
  XOR2_X1 U3373 ( .A(n3424), .B(n3425), .Z(n3337) );
  XOR2_X1 U3374 ( .A(n3426), .B(n3427), .Z(n3425) );
  OR2_X1 U3375 ( .A1(n2256), .A2(n2264), .ZN(n3340) );
  OR2_X1 U3376 ( .A1(n3344), .A2(n3341), .ZN(n3389) );
  XOR2_X1 U3377 ( .A(n3428), .B(n3429), .Z(n3341) );
  XOR2_X1 U3378 ( .A(n3430), .B(n3431), .Z(n3429) );
  OR2_X1 U3379 ( .A1(n2256), .A2(n2259), .ZN(n3344) );
  XOR2_X1 U3380 ( .A(n3432), .B(n3433), .Z(n3345) );
  XOR2_X1 U3381 ( .A(n3434), .B(n3435), .Z(n3433) );
  OR2_X1 U3382 ( .A1(n3351), .A2(n3348), .ZN(n3383) );
  XOR2_X1 U3383 ( .A(n3436), .B(n3437), .Z(n3348) );
  XOR2_X1 U3384 ( .A(n3438), .B(n3439), .Z(n3437) );
  OR2_X1 U3385 ( .A1(n2256), .A2(n2250), .ZN(n3351) );
  XNOR2_X1 U3386 ( .A(n3440), .B(n3441), .ZN(n3352) );
  XNOR2_X1 U3387 ( .A(n2252), .B(n3442), .ZN(n3440) );
  XOR2_X1 U3388 ( .A(n3443), .B(n3444), .Z(n3356) );
  XOR2_X1 U3389 ( .A(n3445), .B(n3446), .Z(n3444) );
  XOR2_X1 U3390 ( .A(n3447), .B(n3448), .Z(n3360) );
  XOR2_X1 U3391 ( .A(n3449), .B(n3450), .Z(n3448) );
  XOR2_X1 U3392 ( .A(n3451), .B(n3452), .Z(n3364) );
  XOR2_X1 U3393 ( .A(n3453), .B(n3454), .Z(n3452) );
  XOR2_X1 U3394 ( .A(n2502), .B(n3455), .Z(n2495) );
  XOR2_X1 U3395 ( .A(n2501), .B(n2500), .Z(n3455) );
  OR2_X1 U3396 ( .A1(n2251), .A2(n2232), .ZN(n2500) );
  OR2_X1 U3397 ( .A1(n3456), .A2(n3457), .ZN(n2501) );
  AND2_X1 U3398 ( .A1(n3454), .A2(n3453), .ZN(n3457) );
  AND2_X1 U3399 ( .A1(n3451), .A2(n3458), .ZN(n3456) );
  OR2_X1 U3400 ( .A1(n3453), .A2(n3454), .ZN(n3458) );
  OR2_X1 U3401 ( .A1(n2237), .A2(n2251), .ZN(n3454) );
  OR2_X1 U3402 ( .A1(n3459), .A2(n3460), .ZN(n3453) );
  AND2_X1 U3403 ( .A1(n3450), .A2(n3449), .ZN(n3460) );
  AND2_X1 U3404 ( .A1(n3447), .A2(n3461), .ZN(n3459) );
  OR2_X1 U3405 ( .A1(n3449), .A2(n3450), .ZN(n3461) );
  OR2_X1 U3406 ( .A1(n2251), .A2(n2241), .ZN(n3450) );
  OR2_X1 U3407 ( .A1(n3462), .A2(n3463), .ZN(n3449) );
  AND2_X1 U3408 ( .A1(n3446), .A2(n3445), .ZN(n3463) );
  AND2_X1 U3409 ( .A1(n3443), .A2(n3464), .ZN(n3462) );
  OR2_X1 U3410 ( .A1(n3445), .A2(n3446), .ZN(n3464) );
  OR2_X1 U3411 ( .A1(n2246), .A2(n2251), .ZN(n3446) );
  OR2_X1 U3412 ( .A1(n3465), .A2(n3466), .ZN(n3445) );
  AND2_X1 U3413 ( .A1(n3442), .A2(n2252), .ZN(n3466) );
  AND2_X1 U3414 ( .A1(n3441), .A2(n3467), .ZN(n3465) );
  OR2_X1 U3415 ( .A1(n2252), .A2(n3442), .ZN(n3467) );
  OR2_X1 U3416 ( .A1(n3468), .A2(n3469), .ZN(n3442) );
  AND2_X1 U3417 ( .A1(n3436), .A2(n3439), .ZN(n3469) );
  AND2_X1 U3418 ( .A1(n3470), .A2(n3438), .ZN(n3468) );
  OR2_X1 U3419 ( .A1(n3471), .A2(n3472), .ZN(n3438) );
  AND2_X1 U3420 ( .A1(n3435), .A2(n3434), .ZN(n3472) );
  AND2_X1 U3421 ( .A1(n3432), .A2(n3473), .ZN(n3471) );
  OR2_X1 U3422 ( .A1(n3434), .A2(n3435), .ZN(n3473) );
  OR2_X1 U3423 ( .A1(n2259), .A2(n2251), .ZN(n3435) );
  OR2_X1 U3424 ( .A1(n3474), .A2(n3475), .ZN(n3434) );
  AND2_X1 U3425 ( .A1(n3428), .A2(n3431), .ZN(n3475) );
  AND2_X1 U3426 ( .A1(n3476), .A2(n3430), .ZN(n3474) );
  OR2_X1 U3427 ( .A1(n3477), .A2(n3478), .ZN(n3430) );
  AND2_X1 U3428 ( .A1(n3424), .A2(n3427), .ZN(n3478) );
  AND2_X1 U3429 ( .A1(n3479), .A2(n3426), .ZN(n3477) );
  OR2_X1 U3430 ( .A1(n3480), .A2(n3481), .ZN(n3426) );
  AND2_X1 U3431 ( .A1(n3420), .A2(n3423), .ZN(n3481) );
  AND2_X1 U3432 ( .A1(n3482), .A2(n3422), .ZN(n3480) );
  OR2_X1 U3433 ( .A1(n3483), .A2(n3484), .ZN(n3422) );
  AND2_X1 U3434 ( .A1(n3416), .A2(n3419), .ZN(n3484) );
  AND2_X1 U3435 ( .A1(n3485), .A2(n3418), .ZN(n3483) );
  OR2_X1 U3436 ( .A1(n3486), .A2(n3487), .ZN(n3418) );
  AND2_X1 U3437 ( .A1(n3412), .A2(n3415), .ZN(n3487) );
  AND2_X1 U3438 ( .A1(n3414), .A2(n3488), .ZN(n3486) );
  OR2_X1 U3439 ( .A1(n3415), .A2(n3412), .ZN(n3488) );
  OR2_X1 U3440 ( .A1(n2281), .A2(n2251), .ZN(n3412) );
  OR3_X1 U3441 ( .A1(n2247), .A2(n2251), .A3(n2596), .ZN(n3415) );
  INV_X1 U3442 ( .A(n3489), .ZN(n3414) );
  OR2_X1 U3443 ( .A1(n3490), .A2(n3491), .ZN(n3489) );
  AND2_X1 U3444 ( .A1(b_5_), .A2(n3492), .ZN(n3491) );
  OR2_X1 U3445 ( .A1(n3493), .A2(n2029), .ZN(n3492) );
  AND2_X1 U3446 ( .A1(a_14_), .A2(n2242), .ZN(n3493) );
  AND2_X1 U3447 ( .A1(b_4_), .A2(n3494), .ZN(n3490) );
  OR2_X1 U3448 ( .A1(n3495), .A2(n2031), .ZN(n3494) );
  AND2_X1 U3449 ( .A1(a_15_), .A2(n2247), .ZN(n3495) );
  OR2_X1 U3450 ( .A1(n3419), .A2(n3416), .ZN(n3485) );
  XNOR2_X1 U3451 ( .A(n3496), .B(n3497), .ZN(n3416) );
  XNOR2_X1 U3452 ( .A(n3498), .B(n3499), .ZN(n3497) );
  OR2_X1 U3453 ( .A1(n2276), .A2(n2251), .ZN(n3419) );
  OR2_X1 U3454 ( .A1(n3423), .A2(n3420), .ZN(n3482) );
  XOR2_X1 U3455 ( .A(n3500), .B(n3501), .Z(n3420) );
  XOR2_X1 U3456 ( .A(n3502), .B(n3503), .Z(n3501) );
  OR2_X1 U3457 ( .A1(n2273), .A2(n2251), .ZN(n3423) );
  OR2_X1 U3458 ( .A1(n3427), .A2(n3424), .ZN(n3479) );
  XOR2_X1 U3459 ( .A(n3504), .B(n3505), .Z(n3424) );
  XOR2_X1 U3460 ( .A(n3506), .B(n3507), .Z(n3505) );
  OR2_X1 U3461 ( .A1(n2268), .A2(n2251), .ZN(n3427) );
  OR2_X1 U3462 ( .A1(n3431), .A2(n3428), .ZN(n3476) );
  XOR2_X1 U3463 ( .A(n3508), .B(n3509), .Z(n3428) );
  XOR2_X1 U3464 ( .A(n3510), .B(n3511), .Z(n3509) );
  OR2_X1 U3465 ( .A1(n2264), .A2(n2251), .ZN(n3431) );
  XOR2_X1 U3466 ( .A(n3512), .B(n3513), .Z(n3432) );
  XOR2_X1 U3467 ( .A(n3514), .B(n3515), .Z(n3513) );
  OR2_X1 U3468 ( .A1(n3439), .A2(n3436), .ZN(n3470) );
  XOR2_X1 U3469 ( .A(n3516), .B(n3517), .Z(n3436) );
  XOR2_X1 U3470 ( .A(n3518), .B(n3519), .Z(n3517) );
  OR2_X1 U3471 ( .A1(n2255), .A2(n2251), .ZN(n3439) );
  INV_X1 U3472 ( .A(n2142), .ZN(n2252) );
  AND2_X1 U3473 ( .A1(a_6_), .A2(b_6_), .ZN(n2142) );
  XOR2_X1 U3474 ( .A(n3520), .B(n3521), .Z(n3441) );
  XOR2_X1 U3475 ( .A(n3522), .B(n3523), .Z(n3521) );
  XOR2_X1 U3476 ( .A(n3524), .B(n3525), .Z(n3443) );
  XOR2_X1 U3477 ( .A(n3526), .B(n3527), .Z(n3525) );
  XOR2_X1 U3478 ( .A(n3528), .B(n3529), .Z(n3447) );
  XOR2_X1 U3479 ( .A(n3530), .B(n2248), .Z(n3529) );
  XOR2_X1 U3480 ( .A(n3531), .B(n3532), .Z(n3451) );
  XOR2_X1 U3481 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR2_X1 U3482 ( .A(n2509), .B(n3535), .Z(n2502) );
  XOR2_X1 U3483 ( .A(n2508), .B(n2507), .Z(n3535) );
  OR2_X1 U3484 ( .A1(n2237), .A2(n2247), .ZN(n2507) );
  OR2_X1 U3485 ( .A1(n3536), .A2(n3537), .ZN(n2508) );
  AND2_X1 U3486 ( .A1(n3534), .A2(n3533), .ZN(n3537) );
  AND2_X1 U3487 ( .A1(n3531), .A2(n3538), .ZN(n3536) );
  OR2_X1 U3488 ( .A1(n3533), .A2(n3534), .ZN(n3538) );
  OR2_X1 U3489 ( .A1(n2247), .A2(n2241), .ZN(n3534) );
  OR2_X1 U3490 ( .A1(n3539), .A2(n3540), .ZN(n3533) );
  AND2_X1 U3491 ( .A1(n2248), .A2(n3530), .ZN(n3540) );
  AND2_X1 U3492 ( .A1(n3528), .A2(n3541), .ZN(n3539) );
  OR2_X1 U3493 ( .A1(n3530), .A2(n2248), .ZN(n3541) );
  OR2_X1 U3494 ( .A1(n2246), .A2(n2247), .ZN(n2248) );
  OR2_X1 U3495 ( .A1(n3542), .A2(n3543), .ZN(n3530) );
  AND2_X1 U3496 ( .A1(n3527), .A2(n3526), .ZN(n3543) );
  AND2_X1 U3497 ( .A1(n3524), .A2(n3544), .ZN(n3542) );
  OR2_X1 U3498 ( .A1(n3526), .A2(n3527), .ZN(n3544) );
  OR2_X1 U3499 ( .A1(n2247), .A2(n2250), .ZN(n3527) );
  OR2_X1 U3500 ( .A1(n3545), .A2(n3546), .ZN(n3526) );
  AND2_X1 U3501 ( .A1(n3523), .A2(n3522), .ZN(n3546) );
  AND2_X1 U3502 ( .A1(n3520), .A2(n3547), .ZN(n3545) );
  OR2_X1 U3503 ( .A1(n3522), .A2(n3523), .ZN(n3547) );
  OR2_X1 U3504 ( .A1(n2247), .A2(n2255), .ZN(n3523) );
  OR2_X1 U3505 ( .A1(n3548), .A2(n3549), .ZN(n3522) );
  AND2_X1 U3506 ( .A1(n3516), .A2(n3519), .ZN(n3549) );
  AND2_X1 U3507 ( .A1(n3550), .A2(n3518), .ZN(n3548) );
  OR2_X1 U3508 ( .A1(n3551), .A2(n3552), .ZN(n3518) );
  AND2_X1 U3509 ( .A1(n3515), .A2(n3514), .ZN(n3552) );
  AND2_X1 U3510 ( .A1(n3512), .A2(n3553), .ZN(n3551) );
  OR2_X1 U3511 ( .A1(n3514), .A2(n3515), .ZN(n3553) );
  OR2_X1 U3512 ( .A1(n2247), .A2(n2264), .ZN(n3515) );
  OR2_X1 U3513 ( .A1(n3554), .A2(n3555), .ZN(n3514) );
  AND2_X1 U3514 ( .A1(n3508), .A2(n3511), .ZN(n3555) );
  AND2_X1 U3515 ( .A1(n3556), .A2(n3510), .ZN(n3554) );
  OR2_X1 U3516 ( .A1(n3557), .A2(n3558), .ZN(n3510) );
  AND2_X1 U3517 ( .A1(n3504), .A2(n3507), .ZN(n3558) );
  AND2_X1 U3518 ( .A1(n3559), .A2(n3506), .ZN(n3557) );
  OR2_X1 U3519 ( .A1(n3560), .A2(n3561), .ZN(n3506) );
  AND2_X1 U3520 ( .A1(n3500), .A2(n3503), .ZN(n3561) );
  AND2_X1 U3521 ( .A1(n3562), .A2(n3502), .ZN(n3560) );
  OR2_X1 U3522 ( .A1(n3563), .A2(n3564), .ZN(n3502) );
  AND2_X1 U3523 ( .A1(n3496), .A2(n3499), .ZN(n3564) );
  AND2_X1 U3524 ( .A1(n3498), .A2(n3565), .ZN(n3563) );
  OR2_X1 U3525 ( .A1(n3499), .A2(n3496), .ZN(n3565) );
  OR2_X1 U3526 ( .A1(n2247), .A2(n2281), .ZN(n3496) );
  OR3_X1 U3527 ( .A1(n2242), .A2(n2247), .A3(n2596), .ZN(n3499) );
  INV_X1 U3528 ( .A(n3566), .ZN(n3498) );
  OR2_X1 U3529 ( .A1(n3567), .A2(n3568), .ZN(n3566) );
  AND2_X1 U3530 ( .A1(b_4_), .A2(n3569), .ZN(n3568) );
  OR2_X1 U3531 ( .A1(n3570), .A2(n2029), .ZN(n3569) );
  AND2_X1 U3532 ( .A1(a_14_), .A2(n2238), .ZN(n3570) );
  AND2_X1 U3533 ( .A1(b_3_), .A2(n3571), .ZN(n3567) );
  OR2_X1 U3534 ( .A1(n3572), .A2(n2031), .ZN(n3571) );
  AND2_X1 U3535 ( .A1(a_15_), .A2(n2242), .ZN(n3572) );
  OR2_X1 U3536 ( .A1(n3503), .A2(n3500), .ZN(n3562) );
  XNOR2_X1 U3537 ( .A(n3573), .B(n3574), .ZN(n3500) );
  XNOR2_X1 U3538 ( .A(n3575), .B(n3576), .ZN(n3574) );
  OR2_X1 U3539 ( .A1(n2247), .A2(n2276), .ZN(n3503) );
  OR2_X1 U3540 ( .A1(n3507), .A2(n3504), .ZN(n3559) );
  XOR2_X1 U3541 ( .A(n3577), .B(n3578), .Z(n3504) );
  XOR2_X1 U3542 ( .A(n3579), .B(n3580), .Z(n3578) );
  OR2_X1 U3543 ( .A1(n2247), .A2(n2273), .ZN(n3507) );
  OR2_X1 U3544 ( .A1(n3511), .A2(n3508), .ZN(n3556) );
  XOR2_X1 U3545 ( .A(n3581), .B(n3582), .Z(n3508) );
  XOR2_X1 U3546 ( .A(n3583), .B(n3584), .Z(n3582) );
  OR2_X1 U3547 ( .A1(n2247), .A2(n2268), .ZN(n3511) );
  XOR2_X1 U3548 ( .A(n3585), .B(n3586), .Z(n3512) );
  XOR2_X1 U3549 ( .A(n3587), .B(n3588), .Z(n3586) );
  OR2_X1 U3550 ( .A1(n3519), .A2(n3516), .ZN(n3550) );
  XOR2_X1 U3551 ( .A(n3589), .B(n3590), .Z(n3516) );
  XOR2_X1 U3552 ( .A(n3591), .B(n3592), .Z(n3590) );
  OR2_X1 U3553 ( .A1(n2247), .A2(n2259), .ZN(n3519) );
  XOR2_X1 U3554 ( .A(n3593), .B(n3594), .Z(n3520) );
  XOR2_X1 U3555 ( .A(n3595), .B(n3596), .Z(n3594) );
  XOR2_X1 U3556 ( .A(n3597), .B(n3598), .Z(n3524) );
  XOR2_X1 U3557 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR2_X1 U3558 ( .A(n3601), .B(n3602), .Z(n3528) );
  XOR2_X1 U3559 ( .A(n3603), .B(n3604), .Z(n3602) );
  XOR2_X1 U3560 ( .A(n3605), .B(n3606), .Z(n3531) );
  XOR2_X1 U3561 ( .A(n3607), .B(n3608), .Z(n3606) );
  XNOR2_X1 U3562 ( .A(n3609), .B(n2515), .ZN(n2509) );
  XOR2_X1 U3563 ( .A(n2522), .B(n3610), .Z(n2515) );
  XOR2_X1 U3564 ( .A(n2521), .B(n2520), .Z(n3610) );
  OR2_X1 U3565 ( .A1(n2238), .A2(n2246), .ZN(n2520) );
  OR2_X1 U3566 ( .A1(n3611), .A2(n3612), .ZN(n2521) );
  AND2_X1 U3567 ( .A1(n3613), .A2(n3614), .ZN(n3612) );
  AND2_X1 U3568 ( .A1(n3615), .A2(n3616), .ZN(n3611) );
  OR2_X1 U3569 ( .A1(n3614), .A2(n3613), .ZN(n3616) );
  XOR2_X1 U3570 ( .A(n3617), .B(n3618), .Z(n2522) );
  XOR2_X1 U3571 ( .A(n3619), .B(n3620), .Z(n3618) );
  XNOR2_X1 U3572 ( .A(n2243), .B(n2514), .ZN(n3609) );
  OR2_X1 U3573 ( .A1(n3621), .A2(n3622), .ZN(n2514) );
  AND2_X1 U3574 ( .A1(n3608), .A2(n3607), .ZN(n3622) );
  AND2_X1 U3575 ( .A1(n3605), .A2(n3623), .ZN(n3621) );
  OR2_X1 U3576 ( .A1(n3607), .A2(n3608), .ZN(n3623) );
  OR2_X1 U3577 ( .A1(n2242), .A2(n2246), .ZN(n3608) );
  OR2_X1 U3578 ( .A1(n3624), .A2(n3625), .ZN(n3607) );
  AND2_X1 U3579 ( .A1(n3604), .A2(n3603), .ZN(n3625) );
  AND2_X1 U3580 ( .A1(n3601), .A2(n3626), .ZN(n3624) );
  OR2_X1 U3581 ( .A1(n3603), .A2(n3604), .ZN(n3626) );
  OR2_X1 U3582 ( .A1(n2242), .A2(n2250), .ZN(n3604) );
  OR2_X1 U3583 ( .A1(n3627), .A2(n3628), .ZN(n3603) );
  AND2_X1 U3584 ( .A1(n3600), .A2(n3599), .ZN(n3628) );
  AND2_X1 U3585 ( .A1(n3597), .A2(n3629), .ZN(n3627) );
  OR2_X1 U3586 ( .A1(n3599), .A2(n3600), .ZN(n3629) );
  OR2_X1 U3587 ( .A1(n2242), .A2(n2255), .ZN(n3600) );
  OR2_X1 U3588 ( .A1(n3630), .A2(n3631), .ZN(n3599) );
  AND2_X1 U3589 ( .A1(n3596), .A2(n3595), .ZN(n3631) );
  AND2_X1 U3590 ( .A1(n3593), .A2(n3632), .ZN(n3630) );
  OR2_X1 U3591 ( .A1(n3595), .A2(n3596), .ZN(n3632) );
  OR2_X1 U3592 ( .A1(n2242), .A2(n2259), .ZN(n3596) );
  OR2_X1 U3593 ( .A1(n3633), .A2(n3634), .ZN(n3595) );
  AND2_X1 U3594 ( .A1(n3589), .A2(n3592), .ZN(n3634) );
  AND2_X1 U3595 ( .A1(n3635), .A2(n3591), .ZN(n3633) );
  OR2_X1 U3596 ( .A1(n3636), .A2(n3637), .ZN(n3591) );
  AND2_X1 U3597 ( .A1(n3588), .A2(n3587), .ZN(n3637) );
  AND2_X1 U3598 ( .A1(n3585), .A2(n3638), .ZN(n3636) );
  OR2_X1 U3599 ( .A1(n3587), .A2(n3588), .ZN(n3638) );
  OR2_X1 U3600 ( .A1(n2242), .A2(n2268), .ZN(n3588) );
  OR2_X1 U3601 ( .A1(n3639), .A2(n3640), .ZN(n3587) );
  AND2_X1 U3602 ( .A1(n3581), .A2(n3584), .ZN(n3640) );
  AND2_X1 U3603 ( .A1(n3641), .A2(n3583), .ZN(n3639) );
  OR2_X1 U3604 ( .A1(n3642), .A2(n3643), .ZN(n3583) );
  AND2_X1 U3605 ( .A1(n3577), .A2(n3580), .ZN(n3643) );
  AND2_X1 U3606 ( .A1(n3644), .A2(n3579), .ZN(n3642) );
  OR2_X1 U3607 ( .A1(n3645), .A2(n3646), .ZN(n3579) );
  AND2_X1 U3608 ( .A1(n3573), .A2(n3576), .ZN(n3646) );
  AND2_X1 U3609 ( .A1(n3575), .A2(n3647), .ZN(n3645) );
  OR2_X1 U3610 ( .A1(n3576), .A2(n3573), .ZN(n3647) );
  OR2_X1 U3611 ( .A1(n2242), .A2(n2281), .ZN(n3573) );
  OR3_X1 U3612 ( .A1(n2238), .A2(n2242), .A3(n2596), .ZN(n3576) );
  INV_X1 U3613 ( .A(n3648), .ZN(n3575) );
  OR2_X1 U3614 ( .A1(n3649), .A2(n3650), .ZN(n3648) );
  AND2_X1 U3615 ( .A1(b_3_), .A2(n3651), .ZN(n3650) );
  OR2_X1 U3616 ( .A1(n3652), .A2(n2029), .ZN(n3651) );
  AND2_X1 U3617 ( .A1(a_14_), .A2(n2233), .ZN(n3652) );
  AND2_X1 U3618 ( .A1(b_2_), .A2(n3653), .ZN(n3649) );
  OR2_X1 U3619 ( .A1(n3654), .A2(n2031), .ZN(n3653) );
  AND2_X1 U3620 ( .A1(a_15_), .A2(n2238), .ZN(n3654) );
  OR2_X1 U3621 ( .A1(n3580), .A2(n3577), .ZN(n3644) );
  XNOR2_X1 U3622 ( .A(n3655), .B(n3656), .ZN(n3577) );
  XNOR2_X1 U3623 ( .A(n3657), .B(n3658), .ZN(n3656) );
  OR2_X1 U3624 ( .A1(n2242), .A2(n2276), .ZN(n3580) );
  OR2_X1 U3625 ( .A1(n3584), .A2(n3581), .ZN(n3641) );
  XOR2_X1 U3626 ( .A(n3659), .B(n3660), .Z(n3581) );
  XOR2_X1 U3627 ( .A(n3661), .B(n3662), .Z(n3660) );
  OR2_X1 U3628 ( .A1(n2242), .A2(n2273), .ZN(n3584) );
  XOR2_X1 U3629 ( .A(n3663), .B(n3664), .Z(n3585) );
  XOR2_X1 U3630 ( .A(n3665), .B(n3666), .Z(n3664) );
  OR2_X1 U3631 ( .A1(n3592), .A2(n3589), .ZN(n3635) );
  XOR2_X1 U3632 ( .A(n3667), .B(n3668), .Z(n3589) );
  XOR2_X1 U3633 ( .A(n3669), .B(n3670), .Z(n3668) );
  OR2_X1 U3634 ( .A1(n2242), .A2(n2264), .ZN(n3592) );
  XOR2_X1 U3635 ( .A(n3671), .B(n3672), .Z(n3593) );
  XOR2_X1 U3636 ( .A(n3673), .B(n3674), .Z(n3672) );
  XOR2_X1 U3637 ( .A(n3675), .B(n3676), .Z(n3597) );
  XOR2_X1 U3638 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR2_X1 U3639 ( .A(n3679), .B(n3680), .Z(n3601) );
  XOR2_X1 U3640 ( .A(n3681), .B(n3682), .Z(n3680) );
  XOR2_X1 U3641 ( .A(n3615), .B(n3683), .Z(n3605) );
  XOR2_X1 U3642 ( .A(n3614), .B(n3613), .Z(n3683) );
  OR2_X1 U3643 ( .A1(n2238), .A2(n2250), .ZN(n3613) );
  OR2_X1 U3644 ( .A1(n3684), .A2(n3685), .ZN(n3614) );
  AND2_X1 U3645 ( .A1(n3682), .A2(n3681), .ZN(n3685) );
  AND2_X1 U3646 ( .A1(n3679), .A2(n3686), .ZN(n3684) );
  OR2_X1 U3647 ( .A1(n3681), .A2(n3682), .ZN(n3686) );
  OR2_X1 U3648 ( .A1(n2238), .A2(n2255), .ZN(n3682) );
  OR2_X1 U3649 ( .A1(n3687), .A2(n3688), .ZN(n3681) );
  AND2_X1 U3650 ( .A1(n3678), .A2(n3677), .ZN(n3688) );
  AND2_X1 U3651 ( .A1(n3675), .A2(n3689), .ZN(n3687) );
  OR2_X1 U3652 ( .A1(n3677), .A2(n3678), .ZN(n3689) );
  OR2_X1 U3653 ( .A1(n2238), .A2(n2259), .ZN(n3678) );
  OR2_X1 U3654 ( .A1(n3690), .A2(n3691), .ZN(n3677) );
  AND2_X1 U3655 ( .A1(n3674), .A2(n3673), .ZN(n3691) );
  AND2_X1 U3656 ( .A1(n3671), .A2(n3692), .ZN(n3690) );
  OR2_X1 U3657 ( .A1(n3673), .A2(n3674), .ZN(n3692) );
  OR2_X1 U3658 ( .A1(n2238), .A2(n2264), .ZN(n3674) );
  OR2_X1 U3659 ( .A1(n3693), .A2(n3694), .ZN(n3673) );
  AND2_X1 U3660 ( .A1(n3667), .A2(n3670), .ZN(n3694) );
  AND2_X1 U3661 ( .A1(n3695), .A2(n3669), .ZN(n3693) );
  OR2_X1 U3662 ( .A1(n3696), .A2(n3697), .ZN(n3669) );
  AND2_X1 U3663 ( .A1(n3666), .A2(n3665), .ZN(n3697) );
  AND2_X1 U3664 ( .A1(n3663), .A2(n3698), .ZN(n3696) );
  OR2_X1 U3665 ( .A1(n3665), .A2(n3666), .ZN(n3698) );
  OR2_X1 U3666 ( .A1(n2238), .A2(n2273), .ZN(n3666) );
  OR2_X1 U3667 ( .A1(n3699), .A2(n3700), .ZN(n3665) );
  AND2_X1 U3668 ( .A1(n3659), .A2(n3662), .ZN(n3700) );
  AND2_X1 U3669 ( .A1(n3701), .A2(n3661), .ZN(n3699) );
  OR2_X1 U3670 ( .A1(n3702), .A2(n3703), .ZN(n3661) );
  AND2_X1 U3671 ( .A1(n3655), .A2(n3658), .ZN(n3703) );
  AND2_X1 U3672 ( .A1(n3657), .A2(n3704), .ZN(n3702) );
  OR2_X1 U3673 ( .A1(n3658), .A2(n3655), .ZN(n3704) );
  OR2_X1 U3674 ( .A1(n2238), .A2(n2281), .ZN(n3655) );
  OR3_X1 U3675 ( .A1(n2238), .A2(n2233), .A3(n2596), .ZN(n3658) );
  INV_X1 U3676 ( .A(n3705), .ZN(n3657) );
  OR2_X1 U3677 ( .A1(n3706), .A2(n3707), .ZN(n3705) );
  AND2_X1 U3678 ( .A1(b_2_), .A2(n3708), .ZN(n3707) );
  OR2_X1 U3679 ( .A1(n3709), .A2(n2029), .ZN(n3708) );
  AND2_X1 U3680 ( .A1(a_14_), .A2(n2229), .ZN(n3709) );
  AND2_X1 U3681 ( .A1(b_1_), .A2(n3710), .ZN(n3706) );
  OR2_X1 U3682 ( .A1(n3711), .A2(n2031), .ZN(n3710) );
  AND2_X1 U3683 ( .A1(a_15_), .A2(n2233), .ZN(n3711) );
  OR2_X1 U3684 ( .A1(n3662), .A2(n3659), .ZN(n3701) );
  XNOR2_X1 U3685 ( .A(n3712), .B(n3713), .ZN(n3659) );
  XNOR2_X1 U3686 ( .A(n3714), .B(n3715), .ZN(n3713) );
  OR2_X1 U3687 ( .A1(n2238), .A2(n2276), .ZN(n3662) );
  XOR2_X1 U3688 ( .A(n3716), .B(n3717), .Z(n3663) );
  XOR2_X1 U3689 ( .A(n3718), .B(n3719), .Z(n3717) );
  OR2_X1 U3690 ( .A1(n3670), .A2(n3667), .ZN(n3695) );
  XOR2_X1 U3691 ( .A(n3720), .B(n3721), .Z(n3667) );
  XOR2_X1 U3692 ( .A(n3722), .B(n3723), .Z(n3721) );
  OR2_X1 U3693 ( .A1(n2238), .A2(n2268), .ZN(n3670) );
  XOR2_X1 U3694 ( .A(n3724), .B(n3725), .Z(n3671) );
  XOR2_X1 U3695 ( .A(n3726), .B(n3727), .Z(n3725) );
  XOR2_X1 U3696 ( .A(n3728), .B(n3729), .Z(n3675) );
  XOR2_X1 U3697 ( .A(n3730), .B(n3731), .Z(n3729) );
  XOR2_X1 U3698 ( .A(n3732), .B(n3733), .Z(n3679) );
  XOR2_X1 U3699 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR2_X1 U3700 ( .A(n3736), .B(n3737), .Z(n3615) );
  XOR2_X1 U3701 ( .A(n3738), .B(n3739), .Z(n3737) );
  INV_X1 U3702 ( .A(n2167), .ZN(n2243) );
  AND2_X1 U3703 ( .A1(b_4_), .A2(a_4_), .ZN(n2167) );
  AND2_X1 U3704 ( .A1(n3740), .A2(b_0_), .ZN(n2336) );
  AND3_X1 U3705 ( .A1(n2176), .A2(n2175), .A3(n2173), .ZN(n2177) );
  INV_X1 U3706 ( .A(n3741), .ZN(n2173) );
  OR2_X1 U3707 ( .A1(n3740), .A2(n2225), .ZN(n3741) );
  OR3_X1 U3708 ( .A1(n3742), .A2(n3743), .A3(n3744), .ZN(n2175) );
  XOR2_X1 U3709 ( .A(n3740), .B(n3745), .Z(n3744) );
  AND2_X1 U3710 ( .A1(b_0_), .A2(a_1_), .ZN(n3745) );
  AND2_X1 U3711 ( .A1(b_1_), .A2(a_0_), .ZN(n3740) );
  INV_X1 U3712 ( .A(n3746), .ZN(n3743) );
  OR2_X1 U3713 ( .A1(n2355), .A2(n3747), .ZN(n2176) );
  AND2_X1 U3714 ( .A1(n2356), .A2(n2353), .ZN(n3747) );
  XOR2_X1 U3715 ( .A(n3748), .B(n3746), .Z(n2353) );
  OR2_X1 U3716 ( .A1(n3749), .A2(n3750), .ZN(n3746) );
  AND2_X1 U3717 ( .A1(n3751), .A2(n3752), .ZN(n3750) );
  AND2_X1 U3718 ( .A1(n3753), .A2(n3754), .ZN(n3749) );
  OR2_X1 U3719 ( .A1(n3752), .A2(n3751), .ZN(n3753) );
  OR2_X1 U3720 ( .A1(n3755), .A2(n3742), .ZN(n3748) );
  AND3_X1 U3721 ( .A1(a_2_), .A2(b_0_), .A3(n3756), .ZN(n3742) );
  AND2_X1 U3722 ( .A1(n3757), .A2(n2230), .ZN(n3755) );
  INV_X1 U3723 ( .A(n3756), .ZN(n2230) );
  AND2_X1 U3724 ( .A1(b_1_), .A2(a_1_), .ZN(n3756) );
  OR2_X1 U3725 ( .A1(n2232), .A2(n2225), .ZN(n3757) );
  AND2_X1 U3726 ( .A1(b_2_), .A2(a_0_), .ZN(n2356) );
  INV_X1 U3727 ( .A(n3758), .ZN(n2355) );
  OR2_X1 U3728 ( .A1(n3759), .A2(n3760), .ZN(n3758) );
  AND2_X1 U3729 ( .A1(n2374), .A2(n2373), .ZN(n3760) );
  AND2_X1 U3730 ( .A1(n2371), .A2(n3761), .ZN(n3759) );
  OR2_X1 U3731 ( .A1(n2373), .A2(n2374), .ZN(n3761) );
  OR2_X1 U3732 ( .A1(n2233), .A2(n2228), .ZN(n2374) );
  OR2_X1 U3733 ( .A1(n3762), .A2(n3763), .ZN(n2373) );
  AND2_X1 U3734 ( .A1(n2406), .A2(n2234), .ZN(n3763) );
  AND2_X1 U3735 ( .A1(n2405), .A2(n3764), .ZN(n3762) );
  OR2_X1 U3736 ( .A1(n2234), .A2(n2406), .ZN(n3764) );
  OR2_X1 U3737 ( .A1(n3765), .A2(n3766), .ZN(n2406) );
  AND2_X1 U3738 ( .A1(n2436), .A2(n2435), .ZN(n3766) );
  AND2_X1 U3739 ( .A1(n2433), .A2(n3767), .ZN(n3765) );
  OR2_X1 U3740 ( .A1(n2435), .A2(n2436), .ZN(n3767) );
  OR2_X1 U3741 ( .A1(n2237), .A2(n2233), .ZN(n2436) );
  OR2_X1 U3742 ( .A1(n3768), .A2(n3769), .ZN(n2435) );
  AND2_X1 U3743 ( .A1(n2483), .A2(n2482), .ZN(n3769) );
  AND2_X1 U3744 ( .A1(n2480), .A2(n3770), .ZN(n3768) );
  OR2_X1 U3745 ( .A1(n2482), .A2(n2483), .ZN(n3770) );
  OR2_X1 U3746 ( .A1(n2241), .A2(n2233), .ZN(n2483) );
  OR2_X1 U3747 ( .A1(n3771), .A2(n3772), .ZN(n2482) );
  AND2_X1 U3748 ( .A1(n2527), .A2(n2526), .ZN(n3772) );
  AND2_X1 U3749 ( .A1(n2524), .A2(n3773), .ZN(n3771) );
  OR2_X1 U3750 ( .A1(n2526), .A2(n2527), .ZN(n3773) );
  OR2_X1 U3751 ( .A1(n2246), .A2(n2233), .ZN(n2527) );
  OR2_X1 U3752 ( .A1(n3774), .A2(n3775), .ZN(n2526) );
  AND2_X1 U3753 ( .A1(n3620), .A2(n3619), .ZN(n3775) );
  AND2_X1 U3754 ( .A1(n3617), .A2(n3776), .ZN(n3774) );
  OR2_X1 U3755 ( .A1(n3619), .A2(n3620), .ZN(n3776) );
  OR2_X1 U3756 ( .A1(n2250), .A2(n2233), .ZN(n3620) );
  OR2_X1 U3757 ( .A1(n3777), .A2(n3778), .ZN(n3619) );
  AND2_X1 U3758 ( .A1(n3739), .A2(n3738), .ZN(n3778) );
  AND2_X1 U3759 ( .A1(n3736), .A2(n3779), .ZN(n3777) );
  OR2_X1 U3760 ( .A1(n3738), .A2(n3739), .ZN(n3779) );
  OR2_X1 U3761 ( .A1(n2255), .A2(n2233), .ZN(n3739) );
  OR2_X1 U3762 ( .A1(n3780), .A2(n3781), .ZN(n3738) );
  AND2_X1 U3763 ( .A1(n3735), .A2(n3734), .ZN(n3781) );
  AND2_X1 U3764 ( .A1(n3732), .A2(n3782), .ZN(n3780) );
  OR2_X1 U3765 ( .A1(n3734), .A2(n3735), .ZN(n3782) );
  OR2_X1 U3766 ( .A1(n2259), .A2(n2233), .ZN(n3735) );
  OR2_X1 U3767 ( .A1(n3783), .A2(n3784), .ZN(n3734) );
  AND2_X1 U3768 ( .A1(n3731), .A2(n3730), .ZN(n3784) );
  AND2_X1 U3769 ( .A1(n3728), .A2(n3785), .ZN(n3783) );
  OR2_X1 U3770 ( .A1(n3730), .A2(n3731), .ZN(n3785) );
  OR2_X1 U3771 ( .A1(n2264), .A2(n2233), .ZN(n3731) );
  OR2_X1 U3772 ( .A1(n3786), .A2(n3787), .ZN(n3730) );
  AND2_X1 U3773 ( .A1(n3727), .A2(n3726), .ZN(n3787) );
  AND2_X1 U3774 ( .A1(n3724), .A2(n3788), .ZN(n3786) );
  OR2_X1 U3775 ( .A1(n3726), .A2(n3727), .ZN(n3788) );
  OR2_X1 U3776 ( .A1(n2268), .A2(n2233), .ZN(n3727) );
  OR2_X1 U3777 ( .A1(n3789), .A2(n3790), .ZN(n3726) );
  AND2_X1 U3778 ( .A1(n3720), .A2(n3723), .ZN(n3790) );
  AND2_X1 U3779 ( .A1(n3791), .A2(n3722), .ZN(n3789) );
  OR2_X1 U3780 ( .A1(n3792), .A2(n3793), .ZN(n3722) );
  AND2_X1 U3781 ( .A1(n3719), .A2(n3718), .ZN(n3793) );
  AND2_X1 U3782 ( .A1(n3716), .A2(n3794), .ZN(n3792) );
  OR2_X1 U3783 ( .A1(n3718), .A2(n3719), .ZN(n3794) );
  OR2_X1 U3784 ( .A1(n2276), .A2(n2233), .ZN(n3719) );
  OR2_X1 U3785 ( .A1(n3795), .A2(n3796), .ZN(n3718) );
  AND2_X1 U3786 ( .A1(n3712), .A2(n3715), .ZN(n3796) );
  AND2_X1 U3787 ( .A1(n3714), .A2(n3797), .ZN(n3795) );
  OR2_X1 U3788 ( .A1(n3715), .A2(n3712), .ZN(n3797) );
  OR2_X1 U3789 ( .A1(n2281), .A2(n2233), .ZN(n3712) );
  OR3_X1 U3790 ( .A1(n2229), .A2(n2233), .A3(n2596), .ZN(n3715) );
  INV_X1 U3791 ( .A(n3798), .ZN(n3714) );
  OR2_X1 U3792 ( .A1(n3799), .A2(n3800), .ZN(n3798) );
  AND2_X1 U3793 ( .A1(b_1_), .A2(n3801), .ZN(n3800) );
  OR2_X1 U3794 ( .A1(n3802), .A2(n2029), .ZN(n3801) );
  AND2_X1 U3795 ( .A1(n2017), .A2(a_14_), .ZN(n2029) );
  INV_X1 U3796 ( .A(a_15_), .ZN(n2017) );
  AND2_X1 U3797 ( .A1(a_14_), .A2(n2225), .ZN(n3802) );
  AND2_X1 U3798 ( .A1(b_0_), .A2(n3803), .ZN(n3799) );
  OR2_X1 U3799 ( .A1(n3804), .A2(n2031), .ZN(n3803) );
  AND2_X1 U3800 ( .A1(n3805), .A2(a_15_), .ZN(n2031) );
  AND2_X1 U3801 ( .A1(a_15_), .A2(n2229), .ZN(n3804) );
  XNOR2_X1 U3802 ( .A(n3806), .B(n3807), .ZN(n3716) );
  OR2_X1 U3803 ( .A1(n3808), .A2(n3809), .ZN(n3806) );
  INV_X1 U3804 ( .A(n3810), .ZN(n3809) );
  AND2_X1 U3805 ( .A1(n3811), .A2(n3812), .ZN(n3808) );
  OR2_X1 U3806 ( .A1(n3805), .A2(n2225), .ZN(n3811) );
  OR2_X1 U3807 ( .A1(n3723), .A2(n3720), .ZN(n3791) );
  XOR2_X1 U3808 ( .A(n3813), .B(n3814), .Z(n3720) );
  XOR2_X1 U3809 ( .A(n3815), .B(n3816), .Z(n3813) );
  OR2_X1 U3810 ( .A1(n2273), .A2(n2233), .ZN(n3723) );
  XNOR2_X1 U3811 ( .A(n3817), .B(n3818), .ZN(n3724) );
  XNOR2_X1 U3812 ( .A(n3819), .B(n3820), .ZN(n3817) );
  XNOR2_X1 U3813 ( .A(n3821), .B(n3822), .ZN(n3728) );
  XNOR2_X1 U3814 ( .A(n3823), .B(n3824), .ZN(n3821) );
  XNOR2_X1 U3815 ( .A(n3825), .B(n3826), .ZN(n3732) );
  XNOR2_X1 U3816 ( .A(n3827), .B(n3828), .ZN(n3825) );
  XOR2_X1 U3817 ( .A(n3829), .B(n3830), .Z(n3736) );
  XOR2_X1 U3818 ( .A(n3831), .B(n3832), .Z(n3830) );
  XOR2_X1 U3819 ( .A(n3833), .B(n3834), .Z(n3617) );
  XOR2_X1 U3820 ( .A(n3835), .B(n3836), .Z(n3834) );
  XOR2_X1 U3821 ( .A(n3837), .B(n3838), .Z(n2524) );
  XOR2_X1 U3822 ( .A(n3839), .B(n3840), .Z(n3838) );
  XOR2_X1 U3823 ( .A(n3841), .B(n3842), .Z(n2480) );
  XOR2_X1 U3824 ( .A(n3843), .B(n3844), .Z(n3842) );
  XOR2_X1 U3825 ( .A(n3845), .B(n3846), .Z(n2433) );
  XOR2_X1 U3826 ( .A(n3847), .B(n3848), .Z(n3846) );
  INV_X1 U3827 ( .A(n2202), .ZN(n2234) );
  AND2_X1 U3828 ( .A1(a_2_), .A2(b_2_), .ZN(n2202) );
  XOR2_X1 U3829 ( .A(n3849), .B(n3850), .Z(n2405) );
  XOR2_X1 U3830 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR2_X1 U3831 ( .A(n3751), .B(n3853), .Z(n2371) );
  XOR2_X1 U3832 ( .A(n3752), .B(n3754), .Z(n3853) );
  OR2_X1 U3833 ( .A1(n2237), .A2(n2225), .ZN(n3754) );
  OR2_X1 U3834 ( .A1(n3854), .A2(n3855), .ZN(n3752) );
  AND2_X1 U3835 ( .A1(n3849), .A2(n3851), .ZN(n3855) );
  AND2_X1 U3836 ( .A1(n3856), .A2(n3852), .ZN(n3854) );
  OR2_X1 U3837 ( .A1(n2241), .A2(n2225), .ZN(n3852) );
  OR2_X1 U3838 ( .A1(n3851), .A2(n3849), .ZN(n3856) );
  OR2_X1 U3839 ( .A1(n2229), .A2(n2237), .ZN(n3849) );
  INV_X1 U3840 ( .A(a_3_), .ZN(n2237) );
  OR2_X1 U3841 ( .A1(n3857), .A2(n3858), .ZN(n3851) );
  AND2_X1 U3842 ( .A1(n3845), .A2(n3847), .ZN(n3858) );
  AND2_X1 U3843 ( .A1(n3859), .A2(n3848), .ZN(n3857) );
  OR2_X1 U3844 ( .A1(n2246), .A2(n2225), .ZN(n3848) );
  OR2_X1 U3845 ( .A1(n3847), .A2(n3845), .ZN(n3859) );
  OR2_X1 U3846 ( .A1(n2229), .A2(n2241), .ZN(n3845) );
  INV_X1 U3847 ( .A(a_4_), .ZN(n2241) );
  OR2_X1 U3848 ( .A1(n3860), .A2(n3861), .ZN(n3847) );
  AND2_X1 U3849 ( .A1(n3841), .A2(n3843), .ZN(n3861) );
  AND2_X1 U3850 ( .A1(n3862), .A2(n3844), .ZN(n3860) );
  OR2_X1 U3851 ( .A1(n2250), .A2(n2225), .ZN(n3844) );
  OR2_X1 U3852 ( .A1(n3843), .A2(n3841), .ZN(n3862) );
  OR2_X1 U3853 ( .A1(n2229), .A2(n2246), .ZN(n3841) );
  INV_X1 U3854 ( .A(a_5_), .ZN(n2246) );
  OR2_X1 U3855 ( .A1(n3863), .A2(n3864), .ZN(n3843) );
  AND2_X1 U3856 ( .A1(n3837), .A2(n3839), .ZN(n3864) );
  AND2_X1 U3857 ( .A1(n3865), .A2(n3840), .ZN(n3863) );
  OR2_X1 U3858 ( .A1(n2255), .A2(n2225), .ZN(n3840) );
  OR2_X1 U3859 ( .A1(n3839), .A2(n3837), .ZN(n3865) );
  OR2_X1 U3860 ( .A1(n2229), .A2(n2250), .ZN(n3837) );
  INV_X1 U3861 ( .A(a_6_), .ZN(n2250) );
  OR2_X1 U3862 ( .A1(n3866), .A2(n3867), .ZN(n3839) );
  AND2_X1 U3863 ( .A1(n3833), .A2(n3835), .ZN(n3867) );
  AND2_X1 U3864 ( .A1(n3868), .A2(n3836), .ZN(n3866) );
  OR2_X1 U3865 ( .A1(n2259), .A2(n2225), .ZN(n3836) );
  OR2_X1 U3866 ( .A1(n3835), .A2(n3833), .ZN(n3868) );
  OR2_X1 U3867 ( .A1(n2229), .A2(n2255), .ZN(n3833) );
  INV_X1 U3868 ( .A(a_7_), .ZN(n2255) );
  OR2_X1 U3869 ( .A1(n3869), .A2(n3870), .ZN(n3835) );
  AND2_X1 U3870 ( .A1(n3829), .A2(n3831), .ZN(n3870) );
  AND2_X1 U3871 ( .A1(n3871), .A2(n3832), .ZN(n3869) );
  OR2_X1 U3872 ( .A1(n2264), .A2(n2225), .ZN(n3832) );
  OR2_X1 U3873 ( .A1(n3831), .A2(n3829), .ZN(n3871) );
  OR2_X1 U3874 ( .A1(n2229), .A2(n2259), .ZN(n3829) );
  INV_X1 U3875 ( .A(a_8_), .ZN(n2259) );
  OR2_X1 U3876 ( .A1(n3872), .A2(n3873), .ZN(n3831) );
  AND2_X1 U3877 ( .A1(n3826), .A2(n3828), .ZN(n3873) );
  AND2_X1 U3878 ( .A1(n3874), .A2(n3827), .ZN(n3872) );
  OR2_X1 U3879 ( .A1(n2268), .A2(n2225), .ZN(n3827) );
  OR2_X1 U3880 ( .A1(n3828), .A2(n3826), .ZN(n3874) );
  OR2_X1 U3881 ( .A1(n2229), .A2(n2264), .ZN(n3826) );
  INV_X1 U3882 ( .A(a_9_), .ZN(n2264) );
  OR2_X1 U3883 ( .A1(n3875), .A2(n3876), .ZN(n3828) );
  AND2_X1 U3884 ( .A1(n3822), .A2(n3824), .ZN(n3876) );
  AND2_X1 U3885 ( .A1(n3877), .A2(n3823), .ZN(n3875) );
  OR2_X1 U3886 ( .A1(n2273), .A2(n2225), .ZN(n3823) );
  OR2_X1 U3887 ( .A1(n3824), .A2(n3822), .ZN(n3877) );
  OR2_X1 U3888 ( .A1(n2229), .A2(n2268), .ZN(n3822) );
  INV_X1 U3889 ( .A(a_10_), .ZN(n2268) );
  OR2_X1 U3890 ( .A1(n3878), .A2(n3879), .ZN(n3824) );
  AND2_X1 U3891 ( .A1(n3818), .A2(n3820), .ZN(n3879) );
  AND2_X1 U3892 ( .A1(n3880), .A2(n3819), .ZN(n3878) );
  OR2_X1 U3893 ( .A1(n2276), .A2(n2225), .ZN(n3819) );
  OR2_X1 U3894 ( .A1(n3820), .A2(n3818), .ZN(n3880) );
  OR2_X1 U3895 ( .A1(n2229), .A2(n2273), .ZN(n3818) );
  INV_X1 U3896 ( .A(a_11_), .ZN(n2273) );
  OR2_X1 U3897 ( .A1(n3881), .A2(n3882), .ZN(n3820) );
  AND2_X1 U3898 ( .A1(n3814), .A2(n3816), .ZN(n3882) );
  AND2_X1 U3899 ( .A1(n3815), .A2(n3883), .ZN(n3881) );
  OR2_X1 U3900 ( .A1(n3816), .A2(n3814), .ZN(n3883) );
  OR2_X1 U3901 ( .A1(n2229), .A2(n2276), .ZN(n3814) );
  INV_X1 U3902 ( .A(a_12_), .ZN(n2276) );
  OR2_X1 U3903 ( .A1(n2281), .A2(n2225), .ZN(n3816) );
  AND2_X1 U3904 ( .A1(n3810), .A2(n3807), .ZN(n3815) );
  OR3_X1 U3905 ( .A1(n2229), .A2(n2225), .A3(n2596), .ZN(n3807) );
  INV_X1 U3906 ( .A(n2288), .ZN(n2596) );
  OR3_X1 U3907 ( .A1(n3805), .A2(n2225), .A3(n3812), .ZN(n3810) );
  OR2_X1 U3908 ( .A1(n2229), .A2(n2281), .ZN(n3812) );
  INV_X1 U3909 ( .A(a_13_), .ZN(n2281) );
  INV_X1 U3910 ( .A(b_0_), .ZN(n2225) );
  INV_X1 U3911 ( .A(a_14_), .ZN(n3805) );
  OR2_X1 U3912 ( .A1(n2229), .A2(n2232), .ZN(n3751) );
  INV_X1 U3913 ( .A(a_2_), .ZN(n2232) );
  INV_X1 U3914 ( .A(n2015), .ZN(n1963) );
  OR2_X1 U3915 ( .A1(n3884), .A2(n3885), .ZN(n2015) );
  AND2_X1 U3916 ( .A1(n3886), .A2(n2364), .ZN(n3885) );
  AND2_X1 U3917 ( .A1(b_0_), .A2(n3887), .ZN(n3884) );
  OR2_X1 U3918 ( .A1(n3886), .A2(n2364), .ZN(n3887) );
  INV_X1 U3919 ( .A(a_0_), .ZN(n2364) );
  AND2_X1 U3920 ( .A1(n3888), .A2(n2214), .ZN(n3886) );
  OR2_X1 U3921 ( .A1(b_1_), .A2(n2228), .ZN(n2214) );
  INV_X1 U3922 ( .A(a_1_), .ZN(n2228) );
  INV_X1 U3923 ( .A(n3889), .ZN(n3888) );
  AND3_X1 U3924 ( .A1(n3890), .A2(n2213), .A3(n3891), .ZN(n3889) );
  OR2_X1 U3925 ( .A1(a_2_), .A2(n2233), .ZN(n3891) );
  OR2_X1 U3926 ( .A1(a_1_), .A2(n2229), .ZN(n2213) );
  INV_X1 U3927 ( .A(b_1_), .ZN(n2229) );
  OR3_X1 U3928 ( .A1(n2190), .A2(n3892), .A3(n3893), .ZN(n3890) );
  AND2_X1 U3929 ( .A1(a_2_), .A2(n2233), .ZN(n3893) );
  INV_X1 U3930 ( .A(b_2_), .ZN(n2233) );
  AND3_X1 U3931 ( .A1(n3894), .A2(n2188), .A3(n3895), .ZN(n3892) );
  OR3_X1 U3932 ( .A1(n2155), .A2(n3896), .A3(n3897), .ZN(n3895) );
  AND2_X1 U3933 ( .A1(a_4_), .A2(n2242), .ZN(n3897) );
  AND3_X1 U3934 ( .A1(n3898), .A2(n2153), .A3(n3899), .ZN(n3896) );
  OR2_X1 U3935 ( .A1(a_6_), .A2(n2251), .ZN(n3899) );
  OR2_X1 U3936 ( .A1(a_5_), .A2(n2247), .ZN(n2153) );
  OR3_X1 U3937 ( .A1(n2130), .A2(n3900), .A3(n3901), .ZN(n3898) );
  AND2_X1 U3938 ( .A1(a_6_), .A2(n2251), .ZN(n3901) );
  INV_X1 U3939 ( .A(b_6_), .ZN(n2251) );
  AND3_X1 U3940 ( .A1(n3902), .A2(n2128), .A3(n3903), .ZN(n3900) );
  OR3_X1 U3941 ( .A1(n2105), .A2(n3904), .A3(n3905), .ZN(n3903) );
  AND2_X1 U3942 ( .A1(a_8_), .A2(n2260), .ZN(n3905) );
  AND3_X1 U3943 ( .A1(n2103), .A2(n3906), .A3(n3907), .ZN(n3904) );
  OR2_X1 U3944 ( .A1(a_10_), .A2(n2269), .ZN(n3907) );
  OR3_X1 U3945 ( .A1(n3908), .A2(n3909), .A3(n3910), .ZN(n3906) );
  AND2_X1 U3946 ( .A1(a_11_), .A2(n2274), .ZN(n3910) );
  AND2_X1 U3947 ( .A1(a_10_), .A2(n2269), .ZN(n3909) );
  INV_X1 U3948 ( .A(b_10_), .ZN(n2269) );
  AND3_X1 U3949 ( .A1(n3911), .A2(n3912), .A3(n2080), .ZN(n3908) );
  OR2_X1 U3950 ( .A1(a_11_), .A2(n2274), .ZN(n2080) );
  INV_X1 U3951 ( .A(b_11_), .ZN(n2274) );
  OR3_X1 U3952 ( .A1(n3913), .A2(n3914), .A3(n3915), .ZN(n3912) );
  AND2_X1 U3953 ( .A1(a_13_), .A2(n2282), .ZN(n3915) );
  AND2_X1 U3954 ( .A1(a_12_), .A2(n2277), .ZN(n3914) );
  AND4_X1 U3955 ( .A1(n2049), .A2(n2287), .A3(n3916), .A4(n3917), .ZN(n3913)
         );
  OR2_X1 U3956 ( .A1(n2288), .A2(n2023), .ZN(n3917) );
  AND2_X1 U3957 ( .A1(a_14_), .A2(a_15_), .ZN(n2288) );
  OR2_X1 U3958 ( .A1(n2014), .A2(a_14_), .ZN(n3916) );
  AND2_X1 U3959 ( .A1(n2595), .A2(a_15_), .ZN(n2014) );
  OR2_X1 U3960 ( .A1(n2023), .A2(n2595), .ZN(n2287) );
  INV_X1 U3961 ( .A(b_15_), .ZN(n2595) );
  INV_X1 U3962 ( .A(b_14_), .ZN(n2023) );
  OR2_X1 U3963 ( .A1(a_13_), .A2(n2282), .ZN(n2049) );
  INV_X1 U3964 ( .A(b_13_), .ZN(n2282) );
  OR2_X1 U3965 ( .A1(a_12_), .A2(n2277), .ZN(n3911) );
  INV_X1 U3966 ( .A(b_12_), .ZN(n2277) );
  OR2_X1 U3967 ( .A1(a_9_), .A2(n2265), .ZN(n2103) );
  AND2_X1 U3968 ( .A1(n2265), .A2(a_9_), .ZN(n2105) );
  INV_X1 U3969 ( .A(b_9_), .ZN(n2265) );
  OR2_X1 U3970 ( .A1(a_7_), .A2(n2256), .ZN(n2128) );
  OR2_X1 U3971 ( .A1(a_8_), .A2(n2260), .ZN(n3902) );
  INV_X1 U3972 ( .A(b_8_), .ZN(n2260) );
  AND2_X1 U3973 ( .A1(n2256), .A2(a_7_), .ZN(n2130) );
  INV_X1 U3974 ( .A(b_7_), .ZN(n2256) );
  AND2_X1 U3975 ( .A1(n2247), .A2(a_5_), .ZN(n2155) );
  INV_X1 U3976 ( .A(b_5_), .ZN(n2247) );
  OR2_X1 U3977 ( .A1(a_3_), .A2(n2238), .ZN(n2188) );
  OR2_X1 U3978 ( .A1(a_4_), .A2(n2242), .ZN(n3894) );
  INV_X1 U3979 ( .A(b_4_), .ZN(n2242) );
  AND2_X1 U3980 ( .A1(n2238), .A2(a_3_), .ZN(n2190) );
  INV_X1 U3981 ( .A(b_3_), .ZN(n2238) );
endmodule

