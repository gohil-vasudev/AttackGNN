module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n595_, new_n614_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n442_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n580_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n301_, new_n169_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n177_, new_n493_, new_n547_, new_n264_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n459_, new_n555_, new_n174_, new_n468_, new_n354_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n417_, new_n591_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n550_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n607_, new_n327_, new_n495_, new_n196_, new_n574_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n195_, new_n576_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n406_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

xnor g000 ( new_n138_, N65, N69 );
xnor g001 ( new_n139_, new_n138_, keyIn_0_5 );
xnor g002 ( new_n140_, N73, N77 );
xnor g003 ( new_n141_, new_n140_, keyIn_0_6 );
xnor g004 ( new_n142_, new_n139_, new_n141_ );
xor g005 ( new_n143_, N81, N85 );
xnor g006 ( new_n144_, N89, N93 );
xnor g007 ( new_n145_, new_n143_, new_n144_ );
xnor g008 ( new_n146_, new_n142_, new_n145_ );
nand g009 ( new_n147_, N129, N137 );
xor g010 ( new_n148_, new_n146_, new_n147_ );
xor g011 ( new_n149_, N1, N17 );
xnor g012 ( new_n150_, N33, N49 );
xnor g013 ( new_n151_, new_n149_, new_n150_ );
not g014 ( new_n152_, new_n151_ );
xnor g015 ( new_n153_, new_n148_, new_n152_ );
not g016 ( new_n154_, keyIn_0_36 );
not g017 ( new_n155_, keyIn_0_23 );
xnor g018 ( new_n156_, N121, N125 );
xnor g019 ( new_n157_, new_n156_, keyIn_0_7 );
xor g020 ( new_n158_, N113, N117 );
xnor g021 ( new_n159_, new_n157_, new_n158_ );
xnor g022 ( new_n160_, new_n159_, keyIn_0_19 );
xnor g023 ( new_n161_, new_n160_, new_n145_ );
nand g024 ( new_n162_, N132, N137 );
xor g025 ( new_n163_, new_n162_, keyIn_0_9 );
xnor g026 ( new_n164_, new_n161_, new_n163_ );
xnor g027 ( new_n165_, new_n164_, new_n155_ );
xnor g028 ( new_n166_, N13, N29 );
xnor g029 ( new_n167_, new_n166_, keyIn_0_14 );
xnor g030 ( new_n168_, N45, N61 );
xnor g031 ( new_n169_, new_n167_, new_n168_ );
xnor g032 ( new_n170_, new_n165_, new_n169_ );
xnor g033 ( new_n171_, N5, N21 );
xnor g034 ( new_n172_, new_n171_, keyIn_0_12 );
xnor g035 ( new_n173_, N37, N53 );
xnor g036 ( new_n174_, new_n173_, keyIn_0_13 );
xnor g037 ( new_n175_, new_n172_, new_n174_ );
not g038 ( new_n176_, keyIn_0_22 );
not g039 ( new_n177_, keyIn_0_19 );
xnor g040 ( new_n178_, new_n159_, new_n177_ );
not g041 ( new_n179_, keyIn_0_18 );
xor g042 ( new_n180_, N97, N101 );
xnor g043 ( new_n181_, N105, N109 );
xnor g044 ( new_n182_, new_n180_, new_n181_ );
xnor g045 ( new_n183_, new_n182_, new_n179_ );
nand g046 ( new_n184_, new_n178_, new_n183_ );
not g047 ( new_n185_, new_n183_ );
nand g048 ( new_n186_, new_n160_, new_n185_ );
nand g049 ( new_n187_, new_n184_, new_n186_ );
xnor g050 ( new_n188_, new_n187_, new_n176_ );
nand g051 ( new_n189_, N130, N137 );
xor g052 ( new_n190_, new_n189_, keyIn_0_8 );
nand g053 ( new_n191_, new_n188_, new_n190_ );
xnor g054 ( new_n192_, new_n187_, keyIn_0_22 );
not g055 ( new_n193_, new_n190_ );
nand g056 ( new_n194_, new_n192_, new_n193_ );
nand g057 ( new_n195_, new_n191_, new_n194_ );
xnor g058 ( new_n196_, new_n195_, new_n175_ );
nor g059 ( new_n197_, new_n196_, new_n153_ );
nand g060 ( new_n198_, new_n197_, new_n170_ );
not g061 ( new_n199_, keyIn_0_24 );
xnor g062 ( new_n200_, new_n183_, new_n142_ );
nand g063 ( new_n201_, N131, N137 );
xnor g064 ( new_n202_, new_n200_, new_n201_ );
xnor g065 ( new_n203_, N9, N25 );
xnor g066 ( new_n204_, N41, N57 );
xnor g067 ( new_n205_, new_n203_, new_n204_ );
not g068 ( new_n206_, new_n205_ );
xnor g069 ( new_n207_, new_n202_, new_n206_ );
xnor g070 ( new_n208_, new_n207_, new_n199_ );
xnor g071 ( new_n209_, new_n208_, keyIn_0_26 );
nor g072 ( new_n210_, new_n198_, new_n209_ );
nand g073 ( new_n211_, new_n210_, new_n154_ );
nor g074 ( new_n212_, new_n210_, new_n154_ );
xnor g075 ( new_n213_, new_n148_, new_n151_ );
xnor g076 ( new_n214_, new_n207_, keyIn_0_24 );
nor g077 ( new_n215_, new_n214_, new_n213_ );
nand g078 ( new_n216_, new_n215_, new_n196_ );
not g079 ( new_n217_, new_n175_ );
xnor g080 ( new_n218_, new_n195_, new_n217_ );
not g081 ( new_n219_, keyIn_0_25 );
nand g082 ( new_n220_, new_n213_, new_n219_ );
nand g083 ( new_n221_, new_n153_, keyIn_0_25 );
nand g084 ( new_n222_, new_n220_, new_n221_ );
nor g085 ( new_n223_, new_n208_, new_n222_ );
nand g086 ( new_n224_, new_n223_, new_n218_ );
nand g087 ( new_n225_, new_n216_, new_n224_ );
nand g088 ( new_n226_, new_n225_, new_n170_ );
not g089 ( new_n227_, new_n170_ );
not g090 ( new_n228_, new_n215_ );
nor g091 ( new_n229_, new_n228_, new_n196_ );
nand g092 ( new_n230_, new_n229_, new_n227_ );
nand g093 ( new_n231_, new_n226_, new_n230_ );
nor g094 ( new_n232_, new_n212_, new_n231_ );
nand g095 ( new_n233_, new_n232_, new_n211_ );
xnor g096 ( new_n234_, N73, N89 );
xnor g097 ( new_n235_, N105, N121 );
xnor g098 ( new_n236_, new_n234_, new_n235_ );
xor g099 ( new_n237_, new_n236_, keyIn_0_20 );
nand g100 ( new_n238_, N135, N137 );
xnor g101 ( new_n239_, new_n238_, keyIn_0_10 );
not g102 ( new_n240_, keyIn_0_21 );
not g103 ( new_n241_, keyIn_0_17 );
not g104 ( new_n242_, keyIn_0_2 );
xnor g105 ( new_n243_, N33, N37 );
xnor g106 ( new_n244_, new_n243_, new_n242_ );
not g107 ( new_n245_, keyIn_0_3 );
xnor g108 ( new_n246_, N41, N45 );
xnor g109 ( new_n247_, new_n246_, new_n245_ );
nand g110 ( new_n248_, new_n244_, new_n247_ );
xnor g111 ( new_n249_, new_n243_, keyIn_0_2 );
nand g112 ( new_n250_, new_n246_, keyIn_0_3 );
nand g113 ( new_n251_, N41, N45 );
not g114 ( new_n252_, new_n251_ );
nor g115 ( new_n253_, N41, N45 );
nor g116 ( new_n254_, new_n252_, new_n253_ );
nand g117 ( new_n255_, new_n254_, new_n245_ );
nand g118 ( new_n256_, new_n255_, new_n250_ );
nand g119 ( new_n257_, new_n249_, new_n256_ );
nand g120 ( new_n258_, new_n248_, new_n257_ );
nand g121 ( new_n259_, new_n258_, new_n241_ );
xnor g122 ( new_n260_, new_n244_, new_n256_ );
nand g123 ( new_n261_, new_n260_, keyIn_0_17 );
nand g124 ( new_n262_, new_n261_, new_n259_ );
not g125 ( new_n263_, keyIn_0_16 );
xnor g126 ( new_n264_, N1, N13 );
xnor g127 ( new_n265_, N5, N9 );
xnor g128 ( new_n266_, new_n264_, new_n265_ );
xnor g129 ( new_n267_, new_n266_, new_n263_ );
nand g130 ( new_n268_, new_n262_, new_n267_ );
xnor g131 ( new_n269_, new_n258_, keyIn_0_17 );
xnor g132 ( new_n270_, new_n266_, keyIn_0_16 );
nand g133 ( new_n271_, new_n269_, new_n270_ );
nand g134 ( new_n272_, new_n271_, new_n268_ );
nand g135 ( new_n273_, new_n272_, new_n240_ );
xnor g136 ( new_n274_, new_n262_, new_n270_ );
nand g137 ( new_n275_, new_n274_, keyIn_0_21 );
nand g138 ( new_n276_, new_n275_, new_n273_ );
nand g139 ( new_n277_, new_n276_, new_n239_ );
not g140 ( new_n278_, new_n239_ );
xnor g141 ( new_n279_, new_n272_, keyIn_0_21 );
nand g142 ( new_n280_, new_n279_, new_n278_ );
nand g143 ( new_n281_, new_n280_, new_n277_ );
xnor g144 ( new_n282_, new_n281_, new_n237_ );
xnor g145 ( new_n283_, N69, N85 );
xnor g146 ( new_n284_, N101, N117 );
xnor g147 ( new_n285_, new_n283_, new_n284_ );
xnor g148 ( new_n286_, N57, N61 );
not g149 ( new_n287_, keyIn_0_4 );
xnor g150 ( new_n288_, N49, N53 );
xnor g151 ( new_n289_, new_n288_, new_n287_ );
xnor g152 ( new_n290_, new_n289_, new_n286_ );
nand g153 ( new_n291_, new_n262_, new_n290_ );
not g154 ( new_n292_, new_n286_ );
xnor g155 ( new_n293_, new_n289_, new_n292_ );
nand g156 ( new_n294_, new_n269_, new_n293_ );
nand g157 ( new_n295_, new_n294_, new_n291_ );
nand g158 ( new_n296_, N134, N137 );
not g159 ( new_n297_, new_n296_ );
xnor g160 ( new_n298_, new_n295_, new_n297_ );
nand g161 ( new_n299_, new_n298_, new_n285_ );
not g162 ( new_n300_, new_n285_ );
xnor g163 ( new_n301_, new_n295_, new_n296_ );
nand g164 ( new_n302_, new_n301_, new_n300_ );
nand g165 ( new_n303_, new_n299_, new_n302_ );
not g166 ( new_n304_, new_n303_ );
xor g167 ( new_n305_, N97, N113 );
xnor g168 ( new_n306_, new_n305_, keyIn_0_15 );
xnor g169 ( new_n307_, N65, N81 );
xnor g170 ( new_n308_, new_n306_, new_n307_ );
not g171 ( new_n309_, new_n308_ );
not g172 ( new_n310_, keyIn_0_1 );
xnor g173 ( new_n311_, N25, N29 );
xnor g174 ( new_n312_, new_n311_, new_n310_ );
not g175 ( new_n313_, keyIn_0_0 );
xnor g176 ( new_n314_, N17, N21 );
xnor g177 ( new_n315_, new_n314_, new_n313_ );
xnor g178 ( new_n316_, new_n312_, new_n315_ );
nand g179 ( new_n317_, new_n267_, new_n316_ );
xnor g180 ( new_n318_, new_n314_, keyIn_0_0 );
nand g181 ( new_n319_, new_n312_, new_n318_ );
xnor g182 ( new_n320_, new_n311_, keyIn_0_1 );
nand g183 ( new_n321_, new_n320_, new_n315_ );
nand g184 ( new_n322_, new_n319_, new_n321_ );
nand g185 ( new_n323_, new_n270_, new_n322_ );
nand g186 ( new_n324_, new_n317_, new_n323_ );
nand g187 ( new_n325_, N133, N137 );
xnor g188 ( new_n326_, new_n324_, new_n325_ );
nand g189 ( new_n327_, new_n326_, new_n309_ );
not g190 ( new_n328_, new_n325_ );
xnor g191 ( new_n329_, new_n324_, new_n328_ );
nand g192 ( new_n330_, new_n329_, new_n308_ );
nand g193 ( new_n331_, new_n330_, new_n327_ );
not g194 ( new_n332_, new_n331_ );
nand g195 ( new_n333_, new_n304_, new_n332_ );
xnor g196 ( new_n334_, N77, N93 );
xnor g197 ( new_n335_, N109, N125 );
xnor g198 ( new_n336_, new_n334_, new_n335_ );
nand g199 ( new_n337_, N136, N137 );
xnor g200 ( new_n338_, new_n337_, keyIn_0_11 );
nand g201 ( new_n339_, new_n290_, new_n322_ );
nand g202 ( new_n340_, new_n316_, new_n293_ );
nand g203 ( new_n341_, new_n340_, new_n339_ );
xnor g204 ( new_n342_, new_n341_, new_n338_ );
nand g205 ( new_n343_, new_n342_, new_n336_ );
not g206 ( new_n344_, new_n336_ );
not g207 ( new_n345_, new_n338_ );
xnor g208 ( new_n346_, new_n341_, new_n345_ );
nand g209 ( new_n347_, new_n346_, new_n344_ );
nand g210 ( new_n348_, new_n347_, new_n343_ );
not g211 ( new_n349_, new_n348_ );
nor g212 ( new_n350_, new_n333_, new_n349_ );
nand g213 ( new_n351_, new_n350_, new_n282_ );
not g214 ( new_n352_, new_n351_ );
nand g215 ( new_n353_, new_n233_, new_n352_ );
nor g216 ( new_n354_, new_n353_, new_n153_ );
xnor g217 ( new_n355_, new_n354_, keyIn_0_41 );
xnor g218 ( N724, new_n355_, N1 );
nor g219 ( new_n357_, new_n353_, new_n218_ );
xnor g220 ( new_n358_, new_n357_, keyIn_0_42 );
xor g221 ( N725, new_n358_, N5 );
not g222 ( new_n360_, new_n353_ );
nand g223 ( new_n361_, new_n360_, new_n214_ );
xnor g224 ( N726, new_n361_, N9 );
nand g225 ( new_n363_, new_n360_, new_n227_ );
xnor g226 ( N727, new_n363_, N13 );
not g227 ( new_n365_, new_n237_ );
nand g228 ( new_n366_, new_n281_, new_n365_ );
xnor g229 ( new_n367_, new_n276_, new_n278_ );
nand g230 ( new_n368_, new_n367_, new_n237_ );
nand g231 ( new_n369_, new_n368_, new_n366_ );
nor g232 ( new_n370_, new_n333_, new_n348_ );
nand g233 ( new_n371_, new_n370_, new_n369_ );
not g234 ( new_n372_, new_n371_ );
nand g235 ( new_n373_, new_n233_, new_n372_ );
nor g236 ( new_n374_, new_n373_, new_n153_ );
xnor g237 ( new_n375_, new_n374_, N17 );
xor g238 ( N728, new_n375_, keyIn_0_54 );
nor g239 ( new_n377_, new_n373_, new_n218_ );
xnor g240 ( new_n378_, new_n377_, N21 );
xor g241 ( N729, new_n378_, keyIn_0_55 );
nor g242 ( new_n380_, new_n373_, new_n208_ );
xor g243 ( N730, new_n380_, N25 );
nor g244 ( new_n382_, new_n373_, new_n170_ );
xnor g245 ( new_n383_, new_n382_, keyIn_0_43 );
xnor g246 ( N731, new_n383_, N29 );
nand g247 ( new_n385_, new_n303_, new_n331_ );
nor g248 ( new_n386_, new_n385_, new_n349_ );
not g249 ( new_n387_, new_n386_ );
nor g250 ( new_n388_, new_n387_, new_n369_ );
nand g251 ( new_n389_, new_n233_, new_n388_ );
nor g252 ( new_n390_, new_n389_, new_n153_ );
xor g253 ( new_n391_, new_n390_, N33 );
xnor g254 ( N732, new_n391_, keyIn_0_56 );
nor g255 ( new_n393_, new_n389_, new_n218_ );
xnor g256 ( new_n394_, new_n393_, N37 );
xnor g257 ( N733, new_n394_, keyIn_0_57 );
nor g258 ( new_n396_, new_n389_, new_n208_ );
xnor g259 ( new_n397_, new_n396_, keyIn_0_44 );
xnor g260 ( N734, new_n397_, N41 );
not g261 ( new_n399_, keyIn_0_58 );
not g262 ( new_n400_, keyIn_0_45 );
nor g263 ( new_n401_, new_n389_, new_n170_ );
xnor g264 ( new_n402_, new_n401_, new_n400_ );
xnor g265 ( new_n403_, new_n402_, N45 );
xnor g266 ( N735, new_n403_, new_n399_ );
not g267 ( new_n405_, keyIn_0_59 );
not g268 ( new_n406_, keyIn_0_39 );
nor g269 ( new_n407_, new_n369_, keyIn_0_27 );
nand g270 ( new_n408_, new_n369_, keyIn_0_27 );
nor g271 ( new_n409_, new_n385_, new_n348_ );
nand g272 ( new_n410_, new_n408_, new_n409_ );
nor g273 ( new_n411_, new_n410_, new_n407_ );
nand g274 ( new_n412_, new_n233_, new_n411_ );
xnor g275 ( new_n413_, new_n412_, new_n406_ );
not g276 ( new_n414_, N49 );
nor g277 ( new_n415_, new_n153_, new_n414_ );
nand g278 ( new_n416_, new_n413_, new_n415_ );
xnor g279 ( new_n417_, new_n412_, keyIn_0_39 );
nor g280 ( new_n418_, new_n409_, new_n406_ );
nor g281 ( new_n419_, new_n417_, new_n418_ );
nand g282 ( new_n420_, new_n419_, new_n213_ );
nand g283 ( new_n421_, new_n420_, new_n414_ );
nand g284 ( new_n422_, new_n421_, new_n416_ );
nand g285 ( new_n423_, new_n422_, new_n405_ );
not g286 ( new_n424_, new_n418_ );
nand g287 ( new_n425_, new_n413_, new_n424_ );
nor g288 ( new_n426_, new_n425_, new_n153_ );
nand g289 ( new_n427_, new_n426_, N49 );
nor g290 ( new_n428_, new_n426_, N49 );
nor g291 ( new_n429_, new_n428_, new_n405_ );
nand g292 ( new_n430_, new_n429_, new_n427_ );
nand g293 ( N736, new_n430_, new_n423_ );
not g294 ( new_n432_, N53 );
not g295 ( new_n433_, keyIn_0_46 );
nor g296 ( new_n434_, new_n218_, new_n433_ );
nand g297 ( new_n435_, new_n413_, new_n434_ );
nand g298 ( new_n436_, new_n419_, new_n196_ );
nand g299 ( new_n437_, new_n436_, new_n433_ );
nand g300 ( new_n438_, new_n437_, new_n435_ );
nand g301 ( new_n439_, new_n438_, new_n432_ );
nor g302 ( new_n440_, new_n425_, new_n218_ );
nand g303 ( new_n441_, new_n440_, keyIn_0_46 );
nor g304 ( new_n442_, new_n440_, keyIn_0_46 );
nor g305 ( new_n443_, new_n442_, new_n432_ );
nand g306 ( new_n444_, new_n443_, new_n441_ );
nand g307 ( N737, new_n444_, new_n439_ );
nand g308 ( new_n446_, new_n419_, new_n214_ );
xnor g309 ( N738, new_n446_, N57 );
nand g310 ( new_n448_, new_n419_, new_n227_ );
xnor g311 ( N739, new_n448_, N61 );
not g312 ( new_n450_, keyIn_0_47 );
nor g313 ( new_n451_, new_n198_, new_n208_ );
nor g314 ( new_n452_, new_n282_, keyIn_0_31 );
not g315 ( new_n453_, new_n452_ );
not g316 ( new_n454_, keyIn_0_31 );
nor g317 ( new_n455_, new_n369_, new_n454_ );
nor g318 ( new_n456_, new_n455_, new_n387_ );
nand g319 ( new_n457_, new_n456_, new_n453_ );
nor g320 ( new_n458_, new_n457_, keyIn_0_37 );
nand g321 ( new_n459_, new_n457_, keyIn_0_37 );
not g322 ( new_n460_, keyIn_0_32 );
nor g323 ( new_n461_, new_n369_, new_n460_ );
nand g324 ( new_n462_, new_n369_, new_n460_ );
xnor g325 ( new_n463_, new_n348_, keyIn_0_33 );
nor g326 ( new_n464_, new_n333_, new_n463_ );
nand g327 ( new_n465_, new_n462_, new_n464_ );
nor g328 ( new_n466_, new_n465_, new_n461_ );
not g329 ( new_n467_, keyIn_0_28 );
nor g330 ( new_n468_, new_n303_, new_n467_ );
nand g331 ( new_n469_, new_n303_, new_n467_ );
nor g332 ( new_n470_, new_n332_, new_n348_ );
nand g333 ( new_n471_, new_n469_, new_n470_ );
nor g334 ( new_n472_, new_n471_, new_n468_ );
nand g335 ( new_n473_, new_n472_, new_n369_ );
not g336 ( new_n474_, keyIn_0_29 );
nand g337 ( new_n475_, new_n331_, new_n474_ );
not g338 ( new_n476_, keyIn_0_30 );
nand g339 ( new_n477_, new_n348_, new_n476_ );
nand g340 ( new_n478_, new_n475_, new_n477_ );
not g341 ( new_n479_, new_n478_ );
nor g342 ( new_n480_, new_n331_, new_n474_ );
nor g343 ( new_n481_, new_n348_, new_n476_ );
nor g344 ( new_n482_, new_n480_, new_n481_ );
nand g345 ( new_n483_, new_n479_, new_n482_ );
nor g346 ( new_n484_, new_n483_, new_n303_ );
nand g347 ( new_n485_, new_n484_, new_n282_ );
nand g348 ( new_n486_, new_n473_, new_n485_ );
nor g349 ( new_n487_, new_n466_, new_n486_ );
nand g350 ( new_n488_, new_n459_, new_n487_ );
nor g351 ( new_n489_, new_n488_, new_n458_ );
nand g352 ( new_n490_, new_n489_, keyIn_0_38 );
not g353 ( new_n491_, keyIn_0_38 );
not g354 ( new_n492_, new_n458_ );
not g355 ( new_n493_, keyIn_0_37 );
nand g356 ( new_n494_, new_n282_, keyIn_0_31 );
nand g357 ( new_n495_, new_n494_, new_n386_ );
nor g358 ( new_n496_, new_n495_, new_n452_ );
nor g359 ( new_n497_, new_n496_, new_n493_ );
not g360 ( new_n498_, new_n461_ );
nor g361 ( new_n499_, new_n282_, keyIn_0_32 );
not g362 ( new_n500_, new_n333_ );
not g363 ( new_n501_, new_n463_ );
nand g364 ( new_n502_, new_n500_, new_n501_ );
nor g365 ( new_n503_, new_n499_, new_n502_ );
nand g366 ( new_n504_, new_n503_, new_n498_ );
not g367 ( new_n505_, new_n486_ );
nand g368 ( new_n506_, new_n505_, new_n504_ );
nor g369 ( new_n507_, new_n506_, new_n497_ );
nand g370 ( new_n508_, new_n507_, new_n492_ );
nand g371 ( new_n509_, new_n508_, new_n491_ );
nand g372 ( new_n510_, new_n509_, new_n490_ );
nand g373 ( new_n511_, new_n510_, new_n451_ );
xnor g374 ( new_n512_, new_n511_, keyIn_0_40 );
nand g375 ( new_n513_, new_n512_, new_n332_ );
nand g376 ( new_n514_, new_n513_, new_n450_ );
not g377 ( new_n515_, keyIn_0_40 );
xnor g378 ( new_n516_, new_n511_, new_n515_ );
nor g379 ( new_n517_, new_n516_, new_n331_ );
nand g380 ( new_n518_, new_n517_, keyIn_0_47 );
nand g381 ( new_n519_, new_n518_, new_n514_ );
nand g382 ( new_n520_, new_n519_, N65 );
not g383 ( new_n521_, N65 );
xnor g384 ( new_n522_, new_n513_, keyIn_0_47 );
nand g385 ( new_n523_, new_n522_, new_n521_ );
nand g386 ( N740, new_n523_, new_n520_ );
not g387 ( new_n525_, keyIn_0_48 );
nand g388 ( new_n526_, new_n512_, new_n303_ );
nand g389 ( new_n527_, new_n526_, new_n525_ );
nor g390 ( new_n528_, new_n516_, new_n304_ );
nand g391 ( new_n529_, new_n528_, keyIn_0_48 );
nand g392 ( new_n530_, new_n529_, new_n527_ );
nand g393 ( new_n531_, new_n530_, N69 );
not g394 ( new_n532_, N69 );
xnor g395 ( new_n533_, new_n526_, keyIn_0_48 );
nand g396 ( new_n534_, new_n533_, new_n532_ );
nand g397 ( N741, new_n534_, new_n531_ );
nand g398 ( new_n536_, new_n512_, new_n282_ );
xnor g399 ( N742, new_n536_, N73 );
not g400 ( new_n538_, keyIn_0_60 );
not g401 ( new_n539_, N77 );
nand g402 ( new_n540_, new_n512_, new_n349_ );
nand g403 ( new_n541_, new_n540_, new_n539_ );
nor g404 ( new_n542_, new_n516_, new_n348_ );
nand g405 ( new_n543_, new_n542_, N77 );
nand g406 ( new_n544_, new_n543_, new_n541_ );
nand g407 ( new_n545_, new_n544_, new_n538_ );
xnor g408 ( new_n546_, new_n540_, N77 );
nand g409 ( new_n547_, new_n546_, keyIn_0_60 );
nand g410 ( N743, new_n547_, new_n545_ );
xnor g411 ( new_n549_, new_n489_, new_n491_ );
not g412 ( new_n550_, keyIn_0_34 );
nor g413 ( new_n551_, new_n218_, new_n550_ );
nor g414 ( new_n552_, new_n196_, keyIn_0_34 );
nor g415 ( new_n553_, new_n214_, new_n153_ );
nand g416 ( new_n554_, new_n227_, new_n553_ );
nor g417 ( new_n555_, new_n554_, new_n552_ );
not g418 ( new_n556_, new_n555_ );
nor g419 ( new_n557_, new_n556_, new_n551_ );
not g420 ( new_n558_, new_n557_ );
nor g421 ( new_n559_, new_n549_, new_n558_ );
nand g422 ( new_n560_, new_n559_, new_n332_ );
xnor g423 ( N744, new_n560_, N81 );
nand g424 ( new_n562_, new_n559_, new_n303_ );
xnor g425 ( new_n563_, new_n562_, keyIn_0_49 );
xnor g426 ( N745, new_n563_, N85 );
nand g427 ( new_n565_, new_n559_, new_n282_ );
xnor g428 ( new_n566_, new_n565_, N89 );
xnor g429 ( N746, new_n566_, keyIn_0_61 );
nand g430 ( new_n568_, new_n559_, new_n349_ );
xnor g431 ( N747, new_n568_, N93 );
xnor g432 ( new_n570_, new_n213_, keyIn_0_35 );
nand g433 ( new_n571_, new_n570_, new_n214_ );
nor g434 ( new_n572_, new_n571_, new_n218_ );
nand g435 ( new_n573_, new_n572_, new_n170_ );
not g436 ( new_n574_, new_n573_ );
nand g437 ( new_n575_, new_n510_, new_n574_ );
not g438 ( new_n576_, new_n575_ );
nand g439 ( new_n577_, new_n576_, new_n332_ );
xnor g440 ( N748, new_n577_, N97 );
nor g441 ( new_n579_, new_n575_, new_n304_ );
xnor g442 ( new_n580_, new_n579_, keyIn_0_50 );
xor g443 ( N749, new_n580_, N101 );
nand g444 ( new_n582_, new_n576_, new_n282_ );
xnor g445 ( N750, new_n582_, N105 );
nand g446 ( new_n584_, new_n576_, new_n349_ );
xnor g447 ( N751, new_n584_, N109 );
nor g448 ( new_n586_, new_n216_, new_n170_ );
not g449 ( new_n587_, new_n586_ );
nor g450 ( new_n588_, new_n549_, new_n587_ );
nand g451 ( new_n589_, new_n588_, new_n332_ );
xnor g452 ( N752, new_n589_, N113 );
nand g453 ( new_n591_, new_n510_, new_n586_ );
nor g454 ( new_n592_, new_n591_, new_n304_ );
xnor g455 ( new_n593_, new_n592_, keyIn_0_51 );
xnor g456 ( N753, new_n593_, N117 );
not g457 ( new_n595_, N121 );
nor g458 ( new_n596_, new_n591_, new_n369_ );
nand g459 ( new_n597_, new_n596_, keyIn_0_52 );
not g460 ( new_n598_, keyIn_0_52 );
nand g461 ( new_n599_, new_n588_, new_n282_ );
nand g462 ( new_n600_, new_n599_, new_n598_ );
nand g463 ( new_n601_, new_n600_, new_n597_ );
nand g464 ( new_n602_, new_n601_, new_n595_ );
xnor g465 ( new_n603_, new_n596_, new_n598_ );
nand g466 ( new_n604_, new_n603_, N121 );
nand g467 ( new_n605_, new_n604_, new_n602_ );
nand g468 ( new_n606_, new_n605_, keyIn_0_62 );
not g469 ( new_n607_, keyIn_0_62 );
xnor g470 ( new_n608_, new_n601_, N121 );
nand g471 ( new_n609_, new_n608_, new_n607_ );
nand g472 ( N754, new_n609_, new_n606_ );
not g473 ( new_n611_, keyIn_0_63 );
not g474 ( new_n612_, keyIn_0_53 );
nor g475 ( new_n613_, new_n591_, new_n348_ );
nand g476 ( new_n614_, new_n613_, new_n612_ );
nand g477 ( new_n615_, new_n588_, new_n349_ );
nand g478 ( new_n616_, new_n615_, keyIn_0_53 );
nand g479 ( new_n617_, new_n616_, new_n614_ );
xnor g480 ( new_n618_, new_n617_, N125 );
nand g481 ( new_n619_, new_n618_, new_n611_ );
not g482 ( new_n620_, N125 );
nand g483 ( new_n621_, new_n617_, new_n620_ );
xnor g484 ( new_n622_, new_n613_, keyIn_0_53 );
nand g485 ( new_n623_, new_n622_, N125 );
nand g486 ( new_n624_, new_n623_, new_n621_ );
nand g487 ( new_n625_, new_n624_, keyIn_0_63 );
nand g488 ( N755, new_n619_, new_n625_ );
endmodule