module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n1359_, new_n595_, new_n445_, new_n1009_, new_n238_, new_n479_, new_n1105_, new_n1215_, new_n1448_, new_n608_, new_n501_, new_n1157_, new_n1442_, new_n1345_, new_n421_, new_n777_, new_n1433_, new_n1575_, new_n1472_, new_n1048_, new_n885_, new_n439_, new_n1532_, new_n283_, new_n223_, new_n390_, new_n743_, new_n1327_, new_n241_, new_n1535_, new_n566_, new_n641_, new_n339_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n1351_, new_n556_, new_n636_, new_n691_, new_n1024_, new_n670_, new_n456_, new_n1125_, new_n246_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n1237_, new_n728_, new_n1479_, new_n1071_, new_n1294_, new_n214_, new_n894_, new_n853_, new_n695_, new_n660_, new_n1311_, new_n526_, new_n908_, new_n552_, new_n678_, new_n342_, new_n706_, new_n649_, new_n1119_, new_n752_, new_n1524_, new_n1045_, new_n1305_, new_n500_, new_n1163_, new_n786_, new_n317_, new_n1188_, new_n1415_, new_n1390_, new_n721_, new_n504_, new_n1414_, new_n742_, new_n892_, new_n1368_, new_n234_, new_n472_, new_n873_, new_n1167_, new_n1530_, new_n1300_, new_n1490_, new_n774_, new_n792_, new_n953_, new_n257_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n449_, new_n580_, new_n639_, new_n484_, new_n766_, new_n272_, new_n282_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n1332_, new_n1447_, new_n635_, new_n685_, new_n326_, new_n648_, new_n903_, new_n983_, new_n822_, new_n1406_, new_n1082_, new_n1018_, new_n606_, new_n796_, new_n1054_, new_n655_, new_n1288_, new_n630_, new_n385_, new_n1049_, new_n1330_, new_n694_, new_n461_, new_n1323_, new_n297_, new_n565_, new_n1196_, new_n1366_, new_n511_, new_n303_, new_n325_, new_n1285_, new_n1031_, new_n1216_, new_n1281_, new_n629_, new_n1214_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n324_, new_n960_, new_n1377_, new_n549_, new_n491_, new_n676_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n1362_, new_n1404_, new_n1443_, new_n1484_, new_n497_, new_n816_, new_n1355_, new_n568_, new_n420_, new_n876_, new_n423_, new_n498_, new_n496_, new_n1217_, new_n1046_, new_n1182_, new_n708_, new_n206_, new_n1463_, new_n429_, new_n1222_, new_n353_, new_n734_, new_n912_, new_n1424_, new_n1062_, new_n680_, new_n981_, new_n506_, new_n872_, new_n1527_, new_n1275_, new_n1277_, new_n1428_, new_n1440_, new_n656_, new_n1127_, new_n388_, new_n1028_, new_n1168_, new_n483_, new_n1004_, new_n1152_, new_n1558_, new_n299_, new_n394_, new_n935_, new_n657_, new_n1150_, new_n652_, new_n582_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n785_, new_n1501_, new_n441_, new_n477_, new_n664_, new_n600_, new_n280_, new_n1041_, new_n1562_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n1576_, new_n301_, new_n1333_, new_n1132_, new_n395_, new_n383_, new_n343_, new_n854_, new_n458_, new_n1106_, new_n207_, new_n267_, new_n1395_, new_n473_, new_n1147_, new_n1373_, new_n1229_, new_n1422_, new_n1523_, new_n1468_, new_n969_, new_n334_, new_n331_, new_n1234_, new_n835_, new_n1360_, new_n378_, new_n1574_, new_n621_, new_n1423_, new_n244_, new_n705_, new_n943_, new_n874_, new_n402_, new_n1321_, new_n1209_, new_n335_, new_n347_, new_n659_, new_n700_, new_n1419_, new_n921_, new_n346_, new_n396_, new_n1315_, new_n1003_, new_n696_, new_n208_, new_n1039_, new_n1439_, new_n1365_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n729_, new_n1111_, new_n1413_, new_n1218_, new_n1385_, new_n1346_, new_n1201_, new_n559_, new_n1282_, new_n762_, new_n1349_, new_n1193_, new_n1547_, new_n1437_, new_n1187_, new_n1205_, new_n1154_, new_n1253_, new_n295_, new_n1453_, new_n1256_, new_n628_, new_n1513_, new_n409_, new_n1090_, new_n745_, new_n1489_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n1171_, new_n867_, new_n954_, new_n1032_, new_n1545_, new_n276_, new_n901_, new_n688_, new_n1255_, new_n410_, new_n985_, new_n851_, new_n1518_, new_n932_, new_n878_, new_n543_, new_n886_, new_n371_, new_n509_, new_n202_, new_n296_, new_n661_, new_n797_, new_n232_, new_n1358_, new_n724_, new_n1070_, new_n1416_, new_n1109_, new_n261_, new_n672_, new_n1496_, new_n616_, new_n529_, new_n323_, new_n914_, new_n884_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n604_, new_n1104_, new_n1511_, new_n571_, new_n1504_, new_n758_, new_n460_, new_n1267_, new_n328_, new_n268_, new_n1466_, new_n1516_, new_n1299_, new_n380_, new_n1477_, new_n1079_, new_n861_, new_n1564_, new_n1252_, new_n352_, new_n1553_, new_n931_, new_n575_, new_n1493_, new_n562_, new_n944_, new_n1542_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n1480_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n963_, new_n1481_, new_n1325_, new_n993_, new_n1191_, new_n1357_, new_n824_, new_n717_, new_n1455_, new_n403_, new_n868_, new_n1242_, new_n475_, new_n237_, new_n858_, new_n1384_, new_n1343_, new_n936_, new_n1459_, new_n1434_, new_n1438_, new_n1016_, new_n411_, new_n673_, new_n1144_, new_n1465_, new_n666_, new_n1290_, new_n407_, new_n1519_, new_n1407_, new_n879_, new_n1417_, new_n736_, new_n513_, new_n558_, new_n219_, new_n382_, new_n313_, new_n1370_, new_n239_, new_n718_, new_n1310_, new_n1398_, new_n1126_, new_n546_, new_n612_, new_n1015_, new_n919_, new_n302_, new_n755_, new_n1040_, new_n1509_, new_n1559_, new_n544_, new_n615_, new_n722_, new_n856_, new_n415_, new_n1324_, new_n1293_, new_n537_, new_n1336_, new_n345_, new_n499_, new_n533_, new_n255_, new_n1130_, new_n795_, new_n459_, new_n1441_, new_n1122_, new_n1240_, new_n1510_, new_n354_, new_n1174_, new_n968_, new_n1464_, new_n613_, new_n1508_, new_n337_, new_n1195_, new_n417_, new_n658_, new_n837_, new_n591_, new_n801_, new_n1458_, new_n631_, new_n453_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n1521_, new_n1334_, new_n531_, new_n593_, new_n1543_, new_n974_, new_n1565_, new_n252_, new_n751_, new_n1038_, new_n372_, new_n852_, new_n1454_, new_n1474_, new_n1328_, new_n978_, new_n1308_, new_n408_, new_n1430_, new_n470_, new_n213_, new_n769_, new_n433_, new_n871_, new_n1450_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n689_, new_n933_, new_n584_, new_n815_, new_n1492_, new_n1367_, new_n278_, new_n304_, new_n1052_, new_n1425_, new_n857_, new_n1379_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n269_, new_n512_, new_n1471_, new_n1220_, new_n989_, new_n1117_, new_n1421_, new_n644_, new_n836_, new_n1116_, new_n904_, new_n1392_, new_n1276_, new_n1444_, new_n913_, new_n327_, new_n681_, new_n594_, new_n561_, new_n495_, new_n927_, new_n431_, new_n1206_, new_n1427_, new_n818_, new_n881_, new_n1268_, new_n1376_, new_n1381_, new_n1566_, new_n1534_, new_n684_, new_n640_, new_n754_, new_n653_, new_n905_, new_n377_, new_n1258_, new_n1539_, new_n375_, new_n962_, new_n760_, new_n627_, new_n1391_, new_n1436_, new_n567_, new_n1353_, new_n1033_, new_n576_, new_n831_, new_n791_, new_n1153_, new_n357_, new_n1339_, new_n320_, new_n984_, new_n780_, new_n1183_, new_n245_, new_n643_, new_n1316_, new_n1194_, new_n1338_, new_n1460_, new_n1230_, new_n1027_, new_n348_, new_n610_, new_n1369_, new_n843_, new_n322_, new_n703_, new_n698_, new_n1165_, new_n1401_, new_n1259_, new_n226_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n1235_, new_n1320_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n686_, new_n293_, new_n934_, new_n1567_, new_n770_, new_n1389_, new_n1400_, new_n757_, new_n1225_, new_n521_, new_n793_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n1089_, new_n1192_, new_n405_, new_n942_, new_n614_, new_n895_, new_n958_, new_n976_, new_n699_, new_n236_, new_n1405_, new_n1249_, new_n1354_, new_n955_, new_n847_, new_n250_, new_n888_, new_n1505_, new_n288_, new_n1340_, new_n798_, new_n817_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1361_, new_n941_, new_n1410_, new_n738_, new_n827_, new_n1356_, new_n1363_, new_n1317_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n365_, new_n859_, new_n1211_, new_n1412_, new_n1207_, new_n1176_, new_n1374_, new_n601_, new_n842_, new_n1552_, new_n1057_, new_n682_, new_n1075_, new_n812_, new_n266_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1397_, new_n220_, new_n1402_, new_n1313_, new_n1172_, new_n419_, new_n624_, new_n534_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n804_, new_n1342_, new_n424_, new_n602_, new_n1210_, new_n1060_, new_n1303_, new_n240_, new_n413_, new_n1544_, new_n1382_, new_n442_, new_n677_, new_n1487_, new_n642_, new_n211_, new_n1418_, new_n462_, new_n603_, new_n564_, new_n1528_, new_n761_, new_n840_, new_n735_, new_n1283_, new_n898_, new_n799_, new_n1304_, new_n1537_, new_n946_, new_n344_, new_n287_, new_n1108_, new_n1469_, new_n862_, new_n427_, new_n532_, new_n393_, new_n418_, new_n746_, new_n1221_, new_n292_, new_n215_, new_n1319_, new_n626_, new_n959_, new_n990_, new_n716_, new_n701_, new_n1058_, new_n1162_, new_n212_, new_n1278_, new_n902_, new_n364_, new_n832_, new_n414_, new_n1101_, new_n1250_, new_n315_, new_n1482_, new_n1050_, new_n554_, new_n230_, new_n1151_, new_n844_, new_n1302_, new_n281_, new_n430_, new_n482_, new_n849_, new_n855_, new_n1037_, new_n589_, new_n248_, new_n350_, new_n759_, new_n1083_, new_n1297_, new_n829_, new_n1257_, new_n1306_, new_n988_, new_n478_, new_n1307_, new_n1228_, new_n710_, new_n971_, new_n1486_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1409_, new_n1429_, new_n463_, new_n1372_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n1292_, new_n1426_, new_n517_, new_n609_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n702_, new_n833_, new_n1560_, new_n715_, new_n811_, new_n1445_, new_n1371_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n970_, new_n466_, new_n262_, new_n218_, new_n845_, new_n768_, new_n773_, new_n305_, new_n1452_, new_n1051_, new_n899_, new_n1053_, new_n1540_, new_n205_, new_n492_, new_n1200_, new_n1533_, new_n650_, new_n750_, new_n887_, new_n254_, new_n355_, new_n926_, new_n432_, new_n925_, new_n875_, new_n256_, new_n1226_, new_n778_, new_n452_, new_n381_, new_n1483_, new_n1219_, new_n920_, new_n1121_, new_n1495_, new_n1341_, new_n820_, new_n1386_, new_n771_, new_n979_, new_n508_, new_n1435_, new_n714_, new_n1280_, new_n1007_, new_n1241_, new_n882_, new_n1145_, new_n1557_, new_n929_, new_n986_, new_n1159_, new_n314_, new_n1337_, new_n216_, new_n1348_, new_n917_, new_n1555_, new_n1322_, new_n1133_, new_n1177_, new_n646_, new_n538_, new_n1026_, new_n541_, new_n210_, new_n447_, new_n1388_, new_n1550_, new_n790_, new_n1081_, new_n311_, new_n587_, new_n1247_, new_n1411_, new_n465_, new_n783_, new_n1380_, new_n739_, new_n263_, new_n341_, new_n996_, new_n1318_, new_n846_, new_n915_, new_n488_, new_n524_, new_n349_, new_n848_, new_n277_, new_n1245_, new_n663_, new_n1499_, new_n1497_, new_n579_, new_n286_, new_n1375_, new_n1254_, new_n438_, new_n1344_, new_n939_, new_n1393_, new_n632_, new_n1335_, new_n1364_, new_n671_, new_n965_, new_n1514_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n1526_, new_n397_, new_n1446_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n945_, new_n870_, new_n805_, new_n1420_, new_n1403_, new_n1115_, new_n1383_, new_n1231_, new_n948_, new_n1520_, new_n1055_, new_n1431_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n457_, new_n1301_, new_n1128_, new_n1002_, new_n1169_, new_n448_, new_n384_, new_n900_, new_n1329_, new_n1161_, new_n924_, new_n775_, new_n454_, new_n1034_, new_n1124_, new_n1000_, new_n308_, new_n633_, new_n784_, new_n1273_, new_n1396_, new_n1491_, new_n1554_, new_n258_, new_n860_, new_n306_, new_n494_, new_n291_, new_n309_, new_n1160_, new_n1166_, new_n259_, new_n654_, new_n1456_, new_n713_, new_n880_, new_n1102_, new_n227_, new_n690_, new_n416_, new_n1043_, new_n222_, new_n744_, new_n400_, new_n1136_, new_n1272_, new_n693_, new_n1287_, new_n505_, new_n1462_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1538_, new_n1561_, new_n1271_, new_n1251_, new_n747_, new_n749_, new_n1091_, new_n1095_, new_n310_, new_n275_, new_n998_, new_n1056_, new_n1331_, new_n1094_, new_n839_, new_n1030_, new_n485_, new_n578_, new_n525_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1284_, new_n1572_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n1387_, new_n719_, new_n869_, new_n1178_, new_n1525_, new_n270_, new_n570_, new_n598_, new_n893_, new_n1063_, new_n520_, new_n1347_, new_n1001_, new_n253_, new_n825_, new_n557_, new_n260_, new_n251_, new_n300_, new_n1503_, new_n507_, new_n741_, new_n806_, new_n605_, new_n1224_, new_n1074_, new_n748_, new_n1137_, new_n1286_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n1326_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n231_, new_n1080_, new_n583_, new_n617_, new_n1279_, new_n1467_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n916_, new_n428_, new_n487_, new_n675_, new_n1155_, new_n360_, new_n1186_, new_n1261_, new_n225_, new_n1246_, new_n1488_, new_n922_, new_n387_, new_n476_, new_n987_, new_n949_, new_n221_, new_n450_, new_n1394_, new_n243_, new_n1179_, new_n298_, new_n1088_, new_n1148_, new_n1146_, new_n569_, new_n555_, new_n468_, new_n977_, new_n1139_, new_n782_, new_n444_, new_n392_, new_n518_, new_n950_, new_n737_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n209_, new_n623_, new_n446_, new_n316_, new_n203_, new_n590_, new_n826_, new_n789_, new_n1476_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n516_, new_n1227_, new_n1352_, new_n733_, new_n1021_, new_n1076_, new_n585_, new_n1350_, new_n312_, new_n535_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n1244_, new_n307_, new_n1378_, new_n1478_, new_n1181_, new_n1093_, new_n597_, new_n1451_, new_n1092_, new_n1143_, new_n1072_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n1164_, new_n1296_, new_n435_, new_n1309_, new_n1010_, new_n776_, new_n687_, new_n1029_, new_n370_, new_n1515_, new_n638_, new_n523_, new_n909_, new_n1571_, new_n217_, new_n788_, new_n841_, new_n1457_, new_n1204_, new_n1470_, new_n1112_, new_n711_, new_n1156_, new_n1298_, new_n731_, new_n599_, new_n930_, new_n1475_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n1529_, new_n645_, new_n1087_, new_n1096_, new_n723_, new_n756_, new_n823_, new_n1549_, new_n1577_, new_n574_, new_n1500_, new_n928_, new_n1548_, new_n319_, new_n1008_, new_n338_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n1134_, new_n336_, new_n1291_, new_n247_, new_n539_, new_n1399_, new_n803_, new_n330_, new_n1270_, new_n727_, new_n1531_, new_n294_, new_n1295_, new_n1173_, new_n704_, new_n1432_, new_n1570_, new_n1189_, new_n1197_, new_n1312_, new_n1502_, new_n474_, new_n1223_, new_n1129_, new_n1013_, new_n467_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n358_, new_n877_, new_n1506_, new_n545_, new_n228_, new_n611_, new_n289_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n1236_, new_n866_, new_n1556_, new_n947_, new_n994_, new_n982_, new_n1494_, new_n964_, new_n1078_, new_n551_, new_n1408_, new_n279_, new_n455_, new_n1569_, new_n618_, new_n1140_, new_n1042_, new_n863_, new_n828_, new_n980_, new_n464_, new_n1498_, new_n204_, new_n573_, new_n765_, new_n1314_, new_n1103_;

not g0000 ( new_n202_, keyIn_0_64 );
not g0001 ( new_n203_, keyIn_0_60 );
not g0002 ( new_n204_, keyIn_0_44 );
not g0003 ( new_n205_, keyIn_0_8 );
not g0004 ( new_n206_, N69 );
nand g0005 ( new_n207_, new_n206_, N65 );
not g0006 ( new_n208_, N65 );
nand g0007 ( new_n209_, new_n208_, N69 );
nand g0008 ( new_n210_, new_n207_, new_n209_ );
nand g0009 ( new_n211_, new_n210_, new_n205_ );
nor g0010 ( new_n212_, new_n210_, new_n205_ );
not g0011 ( new_n213_, new_n212_ );
nand g0012 ( new_n214_, new_n213_, new_n211_ );
not g0013 ( new_n215_, keyIn_0_9 );
not g0014 ( new_n216_, N77 );
nand g0015 ( new_n217_, new_n216_, N73 );
not g0016 ( new_n218_, N73 );
nand g0017 ( new_n219_, new_n218_, N77 );
nand g0018 ( new_n220_, new_n217_, new_n219_ );
nor g0019 ( new_n221_, new_n220_, new_n215_ );
nand g0020 ( new_n222_, new_n220_, new_n215_ );
not g0021 ( new_n223_, new_n222_ );
nor g0022 ( new_n224_, new_n223_, new_n221_ );
nand g0023 ( new_n225_, new_n224_, new_n214_ );
not g0024 ( new_n226_, new_n211_ );
nor g0025 ( new_n227_, new_n226_, new_n212_ );
not g0026 ( new_n228_, new_n221_ );
nand g0027 ( new_n229_, new_n228_, new_n222_ );
nand g0028 ( new_n230_, new_n227_, new_n229_ );
nand g0029 ( new_n231_, new_n225_, new_n230_ );
nand g0030 ( new_n232_, new_n231_, new_n204_ );
not g0031 ( new_n233_, new_n232_ );
nor g0032 ( new_n234_, new_n231_, new_n204_ );
nor g0033 ( new_n235_, new_n233_, new_n234_ );
not g0034 ( new_n236_, keyIn_0_45 );
not g0035 ( new_n237_, keyIn_0_10 );
not g0036 ( new_n238_, N85 );
nand g0037 ( new_n239_, new_n238_, N81 );
not g0038 ( new_n240_, N81 );
nand g0039 ( new_n241_, new_n240_, N85 );
nand g0040 ( new_n242_, new_n239_, new_n241_ );
nand g0041 ( new_n243_, new_n242_, new_n237_ );
nor g0042 ( new_n244_, new_n242_, new_n237_ );
not g0043 ( new_n245_, new_n244_ );
nand g0044 ( new_n246_, new_n245_, new_n243_ );
not g0045 ( new_n247_, N93 );
nand g0046 ( new_n248_, new_n247_, N89 );
not g0047 ( new_n249_, N89 );
nand g0048 ( new_n250_, new_n249_, N93 );
nand g0049 ( new_n251_, new_n248_, new_n250_ );
nand g0050 ( new_n252_, new_n251_, keyIn_0_11 );
not g0051 ( new_n253_, keyIn_0_11 );
not g0052 ( new_n254_, new_n251_ );
nand g0053 ( new_n255_, new_n254_, new_n253_ );
nand g0054 ( new_n256_, new_n255_, new_n252_ );
nand g0055 ( new_n257_, new_n246_, new_n256_ );
not g0056 ( new_n258_, new_n243_ );
nor g0057 ( new_n259_, new_n258_, new_n244_ );
not g0058 ( new_n260_, new_n252_ );
nor g0059 ( new_n261_, new_n251_, keyIn_0_11 );
nor g0060 ( new_n262_, new_n260_, new_n261_ );
nand g0061 ( new_n263_, new_n259_, new_n262_ );
nand g0062 ( new_n264_, new_n263_, new_n257_ );
nand g0063 ( new_n265_, new_n264_, new_n236_ );
not g0064 ( new_n266_, new_n265_ );
nor g0065 ( new_n267_, new_n264_, new_n236_ );
nor g0066 ( new_n268_, new_n266_, new_n267_ );
nand g0067 ( new_n269_, new_n235_, new_n268_ );
not g0068 ( new_n270_, new_n234_ );
nand g0069 ( new_n271_, new_n270_, new_n232_ );
not g0070 ( new_n272_, new_n264_ );
nand g0071 ( new_n273_, new_n272_, keyIn_0_45 );
nand g0072 ( new_n274_, new_n273_, new_n265_ );
nand g0073 ( new_n275_, new_n271_, new_n274_ );
nand g0074 ( new_n276_, new_n269_, new_n275_ );
not g0075 ( new_n277_, new_n276_ );
nand g0076 ( new_n278_, new_n277_, new_n203_ );
nand g0077 ( new_n279_, new_n276_, keyIn_0_60 );
nand g0078 ( new_n280_, new_n278_, new_n279_ );
nand g0079 ( new_n281_, N129, N137 );
nor g0080 ( new_n282_, new_n281_, keyIn_0_16 );
nand g0081 ( new_n283_, new_n281_, keyIn_0_16 );
not g0082 ( new_n284_, new_n283_ );
nor g0083 ( new_n285_, new_n284_, new_n282_ );
not g0084 ( new_n286_, new_n285_ );
nand g0085 ( new_n287_, new_n280_, new_n286_ );
nor g0086 ( new_n288_, new_n276_, keyIn_0_60 );
not g0087 ( new_n289_, new_n279_ );
nor g0088 ( new_n290_, new_n289_, new_n288_ );
nand g0089 ( new_n291_, new_n290_, new_n285_ );
nand g0090 ( new_n292_, new_n291_, new_n287_ );
nand g0091 ( new_n293_, new_n292_, new_n202_ );
nor g0092 ( new_n294_, new_n290_, new_n285_ );
nor g0093 ( new_n295_, new_n280_, new_n286_ );
nor g0094 ( new_n296_, new_n294_, new_n295_ );
nand g0095 ( new_n297_, new_n296_, keyIn_0_64 );
nand g0096 ( new_n298_, new_n297_, new_n293_ );
not g0097 ( new_n299_, N1 );
nor g0098 ( new_n300_, new_n299_, N17 );
not g0099 ( new_n301_, N17 );
nor g0100 ( new_n302_, new_n301_, N1 );
nor g0101 ( new_n303_, new_n300_, new_n302_ );
not g0102 ( new_n304_, new_n303_ );
nand g0103 ( new_n305_, new_n304_, keyIn_0_24 );
not g0104 ( new_n306_, new_n305_ );
nor g0105 ( new_n307_, new_n304_, keyIn_0_24 );
nor g0106 ( new_n308_, new_n306_, new_n307_ );
not g0107 ( new_n309_, N33 );
nor g0108 ( new_n310_, new_n309_, N49 );
not g0109 ( new_n311_, N49 );
nor g0110 ( new_n312_, new_n311_, N33 );
nor g0111 ( new_n313_, new_n310_, new_n312_ );
not g0112 ( new_n314_, new_n313_ );
nand g0113 ( new_n315_, new_n314_, keyIn_0_25 );
not g0114 ( new_n316_, new_n315_ );
nor g0115 ( new_n317_, new_n314_, keyIn_0_25 );
nor g0116 ( new_n318_, new_n316_, new_n317_ );
not g0117 ( new_n319_, new_n318_ );
nor g0118 ( new_n320_, new_n319_, new_n308_ );
nand g0119 ( new_n321_, new_n319_, new_n308_ );
not g0120 ( new_n322_, new_n321_ );
nor g0121 ( new_n323_, new_n322_, new_n320_ );
not g0122 ( new_n324_, new_n323_ );
nand g0123 ( new_n325_, new_n324_, keyIn_0_48 );
not g0124 ( new_n326_, new_n325_ );
nor g0125 ( new_n327_, new_n324_, keyIn_0_48 );
nor g0126 ( new_n328_, new_n326_, new_n327_ );
nand g0127 ( new_n329_, new_n298_, new_n328_ );
not g0128 ( new_n330_, new_n329_ );
nor g0129 ( new_n331_, new_n298_, new_n328_ );
nor g0130 ( new_n332_, new_n330_, new_n331_ );
nand g0131 ( new_n333_, new_n332_, keyIn_0_72 );
not g0132 ( new_n334_, keyIn_0_72 );
not g0133 ( new_n335_, new_n293_ );
nor g0134 ( new_n336_, new_n292_, new_n202_ );
nor g0135 ( new_n337_, new_n335_, new_n336_ );
not g0136 ( new_n338_, new_n328_ );
nand g0137 ( new_n339_, new_n337_, new_n338_ );
nand g0138 ( new_n340_, new_n339_, new_n329_ );
nand g0139 ( new_n341_, new_n340_, new_n334_ );
nand g0140 ( new_n342_, new_n333_, new_n341_ );
not g0141 ( new_n343_, keyIn_0_114 );
not g0142 ( new_n344_, keyIn_0_112 );
not g0143 ( new_n345_, keyIn_0_62 );
not g0144 ( new_n346_, N101 );
nand g0145 ( new_n347_, new_n346_, N97 );
not g0146 ( new_n348_, N97 );
nand g0147 ( new_n349_, new_n348_, N101 );
nand g0148 ( new_n350_, new_n347_, new_n349_ );
nand g0149 ( new_n351_, new_n350_, keyIn_0_12 );
not g0150 ( new_n352_, new_n351_ );
nor g0151 ( new_n353_, new_n350_, keyIn_0_12 );
nor g0152 ( new_n354_, new_n352_, new_n353_ );
not g0153 ( new_n355_, keyIn_0_13 );
not g0154 ( new_n356_, N109 );
nand g0155 ( new_n357_, new_n356_, N105 );
not g0156 ( new_n358_, N105 );
nand g0157 ( new_n359_, new_n358_, N109 );
nand g0158 ( new_n360_, new_n357_, new_n359_ );
nor g0159 ( new_n361_, new_n360_, new_n355_ );
not g0160 ( new_n362_, new_n361_ );
nand g0161 ( new_n363_, new_n360_, new_n355_ );
nand g0162 ( new_n364_, new_n362_, new_n363_ );
nand g0163 ( new_n365_, new_n354_, new_n364_ );
not g0164 ( new_n366_, keyIn_0_12 );
not g0165 ( new_n367_, new_n350_ );
nand g0166 ( new_n368_, new_n367_, new_n366_ );
nand g0167 ( new_n369_, new_n368_, new_n351_ );
not g0168 ( new_n370_, new_n363_ );
nor g0169 ( new_n371_, new_n370_, new_n361_ );
nand g0170 ( new_n372_, new_n371_, new_n369_ );
nand g0171 ( new_n373_, new_n365_, new_n372_ );
nor g0172 ( new_n374_, new_n373_, keyIn_0_46 );
not g0173 ( new_n375_, new_n374_ );
nand g0174 ( new_n376_, new_n373_, keyIn_0_46 );
nand g0175 ( new_n377_, new_n375_, new_n376_ );
nand g0176 ( new_n378_, new_n235_, new_n377_ );
not g0177 ( new_n379_, new_n376_ );
nor g0178 ( new_n380_, new_n379_, new_n374_ );
nand g0179 ( new_n381_, new_n271_, new_n380_ );
nand g0180 ( new_n382_, new_n378_, new_n381_ );
nand g0181 ( new_n383_, new_n382_, new_n345_ );
not g0182 ( new_n384_, new_n382_ );
nand g0183 ( new_n385_, new_n384_, keyIn_0_62 );
nand g0184 ( new_n386_, new_n385_, new_n383_ );
nand g0185 ( new_n387_, N131, N137 );
nor g0186 ( new_n388_, new_n387_, keyIn_0_18 );
nand g0187 ( new_n389_, new_n387_, keyIn_0_18 );
not g0188 ( new_n390_, new_n389_ );
nor g0189 ( new_n391_, new_n390_, new_n388_ );
not g0190 ( new_n392_, new_n391_ );
nand g0191 ( new_n393_, new_n386_, new_n392_ );
not g0192 ( new_n394_, new_n383_ );
nor g0193 ( new_n395_, new_n382_, new_n345_ );
nor g0194 ( new_n396_, new_n394_, new_n395_ );
nand g0195 ( new_n397_, new_n396_, new_n391_ );
nand g0196 ( new_n398_, new_n397_, new_n393_ );
nand g0197 ( new_n399_, new_n398_, keyIn_0_66 );
not g0198 ( new_n400_, keyIn_0_66 );
nor g0199 ( new_n401_, new_n396_, new_n391_ );
nor g0200 ( new_n402_, new_n386_, new_n392_ );
nor g0201 ( new_n403_, new_n401_, new_n402_ );
nand g0202 ( new_n404_, new_n403_, new_n400_ );
nand g0203 ( new_n405_, new_n404_, new_n399_ );
not g0204 ( new_n406_, keyIn_0_50 );
not g0205 ( new_n407_, keyIn_0_28 );
not g0206 ( new_n408_, N9 );
nor g0207 ( new_n409_, new_n408_, N25 );
not g0208 ( new_n410_, N25 );
nor g0209 ( new_n411_, new_n410_, N9 );
nor g0210 ( new_n412_, new_n409_, new_n411_ );
not g0211 ( new_n413_, new_n412_ );
nand g0212 ( new_n414_, new_n413_, new_n407_ );
not g0213 ( new_n415_, new_n414_ );
nor g0214 ( new_n416_, new_n413_, new_n407_ );
nor g0215 ( new_n417_, new_n415_, new_n416_ );
not g0216 ( new_n418_, N41 );
nor g0217 ( new_n419_, new_n418_, N57 );
not g0218 ( new_n420_, N57 );
nor g0219 ( new_n421_, new_n420_, N41 );
nor g0220 ( new_n422_, new_n419_, new_n421_ );
not g0221 ( new_n423_, new_n422_ );
nand g0222 ( new_n424_, new_n423_, keyIn_0_29 );
not g0223 ( new_n425_, new_n424_ );
nor g0224 ( new_n426_, new_n423_, keyIn_0_29 );
nor g0225 ( new_n427_, new_n425_, new_n426_ );
not g0226 ( new_n428_, new_n427_ );
nor g0227 ( new_n429_, new_n428_, new_n417_ );
nand g0228 ( new_n430_, new_n428_, new_n417_ );
not g0229 ( new_n431_, new_n430_ );
nor g0230 ( new_n432_, new_n431_, new_n429_ );
not g0231 ( new_n433_, new_n432_ );
nand g0232 ( new_n434_, new_n433_, new_n406_ );
not g0233 ( new_n435_, new_n434_ );
nor g0234 ( new_n436_, new_n433_, new_n406_ );
nor g0235 ( new_n437_, new_n435_, new_n436_ );
nand g0236 ( new_n438_, new_n405_, new_n437_ );
not g0237 ( new_n439_, new_n438_ );
nor g0238 ( new_n440_, new_n405_, new_n437_ );
nor g0239 ( new_n441_, new_n439_, new_n440_ );
nand g0240 ( new_n442_, new_n441_, keyIn_0_74 );
not g0241 ( new_n443_, keyIn_0_74 );
not g0242 ( new_n444_, new_n399_ );
nor g0243 ( new_n445_, new_n398_, keyIn_0_66 );
nor g0244 ( new_n446_, new_n444_, new_n445_ );
not g0245 ( new_n447_, new_n437_ );
nand g0246 ( new_n448_, new_n446_, new_n447_ );
nand g0247 ( new_n449_, new_n448_, new_n438_ );
nand g0248 ( new_n450_, new_n449_, new_n443_ );
nand g0249 ( new_n451_, new_n442_, new_n450_ );
nor g0250 ( new_n452_, new_n451_, keyIn_0_82 );
not g0251 ( new_n453_, keyIn_0_47 );
not g0252 ( new_n454_, N117 );
nand g0253 ( new_n455_, new_n454_, N113 );
not g0254 ( new_n456_, N113 );
nand g0255 ( new_n457_, new_n456_, N117 );
nand g0256 ( new_n458_, new_n455_, new_n457_ );
nand g0257 ( new_n459_, new_n458_, keyIn_0_14 );
not g0258 ( new_n460_, new_n459_ );
nor g0259 ( new_n461_, new_n458_, keyIn_0_14 );
nor g0260 ( new_n462_, new_n460_, new_n461_ );
not g0261 ( new_n463_, N125 );
nand g0262 ( new_n464_, new_n463_, N121 );
not g0263 ( new_n465_, N121 );
nand g0264 ( new_n466_, new_n465_, N125 );
nand g0265 ( new_n467_, new_n464_, new_n466_ );
nand g0266 ( new_n468_, new_n467_, keyIn_0_15 );
not g0267 ( new_n469_, new_n468_ );
nor g0268 ( new_n470_, new_n467_, keyIn_0_15 );
nor g0269 ( new_n471_, new_n469_, new_n470_ );
nand g0270 ( new_n472_, new_n462_, new_n471_ );
not g0271 ( new_n473_, keyIn_0_14 );
not g0272 ( new_n474_, new_n458_ );
nand g0273 ( new_n475_, new_n474_, new_n473_ );
nand g0274 ( new_n476_, new_n475_, new_n459_ );
not g0275 ( new_n477_, keyIn_0_15 );
not g0276 ( new_n478_, new_n467_ );
nand g0277 ( new_n479_, new_n478_, new_n477_ );
nand g0278 ( new_n480_, new_n479_, new_n468_ );
nand g0279 ( new_n481_, new_n476_, new_n480_ );
nand g0280 ( new_n482_, new_n472_, new_n481_ );
nand g0281 ( new_n483_, new_n482_, new_n453_ );
not g0282 ( new_n484_, new_n483_ );
nor g0283 ( new_n485_, new_n482_, new_n453_ );
nor g0284 ( new_n486_, new_n484_, new_n485_ );
nand g0285 ( new_n487_, new_n268_, new_n486_ );
not g0286 ( new_n488_, new_n482_ );
nand g0287 ( new_n489_, new_n488_, keyIn_0_47 );
nand g0288 ( new_n490_, new_n489_, new_n483_ );
nand g0289 ( new_n491_, new_n274_, new_n490_ );
nand g0290 ( new_n492_, new_n487_, new_n491_ );
not g0291 ( new_n493_, new_n492_ );
nand g0292 ( new_n494_, new_n493_, keyIn_0_63 );
not g0293 ( new_n495_, keyIn_0_63 );
nand g0294 ( new_n496_, new_n492_, new_n495_ );
nand g0295 ( new_n497_, new_n494_, new_n496_ );
nand g0296 ( new_n498_, N132, N137 );
nor g0297 ( new_n499_, new_n498_, keyIn_0_19 );
nand g0298 ( new_n500_, new_n498_, keyIn_0_19 );
not g0299 ( new_n501_, new_n500_ );
nor g0300 ( new_n502_, new_n501_, new_n499_ );
not g0301 ( new_n503_, new_n502_ );
nand g0302 ( new_n504_, new_n497_, new_n503_ );
nor g0303 ( new_n505_, new_n492_, new_n495_ );
not g0304 ( new_n506_, new_n496_ );
nor g0305 ( new_n507_, new_n506_, new_n505_ );
nand g0306 ( new_n508_, new_n507_, new_n502_ );
nand g0307 ( new_n509_, new_n508_, new_n504_ );
nand g0308 ( new_n510_, new_n509_, keyIn_0_67 );
not g0309 ( new_n511_, keyIn_0_67 );
nor g0310 ( new_n512_, new_n507_, new_n502_ );
nor g0311 ( new_n513_, new_n497_, new_n503_ );
nor g0312 ( new_n514_, new_n512_, new_n513_ );
nand g0313 ( new_n515_, new_n514_, new_n511_ );
nand g0314 ( new_n516_, new_n515_, new_n510_ );
not g0315 ( new_n517_, keyIn_0_51 );
not g0316 ( new_n518_, N13 );
nor g0317 ( new_n519_, new_n518_, N29 );
not g0318 ( new_n520_, N29 );
nor g0319 ( new_n521_, new_n520_, N13 );
nor g0320 ( new_n522_, new_n519_, new_n521_ );
not g0321 ( new_n523_, new_n522_ );
nand g0322 ( new_n524_, new_n523_, keyIn_0_30 );
not g0323 ( new_n525_, new_n524_ );
nor g0324 ( new_n526_, new_n523_, keyIn_0_30 );
nor g0325 ( new_n527_, new_n525_, new_n526_ );
not g0326 ( new_n528_, new_n527_ );
not g0327 ( new_n529_, keyIn_0_31 );
not g0328 ( new_n530_, N45 );
nor g0329 ( new_n531_, new_n530_, N61 );
not g0330 ( new_n532_, N61 );
nor g0331 ( new_n533_, new_n532_, N45 );
nor g0332 ( new_n534_, new_n531_, new_n533_ );
not g0333 ( new_n535_, new_n534_ );
nand g0334 ( new_n536_, new_n535_, new_n529_ );
not g0335 ( new_n537_, new_n536_ );
nor g0336 ( new_n538_, new_n535_, new_n529_ );
nor g0337 ( new_n539_, new_n537_, new_n538_ );
not g0338 ( new_n540_, new_n539_ );
nor g0339 ( new_n541_, new_n528_, new_n540_ );
nor g0340 ( new_n542_, new_n527_, new_n539_ );
nor g0341 ( new_n543_, new_n541_, new_n542_ );
not g0342 ( new_n544_, new_n543_ );
nand g0343 ( new_n545_, new_n544_, new_n517_ );
not g0344 ( new_n546_, new_n545_ );
nor g0345 ( new_n547_, new_n544_, new_n517_ );
nor g0346 ( new_n548_, new_n546_, new_n547_ );
nand g0347 ( new_n549_, new_n516_, new_n548_ );
nor g0348 ( new_n550_, new_n514_, new_n511_ );
nor g0349 ( new_n551_, new_n509_, keyIn_0_67 );
nor g0350 ( new_n552_, new_n550_, new_n551_ );
not g0351 ( new_n553_, new_n548_ );
nand g0352 ( new_n554_, new_n552_, new_n553_ );
nand g0353 ( new_n555_, new_n554_, new_n549_ );
nor g0354 ( new_n556_, new_n555_, keyIn_0_75 );
not g0355 ( new_n557_, keyIn_0_75 );
nor g0356 ( new_n558_, new_n552_, new_n553_ );
nor g0357 ( new_n559_, new_n516_, new_n548_ );
nor g0358 ( new_n560_, new_n558_, new_n559_ );
nor g0359 ( new_n561_, new_n560_, new_n557_ );
nor g0360 ( new_n562_, new_n561_, new_n556_ );
nand g0361 ( new_n563_, new_n451_, keyIn_0_82 );
nand g0362 ( new_n564_, new_n563_, new_n562_ );
nor g0363 ( new_n565_, new_n564_, new_n452_ );
not g0364 ( new_n566_, keyIn_0_81 );
not g0365 ( new_n567_, keyIn_0_65 );
not g0366 ( new_n568_, keyIn_0_61 );
nand g0367 ( new_n569_, new_n486_, new_n377_ );
nand g0368 ( new_n570_, new_n380_, new_n490_ );
nand g0369 ( new_n571_, new_n569_, new_n570_ );
nand g0370 ( new_n572_, new_n571_, new_n568_ );
not g0371 ( new_n573_, new_n571_ );
nand g0372 ( new_n574_, new_n573_, keyIn_0_61 );
nand g0373 ( new_n575_, new_n574_, new_n572_ );
nand g0374 ( new_n576_, N130, N137 );
nor g0375 ( new_n577_, new_n576_, keyIn_0_17 );
nand g0376 ( new_n578_, new_n576_, keyIn_0_17 );
not g0377 ( new_n579_, new_n578_ );
nor g0378 ( new_n580_, new_n579_, new_n577_ );
not g0379 ( new_n581_, new_n580_ );
nand g0380 ( new_n582_, new_n575_, new_n581_ );
not g0381 ( new_n583_, new_n572_ );
nor g0382 ( new_n584_, new_n571_, new_n568_ );
nor g0383 ( new_n585_, new_n583_, new_n584_ );
nand g0384 ( new_n586_, new_n585_, new_n580_ );
nand g0385 ( new_n587_, new_n586_, new_n582_ );
nand g0386 ( new_n588_, new_n587_, new_n567_ );
nor g0387 ( new_n589_, new_n585_, new_n580_ );
nor g0388 ( new_n590_, new_n575_, new_n581_ );
nor g0389 ( new_n591_, new_n589_, new_n590_ );
nand g0390 ( new_n592_, new_n591_, keyIn_0_65 );
nand g0391 ( new_n593_, new_n592_, new_n588_ );
not g0392 ( new_n594_, keyIn_0_49 );
not g0393 ( new_n595_, keyIn_0_26 );
not g0394 ( new_n596_, N5 );
nor g0395 ( new_n597_, new_n596_, N21 );
not g0396 ( new_n598_, N21 );
nor g0397 ( new_n599_, new_n598_, N5 );
nor g0398 ( new_n600_, new_n597_, new_n599_ );
not g0399 ( new_n601_, new_n600_ );
nand g0400 ( new_n602_, new_n601_, new_n595_ );
not g0401 ( new_n603_, new_n602_ );
nor g0402 ( new_n604_, new_n601_, new_n595_ );
nor g0403 ( new_n605_, new_n603_, new_n604_ );
not g0404 ( new_n606_, keyIn_0_27 );
not g0405 ( new_n607_, N37 );
nor g0406 ( new_n608_, new_n607_, N53 );
not g0407 ( new_n609_, N53 );
nor g0408 ( new_n610_, new_n609_, N37 );
nor g0409 ( new_n611_, new_n608_, new_n610_ );
not g0410 ( new_n612_, new_n611_ );
nand g0411 ( new_n613_, new_n612_, new_n606_ );
not g0412 ( new_n614_, new_n613_ );
nor g0413 ( new_n615_, new_n612_, new_n606_ );
nor g0414 ( new_n616_, new_n614_, new_n615_ );
not g0415 ( new_n617_, new_n616_ );
nor g0416 ( new_n618_, new_n617_, new_n605_ );
nand g0417 ( new_n619_, new_n617_, new_n605_ );
not g0418 ( new_n620_, new_n619_ );
nor g0419 ( new_n621_, new_n620_, new_n618_ );
not g0420 ( new_n622_, new_n621_ );
nand g0421 ( new_n623_, new_n622_, new_n594_ );
not g0422 ( new_n624_, new_n623_ );
nor g0423 ( new_n625_, new_n622_, new_n594_ );
nor g0424 ( new_n626_, new_n624_, new_n625_ );
nand g0425 ( new_n627_, new_n593_, new_n626_ );
not g0426 ( new_n628_, new_n588_ );
nor g0427 ( new_n629_, new_n587_, new_n567_ );
nor g0428 ( new_n630_, new_n628_, new_n629_ );
not g0429 ( new_n631_, new_n626_ );
nand g0430 ( new_n632_, new_n630_, new_n631_ );
nand g0431 ( new_n633_, new_n632_, new_n627_ );
nand g0432 ( new_n634_, new_n633_, keyIn_0_73 );
not g0433 ( new_n635_, new_n634_ );
nor g0434 ( new_n636_, new_n633_, keyIn_0_73 );
nor g0435 ( new_n637_, new_n635_, new_n636_ );
nand g0436 ( new_n638_, new_n637_, new_n566_ );
not g0437 ( new_n639_, keyIn_0_73 );
not g0438 ( new_n640_, new_n627_ );
nor g0439 ( new_n641_, new_n593_, new_n626_ );
nor g0440 ( new_n642_, new_n640_, new_n641_ );
nand g0441 ( new_n643_, new_n642_, new_n639_ );
nand g0442 ( new_n644_, new_n643_, new_n634_ );
nand g0443 ( new_n645_, new_n644_, keyIn_0_81 );
nand g0444 ( new_n646_, new_n638_, new_n645_ );
not g0445 ( new_n647_, keyIn_0_80 );
nor g0446 ( new_n648_, new_n340_, new_n334_ );
not g0447 ( new_n649_, new_n341_ );
nor g0448 ( new_n650_, new_n649_, new_n648_ );
nand g0449 ( new_n651_, new_n650_, new_n647_ );
nand g0450 ( new_n652_, new_n342_, keyIn_0_80 );
nand g0451 ( new_n653_, new_n651_, new_n652_ );
nand g0452 ( new_n654_, new_n653_, new_n646_ );
not g0453 ( new_n655_, new_n654_ );
nand g0454 ( new_n656_, new_n655_, new_n565_ );
nand g0455 ( new_n657_, new_n656_, keyIn_0_104 );
not g0456 ( new_n658_, keyIn_0_104 );
not g0457 ( new_n659_, new_n565_ );
nor g0458 ( new_n660_, new_n659_, new_n654_ );
nand g0459 ( new_n661_, new_n660_, new_n658_ );
nand g0460 ( new_n662_, new_n657_, new_n661_ );
nor g0461 ( new_n663_, new_n644_, keyIn_0_84 );
nor g0462 ( new_n664_, new_n449_, new_n443_ );
not g0463 ( new_n665_, new_n450_ );
nor g0464 ( new_n666_, new_n665_, new_n664_ );
nand g0465 ( new_n667_, new_n644_, keyIn_0_84 );
nand g0466 ( new_n668_, new_n667_, new_n666_ );
nor g0467 ( new_n669_, new_n668_, new_n663_ );
nand g0468 ( new_n670_, new_n650_, keyIn_0_83 );
not g0469 ( new_n671_, keyIn_0_83 );
nand g0470 ( new_n672_, new_n342_, new_n671_ );
nand g0471 ( new_n673_, new_n670_, new_n672_ );
not g0472 ( new_n674_, keyIn_0_85 );
nand g0473 ( new_n675_, new_n562_, new_n674_ );
nand g0474 ( new_n676_, new_n560_, new_n557_ );
nand g0475 ( new_n677_, new_n555_, keyIn_0_75 );
nand g0476 ( new_n678_, new_n676_, new_n677_ );
nand g0477 ( new_n679_, new_n678_, keyIn_0_85 );
nand g0478 ( new_n680_, new_n675_, new_n679_ );
nand g0479 ( new_n681_, new_n673_, new_n680_ );
not g0480 ( new_n682_, new_n681_ );
nand g0481 ( new_n683_, new_n682_, new_n669_ );
nand g0482 ( new_n684_, new_n683_, keyIn_0_105 );
not g0483 ( new_n685_, keyIn_0_105 );
not g0484 ( new_n686_, new_n669_ );
nor g0485 ( new_n687_, new_n686_, new_n681_ );
nand g0486 ( new_n688_, new_n687_, new_n685_ );
nand g0487 ( new_n689_, new_n684_, new_n688_ );
nor g0488 ( new_n690_, new_n662_, new_n689_ );
nor g0489 ( new_n691_, new_n650_, keyIn_0_86 );
not g0490 ( new_n692_, new_n691_ );
nor g0491 ( new_n693_, new_n451_, keyIn_0_87 );
nand g0492 ( new_n694_, new_n451_, keyIn_0_87 );
not g0493 ( new_n695_, new_n694_ );
nor g0494 ( new_n696_, new_n695_, new_n693_ );
nand g0495 ( new_n697_, new_n696_, new_n692_ );
not g0496 ( new_n698_, keyIn_0_86 );
nor g0497 ( new_n699_, new_n342_, new_n698_ );
nor g0498 ( new_n700_, new_n699_, new_n644_ );
nor g0499 ( new_n701_, new_n678_, keyIn_0_88 );
nand g0500 ( new_n702_, new_n678_, keyIn_0_88 );
not g0501 ( new_n703_, new_n702_ );
nor g0502 ( new_n704_, new_n703_, new_n701_ );
nand g0503 ( new_n705_, new_n704_, new_n700_ );
nor g0504 ( new_n706_, new_n697_, new_n705_ );
nand g0505 ( new_n707_, new_n706_, keyIn_0_106 );
not g0506 ( new_n708_, keyIn_0_106 );
not g0507 ( new_n709_, keyIn_0_87 );
nand g0508 ( new_n710_, new_n666_, new_n709_ );
nand g0509 ( new_n711_, new_n710_, new_n694_ );
nor g0510 ( new_n712_, new_n711_, new_n691_ );
nand g0511 ( new_n713_, new_n650_, keyIn_0_86 );
nand g0512 ( new_n714_, new_n713_, new_n637_ );
not g0513 ( new_n715_, keyIn_0_88 );
nand g0514 ( new_n716_, new_n562_, new_n715_ );
nand g0515 ( new_n717_, new_n716_, new_n702_ );
nor g0516 ( new_n718_, new_n714_, new_n717_ );
nand g0517 ( new_n719_, new_n718_, new_n712_ );
nand g0518 ( new_n720_, new_n719_, new_n708_ );
nand g0519 ( new_n721_, new_n707_, new_n720_ );
not g0520 ( new_n722_, keyIn_0_107 );
nor g0521 ( new_n723_, new_n451_, keyIn_0_90 );
not g0522 ( new_n724_, keyIn_0_89 );
nand g0523 ( new_n725_, new_n644_, new_n724_ );
nand g0524 ( new_n726_, new_n637_, keyIn_0_89 );
nand g0525 ( new_n727_, new_n726_, new_n725_ );
nor g0526 ( new_n728_, new_n727_, new_n723_ );
nand g0527 ( new_n729_, new_n451_, keyIn_0_90 );
nand g0528 ( new_n730_, new_n729_, new_n650_ );
nand g0529 ( new_n731_, new_n562_, keyIn_0_91 );
not g0530 ( new_n732_, keyIn_0_91 );
nand g0531 ( new_n733_, new_n678_, new_n732_ );
nand g0532 ( new_n734_, new_n731_, new_n733_ );
nor g0533 ( new_n735_, new_n734_, new_n730_ );
nand g0534 ( new_n736_, new_n728_, new_n735_ );
nand g0535 ( new_n737_, new_n736_, new_n722_ );
not g0536 ( new_n738_, new_n736_ );
nand g0537 ( new_n739_, new_n738_, keyIn_0_107 );
nand g0538 ( new_n740_, new_n739_, new_n737_ );
nor g0539 ( new_n741_, new_n740_, new_n721_ );
nand g0540 ( new_n742_, new_n690_, new_n741_ );
nor g0541 ( new_n743_, new_n742_, new_n344_ );
nor g0542 ( new_n744_, new_n660_, new_n658_ );
nor g0543 ( new_n745_, new_n656_, keyIn_0_104 );
nor g0544 ( new_n746_, new_n745_, new_n744_ );
nor g0545 ( new_n747_, new_n687_, new_n685_ );
nor g0546 ( new_n748_, new_n683_, keyIn_0_105 );
nor g0547 ( new_n749_, new_n748_, new_n747_ );
nand g0548 ( new_n750_, new_n746_, new_n749_ );
nor g0549 ( new_n751_, new_n719_, new_n708_ );
nor g0550 ( new_n752_, new_n706_, keyIn_0_106 );
nor g0551 ( new_n753_, new_n752_, new_n751_ );
not g0552 ( new_n754_, new_n737_ );
nor g0553 ( new_n755_, new_n736_, new_n722_ );
nor g0554 ( new_n756_, new_n754_, new_n755_ );
nand g0555 ( new_n757_, new_n753_, new_n756_ );
nor g0556 ( new_n758_, new_n750_, new_n757_ );
nor g0557 ( new_n759_, new_n758_, keyIn_0_112 );
nor g0558 ( new_n760_, new_n759_, new_n743_ );
not g0559 ( new_n761_, keyIn_0_56 );
nand g0560 ( new_n762_, new_n596_, N1 );
nand g0561 ( new_n763_, new_n299_, N5 );
nand g0562 ( new_n764_, new_n762_, new_n763_ );
nand g0563 ( new_n765_, new_n764_, keyIn_0_0 );
nor g0564 ( new_n766_, new_n764_, keyIn_0_0 );
not g0565 ( new_n767_, new_n766_ );
nand g0566 ( new_n768_, new_n767_, new_n765_ );
not g0567 ( new_n769_, keyIn_0_1 );
nand g0568 ( new_n770_, new_n518_, N9 );
nand g0569 ( new_n771_, new_n408_, N13 );
nand g0570 ( new_n772_, new_n770_, new_n771_ );
nor g0571 ( new_n773_, new_n772_, new_n769_ );
nand g0572 ( new_n774_, new_n772_, new_n769_ );
not g0573 ( new_n775_, new_n774_ );
nor g0574 ( new_n776_, new_n775_, new_n773_ );
nand g0575 ( new_n777_, new_n776_, new_n768_ );
not g0576 ( new_n778_, new_n765_ );
nor g0577 ( new_n779_, new_n778_, new_n766_ );
not g0578 ( new_n780_, new_n772_ );
nand g0579 ( new_n781_, new_n780_, keyIn_0_1 );
nand g0580 ( new_n782_, new_n781_, new_n774_ );
nand g0581 ( new_n783_, new_n779_, new_n782_ );
nand g0582 ( new_n784_, new_n777_, new_n783_ );
nand g0583 ( new_n785_, new_n784_, keyIn_0_40 );
not g0584 ( new_n786_, new_n785_ );
nor g0585 ( new_n787_, new_n784_, keyIn_0_40 );
nor g0586 ( new_n788_, new_n786_, new_n787_ );
not g0587 ( new_n789_, keyIn_0_41 );
nand g0588 ( new_n790_, new_n598_, N17 );
nand g0589 ( new_n791_, new_n301_, N21 );
nand g0590 ( new_n792_, new_n790_, new_n791_ );
nand g0591 ( new_n793_, new_n792_, keyIn_0_2 );
nor g0592 ( new_n794_, new_n792_, keyIn_0_2 );
not g0593 ( new_n795_, new_n794_ );
nand g0594 ( new_n796_, new_n795_, new_n793_ );
nand g0595 ( new_n797_, new_n520_, N25 );
nand g0596 ( new_n798_, new_n410_, N29 );
nand g0597 ( new_n799_, new_n797_, new_n798_ );
nand g0598 ( new_n800_, new_n799_, keyIn_0_3 );
not g0599 ( new_n801_, keyIn_0_3 );
not g0600 ( new_n802_, new_n799_ );
nand g0601 ( new_n803_, new_n802_, new_n801_ );
nand g0602 ( new_n804_, new_n803_, new_n800_ );
nand g0603 ( new_n805_, new_n796_, new_n804_ );
not g0604 ( new_n806_, new_n793_ );
nor g0605 ( new_n807_, new_n806_, new_n794_ );
not g0606 ( new_n808_, new_n800_ );
nor g0607 ( new_n809_, new_n799_, keyIn_0_3 );
nor g0608 ( new_n810_, new_n808_, new_n809_ );
nand g0609 ( new_n811_, new_n807_, new_n810_ );
nand g0610 ( new_n812_, new_n811_, new_n805_ );
nand g0611 ( new_n813_, new_n812_, new_n789_ );
not g0612 ( new_n814_, new_n813_ );
nor g0613 ( new_n815_, new_n812_, new_n789_ );
nor g0614 ( new_n816_, new_n814_, new_n815_ );
nand g0615 ( new_n817_, new_n788_, new_n816_ );
not g0616 ( new_n818_, new_n787_ );
nand g0617 ( new_n819_, new_n818_, new_n785_ );
not g0618 ( new_n820_, new_n812_ );
nand g0619 ( new_n821_, new_n820_, keyIn_0_41 );
nand g0620 ( new_n822_, new_n821_, new_n813_ );
nand g0621 ( new_n823_, new_n819_, new_n822_ );
nand g0622 ( new_n824_, new_n817_, new_n823_ );
not g0623 ( new_n825_, new_n824_ );
nand g0624 ( new_n826_, new_n825_, new_n761_ );
nand g0625 ( new_n827_, new_n824_, keyIn_0_56 );
nand g0626 ( new_n828_, new_n826_, new_n827_ );
nand g0627 ( new_n829_, N133, N137 );
nor g0628 ( new_n830_, new_n829_, keyIn_0_20 );
nand g0629 ( new_n831_, new_n829_, keyIn_0_20 );
not g0630 ( new_n832_, new_n831_ );
nor g0631 ( new_n833_, new_n832_, new_n830_ );
not g0632 ( new_n834_, new_n833_ );
nand g0633 ( new_n835_, new_n828_, new_n834_ );
nor g0634 ( new_n836_, new_n824_, keyIn_0_56 );
not g0635 ( new_n837_, new_n827_ );
nor g0636 ( new_n838_, new_n837_, new_n836_ );
nand g0637 ( new_n839_, new_n838_, new_n833_ );
nand g0638 ( new_n840_, new_n839_, new_n835_ );
nand g0639 ( new_n841_, new_n840_, keyIn_0_68 );
not g0640 ( new_n842_, keyIn_0_68 );
nor g0641 ( new_n843_, new_n838_, new_n833_ );
nor g0642 ( new_n844_, new_n828_, new_n834_ );
nor g0643 ( new_n845_, new_n843_, new_n844_ );
nand g0644 ( new_n846_, new_n845_, new_n842_ );
nand g0645 ( new_n847_, new_n846_, new_n841_ );
not g0646 ( new_n848_, keyIn_0_52 );
nor g0647 ( new_n849_, new_n208_, N81 );
nor g0648 ( new_n850_, new_n240_, N65 );
nor g0649 ( new_n851_, new_n849_, new_n850_ );
not g0650 ( new_n852_, new_n851_ );
nand g0651 ( new_n853_, new_n852_, keyIn_0_32 );
not g0652 ( new_n854_, new_n853_ );
nor g0653 ( new_n855_, new_n852_, keyIn_0_32 );
nor g0654 ( new_n856_, new_n854_, new_n855_ );
not g0655 ( new_n857_, new_n856_ );
nor g0656 ( new_n858_, new_n348_, N113 );
nor g0657 ( new_n859_, new_n456_, N97 );
nor g0658 ( new_n860_, new_n858_, new_n859_ );
not g0659 ( new_n861_, new_n860_ );
nand g0660 ( new_n862_, new_n861_, keyIn_0_33 );
not g0661 ( new_n863_, new_n862_ );
nor g0662 ( new_n864_, new_n861_, keyIn_0_33 );
nor g0663 ( new_n865_, new_n863_, new_n864_ );
not g0664 ( new_n866_, new_n865_ );
nor g0665 ( new_n867_, new_n857_, new_n866_ );
nor g0666 ( new_n868_, new_n856_, new_n865_ );
nor g0667 ( new_n869_, new_n867_, new_n868_ );
not g0668 ( new_n870_, new_n869_ );
nand g0669 ( new_n871_, new_n870_, new_n848_ );
not g0670 ( new_n872_, new_n871_ );
nor g0671 ( new_n873_, new_n870_, new_n848_ );
nor g0672 ( new_n874_, new_n872_, new_n873_ );
nand g0673 ( new_n875_, new_n847_, new_n874_ );
not g0674 ( new_n876_, new_n875_ );
nor g0675 ( new_n877_, new_n847_, new_n874_ );
nor g0676 ( new_n878_, new_n876_, new_n877_ );
nor g0677 ( new_n879_, new_n878_, keyIn_0_76 );
not g0678 ( new_n880_, keyIn_0_76 );
not g0679 ( new_n881_, new_n841_ );
nor g0680 ( new_n882_, new_n840_, keyIn_0_68 );
nor g0681 ( new_n883_, new_n881_, new_n882_ );
not g0682 ( new_n884_, new_n874_ );
nand g0683 ( new_n885_, new_n883_, new_n884_ );
nand g0684 ( new_n886_, new_n885_, new_n875_ );
nor g0685 ( new_n887_, new_n886_, new_n880_ );
nor g0686 ( new_n888_, new_n879_, new_n887_ );
not g0687 ( new_n889_, keyIn_0_77 );
not g0688 ( new_n890_, keyIn_0_57 );
not g0689 ( new_n891_, keyIn_0_42 );
nand g0690 ( new_n892_, new_n530_, N41 );
nand g0691 ( new_n893_, new_n418_, N45 );
nand g0692 ( new_n894_, new_n892_, new_n893_ );
nand g0693 ( new_n895_, new_n894_, keyIn_0_5 );
nor g0694 ( new_n896_, new_n894_, keyIn_0_5 );
not g0695 ( new_n897_, new_n896_ );
nand g0696 ( new_n898_, new_n897_, new_n895_ );
nand g0697 ( new_n899_, new_n607_, N33 );
nand g0698 ( new_n900_, new_n309_, N37 );
nand g0699 ( new_n901_, new_n899_, new_n900_ );
nor g0700 ( new_n902_, new_n901_, keyIn_0_4 );
nand g0701 ( new_n903_, new_n901_, keyIn_0_4 );
not g0702 ( new_n904_, new_n903_ );
nor g0703 ( new_n905_, new_n904_, new_n902_ );
nand g0704 ( new_n906_, new_n905_, new_n898_ );
not g0705 ( new_n907_, new_n895_ );
nor g0706 ( new_n908_, new_n907_, new_n896_ );
not g0707 ( new_n909_, new_n902_ );
nand g0708 ( new_n910_, new_n909_, new_n903_ );
nand g0709 ( new_n911_, new_n908_, new_n910_ );
nand g0710 ( new_n912_, new_n906_, new_n911_ );
nand g0711 ( new_n913_, new_n912_, new_n891_ );
not g0712 ( new_n914_, new_n913_ );
nor g0713 ( new_n915_, new_n912_, new_n891_ );
nor g0714 ( new_n916_, new_n914_, new_n915_ );
nand g0715 ( new_n917_, new_n532_, N57 );
nand g0716 ( new_n918_, new_n420_, N61 );
nand g0717 ( new_n919_, new_n917_, new_n918_ );
nand g0718 ( new_n920_, new_n919_, keyIn_0_7 );
nor g0719 ( new_n921_, new_n919_, keyIn_0_7 );
not g0720 ( new_n922_, new_n921_ );
nand g0721 ( new_n923_, new_n922_, new_n920_ );
nand g0722 ( new_n924_, new_n609_, N49 );
nand g0723 ( new_n925_, new_n311_, N53 );
nand g0724 ( new_n926_, new_n924_, new_n925_ );
nor g0725 ( new_n927_, new_n926_, keyIn_0_6 );
nand g0726 ( new_n928_, new_n926_, keyIn_0_6 );
not g0727 ( new_n929_, new_n928_ );
nor g0728 ( new_n930_, new_n929_, new_n927_ );
nand g0729 ( new_n931_, new_n930_, new_n923_ );
not g0730 ( new_n932_, new_n920_ );
nor g0731 ( new_n933_, new_n932_, new_n921_ );
not g0732 ( new_n934_, keyIn_0_6 );
not g0733 ( new_n935_, new_n926_ );
nand g0734 ( new_n936_, new_n935_, new_n934_ );
nand g0735 ( new_n937_, new_n936_, new_n928_ );
nand g0736 ( new_n938_, new_n933_, new_n937_ );
nand g0737 ( new_n939_, new_n931_, new_n938_ );
nand g0738 ( new_n940_, new_n939_, keyIn_0_43 );
not g0739 ( new_n941_, new_n940_ );
nor g0740 ( new_n942_, new_n939_, keyIn_0_43 );
nor g0741 ( new_n943_, new_n941_, new_n942_ );
nand g0742 ( new_n944_, new_n916_, new_n943_ );
not g0743 ( new_n945_, new_n912_ );
nand g0744 ( new_n946_, new_n945_, keyIn_0_42 );
nand g0745 ( new_n947_, new_n946_, new_n913_ );
not g0746 ( new_n948_, keyIn_0_43 );
not g0747 ( new_n949_, new_n939_ );
nand g0748 ( new_n950_, new_n949_, new_n948_ );
nand g0749 ( new_n951_, new_n950_, new_n940_ );
nand g0750 ( new_n952_, new_n947_, new_n951_ );
nand g0751 ( new_n953_, new_n944_, new_n952_ );
nor g0752 ( new_n954_, new_n953_, new_n890_ );
nand g0753 ( new_n955_, new_n953_, new_n890_ );
not g0754 ( new_n956_, new_n955_ );
nor g0755 ( new_n957_, new_n956_, new_n954_ );
nand g0756 ( new_n958_, N134, N137 );
nor g0757 ( new_n959_, new_n958_, keyIn_0_21 );
nand g0758 ( new_n960_, new_n958_, keyIn_0_21 );
not g0759 ( new_n961_, new_n960_ );
nor g0760 ( new_n962_, new_n961_, new_n959_ );
nor g0761 ( new_n963_, new_n957_, new_n962_ );
not g0762 ( new_n964_, new_n953_ );
nand g0763 ( new_n965_, new_n964_, keyIn_0_57 );
nand g0764 ( new_n966_, new_n965_, new_n955_ );
not g0765 ( new_n967_, new_n962_ );
nor g0766 ( new_n968_, new_n966_, new_n967_ );
nor g0767 ( new_n969_, new_n963_, new_n968_ );
nor g0768 ( new_n970_, new_n969_, keyIn_0_69 );
not g0769 ( new_n971_, keyIn_0_69 );
nand g0770 ( new_n972_, new_n966_, new_n967_ );
nand g0771 ( new_n973_, new_n957_, new_n962_ );
nand g0772 ( new_n974_, new_n973_, new_n972_ );
nor g0773 ( new_n975_, new_n974_, new_n971_ );
nor g0774 ( new_n976_, new_n970_, new_n975_ );
not g0775 ( new_n977_, keyIn_0_53 );
not g0776 ( new_n978_, keyIn_0_34 );
nor g0777 ( new_n979_, new_n206_, N85 );
nor g0778 ( new_n980_, new_n238_, N69 );
nor g0779 ( new_n981_, new_n979_, new_n980_ );
not g0780 ( new_n982_, new_n981_ );
nand g0781 ( new_n983_, new_n982_, new_n978_ );
not g0782 ( new_n984_, new_n983_ );
nor g0783 ( new_n985_, new_n982_, new_n978_ );
nor g0784 ( new_n986_, new_n984_, new_n985_ );
not g0785 ( new_n987_, new_n986_ );
not g0786 ( new_n988_, keyIn_0_35 );
nor g0787 ( new_n989_, new_n346_, N117 );
nor g0788 ( new_n990_, new_n454_, N101 );
nor g0789 ( new_n991_, new_n989_, new_n990_ );
not g0790 ( new_n992_, new_n991_ );
nand g0791 ( new_n993_, new_n992_, new_n988_ );
not g0792 ( new_n994_, new_n993_ );
nor g0793 ( new_n995_, new_n992_, new_n988_ );
nor g0794 ( new_n996_, new_n994_, new_n995_ );
not g0795 ( new_n997_, new_n996_ );
nor g0796 ( new_n998_, new_n987_, new_n997_ );
nor g0797 ( new_n999_, new_n986_, new_n996_ );
nor g0798 ( new_n1000_, new_n998_, new_n999_ );
not g0799 ( new_n1001_, new_n1000_ );
nand g0800 ( new_n1002_, new_n1001_, new_n977_ );
not g0801 ( new_n1003_, new_n1002_ );
nor g0802 ( new_n1004_, new_n1001_, new_n977_ );
nor g0803 ( new_n1005_, new_n1003_, new_n1004_ );
nor g0804 ( new_n1006_, new_n976_, new_n1005_ );
nand g0805 ( new_n1007_, new_n974_, new_n971_ );
nand g0806 ( new_n1008_, new_n969_, keyIn_0_69 );
nand g0807 ( new_n1009_, new_n1008_, new_n1007_ );
not g0808 ( new_n1010_, new_n1005_ );
nor g0809 ( new_n1011_, new_n1009_, new_n1010_ );
nor g0810 ( new_n1012_, new_n1006_, new_n1011_ );
nand g0811 ( new_n1013_, new_n1012_, new_n889_ );
nand g0812 ( new_n1014_, new_n1009_, new_n1010_ );
nand g0813 ( new_n1015_, new_n976_, new_n1005_ );
nand g0814 ( new_n1016_, new_n1015_, new_n1014_ );
nand g0815 ( new_n1017_, new_n1016_, keyIn_0_77 );
nand g0816 ( new_n1018_, new_n1013_, new_n1017_ );
nor g0817 ( new_n1019_, new_n888_, new_n1018_ );
not g0818 ( new_n1020_, new_n1019_ );
not g0819 ( new_n1021_, keyIn_0_78 );
not g0820 ( new_n1022_, keyIn_0_70 );
nand g0821 ( new_n1023_, new_n916_, new_n819_ );
nand g0822 ( new_n1024_, new_n788_, new_n947_ );
nand g0823 ( new_n1025_, new_n1023_, new_n1024_ );
nand g0824 ( new_n1026_, new_n1025_, keyIn_0_58 );
not g0825 ( new_n1027_, keyIn_0_58 );
not g0826 ( new_n1028_, new_n1025_ );
nand g0827 ( new_n1029_, new_n1028_, new_n1027_ );
nand g0828 ( new_n1030_, new_n1029_, new_n1026_ );
nand g0829 ( new_n1031_, N135, N137 );
nor g0830 ( new_n1032_, new_n1031_, keyIn_0_22 );
nand g0831 ( new_n1033_, new_n1031_, keyIn_0_22 );
not g0832 ( new_n1034_, new_n1033_ );
nor g0833 ( new_n1035_, new_n1034_, new_n1032_ );
not g0834 ( new_n1036_, new_n1035_ );
nand g0835 ( new_n1037_, new_n1030_, new_n1036_ );
not g0836 ( new_n1038_, new_n1026_ );
nor g0837 ( new_n1039_, new_n1025_, keyIn_0_58 );
nor g0838 ( new_n1040_, new_n1038_, new_n1039_ );
nand g0839 ( new_n1041_, new_n1040_, new_n1035_ );
nand g0840 ( new_n1042_, new_n1041_, new_n1037_ );
nand g0841 ( new_n1043_, new_n1042_, new_n1022_ );
nor g0842 ( new_n1044_, new_n1040_, new_n1035_ );
nor g0843 ( new_n1045_, new_n1030_, new_n1036_ );
nor g0844 ( new_n1046_, new_n1044_, new_n1045_ );
nand g0845 ( new_n1047_, new_n1046_, keyIn_0_70 );
nand g0846 ( new_n1048_, new_n1047_, new_n1043_ );
nor g0847 ( new_n1049_, new_n218_, N89 );
nor g0848 ( new_n1050_, new_n249_, N73 );
nor g0849 ( new_n1051_, new_n1049_, new_n1050_ );
not g0850 ( new_n1052_, new_n1051_ );
nand g0851 ( new_n1053_, new_n1052_, keyIn_0_36 );
not g0852 ( new_n1054_, new_n1053_ );
nor g0853 ( new_n1055_, new_n1052_, keyIn_0_36 );
nor g0854 ( new_n1056_, new_n1054_, new_n1055_ );
not g0855 ( new_n1057_, new_n1056_ );
nor g0856 ( new_n1058_, new_n358_, N121 );
nor g0857 ( new_n1059_, new_n465_, N105 );
nor g0858 ( new_n1060_, new_n1058_, new_n1059_ );
not g0859 ( new_n1061_, new_n1060_ );
nand g0860 ( new_n1062_, new_n1061_, keyIn_0_37 );
not g0861 ( new_n1063_, new_n1062_ );
nor g0862 ( new_n1064_, new_n1061_, keyIn_0_37 );
nor g0863 ( new_n1065_, new_n1063_, new_n1064_ );
not g0864 ( new_n1066_, new_n1065_ );
nor g0865 ( new_n1067_, new_n1057_, new_n1066_ );
nor g0866 ( new_n1068_, new_n1056_, new_n1065_ );
nor g0867 ( new_n1069_, new_n1067_, new_n1068_ );
not g0868 ( new_n1070_, new_n1069_ );
nand g0869 ( new_n1071_, new_n1070_, keyIn_0_54 );
not g0870 ( new_n1072_, new_n1071_ );
nor g0871 ( new_n1073_, new_n1070_, keyIn_0_54 );
nor g0872 ( new_n1074_, new_n1072_, new_n1073_ );
not g0873 ( new_n1075_, new_n1074_ );
nand g0874 ( new_n1076_, new_n1048_, new_n1075_ );
not g0875 ( new_n1077_, new_n1076_ );
nor g0876 ( new_n1078_, new_n1048_, new_n1075_ );
nor g0877 ( new_n1079_, new_n1077_, new_n1078_ );
nand g0878 ( new_n1080_, new_n1079_, new_n1021_ );
not g0879 ( new_n1081_, new_n1043_ );
nor g0880 ( new_n1082_, new_n1042_, new_n1022_ );
nor g0881 ( new_n1083_, new_n1081_, new_n1082_ );
nand g0882 ( new_n1084_, new_n1083_, new_n1074_ );
nand g0883 ( new_n1085_, new_n1084_, new_n1076_ );
nand g0884 ( new_n1086_, new_n1085_, keyIn_0_78 );
nand g0885 ( new_n1087_, new_n1080_, new_n1086_ );
not g0886 ( new_n1088_, keyIn_0_79 );
not g0887 ( new_n1089_, keyIn_0_59 );
nand g0888 ( new_n1090_, new_n816_, new_n951_ );
nand g0889 ( new_n1091_, new_n943_, new_n822_ );
nand g0890 ( new_n1092_, new_n1090_, new_n1091_ );
nand g0891 ( new_n1093_, new_n1092_, new_n1089_ );
nor g0892 ( new_n1094_, new_n1092_, new_n1089_ );
not g0893 ( new_n1095_, new_n1094_ );
nand g0894 ( new_n1096_, new_n1095_, new_n1093_ );
nand g0895 ( new_n1097_, N136, N137 );
nor g0896 ( new_n1098_, new_n1097_, keyIn_0_23 );
nand g0897 ( new_n1099_, new_n1097_, keyIn_0_23 );
not g0898 ( new_n1100_, new_n1099_ );
nor g0899 ( new_n1101_, new_n1100_, new_n1098_ );
not g0900 ( new_n1102_, new_n1101_ );
nand g0901 ( new_n1103_, new_n1096_, new_n1102_ );
not g0902 ( new_n1104_, new_n1093_ );
nor g0903 ( new_n1105_, new_n1104_, new_n1094_ );
nand g0904 ( new_n1106_, new_n1105_, new_n1101_ );
nand g0905 ( new_n1107_, new_n1106_, new_n1103_ );
nand g0906 ( new_n1108_, new_n1107_, keyIn_0_71 );
not g0907 ( new_n1109_, new_n1108_ );
nor g0908 ( new_n1110_, new_n1107_, keyIn_0_71 );
nor g0909 ( new_n1111_, new_n1109_, new_n1110_ );
not g0910 ( new_n1112_, keyIn_0_55 );
not g0911 ( new_n1113_, keyIn_0_38 );
nor g0912 ( new_n1114_, new_n216_, N93 );
nor g0913 ( new_n1115_, new_n247_, N77 );
nor g0914 ( new_n1116_, new_n1114_, new_n1115_ );
not g0915 ( new_n1117_, new_n1116_ );
nand g0916 ( new_n1118_, new_n1117_, new_n1113_ );
not g0917 ( new_n1119_, new_n1118_ );
nor g0918 ( new_n1120_, new_n1117_, new_n1113_ );
nor g0919 ( new_n1121_, new_n1119_, new_n1120_ );
not g0920 ( new_n1122_, keyIn_0_39 );
nor g0921 ( new_n1123_, new_n356_, N125 );
nor g0922 ( new_n1124_, new_n463_, N109 );
nor g0923 ( new_n1125_, new_n1123_, new_n1124_ );
not g0924 ( new_n1126_, new_n1125_ );
nand g0925 ( new_n1127_, new_n1126_, new_n1122_ );
not g0926 ( new_n1128_, new_n1127_ );
nor g0927 ( new_n1129_, new_n1126_, new_n1122_ );
nor g0928 ( new_n1130_, new_n1128_, new_n1129_ );
not g0929 ( new_n1131_, new_n1130_ );
nor g0930 ( new_n1132_, new_n1131_, new_n1121_ );
nand g0931 ( new_n1133_, new_n1131_, new_n1121_ );
not g0932 ( new_n1134_, new_n1133_ );
nor g0933 ( new_n1135_, new_n1134_, new_n1132_ );
not g0934 ( new_n1136_, new_n1135_ );
nand g0935 ( new_n1137_, new_n1136_, new_n1112_ );
not g0936 ( new_n1138_, new_n1137_ );
nor g0937 ( new_n1139_, new_n1136_, new_n1112_ );
nor g0938 ( new_n1140_, new_n1138_, new_n1139_ );
nor g0939 ( new_n1141_, new_n1111_, new_n1140_ );
not g0940 ( new_n1142_, keyIn_0_71 );
nor g0941 ( new_n1143_, new_n1105_, new_n1101_ );
nor g0942 ( new_n1144_, new_n1096_, new_n1102_ );
nor g0943 ( new_n1145_, new_n1143_, new_n1144_ );
nand g0944 ( new_n1146_, new_n1145_, new_n1142_ );
nand g0945 ( new_n1147_, new_n1146_, new_n1108_ );
not g0946 ( new_n1148_, new_n1140_ );
nor g0947 ( new_n1149_, new_n1147_, new_n1148_ );
nor g0948 ( new_n1150_, new_n1141_, new_n1149_ );
nand g0949 ( new_n1151_, new_n1150_, new_n1088_ );
nand g0950 ( new_n1152_, new_n1147_, new_n1148_ );
nand g0951 ( new_n1153_, new_n1111_, new_n1140_ );
nand g0952 ( new_n1154_, new_n1153_, new_n1152_ );
nand g0953 ( new_n1155_, new_n1154_, keyIn_0_79 );
nand g0954 ( new_n1156_, new_n1151_, new_n1155_ );
nor g0955 ( new_n1157_, new_n1156_, new_n1087_ );
not g0956 ( new_n1158_, new_n1157_ );
nor g0957 ( new_n1159_, new_n1020_, new_n1158_ );
nand g0958 ( new_n1160_, new_n760_, new_n1159_ );
nor g0959 ( new_n1161_, new_n1160_, new_n343_ );
nand g0960 ( new_n1162_, new_n1160_, new_n343_ );
not g0961 ( new_n1163_, new_n1162_ );
nor g0962 ( new_n1164_, new_n1163_, new_n1161_ );
not g0963 ( new_n1165_, new_n1164_ );
nor g0964 ( new_n1166_, new_n1165_, new_n342_ );
not g0965 ( new_n1167_, new_n1166_ );
nand g0966 ( new_n1168_, new_n1167_, N1 );
nand g0967 ( new_n1169_, new_n1166_, new_n299_ );
nand g0968 ( N724, new_n1168_, new_n1169_ );
nor g0969 ( new_n1171_, new_n1165_, new_n644_ );
not g0970 ( new_n1172_, new_n1171_ );
nand g0971 ( new_n1173_, new_n1172_, N5 );
nand g0972 ( new_n1174_, new_n1171_, new_n596_ );
nand g0973 ( N725, new_n1173_, new_n1174_ );
nor g0974 ( new_n1176_, new_n1165_, new_n451_ );
not g0975 ( new_n1177_, new_n1176_ );
nand g0976 ( new_n1178_, new_n1177_, N9 );
nand g0977 ( new_n1179_, new_n1176_, new_n408_ );
nand g0978 ( N726, new_n1178_, new_n1179_ );
nor g0979 ( new_n1181_, new_n1165_, new_n678_ );
not g0980 ( new_n1182_, new_n1181_ );
nand g0981 ( new_n1183_, new_n1182_, N13 );
nand g0982 ( new_n1184_, new_n1181_, new_n518_ );
nand g0983 ( N727, new_n1183_, new_n1184_ );
nand g0984 ( new_n1186_, new_n1156_, new_n1087_ );
nor g0985 ( new_n1187_, new_n1020_, new_n1186_ );
nand g0986 ( new_n1188_, new_n760_, new_n1187_ );
nor g0987 ( new_n1189_, new_n1188_, keyIn_0_115 );
nand g0988 ( new_n1190_, new_n1188_, keyIn_0_115 );
not g0989 ( new_n1191_, new_n1190_ );
nor g0990 ( new_n1192_, new_n1191_, new_n1189_ );
not g0991 ( new_n1193_, new_n1192_ );
nor g0992 ( new_n1194_, new_n1193_, new_n342_ );
not g0993 ( new_n1195_, new_n1194_ );
nand g0994 ( new_n1196_, new_n1195_, N17 );
nand g0995 ( new_n1197_, new_n1194_, new_n301_ );
nand g0996 ( N728, new_n1196_, new_n1197_ );
nor g0997 ( new_n1199_, new_n1193_, new_n644_ );
not g0998 ( new_n1200_, new_n1199_ );
nand g0999 ( new_n1201_, new_n1200_, N21 );
nand g1000 ( new_n1202_, new_n1199_, new_n598_ );
nand g1001 ( N729, new_n1201_, new_n1202_ );
nor g1002 ( new_n1204_, new_n1193_, new_n451_ );
not g1003 ( new_n1205_, new_n1204_ );
nand g1004 ( new_n1206_, new_n1205_, N25 );
nand g1005 ( new_n1207_, new_n1204_, new_n410_ );
nand g1006 ( N730, new_n1206_, new_n1207_ );
nor g1007 ( new_n1209_, new_n1193_, new_n678_ );
not g1008 ( new_n1210_, new_n1209_ );
nand g1009 ( new_n1211_, new_n1210_, N29 );
nand g1010 ( new_n1212_, new_n1209_, new_n520_ );
nand g1011 ( N731, new_n1211_, new_n1212_ );
not g1012 ( new_n1214_, keyIn_0_116 );
nand g1013 ( new_n1215_, new_n886_, new_n880_ );
nand g1014 ( new_n1216_, new_n878_, keyIn_0_76 );
nand g1015 ( new_n1217_, new_n1216_, new_n1215_ );
nor g1016 ( new_n1218_, new_n1016_, keyIn_0_77 );
not g1017 ( new_n1219_, new_n1017_ );
nor g1018 ( new_n1220_, new_n1219_, new_n1218_ );
nor g1019 ( new_n1221_, new_n1220_, new_n1217_ );
not g1020 ( new_n1222_, new_n1221_ );
nor g1021 ( new_n1223_, new_n1222_, new_n1158_ );
nand g1022 ( new_n1224_, new_n760_, new_n1223_ );
nor g1023 ( new_n1225_, new_n1224_, new_n1214_ );
nand g1024 ( new_n1226_, new_n1224_, new_n1214_ );
not g1025 ( new_n1227_, new_n1226_ );
nor g1026 ( new_n1228_, new_n1227_, new_n1225_ );
nor g1027 ( new_n1229_, new_n1228_, new_n342_ );
not g1028 ( new_n1230_, new_n1229_ );
nand g1029 ( new_n1231_, new_n1230_, N33 );
nand g1030 ( new_n1232_, new_n1229_, new_n309_ );
nand g1031 ( N732, new_n1231_, new_n1232_ );
nor g1032 ( new_n1234_, new_n1228_, new_n644_ );
not g1033 ( new_n1235_, new_n1234_ );
nand g1034 ( new_n1236_, new_n1235_, N37 );
nand g1035 ( new_n1237_, new_n1234_, new_n607_ );
nand g1036 ( N733, new_n1236_, new_n1237_ );
nor g1037 ( new_n1239_, new_n1228_, new_n451_ );
not g1038 ( new_n1240_, new_n1239_ );
nand g1039 ( new_n1241_, new_n1240_, N41 );
nand g1040 ( new_n1242_, new_n1239_, new_n418_ );
nand g1041 ( N734, new_n1241_, new_n1242_ );
nor g1042 ( new_n1244_, new_n1228_, new_n678_ );
not g1043 ( new_n1245_, new_n1244_ );
nand g1044 ( new_n1246_, new_n1245_, N45 );
nand g1045 ( new_n1247_, new_n1244_, new_n530_ );
nand g1046 ( N735, new_n1246_, new_n1247_ );
nand g1047 ( new_n1249_, new_n758_, keyIn_0_112 );
nand g1048 ( new_n1250_, new_n742_, new_n344_ );
nand g1049 ( new_n1251_, new_n1249_, new_n1250_ );
nor g1050 ( new_n1252_, new_n1222_, new_n1186_ );
not g1051 ( new_n1253_, new_n1252_ );
nor g1052 ( new_n1254_, new_n1251_, new_n1253_ );
nor g1053 ( new_n1255_, new_n1254_, keyIn_0_117 );
not g1054 ( new_n1256_, keyIn_0_117 );
nand g1055 ( new_n1257_, new_n760_, new_n1252_ );
nor g1056 ( new_n1258_, new_n1257_, new_n1256_ );
nor g1057 ( new_n1259_, new_n1258_, new_n1255_ );
nor g1058 ( new_n1260_, new_n1259_, new_n342_ );
not g1059 ( new_n1261_, new_n1260_ );
nand g1060 ( new_n1262_, new_n1261_, N49 );
nand g1061 ( new_n1263_, new_n1260_, new_n311_ );
nand g1062 ( N736, new_n1262_, new_n1263_ );
nor g1063 ( new_n1265_, new_n1259_, new_n644_ );
not g1064 ( new_n1266_, new_n1265_ );
nand g1065 ( new_n1267_, new_n1266_, N53 );
nand g1066 ( new_n1268_, new_n1265_, new_n609_ );
nand g1067 ( N737, new_n1267_, new_n1268_ );
nor g1068 ( new_n1270_, new_n1259_, new_n451_ );
not g1069 ( new_n1271_, new_n1270_ );
nand g1070 ( new_n1272_, new_n1271_, N57 );
nand g1071 ( new_n1273_, new_n1270_, new_n420_ );
nand g1072 ( N738, new_n1272_, new_n1273_ );
nand g1073 ( new_n1275_, new_n1257_, new_n1256_ );
nand g1074 ( new_n1276_, new_n1254_, keyIn_0_117 );
nand g1075 ( new_n1277_, new_n1275_, new_n1276_ );
nand g1076 ( new_n1278_, new_n1277_, new_n562_ );
nand g1077 ( new_n1279_, new_n1278_, keyIn_0_122 );
not g1078 ( new_n1280_, keyIn_0_122 );
not g1079 ( new_n1281_, new_n1278_ );
nand g1080 ( new_n1282_, new_n1281_, new_n1280_ );
nand g1081 ( new_n1283_, new_n1282_, new_n1279_ );
nand g1082 ( new_n1284_, new_n1283_, new_n532_ );
not g1083 ( new_n1285_, new_n1279_ );
nor g1084 ( new_n1286_, new_n1278_, keyIn_0_122 );
nor g1085 ( new_n1287_, new_n1285_, new_n1286_ );
nand g1086 ( new_n1288_, new_n1287_, N61 );
nand g1087 ( N739, new_n1288_, new_n1284_ );
not g1088 ( new_n1290_, keyIn_0_118 );
not g1089 ( new_n1291_, keyIn_0_113 );
not g1090 ( new_n1292_, keyIn_0_108 );
nor g1091 ( new_n1293_, new_n888_, keyIn_0_92 );
not g1092 ( new_n1294_, new_n1293_ );
nor g1093 ( new_n1295_, new_n1154_, keyIn_0_79 );
not g1094 ( new_n1296_, new_n1155_ );
nor g1095 ( new_n1297_, new_n1296_, new_n1295_ );
not g1096 ( new_n1298_, keyIn_0_92 );
nor g1097 ( new_n1299_, new_n1217_, new_n1298_ );
nor g1098 ( new_n1300_, new_n1299_, new_n1297_ );
nand g1099 ( new_n1301_, new_n1300_, new_n1294_ );
not g1100 ( new_n1302_, new_n1301_ );
not g1101 ( new_n1303_, keyIn_0_93 );
nand g1102 ( new_n1304_, new_n1220_, new_n1303_ );
nand g1103 ( new_n1305_, new_n1018_, keyIn_0_93 );
nand g1104 ( new_n1306_, new_n1304_, new_n1305_ );
not g1105 ( new_n1307_, keyIn_0_94 );
nor g1106 ( new_n1308_, new_n1085_, keyIn_0_78 );
nor g1107 ( new_n1309_, new_n1079_, new_n1021_ );
nor g1108 ( new_n1310_, new_n1309_, new_n1308_ );
nand g1109 ( new_n1311_, new_n1310_, new_n1307_ );
nand g1110 ( new_n1312_, new_n1087_, keyIn_0_94 );
nand g1111 ( new_n1313_, new_n1311_, new_n1312_ );
nand g1112 ( new_n1314_, new_n1313_, new_n1306_ );
not g1113 ( new_n1315_, new_n1314_ );
nand g1114 ( new_n1316_, new_n1315_, new_n1302_ );
nand g1115 ( new_n1317_, new_n1316_, new_n1292_ );
nor g1116 ( new_n1318_, new_n1314_, new_n1301_ );
nand g1117 ( new_n1319_, new_n1318_, keyIn_0_108 );
nand g1118 ( new_n1320_, new_n1317_, new_n1319_ );
not g1119 ( new_n1321_, keyIn_0_109 );
nor g1120 ( new_n1322_, new_n1156_, keyIn_0_97 );
nand g1121 ( new_n1323_, new_n1156_, keyIn_0_97 );
nand g1122 ( new_n1324_, new_n1323_, new_n1310_ );
nor g1123 ( new_n1325_, new_n1324_, new_n1322_ );
nand g1124 ( new_n1326_, new_n1220_, keyIn_0_96 );
not g1125 ( new_n1327_, keyIn_0_96 );
nand g1126 ( new_n1328_, new_n1018_, new_n1327_ );
nand g1127 ( new_n1329_, new_n1326_, new_n1328_ );
nand g1128 ( new_n1330_, new_n888_, keyIn_0_95 );
not g1129 ( new_n1331_, keyIn_0_95 );
nand g1130 ( new_n1332_, new_n1217_, new_n1331_ );
nand g1131 ( new_n1333_, new_n1330_, new_n1332_ );
nand g1132 ( new_n1334_, new_n1329_, new_n1333_ );
not g1133 ( new_n1335_, new_n1334_ );
nand g1134 ( new_n1336_, new_n1335_, new_n1325_ );
nand g1135 ( new_n1337_, new_n1336_, new_n1321_ );
not g1136 ( new_n1338_, new_n1322_ );
not g1137 ( new_n1339_, new_n1324_ );
nand g1138 ( new_n1340_, new_n1339_, new_n1338_ );
nor g1139 ( new_n1341_, new_n1340_, new_n1334_ );
nand g1140 ( new_n1342_, new_n1341_, keyIn_0_109 );
nand g1141 ( new_n1343_, new_n1337_, new_n1342_ );
nor g1142 ( new_n1344_, new_n1320_, new_n1343_ );
not g1143 ( new_n1345_, keyIn_0_110 );
not g1144 ( new_n1346_, keyIn_0_100 );
nor g1145 ( new_n1347_, new_n1297_, new_n1346_ );
nor g1146 ( new_n1348_, new_n1087_, keyIn_0_99 );
not g1147 ( new_n1349_, new_n1348_ );
nand g1148 ( new_n1350_, new_n1297_, new_n1346_ );
nand g1149 ( new_n1351_, new_n1349_, new_n1350_ );
nor g1150 ( new_n1352_, new_n1351_, new_n1347_ );
not g1151 ( new_n1353_, keyIn_0_98 );
nor g1152 ( new_n1354_, new_n1217_, new_n1353_ );
nand g1153 ( new_n1355_, new_n1217_, new_n1353_ );
not g1154 ( new_n1356_, new_n1355_ );
nor g1155 ( new_n1357_, new_n1356_, new_n1354_ );
nand g1156 ( new_n1358_, new_n1087_, keyIn_0_99 );
nand g1157 ( new_n1359_, new_n1358_, new_n1018_ );
nor g1158 ( new_n1360_, new_n1357_, new_n1359_ );
nand g1159 ( new_n1361_, new_n1352_, new_n1360_ );
nand g1160 ( new_n1362_, new_n1361_, new_n1345_ );
not g1161 ( new_n1363_, new_n1347_ );
nor g1162 ( new_n1364_, new_n1156_, keyIn_0_100 );
nor g1163 ( new_n1365_, new_n1364_, new_n1348_ );
nand g1164 ( new_n1366_, new_n1365_, new_n1363_ );
nand g1165 ( new_n1367_, new_n888_, keyIn_0_98 );
nand g1166 ( new_n1368_, new_n1367_, new_n1355_ );
not g1167 ( new_n1369_, new_n1359_ );
nand g1168 ( new_n1370_, new_n1369_, new_n1368_ );
nor g1169 ( new_n1371_, new_n1370_, new_n1366_ );
nand g1170 ( new_n1372_, new_n1371_, keyIn_0_110 );
nand g1171 ( new_n1373_, new_n1362_, new_n1372_ );
nand g1172 ( new_n1374_, new_n1156_, keyIn_0_103 );
not g1173 ( new_n1375_, new_n1374_ );
not g1174 ( new_n1376_, keyIn_0_103 );
nand g1175 ( new_n1377_, new_n1297_, new_n1376_ );
not g1176 ( new_n1378_, keyIn_0_101 );
nand g1177 ( new_n1379_, new_n1220_, new_n1378_ );
nand g1178 ( new_n1380_, new_n1377_, new_n1379_ );
nor g1179 ( new_n1381_, new_n1380_, new_n1375_ );
not g1180 ( new_n1382_, keyIn_0_102 );
nor g1181 ( new_n1383_, new_n1087_, new_n1382_ );
nor g1182 ( new_n1384_, new_n1310_, keyIn_0_102 );
nor g1183 ( new_n1385_, new_n1384_, new_n1383_ );
nand g1184 ( new_n1386_, new_n1018_, keyIn_0_101 );
nand g1185 ( new_n1387_, new_n1386_, new_n1217_ );
nor g1186 ( new_n1388_, new_n1385_, new_n1387_ );
nand g1187 ( new_n1389_, new_n1388_, new_n1381_ );
nand g1188 ( new_n1390_, new_n1389_, keyIn_0_111 );
not g1189 ( new_n1391_, keyIn_0_111 );
nor g1190 ( new_n1392_, new_n1156_, keyIn_0_103 );
nor g1191 ( new_n1393_, new_n1018_, keyIn_0_101 );
nor g1192 ( new_n1394_, new_n1392_, new_n1393_ );
nand g1193 ( new_n1395_, new_n1394_, new_n1374_ );
nand g1194 ( new_n1396_, new_n1310_, keyIn_0_102 );
nand g1195 ( new_n1397_, new_n1087_, new_n1382_ );
nand g1196 ( new_n1398_, new_n1396_, new_n1397_ );
not g1197 ( new_n1399_, new_n1387_ );
nand g1198 ( new_n1400_, new_n1399_, new_n1398_ );
nor g1199 ( new_n1401_, new_n1400_, new_n1395_ );
nand g1200 ( new_n1402_, new_n1401_, new_n1391_ );
nand g1201 ( new_n1403_, new_n1390_, new_n1402_ );
nor g1202 ( new_n1404_, new_n1373_, new_n1403_ );
nand g1203 ( new_n1405_, new_n1344_, new_n1404_ );
nand g1204 ( new_n1406_, new_n1405_, new_n1291_ );
nor g1205 ( new_n1407_, new_n1318_, keyIn_0_108 );
not g1206 ( new_n1408_, new_n1319_ );
nor g1207 ( new_n1409_, new_n1408_, new_n1407_ );
nor g1208 ( new_n1410_, new_n1341_, keyIn_0_109 );
nor g1209 ( new_n1411_, new_n1336_, new_n1321_ );
nor g1210 ( new_n1412_, new_n1411_, new_n1410_ );
nand g1211 ( new_n1413_, new_n1409_, new_n1412_ );
nor g1212 ( new_n1414_, new_n1371_, keyIn_0_110 );
nor g1213 ( new_n1415_, new_n1361_, new_n1345_ );
nor g1214 ( new_n1416_, new_n1415_, new_n1414_ );
nor g1215 ( new_n1417_, new_n1401_, new_n1391_ );
nor g1216 ( new_n1418_, new_n1389_, keyIn_0_111 );
nor g1217 ( new_n1419_, new_n1418_, new_n1417_ );
nand g1218 ( new_n1420_, new_n1416_, new_n1419_ );
nor g1219 ( new_n1421_, new_n1413_, new_n1420_ );
nand g1220 ( new_n1422_, new_n1421_, keyIn_0_113 );
nand g1221 ( new_n1423_, new_n1422_, new_n1406_ );
nor g1222 ( new_n1424_, new_n637_, new_n342_ );
not g1223 ( new_n1425_, new_n1424_ );
nor g1224 ( new_n1426_, new_n562_, new_n451_ );
not g1225 ( new_n1427_, new_n1426_ );
nor g1226 ( new_n1428_, new_n1425_, new_n1427_ );
not g1227 ( new_n1429_, new_n1428_ );
nor g1228 ( new_n1430_, new_n1423_, new_n1429_ );
nand g1229 ( new_n1431_, new_n1430_, new_n1290_ );
not g1230 ( new_n1432_, new_n1406_ );
nor g1231 ( new_n1433_, new_n1405_, new_n1291_ );
nor g1232 ( new_n1434_, new_n1432_, new_n1433_ );
nand g1233 ( new_n1435_, new_n1434_, new_n1428_ );
nand g1234 ( new_n1436_, new_n1435_, keyIn_0_118 );
nand g1235 ( new_n1437_, new_n1436_, new_n1431_ );
nand g1236 ( new_n1438_, new_n1437_, new_n1217_ );
nand g1237 ( new_n1439_, new_n1438_, keyIn_0_123 );
not g1238 ( new_n1440_, keyIn_0_123 );
not g1239 ( new_n1441_, new_n1438_ );
nand g1240 ( new_n1442_, new_n1441_, new_n1440_ );
nand g1241 ( new_n1443_, new_n1442_, new_n1439_ );
nand g1242 ( new_n1444_, new_n1443_, N65 );
not g1243 ( new_n1445_, new_n1439_ );
nor g1244 ( new_n1446_, new_n1438_, keyIn_0_123 );
nor g1245 ( new_n1447_, new_n1445_, new_n1446_ );
nand g1246 ( new_n1448_, new_n1447_, new_n208_ );
nand g1247 ( N740, new_n1448_, new_n1444_ );
not g1248 ( new_n1450_, keyIn_0_124 );
nand g1249 ( new_n1451_, new_n1437_, new_n1018_ );
nand g1250 ( new_n1452_, new_n1451_, new_n1450_ );
not g1251 ( new_n1453_, new_n1451_ );
nand g1252 ( new_n1454_, new_n1453_, keyIn_0_124 );
nand g1253 ( new_n1455_, new_n1454_, new_n1452_ );
nand g1254 ( new_n1456_, new_n1455_, new_n206_ );
not g1255 ( new_n1457_, new_n1452_ );
nor g1256 ( new_n1458_, new_n1451_, new_n1450_ );
nor g1257 ( new_n1459_, new_n1457_, new_n1458_ );
nand g1258 ( new_n1460_, new_n1459_, N69 );
nand g1259 ( N741, new_n1460_, new_n1456_ );
not g1260 ( new_n1462_, keyIn_0_125 );
nand g1261 ( new_n1463_, new_n1437_, new_n1310_ );
nand g1262 ( new_n1464_, new_n1463_, new_n1462_ );
not g1263 ( new_n1465_, new_n1463_ );
nand g1264 ( new_n1466_, new_n1465_, keyIn_0_125 );
nand g1265 ( new_n1467_, new_n1466_, new_n1464_ );
nand g1266 ( new_n1468_, new_n1467_, N73 );
not g1267 ( new_n1469_, new_n1464_ );
nor g1268 ( new_n1470_, new_n1463_, new_n1462_ );
nor g1269 ( new_n1471_, new_n1469_, new_n1470_ );
nand g1270 ( new_n1472_, new_n1471_, new_n218_ );
nand g1271 ( N742, new_n1472_, new_n1468_ );
not g1272 ( new_n1474_, keyIn_0_126 );
nand g1273 ( new_n1475_, new_n1437_, new_n1156_ );
nand g1274 ( new_n1476_, new_n1475_, new_n1474_ );
not g1275 ( new_n1477_, new_n1475_ );
nand g1276 ( new_n1478_, new_n1477_, keyIn_0_126 );
nand g1277 ( new_n1479_, new_n1478_, new_n1476_ );
nand g1278 ( new_n1480_, new_n1479_, new_n216_ );
not g1279 ( new_n1481_, new_n1476_ );
nor g1280 ( new_n1482_, new_n1475_, new_n1474_ );
nor g1281 ( new_n1483_, new_n1481_, new_n1482_ );
nand g1282 ( new_n1484_, new_n1483_, N77 );
nand g1283 ( N743, new_n1484_, new_n1480_ );
not g1284 ( new_n1486_, keyIn_0_119 );
nor g1285 ( new_n1487_, new_n666_, new_n678_ );
not g1286 ( new_n1488_, new_n1487_ );
nor g1287 ( new_n1489_, new_n1488_, new_n1425_ );
not g1288 ( new_n1490_, new_n1489_ );
nor g1289 ( new_n1491_, new_n1423_, new_n1490_ );
nand g1290 ( new_n1492_, new_n1491_, new_n1486_ );
nand g1291 ( new_n1493_, new_n1434_, new_n1489_ );
nand g1292 ( new_n1494_, new_n1493_, keyIn_0_119 );
nand g1293 ( new_n1495_, new_n1494_, new_n1492_ );
nand g1294 ( new_n1496_, new_n1495_, new_n1217_ );
nand g1295 ( new_n1497_, new_n1496_, keyIn_0_127 );
not g1296 ( new_n1498_, keyIn_0_127 );
not g1297 ( new_n1499_, new_n1496_ );
nand g1298 ( new_n1500_, new_n1499_, new_n1498_ );
nand g1299 ( new_n1501_, new_n1500_, new_n1497_ );
nand g1300 ( new_n1502_, new_n1501_, N81 );
not g1301 ( new_n1503_, new_n1497_ );
nor g1302 ( new_n1504_, new_n1496_, keyIn_0_127 );
nor g1303 ( new_n1505_, new_n1503_, new_n1504_ );
nand g1304 ( new_n1506_, new_n1505_, new_n240_ );
nand g1305 ( N744, new_n1506_, new_n1502_ );
nand g1306 ( new_n1508_, new_n1495_, new_n1018_ );
nand g1307 ( new_n1509_, new_n1508_, N85 );
not g1308 ( new_n1510_, new_n1508_ );
nand g1309 ( new_n1511_, new_n1510_, new_n238_ );
nand g1310 ( N745, new_n1511_, new_n1509_ );
nand g1311 ( new_n1513_, new_n1495_, new_n1310_ );
nand g1312 ( new_n1514_, new_n1513_, N89 );
not g1313 ( new_n1515_, new_n1513_ );
nand g1314 ( new_n1516_, new_n1515_, new_n249_ );
nand g1315 ( N746, new_n1516_, new_n1514_ );
nand g1316 ( new_n1518_, new_n1495_, new_n1156_ );
nand g1317 ( new_n1519_, new_n1518_, N93 );
not g1318 ( new_n1520_, new_n1518_ );
nand g1319 ( new_n1521_, new_n1520_, new_n247_ );
nand g1320 ( N747, new_n1521_, new_n1519_ );
not g1321 ( new_n1523_, keyIn_0_120 );
nor g1322 ( new_n1524_, new_n650_, new_n644_ );
not g1323 ( new_n1525_, new_n1524_ );
nor g1324 ( new_n1526_, new_n1525_, new_n1427_ );
nand g1325 ( new_n1527_, new_n1434_, new_n1526_ );
not g1326 ( new_n1528_, new_n1527_ );
nand g1327 ( new_n1529_, new_n1528_, new_n1523_ );
nand g1328 ( new_n1530_, new_n1527_, keyIn_0_120 );
nand g1329 ( new_n1531_, new_n1529_, new_n1530_ );
nor g1330 ( new_n1532_, new_n1531_, new_n888_ );
not g1331 ( new_n1533_, new_n1532_ );
nand g1332 ( new_n1534_, new_n1533_, N97 );
nand g1333 ( new_n1535_, new_n1532_, new_n348_ );
nand g1334 ( N748, new_n1534_, new_n1535_ );
nor g1335 ( new_n1537_, new_n1531_, new_n1220_ );
not g1336 ( new_n1538_, new_n1537_ );
nand g1337 ( new_n1539_, new_n1538_, N101 );
nand g1338 ( new_n1540_, new_n1537_, new_n346_ );
nand g1339 ( N749, new_n1539_, new_n1540_ );
nor g1340 ( new_n1542_, new_n1531_, new_n1087_ );
not g1341 ( new_n1543_, new_n1542_ );
nand g1342 ( new_n1544_, new_n1543_, N105 );
nand g1343 ( new_n1545_, new_n1542_, new_n358_ );
nand g1344 ( N750, new_n1544_, new_n1545_ );
nor g1345 ( new_n1547_, new_n1531_, new_n1297_ );
not g1346 ( new_n1548_, new_n1547_ );
nand g1347 ( new_n1549_, new_n1548_, N109 );
nand g1348 ( new_n1550_, new_n1547_, new_n356_ );
nand g1349 ( N751, new_n1549_, new_n1550_ );
nor g1350 ( new_n1552_, new_n1488_, new_n1525_ );
nand g1351 ( new_n1553_, new_n1434_, new_n1552_ );
not g1352 ( new_n1554_, new_n1553_ );
nand g1353 ( new_n1555_, new_n1554_, keyIn_0_121 );
not g1354 ( new_n1556_, keyIn_0_121 );
nand g1355 ( new_n1557_, new_n1553_, new_n1556_ );
nand g1356 ( new_n1558_, new_n1555_, new_n1557_ );
nor g1357 ( new_n1559_, new_n1558_, new_n888_ );
not g1358 ( new_n1560_, new_n1559_ );
nand g1359 ( new_n1561_, new_n1560_, N113 );
nand g1360 ( new_n1562_, new_n1559_, new_n456_ );
nand g1361 ( N752, new_n1561_, new_n1562_ );
nor g1362 ( new_n1564_, new_n1558_, new_n1220_ );
not g1363 ( new_n1565_, new_n1564_ );
nand g1364 ( new_n1566_, new_n1565_, N117 );
nand g1365 ( new_n1567_, new_n1564_, new_n454_ );
nand g1366 ( N753, new_n1566_, new_n1567_ );
nor g1367 ( new_n1569_, new_n1558_, new_n1087_ );
not g1368 ( new_n1570_, new_n1569_ );
nand g1369 ( new_n1571_, new_n1570_, N121 );
nand g1370 ( new_n1572_, new_n1569_, new_n465_ );
nand g1371 ( N754, new_n1571_, new_n1572_ );
nor g1372 ( new_n1574_, new_n1558_, new_n1297_ );
not g1373 ( new_n1575_, new_n1574_ );
nand g1374 ( new_n1576_, new_n1575_, N125 );
nand g1375 ( new_n1577_, new_n1574_, new_n463_ );
nand g1376 ( N755, new_n1576_, new_n1577_ );
endmodule