module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n620_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n636_, new_n456_, new_n170_, new_n246_, new_n266_, new_n367_, new_n542_, new_n548_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n117_, new_n630_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n656_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n621_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n559_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n628_, new_n166_, new_n409_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n113_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n633_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n604_, new_n227_, new_n416_, new_n222_, new_n571_, new_n400_, new_n328_, new_n460_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n562_, new_n525_, new_n578_, new_n126_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n625_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n588_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n112_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n115_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n651_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n584_, new_n278_, new_n304_, new_n523_, new_n638_, new_n550_, new_n217_, new_n269_, new_n512_, new_n129_, new_n644_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n574_, new_n319_, new_n640_, new_n338_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n330_, new_n375_, new_n294_, new_n627_, new_n195_, new_n567_, new_n576_, new_n357_, new_n320_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n120_, new_n521_, new_n406_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n405_;

not g000 ( new_n108_, N30 );
or g001 ( new_n109_, new_n108_, N24 );
and g002 ( new_n110_, new_n109_, keyIn_0_8 );
not g003 ( new_n111_, keyIn_0_8 );
not g004 ( new_n112_, N24 );
and g005 ( new_n113_, new_n111_, new_n112_, N30 );
or g006 ( new_n114_, new_n110_, new_n113_ );
not g007 ( new_n115_, N69 );
or g008 ( new_n116_, new_n115_, N63 );
and g009 ( new_n117_, new_n116_, keyIn_0_9 );
not g010 ( new_n118_, keyIn_0_9 );
not g011 ( new_n119_, N63 );
and g012 ( new_n120_, new_n118_, new_n119_, N69 );
or g013 ( new_n121_, new_n117_, new_n120_ );
not g014 ( new_n122_, keyIn_0_7 );
not g015 ( new_n123_, N17 );
or g016 ( new_n124_, new_n123_, N11 );
and g017 ( new_n125_, new_n124_, new_n122_ );
not g018 ( new_n126_, N11 );
and g019 ( new_n127_, new_n126_, keyIn_0_7, N17 );
or g020 ( new_n128_, new_n125_, new_n127_ );
and g021 ( new_n129_, new_n114_, new_n121_, new_n128_ );
and g022 ( new_n130_, keyIn_0_5, N89 );
not g023 ( new_n131_, new_n130_ );
or g024 ( new_n132_, keyIn_0_5, N89 );
and g025 ( new_n133_, new_n131_, N95, new_n132_ );
not g026 ( new_n134_, new_n133_ );
not g027 ( new_n135_, N4 );
or g028 ( new_n136_, new_n135_, N1 );
not g029 ( new_n137_, N82 );
or g030 ( new_n138_, new_n137_, N76 );
not g031 ( new_n139_, N50 );
and g032 ( new_n140_, new_n139_, N56 );
not g033 ( new_n141_, new_n140_ );
and g034 ( new_n142_, new_n141_, new_n136_, new_n138_ );
not g035 ( new_n143_, N43 );
not g036 ( new_n144_, keyIn_0_2 );
and g037 ( new_n145_, new_n144_, N37 );
not g038 ( new_n146_, N37 );
and g039 ( new_n147_, new_n146_, keyIn_0_2 );
or g040 ( new_n148_, new_n145_, new_n147_, new_n143_ );
not g041 ( new_n149_, N108 );
or g042 ( new_n150_, new_n149_, N102 );
and g043 ( new_n151_, new_n150_, keyIn_0_10 );
not g044 ( new_n152_, keyIn_0_10 );
not g045 ( new_n153_, N102 );
and g046 ( new_n154_, new_n152_, new_n153_, N108 );
or g047 ( new_n155_, new_n151_, new_n154_ );
and g048 ( new_n156_, new_n155_, new_n134_, new_n142_, new_n148_ );
and g049 ( new_n157_, new_n156_, new_n129_ );
not g050 ( new_n158_, new_n157_ );
and g051 ( new_n159_, new_n158_, keyIn_0_20 );
not g052 ( new_n160_, keyIn_0_20 );
and g053 ( new_n161_, new_n157_, new_n160_ );
or g054 ( N223, new_n159_, new_n161_ );
not g055 ( new_n163_, keyIn_0_32 );
not g056 ( new_n164_, keyIn_0_21 );
not g057 ( new_n165_, keyIn_0_18 );
not g058 ( new_n166_, new_n128_ );
and g059 ( new_n167_, new_n166_, new_n165_ );
or g060 ( new_n168_, new_n157_, keyIn_0_18 );
and g061 ( new_n169_, new_n156_, new_n129_, keyIn_0_18 );
not g062 ( new_n170_, new_n169_ );
and g063 ( new_n171_, new_n168_, new_n128_, new_n170_ );
or g064 ( new_n172_, new_n171_, new_n167_ );
and g065 ( new_n173_, new_n172_, new_n164_ );
not g066 ( new_n174_, new_n167_ );
not g067 ( new_n175_, new_n171_ );
and g068 ( new_n176_, new_n175_, keyIn_0_21, new_n174_ );
or g069 ( new_n177_, new_n173_, new_n176_, new_n123_, N21 );
and g070 ( new_n178_, new_n177_, keyIn_0_29 );
not g071 ( new_n179_, keyIn_0_29 );
not g072 ( new_n180_, new_n173_ );
not g073 ( new_n181_, N21 );
not g074 ( new_n182_, new_n176_ );
and g075 ( new_n183_, new_n182_, new_n181_ );
and g076 ( new_n184_, new_n183_, new_n179_, N17, new_n180_ );
or g077 ( new_n185_, new_n178_, new_n184_ );
not g078 ( new_n186_, N86 );
not g079 ( new_n187_, new_n138_ );
and g080 ( new_n188_, new_n168_, new_n170_ );
and g081 ( new_n189_, new_n188_, new_n187_ );
not g082 ( new_n190_, new_n189_ );
or g083 ( new_n191_, new_n188_, new_n187_ );
and g084 ( new_n192_, new_n190_, N82, new_n186_, new_n191_ );
not g085 ( new_n193_, new_n192_ );
not g086 ( new_n194_, N73 );
not g087 ( new_n195_, new_n121_ );
and g088 ( new_n196_, new_n188_, new_n195_ );
not g089 ( new_n197_, new_n196_ );
or g090 ( new_n198_, new_n188_, new_n195_ );
and g091 ( new_n199_, keyIn_0_4, N69 );
not g092 ( new_n200_, new_n199_ );
or g093 ( new_n201_, keyIn_0_4, N69 );
and g094 ( new_n202_, new_n200_, new_n201_ );
not g095 ( new_n203_, new_n202_ );
and g096 ( new_n204_, new_n197_, new_n194_, new_n198_, new_n203_ );
not g097 ( new_n205_, new_n204_ );
and g098 ( new_n206_, new_n193_, new_n205_ );
or g099 ( new_n207_, new_n114_, new_n165_ );
not g100 ( new_n208_, new_n114_ );
or g101 ( new_n209_, new_n188_, new_n208_ );
and g102 ( new_n210_, new_n209_, new_n207_ );
not g103 ( new_n211_, N34 );
and g104 ( new_n212_, new_n108_, keyIn_0_1 );
not g105 ( new_n213_, new_n212_ );
or g106 ( new_n214_, new_n108_, keyIn_0_1 );
and g107 ( new_n215_, new_n213_, new_n214_ );
and g108 ( new_n216_, new_n215_, new_n211_ );
and g109 ( new_n217_, new_n210_, new_n216_ );
not g110 ( new_n218_, new_n217_ );
not g111 ( new_n219_, N99 );
and g112 ( new_n220_, new_n188_, new_n133_ );
not g113 ( new_n221_, new_n220_ );
or g114 ( new_n222_, new_n188_, new_n133_ );
and g115 ( new_n223_, new_n221_, new_n222_ );
and g116 ( new_n224_, new_n223_, N95, new_n219_ );
not g117 ( new_n225_, new_n224_ );
and g118 ( new_n226_, new_n188_, new_n140_ );
not g119 ( new_n227_, new_n226_ );
or g120 ( new_n228_, new_n188_, new_n140_ );
not g121 ( new_n229_, N60 );
and g122 ( new_n230_, new_n229_, N56 );
or g123 ( new_n231_, new_n230_, keyIn_0_13 );
not g124 ( new_n232_, keyIn_0_13 );
not g125 ( new_n233_, N56 );
or g126 ( new_n234_, new_n232_, new_n233_, N60 );
and g127 ( new_n235_, new_n231_, new_n234_ );
and g128 ( new_n236_, new_n227_, new_n228_, new_n235_ );
not g129 ( new_n237_, new_n236_ );
and g130 ( new_n238_, new_n153_, N108 );
or g131 ( new_n239_, new_n238_, new_n152_ );
not g132 ( new_n240_, new_n154_ );
and g133 ( new_n241_, new_n239_, new_n240_ );
and g134 ( new_n242_, new_n188_, new_n241_ );
not g135 ( new_n243_, new_n242_ );
or g136 ( new_n244_, new_n188_, new_n241_ );
not g137 ( new_n245_, keyIn_0_17 );
not g138 ( new_n246_, N112 );
and g139 ( new_n247_, new_n246_, N108 );
or g140 ( new_n248_, new_n247_, new_n245_ );
or g141 ( new_n249_, new_n149_, keyIn_0_17, N112 );
and g142 ( new_n250_, new_n248_, new_n249_ );
and g143 ( new_n251_, new_n243_, new_n244_, new_n250_ );
not g144 ( new_n252_, new_n251_ );
and g145 ( new_n253_, new_n237_, new_n252_ );
and g146 ( new_n254_, new_n206_, new_n253_, new_n225_, new_n218_ );
not g147 ( new_n255_, keyIn_0_27 );
and g148 ( new_n256_, new_n188_, new_n136_ );
not g149 ( new_n257_, new_n256_ );
or g150 ( new_n258_, new_n188_, new_n136_ );
and g151 ( new_n259_, new_n257_, new_n258_ );
and g152 ( new_n260_, new_n135_, keyIn_0_0 );
not g153 ( new_n261_, new_n260_ );
or g154 ( new_n262_, new_n135_, keyIn_0_0 );
and g155 ( new_n263_, new_n261_, new_n262_ );
or g156 ( new_n264_, new_n263_, N8 );
not g157 ( new_n265_, new_n264_ );
and g158 ( new_n266_, new_n265_, keyIn_0_6 );
not g159 ( new_n267_, new_n266_ );
or g160 ( new_n268_, new_n265_, keyIn_0_6 );
and g161 ( new_n269_, new_n267_, new_n268_ );
or g162 ( new_n270_, new_n259_, new_n269_ );
and g163 ( new_n271_, new_n270_, new_n255_ );
not g164 ( new_n272_, new_n259_ );
not g165 ( new_n273_, new_n269_ );
and g166 ( new_n274_, new_n272_, keyIn_0_27, new_n273_ );
or g167 ( new_n275_, new_n271_, new_n274_ );
not g168 ( new_n276_, keyIn_0_30 );
and g169 ( new_n277_, new_n188_, new_n148_ );
not g170 ( new_n278_, new_n277_ );
or g171 ( new_n279_, new_n188_, new_n148_ );
and g172 ( new_n280_, new_n278_, new_n279_ );
and g173 ( new_n281_, new_n143_, keyIn_0_3 );
not g174 ( new_n282_, new_n281_ );
or g175 ( new_n283_, new_n143_, keyIn_0_3 );
and g176 ( new_n284_, new_n282_, new_n283_ );
or g177 ( new_n285_, new_n284_, N47 );
not g178 ( new_n286_, new_n285_ );
and g179 ( new_n287_, new_n286_, keyIn_0_12 );
not g180 ( new_n288_, new_n287_ );
or g181 ( new_n289_, new_n286_, keyIn_0_12 );
and g182 ( new_n290_, new_n288_, new_n289_ );
or g183 ( new_n291_, new_n280_, new_n290_ );
and g184 ( new_n292_, new_n291_, new_n276_ );
not g185 ( new_n293_, new_n280_ );
not g186 ( new_n294_, new_n290_ );
and g187 ( new_n295_, new_n293_, keyIn_0_30, new_n294_ );
or g188 ( new_n296_, new_n292_, new_n295_ );
and g189 ( new_n297_, new_n185_, new_n254_, new_n275_, new_n296_ );
not g190 ( new_n298_, new_n297_ );
and g191 ( new_n299_, new_n298_, new_n163_ );
and g192 ( new_n300_, new_n275_, new_n296_ );
and g193 ( new_n301_, new_n300_, keyIn_0_32, new_n185_, new_n254_ );
or g194 ( new_n302_, new_n299_, new_n301_ );
and g195 ( new_n303_, new_n302_, keyIn_0_38 );
not g196 ( new_n304_, keyIn_0_38 );
or g197 ( new_n305_, new_n297_, keyIn_0_32 );
not g198 ( new_n306_, new_n301_ );
and g199 ( new_n307_, new_n306_, new_n305_ );
and g200 ( new_n308_, new_n307_, new_n304_ );
or g201 ( N329, new_n303_, new_n308_ );
not g202 ( new_n310_, keyIn_0_48 );
not g203 ( new_n311_, keyIn_0_46 );
not g204 ( new_n312_, keyIn_0_42 );
and g205 ( new_n313_, new_n302_, keyIn_0_37 );
not g206 ( new_n314_, keyIn_0_37 );
and g207 ( new_n315_, new_n306_, new_n305_, new_n314_ );
or g208 ( new_n316_, new_n313_, new_n315_ );
and g209 ( new_n317_, new_n316_, new_n205_ );
or g210 ( new_n318_, new_n307_, new_n314_ );
not g211 ( new_n319_, new_n315_ );
and g212 ( new_n320_, new_n318_, new_n204_, new_n319_ );
or g213 ( new_n321_, new_n317_, new_n320_ );
and g214 ( new_n322_, new_n321_, new_n312_ );
and g215 ( new_n323_, new_n318_, new_n319_ );
or g216 ( new_n324_, new_n323_, new_n204_ );
not g217 ( new_n325_, new_n320_ );
and g218 ( new_n326_, new_n324_, keyIn_0_42, new_n325_ );
or g219 ( new_n327_, new_n322_, new_n326_ );
not g220 ( new_n328_, keyIn_0_35 );
not g221 ( new_n329_, keyIn_0_14 );
not g222 ( new_n330_, N79 );
and g223 ( new_n331_, new_n203_, new_n330_ );
and g224 ( new_n332_, new_n331_, new_n329_ );
not g225 ( new_n333_, new_n331_ );
and g226 ( new_n334_, new_n333_, keyIn_0_14 );
or g227 ( new_n335_, new_n334_, new_n332_ );
and g228 ( new_n336_, new_n197_, new_n198_, new_n335_ );
and g229 ( new_n337_, new_n336_, new_n328_ );
not g230 ( new_n338_, new_n337_ );
or g231 ( new_n339_, new_n336_, new_n328_ );
and g232 ( new_n340_, new_n338_, new_n339_ );
not g233 ( new_n341_, new_n340_ );
and g234 ( new_n342_, new_n327_, new_n311_, new_n341_ );
not g235 ( new_n343_, new_n342_ );
and g236 ( new_n344_, new_n327_, new_n341_ );
or g237 ( new_n345_, new_n344_, new_n311_ );
not g238 ( new_n346_, keyIn_0_43 );
and g239 ( new_n347_, new_n323_, new_n251_ );
not g240 ( new_n348_, new_n347_ );
or g241 ( new_n349_, new_n323_, new_n251_ );
and g242 ( new_n350_, new_n348_, new_n346_, new_n349_ );
not g243 ( new_n351_, new_n350_ );
not g244 ( new_n352_, keyIn_0_31 );
not g245 ( new_n353_, N115 );
and g246 ( new_n354_, new_n243_, new_n244_ );
and g247 ( new_n355_, new_n354_, N108, new_n353_ );
not g248 ( new_n356_, new_n355_ );
and g249 ( new_n357_, new_n356_, new_n352_ );
and g250 ( new_n358_, new_n355_, keyIn_0_31 );
or g251 ( new_n359_, new_n357_, new_n358_ );
and g252 ( new_n360_, new_n348_, new_n349_ );
or g253 ( new_n361_, new_n360_, new_n346_ );
and g254 ( new_n362_, new_n361_, new_n351_, new_n359_ );
or g255 ( new_n363_, new_n323_, new_n236_ );
and g256 ( new_n364_, new_n323_, new_n236_ );
not g257 ( new_n365_, new_n364_ );
not g258 ( new_n366_, N66 );
and g259 ( new_n367_, new_n227_, N56, new_n366_, new_n228_ );
and g260 ( new_n368_, new_n365_, new_n363_, new_n367_ );
or g261 ( new_n369_, new_n323_, new_n192_ );
not g262 ( new_n370_, N92 );
and g263 ( new_n371_, new_n370_, N82 );
or g264 ( new_n372_, new_n371_, keyIn_0_15 );
not g265 ( new_n373_, keyIn_0_15 );
or g266 ( new_n374_, new_n373_, new_n137_, N92 );
and g267 ( new_n375_, new_n190_, new_n191_, new_n372_, new_n374_ );
and g268 ( new_n376_, new_n375_, keyIn_0_36 );
not g269 ( new_n377_, new_n376_ );
or g270 ( new_n378_, new_n375_, keyIn_0_36 );
and g271 ( new_n379_, new_n377_, new_n378_ );
not g272 ( new_n380_, new_n379_ );
and g273 ( new_n381_, new_n323_, new_n192_ );
not g274 ( new_n382_, new_n381_ );
and g275 ( new_n383_, new_n382_, new_n369_, new_n380_ );
or g276 ( new_n384_, new_n323_, new_n217_ );
not g277 ( new_n385_, N40 );
and g278 ( new_n386_, new_n215_, new_n385_ );
not g279 ( new_n387_, new_n386_ );
and g280 ( new_n388_, new_n387_, keyIn_0_11 );
not g281 ( new_n389_, keyIn_0_11 );
and g282 ( new_n390_, new_n386_, new_n389_ );
or g283 ( new_n391_, new_n388_, new_n390_ );
and g284 ( new_n392_, new_n210_, new_n391_ );
and g285 ( new_n393_, new_n392_, keyIn_0_34 );
not g286 ( new_n394_, new_n393_ );
or g287 ( new_n395_, new_n392_, keyIn_0_34 );
and g288 ( new_n396_, new_n394_, new_n395_ );
not g289 ( new_n397_, new_n396_ );
and g290 ( new_n398_, new_n323_, new_n217_ );
not g291 ( new_n399_, new_n398_ );
and g292 ( new_n400_, new_n399_, new_n384_, new_n397_ );
or g293 ( new_n401_, new_n368_, new_n383_, new_n400_ );
or g294 ( new_n402_, new_n362_, new_n401_ );
not g295 ( new_n403_, new_n402_ );
and g296 ( new_n404_, new_n345_, new_n403_ );
not g297 ( new_n405_, keyIn_0_45 );
not g298 ( new_n406_, keyIn_0_41 );
or g299 ( new_n407_, new_n323_, new_n296_ );
and g300 ( new_n408_, new_n318_, new_n296_, new_n319_ );
not g301 ( new_n409_, new_n408_ );
and g302 ( new_n410_, new_n407_, new_n409_ );
or g303 ( new_n411_, new_n410_, new_n406_ );
and g304 ( new_n412_, new_n407_, new_n406_, new_n409_ );
not g305 ( new_n413_, new_n412_ );
and g306 ( new_n414_, new_n411_, new_n413_ );
or g307 ( new_n415_, new_n280_, N53, new_n284_ );
or g308 ( new_n416_, new_n414_, new_n415_ );
and g309 ( new_n417_, new_n416_, new_n405_ );
not g310 ( new_n418_, new_n414_ );
not g311 ( new_n419_, new_n415_ );
and g312 ( new_n420_, new_n418_, keyIn_0_45, new_n419_ );
or g313 ( new_n421_, new_n417_, new_n420_ );
not g314 ( new_n422_, keyIn_0_40 );
not g315 ( new_n423_, new_n185_ );
and g316 ( new_n424_, new_n323_, new_n423_ );
and g317 ( new_n425_, new_n316_, new_n185_ );
or g318 ( new_n426_, new_n425_, new_n424_ );
and g319 ( new_n427_, new_n426_, new_n422_ );
not g320 ( new_n428_, keyIn_0_33 );
not g321 ( new_n429_, N27 );
and g322 ( new_n430_, new_n180_, N17, new_n429_, new_n182_ );
or g323 ( new_n431_, new_n430_, new_n428_ );
and g324 ( new_n432_, new_n430_, new_n428_ );
not g325 ( new_n433_, new_n432_ );
and g326 ( new_n434_, new_n433_, new_n431_ );
not g327 ( new_n435_, new_n424_ );
not g328 ( new_n436_, new_n425_ );
and g329 ( new_n437_, new_n436_, keyIn_0_40, new_n435_ );
or g330 ( new_n438_, new_n427_, new_n437_, new_n434_ );
or g331 ( new_n439_, new_n323_, new_n275_ );
and g332 ( new_n440_, new_n323_, new_n275_ );
not g333 ( new_n441_, new_n440_ );
and g334 ( new_n442_, new_n441_, new_n439_ );
and g335 ( new_n443_, new_n442_, keyIn_0_39 );
not g336 ( new_n444_, new_n443_ );
not g337 ( new_n445_, keyIn_0_28 );
or g338 ( new_n446_, new_n259_, N14, new_n263_ );
and g339 ( new_n447_, new_n446_, new_n445_ );
not g340 ( new_n448_, new_n446_ );
and g341 ( new_n449_, new_n448_, keyIn_0_28 );
or g342 ( new_n450_, new_n449_, new_n447_ );
or g343 ( new_n451_, new_n442_, keyIn_0_39 );
and g344 ( new_n452_, new_n444_, new_n450_, new_n451_ );
not g345 ( new_n453_, new_n452_ );
not g346 ( new_n454_, keyIn_0_47 );
and g347 ( new_n455_, new_n316_, new_n224_ );
and g348 ( new_n456_, new_n323_, new_n225_ );
or g349 ( new_n457_, new_n455_, new_n456_ );
not g350 ( new_n458_, new_n457_ );
not g351 ( new_n459_, N105 );
and g352 ( new_n460_, new_n459_, N95 );
or g353 ( new_n461_, new_n460_, keyIn_0_16 );
not g354 ( new_n462_, keyIn_0_16 );
not g355 ( new_n463_, N95 );
or g356 ( new_n464_, new_n462_, new_n463_, N105 );
and g357 ( new_n465_, new_n461_, new_n464_ );
and g358 ( new_n466_, new_n223_, new_n465_ );
not g359 ( new_n467_, new_n466_ );
or g360 ( new_n468_, new_n458_, new_n467_ );
and g361 ( new_n469_, new_n468_, new_n454_ );
and g362 ( new_n470_, new_n457_, keyIn_0_47, new_n466_ );
or g363 ( new_n471_, new_n469_, new_n470_ );
and g364 ( new_n472_, new_n471_, new_n453_, new_n438_ );
and g365 ( new_n473_, new_n404_, new_n343_, new_n421_, new_n472_ );
or g366 ( new_n474_, new_n473_, new_n310_ );
and g367 ( new_n475_, new_n324_, new_n325_ );
or g368 ( new_n476_, new_n475_, keyIn_0_42 );
not g369 ( new_n477_, new_n326_ );
and g370 ( new_n478_, new_n476_, new_n477_ );
or g371 ( new_n479_, new_n478_, new_n340_ );
and g372 ( new_n480_, new_n479_, keyIn_0_46 );
or g373 ( new_n481_, new_n480_, new_n342_, new_n402_ );
not g374 ( new_n482_, new_n421_ );
not g375 ( new_n483_, new_n472_ );
or g376 ( new_n484_, new_n482_, new_n483_, new_n481_, keyIn_0_48 );
and g377 ( N370, new_n474_, new_n484_ );
not g378 ( new_n486_, keyIn_0_58 );
not g379 ( new_n487_, keyIn_0_55 );
or g380 ( new_n488_, N370, keyIn_0_49 );
not g381 ( new_n489_, keyIn_0_49 );
not g382 ( new_n490_, new_n473_ );
and g383 ( new_n491_, new_n490_, keyIn_0_48 );
not g384 ( new_n492_, new_n484_ );
or g385 ( new_n493_, new_n491_, new_n492_, new_n489_ );
and g386 ( new_n494_, new_n488_, N105, new_n493_ );
or g387 ( new_n495_, new_n494_, keyIn_0_52 );
and g388 ( new_n496_, new_n488_, keyIn_0_52, N105, new_n493_ );
not g389 ( new_n497_, new_n496_ );
and g390 ( new_n498_, new_n495_, new_n497_ );
and g391 ( new_n499_, new_n307_, N99 );
and g392 ( new_n500_, new_n157_, keyIn_0_19 );
not g393 ( new_n501_, new_n500_ );
or g394 ( new_n502_, new_n157_, keyIn_0_19 );
and g395 ( new_n503_, new_n501_, new_n502_ );
not g396 ( new_n504_, new_n503_ );
and g397 ( new_n505_, new_n504_, N89 );
or g398 ( new_n506_, new_n499_, new_n463_, new_n505_ );
or g399 ( new_n507_, new_n498_, new_n506_ );
and g400 ( new_n508_, new_n507_, new_n487_ );
not g401 ( new_n509_, new_n498_ );
not g402 ( new_n510_, new_n506_ );
and g403 ( new_n511_, new_n509_, keyIn_0_55, new_n510_ );
or g404 ( new_n512_, new_n508_, new_n511_ );
not g405 ( new_n513_, keyIn_0_50 );
and g406 ( new_n514_, new_n488_, N66, new_n493_ );
or g407 ( new_n515_, new_n514_, new_n513_ );
not g408 ( new_n516_, new_n515_ );
and g409 ( new_n517_, new_n514_, new_n513_ );
and g410 ( new_n518_, new_n307_, N60 );
not g411 ( new_n519_, keyIn_0_24 );
and g412 ( new_n520_, new_n504_, N50 );
and g413 ( new_n521_, new_n520_, new_n519_ );
or g414 ( new_n522_, new_n520_, new_n519_ );
not g415 ( new_n523_, new_n522_ );
or g416 ( new_n524_, new_n518_, new_n233_, new_n521_, new_n523_ );
or g417 ( new_n525_, new_n516_, new_n517_, new_n524_ );
and g418 ( new_n526_, new_n488_, new_n493_ );
and g419 ( new_n527_, new_n526_, N53 );
and g420 ( new_n528_, new_n307_, N47 );
and g421 ( new_n529_, new_n504_, N37 );
or g422 ( new_n530_, new_n529_, keyIn_0_23 );
not g423 ( new_n531_, new_n530_ );
and g424 ( new_n532_, new_n529_, keyIn_0_23 );
or g425 ( new_n533_, new_n528_, new_n143_, new_n531_, new_n532_ );
or g426 ( new_n534_, new_n527_, new_n533_ );
and g427 ( new_n535_, new_n525_, new_n534_ );
and g428 ( new_n536_, new_n526_, N40 );
and g429 ( new_n537_, new_n307_, N34 );
and g430 ( new_n538_, new_n504_, N24 );
or g431 ( new_n539_, new_n536_, new_n108_, new_n537_, new_n538_ );
and g432 ( new_n540_, new_n526_, N27 );
and g433 ( new_n541_, new_n307_, N21 );
not g434 ( new_n542_, keyIn_0_22 );
and g435 ( new_n543_, new_n504_, N11 );
and g436 ( new_n544_, new_n543_, new_n542_ );
or g437 ( new_n545_, new_n543_, new_n542_ );
not g438 ( new_n546_, new_n545_ );
or g439 ( new_n547_, new_n541_, new_n123_, new_n544_, new_n546_ );
or g440 ( new_n548_, new_n540_, new_n547_ );
and g441 ( new_n549_, new_n539_, new_n548_ );
and g442 ( new_n550_, new_n488_, N115, new_n493_ );
not g443 ( new_n551_, keyIn_0_44 );
and g444 ( new_n552_, new_n307_, N112 );
and g445 ( new_n553_, new_n552_, new_n551_ );
not g446 ( new_n554_, new_n553_ );
or g447 ( new_n555_, new_n552_, new_n551_ );
or g448 ( new_n556_, new_n503_, new_n153_ );
and g449 ( new_n557_, new_n554_, N108, new_n555_, new_n556_ );
not g450 ( new_n558_, new_n557_ );
or g451 ( new_n559_, new_n550_, new_n558_ );
and g452 ( new_n560_, new_n559_, keyIn_0_56 );
not g453 ( new_n561_, keyIn_0_56 );
not g454 ( new_n562_, new_n550_ );
and g455 ( new_n563_, new_n562_, new_n561_, new_n557_ );
or g456 ( new_n564_, new_n560_, new_n563_ );
and g457 ( new_n565_, new_n488_, N92, new_n493_ );
and g458 ( new_n566_, new_n307_, N86 );
not g459 ( new_n567_, keyIn_0_26 );
and g460 ( new_n568_, new_n504_, N76 );
or g461 ( new_n569_, new_n568_, new_n567_ );
not g462 ( new_n570_, new_n569_ );
and g463 ( new_n571_, new_n568_, new_n567_ );
or g464 ( new_n572_, new_n566_, new_n137_, new_n570_, new_n571_ );
or g465 ( new_n573_, new_n565_, new_n572_ );
and g466 ( new_n574_, new_n573_, keyIn_0_54 );
not g467 ( new_n575_, keyIn_0_54 );
not g468 ( new_n576_, new_n565_ );
not g469 ( new_n577_, new_n572_ );
and g470 ( new_n578_, new_n576_, new_n575_, new_n577_ );
or g471 ( new_n579_, new_n574_, new_n578_ );
not g472 ( new_n580_, keyIn_0_51 );
not g473 ( new_n581_, N370 );
and g474 ( new_n582_, new_n581_, new_n489_ );
and g475 ( new_n583_, N370, keyIn_0_49 );
or g476 ( new_n584_, new_n582_, new_n583_, new_n330_ );
and g477 ( new_n585_, new_n584_, new_n580_ );
and g478 ( new_n586_, new_n526_, keyIn_0_51, N79 );
and g479 ( new_n587_, new_n307_, N73 );
not g480 ( new_n588_, keyIn_0_25 );
and g481 ( new_n589_, new_n504_, N63 );
and g482 ( new_n590_, new_n589_, new_n588_ );
or g483 ( new_n591_, new_n589_, new_n588_ );
not g484 ( new_n592_, new_n591_ );
or g485 ( new_n593_, new_n587_, new_n115_, new_n590_, new_n592_ );
or g486 ( new_n594_, new_n585_, new_n586_, new_n593_ );
and g487 ( new_n595_, new_n579_, new_n594_ );
and g488 ( new_n596_, new_n595_, new_n535_, new_n549_, new_n564_ );
and g489 ( new_n597_, new_n596_, new_n512_ );
not g490 ( new_n598_, new_n597_ );
and g491 ( new_n599_, new_n598_, new_n486_ );
and g492 ( new_n600_, new_n597_, keyIn_0_58 );
or g493 ( new_n601_, new_n599_, new_n600_ );
and g494 ( new_n602_, new_n526_, N14 );
and g495 ( new_n603_, new_n307_, N8 );
and g496 ( new_n604_, new_n504_, N1 );
or g497 ( new_n605_, new_n602_, new_n135_, new_n603_, new_n604_ );
and g498 ( new_n606_, new_n605_, keyIn_0_53 );
not g499 ( new_n607_, new_n606_ );
or g500 ( new_n608_, new_n605_, keyIn_0_53 );
and g501 ( new_n609_, new_n607_, new_n608_ );
not g502 ( new_n610_, new_n609_ );
and g503 ( new_n611_, new_n610_, keyIn_0_57 );
not g504 ( new_n612_, keyIn_0_57 );
and g505 ( new_n613_, new_n609_, new_n612_ );
or g506 ( new_n614_, new_n611_, new_n613_ );
and g507 ( N421, new_n601_, new_n614_ );
not g508 ( new_n616_, new_n517_ );
not g509 ( new_n617_, new_n524_ );
and g510 ( new_n618_, new_n616_, new_n515_, new_n617_ );
not g511 ( new_n619_, new_n549_ );
not g512 ( new_n620_, new_n534_ );
and g513 ( new_n621_, new_n539_, new_n620_ );
not g514 ( new_n622_, new_n621_ );
and g515 ( new_n623_, new_n622_, keyIn_0_60 );
not g516 ( new_n624_, new_n623_ );
or g517 ( new_n625_, new_n622_, keyIn_0_60 );
and g518 ( new_n626_, new_n624_, new_n625_ );
or g519 ( new_n627_, new_n626_, new_n618_, new_n619_ );
and g520 ( new_n628_, new_n627_, keyIn_0_62 );
not g521 ( new_n629_, keyIn_0_62 );
not g522 ( new_n630_, new_n626_ );
and g523 ( new_n631_, new_n630_, new_n629_, new_n525_, new_n549_ );
or g524 ( N430, new_n628_, new_n631_ );
not g525 ( new_n633_, keyIn_0_63 );
not g526 ( new_n634_, keyIn_0_59 );
not g527 ( new_n635_, new_n574_ );
not g528 ( new_n636_, new_n578_ );
and g529 ( new_n637_, new_n635_, new_n634_, new_n636_ );
not g530 ( new_n638_, new_n637_ );
and g531 ( new_n639_, new_n579_, keyIn_0_59 );
not g532 ( new_n640_, new_n639_ );
and g533 ( new_n641_, new_n640_, keyIn_0_61, new_n535_, new_n638_ );
not g534 ( new_n642_, keyIn_0_61 );
or g535 ( new_n643_, new_n618_, new_n620_ );
or g536 ( new_n644_, new_n639_, new_n643_, new_n637_ );
and g537 ( new_n645_, new_n644_, new_n642_ );
not g538 ( new_n646_, new_n594_ );
and g539 ( new_n647_, new_n535_, new_n539_, new_n646_ );
or g540 ( new_n648_, new_n647_, new_n619_ );
or g541 ( new_n649_, new_n645_, new_n641_, new_n648_ );
and g542 ( new_n650_, new_n649_, new_n633_ );
not g543 ( new_n651_, new_n641_ );
not g544 ( new_n652_, new_n645_ );
not g545 ( new_n653_, new_n648_ );
and g546 ( new_n654_, new_n652_, keyIn_0_63, new_n651_, new_n653_ );
or g547 ( N431, new_n650_, new_n654_ );
not g548 ( new_n656_, new_n548_ );
not g549 ( new_n657_, new_n508_ );
not g550 ( new_n658_, new_n511_ );
and g551 ( new_n659_, new_n579_, new_n534_, new_n539_ );
and g552 ( new_n660_, new_n657_, new_n658_, new_n659_ );
or g553 ( N432, new_n626_, new_n656_, new_n647_, new_n660_ );
endmodule