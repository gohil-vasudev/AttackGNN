module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n173_, new_n220_, new_n419_, new_n214_, new_n451_, new_n424_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n317_, new_n344_, new_n287_, new_n427_, new_n234_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n150_, new_n137_, new_n183_, new_n463_, new_n303_, new_n351_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n305_, new_n420_, new_n423_, new_n205_, new_n141_, new_n206_, new_n254_, new_n355_, new_n353_, new_n432_, new_n256_, new_n452_, new_n381_, new_n388_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n314_, new_n363_, new_n165_, new_n477_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n343_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n244_, new_n172_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n371_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n362_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n130_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n310_, new_n144_, new_n275_, new_n352_, new_n177_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n125_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n182_, new_n407_, new_n480_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n360_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n332_, new_n453_, new_n163_, new_n440_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n307_, new_n190_, new_n408_, new_n470_, new_n213_, new_n433_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n129_, new_n412_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n358_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n406_, new_n356_, new_n229_, new_n464_, new_n204_, new_n181_, new_n405_;

nand g000 ( new_n119_, N29, N42, N75 );
not g001 ( N388, new_n119_ );
nand g002 ( new_n121_, N29, N36, N80 );
not g003 ( N389, new_n121_ );
nand g004 ( new_n123_, N29, N36, N42 );
not g005 ( N390, new_n123_ );
nand g006 ( new_n125_, N85, N86 );
not g007 ( N391, new_n125_ );
nand g008 ( new_n127_, N1, N8, N13, N17 );
not g009 ( N418, new_n127_ );
nand g010 ( new_n129_, N1, N26 );
nand g011 ( new_n130_, N13, N17 );
nor g012 ( new_n131_, new_n129_, new_n130_ );
nand g013 ( N419, new_n131_, new_n123_ );
nand g014 ( N420, N59, N75, N80 );
nand g015 ( N421, N36, N59, N80 );
nand g016 ( N422, N36, N42, N59 );
not g017 ( new_n136_, N90 );
nor g018 ( new_n137_, N87, N88 );
nor g019 ( N423, new_n137_, new_n136_ );
nand g020 ( N446, new_n131_, N390 );
nand g021 ( new_n140_, keyIn_0_0, N1, N26, N51 );
not g022 ( new_n141_, keyIn_0_0 );
nand g023 ( new_n142_, N1, N26, N51 );
nand g024 ( new_n143_, new_n142_, new_n141_ );
nand g025 ( new_n144_, new_n143_, new_n140_ );
not g026 ( N447, new_n144_ );
nand g027 ( new_n146_, N1, N8, N13, N55 );
nand g028 ( new_n147_, N29, N68 );
nor g029 ( N448, new_n146_, new_n147_ );
not g030 ( new_n149_, N74 );
nand g031 ( new_n150_, N59, N68 );
nor g032 ( N449, new_n146_, new_n149_, new_n150_ );
not g033 ( new_n152_, N89 );
nor g034 ( N450, new_n137_, new_n152_ );
xor g035 ( new_n154_, N111, N116 );
xnor g036 ( new_n155_, N121, N126 );
xnor g037 ( new_n156_, new_n154_, new_n155_ );
xnor g038 ( new_n157_, new_n156_, N135 );
xnor g039 ( new_n158_, N91, N96 );
xnor g040 ( new_n159_, N101, N106 );
xnor g041 ( new_n160_, new_n158_, new_n159_ );
xnor g042 ( new_n161_, new_n160_, N130 );
xnor g043 ( N767, new_n157_, new_n161_ );
xor g044 ( new_n163_, N183, N189 );
xnor g045 ( new_n164_, N195, N201 );
xnor g046 ( new_n165_, new_n163_, new_n164_ );
xnor g047 ( new_n166_, new_n165_, N207 );
xnor g048 ( new_n167_, N159, N165 );
xnor g049 ( new_n168_, N171, N177 );
xnor g050 ( new_n169_, new_n167_, new_n168_ );
xnor g051 ( new_n170_, new_n169_, N130 );
xnor g052 ( N768, new_n166_, new_n170_ );
not g053 ( new_n172_, keyIn_0_23 );
not g054 ( new_n173_, keyIn_0_21 );
not g055 ( new_n174_, keyIn_0_16 );
not g056 ( new_n175_, keyIn_0_10 );
nand g057 ( new_n176_, new_n144_, keyIn_0_6 );
not g058 ( new_n177_, keyIn_0_6 );
nand g059 ( new_n178_, new_n143_, new_n177_, new_n140_ );
nand g060 ( new_n179_, new_n176_, new_n178_ );
nand g061 ( new_n180_, new_n179_, new_n175_ );
nand g062 ( new_n181_, new_n176_, keyIn_0_10, new_n178_ );
nand g063 ( new_n182_, new_n180_, new_n181_ );
nand g064 ( new_n183_, N59, N156 );
xnor g065 ( new_n184_, new_n183_, keyIn_0_3 );
nand g066 ( new_n185_, new_n182_, new_n184_ );
not g067 ( new_n186_, new_n185_ );
nand g068 ( new_n187_, new_n186_, new_n174_, N17 );
nand g069 ( new_n188_, new_n186_, N17 );
nand g070 ( new_n189_, new_n188_, keyIn_0_16 );
nand g071 ( new_n190_, new_n189_, N1, new_n187_ );
nand g072 ( new_n191_, new_n190_, N153 );
not g073 ( new_n192_, keyIn_0_15 );
not g074 ( new_n193_, new_n183_ );
not g075 ( new_n194_, keyIn_0_4 );
nor g076 ( new_n195_, N17, N42 );
xnor g077 ( new_n196_, new_n195_, new_n194_ );
nand g078 ( new_n197_, N17, N42 );
xnor g079 ( new_n198_, new_n197_, keyIn_0_5 );
nand g080 ( new_n199_, new_n196_, new_n198_ );
nand g081 ( new_n200_, new_n199_, keyIn_0_9 );
not g082 ( new_n201_, keyIn_0_9 );
nand g083 ( new_n202_, new_n196_, new_n201_, new_n198_ );
nand g084 ( new_n203_, new_n200_, new_n202_ );
nand g085 ( new_n204_, new_n182_, new_n192_, new_n193_, new_n203_ );
nand g086 ( new_n205_, new_n182_, new_n193_, new_n203_ );
nand g087 ( new_n206_, new_n205_, keyIn_0_15 );
nand g088 ( new_n207_, new_n206_, new_n204_ );
not g089 ( new_n208_, keyIn_0_11 );
nand g090 ( new_n209_, N42, N59, N75 );
xnor g091 ( new_n210_, new_n209_, keyIn_0_2 );
xnor g092 ( new_n211_, new_n210_, keyIn_0_8 );
not g093 ( new_n212_, keyIn_0_1 );
nand g094 ( new_n213_, N1, N8, N17, N51 );
xnor g095 ( new_n214_, new_n213_, new_n212_ );
xnor g096 ( new_n215_, new_n214_, keyIn_0_7 );
nand g097 ( new_n216_, new_n215_, new_n211_ );
xnor g098 ( new_n217_, new_n216_, new_n208_ );
nand g099 ( new_n218_, new_n207_, new_n217_, keyIn_0_17 );
not g100 ( new_n219_, keyIn_0_17 );
nand g101 ( new_n220_, new_n207_, new_n217_ );
nand g102 ( new_n221_, new_n220_, new_n219_ );
nand g103 ( new_n222_, new_n221_, new_n218_ );
nand g104 ( new_n223_, new_n222_, N126 );
nand g105 ( new_n224_, new_n223_, new_n173_, new_n191_ );
nand g106 ( new_n225_, new_n223_, new_n191_ );
nand g107 ( new_n226_, new_n225_, keyIn_0_21 );
not g108 ( new_n227_, N268 );
not g109 ( new_n228_, keyIn_0_14 );
nand g110 ( new_n229_, N29, N75, N80 );
not g111 ( new_n230_, new_n229_ );
nand g112 ( new_n231_, new_n182_, new_n228_, N55, new_n230_ );
nand g113 ( new_n232_, new_n182_, N55, new_n230_ );
nand g114 ( new_n233_, new_n232_, keyIn_0_14 );
nand g115 ( new_n234_, new_n233_, new_n227_, new_n231_ );
xnor g116 ( new_n235_, new_n234_, keyIn_0_19 );
nand g117 ( new_n236_, new_n226_, new_n224_, new_n235_ );
nand g118 ( new_n237_, new_n236_, new_n172_ );
nand g119 ( new_n238_, new_n226_, keyIn_0_23, new_n224_, new_n235_ );
nand g120 ( new_n239_, new_n237_, new_n238_ );
nand g121 ( new_n240_, new_n239_, N201 );
not g122 ( new_n241_, N201 );
nand g123 ( new_n242_, new_n237_, new_n241_, new_n238_ );
nand g124 ( new_n243_, new_n240_, new_n242_ );
not g125 ( new_n244_, new_n243_ );
nand g126 ( new_n245_, new_n244_, N261 );
not g127 ( new_n246_, N261 );
nand g128 ( new_n247_, new_n243_, new_n246_ );
nand g129 ( new_n248_, new_n245_, new_n247_, N219 );
nand g130 ( new_n249_, new_n244_, N228 );
not g131 ( new_n250_, new_n240_ );
nand g132 ( new_n251_, new_n250_, N237 );
nand g133 ( new_n252_, new_n239_, N246 );
nand g134 ( new_n253_, N42, N72, N73 );
nor g135 ( new_n254_, new_n146_, new_n253_, new_n150_ );
not g136 ( new_n255_, new_n254_ );
nor g137 ( new_n256_, new_n255_, new_n241_ );
nand g138 ( new_n257_, N255, N267 );
nand g139 ( new_n258_, N121, N210 );
nand g140 ( new_n259_, new_n257_, new_n258_ );
nor g141 ( new_n260_, new_n256_, new_n259_ );
nand g142 ( new_n261_, new_n251_, new_n252_, new_n260_ );
not g143 ( new_n262_, new_n261_ );
nand g144 ( new_n263_, new_n248_, new_n249_, new_n262_ );
xor g145 ( N850, new_n263_, keyIn_0_27 );
not g146 ( new_n265_, keyIn_0_25 );
not g147 ( new_n266_, N189 );
nand g148 ( new_n267_, new_n222_, N116 );
nand g149 ( new_n268_, new_n190_, N146 );
nand g150 ( new_n269_, new_n268_, new_n234_ );
not g151 ( new_n270_, new_n269_ );
nand g152 ( new_n271_, new_n270_, new_n266_, new_n267_ );
not g153 ( new_n272_, N195 );
not g154 ( new_n273_, keyIn_0_22 );
not g155 ( new_n274_, keyIn_0_20 );
nand g156 ( new_n275_, new_n222_, N121 );
nand g157 ( new_n276_, new_n190_, N149 );
nand g158 ( new_n277_, new_n275_, new_n274_, new_n276_ );
nand g159 ( new_n278_, new_n275_, new_n276_ );
nand g160 ( new_n279_, new_n278_, keyIn_0_20 );
xor g161 ( new_n280_, new_n234_, keyIn_0_18 );
nand g162 ( new_n281_, new_n279_, new_n273_, new_n277_, new_n280_ );
nand g163 ( new_n282_, new_n279_, new_n277_, new_n280_ );
nand g164 ( new_n283_, new_n282_, keyIn_0_22 );
nand g165 ( new_n284_, new_n283_, new_n272_, new_n281_ );
nand g166 ( new_n285_, new_n250_, new_n265_, new_n271_, new_n284_ );
nand g167 ( new_n286_, new_n284_, new_n239_, N201, new_n271_ );
nand g168 ( new_n287_, new_n286_, keyIn_0_25 );
nand g169 ( new_n288_, new_n285_, new_n287_ );
not g170 ( new_n289_, keyIn_0_24 );
nand g171 ( new_n290_, new_n242_, new_n284_, N261, new_n271_ );
not g172 ( new_n291_, new_n290_ );
nand g173 ( new_n292_, new_n291_, new_n289_ );
nand g174 ( new_n293_, new_n290_, keyIn_0_24 );
nand g175 ( new_n294_, new_n283_, new_n281_ );
nand g176 ( new_n295_, new_n294_, N195, new_n271_ );
nand g177 ( new_n296_, new_n270_, new_n267_ );
nand g178 ( new_n297_, new_n296_, N189 );
nand g179 ( new_n298_, new_n295_, new_n297_ );
not g180 ( new_n299_, new_n298_ );
nand g181 ( new_n300_, new_n299_, new_n293_ );
not g182 ( new_n301_, new_n300_ );
nand g183 ( new_n302_, new_n301_, keyIn_0_26, new_n288_, new_n292_ );
not g184 ( new_n303_, keyIn_0_26 );
nand g185 ( new_n304_, new_n288_, new_n292_, new_n293_, new_n299_ );
nand g186 ( new_n305_, new_n304_, new_n303_ );
nand g187 ( new_n306_, new_n305_, new_n302_ );
nand g188 ( new_n307_, new_n222_, N111 );
nand g189 ( new_n308_, new_n190_, N143 );
nand g190 ( new_n309_, new_n308_, new_n234_ );
not g191 ( new_n310_, new_n309_ );
nand g192 ( new_n311_, new_n310_, new_n307_ );
nand g193 ( new_n312_, new_n311_, N183 );
not g194 ( new_n313_, N183 );
nand g195 ( new_n314_, new_n310_, new_n313_, new_n307_ );
nand g196 ( new_n315_, new_n312_, new_n314_ );
not g197 ( new_n316_, new_n315_ );
nand g198 ( new_n317_, new_n306_, new_n316_ );
nand g199 ( new_n318_, new_n305_, new_n302_, new_n315_ );
nand g200 ( new_n319_, new_n317_, N219, new_n318_ );
nand g201 ( new_n320_, new_n316_, N228 );
nand g202 ( new_n321_, new_n311_, N183, N237 );
nand g203 ( new_n322_, new_n311_, N246 );
nand g204 ( new_n323_, N106, N210 );
nand g205 ( new_n324_, new_n254_, N183 );
nand g206 ( new_n325_, new_n321_, new_n322_, new_n323_, new_n324_ );
not g207 ( new_n326_, new_n325_ );
nand g208 ( N863, new_n319_, new_n320_, new_n326_ );
nand g209 ( new_n328_, new_n294_, N195 );
nand g210 ( new_n329_, new_n242_, N261 );
nand g211 ( new_n330_, new_n329_, new_n240_ );
nand g212 ( new_n331_, new_n330_, new_n284_ );
nand g213 ( new_n332_, new_n331_, new_n328_ );
nand g214 ( new_n333_, new_n297_, new_n271_ );
not g215 ( new_n334_, new_n333_ );
nand g216 ( new_n335_, new_n332_, new_n334_ );
nand g217 ( new_n336_, new_n331_, new_n328_, new_n333_ );
nand g218 ( new_n337_, new_n335_, N219, new_n336_ );
nand g219 ( new_n338_, new_n334_, N228 );
nand g220 ( new_n339_, new_n296_, N189, N237 );
nand g221 ( new_n340_, new_n296_, N246 );
nor g222 ( new_n341_, new_n255_, new_n266_ );
nand g223 ( new_n342_, N255, N259 );
nand g224 ( new_n343_, N111, N210 );
nand g225 ( new_n344_, new_n342_, new_n343_ );
nor g226 ( new_n345_, new_n341_, new_n344_ );
nand g227 ( new_n346_, new_n339_, new_n340_, new_n345_ );
not g228 ( new_n347_, new_n346_ );
nand g229 ( new_n348_, new_n337_, new_n338_, new_n347_ );
xnor g230 ( N864, new_n348_, keyIn_0_30 );
nand g231 ( new_n350_, new_n330_, new_n284_, new_n328_ );
nand g232 ( new_n351_, new_n328_, new_n284_ );
nand g233 ( new_n352_, new_n351_, new_n240_, new_n329_ );
nand g234 ( new_n353_, new_n350_, N219, new_n352_ );
nand g235 ( new_n354_, new_n328_, N228, new_n284_ );
nand g236 ( new_n355_, new_n294_, N195, N237 );
nand g237 ( new_n356_, new_n294_, N246 );
nor g238 ( new_n357_, new_n255_, new_n272_ );
nand g239 ( new_n358_, N255, N260 );
nand g240 ( new_n359_, N116, N210 );
nand g241 ( new_n360_, new_n358_, new_n359_ );
nor g242 ( new_n361_, new_n357_, new_n360_ );
nand g243 ( new_n362_, new_n355_, new_n356_, new_n361_ );
not g244 ( new_n363_, new_n362_ );
nand g245 ( new_n364_, new_n353_, new_n354_, new_n363_ );
xor g246 ( N865, new_n364_, keyIn_0_31 );
nand g247 ( new_n366_, new_n306_, new_n314_ );
nand g248 ( new_n367_, new_n366_, new_n312_ );
not g249 ( new_n368_, N171 );
nand g250 ( new_n369_, new_n222_, N101 );
nand g251 ( new_n370_, new_n186_, N55 );
xnor g252 ( new_n371_, new_n370_, keyIn_0_12 );
nand g253 ( new_n372_, new_n371_, N149 );
nand g254 ( new_n373_, new_n182_, keyIn_0_13, N17, new_n230_ );
not g255 ( new_n374_, keyIn_0_13 );
nand g256 ( new_n375_, new_n182_, N17, new_n230_ );
nand g257 ( new_n376_, new_n375_, new_n374_ );
nand g258 ( new_n377_, new_n376_, new_n227_, new_n373_ );
nand g259 ( new_n378_, N17, N138 );
nand g260 ( new_n379_, new_n372_, new_n377_, new_n378_ );
not g261 ( new_n380_, new_n379_ );
nand g262 ( new_n381_, new_n380_, new_n368_, new_n369_ );
not g263 ( new_n382_, N165 );
nand g264 ( new_n383_, new_n222_, N96 );
nand g265 ( new_n384_, new_n371_, N146 );
nand g266 ( new_n385_, N51, N138 );
nand g267 ( new_n386_, new_n384_, new_n377_, new_n385_ );
not g268 ( new_n387_, new_n386_ );
nand g269 ( new_n388_, new_n387_, new_n382_, new_n383_ );
nand g270 ( new_n389_, new_n381_, new_n388_ );
not g271 ( new_n390_, new_n389_ );
not g272 ( new_n391_, N177 );
nand g273 ( new_n392_, new_n222_, N106 );
nand g274 ( new_n393_, new_n371_, N153 );
nand g275 ( new_n394_, N138, N152 );
nand g276 ( new_n395_, new_n393_, new_n377_, new_n394_ );
not g277 ( new_n396_, new_n395_ );
nand g278 ( new_n397_, new_n396_, new_n391_, new_n392_ );
nand g279 ( new_n398_, new_n390_, new_n397_ );
not g280 ( new_n399_, new_n398_ );
nand g281 ( new_n400_, new_n367_, new_n399_ );
nand g282 ( new_n401_, new_n400_, keyIn_0_28 );
not g283 ( new_n402_, keyIn_0_28 );
nand g284 ( new_n403_, new_n367_, new_n402_, new_n399_ );
nand g285 ( new_n404_, new_n387_, new_n383_ );
nand g286 ( new_n405_, new_n404_, N165 );
nand g287 ( new_n406_, new_n396_, new_n392_ );
nand g288 ( new_n407_, new_n406_, N177 );
nand g289 ( new_n408_, new_n380_, new_n369_ );
nand g290 ( new_n409_, new_n408_, N171 );
nand g291 ( new_n410_, new_n407_, new_n409_ );
nand g292 ( new_n411_, new_n390_, new_n410_ );
nand g293 ( new_n412_, new_n411_, new_n405_ );
not g294 ( new_n413_, new_n412_ );
nand g295 ( new_n414_, new_n401_, keyIn_0_29, new_n403_, new_n413_ );
not g296 ( new_n415_, keyIn_0_29 );
nand g297 ( new_n416_, new_n401_, new_n403_, new_n413_ );
nand g298 ( new_n417_, new_n416_, new_n415_ );
nand g299 ( new_n418_, new_n417_, new_n414_ );
not g300 ( new_n419_, N159 );
nand g301 ( new_n420_, new_n222_, N91 );
nand g302 ( new_n421_, new_n371_, N143 );
nand g303 ( new_n422_, N8, N138 );
nand g304 ( new_n423_, new_n421_, new_n377_, new_n422_ );
not g305 ( new_n424_, new_n423_ );
nand g306 ( new_n425_, new_n424_, new_n419_, new_n420_ );
nand g307 ( new_n426_, new_n418_, new_n425_ );
nand g308 ( new_n427_, new_n424_, new_n420_ );
nand g309 ( new_n428_, new_n427_, N159 );
nand g310 ( N866, new_n426_, new_n428_ );
nand g311 ( new_n430_, new_n367_, new_n397_, new_n407_ );
nand g312 ( new_n431_, new_n407_, new_n397_ );
nand g313 ( new_n432_, new_n366_, new_n312_, new_n431_ );
nand g314 ( new_n433_, new_n430_, N219, new_n432_ );
nand g315 ( new_n434_, new_n407_, N228, new_n397_ );
nand g316 ( new_n435_, new_n406_, N177, N237 );
nand g317 ( new_n436_, new_n406_, N246 );
nand g318 ( new_n437_, N101, N210 );
nand g319 ( new_n438_, new_n254_, N177 );
nand g320 ( new_n439_, new_n435_, new_n436_, new_n437_, new_n438_ );
not g321 ( new_n440_, new_n439_ );
nand g322 ( N874, new_n433_, new_n434_, new_n440_ );
nand g323 ( new_n442_, new_n428_, new_n425_ );
not g324 ( new_n443_, new_n442_ );
nand g325 ( new_n444_, new_n418_, new_n443_ );
nand g326 ( new_n445_, new_n417_, new_n414_, new_n442_ );
nand g327 ( new_n446_, new_n444_, N219, new_n445_ );
nand g328 ( new_n447_, new_n443_, N228 );
not g329 ( new_n448_, new_n447_ );
nand g330 ( new_n449_, new_n427_, N159, N237 );
nand g331 ( new_n450_, new_n427_, N246 );
nand g332 ( new_n451_, new_n254_, N159 );
nand g333 ( new_n452_, N210, N268 );
nand g334 ( new_n453_, new_n449_, new_n450_, new_n451_, new_n452_ );
nor g335 ( new_n454_, new_n448_, new_n453_ );
nand g336 ( N878, new_n446_, new_n454_ );
nand g337 ( new_n456_, new_n367_, new_n397_ );
nand g338 ( new_n457_, new_n456_, new_n407_ );
nand g339 ( new_n458_, new_n457_, new_n381_ );
nand g340 ( new_n459_, new_n458_, new_n409_ );
nand g341 ( new_n460_, new_n405_, new_n388_ );
not g342 ( new_n461_, new_n460_ );
nand g343 ( new_n462_, new_n459_, new_n461_ );
nand g344 ( new_n463_, new_n458_, new_n409_, new_n460_ );
nand g345 ( new_n464_, new_n462_, N219, new_n463_ );
nand g346 ( new_n465_, new_n461_, N228 );
nand g347 ( new_n466_, new_n404_, N165, N237 );
nand g348 ( new_n467_, new_n404_, N246 );
nand g349 ( new_n468_, N91, N210 );
nand g350 ( new_n469_, new_n254_, N165 );
nand g351 ( new_n470_, new_n466_, new_n467_, new_n468_, new_n469_ );
not g352 ( new_n471_, new_n470_ );
nand g353 ( N879, new_n464_, new_n465_, new_n471_ );
nand g354 ( new_n473_, new_n457_, new_n381_, new_n409_ );
nand g355 ( new_n474_, new_n409_, new_n381_ );
nand g356 ( new_n475_, new_n456_, new_n407_, new_n474_ );
nand g357 ( new_n476_, new_n473_, N219, new_n475_ );
nand g358 ( new_n477_, new_n409_, N228, new_n381_ );
nand g359 ( new_n478_, new_n408_, N171, N237 );
nand g360 ( new_n479_, new_n408_, N246 );
nand g361 ( new_n480_, N96, N210 );
nand g362 ( new_n481_, new_n254_, N171 );
nand g363 ( new_n482_, new_n478_, new_n479_, new_n480_, new_n481_ );
not g364 ( new_n483_, new_n482_ );
nand g365 ( N880, new_n476_, new_n477_, new_n483_ );
endmodule