module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n1017_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n172_, keyIn_0_28 );
not g001 ( new_n173_, N108 );
not g002 ( new_n174_, N102 );
and g003 ( new_n175_, new_n174_, keyIn_0_16 );
not g004 ( new_n176_, keyIn_0_16 );
and g005 ( new_n177_, new_n176_, N102 );
or g006 ( new_n178_, new_n175_, new_n177_, new_n173_ );
and g007 ( new_n179_, new_n178_, new_n172_ );
not g008 ( new_n180_, new_n175_ );
not g009 ( new_n181_, new_n177_ );
and g010 ( new_n182_, new_n180_, new_n181_, keyIn_0_28, N108 );
or g011 ( new_n183_, new_n179_, new_n182_ );
not g012 ( new_n184_, keyIn_0_26 );
not g013 ( new_n185_, N76 );
and g014 ( new_n186_, new_n185_, keyIn_0_12 );
not g015 ( new_n187_, new_n186_ );
or g016 ( new_n188_, new_n185_, keyIn_0_12 );
and g017 ( new_n189_, new_n187_, new_n188_, new_n184_, N82 );
not g018 ( new_n190_, N82 );
not g019 ( new_n191_, keyIn_0_12 );
and g020 ( new_n192_, new_n191_, N76 );
or g021 ( new_n193_, new_n186_, new_n192_, new_n190_ );
and g022 ( new_n194_, new_n193_, keyIn_0_26 );
or g023 ( new_n195_, new_n194_, new_n189_ );
not g024 ( new_n196_, keyIn_0_27 );
not g025 ( new_n197_, N95 );
or g026 ( new_n198_, keyIn_0_14, N89 );
not g027 ( new_n199_, new_n198_ );
and g028 ( new_n200_, keyIn_0_14, N89 );
or g029 ( new_n201_, new_n199_, new_n197_, new_n200_ );
and g030 ( new_n202_, new_n201_, new_n196_ );
not g031 ( new_n203_, new_n200_ );
and g032 ( new_n204_, new_n203_, keyIn_0_27, N95, new_n198_ );
or g033 ( new_n205_, new_n202_, new_n204_ );
and g034 ( new_n206_, new_n183_, new_n205_, new_n195_ );
not g035 ( new_n207_, N69 );
not g036 ( new_n208_, N63 );
and g037 ( new_n209_, new_n208_, keyIn_0_10 );
not g038 ( new_n210_, keyIn_0_10 );
and g039 ( new_n211_, new_n210_, N63 );
or g040 ( new_n212_, new_n209_, new_n211_, new_n207_ );
and g041 ( new_n213_, new_n212_, keyIn_0_25 );
not g042 ( new_n214_, keyIn_0_25 );
not g043 ( new_n215_, new_n209_ );
not g044 ( new_n216_, new_n211_ );
and g045 ( new_n217_, new_n215_, new_n216_, new_n214_, N69 );
or g046 ( new_n218_, new_n213_, new_n217_ );
not g047 ( new_n219_, N56 );
not g048 ( new_n220_, N50 );
and g049 ( new_n221_, new_n220_, keyIn_0_8 );
not g050 ( new_n222_, keyIn_0_8 );
and g051 ( new_n223_, new_n222_, N50 );
or g052 ( new_n224_, new_n221_, new_n223_, new_n219_ );
and g053 ( new_n225_, new_n224_, keyIn_0_24 );
not g054 ( new_n226_, keyIn_0_24 );
not g055 ( new_n227_, new_n221_ );
not g056 ( new_n228_, new_n223_ );
and g057 ( new_n229_, new_n227_, new_n228_, new_n226_, N56 );
or g058 ( new_n230_, new_n225_, new_n229_ );
and g059 ( new_n231_, new_n218_, new_n230_ );
not g060 ( new_n232_, N4 );
not g061 ( new_n233_, N1 );
and g062 ( new_n234_, new_n233_, keyIn_0_0 );
not g063 ( new_n235_, keyIn_0_0 );
and g064 ( new_n236_, new_n235_, N1 );
or g065 ( new_n237_, new_n234_, new_n236_, new_n232_ );
and g066 ( new_n238_, new_n237_, keyIn_0_18 );
not g067 ( new_n239_, keyIn_0_18 );
not g068 ( new_n240_, new_n234_ );
not g069 ( new_n241_, new_n236_ );
and g070 ( new_n242_, new_n240_, new_n241_, new_n239_, N4 );
or g071 ( new_n243_, new_n238_, new_n242_ );
not g072 ( new_n244_, keyIn_0_21 );
not g073 ( new_n245_, N17 );
not g074 ( new_n246_, N11 );
and g075 ( new_n247_, new_n246_, keyIn_0_2 );
not g076 ( new_n248_, keyIn_0_2 );
and g077 ( new_n249_, new_n248_, N11 );
or g078 ( new_n250_, new_n247_, new_n249_, new_n245_ );
and g079 ( new_n251_, new_n250_, new_n244_ );
not g080 ( new_n252_, new_n247_ );
not g081 ( new_n253_, new_n249_ );
and g082 ( new_n254_, new_n252_, new_n253_, keyIn_0_21, N17 );
or g083 ( new_n255_, new_n251_, new_n254_ );
and g084 ( new_n256_, new_n243_, new_n255_ );
not g085 ( new_n257_, keyIn_0_22 );
not g086 ( new_n258_, N30 );
not g087 ( new_n259_, N24 );
and g088 ( new_n260_, new_n259_, keyIn_0_4 );
not g089 ( new_n261_, keyIn_0_4 );
and g090 ( new_n262_, new_n261_, N24 );
or g091 ( new_n263_, new_n260_, new_n262_, new_n258_ );
and g092 ( new_n264_, new_n263_, new_n257_ );
not g093 ( new_n265_, new_n260_ );
not g094 ( new_n266_, new_n262_ );
and g095 ( new_n267_, new_n265_, new_n266_, keyIn_0_22, N30 );
or g096 ( new_n268_, new_n264_, new_n267_ );
not g097 ( new_n269_, keyIn_0_23 );
or g098 ( new_n270_, keyIn_0_6, N37 );
and g099 ( new_n271_, keyIn_0_6, N37 );
not g100 ( new_n272_, new_n271_ );
and g101 ( new_n273_, new_n272_, new_n270_ );
not g102 ( new_n274_, new_n273_ );
and g103 ( new_n275_, new_n274_, new_n269_, N43 );
not g104 ( new_n276_, N43 );
or g105 ( new_n277_, new_n273_, new_n276_ );
and g106 ( new_n278_, new_n277_, keyIn_0_23 );
or g107 ( new_n279_, new_n278_, new_n275_ );
and g108 ( new_n280_, new_n279_, new_n268_ );
and g109 ( new_n281_, new_n280_, new_n206_, new_n231_, new_n256_ );
or g110 ( new_n282_, new_n281_, keyIn_0_45 );
and g111 ( new_n283_, new_n279_, new_n243_, new_n255_, new_n268_ );
and g112 ( new_n284_, new_n283_, keyIn_0_45, new_n206_, new_n231_ );
not g113 ( new_n285_, new_n284_ );
and g114 ( new_n286_, new_n282_, new_n285_ );
not g115 ( N223, new_n286_ );
not g116 ( new_n288_, keyIn_0_76 );
not g117 ( new_n289_, keyIn_0_64 );
not g118 ( new_n290_, keyIn_0_53 );
not g119 ( new_n291_, new_n218_ );
and g120 ( new_n292_, new_n282_, keyIn_0_46, new_n285_ );
not g121 ( new_n293_, new_n292_ );
or g122 ( new_n294_, new_n286_, keyIn_0_46 );
and g123 ( new_n295_, new_n294_, new_n291_, new_n293_ );
not g124 ( new_n296_, new_n295_ );
and g125 ( new_n297_, new_n294_, new_n293_ );
or g126 ( new_n298_, new_n297_, new_n291_ );
and g127 ( new_n299_, new_n298_, new_n290_, new_n296_ );
not g128 ( new_n300_, new_n299_ );
and g129 ( new_n301_, new_n298_, new_n296_ );
or g130 ( new_n302_, new_n301_, new_n290_ );
and g131 ( new_n303_, new_n302_, new_n300_ );
not g132 ( new_n304_, keyIn_0_37 );
or g133 ( new_n305_, keyIn_0_11, N69 );
not g134 ( new_n306_, new_n305_ );
and g135 ( new_n307_, keyIn_0_11, N69 );
or g136 ( new_n308_, new_n306_, N73, new_n307_ );
not g137 ( new_n309_, new_n308_ );
and g138 ( new_n310_, new_n309_, new_n304_ );
and g139 ( new_n311_, new_n308_, keyIn_0_37 );
or g140 ( new_n312_, new_n310_, new_n311_ );
not g141 ( new_n313_, new_n312_ );
or g142 ( new_n314_, new_n303_, new_n313_ );
and g143 ( new_n315_, new_n314_, new_n289_ );
not g144 ( new_n316_, new_n303_ );
and g145 ( new_n317_, new_n316_, keyIn_0_64, new_n312_ );
or g146 ( new_n318_, new_n315_, new_n317_ );
not g147 ( new_n319_, keyIn_0_63 );
not g148 ( new_n320_, keyIn_0_52 );
not g149 ( new_n321_, new_n230_ );
and g150 ( new_n322_, new_n294_, new_n321_, new_n293_ );
not g151 ( new_n323_, new_n322_ );
or g152 ( new_n324_, new_n297_, new_n321_ );
and g153 ( new_n325_, new_n324_, new_n320_, new_n323_ );
not g154 ( new_n326_, new_n325_ );
and g155 ( new_n327_, new_n324_, new_n323_ );
or g156 ( new_n328_, new_n327_, new_n320_ );
and g157 ( new_n329_, new_n328_, new_n326_ );
not g158 ( new_n330_, keyIn_0_35 );
or g159 ( new_n331_, keyIn_0_9, N56 );
not g160 ( new_n332_, new_n331_ );
and g161 ( new_n333_, keyIn_0_9, N56 );
or g162 ( new_n334_, new_n332_, N60, new_n333_ );
not g163 ( new_n335_, new_n334_ );
and g164 ( new_n336_, new_n335_, new_n330_ );
and g165 ( new_n337_, new_n334_, keyIn_0_35 );
or g166 ( new_n338_, new_n336_, new_n337_ );
not g167 ( new_n339_, new_n338_ );
or g168 ( new_n340_, new_n329_, new_n339_ );
and g169 ( new_n341_, new_n340_, new_n319_ );
not g170 ( new_n342_, new_n329_ );
and g171 ( new_n343_, new_n342_, keyIn_0_63, new_n338_ );
or g172 ( new_n344_, new_n341_, new_n343_ );
not g173 ( new_n345_, keyIn_0_67 );
not g174 ( new_n346_, keyIn_0_56 );
not g175 ( new_n347_, new_n183_ );
and g176 ( new_n348_, new_n294_, new_n347_, new_n293_ );
not g177 ( new_n349_, new_n348_ );
or g178 ( new_n350_, new_n297_, new_n347_ );
and g179 ( new_n351_, new_n350_, new_n346_, new_n349_ );
not g180 ( new_n352_, new_n351_ );
and g181 ( new_n353_, new_n350_, new_n349_ );
or g182 ( new_n354_, new_n353_, new_n346_ );
and g183 ( new_n355_, new_n354_, new_n352_ );
not g184 ( new_n356_, keyIn_0_43 );
or g185 ( new_n357_, keyIn_0_17, N108 );
and g186 ( new_n358_, keyIn_0_17, N108 );
not g187 ( new_n359_, new_n358_ );
and g188 ( new_n360_, new_n359_, new_n357_ );
or g189 ( new_n361_, new_n360_, N112 );
not g190 ( new_n362_, new_n361_ );
and g191 ( new_n363_, new_n362_, new_n356_ );
and g192 ( new_n364_, new_n361_, keyIn_0_43 );
or g193 ( new_n365_, new_n363_, new_n364_ );
not g194 ( new_n366_, new_n365_ );
or g195 ( new_n367_, new_n355_, new_n366_ );
and g196 ( new_n368_, new_n367_, new_n345_ );
not g197 ( new_n369_, new_n355_ );
and g198 ( new_n370_, new_n369_, keyIn_0_67, new_n365_ );
or g199 ( new_n371_, new_n368_, new_n370_ );
and g200 ( new_n372_, new_n318_, new_n344_, new_n371_ );
not g201 ( new_n373_, keyIn_0_60 );
not g202 ( new_n374_, keyIn_0_49 );
and g203 ( new_n375_, new_n294_, new_n255_, new_n293_ );
not g204 ( new_n376_, new_n375_ );
or g205 ( new_n377_, new_n297_, new_n255_ );
and g206 ( new_n378_, new_n377_, new_n374_, new_n376_ );
not g207 ( new_n379_, new_n378_ );
and g208 ( new_n380_, new_n377_, new_n376_ );
or g209 ( new_n381_, new_n380_, new_n374_ );
and g210 ( new_n382_, new_n381_, new_n379_ );
not g211 ( new_n383_, keyIn_0_29 );
or g212 ( new_n384_, keyIn_0_3, N17 );
and g213 ( new_n385_, keyIn_0_3, N17 );
not g214 ( new_n386_, new_n385_ );
and g215 ( new_n387_, new_n386_, new_n384_ );
or g216 ( new_n388_, new_n387_, N21 );
not g217 ( new_n389_, new_n388_ );
and g218 ( new_n390_, new_n389_, new_n383_ );
and g219 ( new_n391_, new_n388_, keyIn_0_29 );
or g220 ( new_n392_, new_n390_, new_n391_ );
not g221 ( new_n393_, new_n392_ );
or g222 ( new_n394_, new_n382_, new_n393_ );
and g223 ( new_n395_, new_n394_, new_n373_ );
not g224 ( new_n396_, new_n382_ );
and g225 ( new_n397_, new_n396_, keyIn_0_60, new_n392_ );
or g226 ( new_n398_, new_n395_, new_n397_ );
not g227 ( new_n399_, keyIn_0_48 );
not g228 ( new_n400_, new_n243_ );
and g229 ( new_n401_, new_n294_, new_n400_, new_n293_ );
not g230 ( new_n402_, new_n401_ );
or g231 ( new_n403_, new_n297_, new_n400_ );
and g232 ( new_n404_, new_n403_, new_n399_, new_n402_ );
not g233 ( new_n405_, new_n404_ );
and g234 ( new_n406_, new_n403_, new_n402_ );
or g235 ( new_n407_, new_n406_, new_n399_ );
and g236 ( new_n408_, new_n407_, new_n405_ );
not g237 ( new_n409_, keyIn_0_19 );
or g238 ( new_n410_, keyIn_0_1, N4 );
not g239 ( new_n411_, new_n410_ );
and g240 ( new_n412_, keyIn_0_1, N4 );
or g241 ( new_n413_, new_n411_, N8, new_n412_ );
not g242 ( new_n414_, new_n413_ );
and g243 ( new_n415_, new_n414_, new_n409_ );
and g244 ( new_n416_, new_n413_, keyIn_0_19 );
or g245 ( new_n417_, new_n415_, new_n416_ );
not g246 ( new_n418_, new_n417_ );
or g247 ( new_n419_, new_n408_, new_n418_ );
and g248 ( new_n420_, new_n419_, keyIn_0_58 );
not g249 ( new_n421_, keyIn_0_58 );
not g250 ( new_n422_, new_n408_ );
and g251 ( new_n423_, new_n422_, new_n421_, new_n417_ );
or g252 ( new_n424_, new_n420_, new_n423_ );
and g253 ( new_n425_, new_n398_, new_n424_ );
not g254 ( new_n426_, keyIn_0_65 );
not g255 ( new_n427_, new_n195_ );
and g256 ( new_n428_, new_n294_, new_n427_, new_n293_ );
not g257 ( new_n429_, new_n428_ );
or g258 ( new_n430_, new_n297_, new_n427_ );
and g259 ( new_n431_, new_n430_, keyIn_0_54, new_n429_ );
not g260 ( new_n432_, new_n431_ );
and g261 ( new_n433_, new_n430_, new_n429_ );
or g262 ( new_n434_, new_n433_, keyIn_0_54 );
and g263 ( new_n435_, new_n434_, new_n432_ );
not g264 ( new_n436_, keyIn_0_39 );
or g265 ( new_n437_, keyIn_0_13, N82 );
not g266 ( new_n438_, new_n437_ );
and g267 ( new_n439_, keyIn_0_13, N82 );
or g268 ( new_n440_, new_n438_, N86, new_n439_ );
not g269 ( new_n441_, new_n440_ );
and g270 ( new_n442_, new_n441_, new_n436_ );
and g271 ( new_n443_, new_n440_, keyIn_0_39 );
or g272 ( new_n444_, new_n442_, new_n443_ );
not g273 ( new_n445_, new_n444_ );
or g274 ( new_n446_, new_n435_, new_n445_ );
and g275 ( new_n447_, new_n446_, new_n426_ );
not g276 ( new_n448_, new_n435_ );
and g277 ( new_n449_, new_n448_, keyIn_0_65, new_n444_ );
or g278 ( new_n450_, new_n447_, new_n449_ );
and g279 ( new_n451_, new_n294_, new_n205_, new_n293_ );
not g280 ( new_n452_, new_n451_ );
or g281 ( new_n453_, new_n297_, new_n205_ );
and g282 ( new_n454_, new_n453_, keyIn_0_55, new_n452_ );
not g283 ( new_n455_, new_n454_ );
and g284 ( new_n456_, new_n453_, new_n452_ );
or g285 ( new_n457_, new_n456_, keyIn_0_55 );
and g286 ( new_n458_, new_n457_, new_n455_ );
not g287 ( new_n459_, keyIn_0_41 );
or g288 ( new_n460_, keyIn_0_15, N95 );
and g289 ( new_n461_, keyIn_0_15, N95 );
not g290 ( new_n462_, new_n461_ );
and g291 ( new_n463_, new_n462_, new_n460_ );
or g292 ( new_n464_, new_n463_, N99 );
not g293 ( new_n465_, new_n464_ );
and g294 ( new_n466_, new_n465_, new_n459_ );
and g295 ( new_n467_, new_n464_, keyIn_0_41 );
or g296 ( new_n468_, new_n466_, new_n467_ );
not g297 ( new_n469_, new_n468_ );
or g298 ( new_n470_, new_n458_, new_n469_ );
and g299 ( new_n471_, new_n470_, keyIn_0_66 );
not g300 ( new_n472_, keyIn_0_66 );
not g301 ( new_n473_, new_n458_ );
and g302 ( new_n474_, new_n473_, new_n472_, new_n468_ );
or g303 ( new_n475_, new_n471_, new_n474_ );
and g304 ( new_n476_, new_n450_, new_n475_ );
not g305 ( new_n477_, keyIn_0_62 );
not g306 ( new_n478_, new_n279_ );
and g307 ( new_n479_, new_n294_, new_n478_, new_n293_ );
not g308 ( new_n480_, new_n479_ );
or g309 ( new_n481_, new_n297_, new_n478_ );
and g310 ( new_n482_, new_n481_, new_n480_ );
or g311 ( new_n483_, new_n482_, keyIn_0_51 );
and g312 ( new_n484_, new_n481_, keyIn_0_51, new_n480_ );
not g313 ( new_n485_, new_n484_ );
and g314 ( new_n486_, new_n483_, new_n485_ );
not g315 ( new_n487_, new_n486_ );
not g316 ( new_n488_, keyIn_0_33 );
or g317 ( new_n489_, keyIn_0_7, N43 );
and g318 ( new_n490_, keyIn_0_7, N43 );
not g319 ( new_n491_, new_n490_ );
and g320 ( new_n492_, new_n491_, new_n489_ );
or g321 ( new_n493_, new_n492_, N47 );
not g322 ( new_n494_, new_n493_ );
and g323 ( new_n495_, new_n494_, new_n488_ );
and g324 ( new_n496_, new_n493_, keyIn_0_33 );
or g325 ( new_n497_, new_n495_, new_n496_ );
and g326 ( new_n498_, new_n487_, new_n477_, new_n497_ );
not g327 ( new_n499_, new_n497_ );
or g328 ( new_n500_, new_n486_, new_n499_ );
and g329 ( new_n501_, new_n500_, keyIn_0_62 );
or g330 ( new_n502_, new_n501_, new_n498_ );
not g331 ( new_n503_, keyIn_0_61 );
not g332 ( new_n504_, keyIn_0_50 );
not g333 ( new_n505_, new_n268_ );
and g334 ( new_n506_, new_n294_, new_n505_, new_n293_ );
not g335 ( new_n507_, new_n506_ );
or g336 ( new_n508_, new_n297_, new_n505_ );
and g337 ( new_n509_, new_n508_, new_n504_, new_n507_ );
not g338 ( new_n510_, new_n509_ );
and g339 ( new_n511_, new_n508_, new_n507_ );
or g340 ( new_n512_, new_n511_, new_n504_ );
and g341 ( new_n513_, new_n512_, new_n510_ );
not g342 ( new_n514_, keyIn_0_31 );
and g343 ( new_n515_, keyIn_0_5, N30 );
or g344 ( new_n516_, keyIn_0_5, N30 );
not g345 ( new_n517_, new_n516_ );
or g346 ( new_n518_, new_n517_, N34, new_n515_ );
and g347 ( new_n519_, new_n518_, new_n514_ );
not g348 ( new_n520_, new_n519_ );
or g349 ( new_n521_, new_n518_, new_n514_ );
and g350 ( new_n522_, new_n520_, new_n521_ );
or g351 ( new_n523_, new_n513_, new_n522_ );
and g352 ( new_n524_, new_n523_, new_n503_ );
not g353 ( new_n525_, new_n513_ );
not g354 ( new_n526_, new_n522_ );
and g355 ( new_n527_, new_n525_, keyIn_0_61, new_n526_ );
or g356 ( new_n528_, new_n524_, new_n527_ );
and g357 ( new_n529_, new_n502_, new_n528_ );
and g358 ( new_n530_, new_n372_, new_n425_, new_n476_, new_n529_ );
or g359 ( new_n531_, new_n530_, new_n288_ );
and g360 ( new_n532_, new_n450_, new_n475_, new_n502_, new_n528_ );
and g361 ( new_n533_, new_n532_, new_n288_, new_n372_, new_n425_ );
not g362 ( new_n534_, new_n533_ );
and g363 ( N329, new_n531_, new_n534_ );
not g364 ( new_n536_, keyIn_0_100 );
not g365 ( new_n537_, keyIn_0_90 );
not g366 ( new_n538_, keyIn_0_86 );
and g367 ( new_n539_, new_n531_, new_n538_, new_n534_ );
not g368 ( new_n540_, new_n539_ );
or g369 ( new_n541_, N329, new_n538_ );
and g370 ( new_n542_, new_n541_, new_n540_ );
or g371 ( new_n543_, new_n542_, new_n528_ );
and g372 ( new_n544_, new_n541_, new_n528_, new_n540_ );
not g373 ( new_n545_, new_n544_ );
and g374 ( new_n546_, new_n543_, new_n545_ );
not g375 ( new_n547_, new_n546_ );
and g376 ( new_n548_, new_n547_, new_n537_ );
not g377 ( new_n549_, new_n548_ );
and g378 ( new_n550_, new_n543_, keyIn_0_90, new_n545_ );
not g379 ( new_n551_, new_n550_ );
not g380 ( new_n552_, keyIn_0_79 );
not g381 ( new_n553_, keyIn_0_69 );
not g382 ( new_n554_, keyIn_0_32 );
or g383 ( new_n555_, new_n517_, N40, new_n515_ );
and g384 ( new_n556_, new_n555_, new_n554_ );
not g385 ( new_n557_, new_n556_ );
or g386 ( new_n558_, new_n555_, new_n554_ );
and g387 ( new_n559_, new_n557_, new_n558_ );
or g388 ( new_n560_, new_n513_, new_n559_ );
and g389 ( new_n561_, new_n560_, new_n553_ );
not g390 ( new_n562_, new_n561_ );
or g391 ( new_n563_, new_n560_, new_n553_ );
and g392 ( new_n564_, new_n562_, new_n563_ );
not g393 ( new_n565_, new_n564_ );
and g394 ( new_n566_, new_n565_, new_n552_ );
and g395 ( new_n567_, new_n564_, keyIn_0_79 );
or g396 ( new_n568_, new_n566_, new_n567_ );
and g397 ( new_n569_, new_n549_, new_n536_, new_n551_, new_n568_ );
not g398 ( new_n570_, new_n568_ );
or g399 ( new_n571_, new_n550_, new_n570_ );
or g400 ( new_n572_, new_n548_, new_n571_ );
and g401 ( new_n573_, new_n572_, keyIn_0_100 );
or g402 ( new_n574_, new_n573_, new_n569_ );
not g403 ( new_n575_, keyIn_0_98 );
or g404 ( new_n576_, new_n542_, new_n424_ );
and g405 ( new_n577_, new_n541_, new_n424_, new_n540_ );
not g406 ( new_n578_, new_n577_ );
and g407 ( new_n579_, new_n576_, new_n578_ );
not g408 ( new_n580_, new_n579_ );
and g409 ( new_n581_, new_n580_, keyIn_0_88 );
not g410 ( new_n582_, new_n581_ );
not g411 ( new_n583_, keyIn_0_88 );
and g412 ( new_n584_, new_n576_, new_n583_, new_n578_ );
not g413 ( new_n585_, new_n584_ );
not g414 ( new_n586_, keyIn_0_77 );
not g415 ( new_n587_, keyIn_0_59 );
not g416 ( new_n588_, keyIn_0_20 );
or g417 ( new_n589_, new_n411_, N14, new_n412_ );
and g418 ( new_n590_, new_n589_, new_n588_ );
not g419 ( new_n591_, new_n590_ );
or g420 ( new_n592_, new_n589_, new_n588_ );
and g421 ( new_n593_, new_n591_, new_n592_ );
or g422 ( new_n594_, new_n408_, new_n593_ );
not g423 ( new_n595_, new_n594_ );
and g424 ( new_n596_, new_n595_, new_n587_ );
and g425 ( new_n597_, new_n594_, keyIn_0_59 );
or g426 ( new_n598_, new_n596_, new_n597_ );
not g427 ( new_n599_, new_n598_ );
and g428 ( new_n600_, new_n599_, new_n586_ );
and g429 ( new_n601_, new_n598_, keyIn_0_77 );
or g430 ( new_n602_, new_n600_, new_n601_ );
and g431 ( new_n603_, new_n582_, new_n575_, new_n585_, new_n602_ );
not g432 ( new_n604_, new_n602_ );
or g433 ( new_n605_, new_n584_, new_n604_ );
or g434 ( new_n606_, new_n581_, new_n605_ );
and g435 ( new_n607_, new_n606_, keyIn_0_98 );
or g436 ( new_n608_, new_n607_, new_n603_ );
not g437 ( new_n609_, keyIn_0_106 );
not g438 ( new_n610_, new_n371_ );
not g439 ( new_n611_, new_n530_ );
and g440 ( new_n612_, new_n611_, keyIn_0_76 );
or g441 ( new_n613_, new_n612_, new_n533_ );
and g442 ( new_n614_, new_n613_, keyIn_0_86 );
or g443 ( new_n615_, new_n614_, new_n539_ );
and g444 ( new_n616_, new_n615_, new_n610_ );
and g445 ( new_n617_, new_n541_, new_n371_, new_n540_ );
or g446 ( new_n618_, new_n616_, new_n617_ );
and g447 ( new_n619_, new_n618_, keyIn_0_97 );
not g448 ( new_n620_, keyIn_0_97 );
or g449 ( new_n621_, new_n542_, new_n371_ );
not g450 ( new_n622_, new_n617_ );
and g451 ( new_n623_, new_n621_, new_n620_, new_n622_ );
not g452 ( new_n624_, keyIn_0_85 );
not g453 ( new_n625_, keyIn_0_75 );
not g454 ( new_n626_, keyIn_0_44 );
or g455 ( new_n627_, new_n360_, N115 );
not g456 ( new_n628_, new_n627_ );
and g457 ( new_n629_, new_n628_, new_n626_ );
and g458 ( new_n630_, new_n627_, keyIn_0_44 );
or g459 ( new_n631_, new_n629_, new_n630_ );
and g460 ( new_n632_, new_n369_, new_n631_ );
not g461 ( new_n633_, new_n632_ );
and g462 ( new_n634_, new_n633_, new_n625_ );
and g463 ( new_n635_, new_n632_, keyIn_0_75 );
or g464 ( new_n636_, new_n634_, new_n635_ );
and g465 ( new_n637_, new_n636_, new_n624_ );
not g466 ( new_n638_, new_n637_ );
or g467 ( new_n639_, new_n636_, new_n624_ );
and g468 ( new_n640_, new_n638_, new_n639_ );
or g469 ( new_n641_, new_n623_, new_n640_ );
or g470 ( new_n642_, new_n619_, new_n641_ );
and g471 ( new_n643_, new_n642_, new_n609_ );
not g472 ( new_n644_, new_n619_ );
not g473 ( new_n645_, new_n623_ );
not g474 ( new_n646_, new_n640_ );
and g475 ( new_n647_, new_n644_, keyIn_0_106, new_n645_, new_n646_ );
or g476 ( new_n648_, new_n643_, new_n647_ );
and g477 ( new_n649_, new_n574_, new_n608_, new_n648_ );
not g478 ( new_n650_, keyIn_0_102 );
not g479 ( new_n651_, new_n344_ );
and g480 ( new_n652_, new_n542_, new_n651_ );
not g481 ( new_n653_, new_n652_ );
or g482 ( new_n654_, new_n542_, new_n651_ );
and g483 ( new_n655_, new_n653_, new_n654_ );
and g484 ( new_n656_, new_n655_, keyIn_0_92 );
not g485 ( new_n657_, new_n656_ );
or g486 ( new_n658_, new_n655_, keyIn_0_92 );
not g487 ( new_n659_, keyIn_0_71 );
not g488 ( new_n660_, keyIn_0_36 );
or g489 ( new_n661_, new_n332_, N66, new_n333_ );
not g490 ( new_n662_, new_n661_ );
and g491 ( new_n663_, new_n662_, new_n660_ );
and g492 ( new_n664_, new_n661_, keyIn_0_36 );
or g493 ( new_n665_, new_n663_, new_n664_ );
and g494 ( new_n666_, new_n342_, new_n665_ );
not g495 ( new_n667_, new_n666_ );
and g496 ( new_n668_, new_n667_, new_n659_ );
and g497 ( new_n669_, new_n666_, keyIn_0_71 );
or g498 ( new_n670_, new_n668_, new_n669_ );
or g499 ( new_n671_, new_n670_, keyIn_0_81 );
not g500 ( new_n672_, keyIn_0_81 );
not g501 ( new_n673_, new_n670_ );
or g502 ( new_n674_, new_n673_, new_n672_ );
and g503 ( new_n675_, new_n657_, new_n658_, new_n671_, new_n674_ );
or g504 ( new_n676_, new_n675_, new_n650_ );
not g505 ( new_n677_, keyIn_0_91 );
not g506 ( new_n678_, new_n502_ );
and g507 ( new_n679_, new_n541_, new_n678_, new_n540_ );
not g508 ( new_n680_, new_n679_ );
or g509 ( new_n681_, new_n542_, new_n678_ );
and g510 ( new_n682_, new_n681_, new_n680_ );
or g511 ( new_n683_, new_n682_, new_n677_ );
not g512 ( new_n684_, new_n683_ );
and g513 ( new_n685_, new_n681_, new_n677_, new_n680_ );
not g514 ( new_n686_, keyIn_0_80 );
not g515 ( new_n687_, keyIn_0_70 );
not g516 ( new_n688_, keyIn_0_34 );
or g517 ( new_n689_, new_n492_, N53 );
not g518 ( new_n690_, new_n689_ );
and g519 ( new_n691_, new_n690_, new_n688_ );
and g520 ( new_n692_, new_n689_, keyIn_0_34 );
or g521 ( new_n693_, new_n691_, new_n692_ );
and g522 ( new_n694_, new_n487_, new_n693_ );
not g523 ( new_n695_, new_n694_ );
and g524 ( new_n696_, new_n695_, new_n687_ );
and g525 ( new_n697_, new_n694_, keyIn_0_70 );
or g526 ( new_n698_, new_n696_, new_n697_ );
and g527 ( new_n699_, new_n698_, new_n686_ );
or g528 ( new_n700_, new_n698_, new_n686_ );
not g529 ( new_n701_, new_n700_ );
or g530 ( new_n702_, new_n685_, new_n699_, new_n701_ );
or g531 ( new_n703_, new_n684_, new_n702_, keyIn_0_101 );
and g532 ( new_n704_, new_n675_, new_n650_ );
not g533 ( new_n705_, new_n704_ );
and g534 ( new_n706_, new_n705_, new_n676_, new_n703_ );
not g535 ( new_n707_, keyIn_0_99 );
not g536 ( new_n708_, keyIn_0_89 );
not g537 ( new_n709_, new_n398_ );
and g538 ( new_n710_, new_n541_, new_n709_, new_n540_ );
not g539 ( new_n711_, new_n710_ );
or g540 ( new_n712_, new_n542_, new_n709_ );
and g541 ( new_n713_, new_n712_, new_n711_ );
or g542 ( new_n714_, new_n713_, new_n708_ );
and g543 ( new_n715_, new_n712_, new_n708_, new_n711_ );
not g544 ( new_n716_, new_n715_ );
not g545 ( new_n717_, keyIn_0_78 );
not g546 ( new_n718_, keyIn_0_68 );
not g547 ( new_n719_, keyIn_0_30 );
or g548 ( new_n720_, new_n387_, N27 );
and g549 ( new_n721_, new_n720_, new_n719_ );
not g550 ( new_n722_, new_n721_ );
or g551 ( new_n723_, new_n720_, new_n719_ );
and g552 ( new_n724_, new_n722_, new_n723_ );
or g553 ( new_n725_, new_n382_, new_n724_ );
not g554 ( new_n726_, new_n725_ );
and g555 ( new_n727_, new_n726_, new_n718_ );
and g556 ( new_n728_, new_n725_, keyIn_0_68 );
or g557 ( new_n729_, new_n727_, new_n728_ );
and g558 ( new_n730_, new_n729_, new_n717_ );
not g559 ( new_n731_, new_n730_ );
or g560 ( new_n732_, new_n729_, new_n717_ );
and g561 ( new_n733_, new_n731_, new_n732_ );
and g562 ( new_n734_, new_n714_, new_n716_, new_n733_ );
or g563 ( new_n735_, new_n734_, new_n707_ );
not g564 ( new_n736_, keyIn_0_105 );
not g565 ( new_n737_, new_n475_ );
and g566 ( new_n738_, new_n541_, new_n737_, new_n540_ );
not g567 ( new_n739_, new_n738_ );
or g568 ( new_n740_, new_n542_, new_n737_ );
and g569 ( new_n741_, new_n740_, new_n739_ );
or g570 ( new_n742_, new_n741_, keyIn_0_96 );
and g571 ( new_n743_, new_n740_, keyIn_0_96, new_n739_ );
not g572 ( new_n744_, new_n743_ );
not g573 ( new_n745_, keyIn_0_84 );
not g574 ( new_n746_, keyIn_0_74 );
not g575 ( new_n747_, keyIn_0_42 );
or g576 ( new_n748_, new_n463_, N105 );
and g577 ( new_n749_, new_n748_, new_n747_ );
not g578 ( new_n750_, new_n749_ );
or g579 ( new_n751_, new_n748_, new_n747_ );
and g580 ( new_n752_, new_n750_, new_n751_ );
or g581 ( new_n753_, new_n458_, new_n752_ );
and g582 ( new_n754_, new_n753_, new_n746_ );
not g583 ( new_n755_, new_n754_ );
or g584 ( new_n756_, new_n753_, new_n746_ );
and g585 ( new_n757_, new_n755_, new_n756_ );
and g586 ( new_n758_, new_n757_, new_n745_ );
not g587 ( new_n759_, new_n758_ );
or g588 ( new_n760_, new_n757_, new_n745_ );
and g589 ( new_n761_, new_n759_, new_n760_ );
and g590 ( new_n762_, new_n742_, new_n744_, new_n761_ );
or g591 ( new_n763_, new_n762_, new_n736_ );
and g592 ( new_n764_, new_n735_, new_n763_ );
not g593 ( new_n765_, keyIn_0_101 );
not g594 ( new_n766_, new_n685_ );
not g595 ( new_n767_, new_n699_ );
and g596 ( new_n768_, new_n767_, new_n700_ );
and g597 ( new_n769_, new_n683_, new_n766_, new_n768_ );
or g598 ( new_n770_, new_n769_, new_n765_ );
not g599 ( new_n771_, new_n714_ );
not g600 ( new_n772_, new_n732_ );
or g601 ( new_n773_, new_n715_, new_n730_, new_n772_ );
or g602 ( new_n774_, new_n771_, new_n773_, keyIn_0_99 );
and g603 ( new_n775_, new_n770_, new_n774_ );
or g604 ( new_n776_, new_n542_, new_n318_ );
and g605 ( new_n777_, new_n541_, new_n318_, new_n540_ );
not g606 ( new_n778_, new_n777_ );
and g607 ( new_n779_, new_n776_, new_n778_ );
or g608 ( new_n780_, new_n779_, keyIn_0_93 );
and g609 ( new_n781_, new_n776_, keyIn_0_93, new_n778_ );
not g610 ( new_n782_, new_n781_ );
not g611 ( new_n783_, keyIn_0_82 );
not g612 ( new_n784_, keyIn_0_72 );
not g613 ( new_n785_, keyIn_0_38 );
or g614 ( new_n786_, new_n306_, N79, new_n307_ );
not g615 ( new_n787_, new_n786_ );
and g616 ( new_n788_, new_n787_, new_n785_ );
and g617 ( new_n789_, new_n786_, keyIn_0_38 );
or g618 ( new_n790_, new_n788_, new_n789_ );
and g619 ( new_n791_, new_n316_, new_n790_ );
not g620 ( new_n792_, new_n791_ );
and g621 ( new_n793_, new_n792_, new_n784_ );
and g622 ( new_n794_, new_n791_, keyIn_0_72 );
or g623 ( new_n795_, new_n793_, new_n794_ );
not g624 ( new_n796_, new_n795_ );
and g625 ( new_n797_, new_n796_, new_n783_ );
not g626 ( new_n798_, new_n797_ );
and g627 ( new_n799_, new_n795_, keyIn_0_82 );
not g628 ( new_n800_, new_n799_ );
and g629 ( new_n801_, new_n798_, new_n800_ );
and g630 ( new_n802_, new_n780_, new_n782_, new_n801_ );
or g631 ( new_n803_, new_n802_, keyIn_0_103 );
not g632 ( new_n804_, keyIn_0_104 );
not g633 ( new_n805_, keyIn_0_94 );
not g634 ( new_n806_, new_n450_ );
and g635 ( new_n807_, new_n541_, new_n806_, new_n540_ );
not g636 ( new_n808_, new_n807_ );
or g637 ( new_n809_, new_n542_, new_n806_ );
and g638 ( new_n810_, new_n809_, new_n805_, new_n808_ );
not g639 ( new_n811_, keyIn_0_83 );
not g640 ( new_n812_, keyIn_0_73 );
not g641 ( new_n813_, keyIn_0_40 );
or g642 ( new_n814_, new_n438_, N92, new_n439_ );
not g643 ( new_n815_, new_n814_ );
and g644 ( new_n816_, new_n815_, new_n813_ );
and g645 ( new_n817_, new_n814_, keyIn_0_40 );
or g646 ( new_n818_, new_n816_, new_n817_ );
and g647 ( new_n819_, new_n448_, new_n818_ );
not g648 ( new_n820_, new_n819_ );
and g649 ( new_n821_, new_n820_, new_n812_ );
and g650 ( new_n822_, new_n819_, keyIn_0_73 );
or g651 ( new_n823_, new_n821_, new_n822_ );
not g652 ( new_n824_, new_n823_ );
and g653 ( new_n825_, new_n824_, new_n811_ );
and g654 ( new_n826_, new_n823_, keyIn_0_83 );
or g655 ( new_n827_, new_n810_, new_n825_, new_n826_ );
and g656 ( new_n828_, new_n809_, new_n808_ );
or g657 ( new_n829_, new_n828_, new_n805_ );
not g658 ( new_n830_, new_n829_ );
or g659 ( new_n831_, new_n830_, new_n827_, new_n804_ );
not g660 ( new_n832_, new_n742_ );
not g661 ( new_n833_, new_n760_ );
or g662 ( new_n834_, new_n743_, new_n758_, new_n833_ );
or g663 ( new_n835_, new_n832_, new_n834_, keyIn_0_105 );
and g664 ( new_n836_, new_n803_, new_n831_, new_n835_ );
not g665 ( new_n837_, keyIn_0_103 );
not g666 ( new_n838_, new_n780_ );
or g667 ( new_n839_, new_n781_, new_n797_, new_n799_ );
or g668 ( new_n840_, new_n838_, new_n839_, new_n837_ );
not g669 ( new_n841_, new_n810_ );
not g670 ( new_n842_, new_n825_ );
not g671 ( new_n843_, new_n826_ );
and g672 ( new_n844_, new_n842_, new_n843_ );
and g673 ( new_n845_, new_n829_, new_n841_, new_n844_ );
or g674 ( new_n846_, new_n845_, keyIn_0_104 );
and g675 ( new_n847_, new_n846_, new_n840_ );
and g676 ( new_n848_, new_n836_, new_n764_, new_n775_, new_n847_ );
and g677 ( new_n849_, new_n649_, new_n848_, new_n706_ );
or g678 ( new_n850_, new_n849_, keyIn_0_107 );
and g679 ( new_n851_, new_n649_, new_n848_, new_n706_, keyIn_0_107 );
not g680 ( new_n852_, new_n851_ );
and g681 ( new_n853_, new_n850_, new_n852_ );
not g682 ( N370, new_n853_ );
not g683 ( new_n855_, keyIn_0_120 );
not g684 ( new_n856_, keyIn_0_119 );
not g685 ( new_n857_, keyIn_0_108 );
and g686 ( new_n858_, new_n850_, new_n857_, new_n852_ );
not g687 ( new_n859_, new_n858_ );
or g688 ( new_n860_, new_n853_, new_n857_ );
and g689 ( new_n861_, new_n860_, N53, new_n859_ );
or g690 ( new_n862_, new_n861_, keyIn_0_109 );
and g691 ( new_n863_, new_n860_, keyIn_0_109, N53, new_n859_ );
not g692 ( new_n864_, new_n863_ );
not g693 ( new_n865_, keyIn_0_95 );
not g694 ( new_n866_, keyIn_0_87 );
and g695 ( new_n867_, N329, new_n866_ );
not g696 ( new_n868_, new_n867_ );
or g697 ( new_n869_, N329, new_n866_ );
and g698 ( new_n870_, new_n868_, new_n869_ );
and g699 ( new_n871_, new_n870_, N47 );
or g700 ( new_n872_, new_n871_, new_n865_ );
not g701 ( new_n873_, new_n872_ );
and g702 ( new_n874_, new_n871_, new_n865_ );
not g703 ( new_n875_, keyIn_0_57 );
or g704 ( new_n876_, new_n286_, keyIn_0_47 );
and g705 ( new_n877_, new_n286_, keyIn_0_47 );
not g706 ( new_n878_, new_n877_ );
and g707 ( new_n879_, new_n878_, new_n876_ );
not g708 ( new_n880_, new_n879_ );
and g709 ( new_n881_, new_n880_, N37 );
and g710 ( new_n882_, new_n881_, new_n875_ );
not g711 ( new_n883_, new_n882_ );
or g712 ( new_n884_, new_n881_, new_n875_ );
and g713 ( new_n885_, new_n883_, new_n884_ );
or g714 ( new_n886_, new_n873_, new_n874_, new_n276_, new_n885_ );
not g715 ( new_n887_, new_n886_ );
and g716 ( new_n888_, new_n862_, new_n864_, new_n887_ );
or g717 ( new_n889_, new_n888_, keyIn_0_113 );
not g718 ( new_n890_, keyIn_0_113 );
not g719 ( new_n891_, keyIn_0_109 );
not g720 ( new_n892_, new_n861_ );
and g721 ( new_n893_, new_n892_, new_n891_ );
or g722 ( new_n894_, new_n863_, new_n886_ );
or g723 ( new_n895_, new_n893_, new_n894_, new_n890_ );
and g724 ( new_n896_, new_n889_, new_n895_ );
not g725 ( new_n897_, keyIn_0_114 );
and g726 ( new_n898_, new_n860_, N66, new_n859_ );
and g727 ( new_n899_, new_n870_, N60 );
and g728 ( new_n900_, new_n880_, N50 );
or g729 ( new_n901_, new_n899_, new_n219_, new_n900_ );
or g730 ( new_n902_, new_n898_, new_n901_ );
not g731 ( new_n903_, new_n902_ );
and g732 ( new_n904_, new_n903_, new_n897_ );
and g733 ( new_n905_, new_n902_, keyIn_0_114 );
or g734 ( new_n906_, new_n904_, new_n905_ );
not g735 ( new_n907_, new_n906_ );
or g736 ( new_n908_, new_n896_, new_n907_ );
not g737 ( new_n909_, keyIn_0_111 );
and g738 ( new_n910_, new_n860_, new_n859_ );
and g739 ( new_n911_, new_n910_, N27 );
not g740 ( new_n912_, new_n911_ );
and g741 ( new_n913_, new_n870_, N21 );
and g742 ( new_n914_, new_n880_, N11 );
or g743 ( new_n915_, new_n913_, new_n245_, new_n914_ );
not g744 ( new_n916_, new_n915_ );
and g745 ( new_n917_, new_n912_, new_n909_, new_n916_ );
or g746 ( new_n918_, new_n911_, new_n915_ );
and g747 ( new_n919_, new_n918_, keyIn_0_111 );
or g748 ( new_n920_, new_n919_, new_n917_ );
not g749 ( new_n921_, keyIn_0_112 );
and g750 ( new_n922_, new_n860_, N40, new_n859_ );
and g751 ( new_n923_, new_n870_, N34 );
and g752 ( new_n924_, new_n880_, N24 );
or g753 ( new_n925_, new_n923_, new_n258_, new_n924_ );
or g754 ( new_n926_, new_n922_, new_n925_ );
and g755 ( new_n927_, new_n926_, new_n921_ );
not g756 ( new_n928_, new_n922_ );
not g757 ( new_n929_, new_n925_ );
and g758 ( new_n930_, new_n928_, keyIn_0_112, new_n929_ );
or g759 ( new_n931_, new_n927_, new_n930_ );
and g760 ( new_n932_, new_n920_, new_n931_ );
not g761 ( new_n933_, new_n932_ );
not g762 ( new_n934_, keyIn_0_117 );
and g763 ( new_n935_, new_n860_, N105, new_n859_ );
and g764 ( new_n936_, new_n870_, N99 );
and g765 ( new_n937_, new_n880_, N89 );
or g766 ( new_n938_, new_n936_, new_n197_, new_n937_ );
or g767 ( new_n939_, new_n935_, new_n938_ );
and g768 ( new_n940_, new_n939_, new_n934_ );
or g769 ( new_n941_, new_n939_, new_n934_ );
not g770 ( new_n942_, new_n941_ );
or g771 ( new_n943_, new_n942_, new_n940_ );
not g772 ( new_n944_, keyIn_0_118 );
and g773 ( new_n945_, new_n860_, N115, new_n859_ );
and g774 ( new_n946_, new_n870_, N112 );
and g775 ( new_n947_, new_n880_, N102 );
or g776 ( new_n948_, new_n945_, new_n173_, new_n946_, new_n947_ );
and g777 ( new_n949_, new_n948_, new_n944_ );
not g778 ( new_n950_, new_n945_ );
not g779 ( new_n951_, new_n946_ );
not g780 ( new_n952_, new_n947_ );
and g781 ( new_n953_, new_n951_, N108, new_n952_ );
and g782 ( new_n954_, new_n950_, keyIn_0_118, new_n953_ );
or g783 ( new_n955_, new_n949_, new_n954_ );
not g784 ( new_n956_, keyIn_0_115 );
and g785 ( new_n957_, new_n860_, N79, new_n859_ );
and g786 ( new_n958_, new_n870_, N73 );
and g787 ( new_n959_, new_n880_, N63 );
or g788 ( new_n960_, new_n958_, new_n207_, new_n959_ );
or g789 ( new_n961_, new_n957_, new_n960_ );
and g790 ( new_n962_, new_n961_, new_n956_ );
or g791 ( new_n963_, new_n961_, new_n956_ );
not g792 ( new_n964_, new_n963_ );
or g793 ( new_n965_, new_n964_, new_n962_ );
not g794 ( new_n966_, keyIn_0_116 );
and g795 ( new_n967_, new_n860_, N92, new_n859_ );
and g796 ( new_n968_, new_n870_, N86 );
and g797 ( new_n969_, new_n880_, N76 );
or g798 ( new_n970_, new_n968_, new_n190_, new_n969_ );
or g799 ( new_n971_, new_n967_, new_n970_ );
and g800 ( new_n972_, new_n971_, new_n966_ );
not g801 ( new_n973_, new_n967_ );
not g802 ( new_n974_, new_n970_ );
and g803 ( new_n975_, new_n973_, keyIn_0_116, new_n974_ );
or g804 ( new_n976_, new_n972_, new_n975_ );
and g805 ( new_n977_, new_n943_, new_n965_, new_n955_, new_n976_ );
not g806 ( new_n978_, new_n977_ );
or g807 ( new_n979_, new_n978_, new_n933_, new_n908_, new_n856_ );
or g808 ( new_n980_, new_n893_, new_n894_ );
and g809 ( new_n981_, new_n980_, new_n890_ );
not g810 ( new_n982_, new_n895_ );
or g811 ( new_n983_, new_n981_, new_n982_ );
and g812 ( new_n984_, new_n977_, new_n932_, new_n983_, new_n906_ );
or g813 ( new_n985_, new_n984_, keyIn_0_119 );
not g814 ( new_n986_, keyIn_0_110 );
and g815 ( new_n987_, new_n910_, N14 );
and g816 ( new_n988_, new_n870_, N8 );
and g817 ( new_n989_, new_n880_, N1 );
or g818 ( new_n990_, new_n987_, new_n232_, new_n988_, new_n989_ );
and g819 ( new_n991_, new_n990_, new_n986_ );
not g820 ( new_n992_, new_n990_ );
and g821 ( new_n993_, new_n992_, keyIn_0_110 );
or g822 ( new_n994_, new_n993_, new_n991_ );
and g823 ( new_n995_, new_n985_, new_n979_, new_n994_ );
not g824 ( new_n996_, new_n995_ );
and g825 ( new_n997_, new_n996_, new_n855_ );
and g826 ( new_n998_, new_n995_, keyIn_0_120 );
or g827 ( N421, new_n997_, new_n998_ );
not g828 ( new_n1000_, keyIn_0_125 );
and g829 ( new_n1001_, new_n889_, new_n895_, new_n931_ );
or g830 ( new_n1002_, new_n1001_, keyIn_0_121 );
and g831 ( new_n1003_, new_n889_, new_n931_, keyIn_0_121, new_n895_ );
not g832 ( new_n1004_, new_n1003_ );
and g833 ( new_n1005_, new_n1002_, new_n1004_ );
or g834 ( new_n1006_, new_n1005_, new_n907_, new_n933_ );
and g835 ( new_n1007_, new_n1006_, new_n1000_ );
not g836 ( new_n1008_, new_n1005_ );
and g837 ( new_n1009_, new_n1008_, keyIn_0_125, new_n906_, new_n932_ );
or g838 ( N430, new_n1007_, new_n1009_ );
not g839 ( new_n1011_, keyIn_0_126 );
not g840 ( new_n1012_, new_n962_ );
and g841 ( new_n1013_, new_n906_, new_n1012_, new_n963_ );
and g842 ( new_n1014_, new_n1013_, new_n983_, new_n931_ );
or g843 ( new_n1015_, new_n1014_, keyIn_0_122 );
not g844 ( new_n1016_, keyIn_0_122 );
not g845 ( new_n1017_, new_n931_ );
or g846 ( new_n1018_, new_n896_, new_n1017_ );
not g847 ( new_n1019_, new_n1013_ );
or g848 ( new_n1020_, new_n1018_, new_n1019_, new_n1016_ );
and g849 ( new_n1021_, new_n1015_, new_n1020_ );
not g850 ( new_n1022_, keyIn_0_123 );
not g851 ( new_n1023_, new_n976_ );
and g852 ( new_n1024_, new_n983_, new_n906_, new_n1023_ );
or g853 ( new_n1025_, new_n1024_, new_n1022_ );
or g854 ( new_n1026_, new_n908_, keyIn_0_123, new_n976_ );
and g855 ( new_n1027_, new_n1025_, new_n1026_ );
or g856 ( new_n1028_, new_n1021_, new_n1027_, new_n933_ );
and g857 ( new_n1029_, new_n1028_, new_n1011_ );
not g858 ( new_n1030_, new_n1021_ );
not g859 ( new_n1031_, new_n1027_ );
and g860 ( new_n1032_, new_n1030_, new_n1031_, keyIn_0_126, new_n932_ );
or g861 ( N431, new_n1029_, new_n1032_ );
not g862 ( new_n1034_, new_n940_ );
and g863 ( new_n1035_, new_n976_, new_n1034_, new_n941_ );
not g864 ( new_n1036_, new_n1035_ );
or g865 ( new_n1037_, new_n1018_, keyIn_0_124, new_n1036_ );
not g866 ( new_n1038_, keyIn_0_124 );
and g867 ( new_n1039_, new_n983_, new_n931_, new_n1035_ );
or g868 ( new_n1040_, new_n1039_, new_n1038_ );
and g869 ( new_n1041_, new_n1040_, new_n1037_ );
not g870 ( new_n1042_, new_n920_ );
or g871 ( new_n1043_, new_n1005_, new_n1042_ );
or g872 ( new_n1044_, new_n1021_, new_n1041_, new_n1043_ );
and g873 ( new_n1045_, new_n1044_, keyIn_0_127 );
not g874 ( new_n1046_, keyIn_0_127 );
not g875 ( new_n1047_, new_n1041_ );
not g876 ( new_n1048_, new_n1043_ );
and g877 ( new_n1049_, new_n1030_, new_n1047_, new_n1046_, new_n1048_ );
or g878 ( N432, new_n1045_, new_n1049_ );
endmodule