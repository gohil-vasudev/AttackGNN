module add_mul_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, 
        b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, 
        b_15_, operation, Result_0_, Result_1_, Result_2_, Result_3_, 
        Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, 
        Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, 
        Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, 
        Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, 
        Result_28_, Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013;

  NOR2_X2 U1943 ( .A1(n2208), .A2(a_14_), .ZN(n2380) );
  NOR2_X2 U1944 ( .A1(n2499), .A2(a_15_), .ZN(n2383) );
  INV_X2 U1945 ( .A(operation), .ZN(n1911) );
  NOR2_X1 U1946 ( .A1(n1911), .A2(n1912), .ZN(Result_9_) );
  XOR2_X1 U1947 ( .A(n1913), .B(n1914), .Z(n1912) );
  NAND2_X1 U1948 ( .A1(n1915), .A2(n1916), .ZN(n1914) );
  NOR2_X1 U1949 ( .A1(n1911), .A2(n1917), .ZN(Result_8_) );
  XOR2_X1 U1950 ( .A(n1918), .B(n1919), .Z(n1917) );
  NAND2_X1 U1951 ( .A1(n1920), .A2(n1921), .ZN(n1919) );
  NOR2_X1 U1952 ( .A1(n1911), .A2(n1922), .ZN(Result_7_) );
  XOR2_X1 U1953 ( .A(n1923), .B(n1924), .Z(n1922) );
  NAND2_X1 U1954 ( .A1(n1925), .A2(n1926), .ZN(n1924) );
  NOR2_X1 U1955 ( .A1(n1911), .A2(n1927), .ZN(Result_6_) );
  XOR2_X1 U1956 ( .A(n1928), .B(n1929), .Z(n1927) );
  NAND2_X1 U1957 ( .A1(n1930), .A2(n1931), .ZN(n1929) );
  NOR2_X1 U1958 ( .A1(n1911), .A2(n1932), .ZN(Result_5_) );
  XOR2_X1 U1959 ( .A(n1933), .B(n1934), .Z(n1932) );
  NAND2_X1 U1960 ( .A1(n1935), .A2(n1936), .ZN(n1934) );
  NOR2_X1 U1961 ( .A1(n1911), .A2(n1937), .ZN(Result_4_) );
  XOR2_X1 U1962 ( .A(n1938), .B(n1939), .Z(n1937) );
  NAND2_X1 U1963 ( .A1(n1940), .A2(n1941), .ZN(n1939) );
  NOR2_X1 U1964 ( .A1(n1911), .A2(n1942), .ZN(Result_3_) );
  XOR2_X1 U1965 ( .A(n1943), .B(n1944), .Z(n1942) );
  NAND2_X1 U1966 ( .A1(n1945), .A2(n1946), .ZN(n1944) );
  NAND2_X1 U1967 ( .A1(n1947), .A2(n1948), .ZN(Result_31_) );
  NAND2_X1 U1968 ( .A1(n1949), .A2(n1911), .ZN(n1948) );
  XNOR2_X1 U1969 ( .A(n1950), .B(a_15_), .ZN(n1949) );
  NAND2_X1 U1970 ( .A1(n1951), .A2(operation), .ZN(n1947) );
  NAND2_X1 U1971 ( .A1(n1952), .A2(n1953), .ZN(Result_30_) );
  NAND2_X1 U1972 ( .A1(operation), .A2(n1954), .ZN(n1953) );
  NAND2_X1 U1973 ( .A1(n1955), .A2(n1956), .ZN(n1954) );
  NAND2_X1 U1974 ( .A1(b_14_), .A2(n1957), .ZN(n1956) );
  NAND2_X1 U1975 ( .A1(n1958), .A2(n1959), .ZN(n1957) );
  NAND2_X1 U1976 ( .A1(a_15_), .A2(n1950), .ZN(n1959) );
  NAND2_X1 U1977 ( .A1(b_15_), .A2(n1960), .ZN(n1955) );
  NAND2_X1 U1978 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
  NAND2_X1 U1979 ( .A1(a_14_), .A2(n1963), .ZN(n1962) );
  NAND2_X1 U1980 ( .A1(n1964), .A2(n1911), .ZN(n1952) );
  XNOR2_X1 U1981 ( .A(n1951), .B(n1965), .ZN(n1964) );
  XNOR2_X1 U1982 ( .A(a_14_), .B(b_14_), .ZN(n1965) );
  NOR2_X1 U1983 ( .A1(n1911), .A2(n1966), .ZN(Result_2_) );
  XOR2_X1 U1984 ( .A(n1967), .B(n1968), .Z(n1966) );
  NAND2_X1 U1985 ( .A1(n1969), .A2(n1970), .ZN(n1968) );
  NAND2_X1 U1986 ( .A1(n1971), .A2(n1972), .ZN(Result_29_) );
  NAND2_X1 U1987 ( .A1(n1973), .A2(n1911), .ZN(n1972) );
  NAND2_X1 U1988 ( .A1(n1974), .A2(n1975), .ZN(n1973) );
  NAND2_X1 U1989 ( .A1(n1976), .A2(n1977), .ZN(n1975) );
  NOR2_X1 U1990 ( .A1(n1978), .A2(n1979), .ZN(n1974) );
  NOR2_X1 U1991 ( .A1(b_13_), .A2(n1980), .ZN(n1979) );
  XNOR2_X1 U1992 ( .A(a_13_), .B(n1977), .ZN(n1980) );
  NOR2_X1 U1993 ( .A1(n1981), .A2(n1982), .ZN(n1978) );
  OR2_X1 U1994 ( .A1(n1977), .A2(a_13_), .ZN(n1982) );
  NAND2_X1 U1995 ( .A1(n1983), .A2(operation), .ZN(n1971) );
  XOR2_X1 U1996 ( .A(n1984), .B(n1985), .Z(n1983) );
  XNOR2_X1 U1997 ( .A(n1986), .B(n1987), .ZN(n1985) );
  NAND2_X1 U1998 ( .A1(b_15_), .A2(a_13_), .ZN(n1984) );
  NAND2_X1 U1999 ( .A1(n1988), .A2(n1989), .ZN(Result_28_) );
  NAND2_X1 U2000 ( .A1(n1990), .A2(n1911), .ZN(n1989) );
  XOR2_X1 U2001 ( .A(n1991), .B(n1992), .Z(n1990) );
  AND2_X1 U2002 ( .A1(n1993), .A2(n1994), .ZN(n1992) );
  NAND2_X1 U2003 ( .A1(n1995), .A2(operation), .ZN(n1988) );
  XNOR2_X1 U2004 ( .A(n1996), .B(n1997), .ZN(n1995) );
  XNOR2_X1 U2005 ( .A(n1998), .B(n1999), .ZN(n1997) );
  NOR2_X1 U2006 ( .A1(n2000), .A2(n1950), .ZN(n1999) );
  NAND2_X1 U2007 ( .A1(n2001), .A2(n2002), .ZN(Result_27_) );
  NAND2_X1 U2008 ( .A1(n2003), .A2(n1911), .ZN(n2002) );
  NAND2_X1 U2009 ( .A1(n2004), .A2(n2005), .ZN(n2003) );
  NAND2_X1 U2010 ( .A1(n2006), .A2(n2007), .ZN(n2005) );
  NOR2_X1 U2011 ( .A1(n2008), .A2(n2009), .ZN(n2004) );
  NOR2_X1 U2012 ( .A1(b_11_), .A2(n2010), .ZN(n2009) );
  XNOR2_X1 U2013 ( .A(a_11_), .B(n2007), .ZN(n2010) );
  NOR2_X1 U2014 ( .A1(n2011), .A2(n2012), .ZN(n2008) );
  OR2_X1 U2015 ( .A1(n2007), .A2(a_11_), .ZN(n2012) );
  NAND2_X1 U2016 ( .A1(n2013), .A2(operation), .ZN(n2001) );
  XNOR2_X1 U2017 ( .A(n2014), .B(n2015), .ZN(n2013) );
  XOR2_X1 U2018 ( .A(n2016), .B(n2017), .Z(n2015) );
  NAND2_X1 U2019 ( .A1(b_15_), .A2(a_11_), .ZN(n2017) );
  NAND2_X1 U2020 ( .A1(n2018), .A2(n2019), .ZN(Result_26_) );
  NAND2_X1 U2021 ( .A1(n2020), .A2(n1911), .ZN(n2019) );
  XOR2_X1 U2022 ( .A(n2021), .B(n2022), .Z(n2020) );
  AND2_X1 U2023 ( .A1(n2023), .A2(n2024), .ZN(n2022) );
  NAND2_X1 U2024 ( .A1(n2025), .A2(operation), .ZN(n2018) );
  XNOR2_X1 U2025 ( .A(n2026), .B(n2027), .ZN(n2025) );
  NAND2_X1 U2026 ( .A1(n2028), .A2(n2029), .ZN(n2026) );
  NAND2_X1 U2027 ( .A1(n2030), .A2(n2031), .ZN(Result_25_) );
  NAND2_X1 U2028 ( .A1(n2032), .A2(n1911), .ZN(n2031) );
  NAND2_X1 U2029 ( .A1(n2033), .A2(n2034), .ZN(n2032) );
  NAND2_X1 U2030 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  NOR2_X1 U2031 ( .A1(n2037), .A2(n2038), .ZN(n2033) );
  NOR2_X1 U2032 ( .A1(b_9_), .A2(n2039), .ZN(n2038) );
  XNOR2_X1 U2033 ( .A(a_9_), .B(n2036), .ZN(n2039) );
  NOR2_X1 U2034 ( .A1(n2040), .A2(n2041), .ZN(n2037) );
  OR2_X1 U2035 ( .A1(n2036), .A2(a_9_), .ZN(n2041) );
  NAND2_X1 U2036 ( .A1(n2042), .A2(operation), .ZN(n2030) );
  XNOR2_X1 U2037 ( .A(n2043), .B(n2044), .ZN(n2042) );
  NAND2_X1 U2038 ( .A1(n2045), .A2(n2046), .ZN(n2043) );
  NAND2_X1 U2039 ( .A1(n2047), .A2(n2048), .ZN(Result_24_) );
  NAND2_X1 U2040 ( .A1(n2049), .A2(n1911), .ZN(n2048) );
  XNOR2_X1 U2041 ( .A(n2050), .B(n2051), .ZN(n2049) );
  NOR2_X1 U2042 ( .A1(n2052), .A2(n2053), .ZN(n2051) );
  NAND2_X1 U2043 ( .A1(n2054), .A2(operation), .ZN(n2047) );
  XOR2_X1 U2044 ( .A(n2055), .B(n2056), .Z(n2054) );
  XOR2_X1 U2045 ( .A(n2057), .B(n2058), .Z(n2055) );
  NOR2_X1 U2046 ( .A1(n2059), .A2(n1950), .ZN(n2058) );
  NAND2_X1 U2047 ( .A1(n2060), .A2(n2061), .ZN(Result_23_) );
  NAND2_X1 U2048 ( .A1(n2062), .A2(n1911), .ZN(n2061) );
  NAND2_X1 U2049 ( .A1(n2063), .A2(n2064), .ZN(n2062) );
  NAND2_X1 U2050 ( .A1(n2065), .A2(n2066), .ZN(n2064) );
  NOR2_X1 U2051 ( .A1(n2067), .A2(n2068), .ZN(n2063) );
  NOR2_X1 U2052 ( .A1(b_7_), .A2(n2069), .ZN(n2068) );
  XNOR2_X1 U2053 ( .A(a_7_), .B(n2066), .ZN(n2069) );
  NOR2_X1 U2054 ( .A1(n2070), .A2(n2071), .ZN(n2067) );
  NAND2_X1 U2055 ( .A1(n2072), .A2(n2073), .ZN(n2071) );
  NAND2_X1 U2056 ( .A1(n2074), .A2(operation), .ZN(n2060) );
  XNOR2_X1 U2057 ( .A(n2075), .B(n2076), .ZN(n2074) );
  XOR2_X1 U2058 ( .A(n2077), .B(n2078), .Z(n2076) );
  NAND2_X1 U2059 ( .A1(b_15_), .A2(a_7_), .ZN(n2078) );
  NAND2_X1 U2060 ( .A1(n2079), .A2(n2080), .ZN(Result_22_) );
  NAND2_X1 U2061 ( .A1(n2081), .A2(n1911), .ZN(n2080) );
  XOR2_X1 U2062 ( .A(n2082), .B(n2083), .Z(n2081) );
  AND2_X1 U2063 ( .A1(n2084), .A2(n2085), .ZN(n2083) );
  NAND2_X1 U2064 ( .A1(n2086), .A2(operation), .ZN(n2079) );
  XNOR2_X1 U2065 ( .A(n2087), .B(n2088), .ZN(n2086) );
  XOR2_X1 U2066 ( .A(n2089), .B(n2090), .Z(n2088) );
  NAND2_X1 U2067 ( .A1(b_15_), .A2(a_6_), .ZN(n2090) );
  NAND2_X1 U2068 ( .A1(n2091), .A2(n2092), .ZN(Result_21_) );
  NAND2_X1 U2069 ( .A1(n2093), .A2(n1911), .ZN(n2092) );
  NAND2_X1 U2070 ( .A1(n2094), .A2(n2095), .ZN(n2093) );
  NAND2_X1 U2071 ( .A1(n2096), .A2(n2097), .ZN(n2095) );
  NOR2_X1 U2072 ( .A1(n2098), .A2(n2099), .ZN(n2094) );
  NOR2_X1 U2073 ( .A1(b_5_), .A2(n2100), .ZN(n2099) );
  XNOR2_X1 U2074 ( .A(a_5_), .B(n2097), .ZN(n2100) );
  NOR2_X1 U2075 ( .A1(n2101), .A2(n2102), .ZN(n2098) );
  OR2_X1 U2076 ( .A1(n2097), .A2(a_5_), .ZN(n2102) );
  NAND2_X1 U2077 ( .A1(n2103), .A2(operation), .ZN(n2091) );
  XOR2_X1 U2078 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR2_X1 U2079 ( .A(n2106), .B(n2107), .Z(n2104) );
  NOR2_X1 U2080 ( .A1(n2108), .A2(n1950), .ZN(n2107) );
  NAND2_X1 U2081 ( .A1(n2109), .A2(n2110), .ZN(Result_20_) );
  NAND2_X1 U2082 ( .A1(n2111), .A2(n1911), .ZN(n2110) );
  XOR2_X1 U2083 ( .A(n2112), .B(n2113), .Z(n2111) );
  AND2_X1 U2084 ( .A1(n2114), .A2(n2115), .ZN(n2113) );
  NAND2_X1 U2085 ( .A1(n2116), .A2(operation), .ZN(n2109) );
  XNOR2_X1 U2086 ( .A(n2117), .B(n2118), .ZN(n2116) );
  XOR2_X1 U2087 ( .A(n2119), .B(n2120), .Z(n2118) );
  NAND2_X1 U2088 ( .A1(b_15_), .A2(a_4_), .ZN(n2120) );
  NOR2_X1 U2089 ( .A1(n1911), .A2(n2121), .ZN(Result_1_) );
  XOR2_X1 U2090 ( .A(n2122), .B(n2123), .Z(n2121) );
  NAND2_X1 U2091 ( .A1(n2124), .A2(n2125), .ZN(n2123) );
  NAND2_X1 U2092 ( .A1(n2126), .A2(n2127), .ZN(Result_19_) );
  NAND2_X1 U2093 ( .A1(n2128), .A2(n1911), .ZN(n2127) );
  NAND2_X1 U2094 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
  NAND2_X1 U2095 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
  NOR2_X1 U2096 ( .A1(n2133), .A2(n2134), .ZN(n2129) );
  NOR2_X1 U2097 ( .A1(b_3_), .A2(n2135), .ZN(n2134) );
  XNOR2_X1 U2098 ( .A(a_3_), .B(n2132), .ZN(n2135) );
  NOR2_X1 U2099 ( .A1(n2136), .A2(n2137), .ZN(n2133) );
  OR2_X1 U2100 ( .A1(n2132), .A2(a_3_), .ZN(n2137) );
  NAND2_X1 U2101 ( .A1(n2138), .A2(operation), .ZN(n2126) );
  XOR2_X1 U2102 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR2_X1 U2103 ( .A(n2141), .B(n2142), .Z(n2139) );
  NOR2_X1 U2104 ( .A1(n2143), .A2(n1950), .ZN(n2142) );
  NAND2_X1 U2105 ( .A1(n2144), .A2(n2145), .ZN(Result_18_) );
  NAND2_X1 U2106 ( .A1(n2146), .A2(n1911), .ZN(n2145) );
  XOR2_X1 U2107 ( .A(n2147), .B(n2148), .Z(n2146) );
  AND2_X1 U2108 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
  NAND2_X1 U2109 ( .A1(n2151), .A2(operation), .ZN(n2144) );
  XNOR2_X1 U2110 ( .A(n2152), .B(n2153), .ZN(n2151) );
  XOR2_X1 U2111 ( .A(n2154), .B(n2155), .Z(n2153) );
  NAND2_X1 U2112 ( .A1(b_15_), .A2(a_2_), .ZN(n2155) );
  NAND2_X1 U2113 ( .A1(n2156), .A2(n2157), .ZN(Result_17_) );
  NAND2_X1 U2114 ( .A1(n2158), .A2(n1911), .ZN(n2157) );
  NAND2_X1 U2115 ( .A1(n2159), .A2(n2160), .ZN(n2158) );
  NAND2_X1 U2116 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
  OR2_X1 U2117 ( .A1(n2163), .A2(n2164), .ZN(n2161) );
  NAND2_X1 U2118 ( .A1(n2165), .A2(n2166), .ZN(n2159) );
  INV_X1 U2119 ( .A(n2162), .ZN(n2166) );
  XNOR2_X1 U2120 ( .A(n2167), .B(a_1_), .ZN(n2165) );
  NAND2_X1 U2121 ( .A1(n2168), .A2(operation), .ZN(n2156) );
  XNOR2_X1 U2122 ( .A(n2169), .B(n2170), .ZN(n2168) );
  XOR2_X1 U2123 ( .A(n2171), .B(n2172), .Z(n2170) );
  NAND2_X1 U2124 ( .A1(b_15_), .A2(a_1_), .ZN(n2172) );
  NAND2_X1 U2125 ( .A1(n2173), .A2(n2174), .ZN(Result_16_) );
  NAND2_X1 U2126 ( .A1(n2175), .A2(n1911), .ZN(n2174) );
  XOR2_X1 U2127 ( .A(n2176), .B(n2177), .Z(n2175) );
  NOR2_X1 U2128 ( .A1(n2178), .A2(n2179), .ZN(n2177) );
  NOR2_X1 U2129 ( .A1(b_0_), .A2(a_0_), .ZN(n2178) );
  NOR2_X1 U2130 ( .A1(n2164), .A2(n2180), .ZN(n2176) );
  NOR2_X1 U2131 ( .A1(n2163), .A2(n2162), .ZN(n2180) );
  NAND2_X1 U2132 ( .A1(n2150), .A2(n2181), .ZN(n2162) );
  NAND2_X1 U2133 ( .A1(n2149), .A2(n2147), .ZN(n2181) );
  NAND2_X1 U2134 ( .A1(n2182), .A2(n2183), .ZN(n2147) );
  NAND2_X1 U2135 ( .A1(n2184), .A2(n2132), .ZN(n2183) );
  NAND2_X1 U2136 ( .A1(n2115), .A2(n2185), .ZN(n2132) );
  NAND2_X1 U2137 ( .A1(n2114), .A2(n2112), .ZN(n2185) );
  NAND2_X1 U2138 ( .A1(n2186), .A2(n2187), .ZN(n2112) );
  NAND2_X1 U2139 ( .A1(n2188), .A2(n2097), .ZN(n2187) );
  NAND2_X1 U2140 ( .A1(n2085), .A2(n2189), .ZN(n2097) );
  NAND2_X1 U2141 ( .A1(n2084), .A2(n2082), .ZN(n2189) );
  NAND2_X1 U2142 ( .A1(n2190), .A2(n2191), .ZN(n2082) );
  NAND2_X1 U2143 ( .A1(n2192), .A2(n2066), .ZN(n2191) );
  INV_X1 U2144 ( .A(n2072), .ZN(n2066) );
  NOR2_X1 U2145 ( .A1(n2053), .A2(n2193), .ZN(n2072) );
  NOR2_X1 U2146 ( .A1(n2052), .A2(n2050), .ZN(n2193) );
  AND2_X1 U2147 ( .A1(n2194), .A2(n2195), .ZN(n2050) );
  NAND2_X1 U2148 ( .A1(n2196), .A2(n2036), .ZN(n2195) );
  NAND2_X1 U2149 ( .A1(n2024), .A2(n2197), .ZN(n2036) );
  NAND2_X1 U2150 ( .A1(n2023), .A2(n2021), .ZN(n2197) );
  NAND2_X1 U2151 ( .A1(n2198), .A2(n2199), .ZN(n2021) );
  NAND2_X1 U2152 ( .A1(n2200), .A2(n2007), .ZN(n2199) );
  NAND2_X1 U2153 ( .A1(n1994), .A2(n2201), .ZN(n2007) );
  NAND2_X1 U2154 ( .A1(n1993), .A2(n1991), .ZN(n2201) );
  NAND2_X1 U2155 ( .A1(n2202), .A2(n2203), .ZN(n1991) );
  NAND2_X1 U2156 ( .A1(n2204), .A2(n1977), .ZN(n2203) );
  NAND2_X1 U2157 ( .A1(n2205), .A2(n2206), .ZN(n1977) );
  NAND2_X1 U2158 ( .A1(b_14_), .A2(n2207), .ZN(n2206) );
  OR2_X1 U2159 ( .A1(a_14_), .A2(n1951), .ZN(n2207) );
  NOR2_X1 U2160 ( .A1(n1950), .A2(n2208), .ZN(n1951) );
  NAND2_X1 U2161 ( .A1(b_15_), .A2(n2209), .ZN(n2205) );
  NAND2_X1 U2162 ( .A1(n1981), .A2(n2210), .ZN(n2204) );
  NAND2_X1 U2163 ( .A1(n2211), .A2(n2000), .ZN(n1993) );
  NAND2_X1 U2164 ( .A1(n2011), .A2(n2212), .ZN(n2200) );
  INV_X1 U2165 ( .A(n2006), .ZN(n2198) );
  NAND2_X1 U2166 ( .A1(n2213), .A2(n2214), .ZN(n2023) );
  NAND2_X1 U2167 ( .A1(n2040), .A2(n2215), .ZN(n2196) );
  NOR2_X1 U2168 ( .A1(b_8_), .A2(a_8_), .ZN(n2052) );
  NAND2_X1 U2169 ( .A1(n2070), .A2(n2073), .ZN(n2192) );
  NAND2_X1 U2170 ( .A1(n2216), .A2(n2217), .ZN(n2084) );
  INV_X1 U2171 ( .A(n2218), .ZN(n2085) );
  NAND2_X1 U2172 ( .A1(n2101), .A2(n2108), .ZN(n2188) );
  INV_X1 U2173 ( .A(n2096), .ZN(n2186) );
  NAND2_X1 U2174 ( .A1(n2219), .A2(n2220), .ZN(n2114) );
  NAND2_X1 U2175 ( .A1(n2136), .A2(n2143), .ZN(n2184) );
  NAND2_X1 U2176 ( .A1(n2221), .A2(n2222), .ZN(n2149) );
  NOR2_X1 U2177 ( .A1(b_1_), .A2(a_1_), .ZN(n2164) );
  NAND2_X1 U2178 ( .A1(n2223), .A2(operation), .ZN(n2173) );
  XOR2_X1 U2179 ( .A(n2224), .B(n2225), .Z(n2223) );
  XOR2_X1 U2180 ( .A(n2226), .B(n2227), .Z(n2224) );
  NOR2_X1 U2181 ( .A1(n2228), .A2(n1950), .ZN(n2227) );
  INV_X1 U2182 ( .A(b_15_), .ZN(n1950) );
  NOR2_X1 U2183 ( .A1(n1911), .A2(n2229), .ZN(Result_15_) );
  XNOR2_X1 U2184 ( .A(n2230), .B(n2231), .ZN(n2229) );
  NOR2_X1 U2185 ( .A1(n1911), .A2(n2232), .ZN(Result_14_) );
  NAND2_X1 U2186 ( .A1(n2233), .A2(n2234), .ZN(n2232) );
  NAND2_X1 U2187 ( .A1(n2235), .A2(n2236), .ZN(n2233) );
  NAND2_X1 U2188 ( .A1(n2231), .A2(n2230), .ZN(n2236) );
  XNOR2_X1 U2189 ( .A(n2237), .B(n2238), .ZN(n2235) );
  NOR2_X1 U2190 ( .A1(n1911), .A2(n2239), .ZN(Result_13_) );
  NAND2_X1 U2191 ( .A1(n2240), .A2(n2241), .ZN(n2239) );
  NAND2_X1 U2192 ( .A1(n2242), .A2(n2234), .ZN(n2241) );
  NAND2_X1 U2193 ( .A1(n2243), .A2(n2244), .ZN(n2242) );
  OR2_X1 U2194 ( .A1(n2245), .A2(n2246), .ZN(n2243) );
  NAND2_X1 U2195 ( .A1(n2247), .A2(n2244), .ZN(n2240) );
  NAND2_X1 U2196 ( .A1(n2245), .A2(n2246), .ZN(n2244) );
  INV_X1 U2197 ( .A(n2234), .ZN(n2247) );
  NOR2_X1 U2198 ( .A1(n2248), .A2(n1911), .ZN(Result_12_) );
  XNOR2_X1 U2199 ( .A(n2249), .B(n2250), .ZN(n2248) );
  NOR2_X1 U2200 ( .A1(n2251), .A2(n1911), .ZN(Result_11_) );
  XNOR2_X1 U2201 ( .A(n2252), .B(n2253), .ZN(n2251) );
  NOR2_X1 U2202 ( .A1(n2254), .A2(n2255), .ZN(n2253) );
  NOR2_X1 U2203 ( .A1(n2256), .A2(n2257), .ZN(n2255) );
  INV_X1 U2204 ( .A(n2258), .ZN(n2254) );
  NOR2_X1 U2205 ( .A1(n1911), .A2(n2259), .ZN(Result_10_) );
  XNOR2_X1 U2206 ( .A(n2260), .B(n2261), .ZN(n2259) );
  NOR2_X1 U2207 ( .A1(n2262), .A2(n2263), .ZN(n2261) );
  AND2_X1 U2208 ( .A1(n2264), .A2(n2265), .ZN(n2263) );
  NOR2_X1 U2209 ( .A1(n2266), .A2(n1911), .ZN(Result_0_) );
  NOR2_X1 U2210 ( .A1(n2267), .A2(n2268), .ZN(n2266) );
  NAND2_X1 U2211 ( .A1(n2269), .A2(n2125), .ZN(n2268) );
  NAND2_X1 U2212 ( .A1(n2270), .A2(n2271), .ZN(n2125) );
  NOR2_X1 U2213 ( .A1(n2272), .A2(n2273), .ZN(n2271) );
  NOR2_X1 U2214 ( .A1(n2274), .A2(n2275), .ZN(n2270) );
  INV_X1 U2215 ( .A(n2179), .ZN(n2274) );
  NAND2_X1 U2216 ( .A1(n2124), .A2(n2122), .ZN(n2269) );
  NAND2_X1 U2217 ( .A1(n1969), .A2(n2276), .ZN(n2122) );
  NAND2_X1 U2218 ( .A1(n1970), .A2(n1967), .ZN(n2276) );
  NAND2_X1 U2219 ( .A1(n1945), .A2(n2277), .ZN(n1967) );
  NAND2_X1 U2220 ( .A1(n1946), .A2(n1943), .ZN(n2277) );
  NAND2_X1 U2221 ( .A1(n1940), .A2(n2278), .ZN(n1943) );
  NAND2_X1 U2222 ( .A1(n1941), .A2(n1938), .ZN(n2278) );
  NAND2_X1 U2223 ( .A1(n1935), .A2(n2279), .ZN(n1938) );
  NAND2_X1 U2224 ( .A1(n1936), .A2(n1933), .ZN(n2279) );
  NAND2_X1 U2225 ( .A1(n1930), .A2(n2280), .ZN(n1933) );
  NAND2_X1 U2226 ( .A1(n1931), .A2(n1928), .ZN(n2280) );
  NAND2_X1 U2227 ( .A1(n1925), .A2(n2281), .ZN(n1928) );
  NAND2_X1 U2228 ( .A1(n1926), .A2(n1923), .ZN(n2281) );
  NAND2_X1 U2229 ( .A1(n1920), .A2(n2282), .ZN(n1923) );
  NAND2_X1 U2230 ( .A1(n1921), .A2(n1918), .ZN(n2282) );
  NAND2_X1 U2231 ( .A1(n1915), .A2(n2283), .ZN(n1918) );
  NAND2_X1 U2232 ( .A1(n1916), .A2(n1913), .ZN(n2283) );
  NAND2_X1 U2233 ( .A1(n2284), .A2(n2285), .ZN(n1913) );
  NAND2_X1 U2234 ( .A1(n2265), .A2(n2264), .ZN(n2285) );
  NAND2_X1 U2235 ( .A1(n2260), .A2(n2286), .ZN(n2284) );
  INV_X1 U2236 ( .A(n2262), .ZN(n2286) );
  NOR2_X1 U2237 ( .A1(n2264), .A2(n2265), .ZN(n2262) );
  XOR2_X1 U2238 ( .A(n2287), .B(n2288), .Z(n2264) );
  NAND2_X1 U2239 ( .A1(n2289), .A2(n2258), .ZN(n2260) );
  NAND2_X1 U2240 ( .A1(n2257), .A2(n2256), .ZN(n2258) );
  AND2_X1 U2241 ( .A1(n2290), .A2(n2291), .ZN(n2256) );
  NAND2_X1 U2242 ( .A1(n2252), .A2(n2257), .ZN(n2289) );
  NOR2_X1 U2243 ( .A1(n2265), .A2(n2292), .ZN(n2257) );
  AND2_X1 U2244 ( .A1(n2293), .A2(n2294), .ZN(n2292) );
  NOR2_X1 U2245 ( .A1(n2294), .A2(n2293), .ZN(n2265) );
  XOR2_X1 U2246 ( .A(n2295), .B(n2296), .Z(n2293) );
  NAND2_X1 U2247 ( .A1(n2297), .A2(n2298), .ZN(n2295) );
  NAND2_X1 U2248 ( .A1(n2299), .A2(n2300), .ZN(n2294) );
  NAND2_X1 U2249 ( .A1(n2301), .A2(n2302), .ZN(n2300) );
  NAND2_X1 U2250 ( .A1(n2303), .A2(n2304), .ZN(n2302) );
  OR2_X1 U2251 ( .A1(n2304), .A2(n2303), .ZN(n2299) );
  NOR2_X1 U2252 ( .A1(n2250), .A2(n2249), .ZN(n2252) );
  AND2_X1 U2253 ( .A1(n2305), .A2(n2306), .ZN(n2249) );
  NAND2_X1 U2254 ( .A1(n2307), .A2(n2308), .ZN(n2305) );
  NAND2_X1 U2255 ( .A1(n2234), .A2(n2245), .ZN(n2308) );
  NAND2_X1 U2256 ( .A1(n2309), .A2(n2310), .ZN(n2234) );
  AND2_X1 U2257 ( .A1(n2230), .A2(n2245), .ZN(n2310) );
  NAND2_X1 U2258 ( .A1(n2237), .A2(n2238), .ZN(n2245) );
  NAND2_X1 U2259 ( .A1(n2311), .A2(n2312), .ZN(n2230) );
  NAND2_X1 U2260 ( .A1(n2313), .A2(b_15_), .ZN(n2312) );
  NOR2_X1 U2261 ( .A1(n2314), .A2(n2228), .ZN(n2313) );
  NOR2_X1 U2262 ( .A1(n2225), .A2(n2226), .ZN(n2314) );
  NAND2_X1 U2263 ( .A1(n2225), .A2(n2226), .ZN(n2311) );
  NAND2_X1 U2264 ( .A1(n2315), .A2(n2316), .ZN(n2226) );
  NAND2_X1 U2265 ( .A1(n2317), .A2(b_15_), .ZN(n2316) );
  NOR2_X1 U2266 ( .A1(n2318), .A2(n2319), .ZN(n2317) );
  NOR2_X1 U2267 ( .A1(n2169), .A2(n2171), .ZN(n2318) );
  NAND2_X1 U2268 ( .A1(n2169), .A2(n2171), .ZN(n2315) );
  NAND2_X1 U2269 ( .A1(n2320), .A2(n2321), .ZN(n2171) );
  NAND2_X1 U2270 ( .A1(n2322), .A2(b_15_), .ZN(n2321) );
  NOR2_X1 U2271 ( .A1(n2323), .A2(n2222), .ZN(n2322) );
  NOR2_X1 U2272 ( .A1(n2152), .A2(n2154), .ZN(n2323) );
  NAND2_X1 U2273 ( .A1(n2152), .A2(n2154), .ZN(n2320) );
  NAND2_X1 U2274 ( .A1(n2324), .A2(n2325), .ZN(n2154) );
  NAND2_X1 U2275 ( .A1(n2326), .A2(b_15_), .ZN(n2325) );
  NOR2_X1 U2276 ( .A1(n2327), .A2(n2143), .ZN(n2326) );
  NOR2_X1 U2277 ( .A1(n2140), .A2(n2141), .ZN(n2327) );
  NAND2_X1 U2278 ( .A1(n2140), .A2(n2141), .ZN(n2324) );
  NAND2_X1 U2279 ( .A1(n2328), .A2(n2329), .ZN(n2141) );
  NAND2_X1 U2280 ( .A1(n2330), .A2(b_15_), .ZN(n2329) );
  NOR2_X1 U2281 ( .A1(n2331), .A2(n2220), .ZN(n2330) );
  NOR2_X1 U2282 ( .A1(n2117), .A2(n2119), .ZN(n2331) );
  NAND2_X1 U2283 ( .A1(n2117), .A2(n2119), .ZN(n2328) );
  NAND2_X1 U2284 ( .A1(n2332), .A2(n2333), .ZN(n2119) );
  NAND2_X1 U2285 ( .A1(n2334), .A2(b_15_), .ZN(n2333) );
  NOR2_X1 U2286 ( .A1(n2335), .A2(n2108), .ZN(n2334) );
  NOR2_X1 U2287 ( .A1(n2105), .A2(n2106), .ZN(n2335) );
  NAND2_X1 U2288 ( .A1(n2105), .A2(n2106), .ZN(n2332) );
  NAND2_X1 U2289 ( .A1(n2336), .A2(n2337), .ZN(n2106) );
  NAND2_X1 U2290 ( .A1(n2338), .A2(b_15_), .ZN(n2337) );
  NOR2_X1 U2291 ( .A1(n2339), .A2(n2217), .ZN(n2338) );
  NOR2_X1 U2292 ( .A1(n2087), .A2(n2089), .ZN(n2339) );
  NAND2_X1 U2293 ( .A1(n2087), .A2(n2089), .ZN(n2336) );
  NAND2_X1 U2294 ( .A1(n2340), .A2(n2341), .ZN(n2089) );
  NAND2_X1 U2295 ( .A1(n2342), .A2(b_15_), .ZN(n2341) );
  NOR2_X1 U2296 ( .A1(n2343), .A2(n2073), .ZN(n2342) );
  NOR2_X1 U2297 ( .A1(n2075), .A2(n2077), .ZN(n2343) );
  NAND2_X1 U2298 ( .A1(n2075), .A2(n2077), .ZN(n2340) );
  NAND2_X1 U2299 ( .A1(n2344), .A2(n2345), .ZN(n2077) );
  NAND2_X1 U2300 ( .A1(n2346), .A2(b_15_), .ZN(n2345) );
  NOR2_X1 U2301 ( .A1(n2347), .A2(n2059), .ZN(n2346) );
  NOR2_X1 U2302 ( .A1(n2056), .A2(n2057), .ZN(n2347) );
  NAND2_X1 U2303 ( .A1(n2056), .A2(n2057), .ZN(n2344) );
  NAND2_X1 U2304 ( .A1(n2045), .A2(n2348), .ZN(n2057) );
  NAND2_X1 U2305 ( .A1(n2044), .A2(n2046), .ZN(n2348) );
  NAND2_X1 U2306 ( .A1(n2349), .A2(n2350), .ZN(n2046) );
  NAND2_X1 U2307 ( .A1(b_15_), .A2(a_9_), .ZN(n2350) );
  INV_X1 U2308 ( .A(n2351), .ZN(n2349) );
  XNOR2_X1 U2309 ( .A(n2352), .B(n2353), .ZN(n2044) );
  XOR2_X1 U2310 ( .A(n2354), .B(n2355), .Z(n2353) );
  NAND2_X1 U2311 ( .A1(b_14_), .A2(a_10_), .ZN(n2355) );
  NAND2_X1 U2312 ( .A1(a_9_), .A2(n2351), .ZN(n2045) );
  NAND2_X1 U2313 ( .A1(n2028), .A2(n2356), .ZN(n2351) );
  NAND2_X1 U2314 ( .A1(n2027), .A2(n2029), .ZN(n2356) );
  NAND2_X1 U2315 ( .A1(n2357), .A2(n2358), .ZN(n2029) );
  NAND2_X1 U2316 ( .A1(b_15_), .A2(a_10_), .ZN(n2358) );
  INV_X1 U2317 ( .A(n2359), .ZN(n2357) );
  XNOR2_X1 U2318 ( .A(n2360), .B(n2361), .ZN(n2027) );
  XNOR2_X1 U2319 ( .A(n2362), .B(n2363), .ZN(n2360) );
  NAND2_X1 U2320 ( .A1(a_10_), .A2(n2359), .ZN(n2028) );
  NAND2_X1 U2321 ( .A1(n2364), .A2(n2365), .ZN(n2359) );
  NAND2_X1 U2322 ( .A1(n2366), .A2(b_15_), .ZN(n2365) );
  NOR2_X1 U2323 ( .A1(n2367), .A2(n2212), .ZN(n2366) );
  NOR2_X1 U2324 ( .A1(n2014), .A2(n2016), .ZN(n2367) );
  NAND2_X1 U2325 ( .A1(n2014), .A2(n2016), .ZN(n2364) );
  NAND2_X1 U2326 ( .A1(n2368), .A2(n2369), .ZN(n2016) );
  NAND2_X1 U2327 ( .A1(n2370), .A2(b_15_), .ZN(n2369) );
  NOR2_X1 U2328 ( .A1(n2371), .A2(n2000), .ZN(n2370) );
  NOR2_X1 U2329 ( .A1(n1996), .A2(n1998), .ZN(n2371) );
  NAND2_X1 U2330 ( .A1(n1996), .A2(n1998), .ZN(n2368) );
  NAND2_X1 U2331 ( .A1(n2372), .A2(n2373), .ZN(n1998) );
  NAND2_X1 U2332 ( .A1(n2374), .A2(b_15_), .ZN(n2373) );
  NOR2_X1 U2333 ( .A1(n2375), .A2(n2210), .ZN(n2374) );
  NOR2_X1 U2334 ( .A1(n1986), .A2(n1987), .ZN(n2375) );
  NAND2_X1 U2335 ( .A1(n1986), .A2(n1987), .ZN(n2372) );
  NAND2_X1 U2336 ( .A1(n2376), .A2(n2377), .ZN(n1987) );
  NAND2_X1 U2337 ( .A1(b_13_), .A2(n2378), .ZN(n2377) );
  NAND2_X1 U2338 ( .A1(n1958), .A2(n2379), .ZN(n2378) );
  NAND2_X1 U2339 ( .A1(a_15_), .A2(n1963), .ZN(n2379) );
  INV_X1 U2340 ( .A(n2380), .ZN(n1958) );
  NAND2_X1 U2341 ( .A1(b_14_), .A2(n2381), .ZN(n2376) );
  NAND2_X1 U2342 ( .A1(n1961), .A2(n2382), .ZN(n2381) );
  NAND2_X1 U2343 ( .A1(a_14_), .A2(n1981), .ZN(n2382) );
  INV_X1 U2344 ( .A(n2383), .ZN(n1961) );
  AND2_X1 U2345 ( .A1(n2384), .A2(b_15_), .ZN(n1986) );
  NOR2_X1 U2346 ( .A1(n2385), .A2(n1963), .ZN(n2384) );
  XOR2_X1 U2347 ( .A(n2386), .B(n2387), .Z(n1996) );
  NOR2_X1 U2348 ( .A1(n2210), .A2(n1963), .ZN(n2387) );
  XOR2_X1 U2349 ( .A(n2388), .B(n2389), .Z(n2386) );
  XNOR2_X1 U2350 ( .A(n2390), .B(n2391), .ZN(n2014) );
  NAND2_X1 U2351 ( .A1(n2392), .A2(n2393), .ZN(n2390) );
  XNOR2_X1 U2352 ( .A(n2394), .B(n2395), .ZN(n2056) );
  XNOR2_X1 U2353 ( .A(n2396), .B(n2397), .ZN(n2394) );
  XOR2_X1 U2354 ( .A(n2398), .B(n2399), .Z(n2075) );
  XOR2_X1 U2355 ( .A(n2400), .B(n2401), .Z(n2398) );
  NOR2_X1 U2356 ( .A1(n2059), .A2(n1963), .ZN(n2401) );
  XNOR2_X1 U2357 ( .A(n2402), .B(n2403), .ZN(n2087) );
  XNOR2_X1 U2358 ( .A(n2404), .B(n2405), .ZN(n2403) );
  XOR2_X1 U2359 ( .A(n2406), .B(n2407), .Z(n2105) );
  XOR2_X1 U2360 ( .A(n2408), .B(n2409), .Z(n2406) );
  NOR2_X1 U2361 ( .A1(n2217), .A2(n1963), .ZN(n2409) );
  XOR2_X1 U2362 ( .A(n2410), .B(n2411), .Z(n2117) );
  XOR2_X1 U2363 ( .A(n2412), .B(n2413), .Z(n2410) );
  XNOR2_X1 U2364 ( .A(n2414), .B(n2415), .ZN(n2140) );
  XOR2_X1 U2365 ( .A(n2416), .B(n2417), .Z(n2415) );
  NAND2_X1 U2366 ( .A1(b_14_), .A2(a_4_), .ZN(n2417) );
  XOR2_X1 U2367 ( .A(n2418), .B(n2419), .Z(n2152) );
  XOR2_X1 U2368 ( .A(n2420), .B(n2421), .Z(n2418) );
  XOR2_X1 U2369 ( .A(n2422), .B(n2423), .Z(n2169) );
  XOR2_X1 U2370 ( .A(n2424), .B(n2425), .Z(n2422) );
  NOR2_X1 U2371 ( .A1(n2222), .A2(n1963), .ZN(n2425) );
  XNOR2_X1 U2372 ( .A(n2426), .B(n2427), .ZN(n2225) );
  NAND2_X1 U2373 ( .A1(n2428), .A2(n2429), .ZN(n2426) );
  NOR2_X1 U2374 ( .A1(n2430), .A2(n2431), .ZN(n2309) );
  INV_X1 U2375 ( .A(n2231), .ZN(n2431) );
  XNOR2_X1 U2376 ( .A(n2432), .B(n2433), .ZN(n2231) );
  XNOR2_X1 U2377 ( .A(n2434), .B(n2435), .ZN(n2432) );
  NOR2_X1 U2378 ( .A1(n2237), .A2(n2238), .ZN(n2430) );
  NAND2_X1 U2379 ( .A1(n2436), .A2(n2437), .ZN(n2238) );
  NAND2_X1 U2380 ( .A1(n2435), .A2(n2438), .ZN(n2437) );
  NAND2_X1 U2381 ( .A1(n2434), .A2(n2433), .ZN(n2438) );
  NOR2_X1 U2382 ( .A1(n1963), .A2(n2228), .ZN(n2435) );
  OR2_X1 U2383 ( .A1(n2433), .A2(n2434), .ZN(n2436) );
  AND2_X1 U2384 ( .A1(n2428), .A2(n2439), .ZN(n2434) );
  NAND2_X1 U2385 ( .A1(n2427), .A2(n2429), .ZN(n2439) );
  NAND2_X1 U2386 ( .A1(n2440), .A2(n2441), .ZN(n2429) );
  NAND2_X1 U2387 ( .A1(b_14_), .A2(a_1_), .ZN(n2441) );
  INV_X1 U2388 ( .A(n2442), .ZN(n2440) );
  XNOR2_X1 U2389 ( .A(n2443), .B(n2444), .ZN(n2427) );
  XNOR2_X1 U2390 ( .A(n2445), .B(n2446), .ZN(n2443) );
  NAND2_X1 U2391 ( .A1(a_1_), .A2(n2442), .ZN(n2428) );
  NAND2_X1 U2392 ( .A1(n2447), .A2(n2448), .ZN(n2442) );
  NAND2_X1 U2393 ( .A1(n2449), .A2(b_14_), .ZN(n2448) );
  NOR2_X1 U2394 ( .A1(n2450), .A2(n2222), .ZN(n2449) );
  NOR2_X1 U2395 ( .A1(n2423), .A2(n2424), .ZN(n2450) );
  NAND2_X1 U2396 ( .A1(n2423), .A2(n2424), .ZN(n2447) );
  NAND2_X1 U2397 ( .A1(n2451), .A2(n2452), .ZN(n2424) );
  NAND2_X1 U2398 ( .A1(n2421), .A2(n2453), .ZN(n2452) );
  OR2_X1 U2399 ( .A1(n2420), .A2(n2419), .ZN(n2453) );
  NOR2_X1 U2400 ( .A1(n1963), .A2(n2143), .ZN(n2421) );
  NAND2_X1 U2401 ( .A1(n2419), .A2(n2420), .ZN(n2451) );
  NAND2_X1 U2402 ( .A1(n2454), .A2(n2455), .ZN(n2420) );
  NAND2_X1 U2403 ( .A1(n2456), .A2(b_14_), .ZN(n2455) );
  NOR2_X1 U2404 ( .A1(n2457), .A2(n2220), .ZN(n2456) );
  NOR2_X1 U2405 ( .A1(n2414), .A2(n2416), .ZN(n2457) );
  NAND2_X1 U2406 ( .A1(n2414), .A2(n2416), .ZN(n2454) );
  NAND2_X1 U2407 ( .A1(n2458), .A2(n2459), .ZN(n2416) );
  NAND2_X1 U2408 ( .A1(n2413), .A2(n2460), .ZN(n2459) );
  OR2_X1 U2409 ( .A1(n2412), .A2(n2411), .ZN(n2460) );
  NOR2_X1 U2410 ( .A1(n1963), .A2(n2108), .ZN(n2413) );
  NAND2_X1 U2411 ( .A1(n2411), .A2(n2412), .ZN(n2458) );
  NAND2_X1 U2412 ( .A1(n2461), .A2(n2462), .ZN(n2412) );
  NAND2_X1 U2413 ( .A1(n2463), .A2(b_14_), .ZN(n2462) );
  NOR2_X1 U2414 ( .A1(n2464), .A2(n2217), .ZN(n2463) );
  NOR2_X1 U2415 ( .A1(n2407), .A2(n2408), .ZN(n2464) );
  NAND2_X1 U2416 ( .A1(n2407), .A2(n2408), .ZN(n2461) );
  NAND2_X1 U2417 ( .A1(n2465), .A2(n2466), .ZN(n2408) );
  NAND2_X1 U2418 ( .A1(n2405), .A2(n2467), .ZN(n2466) );
  OR2_X1 U2419 ( .A1(n2404), .A2(n2402), .ZN(n2467) );
  NOR2_X1 U2420 ( .A1(n1963), .A2(n2073), .ZN(n2405) );
  NAND2_X1 U2421 ( .A1(n2402), .A2(n2404), .ZN(n2465) );
  NAND2_X1 U2422 ( .A1(n2468), .A2(n2469), .ZN(n2404) );
  NAND2_X1 U2423 ( .A1(n2470), .A2(b_14_), .ZN(n2469) );
  NOR2_X1 U2424 ( .A1(n2471), .A2(n2059), .ZN(n2470) );
  NOR2_X1 U2425 ( .A1(n2399), .A2(n2400), .ZN(n2471) );
  NAND2_X1 U2426 ( .A1(n2399), .A2(n2400), .ZN(n2468) );
  NAND2_X1 U2427 ( .A1(n2472), .A2(n2473), .ZN(n2400) );
  NAND2_X1 U2428 ( .A1(n2397), .A2(n2474), .ZN(n2473) );
  NAND2_X1 U2429 ( .A1(n2396), .A2(n2395), .ZN(n2474) );
  NOR2_X1 U2430 ( .A1(n1963), .A2(n2215), .ZN(n2397) );
  OR2_X1 U2431 ( .A1(n2395), .A2(n2396), .ZN(n2472) );
  AND2_X1 U2432 ( .A1(n2475), .A2(n2476), .ZN(n2396) );
  NAND2_X1 U2433 ( .A1(n2477), .A2(b_14_), .ZN(n2476) );
  NOR2_X1 U2434 ( .A1(n2478), .A2(n2214), .ZN(n2477) );
  NOR2_X1 U2435 ( .A1(n2352), .A2(n2354), .ZN(n2478) );
  NAND2_X1 U2436 ( .A1(n2352), .A2(n2354), .ZN(n2475) );
  NAND2_X1 U2437 ( .A1(n2479), .A2(n2480), .ZN(n2354) );
  NAND2_X1 U2438 ( .A1(n2363), .A2(n2481), .ZN(n2480) );
  NAND2_X1 U2439 ( .A1(n2362), .A2(n2361), .ZN(n2481) );
  NOR2_X1 U2440 ( .A1(n1963), .A2(n2212), .ZN(n2363) );
  INV_X1 U2441 ( .A(b_14_), .ZN(n1963) );
  OR2_X1 U2442 ( .A1(n2361), .A2(n2362), .ZN(n2479) );
  AND2_X1 U2443 ( .A1(n2392), .A2(n2482), .ZN(n2362) );
  NAND2_X1 U2444 ( .A1(n2391), .A2(n2393), .ZN(n2482) );
  NAND2_X1 U2445 ( .A1(n2483), .A2(n2484), .ZN(n2393) );
  NAND2_X1 U2446 ( .A1(b_14_), .A2(a_12_), .ZN(n2484) );
  INV_X1 U2447 ( .A(n2485), .ZN(n2483) );
  XOR2_X1 U2448 ( .A(n2486), .B(n2487), .Z(n2391) );
  XNOR2_X1 U2449 ( .A(n1976), .B(n2488), .ZN(n2486) );
  NAND2_X1 U2450 ( .A1(a_12_), .A2(n2485), .ZN(n2392) );
  NAND2_X1 U2451 ( .A1(n2489), .A2(n2490), .ZN(n2485) );
  NAND2_X1 U2452 ( .A1(n2491), .A2(b_14_), .ZN(n2490) );
  NOR2_X1 U2453 ( .A1(n2492), .A2(n2210), .ZN(n2491) );
  NOR2_X1 U2454 ( .A1(n2388), .A2(n2389), .ZN(n2492) );
  NAND2_X1 U2455 ( .A1(n2388), .A2(n2389), .ZN(n2489) );
  NAND2_X1 U2456 ( .A1(n2493), .A2(n2494), .ZN(n2389) );
  NAND2_X1 U2457 ( .A1(n2495), .A2(b_12_), .ZN(n2494) );
  NOR2_X1 U2458 ( .A1(n2496), .A2(n2208), .ZN(n2495) );
  NOR2_X1 U2459 ( .A1(n2380), .A2(n1981), .ZN(n2496) );
  NAND2_X1 U2460 ( .A1(n2497), .A2(b_13_), .ZN(n2493) );
  NOR2_X1 U2461 ( .A1(n2498), .A2(n2499), .ZN(n2497) );
  NOR2_X1 U2462 ( .A1(n2383), .A2(n2211), .ZN(n2498) );
  AND2_X1 U2463 ( .A1(n2500), .A2(b_14_), .ZN(n2388) );
  NOR2_X1 U2464 ( .A1(n2385), .A2(n1981), .ZN(n2500) );
  XOR2_X1 U2465 ( .A(n2501), .B(n2502), .Z(n2361) );
  NAND2_X1 U2466 ( .A1(n2503), .A2(n2504), .ZN(n2501) );
  XOR2_X1 U2467 ( .A(n2505), .B(n2506), .Z(n2352) );
  XOR2_X1 U2468 ( .A(n2507), .B(n2508), .Z(n2505) );
  XOR2_X1 U2469 ( .A(n2509), .B(n2510), .Z(n2395) );
  XOR2_X1 U2470 ( .A(n2511), .B(n2512), .Z(n2510) );
  NAND2_X1 U2471 ( .A1(b_13_), .A2(a_10_), .ZN(n2512) );
  XNOR2_X1 U2472 ( .A(n2513), .B(n2514), .ZN(n2399) );
  XOR2_X1 U2473 ( .A(n2515), .B(n2516), .Z(n2514) );
  NAND2_X1 U2474 ( .A1(b_13_), .A2(a_9_), .ZN(n2516) );
  XNOR2_X1 U2475 ( .A(n2517), .B(n2518), .ZN(n2402) );
  NAND2_X1 U2476 ( .A1(n2519), .A2(n2520), .ZN(n2517) );
  XOR2_X1 U2477 ( .A(n2521), .B(n2522), .Z(n2407) );
  XOR2_X1 U2478 ( .A(n2523), .B(n2524), .Z(n2521) );
  XOR2_X1 U2479 ( .A(n2525), .B(n2526), .Z(n2411) );
  XOR2_X1 U2480 ( .A(n2527), .B(n2528), .Z(n2525) );
  NOR2_X1 U2481 ( .A1(n2217), .A2(n1981), .ZN(n2528) );
  XOR2_X1 U2482 ( .A(n2529), .B(n2530), .Z(n2414) );
  XOR2_X1 U2483 ( .A(n2531), .B(n2532), .Z(n2529) );
  XNOR2_X1 U2484 ( .A(n2533), .B(n2534), .ZN(n2419) );
  XOR2_X1 U2485 ( .A(n2535), .B(n2536), .Z(n2534) );
  NAND2_X1 U2486 ( .A1(b_13_), .A2(a_4_), .ZN(n2536) );
  XNOR2_X1 U2487 ( .A(n2537), .B(n2538), .ZN(n2423) );
  XNOR2_X1 U2488 ( .A(n2539), .B(n2540), .ZN(n2537) );
  XOR2_X1 U2489 ( .A(n2541), .B(n2542), .Z(n2433) );
  NAND2_X1 U2490 ( .A1(n2543), .A2(n2544), .ZN(n2541) );
  XOR2_X1 U2491 ( .A(n2545), .B(n2546), .Z(n2237) );
  XNOR2_X1 U2492 ( .A(n2547), .B(n2548), .ZN(n2545) );
  INV_X1 U2493 ( .A(n2246), .ZN(n2307) );
  NAND2_X1 U2494 ( .A1(n2549), .A2(n2306), .ZN(n2246) );
  NAND2_X1 U2495 ( .A1(n2550), .A2(n2551), .ZN(n2306) );
  OR2_X1 U2496 ( .A1(n2551), .A2(n2550), .ZN(n2549) );
  AND2_X1 U2497 ( .A1(n2552), .A2(n2553), .ZN(n2550) );
  NAND2_X1 U2498 ( .A1(n2547), .A2(n2554), .ZN(n2553) );
  NAND2_X1 U2499 ( .A1(n2548), .A2(n2546), .ZN(n2554) );
  AND2_X1 U2500 ( .A1(n2543), .A2(n2555), .ZN(n2547) );
  NAND2_X1 U2501 ( .A1(n2542), .A2(n2544), .ZN(n2555) );
  NAND2_X1 U2502 ( .A1(n2556), .A2(n2557), .ZN(n2544) );
  NAND2_X1 U2503 ( .A1(b_13_), .A2(a_1_), .ZN(n2557) );
  INV_X1 U2504 ( .A(n2558), .ZN(n2556) );
  XOR2_X1 U2505 ( .A(n2559), .B(n2560), .Z(n2542) );
  XOR2_X1 U2506 ( .A(n2561), .B(n2562), .Z(n2559) );
  NAND2_X1 U2507 ( .A1(a_1_), .A2(n2558), .ZN(n2543) );
  NAND2_X1 U2508 ( .A1(n2563), .A2(n2564), .ZN(n2558) );
  NAND2_X1 U2509 ( .A1(n2446), .A2(n2565), .ZN(n2564) );
  NAND2_X1 U2510 ( .A1(n2445), .A2(n2444), .ZN(n2565) );
  NOR2_X1 U2511 ( .A1(n1981), .A2(n2222), .ZN(n2446) );
  OR2_X1 U2512 ( .A1(n2444), .A2(n2445), .ZN(n2563) );
  AND2_X1 U2513 ( .A1(n2566), .A2(n2567), .ZN(n2445) );
  NAND2_X1 U2514 ( .A1(n2540), .A2(n2568), .ZN(n2567) );
  NAND2_X1 U2515 ( .A1(n2539), .A2(n2538), .ZN(n2568) );
  NOR2_X1 U2516 ( .A1(n1981), .A2(n2143), .ZN(n2540) );
  OR2_X1 U2517 ( .A1(n2538), .A2(n2539), .ZN(n2566) );
  AND2_X1 U2518 ( .A1(n2569), .A2(n2570), .ZN(n2539) );
  NAND2_X1 U2519 ( .A1(n2571), .A2(b_13_), .ZN(n2570) );
  NOR2_X1 U2520 ( .A1(n2572), .A2(n2220), .ZN(n2571) );
  NOR2_X1 U2521 ( .A1(n2533), .A2(n2535), .ZN(n2572) );
  NAND2_X1 U2522 ( .A1(n2533), .A2(n2535), .ZN(n2569) );
  NAND2_X1 U2523 ( .A1(n2573), .A2(n2574), .ZN(n2535) );
  NAND2_X1 U2524 ( .A1(n2532), .A2(n2575), .ZN(n2574) );
  OR2_X1 U2525 ( .A1(n2531), .A2(n2530), .ZN(n2575) );
  NOR2_X1 U2526 ( .A1(n1981), .A2(n2108), .ZN(n2532) );
  NAND2_X1 U2527 ( .A1(n2530), .A2(n2531), .ZN(n2573) );
  NAND2_X1 U2528 ( .A1(n2576), .A2(n2577), .ZN(n2531) );
  NAND2_X1 U2529 ( .A1(n2578), .A2(b_13_), .ZN(n2577) );
  NOR2_X1 U2530 ( .A1(n2579), .A2(n2217), .ZN(n2578) );
  NOR2_X1 U2531 ( .A1(n2526), .A2(n2527), .ZN(n2579) );
  NAND2_X1 U2532 ( .A1(n2526), .A2(n2527), .ZN(n2576) );
  NAND2_X1 U2533 ( .A1(n2580), .A2(n2581), .ZN(n2527) );
  NAND2_X1 U2534 ( .A1(n2524), .A2(n2582), .ZN(n2581) );
  OR2_X1 U2535 ( .A1(n2523), .A2(n2522), .ZN(n2582) );
  NOR2_X1 U2536 ( .A1(n1981), .A2(n2073), .ZN(n2524) );
  NAND2_X1 U2537 ( .A1(n2522), .A2(n2523), .ZN(n2580) );
  NAND2_X1 U2538 ( .A1(n2519), .A2(n2583), .ZN(n2523) );
  NAND2_X1 U2539 ( .A1(n2518), .A2(n2520), .ZN(n2583) );
  NAND2_X1 U2540 ( .A1(n2584), .A2(n2585), .ZN(n2520) );
  NAND2_X1 U2541 ( .A1(b_13_), .A2(a_8_), .ZN(n2585) );
  INV_X1 U2542 ( .A(n2586), .ZN(n2584) );
  XOR2_X1 U2543 ( .A(n2587), .B(n2588), .Z(n2518) );
  XOR2_X1 U2544 ( .A(n2589), .B(n2590), .Z(n2587) );
  NOR2_X1 U2545 ( .A1(n2215), .A2(n2211), .ZN(n2590) );
  NAND2_X1 U2546 ( .A1(a_8_), .A2(n2586), .ZN(n2519) );
  NAND2_X1 U2547 ( .A1(n2591), .A2(n2592), .ZN(n2586) );
  NAND2_X1 U2548 ( .A1(n2593), .A2(b_13_), .ZN(n2592) );
  NOR2_X1 U2549 ( .A1(n2594), .A2(n2215), .ZN(n2593) );
  NOR2_X1 U2550 ( .A1(n2513), .A2(n2515), .ZN(n2594) );
  NAND2_X1 U2551 ( .A1(n2513), .A2(n2515), .ZN(n2591) );
  NAND2_X1 U2552 ( .A1(n2595), .A2(n2596), .ZN(n2515) );
  NAND2_X1 U2553 ( .A1(n2597), .A2(b_13_), .ZN(n2596) );
  NOR2_X1 U2554 ( .A1(n2598), .A2(n2214), .ZN(n2597) );
  NOR2_X1 U2555 ( .A1(n2509), .A2(n2511), .ZN(n2598) );
  NAND2_X1 U2556 ( .A1(n2509), .A2(n2511), .ZN(n2595) );
  NAND2_X1 U2557 ( .A1(n2599), .A2(n2600), .ZN(n2511) );
  NAND2_X1 U2558 ( .A1(n2508), .A2(n2601), .ZN(n2600) );
  OR2_X1 U2559 ( .A1(n2507), .A2(n2506), .ZN(n2601) );
  NOR2_X1 U2560 ( .A1(n1981), .A2(n2212), .ZN(n2508) );
  NAND2_X1 U2561 ( .A1(n2506), .A2(n2507), .ZN(n2599) );
  NAND2_X1 U2562 ( .A1(n2503), .A2(n2602), .ZN(n2507) );
  NAND2_X1 U2563 ( .A1(n2502), .A2(n2504), .ZN(n2602) );
  NAND2_X1 U2564 ( .A1(n2603), .A2(n2604), .ZN(n2504) );
  NAND2_X1 U2565 ( .A1(b_13_), .A2(a_12_), .ZN(n2604) );
  INV_X1 U2566 ( .A(n2605), .ZN(n2603) );
  XOR2_X1 U2567 ( .A(n2606), .B(n2607), .Z(n2502) );
  NOR2_X1 U2568 ( .A1(n2210), .A2(n2211), .ZN(n2607) );
  XOR2_X1 U2569 ( .A(n2608), .B(n2609), .Z(n2606) );
  NAND2_X1 U2570 ( .A1(a_12_), .A2(n2605), .ZN(n2503) );
  NAND2_X1 U2571 ( .A1(n2610), .A2(n2611), .ZN(n2605) );
  NAND2_X1 U2572 ( .A1(n2487), .A2(n2612), .ZN(n2611) );
  NAND2_X1 U2573 ( .A1(n2488), .A2(n2202), .ZN(n2612) );
  INV_X1 U2574 ( .A(n1976), .ZN(n2202) );
  INV_X1 U2575 ( .A(n2613), .ZN(n2488) );
  AND2_X1 U2576 ( .A1(n2614), .A2(b_13_), .ZN(n2487) );
  NOR2_X1 U2577 ( .A1(n2385), .A2(n2211), .ZN(n2614) );
  NAND2_X1 U2578 ( .A1(n1976), .A2(n2613), .ZN(n2610) );
  NAND2_X1 U2579 ( .A1(n2615), .A2(n2616), .ZN(n2613) );
  NAND2_X1 U2580 ( .A1(n2617), .A2(a_15_), .ZN(n2616) );
  NOR2_X1 U2581 ( .A1(n2618), .A2(n2011), .ZN(n2617) );
  NOR2_X1 U2582 ( .A1(n2380), .A2(n2211), .ZN(n2618) );
  NAND2_X1 U2583 ( .A1(n2619), .A2(b_12_), .ZN(n2615) );
  NOR2_X1 U2584 ( .A1(n2620), .A2(n2499), .ZN(n2619) );
  NOR2_X1 U2585 ( .A1(n2383), .A2(n2011), .ZN(n2620) );
  NOR2_X1 U2586 ( .A1(n1981), .A2(n2210), .ZN(n1976) );
  XOR2_X1 U2587 ( .A(n2621), .B(n2622), .Z(n2506) );
  XNOR2_X1 U2588 ( .A(n2623), .B(n2624), .ZN(n2621) );
  XNOR2_X1 U2589 ( .A(n2625), .B(n2626), .ZN(n2509) );
  XNOR2_X1 U2590 ( .A(n2627), .B(n2628), .ZN(n2625) );
  XOR2_X1 U2591 ( .A(n2629), .B(n2630), .Z(n2513) );
  XNOR2_X1 U2592 ( .A(n2631), .B(n2632), .ZN(n2629) );
  NAND2_X1 U2593 ( .A1(b_12_), .A2(a_10_), .ZN(n2631) );
  XNOR2_X1 U2594 ( .A(n2633), .B(n2634), .ZN(n2522) );
  NAND2_X1 U2595 ( .A1(n2635), .A2(n2636), .ZN(n2633) );
  XOR2_X1 U2596 ( .A(n2637), .B(n2638), .Z(n2526) );
  XOR2_X1 U2597 ( .A(n2639), .B(n2640), .Z(n2637) );
  XOR2_X1 U2598 ( .A(n2641), .B(n2642), .Z(n2530) );
  XOR2_X1 U2599 ( .A(n2643), .B(n2644), .Z(n2641) );
  NOR2_X1 U2600 ( .A1(n2217), .A2(n2211), .ZN(n2644) );
  XOR2_X1 U2601 ( .A(n2645), .B(n2646), .Z(n2533) );
  XOR2_X1 U2602 ( .A(n2647), .B(n2648), .Z(n2645) );
  XOR2_X1 U2603 ( .A(n2649), .B(n2650), .Z(n2538) );
  XOR2_X1 U2604 ( .A(n2651), .B(n2652), .Z(n2650) );
  NAND2_X1 U2605 ( .A1(b_12_), .A2(a_4_), .ZN(n2652) );
  XNOR2_X1 U2606 ( .A(n2653), .B(n2654), .ZN(n2444) );
  XOR2_X1 U2607 ( .A(n2655), .B(n2656), .Z(n2653) );
  NOR2_X1 U2608 ( .A1(n2143), .A2(n2211), .ZN(n2656) );
  OR2_X1 U2609 ( .A1(n2546), .A2(n2548), .ZN(n2552) );
  NOR2_X1 U2610 ( .A1(n1981), .A2(n2228), .ZN(n2548) );
  INV_X1 U2611 ( .A(b_13_), .ZN(n1981) );
  XNOR2_X1 U2612 ( .A(n2657), .B(n2658), .ZN(n2546) );
  XNOR2_X1 U2613 ( .A(n2659), .B(n2660), .ZN(n2657) );
  XOR2_X1 U2614 ( .A(n2661), .B(n2662), .Z(n2551) );
  XOR2_X1 U2615 ( .A(n2663), .B(n2664), .Z(n2661) );
  NOR2_X1 U2616 ( .A1(n2228), .A2(n2211), .ZN(n2664) );
  XNOR2_X1 U2617 ( .A(n2290), .B(n2291), .ZN(n2250) );
  NAND2_X1 U2618 ( .A1(n2665), .A2(n2666), .ZN(n2291) );
  NAND2_X1 U2619 ( .A1(n2667), .A2(b_12_), .ZN(n2666) );
  NOR2_X1 U2620 ( .A1(n2668), .A2(n2228), .ZN(n2667) );
  NOR2_X1 U2621 ( .A1(n2662), .A2(n2663), .ZN(n2668) );
  NAND2_X1 U2622 ( .A1(n2662), .A2(n2663), .ZN(n2665) );
  NAND2_X1 U2623 ( .A1(n2669), .A2(n2670), .ZN(n2663) );
  NAND2_X1 U2624 ( .A1(n2660), .A2(n2671), .ZN(n2670) );
  NAND2_X1 U2625 ( .A1(n2659), .A2(n2658), .ZN(n2671) );
  NOR2_X1 U2626 ( .A1(n2211), .A2(n2319), .ZN(n2660) );
  OR2_X1 U2627 ( .A1(n2658), .A2(n2659), .ZN(n2669) );
  AND2_X1 U2628 ( .A1(n2672), .A2(n2673), .ZN(n2659) );
  NAND2_X1 U2629 ( .A1(n2562), .A2(n2674), .ZN(n2673) );
  OR2_X1 U2630 ( .A1(n2561), .A2(n2560), .ZN(n2674) );
  NOR2_X1 U2631 ( .A1(n2211), .A2(n2222), .ZN(n2562) );
  NAND2_X1 U2632 ( .A1(n2560), .A2(n2561), .ZN(n2672) );
  NAND2_X1 U2633 ( .A1(n2675), .A2(n2676), .ZN(n2561) );
  NAND2_X1 U2634 ( .A1(n2677), .A2(b_12_), .ZN(n2676) );
  NOR2_X1 U2635 ( .A1(n2678), .A2(n2143), .ZN(n2677) );
  NOR2_X1 U2636 ( .A1(n2654), .A2(n2655), .ZN(n2678) );
  NAND2_X1 U2637 ( .A1(n2654), .A2(n2655), .ZN(n2675) );
  NAND2_X1 U2638 ( .A1(n2679), .A2(n2680), .ZN(n2655) );
  NAND2_X1 U2639 ( .A1(n2681), .A2(b_12_), .ZN(n2680) );
  NOR2_X1 U2640 ( .A1(n2682), .A2(n2220), .ZN(n2681) );
  NOR2_X1 U2641 ( .A1(n2649), .A2(n2651), .ZN(n2682) );
  NAND2_X1 U2642 ( .A1(n2649), .A2(n2651), .ZN(n2679) );
  NAND2_X1 U2643 ( .A1(n2683), .A2(n2684), .ZN(n2651) );
  NAND2_X1 U2644 ( .A1(n2648), .A2(n2685), .ZN(n2684) );
  OR2_X1 U2645 ( .A1(n2647), .A2(n2646), .ZN(n2685) );
  NOR2_X1 U2646 ( .A1(n2211), .A2(n2108), .ZN(n2648) );
  NAND2_X1 U2647 ( .A1(n2646), .A2(n2647), .ZN(n2683) );
  NAND2_X1 U2648 ( .A1(n2686), .A2(n2687), .ZN(n2647) );
  NAND2_X1 U2649 ( .A1(n2688), .A2(b_12_), .ZN(n2687) );
  NOR2_X1 U2650 ( .A1(n2689), .A2(n2217), .ZN(n2688) );
  NOR2_X1 U2651 ( .A1(n2642), .A2(n2643), .ZN(n2689) );
  NAND2_X1 U2652 ( .A1(n2642), .A2(n2643), .ZN(n2686) );
  NAND2_X1 U2653 ( .A1(n2690), .A2(n2691), .ZN(n2643) );
  NAND2_X1 U2654 ( .A1(n2640), .A2(n2692), .ZN(n2691) );
  OR2_X1 U2655 ( .A1(n2639), .A2(n2638), .ZN(n2692) );
  NOR2_X1 U2656 ( .A1(n2211), .A2(n2073), .ZN(n2640) );
  NAND2_X1 U2657 ( .A1(n2638), .A2(n2639), .ZN(n2690) );
  NAND2_X1 U2658 ( .A1(n2635), .A2(n2693), .ZN(n2639) );
  NAND2_X1 U2659 ( .A1(n2634), .A2(n2636), .ZN(n2693) );
  NAND2_X1 U2660 ( .A1(n2694), .A2(n2695), .ZN(n2636) );
  NAND2_X1 U2661 ( .A1(b_12_), .A2(a_8_), .ZN(n2695) );
  INV_X1 U2662 ( .A(n2696), .ZN(n2694) );
  XOR2_X1 U2663 ( .A(n2697), .B(n2698), .Z(n2634) );
  XOR2_X1 U2664 ( .A(n2699), .B(n2700), .Z(n2697) );
  NOR2_X1 U2665 ( .A1(n2011), .A2(n2215), .ZN(n2700) );
  NAND2_X1 U2666 ( .A1(a_8_), .A2(n2696), .ZN(n2635) );
  NAND2_X1 U2667 ( .A1(n2701), .A2(n2702), .ZN(n2696) );
  NAND2_X1 U2668 ( .A1(n2703), .A2(b_12_), .ZN(n2702) );
  NOR2_X1 U2669 ( .A1(n2704), .A2(n2215), .ZN(n2703) );
  NOR2_X1 U2670 ( .A1(n2588), .A2(n2589), .ZN(n2704) );
  NAND2_X1 U2671 ( .A1(n2588), .A2(n2589), .ZN(n2701) );
  NAND2_X1 U2672 ( .A1(n2705), .A2(n2706), .ZN(n2589) );
  NAND2_X1 U2673 ( .A1(n2707), .A2(b_12_), .ZN(n2706) );
  NOR2_X1 U2674 ( .A1(n2708), .A2(n2214), .ZN(n2707) );
  NOR2_X1 U2675 ( .A1(n2630), .A2(n2632), .ZN(n2708) );
  NAND2_X1 U2676 ( .A1(n2630), .A2(n2632), .ZN(n2705) );
  NAND2_X1 U2677 ( .A1(n2709), .A2(n2710), .ZN(n2632) );
  NAND2_X1 U2678 ( .A1(n2628), .A2(n2711), .ZN(n2710) );
  NAND2_X1 U2679 ( .A1(n2627), .A2(n2626), .ZN(n2711) );
  NOR2_X1 U2680 ( .A1(n2211), .A2(n2212), .ZN(n2628) );
  OR2_X1 U2681 ( .A1(n2626), .A2(n2627), .ZN(n2709) );
  AND2_X1 U2682 ( .A1(n2712), .A2(n2713), .ZN(n2627) );
  NAND2_X1 U2683 ( .A1(n2622), .A2(n2714), .ZN(n2713) );
  NAND2_X1 U2684 ( .A1(n2624), .A2(n1994), .ZN(n2714) );
  INV_X1 U2685 ( .A(n2623), .ZN(n1994) );
  INV_X1 U2686 ( .A(n2715), .ZN(n2624) );
  XOR2_X1 U2687 ( .A(n2716), .B(n2717), .Z(n2622) );
  NOR2_X1 U2688 ( .A1(n2011), .A2(n2210), .ZN(n2717) );
  XOR2_X1 U2689 ( .A(n2718), .B(n2719), .Z(n2716) );
  NAND2_X1 U2690 ( .A1(n2623), .A2(n2715), .ZN(n2712) );
  NAND2_X1 U2691 ( .A1(n2720), .A2(n2721), .ZN(n2715) );
  NAND2_X1 U2692 ( .A1(n2722), .A2(b_12_), .ZN(n2721) );
  NOR2_X1 U2693 ( .A1(n2723), .A2(n2210), .ZN(n2722) );
  NOR2_X1 U2694 ( .A1(n2608), .A2(n2609), .ZN(n2723) );
  NAND2_X1 U2695 ( .A1(n2608), .A2(n2609), .ZN(n2720) );
  NAND2_X1 U2696 ( .A1(n2724), .A2(n2725), .ZN(n2609) );
  NAND2_X1 U2697 ( .A1(n2726), .A2(a_15_), .ZN(n2725) );
  NOR2_X1 U2698 ( .A1(n2727), .A2(n2213), .ZN(n2726) );
  NOR2_X1 U2699 ( .A1(n2380), .A2(n2011), .ZN(n2727) );
  NAND2_X1 U2700 ( .A1(n2728), .A2(a_14_), .ZN(n2724) );
  NOR2_X1 U2701 ( .A1(n2729), .A2(n2011), .ZN(n2728) );
  NOR2_X1 U2702 ( .A1(n2383), .A2(n2213), .ZN(n2729) );
  AND2_X1 U2703 ( .A1(n2730), .A2(b_12_), .ZN(n2608) );
  NOR2_X1 U2704 ( .A1(n2011), .A2(n2385), .ZN(n2730) );
  NOR2_X1 U2705 ( .A1(n2211), .A2(n2000), .ZN(n2623) );
  INV_X1 U2706 ( .A(b_12_), .ZN(n2211) );
  XOR2_X1 U2707 ( .A(n2731), .B(n2732), .Z(n2626) );
  NAND2_X1 U2708 ( .A1(n2733), .A2(n2734), .ZN(n2731) );
  XNOR2_X1 U2709 ( .A(n2735), .B(n2736), .ZN(n2630) );
  XNOR2_X1 U2710 ( .A(n2737), .B(n2006), .ZN(n2735) );
  XOR2_X1 U2711 ( .A(n2738), .B(n2739), .Z(n2588) );
  XNOR2_X1 U2712 ( .A(n2740), .B(n2741), .ZN(n2738) );
  NAND2_X1 U2713 ( .A1(a_10_), .A2(b_11_), .ZN(n2740) );
  XNOR2_X1 U2714 ( .A(n2742), .B(n2743), .ZN(n2638) );
  NAND2_X1 U2715 ( .A1(n2744), .A2(n2745), .ZN(n2742) );
  XOR2_X1 U2716 ( .A(n2746), .B(n2747), .Z(n2642) );
  XOR2_X1 U2717 ( .A(n2748), .B(n2749), .Z(n2746) );
  XOR2_X1 U2718 ( .A(n2750), .B(n2751), .Z(n2646) );
  XOR2_X1 U2719 ( .A(n2752), .B(n2753), .Z(n2750) );
  NOR2_X1 U2720 ( .A1(n2011), .A2(n2217), .ZN(n2753) );
  XNOR2_X1 U2721 ( .A(n2754), .B(n2755), .ZN(n2649) );
  XNOR2_X1 U2722 ( .A(n2756), .B(n2757), .ZN(n2754) );
  XNOR2_X1 U2723 ( .A(n2758), .B(n2759), .ZN(n2654) );
  XNOR2_X1 U2724 ( .A(n2760), .B(n2761), .ZN(n2758) );
  XOR2_X1 U2725 ( .A(n2762), .B(n2763), .Z(n2560) );
  XOR2_X1 U2726 ( .A(n2764), .B(n2765), .Z(n2762) );
  NOR2_X1 U2727 ( .A1(n2011), .A2(n2143), .ZN(n2765) );
  XOR2_X1 U2728 ( .A(n2766), .B(n2767), .Z(n2658) );
  NAND2_X1 U2729 ( .A1(n2768), .A2(n2769), .ZN(n2766) );
  XOR2_X1 U2730 ( .A(n2770), .B(n2771), .Z(n2662) );
  XOR2_X1 U2731 ( .A(n2772), .B(n2773), .Z(n2770) );
  NOR2_X1 U2732 ( .A1(n2011), .A2(n2319), .ZN(n2773) );
  XNOR2_X1 U2733 ( .A(n2774), .B(n2301), .ZN(n2290) );
  XOR2_X1 U2734 ( .A(n2775), .B(n2776), .Z(n2301) );
  XNOR2_X1 U2735 ( .A(n2777), .B(n2778), .ZN(n2776) );
  XOR2_X1 U2736 ( .A(n2304), .B(n2303), .Z(n2774) );
  NOR2_X1 U2737 ( .A1(n2228), .A2(n2011), .ZN(n2303) );
  NAND2_X1 U2738 ( .A1(n2779), .A2(n2780), .ZN(n2304) );
  NAND2_X1 U2739 ( .A1(n2781), .A2(a_1_), .ZN(n2780) );
  NOR2_X1 U2740 ( .A1(n2782), .A2(n2011), .ZN(n2781) );
  NOR2_X1 U2741 ( .A1(n2771), .A2(n2772), .ZN(n2782) );
  NAND2_X1 U2742 ( .A1(n2771), .A2(n2772), .ZN(n2779) );
  NAND2_X1 U2743 ( .A1(n2768), .A2(n2783), .ZN(n2772) );
  NAND2_X1 U2744 ( .A1(n2767), .A2(n2769), .ZN(n2783) );
  NAND2_X1 U2745 ( .A1(n2784), .A2(n2785), .ZN(n2769) );
  NAND2_X1 U2746 ( .A1(a_2_), .A2(b_11_), .ZN(n2785) );
  INV_X1 U2747 ( .A(n2786), .ZN(n2784) );
  XOR2_X1 U2748 ( .A(n2787), .B(n2788), .Z(n2767) );
  XOR2_X1 U2749 ( .A(n2789), .B(n2790), .Z(n2787) );
  NAND2_X1 U2750 ( .A1(a_2_), .A2(n2786), .ZN(n2768) );
  NAND2_X1 U2751 ( .A1(n2791), .A2(n2792), .ZN(n2786) );
  NAND2_X1 U2752 ( .A1(n2793), .A2(a_3_), .ZN(n2792) );
  NOR2_X1 U2753 ( .A1(n2794), .A2(n2011), .ZN(n2793) );
  NOR2_X1 U2754 ( .A1(n2763), .A2(n2764), .ZN(n2794) );
  NAND2_X1 U2755 ( .A1(n2763), .A2(n2764), .ZN(n2791) );
  NAND2_X1 U2756 ( .A1(n2795), .A2(n2796), .ZN(n2764) );
  NAND2_X1 U2757 ( .A1(n2761), .A2(n2797), .ZN(n2796) );
  NAND2_X1 U2758 ( .A1(n2760), .A2(n2759), .ZN(n2797) );
  NOR2_X1 U2759 ( .A1(n2011), .A2(n2220), .ZN(n2761) );
  OR2_X1 U2760 ( .A1(n2759), .A2(n2760), .ZN(n2795) );
  AND2_X1 U2761 ( .A1(n2798), .A2(n2799), .ZN(n2760) );
  NAND2_X1 U2762 ( .A1(n2757), .A2(n2800), .ZN(n2799) );
  NAND2_X1 U2763 ( .A1(n2756), .A2(n2755), .ZN(n2800) );
  NOR2_X1 U2764 ( .A1(n2108), .A2(n2011), .ZN(n2757) );
  OR2_X1 U2765 ( .A1(n2755), .A2(n2756), .ZN(n2798) );
  AND2_X1 U2766 ( .A1(n2801), .A2(n2802), .ZN(n2756) );
  NAND2_X1 U2767 ( .A1(n2803), .A2(a_6_), .ZN(n2802) );
  NOR2_X1 U2768 ( .A1(n2804), .A2(n2011), .ZN(n2803) );
  NOR2_X1 U2769 ( .A1(n2751), .A2(n2752), .ZN(n2804) );
  NAND2_X1 U2770 ( .A1(n2751), .A2(n2752), .ZN(n2801) );
  NAND2_X1 U2771 ( .A1(n2805), .A2(n2806), .ZN(n2752) );
  NAND2_X1 U2772 ( .A1(n2749), .A2(n2807), .ZN(n2806) );
  OR2_X1 U2773 ( .A1(n2748), .A2(n2747), .ZN(n2807) );
  NOR2_X1 U2774 ( .A1(n2073), .A2(n2011), .ZN(n2749) );
  NAND2_X1 U2775 ( .A1(n2747), .A2(n2748), .ZN(n2805) );
  NAND2_X1 U2776 ( .A1(n2744), .A2(n2808), .ZN(n2748) );
  NAND2_X1 U2777 ( .A1(n2743), .A2(n2745), .ZN(n2808) );
  NAND2_X1 U2778 ( .A1(n2809), .A2(n2810), .ZN(n2745) );
  NAND2_X1 U2779 ( .A1(a_8_), .A2(b_11_), .ZN(n2810) );
  INV_X1 U2780 ( .A(n2811), .ZN(n2809) );
  XOR2_X1 U2781 ( .A(n2812), .B(n2813), .Z(n2743) );
  XOR2_X1 U2782 ( .A(n2814), .B(n2815), .Z(n2812) );
  NOR2_X1 U2783 ( .A1(n2213), .A2(n2215), .ZN(n2815) );
  NAND2_X1 U2784 ( .A1(a_8_), .A2(n2811), .ZN(n2744) );
  NAND2_X1 U2785 ( .A1(n2816), .A2(n2817), .ZN(n2811) );
  NAND2_X1 U2786 ( .A1(n2818), .A2(a_9_), .ZN(n2817) );
  NOR2_X1 U2787 ( .A1(n2819), .A2(n2011), .ZN(n2818) );
  NOR2_X1 U2788 ( .A1(n2698), .A2(n2699), .ZN(n2819) );
  NAND2_X1 U2789 ( .A1(n2698), .A2(n2699), .ZN(n2816) );
  NAND2_X1 U2790 ( .A1(n2820), .A2(n2821), .ZN(n2699) );
  NAND2_X1 U2791 ( .A1(n2822), .A2(a_10_), .ZN(n2821) );
  NOR2_X1 U2792 ( .A1(n2823), .A2(n2011), .ZN(n2822) );
  NOR2_X1 U2793 ( .A1(n2739), .A2(n2741), .ZN(n2823) );
  NAND2_X1 U2794 ( .A1(n2739), .A2(n2741), .ZN(n2820) );
  NAND2_X1 U2795 ( .A1(n2824), .A2(n2825), .ZN(n2741) );
  NAND2_X1 U2796 ( .A1(n2006), .A2(n2826), .ZN(n2825) );
  NAND2_X1 U2797 ( .A1(n2737), .A2(n2736), .ZN(n2826) );
  NOR2_X1 U2798 ( .A1(n2212), .A2(n2011), .ZN(n2006) );
  OR2_X1 U2799 ( .A1(n2736), .A2(n2737), .ZN(n2824) );
  AND2_X1 U2800 ( .A1(n2733), .A2(n2827), .ZN(n2737) );
  NAND2_X1 U2801 ( .A1(n2732), .A2(n2734), .ZN(n2827) );
  NAND2_X1 U2802 ( .A1(n2828), .A2(n2829), .ZN(n2734) );
  NAND2_X1 U2803 ( .A1(a_12_), .A2(b_11_), .ZN(n2829) );
  INV_X1 U2804 ( .A(n2830), .ZN(n2828) );
  XOR2_X1 U2805 ( .A(n2831), .B(n2832), .Z(n2732) );
  NOR2_X1 U2806 ( .A1(n2213), .A2(n2210), .ZN(n2832) );
  XOR2_X1 U2807 ( .A(n2833), .B(n2834), .Z(n2831) );
  NAND2_X1 U2808 ( .A1(a_12_), .A2(n2830), .ZN(n2733) );
  NAND2_X1 U2809 ( .A1(n2835), .A2(n2836), .ZN(n2830) );
  NAND2_X1 U2810 ( .A1(n2837), .A2(a_13_), .ZN(n2836) );
  NOR2_X1 U2811 ( .A1(n2838), .A2(n2011), .ZN(n2837) );
  NOR2_X1 U2812 ( .A1(n2718), .A2(n2719), .ZN(n2838) );
  NAND2_X1 U2813 ( .A1(n2718), .A2(n2719), .ZN(n2835) );
  NAND2_X1 U2814 ( .A1(n2839), .A2(n2840), .ZN(n2719) );
  NAND2_X1 U2815 ( .A1(n2841), .A2(b_10_), .ZN(n2840) );
  NOR2_X1 U2816 ( .A1(n2842), .A2(n2499), .ZN(n2841) );
  NOR2_X1 U2817 ( .A1(n2383), .A2(n2040), .ZN(n2842) );
  NAND2_X1 U2818 ( .A1(n2843), .A2(a_15_), .ZN(n2839) );
  NOR2_X1 U2819 ( .A1(n2844), .A2(n2040), .ZN(n2843) );
  NOR2_X1 U2820 ( .A1(n2380), .A2(n2213), .ZN(n2844) );
  AND2_X1 U2821 ( .A1(n2845), .A2(n2209), .ZN(n2718) );
  NOR2_X1 U2822 ( .A1(n2011), .A2(n2213), .ZN(n2845) );
  INV_X1 U2823 ( .A(b_11_), .ZN(n2011) );
  XOR2_X1 U2824 ( .A(n2846), .B(n2847), .Z(n2736) );
  NAND2_X1 U2825 ( .A1(n2848), .A2(n2849), .ZN(n2846) );
  XNOR2_X1 U2826 ( .A(n2850), .B(n2851), .ZN(n2739) );
  XNOR2_X1 U2827 ( .A(n2852), .B(n2853), .ZN(n2850) );
  XOR2_X1 U2828 ( .A(n2854), .B(n2855), .Z(n2698) );
  XNOR2_X1 U2829 ( .A(n2856), .B(n2857), .ZN(n2854) );
  XNOR2_X1 U2830 ( .A(n2858), .B(n2859), .ZN(n2747) );
  NAND2_X1 U2831 ( .A1(n2860), .A2(n2861), .ZN(n2858) );
  XOR2_X1 U2832 ( .A(n2862), .B(n2863), .Z(n2751) );
  XOR2_X1 U2833 ( .A(n2864), .B(n2865), .Z(n2862) );
  XNOR2_X1 U2834 ( .A(n2866), .B(n2867), .ZN(n2755) );
  XOR2_X1 U2835 ( .A(n2868), .B(n2869), .Z(n2866) );
  NOR2_X1 U2836 ( .A1(n2213), .A2(n2217), .ZN(n2869) );
  XOR2_X1 U2837 ( .A(n2870), .B(n2871), .Z(n2759) );
  NAND2_X1 U2838 ( .A1(n2872), .A2(n2873), .ZN(n2870) );
  XOR2_X1 U2839 ( .A(n2874), .B(n2875), .Z(n2763) );
  XOR2_X1 U2840 ( .A(n2876), .B(n2877), .Z(n2874) );
  XNOR2_X1 U2841 ( .A(n2878), .B(n2879), .ZN(n2771) );
  XNOR2_X1 U2842 ( .A(n2880), .B(n2881), .ZN(n2878) );
  NAND2_X1 U2843 ( .A1(n2882), .A2(n2883), .ZN(n1916) );
  NAND2_X1 U2844 ( .A1(n2287), .A2(n2288), .ZN(n2883) );
  XNOR2_X1 U2845 ( .A(n2884), .B(n2885), .ZN(n2882) );
  NAND2_X1 U2846 ( .A1(n2886), .A2(n2887), .ZN(n1915) );
  XOR2_X1 U2847 ( .A(n2884), .B(n2885), .Z(n2887) );
  AND2_X1 U2848 ( .A1(n2288), .A2(n2287), .ZN(n2886) );
  XOR2_X1 U2849 ( .A(n2888), .B(n2889), .Z(n2287) );
  XOR2_X1 U2850 ( .A(n2890), .B(n2891), .Z(n2888) );
  NOR2_X1 U2851 ( .A1(n2040), .A2(n2228), .ZN(n2891) );
  NAND2_X1 U2852 ( .A1(n2297), .A2(n2892), .ZN(n2288) );
  NAND2_X1 U2853 ( .A1(n2296), .A2(n2298), .ZN(n2892) );
  NAND2_X1 U2854 ( .A1(n2893), .A2(n2894), .ZN(n2298) );
  NAND2_X1 U2855 ( .A1(a_0_), .A2(b_10_), .ZN(n2894) );
  INV_X1 U2856 ( .A(n2895), .ZN(n2893) );
  XNOR2_X1 U2857 ( .A(n2896), .B(n2897), .ZN(n2296) );
  XOR2_X1 U2858 ( .A(n2898), .B(n2899), .Z(n2897) );
  NAND2_X1 U2859 ( .A1(a_1_), .A2(b_9_), .ZN(n2899) );
  NAND2_X1 U2860 ( .A1(a_0_), .A2(n2895), .ZN(n2297) );
  NAND2_X1 U2861 ( .A1(n2900), .A2(n2901), .ZN(n2895) );
  NAND2_X1 U2862 ( .A1(n2778), .A2(n2902), .ZN(n2901) );
  OR2_X1 U2863 ( .A1(n2775), .A2(n2777), .ZN(n2902) );
  NOR2_X1 U2864 ( .A1(n2319), .A2(n2213), .ZN(n2778) );
  NAND2_X1 U2865 ( .A1(n2775), .A2(n2777), .ZN(n2900) );
  NAND2_X1 U2866 ( .A1(n2903), .A2(n2904), .ZN(n2777) );
  NAND2_X1 U2867 ( .A1(n2881), .A2(n2905), .ZN(n2904) );
  NAND2_X1 U2868 ( .A1(n2880), .A2(n2879), .ZN(n2905) );
  NOR2_X1 U2869 ( .A1(n2222), .A2(n2213), .ZN(n2881) );
  OR2_X1 U2870 ( .A1(n2879), .A2(n2880), .ZN(n2903) );
  AND2_X1 U2871 ( .A1(n2906), .A2(n2907), .ZN(n2880) );
  NAND2_X1 U2872 ( .A1(n2790), .A2(n2908), .ZN(n2907) );
  OR2_X1 U2873 ( .A1(n2788), .A2(n2789), .ZN(n2908) );
  NOR2_X1 U2874 ( .A1(n2143), .A2(n2213), .ZN(n2790) );
  NAND2_X1 U2875 ( .A1(n2788), .A2(n2789), .ZN(n2906) );
  NAND2_X1 U2876 ( .A1(n2909), .A2(n2910), .ZN(n2789) );
  NAND2_X1 U2877 ( .A1(n2877), .A2(n2911), .ZN(n2910) );
  OR2_X1 U2878 ( .A1(n2875), .A2(n2876), .ZN(n2911) );
  NOR2_X1 U2879 ( .A1(n2213), .A2(n2220), .ZN(n2877) );
  NAND2_X1 U2880 ( .A1(n2875), .A2(n2876), .ZN(n2909) );
  NAND2_X1 U2881 ( .A1(n2872), .A2(n2912), .ZN(n2876) );
  NAND2_X1 U2882 ( .A1(n2871), .A2(n2873), .ZN(n2912) );
  NAND2_X1 U2883 ( .A1(n2913), .A2(n2914), .ZN(n2873) );
  NAND2_X1 U2884 ( .A1(b_10_), .A2(a_5_), .ZN(n2914) );
  INV_X1 U2885 ( .A(n2915), .ZN(n2913) );
  XNOR2_X1 U2886 ( .A(n2916), .B(n2917), .ZN(n2871) );
  XOR2_X1 U2887 ( .A(n2918), .B(n2919), .Z(n2917) );
  NAND2_X1 U2888 ( .A1(a_6_), .A2(b_9_), .ZN(n2919) );
  NAND2_X1 U2889 ( .A1(a_5_), .A2(n2915), .ZN(n2872) );
  NAND2_X1 U2890 ( .A1(n2920), .A2(n2921), .ZN(n2915) );
  NAND2_X1 U2891 ( .A1(n2922), .A2(a_6_), .ZN(n2921) );
  NOR2_X1 U2892 ( .A1(n2923), .A2(n2213), .ZN(n2922) );
  NOR2_X1 U2893 ( .A1(n2868), .A2(n2867), .ZN(n2923) );
  NAND2_X1 U2894 ( .A1(n2867), .A2(n2868), .ZN(n2920) );
  NAND2_X1 U2895 ( .A1(n2924), .A2(n2925), .ZN(n2868) );
  NAND2_X1 U2896 ( .A1(n2865), .A2(n2926), .ZN(n2925) );
  OR2_X1 U2897 ( .A1(n2863), .A2(n2864), .ZN(n2926) );
  NOR2_X1 U2898 ( .A1(n2213), .A2(n2073), .ZN(n2865) );
  NAND2_X1 U2899 ( .A1(n2863), .A2(n2864), .ZN(n2924) );
  NAND2_X1 U2900 ( .A1(n2860), .A2(n2927), .ZN(n2864) );
  NAND2_X1 U2901 ( .A1(n2859), .A2(n2861), .ZN(n2927) );
  NAND2_X1 U2902 ( .A1(n2928), .A2(n2929), .ZN(n2861) );
  NAND2_X1 U2903 ( .A1(a_8_), .A2(b_10_), .ZN(n2929) );
  INV_X1 U2904 ( .A(n2930), .ZN(n2928) );
  XOR2_X1 U2905 ( .A(n2931), .B(n2932), .Z(n2859) );
  XNOR2_X1 U2906 ( .A(n2933), .B(n2194), .ZN(n2931) );
  INV_X1 U2907 ( .A(n2035), .ZN(n2194) );
  NAND2_X1 U2908 ( .A1(a_8_), .A2(n2930), .ZN(n2860) );
  NAND2_X1 U2909 ( .A1(n2934), .A2(n2935), .ZN(n2930) );
  NAND2_X1 U2910 ( .A1(n2936), .A2(a_9_), .ZN(n2935) );
  NOR2_X1 U2911 ( .A1(n2937), .A2(n2213), .ZN(n2936) );
  NOR2_X1 U2912 ( .A1(n2813), .A2(n2814), .ZN(n2937) );
  NAND2_X1 U2913 ( .A1(n2813), .A2(n2814), .ZN(n2934) );
  NAND2_X1 U2914 ( .A1(n2938), .A2(n2939), .ZN(n2814) );
  NAND2_X1 U2915 ( .A1(n2855), .A2(n2940), .ZN(n2939) );
  NAND2_X1 U2916 ( .A1(n2857), .A2(n2024), .ZN(n2940) );
  INV_X1 U2917 ( .A(n2856), .ZN(n2024) );
  INV_X1 U2918 ( .A(n2941), .ZN(n2857) );
  XNOR2_X1 U2919 ( .A(n2942), .B(n2943), .ZN(n2855) );
  XNOR2_X1 U2920 ( .A(n2944), .B(n2945), .ZN(n2942) );
  NAND2_X1 U2921 ( .A1(n2856), .A2(n2941), .ZN(n2938) );
  NAND2_X1 U2922 ( .A1(n2946), .A2(n2947), .ZN(n2941) );
  NAND2_X1 U2923 ( .A1(n2853), .A2(n2948), .ZN(n2947) );
  NAND2_X1 U2924 ( .A1(n2852), .A2(n2851), .ZN(n2948) );
  NOR2_X1 U2925 ( .A1(n2213), .A2(n2212), .ZN(n2853) );
  OR2_X1 U2926 ( .A1(n2851), .A2(n2852), .ZN(n2946) );
  AND2_X1 U2927 ( .A1(n2848), .A2(n2949), .ZN(n2852) );
  NAND2_X1 U2928 ( .A1(n2847), .A2(n2849), .ZN(n2949) );
  NAND2_X1 U2929 ( .A1(n2950), .A2(n2951), .ZN(n2849) );
  NAND2_X1 U2930 ( .A1(a_12_), .A2(b_10_), .ZN(n2951) );
  INV_X1 U2931 ( .A(n2952), .ZN(n2950) );
  XOR2_X1 U2932 ( .A(n2953), .B(n2954), .Z(n2847) );
  NOR2_X1 U2933 ( .A1(n2040), .A2(n2210), .ZN(n2954) );
  XOR2_X1 U2934 ( .A(n2955), .B(n2956), .Z(n2953) );
  NAND2_X1 U2935 ( .A1(a_12_), .A2(n2952), .ZN(n2848) );
  NAND2_X1 U2936 ( .A1(n2957), .A2(n2958), .ZN(n2952) );
  NAND2_X1 U2937 ( .A1(n2959), .A2(a_13_), .ZN(n2958) );
  NOR2_X1 U2938 ( .A1(n2960), .A2(n2213), .ZN(n2959) );
  NOR2_X1 U2939 ( .A1(n2833), .A2(n2834), .ZN(n2960) );
  NAND2_X1 U2940 ( .A1(n2833), .A2(n2834), .ZN(n2957) );
  NAND2_X1 U2941 ( .A1(n2961), .A2(n2962), .ZN(n2834) );
  NAND2_X1 U2942 ( .A1(n2963), .A2(b_8_), .ZN(n2962) );
  NOR2_X1 U2943 ( .A1(n2964), .A2(n2208), .ZN(n2963) );
  NOR2_X1 U2944 ( .A1(n2380), .A2(n2040), .ZN(n2964) );
  NAND2_X1 U2945 ( .A1(n2965), .A2(b_9_), .ZN(n2961) );
  NOR2_X1 U2946 ( .A1(n2966), .A2(n2499), .ZN(n2965) );
  NOR2_X1 U2947 ( .A1(n2383), .A2(n2967), .ZN(n2966) );
  AND2_X1 U2948 ( .A1(n2968), .A2(n2209), .ZN(n2833) );
  NOR2_X1 U2949 ( .A1(n2040), .A2(n2213), .ZN(n2968) );
  XOR2_X1 U2950 ( .A(n2969), .B(n2970), .Z(n2851) );
  NAND2_X1 U2951 ( .A1(n2971), .A2(n2972), .ZN(n2969) );
  NOR2_X1 U2952 ( .A1(n2214), .A2(n2213), .ZN(n2856) );
  INV_X1 U2953 ( .A(b_10_), .ZN(n2213) );
  XOR2_X1 U2954 ( .A(n2973), .B(n2974), .Z(n2813) );
  XNOR2_X1 U2955 ( .A(n2975), .B(n2976), .ZN(n2973) );
  NAND2_X1 U2956 ( .A1(a_10_), .A2(b_9_), .ZN(n2975) );
  XNOR2_X1 U2957 ( .A(n2977), .B(n2978), .ZN(n2863) );
  NAND2_X1 U2958 ( .A1(n2979), .A2(n2980), .ZN(n2977) );
  XNOR2_X1 U2959 ( .A(n2981), .B(n2982), .ZN(n2867) );
  XNOR2_X1 U2960 ( .A(n2983), .B(n2984), .ZN(n2981) );
  XNOR2_X1 U2961 ( .A(n2985), .B(n2986), .ZN(n2875) );
  NAND2_X1 U2962 ( .A1(n2987), .A2(n2988), .ZN(n2985) );
  XNOR2_X1 U2963 ( .A(n2989), .B(n2990), .ZN(n2788) );
  XOR2_X1 U2964 ( .A(n2991), .B(n2992), .Z(n2990) );
  NAND2_X1 U2965 ( .A1(b_9_), .A2(a_4_), .ZN(n2992) );
  XNOR2_X1 U2966 ( .A(n2993), .B(n2994), .ZN(n2879) );
  XOR2_X1 U2967 ( .A(n2995), .B(n2996), .Z(n2993) );
  NOR2_X1 U2968 ( .A1(n2040), .A2(n2143), .ZN(n2996) );
  XOR2_X1 U2969 ( .A(n2997), .B(n2998), .Z(n2775) );
  XOR2_X1 U2970 ( .A(n2999), .B(n3000), .Z(n2997) );
  NOR2_X1 U2971 ( .A1(n2040), .A2(n2222), .ZN(n3000) );
  NAND2_X1 U2972 ( .A1(n3001), .A2(n3002), .ZN(n1921) );
  NAND2_X1 U2973 ( .A1(n2885), .A2(n2884), .ZN(n3002) );
  XNOR2_X1 U2974 ( .A(n3003), .B(n3004), .ZN(n3001) );
  NAND2_X1 U2975 ( .A1(n3005), .A2(n3006), .ZN(n1920) );
  XNOR2_X1 U2976 ( .A(n3007), .B(n3003), .ZN(n3006) );
  AND2_X1 U2977 ( .A1(n2884), .A2(n2885), .ZN(n3005) );
  XOR2_X1 U2978 ( .A(n3008), .B(n3009), .Z(n2885) );
  XOR2_X1 U2979 ( .A(n3010), .B(n3011), .Z(n3009) );
  NAND2_X1 U2980 ( .A1(n3012), .A2(n3013), .ZN(n2884) );
  NAND2_X1 U2981 ( .A1(n3014), .A2(a_0_), .ZN(n3013) );
  NOR2_X1 U2982 ( .A1(n3015), .A2(n2040), .ZN(n3014) );
  NOR2_X1 U2983 ( .A1(n2890), .A2(n2889), .ZN(n3015) );
  NAND2_X1 U2984 ( .A1(n2889), .A2(n2890), .ZN(n3012) );
  NAND2_X1 U2985 ( .A1(n3016), .A2(n3017), .ZN(n2890) );
  NAND2_X1 U2986 ( .A1(n3018), .A2(a_1_), .ZN(n3017) );
  NOR2_X1 U2987 ( .A1(n3019), .A2(n2040), .ZN(n3018) );
  NOR2_X1 U2988 ( .A1(n2896), .A2(n2898), .ZN(n3019) );
  NAND2_X1 U2989 ( .A1(n2896), .A2(n2898), .ZN(n3016) );
  NAND2_X1 U2990 ( .A1(n3020), .A2(n3021), .ZN(n2898) );
  NAND2_X1 U2991 ( .A1(n3022), .A2(a_2_), .ZN(n3021) );
  NOR2_X1 U2992 ( .A1(n3023), .A2(n2040), .ZN(n3022) );
  NOR2_X1 U2993 ( .A1(n2998), .A2(n2999), .ZN(n3023) );
  NAND2_X1 U2994 ( .A1(n2998), .A2(n2999), .ZN(n3020) );
  NAND2_X1 U2995 ( .A1(n3024), .A2(n3025), .ZN(n2999) );
  NAND2_X1 U2996 ( .A1(n3026), .A2(a_3_), .ZN(n3025) );
  NOR2_X1 U2997 ( .A1(n3027), .A2(n2040), .ZN(n3026) );
  NOR2_X1 U2998 ( .A1(n2995), .A2(n2994), .ZN(n3027) );
  NAND2_X1 U2999 ( .A1(n2994), .A2(n2995), .ZN(n3024) );
  NAND2_X1 U3000 ( .A1(n3028), .A2(n3029), .ZN(n2995) );
  NAND2_X1 U3001 ( .A1(n3030), .A2(b_9_), .ZN(n3029) );
  NOR2_X1 U3002 ( .A1(n3031), .A2(n2220), .ZN(n3030) );
  NOR2_X1 U3003 ( .A1(n2989), .A2(n2991), .ZN(n3031) );
  NAND2_X1 U3004 ( .A1(n2989), .A2(n2991), .ZN(n3028) );
  NAND2_X1 U3005 ( .A1(n2987), .A2(n3032), .ZN(n2991) );
  NAND2_X1 U3006 ( .A1(n2986), .A2(n2988), .ZN(n3032) );
  NAND2_X1 U3007 ( .A1(n3033), .A2(n3034), .ZN(n2988) );
  NAND2_X1 U3008 ( .A1(b_9_), .A2(a_5_), .ZN(n3034) );
  INV_X1 U3009 ( .A(n3035), .ZN(n3033) );
  XNOR2_X1 U3010 ( .A(n3036), .B(n3037), .ZN(n2986) );
  XNOR2_X1 U3011 ( .A(n3038), .B(n3039), .ZN(n3037) );
  NAND2_X1 U3012 ( .A1(a_5_), .A2(n3035), .ZN(n2987) );
  NAND2_X1 U3013 ( .A1(n3040), .A2(n3041), .ZN(n3035) );
  NAND2_X1 U3014 ( .A1(n3042), .A2(a_6_), .ZN(n3041) );
  NOR2_X1 U3015 ( .A1(n3043), .A2(n2040), .ZN(n3042) );
  NOR2_X1 U3016 ( .A1(n2918), .A2(n2916), .ZN(n3043) );
  NAND2_X1 U3017 ( .A1(n2916), .A2(n2918), .ZN(n3040) );
  NAND2_X1 U3018 ( .A1(n3044), .A2(n3045), .ZN(n2918) );
  NAND2_X1 U3019 ( .A1(n2984), .A2(n3046), .ZN(n3045) );
  NAND2_X1 U3020 ( .A1(n2983), .A2(n2982), .ZN(n3046) );
  NOR2_X1 U3021 ( .A1(n2040), .A2(n2073), .ZN(n2984) );
  OR2_X1 U3022 ( .A1(n2982), .A2(n2983), .ZN(n3044) );
  AND2_X1 U3023 ( .A1(n2979), .A2(n3047), .ZN(n2983) );
  NAND2_X1 U3024 ( .A1(n2978), .A2(n2980), .ZN(n3047) );
  NAND2_X1 U3025 ( .A1(n3048), .A2(n3049), .ZN(n2980) );
  NAND2_X1 U3026 ( .A1(a_8_), .A2(b_9_), .ZN(n3049) );
  INV_X1 U3027 ( .A(n3050), .ZN(n3048) );
  XNOR2_X1 U3028 ( .A(n3051), .B(n3052), .ZN(n2978) );
  XOR2_X1 U3029 ( .A(n3053), .B(n3054), .Z(n3052) );
  NAND2_X1 U3030 ( .A1(a_9_), .A2(b_8_), .ZN(n3054) );
  NAND2_X1 U3031 ( .A1(a_8_), .A2(n3050), .ZN(n2979) );
  NAND2_X1 U3032 ( .A1(n3055), .A2(n3056), .ZN(n3050) );
  NAND2_X1 U3033 ( .A1(n2932), .A2(n3057), .ZN(n3056) );
  OR2_X1 U3034 ( .A1(n2933), .A2(n2035), .ZN(n3057) );
  XOR2_X1 U3035 ( .A(n3058), .B(n3059), .Z(n2932) );
  XNOR2_X1 U3036 ( .A(n3060), .B(n3061), .ZN(n3058) );
  NAND2_X1 U3037 ( .A1(a_10_), .A2(b_8_), .ZN(n3060) );
  NAND2_X1 U3038 ( .A1(n2035), .A2(n2933), .ZN(n3055) );
  NAND2_X1 U3039 ( .A1(n3062), .A2(n3063), .ZN(n2933) );
  NAND2_X1 U3040 ( .A1(n3064), .A2(a_10_), .ZN(n3063) );
  NOR2_X1 U3041 ( .A1(n3065), .A2(n2040), .ZN(n3064) );
  NOR2_X1 U3042 ( .A1(n2976), .A2(n2974), .ZN(n3065) );
  NAND2_X1 U3043 ( .A1(n2974), .A2(n2976), .ZN(n3062) );
  NAND2_X1 U3044 ( .A1(n3066), .A2(n3067), .ZN(n2976) );
  NAND2_X1 U3045 ( .A1(n2945), .A2(n3068), .ZN(n3067) );
  NAND2_X1 U3046 ( .A1(n2944), .A2(n2943), .ZN(n3068) );
  NOR2_X1 U3047 ( .A1(n2040), .A2(n2212), .ZN(n2945) );
  OR2_X1 U3048 ( .A1(n2943), .A2(n2944), .ZN(n3066) );
  AND2_X1 U3049 ( .A1(n2971), .A2(n3069), .ZN(n2944) );
  NAND2_X1 U3050 ( .A1(n2970), .A2(n2972), .ZN(n3069) );
  NAND2_X1 U3051 ( .A1(n3070), .A2(n3071), .ZN(n2972) );
  NAND2_X1 U3052 ( .A1(a_12_), .A2(b_9_), .ZN(n3071) );
  INV_X1 U3053 ( .A(n3072), .ZN(n3070) );
  XOR2_X1 U3054 ( .A(n3073), .B(n3074), .Z(n2970) );
  NOR2_X1 U3055 ( .A1(n2210), .A2(n2967), .ZN(n3074) );
  XOR2_X1 U3056 ( .A(n3075), .B(n3076), .Z(n3073) );
  NAND2_X1 U3057 ( .A1(a_12_), .A2(n3072), .ZN(n2971) );
  NAND2_X1 U3058 ( .A1(n3077), .A2(n3078), .ZN(n3072) );
  NAND2_X1 U3059 ( .A1(n3079), .A2(a_13_), .ZN(n3078) );
  NOR2_X1 U3060 ( .A1(n3080), .A2(n2040), .ZN(n3079) );
  NOR2_X1 U3061 ( .A1(n2955), .A2(n2956), .ZN(n3080) );
  NAND2_X1 U3062 ( .A1(n2955), .A2(n2956), .ZN(n3077) );
  NAND2_X1 U3063 ( .A1(n3081), .A2(n3082), .ZN(n2956) );
  NAND2_X1 U3064 ( .A1(n3083), .A2(b_7_), .ZN(n3082) );
  NOR2_X1 U3065 ( .A1(n3084), .A2(n2208), .ZN(n3083) );
  NOR2_X1 U3066 ( .A1(n2380), .A2(n2967), .ZN(n3084) );
  NAND2_X1 U3067 ( .A1(n3085), .A2(b_8_), .ZN(n3081) );
  NOR2_X1 U3068 ( .A1(n3086), .A2(n2499), .ZN(n3085) );
  NOR2_X1 U3069 ( .A1(n2383), .A2(n2070), .ZN(n3086) );
  AND2_X1 U3070 ( .A1(n3087), .A2(b_8_), .ZN(n2955) );
  NOR2_X1 U3071 ( .A1(n2040), .A2(n2385), .ZN(n3087) );
  XOR2_X1 U3072 ( .A(n3088), .B(n3089), .Z(n2943) );
  NAND2_X1 U3073 ( .A1(n3090), .A2(n3091), .ZN(n3088) );
  XNOR2_X1 U3074 ( .A(n3092), .B(n3093), .ZN(n2974) );
  XNOR2_X1 U3075 ( .A(n3094), .B(n3095), .ZN(n3092) );
  NOR2_X1 U3076 ( .A1(n2215), .A2(n2040), .ZN(n2035) );
  INV_X1 U3077 ( .A(b_9_), .ZN(n2040) );
  XOR2_X1 U3078 ( .A(n3096), .B(n3097), .Z(n2982) );
  XNOR2_X1 U3079 ( .A(n3098), .B(n2053), .ZN(n3097) );
  XOR2_X1 U3080 ( .A(n3099), .B(n3100), .Z(n2916) );
  XOR2_X1 U3081 ( .A(n3101), .B(n3102), .Z(n3099) );
  NOR2_X1 U3082 ( .A1(n2073), .A2(n2967), .ZN(n3102) );
  XOR2_X1 U3083 ( .A(n3103), .B(n3104), .Z(n2989) );
  XOR2_X1 U3084 ( .A(n3105), .B(n3106), .Z(n3103) );
  NOR2_X1 U3085 ( .A1(n2108), .A2(n2967), .ZN(n3106) );
  XNOR2_X1 U3086 ( .A(n3107), .B(n3108), .ZN(n2994) );
  XOR2_X1 U3087 ( .A(n3109), .B(n3110), .Z(n3108) );
  NAND2_X1 U3088 ( .A1(b_8_), .A2(a_4_), .ZN(n3110) );
  XNOR2_X1 U3089 ( .A(n3111), .B(n3112), .ZN(n2998) );
  XNOR2_X1 U3090 ( .A(n3113), .B(n3114), .ZN(n3111) );
  XOR2_X1 U3091 ( .A(n3115), .B(n3116), .Z(n2896) );
  XOR2_X1 U3092 ( .A(n3117), .B(n3118), .Z(n3115) );
  XNOR2_X1 U3093 ( .A(n3119), .B(n3120), .ZN(n2889) );
  XNOR2_X1 U3094 ( .A(n3121), .B(n3122), .ZN(n3119) );
  NAND2_X1 U3095 ( .A1(n3123), .A2(n3124), .ZN(n1926) );
  NAND2_X1 U3096 ( .A1(n3125), .A2(n3007), .ZN(n3124) );
  NAND2_X1 U3097 ( .A1(n3126), .A2(n3125), .ZN(n1925) );
  INV_X1 U3098 ( .A(n3003), .ZN(n3125) );
  XOR2_X1 U3099 ( .A(n3127), .B(n3128), .Z(n3003) );
  XOR2_X1 U3100 ( .A(n3129), .B(n3130), .Z(n3128) );
  NAND2_X1 U3101 ( .A1(a_0_), .A2(b_7_), .ZN(n3130) );
  NOR2_X1 U3102 ( .A1(n3004), .A2(n3123), .ZN(n3126) );
  XNOR2_X1 U3103 ( .A(n3131), .B(n3132), .ZN(n3123) );
  INV_X1 U3104 ( .A(n3007), .ZN(n3004) );
  NAND2_X1 U3105 ( .A1(n3133), .A2(n3134), .ZN(n3007) );
  NAND2_X1 U3106 ( .A1(n3011), .A2(n3135), .ZN(n3134) );
  NAND2_X1 U3107 ( .A1(n3010), .A2(n3008), .ZN(n3135) );
  NOR2_X1 U3108 ( .A1(n2228), .A2(n2967), .ZN(n3011) );
  OR2_X1 U3109 ( .A1(n3008), .A2(n3010), .ZN(n3133) );
  AND2_X1 U3110 ( .A1(n3136), .A2(n3137), .ZN(n3010) );
  NAND2_X1 U3111 ( .A1(n3122), .A2(n3138), .ZN(n3137) );
  NAND2_X1 U3112 ( .A1(n3121), .A2(n3120), .ZN(n3138) );
  NOR2_X1 U3113 ( .A1(n2319), .A2(n2967), .ZN(n3122) );
  OR2_X1 U3114 ( .A1(n3120), .A2(n3121), .ZN(n3136) );
  AND2_X1 U3115 ( .A1(n3139), .A2(n3140), .ZN(n3121) );
  NAND2_X1 U3116 ( .A1(n3118), .A2(n3141), .ZN(n3140) );
  OR2_X1 U3117 ( .A1(n3116), .A2(n3117), .ZN(n3141) );
  NOR2_X1 U3118 ( .A1(n2222), .A2(n2967), .ZN(n3118) );
  NAND2_X1 U3119 ( .A1(n3116), .A2(n3117), .ZN(n3139) );
  NAND2_X1 U3120 ( .A1(n3142), .A2(n3143), .ZN(n3117) );
  NAND2_X1 U3121 ( .A1(n3114), .A2(n3144), .ZN(n3143) );
  NAND2_X1 U3122 ( .A1(n3112), .A2(n3113), .ZN(n3144) );
  NOR2_X1 U3123 ( .A1(n2143), .A2(n2967), .ZN(n3114) );
  OR2_X1 U3124 ( .A1(n3112), .A2(n3113), .ZN(n3142) );
  AND2_X1 U3125 ( .A1(n3145), .A2(n3146), .ZN(n3113) );
  NAND2_X1 U3126 ( .A1(n3147), .A2(b_8_), .ZN(n3146) );
  NOR2_X1 U3127 ( .A1(n3148), .A2(n2220), .ZN(n3147) );
  NOR2_X1 U3128 ( .A1(n3107), .A2(n3109), .ZN(n3148) );
  NAND2_X1 U3129 ( .A1(n3107), .A2(n3109), .ZN(n3145) );
  NAND2_X1 U3130 ( .A1(n3149), .A2(n3150), .ZN(n3109) );
  NAND2_X1 U3131 ( .A1(n3151), .A2(b_8_), .ZN(n3150) );
  NOR2_X1 U3132 ( .A1(n3152), .A2(n2108), .ZN(n3151) );
  NOR2_X1 U3133 ( .A1(n3105), .A2(n3104), .ZN(n3152) );
  NAND2_X1 U3134 ( .A1(n3104), .A2(n3105), .ZN(n3149) );
  NAND2_X1 U3135 ( .A1(n3153), .A2(n3154), .ZN(n3105) );
  NAND2_X1 U3136 ( .A1(n3039), .A2(n3155), .ZN(n3154) );
  OR2_X1 U3137 ( .A1(n3038), .A2(n3036), .ZN(n3155) );
  NOR2_X1 U3138 ( .A1(n2217), .A2(n2967), .ZN(n3039) );
  NAND2_X1 U3139 ( .A1(n3036), .A2(n3038), .ZN(n3153) );
  NAND2_X1 U3140 ( .A1(n3156), .A2(n3157), .ZN(n3038) );
  NAND2_X1 U3141 ( .A1(n3158), .A2(b_8_), .ZN(n3157) );
  NOR2_X1 U3142 ( .A1(n3159), .A2(n2073), .ZN(n3158) );
  NOR2_X1 U3143 ( .A1(n3100), .A2(n3101), .ZN(n3159) );
  NAND2_X1 U3144 ( .A1(n3100), .A2(n3101), .ZN(n3156) );
  NAND2_X1 U3145 ( .A1(n3160), .A2(n3161), .ZN(n3101) );
  NAND2_X1 U3146 ( .A1(n3096), .A2(n3162), .ZN(n3161) );
  OR2_X1 U3147 ( .A1(n3098), .A2(n2053), .ZN(n3162) );
  XNOR2_X1 U3148 ( .A(n3163), .B(n3164), .ZN(n3096) );
  XOR2_X1 U3149 ( .A(n3165), .B(n3166), .Z(n3164) );
  NAND2_X1 U3150 ( .A1(a_9_), .A2(b_7_), .ZN(n3166) );
  NAND2_X1 U3151 ( .A1(n2053), .A2(n3098), .ZN(n3160) );
  NAND2_X1 U3152 ( .A1(n3167), .A2(n3168), .ZN(n3098) );
  NAND2_X1 U3153 ( .A1(n3169), .A2(a_9_), .ZN(n3168) );
  NOR2_X1 U3154 ( .A1(n3170), .A2(n2967), .ZN(n3169) );
  NOR2_X1 U3155 ( .A1(n3051), .A2(n3053), .ZN(n3170) );
  NAND2_X1 U3156 ( .A1(n3051), .A2(n3053), .ZN(n3167) );
  NAND2_X1 U3157 ( .A1(n3171), .A2(n3172), .ZN(n3053) );
  NAND2_X1 U3158 ( .A1(n3173), .A2(a_10_), .ZN(n3172) );
  NOR2_X1 U3159 ( .A1(n3174), .A2(n2967), .ZN(n3173) );
  NOR2_X1 U3160 ( .A1(n3061), .A2(n3059), .ZN(n3174) );
  NAND2_X1 U3161 ( .A1(n3059), .A2(n3061), .ZN(n3171) );
  NAND2_X1 U3162 ( .A1(n3175), .A2(n3176), .ZN(n3061) );
  NAND2_X1 U3163 ( .A1(n3095), .A2(n3177), .ZN(n3176) );
  NAND2_X1 U3164 ( .A1(n3094), .A2(n3093), .ZN(n3177) );
  NOR2_X1 U3165 ( .A1(n2967), .A2(n2212), .ZN(n3095) );
  OR2_X1 U3166 ( .A1(n3093), .A2(n3094), .ZN(n3175) );
  AND2_X1 U3167 ( .A1(n3090), .A2(n3178), .ZN(n3094) );
  NAND2_X1 U3168 ( .A1(n3089), .A2(n3091), .ZN(n3178) );
  NAND2_X1 U3169 ( .A1(n3179), .A2(n3180), .ZN(n3091) );
  NAND2_X1 U3170 ( .A1(b_8_), .A2(a_12_), .ZN(n3180) );
  INV_X1 U3171 ( .A(n3181), .ZN(n3179) );
  XOR2_X1 U3172 ( .A(n3182), .B(n3183), .Z(n3089) );
  NOR2_X1 U3173 ( .A1(n2210), .A2(n2070), .ZN(n3183) );
  XOR2_X1 U3174 ( .A(n3184), .B(n3185), .Z(n3182) );
  NAND2_X1 U3175 ( .A1(a_12_), .A2(n3181), .ZN(n3090) );
  NAND2_X1 U3176 ( .A1(n3186), .A2(n3187), .ZN(n3181) );
  NAND2_X1 U3177 ( .A1(n3188), .A2(b_8_), .ZN(n3187) );
  NOR2_X1 U3178 ( .A1(n3189), .A2(n2210), .ZN(n3188) );
  NOR2_X1 U3179 ( .A1(n3075), .A2(n3076), .ZN(n3189) );
  NAND2_X1 U3180 ( .A1(n3075), .A2(n3076), .ZN(n3186) );
  NAND2_X1 U3181 ( .A1(n3190), .A2(n3191), .ZN(n3076) );
  NAND2_X1 U3182 ( .A1(n3192), .A2(b_6_), .ZN(n3191) );
  NOR2_X1 U3183 ( .A1(n3193), .A2(n2208), .ZN(n3192) );
  NOR2_X1 U3184 ( .A1(n2380), .A2(n2070), .ZN(n3193) );
  NAND2_X1 U3185 ( .A1(n3194), .A2(b_7_), .ZN(n3190) );
  NOR2_X1 U3186 ( .A1(n3195), .A2(n2499), .ZN(n3194) );
  NOR2_X1 U3187 ( .A1(n2383), .A2(n2216), .ZN(n3195) );
  AND2_X1 U3188 ( .A1(n3196), .A2(b_7_), .ZN(n3075) );
  NOR2_X1 U3189 ( .A1(n2385), .A2(n2967), .ZN(n3196) );
  XOR2_X1 U3190 ( .A(n3197), .B(n3198), .Z(n3093) );
  NAND2_X1 U3191 ( .A1(n3199), .A2(n3200), .ZN(n3197) );
  XNOR2_X1 U3192 ( .A(n3201), .B(n3202), .ZN(n3059) );
  XNOR2_X1 U3193 ( .A(n3203), .B(n3204), .ZN(n3201) );
  XOR2_X1 U3194 ( .A(n3205), .B(n3206), .Z(n3051) );
  XNOR2_X1 U3195 ( .A(n3207), .B(n3208), .ZN(n3205) );
  NAND2_X1 U3196 ( .A1(a_10_), .A2(b_7_), .ZN(n3207) );
  NOR2_X1 U3197 ( .A1(n2059), .A2(n2967), .ZN(n2053) );
  INV_X1 U3198 ( .A(b_8_), .ZN(n2967) );
  XNOR2_X1 U3199 ( .A(n3209), .B(n3210), .ZN(n3100) );
  XNOR2_X1 U3200 ( .A(n3211), .B(n3212), .ZN(n3210) );
  XOR2_X1 U3201 ( .A(n3213), .B(n3214), .Z(n3036) );
  XNOR2_X1 U3202 ( .A(n3215), .B(n2190), .ZN(n3213) );
  INV_X1 U3203 ( .A(n2065), .ZN(n2190) );
  XNOR2_X1 U3204 ( .A(n3216), .B(n3217), .ZN(n3104) );
  XOR2_X1 U3205 ( .A(n3218), .B(n3219), .Z(n3217) );
  NAND2_X1 U3206 ( .A1(a_6_), .A2(b_7_), .ZN(n3219) );
  XOR2_X1 U3207 ( .A(n3220), .B(n3221), .Z(n3107) );
  XOR2_X1 U3208 ( .A(n3222), .B(n3223), .Z(n3220) );
  NOR2_X1 U3209 ( .A1(n2108), .A2(n2070), .ZN(n3223) );
  XOR2_X1 U3210 ( .A(n3224), .B(n3225), .Z(n3112) );
  XOR2_X1 U3211 ( .A(n3226), .B(n3227), .Z(n3225) );
  NAND2_X1 U3212 ( .A1(b_7_), .A2(a_4_), .ZN(n3227) );
  XNOR2_X1 U3213 ( .A(n3228), .B(n3229), .ZN(n3116) );
  XOR2_X1 U3214 ( .A(n3230), .B(n3231), .Z(n3229) );
  NAND2_X1 U3215 ( .A1(a_3_), .A2(b_7_), .ZN(n3231) );
  XNOR2_X1 U3216 ( .A(n3232), .B(n3233), .ZN(n3120) );
  XOR2_X1 U3217 ( .A(n3234), .B(n3235), .Z(n3232) );
  NOR2_X1 U3218 ( .A1(n2070), .A2(n2222), .ZN(n3235) );
  XNOR2_X1 U3219 ( .A(n3236), .B(n3237), .ZN(n3008) );
  XOR2_X1 U3220 ( .A(n3238), .B(n3239), .Z(n3236) );
  NOR2_X1 U3221 ( .A1(n2070), .A2(n2319), .ZN(n3239) );
  NAND2_X1 U3222 ( .A1(n3240), .A2(n3241), .ZN(n1931) );
  NAND2_X1 U3223 ( .A1(n3131), .A2(n3132), .ZN(n3241) );
  NAND2_X1 U3224 ( .A1(n3242), .A2(n3131), .ZN(n1930) );
  XOR2_X1 U3225 ( .A(n3243), .B(n3244), .Z(n3131) );
  XOR2_X1 U3226 ( .A(n3245), .B(n3246), .Z(n3243) );
  NOR2_X1 U3227 ( .A1(n2216), .A2(n2228), .ZN(n3246) );
  NOR2_X1 U3228 ( .A1(n3247), .A2(n3240), .ZN(n3242) );
  XNOR2_X1 U3229 ( .A(n3248), .B(n3249), .ZN(n3240) );
  INV_X1 U3230 ( .A(n3132), .ZN(n3247) );
  NAND2_X1 U3231 ( .A1(n3250), .A2(n3251), .ZN(n3132) );
  NAND2_X1 U3232 ( .A1(n3252), .A2(a_0_), .ZN(n3251) );
  NOR2_X1 U3233 ( .A1(n3253), .A2(n2070), .ZN(n3252) );
  NOR2_X1 U3234 ( .A1(n3129), .A2(n3127), .ZN(n3253) );
  NAND2_X1 U3235 ( .A1(n3127), .A2(n3129), .ZN(n3250) );
  NAND2_X1 U3236 ( .A1(n3254), .A2(n3255), .ZN(n3129) );
  NAND2_X1 U3237 ( .A1(n3256), .A2(a_1_), .ZN(n3255) );
  NOR2_X1 U3238 ( .A1(n3257), .A2(n2070), .ZN(n3256) );
  NOR2_X1 U3239 ( .A1(n3238), .A2(n3237), .ZN(n3257) );
  NAND2_X1 U3240 ( .A1(n3237), .A2(n3238), .ZN(n3254) );
  NAND2_X1 U3241 ( .A1(n3258), .A2(n3259), .ZN(n3238) );
  NAND2_X1 U3242 ( .A1(n3260), .A2(a_2_), .ZN(n3259) );
  NOR2_X1 U3243 ( .A1(n3261), .A2(n2070), .ZN(n3260) );
  NOR2_X1 U3244 ( .A1(n3234), .A2(n3233), .ZN(n3261) );
  NAND2_X1 U3245 ( .A1(n3233), .A2(n3234), .ZN(n3258) );
  NAND2_X1 U3246 ( .A1(n3262), .A2(n3263), .ZN(n3234) );
  NAND2_X1 U3247 ( .A1(n3264), .A2(a_3_), .ZN(n3263) );
  NOR2_X1 U3248 ( .A1(n3265), .A2(n2070), .ZN(n3264) );
  NOR2_X1 U3249 ( .A1(n3228), .A2(n3230), .ZN(n3265) );
  NAND2_X1 U3250 ( .A1(n3228), .A2(n3230), .ZN(n3262) );
  NAND2_X1 U3251 ( .A1(n3266), .A2(n3267), .ZN(n3230) );
  NAND2_X1 U3252 ( .A1(n3268), .A2(b_7_), .ZN(n3267) );
  NOR2_X1 U3253 ( .A1(n3269), .A2(n2220), .ZN(n3268) );
  NOR2_X1 U3254 ( .A1(n3224), .A2(n3226), .ZN(n3269) );
  NAND2_X1 U3255 ( .A1(n3224), .A2(n3226), .ZN(n3266) );
  NAND2_X1 U3256 ( .A1(n3270), .A2(n3271), .ZN(n3226) );
  NAND2_X1 U3257 ( .A1(n3272), .A2(b_7_), .ZN(n3271) );
  NOR2_X1 U3258 ( .A1(n3273), .A2(n2108), .ZN(n3272) );
  NOR2_X1 U3259 ( .A1(n3222), .A2(n3221), .ZN(n3273) );
  NAND2_X1 U3260 ( .A1(n3221), .A2(n3222), .ZN(n3270) );
  NAND2_X1 U3261 ( .A1(n3274), .A2(n3275), .ZN(n3222) );
  NAND2_X1 U3262 ( .A1(n3276), .A2(a_6_), .ZN(n3275) );
  NOR2_X1 U3263 ( .A1(n3277), .A2(n2070), .ZN(n3276) );
  NOR2_X1 U3264 ( .A1(n3216), .A2(n3218), .ZN(n3277) );
  NAND2_X1 U3265 ( .A1(n3216), .A2(n3218), .ZN(n3274) );
  NAND2_X1 U3266 ( .A1(n3278), .A2(n3279), .ZN(n3218) );
  NAND2_X1 U3267 ( .A1(n3214), .A2(n3280), .ZN(n3279) );
  OR2_X1 U3268 ( .A1(n3215), .A2(n2065), .ZN(n3280) );
  XNOR2_X1 U3269 ( .A(n3281), .B(n3282), .ZN(n3214) );
  NAND2_X1 U3270 ( .A1(n3283), .A2(n3284), .ZN(n3281) );
  NAND2_X1 U3271 ( .A1(n2065), .A2(n3215), .ZN(n3278) );
  NAND2_X1 U3272 ( .A1(n3285), .A2(n3286), .ZN(n3215) );
  NAND2_X1 U3273 ( .A1(n3212), .A2(n3287), .ZN(n3286) );
  OR2_X1 U3274 ( .A1(n3209), .A2(n3211), .ZN(n3287) );
  NOR2_X1 U3275 ( .A1(n2059), .A2(n2070), .ZN(n3212) );
  NAND2_X1 U3276 ( .A1(n3209), .A2(n3211), .ZN(n3285) );
  NAND2_X1 U3277 ( .A1(n3288), .A2(n3289), .ZN(n3211) );
  NAND2_X1 U3278 ( .A1(n3290), .A2(a_9_), .ZN(n3289) );
  NOR2_X1 U3279 ( .A1(n3291), .A2(n2070), .ZN(n3290) );
  NOR2_X1 U3280 ( .A1(n3163), .A2(n3165), .ZN(n3291) );
  NAND2_X1 U3281 ( .A1(n3163), .A2(n3165), .ZN(n3288) );
  NAND2_X1 U3282 ( .A1(n3292), .A2(n3293), .ZN(n3165) );
  NAND2_X1 U3283 ( .A1(n3294), .A2(a_10_), .ZN(n3293) );
  NOR2_X1 U3284 ( .A1(n3295), .A2(n2070), .ZN(n3294) );
  NOR2_X1 U3285 ( .A1(n3208), .A2(n3206), .ZN(n3295) );
  NAND2_X1 U3286 ( .A1(n3206), .A2(n3208), .ZN(n3292) );
  NAND2_X1 U3287 ( .A1(n3296), .A2(n3297), .ZN(n3208) );
  NAND2_X1 U3288 ( .A1(n3204), .A2(n3298), .ZN(n3297) );
  NAND2_X1 U3289 ( .A1(n3203), .A2(n3202), .ZN(n3298) );
  NOR2_X1 U3290 ( .A1(n2070), .A2(n2212), .ZN(n3204) );
  OR2_X1 U3291 ( .A1(n3202), .A2(n3203), .ZN(n3296) );
  AND2_X1 U3292 ( .A1(n3199), .A2(n3299), .ZN(n3203) );
  NAND2_X1 U3293 ( .A1(n3198), .A2(n3200), .ZN(n3299) );
  NAND2_X1 U3294 ( .A1(n3300), .A2(n3301), .ZN(n3200) );
  NAND2_X1 U3295 ( .A1(b_7_), .A2(a_12_), .ZN(n3301) );
  INV_X1 U3296 ( .A(n3302), .ZN(n3300) );
  XOR2_X1 U3297 ( .A(n3303), .B(n3304), .Z(n3198) );
  NOR2_X1 U3298 ( .A1(n2210), .A2(n2216), .ZN(n3304) );
  XOR2_X1 U3299 ( .A(n3305), .B(n3306), .Z(n3303) );
  NAND2_X1 U3300 ( .A1(a_12_), .A2(n3302), .ZN(n3199) );
  NAND2_X1 U3301 ( .A1(n3307), .A2(n3308), .ZN(n3302) );
  NAND2_X1 U3302 ( .A1(n3309), .A2(b_7_), .ZN(n3308) );
  NOR2_X1 U3303 ( .A1(n3310), .A2(n2210), .ZN(n3309) );
  NOR2_X1 U3304 ( .A1(n3184), .A2(n3185), .ZN(n3310) );
  NAND2_X1 U3305 ( .A1(n3184), .A2(n3185), .ZN(n3307) );
  NAND2_X1 U3306 ( .A1(n3311), .A2(n3312), .ZN(n3185) );
  NAND2_X1 U3307 ( .A1(n3313), .A2(b_5_), .ZN(n3312) );
  NOR2_X1 U3308 ( .A1(n3314), .A2(n2208), .ZN(n3313) );
  NOR2_X1 U3309 ( .A1(n2380), .A2(n2216), .ZN(n3314) );
  NAND2_X1 U3310 ( .A1(n3315), .A2(b_6_), .ZN(n3311) );
  NOR2_X1 U3311 ( .A1(n3316), .A2(n2499), .ZN(n3315) );
  NOR2_X1 U3312 ( .A1(n2383), .A2(n2101), .ZN(n3316) );
  AND2_X1 U3313 ( .A1(n3317), .A2(b_6_), .ZN(n3184) );
  NOR2_X1 U3314 ( .A1(n2385), .A2(n2070), .ZN(n3317) );
  XOR2_X1 U3315 ( .A(n3318), .B(n3319), .Z(n3202) );
  NAND2_X1 U3316 ( .A1(n3320), .A2(n3321), .ZN(n3318) );
  XNOR2_X1 U3317 ( .A(n3322), .B(n3323), .ZN(n3206) );
  XNOR2_X1 U3318 ( .A(n3324), .B(n3325), .ZN(n3322) );
  XOR2_X1 U3319 ( .A(n3326), .B(n3327), .Z(n3163) );
  XNOR2_X1 U3320 ( .A(n3328), .B(n3329), .ZN(n3326) );
  NAND2_X1 U3321 ( .A1(a_10_), .A2(b_6_), .ZN(n3328) );
  XNOR2_X1 U3322 ( .A(n3330), .B(n3331), .ZN(n3209) );
  XOR2_X1 U3323 ( .A(n3332), .B(n3333), .Z(n3331) );
  NAND2_X1 U3324 ( .A1(a_9_), .A2(b_6_), .ZN(n3333) );
  NOR2_X1 U3325 ( .A1(n2070), .A2(n2073), .ZN(n2065) );
  INV_X1 U3326 ( .A(b_7_), .ZN(n2070) );
  XOR2_X1 U3327 ( .A(n3334), .B(n3335), .Z(n3216) );
  XOR2_X1 U3328 ( .A(n3336), .B(n3337), .Z(n3334) );
  NOR2_X1 U3329 ( .A1(n2073), .A2(n2216), .ZN(n3337) );
  XOR2_X1 U3330 ( .A(n3338), .B(n3339), .Z(n3221) );
  XNOR2_X1 U3331 ( .A(n3340), .B(n2218), .ZN(n3339) );
  XOR2_X1 U3332 ( .A(n3341), .B(n3342), .Z(n3224) );
  XOR2_X1 U3333 ( .A(n3343), .B(n3344), .Z(n3341) );
  XOR2_X1 U3334 ( .A(n3345), .B(n3346), .Z(n3228) );
  XOR2_X1 U3335 ( .A(n3347), .B(n3348), .Z(n3345) );
  XNOR2_X1 U3336 ( .A(n3349), .B(n3350), .ZN(n3233) );
  XNOR2_X1 U3337 ( .A(n3351), .B(n3352), .ZN(n3349) );
  XNOR2_X1 U3338 ( .A(n3353), .B(n3354), .ZN(n3237) );
  NAND2_X1 U3339 ( .A1(n3355), .A2(n3356), .ZN(n3353) );
  XNOR2_X1 U3340 ( .A(n3357), .B(n3358), .ZN(n3127) );
  XOR2_X1 U3341 ( .A(n3359), .B(n3360), .Z(n3358) );
  NAND2_X1 U3342 ( .A1(a_1_), .A2(b_6_), .ZN(n3360) );
  NAND2_X1 U3343 ( .A1(n3361), .A2(n3362), .ZN(n1936) );
  OR2_X1 U3344 ( .A1(n3249), .A2(n3248), .ZN(n3362) );
  XNOR2_X1 U3345 ( .A(n3363), .B(n3364), .ZN(n3361) );
  NAND2_X1 U3346 ( .A1(n3365), .A2(n3366), .ZN(n1935) );
  XNOR2_X1 U3347 ( .A(n3363), .B(n3367), .ZN(n3366) );
  INV_X1 U3348 ( .A(n3364), .ZN(n3367) );
  NOR2_X1 U3349 ( .A1(n3248), .A2(n3249), .ZN(n3365) );
  XNOR2_X1 U3350 ( .A(n3368), .B(n3369), .ZN(n3249) );
  XOR2_X1 U3351 ( .A(n3370), .B(n3371), .Z(n3368) );
  NOR2_X1 U3352 ( .A1(n2101), .A2(n2228), .ZN(n3371) );
  AND2_X1 U3353 ( .A1(n3372), .A2(n3373), .ZN(n3248) );
  NAND2_X1 U3354 ( .A1(n3374), .A2(a_0_), .ZN(n3373) );
  NOR2_X1 U3355 ( .A1(n3375), .A2(n2216), .ZN(n3374) );
  NOR2_X1 U3356 ( .A1(n3245), .A2(n3244), .ZN(n3375) );
  NAND2_X1 U3357 ( .A1(n3244), .A2(n3245), .ZN(n3372) );
  NAND2_X1 U3358 ( .A1(n3376), .A2(n3377), .ZN(n3245) );
  NAND2_X1 U3359 ( .A1(n3378), .A2(a_1_), .ZN(n3377) );
  NOR2_X1 U3360 ( .A1(n3379), .A2(n2216), .ZN(n3378) );
  NOR2_X1 U3361 ( .A1(n3357), .A2(n3359), .ZN(n3379) );
  NAND2_X1 U3362 ( .A1(n3357), .A2(n3359), .ZN(n3376) );
  NAND2_X1 U3363 ( .A1(n3355), .A2(n3380), .ZN(n3359) );
  NAND2_X1 U3364 ( .A1(n3354), .A2(n3356), .ZN(n3380) );
  NAND2_X1 U3365 ( .A1(n3381), .A2(n3382), .ZN(n3356) );
  NAND2_X1 U3366 ( .A1(a_2_), .A2(b_6_), .ZN(n3382) );
  INV_X1 U3367 ( .A(n3383), .ZN(n3381) );
  XOR2_X1 U3368 ( .A(n3384), .B(n3385), .Z(n3354) );
  XNOR2_X1 U3369 ( .A(n3386), .B(n3387), .ZN(n3384) );
  NAND2_X1 U3370 ( .A1(a_3_), .A2(b_5_), .ZN(n3386) );
  NAND2_X1 U3371 ( .A1(a_2_), .A2(n3383), .ZN(n3355) );
  NAND2_X1 U3372 ( .A1(n3388), .A2(n3389), .ZN(n3383) );
  NAND2_X1 U3373 ( .A1(n3352), .A2(n3390), .ZN(n3389) );
  NAND2_X1 U3374 ( .A1(n3351), .A2(n3350), .ZN(n3390) );
  NOR2_X1 U3375 ( .A1(n2143), .A2(n2216), .ZN(n3352) );
  OR2_X1 U3376 ( .A1(n3350), .A2(n3351), .ZN(n3388) );
  AND2_X1 U3377 ( .A1(n3391), .A2(n3392), .ZN(n3351) );
  NAND2_X1 U3378 ( .A1(n3348), .A2(n3393), .ZN(n3392) );
  OR2_X1 U3379 ( .A1(n3346), .A2(n3347), .ZN(n3393) );
  NOR2_X1 U3380 ( .A1(n2216), .A2(n2220), .ZN(n3348) );
  NAND2_X1 U3381 ( .A1(n3346), .A2(n3347), .ZN(n3391) );
  NAND2_X1 U3382 ( .A1(n3394), .A2(n3395), .ZN(n3347) );
  NAND2_X1 U3383 ( .A1(n3344), .A2(n3396), .ZN(n3395) );
  NAND2_X1 U3384 ( .A1(n3342), .A2(n3343), .ZN(n3396) );
  NOR2_X1 U3385 ( .A1(n2216), .A2(n2108), .ZN(n3344) );
  OR2_X1 U3386 ( .A1(n3342), .A2(n3343), .ZN(n3394) );
  NAND2_X1 U3387 ( .A1(n3397), .A2(n3398), .ZN(n3343) );
  NAND2_X1 U3388 ( .A1(n3338), .A2(n3399), .ZN(n3398) );
  NAND2_X1 U3389 ( .A1(n2218), .A2(n3340), .ZN(n3399) );
  XNOR2_X1 U3390 ( .A(n3400), .B(n3401), .ZN(n3338) );
  XOR2_X1 U3391 ( .A(n3402), .B(n3403), .Z(n3400) );
  NOR2_X1 U3392 ( .A1(n2073), .A2(n2101), .ZN(n3403) );
  OR2_X1 U3393 ( .A1(n3340), .A2(n2218), .ZN(n3397) );
  NOR2_X1 U3394 ( .A1(n2217), .A2(n2216), .ZN(n2218) );
  NAND2_X1 U3395 ( .A1(n3404), .A2(n3405), .ZN(n3340) );
  NAND2_X1 U3396 ( .A1(n3406), .A2(b_6_), .ZN(n3405) );
  NOR2_X1 U3397 ( .A1(n3407), .A2(n2073), .ZN(n3406) );
  NOR2_X1 U3398 ( .A1(n3336), .A2(n3335), .ZN(n3407) );
  NAND2_X1 U3399 ( .A1(n3335), .A2(n3336), .ZN(n3404) );
  NAND2_X1 U3400 ( .A1(n3283), .A2(n3408), .ZN(n3336) );
  NAND2_X1 U3401 ( .A1(n3282), .A2(n3284), .ZN(n3408) );
  NAND2_X1 U3402 ( .A1(n3409), .A2(n3410), .ZN(n3284) );
  NAND2_X1 U3403 ( .A1(a_8_), .A2(b_6_), .ZN(n3410) );
  INV_X1 U3404 ( .A(n3411), .ZN(n3409) );
  XOR2_X1 U3405 ( .A(n3412), .B(n3413), .Z(n3282) );
  XOR2_X1 U3406 ( .A(n3414), .B(n3415), .Z(n3412) );
  NOR2_X1 U3407 ( .A1(n2101), .A2(n2215), .ZN(n3415) );
  NAND2_X1 U3408 ( .A1(a_8_), .A2(n3411), .ZN(n3283) );
  NAND2_X1 U3409 ( .A1(n3416), .A2(n3417), .ZN(n3411) );
  NAND2_X1 U3410 ( .A1(n3418), .A2(a_9_), .ZN(n3417) );
  NOR2_X1 U3411 ( .A1(n3419), .A2(n2216), .ZN(n3418) );
  NOR2_X1 U3412 ( .A1(n3330), .A2(n3332), .ZN(n3419) );
  NAND2_X1 U3413 ( .A1(n3330), .A2(n3332), .ZN(n3416) );
  NAND2_X1 U3414 ( .A1(n3420), .A2(n3421), .ZN(n3332) );
  NAND2_X1 U3415 ( .A1(n3422), .A2(a_10_), .ZN(n3421) );
  NOR2_X1 U3416 ( .A1(n3423), .A2(n2216), .ZN(n3422) );
  NOR2_X1 U3417 ( .A1(n3329), .A2(n3327), .ZN(n3423) );
  NAND2_X1 U3418 ( .A1(n3327), .A2(n3329), .ZN(n3420) );
  NAND2_X1 U3419 ( .A1(n3424), .A2(n3425), .ZN(n3329) );
  NAND2_X1 U3420 ( .A1(n3325), .A2(n3426), .ZN(n3425) );
  NAND2_X1 U3421 ( .A1(n3324), .A2(n3323), .ZN(n3426) );
  NOR2_X1 U3422 ( .A1(n2216), .A2(n2212), .ZN(n3325) );
  OR2_X1 U3423 ( .A1(n3323), .A2(n3324), .ZN(n3424) );
  AND2_X1 U3424 ( .A1(n3320), .A2(n3427), .ZN(n3324) );
  NAND2_X1 U3425 ( .A1(n3319), .A2(n3321), .ZN(n3427) );
  NAND2_X1 U3426 ( .A1(n3428), .A2(n3429), .ZN(n3321) );
  NAND2_X1 U3427 ( .A1(b_6_), .A2(a_12_), .ZN(n3429) );
  INV_X1 U3428 ( .A(n3430), .ZN(n3428) );
  XOR2_X1 U3429 ( .A(n3431), .B(n3432), .Z(n3319) );
  NOR2_X1 U3430 ( .A1(n2210), .A2(n2101), .ZN(n3432) );
  XOR2_X1 U3431 ( .A(n3433), .B(n3434), .Z(n3431) );
  NAND2_X1 U3432 ( .A1(a_12_), .A2(n3430), .ZN(n3320) );
  NAND2_X1 U3433 ( .A1(n3435), .A2(n3436), .ZN(n3430) );
  NAND2_X1 U3434 ( .A1(n3437), .A2(b_6_), .ZN(n3436) );
  NOR2_X1 U3435 ( .A1(n3438), .A2(n2210), .ZN(n3437) );
  NOR2_X1 U3436 ( .A1(n3305), .A2(n3306), .ZN(n3438) );
  NAND2_X1 U3437 ( .A1(n3305), .A2(n3306), .ZN(n3435) );
  NAND2_X1 U3438 ( .A1(n3439), .A2(n3440), .ZN(n3306) );
  NAND2_X1 U3439 ( .A1(n3441), .A2(b_4_), .ZN(n3440) );
  NOR2_X1 U3440 ( .A1(n3442), .A2(n2208), .ZN(n3441) );
  NOR2_X1 U3441 ( .A1(n2380), .A2(n2101), .ZN(n3442) );
  NAND2_X1 U3442 ( .A1(n3443), .A2(b_5_), .ZN(n3439) );
  NOR2_X1 U3443 ( .A1(n3444), .A2(n2499), .ZN(n3443) );
  NOR2_X1 U3444 ( .A1(n2383), .A2(n2219), .ZN(n3444) );
  AND2_X1 U3445 ( .A1(n3445), .A2(b_5_), .ZN(n3305) );
  NOR2_X1 U3446 ( .A1(n2385), .A2(n2216), .ZN(n3445) );
  INV_X1 U3447 ( .A(b_6_), .ZN(n2216) );
  XOR2_X1 U3448 ( .A(n3446), .B(n3447), .Z(n3323) );
  NAND2_X1 U3449 ( .A1(n3448), .A2(n3449), .ZN(n3446) );
  XNOR2_X1 U3450 ( .A(n3450), .B(n3451), .ZN(n3327) );
  XNOR2_X1 U3451 ( .A(n3452), .B(n3453), .ZN(n3450) );
  XOR2_X1 U3452 ( .A(n3454), .B(n3455), .Z(n3330) );
  XNOR2_X1 U3453 ( .A(n3456), .B(n3457), .ZN(n3454) );
  NAND2_X1 U3454 ( .A1(b_5_), .A2(a_10_), .ZN(n3456) );
  XNOR2_X1 U3455 ( .A(n3458), .B(n3459), .ZN(n3335) );
  NAND2_X1 U3456 ( .A1(n3460), .A2(n3461), .ZN(n3458) );
  XOR2_X1 U3457 ( .A(n3462), .B(n3463), .Z(n3342) );
  XOR2_X1 U3458 ( .A(n3464), .B(n3465), .Z(n3463) );
  NAND2_X1 U3459 ( .A1(a_6_), .A2(b_5_), .ZN(n3465) );
  XNOR2_X1 U3460 ( .A(n3466), .B(n3467), .ZN(n3346) );
  XNOR2_X1 U3461 ( .A(n2096), .B(n3468), .ZN(n3467) );
  XNOR2_X1 U3462 ( .A(n3469), .B(n3470), .ZN(n3350) );
  XNOR2_X1 U3463 ( .A(n3471), .B(n3472), .ZN(n3469) );
  NAND2_X1 U3464 ( .A1(b_5_), .A2(a_4_), .ZN(n3471) );
  XOR2_X1 U3465 ( .A(n3473), .B(n3474), .Z(n3357) );
  XOR2_X1 U3466 ( .A(n3475), .B(n3476), .Z(n3473) );
  NOR2_X1 U3467 ( .A1(n2101), .A2(n2222), .ZN(n3476) );
  XOR2_X1 U3468 ( .A(n3477), .B(n3478), .Z(n3244) );
  XOR2_X1 U3469 ( .A(n3479), .B(n3480), .Z(n3477) );
  NOR2_X1 U3470 ( .A1(n2101), .A2(n2319), .ZN(n3480) );
  NAND2_X1 U3471 ( .A1(n3481), .A2(n3482), .ZN(n1941) );
  NAND2_X1 U3472 ( .A1(n3364), .A2(n3363), .ZN(n3482) );
  XNOR2_X1 U3473 ( .A(n3483), .B(n3484), .ZN(n3481) );
  NAND2_X1 U3474 ( .A1(n3485), .A2(n3486), .ZN(n1940) );
  XNOR2_X1 U3475 ( .A(n3487), .B(n3484), .ZN(n3486) );
  AND2_X1 U3476 ( .A1(n3363), .A2(n3364), .ZN(n3485) );
  XNOR2_X1 U3477 ( .A(n3488), .B(n3489), .ZN(n3364) );
  XOR2_X1 U3478 ( .A(n3490), .B(n3491), .Z(n3489) );
  NAND2_X1 U3479 ( .A1(a_0_), .A2(b_4_), .ZN(n3491) );
  NAND2_X1 U3480 ( .A1(n3492), .A2(n3493), .ZN(n3363) );
  NAND2_X1 U3481 ( .A1(n3494), .A2(a_0_), .ZN(n3493) );
  NOR2_X1 U3482 ( .A1(n3495), .A2(n2101), .ZN(n3494) );
  NOR2_X1 U3483 ( .A1(n3370), .A2(n3369), .ZN(n3495) );
  NAND2_X1 U3484 ( .A1(n3369), .A2(n3370), .ZN(n3492) );
  NAND2_X1 U3485 ( .A1(n3496), .A2(n3497), .ZN(n3370) );
  NAND2_X1 U3486 ( .A1(n3498), .A2(a_1_), .ZN(n3497) );
  NOR2_X1 U3487 ( .A1(n3499), .A2(n2101), .ZN(n3498) );
  NOR2_X1 U3488 ( .A1(n3478), .A2(n3479), .ZN(n3499) );
  NAND2_X1 U3489 ( .A1(n3478), .A2(n3479), .ZN(n3496) );
  NAND2_X1 U3490 ( .A1(n3500), .A2(n3501), .ZN(n3479) );
  NAND2_X1 U3491 ( .A1(n3502), .A2(a_2_), .ZN(n3501) );
  NOR2_X1 U3492 ( .A1(n3503), .A2(n2101), .ZN(n3502) );
  NOR2_X1 U3493 ( .A1(n3475), .A2(n3474), .ZN(n3503) );
  NAND2_X1 U3494 ( .A1(n3474), .A2(n3475), .ZN(n3500) );
  NAND2_X1 U3495 ( .A1(n3504), .A2(n3505), .ZN(n3475) );
  NAND2_X1 U3496 ( .A1(n3506), .A2(a_3_), .ZN(n3505) );
  NOR2_X1 U3497 ( .A1(n3507), .A2(n2101), .ZN(n3506) );
  NOR2_X1 U3498 ( .A1(n3385), .A2(n3387), .ZN(n3507) );
  NAND2_X1 U3499 ( .A1(n3385), .A2(n3387), .ZN(n3504) );
  NAND2_X1 U3500 ( .A1(n3508), .A2(n3509), .ZN(n3387) );
  NAND2_X1 U3501 ( .A1(n3510), .A2(b_5_), .ZN(n3509) );
  NOR2_X1 U3502 ( .A1(n3511), .A2(n2220), .ZN(n3510) );
  NOR2_X1 U3503 ( .A1(n3472), .A2(n3470), .ZN(n3511) );
  NAND2_X1 U3504 ( .A1(n3470), .A2(n3472), .ZN(n3508) );
  NAND2_X1 U3505 ( .A1(n3512), .A2(n3513), .ZN(n3472) );
  NAND2_X1 U3506 ( .A1(n3466), .A2(n3514), .ZN(n3513) );
  OR2_X1 U3507 ( .A1(n3468), .A2(n2096), .ZN(n3514) );
  XOR2_X1 U3508 ( .A(n3515), .B(n3516), .Z(n3466) );
  XOR2_X1 U3509 ( .A(n3517), .B(n3518), .Z(n3515) );
  NOR2_X1 U3510 ( .A1(n2219), .A2(n2217), .ZN(n3518) );
  NAND2_X1 U3511 ( .A1(n2096), .A2(n3468), .ZN(n3512) );
  NAND2_X1 U3512 ( .A1(n3519), .A2(n3520), .ZN(n3468) );
  NAND2_X1 U3513 ( .A1(n3521), .A2(a_6_), .ZN(n3520) );
  NOR2_X1 U3514 ( .A1(n3522), .A2(n2101), .ZN(n3521) );
  NOR2_X1 U3515 ( .A1(n3464), .A2(n3462), .ZN(n3522) );
  NAND2_X1 U3516 ( .A1(n3462), .A2(n3464), .ZN(n3519) );
  NAND2_X1 U3517 ( .A1(n3523), .A2(n3524), .ZN(n3464) );
  NAND2_X1 U3518 ( .A1(n3525), .A2(b_5_), .ZN(n3524) );
  NOR2_X1 U3519 ( .A1(n3526), .A2(n2073), .ZN(n3525) );
  NOR2_X1 U3520 ( .A1(n3402), .A2(n3401), .ZN(n3526) );
  NAND2_X1 U3521 ( .A1(n3401), .A2(n3402), .ZN(n3523) );
  NAND2_X1 U3522 ( .A1(n3460), .A2(n3527), .ZN(n3402) );
  NAND2_X1 U3523 ( .A1(n3459), .A2(n3461), .ZN(n3527) );
  NAND2_X1 U3524 ( .A1(n3528), .A2(n3529), .ZN(n3461) );
  NAND2_X1 U3525 ( .A1(a_8_), .A2(b_5_), .ZN(n3529) );
  INV_X1 U3526 ( .A(n3530), .ZN(n3528) );
  XNOR2_X1 U3527 ( .A(n3531), .B(n3532), .ZN(n3459) );
  XNOR2_X1 U3528 ( .A(n3533), .B(n3534), .ZN(n3531) );
  NAND2_X1 U3529 ( .A1(a_8_), .A2(n3530), .ZN(n3460) );
  NAND2_X1 U3530 ( .A1(n3535), .A2(n3536), .ZN(n3530) );
  NAND2_X1 U3531 ( .A1(n3537), .A2(a_9_), .ZN(n3536) );
  NOR2_X1 U3532 ( .A1(n3538), .A2(n2101), .ZN(n3537) );
  NOR2_X1 U3533 ( .A1(n3413), .A2(n3414), .ZN(n3538) );
  NAND2_X1 U3534 ( .A1(n3413), .A2(n3414), .ZN(n3535) );
  NAND2_X1 U3535 ( .A1(n3539), .A2(n3540), .ZN(n3414) );
  NAND2_X1 U3536 ( .A1(n3541), .A2(b_5_), .ZN(n3540) );
  NOR2_X1 U3537 ( .A1(n3542), .A2(n2214), .ZN(n3541) );
  NOR2_X1 U3538 ( .A1(n3457), .A2(n3455), .ZN(n3542) );
  NAND2_X1 U3539 ( .A1(n3455), .A2(n3457), .ZN(n3539) );
  NAND2_X1 U3540 ( .A1(n3543), .A2(n3544), .ZN(n3457) );
  NAND2_X1 U3541 ( .A1(n3453), .A2(n3545), .ZN(n3544) );
  NAND2_X1 U3542 ( .A1(n3452), .A2(n3451), .ZN(n3545) );
  NOR2_X1 U3543 ( .A1(n2101), .A2(n2212), .ZN(n3453) );
  OR2_X1 U3544 ( .A1(n3451), .A2(n3452), .ZN(n3543) );
  AND2_X1 U3545 ( .A1(n3448), .A2(n3546), .ZN(n3452) );
  NAND2_X1 U3546 ( .A1(n3447), .A2(n3449), .ZN(n3546) );
  NAND2_X1 U3547 ( .A1(n3547), .A2(n3548), .ZN(n3449) );
  NAND2_X1 U3548 ( .A1(b_5_), .A2(a_12_), .ZN(n3548) );
  INV_X1 U3549 ( .A(n3549), .ZN(n3547) );
  XOR2_X1 U3550 ( .A(n3550), .B(n3551), .Z(n3447) );
  NOR2_X1 U3551 ( .A1(n2210), .A2(n2219), .ZN(n3551) );
  XOR2_X1 U3552 ( .A(n3552), .B(n3553), .Z(n3550) );
  NAND2_X1 U3553 ( .A1(a_12_), .A2(n3549), .ZN(n3448) );
  NAND2_X1 U3554 ( .A1(n3554), .A2(n3555), .ZN(n3549) );
  NAND2_X1 U3555 ( .A1(n3556), .A2(b_5_), .ZN(n3555) );
  NOR2_X1 U3556 ( .A1(n3557), .A2(n2210), .ZN(n3556) );
  NOR2_X1 U3557 ( .A1(n3433), .A2(n3434), .ZN(n3557) );
  NAND2_X1 U3558 ( .A1(n3433), .A2(n3434), .ZN(n3554) );
  NAND2_X1 U3559 ( .A1(n3558), .A2(n3559), .ZN(n3434) );
  NAND2_X1 U3560 ( .A1(n3560), .A2(b_3_), .ZN(n3559) );
  NOR2_X1 U3561 ( .A1(n3561), .A2(n2208), .ZN(n3560) );
  NOR2_X1 U3562 ( .A1(n2380), .A2(n2219), .ZN(n3561) );
  NAND2_X1 U3563 ( .A1(n3562), .A2(b_4_), .ZN(n3558) );
  NOR2_X1 U3564 ( .A1(n3563), .A2(n2499), .ZN(n3562) );
  NOR2_X1 U3565 ( .A1(n2383), .A2(n2136), .ZN(n3563) );
  AND2_X1 U3566 ( .A1(n3564), .A2(b_4_), .ZN(n3433) );
  NOR2_X1 U3567 ( .A1(n2385), .A2(n2101), .ZN(n3564) );
  XOR2_X1 U3568 ( .A(n3565), .B(n3566), .Z(n3451) );
  NAND2_X1 U3569 ( .A1(n3567), .A2(n3568), .ZN(n3565) );
  XOR2_X1 U3570 ( .A(n3569), .B(n3570), .Z(n3455) );
  XOR2_X1 U3571 ( .A(n3571), .B(n3572), .Z(n3569) );
  NOR2_X1 U3572 ( .A1(n2212), .A2(n2219), .ZN(n3572) );
  XOR2_X1 U3573 ( .A(n3573), .B(n3574), .Z(n3413) );
  XOR2_X1 U3574 ( .A(n3575), .B(n3576), .Z(n3573) );
  NOR2_X1 U3575 ( .A1(n2214), .A2(n2219), .ZN(n3576) );
  XNOR2_X1 U3576 ( .A(n3577), .B(n3578), .ZN(n3401) );
  NAND2_X1 U3577 ( .A1(n3579), .A2(n3580), .ZN(n3577) );
  XOR2_X1 U3578 ( .A(n3581), .B(n3582), .Z(n3462) );
  XOR2_X1 U3579 ( .A(n3583), .B(n3584), .Z(n3581) );
  NOR2_X1 U3580 ( .A1(n2073), .A2(n2219), .ZN(n3584) );
  NOR2_X1 U3581 ( .A1(n2101), .A2(n2108), .ZN(n2096) );
  INV_X1 U3582 ( .A(b_5_), .ZN(n2101) );
  XOR2_X1 U3583 ( .A(n3585), .B(n3586), .Z(n3470) );
  XOR2_X1 U3584 ( .A(n3587), .B(n3588), .Z(n3585) );
  NOR2_X1 U3585 ( .A1(n2108), .A2(n2219), .ZN(n3588) );
  XOR2_X1 U3586 ( .A(n3589), .B(n3590), .Z(n3385) );
  XNOR2_X1 U3587 ( .A(n3591), .B(n2115), .ZN(n3589) );
  INV_X1 U3588 ( .A(n3592), .ZN(n2115) );
  XOR2_X1 U3589 ( .A(n3593), .B(n3594), .Z(n3474) );
  XOR2_X1 U3590 ( .A(n3595), .B(n3596), .Z(n3593) );
  NOR2_X1 U3591 ( .A1(n2219), .A2(n2143), .ZN(n3596) );
  XOR2_X1 U3592 ( .A(n3597), .B(n3598), .Z(n3478) );
  XOR2_X1 U3593 ( .A(n3599), .B(n3600), .Z(n3597) );
  NOR2_X1 U3594 ( .A1(n2219), .A2(n2222), .ZN(n3600) );
  XOR2_X1 U3595 ( .A(n3601), .B(n3602), .Z(n3369) );
  XOR2_X1 U3596 ( .A(n3603), .B(n3604), .Z(n3601) );
  NOR2_X1 U3597 ( .A1(n2219), .A2(n2319), .ZN(n3604) );
  NAND2_X1 U3598 ( .A1(n3605), .A2(n3606), .ZN(n1946) );
  NAND2_X1 U3599 ( .A1(n3484), .A2(n3483), .ZN(n3606) );
  NAND2_X1 U3600 ( .A1(n3607), .A2(n3484), .ZN(n1945) );
  XOR2_X1 U3601 ( .A(n3608), .B(n3609), .Z(n3484) );
  XOR2_X1 U3602 ( .A(n3610), .B(n3611), .Z(n3608) );
  NOR2_X1 U3603 ( .A1(n2136), .A2(n2228), .ZN(n3611) );
  NOR2_X1 U3604 ( .A1(n3487), .A2(n3605), .ZN(n3607) );
  XNOR2_X1 U3605 ( .A(n3612), .B(n3613), .ZN(n3605) );
  INV_X1 U3606 ( .A(n3483), .ZN(n3487) );
  NAND2_X1 U3607 ( .A1(n3614), .A2(n3615), .ZN(n3483) );
  NAND2_X1 U3608 ( .A1(n3616), .A2(a_0_), .ZN(n3615) );
  NOR2_X1 U3609 ( .A1(n3617), .A2(n2219), .ZN(n3616) );
  NOR2_X1 U3610 ( .A1(n3488), .A2(n3490), .ZN(n3617) );
  NAND2_X1 U3611 ( .A1(n3488), .A2(n3490), .ZN(n3614) );
  NAND2_X1 U3612 ( .A1(n3618), .A2(n3619), .ZN(n3490) );
  NAND2_X1 U3613 ( .A1(n3620), .A2(a_1_), .ZN(n3619) );
  NOR2_X1 U3614 ( .A1(n3621), .A2(n2219), .ZN(n3620) );
  NOR2_X1 U3615 ( .A1(n3602), .A2(n3603), .ZN(n3621) );
  NAND2_X1 U3616 ( .A1(n3602), .A2(n3603), .ZN(n3618) );
  NAND2_X1 U3617 ( .A1(n3622), .A2(n3623), .ZN(n3603) );
  NAND2_X1 U3618 ( .A1(n3624), .A2(a_2_), .ZN(n3623) );
  NOR2_X1 U3619 ( .A1(n3625), .A2(n2219), .ZN(n3624) );
  NOR2_X1 U3620 ( .A1(n3599), .A2(n3598), .ZN(n3625) );
  NAND2_X1 U3621 ( .A1(n3598), .A2(n3599), .ZN(n3622) );
  NAND2_X1 U3622 ( .A1(n3626), .A2(n3627), .ZN(n3599) );
  NAND2_X1 U3623 ( .A1(n3628), .A2(a_3_), .ZN(n3627) );
  NOR2_X1 U3624 ( .A1(n3629), .A2(n2219), .ZN(n3628) );
  NOR2_X1 U3625 ( .A1(n3594), .A2(n3595), .ZN(n3629) );
  NAND2_X1 U3626 ( .A1(n3594), .A2(n3595), .ZN(n3626) );
  NAND2_X1 U3627 ( .A1(n3630), .A2(n3631), .ZN(n3595) );
  NAND2_X1 U3628 ( .A1(n3590), .A2(n3632), .ZN(n3631) );
  OR2_X1 U3629 ( .A1(n3591), .A2(n3592), .ZN(n3632) );
  XOR2_X1 U3630 ( .A(n3633), .B(n3634), .Z(n3590) );
  XOR2_X1 U3631 ( .A(n3635), .B(n3636), .Z(n3633) );
  NOR2_X1 U3632 ( .A1(n2108), .A2(n2136), .ZN(n3636) );
  NAND2_X1 U3633 ( .A1(n3592), .A2(n3591), .ZN(n3630) );
  NAND2_X1 U3634 ( .A1(n3637), .A2(n3638), .ZN(n3591) );
  NAND2_X1 U3635 ( .A1(n3639), .A2(b_4_), .ZN(n3638) );
  NOR2_X1 U3636 ( .A1(n3640), .A2(n2108), .ZN(n3639) );
  NOR2_X1 U3637 ( .A1(n3586), .A2(n3587), .ZN(n3640) );
  NAND2_X1 U3638 ( .A1(n3586), .A2(n3587), .ZN(n3637) );
  NAND2_X1 U3639 ( .A1(n3641), .A2(n3642), .ZN(n3587) );
  NAND2_X1 U3640 ( .A1(n3643), .A2(a_6_), .ZN(n3642) );
  NOR2_X1 U3641 ( .A1(n3644), .A2(n2219), .ZN(n3643) );
  NOR2_X1 U3642 ( .A1(n3517), .A2(n3516), .ZN(n3644) );
  NAND2_X1 U3643 ( .A1(n3516), .A2(n3517), .ZN(n3641) );
  NAND2_X1 U3644 ( .A1(n3645), .A2(n3646), .ZN(n3517) );
  NAND2_X1 U3645 ( .A1(n3647), .A2(b_4_), .ZN(n3646) );
  NOR2_X1 U3646 ( .A1(n3648), .A2(n2073), .ZN(n3647) );
  NOR2_X1 U3647 ( .A1(n3582), .A2(n3583), .ZN(n3648) );
  NAND2_X1 U3648 ( .A1(n3582), .A2(n3583), .ZN(n3645) );
  NAND2_X1 U3649 ( .A1(n3579), .A2(n3649), .ZN(n3583) );
  NAND2_X1 U3650 ( .A1(n3578), .A2(n3580), .ZN(n3649) );
  NAND2_X1 U3651 ( .A1(n3650), .A2(n3651), .ZN(n3580) );
  NAND2_X1 U3652 ( .A1(b_4_), .A2(a_8_), .ZN(n3651) );
  INV_X1 U3653 ( .A(n3652), .ZN(n3650) );
  XOR2_X1 U3654 ( .A(n3653), .B(n3654), .Z(n3578) );
  XOR2_X1 U3655 ( .A(n3655), .B(n3656), .Z(n3653) );
  NOR2_X1 U3656 ( .A1(n2215), .A2(n2136), .ZN(n3656) );
  NAND2_X1 U3657 ( .A1(a_8_), .A2(n3652), .ZN(n3579) );
  NAND2_X1 U3658 ( .A1(n3657), .A2(n3658), .ZN(n3652) );
  NAND2_X1 U3659 ( .A1(n3533), .A2(n3659), .ZN(n3658) );
  NAND2_X1 U3660 ( .A1(n3534), .A2(n3532), .ZN(n3659) );
  NOR2_X1 U3661 ( .A1(n2219), .A2(n2215), .ZN(n3533) );
  OR2_X1 U3662 ( .A1(n3532), .A2(n3534), .ZN(n3657) );
  AND2_X1 U3663 ( .A1(n3660), .A2(n3661), .ZN(n3534) );
  NAND2_X1 U3664 ( .A1(n3662), .A2(b_4_), .ZN(n3661) );
  NOR2_X1 U3665 ( .A1(n3663), .A2(n2214), .ZN(n3662) );
  NOR2_X1 U3666 ( .A1(n3575), .A2(n3574), .ZN(n3663) );
  NAND2_X1 U3667 ( .A1(n3574), .A2(n3575), .ZN(n3660) );
  NAND2_X1 U3668 ( .A1(n3664), .A2(n3665), .ZN(n3575) );
  NAND2_X1 U3669 ( .A1(n3666), .A2(b_4_), .ZN(n3665) );
  NOR2_X1 U3670 ( .A1(n3667), .A2(n2212), .ZN(n3666) );
  NOR2_X1 U3671 ( .A1(n3570), .A2(n3571), .ZN(n3667) );
  NAND2_X1 U3672 ( .A1(n3570), .A2(n3571), .ZN(n3664) );
  NAND2_X1 U3673 ( .A1(n3567), .A2(n3668), .ZN(n3571) );
  NAND2_X1 U3674 ( .A1(n3566), .A2(n3568), .ZN(n3668) );
  NAND2_X1 U3675 ( .A1(n3669), .A2(n3670), .ZN(n3568) );
  NAND2_X1 U3676 ( .A1(b_4_), .A2(a_12_), .ZN(n3670) );
  INV_X1 U3677 ( .A(n3671), .ZN(n3669) );
  XOR2_X1 U3678 ( .A(n3672), .B(n3673), .Z(n3566) );
  XOR2_X1 U3679 ( .A(n3674), .B(n3675), .Z(n3672) );
  NAND2_X1 U3680 ( .A1(a_12_), .A2(n3671), .ZN(n3567) );
  NAND2_X1 U3681 ( .A1(n3676), .A2(n3677), .ZN(n3671) );
  NAND2_X1 U3682 ( .A1(n3678), .A2(b_4_), .ZN(n3677) );
  NOR2_X1 U3683 ( .A1(n3679), .A2(n2210), .ZN(n3678) );
  NOR2_X1 U3684 ( .A1(n3552), .A2(n3553), .ZN(n3679) );
  NAND2_X1 U3685 ( .A1(n3552), .A2(n3553), .ZN(n3676) );
  NAND2_X1 U3686 ( .A1(n3680), .A2(n3681), .ZN(n3553) );
  NAND2_X1 U3687 ( .A1(n3682), .A2(b_2_), .ZN(n3681) );
  NOR2_X1 U3688 ( .A1(n3683), .A2(n2208), .ZN(n3682) );
  NOR2_X1 U3689 ( .A1(n2380), .A2(n2136), .ZN(n3683) );
  NAND2_X1 U3690 ( .A1(n3684), .A2(b_3_), .ZN(n3680) );
  NOR2_X1 U3691 ( .A1(n3685), .A2(n2499), .ZN(n3684) );
  NOR2_X1 U3692 ( .A1(n2383), .A2(n2221), .ZN(n3685) );
  AND2_X1 U3693 ( .A1(n3686), .A2(b_3_), .ZN(n3552) );
  NOR2_X1 U3694 ( .A1(n2385), .A2(n2219), .ZN(n3686) );
  XNOR2_X1 U3695 ( .A(n3687), .B(n3688), .ZN(n3570) );
  NAND2_X1 U3696 ( .A1(n3689), .A2(n3690), .ZN(n3687) );
  XOR2_X1 U3697 ( .A(n3691), .B(n3692), .Z(n3574) );
  XOR2_X1 U3698 ( .A(n3693), .B(n3694), .Z(n3691) );
  NOR2_X1 U3699 ( .A1(n2212), .A2(n2136), .ZN(n3694) );
  XNOR2_X1 U3700 ( .A(n3695), .B(n3696), .ZN(n3532) );
  XOR2_X1 U3701 ( .A(n3697), .B(n3698), .Z(n3695) );
  NOR2_X1 U3702 ( .A1(n2214), .A2(n2136), .ZN(n3698) );
  XOR2_X1 U3703 ( .A(n3699), .B(n3700), .Z(n3582) );
  XOR2_X1 U3704 ( .A(n3701), .B(n3702), .Z(n3699) );
  NOR2_X1 U3705 ( .A1(n2059), .A2(n2136), .ZN(n3702) );
  XOR2_X1 U3706 ( .A(n3703), .B(n3704), .Z(n3516) );
  XOR2_X1 U3707 ( .A(n3705), .B(n3706), .Z(n3703) );
  NOR2_X1 U3708 ( .A1(n2073), .A2(n2136), .ZN(n3706) );
  XOR2_X1 U3709 ( .A(n3707), .B(n3708), .Z(n3586) );
  XOR2_X1 U3710 ( .A(n3709), .B(n3710), .Z(n3707) );
  NOR2_X1 U3711 ( .A1(n2136), .A2(n2217), .ZN(n3710) );
  NOR2_X1 U3712 ( .A1(n2219), .A2(n2220), .ZN(n3592) );
  INV_X1 U3713 ( .A(b_4_), .ZN(n2219) );
  XOR2_X1 U3714 ( .A(n3711), .B(n3712), .Z(n3594) );
  XOR2_X1 U3715 ( .A(n3713), .B(n3714), .Z(n3711) );
  NOR2_X1 U3716 ( .A1(n2220), .A2(n2136), .ZN(n3714) );
  XOR2_X1 U3717 ( .A(n3715), .B(n3716), .Z(n3598) );
  XNOR2_X1 U3718 ( .A(n3717), .B(n2182), .ZN(n3715) );
  INV_X1 U3719 ( .A(n2131), .ZN(n2182) );
  XOR2_X1 U3720 ( .A(n3718), .B(n3719), .Z(n3602) );
  XNOR2_X1 U3721 ( .A(n3720), .B(n3721), .ZN(n3718) );
  NAND2_X1 U3722 ( .A1(a_2_), .A2(b_3_), .ZN(n3720) );
  XOR2_X1 U3723 ( .A(n3722), .B(n3723), .Z(n3488) );
  XOR2_X1 U3724 ( .A(n3724), .B(n3725), .Z(n3722) );
  NOR2_X1 U3725 ( .A1(n2136), .A2(n2319), .ZN(n3725) );
  NAND2_X1 U3726 ( .A1(n3726), .A2(n3727), .ZN(n1970) );
  NAND2_X1 U3727 ( .A1(n3728), .A2(n3729), .ZN(n3727) );
  NAND2_X1 U3728 ( .A1(n3730), .A2(n3728), .ZN(n1969) );
  INV_X1 U3729 ( .A(n3613), .ZN(n3728) );
  XOR2_X1 U3730 ( .A(n3731), .B(n3732), .Z(n3613) );
  NAND2_X1 U3731 ( .A1(n3733), .A2(n3734), .ZN(n3731) );
  NOR2_X1 U3732 ( .A1(n3612), .A2(n3726), .ZN(n3730) );
  XNOR2_X1 U3733 ( .A(n2272), .B(n2273), .ZN(n3726) );
  INV_X1 U3734 ( .A(n3729), .ZN(n3612) );
  NAND2_X1 U3735 ( .A1(n3735), .A2(n3736), .ZN(n3729) );
  NAND2_X1 U3736 ( .A1(n3737), .A2(a_0_), .ZN(n3736) );
  NOR2_X1 U3737 ( .A1(n3738), .A2(n2136), .ZN(n3737) );
  NOR2_X1 U3738 ( .A1(n3610), .A2(n3609), .ZN(n3738) );
  NAND2_X1 U3739 ( .A1(n3609), .A2(n3610), .ZN(n3735) );
  NAND2_X1 U3740 ( .A1(n3739), .A2(n3740), .ZN(n3610) );
  NAND2_X1 U3741 ( .A1(n3741), .A2(a_1_), .ZN(n3740) );
  NOR2_X1 U3742 ( .A1(n3742), .A2(n2136), .ZN(n3741) );
  NOR2_X1 U3743 ( .A1(n3724), .A2(n3723), .ZN(n3742) );
  NAND2_X1 U3744 ( .A1(n3723), .A2(n3724), .ZN(n3739) );
  NAND2_X1 U3745 ( .A1(n3743), .A2(n3744), .ZN(n3724) );
  NAND2_X1 U3746 ( .A1(n3745), .A2(a_2_), .ZN(n3744) );
  NOR2_X1 U3747 ( .A1(n3746), .A2(n2136), .ZN(n3745) );
  NOR2_X1 U3748 ( .A1(n3721), .A2(n3719), .ZN(n3746) );
  NAND2_X1 U3749 ( .A1(n3719), .A2(n3721), .ZN(n3743) );
  NAND2_X1 U3750 ( .A1(n3747), .A2(n3748), .ZN(n3721) );
  NAND2_X1 U3751 ( .A1(n3716), .A2(n3749), .ZN(n3748) );
  OR2_X1 U3752 ( .A1(n3717), .A2(n2131), .ZN(n3749) );
  XNOR2_X1 U3753 ( .A(n3750), .B(n3751), .ZN(n3716) );
  NAND2_X1 U3754 ( .A1(n3752), .A2(n3753), .ZN(n3750) );
  NAND2_X1 U3755 ( .A1(n2131), .A2(n3717), .ZN(n3747) );
  NAND2_X1 U3756 ( .A1(n3754), .A2(n3755), .ZN(n3717) );
  NAND2_X1 U3757 ( .A1(n3756), .A2(b_3_), .ZN(n3755) );
  NOR2_X1 U3758 ( .A1(n3757), .A2(n2220), .ZN(n3756) );
  NOR2_X1 U3759 ( .A1(n3713), .A2(n3712), .ZN(n3757) );
  NAND2_X1 U3760 ( .A1(n3712), .A2(n3713), .ZN(n3754) );
  NAND2_X1 U3761 ( .A1(n3758), .A2(n3759), .ZN(n3713) );
  NAND2_X1 U3762 ( .A1(n3760), .A2(b_3_), .ZN(n3759) );
  NOR2_X1 U3763 ( .A1(n3761), .A2(n2108), .ZN(n3760) );
  NOR2_X1 U3764 ( .A1(n3634), .A2(n3635), .ZN(n3761) );
  NAND2_X1 U3765 ( .A1(n3634), .A2(n3635), .ZN(n3758) );
  NAND2_X1 U3766 ( .A1(n3762), .A2(n3763), .ZN(n3635) );
  NAND2_X1 U3767 ( .A1(n3764), .A2(a_6_), .ZN(n3763) );
  NOR2_X1 U3768 ( .A1(n3765), .A2(n2136), .ZN(n3764) );
  NOR2_X1 U3769 ( .A1(n3709), .A2(n3708), .ZN(n3765) );
  NAND2_X1 U3770 ( .A1(n3708), .A2(n3709), .ZN(n3762) );
  NAND2_X1 U3771 ( .A1(n3766), .A2(n3767), .ZN(n3709) );
  NAND2_X1 U3772 ( .A1(n3768), .A2(b_3_), .ZN(n3767) );
  NOR2_X1 U3773 ( .A1(n3769), .A2(n2073), .ZN(n3768) );
  NOR2_X1 U3774 ( .A1(n3704), .A2(n3705), .ZN(n3769) );
  NAND2_X1 U3775 ( .A1(n3704), .A2(n3705), .ZN(n3766) );
  NAND2_X1 U3776 ( .A1(n3770), .A2(n3771), .ZN(n3705) );
  NAND2_X1 U3777 ( .A1(n3772), .A2(b_3_), .ZN(n3771) );
  NOR2_X1 U3778 ( .A1(n3773), .A2(n2059), .ZN(n3772) );
  NOR2_X1 U3779 ( .A1(n3701), .A2(n3700), .ZN(n3773) );
  NAND2_X1 U3780 ( .A1(n3700), .A2(n3701), .ZN(n3770) );
  NAND2_X1 U3781 ( .A1(n3774), .A2(n3775), .ZN(n3701) );
  NAND2_X1 U3782 ( .A1(n3776), .A2(b_3_), .ZN(n3775) );
  NOR2_X1 U3783 ( .A1(n3777), .A2(n2215), .ZN(n3776) );
  NOR2_X1 U3784 ( .A1(n3654), .A2(n3655), .ZN(n3777) );
  NAND2_X1 U3785 ( .A1(n3654), .A2(n3655), .ZN(n3774) );
  NAND2_X1 U3786 ( .A1(n3778), .A2(n3779), .ZN(n3655) );
  NAND2_X1 U3787 ( .A1(n3780), .A2(b_3_), .ZN(n3779) );
  NOR2_X1 U3788 ( .A1(n3781), .A2(n2214), .ZN(n3780) );
  NOR2_X1 U3789 ( .A1(n3697), .A2(n3696), .ZN(n3781) );
  NAND2_X1 U3790 ( .A1(n3696), .A2(n3697), .ZN(n3778) );
  NAND2_X1 U3791 ( .A1(n3782), .A2(n3783), .ZN(n3697) );
  NAND2_X1 U3792 ( .A1(n3784), .A2(b_3_), .ZN(n3783) );
  NOR2_X1 U3793 ( .A1(n3785), .A2(n2212), .ZN(n3784) );
  NOR2_X1 U3794 ( .A1(n3692), .A2(n3693), .ZN(n3785) );
  NAND2_X1 U3795 ( .A1(n3692), .A2(n3693), .ZN(n3782) );
  NAND2_X1 U3796 ( .A1(n3689), .A2(n3786), .ZN(n3693) );
  NAND2_X1 U3797 ( .A1(n3688), .A2(n3690), .ZN(n3786) );
  NAND2_X1 U3798 ( .A1(n3787), .A2(n3788), .ZN(n3690) );
  NAND2_X1 U3799 ( .A1(b_3_), .A2(a_12_), .ZN(n3788) );
  INV_X1 U3800 ( .A(n3789), .ZN(n3787) );
  XOR2_X1 U3801 ( .A(n3790), .B(n3791), .Z(n3688) );
  NOR2_X1 U3802 ( .A1(n2210), .A2(n2221), .ZN(n3791) );
  XOR2_X1 U3803 ( .A(n3792), .B(n3793), .Z(n3790) );
  NAND2_X1 U3804 ( .A1(a_12_), .A2(n3789), .ZN(n3689) );
  NAND2_X1 U3805 ( .A1(n3794), .A2(n3795), .ZN(n3789) );
  NAND2_X1 U3806 ( .A1(n3673), .A2(n3796), .ZN(n3795) );
  NAND2_X1 U3807 ( .A1(n3675), .A2(n3674), .ZN(n3796) );
  NOR2_X1 U3808 ( .A1(n2136), .A2(n2210), .ZN(n3673) );
  OR2_X1 U3809 ( .A1(n3674), .A2(n3675), .ZN(n3794) );
  AND2_X1 U3810 ( .A1(n3797), .A2(n3798), .ZN(n3675) );
  NAND2_X1 U3811 ( .A1(n3799), .A2(b_1_), .ZN(n3798) );
  NOR2_X1 U3812 ( .A1(n3800), .A2(n2208), .ZN(n3799) );
  NOR2_X1 U3813 ( .A1(n2380), .A2(n2221), .ZN(n3800) );
  NAND2_X1 U3814 ( .A1(n3801), .A2(b_2_), .ZN(n3797) );
  NOR2_X1 U3815 ( .A1(n3802), .A2(n2499), .ZN(n3801) );
  NOR2_X1 U3816 ( .A1(n2383), .A2(n2167), .ZN(n3802) );
  NAND2_X1 U3817 ( .A1(n3803), .A2(b_2_), .ZN(n3674) );
  NOR2_X1 U3818 ( .A1(n2385), .A2(n2136), .ZN(n3803) );
  XOR2_X1 U3819 ( .A(n3804), .B(n3805), .Z(n3692) );
  XOR2_X1 U3820 ( .A(n3806), .B(n3807), .Z(n3804) );
  XNOR2_X1 U3821 ( .A(n3808), .B(n3809), .ZN(n3696) );
  XNOR2_X1 U3822 ( .A(n3810), .B(n3811), .ZN(n3809) );
  XNOR2_X1 U3823 ( .A(n3812), .B(n3813), .ZN(n3654) );
  NAND2_X1 U3824 ( .A1(n3814), .A2(n3815), .ZN(n3812) );
  XNOR2_X1 U3825 ( .A(n3816), .B(n3817), .ZN(n3700) );
  XNOR2_X1 U3826 ( .A(n3818), .B(n3819), .ZN(n3816) );
  XNOR2_X1 U3827 ( .A(n3820), .B(n3821), .ZN(n3704) );
  NAND2_X1 U3828 ( .A1(n3822), .A2(n3823), .ZN(n3820) );
  XNOR2_X1 U3829 ( .A(n3824), .B(n3825), .ZN(n3708) );
  XNOR2_X1 U3830 ( .A(n3826), .B(n3827), .ZN(n3824) );
  XNOR2_X1 U3831 ( .A(n3828), .B(n3829), .ZN(n3634) );
  NAND2_X1 U3832 ( .A1(n3830), .A2(n3831), .ZN(n3828) );
  XNOR2_X1 U3833 ( .A(n3832), .B(n3833), .ZN(n3712) );
  XNOR2_X1 U3834 ( .A(n3834), .B(n3835), .ZN(n3832) );
  NOR2_X1 U3835 ( .A1(n2143), .A2(n2136), .ZN(n2131) );
  INV_X1 U3836 ( .A(b_3_), .ZN(n2136) );
  XNOR2_X1 U3837 ( .A(n3836), .B(n3837), .ZN(n3719) );
  XNOR2_X1 U3838 ( .A(n3838), .B(n3839), .ZN(n3836) );
  XOR2_X1 U3839 ( .A(n3840), .B(n3841), .Z(n3723) );
  XNOR2_X1 U3840 ( .A(n3842), .B(n2150), .ZN(n3840) );
  INV_X1 U3841 ( .A(n3843), .ZN(n2150) );
  XNOR2_X1 U3842 ( .A(n3844), .B(n3845), .ZN(n3609) );
  XNOR2_X1 U3843 ( .A(n3846), .B(n3847), .ZN(n3844) );
  NAND2_X1 U3844 ( .A1(n3848), .A2(n3849), .ZN(n2124) );
  OR2_X1 U3845 ( .A1(n2273), .A2(n2272), .ZN(n3849) );
  AND2_X1 U3846 ( .A1(n3733), .A2(n3850), .ZN(n2272) );
  NAND2_X1 U3847 ( .A1(n3732), .A2(n3734), .ZN(n3850) );
  NAND2_X1 U3848 ( .A1(n3851), .A2(n3852), .ZN(n3734) );
  NAND2_X1 U3849 ( .A1(a_0_), .A2(b_2_), .ZN(n3852) );
  INV_X1 U3850 ( .A(n3853), .ZN(n3851) );
  XOR2_X1 U3851 ( .A(n3854), .B(n3855), .Z(n3732) );
  NOR2_X1 U3852 ( .A1(n3856), .A2(n2222), .ZN(n3855) );
  XOR2_X1 U3853 ( .A(n3857), .B(n2163), .Z(n3854) );
  NAND2_X1 U3854 ( .A1(a_0_), .A2(n3853), .ZN(n3733) );
  NAND2_X1 U3855 ( .A1(n3858), .A2(n3859), .ZN(n3853) );
  NAND2_X1 U3856 ( .A1(n3847), .A2(n3860), .ZN(n3859) );
  NAND2_X1 U3857 ( .A1(n3846), .A2(n3845), .ZN(n3860) );
  NOR2_X1 U3858 ( .A1(n2319), .A2(n2221), .ZN(n3847) );
  OR2_X1 U3859 ( .A1(n3845), .A2(n3846), .ZN(n3858) );
  AND2_X1 U3860 ( .A1(n3861), .A2(n3862), .ZN(n3846) );
  NAND2_X1 U3861 ( .A1(n3841), .A2(n3863), .ZN(n3862) );
  OR2_X1 U3862 ( .A1(n3842), .A2(n3843), .ZN(n3863) );
  XOR2_X1 U3863 ( .A(n3864), .B(n3865), .Z(n3841) );
  NOR2_X1 U3864 ( .A1(n2167), .A2(n2143), .ZN(n3865) );
  XOR2_X1 U3865 ( .A(n3866), .B(n3867), .Z(n3864) );
  NAND2_X1 U3866 ( .A1(n3843), .A2(n3842), .ZN(n3861) );
  NAND2_X1 U3867 ( .A1(n3868), .A2(n3869), .ZN(n3842) );
  NAND2_X1 U3868 ( .A1(n3839), .A2(n3870), .ZN(n3869) );
  NAND2_X1 U3869 ( .A1(n3838), .A2(n3837), .ZN(n3870) );
  NOR2_X1 U3870 ( .A1(n2143), .A2(n2221), .ZN(n3839) );
  OR2_X1 U3871 ( .A1(n3837), .A2(n3838), .ZN(n3868) );
  AND2_X1 U3872 ( .A1(n3752), .A2(n3871), .ZN(n3838) );
  NAND2_X1 U3873 ( .A1(n3751), .A2(n3753), .ZN(n3871) );
  NAND2_X1 U3874 ( .A1(n3872), .A2(n3873), .ZN(n3753) );
  NAND2_X1 U3875 ( .A1(b_2_), .A2(a_4_), .ZN(n3873) );
  INV_X1 U3876 ( .A(n3874), .ZN(n3872) );
  XOR2_X1 U3877 ( .A(n3875), .B(n3876), .Z(n3751) );
  NOR2_X1 U3878 ( .A1(n2108), .A2(n2167), .ZN(n3876) );
  XOR2_X1 U3879 ( .A(n3877), .B(n3878), .Z(n3875) );
  NAND2_X1 U3880 ( .A1(a_4_), .A2(n3874), .ZN(n3752) );
  NAND2_X1 U3881 ( .A1(n3879), .A2(n3880), .ZN(n3874) );
  NAND2_X1 U3882 ( .A1(n3835), .A2(n3881), .ZN(n3880) );
  NAND2_X1 U3883 ( .A1(n3834), .A2(n3833), .ZN(n3881) );
  NOR2_X1 U3884 ( .A1(n2221), .A2(n2108), .ZN(n3835) );
  OR2_X1 U3885 ( .A1(n3833), .A2(n3834), .ZN(n3879) );
  AND2_X1 U3886 ( .A1(n3830), .A2(n3882), .ZN(n3834) );
  NAND2_X1 U3887 ( .A1(n3829), .A2(n3831), .ZN(n3882) );
  NAND2_X1 U3888 ( .A1(n3883), .A2(n3884), .ZN(n3831) );
  NAND2_X1 U3889 ( .A1(a_6_), .A2(b_2_), .ZN(n3884) );
  INV_X1 U3890 ( .A(n3885), .ZN(n3883) );
  XOR2_X1 U3891 ( .A(n3886), .B(n3887), .Z(n3829) );
  NOR2_X1 U3892 ( .A1(n2073), .A2(n2167), .ZN(n3887) );
  XOR2_X1 U3893 ( .A(n3888), .B(n3889), .Z(n3886) );
  NAND2_X1 U3894 ( .A1(a_6_), .A2(n3885), .ZN(n3830) );
  NAND2_X1 U3895 ( .A1(n3890), .A2(n3891), .ZN(n3885) );
  NAND2_X1 U3896 ( .A1(n3827), .A2(n3892), .ZN(n3891) );
  NAND2_X1 U3897 ( .A1(n3826), .A2(n3825), .ZN(n3892) );
  NOR2_X1 U3898 ( .A1(n2221), .A2(n2073), .ZN(n3827) );
  OR2_X1 U3899 ( .A1(n3825), .A2(n3826), .ZN(n3890) );
  AND2_X1 U3900 ( .A1(n3822), .A2(n3893), .ZN(n3826) );
  NAND2_X1 U3901 ( .A1(n3821), .A2(n3823), .ZN(n3893) );
  NAND2_X1 U3902 ( .A1(n3894), .A2(n3895), .ZN(n3823) );
  NAND2_X1 U3903 ( .A1(b_2_), .A2(a_8_), .ZN(n3895) );
  INV_X1 U3904 ( .A(n3896), .ZN(n3894) );
  XOR2_X1 U3905 ( .A(n3897), .B(n3898), .Z(n3821) );
  XNOR2_X1 U3906 ( .A(n3899), .B(n3900), .ZN(n3898) );
  NAND2_X1 U3907 ( .A1(b_1_), .A2(a_9_), .ZN(n3897) );
  NAND2_X1 U3908 ( .A1(a_8_), .A2(n3896), .ZN(n3822) );
  NAND2_X1 U3909 ( .A1(n3901), .A2(n3902), .ZN(n3896) );
  NAND2_X1 U3910 ( .A1(n3819), .A2(n3903), .ZN(n3902) );
  NAND2_X1 U3911 ( .A1(n3818), .A2(n3817), .ZN(n3903) );
  NOR2_X1 U3912 ( .A1(n2221), .A2(n2215), .ZN(n3819) );
  OR2_X1 U3913 ( .A1(n3817), .A2(n3818), .ZN(n3901) );
  AND2_X1 U3914 ( .A1(n3814), .A2(n3904), .ZN(n3818) );
  NAND2_X1 U3915 ( .A1(n3813), .A2(n3815), .ZN(n3904) );
  NAND2_X1 U3916 ( .A1(n3905), .A2(n3906), .ZN(n3815) );
  NAND2_X1 U3917 ( .A1(b_2_), .A2(a_10_), .ZN(n3906) );
  INV_X1 U3918 ( .A(n3907), .ZN(n3905) );
  XOR2_X1 U3919 ( .A(n3908), .B(n3909), .Z(n3813) );
  NOR2_X1 U3920 ( .A1(n2212), .A2(n2167), .ZN(n3909) );
  XOR2_X1 U3921 ( .A(n3910), .B(n3911), .Z(n3908) );
  NAND2_X1 U3922 ( .A1(a_10_), .A2(n3907), .ZN(n3814) );
  NAND2_X1 U3923 ( .A1(n3912), .A2(n3913), .ZN(n3907) );
  NAND2_X1 U3924 ( .A1(n3811), .A2(n3914), .ZN(n3913) );
  OR2_X1 U3925 ( .A1(n3810), .A2(n3808), .ZN(n3914) );
  NOR2_X1 U3926 ( .A1(n2221), .A2(n2212), .ZN(n3811) );
  NAND2_X1 U3927 ( .A1(n3808), .A2(n3810), .ZN(n3912) );
  NAND2_X1 U3928 ( .A1(n3915), .A2(n3916), .ZN(n3810) );
  NAND2_X1 U3929 ( .A1(n3806), .A2(n3917), .ZN(n3916) );
  OR2_X1 U3930 ( .A1(n3805), .A2(n3807), .ZN(n3917) );
  NOR2_X1 U3931 ( .A1(n2221), .A2(n2000), .ZN(n3806) );
  NAND2_X1 U3932 ( .A1(n3805), .A2(n3807), .ZN(n3915) );
  NAND2_X1 U3933 ( .A1(n3918), .A2(n3919), .ZN(n3807) );
  NAND2_X1 U3934 ( .A1(n3920), .A2(b_2_), .ZN(n3919) );
  NOR2_X1 U3935 ( .A1(n3921), .A2(n2210), .ZN(n3920) );
  NOR2_X1 U3936 ( .A1(n3792), .A2(n3793), .ZN(n3921) );
  NAND2_X1 U3937 ( .A1(n3792), .A2(n3793), .ZN(n3918) );
  NAND2_X1 U3938 ( .A1(n3922), .A2(n3923), .ZN(n3793) );
  NAND2_X1 U3939 ( .A1(n3924), .A2(b_0_), .ZN(n3923) );
  NOR2_X1 U3940 ( .A1(n3925), .A2(n2208), .ZN(n3924) );
  NOR2_X1 U3941 ( .A1(n2380), .A2(n2167), .ZN(n3925) );
  NAND2_X1 U3942 ( .A1(n3926), .A2(b_1_), .ZN(n3922) );
  NOR2_X1 U3943 ( .A1(n3927), .A2(n2499), .ZN(n3926) );
  NOR2_X1 U3944 ( .A1(n2383), .A2(n3856), .ZN(n3927) );
  AND2_X1 U3945 ( .A1(n3928), .A2(b_1_), .ZN(n3792) );
  NOR2_X1 U3946 ( .A1(n2385), .A2(n2221), .ZN(n3928) );
  XOR2_X1 U3947 ( .A(n3929), .B(n3930), .Z(n3805) );
  XNOR2_X1 U3948 ( .A(n3931), .B(n3932), .ZN(n3930) );
  XOR2_X1 U3949 ( .A(n3933), .B(n3934), .Z(n3808) );
  XOR2_X1 U3950 ( .A(n3935), .B(n3936), .Z(n3933) );
  XNOR2_X1 U3951 ( .A(n3937), .B(n3938), .ZN(n3817) );
  XOR2_X1 U3952 ( .A(n3939), .B(n3940), .Z(n3937) );
  XOR2_X1 U3953 ( .A(n3941), .B(n3942), .Z(n3825) );
  XNOR2_X1 U3954 ( .A(n3943), .B(n3944), .ZN(n3942) );
  XOR2_X1 U3955 ( .A(n3945), .B(n3946), .Z(n3833) );
  XNOR2_X1 U3956 ( .A(n3947), .B(n3948), .ZN(n3946) );
  XNOR2_X1 U3957 ( .A(n3949), .B(n3950), .ZN(n3837) );
  XOR2_X1 U3958 ( .A(n3951), .B(n3952), .Z(n3949) );
  NOR2_X1 U3959 ( .A1(n2222), .A2(n2221), .ZN(n3843) );
  INV_X1 U3960 ( .A(b_2_), .ZN(n2221) );
  XNOR2_X1 U3961 ( .A(n3953), .B(n3954), .ZN(n3845) );
  NOR2_X1 U3962 ( .A1(n3955), .A2(n3956), .ZN(n3954) );
  INV_X1 U3963 ( .A(n3957), .ZN(n3956) );
  NOR2_X1 U3964 ( .A1(n3958), .A2(n3959), .ZN(n3955) );
  XNOR2_X1 U3965 ( .A(n3960), .B(n3961), .ZN(n2273) );
  NOR2_X1 U3966 ( .A1(n3962), .A2(n3963), .ZN(n3961) );
  INV_X1 U3967 ( .A(n3964), .ZN(n3963) );
  NOR2_X1 U3968 ( .A1(n3965), .A2(n3966), .ZN(n3962) );
  XNOR2_X1 U3969 ( .A(n2275), .B(n2179), .ZN(n3848) );
  NOR2_X1 U3970 ( .A1(n2228), .A2(n3856), .ZN(n2179) );
  AND2_X1 U3971 ( .A1(n2275), .A2(a_0_), .ZN(n2267) );
  NAND2_X1 U3972 ( .A1(n3964), .A2(n3967), .ZN(n2275) );
  NAND2_X1 U3973 ( .A1(n3968), .A2(n3960), .ZN(n3967) );
  NAND2_X1 U3974 ( .A1(n3969), .A2(n3970), .ZN(n3960) );
  NAND2_X1 U3975 ( .A1(n3971), .A2(a_2_), .ZN(n3970) );
  NOR2_X1 U3976 ( .A1(n3972), .A2(n3856), .ZN(n3971) );
  NOR2_X1 U3977 ( .A1(n2163), .A2(n3857), .ZN(n3972) );
  NAND2_X1 U3978 ( .A1(n2163), .A2(n3857), .ZN(n3969) );
  NAND2_X1 U3979 ( .A1(n3957), .A2(n3973), .ZN(n3857) );
  NAND2_X1 U3980 ( .A1(n3974), .A2(n3953), .ZN(n3973) );
  NAND2_X1 U3981 ( .A1(n3975), .A2(n3976), .ZN(n3953) );
  NAND2_X1 U3982 ( .A1(n3977), .A2(a_3_), .ZN(n3976) );
  NOR2_X1 U3983 ( .A1(n3978), .A2(n2167), .ZN(n3977) );
  NOR2_X1 U3984 ( .A1(n3866), .A2(n3867), .ZN(n3978) );
  NAND2_X1 U3985 ( .A1(n3866), .A2(n3867), .ZN(n3975) );
  NAND2_X1 U3986 ( .A1(n3979), .A2(n3980), .ZN(n3867) );
  NAND2_X1 U3987 ( .A1(n3950), .A2(n3981), .ZN(n3980) );
  OR2_X1 U3988 ( .A1(n3951), .A2(n3952), .ZN(n3981) );
  NOR2_X1 U3989 ( .A1(n2167), .A2(n2220), .ZN(n3950) );
  NAND2_X1 U3990 ( .A1(n3952), .A2(n3951), .ZN(n3979) );
  NAND2_X1 U3991 ( .A1(n3982), .A2(n3983), .ZN(n3951) );
  NAND2_X1 U3992 ( .A1(n3984), .A2(b_1_), .ZN(n3983) );
  NOR2_X1 U3993 ( .A1(n3985), .A2(n2108), .ZN(n3984) );
  NOR2_X1 U3994 ( .A1(n3878), .A2(n3877), .ZN(n3985) );
  NAND2_X1 U3995 ( .A1(n3878), .A2(n3877), .ZN(n3982) );
  NAND2_X1 U3996 ( .A1(n3986), .A2(n3987), .ZN(n3877) );
  NAND2_X1 U3997 ( .A1(n3945), .A2(n3988), .ZN(n3987) );
  NAND2_X1 U3998 ( .A1(n3948), .A2(n3947), .ZN(n3988) );
  INV_X1 U3999 ( .A(n3989), .ZN(n3947) );
  INV_X1 U4000 ( .A(n3990), .ZN(n3948) );
  NOR2_X1 U4001 ( .A1(n2167), .A2(n2217), .ZN(n3945) );
  NAND2_X1 U4002 ( .A1(n3989), .A2(n3990), .ZN(n3986) );
  NAND2_X1 U4003 ( .A1(n3991), .A2(n3992), .ZN(n3990) );
  NAND2_X1 U4004 ( .A1(n3993), .A2(b_1_), .ZN(n3992) );
  NOR2_X1 U4005 ( .A1(n3994), .A2(n2073), .ZN(n3993) );
  NOR2_X1 U4006 ( .A1(n3888), .A2(n3889), .ZN(n3994) );
  NAND2_X1 U4007 ( .A1(n3888), .A2(n3889), .ZN(n3991) );
  NAND2_X1 U4008 ( .A1(n3995), .A2(n3996), .ZN(n3889) );
  NAND2_X1 U4009 ( .A1(n3941), .A2(n3997), .ZN(n3996) );
  OR2_X1 U4010 ( .A1(n3944), .A2(n3943), .ZN(n3997) );
  NOR2_X1 U4011 ( .A1(n2167), .A2(n2059), .ZN(n3941) );
  NAND2_X1 U4012 ( .A1(n3943), .A2(n3944), .ZN(n3995) );
  NAND2_X1 U4013 ( .A1(n3998), .A2(n3999), .ZN(n3944) );
  NAND2_X1 U4014 ( .A1(n4000), .A2(b_1_), .ZN(n3999) );
  NOR2_X1 U4015 ( .A1(n4001), .A2(n2215), .ZN(n4000) );
  NOR2_X1 U4016 ( .A1(n3900), .A2(n3899), .ZN(n4001) );
  NAND2_X1 U4017 ( .A1(n3900), .A2(n3899), .ZN(n3998) );
  NAND2_X1 U4018 ( .A1(n4002), .A2(n4003), .ZN(n3899) );
  NAND2_X1 U4019 ( .A1(n3938), .A2(n4004), .ZN(n4003) );
  OR2_X1 U4020 ( .A1(n3940), .A2(n3939), .ZN(n4004) );
  NOR2_X1 U4021 ( .A1(n2167), .A2(n2214), .ZN(n3938) );
  NAND2_X1 U4022 ( .A1(n3939), .A2(n3940), .ZN(n4002) );
  NAND2_X1 U4023 ( .A1(n4005), .A2(n4006), .ZN(n3940) );
  NAND2_X1 U4024 ( .A1(n4007), .A2(b_1_), .ZN(n4006) );
  NOR2_X1 U4025 ( .A1(n4008), .A2(n2212), .ZN(n4007) );
  NOR2_X1 U4026 ( .A1(n3910), .A2(n3911), .ZN(n4008) );
  NAND2_X1 U4027 ( .A1(n3910), .A2(n3911), .ZN(n4005) );
  NAND2_X1 U4028 ( .A1(n4009), .A2(n4010), .ZN(n3911) );
  NAND2_X1 U4029 ( .A1(n3934), .A2(n4011), .ZN(n4010) );
  OR2_X1 U4030 ( .A1(n3935), .A2(n3936), .ZN(n4011) );
  NOR2_X1 U4031 ( .A1(n2167), .A2(n2000), .ZN(n3934) );
  NAND2_X1 U4032 ( .A1(n3936), .A2(n3935), .ZN(n4009) );
  NAND2_X1 U4033 ( .A1(n4012), .A2(n3932), .ZN(n3935) );
  NAND2_X1 U4034 ( .A1(n4013), .A2(b_0_), .ZN(n3932) );
  NOR2_X1 U4035 ( .A1(n2385), .A2(n2167), .ZN(n4013) );
  INV_X1 U4036 ( .A(n2209), .ZN(n2385) );
  NOR2_X1 U4037 ( .A1(n2208), .A2(n2499), .ZN(n2209) );
  INV_X1 U4038 ( .A(a_15_), .ZN(n2208) );
  NAND2_X1 U4039 ( .A1(n3929), .A2(n3931), .ZN(n4012) );
  NOR2_X1 U4040 ( .A1(n2167), .A2(n2210), .ZN(n3931) );
  NOR2_X1 U4041 ( .A1(n3856), .A2(n2499), .ZN(n3929) );
  INV_X1 U4042 ( .A(a_14_), .ZN(n2499) );
  NOR2_X1 U4043 ( .A1(n3856), .A2(n2210), .ZN(n3936) );
  INV_X1 U4044 ( .A(a_13_), .ZN(n2210) );
  NOR2_X1 U4045 ( .A1(n3856), .A2(n2000), .ZN(n3910) );
  INV_X1 U4046 ( .A(a_12_), .ZN(n2000) );
  NOR2_X1 U4047 ( .A1(n3856), .A2(n2212), .ZN(n3939) );
  INV_X1 U4048 ( .A(a_11_), .ZN(n2212) );
  NOR2_X1 U4049 ( .A1(n3856), .A2(n2214), .ZN(n3900) );
  INV_X1 U4050 ( .A(a_10_), .ZN(n2214) );
  NOR2_X1 U4051 ( .A1(n3856), .A2(n2215), .ZN(n3943) );
  INV_X1 U4052 ( .A(a_9_), .ZN(n2215) );
  NOR2_X1 U4053 ( .A1(n3856), .A2(n2059), .ZN(n3888) );
  INV_X1 U4054 ( .A(a_8_), .ZN(n2059) );
  NOR2_X1 U4055 ( .A1(n3856), .A2(n2073), .ZN(n3989) );
  INV_X1 U4056 ( .A(a_7_), .ZN(n2073) );
  NOR2_X1 U4057 ( .A1(n3856), .A2(n2217), .ZN(n3878) );
  INV_X1 U4058 ( .A(a_6_), .ZN(n2217) );
  NOR2_X1 U4059 ( .A1(n3856), .A2(n2108), .ZN(n3952) );
  INV_X1 U4060 ( .A(a_5_), .ZN(n2108) );
  NOR2_X1 U4061 ( .A1(n3856), .A2(n2220), .ZN(n3866) );
  INV_X1 U4062 ( .A(a_4_), .ZN(n2220) );
  OR2_X1 U4063 ( .A1(n3958), .A2(a_2_), .ZN(n3974) );
  NAND2_X1 U4064 ( .A1(n3959), .A2(n3958), .ZN(n3957) );
  NOR2_X1 U4065 ( .A1(n2143), .A2(n3856), .ZN(n3958) );
  INV_X1 U4066 ( .A(a_3_), .ZN(n2143) );
  NOR2_X1 U4067 ( .A1(n2167), .A2(n2222), .ZN(n3959) );
  INV_X1 U4068 ( .A(a_2_), .ZN(n2222) );
  NOR2_X1 U4069 ( .A1(n2319), .A2(n2167), .ZN(n2163) );
  OR2_X1 U4070 ( .A1(n3965), .A2(a_0_), .ZN(n3968) );
  NAND2_X1 U4071 ( .A1(n3966), .A2(n3965), .ZN(n3964) );
  NOR2_X1 U4072 ( .A1(n2319), .A2(n3856), .ZN(n3965) );
  INV_X1 U4073 ( .A(b_0_), .ZN(n3856) );
  INV_X1 U4074 ( .A(a_1_), .ZN(n2319) );
  NOR2_X1 U4075 ( .A1(n2167), .A2(n2228), .ZN(n3966) );
  INV_X1 U4076 ( .A(a_0_), .ZN(n2228) );
  INV_X1 U4077 ( .A(b_1_), .ZN(n2167) );
endmodule

