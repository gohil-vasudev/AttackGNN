module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX647, n3527, WX649, n3525,
         WX653, n3521, WX655, n3519, WX657, n3517, WX658, WX659, n3515, WX661,
         n3513, WX663, n3511, WX665, n3509, WX666, WX667, n3507, WX669, n3505,
         WX671, n3503, WX673, n3501, WX674, WX675, n3499, WX677, n3497, WX679,
         n3495, WX681, n3493, WX683, n3491, WX685, n3489, WX686, WX689, n3485,
         WX691, n3483, WX693, n3481, WX695, n3479, WX697, n3477, WX699, n3475,
         WX701, n3473, WX703, n3471, WX705, n3469, WX707, n3467, WX708, WX709,
         WX710, WX711, WX712, WX713, WX714, WX715, WX716, WX717, WX718, WX719,
         WX720, WX721, WX722, WX724, WX725, WX726, WX727, WX728, WX729, WX730,
         WX731, WX732, WX733, WX734, WX735, WX736, WX737, WX738, WX739, WX740,
         WX741, WX742, WX743, WX744, WX745, WX746, WX747, WX748, WX749, WX750,
         WX751, WX752, WX753, WX754, WX755, WX756, WX757, WX758, WX760, WX761,
         WX762, WX763, WX764, WX765, WX766, WX767, WX768, WX769, WX770, WX771,
         WX772, WX773, WX774, WX775, WX776, WX777, WX778, WX779, WX780, WX781,
         WX782, WX783, WX784, WX785, WX786, WX787, WX788, WX789, WX790, WX791,
         WX792, WX793, WX794, WX796, WX797, WX798, WX799, WX800, WX801, WX802,
         WX803, WX804, WX805, WX806, WX807, WX808, WX809, WX810, WX811, WX812,
         WX813, WX814, WX815, WX816, WX817, WX818, WX819, WX820, WX821, WX822,
         WX823, WX824, WX825, WX826, WX827, WX828, WX829, WX830, WX832, WX833,
         WX834, WX835, WX836, WX837, WX838, WX839, WX840, WX841, WX842, WX843,
         WX844, WX845, WX846, WX847, WX848, WX849, WX850, WX851, WX852, WX853,
         WX854, WX855, WX856, WX857, WX858, WX859, WX860, WX861, WX862, WX863,
         WX864, WX865, WX866, WX868, WX869, WX870, WX871, WX872, WX873, WX874,
         WX875, WX876, WX877, WX878, WX879, WX880, WX881, WX882, WX883, WX884,
         WX885, WX886, WX887, WX888, WX889, WX890, WX891, WX892, WX893, WX894,
         WX895, WX896, WX897, WX898, WX899, WX1264, DFF_160_n1, WX1266, WX1268,
         DFF_162_n1, WX1270, WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276,
         DFF_166_n1, WX1278, DFF_167_n1, WX1280, DFF_168_n1, WX1282,
         DFF_169_n1, WX1284, WX1286, DFF_171_n1, WX1288, DFF_172_n1, WX1290,
         DFF_173_n1, WX1292, DFF_174_n1, WX1294, DFF_175_n1, WX1296,
         DFF_176_n1, WX1298, DFF_177_n1, WX1300, DFF_178_n1, WX1302, WX1304,
         DFF_180_n1, WX1306, DFF_181_n1, WX1308, DFF_182_n1, WX1310,
         DFF_183_n1, WX1312, DFF_184_n1, WX1314, DFF_185_n1, WX1316,
         DFF_186_n1, WX1318, DFF_187_n1, WX1320, DFF_188_n1, WX1322,
         DFF_189_n1, WX1324, DFF_190_n1, WX1326, DFF_191_n1, WX1778, n8702,
         n8701, n8700, n8699, n8696, n8695, n8694, n8693, n8692, n8691, n8690,
         n8689, n8688, n8687, n8686, n8685, n8684, n8683, n8682, n8681, n8680,
         n8677, n8676, n8675, n8674, n8673, n8672, n8671, WX1839, n8670,
         WX1937, n8669, WX1939, n8668, WX1941, n8667, WX1943, n8666, WX1945,
         n8665, WX1947, n8664, WX1949, n8663, WX1951, n8662, WX1953, n8661,
         WX1955, WX1957, n8658, WX1959, n8657, WX1961, n8656, WX1963, n8655,
         WX1965, n8654, WX1967, n8653, WX1969, WX1970, WX1971, WX1972, WX1973,
         WX1974, WX1975, WX1976, WX1977, WX1978, WX1979, WX1980, WX1981,
         WX1982, WX1983, WX1984, WX1985, WX1986, WX1987, WX1988, WX1989,
         WX1990, WX1991, WX1993, WX1994, WX1995, WX1996, WX1997, WX1998,
         WX1999, WX2000, WX2001, WX2002, WX2003, WX2004, WX2005, WX2006,
         WX2007, WX2008, WX2009, WX2010, WX2011, WX2012, WX2013, WX2014,
         WX2015, WX2016, WX2017, WX2018, WX2019, WX2020, WX2021, WX2022,
         WX2023, WX2024, WX2025, WX2026, WX2027, WX2029, WX2030, WX2031,
         WX2032, WX2033, WX2034, WX2035, WX2036, WX2037, WX2038, WX2039,
         WX2040, WX2041, WX2042, WX2043, WX2044, WX2045, WX2046, WX2047,
         WX2048, WX2049, WX2050, WX2051, WX2052, WX2053, WX2054, WX2055,
         WX2056, WX2057, WX2058, WX2059, WX2060, WX2061, WX2062, WX2063,
         WX2065, WX2066, WX2067, WX2068, WX2069, WX2070, WX2071, WX2072,
         WX2073, WX2074, WX2075, WX2076, WX2077, WX2078, WX2079, WX2080,
         WX2081, WX2082, WX2083, WX2084, WX2085, WX2086, WX2087, WX2088,
         WX2089, WX2090, WX2091, WX2092, WX2093, WX2094, WX2095, WX2096,
         WX2097, WX2098, WX2099, WX2101, WX2102, WX2103, WX2104, WX2105,
         WX2106, WX2107, WX2108, WX2109, WX2110, WX2111, WX2112, WX2113,
         WX2114, WX2115, WX2116, WX2117, WX2118, WX2119, WX2120, WX2121,
         WX2122, WX2123, WX2124, WX2125, WX2126, WX2127, WX2128, WX2129,
         WX2130, WX2131, WX2132, WX2133, WX2134, WX2135, WX2137, WX2138,
         WX2139, WX2140, WX2141, WX2142, WX2143, WX2144, WX2145, WX2146,
         WX2147, WX2148, WX2149, WX2150, WX2151, WX2152, WX2153, WX2154,
         WX2155, WX2156, WX2157, WX2158, WX2159, WX2160, WX2161, WX2162,
         WX2163, WX2164, WX2165, WX2166, WX2167, WX2168, WX2169, WX2170,
         WX2171, WX2173, WX2174, WX2175, WX2176, WX2177, WX2178, WX2179,
         WX2180, WX2181, WX2182, WX2183, WX2184, WX2185, WX2186, WX2187,
         WX2188, WX2189, WX2190, WX2191, WX2192, WX2557, DFF_352_n1, WX2559,
         DFF_353_n1, WX2561, DFF_354_n1, WX2563, DFF_355_n1, WX2565,
         DFF_356_n1, WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571, WX2573,
         DFF_360_n1, WX2575, DFF_361_n1, WX2577, DFF_362_n1, WX2579,
         DFF_363_n1, WX2581, DFF_364_n1, WX2583, DFF_365_n1, WX2585,
         DFF_366_n1, WX2587, DFF_367_n1, WX2589, DFF_368_n1, WX2591,
         DFF_369_n1, WX2593, DFF_370_n1, WX2595, DFF_371_n1, WX2597,
         DFF_372_n1, WX2599, DFF_373_n1, WX2601, DFF_374_n1, WX2603,
         DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609, DFF_378_n1, WX2611,
         DFF_379_n1, WX2613, DFF_380_n1, WX2615, DFF_381_n1, WX2617,
         DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644, n8643, n8642, n8641,
         n8640, n8639, n8638, n8637, n8636, n8635, n8632, n8631, n8630, n8629,
         n8628, n8627, n8626, n8625, n8624, n8623, n8622, n8621, n8620, n8619,
         n8618, n8617, n8616, n8613, WX3132, n8612, WX3230, n8611, WX3232,
         n8610, WX3234, n8609, WX3236, n8608, WX3238, n8607, WX3240, n8606,
         WX3242, n8605, WX3244, n8604, WX3246, n8603, WX3248, n8602, WX3250,
         n8601, WX3252, n8600, WX3254, n8599, WX3256, n8598, WX3258, n8597,
         WX3260, WX3262, WX3263, WX3264, WX3265, WX3266, WX3267, WX3268,
         WX3269, WX3270, WX3271, WX3272, WX3273, WX3274, WX3275, WX3276,
         WX3277, WX3278, WX3279, WX3280, WX3281, WX3282, WX3283, WX3284,
         WX3285, WX3286, WX3287, WX3288, WX3289, WX3290, WX3291, WX3292,
         WX3293, WX3294, WX3295, WX3296, WX3298, WX3299, WX3300, WX3301,
         WX3302, WX3303, WX3304, WX3305, WX3306, WX3307, WX3308, WX3309,
         WX3310, WX3311, WX3312, WX3313, WX3314, WX3315, WX3316, WX3317,
         WX3318, WX3319, WX3320, WX3321, WX3322, WX3323, WX3324, WX3325,
         WX3326, WX3327, WX3328, WX3329, WX3330, WX3331, WX3332, WX3334,
         WX3335, WX3336, WX3337, WX3338, WX3339, WX3340, WX3341, WX3342,
         WX3343, WX3344, WX3345, WX3346, WX3347, WX3348, WX3349, WX3350,
         WX3351, WX3352, WX3353, WX3354, WX3355, WX3356, WX3357, WX3358,
         WX3359, WX3360, WX3361, WX3362, WX3363, WX3364, WX3365, WX3366,
         WX3367, WX3368, WX3370, WX3371, WX3372, WX3373, WX3374, WX3375,
         WX3376, WX3377, WX3378, WX3379, WX3380, WX3381, WX3382, WX3383,
         WX3384, WX3385, WX3386, WX3387, WX3388, WX3389, WX3390, WX3391,
         WX3392, WX3393, WX3394, WX3395, WX3396, WX3397, WX3398, WX3399,
         WX3400, WX3401, WX3402, WX3403, WX3404, WX3406, WX3407, WX3408,
         WX3409, WX3410, WX3411, WX3412, WX3413, WX3414, WX3415, WX3416,
         WX3417, WX3418, WX3419, WX3420, WX3421, WX3422, WX3423, WX3424,
         WX3425, WX3426, WX3427, WX3428, WX3429, WX3430, WX3431, WX3432,
         WX3433, WX3434, WX3435, WX3436, WX3437, WX3438, WX3440, WX3441,
         WX3442, WX3443, WX3444, WX3445, WX3446, WX3447, WX3448, WX3449,
         WX3450, WX3451, WX3452, WX3453, WX3454, WX3455, WX3456, WX3457,
         WX3458, WX3459, WX3460, WX3461, WX3462, WX3463, WX3464, WX3465,
         WX3466, WX3467, WX3468, WX3469, WX3470, WX3471, WX3472, WX3474,
         WX3475, WX3476, WX3477, WX3478, WX3479, WX3480, WX3481, WX3482,
         WX3483, WX3484, WX3485, WX3850, DFF_544_n1, WX3852, DFF_545_n1,
         WX3854, DFF_546_n1, WX3856, DFF_547_n1, WX3858, DFF_548_n1, WX3860,
         DFF_549_n1, WX3862, DFF_550_n1, WX3864, DFF_551_n1, WX3866,
         DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872, DFF_555_n1, WX3874,
         DFF_556_n1, WX3876, DFF_557_n1, WX3878, DFF_558_n1, WX3880,
         DFF_559_n1, WX3882, DFF_560_n1, WX3884, DFF_561_n1, WX3886,
         DFF_562_n1, WX3888, DFF_563_n1, WX3890, DFF_564_n1, WX3892,
         DFF_565_n1, WX3894, DFF_566_n1, WX3896, DFF_567_n1, WX3898,
         DFF_568_n1, WX3900, DFF_569_n1, WX3902, DFF_570_n1, WX3904, WX3906,
         DFF_572_n1, WX3908, DFF_573_n1, WX3910, DFF_574_n1, WX3912,
         DFF_575_n1, WX4364, n8586, n8585, n8584, n8583, n8582, n8581, n8580,
         n8579, n8578, n8577, n8576, n8573, n8572, n8571, n8570, n8569, n8568,
         n8567, n8566, n8565, n8564, n8563, n8562, n8561, n8560, n8559, n8558,
         n8555, WX4425, n8554, WX4523, n8553, WX4525, n8552, WX4527, n8551,
         WX4529, n8550, WX4531, n8549, WX4533, n8548, WX4535, n8547, WX4537,
         n8546, WX4539, n8545, WX4541, n8544, WX4543, n8543, WX4545, n8542,
         WX4547, n8541, WX4549, n8540, WX4551, WX4553, n8537, WX4555, WX4556,
         WX4557, WX4558, WX4559, WX4560, WX4561, WX4562, WX4563, WX4564,
         WX4565, WX4566, WX4567, WX4568, WX4569, WX4570, WX4571, WX4572,
         WX4573, WX4574, WX4575, WX4576, WX4577, WX4578, WX4579, WX4580,
         WX4581, WX4582, WX4583, WX4584, WX4585, WX4587, WX4588, WX4589,
         WX4590, WX4591, WX4592, WX4593, WX4594, WX4595, WX4596, WX4597,
         WX4598, WX4599, WX4600, WX4601, WX4602, WX4603, WX4604, WX4605,
         WX4606, WX4607, WX4608, WX4609, WX4610, WX4611, WX4612, WX4613,
         WX4614, WX4615, WX4616, WX4617, WX4618, WX4619, WX4621, WX4622,
         WX4623, WX4624, WX4625, WX4626, WX4627, WX4628, WX4629, WX4630,
         WX4631, WX4632, WX4633, WX4634, WX4635, WX4636, WX4637, WX4638,
         WX4639, WX4640, WX4641, WX4642, WX4643, WX4644, WX4645, WX4646,
         WX4647, WX4648, WX4649, WX4650, WX4651, WX4652, WX4653, WX4655,
         WX4656, WX4657, WX4658, WX4659, WX4660, WX4661, WX4662, WX4663,
         WX4664, WX4665, WX4666, WX4667, WX4668, WX4669, WX4670, WX4671,
         WX4672, WX4673, WX4674, WX4675, WX4676, WX4677, WX4678, WX4679,
         WX4680, WX4681, WX4682, WX4683, WX4684, WX4685, WX4686, WX4687,
         WX4689, WX4690, WX4691, WX4692, WX4693, WX4694, WX4695, WX4696,
         WX4697, WX4698, WX4699, WX4700, WX4701, WX4702, WX4703, WX4704,
         WX4705, WX4706, WX4707, WX4708, WX4709, WX4710, WX4711, WX4712,
         WX4713, WX4714, WX4715, WX4716, WX4717, WX4718, WX4719, WX4720,
         WX4721, WX4723, WX4724, WX4725, WX4726, WX4727, WX4728, WX4729,
         WX4730, WX4731, WX4732, WX4733, WX4734, WX4735, WX4736, WX4737,
         WX4738, WX4739, WX4740, WX4741, WX4742, WX4743, WX4744, WX4745,
         WX4746, WX4747, WX4748, WX4749, WX4750, WX4751, WX4752, WX4753,
         WX4754, WX4755, WX4757, WX4758, WX4759, WX4760, WX4761, WX4762,
         WX4763, WX4764, WX4765, WX4766, WX4767, WX4768, WX4769, WX4770,
         WX4771, WX4772, WX4773, WX4774, WX4775, WX4776, WX4777, WX4778,
         WX5143, DFF_736_n1, WX5145, DFF_737_n1, WX5147, DFF_738_n1, WX5149,
         DFF_739_n1, WX5151, DFF_740_n1, WX5153, WX5155, DFF_742_n1, WX5157,
         DFF_743_n1, WX5159, DFF_744_n1, WX5161, DFF_745_n1, WX5163,
         DFF_746_n1, WX5165, DFF_747_n1, WX5167, DFF_748_n1, WX5169,
         DFF_749_n1, WX5171, DFF_750_n1, WX5173, DFF_751_n1, WX5175,
         DFF_752_n1, WX5177, DFF_753_n1, WX5179, DFF_754_n1, WX5181,
         DFF_755_n1, WX5183, DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189,
         DFF_759_n1, WX5191, DFF_760_n1, WX5193, DFF_761_n1, WX5195,
         DFF_762_n1, WX5197, DFF_763_n1, WX5199, DFF_764_n1, WX5201,
         DFF_765_n1, WX5203, DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528,
         n8527, n8526, n8525, n8524, n8523, n8520, n8519, n8518, n8517, n8516,
         n8515, n8514, n8513, n8512, n8511, n8510, n8509, n8508, n8507, n8506,
         n8505, n8502, n8501, n8500, n8499, n8498, n8497, WX5718, n8496,
         WX5816, n8495, WX5818, n8494, WX5820, n8493, WX5822, n8492, WX5824,
         n8491, WX5826, n8490, WX5828, n8489, WX5830, n8488, WX5832, n8487,
         WX5834, WX5836, n8484, WX5838, n8483, WX5840, n8482, WX5842, n8481,
         WX5844, n8480, WX5846, n8479, WX5848, WX5849, WX5850, WX5851, WX5852,
         WX5853, WX5854, WX5855, WX5856, WX5857, WX5858, WX5859, WX5860,
         WX5861, WX5862, WX5863, WX5864, WX5865, WX5866, WX5867, WX5868,
         WX5870, WX5871, WX5872, WX5873, WX5874, WX5875, WX5876, WX5877,
         WX5878, WX5879, WX5880, WX5881, WX5882, WX5883, WX5884, WX5885,
         WX5886, WX5887, WX5888, WX5889, WX5890, WX5891, WX5892, WX5893,
         WX5894, WX5895, WX5896, WX5897, WX5898, WX5899, WX5900, WX5901,
         WX5902, WX5904, WX5905, WX5906, WX5907, WX5908, WX5909, WX5910,
         WX5911, WX5912, WX5913, WX5914, WX5915, WX5916, WX5917, WX5918,
         WX5919, WX5920, WX5921, WX5922, WX5923, WX5924, WX5925, WX5926,
         WX5927, WX5928, WX5929, WX5930, WX5931, WX5932, WX5933, WX5934,
         WX5935, WX5936, WX5938, WX5939, WX5940, WX5941, WX5942, WX5943,
         WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950, WX5951,
         WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958, WX5959,
         WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966, WX5967,
         WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975, WX5976,
         WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983, WX5984,
         WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991, WX5992,
         WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999, WX6000,
         WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008, WX6009,
         WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016, WX6017,
         WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024, WX6025,
         WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032, WX6033,
         WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041, WX6042,
         WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049, WX6050,
         WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057, WX6058,
         WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065, WX6066,
         WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438, DFF_929_n1,
         WX6440, DFF_930_n1, WX6442, DFF_931_n1, WX6444, DFF_932_n1, WX6446,
         DFF_933_n1, WX6448, DFF_934_n1, WX6450, DFF_935_n1, WX6452,
         DFF_936_n1, WX6454, DFF_937_n1, WX6456, DFF_938_n1, WX6458,
         DFF_939_n1, WX6460, DFF_940_n1, WX6462, DFF_941_n1, WX6464,
         DFF_942_n1, WX6466, DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472,
         DFF_946_n1, WX6474, DFF_947_n1, WX6476, DFF_948_n1, WX6478,
         DFF_949_n1, WX6480, DFF_950_n1, WX6482, DFF_951_n1, WX6484,
         DFF_952_n1, WX6486, DFF_953_n1, WX6488, DFF_954_n1, WX6490,
         DFF_955_n1, WX6492, DFF_956_n1, WX6494, DFF_957_n1, WX6496,
         DFF_958_n1, WX6498, DFF_959_n1, WX6950, n8470, n8467, n8466, n8465,
         n8464, n8463, n8462, n8461, n8460, n8459, n8458, n8457, n8456, n8455,
         n8454, n8453, n8452, n8449, n8448, n8447, n8446, n8445, n8444, n8443,
         n8442, n8441, n8440, n8439, WX7011, n8438, WX7109, n8437, WX7111,
         n8436, WX7113, n8435, WX7115, n8434, WX7117, WX7119, n8431, WX7121,
         n8430, WX7123, n8429, WX7125, n8428, WX7127, n8427, WX7129, n8426,
         WX7131, n8425, WX7133, n8424, WX7135, n8423, WX7137, n8422, WX7139,
         n8421, WX7141, WX7142, WX7143, WX7144, WX7145, WX7146, WX7147, WX7148,
         WX7149, WX7150, WX7151, WX7153, WX7154, WX7155, WX7156, WX7157,
         WX7158, WX7159, WX7160, WX7161, WX7162, WX7163, WX7164, WX7165,
         WX7166, WX7167, WX7168, WX7169, WX7170, WX7171, WX7172, WX7173,
         WX7174, WX7175, WX7176, WX7177, WX7178, WX7179, WX7180, WX7181,
         WX7182, WX7183, WX7184, WX7185, WX7187, WX7188, WX7189, WX7190,
         WX7191, WX7192, WX7193, WX7194, WX7195, WX7196, WX7197, WX7198,
         WX7199, WX7200, WX7201, WX7202, WX7203, WX7204, WX7205, WX7206,
         WX7207, WX7208, WX7209, WX7210, WX7211, WX7212, WX7213, WX7214,
         WX7215, WX7216, WX7217, WX7218, WX7219, WX7221, WX7222, WX7223,
         WX7224, WX7225, WX7226, WX7227, WX7228, WX7229, WX7230, WX7231,
         WX7232, WX7233, WX7234, WX7235, WX7236, WX7237, WX7238, WX7239,
         WX7240, WX7241, WX7242, WX7243, WX7244, WX7245, WX7246, WX7247,
         WX7248, WX7249, WX7250, WX7251, WX7252, WX7253, WX7255, WX7256,
         WX7257, WX7258, WX7259, WX7260, WX7261, WX7262, WX7263, WX7264,
         WX7265, WX7266, WX7267, WX7268, WX7269, WX7270, WX7271, WX7272,
         WX7273, WX7274, WX7275, WX7276, WX7277, WX7278, WX7279, WX7280,
         WX7281, WX7282, WX7283, WX7284, WX7285, WX7286, WX7287, WX7289,
         WX7290, WX7291, WX7292, WX7293, WX7294, WX7295, WX7296, WX7297,
         WX7298, WX7299, WX7300, WX7301, WX7302, WX7303, WX7304, WX7305,
         WX7306, WX7307, WX7308, WX7309, WX7310, WX7311, WX7312, WX7313,
         WX7314, WX7315, WX7316, WX7317, WX7318, WX7319, WX7320, WX7321,
         WX7323, WX7324, WX7325, WX7326, WX7327, WX7328, WX7329, WX7330,
         WX7331, WX7332, WX7333, WX7334, WX7335, WX7336, WX7337, WX7338,
         WX7339, WX7340, WX7341, WX7342, WX7343, WX7344, WX7345, WX7346,
         WX7347, WX7348, WX7349, WX7350, WX7351, WX7352, WX7353, WX7354,
         WX7355, WX7357, WX7358, WX7359, WX7360, WX7361, WX7362, WX7363,
         WX7364, WX7729, DFF_1120_n1, WX7731, DFF_1121_n1, WX7733, DFF_1122_n1,
         WX7735, DFF_1123_n1, WX7737, DFF_1124_n1, WX7739, DFF_1125_n1, WX7741,
         DFF_1126_n1, WX7743, DFF_1127_n1, WX7745, DFF_1128_n1, WX7747,
         DFF_1129_n1, WX7749, DFF_1130_n1, WX7751, DFF_1131_n1, WX7753, WX7755,
         DFF_1133_n1, WX7757, DFF_1134_n1, WX7759, DFF_1135_n1, WX7761,
         DFF_1136_n1, WX7763, DFF_1137_n1, WX7765, DFF_1138_n1, WX7767,
         DFF_1139_n1, WX7769, DFF_1140_n1, WX7771, DFF_1141_n1, WX7773,
         DFF_1142_n1, WX7775, DFF_1143_n1, WX7777, DFF_1144_n1, WX7779,
         DFF_1145_n1, WX7781, DFF_1146_n1, WX7783, DFF_1147_n1, WX7785,
         DFF_1148_n1, WX7787, WX7789, DFF_1150_n1, WX7791, DFF_1151_n1, WX8243,
         n8411, n8410, n8409, n8408, n8407, n8406, n8405, n8404, n8403, n8402,
         n8401, n8400, n8399, n8396, n8395, n8394, n8393, n8392, n8391, n8390,
         n8389, n8388, n8387, n8386, n8385, n8384, n8383, n8382, n8381, WX8304,
         WX8402, n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410,
         n8374, WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370,
         WX8420, n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428,
         n8365, WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438,
         WX8439, WX8440, WX8441, WX8442, WX8443, WX8444, WX8445, WX8446,
         WX8447, WX8448, WX8449, WX8450, WX8451, WX8452, WX8453, WX8454,
         WX8455, WX8456, WX8457, WX8458, WX8459, WX8460, WX8461, WX8462,
         WX8463, WX8464, WX8465, WX8466, WX8467, WX8468, WX8470, WX8471,
         WX8472, WX8473, WX8474, WX8475, WX8476, WX8477, WX8478, WX8479,
         WX8480, WX8481, WX8482, WX8483, WX8484, WX8485, WX8486, WX8487,
         WX8488, WX8489, WX8490, WX8491, WX8492, WX8493, WX8494, WX8495,
         WX8496, WX8497, WX8498, WX8499, WX8500, WX8501, WX8502, WX8504,
         WX8505, WX8506, WX8507, WX8508, WX8509, WX8510, WX8511, WX8512,
         WX8513, WX8514, WX8515, WX8516, WX8517, WX8518, WX8519, WX8520,
         WX8521, WX8522, WX8523, WX8524, WX8525, WX8526, WX8527, WX8528,
         WX8529, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535, WX8536,
         WX8538, WX8539, WX8540, WX8541, WX8542, WX8543, WX8544, WX8545,
         WX8546, WX8547, WX8548, WX8549, WX8550, WX8551, WX8552, WX8553,
         WX8554, WX8555, WX8556, WX8557, WX8558, WX8559, WX8560, WX8561,
         WX8562, WX8563, WX8564, WX8565, WX8566, WX8567, WX8568, WX8569,
         WX8570, WX8572, WX8573, WX8574, WX8575, WX8576, WX8577, WX8578,
         WX8579, WX8580, WX8581, WX8582, WX8583, WX8584, WX8585, WX8586,
         WX8587, WX8588, WX8589, WX8590, WX8591, WX8592, WX8593, WX8594,
         WX8595, WX8596, WX8597, WX8598, WX8599, WX8600, WX8601, WX8602,
         WX8603, WX8604, WX8606, WX8607, WX8608, WX8609, WX8610, WX8611,
         WX8612, WX8613, WX8614, WX8615, WX8616, WX8617, WX8618, WX8619,
         WX8620, WX8621, WX8622, WX8623, WX8624, WX8625, WX8626, WX8627,
         WX8628, WX8629, WX8630, WX8631, WX8632, WX8633, WX8634, WX8635,
         WX8636, WX8637, WX8638, WX8640, WX8641, WX8642, WX8643, WX8644,
         WX8645, WX8646, WX8647, WX8648, WX8649, WX8650, WX8651, WX8652,
         WX8653, WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1, WX9024,
         DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, DFF_1315_n1, WX9030,
         DFF_1316_n1, WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038,
         DFF_1320_n1, WX9040, DFF_1321_n1, WX9042, DFF_1322_n1, WX9044,
         DFF_1323_n1, WX9046, DFF_1324_n1, WX9048, DFF_1325_n1, WX9050,
         DFF_1326_n1, WX9052, DFF_1327_n1, WX9054, DFF_1328_n1, WX9056,
         DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n8352, n8351, n8350,
         n8349, n8348, n8347, n8346, n8343, n8342, n8341, n8340, n8339, n8338,
         n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328,
         n8325, n8324, n8323, n8322, WX9597, n8321, WX9695, n8320, WX9697,
         n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705, n8315,
         WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311, WX9715,
         n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305, WX9725,
         n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733, WX9734,
         WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741, WX9742,
         WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749, WX9750,
         WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758, WX9759,
         WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766, WX9767,
         WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774, WX9775,
         WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782, WX9783,
         WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791, WX9792,
         WX9793, WX9794, WX9795, WX9796, WX9797, WX9798, WX9799, WX9800,
         WX9801, WX9802, WX9803, WX9804, WX9805, WX9806, WX9807, WX9808,
         WX9809, WX9810, WX9811, WX9812, WX9813, WX9814, WX9815, WX9816,
         WX9817, WX9818, WX9819, WX9821, WX9822, WX9823, WX9824, WX9825,
         WX9826, WX9827, WX9828, WX9829, WX9830, WX9831, WX9832, WX9833,
         WX9834, WX9835, WX9836, WX9837, WX9838, WX9839, WX9840, WX9841,
         WX9842, WX9843, WX9844, WX9845, WX9846, WX9847, WX9848, WX9849,
         WX9850, WX9851, WX9852, WX9853, WX9855, WX9856, WX9857, WX9858,
         WX9859, WX9860, WX9861, WX9862, WX9863, WX9864, WX9865, WX9866,
         WX9867, WX9868, WX9869, WX9870, WX9871, WX9872, WX9873, WX9874,
         WX9875, WX9876, WX9877, WX9878, WX9879, WX9880, WX9881, WX9882,
         WX9883, WX9884, WX9885, WX9886, WX9887, WX9889, WX9890, WX9891,
         WX9892, WX9893, WX9894, WX9895, WX9896, WX9897, WX9898, WX9899,
         WX9900, WX9901, WX9902, WX9903, WX9904, WX9905, WX9906, WX9907,
         WX9908, WX9909, WX9910, WX9911, WX9912, WX9913, WX9914, WX9915,
         WX9916, WX9917, WX9918, WX9919, WX9920, WX9921, WX9923, WX9924,
         WX9925, WX9926, WX9927, WX9928, WX9929, WX9930, WX9931, WX9932,
         WX9933, WX9934, WX9935, WX9936, WX9937, WX9938, WX9939, WX9940,
         WX9941, WX9942, WX9943, WX9944, WX9945, WX9946, WX9947, WX9948,
         WX9949, WX9950, WX10315, DFF_1504_n1, WX10317, DFF_1505_n1, WX10319,
         WX10321, DFF_1507_n1, WX10323, DFF_1508_n1, WX10325, DFF_1509_n1,
         WX10327, DFF_1510_n1, WX10329, DFF_1511_n1, WX10331, DFF_1512_n1,
         WX10333, DFF_1513_n1, WX10335, DFF_1514_n1, WX10337, DFF_1515_n1,
         WX10339, DFF_1516_n1, WX10341, DFF_1517_n1, WX10343, DFF_1518_n1,
         WX10345, DFF_1519_n1, WX10347, DFF_1520_n1, WX10349, DFF_1521_n1,
         WX10351, DFF_1522_n1, WX10353, WX10355, DFF_1524_n1, WX10357,
         DFF_1525_n1, WX10359, DFF_1526_n1, WX10361, DFF_1527_n1, WX10363,
         DFF_1528_n1, WX10365, DFF_1529_n1, WX10367, DFF_1530_n1, WX10369,
         DFF_1531_n1, WX10371, DFF_1532_n1, WX10373, DFF_1533_n1, WX10375,
         DFF_1534_n1, WX10377, DFF_1535_n1, WX10829, n8295, n8294, n8293,
         n8290, n8289, n8288, n8287, n8286, n8285, n8284, n8283, n8282, n8281,
         n8280, n8279, n8278, n8277, n8276, n8275, n8272, n8271, n8270, n8269,
         n8268, n8267, n8266, n8265, n8264, WX10890, n8263, n8262, n8261,
         n8260, n8259, n8258, n8257, n8254, n8253, n8252, n8251, n8250, n8249,
         n8248, n8247, n8246, WX11021, WX11023, WX11025, WX11027, WX11029,
         WX11031, WX11033, WX11037, WX11039, WX11041, WX11043, WX11045,
         WX11047, WX11049, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, WX11086, WX11087, WX11088, WX11089, WX11090, WX11091,
         WX11092, WX11093, WX11094, WX11095, WX11096, WX11097, WX11098,
         WX11099, WX11100, WX11101, WX11102, WX11104, WX11105, WX11106,
         WX11107, WX11108, WX11109, WX11110, WX11111, WX11112, WX11113,
         WX11114, WX11115, WX11116, WX11117, WX11118, WX11119, WX11120,
         WX11121, WX11122, WX11123, WX11124, WX11125, WX11126, WX11127,
         WX11128, WX11129, WX11130, WX11131, WX11132, WX11133, WX11134,
         WX11135, WX11136, WX11138, WX11139, WX11140, WX11141, WX11142,
         WX11143, WX11144, WX11145, WX11146, WX11147, WX11148, WX11149,
         WX11150, WX11151, WX11152, WX11153, WX11154, WX11155, WX11156,
         WX11157, WX11158, WX11159, WX11160, WX11161, WX11162, WX11163,
         WX11164, WX11165, WX11166, WX11167, WX11168, WX11169, WX11170,
         WX11172, WX11173, WX11174, WX11175, WX11176, WX11177, WX11178,
         WX11179, WX11180, WX11181, WX11182, WX11183, WX11184, WX11185,
         WX11186, WX11187, WX11188, WX11189, WX11190, WX11191, WX11192,
         WX11193, WX11194, WX11195, WX11196, WX11197, WX11198, WX11199,
         WX11200, WX11201, WX11202, WX11203, WX11204, WX11206, WX11207,
         WX11208, WX11209, WX11210, WX11211, WX11212, WX11213, WX11214,
         WX11215, WX11216, WX11217, WX11218, WX11219, WX11220, WX11221,
         WX11222, WX11223, WX11224, WX11225, WX11226, WX11227, WX11228,
         WX11229, WX11230, WX11231, WX11232, WX11233, WX11234, WX11235,
         WX11236, WX11237, WX11238, WX11240, WX11241, WX11242, WX11243,
         WX11608, DFF_1696_n1, WX11610, WX11612, DFF_1698_n1, WX11614,
         DFF_1699_n1, WX11616, DFF_1700_n1, WX11618, DFF_1701_n1, WX11620,
         DFF_1702_n1, WX11622, DFF_1703_n1, WX11624, DFF_1704_n1, WX11626,
         DFF_1705_n1, WX11628, DFF_1706_n1, WX11630, DFF_1707_n1, WX11632,
         DFF_1708_n1, WX11634, DFF_1709_n1, WX11636, WX11638, DFF_1711_n1,
         WX11640, DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, WX11646,
         DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1, WX11652,
         DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1, WX11658,
         DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1, WX11664,
         DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1, WX11670,
         n2245, n2153, n3278, n2152, Tj_Trigger, Tj_OUT1, Tj_OUT2, Tj_OUT3,
         Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n432, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n583, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4146, n4148, n4150, n4152, n4155, n4158, n4161,
         n4163, n4165, n4167, n4169, n4171, n4173, n4175, n4178, n4181, n4183,
         n4185, n4187, n4189, n4191, n4193, n4195, n4197, n4199, n4201, n4203,
         n4205, n4207, n4209, n4211, n4213, n4215, n4217, n4219, n4221, n4223,
         n4225, n4228, n4231, n4234, n4236, n4238, n4240, n4242, n4244, n4247,
         n4250, n4253, n4255, n4257, n4259, n4261, n4263, n4266, n4269, n4272,
         n4274, n4276, n4278, n4280, n4282, n4284, n4286, n4288, n4290, n4293,
         n4295, n4297, n4299, n4301, n4303, n4305, n4307, n4309, n4311, n4313,
         n4315, n4318, n4321, n4323, n4325, n4327, n4329, n4331, n4333, n4335,
         n4338, n4340, n4342, n4345, n4347, n4349, n4352, n4354, n4356, n4359,
         n4361, n4363, n4365, n4367, n4369, n4371, n4373, n4375, n4378, n4379,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8255, n8256, n8273, n8274, n8291, n8292, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8308, n8309, n8326, n8327, n8344, n8345,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8379,
         n8380, n8397, n8398, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8432, n8433, n8450, n8451, n8468, n8469, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8485, n8486, n8503, n8504,
         n8521, n8522, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8538, n8539, n8556, n8557, n8574, n8575, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8614, n8615, n8633, n8634,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8659, n8660,
         n8678, n8679, n8697, n8698, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1, U5719_n1,
         U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1, U5726_n1,
         U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1, U5733_n1,
         U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1, U5740_n1,
         U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1, U5747_n1,
         U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1,
         U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1,
         U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1, U5768_n1,
         U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1, U5775_n1,
         U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1, U5782_n1,
         U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1, U5789_n1,
         U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1, U5796_n1,
         U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1, U5803_n1,
         U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1, U5810_n1,
         U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1, U5817_n1,
         U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1, U5824_n1,
         U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1, U5831_n1,
         U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1, U5838_n1,
         U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1, U5845_n1,
         U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1, U5852_n1,
         U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1, U5859_n1,
         U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1, U5866_n1,
         U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1, U5873_n1,
         U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1, U5880_n1,
         U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1, U5887_n1,
         U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1, U5894_n1,
         U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1, U5901_n1,
         U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1, U5908_n1,
         U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1, U5915_n1,
         U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1, U5922_n1,
         U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1, U5929_n1,
         U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1, U5936_n1,
         U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U5943_n1,
         U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1, U5950_n1,
         U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1, U5957_n1,
         U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1, U5964_n1,
         U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1, U5971_n1,
         U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1, U5978_n1,
         U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1, U5985_n1,
         U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1, U5992_n1,
         U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1, U5999_n1,
         U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1, U6006_n1,
         U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1, U6013_n1,
         U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1, U6020_n1,
         U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1, U6027_n1,
         U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1, U6034_n1,
         U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1, U6041_n1,
         U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1, U6048_n1,
         U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1, U6055_n1,
         U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1, U6062_n1,
         U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1, U6069_n1,
         U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1, U6076_n1,
         U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1, U6083_n1,
         U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1, U6090_n1,
         U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1, U6097_n1,
         U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1, U6104_n1,
         U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1, U6111_n1,
         U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1, U6118_n1,
         U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1, U6125_n1,
         U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1, U6132_n1,
         U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1, U6139_n1,
         U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1, U6146_n1,
         U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1, U6153_n1,
         U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1, U6160_n1,
         U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1, U6167_n1,
         U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1, U6174_n1,
         U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1, U6181_n1,
         U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1, U6188_n1,
         U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1, U6195_n1,
         U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1, U6202_n1,
         U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1, U6209_n1,
         U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1, U6216_n1,
         U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1, U6223_n1,
         U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1, U6230_n1,
         U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1, U6237_n1,
         U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1, U6244_n1,
         U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1, U6251_n1,
         U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1, U6258_n1,
         U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1, U6265_n1,
         U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1, U6272_n1,
         U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1, U6279_n1,
         U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1, U6286_n1,
         U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1, U6293_n1,
         U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1, U6300_n1,
         U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1, U6307_n1,
         U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1, U6314_n1,
         U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1, U6321_n1,
         U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1, U6328_n1,
         U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1, U6335_n1,
         U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1, U6342_n1,
         U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1, U6349_n1,
         U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1, U6356_n1,
         U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1, U6363_n1,
         U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1, U6370_n1,
         U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1, U6377_n1,
         U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1, U6384_n1,
         U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1, U6391_n1,
         U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1, U6398_n1,
         U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1, U6405_n1,
         U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1, U6412_n1,
         U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1, U6419_n1,
         U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1, U6426_n1,
         U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1, U6433_n1,
         U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1, U6440_n1,
         U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1, U6447_n1,
         U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1, U6454_n1,
         U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1, U6461_n1,
         U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1, U6468_n1,
         U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1, U6475_n1,
         U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n5101), .CLK(n5442), .Q(
        WX485), .QN(n4379) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n5096), .CLK(n5444), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n5096), .CLK(n5444), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n5097), .CLK(n5444), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n5097), .CLK(n5444), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n5097), .CLK(n5444), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n5097), .CLK(n5444), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n5097), .CLK(n5444), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n5097), .CLK(n5444), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n5098), .CLK(n5443), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n5098), .CLK(n5443), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n5098), .CLK(n5443), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n5098), .CLK(n5443), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n5098), .CLK(n5443), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n5098), .CLK(n5443), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n5099), .CLK(n5443), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n5099), .CLK(n5443), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n5099), .CLK(n5443), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n5099), .CLK(n5443), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n5099), .CLK(n5443), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n5099), .CLK(n5443), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n5100), .CLK(n5442), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n5100), .CLK(n5442), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n5100), .CLK(n5442), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n5100), .CLK(n5442), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n5100), .CLK(n5442), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n5100), .CLK(n5442), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n5101), .CLK(n5442), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n5101), .CLK(n5442), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n5101), .CLK(n5442), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n5101), .CLK(n5442), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n5101), .CLK(n5442), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n5096), .CLK(n5444), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(n2), .SI(WX645), .SE(n5096), .CLK(n5444), .Q(WX647), 
        .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(n3), .SI(WX647), .SE(n5096), .CLK(n5444), .Q(WX649), 
        .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(n4), .SI(WX649), .SE(n5096), .CLK(n5444), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(n5), .SI(test_si3), .SE(n5095), .CLK(n5445), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(n6), .SI(WX653), .SE(n5095), .CLK(n5445), .Q(WX655), 
        .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(n7), .SI(WX655), .SE(n5095), .CLK(n5445), .Q(WX657), 
        .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n5094), .CLK(n5445), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(n8), .SI(WX659), .SE(n5094), .CLK(n5445), .Q(WX661), 
        .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(n9), .SI(WX661), .SE(n5094), .CLK(n5445), .Q(WX663), 
        .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(n10), .SI(WX663), .SE(n5093), .CLK(n5446), .Q(WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n5093), .CLK(n5446), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(n11), .SI(WX667), .SE(n5093), .CLK(n5446), .Q(WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(n12), .SI(WX669), .SE(n5092), .CLK(n5446), .Q(WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(n13), .SI(WX671), .SE(n5092), .CLK(n5446), .Q(WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n5091), .CLK(n5447), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(n14), .SI(WX675), .SE(n5091), .CLK(n5447), .Q(WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(n15), .SI(WX677), .SE(n5090), .CLK(n5447), .Q(WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(n16), .SI(WX679), .SE(n5089), .CLK(n5448), .Q(WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(n17), .SI(WX681), .SE(n5089), .CLK(n5448), .Q(WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(n18), .SI(WX683), .SE(n5088), .CLK(n5448), .Q(WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n5087), .CLK(n5449), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(n19), .SI(test_si4), .SE(n4815), .CLK(n5585), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(n20), .SI(WX689), .SE(n5086), .CLK(n5449), .Q(WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(n21), .SI(WX691), .SE(n5085), .CLK(n5450), .Q(WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(n22), .SI(WX693), .SE(n5085), .CLK(n5450), .Q(WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(n23), .SI(WX695), .SE(n5084), .CLK(n5450), .Q(WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(n24), .SI(WX697), .SE(n5083), .CLK(n5451), .Q(WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(n25), .SI(WX699), .SE(n5083), .CLK(n5451), .Q(WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(n26), .SI(WX701), .SE(n5082), .CLK(n5451), .Q(WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(n27), .SI(WX703), .SE(n5081), .CLK(n5452), .Q(WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(n28), .SI(WX705), .SE(n5081), .CLK(n5452), .Q(WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n5080), .CLK(n5452), .Q(
        WX709) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n5080), .CLK(n5452), .Q(
        WX711), .QN(n4629) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n5079), .CLK(n5453), .Q(
        WX713), .QN(n9736) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n5095), .CLK(n5445), .Q(
        WX715), .QN(n4638) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n5095), .CLK(n5445), .Q(
        WX717), .QN(n9737) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n5095), .CLK(n5445), .Q(
        WX719), .QN(n9738) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n5094), .CLK(n5445), .Q(
        WX721), .QN(n9739) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n5094), .CLK(n5445), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n5094), .CLK(n5445), .Q(
        WX725), .QN(n9740) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n5093), .CLK(n5446), .Q(
        WX727), .QN(n4655) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n5093), .CLK(n5446), .Q(
        WX729), .QN(n4659) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n5093), .CLK(n5446), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n5092), .CLK(n5446), .Q(
        WX733), .QN(n9741) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n5092), .CLK(n5446), .Q(
        WX735), .QN(n9742) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n5091), .CLK(n5447), .Q(
        WX737), .QN(n9743) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n5091), .CLK(n5447), .Q(
        WX739) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n5090), .CLK(n5447), .Q(
        WX741), .QN(n4657) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n5090), .CLK(n5447), .Q(
        WX743), .QN(n9744) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n5089), .CLK(n5448), .Q(
        WX745), .QN(n9745) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n5088), .CLK(n5448), .Q(
        WX747), .QN(n9746) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n5088), .CLK(n5448), .Q(
        WX749), .QN(n9747) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n5087), .CLK(n5449), .Q(
        WX751), .QN(n4643) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n5087), .CLK(n5449), .Q(
        WX753) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n5086), .CLK(n5449), .Q(
        WX755), .QN(n9731) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n5085), .CLK(n5450), .Q(
        WX757), .QN(n4667) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n5085), .CLK(n5450), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n5084), .CLK(n5450), .Q(
        WX761), .QN(n9732) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n5083), .CLK(n5451), .Q(
        WX763), .QN(n9733) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n5083), .CLK(n5451), .Q(
        WX765), .QN(n9735) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n5082), .CLK(n5451), .Q(
        WX767) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n5081), .CLK(n5452), .Q(
        WX769), .QN(n9748) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n5081), .CLK(n5452), .Q(
        WX771), .QN(n4670) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n5080), .CLK(n5452), .Q(
        WX773), .QN(n9734) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n5079), .CLK(n5453), .Q(
        WX775) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n5079), .CLK(n5453), .Q(
        WX777) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n5079), .CLK(n5453), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n5078), .CLK(n5453), .Q(
        WX781) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n5078), .CLK(n5453), .Q(
        WX783) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n5078), .CLK(n5453), .Q(
        WX785) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n5077), .CLK(n5454), .Q(
        WX787) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n5077), .CLK(n5454), .Q(
        WX789) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n5077), .CLK(n5454), .Q(
        WX791) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n5076), .CLK(n5454), .Q(
        WX793) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n5076), .CLK(n5454), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n5092), .CLK(n5446), 
        .Q(WX797) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n5092), .CLK(n5446), .Q(
        WX799) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n5091), .CLK(n5447), .Q(
        WX801) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n5091), .CLK(n5447), .Q(
        WX803), .QN(n4651) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n5090), .CLK(n5447), .Q(
        WX805) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n5090), .CLK(n5447), .Q(
        WX807) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n5089), .CLK(n5448), .Q(
        WX809) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n5088), .CLK(n5448), .Q(
        WX811) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n5088), .CLK(n5448), .Q(
        WX813) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n5087), .CLK(n5449), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n5086), .CLK(n5449), .Q(
        WX817), .QN(n9730) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n5086), .CLK(n5449), .Q(
        WX819) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n5085), .CLK(n5450), .Q(
        WX821) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n5084), .CLK(n5450), .Q(
        WX823) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n5084), .CLK(n5450), .Q(
        WX825) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n5083), .CLK(n5451), .Q(
        WX827) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n5082), .CLK(n5451), .Q(
        WX829) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n5082), .CLK(n5451), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n5081), .CLK(n5452), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n5080), .CLK(n5452), .Q(
        WX835) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n5080), .CLK(n5452), .Q(
        WX837), .QN(n4664) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n5079), .CLK(n5453), .Q(
        WX839), .QN(n4630) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n5079), .CLK(n5453), .Q(
        WX841), .QN(n4633) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n5078), .CLK(n5453), .Q(
        WX843), .QN(n4637) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n5078), .CLK(n5453), .Q(
        WX845), .QN(n4640) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n5078), .CLK(n5453), .Q(
        WX847), .QN(n4641) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n5077), .CLK(n5454), .Q(
        WX849), .QN(n4645) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n5077), .CLK(n5454), .Q(
        WX851), .QN(n4648) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n5077), .CLK(n5454), .Q(
        WX853), .QN(n4650) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n5076), .CLK(n5454), .Q(
        WX855), .QN(n4656) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n5076), .CLK(n5454), .Q(
        WX857), .QN(n4660) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n5076), .CLK(n5454), .Q(
        WX859), .QN(n4662) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n5076), .CLK(n5454), .Q(
        WX861), .QN(n4632) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n5075), .CLK(n5455), .Q(
        WX863), .QN(n4639) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n5075), .CLK(n5455), .Q(
        WX865), .QN(n4644) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n5075), .CLK(n5455), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n5090), .CLK(n5447), 
        .Q(WX869), .QN(n4658) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n5089), .CLK(n5448), .Q(
        WX871), .QN(n4665) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n5089), .CLK(n5448), .Q(
        WX873), .QN(n4634) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n5088), .CLK(n5448), .Q(
        WX875), .QN(n4646) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n5087), .CLK(n5449), .Q(
        WX877), .QN(n4669) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n5087), .CLK(n5449), .Q(
        WX879), .QN(n4642) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n5086), .CLK(n5449), .Q(
        WX881), .QN(n4647) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n5086), .CLK(n5449), .Q(
        WX883), .QN(n4652) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n5085), .CLK(n5450), .Q(
        WX885), .QN(n4668) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n5084), .CLK(n5450), .Q(
        WX887), .QN(n4661) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n5084), .CLK(n5450), .Q(
        WX889), .QN(n4653) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n5083), .CLK(n5451), .Q(
        WX891), .QN(n4654) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n5082), .CLK(n5451), .Q(
        WX893), .QN(n4631) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n5082), .CLK(n5451), .Q(
        WX895), .QN(n4666) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n5081), .CLK(n5452), .Q(
        WX897), .QN(n4635) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n5080), .CLK(n5452), .Q(
        WX899), .QN(n4671) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n4817), .CLK(n5584), .Q(
        CRC_OUT_9_0), .QN(DFF_160_n1) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n4817), .CLK(n5584), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n4817), .CLK(n5584), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_3) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n4816), .CLK(n5584), 
        .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n4815), .CLK(n5585), 
        .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n4815), .CLK(n5585), 
        .Q(CRC_OUT_9_10) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n4815), .CLK(n5585), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n4815), .CLK(n5585), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n4815), .CLK(n5585), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n4814), .CLK(n5585), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n4814), .CLK(n5585), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n4814), .CLK(n5585), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n4814), .CLK(n5585), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n4814), .CLK(n5585), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n4814), .CLK(n5585), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n5075), .CLK(n5455), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n5075), .CLK(n5455), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n5075), .CLK(n5455), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n5074), .CLK(n5455), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n5073), .CLK(n5456), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n5073), .CLK(n5456), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n5073), .CLK(n5456), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n55), .SI(CRC_OUT_9_31), .SE(n5073), .CLK(n5456), 
        .Q(WX1778), .QN(n4387) );
  SDFFX1 DFF_193_Q_reg ( .D(n56), .SI(WX1778), .SE(n5068), .CLK(n5458), .Q(
        n8702) );
  SDFFX1 DFF_194_Q_reg ( .D(n57), .SI(n8702), .SE(n5068), .CLK(n5458), .Q(
        n8701) );
  SDFFX1 DFF_195_Q_reg ( .D(n58), .SI(n8701), .SE(n5068), .CLK(n5458), .Q(
        n8700) );
  SDFFX1 DFF_196_Q_reg ( .D(n59), .SI(n8700), .SE(n5068), .CLK(n5458), .Q(
        n8699) );
  SDFFX1 DFF_197_Q_reg ( .D(n60), .SI(n8699), .SE(n5068), .CLK(n5458), .Q(
        test_so11) );
  SDFFX1 DFF_198_Q_reg ( .D(n61), .SI(test_si12), .SE(n5069), .CLK(n5458), .Q(
        n8696) );
  SDFFX1 DFF_199_Q_reg ( .D(n62), .SI(n8696), .SE(n5069), .CLK(n5458), .Q(
        n8695) );
  SDFFX1 DFF_200_Q_reg ( .D(n63), .SI(n8695), .SE(n5069), .CLK(n5458), .Q(
        n8694) );
  SDFFX1 DFF_201_Q_reg ( .D(n64), .SI(n8694), .SE(n5069), .CLK(n5458), .Q(
        n8693) );
  SDFFX1 DFF_202_Q_reg ( .D(n65), .SI(n8693), .SE(n5069), .CLK(n5458), .Q(
        n8692) );
  SDFFX1 DFF_203_Q_reg ( .D(n66), .SI(n8692), .SE(n5069), .CLK(n5458), .Q(
        n8691) );
  SDFFX1 DFF_204_Q_reg ( .D(n67), .SI(n8691), .SE(n5070), .CLK(n5457), .Q(
        n8690) );
  SDFFX1 DFF_205_Q_reg ( .D(n68), .SI(n8690), .SE(n5070), .CLK(n5457), .Q(
        n8689) );
  SDFFX1 DFF_206_Q_reg ( .D(n69), .SI(n8689), .SE(n5070), .CLK(n5457), .Q(
        n8688) );
  SDFFX1 DFF_207_Q_reg ( .D(n70), .SI(n8688), .SE(n5070), .CLK(n5457), .Q(
        n8687) );
  SDFFX1 DFF_208_Q_reg ( .D(n71), .SI(n8687), .SE(n5070), .CLK(n5457), .Q(
        n8686) );
  SDFFX1 DFF_209_Q_reg ( .D(n72), .SI(n8686), .SE(n5070), .CLK(n5457), .Q(
        n8685) );
  SDFFX1 DFF_210_Q_reg ( .D(n73), .SI(n8685), .SE(n5071), .CLK(n5457), .Q(
        n8684) );
  SDFFX1 DFF_211_Q_reg ( .D(n74), .SI(n8684), .SE(n5071), .CLK(n5457), .Q(
        n8683) );
  SDFFX1 DFF_212_Q_reg ( .D(n75), .SI(n8683), .SE(n5071), .CLK(n5457), .Q(
        n8682) );
  SDFFX1 DFF_213_Q_reg ( .D(n76), .SI(n8682), .SE(n5071), .CLK(n5457), .Q(
        n8681) );
  SDFFX1 DFF_214_Q_reg ( .D(n77), .SI(n8681), .SE(n5071), .CLK(n5457), .Q(
        n8680) );
  SDFFX1 DFF_215_Q_reg ( .D(n78), .SI(n8680), .SE(n5071), .CLK(n5457), .Q(
        test_so12) );
  SDFFX1 DFF_216_Q_reg ( .D(n79), .SI(test_si13), .SE(n5072), .CLK(n5456), .Q(
        n8677) );
  SDFFX1 DFF_217_Q_reg ( .D(n80), .SI(n8677), .SE(n5072), .CLK(n5456), .Q(
        n8676) );
  SDFFX1 DFF_218_Q_reg ( .D(n81), .SI(n8676), .SE(n5072), .CLK(n5456), .Q(
        n8675) );
  SDFFX1 DFF_219_Q_reg ( .D(n82), .SI(n8675), .SE(n5072), .CLK(n5456), .Q(
        n8674) );
  SDFFX1 DFF_220_Q_reg ( .D(n83), .SI(n8674), .SE(n5072), .CLK(n5456), .Q(
        n8673) );
  SDFFX1 DFF_221_Q_reg ( .D(n84), .SI(n8673), .SE(n5072), .CLK(n5456), .Q(
        n8672) );
  SDFFX1 DFF_222_Q_reg ( .D(n85), .SI(n8672), .SE(n5073), .CLK(n5456), .Q(
        n8671) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n5073), .CLK(n5456), .Q(
        n8670) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n5068), .CLK(n5458), .Q(
        n8669), .QN(n9694) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n5067), .CLK(n5459), .Q(
        n8668), .QN(n9689) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n5067), .CLK(n5459), .Q(
        n8667), .QN(n9687) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n4824), .CLK(n5580), .Q(
        n8666), .QN(n9685) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n5065), .CLK(n5460), .Q(
        n8665), .QN(n9683) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n5065), .CLK(n5460), .Q(
        n8664), .QN(n9679) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n5064), .CLK(n5460), .Q(
        n8663), .QN(n9677) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n5064), .CLK(n5460), .Q(
        n8662), .QN(n9675) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n5063), .CLK(n5461), .Q(
        n8661), .QN(n9673) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n5062), .CLK(n5461), .Q(
        test_so13), .QN(n4711) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n5061), .CLK(n5462), 
        .Q(n8658), .QN(n9670) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n5061), .CLK(n5462), .Q(
        n8657), .QN(n9668) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n5060), .CLK(n5462), .Q(
        n8656), .QN(n9666) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n5060), .CLK(n5462), .Q(
        n8655), .QN(n9662) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n4824), .CLK(n5580), .Q(
        n8654), .QN(n9660) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n4824), .CLK(n5580), .Q(
        n8653), .QN(n9659) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n5058), .CLK(n5463), .Q(
        WX1970) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n5058), .CLK(n5463), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n5058), .CLK(n5463), .Q(
        WX1974) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n5058), .CLK(n5463), .Q(
        WX1976) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n5057), .CLK(n5464), .Q(
        WX1978) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n5057), .CLK(n5464), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n5057), .CLK(n5464), .Q(
        WX1982) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n5057), .CLK(n5464), .Q(
        WX1984) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n5057), .CLK(n5464), .Q(
        WX1986) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n5057), .CLK(n5464), .Q(
        WX1988) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n5056), .CLK(n5464), .Q(
        WX1990) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n5056), .CLK(n5464), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n5056), .CLK(n5464), 
        .Q(WX1994) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n5056), .CLK(n5464), .Q(
        WX1996) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n5055), .CLK(n5465), .Q(
        WX1998) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n5055), .CLK(n5465), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n5067), .CLK(n5459), .Q(
        WX2002), .QN(n4038) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n5067), .CLK(n5459), .Q(
        WX2004), .QN(n4144) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n5066), .CLK(n5459), .Q(
        WX2006), .QN(n4143) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n5066), .CLK(n5459), .Q(
        WX2008) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n5066), .CLK(n5459), .Q(
        WX2010), .QN(n4141) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n5065), .CLK(n5460), .Q(
        WX2012), .QN(n4140) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n5064), .CLK(n5460), .Q(
        WX2014), .QN(n4139) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n5064), .CLK(n5460), .Q(
        WX2016), .QN(n4138) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n5063), .CLK(n5461), .Q(
        WX2018), .QN(n4137) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n5062), .CLK(n5461), .Q(
        WX2020) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n5062), .CLK(n5461), .Q(
        WX2022), .QN(n4135) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n5061), .CLK(n5462), .Q(
        WX2024), .QN(n4134) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n5060), .CLK(n5462), .Q(
        WX2026), .QN(n4133) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n5060), .CLK(n5462), .Q(
        test_so15), .QN(n9663) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n4824), .CLK(n5580), 
        .Q(WX2030), .QN(n4132) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n4824), .CLK(n5580), .Q(
        WX2032), .QN(n4131) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n4824), .CLK(n5580), .Q(
        WX2034), .QN(n9657) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n4823), .CLK(n5581), .Q(
        WX2036), .QN(n9655) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n4823), .CLK(n5581), .Q(
        WX2038), .QN(n9653) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n4822), .CLK(n5581), .Q(
        WX2040), .QN(n9651) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n4822), .CLK(n5581), .Q(
        WX2042), .QN(n9649) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n4821), .CLK(n5582), .Q(
        WX2044), .QN(n9647) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n4821), .CLK(n5582), .Q(
        WX2046), .QN(n9645) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n4820), .CLK(n5582), .Q(
        WX2048), .QN(n9643) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n4820), .CLK(n5582), .Q(
        WX2050), .QN(n9641) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n4819), .CLK(n5583), .Q(
        WX2052), .QN(n9639) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n4819), .CLK(n5583), .Q(
        WX2054), .QN(n9637) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n5056), .CLK(n5464), .Q(
        WX2056), .QN(n9635) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n5056), .CLK(n5464), .Q(
        WX2058), .QN(n9633) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n5055), .CLK(n5465), .Q(
        WX2060), .QN(n9631) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n5055), .CLK(n5465), .Q(
        WX2062), .QN(n9629) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n5055), .CLK(n5465), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n5067), .CLK(n5459), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n5067), .CLK(n5459), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n5066), .CLK(n5459), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n5066), .CLK(n5459), .Q(
        WX2072), .QN(n4142) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n5066), .CLK(n5459), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n5065), .CLK(n5460), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n5064), .CLK(n5460), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n5063), .CLK(n5461), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n5063), .CLK(n5461), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n5062), .CLK(n5461), .Q(
        WX2084), .QN(n4136) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n5062), .CLK(n5461), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n5061), .CLK(n5462), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n5060), .CLK(n5462), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n5059), .CLK(n5463), .Q(
        WX2092), .QN(n9664) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n5059), .CLK(n5463), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n5059), .CLK(n5463), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n5058), .CLK(n5463), .Q(
        WX2098), .QN(n4378) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n4823), .CLK(n5581), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n4823), .CLK(n5581), 
        .Q(WX2102), .QN(n4375) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n4822), .CLK(n5581), .Q(
        WX2104), .QN(n4373) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n4822), .CLK(n5581), .Q(
        WX2106), .QN(n4371) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n4821), .CLK(n5582), .Q(
        WX2108), .QN(n4369) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n4821), .CLK(n5582), .Q(
        WX2110), .QN(n4367) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n4820), .CLK(n5582), .Q(
        WX2112), .QN(n4365) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n4820), .CLK(n5582), .Q(
        WX2114), .QN(n4363) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n4819), .CLK(n5583), .Q(
        WX2116), .QN(n4361) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n4819), .CLK(n5583), .Q(
        WX2118), .QN(n4359) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n4818), .CLK(n5583), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n4818), .CLK(n5583), .Q(
        WX2122), .QN(n4356) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n4818), .CLK(n5583), .Q(
        WX2124), .QN(n4354) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n4817), .CLK(n5584), .Q(
        WX2126), .QN(n4352) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n5055), .CLK(n5465), .Q(
        WX2128), .QN(n9627) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n5054), .CLK(n5465), .Q(
        WX2130), .QN(n4603) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n5054), .CLK(n5465), .Q(
        WX2132), .QN(n4604) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n5054), .CLK(n5465), .Q(
        WX2134), .QN(n4605) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n5054), .CLK(n5465), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n5065), .CLK(n5460), 
        .Q(WX2138), .QN(n4606) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n5065), .CLK(n5460), .Q(
        WX2140), .QN(n4607) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n5064), .CLK(n5460), .Q(
        WX2142), .QN(n4608) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n5063), .CLK(n5461), .Q(
        WX2144), .QN(n4609) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n5063), .CLK(n5461), .Q(
        WX2146), .QN(n4610) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n5062), .CLK(n5461), .Q(
        WX2148), .QN(n4611) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n5061), .CLK(n5462), .Q(
        WX2150), .QN(n4612) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n5061), .CLK(n5462), .Q(
        WX2152), .QN(n4613) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n5060), .CLK(n5462), .Q(
        WX2154), .QN(n4614) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n5059), .CLK(n5463), .Q(
        WX2156), .QN(n4615) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n5059), .CLK(n5463), .Q(
        WX2158), .QN(n4616) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n5059), .CLK(n5463), .Q(
        WX2160), .QN(n4406) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n5058), .CLK(n5463), .Q(
        WX2162), .QN(n4617) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n4823), .CLK(n5581), .Q(
        WX2164), .QN(n4618) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n4823), .CLK(n5581), .Q(
        WX2166), .QN(n4619) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n4822), .CLK(n5581), .Q(
        WX2168), .QN(n4620) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n4822), .CLK(n5581), .Q(
        WX2170), .QN(n4407) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n4821), .CLK(n5582), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n4821), .CLK(n5582), 
        .Q(WX2174), .QN(n4621) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n4820), .CLK(n5582), .Q(
        WX2176), .QN(n4622) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n4820), .CLK(n5582), .Q(
        WX2178), .QN(n4623) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n4819), .CLK(n5583), .Q(
        WX2180), .QN(n4624) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n4819), .CLK(n5583), .Q(
        WX2182), .QN(n4625) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n4818), .CLK(n5583), .Q(
        WX2184), .QN(n4408) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n4818), .CLK(n5583), .Q(
        WX2186), .QN(n4626) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n4818), .CLK(n5583), .Q(
        WX2188), .QN(n4627) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n4817), .CLK(n5584), .Q(
        WX2190), .QN(n4628) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n4817), .CLK(n5584), .Q(
        WX2192), .QN(n4416) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n4830), .CLK(n5577), .Q(
        CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n4829), .CLK(n5578), 
        .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n4828), .CLK(n5578), 
        .Q(test_so20), .QN(n4703) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n4828), .CLK(n5578), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n4828), .CLK(n5578), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n4828), .CLK(n5578), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n4828), .CLK(n5578), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n4828), .CLK(n5578), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n4827), .CLK(n5579), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n4826), .CLK(n5579), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n4825), .CLK(n5580), .Q(test_so21), .QN(n4704) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n4825), .CLK(n5580), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n4825), .CLK(n5580), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n4825), .CLK(n5580), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n4825), .CLK(n5580), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n4825), .CLK(n5580), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n5054), .CLK(n5465), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n132), .SI(CRC_OUT_8_31), .SE(n5054), .CLK(n5465), 
        .Q(WX3071), .QN(n4386) );
  SDFFX1 DFF_385_Q_reg ( .D(n133), .SI(WX3071), .SE(n5048), .CLK(n5468), .Q(
        n8644) );
  SDFFX1 DFF_386_Q_reg ( .D(n134), .SI(n8644), .SE(n5049), .CLK(n5468), .Q(
        n8643) );
  SDFFX1 DFF_387_Q_reg ( .D(n135), .SI(n8643), .SE(n5049), .CLK(n5468), .Q(
        n8642) );
  SDFFX1 DFF_388_Q_reg ( .D(n136), .SI(n8642), .SE(n5049), .CLK(n5468), .Q(
        n8641) );
  SDFFX1 DFF_389_Q_reg ( .D(n137), .SI(n8641), .SE(n5049), .CLK(n5468), .Q(
        n8640) );
  SDFFX1 DFF_390_Q_reg ( .D(n138), .SI(n8640), .SE(n5049), .CLK(n5468), .Q(
        n8639) );
  SDFFX1 DFF_391_Q_reg ( .D(n139), .SI(n8639), .SE(n5049), .CLK(n5468), .Q(
        n8638) );
  SDFFX1 DFF_392_Q_reg ( .D(n140), .SI(n8638), .SE(n5050), .CLK(n5467), .Q(
        n8637) );
  SDFFX1 DFF_393_Q_reg ( .D(n141), .SI(n8637), .SE(n5050), .CLK(n5467), .Q(
        n8636) );
  SDFFX1 DFF_394_Q_reg ( .D(n142), .SI(n8636), .SE(n5050), .CLK(n5467), .Q(
        n8635) );
  SDFFX1 DFF_395_Q_reg ( .D(n143), .SI(n8635), .SE(n5050), .CLK(n5467), .Q(
        test_so22) );
  SDFFX1 DFF_396_Q_reg ( .D(n144), .SI(test_si23), .SE(n5050), .CLK(n5467), 
        .Q(n8632) );
  SDFFX1 DFF_397_Q_reg ( .D(n145), .SI(n8632), .SE(n5050), .CLK(n5467), .Q(
        n8631) );
  SDFFX1 DFF_398_Q_reg ( .D(n146), .SI(n8631), .SE(n5051), .CLK(n5467), .Q(
        n8630) );
  SDFFX1 DFF_399_Q_reg ( .D(n147), .SI(n8630), .SE(n5051), .CLK(n5467), .Q(
        n8629) );
  SDFFX1 DFF_400_Q_reg ( .D(n151), .SI(n8629), .SE(n5051), .CLK(n5467), .Q(
        n8628) );
  SDFFX1 DFF_401_Q_reg ( .D(n152), .SI(n8628), .SE(n5051), .CLK(n5467), .Q(
        n8627) );
  SDFFX1 DFF_402_Q_reg ( .D(n153), .SI(n8627), .SE(n5051), .CLK(n5467), .Q(
        n8626) );
  SDFFX1 DFF_403_Q_reg ( .D(n154), .SI(n8626), .SE(n5051), .CLK(n5467), .Q(
        n8625) );
  SDFFX1 DFF_404_Q_reg ( .D(n155), .SI(n8625), .SE(n5052), .CLK(n5466), .Q(
        n8624) );
  SDFFX1 DFF_405_Q_reg ( .D(n156), .SI(n8624), .SE(n5052), .CLK(n5466), .Q(
        n8623) );
  SDFFX1 DFF_406_Q_reg ( .D(n157), .SI(n8623), .SE(n5052), .CLK(n5466), .Q(
        n8622) );
  SDFFX1 DFF_407_Q_reg ( .D(n158), .SI(n8622), .SE(n5052), .CLK(n5466), .Q(
        n8621) );
  SDFFX1 DFF_408_Q_reg ( .D(n159), .SI(n8621), .SE(n5052), .CLK(n5466), .Q(
        n8620) );
  SDFFX1 DFF_409_Q_reg ( .D(n160), .SI(n8620), .SE(n5052), .CLK(n5466), .Q(
        n8619) );
  SDFFX1 DFF_410_Q_reg ( .D(n161), .SI(n8619), .SE(n5053), .CLK(n5466), .Q(
        n8618) );
  SDFFX1 DFF_411_Q_reg ( .D(n162), .SI(n8618), .SE(n5053), .CLK(n5466), .Q(
        n8617) );
  SDFFX1 DFF_412_Q_reg ( .D(n163), .SI(n8617), .SE(n5053), .CLK(n5466), .Q(
        n8616) );
  SDFFX1 DFF_413_Q_reg ( .D(n164), .SI(n8616), .SE(n5053), .CLK(n5466), .Q(
        test_so23) );
  SDFFX1 DFF_414_Q_reg ( .D(n165), .SI(test_si24), .SE(n5053), .CLK(n5466), 
        .Q(n8613) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n5053), .CLK(n5466), .Q(
        n8612) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n5048), .CLK(n5468), .Q(
        n8611), .QN(n9693) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n5048), .CLK(n5468), .Q(
        n8610), .QN(n9690) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n5048), .CLK(n5468), .Q(
        n8609), .QN(n9688) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n5047), .CLK(n5469), .Q(
        n8608), .QN(n9686) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n5047), .CLK(n5469), .Q(
        n8607), .QN(n9684) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n5046), .CLK(n5469), .Q(
        n8606), .QN(n9680) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n5046), .CLK(n5469), .Q(
        n8605), .QN(n9678) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n5045), .CLK(n5470), .Q(
        n8604), .QN(n9676) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n5045), .CLK(n5470), .Q(
        n8603), .QN(n9674) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n5044), .CLK(n5470), .Q(
        n8602), .QN(n9672) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n5044), .CLK(n5470), .Q(
        n8601), .QN(n9671) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n5043), .CLK(n5471), .Q(
        n8600), .QN(n9669) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n5043), .CLK(n5471), .Q(
        n8599), .QN(n9667) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n5042), .CLK(n5471), .Q(
        n8598), .QN(n9665) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n5041), .CLK(n5472), .Q(
        n8597), .QN(n9661) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n5016), .CLK(n5484), .Q(
        test_so24), .QN(n4710) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n5040), .CLK(n5472), 
        .Q(WX3263) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n5040), .CLK(n5472), .Q(
        WX3265) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n5039), .CLK(n5473), .Q(
        WX3267) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n5038), .CLK(n5473), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n5038), .CLK(n5473), .Q(
        WX3271) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n5037), .CLK(n5474), .Q(
        WX3273) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n5036), .CLK(n5474), .Q(
        WX3275) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n5036), .CLK(n5474), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n5035), .CLK(n5475), .Q(
        WX3279) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n5034), .CLK(n5475), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n5034), .CLK(n5475), .Q(
        WX3283) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n5033), .CLK(n5476), .Q(
        WX3285) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n5032), .CLK(n5476), .Q(
        WX3287) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n5032), .CLK(n5476), .Q(
        WX3289) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n5031), .CLK(n5477), .Q(
        WX3291) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n5030), .CLK(n5477), .Q(
        WX3293) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n5048), .CLK(n5468), .Q(
        WX3295), .QN(n4037) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n5048), .CLK(n5468), .Q(
        test_so25), .QN(n9691) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n5047), .CLK(n5469), 
        .Q(WX3299), .QN(n4130) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n5047), .CLK(n5469), .Q(
        WX3301), .QN(n4129) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n5047), .CLK(n5469), .Q(
        WX3303), .QN(n4128) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n5047), .CLK(n5469), .Q(
        WX3305), .QN(n9682) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n5046), .CLK(n5469), .Q(
        WX3307), .QN(n4127) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n5046), .CLK(n5469), .Q(
        WX3309), .QN(n4126) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n5045), .CLK(n5470), .Q(
        WX3311) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n5045), .CLK(n5470), .Q(
        WX3313), .QN(n4124) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n5044), .CLK(n5470), .Q(
        WX3315), .QN(n4123) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n5043), .CLK(n5471), .Q(
        WX3317), .QN(n4122) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n5043), .CLK(n5471), .Q(
        WX3319), .QN(n4121) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n5042), .CLK(n5471), .Q(
        WX3321), .QN(n4120) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n5041), .CLK(n5472), .Q(
        WX3323), .QN(n4119) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n5041), .CLK(n5472), .Q(
        WX3325) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n5040), .CLK(n5472), .Q(
        WX3327), .QN(n9658) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n5039), .CLK(n5473), .Q(
        WX3329), .QN(n9656) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n5039), .CLK(n5473), .Q(
        WX3331), .QN(n9654) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n5038), .CLK(n5473), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n5037), .CLK(n5474), 
        .Q(WX3335), .QN(n9650) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n5037), .CLK(n5474), .Q(
        WX3337), .QN(n9648) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n5036), .CLK(n5474), .Q(
        WX3339), .QN(n9646) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n5035), .CLK(n5475), .Q(
        WX3341), .QN(n9644) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n5035), .CLK(n5475), .Q(
        WX3343), .QN(n9642) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n5034), .CLK(n5475), .Q(
        WX3345), .QN(n9640) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n5033), .CLK(n5476), .Q(
        WX3347), .QN(n9638) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n5033), .CLK(n5476), .Q(
        WX3349), .QN(n9636) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n5032), .CLK(n5476), .Q(
        WX3351), .QN(n9634) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n5031), .CLK(n5477), .Q(
        WX3353), .QN(n9632) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n5031), .CLK(n5477), .Q(
        WX3355), .QN(n9630) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n5030), .CLK(n5477), .Q(
        WX3357), .QN(n9628) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n5030), .CLK(n5477), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n5029), .CLK(n5478), .Q(
        WX3361), .QN(n9692) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n5029), .CLK(n5478), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n5029), .CLK(n5478), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n5028), .CLK(n5478), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n5028), .CLK(n5478), .Q(
        test_so27), .QN(n9681) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n5046), .CLK(n5469), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n5046), .CLK(n5469), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n5045), .CLK(n5470), .Q(
        WX3375), .QN(n4125) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n5045), .CLK(n5470), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n5044), .CLK(n5470), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n5043), .CLK(n5471), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n5042), .CLK(n5471), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n5042), .CLK(n5471), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n5041), .CLK(n5472), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n5041), .CLK(n5472), .Q(
        WX3389), .QN(n4118) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n5040), .CLK(n5472), .Q(
        WX3391), .QN(n4349) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n5039), .CLK(n5473), .Q(
        WX3393), .QN(n4347) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n5039), .CLK(n5473), .Q(
        WX3395), .QN(n4345) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n5038), .CLK(n5473), .Q(
        WX3397), .QN(n9652) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n5037), .CLK(n5474), .Q(
        WX3399), .QN(n4342) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n5037), .CLK(n5474), .Q(
        WX3401), .QN(n4340) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n5036), .CLK(n5474), .Q(
        WX3403), .QN(n4338) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n5035), .CLK(n5475), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n5035), .CLK(n5475), 
        .Q(WX3407), .QN(n4335) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n5034), .CLK(n5475), .Q(
        WX3409), .QN(n4333) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n5033), .CLK(n5476), .Q(
        WX3411), .QN(n4331) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n5033), .CLK(n5476), .Q(
        WX3413), .QN(n4329) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n5032), .CLK(n5476), .Q(
        WX3415), .QN(n4327) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n5031), .CLK(n5477), .Q(
        WX3417), .QN(n4325) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n5031), .CLK(n5477), .Q(
        WX3419), .QN(n4323) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n5030), .CLK(n5477), .Q(
        WX3421), .QN(n4321) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n5029), .CLK(n5478), .Q(
        WX3423), .QN(n4577) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n5029), .CLK(n5478), .Q(
        WX3425), .QN(n4578) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n5029), .CLK(n5478), .Q(
        WX3427), .QN(n4579) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n5028), .CLK(n5478), .Q(
        WX3429), .QN(n4580) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n5028), .CLK(n5478), .Q(
        WX3431), .QN(n4581) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n5028), .CLK(n5478), .Q(
        WX3433), .QN(n4582) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n5028), .CLK(n5478), .Q(
        WX3435), .QN(n4583) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n5027), .CLK(n5479), .Q(
        WX3437), .QN(n4584) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n5027), .CLK(n5479), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n5044), .CLK(n5470), 
        .Q(WX3441), .QN(n4585) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n5044), .CLK(n5470), .Q(
        WX3443), .QN(n4586) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n5043), .CLK(n5471), .Q(
        WX3445), .QN(n4587) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n5042), .CLK(n5471), .Q(
        WX3447), .QN(n4588) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n5042), .CLK(n5471), .Q(
        WX3449), .QN(n4589) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n5041), .CLK(n5472), .Q(
        WX3451), .QN(n4590) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n5040), .CLK(n5472), .Q(
        WX3453), .QN(n4403) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n5040), .CLK(n5472), .Q(
        WX3455), .QN(n4591) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n5039), .CLK(n5473), .Q(
        WX3457), .QN(n4592) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n5038), .CLK(n5473), .Q(
        WX3459), .QN(n4593) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n5038), .CLK(n5473), .Q(
        WX3461), .QN(n4594) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n5037), .CLK(n5474), .Q(
        WX3463), .QN(n4404) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n5036), .CLK(n5474), .Q(
        WX3465), .QN(n4595) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n5036), .CLK(n5474), .Q(
        WX3467), .QN(n4596) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n5035), .CLK(n5475), .Q(
        WX3469), .QN(n4597) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n5034), .CLK(n5475), .Q(
        WX3471), .QN(n4598) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n5034), .CLK(n5475), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n5033), .CLK(n5476), 
        .Q(WX3475), .QN(n4599) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n5032), .CLK(n5476), .Q(
        WX3477), .QN(n4405) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n5032), .CLK(n5476), .Q(
        WX3479), .QN(n4600) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n5031), .CLK(n5477), .Q(
        WX3481), .QN(n4601) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n5030), .CLK(n5477), .Q(
        WX3483), .QN(n4602) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n5030), .CLK(n5477), .Q(
        WX3485), .QN(n4415) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n5021), .CLK(n5482), .Q(
        CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n5021), .CLK(n5482), 
        .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n5020), .CLK(n5482), 
        .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n5019), .CLK(n5483), 
        .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n5019), .CLK(n5483), 
        .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n5019), .CLK(n5483), 
        .Q(test_so31), .QN(n4705) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n5019), .CLK(n5483), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n5019), .CLK(n5483), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n5019), .CLK(n5483), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n5018), .CLK(n5483), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n5017), .CLK(n5484), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n5027), .CLK(n5479), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n5027), .CLK(n5479), .Q(test_so32), .QN(n4702) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n5027), .CLK(n5479), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n5027), .CLK(n5479), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n5026), .CLK(n5479), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n5026), .CLK(n5479), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n185), .SI(CRC_OUT_7_31), .SE(n5026), .CLK(n5479), 
        .Q(WX4364), .QN(n4385) );
  SDFFX1 DFF_577_Q_reg ( .D(n186), .SI(WX4364), .SE(n5021), .CLK(n5482), .Q(
        n8586) );
  SDFFX1 DFF_578_Q_reg ( .D(n187), .SI(n8586), .SE(n5021), .CLK(n5482), .Q(
        n8585) );
  SDFFX1 DFF_579_Q_reg ( .D(n188), .SI(n8585), .SE(n5021), .CLK(n5482), .Q(
        n8584) );
  SDFFX1 DFF_580_Q_reg ( .D(n189), .SI(n8584), .SE(n5021), .CLK(n5482), .Q(
        n8583) );
  SDFFX1 DFF_581_Q_reg ( .D(n190), .SI(n8583), .SE(n5022), .CLK(n5481), .Q(
        n8582) );
  SDFFX1 DFF_582_Q_reg ( .D(n191), .SI(n8582), .SE(n5022), .CLK(n5481), .Q(
        n8581) );
  SDFFX1 DFF_583_Q_reg ( .D(n192), .SI(n8581), .SE(n5022), .CLK(n5481), .Q(
        n8580) );
  SDFFX1 DFF_584_Q_reg ( .D(n193), .SI(n8580), .SE(n5022), .CLK(n5481), .Q(
        n8579) );
  SDFFX1 DFF_585_Q_reg ( .D(n194), .SI(n8579), .SE(n5022), .CLK(n5481), .Q(
        n8578) );
  SDFFX1 DFF_586_Q_reg ( .D(n195), .SI(n8578), .SE(n5022), .CLK(n5481), .Q(
        n8577) );
  SDFFX1 DFF_587_Q_reg ( .D(n196), .SI(n8577), .SE(n5023), .CLK(n5481), .Q(
        n8576) );
  SDFFX1 DFF_588_Q_reg ( .D(n197), .SI(n8576), .SE(n5023), .CLK(n5481), .Q(
        test_so33) );
  SDFFX1 DFF_589_Q_reg ( .D(n198), .SI(test_si34), .SE(n5023), .CLK(n5481), 
        .Q(n8573) );
  SDFFX1 DFF_590_Q_reg ( .D(n199), .SI(n8573), .SE(n5023), .CLK(n5481), .Q(
        n8572) );
  SDFFX1 DFF_591_Q_reg ( .D(n200), .SI(n8572), .SE(n5023), .CLK(n5481), .Q(
        n8571) );
  SDFFX1 DFF_592_Q_reg ( .D(n201), .SI(n8571), .SE(n5023), .CLK(n5481), .Q(
        n8570) );
  SDFFX1 DFF_593_Q_reg ( .D(n202), .SI(n8570), .SE(n5024), .CLK(n5480), .Q(
        n8569) );
  SDFFX1 DFF_594_Q_reg ( .D(n203), .SI(n8569), .SE(n5024), .CLK(n5480), .Q(
        n8568) );
  SDFFX1 DFF_595_Q_reg ( .D(n204), .SI(n8568), .SE(n5024), .CLK(n5480), .Q(
        n8567) );
  SDFFX1 DFF_596_Q_reg ( .D(n205), .SI(n8567), .SE(n5024), .CLK(n5480), .Q(
        n8566) );
  SDFFX1 DFF_597_Q_reg ( .D(n206), .SI(n8566), .SE(n5024), .CLK(n5480), .Q(
        n8565) );
  SDFFX1 DFF_598_Q_reg ( .D(n207), .SI(n8565), .SE(n5024), .CLK(n5480), .Q(
        n8564) );
  SDFFX1 DFF_599_Q_reg ( .D(n208), .SI(n8564), .SE(n5025), .CLK(n5480), .Q(
        n8563) );
  SDFFX1 DFF_600_Q_reg ( .D(n209), .SI(n8563), .SE(n5025), .CLK(n5480), .Q(
        n8562) );
  SDFFX1 DFF_601_Q_reg ( .D(n210), .SI(n8562), .SE(n5025), .CLK(n5480), .Q(
        n8561) );
  SDFFX1 DFF_602_Q_reg ( .D(n211), .SI(n8561), .SE(n5025), .CLK(n5480), .Q(
        n8560) );
  SDFFX1 DFF_603_Q_reg ( .D(n212), .SI(n8560), .SE(n5025), .CLK(n5480), .Q(
        n8559) );
  SDFFX1 DFF_604_Q_reg ( .D(n213), .SI(n8559), .SE(n5025), .CLK(n5480), .Q(
        n8558) );
  SDFFX1 DFF_605_Q_reg ( .D(n214), .SI(n8558), .SE(n5026), .CLK(n5479), .Q(
        test_so34) );
  SDFFX1 DFF_606_Q_reg ( .D(n215), .SI(test_si35), .SE(n5026), .CLK(n5479), 
        .Q(n8555) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n5026), .CLK(n5479), .Q(
        n8554) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n4830), .CLK(n5577), .Q(
        n8553), .QN(n9626) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n5005), .CLK(n5490), .Q(
        n8552), .QN(n9623) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n5004), .CLK(n5490), .Q(
        n8551), .QN(n9622) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n5004), .CLK(n5490), .Q(
        n8550), .QN(n9621) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n5002), .CLK(n5491), .Q(
        n8549), .QN(n9620) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n5002), .CLK(n5491), .Q(
        n8548), .QN(n9619) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n5001), .CLK(n5492), .Q(
        n8547), .QN(n9618) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n5001), .CLK(n5492), .Q(
        n8546), .QN(n9617) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n5000), .CLK(n5492), .Q(
        n8545), .QN(n9616) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n5000), .CLK(n5492), .Q(
        n8544), .QN(n9615) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n4998), .CLK(n5493), .Q(
        n8543), .QN(n9614) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n4998), .CLK(n5493), .Q(
        n8542), .QN(n9613) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n4997), .CLK(n5494), .Q(
        n8541), .QN(n9612) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n4997), .CLK(n5494), .Q(
        n8540), .QN(n9611) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n5015), .CLK(n5485), .Q(
        test_so35), .QN(n4709) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n5015), .CLK(n5485), 
        .Q(n8537), .QN(n9610) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n5015), .CLK(n5485), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n5014), .CLK(n5485), .Q(
        WX4558) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n5014), .CLK(n5485), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n5014), .CLK(n5485), .Q(
        WX4562) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n5013), .CLK(n5486), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n5013), .CLK(n5486), .Q(
        WX4566) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n5012), .CLK(n5486), .Q(
        WX4568) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n5011), .CLK(n5487), .Q(
        WX4570) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n5011), .CLK(n5487), .Q(
        WX4572) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n5010), .CLK(n5487), .Q(
        WX4574) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n5009), .CLK(n5488), .Q(
        WX4576) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n5009), .CLK(n5488), .Q(
        WX4578) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n5008), .CLK(n5488), .Q(
        WX4580) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n5007), .CLK(n5489), .Q(
        WX4582) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n5007), .CLK(n5489), .Q(
        WX4584) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n5006), .CLK(n5489), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n4830), .CLK(n5577), 
        .Q(WX4588), .QN(n4036) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n5004), .CLK(n5490), .Q(
        WX4590), .QN(n9625) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n5004), .CLK(n5490), .Q(
        WX4592), .QN(n4117) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n5003), .CLK(n5491), .Q(
        WX4594) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n5003), .CLK(n5491), .Q(
        WX4596), .QN(n4115) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n5002), .CLK(n5491), .Q(
        WX4598), .QN(n4114) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n5002), .CLK(n5491), .Q(
        WX4600), .QN(n4113) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n5001), .CLK(n5492), .Q(
        WX4602), .QN(n4112) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n5000), .CLK(n5492), .Q(
        WX4604), .QN(n4111) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n4999), .CLK(n5493), .Q(
        WX4606), .QN(n4110) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n4999), .CLK(n5493), .Q(
        WX4608), .QN(n4109) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n4998), .CLK(n5493), .Q(
        WX4610), .QN(n4108) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n4998), .CLK(n5493), .Q(
        WX4612), .QN(n4107) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n4997), .CLK(n5494), .Q(
        WX4614), .QN(n4106) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n5015), .CLK(n5485), .Q(
        WX4616) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n5015), .CLK(n5485), .Q(
        WX4618), .QN(n4104) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n5014), .CLK(n5485), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n5014), .CLK(n5485), 
        .Q(WX4622), .QN(n9608) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n5014), .CLK(n5485), .Q(
        WX4624), .QN(n9607) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n5013), .CLK(n5486), .Q(
        WX4626), .QN(n9606) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n5013), .CLK(n5486), .Q(
        WX4628), .QN(n9605) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n5012), .CLK(n5486), .Q(
        WX4630), .QN(n9604) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n5012), .CLK(n5486), .Q(
        WX4632), .QN(n9603) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n5011), .CLK(n5487), .Q(
        WX4634), .QN(n9602) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n5010), .CLK(n5487), .Q(
        WX4636), .QN(n9601) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n5010), .CLK(n5487), .Q(
        WX4638), .QN(n9600) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n5009), .CLK(n5488), .Q(
        WX4640), .QN(n9599) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n5008), .CLK(n5488), .Q(
        WX4642), .QN(n9598) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n5008), .CLK(n5488), .Q(
        WX4644), .QN(n9597) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n5007), .CLK(n5489), .Q(
        WX4646), .QN(n9596) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n5006), .CLK(n5489), .Q(
        WX4648), .QN(n9595) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n5006), .CLK(n5489), .Q(
        WX4650), .QN(n9594) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n5005), .CLK(n5490), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n5005), .CLK(n5490), .Q(
        test_so38), .QN(n9624) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n5004), .CLK(n5490), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n5003), .CLK(n5491), .Q(
        WX4658), .QN(n4116) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n5003), .CLK(n5491), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n5002), .CLK(n5491), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n5001), .CLK(n5492), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n5001), .CLK(n5492), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n5000), .CLK(n5492), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n4999), .CLK(n5493), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n4999), .CLK(n5493), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n4998), .CLK(n5493), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n4997), .CLK(n5494), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n4997), .CLK(n5494), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n4996), .CLK(n5494), .Q(
        WX4680), .QN(n4105) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n4996), .CLK(n5494), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n4996), .CLK(n5494), .Q(
        WX4684), .QN(n9609) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n4995), .CLK(n5495), .Q(
        WX4686), .QN(n4318) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n4995), .CLK(n5495), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n5013), .CLK(n5486), 
        .Q(WX4690), .QN(n4315) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n5013), .CLK(n5486), .Q(
        WX4692), .QN(n4313) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n5012), .CLK(n5486), .Q(
        WX4694), .QN(n4311) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n5012), .CLK(n5486), .Q(
        WX4696), .QN(n4309) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n5011), .CLK(n5487), .Q(
        WX4698), .QN(n4307) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n5010), .CLK(n5487), .Q(
        WX4700), .QN(n4305) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n5010), .CLK(n5487), .Q(
        WX4702), .QN(n4303) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n5009), .CLK(n5488), .Q(
        WX4704), .QN(n4301) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n5008), .CLK(n5488), .Q(
        WX4706), .QN(n4299) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n5008), .CLK(n5488), .Q(
        WX4708), .QN(n4297) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n5007), .CLK(n5489), .Q(
        WX4710), .QN(n4295) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n5006), .CLK(n5489), .Q(
        WX4712), .QN(n4293) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n5006), .CLK(n5489), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n5005), .CLK(n5490), .Q(
        WX4716), .QN(n4550) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n5005), .CLK(n5490), .Q(
        WX4718), .QN(n4551) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n5004), .CLK(n5490), .Q(
        WX4720), .QN(n4552) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n5003), .CLK(n5491), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n5003), .CLK(n5491), 
        .Q(WX4724), .QN(n4553) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n5002), .CLK(n5491), .Q(
        WX4726), .QN(n4554) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n5001), .CLK(n5492), .Q(
        WX4728), .QN(n4555) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n5000), .CLK(n5492), .Q(
        WX4730), .QN(n4556) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n5000), .CLK(n5492), .Q(
        WX4732), .QN(n4557) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n4999), .CLK(n5493), .Q(
        WX4734), .QN(n4558) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n4999), .CLK(n5493), .Q(
        WX4736), .QN(n4559) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n4998), .CLK(n5493), .Q(
        WX4738), .QN(n4560) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n4997), .CLK(n5494), .Q(
        WX4740), .QN(n4561) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n4996), .CLK(n5494), .Q(
        WX4742), .QN(n4562) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n4996), .CLK(n5494), .Q(
        WX4744), .QN(n4563) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n4996), .CLK(n5494), .Q(
        WX4746), .QN(n4401) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n4995), .CLK(n5495), .Q(
        WX4748), .QN(n4564) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n4995), .CLK(n5495), .Q(
        WX4750), .QN(n4565) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n4995), .CLK(n5495), .Q(
        WX4752), .QN(n4566) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n4995), .CLK(n5495), .Q(
        WX4754), .QN(n4567) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n4994), .CLK(n5495), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n5012), .CLK(n5486), 
        .Q(WX4758), .QN(n4568) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n5011), .CLK(n5487), .Q(
        WX4760), .QN(n4569) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n5011), .CLK(n5487), .Q(
        WX4762), .QN(n4570) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n5010), .CLK(n5487), .Q(
        WX4764), .QN(n4571) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n5009), .CLK(n5488), .Q(
        WX4766), .QN(n4572) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n5009), .CLK(n5488), .Q(
        WX4768), .QN(n4573) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n5008), .CLK(n5488), .Q(
        WX4770), .QN(n4402) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n5007), .CLK(n5489), .Q(
        WX4772), .QN(n4574) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n5007), .CLK(n5489), .Q(
        WX4774), .QN(n4575) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n5006), .CLK(n5489), .Q(
        WX4776), .QN(n4576) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n5005), .CLK(n5490), .Q(
        WX4778), .QN(n4414) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n4832), .CLK(n5576), .Q(
        CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n4832), .CLK(n5576), 
        .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n4832), .CLK(n5576), 
        .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n4832), .CLK(n5576), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n4831), .CLK(n5577), 
        .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n4831), .CLK(n5577), 
        .Q(test_so42), .QN(n4700) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n4831), .CLK(n5577), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n4831), .CLK(n5577), 
        .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n4831), .CLK(n5577), 
        .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n4831), .CLK(n5577), 
        .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n4830), .CLK(n5577), 
        .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n4830), .CLK(n5577), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n4830), .CLK(n5577), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n4994), .CLK(n5495), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n4994), .CLK(n5495), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n4994), .CLK(n5495), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n4994), .CLK(n5495), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n4994), .CLK(n5495), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n4993), .CLK(n5496), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n4993), .CLK(n5496), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n4993), .CLK(n5496), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n4993), .CLK(n5496), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n4993), .CLK(n5496), .Q(test_so43), .QN(n4701) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n4993), .CLK(n5496), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n4992), .CLK(n5496), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n4991), .CLK(n5497), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n4991), .CLK(n5497), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n235), .SI(CRC_OUT_6_31), .SE(n4991), .CLK(n5497), 
        .Q(WX5657), .QN(n4384) );
  SDFFX1 DFF_769_Q_reg ( .D(n236), .SI(WX5657), .SE(n4986), .CLK(n5499), .Q(
        n8528) );
  SDFFX1 DFF_770_Q_reg ( .D(n237), .SI(n8528), .SE(n4986), .CLK(n5499), .Q(
        n8527) );
  SDFFX1 DFF_771_Q_reg ( .D(n238), .SI(n8527), .SE(n4986), .CLK(n5499), .Q(
        n8526) );
  SDFFX1 DFF_772_Q_reg ( .D(n239), .SI(n8526), .SE(n4986), .CLK(n5499), .Q(
        n8525) );
  SDFFX1 DFF_773_Q_reg ( .D(n240), .SI(n8525), .SE(n4987), .CLK(n5499), .Q(
        n8524) );
  SDFFX1 DFF_774_Q_reg ( .D(n241), .SI(n8524), .SE(n4987), .CLK(n5499), .Q(
        n8523) );
  SDFFX1 DFF_775_Q_reg ( .D(n242), .SI(n8523), .SE(n4987), .CLK(n5499), .Q(
        test_so44) );
  SDFFX1 DFF_776_Q_reg ( .D(n243), .SI(test_si45), .SE(n4987), .CLK(n5499), 
        .Q(n8520) );
  SDFFX1 DFF_777_Q_reg ( .D(n244), .SI(n8520), .SE(n4987), .CLK(n5499), .Q(
        n8519) );
  SDFFX1 DFF_778_Q_reg ( .D(n245), .SI(n8519), .SE(n4987), .CLK(n5499), .Q(
        n8518) );
  SDFFX1 DFF_779_Q_reg ( .D(n246), .SI(n8518), .SE(n4988), .CLK(n5498), .Q(
        n8517) );
  SDFFX1 DFF_780_Q_reg ( .D(n247), .SI(n8517), .SE(n4988), .CLK(n5498), .Q(
        n8516) );
  SDFFX1 DFF_781_Q_reg ( .D(n248), .SI(n8516), .SE(n4988), .CLK(n5498), .Q(
        n8515) );
  SDFFX1 DFF_782_Q_reg ( .D(n249), .SI(n8515), .SE(n4988), .CLK(n5498), .Q(
        n8514) );
  SDFFX1 DFF_783_Q_reg ( .D(n250), .SI(n8514), .SE(n4988), .CLK(n5498), .Q(
        n8513) );
  SDFFX1 DFF_784_Q_reg ( .D(n251), .SI(n8513), .SE(n4988), .CLK(n5498), .Q(
        n8512) );
  SDFFX1 DFF_785_Q_reg ( .D(n252), .SI(n8512), .SE(n4989), .CLK(n5498), .Q(
        n8511) );
  SDFFX1 DFF_786_Q_reg ( .D(n253), .SI(n8511), .SE(n4989), .CLK(n5498), .Q(
        n8510) );
  SDFFX1 DFF_787_Q_reg ( .D(n254), .SI(n8510), .SE(n4989), .CLK(n5498), .Q(
        n8509) );
  SDFFX1 DFF_788_Q_reg ( .D(n255), .SI(n8509), .SE(n4989), .CLK(n5498), .Q(
        n8508) );
  SDFFX1 DFF_789_Q_reg ( .D(n256), .SI(n8508), .SE(n4989), .CLK(n5498), .Q(
        n8507) );
  SDFFX1 DFF_790_Q_reg ( .D(n257), .SI(n8507), .SE(n4989), .CLK(n5498), .Q(
        n8506) );
  SDFFX1 DFF_791_Q_reg ( .D(n258), .SI(n8506), .SE(n4990), .CLK(n5497), .Q(
        n8505) );
  SDFFX1 DFF_792_Q_reg ( .D(n259), .SI(n8505), .SE(n4990), .CLK(n5497), .Q(
        test_so45) );
  SDFFX1 DFF_793_Q_reg ( .D(n260), .SI(test_si46), .SE(n4990), .CLK(n5497), 
        .Q(n8502) );
  SDFFX1 DFF_794_Q_reg ( .D(n261), .SI(n8502), .SE(n4990), .CLK(n5497), .Q(
        n8501) );
  SDFFX1 DFF_795_Q_reg ( .D(n262), .SI(n8501), .SE(n4990), .CLK(n5497), .Q(
        n8500) );
  SDFFX1 DFF_796_Q_reg ( .D(n263), .SI(n8500), .SE(n4990), .CLK(n5497), .Q(
        n8499) );
  SDFFX1 DFF_797_Q_reg ( .D(n264), .SI(n8499), .SE(n4991), .CLK(n5497), .Q(
        n8498) );
  SDFFX1 DFF_798_Q_reg ( .D(n265), .SI(n8498), .SE(n4991), .CLK(n5497), .Q(
        n8497) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n4991), .CLK(n5497), .Q(
        n8496) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n4986), .CLK(n5499), .Q(
        n8495), .QN(n9593) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n4985), .CLK(n5500), .Q(
        n8494), .QN(n9592) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n4985), .CLK(n5500), .Q(
        n8493), .QN(n9591) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n4985), .CLK(n5500), .Q(
        n8492), .QN(n9590) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n4984), .CLK(n5500), .Q(
        n8491), .QN(n9589) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n4984), .CLK(n5500), .Q(
        n8490), .QN(n9588) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n4984), .CLK(n5500), .Q(
        n8489), .QN(n9587) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n4983), .CLK(n5501), .Q(
        n8488), .QN(n9586) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n4983), .CLK(n5501), .Q(
        n8487), .QN(n9585) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n4832), .CLK(n5576), .Q(
        test_so46), .QN(n4708) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n4982), .CLK(n5501), 
        .Q(n8484), .QN(n9584) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n4982), .CLK(n5501), .Q(
        n8483), .QN(n9581) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n4833), .CLK(n5576), .Q(
        n8482), .QN(n9580) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n4981), .CLK(n5502), .Q(
        n8481), .QN(n9577) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n5015), .CLK(n5485), .Q(
        n8480), .QN(n9576) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n4832), .CLK(n5576), .Q(
        n8479), .QN(n9575) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n4980), .CLK(n5502), .Q(
        WX5849) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n4980), .CLK(n5502), .Q(
        WX5851) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n4979), .CLK(n5503), .Q(
        WX5853) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n4978), .CLK(n5503), .Q(
        WX5855) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n4978), .CLK(n5503), .Q(
        WX5857) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n4977), .CLK(n5504), .Q(
        WX5859) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n4976), .CLK(n5504), .Q(
        WX5861) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n4976), .CLK(n5504), .Q(
        WX5863) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n4975), .CLK(n5505), .Q(
        WX5865) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n4974), .CLK(n5505), .Q(
        WX5867) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n4974), .CLK(n5505), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n4973), .CLK(n5506), 
        .Q(WX5871) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n4972), .CLK(n5506), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n4972), .CLK(n5506), .Q(
        WX5875) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n4971), .CLK(n5507), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n4970), .CLK(n5507), .Q(
        WX5879) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n4986), .CLK(n5499), .Q(
        WX5881), .QN(n4035) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n4985), .CLK(n5500), .Q(
        WX5883), .QN(n4103) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n4985), .CLK(n5500), .Q(
        WX5885), .QN(n4102) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n4985), .CLK(n5500), .Q(
        WX5887), .QN(n4101) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n4984), .CLK(n5500), .Q(
        WX5889), .QN(n4100) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n4984), .CLK(n5500), .Q(
        WX5891), .QN(n4099) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n4984), .CLK(n5500), .Q(
        WX5893), .QN(n4098) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n4983), .CLK(n5501), .Q(
        WX5895), .QN(n4097) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n4983), .CLK(n5501), .Q(
        WX5897), .QN(n4096) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n4983), .CLK(n5501), .Q(
        WX5899) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n4983), .CLK(n5501), .Q(
        WX5901), .QN(n4094) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n4982), .CLK(n5501), .Q(
        test_so48), .QN(n9582) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n4833), .CLK(n5576), 
        .Q(WX5905), .QN(n4093) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n4981), .CLK(n5502), .Q(
        WX5907), .QN(n9579) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n4981), .CLK(n5502), .Q(
        WX5909), .QN(n4092) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n4981), .CLK(n5502), .Q(
        WX5911) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n4980), .CLK(n5502), .Q(
        WX5913), .QN(n9574) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n4980), .CLK(n5502), .Q(
        WX5915), .QN(n9573) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n4979), .CLK(n5503), .Q(
        WX5917), .QN(n9572) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n4978), .CLK(n5503), .Q(
        WX5919), .QN(n9571) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n4978), .CLK(n5503), .Q(
        WX5921), .QN(n9570) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n4977), .CLK(n5504), .Q(
        WX5923), .QN(n9569) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n4976), .CLK(n5504), .Q(
        WX5925), .QN(n9568) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n4976), .CLK(n5504), .Q(
        WX5927), .QN(n9567) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n4975), .CLK(n5505), .Q(
        WX5929), .QN(n9566) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n4974), .CLK(n5505), .Q(
        WX5931), .QN(n9565) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n4974), .CLK(n5505), .Q(
        WX5933), .QN(n9564) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n4973), .CLK(n5506), .Q(
        WX5935), .QN(n9563) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n4972), .CLK(n5506), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n4972), .CLK(n5506), 
        .Q(WX5939), .QN(n9561) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n4971), .CLK(n5507), .Q(
        WX5941), .QN(n9560) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n4970), .CLK(n5507), .Q(
        WX5943), .QN(n9559) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n4970), .CLK(n5507), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n4969), .CLK(n5508), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n4969), .CLK(n5508), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n4969), .CLK(n5508), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n4968), .CLK(n5508), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n4968), .CLK(n5508), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n4968), .CLK(n5508), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n4967), .CLK(n5509), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n4967), .CLK(n5509), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n4967), .CLK(n5509), .Q(
        WX5963), .QN(n4095) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n4966), .CLK(n5509), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n4982), .CLK(n5501), .Q(
        WX5967), .QN(n9583) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n4982), .CLK(n5501), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n4982), .CLK(n5501), .Q(
        test_so50), .QN(n9578) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n4981), .CLK(n5502), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n4981), .CLK(n5502), .Q(
        WX5975), .QN(n4091) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n4980), .CLK(n5502), .Q(
        WX5977), .QN(n4290) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n4979), .CLK(n5503), .Q(
        WX5979), .QN(n4288) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n4979), .CLK(n5503), .Q(
        WX5981), .QN(n4286) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n4978), .CLK(n5503), .Q(
        WX5983), .QN(n4284) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n4977), .CLK(n5504), .Q(
        WX5985), .QN(n4282) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n4977), .CLK(n5504), .Q(
        WX5987), .QN(n4280) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n4976), .CLK(n5504), .Q(
        WX5989), .QN(n4278) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n4975), .CLK(n5505), .Q(
        WX5991), .QN(n4276) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n4975), .CLK(n5505), .Q(
        WX5993), .QN(n4274) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n4974), .CLK(n5505), .Q(
        WX5995), .QN(n4272) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n4973), .CLK(n5506), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n4973), .CLK(n5506), .Q(
        WX5999), .QN(n4269) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n4972), .CLK(n5506), .Q(
        WX6001), .QN(n9562) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n4971), .CLK(n5507), .Q(
        WX6003), .QN(n4266) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n4971), .CLK(n5507), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n4970), .CLK(n5507), 
        .Q(WX6007), .QN(n4263) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n4970), .CLK(n5507), .Q(
        WX6009), .QN(n4522) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n4969), .CLK(n5508), .Q(
        WX6011), .QN(n4523) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n4969), .CLK(n5508), .Q(
        WX6013), .QN(n4524) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n4969), .CLK(n5508), .Q(
        WX6015), .QN(n4525) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n4968), .CLK(n5508), .Q(
        WX6017), .QN(n4526) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n4968), .CLK(n5508), .Q(
        WX6019), .QN(n4527) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n4968), .CLK(n5508), .Q(
        WX6021), .QN(n4528) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n4967), .CLK(n5509), .Q(
        WX6023), .QN(n4529) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n4967), .CLK(n5509), .Q(
        WX6025), .QN(n4530) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n4967), .CLK(n5509), .Q(
        WX6027), .QN(n4531) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n4966), .CLK(n5509), .Q(
        WX6029), .QN(n4532) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n4966), .CLK(n5509), .Q(
        WX6031), .QN(n4533) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n4966), .CLK(n5509), .Q(
        WX6033), .QN(n4534) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n4966), .CLK(n5509), .Q(
        WX6035), .QN(n4535) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n4966), .CLK(n5509), .Q(
        WX6037), .QN(n4536) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n4965), .CLK(n5510), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n4980), .CLK(n5502), 
        .Q(WX6041), .QN(n4537) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n4979), .CLK(n5503), .Q(
        WX6043), .QN(n4538) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n4979), .CLK(n5503), .Q(
        WX6045), .QN(n4539) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n4978), .CLK(n5503), .Q(
        WX6047), .QN(n4540) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n4977), .CLK(n5504), .Q(
        WX6049), .QN(n4399) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n4977), .CLK(n5504), .Q(
        WX6051), .QN(n4541) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n4976), .CLK(n5504), .Q(
        WX6053), .QN(n4542) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n4975), .CLK(n5505), .Q(
        WX6055), .QN(n4543) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n4975), .CLK(n5505), .Q(
        WX6057), .QN(n4544) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n4974), .CLK(n5505), .Q(
        WX6059), .QN(n4545) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n4973), .CLK(n5506), .Q(
        WX6061), .QN(n4546) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n4973), .CLK(n5506), .Q(
        WX6063), .QN(n4400) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n4972), .CLK(n5506), .Q(
        WX6065), .QN(n4547) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n4971), .CLK(n5507), .Q(
        WX6067), .QN(n4548) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n4971), .CLK(n5507), .Q(
        WX6069), .QN(n4549) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n4970), .CLK(n5507), .Q(
        WX6071), .QN(n4413) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n4836), .CLK(n5574), .Q(
        test_so53), .QN(n4698) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n4836), .CLK(n5574), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n4836), .CLK(n5574), 
        .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n4836), .CLK(n5574), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n4836), .CLK(n5574), 
        .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n4835), .CLK(n5575), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n4834), .CLK(n5575), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n4833), .CLK(n5576), .Q(test_so54), .QN(n4699) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n4833), .CLK(n5576), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n4833), .CLK(n5576), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n4833), .CLK(n5576), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n4965), .CLK(n5510), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n4965), .CLK(n5510), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n4965), .CLK(n5510), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n4965), .CLK(n5510), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n4965), .CLK(n5510), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n4964), .CLK(n5510), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n285), .SI(CRC_OUT_5_31), .SE(n4963), .CLK(n5511), 
        .Q(WX6950), .QN(n4383) );
  SDFFX1 DFF_961_Q_reg ( .D(n286), .SI(WX6950), .SE(n4958), .CLK(n5513), .Q(
        n8470) );
  SDFFX1 DFF_962_Q_reg ( .D(n287), .SI(n8470), .SE(n4958), .CLK(n5513), .Q(
        test_so55) );
  SDFFX1 DFF_963_Q_reg ( .D(n288), .SI(test_si56), .SE(n4959), .CLK(n5513), 
        .Q(n8467) );
  SDFFX1 DFF_964_Q_reg ( .D(n289), .SI(n8467), .SE(n4959), .CLK(n5513), .Q(
        n8466) );
  SDFFX1 DFF_965_Q_reg ( .D(n290), .SI(n8466), .SE(n4959), .CLK(n5513), .Q(
        n8465) );
  SDFFX1 DFF_966_Q_reg ( .D(n291), .SI(n8465), .SE(n4959), .CLK(n5513), .Q(
        n8464) );
  SDFFX1 DFF_967_Q_reg ( .D(n292), .SI(n8464), .SE(n4959), .CLK(n5513), .Q(
        n8463) );
  SDFFX1 DFF_968_Q_reg ( .D(n293), .SI(n8463), .SE(n4959), .CLK(n5513), .Q(
        n8462) );
  SDFFX1 DFF_969_Q_reg ( .D(n294), .SI(n8462), .SE(n4960), .CLK(n5512), .Q(
        n8461) );
  SDFFX1 DFF_970_Q_reg ( .D(n295), .SI(n8461), .SE(n4960), .CLK(n5512), .Q(
        n8460) );
  SDFFX1 DFF_971_Q_reg ( .D(n296), .SI(n8460), .SE(n4960), .CLK(n5512), .Q(
        n8459) );
  SDFFX1 DFF_972_Q_reg ( .D(n297), .SI(n8459), .SE(n4960), .CLK(n5512), .Q(
        n8458) );
  SDFFX1 DFF_973_Q_reg ( .D(n298), .SI(n8458), .SE(n4960), .CLK(n5512), .Q(
        n8457) );
  SDFFX1 DFF_974_Q_reg ( .D(n299), .SI(n8457), .SE(n4960), .CLK(n5512), .Q(
        n8456) );
  SDFFX1 DFF_975_Q_reg ( .D(n300), .SI(n8456), .SE(n4961), .CLK(n5512), .Q(
        n8455) );
  SDFFX1 DFF_976_Q_reg ( .D(n301), .SI(n8455), .SE(n4961), .CLK(n5512), .Q(
        n8454) );
  SDFFX1 DFF_977_Q_reg ( .D(n302), .SI(n8454), .SE(n4961), .CLK(n5512), .Q(
        n8453) );
  SDFFX1 DFF_978_Q_reg ( .D(n303), .SI(n8453), .SE(n4961), .CLK(n5512), .Q(
        n8452) );
  SDFFX1 DFF_979_Q_reg ( .D(n304), .SI(n8452), .SE(n4961), .CLK(n5512), .Q(
        test_so56) );
  SDFFX1 DFF_980_Q_reg ( .D(n305), .SI(test_si57), .SE(n4961), .CLK(n5512), 
        .Q(n8449) );
  SDFFX1 DFF_981_Q_reg ( .D(n306), .SI(n8449), .SE(n4962), .CLK(n5511), .Q(
        n8448) );
  SDFFX1 DFF_982_Q_reg ( .D(n307), .SI(n8448), .SE(n4962), .CLK(n5511), .Q(
        n8447) );
  SDFFX1 DFF_983_Q_reg ( .D(n308), .SI(n8447), .SE(n4962), .CLK(n5511), .Q(
        n8446) );
  SDFFX1 DFF_984_Q_reg ( .D(n309), .SI(n8446), .SE(n4962), .CLK(n5511), .Q(
        n8445) );
  SDFFX1 DFF_985_Q_reg ( .D(n149), .SI(n8445), .SE(n4962), .CLK(n5511), .Q(
        n8444) );
  SDFFX1 DFF_986_Q_reg ( .D(n310), .SI(n8444), .SE(n4962), .CLK(n5511), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(n311), .SI(n8443), .SE(n4963), .CLK(n5511), .Q(
        n8442) );
  SDFFX1 DFF_988_Q_reg ( .D(n312), .SI(n8442), .SE(n4963), .CLK(n5511), .Q(
        n8441) );
  SDFFX1 DFF_989_Q_reg ( .D(n313), .SI(n8441), .SE(n4963), .CLK(n5511), .Q(
        n8440) );
  SDFFX1 DFF_990_Q_reg ( .D(n314), .SI(n8440), .SE(n4963), .CLK(n5511), .Q(
        n8439) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n4963), .CLK(n5511), .Q(
        n8438) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n4958), .CLK(n5513), .Q(
        n8437), .QN(n9558) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n4958), .CLK(n5513), .Q(
        n8436), .QN(n9557) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n4957), .CLK(n5514), .Q(
        n8435), .QN(n9556) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n4957), .CLK(n5514), .Q(
        n8434), .QN(n9555) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n4957), .CLK(n5514), .Q(
        test_so57), .QN(n4707) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n4956), .CLK(n5514), 
        .Q(n8431), .QN(n9554) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n4956), .CLK(n5514), .Q(
        n8430), .QN(n9551) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n4837), .CLK(n5574), .Q(
        n8429), .QN(n9550) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n4955), .CLK(n5515), .Q(
        n8428), .QN(n9547) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n4955), .CLK(n5515), .Q(
        n8427), .QN(n9546) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n4954), .CLK(n5515), .Q(
        n8426), .QN(n9545) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n4953), .CLK(n5516), .Q(
        n8425), .QN(n9544) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n4953), .CLK(n5516), .Q(
        n8424), .QN(n9543) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n4836), .CLK(n5574), .Q(
        n8423), .QN(n9542) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n5016), .CLK(n5484), .Q(
        n8422), .QN(n9541) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n4951), .CLK(n5517), .Q(
        n8421), .QN(n9540) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n4951), .CLK(n5517), .Q(
        WX7142) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n4950), .CLK(n5517), 
        .Q(WX7144) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n4950), .CLK(n5517), 
        .Q(WX7146) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n4949), .CLK(n5518), 
        .Q(WX7148) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n4948), .CLK(n5518), 
        .Q(WX7150) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n4948), .CLK(n5518), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n4946), .CLK(n5519), 
        .Q(WX7154) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n4946), .CLK(n5519), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n4946), .CLK(n5519), 
        .Q(WX7158) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n4945), .CLK(n5520), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n4944), .CLK(n5520), 
        .Q(WX7162) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n4944), .CLK(n5520), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n4943), .CLK(n5521), 
        .Q(WX7166) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n4942), .CLK(n5521), 
        .Q(WX7168) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n4942), .CLK(n5521), 
        .Q(WX7170) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n4941), .CLK(n5522), 
        .Q(WX7172) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n4958), .CLK(n5513), 
        .Q(WX7174), .QN(n4034) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n4958), .CLK(n5513), 
        .Q(WX7176), .QN(n4090) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n4957), .CLK(n5514), 
        .Q(WX7178), .QN(n4089) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n4957), .CLK(n5514), 
        .Q(WX7180), .QN(n4088) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n4957), .CLK(n5514), 
        .Q(WX7182) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n4956), .CLK(n5514), 
        .Q(WX7184), .QN(n4086) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n4956), .CLK(n5514), 
        .Q(test_so59), .QN(n9552) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n4837), .CLK(n5574), 
        .Q(WX7188), .QN(n4085) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n4955), .CLK(n5515), 
        .Q(WX7190), .QN(n9549) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n4955), .CLK(n5515), 
        .Q(WX7192), .QN(n4084) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n4954), .CLK(n5515), 
        .Q(WX7194) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n4954), .CLK(n5515), 
        .Q(WX7196), .QN(n4082) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n4953), .CLK(n5516), 
        .Q(WX7198), .QN(n4081) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n4953), .CLK(n5516), 
        .Q(WX7200), .QN(n4080) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n4952), .CLK(n5516), 
        .Q(WX7202), .QN(n4079) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n4952), .CLK(n5516), 
        .Q(WX7204), .QN(n4078) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n4951), .CLK(n5517), 
        .Q(WX7206), .QN(n9539) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n4950), .CLK(n5517), 
        .Q(WX7208), .QN(n9538) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n4949), .CLK(n5518), 
        .Q(WX7210), .QN(n9537) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n4949), .CLK(n5518), 
        .Q(WX7212), .QN(n9536) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n4948), .CLK(n5518), 
        .Q(WX7214), .QN(n9535) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n4947), .CLK(n5519), 
        .Q(WX7216), .QN(n9534) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n4947), .CLK(n5519), 
        .Q(WX7218), .QN(n9533) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n4946), .CLK(n5519), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n4945), .CLK(n5520), 
        .Q(WX7222), .QN(n9531) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n4945), .CLK(n5520), 
        .Q(WX7224), .QN(n9530) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n4944), .CLK(n5520), 
        .Q(WX7226), .QN(n9529) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n4943), .CLK(n5521), 
        .Q(WX7228), .QN(n9528) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n4943), .CLK(n5521), 
        .Q(WX7230), .QN(n9527) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n4942), .CLK(n5521), 
        .Q(WX7232), .QN(n9526) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n4941), .CLK(n5522), 
        .Q(WX7234), .QN(n9525) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n4941), .CLK(n5522), 
        .Q(WX7236), .QN(n9524) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n4940), .CLK(n5522), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n4940), .CLK(n5522), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n4940), .CLK(n5522), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n4939), .CLK(n5523), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n4939), .CLK(n5523), 
        .Q(WX7246), .QN(n4087) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n4939), .CLK(n5523), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n4956), .CLK(n5514), 
        .Q(WX7250), .QN(n9553) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n4956), .CLK(n5514), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n4955), .CLK(n5515), 
        .Q(test_so61), .QN(n9548) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n4955), .CLK(n5515), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n4954), .CLK(n5515), 
        .Q(WX7258), .QN(n4083) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n4954), .CLK(n5515), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n4953), .CLK(n5516), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n4952), .CLK(n5516), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n4952), .CLK(n5516), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n4951), .CLK(n5517), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n4951), .CLK(n5517), 
        .Q(WX7270), .QN(n4261) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n4950), .CLK(n5517), 
        .Q(WX7272), .QN(n4259) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n4949), .CLK(n5518), 
        .Q(WX7274), .QN(n4257) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n4949), .CLK(n5518), 
        .Q(WX7276), .QN(n4255) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n4948), .CLK(n5518), 
        .Q(WX7278), .QN(n4253) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n4947), .CLK(n5519), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n4947), .CLK(n5519), 
        .Q(WX7282), .QN(n4250) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n4946), .CLK(n5519), 
        .Q(WX7284), .QN(n9532) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n4945), .CLK(n5520), 
        .Q(WX7286), .QN(n4247) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n4945), .CLK(n5520), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n4944), .CLK(n5520), 
        .Q(WX7290), .QN(n4244) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n4943), .CLK(n5521), 
        .Q(WX7292), .QN(n4242) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n4943), .CLK(n5521), 
        .Q(WX7294), .QN(n4240) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n4942), .CLK(n5521), 
        .Q(WX7296), .QN(n4238) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n4941), .CLK(n5522), 
        .Q(WX7298), .QN(n4236) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n4941), .CLK(n5522), 
        .Q(WX7300), .QN(n4234) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n4940), .CLK(n5522), 
        .Q(WX7302), .QN(n4495) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n4940), .CLK(n5522), 
        .Q(WX7304), .QN(n4496) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n4939), .CLK(n5523), 
        .Q(WX7306), .QN(n4497) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n4939), .CLK(n5523), 
        .Q(WX7308), .QN(n4498) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n4939), .CLK(n5523), 
        .Q(WX7310), .QN(n4499) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n4938), .CLK(n5523), 
        .Q(WX7312), .QN(n4500) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n4938), .CLK(n5523), 
        .Q(WX7314), .QN(n4501) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n4938), .CLK(n5523), 
        .Q(WX7316), .QN(n4502) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n4938), .CLK(n5523), 
        .Q(WX7318), .QN(n4503) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n4938), .CLK(n5523), 
        .Q(WX7320), .QN(n4504) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n4938), .CLK(n5523), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n4954), .CLK(n5515), 
        .Q(WX7324), .QN(n4505) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n4953), .CLK(n5516), 
        .Q(WX7326), .QN(n4506) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n4952), .CLK(n5516), 
        .Q(WX7328), .QN(n4507) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n4952), .CLK(n5516), 
        .Q(WX7330), .QN(n4508) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n4951), .CLK(n5517), 
        .Q(WX7332), .QN(n4397) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n4950), .CLK(n5517), 
        .Q(WX7334), .QN(n4509) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n4950), .CLK(n5517), 
        .Q(WX7336), .QN(n4510) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n4949), .CLK(n5518), 
        .Q(WX7338), .QN(n4511) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n4948), .CLK(n5518), 
        .Q(WX7340), .QN(n4512) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n4948), .CLK(n5518), 
        .Q(WX7342), .QN(n4398) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n4947), .CLK(n5519), 
        .Q(WX7344), .QN(n4513) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n4947), .CLK(n5519), 
        .Q(WX7346), .QN(n4514) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n4946), .CLK(n5519), 
        .Q(WX7348), .QN(n4515) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n4945), .CLK(n5520), 
        .Q(WX7350), .QN(n4516) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n4944), .CLK(n5520), 
        .Q(WX7352), .QN(n4517) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n4944), .CLK(n5520), 
        .Q(WX7354), .QN(n4518) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n4943), .CLK(n5521), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n4942), .CLK(n5521), 
        .Q(WX7358), .QN(n4519) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n4942), .CLK(n5521), 
        .Q(WX7360), .QN(n4520) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n4941), .CLK(n5522), 
        .Q(WX7362), .QN(n4521) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n4940), .CLK(n5522), 
        .Q(WX7364), .QN(n4412) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n4841), .CLK(n5572), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n4841), .CLK(n5572), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n4841), .CLK(n5572), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n4841), .CLK(n5572), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n4840), .CLK(n5572), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n4839), .CLK(n5573), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n4839), .CLK(
        n5573), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n4839), .CLK(
        n5573), .Q(test_so65), .QN(n4696) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n4839), .CLK(n5573), 
        .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n4839), .CLK(
        n5573), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n4839), .CLK(
        n5573), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n4838), .CLK(
        n5573), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n4837), .CLK(
        n5574), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n4837), .CLK(
        n5574), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n4837), .CLK(
        n5574), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n4837), .CLK(
        n5574), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n4937), .CLK(
        n5524), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n4937), .CLK(
        n5524), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n4937), .CLK(
        n5524), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n4937), .CLK(
        n5524), .Q(test_so66), .QN(n4697) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n4937), .CLK(n5524), 
        .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n4937), .CLK(
        n5524), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n334), .SI(CRC_OUT_4_31), .SE(n4936), .CLK(n5524), 
        .Q(WX8243), .QN(n4382) );
  SDFFX1 DFF_1153_Q_reg ( .D(n335), .SI(WX8243), .SE(n4936), .CLK(n5524), .Q(
        n8411) );
  SDFFX1 DFF_1154_Q_reg ( .D(n336), .SI(n8411), .SE(n4936), .CLK(n5524), .Q(
        n8410) );
  SDFFX1 DFF_1155_Q_reg ( .D(n337), .SI(n8410), .SE(n4936), .CLK(n5524), .Q(
        n8409) );
  SDFFX1 DFF_1156_Q_reg ( .D(n338), .SI(n8409), .SE(n4936), .CLK(n5524), .Q(
        n8408) );
  SDFFX1 DFF_1157_Q_reg ( .D(n339), .SI(n8408), .SE(n4936), .CLK(n5524), .Q(
        n8407) );
  SDFFX1 DFF_1158_Q_reg ( .D(n340), .SI(n8407), .SE(n4935), .CLK(n5525), .Q(
        n8406) );
  SDFFX1 DFF_1159_Q_reg ( .D(n341), .SI(n8406), .SE(n4935), .CLK(n5525), .Q(
        n8405) );
  SDFFX1 DFF_1160_Q_reg ( .D(n342), .SI(n8405), .SE(n4935), .CLK(n5525), .Q(
        n8404) );
  SDFFX1 DFF_1161_Q_reg ( .D(n343), .SI(n8404), .SE(n4935), .CLK(n5525), .Q(
        n8403) );
  SDFFX1 DFF_1162_Q_reg ( .D(n344), .SI(n8403), .SE(n4935), .CLK(n5525), .Q(
        n8402) );
  SDFFX1 DFF_1163_Q_reg ( .D(n345), .SI(n8402), .SE(n4935), .CLK(n5525), .Q(
        n8401) );
  SDFFX1 DFF_1164_Q_reg ( .D(n150), .SI(n8401), .SE(n5016), .CLK(n5484), .Q(
        n8400) );
  SDFFX1 DFF_1165_Q_reg ( .D(n346), .SI(n8400), .SE(n5016), .CLK(n5484), .Q(
        n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(n347), .SI(n8399), .SE(n5016), .CLK(n5484), .Q(
        test_so67) );
  SDFFX1 DFF_1167_Q_reg ( .D(n348), .SI(test_si68), .SE(n4932), .CLK(n5526), 
        .Q(n8396) );
  SDFFX1 DFF_1168_Q_reg ( .D(n349), .SI(n8396), .SE(n4932), .CLK(n5526), .Q(
        n8395) );
  SDFFX1 DFF_1169_Q_reg ( .D(n350), .SI(n8395), .SE(n4932), .CLK(n5526), .Q(
        n8394) );
  SDFFX1 DFF_1170_Q_reg ( .D(n351), .SI(n8394), .SE(n4932), .CLK(n5526), .Q(
        n8393) );
  SDFFX1 DFF_1171_Q_reg ( .D(n352), .SI(n8393), .SE(n4932), .CLK(n5526), .Q(
        n8392) );
  SDFFX1 DFF_1172_Q_reg ( .D(n353), .SI(n8392), .SE(n4933), .CLK(n5526), .Q(
        n8391) );
  SDFFX1 DFF_1173_Q_reg ( .D(n354), .SI(n8391), .SE(n4933), .CLK(n5526), .Q(
        n8390) );
  SDFFX1 DFF_1174_Q_reg ( .D(n355), .SI(n8390), .SE(n4933), .CLK(n5526), .Q(
        n8389) );
  SDFFX1 DFF_1175_Q_reg ( .D(n356), .SI(n8389), .SE(n4933), .CLK(n5526), .Q(
        n8388) );
  SDFFX1 DFF_1176_Q_reg ( .D(n357), .SI(n8388), .SE(n4933), .CLK(n5526), .Q(
        n8387) );
  SDFFX1 DFF_1177_Q_reg ( .D(n358), .SI(n8387), .SE(n4933), .CLK(n5526), .Q(
        n8386) );
  SDFFX1 DFF_1178_Q_reg ( .D(n359), .SI(n8386), .SE(n4934), .CLK(n5525), .Q(
        n8385) );
  SDFFX1 DFF_1179_Q_reg ( .D(n360), .SI(n8385), .SE(n4934), .CLK(n5525), .Q(
        n8384) );
  SDFFX1 DFF_1180_Q_reg ( .D(n361), .SI(n8384), .SE(n4934), .CLK(n5525), .Q(
        n8383) );
  SDFFX1 DFF_1181_Q_reg ( .D(n362), .SI(n8383), .SE(n4934), .CLK(n5525), .Q(
        n8382) );
  SDFFX1 DFF_1182_Q_reg ( .D(n363), .SI(n8382), .SE(n4934), .CLK(n5525), .Q(
        n8381) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n4934), .CLK(n5525), .Q(
        test_so68) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n4922), .CLK(n5531), 
        .Q(n8378), .QN(n9523) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n4922), .CLK(n5531), .Q(
        n8377), .QN(n9520) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n4842), .CLK(n5571), .Q(
        n8376), .QN(n9519) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n4921), .CLK(n5532), .Q(
        n8375), .QN(n9516) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n4920), .CLK(n5532), .Q(
        n8374), .QN(n9515) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n4920), .CLK(n5532), .Q(
        n8373), .QN(n9514) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n4919), .CLK(n5533), .Q(
        n8372), .QN(n9513) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n4918), .CLK(n5533), .Q(
        n8371), .QN(n9512) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n4917), .CLK(n5534), .Q(
        n8370), .QN(n9511) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n4917), .CLK(n5534), .Q(
        n8369), .QN(n9510) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n4916), .CLK(n5534), .Q(
        n8368), .QN(n9509) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n4916), .CLK(n5534), .Q(
        n8367), .QN(n9508) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n4915), .CLK(n5535), .Q(
        n8366), .QN(n9507) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n4914), .CLK(n5535), .Q(
        n8365), .QN(n9506) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n5016), .CLK(n5484), .Q(
        n8364), .QN(n9505) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n4932), .CLK(n5526), .Q(
        n8363), .QN(n9504) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n4841), .CLK(n5572), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n4931), .CLK(n5527), 
        .Q(WX8437) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n4931), .CLK(n5527), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n4930), .CLK(n5527), 
        .Q(WX8441) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n4930), .CLK(n5527), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n4930), .CLK(n5527), 
        .Q(WX8445) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n4929), .CLK(n5528), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n4929), .CLK(n5528), 
        .Q(WX8449) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n4928), .CLK(n5528), 
        .Q(WX8451) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n4927), .CLK(n5529), 
        .Q(WX8453) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n4927), .CLK(n5529), 
        .Q(WX8455) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n4926), .CLK(n5529), 
        .Q(WX8457) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n4925), .CLK(n5530), 
        .Q(WX8459) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n4925), .CLK(n5530), 
        .Q(WX8461) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n4924), .CLK(n5530), 
        .Q(WX8463) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n4923), .CLK(n5531), 
        .Q(WX8465) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n4923), .CLK(n5531), 
        .Q(WX8467), .QN(n4033) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n4922), .CLK(n5531), 
        .Q(test_so70), .QN(n9521) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n4841), .CLK(n5572), 
        .Q(WX8471), .QN(n4077) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n4921), .CLK(n5532), 
        .Q(WX8473), .QN(n9518) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n4920), .CLK(n5532), 
        .Q(WX8475), .QN(n4076) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n4920), .CLK(n5532), 
        .Q(WX8477) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n4919), .CLK(n5533), 
        .Q(WX8479), .QN(n4074) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n4918), .CLK(n5533), 
        .Q(WX8481), .QN(n4073) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n4918), .CLK(n5533), 
        .Q(WX8483), .QN(n4072) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n4917), .CLK(n5534), 
        .Q(WX8485), .QN(n4071) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n4916), .CLK(n5534), 
        .Q(WX8487), .QN(n4070) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n4916), .CLK(n5534), 
        .Q(WX8489), .QN(n4069) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n4915), .CLK(n5535), 
        .Q(WX8491), .QN(n4068) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n4914), .CLK(n5535), 
        .Q(WX8493), .QN(n4067) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n4914), .CLK(n5535), 
        .Q(WX8495), .QN(n4066) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n4931), .CLK(n5527), 
        .Q(WX8497), .QN(n4065) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n4931), .CLK(n5527), 
        .Q(WX8499), .QN(n9503) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n4931), .CLK(n5527), 
        .Q(WX8501), .QN(n9502) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n4931), .CLK(n5527), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n4930), .CLK(n5527), 
        .Q(WX8505), .QN(n9500) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n4930), .CLK(n5527), 
        .Q(WX8507), .QN(n9499) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n4930), .CLK(n5527), 
        .Q(WX8509), .QN(n9498) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n4929), .CLK(n5528), 
        .Q(WX8511), .QN(n9497) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n4929), .CLK(n5528), 
        .Q(WX8513), .QN(n9496) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n4928), .CLK(n5528), 
        .Q(WX8515), .QN(n9495) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n4927), .CLK(n5529), 
        .Q(WX8517), .QN(n9494) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n4927), .CLK(n5529), 
        .Q(WX8519), .QN(n9493) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n4926), .CLK(n5529), 
        .Q(WX8521), .QN(n9492) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n4925), .CLK(n5530), 
        .Q(WX8523), .QN(n9491) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n4925), .CLK(n5530), 
        .Q(WX8525), .QN(n9490) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n4924), .CLK(n5530), 
        .Q(WX8527), .QN(n9489) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n4923), .CLK(n5531), 
        .Q(WX8529), .QN(n9488) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n4923), .CLK(n5531), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n4922), .CLK(n5531), 
        .Q(WX8533), .QN(n9522) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n4921), .CLK(n5532), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n4921), .CLK(n5532), 
        .Q(test_so72), .QN(n9517) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n4920), .CLK(n5532), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n4919), .CLK(n5533), 
        .Q(WX8541), .QN(n4075) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n4919), .CLK(n5533), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n4918), .CLK(n5533), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n4918), .CLK(n5533), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n4917), .CLK(n5534), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n4916), .CLK(n5534), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n4915), .CLK(n5535), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n4915), .CLK(n5535), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n4914), .CLK(n5535), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n4914), .CLK(n5535), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n4913), .CLK(n5536), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n4913), .CLK(n5536), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n4913), .CLK(n5536), 
        .Q(WX8565), .QN(n4231) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n4912), .CLK(n5536), 
        .Q(WX8567), .QN(n9501) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n4912), .CLK(n5536), 
        .Q(WX8569), .QN(n4228) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n4912), .CLK(n5536), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n4929), .CLK(n5528), 
        .Q(WX8573), .QN(n4225) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n4929), .CLK(n5528), 
        .Q(WX8575), .QN(n4223) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n4928), .CLK(n5528), 
        .Q(WX8577), .QN(n4221) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n4928), .CLK(n5528), 
        .Q(WX8579), .QN(n4219) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n4927), .CLK(n5529), 
        .Q(WX8581), .QN(n4217) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n4926), .CLK(n5529), 
        .Q(WX8583), .QN(n4215) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n4926), .CLK(n5529), 
        .Q(WX8585), .QN(n4213) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n4925), .CLK(n5530), 
        .Q(WX8587), .QN(n4211) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n4924), .CLK(n5530), 
        .Q(WX8589), .QN(n4209) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n4924), .CLK(n5530), 
        .Q(WX8591), .QN(n4207) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n4923), .CLK(n5531), 
        .Q(WX8593), .QN(n4205) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n4922), .CLK(n5531), 
        .Q(WX8595), .QN(n4469) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n4922), .CLK(n5531), 
        .Q(WX8597), .QN(n4470) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n4921), .CLK(n5532), 
        .Q(WX8599), .QN(n4471) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n4921), .CLK(n5532), 
        .Q(WX8601), .QN(n4472) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n4920), .CLK(n5532), 
        .Q(WX8603), .QN(n4473) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n4919), .CLK(n5533), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n4919), .CLK(n5533), 
        .Q(WX8607), .QN(n4474) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n4918), .CLK(n5533), 
        .Q(WX8609), .QN(n4475) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n4917), .CLK(n5534), 
        .Q(WX8611), .QN(n4476) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n4917), .CLK(n5534), 
        .Q(WX8613), .QN(n4477) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n4916), .CLK(n5534), 
        .Q(WX8615), .QN(n4478) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n4915), .CLK(n5535), 
        .Q(WX8617), .QN(n4479) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n4915), .CLK(n5535), 
        .Q(WX8619), .QN(n4480) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n4914), .CLK(n5535), 
        .Q(WX8621), .QN(n4481) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n4913), .CLK(n5536), 
        .Q(WX8623), .QN(n4482) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n4913), .CLK(n5536), 
        .Q(WX8625), .QN(n4394) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n4913), .CLK(n5536), 
        .Q(WX8627), .QN(n4483) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n4912), .CLK(n5536), 
        .Q(WX8629), .QN(n4484) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n4912), .CLK(n5536), 
        .Q(WX8631), .QN(n4485) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n4912), .CLK(n5536), 
        .Q(WX8633), .QN(n4486) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n4911), .CLK(n5537), 
        .Q(WX8635), .QN(n4395) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n4911), .CLK(n5537), 
        .Q(WX8637), .QN(n4487) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n4911), .CLK(n5537), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n4928), .CLK(n5528), 
        .Q(WX8641), .QN(n4488) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n4928), .CLK(n5528), 
        .Q(WX8643), .QN(n4489) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n4927), .CLK(n5529), 
        .Q(WX8645), .QN(n4490) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n4926), .CLK(n5529), 
        .Q(WX8647), .QN(n4491) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n4926), .CLK(n5529), 
        .Q(WX8649), .QN(n4396) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n4925), .CLK(n5530), 
        .Q(WX8651), .QN(n4492) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n4924), .CLK(n5530), 
        .Q(WX8653), .QN(n4493) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n4924), .CLK(n5530), 
        .Q(WX8655), .QN(n4494) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n4923), .CLK(n5531), 
        .Q(WX8657), .QN(n4411) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n4843), .CLK(n5571), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n4843), .CLK(n5571), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n4843), .CLK(n5571), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n4843), .CLK(n5571), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n4843), .CLK(n5571), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n4843), .CLK(n5571), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n4842), .CLK(n5571), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n4842), .CLK(n5571), .Q(test_so76), .QN(n4694) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n4842), .CLK(n5571), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n4842), .CLK(n5571), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n4842), .CLK(n5571), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n4911), .CLK(
        n5537), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n4911), .CLK(
        n5537), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n4911), .CLK(
        n5537), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n4910), .CLK(
        n5537), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n4909), .CLK(
        n5538), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n4909), .CLK(
        n5538), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n4909), .CLK(
        n5538), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n4909), .CLK(
        n5538), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n4909), .CLK(
        n5538), .Q(test_so77), .QN(n4695) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n4909), .CLK(n5538), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n4908), .CLK(
        n5538), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n383), .SI(CRC_OUT_3_31), .SE(n4907), .CLK(n5539), 
        .Q(WX9536), .QN(n4381) );
  SDFFX1 DFF_1345_Q_reg ( .D(n384), .SI(WX9536), .SE(n4902), .CLK(n5541), .Q(
        n8353) );
  SDFFX1 DFF_1346_Q_reg ( .D(n385), .SI(n8353), .SE(n4902), .CLK(n5541), .Q(
        n8352) );
  SDFFX1 DFF_1347_Q_reg ( .D(n386), .SI(n8352), .SE(n4903), .CLK(n5541), .Q(
        n8351) );
  SDFFX1 DFF_1348_Q_reg ( .D(n387), .SI(n8351), .SE(n4903), .CLK(n5541), .Q(
        n8350) );
  SDFFX1 DFF_1349_Q_reg ( .D(n388), .SI(n8350), .SE(n4903), .CLK(n5541), .Q(
        n8349) );
  SDFFX1 DFF_1350_Q_reg ( .D(n389), .SI(n8349), .SE(n4903), .CLK(n5541), .Q(
        n8348) );
  SDFFX1 DFF_1351_Q_reg ( .D(n390), .SI(n8348), .SE(n4903), .CLK(n5541), .Q(
        n8347) );
  SDFFX1 DFF_1352_Q_reg ( .D(n391), .SI(n8347), .SE(n4903), .CLK(n5541), .Q(
        n8346) );
  SDFFX1 DFF_1353_Q_reg ( .D(n392), .SI(n8346), .SE(n4904), .CLK(n5540), .Q(
        test_so78) );
  SDFFX1 DFF_1354_Q_reg ( .D(n393), .SI(test_si79), .SE(n4904), .CLK(n5540), 
        .Q(n8343) );
  SDFFX1 DFF_1355_Q_reg ( .D(n394), .SI(n8343), .SE(n4904), .CLK(n5540), .Q(
        n8342) );
  SDFFX1 DFF_1356_Q_reg ( .D(n395), .SI(n8342), .SE(n4904), .CLK(n5540), .Q(
        n8341) );
  SDFFX1 DFF_1357_Q_reg ( .D(n396), .SI(n8341), .SE(n4904), .CLK(n5540), .Q(
        n8340) );
  SDFFX1 DFF_1358_Q_reg ( .D(n397), .SI(n8340), .SE(n4904), .CLK(n5540), .Q(
        n8339) );
  SDFFX1 DFF_1359_Q_reg ( .D(n398), .SI(n8339), .SE(n4905), .CLK(n5540), .Q(
        n8338) );
  SDFFX1 DFF_1360_Q_reg ( .D(n399), .SI(n8338), .SE(n4905), .CLK(n5540), .Q(
        n8337) );
  SDFFX1 DFF_1361_Q_reg ( .D(n400), .SI(n8337), .SE(n4905), .CLK(n5540), .Q(
        n8336) );
  SDFFX1 DFF_1362_Q_reg ( .D(n401), .SI(n8336), .SE(n4905), .CLK(n5540), .Q(
        n8335) );
  SDFFX1 DFF_1363_Q_reg ( .D(n402), .SI(n8335), .SE(n4905), .CLK(n5540), .Q(
        n8334) );
  SDFFX1 DFF_1364_Q_reg ( .D(n403), .SI(n8334), .SE(n4905), .CLK(n5540), .Q(
        n8333) );
  SDFFX1 DFF_1365_Q_reg ( .D(n404), .SI(n8333), .SE(n4906), .CLK(n5539), .Q(
        n8332) );
  SDFFX1 DFF_1366_Q_reg ( .D(n405), .SI(n8332), .SE(n4906), .CLK(n5539), .Q(
        n8331) );
  SDFFX1 DFF_1367_Q_reg ( .D(n406), .SI(n8331), .SE(n4906), .CLK(n5539), .Q(
        n8330) );
  SDFFX1 DFF_1368_Q_reg ( .D(n407), .SI(n8330), .SE(n4906), .CLK(n5539), .Q(
        n8329) );
  SDFFX1 DFF_1369_Q_reg ( .D(n408), .SI(n8329), .SE(n4906), .CLK(n5539), .Q(
        n8328) );
  SDFFX1 DFF_1370_Q_reg ( .D(n409), .SI(n8328), .SE(n4906), .CLK(n5539), .Q(
        test_so79) );
  SDFFX1 DFF_1371_Q_reg ( .D(n410), .SI(test_si80), .SE(n4907), .CLK(n5539), 
        .Q(n8325) );
  SDFFX1 DFF_1372_Q_reg ( .D(n411), .SI(n8325), .SE(n4907), .CLK(n5539), .Q(
        n8324) );
  SDFFX1 DFF_1373_Q_reg ( .D(n412), .SI(n8324), .SE(n4907), .CLK(n5539), .Q(
        n8323) );
  SDFFX1 DFF_1374_Q_reg ( .D(n413), .SI(n8323), .SE(n4907), .CLK(n5539), .Q(
        n8322) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n4907), .CLK(n5539), .Q(
        n8321) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n4902), .CLK(n5541), .Q(
        n8320), .QN(n9487) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n4902), .CLK(n5541), .Q(
        n8319), .QN(n9486) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n4901), .CLK(n5542), .Q(
        n8318), .QN(n9485) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n4901), .CLK(n5542), .Q(
        n8317), .QN(n9484) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n4901), .CLK(n5542), .Q(
        n8316), .QN(n9483) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n4900), .CLK(n5542), .Q(
        n8315), .QN(n9482) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n4900), .CLK(n5542), .Q(
        n8314), .QN(n9481) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n4900), .CLK(n5542), .Q(
        n8313), .QN(n9480) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n4899), .CLK(n5543), .Q(
        n8312), .QN(n9479) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n4899), .CLK(n5543), .Q(
        n8311), .QN(n9478) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n4899), .CLK(n5543), .Q(
        n8310), .QN(n9477) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n4844), .CLK(n5570), .Q(
        test_so80), .QN(n4706) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n4898), .CLK(n5543), 
        .Q(n8307), .QN(n9476) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n4898), .CLK(n5543), .Q(
        n8306), .QN(n9473) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n4844), .CLK(n5570), .Q(
        n8305), .QN(n9472) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n4897), .CLK(n5544), .Q(
        n8304), .QN(n9469) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n4896), .CLK(n5544), .Q(
        WX9728) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n4896), .CLK(n5544), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n4896), .CLK(n5544), 
        .Q(WX9732) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n4895), .CLK(n5545), 
        .Q(WX9734) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n4894), .CLK(n5545), 
        .Q(WX9736) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n4894), .CLK(n5545), 
        .Q(WX9738) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n4893), .CLK(n5546), 
        .Q(WX9740) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n4892), .CLK(n5546), 
        .Q(WX9742) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n4892), .CLK(n5546), 
        .Q(WX9744) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n4891), .CLK(n5547), 
        .Q(WX9746) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n4890), .CLK(n5547), 
        .Q(WX9748) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n4890), .CLK(n5547), 
        .Q(WX9750) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n4889), .CLK(n5548), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n4888), .CLK(n5548), 
        .Q(WX9754) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n4888), .CLK(n5548), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n4887), .CLK(n5549), 
        .Q(WX9758) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n4902), .CLK(n5541), 
        .Q(WX9760) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n4902), .CLK(n5541), 
        .Q(WX9762), .QN(n4064) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n4901), .CLK(n5542), 
        .Q(WX9764), .QN(n4063) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n4901), .CLK(n5542), 
        .Q(WX9766), .QN(n4062) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n4901), .CLK(n5542), 
        .Q(WX9768), .QN(n4061) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n4900), .CLK(n5542), 
        .Q(WX9770), .QN(n4060) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n4900), .CLK(n5542), 
        .Q(WX9772), .QN(n4059) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n4900), .CLK(n5542), 
        .Q(WX9774), .QN(n4058) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n4899), .CLK(n5543), 
        .Q(WX9776), .QN(n4057) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n4899), .CLK(n5543), 
        .Q(WX9778), .QN(n4056) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n4899), .CLK(n5543), 
        .Q(WX9780), .QN(n4055) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n4898), .CLK(n5543), 
        .Q(WX9782) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n4898), .CLK(n5543), 
        .Q(WX9784), .QN(n4053) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n4898), .CLK(n5543), 
        .Q(test_so82), .QN(n9474) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n4844), .CLK(n5570), 
        .Q(WX9788), .QN(n4052) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n4897), .CLK(n5544), 
        .Q(WX9790), .QN(n9471) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n4897), .CLK(n5544), 
        .Q(WX9792), .QN(n9468) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n4896), .CLK(n5544), 
        .Q(WX9794), .QN(n9467) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n4896), .CLK(n5544), 
        .Q(WX9796), .QN(n9466) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n4895), .CLK(n5545), 
        .Q(WX9798), .QN(n9465) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n4894), .CLK(n5545), 
        .Q(WX9800), .QN(n9464) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n4894), .CLK(n5545), 
        .Q(WX9802), .QN(n9463) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n4893), .CLK(n5546), 
        .Q(WX9804), .QN(n9462) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n4892), .CLK(n5546), 
        .Q(WX9806), .QN(n9461) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n4892), .CLK(n5546), 
        .Q(WX9808), .QN(n9460) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n4891), .CLK(n5547), 
        .Q(WX9810), .QN(n9459) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n4890), .CLK(n5547), 
        .Q(WX9812), .QN(n9458) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n4890), .CLK(n5547), 
        .Q(WX9814), .QN(n9457) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n4889), .CLK(n5548), 
        .Q(WX9816), .QN(n9456) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n4888), .CLK(n5548), 
        .Q(WX9818), .QN(n9455) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n4888), .CLK(n5548), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n4887), .CLK(n5549), 
        .Q(WX9822), .QN(n9453) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n4886), .CLK(n5549), 
        .Q(WX9824), .QN(n4032) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n4886), .CLK(n5549), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n4886), .CLK(n5549), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n4885), .CLK(n5550), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n4885), .CLK(n5550), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n4885), .CLK(n5550), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n4884), .CLK(n5550), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n4884), .CLK(n5550), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n4884), .CLK(n5550), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n4883), .CLK(n5551), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n4883), .CLK(n5551), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n4883), .CLK(n5551), 
        .Q(WX9846), .QN(n4054) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n4882), .CLK(n5551), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n4898), .CLK(n5543), 
        .Q(WX9850), .QN(n9475) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n4897), .CLK(n5544), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n4897), .CLK(n5544), 
        .Q(test_so84), .QN(n9470) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n4897), .CLK(n5544), 
        .Q(WX9856), .QN(n4203) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n4896), .CLK(n5544), 
        .Q(WX9858), .QN(n4201) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n4895), .CLK(n5545), 
        .Q(WX9860), .QN(n4199) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n4895), .CLK(n5545), 
        .Q(WX9862), .QN(n4197) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n4894), .CLK(n5545), 
        .Q(WX9864), .QN(n4195) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n4893), .CLK(n5546), 
        .Q(WX9866), .QN(n4193) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n4893), .CLK(n5546), 
        .Q(WX9868), .QN(n4191) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n4892), .CLK(n5546), 
        .Q(WX9870), .QN(n4189) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n4891), .CLK(n5547), 
        .Q(WX9872), .QN(n4187) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n4891), .CLK(n5547), 
        .Q(WX9874), .QN(n4185) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n4890), .CLK(n5547), 
        .Q(WX9876), .QN(n4183) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n4889), .CLK(n5548), 
        .Q(WX9878), .QN(n4181) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n4889), .CLK(n5548), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n4888), .CLK(n5548), 
        .Q(WX9882), .QN(n4178) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n4887), .CLK(n5549), 
        .Q(WX9884), .QN(n9454) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n4887), .CLK(n5549), 
        .Q(WX9886), .QN(n4175) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n4886), .CLK(n5549), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n4886), .CLK(n5549), 
        .Q(WX9890), .QN(n4443) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n4886), .CLK(n5549), 
        .Q(WX9892), .QN(n4444) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n4885), .CLK(n5550), 
        .Q(WX9894), .QN(n4445) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n4885), .CLK(n5550), 
        .Q(WX9896), .QN(n4446) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n4885), .CLK(n5550), 
        .Q(WX9898), .QN(n4447) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n4884), .CLK(n5550), 
        .Q(WX9900), .QN(n4448) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n4884), .CLK(n5550), 
        .Q(WX9902), .QN(n4449) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n4884), .CLK(n5550), 
        .Q(WX9904), .QN(n4450) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n4883), .CLK(n5551), 
        .Q(WX9906), .QN(n4451) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n4883), .CLK(n5551), 
        .Q(WX9908), .QN(n4452) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n4883), .CLK(n5551), 
        .Q(WX9910), .QN(n4453) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n4882), .CLK(n5551), 
        .Q(WX9912), .QN(n4454) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n4882), .CLK(n5551), 
        .Q(WX9914), .QN(n4455) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n4882), .CLK(n5551), 
        .Q(WX9916), .QN(n4456) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n4882), .CLK(n5551), 
        .Q(WX9918), .QN(n4391) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n4882), .CLK(n5551), 
        .Q(WX9920), .QN(n4457) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n4881), .CLK(n5552), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n4895), .CLK(n5545), 
        .Q(WX9924), .QN(n4458) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n4895), .CLK(n5545), 
        .Q(WX9926), .QN(n4459) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n4894), .CLK(n5545), 
        .Q(WX9928), .QN(n4392) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n4893), .CLK(n5546), 
        .Q(WX9930), .QN(n4460) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n4893), .CLK(n5546), 
        .Q(WX9932), .QN(n4461) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n4892), .CLK(n5546), 
        .Q(WX9934), .QN(n4462) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n4891), .CLK(n5547), 
        .Q(WX9936), .QN(n4463) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n4891), .CLK(n5547), 
        .Q(WX9938), .QN(n4464) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n4890), .CLK(n5547), 
        .Q(WX9940), .QN(n4465) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n4889), .CLK(n5548), 
        .Q(WX9942), .QN(n4393) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n4889), .CLK(n5548), 
        .Q(WX9944), .QN(n4466) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n4888), .CLK(n5548), 
        .Q(WX9946), .QN(n4467) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n4887), .CLK(n5549), 
        .Q(WX9948), .QN(n4468) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n4887), .CLK(n5549), 
        .Q(WX9950), .QN(n4410) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n4847), .CLK(n5569), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n4847), .CLK(
        n5569), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n4847), .CLK(
        n5569), .Q(test_so87), .QN(n4713) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n4847), .CLK(n5569), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n4846), .CLK(
        n5569), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n4845), .CLK(
        n5570), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n4844), .CLK(
        n5570), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n4844), .CLK(
        n5570), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n4844), .CLK(
        n5570), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n4881), .CLK(
        n5552), .Q(test_so88), .QN(n4714) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n4881), .CLK(n5552), 
        .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n4881), .CLK(
        n5552), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n4881), .CLK(
        n5552), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n4881), .CLK(
        n5552), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n4880), .CLK(
        n5552), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n4879), .CLK(
        n5553), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n4879), .CLK(
        n5553), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n435), .SI(CRC_OUT_2_31), .SE(n4879), .CLK(n5553), 
        .Q(WX10829) );
  SDFFX1 DFF_1537_Q_reg ( .D(n437), .SI(WX10829), .SE(n4874), .CLK(n5555), .Q(
        n8295) );
  SDFFX1 DFF_1538_Q_reg ( .D(n439), .SI(n8295), .SE(n4874), .CLK(n5555), .Q(
        n8294) );
  SDFFX1 DFF_1539_Q_reg ( .D(n441), .SI(n8294), .SE(n4874), .CLK(n5555), .Q(
        n8293) );
  SDFFX1 DFF_1540_Q_reg ( .D(n443), .SI(n8293), .SE(n4874), .CLK(n5555), .Q(
        test_so89) );
  SDFFX1 DFF_1541_Q_reg ( .D(n445), .SI(test_si90), .SE(n4875), .CLK(n5555), 
        .Q(n8290) );
  SDFFX1 DFF_1542_Q_reg ( .D(n447), .SI(n8290), .SE(n4875), .CLK(n5555), .Q(
        n8289) );
  SDFFX1 DFF_1543_Q_reg ( .D(n449), .SI(n8289), .SE(n4875), .CLK(n5555), .Q(
        n8288) );
  SDFFX1 DFF_1544_Q_reg ( .D(n451), .SI(n8288), .SE(n4875), .CLK(n5555), .Q(
        n8287) );
  SDFFX1 DFF_1545_Q_reg ( .D(n453), .SI(n8287), .SE(n4875), .CLK(n5555), .Q(
        n8286) );
  SDFFX1 DFF_1546_Q_reg ( .D(n455), .SI(n8286), .SE(n4875), .CLK(n5555), .Q(
        n8285) );
  SDFFX1 DFF_1547_Q_reg ( .D(n457), .SI(n8285), .SE(n4876), .CLK(n5554), .Q(
        n8284) );
  SDFFX1 DFF_1548_Q_reg ( .D(n459), .SI(n8284), .SE(n4876), .CLK(n5554), .Q(
        n8283) );
  SDFFX1 DFF_1549_Q_reg ( .D(n461), .SI(n8283), .SE(n4876), .CLK(n5554), .Q(
        n8282) );
  SDFFX1 DFF_1550_Q_reg ( .D(n463), .SI(n8282), .SE(n4876), .CLK(n5554), .Q(
        n8281) );
  SDFFX1 DFF_1551_Q_reg ( .D(n465), .SI(n8281), .SE(n4876), .CLK(n5554), .Q(
        n8280) );
  SDFFX1 DFF_1552_Q_reg ( .D(n467), .SI(n8280), .SE(n4876), .CLK(n5554), .Q(
        n8279) );
  SDFFX1 DFF_1553_Q_reg ( .D(n469), .SI(n8279), .SE(n4877), .CLK(n5554), .Q(
        n8278) );
  SDFFX1 DFF_1554_Q_reg ( .D(n471), .SI(n8278), .SE(n4877), .CLK(n5554), .Q(
        n8277) );
  SDFFX1 DFF_1555_Q_reg ( .D(n473), .SI(n8277), .SE(n4877), .CLK(n5554), .Q(
        n8276) );
  SDFFX1 DFF_1556_Q_reg ( .D(n475), .SI(n8276), .SE(n4877), .CLK(n5554), .Q(
        n8275) );
  SDFFX1 DFF_1557_Q_reg ( .D(n477), .SI(n8275), .SE(n4877), .CLK(n5554), .Q(
        test_so90) );
  SDFFX1 DFF_1558_Q_reg ( .D(n479), .SI(test_si91), .SE(n4877), .CLK(n5554), 
        .Q(n8272) );
  SDFFX1 DFF_1559_Q_reg ( .D(n481), .SI(n8272), .SE(n4878), .CLK(n5553), .Q(
        n8271) );
  SDFFX1 DFF_1560_Q_reg ( .D(n483), .SI(n8271), .SE(n4878), .CLK(n5553), .Q(
        n8270) );
  SDFFX1 DFF_1561_Q_reg ( .D(n485), .SI(n8270), .SE(n4878), .CLK(n5553), .Q(
        n8269) );
  SDFFX1 DFF_1562_Q_reg ( .D(n487), .SI(n8269), .SE(n4878), .CLK(n5553), .Q(
        n8268) );
  SDFFX1 DFF_1563_Q_reg ( .D(n489), .SI(n8268), .SE(n4878), .CLK(n5553), .Q(
        n8267) );
  SDFFX1 DFF_1564_Q_reg ( .D(n491), .SI(n8267), .SE(n4878), .CLK(n5553), .Q(
        n8266) );
  SDFFX1 DFF_1565_Q_reg ( .D(n493), .SI(n8266), .SE(n4879), .CLK(n5553), .Q(
        n8265) );
  SDFFX1 DFF_1566_Q_reg ( .D(n495), .SI(n8265), .SE(n4879), .CLK(n5553), .Q(
        n8264) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n4879), .CLK(n5553), 
        .Q(n8263) );
  SDFFX1 DFF_1568_Q_reg ( .D(n432), .SI(n8263), .SE(n4874), .CLK(n5555), .Q(
        n8262), .QN(n9729) );
  SDFFX1 DFF_1569_Q_reg ( .D(n434), .SI(n8262), .SE(n4873), .CLK(n5556), .Q(
        n8261), .QN(n9728) );
  SDFFX1 DFF_1570_Q_reg ( .D(n436), .SI(n8261), .SE(n4873), .CLK(n5556), .Q(
        n8260), .QN(n9727) );
  SDFFX1 DFF_1571_Q_reg ( .D(n438), .SI(n8260), .SE(n4873), .CLK(n5556), .Q(
        n8259), .QN(n9726) );
  SDFFX1 DFF_1572_Q_reg ( .D(n440), .SI(n8259), .SE(n4872), .CLK(n5556), .Q(
        n8258), .QN(n9725) );
  SDFFX1 DFF_1573_Q_reg ( .D(n442), .SI(n8258), .SE(n4872), .CLK(n5556), .Q(
        n8257), .QN(n9724) );
  SDFFX1 DFF_1574_Q_reg ( .D(n444), .SI(n8257), .SE(n4872), .CLK(n5556), .Q(
        test_so91), .QN(n4712) );
  SDFFX1 DFF_1575_Q_reg ( .D(n446), .SI(test_si92), .SE(n4871), .CLK(n5557), 
        .Q(n8254), .QN(n9723) );
  SDFFX1 DFF_1576_Q_reg ( .D(n448), .SI(n8254), .SE(n4871), .CLK(n5557), .Q(
        n8253), .QN(n9720) );
  SDFFX1 DFF_1577_Q_reg ( .D(n450), .SI(n8253), .SE(n4848), .CLK(n5568), .Q(
        n8252), .QN(n9719) );
  SDFFX1 DFF_1578_Q_reg ( .D(n452), .SI(n8252), .SE(n4870), .CLK(n5557), .Q(
        n8251), .QN(n9716) );
  SDFFX1 DFF_1579_Q_reg ( .D(n454), .SI(n8251), .SE(n4870), .CLK(n5557), .Q(
        n8250), .QN(n9715) );
  SDFFX1 DFF_1580_Q_reg ( .D(n456), .SI(n8250), .SE(n4869), .CLK(n5558), .Q(
        n8249), .QN(n9714) );
  SDFFX1 DFF_1581_Q_reg ( .D(n458), .SI(n8249), .SE(n4868), .CLK(n5558), .Q(
        n8248), .QN(n9713) );
  SDFFX1 DFF_1582_Q_reg ( .D(n460), .SI(n8248), .SE(n4868), .CLK(n5558), .Q(
        n8247), .QN(n9712) );
  SDFFX1 DFF_1583_Q_reg ( .D(n462), .SI(n8247), .SE(n4867), .CLK(n5559), .Q(
        n8246), .QN(n9711) );
  SDFFX1 DFF_1584_Q_reg ( .D(n464), .SI(n8246), .SE(n4867), .CLK(n5559), .Q(
        WX11021) );
  SDFFX1 DFF_1585_Q_reg ( .D(n466), .SI(WX11021), .SE(n4866), .CLK(n5559), .Q(
        WX11023) );
  SDFFX1 DFF_1586_Q_reg ( .D(n468), .SI(WX11023), .SE(n4866), .CLK(n5559), .Q(
        WX11025) );
  SDFFX1 DFF_1587_Q_reg ( .D(n470), .SI(WX11025), .SE(n4865), .CLK(n5560), .Q(
        WX11027) );
  SDFFX1 DFF_1588_Q_reg ( .D(n472), .SI(WX11027), .SE(n4864), .CLK(n5560), .Q(
        WX11029) );
  SDFFX1 DFF_1589_Q_reg ( .D(n474), .SI(WX11029), .SE(n4864), .CLK(n5560), .Q(
        WX11031) );
  SDFFX1 DFF_1590_Q_reg ( .D(n476), .SI(WX11031), .SE(n4863), .CLK(n5561), .Q(
        WX11033) );
  SDFFX1 DFF_1591_Q_reg ( .D(n478), .SI(WX11033), .SE(n4862), .CLK(n5561), .Q(
        test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(n480), .SI(test_si93), .SE(n4861), .CLK(n5562), 
        .Q(WX11037) );
  SDFFX1 DFF_1593_Q_reg ( .D(n482), .SI(WX11037), .SE(n4861), .CLK(n5562), .Q(
        WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(n484), .SI(WX11039), .SE(n4860), .CLK(n5562), .Q(
        WX11041) );
  SDFFX1 DFF_1595_Q_reg ( .D(n486), .SI(WX11041), .SE(n4860), .CLK(n5562), .Q(
        WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(n488), .SI(WX11043), .SE(n4859), .CLK(n5563), .Q(
        WX11045) );
  SDFFX1 DFF_1597_Q_reg ( .D(n490), .SI(WX11045), .SE(n4858), .CLK(n5563), .Q(
        WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(n492), .SI(WX11047), .SE(n4858), .CLK(n5563), .Q(
        WX11049) );
  SDFFX1 DFF_1599_Q_reg ( .D(n494), .SI(WX11049), .SE(n4857), .CLK(n5564), .Q(
        WX11051) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n4874), .CLK(n5555), 
        .Q(WX11053), .QN(n4031) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n4873), .CLK(n5556), 
        .Q(WX11055), .QN(n4051) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n4873), .CLK(n5556), 
        .Q(WX11057), .QN(n4050) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n4873), .CLK(n5556), 
        .Q(WX11059), .QN(n4049) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n4872), .CLK(n5556), 
        .Q(WX11061), .QN(n4048) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n4872), .CLK(n5556), 
        .Q(WX11063), .QN(n4047) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n4872), .CLK(n5556), 
        .Q(WX11065) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n4871), .CLK(n5557), 
        .Q(WX11067), .QN(n4045) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n4871), .CLK(n5557), 
        .Q(test_so93), .QN(n9721) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n4847), .CLK(n5569), 
        .Q(WX11071), .QN(n4044) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n4870), .CLK(n5557), 
        .Q(WX11073), .QN(n9718) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n4870), .CLK(n5557), 
        .Q(WX11075), .QN(n4043) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n4869), .CLK(n5558), 
        .Q(WX11077) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n4869), .CLK(n5558), 
        .Q(WX11079), .QN(n4041) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n4868), .CLK(n5558), 
        .Q(WX11081), .QN(n4040) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n4868), .CLK(n5558), 
        .Q(WX11083), .QN(n4039) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n4867), .CLK(n5559), 
        .Q(WX11085), .QN(n9710) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n4866), .CLK(n5559), 
        .Q(WX11087), .QN(n9709) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n4865), .CLK(n5560), 
        .Q(WX11089), .QN(n9708) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n4865), .CLK(n5560), 
        .Q(WX11091), .QN(n9707) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n4864), .CLK(n5560), 
        .Q(WX11093), .QN(n9706) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n4863), .CLK(n5561), 
        .Q(WX11095), .QN(n9705) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n4863), .CLK(n5561), 
        .Q(WX11097), .QN(n9704) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n4862), .CLK(n5561), 
        .Q(WX11099), .QN(n9703) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n4862), .CLK(n5561), 
        .Q(WX11101), .QN(n9702) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n4861), .CLK(n5562), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n4860), .CLK(n5562), 
        .Q(WX11105), .QN(n9700) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n4859), .CLK(n5563), 
        .Q(WX11107), .QN(n9699) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n4859), .CLK(n5563), 
        .Q(WX11109), .QN(n9698) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n4858), .CLK(n5563), 
        .Q(WX11111), .QN(n9697) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n4857), .CLK(n5564), 
        .Q(WX11113), .QN(n9696) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n4857), .CLK(n5564), 
        .Q(WX11115), .QN(n9695) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n4856), .CLK(n5564), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n4856), .CLK(n5564), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n4856), .CLK(n5564), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n4855), .CLK(n5565), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n4855), .CLK(n5565), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n4855), .CLK(n5565), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n4854), .CLK(n5565), 
        .Q(WX11129), .QN(n4046) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n4854), .CLK(n5565), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n4871), .CLK(n5557), 
        .Q(WX11133), .QN(n9722) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n4871), .CLK(n5557), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n4870), .CLK(n5557), 
        .Q(test_so95), .QN(n9717) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n4870), .CLK(n5557), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n4869), .CLK(n5558), 
        .Q(WX11141), .QN(n4042) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n4869), .CLK(n5558), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n4868), .CLK(n5558), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n4867), .CLK(n5559), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n4867), .CLK(n5559), 
        .Q(WX11149), .QN(n4173) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n4866), .CLK(n5559), 
        .Q(WX11151), .QN(n4171) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n4865), .CLK(n5560), 
        .Q(WX11153), .QN(n4169) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n4865), .CLK(n5560), 
        .Q(WX11155), .QN(n4167) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n4864), .CLK(n5560), 
        .Q(WX11157), .QN(n4165) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n4863), .CLK(n5561), 
        .Q(WX11159), .QN(n4163) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n4863), .CLK(n5561), 
        .Q(WX11161), .QN(n4161) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n4862), .CLK(n5561), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n4861), .CLK(n5562), 
        .Q(WX11165), .QN(n4158) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n4861), .CLK(n5562), 
        .Q(WX11167), .QN(n9701) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n4860), .CLK(n5562), 
        .Q(WX11169), .QN(n4155) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n4859), .CLK(n5563), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n4859), .CLK(n5563), 
        .Q(WX11173), .QN(n4152) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n4858), .CLK(n5563), 
        .Q(WX11175), .QN(n4150) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n4857), .CLK(n5564), 
        .Q(WX11177), .QN(n4148) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n4857), .CLK(n5564), 
        .Q(WX11179), .QN(n4146) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n4856), .CLK(n5564), 
        .Q(WX11181), .QN(n4417) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n4856), .CLK(n5564), 
        .Q(WX11183), .QN(n4418) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n4855), .CLK(n5565), 
        .Q(WX11185), .QN(n4419) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n4855), .CLK(n5565), 
        .Q(WX11187), .QN(n4420) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n4855), .CLK(n5565), 
        .Q(WX11189), .QN(n4421) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n4854), .CLK(n5565), 
        .Q(WX11191), .QN(n4422) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n4854), .CLK(n5565), 
        .Q(WX11193), .QN(n4423) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n4854), .CLK(n5565), 
        .Q(WX11195), .QN(n4424) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n4854), .CLK(n5565), 
        .Q(WX11197), .QN(n4425) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n4853), .CLK(n5566), 
        .Q(WX11199), .QN(n4426) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n4853), .CLK(n5566), 
        .Q(WX11201), .QN(n4427) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n4853), .CLK(n5566), 
        .Q(WX11203), .QN(n4428) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n4853), .CLK(n5566), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n4869), .CLK(n5558), 
        .Q(WX11207), .QN(n4429) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n4868), .CLK(n5558), 
        .Q(WX11209), .QN(n4430) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n4867), .CLK(n5559), 
        .Q(WX11211), .QN(n4388) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n4866), .CLK(n5559), 
        .Q(WX11213), .QN(n4431) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n4866), .CLK(n5559), 
        .Q(WX11215), .QN(n4432) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n4865), .CLK(n5560), 
        .Q(WX11217), .QN(n4433) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n4864), .CLK(n5560), 
        .Q(WX11219), .QN(n4434) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n4864), .CLK(n5560), 
        .Q(WX11221), .QN(n4389) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n4863), .CLK(n5561), 
        .Q(WX11223), .QN(n4435) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n4862), .CLK(n5561), 
        .Q(WX11225), .QN(n4436) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n4862), .CLK(n5561), 
        .Q(WX11227), .QN(n4437) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n4861), .CLK(n5562), 
        .Q(WX11229), .QN(n4438) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n4860), .CLK(n5562), 
        .Q(WX11231), .QN(n4439) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n4860), .CLK(n5562), 
        .Q(WX11233), .QN(n4440) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n4859), .CLK(n5563), 
        .Q(WX11235), .QN(n4390) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n4858), .CLK(n5563), 
        .Q(WX11237), .QN(n4441) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n4858), .CLK(n5563), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n4857), .CLK(n5564), 
        .Q(WX11241), .QN(n4442) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n4856), .CLK(n5564), 
        .Q(WX11243), .QN(n4409) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n4851), .CLK(n5567), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n4851), .CLK(
        n5567), .Q(CRC_OUT_1_1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n4851), .CLK(
        n5567), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n4851), .CLK(
        n5567), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n4851), .CLK(
        n5567), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n4851), .CLK(
        n5567), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n4850), .CLK(
        n5567), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n4849), .CLK(
        n5568), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n4849), .CLK(
        n5568), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n4849), .CLK(
        n5568), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n4849), .CLK(n5568), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n4849), .CLK(
        n5568), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n4849), .CLK(
        n5568), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n4848), .CLK(
        n5568), .Q(CRC_OUT_1_18) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n4848), .CLK(
        n5568), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n4848), .CLK(
        n5568), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n4848), .CLK(
        n5568), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n4848), .CLK(
        n5568), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n4847), .CLK(
        n5569), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n4853), .CLK(
        n5566), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n4853), .CLK(
        n5566), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n4852), .CLK(
        n5566), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n4852), .CLK(
        n5566), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n4852), .CLK(
        n5566), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n4852), .CLK(
        n5566), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n4852), .CLK(
        n5566), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n4852), .CLK(
        n5566), .Q(test_so100) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n151), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n163), .IN2(n155), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n469), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  INVX0 TrojanINVtest_se ( .INP(n5231), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  NBUFFX2 U4685 ( .INP(n5614), .Z(n5445) );
  NBUFFX2 U4686 ( .INP(n5614), .Z(n5443) );
  NBUFFX2 U4687 ( .INP(n5614), .Z(n5444) );
  NBUFFX2 U4688 ( .INP(n5614), .Z(n5442) );
  NBUFFX2 U4689 ( .INP(n5589), .Z(n5567) );
  NBUFFX2 U4690 ( .INP(n5589), .Z(n5566) );
  NBUFFX2 U4691 ( .INP(n5590), .Z(n5565) );
  NBUFFX2 U4692 ( .INP(n5590), .Z(n5564) );
  NBUFFX2 U4693 ( .INP(n5590), .Z(n5563) );
  NBUFFX2 U4694 ( .INP(n5590), .Z(n5562) );
  NBUFFX2 U4695 ( .INP(n5590), .Z(n5561) );
  NBUFFX2 U4696 ( .INP(n5591), .Z(n5560) );
  NBUFFX2 U4697 ( .INP(n5591), .Z(n5559) );
  NBUFFX2 U4698 ( .INP(n5591), .Z(n5558) );
  NBUFFX2 U4699 ( .INP(n5589), .Z(n5568) );
  NBUFFX2 U4700 ( .INP(n5591), .Z(n5557) );
  NBUFFX2 U4701 ( .INP(n5591), .Z(n5556) );
  NBUFFX2 U4702 ( .INP(n5592), .Z(n5554) );
  NBUFFX2 U4703 ( .INP(n5592), .Z(n5555) );
  NBUFFX2 U4704 ( .INP(n5592), .Z(n5553) );
  NBUFFX2 U4705 ( .INP(n5589), .Z(n5569) );
  NBUFFX2 U4706 ( .INP(n5592), .Z(n5552) );
  NBUFFX2 U4707 ( .INP(n5592), .Z(n5551) );
  NBUFFX2 U4708 ( .INP(n5593), .Z(n5550) );
  NBUFFX2 U4709 ( .INP(n5593), .Z(n5549) );
  NBUFFX2 U4710 ( .INP(n5593), .Z(n5548) );
  NBUFFX2 U4711 ( .INP(n5593), .Z(n5547) );
  NBUFFX2 U4712 ( .INP(n5593), .Z(n5546) );
  NBUFFX2 U4713 ( .INP(n5594), .Z(n5545) );
  NBUFFX2 U4714 ( .INP(n5594), .Z(n5544) );
  NBUFFX2 U4715 ( .INP(n5589), .Z(n5570) );
  NBUFFX2 U4716 ( .INP(n5594), .Z(n5543) );
  NBUFFX2 U4717 ( .INP(n5594), .Z(n5542) );
  NBUFFX2 U4718 ( .INP(n5595), .Z(n5540) );
  NBUFFX2 U4719 ( .INP(n5594), .Z(n5541) );
  NBUFFX2 U4720 ( .INP(n5595), .Z(n5539) );
  NBUFFX2 U4721 ( .INP(n5595), .Z(n5538) );
  NBUFFX2 U4722 ( .INP(n5595), .Z(n5537) );
  NBUFFX2 U4723 ( .INP(n5595), .Z(n5536) );
  NBUFFX2 U4724 ( .INP(n5597), .Z(n5530) );
  NBUFFX2 U4725 ( .INP(n5597), .Z(n5529) );
  NBUFFX2 U4726 ( .INP(n5597), .Z(n5528) );
  NBUFFX2 U4727 ( .INP(n5597), .Z(n5527) );
  NBUFFX2 U4728 ( .INP(n5596), .Z(n5535) );
  NBUFFX2 U4729 ( .INP(n5596), .Z(n5534) );
  NBUFFX2 U4730 ( .INP(n5596), .Z(n5533) );
  NBUFFX2 U4731 ( .INP(n5596), .Z(n5532) );
  NBUFFX2 U4732 ( .INP(n5588), .Z(n5571) );
  NBUFFX2 U4733 ( .INP(n5596), .Z(n5531) );
  NBUFFX2 U4734 ( .INP(n5597), .Z(n5526) );
  NBUFFX2 U4735 ( .INP(n5598), .Z(n5525) );
  NBUFFX2 U4736 ( .INP(n5598), .Z(n5524) );
  NBUFFX2 U4737 ( .INP(n5588), .Z(n5573) );
  NBUFFX2 U4738 ( .INP(n5588), .Z(n5572) );
  NBUFFX2 U4739 ( .INP(n5598), .Z(n5523) );
  NBUFFX2 U4740 ( .INP(n5598), .Z(n5522) );
  NBUFFX2 U4741 ( .INP(n5598), .Z(n5521) );
  NBUFFX2 U4742 ( .INP(n5599), .Z(n5520) );
  NBUFFX2 U4743 ( .INP(n5599), .Z(n5519) );
  NBUFFX2 U4744 ( .INP(n5599), .Z(n5518) );
  NBUFFX2 U4745 ( .INP(n5599), .Z(n5517) );
  NBUFFX2 U4746 ( .INP(n5599), .Z(n5516) );
  NBUFFX2 U4747 ( .INP(n5600), .Z(n5515) );
  NBUFFX2 U4748 ( .INP(n5600), .Z(n5514) );
  NBUFFX2 U4749 ( .INP(n5600), .Z(n5512) );
  NBUFFX2 U4750 ( .INP(n5600), .Z(n5513) );
  NBUFFX2 U4751 ( .INP(n5600), .Z(n5511) );
  NBUFFX2 U4752 ( .INP(n5588), .Z(n5575) );
  NBUFFX2 U4753 ( .INP(n5588), .Z(n5574) );
  NBUFFX2 U4754 ( .INP(n5601), .Z(n5510) );
  NBUFFX2 U4755 ( .INP(n5601), .Z(n5509) );
  NBUFFX2 U4756 ( .INP(n5601), .Z(n5508) );
  NBUFFX2 U4757 ( .INP(n5601), .Z(n5507) );
  NBUFFX2 U4758 ( .INP(n5601), .Z(n5506) );
  NBUFFX2 U4759 ( .INP(n5602), .Z(n5505) );
  NBUFFX2 U4760 ( .INP(n5602), .Z(n5504) );
  NBUFFX2 U4761 ( .INP(n5602), .Z(n5503) );
  NBUFFX2 U4762 ( .INP(n5602), .Z(n5502) );
  NBUFFX2 U4763 ( .INP(n5602), .Z(n5501) );
  NBUFFX2 U4764 ( .INP(n5603), .Z(n5500) );
  NBUFFX2 U4765 ( .INP(n5603), .Z(n5498) );
  NBUFFX2 U4766 ( .INP(n5603), .Z(n5499) );
  NBUFFX2 U4767 ( .INP(n5603), .Z(n5497) );
  NBUFFX2 U4768 ( .INP(n5603), .Z(n5496) );
  NBUFFX2 U4769 ( .INP(n5587), .Z(n5576) );
  NBUFFX2 U4770 ( .INP(n5604), .Z(n5495) );
  NBUFFX2 U4771 ( .INP(n5605), .Z(n5489) );
  NBUFFX2 U4772 ( .INP(n5605), .Z(n5488) );
  NBUFFX2 U4773 ( .INP(n5605), .Z(n5487) );
  NBUFFX2 U4774 ( .INP(n5605), .Z(n5486) );
  NBUFFX2 U4775 ( .INP(n5606), .Z(n5485) );
  NBUFFX2 U4776 ( .INP(n5604), .Z(n5494) );
  NBUFFX2 U4777 ( .INP(n5604), .Z(n5493) );
  NBUFFX2 U4778 ( .INP(n5604), .Z(n5492) );
  NBUFFX2 U4779 ( .INP(n5604), .Z(n5491) );
  NBUFFX2 U4780 ( .INP(n5605), .Z(n5490) );
  NBUFFX2 U4781 ( .INP(n5607), .Z(n5480) );
  NBUFFX2 U4782 ( .INP(n5606), .Z(n5481) );
  NBUFFX2 U4783 ( .INP(n5606), .Z(n5483) );
  NBUFFX2 U4784 ( .INP(n5606), .Z(n5482) );
  NBUFFX2 U4785 ( .INP(n5607), .Z(n5479) );
  NBUFFX2 U4786 ( .INP(n5607), .Z(n5478) );
  NBUFFX2 U4787 ( .INP(n5607), .Z(n5477) );
  NBUFFX2 U4788 ( .INP(n5607), .Z(n5476) );
  NBUFFX2 U4789 ( .INP(n5608), .Z(n5475) );
  NBUFFX2 U4790 ( .INP(n5608), .Z(n5474) );
  NBUFFX2 U4791 ( .INP(n5608), .Z(n5473) );
  NBUFFX2 U4792 ( .INP(n5606), .Z(n5484) );
  NBUFFX2 U4793 ( .INP(n5608), .Z(n5472) );
  NBUFFX2 U4794 ( .INP(n5608), .Z(n5471) );
  NBUFFX2 U4795 ( .INP(n5609), .Z(n5470) );
  NBUFFX2 U4796 ( .INP(n5609), .Z(n5469) );
  NBUFFX2 U4797 ( .INP(n5609), .Z(n5466) );
  NBUFFX2 U4798 ( .INP(n5609), .Z(n5467) );
  NBUFFX2 U4799 ( .INP(n5609), .Z(n5468) );
  NBUFFX2 U4800 ( .INP(n5587), .Z(n5579) );
  NBUFFX2 U4801 ( .INP(n5587), .Z(n5578) );
  NBUFFX2 U4802 ( .INP(n5587), .Z(n5577) );
  NBUFFX2 U4803 ( .INP(n5586), .Z(n5583) );
  NBUFFX2 U4804 ( .INP(n5586), .Z(n5582) );
  NBUFFX2 U4805 ( .INP(n5586), .Z(n5581) );
  NBUFFX2 U4806 ( .INP(n5610), .Z(n5465) );
  NBUFFX2 U4807 ( .INP(n5610), .Z(n5464) );
  NBUFFX2 U4808 ( .INP(n5610), .Z(n5463) );
  NBUFFX2 U4809 ( .INP(n5610), .Z(n5462) );
  NBUFFX2 U4810 ( .INP(n5610), .Z(n5461) );
  NBUFFX2 U4811 ( .INP(n5611), .Z(n5460) );
  NBUFFX2 U4812 ( .INP(n5587), .Z(n5580) );
  NBUFFX2 U4813 ( .INP(n5611), .Z(n5459) );
  NBUFFX2 U4814 ( .INP(n5611), .Z(n5457) );
  NBUFFX2 U4815 ( .INP(n5611), .Z(n5458) );
  NBUFFX2 U4816 ( .INP(n5611), .Z(n5456) );
  NBUFFX2 U4817 ( .INP(n5586), .Z(n5584) );
  NBUFFX2 U4818 ( .INP(n5612), .Z(n5455) );
  NBUFFX2 U4819 ( .INP(n5612), .Z(n5454) );
  NBUFFX2 U4820 ( .INP(n5612), .Z(n5453) );
  NBUFFX2 U4821 ( .INP(n5612), .Z(n5452) );
  NBUFFX2 U4822 ( .INP(n5612), .Z(n5451) );
  NBUFFX2 U4823 ( .INP(n5613), .Z(n5450) );
  NBUFFX2 U4824 ( .INP(n5586), .Z(n5585) );
  NBUFFX2 U4825 ( .INP(n5613), .Z(n5449) );
  NBUFFX2 U4826 ( .INP(n5613), .Z(n5448) );
  NBUFFX2 U4827 ( .INP(n5613), .Z(n5447) );
  NBUFFX2 U4828 ( .INP(n5613), .Z(n5446) );
  NBUFFX2 U4829 ( .INP(n4769), .Z(n4786) );
  NBUFFX2 U4830 ( .INP(n4769), .Z(n4785) );
  NBUFFX2 U4831 ( .INP(n4769), .Z(n4787) );
  NBUFFX2 U4832 ( .INP(n4746), .Z(n4765) );
  NBUFFX2 U4833 ( .INP(n4746), .Z(n4764) );
  NBUFFX2 U4834 ( .INP(n4768), .Z(n4784) );
  NBUFFX2 U4835 ( .INP(n4744), .Z(n4755) );
  NBUFFX2 U4836 ( .INP(n4744), .Z(n4754) );
  NBUFFX2 U4837 ( .INP(n4766), .Z(n4771) );
  NBUFFX2 U4838 ( .INP(n4744), .Z(n4753) );
  NBUFFX2 U4839 ( .INP(n4766), .Z(n4772) );
  NBUFFX2 U4840 ( .INP(n4744), .Z(n4752) );
  NBUFFX2 U4841 ( .INP(n4766), .Z(n4773) );
  NBUFFX2 U4842 ( .INP(n4766), .Z(n4774) );
  NBUFFX2 U4843 ( .INP(n4743), .Z(n4750) );
  NBUFFX2 U4844 ( .INP(n4743), .Z(n4749) );
  NBUFFX2 U4845 ( .INP(n4767), .Z(n4775) );
  NBUFFX2 U4846 ( .INP(n4743), .Z(n4751) );
  NBUFFX2 U4847 ( .INP(n4767), .Z(n4777) );
  NBUFFX2 U4848 ( .INP(n4746), .Z(n4763) );
  NBUFFX2 U4849 ( .INP(n4746), .Z(n4762) );
  NBUFFX2 U4850 ( .INP(n4745), .Z(n4761) );
  NBUFFX2 U4851 ( .INP(n4745), .Z(n4759) );
  NBUFFX2 U4852 ( .INP(n4745), .Z(n4758) );
  NBUFFX2 U4853 ( .INP(n4768), .Z(n4783) );
  NBUFFX2 U4854 ( .INP(n4768), .Z(n4782) );
  NBUFFX2 U4855 ( .INP(n4768), .Z(n4781) );
  NBUFFX2 U4856 ( .INP(n4745), .Z(n4757) );
  NBUFFX2 U4857 ( .INP(n4768), .Z(n4780) );
  NBUFFX2 U4858 ( .INP(n4767), .Z(n4779) );
  NBUFFX2 U4859 ( .INP(n4744), .Z(n4756) );
  NBUFFX2 U4860 ( .INP(n4745), .Z(n4760) );
  NBUFFX2 U4861 ( .INP(n4743), .Z(n4747) );
  NBUFFX2 U4862 ( .INP(n4766), .Z(n4770) );
  NBUFFX2 U4863 ( .INP(n4767), .Z(n4778) );
  NBUFFX2 U4864 ( .INP(n4743), .Z(n4748) );
  NBUFFX2 U4865 ( .INP(n4767), .Z(n4776) );
  NBUFFX2 U4866 ( .INP(n4769), .Z(n4788) );
  NBUFFX2 U4867 ( .INP(n5332), .Z(n5288) );
  NBUFFX2 U4868 ( .INP(n5332), .Z(n5287) );
  NBUFFX2 U4869 ( .INP(n5332), .Z(n5286) );
  NBUFFX2 U4870 ( .INP(n5332), .Z(n5285) );
  NBUFFX2 U4871 ( .INP(n5333), .Z(n5284) );
  NBUFFX2 U4872 ( .INP(n5332), .Z(n5289) );
  NBUFFX2 U4873 ( .INP(n5326), .Z(n5319) );
  NBUFFX2 U4874 ( .INP(n5326), .Z(n5318) );
  NBUFFX2 U4875 ( .INP(n5326), .Z(n5317) );
  NBUFFX2 U4876 ( .INP(n5326), .Z(n5316) );
  NBUFFX2 U4877 ( .INP(n5326), .Z(n5315) );
  NBUFFX2 U4878 ( .INP(n5327), .Z(n5314) );
  NBUFFX2 U4879 ( .INP(n5327), .Z(n5313) );
  NBUFFX2 U4880 ( .INP(n5327), .Z(n5312) );
  NBUFFX2 U4881 ( .INP(n5327), .Z(n5311) );
  NBUFFX2 U4882 ( .INP(n5327), .Z(n5310) );
  NBUFFX2 U4883 ( .INP(n5328), .Z(n5308) );
  NBUFFX2 U4884 ( .INP(n5328), .Z(n5307) );
  NBUFFX2 U4885 ( .INP(n5328), .Z(n5306) );
  NBUFFX2 U4886 ( .INP(n5328), .Z(n5305) );
  NBUFFX2 U4887 ( .INP(n5329), .Z(n5304) );
  NBUFFX2 U4888 ( .INP(n5329), .Z(n5303) );
  NBUFFX2 U4889 ( .INP(n5329), .Z(n5302) );
  NBUFFX2 U4890 ( .INP(n5329), .Z(n5301) );
  NBUFFX2 U4891 ( .INP(n5329), .Z(n5300) );
  NBUFFX2 U4892 ( .INP(n5330), .Z(n5299) );
  NBUFFX2 U4893 ( .INP(n5330), .Z(n5298) );
  NBUFFX2 U4894 ( .INP(n5330), .Z(n5297) );
  NBUFFX2 U4895 ( .INP(n5330), .Z(n5296) );
  NBUFFX2 U4896 ( .INP(n5328), .Z(n5309) );
  NBUFFX2 U4897 ( .INP(n5330), .Z(n5295) );
  NBUFFX2 U4898 ( .INP(n5331), .Z(n5294) );
  NBUFFX2 U4899 ( .INP(n5331), .Z(n5293) );
  NBUFFX2 U4900 ( .INP(n5331), .Z(n5292) );
  NBUFFX2 U4901 ( .INP(n5331), .Z(n5291) );
  NBUFFX2 U4902 ( .INP(n5331), .Z(n5290) );
  NBUFFX2 U4903 ( .INP(n5337), .Z(n5263) );
  NBUFFX2 U4904 ( .INP(n5337), .Z(n5264) );
  NBUFFX2 U4905 ( .INP(n5335), .Z(n5271) );
  NBUFFX2 U4906 ( .INP(n5333), .Z(n5281) );
  NBUFFX2 U4907 ( .INP(n5334), .Z(n5278) );
  NBUFFX2 U4908 ( .INP(n5334), .Z(n5277) );
  NBUFFX2 U4909 ( .INP(n5334), .Z(n5276) );
  NBUFFX2 U4910 ( .INP(n5336), .Z(n5267) );
  NBUFFX2 U4911 ( .INP(n5336), .Z(n5265) );
  NBUFFX2 U4912 ( .INP(n5336), .Z(n5266) );
  NBUFFX2 U4913 ( .INP(n5334), .Z(n5279) );
  NBUFFX2 U4914 ( .INP(n5333), .Z(n5280) );
  NBUFFX2 U4915 ( .INP(n5336), .Z(n5268) );
  NBUFFX2 U4916 ( .INP(n5336), .Z(n5269) );
  NBUFFX2 U4917 ( .INP(n5333), .Z(n5282) );
  NBUFFX2 U4918 ( .INP(n5334), .Z(n5275) );
  NBUFFX2 U4919 ( .INP(n5335), .Z(n5270) );
  NBUFFX2 U4920 ( .INP(n5335), .Z(n5274) );
  NBUFFX2 U4921 ( .INP(n5335), .Z(n5272) );
  NBUFFX2 U4922 ( .INP(n5335), .Z(n5273) );
  NBUFFX2 U4923 ( .INP(n5333), .Z(n5283) );
  NBUFFX2 U4924 ( .INP(n5262), .Z(n5248) );
  NBUFFX2 U4925 ( .INP(n5262), .Z(n5249) );
  NBUFFX2 U4926 ( .INP(n5262), .Z(n5247) );
  NBUFFX2 U4927 ( .INP(n5261), .Z(n5250) );
  NBUFFX2 U4928 ( .INP(n5261), .Z(n5251) );
  NBUFFX2 U4929 ( .INP(n5261), .Z(n5252) );
  NBUFFX2 U4930 ( .INP(n5261), .Z(n5253) );
  NBUFFX2 U4931 ( .INP(n5261), .Z(n5254) );
  NBUFFX2 U4932 ( .INP(n5260), .Z(n5255) );
  NBUFFX2 U4933 ( .INP(n5260), .Z(n5256) );
  NBUFFX2 U4934 ( .INP(n5260), .Z(n5258) );
  NBUFFX2 U4935 ( .INP(n5260), .Z(n5257) );
  INVX0 U4936 ( .INP(n6016), .ZN(n4742) );
  INVX0 U4937 ( .INP(n6023), .ZN(n4813) );
  NBUFFX2 U4938 ( .INP(n5325), .Z(n5321) );
  NBUFFX2 U4939 ( .INP(n5325), .Z(n5320) );
  NBUFFX2 U4940 ( .INP(n5325), .Z(n5322) );
  NBUFFX2 U4941 ( .INP(n5325), .Z(n5323) );
  NBUFFX2 U4942 ( .INP(n5325), .Z(n5324) );
  NBUFFX2 U4943 ( .INP(n5260), .Z(n5259) );
  INVX0 U4944 ( .INP(n4735), .ZN(n4715) );
  INVX0 U4945 ( .INP(n4735), .ZN(n4716) );
  INVX0 U4946 ( .INP(n4735), .ZN(n4717) );
  INVX0 U4947 ( .INP(n4734), .ZN(n4718) );
  INVX0 U4948 ( .INP(n4734), .ZN(n4719) );
  INVX0 U4949 ( .INP(n4734), .ZN(n4720) );
  INVX0 U4950 ( .INP(n4734), .ZN(n4721) );
  INVX0 U4951 ( .INP(n4734), .ZN(n4722) );
  INVX0 U4952 ( .INP(n4734), .ZN(n4723) );
  INVX0 U4953 ( .INP(n4734), .ZN(n4724) );
  INVX0 U4954 ( .INP(n4733), .ZN(n4725) );
  INVX0 U4955 ( .INP(n4733), .ZN(n4726) );
  INVX0 U4956 ( .INP(n4733), .ZN(n4727) );
  INVX0 U4957 ( .INP(n4733), .ZN(n4728) );
  INVX0 U4958 ( .INP(n4733), .ZN(n4729) );
  INVX0 U4959 ( .INP(n4733), .ZN(n4730) );
  INVX0 U4960 ( .INP(n4733), .ZN(n4731) );
  INVX0 U4961 ( .INP(n4733), .ZN(n4732) );
  NBUFFX2 U4962 ( .INP(n4741), .Z(n4733) );
  NBUFFX2 U4963 ( .INP(n4741), .Z(n4734) );
  NBUFFX2 U4964 ( .INP(n4739), .Z(n4735) );
  NBUFFX2 U4965 ( .INP(n4742), .Z(n4736) );
  NBUFFX2 U4966 ( .INP(n4742), .Z(n4737) );
  NBUFFX2 U4967 ( .INP(n4742), .Z(n4738) );
  NBUFFX2 U4968 ( .INP(n4742), .Z(n4739) );
  NBUFFX2 U4969 ( .INP(n4741), .Z(n4740) );
  NBUFFX2 U4970 ( .INP(n4742), .Z(n4741) );
  NBUFFX2 U4971 ( .INP(n6017), .Z(n4743) );
  NBUFFX2 U4972 ( .INP(n6017), .Z(n4744) );
  NBUFFX2 U4973 ( .INP(n6017), .Z(n4745) );
  NBUFFX2 U4974 ( .INP(n6017), .Z(n4746) );
  NBUFFX2 U4975 ( .INP(n6021), .Z(n4766) );
  NBUFFX2 U4976 ( .INP(n6021), .Z(n4767) );
  NBUFFX2 U4977 ( .INP(n6021), .Z(n4768) );
  NBUFFX2 U4978 ( .INP(n6021), .Z(n4769) );
  INVX0 U4979 ( .INP(n4807), .ZN(n4789) );
  INVX0 U4980 ( .INP(n4806), .ZN(n4790) );
  INVX0 U4981 ( .INP(n4807), .ZN(n4791) );
  INVX0 U4982 ( .INP(n4806), .ZN(n4792) );
  INVX0 U4983 ( .INP(n4806), .ZN(n4793) );
  INVX0 U4984 ( .INP(n4806), .ZN(n4794) );
  INVX0 U4985 ( .INP(n4806), .ZN(n4795) );
  INVX0 U4986 ( .INP(n4806), .ZN(n4796) );
  INVX0 U4987 ( .INP(n4806), .ZN(n4797) );
  INVX0 U4988 ( .INP(n4805), .ZN(n4798) );
  INVX0 U4989 ( .INP(n4806), .ZN(n4799) );
  INVX0 U4990 ( .INP(n4805), .ZN(n4800) );
  INVX0 U4991 ( .INP(n4805), .ZN(n4801) );
  INVX0 U4992 ( .INP(n4805), .ZN(n4802) );
  INVX0 U4993 ( .INP(n4805), .ZN(n4803) );
  INVX0 U4994 ( .INP(n4805), .ZN(n4804) );
  NBUFFX2 U4995 ( .INP(n4813), .Z(n4805) );
  NBUFFX2 U4996 ( .INP(n4813), .Z(n4806) );
  NBUFFX2 U4997 ( .INP(n4813), .Z(n4807) );
  NBUFFX2 U4998 ( .INP(n4813), .Z(n4808) );
  NBUFFX2 U4999 ( .INP(n4813), .Z(n4809) );
  NBUFFX2 U5000 ( .INP(n4807), .Z(n4810) );
  NBUFFX2 U5001 ( .INP(n4806), .Z(n4811) );
  NBUFFX2 U5002 ( .INP(n4808), .Z(n4812) );
  NBUFFX2 U5003 ( .INP(n5198), .Z(n4814) );
  NBUFFX2 U5004 ( .INP(n5197), .Z(n4815) );
  NBUFFX2 U5005 ( .INP(n5197), .Z(n4816) );
  NBUFFX2 U5006 ( .INP(n5197), .Z(n4817) );
  NBUFFX2 U5007 ( .INP(n5196), .Z(n4818) );
  NBUFFX2 U5008 ( .INP(n5196), .Z(n4819) );
  NBUFFX2 U5009 ( .INP(n5196), .Z(n4820) );
  NBUFFX2 U5010 ( .INP(n5195), .Z(n4821) );
  NBUFFX2 U5011 ( .INP(n5195), .Z(n4822) );
  NBUFFX2 U5012 ( .INP(n5195), .Z(n4823) );
  NBUFFX2 U5013 ( .INP(n5194), .Z(n4824) );
  NBUFFX2 U5014 ( .INP(n5194), .Z(n4825) );
  NBUFFX2 U5015 ( .INP(n5194), .Z(n4826) );
  NBUFFX2 U5016 ( .INP(n5193), .Z(n4827) );
  NBUFFX2 U5017 ( .INP(n5193), .Z(n4828) );
  NBUFFX2 U5018 ( .INP(n5193), .Z(n4829) );
  NBUFFX2 U5019 ( .INP(n5192), .Z(n4830) );
  NBUFFX2 U5020 ( .INP(n5192), .Z(n4831) );
  NBUFFX2 U5021 ( .INP(n5192), .Z(n4832) );
  NBUFFX2 U5022 ( .INP(n5191), .Z(n4833) );
  NBUFFX2 U5023 ( .INP(n5191), .Z(n4834) );
  NBUFFX2 U5024 ( .INP(n5191), .Z(n4835) );
  NBUFFX2 U5025 ( .INP(n5190), .Z(n4836) );
  NBUFFX2 U5026 ( .INP(n5190), .Z(n4837) );
  NBUFFX2 U5027 ( .INP(n5190), .Z(n4838) );
  NBUFFX2 U5028 ( .INP(n5189), .Z(n4839) );
  NBUFFX2 U5029 ( .INP(n5189), .Z(n4840) );
  NBUFFX2 U5030 ( .INP(n5189), .Z(n4841) );
  NBUFFX2 U5031 ( .INP(n5188), .Z(n4842) );
  NBUFFX2 U5032 ( .INP(n5188), .Z(n4843) );
  NBUFFX2 U5033 ( .INP(n5188), .Z(n4844) );
  NBUFFX2 U5034 ( .INP(n5187), .Z(n4845) );
  NBUFFX2 U5035 ( .INP(n5187), .Z(n4846) );
  NBUFFX2 U5036 ( .INP(n5187), .Z(n4847) );
  NBUFFX2 U5037 ( .INP(n5186), .Z(n4848) );
  NBUFFX2 U5038 ( .INP(n5186), .Z(n4849) );
  NBUFFX2 U5039 ( .INP(n5186), .Z(n4850) );
  NBUFFX2 U5040 ( .INP(n5185), .Z(n4851) );
  NBUFFX2 U5041 ( .INP(n5185), .Z(n4852) );
  NBUFFX2 U5042 ( .INP(n5185), .Z(n4853) );
  NBUFFX2 U5043 ( .INP(n5184), .Z(n4854) );
  NBUFFX2 U5044 ( .INP(n5184), .Z(n4855) );
  NBUFFX2 U5045 ( .INP(n5184), .Z(n4856) );
  NBUFFX2 U5046 ( .INP(n5183), .Z(n4857) );
  NBUFFX2 U5047 ( .INP(n5183), .Z(n4858) );
  NBUFFX2 U5048 ( .INP(n5183), .Z(n4859) );
  NBUFFX2 U5049 ( .INP(n5182), .Z(n4860) );
  NBUFFX2 U5050 ( .INP(n5182), .Z(n4861) );
  NBUFFX2 U5051 ( .INP(n5182), .Z(n4862) );
  NBUFFX2 U5052 ( .INP(n5181), .Z(n4863) );
  NBUFFX2 U5053 ( .INP(n5181), .Z(n4864) );
  NBUFFX2 U5054 ( .INP(n5181), .Z(n4865) );
  NBUFFX2 U5055 ( .INP(n5180), .Z(n4866) );
  NBUFFX2 U5056 ( .INP(n5180), .Z(n4867) );
  NBUFFX2 U5057 ( .INP(n5180), .Z(n4868) );
  NBUFFX2 U5058 ( .INP(n5179), .Z(n4869) );
  NBUFFX2 U5059 ( .INP(n5179), .Z(n4870) );
  NBUFFX2 U5060 ( .INP(n5179), .Z(n4871) );
  NBUFFX2 U5061 ( .INP(n5178), .Z(n4872) );
  NBUFFX2 U5062 ( .INP(n5178), .Z(n4873) );
  NBUFFX2 U5063 ( .INP(n5178), .Z(n4874) );
  NBUFFX2 U5064 ( .INP(n5177), .Z(n4875) );
  NBUFFX2 U5065 ( .INP(n5177), .Z(n4876) );
  NBUFFX2 U5066 ( .INP(n5177), .Z(n4877) );
  NBUFFX2 U5067 ( .INP(n5176), .Z(n4878) );
  NBUFFX2 U5068 ( .INP(n5176), .Z(n4879) );
  NBUFFX2 U5069 ( .INP(n5176), .Z(n4880) );
  NBUFFX2 U5070 ( .INP(n5175), .Z(n4881) );
  NBUFFX2 U5071 ( .INP(n5175), .Z(n4882) );
  NBUFFX2 U5072 ( .INP(n5175), .Z(n4883) );
  NBUFFX2 U5073 ( .INP(n5174), .Z(n4884) );
  NBUFFX2 U5074 ( .INP(n5174), .Z(n4885) );
  NBUFFX2 U5075 ( .INP(n5174), .Z(n4886) );
  NBUFFX2 U5076 ( .INP(n5173), .Z(n4887) );
  NBUFFX2 U5077 ( .INP(n5173), .Z(n4888) );
  NBUFFX2 U5078 ( .INP(n5173), .Z(n4889) );
  NBUFFX2 U5079 ( .INP(n5172), .Z(n4890) );
  NBUFFX2 U5080 ( .INP(n5172), .Z(n4891) );
  NBUFFX2 U5081 ( .INP(n5172), .Z(n4892) );
  NBUFFX2 U5082 ( .INP(n5171), .Z(n4893) );
  NBUFFX2 U5083 ( .INP(n5171), .Z(n4894) );
  NBUFFX2 U5084 ( .INP(n5171), .Z(n4895) );
  NBUFFX2 U5085 ( .INP(n5170), .Z(n4896) );
  NBUFFX2 U5086 ( .INP(n5170), .Z(n4897) );
  NBUFFX2 U5087 ( .INP(n5170), .Z(n4898) );
  NBUFFX2 U5088 ( .INP(n5169), .Z(n4899) );
  NBUFFX2 U5089 ( .INP(n5169), .Z(n4900) );
  NBUFFX2 U5090 ( .INP(n5169), .Z(n4901) );
  NBUFFX2 U5091 ( .INP(n5168), .Z(n4902) );
  NBUFFX2 U5092 ( .INP(n5168), .Z(n4903) );
  NBUFFX2 U5093 ( .INP(n5168), .Z(n4904) );
  NBUFFX2 U5094 ( .INP(n5167), .Z(n4905) );
  NBUFFX2 U5095 ( .INP(n5167), .Z(n4906) );
  NBUFFX2 U5096 ( .INP(n5167), .Z(n4907) );
  NBUFFX2 U5097 ( .INP(n5166), .Z(n4908) );
  NBUFFX2 U5098 ( .INP(n5166), .Z(n4909) );
  NBUFFX2 U5099 ( .INP(n5166), .Z(n4910) );
  NBUFFX2 U5100 ( .INP(n5165), .Z(n4911) );
  NBUFFX2 U5101 ( .INP(n5165), .Z(n4912) );
  NBUFFX2 U5102 ( .INP(n5165), .Z(n4913) );
  NBUFFX2 U5103 ( .INP(n5164), .Z(n4914) );
  NBUFFX2 U5104 ( .INP(n5164), .Z(n4915) );
  NBUFFX2 U5105 ( .INP(n5164), .Z(n4916) );
  NBUFFX2 U5106 ( .INP(n5163), .Z(n4917) );
  NBUFFX2 U5107 ( .INP(n5163), .Z(n4918) );
  NBUFFX2 U5108 ( .INP(n5163), .Z(n4919) );
  NBUFFX2 U5109 ( .INP(n5162), .Z(n4920) );
  NBUFFX2 U5110 ( .INP(n5162), .Z(n4921) );
  NBUFFX2 U5111 ( .INP(n5162), .Z(n4922) );
  NBUFFX2 U5112 ( .INP(n5161), .Z(n4923) );
  NBUFFX2 U5113 ( .INP(n5161), .Z(n4924) );
  NBUFFX2 U5114 ( .INP(n5161), .Z(n4925) );
  NBUFFX2 U5115 ( .INP(n5160), .Z(n4926) );
  NBUFFX2 U5116 ( .INP(n5160), .Z(n4927) );
  NBUFFX2 U5117 ( .INP(n5160), .Z(n4928) );
  NBUFFX2 U5118 ( .INP(n5159), .Z(n4929) );
  NBUFFX2 U5119 ( .INP(n5159), .Z(n4930) );
  NBUFFX2 U5120 ( .INP(n5159), .Z(n4931) );
  NBUFFX2 U5121 ( .INP(n5158), .Z(n4932) );
  NBUFFX2 U5122 ( .INP(n5158), .Z(n4933) );
  NBUFFX2 U5123 ( .INP(n5158), .Z(n4934) );
  NBUFFX2 U5124 ( .INP(n5157), .Z(n4935) );
  NBUFFX2 U5125 ( .INP(n5157), .Z(n4936) );
  NBUFFX2 U5126 ( .INP(n5157), .Z(n4937) );
  NBUFFX2 U5127 ( .INP(n5156), .Z(n4938) );
  NBUFFX2 U5128 ( .INP(n5156), .Z(n4939) );
  NBUFFX2 U5129 ( .INP(n5156), .Z(n4940) );
  NBUFFX2 U5130 ( .INP(n5155), .Z(n4941) );
  NBUFFX2 U5131 ( .INP(n5155), .Z(n4942) );
  NBUFFX2 U5132 ( .INP(n5155), .Z(n4943) );
  NBUFFX2 U5133 ( .INP(n5154), .Z(n4944) );
  NBUFFX2 U5134 ( .INP(n5154), .Z(n4945) );
  NBUFFX2 U5135 ( .INP(n5154), .Z(n4946) );
  NBUFFX2 U5136 ( .INP(n5153), .Z(n4947) );
  NBUFFX2 U5137 ( .INP(n5153), .Z(n4948) );
  NBUFFX2 U5138 ( .INP(n5153), .Z(n4949) );
  NBUFFX2 U5139 ( .INP(n5152), .Z(n4950) );
  NBUFFX2 U5140 ( .INP(n5152), .Z(n4951) );
  NBUFFX2 U5141 ( .INP(n5152), .Z(n4952) );
  NBUFFX2 U5142 ( .INP(n5151), .Z(n4953) );
  NBUFFX2 U5143 ( .INP(n5151), .Z(n4954) );
  NBUFFX2 U5144 ( .INP(n5151), .Z(n4955) );
  NBUFFX2 U5145 ( .INP(n5150), .Z(n4956) );
  NBUFFX2 U5146 ( .INP(n5150), .Z(n4957) );
  NBUFFX2 U5147 ( .INP(n5150), .Z(n4958) );
  NBUFFX2 U5148 ( .INP(n5149), .Z(n4959) );
  NBUFFX2 U5149 ( .INP(n5149), .Z(n4960) );
  NBUFFX2 U5150 ( .INP(n5149), .Z(n4961) );
  NBUFFX2 U5151 ( .INP(n5148), .Z(n4962) );
  NBUFFX2 U5152 ( .INP(n5148), .Z(n4963) );
  NBUFFX2 U5153 ( .INP(n5148), .Z(n4964) );
  NBUFFX2 U5154 ( .INP(n5147), .Z(n4965) );
  NBUFFX2 U5155 ( .INP(n5147), .Z(n4966) );
  NBUFFX2 U5156 ( .INP(n5147), .Z(n4967) );
  NBUFFX2 U5157 ( .INP(n5146), .Z(n4968) );
  NBUFFX2 U5158 ( .INP(n5146), .Z(n4969) );
  NBUFFX2 U5159 ( .INP(n5146), .Z(n4970) );
  NBUFFX2 U5160 ( .INP(n5145), .Z(n4971) );
  NBUFFX2 U5161 ( .INP(n5145), .Z(n4972) );
  NBUFFX2 U5162 ( .INP(n5145), .Z(n4973) );
  NBUFFX2 U5163 ( .INP(n5144), .Z(n4974) );
  NBUFFX2 U5164 ( .INP(n5144), .Z(n4975) );
  NBUFFX2 U5165 ( .INP(n5144), .Z(n4976) );
  NBUFFX2 U5166 ( .INP(n5143), .Z(n4977) );
  NBUFFX2 U5167 ( .INP(n5143), .Z(n4978) );
  NBUFFX2 U5168 ( .INP(n5143), .Z(n4979) );
  NBUFFX2 U5169 ( .INP(n5142), .Z(n4980) );
  NBUFFX2 U5170 ( .INP(n5142), .Z(n4981) );
  NBUFFX2 U5171 ( .INP(n5142), .Z(n4982) );
  NBUFFX2 U5172 ( .INP(n5141), .Z(n4983) );
  NBUFFX2 U5173 ( .INP(n5141), .Z(n4984) );
  NBUFFX2 U5174 ( .INP(n5141), .Z(n4985) );
  NBUFFX2 U5175 ( .INP(n5140), .Z(n4986) );
  NBUFFX2 U5176 ( .INP(n5140), .Z(n4987) );
  NBUFFX2 U5177 ( .INP(n5140), .Z(n4988) );
  NBUFFX2 U5178 ( .INP(n5139), .Z(n4989) );
  NBUFFX2 U5179 ( .INP(n5139), .Z(n4990) );
  NBUFFX2 U5180 ( .INP(n5139), .Z(n4991) );
  NBUFFX2 U5181 ( .INP(n5138), .Z(n4992) );
  NBUFFX2 U5182 ( .INP(n5138), .Z(n4993) );
  NBUFFX2 U5183 ( .INP(n5138), .Z(n4994) );
  NBUFFX2 U5184 ( .INP(n5137), .Z(n4995) );
  NBUFFX2 U5185 ( .INP(n5137), .Z(n4996) );
  NBUFFX2 U5186 ( .INP(n5137), .Z(n4997) );
  NBUFFX2 U5187 ( .INP(n5136), .Z(n4998) );
  NBUFFX2 U5188 ( .INP(n5136), .Z(n4999) );
  NBUFFX2 U5189 ( .INP(n5136), .Z(n5000) );
  NBUFFX2 U5190 ( .INP(n5135), .Z(n5001) );
  NBUFFX2 U5191 ( .INP(n5135), .Z(n5002) );
  NBUFFX2 U5192 ( .INP(n5135), .Z(n5003) );
  NBUFFX2 U5193 ( .INP(n5134), .Z(n5004) );
  NBUFFX2 U5194 ( .INP(n5134), .Z(n5005) );
  NBUFFX2 U5195 ( .INP(n5134), .Z(n5006) );
  NBUFFX2 U5196 ( .INP(n5133), .Z(n5007) );
  NBUFFX2 U5197 ( .INP(n5133), .Z(n5008) );
  NBUFFX2 U5198 ( .INP(n5133), .Z(n5009) );
  NBUFFX2 U5199 ( .INP(n5132), .Z(n5010) );
  NBUFFX2 U5200 ( .INP(n5132), .Z(n5011) );
  NBUFFX2 U5201 ( .INP(n5132), .Z(n5012) );
  NBUFFX2 U5202 ( .INP(n5131), .Z(n5013) );
  NBUFFX2 U5203 ( .INP(n5131), .Z(n5014) );
  NBUFFX2 U5204 ( .INP(n5131), .Z(n5015) );
  NBUFFX2 U5205 ( .INP(n5130), .Z(n5016) );
  NBUFFX2 U5206 ( .INP(n5130), .Z(n5017) );
  NBUFFX2 U5207 ( .INP(n5130), .Z(n5018) );
  NBUFFX2 U5208 ( .INP(n5129), .Z(n5019) );
  NBUFFX2 U5209 ( .INP(n5129), .Z(n5020) );
  NBUFFX2 U5210 ( .INP(n5129), .Z(n5021) );
  NBUFFX2 U5211 ( .INP(n5128), .Z(n5022) );
  NBUFFX2 U5212 ( .INP(n5128), .Z(n5023) );
  NBUFFX2 U5213 ( .INP(n5128), .Z(n5024) );
  NBUFFX2 U5214 ( .INP(n5127), .Z(n5025) );
  NBUFFX2 U5215 ( .INP(n5127), .Z(n5026) );
  NBUFFX2 U5216 ( .INP(n5127), .Z(n5027) );
  NBUFFX2 U5217 ( .INP(n5126), .Z(n5028) );
  NBUFFX2 U5218 ( .INP(n5126), .Z(n5029) );
  NBUFFX2 U5219 ( .INP(n5126), .Z(n5030) );
  NBUFFX2 U5220 ( .INP(n5125), .Z(n5031) );
  NBUFFX2 U5221 ( .INP(n5125), .Z(n5032) );
  NBUFFX2 U5222 ( .INP(n5125), .Z(n5033) );
  NBUFFX2 U5223 ( .INP(n5124), .Z(n5034) );
  NBUFFX2 U5224 ( .INP(n5124), .Z(n5035) );
  NBUFFX2 U5225 ( .INP(n5124), .Z(n5036) );
  NBUFFX2 U5226 ( .INP(n5123), .Z(n5037) );
  NBUFFX2 U5227 ( .INP(n5123), .Z(n5038) );
  NBUFFX2 U5228 ( .INP(n5123), .Z(n5039) );
  NBUFFX2 U5229 ( .INP(n5122), .Z(n5040) );
  NBUFFX2 U5230 ( .INP(n5122), .Z(n5041) );
  NBUFFX2 U5231 ( .INP(n5122), .Z(n5042) );
  NBUFFX2 U5232 ( .INP(n5121), .Z(n5043) );
  NBUFFX2 U5233 ( .INP(n5121), .Z(n5044) );
  NBUFFX2 U5234 ( .INP(n5121), .Z(n5045) );
  NBUFFX2 U5235 ( .INP(n5120), .Z(n5046) );
  NBUFFX2 U5236 ( .INP(n5120), .Z(n5047) );
  NBUFFX2 U5237 ( .INP(n5120), .Z(n5048) );
  NBUFFX2 U5238 ( .INP(n5119), .Z(n5049) );
  NBUFFX2 U5239 ( .INP(n5119), .Z(n5050) );
  NBUFFX2 U5240 ( .INP(n5119), .Z(n5051) );
  NBUFFX2 U5241 ( .INP(n5118), .Z(n5052) );
  NBUFFX2 U5242 ( .INP(n5118), .Z(n5053) );
  NBUFFX2 U5243 ( .INP(n5118), .Z(n5054) );
  NBUFFX2 U5244 ( .INP(n5117), .Z(n5055) );
  NBUFFX2 U5245 ( .INP(n5117), .Z(n5056) );
  NBUFFX2 U5246 ( .INP(n5117), .Z(n5057) );
  NBUFFX2 U5247 ( .INP(n5116), .Z(n5058) );
  NBUFFX2 U5248 ( .INP(n5116), .Z(n5059) );
  NBUFFX2 U5249 ( .INP(n5116), .Z(n5060) );
  NBUFFX2 U5250 ( .INP(n5115), .Z(n5061) );
  NBUFFX2 U5251 ( .INP(n5115), .Z(n5062) );
  NBUFFX2 U5252 ( .INP(n5115), .Z(n5063) );
  NBUFFX2 U5253 ( .INP(n5114), .Z(n5064) );
  NBUFFX2 U5254 ( .INP(n5114), .Z(n5065) );
  NBUFFX2 U5255 ( .INP(n5114), .Z(n5066) );
  NBUFFX2 U5256 ( .INP(n5113), .Z(n5067) );
  NBUFFX2 U5257 ( .INP(n5113), .Z(n5068) );
  NBUFFX2 U5258 ( .INP(n5113), .Z(n5069) );
  NBUFFX2 U5259 ( .INP(n5112), .Z(n5070) );
  NBUFFX2 U5260 ( .INP(n5112), .Z(n5071) );
  NBUFFX2 U5261 ( .INP(n5112), .Z(n5072) );
  NBUFFX2 U5262 ( .INP(n5111), .Z(n5073) );
  NBUFFX2 U5263 ( .INP(n5111), .Z(n5074) );
  NBUFFX2 U5264 ( .INP(n5111), .Z(n5075) );
  NBUFFX2 U5265 ( .INP(n5110), .Z(n5076) );
  NBUFFX2 U5266 ( .INP(n5110), .Z(n5077) );
  NBUFFX2 U5267 ( .INP(n5110), .Z(n5078) );
  NBUFFX2 U5268 ( .INP(n5109), .Z(n5079) );
  NBUFFX2 U5269 ( .INP(n5109), .Z(n5080) );
  NBUFFX2 U5270 ( .INP(n5109), .Z(n5081) );
  NBUFFX2 U5271 ( .INP(n5108), .Z(n5082) );
  NBUFFX2 U5272 ( .INP(n5108), .Z(n5083) );
  NBUFFX2 U5273 ( .INP(n5108), .Z(n5084) );
  NBUFFX2 U5274 ( .INP(n5107), .Z(n5085) );
  NBUFFX2 U5275 ( .INP(n5107), .Z(n5086) );
  NBUFFX2 U5276 ( .INP(n5107), .Z(n5087) );
  NBUFFX2 U5277 ( .INP(n5106), .Z(n5088) );
  NBUFFX2 U5278 ( .INP(n5106), .Z(n5089) );
  NBUFFX2 U5279 ( .INP(n5106), .Z(n5090) );
  NBUFFX2 U5280 ( .INP(n5105), .Z(n5091) );
  NBUFFX2 U5281 ( .INP(n5105), .Z(n5092) );
  NBUFFX2 U5282 ( .INP(n5105), .Z(n5093) );
  NBUFFX2 U5283 ( .INP(n5104), .Z(n5094) );
  NBUFFX2 U5284 ( .INP(n5104), .Z(n5095) );
  NBUFFX2 U5285 ( .INP(n5104), .Z(n5096) );
  NBUFFX2 U5286 ( .INP(n5103), .Z(n5097) );
  NBUFFX2 U5287 ( .INP(n5103), .Z(n5098) );
  NBUFFX2 U5288 ( .INP(n5103), .Z(n5099) );
  NBUFFX2 U5289 ( .INP(n5102), .Z(n5100) );
  NBUFFX2 U5290 ( .INP(n5102), .Z(n5101) );
  NBUFFX2 U5291 ( .INP(n5231), .Z(n5102) );
  NBUFFX2 U5292 ( .INP(n5230), .Z(n5103) );
  NBUFFX2 U5293 ( .INP(n5230), .Z(n5104) );
  NBUFFX2 U5294 ( .INP(n5230), .Z(n5105) );
  NBUFFX2 U5295 ( .INP(n5229), .Z(n5106) );
  NBUFFX2 U5296 ( .INP(n5229), .Z(n5107) );
  NBUFFX2 U5297 ( .INP(n5229), .Z(n5108) );
  NBUFFX2 U5298 ( .INP(n5228), .Z(n5109) );
  NBUFFX2 U5299 ( .INP(n5228), .Z(n5110) );
  NBUFFX2 U5300 ( .INP(n5228), .Z(n5111) );
  NBUFFX2 U5301 ( .INP(n5227), .Z(n5112) );
  NBUFFX2 U5302 ( .INP(n5227), .Z(n5113) );
  NBUFFX2 U5303 ( .INP(n5227), .Z(n5114) );
  NBUFFX2 U5304 ( .INP(n5226), .Z(n5115) );
  NBUFFX2 U5305 ( .INP(n5226), .Z(n5116) );
  NBUFFX2 U5306 ( .INP(n5226), .Z(n5117) );
  NBUFFX2 U5307 ( .INP(n5225), .Z(n5118) );
  NBUFFX2 U5308 ( .INP(n5225), .Z(n5119) );
  NBUFFX2 U5309 ( .INP(n5225), .Z(n5120) );
  NBUFFX2 U5310 ( .INP(n5224), .Z(n5121) );
  NBUFFX2 U5311 ( .INP(n5224), .Z(n5122) );
  NBUFFX2 U5312 ( .INP(n5224), .Z(n5123) );
  NBUFFX2 U5313 ( .INP(n5223), .Z(n5124) );
  NBUFFX2 U5314 ( .INP(n5223), .Z(n5125) );
  NBUFFX2 U5315 ( .INP(n5223), .Z(n5126) );
  NBUFFX2 U5316 ( .INP(n5222), .Z(n5127) );
  NBUFFX2 U5317 ( .INP(n5222), .Z(n5128) );
  NBUFFX2 U5318 ( .INP(n5222), .Z(n5129) );
  NBUFFX2 U5319 ( .INP(n5221), .Z(n5130) );
  NBUFFX2 U5320 ( .INP(n5221), .Z(n5131) );
  NBUFFX2 U5321 ( .INP(n5221), .Z(n5132) );
  NBUFFX2 U5322 ( .INP(n5220), .Z(n5133) );
  NBUFFX2 U5323 ( .INP(n5220), .Z(n5134) );
  NBUFFX2 U5324 ( .INP(n5220), .Z(n5135) );
  NBUFFX2 U5325 ( .INP(n5219), .Z(n5136) );
  NBUFFX2 U5326 ( .INP(n5219), .Z(n5137) );
  NBUFFX2 U5327 ( .INP(n5219), .Z(n5138) );
  NBUFFX2 U5328 ( .INP(n5218), .Z(n5139) );
  NBUFFX2 U5329 ( .INP(n5218), .Z(n5140) );
  NBUFFX2 U5330 ( .INP(n5218), .Z(n5141) );
  NBUFFX2 U5331 ( .INP(n5217), .Z(n5142) );
  NBUFFX2 U5332 ( .INP(n5217), .Z(n5143) );
  NBUFFX2 U5333 ( .INP(n5217), .Z(n5144) );
  NBUFFX2 U5334 ( .INP(n5216), .Z(n5145) );
  NBUFFX2 U5335 ( .INP(n5216), .Z(n5146) );
  NBUFFX2 U5336 ( .INP(n5216), .Z(n5147) );
  NBUFFX2 U5337 ( .INP(n5215), .Z(n5148) );
  NBUFFX2 U5338 ( .INP(n5215), .Z(n5149) );
  NBUFFX2 U5339 ( .INP(n5215), .Z(n5150) );
  NBUFFX2 U5340 ( .INP(n5214), .Z(n5151) );
  NBUFFX2 U5341 ( .INP(n5214), .Z(n5152) );
  NBUFFX2 U5342 ( .INP(n5214), .Z(n5153) );
  NBUFFX2 U5343 ( .INP(n5213), .Z(n5154) );
  NBUFFX2 U5344 ( .INP(n5213), .Z(n5155) );
  NBUFFX2 U5345 ( .INP(n5213), .Z(n5156) );
  NBUFFX2 U5346 ( .INP(n5212), .Z(n5157) );
  NBUFFX2 U5347 ( .INP(n5212), .Z(n5158) );
  NBUFFX2 U5348 ( .INP(n5212), .Z(n5159) );
  NBUFFX2 U5349 ( .INP(n5211), .Z(n5160) );
  NBUFFX2 U5350 ( .INP(n5211), .Z(n5161) );
  NBUFFX2 U5351 ( .INP(n5211), .Z(n5162) );
  NBUFFX2 U5352 ( .INP(n5210), .Z(n5163) );
  NBUFFX2 U5353 ( .INP(n5210), .Z(n5164) );
  NBUFFX2 U5354 ( .INP(n5210), .Z(n5165) );
  NBUFFX2 U5355 ( .INP(n5209), .Z(n5166) );
  NBUFFX2 U5356 ( .INP(n5209), .Z(n5167) );
  NBUFFX2 U5357 ( .INP(n5209), .Z(n5168) );
  NBUFFX2 U5358 ( .INP(n5208), .Z(n5169) );
  NBUFFX2 U5359 ( .INP(n5208), .Z(n5170) );
  NBUFFX2 U5360 ( .INP(n5208), .Z(n5171) );
  NBUFFX2 U5361 ( .INP(n5207), .Z(n5172) );
  NBUFFX2 U5362 ( .INP(n5207), .Z(n5173) );
  NBUFFX2 U5363 ( .INP(n5207), .Z(n5174) );
  NBUFFX2 U5364 ( .INP(n5206), .Z(n5175) );
  NBUFFX2 U5365 ( .INP(n5206), .Z(n5176) );
  NBUFFX2 U5366 ( .INP(n5206), .Z(n5177) );
  NBUFFX2 U5367 ( .INP(n5205), .Z(n5178) );
  NBUFFX2 U5368 ( .INP(n5205), .Z(n5179) );
  NBUFFX2 U5369 ( .INP(n5205), .Z(n5180) );
  NBUFFX2 U5370 ( .INP(n5204), .Z(n5181) );
  NBUFFX2 U5371 ( .INP(n5204), .Z(n5182) );
  NBUFFX2 U5372 ( .INP(n5204), .Z(n5183) );
  NBUFFX2 U5373 ( .INP(n5203), .Z(n5184) );
  NBUFFX2 U5374 ( .INP(n5203), .Z(n5185) );
  NBUFFX2 U5375 ( .INP(n5203), .Z(n5186) );
  NBUFFX2 U5376 ( .INP(n5202), .Z(n5187) );
  NBUFFX2 U5377 ( .INP(n5202), .Z(n5188) );
  NBUFFX2 U5378 ( .INP(n5202), .Z(n5189) );
  NBUFFX2 U5379 ( .INP(n5201), .Z(n5190) );
  NBUFFX2 U5380 ( .INP(n5201), .Z(n5191) );
  NBUFFX2 U5381 ( .INP(n5201), .Z(n5192) );
  NBUFFX2 U5382 ( .INP(n5200), .Z(n5193) );
  NBUFFX2 U5383 ( .INP(n5200), .Z(n5194) );
  NBUFFX2 U5384 ( .INP(n5200), .Z(n5195) );
  NBUFFX2 U5385 ( .INP(n5199), .Z(n5196) );
  NBUFFX2 U5386 ( .INP(n5199), .Z(n5197) );
  NBUFFX2 U5387 ( .INP(n5199), .Z(n5198) );
  NBUFFX2 U5388 ( .INP(n5242), .Z(n5199) );
  NBUFFX2 U5389 ( .INP(n5242), .Z(n5200) );
  NBUFFX2 U5390 ( .INP(n5242), .Z(n5201) );
  NBUFFX2 U5391 ( .INP(n5241), .Z(n5202) );
  NBUFFX2 U5392 ( .INP(n5241), .Z(n5203) );
  NBUFFX2 U5393 ( .INP(n5241), .Z(n5204) );
  NBUFFX2 U5394 ( .INP(n5240), .Z(n5205) );
  NBUFFX2 U5395 ( .INP(n5240), .Z(n5206) );
  NBUFFX2 U5396 ( .INP(n5240), .Z(n5207) );
  NBUFFX2 U5397 ( .INP(n5239), .Z(n5208) );
  NBUFFX2 U5398 ( .INP(n5239), .Z(n5209) );
  NBUFFX2 U5399 ( .INP(n5239), .Z(n5210) );
  NBUFFX2 U5400 ( .INP(n5238), .Z(n5211) );
  NBUFFX2 U5401 ( .INP(n5238), .Z(n5212) );
  NBUFFX2 U5402 ( .INP(n5238), .Z(n5213) );
  NBUFFX2 U5403 ( .INP(n5237), .Z(n5214) );
  NBUFFX2 U5404 ( .INP(n5237), .Z(n5215) );
  NBUFFX2 U5405 ( .INP(n5237), .Z(n5216) );
  NBUFFX2 U5406 ( .INP(n5236), .Z(n5217) );
  NBUFFX2 U5407 ( .INP(n5236), .Z(n5218) );
  NBUFFX2 U5408 ( .INP(n5236), .Z(n5219) );
  NBUFFX2 U5409 ( .INP(n5235), .Z(n5220) );
  NBUFFX2 U5410 ( .INP(n5235), .Z(n5221) );
  NBUFFX2 U5411 ( .INP(n5235), .Z(n5222) );
  NBUFFX2 U5412 ( .INP(n5234), .Z(n5223) );
  NBUFFX2 U5413 ( .INP(n5234), .Z(n5224) );
  NBUFFX2 U5414 ( .INP(n5234), .Z(n5225) );
  NBUFFX2 U5415 ( .INP(n5233), .Z(n5226) );
  NBUFFX2 U5416 ( .INP(n5233), .Z(n5227) );
  NBUFFX2 U5417 ( .INP(n5233), .Z(n5228) );
  NBUFFX2 U5418 ( .INP(n5232), .Z(n5229) );
  NBUFFX2 U5419 ( .INP(n5232), .Z(n5230) );
  NBUFFX2 U5420 ( .INP(n5232), .Z(n5231) );
  NBUFFX2 U5421 ( .INP(n5246), .Z(n5232) );
  NBUFFX2 U5422 ( .INP(n5246), .Z(n5233) );
  NBUFFX2 U5423 ( .INP(n5245), .Z(n5234) );
  NBUFFX2 U5424 ( .INP(n5245), .Z(n5235) );
  NBUFFX2 U5425 ( .INP(n5245), .Z(n5236) );
  NBUFFX2 U5426 ( .INP(n5244), .Z(n5237) );
  NBUFFX2 U5427 ( .INP(n5244), .Z(n5238) );
  NBUFFX2 U5428 ( .INP(n5244), .Z(n5239) );
  NBUFFX2 U5429 ( .INP(n5243), .Z(n5240) );
  NBUFFX2 U5430 ( .INP(n5243), .Z(n5241) );
  NBUFFX2 U5431 ( .INP(n5243), .Z(n5242) );
  NBUFFX2 U5432 ( .INP(test_se), .Z(n5243) );
  NBUFFX2 U5433 ( .INP(test_se), .Z(n5244) );
  NBUFFX2 U5434 ( .INP(test_se), .Z(n5245) );
  NBUFFX2 U5435 ( .INP(test_se), .Z(n5246) );
  NBUFFX2 U5436 ( .INP(TM1), .Z(n5260) );
  NBUFFX2 U5437 ( .INP(TM1), .Z(n5261) );
  NBUFFX2 U5438 ( .INP(TM1), .Z(n5262) );
  NBUFFX2 U5439 ( .INP(n5342), .Z(n5325) );
  NBUFFX2 U5440 ( .INP(n5341), .Z(n5326) );
  NBUFFX2 U5441 ( .INP(n5341), .Z(n5327) );
  NBUFFX2 U5442 ( .INP(n5341), .Z(n5328) );
  NBUFFX2 U5443 ( .INP(n5340), .Z(n5329) );
  NBUFFX2 U5444 ( .INP(n5340), .Z(n5330) );
  NBUFFX2 U5445 ( .INP(n5340), .Z(n5331) );
  NBUFFX2 U5446 ( .INP(n5339), .Z(n5332) );
  NBUFFX2 U5447 ( .INP(n5339), .Z(n5333) );
  NBUFFX2 U5448 ( .INP(n5339), .Z(n5334) );
  NBUFFX2 U5449 ( .INP(n5338), .Z(n5335) );
  NBUFFX2 U5450 ( .INP(n5338), .Z(n5336) );
  NBUFFX2 U5451 ( .INP(n5338), .Z(n5337) );
  NBUFFX2 U5452 ( .INP(RESET), .Z(n5338) );
  NBUFFX2 U5453 ( .INP(RESET), .Z(n5339) );
  NBUFFX2 U5454 ( .INP(RESET), .Z(n5340) );
  NBUFFX2 U5455 ( .INP(RESET), .Z(n5341) );
  NBUFFX2 U5456 ( .INP(RESET), .Z(n5342) );
  INVX0 U5457 ( .INP(n5263), .ZN(n5343) );
  INVX0 U5458 ( .INP(n5263), .ZN(n5344) );
  INVX0 U5459 ( .INP(n5263), .ZN(n5345) );
  INVX0 U5460 ( .INP(n5263), .ZN(n5346) );
  INVX0 U5461 ( .INP(n5263), .ZN(n5347) );
  INVX0 U5462 ( .INP(n5264), .ZN(n5348) );
  INVX0 U5463 ( .INP(n5264), .ZN(n5349) );
  INVX0 U5464 ( .INP(n5264), .ZN(n5350) );
  INVX0 U5465 ( .INP(n5264), .ZN(n5351) );
  INVX0 U5466 ( .INP(n5264), .ZN(n5352) );
  INVX0 U5467 ( .INP(n5265), .ZN(n5353) );
  INVX0 U5468 ( .INP(n5266), .ZN(n5354) );
  INVX0 U5469 ( .INP(n5266), .ZN(n5355) );
  INVX0 U5470 ( .INP(n5266), .ZN(n5356) );
  INVX0 U5471 ( .INP(n5266), .ZN(n5357) );
  INVX0 U5472 ( .INP(n5266), .ZN(n5358) );
  INVX0 U5473 ( .INP(n5267), .ZN(n5359) );
  INVX0 U5474 ( .INP(n5267), .ZN(n5360) );
  INVX0 U5475 ( .INP(n5267), .ZN(n5361) );
  INVX0 U5476 ( .INP(n5267), .ZN(n5362) );
  INVX0 U5477 ( .INP(n5267), .ZN(n5363) );
  INVX0 U5478 ( .INP(n5268), .ZN(n5364) );
  INVX0 U5479 ( .INP(n5268), .ZN(n5365) );
  INVX0 U5480 ( .INP(n5268), .ZN(n5366) );
  INVX0 U5481 ( .INP(n5268), .ZN(n5367) );
  INVX0 U5482 ( .INP(n5268), .ZN(n5368) );
  INVX0 U5483 ( .INP(n5269), .ZN(n5369) );
  INVX0 U5484 ( .INP(n5269), .ZN(n5370) );
  INVX0 U5485 ( .INP(n5269), .ZN(n5371) );
  INVX0 U5486 ( .INP(n5269), .ZN(n5372) );
  INVX0 U5487 ( .INP(n5269), .ZN(n5373) );
  INVX0 U5488 ( .INP(n5270), .ZN(n5374) );
  INVX0 U5489 ( .INP(n5270), .ZN(n5375) );
  INVX0 U5490 ( .INP(n5270), .ZN(n5376) );
  INVX0 U5491 ( .INP(n5270), .ZN(n5377) );
  INVX0 U5492 ( .INP(n5270), .ZN(n5378) );
  INVX0 U5493 ( .INP(n5271), .ZN(n5379) );
  INVX0 U5494 ( .INP(n5271), .ZN(n5380) );
  INVX0 U5495 ( .INP(n5271), .ZN(n5381) );
  INVX0 U5496 ( .INP(n5271), .ZN(n5382) );
  INVX0 U5497 ( .INP(n5271), .ZN(n5383) );
  INVX0 U5498 ( .INP(n5272), .ZN(n5384) );
  INVX0 U5499 ( .INP(n5272), .ZN(n5385) );
  INVX0 U5500 ( .INP(n5272), .ZN(n5386) );
  INVX0 U5501 ( .INP(n5272), .ZN(n5387) );
  INVX0 U5502 ( .INP(n5272), .ZN(n5388) );
  INVX0 U5503 ( .INP(n5273), .ZN(n5389) );
  INVX0 U5504 ( .INP(n5273), .ZN(n5390) );
  INVX0 U5505 ( .INP(n5273), .ZN(n5391) );
  INVX0 U5506 ( .INP(n5273), .ZN(n5392) );
  INVX0 U5507 ( .INP(n5274), .ZN(n5393) );
  INVX0 U5508 ( .INP(n5274), .ZN(n5394) );
  INVX0 U5509 ( .INP(n5274), .ZN(n5395) );
  INVX0 U5510 ( .INP(n5274), .ZN(n5396) );
  INVX0 U5511 ( .INP(n5274), .ZN(n5397) );
  INVX0 U5512 ( .INP(n5275), .ZN(n5398) );
  INVX0 U5513 ( .INP(n5275), .ZN(n5399) );
  INVX0 U5514 ( .INP(n5275), .ZN(n5400) );
  INVX0 U5515 ( .INP(n5275), .ZN(n5401) );
  INVX0 U5516 ( .INP(n5275), .ZN(n5402) );
  INVX0 U5517 ( .INP(n5276), .ZN(n5403) );
  INVX0 U5518 ( .INP(n5276), .ZN(n5404) );
  INVX0 U5519 ( .INP(n5276), .ZN(n5405) );
  INVX0 U5520 ( .INP(n5276), .ZN(n5406) );
  INVX0 U5521 ( .INP(n5276), .ZN(n5407) );
  INVX0 U5522 ( .INP(n5277), .ZN(n5408) );
  INVX0 U5523 ( .INP(n5277), .ZN(n5409) );
  INVX0 U5524 ( .INP(n5277), .ZN(n5410) );
  INVX0 U5525 ( .INP(n5277), .ZN(n5411) );
  INVX0 U5526 ( .INP(n5277), .ZN(n5412) );
  INVX0 U5527 ( .INP(n5278), .ZN(n5413) );
  INVX0 U5528 ( .INP(n5278), .ZN(n5414) );
  INVX0 U5529 ( .INP(n5278), .ZN(n5415) );
  INVX0 U5530 ( .INP(n5278), .ZN(n5416) );
  INVX0 U5531 ( .INP(n5278), .ZN(n5417) );
  INVX0 U5532 ( .INP(n5279), .ZN(n5418) );
  INVX0 U5533 ( .INP(n5279), .ZN(n5419) );
  INVX0 U5534 ( .INP(n5279), .ZN(n5420) );
  INVX0 U5535 ( .INP(n5279), .ZN(n5421) );
  INVX0 U5536 ( .INP(n5279), .ZN(n5422) );
  INVX0 U5537 ( .INP(n5280), .ZN(n5423) );
  INVX0 U5538 ( .INP(n5280), .ZN(n5424) );
  INVX0 U5539 ( .INP(n5280), .ZN(n5425) );
  INVX0 U5540 ( .INP(n5280), .ZN(n5426) );
  INVX0 U5541 ( .INP(n5280), .ZN(n5427) );
  INVX0 U5542 ( .INP(n5281), .ZN(n5428) );
  INVX0 U5543 ( .INP(n5281), .ZN(n5429) );
  INVX0 U5544 ( .INP(n5281), .ZN(n5430) );
  INVX0 U5545 ( .INP(n5281), .ZN(n5431) );
  INVX0 U5546 ( .INP(n5281), .ZN(n5432) );
  INVX0 U5547 ( .INP(n5282), .ZN(n5433) );
  INVX0 U5548 ( .INP(n5282), .ZN(n5434) );
  INVX0 U5549 ( .INP(n5282), .ZN(n5435) );
  INVX0 U5550 ( .INP(n5282), .ZN(n5436) );
  INVX0 U5551 ( .INP(n5282), .ZN(n5437) );
  INVX0 U5552 ( .INP(n5283), .ZN(n5438) );
  INVX0 U5553 ( .INP(n5283), .ZN(n5439) );
  INVX0 U5554 ( .INP(n5283), .ZN(n5440) );
  INVX0 U5555 ( .INP(n5283), .ZN(n5441) );
  NBUFFX2 U5556 ( .INP(n5624), .Z(n5586) );
  NBUFFX2 U5557 ( .INP(n5624), .Z(n5587) );
  NBUFFX2 U5558 ( .INP(n5623), .Z(n5588) );
  NBUFFX2 U5559 ( .INP(n5623), .Z(n5589) );
  NBUFFX2 U5560 ( .INP(n5623), .Z(n5590) );
  NBUFFX2 U5561 ( .INP(n5622), .Z(n5591) );
  NBUFFX2 U5562 ( .INP(n5622), .Z(n5592) );
  NBUFFX2 U5563 ( .INP(n5622), .Z(n5593) );
  NBUFFX2 U5564 ( .INP(n5621), .Z(n5594) );
  NBUFFX2 U5565 ( .INP(n5621), .Z(n5595) );
  NBUFFX2 U5566 ( .INP(n5621), .Z(n5596) );
  NBUFFX2 U5567 ( .INP(n5620), .Z(n5597) );
  NBUFFX2 U5568 ( .INP(n5620), .Z(n5598) );
  NBUFFX2 U5569 ( .INP(n5620), .Z(n5599) );
  NBUFFX2 U5570 ( .INP(n5619), .Z(n5600) );
  NBUFFX2 U5571 ( .INP(n5619), .Z(n5601) );
  NBUFFX2 U5572 ( .INP(n5619), .Z(n5602) );
  NBUFFX2 U5573 ( .INP(n5618), .Z(n5603) );
  NBUFFX2 U5574 ( .INP(n5618), .Z(n5604) );
  NBUFFX2 U5575 ( .INP(n5618), .Z(n5605) );
  NBUFFX2 U5576 ( .INP(n5617), .Z(n5606) );
  NBUFFX2 U5577 ( .INP(n5617), .Z(n5607) );
  NBUFFX2 U5578 ( .INP(n5617), .Z(n5608) );
  NBUFFX2 U5579 ( .INP(n5616), .Z(n5609) );
  NBUFFX2 U5580 ( .INP(n5616), .Z(n5610) );
  NBUFFX2 U5581 ( .INP(n5616), .Z(n5611) );
  NBUFFX2 U5582 ( .INP(n5615), .Z(n5612) );
  NBUFFX2 U5583 ( .INP(n5615), .Z(n5613) );
  NBUFFX2 U5584 ( .INP(n5615), .Z(n5614) );
  NBUFFX2 U5585 ( .INP(CK), .Z(n5615) );
  NBUFFX2 U5586 ( .INP(CK), .Z(n5616) );
  NBUFFX2 U5587 ( .INP(n5624), .Z(n5617) );
  NBUFFX2 U5588 ( .INP(CK), .Z(n5618) );
  NBUFFX2 U5589 ( .INP(n5620), .Z(n5619) );
  NBUFFX2 U5590 ( .INP(CK), .Z(n5620) );
  NBUFFX2 U5591 ( .INP(n5615), .Z(n5621) );
  NBUFFX2 U5592 ( .INP(n5616), .Z(n5622) );
  NBUFFX2 U5593 ( .INP(n5618), .Z(n5623) );
  NBUFFX2 U5594 ( .INP(n5455), .Z(n5624) );
  INVX0 U5595 ( .INP(n5625), .ZN(n9) );
  NOR2X0 U5596 ( .IN1(n5626), .IN2(n5627), .QN(n5625) );
  NAND2X0 U5597 ( .IN1(n5628), .IN2(n5629), .QN(n5627) );
  NAND2X0 U5598 ( .IN1(n4738), .IN2(n5630), .QN(n5629) );
  NAND2X0 U5599 ( .IN1(n2152), .IN2(CRC_OUT_9_22), .QN(n5628) );
  NAND2X0 U5600 ( .IN1(n5631), .IN2(n5632), .QN(n5626) );
  NAND2X0 U5601 ( .IN1(n2153), .IN2(n5633), .QN(n5632) );
  INVX0 U5602 ( .INP(n5634), .ZN(n5633) );
  NAND2X0 U5603 ( .IN1(WX500), .IN2(n4807), .QN(n5631) );
  INVX0 U5604 ( .INP(n5635), .ZN(n85) );
  INVX0 U5605 ( .INP(n5636), .ZN(n84) );
  INVX0 U5606 ( .INP(n5637), .ZN(n83) );
  INVX0 U5607 ( .INP(n5638), .ZN(n82) );
  INVX0 U5608 ( .INP(n5639), .ZN(n81) );
  INVX0 U5609 ( .INP(n5640), .ZN(n80) );
  INVX0 U5610 ( .INP(n5641), .ZN(n8) );
  NOR2X0 U5611 ( .IN1(n5642), .IN2(n5643), .QN(n5641) );
  NAND2X0 U5612 ( .IN1(n5644), .IN2(n5645), .QN(n5643) );
  NAND2X0 U5613 ( .IN1(n4735), .IN2(n5646), .QN(n5645) );
  NAND2X0 U5614 ( .IN1(n2152), .IN2(CRC_OUT_9_23), .QN(n5644) );
  NAND2X0 U5615 ( .IN1(n5647), .IN2(n5648), .QN(n5642) );
  NAND2X0 U5616 ( .IN1(n2153), .IN2(n5649), .QN(n5648) );
  NAND2X0 U5617 ( .IN1(WX498), .IN2(n4812), .QN(n5647) );
  INVX0 U5618 ( .INP(n5650), .ZN(n79) );
  INVX0 U5619 ( .INP(n5651), .ZN(n78) );
  INVX0 U5620 ( .INP(n5652), .ZN(n77) );
  INVX0 U5621 ( .INP(n5653), .ZN(n76) );
  INVX0 U5622 ( .INP(n5654), .ZN(n75) );
  INVX0 U5623 ( .INP(n5655), .ZN(n74) );
  INVX0 U5624 ( .INP(n5656), .ZN(n73) );
  INVX0 U5625 ( .INP(n5657), .ZN(n72) );
  INVX0 U5626 ( .INP(n5658), .ZN(n71) );
  INVX0 U5627 ( .INP(n5659), .ZN(n70) );
  INVX0 U5628 ( .INP(n5660), .ZN(n7) );
  NOR2X0 U5629 ( .IN1(n5661), .IN2(n5662), .QN(n5660) );
  NAND2X0 U5630 ( .IN1(n5663), .IN2(n5664), .QN(n5662) );
  NAND2X0 U5631 ( .IN1(n4735), .IN2(n5665), .QN(n5664) );
  NAND2X0 U5632 ( .IN1(n2152), .IN2(CRC_OUT_9_25), .QN(n5663) );
  NAND2X0 U5633 ( .IN1(n5666), .IN2(n5667), .QN(n5661) );
  NAND2X0 U5634 ( .IN1(n2153), .IN2(n5668), .QN(n5667) );
  NAND2X0 U5635 ( .IN1(WX494), .IN2(n4812), .QN(n5666) );
  INVX0 U5636 ( .INP(n5669), .ZN(n69) );
  INVX0 U5637 ( .INP(n5670), .ZN(n68) );
  INVX0 U5638 ( .INP(n5671), .ZN(n67) );
  INVX0 U5639 ( .INP(n5672), .ZN(n66) );
  INVX0 U5640 ( .INP(n5673), .ZN(n65) );
  INVX0 U5641 ( .INP(n5674), .ZN(n64) );
  INVX0 U5642 ( .INP(n5675), .ZN(n63) );
  INVX0 U5643 ( .INP(n5676), .ZN(n62) );
  INVX0 U5644 ( .INP(n5677), .ZN(n61) );
  INVX0 U5645 ( .INP(n5678), .ZN(n60) );
  INVX0 U5646 ( .INP(n5679), .ZN(n6) );
  NOR2X0 U5647 ( .IN1(n5680), .IN2(n5681), .QN(n5679) );
  NAND2X0 U5648 ( .IN1(n5682), .IN2(n5683), .QN(n5681) );
  NAND2X0 U5649 ( .IN1(n4735), .IN2(n5684), .QN(n5683) );
  NAND2X0 U5650 ( .IN1(n2152), .IN2(CRC_OUT_9_26), .QN(n5682) );
  NAND2X0 U5651 ( .IN1(n5685), .IN2(n5686), .QN(n5680) );
  NAND2X0 U5652 ( .IN1(n2153), .IN2(n5687), .QN(n5686) );
  NAND2X0 U5653 ( .IN1(WX492), .IN2(n4812), .QN(n5685) );
  INVX0 U5654 ( .INP(n5688), .ZN(n59) );
  INVX0 U5655 ( .INP(TM0), .ZN(n583) );
  INVX0 U5656 ( .INP(n5689), .ZN(n58) );
  INVX0 U5657 ( .INP(n5690), .ZN(n57) );
  INVX0 U5658 ( .INP(n5691), .ZN(n56) );
  INVX0 U5659 ( .INP(n5692), .ZN(n55) );
  INVX0 U5660 ( .INP(n5693), .ZN(n5) );
  NOR2X0 U5661 ( .IN1(n5694), .IN2(n5695), .QN(n5693) );
  NAND2X0 U5662 ( .IN1(n5696), .IN2(n5697), .QN(n5695) );
  NAND2X0 U5663 ( .IN1(n4735), .IN2(n5698), .QN(n5697) );
  NAND2X0 U5664 ( .IN1(n2152), .IN2(CRC_OUT_9_27), .QN(n5696) );
  NAND2X0 U5665 ( .IN1(n5699), .IN2(n5700), .QN(n5694) );
  NAND2X0 U5666 ( .IN1(n2153), .IN2(n5701), .QN(n5700) );
  NAND2X0 U5667 ( .IN1(WX490), .IN2(n4812), .QN(n5699) );
  INVX0 U5668 ( .INP(n5702), .ZN(n494) );
  NOR2X0 U5669 ( .IN1(n5703), .IN2(n5704), .QN(n5702) );
  NAND2X0 U5670 ( .IN1(n5705), .IN2(n5706), .QN(n5704) );
  NAND2X0 U5671 ( .IN1(DATA_0_0), .IN2(n2153), .QN(n5706) );
  NAND2X0 U5672 ( .IN1(n2152), .IN2(CRC_OUT_1_0), .QN(n5705) );
  NAND2X0 U5673 ( .IN1(n5707), .IN2(n5708), .QN(n5703) );
  NAND2X0 U5674 ( .IN1(n4735), .IN2(n5709), .QN(n5708) );
  NAND2X0 U5675 ( .IN1(n495), .IN2(n4812), .QN(n5707) );
  INVX0 U5676 ( .INP(n5710), .ZN(n495) );
  NAND2X0 U5677 ( .IN1(n5295), .IN2(n8263), .QN(n5710) );
  INVX0 U5678 ( .INP(n5711), .ZN(n492) );
  NOR2X0 U5679 ( .IN1(n5712), .IN2(n5713), .QN(n5711) );
  NAND2X0 U5680 ( .IN1(n5714), .IN2(n5715), .QN(n5713) );
  NAND2X0 U5681 ( .IN1(DATA_0_1), .IN2(n2153), .QN(n5715) );
  NAND2X0 U5682 ( .IN1(n2152), .IN2(CRC_OUT_1_1), .QN(n5714) );
  NAND2X0 U5683 ( .IN1(n5716), .IN2(n5717), .QN(n5712) );
  NAND2X0 U5684 ( .IN1(n4735), .IN2(n5718), .QN(n5717) );
  NAND2X0 U5685 ( .IN1(n493), .IN2(n4812), .QN(n5716) );
  INVX0 U5686 ( .INP(n5719), .ZN(n493) );
  NAND2X0 U5687 ( .IN1(n5295), .IN2(n8264), .QN(n5719) );
  INVX0 U5688 ( .INP(n5720), .ZN(n490) );
  NOR2X0 U5689 ( .IN1(n5721), .IN2(n5722), .QN(n5720) );
  NAND2X0 U5690 ( .IN1(n5723), .IN2(n5724), .QN(n5722) );
  NAND2X0 U5691 ( .IN1(DATA_0_2), .IN2(n2153), .QN(n5724) );
  NAND2X0 U5692 ( .IN1(n2152), .IN2(CRC_OUT_1_2), .QN(n5723) );
  NAND2X0 U5693 ( .IN1(n5725), .IN2(n5726), .QN(n5721) );
  NAND2X0 U5694 ( .IN1(n5727), .IN2(n4741), .QN(n5726) );
  INVX0 U5695 ( .INP(n5728), .ZN(n5727) );
  NAND2X0 U5696 ( .IN1(n491), .IN2(n4812), .QN(n5725) );
  INVX0 U5697 ( .INP(n5729), .ZN(n491) );
  NAND2X0 U5698 ( .IN1(n5294), .IN2(n8265), .QN(n5729) );
  INVX0 U5699 ( .INP(n5730), .ZN(n488) );
  NOR2X0 U5700 ( .IN1(n5731), .IN2(n5732), .QN(n5730) );
  NAND2X0 U5701 ( .IN1(n5733), .IN2(n5734), .QN(n5732) );
  NAND2X0 U5702 ( .IN1(DATA_0_3), .IN2(n2153), .QN(n5734) );
  NAND2X0 U5703 ( .IN1(n2152), .IN2(CRC_OUT_1_3), .QN(n5733) );
  NAND2X0 U5704 ( .IN1(n5735), .IN2(n5736), .QN(n5731) );
  NAND2X0 U5705 ( .IN1(n4736), .IN2(n5737), .QN(n5736) );
  NAND2X0 U5706 ( .IN1(n489), .IN2(n4812), .QN(n5735) );
  INVX0 U5707 ( .INP(n5738), .ZN(n489) );
  NAND2X0 U5708 ( .IN1(n5294), .IN2(n8266), .QN(n5738) );
  INVX0 U5709 ( .INP(n5739), .ZN(n486) );
  NOR2X0 U5710 ( .IN1(n5740), .IN2(n5741), .QN(n5739) );
  NAND2X0 U5711 ( .IN1(n5742), .IN2(n5743), .QN(n5741) );
  NAND2X0 U5712 ( .IN1(DATA_0_4), .IN2(n2153), .QN(n5743) );
  NAND2X0 U5713 ( .IN1(n2152), .IN2(CRC_OUT_1_4), .QN(n5742) );
  NAND2X0 U5714 ( .IN1(n5744), .IN2(n5745), .QN(n5740) );
  NAND2X0 U5715 ( .IN1(n5746), .IN2(n4740), .QN(n5745) );
  INVX0 U6483 ( .INP(n5747), .ZN(n5746) );
  NAND2X0 U6484 ( .IN1(n487), .IN2(n4812), .QN(n5744) );
  INVX0 U6485 ( .INP(n5748), .ZN(n487) );
  NAND2X0 U6486 ( .IN1(n5294), .IN2(n8267), .QN(n5748) );
  INVX0 U6487 ( .INP(n5749), .ZN(n484) );
  NOR2X0 U6488 ( .IN1(n5750), .IN2(n5751), .QN(n5749) );
  NAND2X0 U6489 ( .IN1(n5752), .IN2(n5753), .QN(n5751) );
  NAND2X0 U6490 ( .IN1(DATA_0_5), .IN2(n2153), .QN(n5753) );
  NAND2X0 U6491 ( .IN1(n2152), .IN2(CRC_OUT_1_5), .QN(n5752) );
  NAND2X0 U6492 ( .IN1(n5754), .IN2(n5755), .QN(n5750) );
  NAND2X0 U6493 ( .IN1(n4736), .IN2(n5756), .QN(n5755) );
  NAND2X0 U6494 ( .IN1(n485), .IN2(n4812), .QN(n5754) );
  INVX0 U6495 ( .INP(n5757), .ZN(n485) );
  NAND2X0 U6496 ( .IN1(n5294), .IN2(n8268), .QN(n5757) );
  INVX0 U6497 ( .INP(n5758), .ZN(n482) );
  NOR2X0 U6498 ( .IN1(n5759), .IN2(n5760), .QN(n5758) );
  NAND2X0 U6499 ( .IN1(n5761), .IN2(n5762), .QN(n5760) );
  NAND2X0 U6500 ( .IN1(DATA_0_6), .IN2(n2153), .QN(n5762) );
  NAND2X0 U6501 ( .IN1(n2152), .IN2(CRC_OUT_1_6), .QN(n5761) );
  NAND2X0 U6502 ( .IN1(n5763), .IN2(n5764), .QN(n5759) );
  NAND2X0 U6503 ( .IN1(n5765), .IN2(n4740), .QN(n5764) );
  INVX0 U6504 ( .INP(n5766), .ZN(n5765) );
  NAND2X0 U6505 ( .IN1(n483), .IN2(n4811), .QN(n5763) );
  INVX0 U6506 ( .INP(n5767), .ZN(n483) );
  NAND2X0 U6507 ( .IN1(n5294), .IN2(n8269), .QN(n5767) );
  INVX0 U6508 ( .INP(n5768), .ZN(n480) );
  NOR2X0 U6509 ( .IN1(n5769), .IN2(n5770), .QN(n5768) );
  NAND2X0 U6510 ( .IN1(n5771), .IN2(n5772), .QN(n5770) );
  NAND2X0 U6511 ( .IN1(DATA_0_7), .IN2(n2153), .QN(n5772) );
  NAND2X0 U6512 ( .IN1(n2152), .IN2(CRC_OUT_1_7), .QN(n5771) );
  NAND2X0 U6513 ( .IN1(n5773), .IN2(n5774), .QN(n5769) );
  NAND2X0 U6514 ( .IN1(n4736), .IN2(n5775), .QN(n5774) );
  NAND2X0 U6515 ( .IN1(n481), .IN2(n4811), .QN(n5773) );
  INVX0 U6516 ( .INP(n5776), .ZN(n481) );
  NAND2X0 U6517 ( .IN1(n5294), .IN2(n8270), .QN(n5776) );
  INVX0 U6518 ( .INP(n5777), .ZN(n478) );
  NOR2X0 U6519 ( .IN1(n5778), .IN2(n5779), .QN(n5777) );
  NAND2X0 U6520 ( .IN1(n5780), .IN2(n5781), .QN(n5779) );
  NAND2X0 U6521 ( .IN1(DATA_0_8), .IN2(n2153), .QN(n5781) );
  NAND2X0 U6522 ( .IN1(n2152), .IN2(CRC_OUT_1_8), .QN(n5780) );
  NAND2X0 U6523 ( .IN1(n5782), .IN2(n5783), .QN(n5778) );
  NAND2X0 U6524 ( .IN1(n5784), .IN2(n4740), .QN(n5783) );
  INVX0 U6525 ( .INP(n5785), .ZN(n5784) );
  NAND2X0 U6526 ( .IN1(n479), .IN2(n4811), .QN(n5782) );
  INVX0 U6527 ( .INP(n5786), .ZN(n479) );
  NAND2X0 U6528 ( .IN1(n5293), .IN2(n8271), .QN(n5786) );
  INVX0 U6529 ( .INP(n5787), .ZN(n476) );
  NOR2X0 U6530 ( .IN1(n5788), .IN2(n5789), .QN(n5787) );
  NAND2X0 U6531 ( .IN1(n5790), .IN2(n5791), .QN(n5789) );
  NAND2X0 U6532 ( .IN1(DATA_0_9), .IN2(n2153), .QN(n5791) );
  NAND2X0 U6533 ( .IN1(n2152), .IN2(CRC_OUT_1_9), .QN(n5790) );
  NAND2X0 U6534 ( .IN1(n5792), .IN2(n5793), .QN(n5788) );
  NAND2X0 U6535 ( .IN1(n4736), .IN2(n5794), .QN(n5793) );
  NAND2X0 U6536 ( .IN1(n477), .IN2(n4811), .QN(n5792) );
  INVX0 U6537 ( .INP(n5795), .ZN(n477) );
  NAND2X0 U6538 ( .IN1(n5293), .IN2(n8272), .QN(n5795) );
  INVX0 U6539 ( .INP(n5796), .ZN(n474) );
  NOR2X0 U6540 ( .IN1(n5797), .IN2(n5798), .QN(n5796) );
  NAND2X0 U6541 ( .IN1(n5799), .IN2(n5800), .QN(n5798) );
  NAND2X0 U6542 ( .IN1(DATA_0_10), .IN2(n2153), .QN(n5800) );
  NAND2X0 U6543 ( .IN1(n2152), .IN2(CRC_OUT_1_10), .QN(n5799) );
  NAND2X0 U6544 ( .IN1(n5801), .IN2(n5802), .QN(n5797) );
  NAND2X0 U6545 ( .IN1(n4736), .IN2(n5803), .QN(n5802) );
  NAND2X0 U6546 ( .IN1(n475), .IN2(n4811), .QN(n5801) );
  INVX0 U6547 ( .INP(n5804), .ZN(n475) );
  NAND2X0 U6548 ( .IN1(test_so90), .IN2(n5322), .QN(n5804) );
  INVX0 U6549 ( .INP(n5805), .ZN(n472) );
  NOR2X0 U6550 ( .IN1(n5806), .IN2(n5807), .QN(n5805) );
  NAND2X0 U6551 ( .IN1(n5808), .IN2(n5809), .QN(n5807) );
  NAND2X0 U6552 ( .IN1(DATA_0_11), .IN2(n2153), .QN(n5809) );
  NAND2X0 U6553 ( .IN1(n2152), .IN2(CRC_OUT_1_11), .QN(n5808) );
  NAND2X0 U6554 ( .IN1(n5810), .IN2(n5811), .QN(n5806) );
  NAND2X0 U6555 ( .IN1(n4736), .IN2(n5812), .QN(n5811) );
  NAND2X0 U6556 ( .IN1(n473), .IN2(n4811), .QN(n5810) );
  INVX0 U6557 ( .INP(n5813), .ZN(n473) );
  NAND2X0 U6558 ( .IN1(n5293), .IN2(n8275), .QN(n5813) );
  INVX0 U6559 ( .INP(n5814), .ZN(n470) );
  NOR2X0 U6560 ( .IN1(n5815), .IN2(n5816), .QN(n5814) );
  NAND2X0 U6561 ( .IN1(n5817), .IN2(n5818), .QN(n5816) );
  NAND2X0 U6562 ( .IN1(DATA_0_12), .IN2(n2153), .QN(n5818) );
  NAND2X0 U6563 ( .IN1(n2152), .IN2(CRC_OUT_1_12), .QN(n5817) );
  NAND2X0 U6564 ( .IN1(n5819), .IN2(n5820), .QN(n5815) );
  NAND2X0 U6565 ( .IN1(n4736), .IN2(n5821), .QN(n5820) );
  NAND2X0 U6566 ( .IN1(n471), .IN2(n4811), .QN(n5819) );
  INVX0 U6567 ( .INP(n5822), .ZN(n471) );
  NAND2X0 U6568 ( .IN1(n5293), .IN2(n8276), .QN(n5822) );
  INVX0 U6569 ( .INP(n5823), .ZN(n468) );
  NOR2X0 U6570 ( .IN1(n5824), .IN2(n5825), .QN(n5823) );
  NAND2X0 U6571 ( .IN1(n5826), .IN2(n5827), .QN(n5825) );
  NAND2X0 U6572 ( .IN1(DATA_0_13), .IN2(n2153), .QN(n5827) );
  NAND2X0 U6573 ( .IN1(n2152), .IN2(CRC_OUT_1_13), .QN(n5826) );
  NAND2X0 U6574 ( .IN1(n5828), .IN2(n5829), .QN(n5824) );
  NAND2X0 U6575 ( .IN1(n4736), .IN2(n5830), .QN(n5829) );
  NAND2X0 U6576 ( .IN1(n469), .IN2(n4811), .QN(n5828) );
  INVX0 U6577 ( .INP(n5831), .ZN(n469) );
  NAND2X0 U6578 ( .IN1(n5293), .IN2(n8277), .QN(n5831) );
  INVX0 U6579 ( .INP(n5832), .ZN(n466) );
  NOR2X0 U6580 ( .IN1(n5833), .IN2(n5834), .QN(n5832) );
  NAND2X0 U6581 ( .IN1(n5835), .IN2(n5836), .QN(n5834) );
  NAND2X0 U6582 ( .IN1(DATA_0_14), .IN2(n2153), .QN(n5836) );
  NAND2X0 U6583 ( .IN1(test_so99), .IN2(n2152), .QN(n5835) );
  NAND2X0 U6584 ( .IN1(n5837), .IN2(n5838), .QN(n5833) );
  NAND2X0 U6585 ( .IN1(n4736), .IN2(n5839), .QN(n5838) );
  NAND2X0 U6586 ( .IN1(n467), .IN2(n4811), .QN(n5837) );
  INVX0 U6587 ( .INP(n5840), .ZN(n467) );
  NAND2X0 U6588 ( .IN1(n5293), .IN2(n8278), .QN(n5840) );
  INVX0 U6589 ( .INP(n5841), .ZN(n464) );
  NOR2X0 U6590 ( .IN1(n5842), .IN2(n5843), .QN(n5841) );
  NAND2X0 U6591 ( .IN1(n5844), .IN2(n5845), .QN(n5843) );
  NAND2X0 U6592 ( .IN1(DATA_0_15), .IN2(n2153), .QN(n5845) );
  NAND2X0 U6593 ( .IN1(n2152), .IN2(CRC_OUT_1_15), .QN(n5844) );
  NAND2X0 U6594 ( .IN1(n5846), .IN2(n5847), .QN(n5842) );
  NAND2X0 U6595 ( .IN1(n4737), .IN2(n5848), .QN(n5847) );
  NAND2X0 U6596 ( .IN1(n465), .IN2(n4811), .QN(n5846) );
  INVX0 U6597 ( .INP(n5849), .ZN(n465) );
  NAND2X0 U6598 ( .IN1(n5292), .IN2(n8279), .QN(n5849) );
  INVX0 U6599 ( .INP(n5850), .ZN(n462) );
  NOR2X0 U6600 ( .IN1(n5851), .IN2(n5852), .QN(n5850) );
  NAND2X0 U6601 ( .IN1(n5853), .IN2(n5854), .QN(n5852) );
  NAND2X0 U6602 ( .IN1(DATA_0_16), .IN2(n2153), .QN(n5854) );
  NAND2X0 U6603 ( .IN1(n2152), .IN2(CRC_OUT_1_16), .QN(n5853) );
  NAND2X0 U6604 ( .IN1(n5855), .IN2(n5856), .QN(n5851) );
  NAND2X0 U6605 ( .IN1(n4737), .IN2(n5857), .QN(n5856) );
  NAND2X0 U6606 ( .IN1(n463), .IN2(n4810), .QN(n5855) );
  INVX0 U6607 ( .INP(n5858), .ZN(n463) );
  NAND2X0 U6608 ( .IN1(n5292), .IN2(n8280), .QN(n5858) );
  INVX0 U6609 ( .INP(n5859), .ZN(n460) );
  NOR2X0 U6610 ( .IN1(n5860), .IN2(n5861), .QN(n5859) );
  NAND2X0 U6611 ( .IN1(n5862), .IN2(n5863), .QN(n5861) );
  NAND2X0 U6612 ( .IN1(DATA_0_17), .IN2(n2153), .QN(n5863) );
  NAND2X0 U6613 ( .IN1(n2152), .IN2(CRC_OUT_1_17), .QN(n5862) );
  NAND2X0 U6614 ( .IN1(n5864), .IN2(n5865), .QN(n5860) );
  NAND2X0 U6615 ( .IN1(n4737), .IN2(n5866), .QN(n5865) );
  NAND2X0 U6616 ( .IN1(n461), .IN2(n4810), .QN(n5864) );
  INVX0 U6617 ( .INP(n5867), .ZN(n461) );
  NAND2X0 U6618 ( .IN1(n5292), .IN2(n8281), .QN(n5867) );
  INVX0 U6619 ( .INP(n5868), .ZN(n458) );
  NOR2X0 U6620 ( .IN1(n5869), .IN2(n5870), .QN(n5868) );
  NAND2X0 U6621 ( .IN1(n5871), .IN2(n5872), .QN(n5870) );
  NAND2X0 U6622 ( .IN1(DATA_0_18), .IN2(n2153), .QN(n5872) );
  NAND2X0 U6623 ( .IN1(n2152), .IN2(CRC_OUT_1_18), .QN(n5871) );
  NAND2X0 U6624 ( .IN1(n5873), .IN2(n5874), .QN(n5869) );
  NAND2X0 U6625 ( .IN1(n4737), .IN2(n5875), .QN(n5874) );
  NAND2X0 U6626 ( .IN1(n459), .IN2(n4810), .QN(n5873) );
  INVX0 U6627 ( .INP(n5876), .ZN(n459) );
  NAND2X0 U6628 ( .IN1(n5292), .IN2(n8282), .QN(n5876) );
  INVX0 U6629 ( .INP(n5877), .ZN(n456) );
  NOR2X0 U6630 ( .IN1(n5878), .IN2(n5879), .QN(n5877) );
  NAND2X0 U6631 ( .IN1(n5880), .IN2(n5881), .QN(n5879) );
  NAND2X0 U6632 ( .IN1(DATA_0_19), .IN2(n2153), .QN(n5881) );
  NAND2X0 U6633 ( .IN1(n2152), .IN2(CRC_OUT_1_19), .QN(n5880) );
  NAND2X0 U6634 ( .IN1(n5882), .IN2(n5883), .QN(n5878) );
  NAND2X0 U6635 ( .IN1(n5884), .IN2(n4741), .QN(n5883) );
  INVX0 U6636 ( .INP(n5885), .ZN(n5884) );
  NAND2X0 U6637 ( .IN1(n457), .IN2(n4810), .QN(n5882) );
  INVX0 U6638 ( .INP(n5886), .ZN(n457) );
  NAND2X0 U6639 ( .IN1(n5292), .IN2(n8283), .QN(n5886) );
  INVX0 U6640 ( .INP(n5887), .ZN(n454) );
  NOR2X0 U6641 ( .IN1(n5888), .IN2(n5889), .QN(n5887) );
  NAND2X0 U6642 ( .IN1(n5890), .IN2(n5891), .QN(n5889) );
  NAND2X0 U6643 ( .IN1(DATA_0_20), .IN2(n2153), .QN(n5891) );
  NAND2X0 U6644 ( .IN1(n2152), .IN2(CRC_OUT_1_20), .QN(n5890) );
  NAND2X0 U6645 ( .IN1(n5892), .IN2(n5893), .QN(n5888) );
  NAND2X0 U6646 ( .IN1(n4737), .IN2(n5894), .QN(n5893) );
  NAND2X0 U6647 ( .IN1(n455), .IN2(n4810), .QN(n5892) );
  INVX0 U6648 ( .INP(n5895), .ZN(n455) );
  NAND2X0 U6649 ( .IN1(n5292), .IN2(n8284), .QN(n5895) );
  INVX0 U6650 ( .INP(n5896), .ZN(n452) );
  NOR2X0 U6651 ( .IN1(n5897), .IN2(n5898), .QN(n5896) );
  NAND2X0 U6652 ( .IN1(n5899), .IN2(n5900), .QN(n5898) );
  NAND2X0 U6653 ( .IN1(DATA_0_21), .IN2(n2153), .QN(n5900) );
  NAND2X0 U6654 ( .IN1(n2152), .IN2(CRC_OUT_1_21), .QN(n5899) );
  NAND2X0 U6655 ( .IN1(n5901), .IN2(n5902), .QN(n5897) );
  NAND2X0 U6656 ( .IN1(n5903), .IN2(n4740), .QN(n5902) );
  INVX0 U6657 ( .INP(n5904), .ZN(n5903) );
  NAND2X0 U6658 ( .IN1(n453), .IN2(n4810), .QN(n5901) );
  INVX0 U6659 ( .INP(n5905), .ZN(n453) );
  NAND2X0 U6660 ( .IN1(n5291), .IN2(n8285), .QN(n5905) );
  INVX0 U6661 ( .INP(n5906), .ZN(n450) );
  NOR2X0 U6662 ( .IN1(n5907), .IN2(n5908), .QN(n5906) );
  NAND2X0 U6663 ( .IN1(n5909), .IN2(n5910), .QN(n5908) );
  NAND2X0 U6664 ( .IN1(DATA_0_22), .IN2(n2153), .QN(n5910) );
  NAND2X0 U6665 ( .IN1(n2152), .IN2(CRC_OUT_1_22), .QN(n5909) );
  NAND2X0 U6666 ( .IN1(n5911), .IN2(n5912), .QN(n5907) );
  NAND2X0 U6667 ( .IN1(n4737), .IN2(n5913), .QN(n5912) );
  NAND2X0 U6668 ( .IN1(n451), .IN2(n4810), .QN(n5911) );
  INVX0 U6669 ( .INP(n5914), .ZN(n451) );
  NAND2X0 U6670 ( .IN1(n5291), .IN2(n8286), .QN(n5914) );
  INVX0 U6671 ( .INP(n5915), .ZN(n448) );
  NOR2X0 U6672 ( .IN1(n5916), .IN2(n5917), .QN(n5915) );
  NAND2X0 U6673 ( .IN1(n5918), .IN2(n5919), .QN(n5917) );
  NAND2X0 U6674 ( .IN1(DATA_0_23), .IN2(n2153), .QN(n5919) );
  NAND2X0 U6675 ( .IN1(n2152), .IN2(CRC_OUT_1_23), .QN(n5918) );
  NAND2X0 U6676 ( .IN1(n5920), .IN2(n5921), .QN(n5916) );
  NAND2X0 U6677 ( .IN1(n5922), .IN2(n4741), .QN(n5921) );
  INVX0 U6678 ( .INP(n5923), .ZN(n5922) );
  NAND2X0 U6679 ( .IN1(n449), .IN2(n4810), .QN(n5920) );
  INVX0 U6680 ( .INP(n5924), .ZN(n449) );
  NAND2X0 U6681 ( .IN1(n5291), .IN2(n8287), .QN(n5924) );
  INVX0 U6682 ( .INP(n5925), .ZN(n446) );
  NOR2X0 U6683 ( .IN1(n5926), .IN2(n5927), .QN(n5925) );
  NAND2X0 U6684 ( .IN1(n5928), .IN2(n5929), .QN(n5927) );
  NAND2X0 U6685 ( .IN1(DATA_0_24), .IN2(n2153), .QN(n5929) );
  NAND2X0 U6686 ( .IN1(n2152), .IN2(CRC_OUT_1_24), .QN(n5928) );
  NAND2X0 U6687 ( .IN1(n5930), .IN2(n5931), .QN(n5926) );
  NAND2X0 U6688 ( .IN1(n4737), .IN2(n5932), .QN(n5931) );
  NAND2X0 U6689 ( .IN1(n447), .IN2(n4810), .QN(n5930) );
  INVX0 U6690 ( .INP(n5933), .ZN(n447) );
  NAND2X0 U6691 ( .IN1(n5291), .IN2(n8288), .QN(n5933) );
  INVX0 U6692 ( .INP(n5934), .ZN(n444) );
  NOR2X0 U6693 ( .IN1(n5935), .IN2(n5936), .QN(n5934) );
  NAND2X0 U6694 ( .IN1(n5937), .IN2(n5938), .QN(n5936) );
  NAND2X0 U6695 ( .IN1(DATA_0_25), .IN2(n2153), .QN(n5938) );
  NAND2X0 U6696 ( .IN1(n2152), .IN2(CRC_OUT_1_25), .QN(n5937) );
  NAND2X0 U6697 ( .IN1(n5939), .IN2(n5940), .QN(n5935) );
  NAND2X0 U6698 ( .IN1(n5941), .IN2(n4741), .QN(n5940) );
  INVX0 U6699 ( .INP(n5942), .ZN(n5941) );
  NAND2X0 U6700 ( .IN1(n445), .IN2(n4809), .QN(n5939) );
  INVX0 U6701 ( .INP(n5943), .ZN(n445) );
  NAND2X0 U6702 ( .IN1(n5291), .IN2(n8289), .QN(n5943) );
  INVX0 U6703 ( .INP(n5944), .ZN(n442) );
  NOR2X0 U6704 ( .IN1(n5945), .IN2(n5946), .QN(n5944) );
  NAND2X0 U6705 ( .IN1(n5947), .IN2(n5948), .QN(n5946) );
  NAND2X0 U6706 ( .IN1(DATA_0_26), .IN2(n2153), .QN(n5948) );
  NAND2X0 U6707 ( .IN1(n2152), .IN2(CRC_OUT_1_26), .QN(n5947) );
  NAND2X0 U6708 ( .IN1(n5949), .IN2(n5950), .QN(n5945) );
  NAND2X0 U6709 ( .IN1(n4737), .IN2(n5951), .QN(n5950) );
  NAND2X0 U6710 ( .IN1(n443), .IN2(n4809), .QN(n5949) );
  INVX0 U6711 ( .INP(n5952), .ZN(n443) );
  NAND2X0 U6712 ( .IN1(n5291), .IN2(n8290), .QN(n5952) );
  INVX0 U6713 ( .INP(n5953), .ZN(n440) );
  NOR2X0 U6714 ( .IN1(n5954), .IN2(n5955), .QN(n5953) );
  NAND2X0 U6715 ( .IN1(n5956), .IN2(n5957), .QN(n5955) );
  NAND2X0 U6716 ( .IN1(DATA_0_27), .IN2(n2153), .QN(n5957) );
  NAND2X0 U6717 ( .IN1(n2152), .IN2(CRC_OUT_1_27), .QN(n5956) );
  NAND2X0 U6718 ( .IN1(n5958), .IN2(n5959), .QN(n5954) );
  NAND2X0 U6719 ( .IN1(n4737), .IN2(n5960), .QN(n5959) );
  NAND2X0 U6720 ( .IN1(n441), .IN2(n4809), .QN(n5958) );
  INVX0 U6721 ( .INP(n5961), .ZN(n441) );
  NAND2X0 U6722 ( .IN1(test_so89), .IN2(n5322), .QN(n5961) );
  INVX0 U6723 ( .INP(n5962), .ZN(n438) );
  NOR2X0 U6724 ( .IN1(n5963), .IN2(n5964), .QN(n5962) );
  NAND2X0 U6725 ( .IN1(n5965), .IN2(n5966), .QN(n5964) );
  NAND2X0 U6726 ( .IN1(DATA_0_28), .IN2(n2153), .QN(n5966) );
  NAND2X0 U6727 ( .IN1(n2152), .IN2(CRC_OUT_1_28), .QN(n5965) );
  NAND2X0 U6728 ( .IN1(n5967), .IN2(n5968), .QN(n5963) );
  NAND2X0 U6729 ( .IN1(n4738), .IN2(n5969), .QN(n5968) );
  NAND2X0 U6730 ( .IN1(n439), .IN2(n4809), .QN(n5967) );
  INVX0 U6731 ( .INP(n5970), .ZN(n439) );
  NAND2X0 U6732 ( .IN1(n5290), .IN2(n8293), .QN(n5970) );
  INVX0 U6733 ( .INP(n5971), .ZN(n436) );
  NOR2X0 U6734 ( .IN1(n5972), .IN2(n5973), .QN(n5971) );
  NAND2X0 U6735 ( .IN1(n5974), .IN2(n5975), .QN(n5973) );
  NAND2X0 U6736 ( .IN1(DATA_0_29), .IN2(n2153), .QN(n5975) );
  NAND2X0 U6737 ( .IN1(n2152), .IN2(CRC_OUT_1_29), .QN(n5974) );
  NAND2X0 U6738 ( .IN1(n5976), .IN2(n5977), .QN(n5972) );
  NAND2X0 U6739 ( .IN1(n4738), .IN2(n5978), .QN(n5977) );
  NAND2X0 U6740 ( .IN1(n437), .IN2(n4809), .QN(n5976) );
  INVX0 U6741 ( .INP(n5979), .ZN(n437) );
  NAND2X0 U6742 ( .IN1(n5290), .IN2(n8294), .QN(n5979) );
  INVX0 U6743 ( .INP(n5980), .ZN(n434) );
  NOR2X0 U6744 ( .IN1(n5981), .IN2(n5982), .QN(n5980) );
  NAND2X0 U6745 ( .IN1(n5983), .IN2(n5984), .QN(n5982) );
  NAND2X0 U6746 ( .IN1(DATA_0_30), .IN2(n2153), .QN(n5984) );
  NAND2X0 U6747 ( .IN1(n2152), .IN2(CRC_OUT_1_30), .QN(n5983) );
  NAND2X0 U6748 ( .IN1(n5985), .IN2(n5986), .QN(n5981) );
  NAND2X0 U6749 ( .IN1(n4738), .IN2(n5987), .QN(n5986) );
  NAND2X0 U6750 ( .IN1(n435), .IN2(n4809), .QN(n5985) );
  INVX0 U6751 ( .INP(n5988), .ZN(n435) );
  NAND2X0 U6752 ( .IN1(n5290), .IN2(n8295), .QN(n5988) );
  INVX0 U6753 ( .INP(n5989), .ZN(n432) );
  NOR2X0 U6754 ( .IN1(n5990), .IN2(n5991), .QN(n5989) );
  NAND2X0 U6755 ( .IN1(n5992), .IN2(n5993), .QN(n5991) );
  NAND2X0 U6756 ( .IN1(test_so100), .IN2(n2152), .QN(n5993) );
  NAND2X0 U6757 ( .IN1(n2245), .IN2(WX10829), .QN(n5992) );
  NAND2X0 U6758 ( .IN1(n5994), .IN2(n5995), .QN(n5990) );
  NAND2X0 U6759 ( .IN1(n4738), .IN2(n5996), .QN(n5995) );
  NAND2X0 U6760 ( .IN1(DATA_0_31), .IN2(n2153), .QN(n5994) );
  INVX0 U6761 ( .INP(n5997), .ZN(n413) );
  INVX0 U6762 ( .INP(n5998), .ZN(n412) );
  INVX0 U6763 ( .INP(n5999), .ZN(n411) );
  INVX0 U6764 ( .INP(n6000), .ZN(n410) );
  INVX0 U6765 ( .INP(n6001), .ZN(n409) );
  INVX0 U6766 ( .INP(n6002), .ZN(n408) );
  INVX0 U6767 ( .INP(n6003), .ZN(n407) );
  INVX0 U6768 ( .INP(n6004), .ZN(n406) );
  INVX0 U6769 ( .INP(n6005), .ZN(n405) );
  INVX0 U6770 ( .INP(n6006), .ZN(n404) );
  INVX0 U6771 ( .INP(n6007), .ZN(n403) );
  INVX0 U6772 ( .INP(n6008), .ZN(n402) );
  INVX0 U6773 ( .INP(n6009), .ZN(n401) );
  INVX0 U6774 ( .INP(n6010), .ZN(n400) );
  NAND2X0 U6775 ( .IN1(n6011), .IN2(n6012), .QN(n4) );
  NOR2X0 U6776 ( .IN1(n6013), .IN2(n6014), .QN(n6012) );
  NOR2X0 U6777 ( .IN1(n6015), .IN2(n4723), .QN(n6014) );
  NOR2X0 U6778 ( .IN1(n4765), .IN2(DFF_188_n1), .QN(n6013) );
  NOR2X0 U6779 ( .IN1(n6018), .IN2(n6019), .QN(n6011) );
  NOR2X0 U6780 ( .IN1(n6020), .IN2(n4778), .QN(n6019) );
  NOR2X0 U6781 ( .IN1(n6022), .IN2(n6023), .QN(n6018) );
  INVX0 U6782 ( .INP(WX488), .ZN(n6022) );
  INVX0 U6783 ( .INP(n6024), .ZN(n399) );
  INVX0 U6784 ( .INP(n6025), .ZN(n398) );
  INVX0 U6785 ( .INP(n6026), .ZN(n397) );
  INVX0 U6786 ( .INP(n6027), .ZN(n396) );
  INVX0 U6787 ( .INP(n6028), .ZN(n395) );
  INVX0 U6788 ( .INP(n6029), .ZN(n394) );
  INVX0 U6789 ( .INP(n6030), .ZN(n393) );
  INVX0 U6790 ( .INP(n6031), .ZN(n392) );
  INVX0 U6791 ( .INP(n6032), .ZN(n391) );
  INVX0 U6792 ( .INP(n6033), .ZN(n390) );
  INVX0 U6793 ( .INP(n6034), .ZN(n389) );
  INVX0 U6794 ( .INP(n6035), .ZN(n388) );
  INVX0 U6795 ( .INP(n6036), .ZN(n387) );
  INVX0 U6796 ( .INP(n6037), .ZN(n386) );
  INVX0 U6797 ( .INP(n6038), .ZN(n385) );
  INVX0 U6798 ( .INP(n6039), .ZN(n384) );
  INVX0 U6799 ( .INP(n6040), .ZN(n383) );
  INVX0 U6800 ( .INP(n6041), .ZN(n363) );
  INVX0 U6801 ( .INP(n6042), .ZN(n362) );
  INVX0 U6802 ( .INP(n6043), .ZN(n361) );
  INVX0 U6803 ( .INP(n6044), .ZN(n360) );
  INVX0 U6804 ( .INP(n6045), .ZN(n359) );
  INVX0 U6805 ( .INP(n6046), .ZN(n358) );
  INVX0 U6806 ( .INP(n6047), .ZN(n357) );
  INVX0 U6807 ( .INP(n6048), .ZN(n356) );
  INVX0 U6808 ( .INP(n6049), .ZN(n355) );
  INVX0 U6809 ( .INP(n6050), .ZN(n354) );
  INVX0 U6810 ( .INP(n6051), .ZN(n353) );
  INVX0 U6811 ( .INP(n6052), .ZN(n352) );
  INVX0 U6812 ( .INP(n6053), .ZN(n351) );
  INVX0 U6813 ( .INP(n6054), .ZN(n350) );
  INVX0 U6814 ( .INP(n6055), .ZN(n349) );
  INVX0 U6815 ( .INP(n6056), .ZN(n348) );
  INVX0 U6816 ( .INP(n6057), .ZN(n347) );
  INVX0 U6817 ( .INP(n6058), .ZN(n346) );
  INVX0 U6818 ( .INP(n6059), .ZN(n345) );
  INVX0 U6819 ( .INP(n6060), .ZN(n344) );
  INVX0 U6820 ( .INP(n6061), .ZN(n343) );
  INVX0 U6821 ( .INP(n6062), .ZN(n342) );
  INVX0 U6822 ( .INP(n6063), .ZN(n341) );
  INVX0 U6823 ( .INP(n6064), .ZN(n340) );
  INVX0 U6824 ( .INP(n6065), .ZN(n339) );
  INVX0 U6825 ( .INP(n6066), .ZN(n338) );
  INVX0 U6826 ( .INP(n6067), .ZN(n337) );
  INVX0 U6827 ( .INP(n6068), .ZN(n336) );
  INVX0 U6828 ( .INP(n6069), .ZN(n335) );
  INVX0 U6829 ( .INP(n6070), .ZN(n334) );
  NOR2X0 U6830 ( .IN1(n5259), .IN2(n5343), .QN(n3278) );
  INVX0 U6831 ( .INP(n6071), .ZN(n314) );
  INVX0 U6832 ( .INP(n6072), .ZN(n313) );
  INVX0 U6833 ( .INP(n6073), .ZN(n312) );
  INVX0 U6834 ( .INP(n6074), .ZN(n311) );
  INVX0 U6835 ( .INP(n6075), .ZN(n310) );
  INVX0 U6836 ( .INP(n6076), .ZN(n309) );
  INVX0 U6837 ( .INP(n6077), .ZN(n308) );
  INVX0 U6838 ( .INP(n6078), .ZN(n307) );
  INVX0 U6839 ( .INP(n6079), .ZN(n306) );
  INVX0 U6840 ( .INP(n6080), .ZN(n305) );
  INVX0 U6841 ( .INP(n6081), .ZN(n304) );
  INVX0 U6842 ( .INP(n6082), .ZN(n303) );
  INVX0 U6843 ( .INP(n6083), .ZN(n302) );
  INVX0 U6844 ( .INP(n6084), .ZN(n301) );
  INVX0 U6845 ( .INP(n6085), .ZN(n300) );
  INVX0 U6846 ( .INP(n6086), .ZN(n3) );
  NOR2X0 U6847 ( .IN1(n6087), .IN2(n6088), .QN(n6086) );
  NAND2X0 U6848 ( .IN1(n6089), .IN2(n6090), .QN(n6088) );
  NAND2X0 U6849 ( .IN1(n4739), .IN2(n6091), .QN(n6090) );
  NAND2X0 U6850 ( .IN1(n2152), .IN2(CRC_OUT_9_29), .QN(n6089) );
  NAND2X0 U6851 ( .IN1(n6092), .IN2(n6093), .QN(n6087) );
  NAND2X0 U6852 ( .IN1(n2153), .IN2(n6094), .QN(n6093) );
  NAND2X0 U6853 ( .IN1(WX486), .IN2(n4809), .QN(n6092) );
  INVX0 U6854 ( .INP(n6095), .ZN(n299) );
  INVX0 U6855 ( .INP(n6096), .ZN(n298) );
  INVX0 U6856 ( .INP(n6097), .ZN(n297) );
  INVX0 U6857 ( .INP(n6098), .ZN(n296) );
  INVX0 U6858 ( .INP(n6099), .ZN(n295) );
  INVX0 U6859 ( .INP(n6100), .ZN(n294) );
  INVX0 U6860 ( .INP(n6101), .ZN(n293) );
  INVX0 U6861 ( .INP(n6102), .ZN(n292) );
  INVX0 U6862 ( .INP(n6103), .ZN(n291) );
  INVX0 U6863 ( .INP(n6104), .ZN(n290) );
  INVX0 U6864 ( .INP(n6105), .ZN(n289) );
  INVX0 U6865 ( .INP(n6106), .ZN(n288) );
  INVX0 U6866 ( .INP(n6107), .ZN(n287) );
  INVX0 U6867 ( .INP(n6108), .ZN(n286) );
  INVX0 U6868 ( .INP(n6109), .ZN(n285) );
  INVX0 U6869 ( .INP(n6110), .ZN(n28) );
  NOR2X0 U6870 ( .IN1(n6111), .IN2(n6112), .QN(n6110) );
  NAND2X0 U6871 ( .IN1(n6113), .IN2(n6114), .QN(n6112) );
  NAND2X0 U6872 ( .IN1(n4738), .IN2(n6115), .QN(n6114) );
  NAND2X0 U6873 ( .IN1(n2152), .IN2(CRC_OUT_9_0), .QN(n6113) );
  NAND2X0 U6874 ( .IN1(n6116), .IN2(n6117), .QN(n6111) );
  NAND2X0 U6875 ( .IN1(n6118), .IN2(n2153), .QN(n6117) );
  INVX0 U6876 ( .INP(n6119), .ZN(n6118) );
  NAND2X0 U6877 ( .IN1(WX544), .IN2(n4809), .QN(n6116) );
  INVX0 U6878 ( .INP(n6120), .ZN(n27) );
  NOR2X0 U6879 ( .IN1(n6121), .IN2(n6122), .QN(n6120) );
  NAND2X0 U6880 ( .IN1(n6123), .IN2(n6124), .QN(n6122) );
  NAND2X0 U6881 ( .IN1(n4739), .IN2(n6125), .QN(n6124) );
  NAND2X0 U6882 ( .IN1(test_so9), .IN2(n2152), .QN(n6123) );
  NAND2X0 U6883 ( .IN1(n6126), .IN2(n6127), .QN(n6121) );
  NAND2X0 U6884 ( .IN1(n2153), .IN2(n6128), .QN(n6127) );
  NAND2X0 U6885 ( .IN1(WX542), .IN2(n4809), .QN(n6126) );
  INVX0 U6886 ( .INP(n6129), .ZN(n265) );
  INVX0 U6887 ( .INP(n6130), .ZN(n264) );
  INVX0 U6888 ( .INP(n6131), .ZN(n263) );
  INVX0 U6889 ( .INP(n6132), .ZN(n262) );
  INVX0 U6890 ( .INP(n6133), .ZN(n261) );
  INVX0 U6891 ( .INP(n6134), .ZN(n260) );
  NAND2X0 U6892 ( .IN1(n6135), .IN2(n6136), .QN(n26) );
  NOR2X0 U6893 ( .IN1(n6137), .IN2(n6138), .QN(n6136) );
  NOR2X0 U6894 ( .IN1(n6139), .IN2(n4723), .QN(n6138) );
  NOR2X0 U6895 ( .IN1(n4765), .IN2(DFF_162_n1), .QN(n6137) );
  NOR2X0 U6896 ( .IN1(n6140), .IN2(n6141), .QN(n6135) );
  NOR2X0 U6897 ( .IN1(n4785), .IN2(n6142), .QN(n6141) );
  NOR2X0 U6898 ( .IN1(n6143), .IN2(n6023), .QN(n6140) );
  INVX0 U6899 ( .INP(WX540), .ZN(n6143) );
  INVX0 U6900 ( .INP(n6144), .ZN(n259) );
  INVX0 U6901 ( .INP(n6145), .ZN(n258) );
  INVX0 U6902 ( .INP(n6146), .ZN(n257) );
  INVX0 U6903 ( .INP(n6147), .ZN(n256) );
  INVX0 U6904 ( .INP(n6148), .ZN(n255) );
  INVX0 U6905 ( .INP(n6149), .ZN(n254) );
  INVX0 U6906 ( .INP(n6150), .ZN(n253) );
  INVX0 U6907 ( .INP(n6151), .ZN(n252) );
  INVX0 U6908 ( .INP(n6152), .ZN(n251) );
  INVX0 U6909 ( .INP(n6153), .ZN(n250) );
  INVX0 U6910 ( .INP(n6154), .ZN(n25) );
  NOR2X0 U6911 ( .IN1(n6155), .IN2(n6156), .QN(n6154) );
  NAND2X0 U6912 ( .IN1(n6157), .IN2(n6158), .QN(n6156) );
  NAND2X0 U6913 ( .IN1(n4739), .IN2(n6159), .QN(n6158) );
  NAND2X0 U6914 ( .IN1(n2152), .IN2(CRC_OUT_9_3), .QN(n6157) );
  NAND2X0 U6915 ( .IN1(n6160), .IN2(n6161), .QN(n6155) );
  NAND2X0 U6916 ( .IN1(n2153), .IN2(n6162), .QN(n6161) );
  NAND2X0 U6917 ( .IN1(WX538), .IN2(n4809), .QN(n6160) );
  INVX0 U6918 ( .INP(n6163), .ZN(n249) );
  INVX0 U6919 ( .INP(n6164), .ZN(n248) );
  INVX0 U6920 ( .INP(n6165), .ZN(n247) );
  INVX0 U6921 ( .INP(n6166), .ZN(n246) );
  INVX0 U6922 ( .INP(n6167), .ZN(n245) );
  INVX0 U6923 ( .INP(n6168), .ZN(n244) );
  INVX0 U6924 ( .INP(n6169), .ZN(n243) );
  INVX0 U6925 ( .INP(n6170), .ZN(n242) );
  INVX0 U6926 ( .INP(n6171), .ZN(n241) );
  INVX0 U6927 ( .INP(n6172), .ZN(n240) );
  INVX0 U6928 ( .INP(n6173), .ZN(n24) );
  NOR2X0 U6929 ( .IN1(n6174), .IN2(n6175), .QN(n6173) );
  NAND2X0 U6930 ( .IN1(n6176), .IN2(n6177), .QN(n6175) );
  NAND2X0 U6931 ( .IN1(n4739), .IN2(n6178), .QN(n6177) );
  NAND2X0 U6932 ( .IN1(n2152), .IN2(CRC_OUT_9_4), .QN(n6176) );
  NAND2X0 U6933 ( .IN1(n6179), .IN2(n6180), .QN(n6174) );
  NAND2X0 U6934 ( .IN1(n6181), .IN2(n2153), .QN(n6180) );
  INVX0 U6935 ( .INP(n6182), .ZN(n6181) );
  NAND2X0 U6936 ( .IN1(WX536), .IN2(n4808), .QN(n6179) );
  INVX0 U6937 ( .INP(n6183), .ZN(n239) );
  INVX0 U6938 ( .INP(n6184), .ZN(n238) );
  INVX0 U6939 ( .INP(n6185), .ZN(n237) );
  INVX0 U6940 ( .INP(n6186), .ZN(n236) );
  INVX0 U6941 ( .INP(n6187), .ZN(n235) );
  INVX0 U6942 ( .INP(n6188), .ZN(n23) );
  NOR2X0 U6943 ( .IN1(n6189), .IN2(n6190), .QN(n6188) );
  NAND2X0 U6944 ( .IN1(n6191), .IN2(n6192), .QN(n6190) );
  NAND2X0 U6945 ( .IN1(n4738), .IN2(n6193), .QN(n6192) );
  NAND2X0 U6946 ( .IN1(n2152), .IN2(CRC_OUT_9_5), .QN(n6191) );
  NAND2X0 U6947 ( .IN1(n6194), .IN2(n6195), .QN(n6189) );
  NAND2X0 U6948 ( .IN1(n2153), .IN2(n6196), .QN(n6195) );
  NAND2X0 U6949 ( .IN1(WX534), .IN2(n4808), .QN(n6194) );
  NAND2X0 U6950 ( .IN1(n6197), .IN2(n6198), .QN(n22) );
  NOR2X0 U6951 ( .IN1(n6199), .IN2(n6200), .QN(n6198) );
  NOR2X0 U6952 ( .IN1(n6201), .IN2(n4723), .QN(n6200) );
  NOR2X0 U6953 ( .IN1(n4765), .IN2(DFF_166_n1), .QN(n6199) );
  NOR2X0 U6954 ( .IN1(n6202), .IN2(n6203), .QN(n6197) );
  NOR2X0 U6955 ( .IN1(n4785), .IN2(n6204), .QN(n6203) );
  NOR2X0 U6956 ( .IN1(n6205), .IN2(n6023), .QN(n6202) );
  INVX0 U6957 ( .INP(WX532), .ZN(n6205) );
  INVX0 U6958 ( .INP(n6206), .ZN(n215) );
  INVX0 U6959 ( .INP(n6207), .ZN(n214) );
  INVX0 U6960 ( .INP(n6208), .ZN(n213) );
  INVX0 U6961 ( .INP(n6209), .ZN(n212) );
  INVX0 U6962 ( .INP(n6210), .ZN(n211) );
  INVX0 U6963 ( .INP(n6211), .ZN(n210) );
  INVX0 U6964 ( .INP(n6212), .ZN(n21) );
  NOR2X0 U6965 ( .IN1(n6213), .IN2(n6214), .QN(n6212) );
  NAND2X0 U6966 ( .IN1(n6215), .IN2(n6216), .QN(n6214) );
  NAND2X0 U6967 ( .IN1(n4739), .IN2(n6217), .QN(n6216) );
  NAND2X0 U6968 ( .IN1(n2152), .IN2(CRC_OUT_9_7), .QN(n6215) );
  NAND2X0 U6969 ( .IN1(n6218), .IN2(n6219), .QN(n6213) );
  NAND2X0 U6970 ( .IN1(n2153), .IN2(n6220), .QN(n6219) );
  NAND2X0 U6971 ( .IN1(WX530), .IN2(n4808), .QN(n6218) );
  INVX0 U6972 ( .INP(n6221), .ZN(n209) );
  INVX0 U6973 ( .INP(n6222), .ZN(n208) );
  INVX0 U6974 ( .INP(n6223), .ZN(n207) );
  INVX0 U6975 ( .INP(n6224), .ZN(n206) );
  INVX0 U6976 ( .INP(n6225), .ZN(n205) );
  INVX0 U6977 ( .INP(n6226), .ZN(n204) );
  INVX0 U6978 ( .INP(n6227), .ZN(n203) );
  INVX0 U6979 ( .INP(n6228), .ZN(n202) );
  INVX0 U6980 ( .INP(n6229), .ZN(n201) );
  INVX0 U6981 ( .INP(n6230), .ZN(n200) );
  INVX0 U6982 ( .INP(n6231), .ZN(n20) );
  NOR2X0 U6983 ( .IN1(n6232), .IN2(n6233), .QN(n6231) );
  NAND2X0 U6984 ( .IN1(n6234), .IN2(n6235), .QN(n6233) );
  NAND2X0 U6985 ( .IN1(n4739), .IN2(n6236), .QN(n6235) );
  NAND2X0 U6986 ( .IN1(n2152), .IN2(CRC_OUT_9_8), .QN(n6234) );
  NAND2X0 U6987 ( .IN1(n6237), .IN2(n6238), .QN(n6232) );
  NAND2X0 U6988 ( .IN1(n2153), .IN2(n6239), .QN(n6238) );
  NAND2X0 U6989 ( .IN1(WX528), .IN2(n4808), .QN(n6237) );
  INVX0 U6990 ( .INP(n6240), .ZN(n2) );
  NOR2X0 U6991 ( .IN1(n6241), .IN2(n6242), .QN(n6240) );
  NAND2X0 U6992 ( .IN1(n6243), .IN2(n6244), .QN(n6242) );
  NAND2X0 U6993 ( .IN1(n4739), .IN2(n6245), .QN(n6244) );
  NAND2X0 U6994 ( .IN1(n2152), .IN2(CRC_OUT_9_30), .QN(n6243) );
  NAND2X0 U6995 ( .IN1(n6246), .IN2(n6247), .QN(n6241) );
  NAND2X0 U6996 ( .IN1(n2153), .IN2(n6248), .QN(n6247) );
  NAND2X0 U6997 ( .IN1(WX484), .IN2(n4808), .QN(n6246) );
  INVX0 U6998 ( .INP(n6249), .ZN(n199) );
  INVX0 U6999 ( .INP(n6250), .ZN(n198) );
  INVX0 U7000 ( .INP(n6251), .ZN(n197) );
  INVX0 U7001 ( .INP(n6252), .ZN(n196) );
  INVX0 U7002 ( .INP(n6253), .ZN(n195) );
  INVX0 U7003 ( .INP(n6254), .ZN(n194) );
  INVX0 U7004 ( .INP(n6255), .ZN(n193) );
  INVX0 U7005 ( .INP(n6256), .ZN(n192) );
  INVX0 U7006 ( .INP(n6257), .ZN(n191) );
  INVX0 U7007 ( .INP(n6258), .ZN(n190) );
  INVX0 U7008 ( .INP(n6259), .ZN(n19) );
  NOR2X0 U7009 ( .IN1(n6260), .IN2(n6261), .QN(n6259) );
  NAND2X0 U7010 ( .IN1(n6262), .IN2(n6263), .QN(n6261) );
  NAND2X0 U7011 ( .IN1(n4738), .IN2(n6264), .QN(n6263) );
  NAND2X0 U7012 ( .IN1(n2152), .IN2(CRC_OUT_9_9), .QN(n6262) );
  NAND2X0 U7013 ( .IN1(n6265), .IN2(n6266), .QN(n6260) );
  NAND2X0 U7014 ( .IN1(n2153), .IN2(n6267), .QN(n6266) );
  NAND2X0 U7015 ( .IN1(WX526), .IN2(n4808), .QN(n6265) );
  INVX0 U7016 ( .INP(n6268), .ZN(n189) );
  INVX0 U7017 ( .INP(n6269), .ZN(n188) );
  INVX0 U7018 ( .INP(n6270), .ZN(n187) );
  INVX0 U7019 ( .INP(n6271), .ZN(n186) );
  INVX0 U7020 ( .INP(n6272), .ZN(n185) );
  INVX0 U7021 ( .INP(n6273), .ZN(n18) );
  NOR2X0 U7022 ( .IN1(n6274), .IN2(n6275), .QN(n6273) );
  NAND2X0 U7023 ( .IN1(n6276), .IN2(n6277), .QN(n6275) );
  NAND2X0 U7024 ( .IN1(n4738), .IN2(n6278), .QN(n6277) );
  NAND2X0 U7025 ( .IN1(n2152), .IN2(CRC_OUT_9_11), .QN(n6276) );
  NAND2X0 U7026 ( .IN1(n6279), .IN2(n6280), .QN(n6274) );
  NAND2X0 U7027 ( .IN1(n2153), .IN2(n6281), .QN(n6280) );
  NAND2X0 U7028 ( .IN1(WX522), .IN2(n4808), .QN(n6279) );
  INVX0 U7029 ( .INP(n6282), .ZN(n17) );
  NOR2X0 U7030 ( .IN1(n6283), .IN2(n6284), .QN(n6282) );
  NAND2X0 U7031 ( .IN1(n6285), .IN2(n6286), .QN(n6284) );
  NAND2X0 U7032 ( .IN1(n4739), .IN2(n6287), .QN(n6286) );
  NAND2X0 U7033 ( .IN1(n2152), .IN2(CRC_OUT_9_12), .QN(n6285) );
  NAND2X0 U7034 ( .IN1(n6288), .IN2(n6289), .QN(n6283) );
  NAND2X0 U7035 ( .IN1(n2153), .IN2(n6290), .QN(n6289) );
  NAND2X0 U7036 ( .IN1(WX520), .IN2(n4808), .QN(n6288) );
  INVX0 U7037 ( .INP(n6291), .ZN(n165) );
  INVX0 U7038 ( .INP(n6292), .ZN(n164) );
  INVX0 U7039 ( .INP(n6293), .ZN(n163) );
  INVX0 U7040 ( .INP(n6294), .ZN(n162) );
  INVX0 U7041 ( .INP(n6295), .ZN(n161) );
  INVX0 U7042 ( .INP(n6296), .ZN(n160) );
  INVX0 U7043 ( .INP(n6297), .ZN(n16) );
  NOR2X0 U7044 ( .IN1(n6298), .IN2(n6299), .QN(n6297) );
  NAND2X0 U7045 ( .IN1(n6300), .IN2(n6301), .QN(n6299) );
  NAND2X0 U7046 ( .IN1(n4740), .IN2(n6302), .QN(n6301) );
  NAND2X0 U7047 ( .IN1(n2152), .IN2(CRC_OUT_9_13), .QN(n6300) );
  NAND2X0 U7048 ( .IN1(n6303), .IN2(n6304), .QN(n6298) );
  NAND2X0 U7049 ( .IN1(n2153), .IN2(n6305), .QN(n6304) );
  NAND2X0 U7050 ( .IN1(WX518), .IN2(n4808), .QN(n6303) );
  INVX0 U7051 ( .INP(n6306), .ZN(n159) );
  INVX0 U7052 ( .INP(n6307), .ZN(n158) );
  INVX0 U7053 ( .INP(n6308), .ZN(n157) );
  INVX0 U7054 ( .INP(n6309), .ZN(n156) );
  INVX0 U7055 ( .INP(n6310), .ZN(n155) );
  INVX0 U7056 ( .INP(n6311), .ZN(n154) );
  INVX0 U7057 ( .INP(n6312), .ZN(n153) );
  INVX0 U7058 ( .INP(n6313), .ZN(n152) );
  INVX0 U7059 ( .INP(n6314), .ZN(n151) );
  INVX0 U7060 ( .INP(n6315), .ZN(n150) );
  INVX0 U7061 ( .INP(n6316), .ZN(n15) );
  NOR2X0 U7062 ( .IN1(n6317), .IN2(n6318), .QN(n6316) );
  NAND2X0 U7063 ( .IN1(n6319), .IN2(n6320), .QN(n6318) );
  NAND2X0 U7064 ( .IN1(n4739), .IN2(n6321), .QN(n6320) );
  NAND2X0 U7065 ( .IN1(n2152), .IN2(CRC_OUT_9_14), .QN(n6319) );
  NAND2X0 U7066 ( .IN1(n6322), .IN2(n6323), .QN(n6317) );
  NAND2X0 U7067 ( .IN1(n6324), .IN2(n2153), .QN(n6323) );
  INVX0 U7068 ( .INP(n6325), .ZN(n6324) );
  NAND2X0 U7069 ( .IN1(WX516), .IN2(n4808), .QN(n6322) );
  INVX0 U7070 ( .INP(n6326), .ZN(n149) );
  INVX0 U7071 ( .INP(n6327), .ZN(n147) );
  INVX0 U7072 ( .INP(n6328), .ZN(n146) );
  INVX0 U7073 ( .INP(n6329), .ZN(n145) );
  INVX0 U7074 ( .INP(n6330), .ZN(n144) );
  INVX0 U7075 ( .INP(n6331), .ZN(n143) );
  INVX0 U7076 ( .INP(n6332), .ZN(n142) );
  INVX0 U7077 ( .INP(n6333), .ZN(n141) );
  INVX0 U7078 ( .INP(n6334), .ZN(n140) );
  INVX0 U7079 ( .INP(n6335), .ZN(n14) );
  NOR2X0 U7080 ( .IN1(n6336), .IN2(n6337), .QN(n6335) );
  NAND2X0 U7081 ( .IN1(n6338), .IN2(n6339), .QN(n6337) );
  NAND2X0 U7082 ( .IN1(n4740), .IN2(n6340), .QN(n6339) );
  NAND2X0 U7083 ( .IN1(n2152), .IN2(CRC_OUT_9_15), .QN(n6338) );
  NAND2X0 U7084 ( .IN1(n6341), .IN2(n6342), .QN(n6336) );
  NAND2X0 U7085 ( .IN1(n2153), .IN2(n6343), .QN(n6342) );
  NAND2X0 U7086 ( .IN1(WX514), .IN2(n4807), .QN(n6341) );
  INVX0 U7087 ( .INP(n6344), .ZN(n139) );
  INVX0 U7088 ( .INP(n6345), .ZN(n138) );
  INVX0 U7089 ( .INP(n6346), .ZN(n137) );
  INVX0 U7090 ( .INP(n6347), .ZN(n136) );
  INVX0 U7091 ( .INP(n6348), .ZN(n135) );
  INVX0 U7092 ( .INP(n6349), .ZN(n134) );
  INVX0 U7093 ( .INP(n6350), .ZN(n133) );
  INVX0 U7094 ( .INP(n6351), .ZN(n132) );
  INVX0 U7095 ( .INP(n6352), .ZN(n13) );
  NOR2X0 U7096 ( .IN1(n6353), .IN2(n6354), .QN(n6352) );
  NAND2X0 U7097 ( .IN1(n6355), .IN2(n6356), .QN(n6354) );
  NAND2X0 U7098 ( .IN1(n4740), .IN2(n6357), .QN(n6356) );
  NAND2X0 U7099 ( .IN1(n2152), .IN2(CRC_OUT_9_17), .QN(n6355) );
  NAND2X0 U7100 ( .IN1(n6358), .IN2(n6359), .QN(n6353) );
  NAND2X0 U7101 ( .IN1(n2153), .IN2(n6360), .QN(n6359) );
  NAND2X0 U7102 ( .IN1(WX510), .IN2(n4807), .QN(n6358) );
  INVX0 U7103 ( .INP(n6361), .ZN(n12) );
  NOR2X0 U7104 ( .IN1(n6362), .IN2(n6363), .QN(n6361) );
  NAND2X0 U7105 ( .IN1(n6364), .IN2(n6365), .QN(n6363) );
  NAND2X0 U7106 ( .IN1(n4740), .IN2(n6366), .QN(n6365) );
  NAND2X0 U7107 ( .IN1(n2152), .IN2(CRC_OUT_9_18), .QN(n6364) );
  NAND2X0 U7108 ( .IN1(n6367), .IN2(n6368), .QN(n6362) );
  NAND2X0 U7109 ( .IN1(n6369), .IN2(n2153), .QN(n6368) );
  INVX0 U7110 ( .INP(n6370), .ZN(n6369) );
  NAND2X0 U7111 ( .IN1(WX508), .IN2(n4807), .QN(n6367) );
  INVX0 U7112 ( .INP(n6371), .ZN(n11) );
  NOR2X0 U7113 ( .IN1(n6372), .IN2(n6373), .QN(n6371) );
  NAND2X0 U7114 ( .IN1(n6374), .IN2(n6375), .QN(n6373) );
  NAND2X0 U7115 ( .IN1(n4740), .IN2(n6376), .QN(n6375) );
  NAND2X0 U7116 ( .IN1(test_so10), .IN2(n2152), .QN(n6374) );
  NAND2X0 U7117 ( .IN1(n6377), .IN2(n6378), .QN(n6372) );
  NAND2X0 U7118 ( .IN1(n2153), .IN2(n6379), .QN(n6378) );
  NAND2X0 U7119 ( .IN1(WX506), .IN2(n4807), .QN(n6377) );
  INVX0 U7120 ( .INP(n6380), .ZN(n10) );
  NOR2X0 U7121 ( .IN1(n6381), .IN2(n6382), .QN(n6380) );
  NAND2X0 U7122 ( .IN1(n6383), .IN2(n6384), .QN(n6382) );
  NAND2X0 U7123 ( .IN1(n4740), .IN2(n6385), .QN(n6384) );
  NAND2X0 U7124 ( .IN1(n2152), .IN2(CRC_OUT_9_21), .QN(n6383) );
  NAND2X0 U7125 ( .IN1(n6386), .IN2(n6387), .QN(n6381) );
  NAND2X0 U7126 ( .IN1(n2153), .IN2(n6388), .QN(n6387) );
  NAND2X0 U7127 ( .IN1(WX502), .IN2(n4807), .QN(n6386) );
  NOR2X0 U7128 ( .IN1(n9469), .IN2(n5343), .QN(WX9789) );
  NOR2X0 U7129 ( .IN1(n9472), .IN2(n5343), .QN(WX9787) );
  NOR2X0 U7130 ( .IN1(n9473), .IN2(n5343), .QN(WX9785) );
  NOR2X0 U7131 ( .IN1(n9476), .IN2(n5343), .QN(WX9783) );
  NOR2X0 U7132 ( .IN1(n5426), .IN2(n4706), .QN(WX9781) );
  NOR2X0 U7133 ( .IN1(n9477), .IN2(n5343), .QN(WX9779) );
  NOR2X0 U7134 ( .IN1(n9478), .IN2(n5343), .QN(WX9777) );
  NOR2X0 U7135 ( .IN1(n9479), .IN2(n5343), .QN(WX9775) );
  NOR2X0 U7136 ( .IN1(n9480), .IN2(n5343), .QN(WX9773) );
  NOR2X0 U7137 ( .IN1(n9481), .IN2(n5343), .QN(WX9771) );
  NOR2X0 U7138 ( .IN1(n9482), .IN2(n5343), .QN(WX9769) );
  NOR2X0 U7139 ( .IN1(n9483), .IN2(n5343), .QN(WX9767) );
  NOR2X0 U7140 ( .IN1(n9484), .IN2(n5344), .QN(WX9765) );
  NOR2X0 U7141 ( .IN1(n9485), .IN2(n5344), .QN(WX9763) );
  NOR2X0 U7142 ( .IN1(n9486), .IN2(n5344), .QN(WX9761) );
  NOR2X0 U7143 ( .IN1(n9487), .IN2(n5344), .QN(WX9759) );
  NAND2X0 U7144 ( .IN1(n6389), .IN2(n6390), .QN(WX9757) );
  NOR2X0 U7145 ( .IN1(n6391), .IN2(n6392), .QN(n6390) );
  NOR2X0 U7146 ( .IN1(n6393), .IN2(n4723), .QN(n6392) );
  NOR2X0 U7147 ( .IN1(n6394), .IN2(n4770), .QN(n6391) );
  INVX0 U7148 ( .INP(n5709), .ZN(n6394) );
  XNOR2X1 U7149 ( .IN1(n6395), .IN2(n6396), .Q(n5709) );
  XOR2X1 U7150 ( .IN1(n9695), .IN2(n4409), .Q(n6396) );
  XOR2X1 U7151 ( .IN1(WX11051), .IN2(n4146), .Q(n6395) );
  NOR2X0 U7152 ( .IN1(n6397), .IN2(n6398), .QN(n6389) );
  NOR2X0 U7153 ( .IN1(DFF_1504_n1), .IN2(n4755), .QN(n6398) );
  NOR2X0 U7154 ( .IN1(n4796), .IN2(n5997), .QN(n6397) );
  NAND2X0 U7155 ( .IN1(n5290), .IN2(n8321), .QN(n5997) );
  NAND2X0 U7156 ( .IN1(n6399), .IN2(n6400), .QN(WX9755) );
  NOR2X0 U7157 ( .IN1(n6401), .IN2(n6402), .QN(n6400) );
  NOR2X0 U7158 ( .IN1(n4732), .IN2(n6403), .QN(n6402) );
  NOR2X0 U7159 ( .IN1(n6404), .IN2(n4770), .QN(n6401) );
  INVX0 U7160 ( .INP(n5718), .ZN(n6404) );
  XNOR2X1 U7161 ( .IN1(n6405), .IN2(n6406), .Q(n5718) );
  XOR2X1 U7162 ( .IN1(n9696), .IN2(n4442), .Q(n6406) );
  XOR2X1 U7163 ( .IN1(WX11049), .IN2(n4148), .Q(n6405) );
  NOR2X0 U7164 ( .IN1(n6407), .IN2(n6408), .QN(n6399) );
  NOR2X0 U7165 ( .IN1(DFF_1505_n1), .IN2(n4755), .QN(n6408) );
  NOR2X0 U7166 ( .IN1(n4796), .IN2(n5998), .QN(n6407) );
  NAND2X0 U7167 ( .IN1(n5290), .IN2(n8322), .QN(n5998) );
  NAND2X0 U7168 ( .IN1(n6409), .IN2(n6410), .QN(WX9753) );
  NOR2X0 U7169 ( .IN1(n6411), .IN2(n6412), .QN(n6410) );
  NOR2X0 U7170 ( .IN1(n6413), .IN2(n4723), .QN(n6412) );
  NOR2X0 U7171 ( .IN1(n4785), .IN2(n5728), .QN(n6411) );
  XNOR2X1 U7172 ( .IN1(n6414), .IN2(n6415), .Q(n5728) );
  XOR2X1 U7173 ( .IN1(test_so98), .IN2(n9697), .Q(n6415) );
  XOR2X1 U7174 ( .IN1(WX11047), .IN2(n4150), .Q(n6414) );
  NOR2X0 U7175 ( .IN1(n6416), .IN2(n6417), .QN(n6409) );
  NOR2X0 U7176 ( .IN1(n4765), .IN2(n4713), .QN(n6417) );
  NOR2X0 U7177 ( .IN1(n4796), .IN2(n5999), .QN(n6416) );
  NAND2X0 U7178 ( .IN1(n5290), .IN2(n8323), .QN(n5999) );
  NAND2X0 U7179 ( .IN1(n6418), .IN2(n6419), .QN(WX9751) );
  NOR2X0 U7180 ( .IN1(n6420), .IN2(n6421), .QN(n6419) );
  NOR2X0 U7181 ( .IN1(n4732), .IN2(n6422), .QN(n6421) );
  NOR2X0 U7182 ( .IN1(n6423), .IN2(n4770), .QN(n6420) );
  INVX0 U7183 ( .INP(n5737), .ZN(n6423) );
  XNOR2X1 U7184 ( .IN1(n6424), .IN2(n6425), .Q(n5737) );
  XOR2X1 U7185 ( .IN1(n9698), .IN2(n4441), .Q(n6425) );
  XOR2X1 U7186 ( .IN1(WX11045), .IN2(n4152), .Q(n6424) );
  NOR2X0 U7187 ( .IN1(n6426), .IN2(n6427), .QN(n6418) );
  NOR2X0 U7188 ( .IN1(DFF_1507_n1), .IN2(n4755), .QN(n6427) );
  NOR2X0 U7189 ( .IN1(n4796), .IN2(n6000), .QN(n6426) );
  NAND2X0 U7190 ( .IN1(n5289), .IN2(n8324), .QN(n6000) );
  NAND2X0 U7191 ( .IN1(n6428), .IN2(n6429), .QN(WX9749) );
  NOR2X0 U7192 ( .IN1(n6430), .IN2(n6431), .QN(n6429) );
  NOR2X0 U7193 ( .IN1(n6432), .IN2(n4723), .QN(n6431) );
  NOR2X0 U7194 ( .IN1(n4785), .IN2(n5747), .QN(n6430) );
  XNOR2X1 U7195 ( .IN1(n6433), .IN2(n6434), .Q(n5747) );
  XOR2X1 U7196 ( .IN1(test_so96), .IN2(n9699), .Q(n6434) );
  XOR2X1 U7197 ( .IN1(WX11043), .IN2(n4390), .Q(n6433) );
  NOR2X0 U7198 ( .IN1(n6435), .IN2(n6436), .QN(n6428) );
  NOR2X0 U7199 ( .IN1(DFF_1508_n1), .IN2(n4755), .QN(n6436) );
  NOR2X0 U7200 ( .IN1(n4796), .IN2(n6001), .QN(n6435) );
  NAND2X0 U7201 ( .IN1(n5289), .IN2(n8325), .QN(n6001) );
  NAND2X0 U7202 ( .IN1(n6437), .IN2(n6438), .QN(WX9747) );
  NOR2X0 U7203 ( .IN1(n6439), .IN2(n6440), .QN(n6438) );
  NOR2X0 U7204 ( .IN1(n6441), .IN2(n4722), .QN(n6440) );
  NOR2X0 U7205 ( .IN1(n6442), .IN2(n4770), .QN(n6439) );
  INVX0 U7206 ( .INP(n5756), .ZN(n6442) );
  XNOR2X1 U7207 ( .IN1(n6443), .IN2(n6444), .Q(n5756) );
  XOR2X1 U7208 ( .IN1(n9700), .IN2(n4440), .Q(n6444) );
  XOR2X1 U7209 ( .IN1(WX11041), .IN2(n4155), .Q(n6443) );
  NOR2X0 U7210 ( .IN1(n6445), .IN2(n6446), .QN(n6437) );
  NOR2X0 U7211 ( .IN1(DFF_1509_n1), .IN2(n4755), .QN(n6446) );
  NOR2X0 U7212 ( .IN1(n4796), .IN2(n6002), .QN(n6445) );
  NAND2X0 U7213 ( .IN1(test_so79), .IN2(n5322), .QN(n6002) );
  NAND2X0 U7214 ( .IN1(n6447), .IN2(n6448), .QN(WX9745) );
  NOR2X0 U7215 ( .IN1(n6449), .IN2(n6450), .QN(n6448) );
  NOR2X0 U7216 ( .IN1(n6451), .IN2(n4722), .QN(n6450) );
  NOR2X0 U7217 ( .IN1(n4784), .IN2(n5766), .QN(n6449) );
  XNOR2X1 U7218 ( .IN1(n6452), .IN2(n6453), .Q(n5766) );
  XOR2X1 U7219 ( .IN1(test_so94), .IN2(n9701), .Q(n6453) );
  XOR2X1 U7220 ( .IN1(WX11039), .IN2(n4439), .Q(n6452) );
  NOR2X0 U7221 ( .IN1(n6454), .IN2(n6455), .QN(n6447) );
  NOR2X0 U7222 ( .IN1(DFF_1510_n1), .IN2(n4755), .QN(n6455) );
  NOR2X0 U7223 ( .IN1(n4796), .IN2(n6003), .QN(n6454) );
  NAND2X0 U7224 ( .IN1(n5289), .IN2(n8328), .QN(n6003) );
  NAND2X0 U7225 ( .IN1(n6456), .IN2(n6457), .QN(WX9743) );
  NOR2X0 U7226 ( .IN1(n6458), .IN2(n6459), .QN(n6457) );
  NOR2X0 U7227 ( .IN1(n6460), .IN2(n4722), .QN(n6459) );
  NOR2X0 U7228 ( .IN1(n6461), .IN2(n4770), .QN(n6458) );
  INVX0 U7229 ( .INP(n5775), .ZN(n6461) );
  XNOR2X1 U7230 ( .IN1(n6462), .IN2(n6463), .Q(n5775) );
  XOR2X1 U7231 ( .IN1(n9702), .IN2(n4438), .Q(n6463) );
  XOR2X1 U7232 ( .IN1(WX11037), .IN2(n4158), .Q(n6462) );
  NOR2X0 U7233 ( .IN1(n6464), .IN2(n6465), .QN(n6456) );
  NOR2X0 U7234 ( .IN1(DFF_1511_n1), .IN2(n4755), .QN(n6465) );
  NOR2X0 U7235 ( .IN1(n4795), .IN2(n6004), .QN(n6464) );
  NAND2X0 U7236 ( .IN1(n5289), .IN2(n8329), .QN(n6004) );
  NAND2X0 U7237 ( .IN1(n6466), .IN2(n6467), .QN(WX9741) );
  NOR2X0 U7238 ( .IN1(n6468), .IN2(n6469), .QN(n6467) );
  NOR2X0 U7239 ( .IN1(n6470), .IN2(n4722), .QN(n6469) );
  NOR2X0 U7240 ( .IN1(n4784), .IN2(n5785), .QN(n6468) );
  XNOR2X1 U7241 ( .IN1(n6471), .IN2(n6472), .Q(n5785) );
  XOR2X1 U7242 ( .IN1(test_so92), .IN2(n9703), .Q(n6472) );
  XOR2X1 U7243 ( .IN1(WX11163), .IN2(n4437), .Q(n6471) );
  NOR2X0 U7244 ( .IN1(n6473), .IN2(n6474), .QN(n6466) );
  NOR2X0 U7245 ( .IN1(DFF_1512_n1), .IN2(n4755), .QN(n6474) );
  NOR2X0 U7246 ( .IN1(n4795), .IN2(n6005), .QN(n6473) );
  NAND2X0 U7247 ( .IN1(n5289), .IN2(n8330), .QN(n6005) );
  NAND2X0 U7248 ( .IN1(n6475), .IN2(n6476), .QN(WX9739) );
  NOR2X0 U7249 ( .IN1(n6477), .IN2(n6478), .QN(n6476) );
  NOR2X0 U7250 ( .IN1(n6479), .IN2(n4722), .QN(n6478) );
  NOR2X0 U7251 ( .IN1(n6480), .IN2(n4770), .QN(n6477) );
  INVX0 U7252 ( .INP(n5794), .ZN(n6480) );
  XNOR2X1 U7253 ( .IN1(n6481), .IN2(n6482), .Q(n5794) );
  XOR2X1 U7254 ( .IN1(n9704), .IN2(n4436), .Q(n6482) );
  XOR2X1 U7255 ( .IN1(WX11033), .IN2(n4161), .Q(n6481) );
  NOR2X0 U7256 ( .IN1(n6483), .IN2(n6484), .QN(n6475) );
  NOR2X0 U7257 ( .IN1(DFF_1513_n1), .IN2(n4755), .QN(n6484) );
  NOR2X0 U7258 ( .IN1(n4795), .IN2(n6006), .QN(n6483) );
  NAND2X0 U7259 ( .IN1(n5288), .IN2(n8331), .QN(n6006) );
  NAND2X0 U7260 ( .IN1(n6485), .IN2(n6486), .QN(WX9737) );
  NOR2X0 U7261 ( .IN1(n6487), .IN2(n6488), .QN(n6486) );
  NOR2X0 U7262 ( .IN1(n6489), .IN2(n4722), .QN(n6488) );
  NOR2X0 U7263 ( .IN1(n6490), .IN2(n4770), .QN(n6487) );
  INVX0 U7264 ( .INP(n5803), .ZN(n6490) );
  XNOR2X1 U7265 ( .IN1(n6491), .IN2(n6492), .Q(n5803) );
  XOR2X1 U7266 ( .IN1(n9705), .IN2(n4435), .Q(n6492) );
  XOR2X1 U7267 ( .IN1(WX11031), .IN2(n4163), .Q(n6491) );
  NOR2X0 U7268 ( .IN1(n6493), .IN2(n6494), .QN(n6485) );
  NOR2X0 U7269 ( .IN1(DFF_1514_n1), .IN2(n4755), .QN(n6494) );
  NOR2X0 U7270 ( .IN1(n4795), .IN2(n6007), .QN(n6493) );
  NAND2X0 U7271 ( .IN1(n5288), .IN2(n8332), .QN(n6007) );
  NAND2X0 U7272 ( .IN1(n6495), .IN2(n6496), .QN(WX9735) );
  NOR2X0 U7273 ( .IN1(n6497), .IN2(n6498), .QN(n6496) );
  NOR2X0 U7274 ( .IN1(n6499), .IN2(n4722), .QN(n6498) );
  NOR2X0 U7275 ( .IN1(n6500), .IN2(n4770), .QN(n6497) );
  INVX0 U7276 ( .INP(n5812), .ZN(n6500) );
  XNOR2X1 U7277 ( .IN1(n6501), .IN2(n6502), .Q(n5812) );
  XOR2X1 U7278 ( .IN1(n9706), .IN2(n4389), .Q(n6502) );
  XOR2X1 U7279 ( .IN1(WX11029), .IN2(n4165), .Q(n6501) );
  NOR2X0 U7280 ( .IN1(n6503), .IN2(n6504), .QN(n6495) );
  NOR2X0 U7281 ( .IN1(DFF_1515_n1), .IN2(n4755), .QN(n6504) );
  NOR2X0 U7282 ( .IN1(n4795), .IN2(n6008), .QN(n6503) );
  NAND2X0 U7283 ( .IN1(n5288), .IN2(n8333), .QN(n6008) );
  NAND2X0 U7284 ( .IN1(n6505), .IN2(n6506), .QN(WX9733) );
  NOR2X0 U7285 ( .IN1(n6507), .IN2(n6508), .QN(n6506) );
  NOR2X0 U7286 ( .IN1(n6509), .IN2(n4722), .QN(n6508) );
  NOR2X0 U7287 ( .IN1(n6510), .IN2(n4770), .QN(n6507) );
  INVX0 U7288 ( .INP(n5821), .ZN(n6510) );
  XNOR2X1 U7289 ( .IN1(n6511), .IN2(n6512), .Q(n5821) );
  XOR2X1 U7290 ( .IN1(n9707), .IN2(n4434), .Q(n6512) );
  XOR2X1 U7291 ( .IN1(WX11027), .IN2(n4167), .Q(n6511) );
  NOR2X0 U7292 ( .IN1(n6513), .IN2(n6514), .QN(n6505) );
  NOR2X0 U7293 ( .IN1(DFF_1516_n1), .IN2(n4755), .QN(n6514) );
  NOR2X0 U7294 ( .IN1(n4795), .IN2(n6009), .QN(n6513) );
  NAND2X0 U7295 ( .IN1(n5288), .IN2(n8334), .QN(n6009) );
  NAND2X0 U7296 ( .IN1(n6515), .IN2(n6516), .QN(WX9731) );
  NOR2X0 U7297 ( .IN1(n6517), .IN2(n6518), .QN(n6516) );
  NOR2X0 U7298 ( .IN1(n6519), .IN2(n4722), .QN(n6518) );
  NOR2X0 U7299 ( .IN1(n6520), .IN2(n4770), .QN(n6517) );
  INVX0 U7300 ( .INP(n5830), .ZN(n6520) );
  XNOR2X1 U7301 ( .IN1(n6521), .IN2(n6522), .Q(n5830) );
  XOR2X1 U7302 ( .IN1(n9708), .IN2(n4433), .Q(n6522) );
  XOR2X1 U7303 ( .IN1(WX11025), .IN2(n4169), .Q(n6521) );
  NOR2X0 U7304 ( .IN1(n6523), .IN2(n6524), .QN(n6515) );
  NOR2X0 U7305 ( .IN1(DFF_1517_n1), .IN2(n4754), .QN(n6524) );
  NOR2X0 U7306 ( .IN1(n4795), .IN2(n6010), .QN(n6523) );
  NAND2X0 U7307 ( .IN1(n5288), .IN2(n8335), .QN(n6010) );
  NAND2X0 U7308 ( .IN1(n6525), .IN2(n6526), .QN(WX9729) );
  NOR2X0 U7309 ( .IN1(n6527), .IN2(n6528), .QN(n6526) );
  NOR2X0 U7310 ( .IN1(n4731), .IN2(n6529), .QN(n6528) );
  NOR2X0 U7311 ( .IN1(n6530), .IN2(n4770), .QN(n6527) );
  INVX0 U7312 ( .INP(n5839), .ZN(n6530) );
  XNOR2X1 U7313 ( .IN1(n6531), .IN2(n6532), .Q(n5839) );
  XOR2X1 U7314 ( .IN1(n9709), .IN2(n4432), .Q(n6532) );
  XOR2X1 U7315 ( .IN1(WX11023), .IN2(n4171), .Q(n6531) );
  NOR2X0 U7316 ( .IN1(n6533), .IN2(n6534), .QN(n6525) );
  NOR2X0 U7317 ( .IN1(DFF_1518_n1), .IN2(n4754), .QN(n6534) );
  NOR2X0 U7318 ( .IN1(n4795), .IN2(n6024), .QN(n6533) );
  NAND2X0 U7319 ( .IN1(n5288), .IN2(n8336), .QN(n6024) );
  NAND2X0 U7320 ( .IN1(n6535), .IN2(n6536), .QN(WX9727) );
  NOR2X0 U7321 ( .IN1(n6537), .IN2(n6538), .QN(n6536) );
  NOR2X0 U7322 ( .IN1(n6539), .IN2(n4722), .QN(n6538) );
  NOR2X0 U7323 ( .IN1(n6540), .IN2(n4771), .QN(n6537) );
  INVX0 U7324 ( .INP(n5848), .ZN(n6540) );
  XNOR2X1 U7325 ( .IN1(n6541), .IN2(n6542), .Q(n5848) );
  XOR2X1 U7326 ( .IN1(n9710), .IN2(n4431), .Q(n6542) );
  XOR2X1 U7327 ( .IN1(WX11021), .IN2(n4173), .Q(n6541) );
  NOR2X0 U7328 ( .IN1(n6543), .IN2(n6544), .QN(n6535) );
  NOR2X0 U7329 ( .IN1(DFF_1519_n1), .IN2(n4754), .QN(n6544) );
  NOR2X0 U7330 ( .IN1(n4795), .IN2(n6025), .QN(n6543) );
  NAND2X0 U7331 ( .IN1(n5287), .IN2(n8337), .QN(n6025) );
  NAND2X0 U7332 ( .IN1(n6545), .IN2(n6546), .QN(WX9725) );
  NOR2X0 U7333 ( .IN1(n6547), .IN2(n6548), .QN(n6546) );
  NOR2X0 U7334 ( .IN1(n4731), .IN2(n6549), .QN(n6548) );
  NOR2X0 U7335 ( .IN1(n6550), .IN2(n4771), .QN(n6547) );
  INVX0 U7336 ( .INP(n5857), .ZN(n6550) );
  XNOR2X1 U7337 ( .IN1(n6551), .IN2(n6552), .Q(n5857) );
  XOR2X1 U7338 ( .IN1(n4039), .IN2(n5247), .Q(n6552) );
  XOR2X1 U7339 ( .IN1(n6553), .IN2(n4388), .Q(n6551) );
  XOR2X1 U7340 ( .IN1(WX11147), .IN2(n9711), .Q(n6553) );
  NOR2X0 U7341 ( .IN1(n6554), .IN2(n6555), .QN(n6545) );
  NOR2X0 U7342 ( .IN1(DFF_1520_n1), .IN2(n4754), .QN(n6555) );
  NOR2X0 U7343 ( .IN1(n4795), .IN2(n6026), .QN(n6554) );
  NAND2X0 U7344 ( .IN1(n5287), .IN2(n8338), .QN(n6026) );
  NAND2X0 U7345 ( .IN1(n6556), .IN2(n6557), .QN(WX9723) );
  NOR2X0 U7346 ( .IN1(n6558), .IN2(n6559), .QN(n6557) );
  NOR2X0 U7347 ( .IN1(n6560), .IN2(n4722), .QN(n6559) );
  NOR2X0 U7348 ( .IN1(n6561), .IN2(n4771), .QN(n6558) );
  INVX0 U7349 ( .INP(n5866), .ZN(n6561) );
  XNOR2X1 U7350 ( .IN1(n6562), .IN2(n6563), .Q(n5866) );
  XOR2X1 U7351 ( .IN1(n4040), .IN2(n5247), .Q(n6563) );
  XOR2X1 U7352 ( .IN1(n6564), .IN2(n4430), .Q(n6562) );
  XOR2X1 U7353 ( .IN1(WX11145), .IN2(n9712), .Q(n6564) );
  NOR2X0 U7354 ( .IN1(n6565), .IN2(n6566), .QN(n6556) );
  NOR2X0 U7355 ( .IN1(DFF_1521_n1), .IN2(n4754), .QN(n6566) );
  NOR2X0 U7356 ( .IN1(n4795), .IN2(n6027), .QN(n6565) );
  NAND2X0 U7357 ( .IN1(n5287), .IN2(n8339), .QN(n6027) );
  NAND2X0 U7358 ( .IN1(n6567), .IN2(n6568), .QN(WX9721) );
  NOR2X0 U7359 ( .IN1(n6569), .IN2(n6570), .QN(n6568) );
  NOR2X0 U7360 ( .IN1(n4731), .IN2(n6571), .QN(n6570) );
  NOR2X0 U7361 ( .IN1(n6572), .IN2(n4771), .QN(n6569) );
  INVX0 U7362 ( .INP(n5875), .ZN(n6572) );
  XNOR2X1 U7363 ( .IN1(n6573), .IN2(n6574), .Q(n5875) );
  XOR2X1 U7364 ( .IN1(n4041), .IN2(n5247), .Q(n6574) );
  XOR2X1 U7365 ( .IN1(n6575), .IN2(n4429), .Q(n6573) );
  XOR2X1 U7366 ( .IN1(WX11143), .IN2(n9713), .Q(n6575) );
  NOR2X0 U7367 ( .IN1(n6576), .IN2(n6577), .QN(n6567) );
  NOR2X0 U7368 ( .IN1(DFF_1522_n1), .IN2(n4754), .QN(n6577) );
  NOR2X0 U7369 ( .IN1(n4795), .IN2(n6028), .QN(n6576) );
  NAND2X0 U7370 ( .IN1(n5287), .IN2(n8340), .QN(n6028) );
  NAND2X0 U7371 ( .IN1(n6578), .IN2(n6579), .QN(WX9719) );
  NOR2X0 U7372 ( .IN1(n6580), .IN2(n6581), .QN(n6579) );
  NOR2X0 U7373 ( .IN1(n6582), .IN2(n4722), .QN(n6581) );
  NOR2X0 U7374 ( .IN1(n4784), .IN2(n5885), .QN(n6580) );
  XNOR2X1 U7375 ( .IN1(n6583), .IN2(n6584), .Q(n5885) );
  XOR2X1 U7376 ( .IN1(n4042), .IN2(n5247), .Q(n6584) );
  XOR2X1 U7377 ( .IN1(WX11077), .IN2(n6585), .Q(n6583) );
  XOR2X1 U7378 ( .IN1(test_so97), .IN2(n9714), .Q(n6585) );
  NOR2X0 U7379 ( .IN1(n6586), .IN2(n6587), .QN(n6578) );
  NOR2X0 U7380 ( .IN1(n4765), .IN2(n4714), .QN(n6587) );
  NOR2X0 U7381 ( .IN1(n4795), .IN2(n6029), .QN(n6586) );
  NAND2X0 U7382 ( .IN1(n5287), .IN2(n8341), .QN(n6029) );
  NAND2X0 U7383 ( .IN1(n6588), .IN2(n6589), .QN(WX9717) );
  NOR2X0 U7384 ( .IN1(n6590), .IN2(n6591), .QN(n6589) );
  NOR2X0 U7385 ( .IN1(n4731), .IN2(n6592), .QN(n6591) );
  NOR2X0 U7386 ( .IN1(n6593), .IN2(n4771), .QN(n6590) );
  INVX0 U7387 ( .INP(n5894), .ZN(n6593) );
  XNOR2X1 U7388 ( .IN1(n6594), .IN2(n6595), .Q(n5894) );
  XOR2X1 U7389 ( .IN1(n4043), .IN2(n5247), .Q(n6595) );
  XOR2X1 U7390 ( .IN1(n6596), .IN2(n4428), .Q(n6594) );
  XOR2X1 U7391 ( .IN1(WX11139), .IN2(n9715), .Q(n6596) );
  NOR2X0 U7392 ( .IN1(n6597), .IN2(n6598), .QN(n6588) );
  NOR2X0 U7393 ( .IN1(DFF_1524_n1), .IN2(n4754), .QN(n6598) );
  NOR2X0 U7394 ( .IN1(n4794), .IN2(n6030), .QN(n6597) );
  NAND2X0 U7395 ( .IN1(n5287), .IN2(n8342), .QN(n6030) );
  NAND2X0 U7396 ( .IN1(n6599), .IN2(n6600), .QN(WX9715) );
  NOR2X0 U7397 ( .IN1(n6601), .IN2(n6602), .QN(n6600) );
  NOR2X0 U7398 ( .IN1(n6603), .IN2(n4721), .QN(n6602) );
  NOR2X0 U7399 ( .IN1(n4785), .IN2(n5904), .QN(n6601) );
  XNOR2X1 U7400 ( .IN1(n6604), .IN2(n6605), .Q(n5904) );
  XOR2X1 U7401 ( .IN1(n4427), .IN2(n5247), .Q(n6605) );
  XOR2X1 U7402 ( .IN1(n6606), .IN2(n9718), .Q(n6604) );
  XOR2X1 U7403 ( .IN1(n9717), .IN2(n9716), .Q(n6606) );
  NOR2X0 U7404 ( .IN1(n6607), .IN2(n6608), .QN(n6599) );
  NOR2X0 U7405 ( .IN1(DFF_1525_n1), .IN2(n4754), .QN(n6608) );
  NOR2X0 U7406 ( .IN1(n4794), .IN2(n6031), .QN(n6607) );
  NAND2X0 U7407 ( .IN1(n5286), .IN2(n8343), .QN(n6031) );
  NAND2X0 U7408 ( .IN1(n6609), .IN2(n6610), .QN(WX9713) );
  NOR2X0 U7409 ( .IN1(n6611), .IN2(n6612), .QN(n6610) );
  NOR2X0 U7410 ( .IN1(n6613), .IN2(n4721), .QN(n6612) );
  NOR2X0 U7411 ( .IN1(n6614), .IN2(n4771), .QN(n6611) );
  INVX0 U7412 ( .INP(n5913), .ZN(n6614) );
  XNOR2X1 U7413 ( .IN1(n6615), .IN2(n6616), .Q(n5913) );
  XOR2X1 U7414 ( .IN1(n4044), .IN2(n5247), .Q(n6616) );
  XOR2X1 U7415 ( .IN1(n6617), .IN2(n4426), .Q(n6615) );
  XOR2X1 U7416 ( .IN1(WX11135), .IN2(n9719), .Q(n6617) );
  NOR2X0 U7417 ( .IN1(n6618), .IN2(n6619), .QN(n6609) );
  NOR2X0 U7418 ( .IN1(DFF_1526_n1), .IN2(n4754), .QN(n6619) );
  NOR2X0 U7419 ( .IN1(n4794), .IN2(n6032), .QN(n6618) );
  NAND2X0 U7420 ( .IN1(test_so78), .IN2(n5323), .QN(n6032) );
  NAND2X0 U7421 ( .IN1(n6620), .IN2(n6621), .QN(WX9711) );
  NOR2X0 U7422 ( .IN1(n6622), .IN2(n6623), .QN(n6621) );
  NOR2X0 U7423 ( .IN1(n6624), .IN2(n4721), .QN(n6623) );
  NOR2X0 U7424 ( .IN1(n4785), .IN2(n5923), .QN(n6622) );
  XNOR2X1 U7425 ( .IN1(n6625), .IN2(n6626), .Q(n5923) );
  XOR2X1 U7426 ( .IN1(n4425), .IN2(n5247), .Q(n6626) );
  XOR2X1 U7427 ( .IN1(n6627), .IN2(n9722), .Q(n6625) );
  XOR2X1 U7428 ( .IN1(n9721), .IN2(n9720), .Q(n6627) );
  NOR2X0 U7429 ( .IN1(n6628), .IN2(n6629), .QN(n6620) );
  NOR2X0 U7430 ( .IN1(DFF_1527_n1), .IN2(n4754), .QN(n6629) );
  NOR2X0 U7431 ( .IN1(n4794), .IN2(n6033), .QN(n6628) );
  NAND2X0 U7432 ( .IN1(n5286), .IN2(n8346), .QN(n6033) );
  NAND2X0 U7433 ( .IN1(n6630), .IN2(n6631), .QN(WX9709) );
  NOR2X0 U7434 ( .IN1(n6632), .IN2(n6633), .QN(n6631) );
  NOR2X0 U7435 ( .IN1(n6634), .IN2(n4721), .QN(n6633) );
  NOR2X0 U7436 ( .IN1(n6635), .IN2(n4771), .QN(n6632) );
  INVX0 U7437 ( .INP(n5932), .ZN(n6635) );
  XNOR2X1 U7438 ( .IN1(n6636), .IN2(n6637), .Q(n5932) );
  XOR2X1 U7439 ( .IN1(n4045), .IN2(n5247), .Q(n6637) );
  XOR2X1 U7440 ( .IN1(n6638), .IN2(n4424), .Q(n6636) );
  XOR2X1 U7441 ( .IN1(WX11131), .IN2(n9723), .Q(n6638) );
  NOR2X0 U7442 ( .IN1(n6639), .IN2(n6640), .QN(n6630) );
  NOR2X0 U7443 ( .IN1(DFF_1528_n1), .IN2(n4754), .QN(n6640) );
  NOR2X0 U7444 ( .IN1(n4794), .IN2(n6034), .QN(n6639) );
  NAND2X0 U7445 ( .IN1(n5286), .IN2(n8347), .QN(n6034) );
  NAND2X0 U7446 ( .IN1(n6641), .IN2(n6642), .QN(WX9707) );
  NOR2X0 U7447 ( .IN1(n6643), .IN2(n6644), .QN(n6642) );
  NOR2X0 U7448 ( .IN1(n6645), .IN2(n4721), .QN(n6644) );
  NOR2X0 U7449 ( .IN1(n4785), .IN2(n5942), .QN(n6643) );
  XNOR2X1 U7450 ( .IN1(n6646), .IN2(n6647), .Q(n5942) );
  XOR2X1 U7451 ( .IN1(n4046), .IN2(n5247), .Q(n6647) );
  XOR2X1 U7452 ( .IN1(n6648), .IN2(n4423), .Q(n6646) );
  XOR2X1 U7453 ( .IN1(WX11065), .IN2(test_so91), .Q(n6648) );
  NOR2X0 U7454 ( .IN1(n6649), .IN2(n6650), .QN(n6641) );
  NOR2X0 U7455 ( .IN1(DFF_1529_n1), .IN2(n4754), .QN(n6650) );
  NOR2X0 U7456 ( .IN1(n4794), .IN2(n6035), .QN(n6649) );
  NAND2X0 U7457 ( .IN1(n5286), .IN2(n8348), .QN(n6035) );
  NAND2X0 U7458 ( .IN1(n6651), .IN2(n6652), .QN(WX9705) );
  NOR2X0 U7459 ( .IN1(n6653), .IN2(n6654), .QN(n6652) );
  NOR2X0 U7460 ( .IN1(n6655), .IN2(n4721), .QN(n6654) );
  NOR2X0 U7461 ( .IN1(n6656), .IN2(n4771), .QN(n6653) );
  INVX0 U7462 ( .INP(n5951), .ZN(n6656) );
  XNOR2X1 U7463 ( .IN1(n6657), .IN2(n6658), .Q(n5951) );
  XOR2X1 U7464 ( .IN1(n4047), .IN2(n5247), .Q(n6658) );
  XOR2X1 U7465 ( .IN1(n6659), .IN2(n4422), .Q(n6657) );
  XOR2X1 U7466 ( .IN1(WX11127), .IN2(n9724), .Q(n6659) );
  NOR2X0 U7467 ( .IN1(n6660), .IN2(n6661), .QN(n6651) );
  NOR2X0 U7468 ( .IN1(DFF_1530_n1), .IN2(n4753), .QN(n6661) );
  NOR2X0 U7469 ( .IN1(n4794), .IN2(n6036), .QN(n6660) );
  NAND2X0 U7470 ( .IN1(n5286), .IN2(n8349), .QN(n6036) );
  NAND2X0 U7471 ( .IN1(n6662), .IN2(n6663), .QN(WX9703) );
  NOR2X0 U7472 ( .IN1(n6664), .IN2(n6665), .QN(n6663) );
  NOR2X0 U7473 ( .IN1(n6666), .IN2(n4721), .QN(n6665) );
  NOR2X0 U7474 ( .IN1(n6667), .IN2(n4771), .QN(n6664) );
  INVX0 U7475 ( .INP(n5960), .ZN(n6667) );
  XNOR2X1 U7476 ( .IN1(n6668), .IN2(n6669), .Q(n5960) );
  XOR2X1 U7477 ( .IN1(n4048), .IN2(n5248), .Q(n6669) );
  XOR2X1 U7478 ( .IN1(n6670), .IN2(n4421), .Q(n6668) );
  XOR2X1 U7479 ( .IN1(WX11125), .IN2(n9725), .Q(n6670) );
  NOR2X0 U7480 ( .IN1(n6671), .IN2(n6672), .QN(n6662) );
  NOR2X0 U7481 ( .IN1(DFF_1531_n1), .IN2(n4753), .QN(n6672) );
  NOR2X0 U7482 ( .IN1(n4794), .IN2(n6037), .QN(n6671) );
  NAND2X0 U7483 ( .IN1(n5286), .IN2(n8350), .QN(n6037) );
  NAND2X0 U7484 ( .IN1(n6673), .IN2(n6674), .QN(WX9701) );
  NOR2X0 U7485 ( .IN1(n6675), .IN2(n6676), .QN(n6674) );
  NOR2X0 U7486 ( .IN1(n6677), .IN2(n4721), .QN(n6676) );
  NOR2X0 U7487 ( .IN1(n6678), .IN2(n4771), .QN(n6675) );
  INVX0 U7488 ( .INP(n5969), .ZN(n6678) );
  XNOR2X1 U7489 ( .IN1(n6679), .IN2(n6680), .Q(n5969) );
  XOR2X1 U7490 ( .IN1(n4049), .IN2(n5248), .Q(n6680) );
  XOR2X1 U7491 ( .IN1(n6681), .IN2(n4420), .Q(n6679) );
  XOR2X1 U7492 ( .IN1(WX11123), .IN2(n9726), .Q(n6681) );
  NOR2X0 U7493 ( .IN1(n6682), .IN2(n6683), .QN(n6673) );
  NOR2X0 U7494 ( .IN1(DFF_1532_n1), .IN2(n4753), .QN(n6683) );
  NOR2X0 U7495 ( .IN1(n4794), .IN2(n6038), .QN(n6682) );
  NAND2X0 U7496 ( .IN1(n5285), .IN2(n8351), .QN(n6038) );
  NAND2X0 U7497 ( .IN1(n6684), .IN2(n6685), .QN(WX9699) );
  NOR2X0 U7498 ( .IN1(n6686), .IN2(n6687), .QN(n6685) );
  NOR2X0 U7499 ( .IN1(n6688), .IN2(n4721), .QN(n6687) );
  NOR2X0 U7500 ( .IN1(n6689), .IN2(n4771), .QN(n6686) );
  INVX0 U7501 ( .INP(n5978), .ZN(n6689) );
  XNOR2X1 U7502 ( .IN1(n6690), .IN2(n6691), .Q(n5978) );
  XOR2X1 U7503 ( .IN1(n4050), .IN2(n5248), .Q(n6691) );
  XOR2X1 U7504 ( .IN1(n6692), .IN2(n4419), .Q(n6690) );
  XOR2X1 U7505 ( .IN1(WX11121), .IN2(n9727), .Q(n6692) );
  NOR2X0 U7506 ( .IN1(n6693), .IN2(n6694), .QN(n6684) );
  NOR2X0 U7507 ( .IN1(DFF_1533_n1), .IN2(n4753), .QN(n6694) );
  NOR2X0 U7508 ( .IN1(n4794), .IN2(n6039), .QN(n6693) );
  NAND2X0 U7509 ( .IN1(n5285), .IN2(n8352), .QN(n6039) );
  NAND2X0 U7510 ( .IN1(n6695), .IN2(n6696), .QN(WX9697) );
  NOR2X0 U7511 ( .IN1(n6697), .IN2(n6698), .QN(n6696) );
  NOR2X0 U7512 ( .IN1(n6699), .IN2(n4721), .QN(n6698) );
  NOR2X0 U7513 ( .IN1(n6700), .IN2(n4771), .QN(n6697) );
  INVX0 U7514 ( .INP(n5987), .ZN(n6700) );
  XNOR2X1 U7515 ( .IN1(n6701), .IN2(n6702), .Q(n5987) );
  XOR2X1 U7516 ( .IN1(n4051), .IN2(n5248), .Q(n6702) );
  XOR2X1 U7517 ( .IN1(n6703), .IN2(n4418), .Q(n6701) );
  XOR2X1 U7518 ( .IN1(WX11119), .IN2(n9728), .Q(n6703) );
  NOR2X0 U7519 ( .IN1(n6704), .IN2(n6705), .QN(n6695) );
  NOR2X0 U7520 ( .IN1(DFF_1534_n1), .IN2(n4753), .QN(n6705) );
  NOR2X0 U7521 ( .IN1(n4794), .IN2(n6040), .QN(n6704) );
  NAND2X0 U7522 ( .IN1(n5285), .IN2(n8353), .QN(n6040) );
  NAND2X0 U7523 ( .IN1(n6706), .IN2(n6707), .QN(WX9695) );
  NOR2X0 U7524 ( .IN1(n6708), .IN2(n6709), .QN(n6707) );
  NOR2X0 U7525 ( .IN1(n4730), .IN2(n6710), .QN(n6709) );
  NOR2X0 U7526 ( .IN1(n6711), .IN2(n4772), .QN(n6708) );
  INVX0 U7527 ( .INP(n5996), .ZN(n6711) );
  XNOR2X1 U7528 ( .IN1(n6712), .IN2(n6713), .Q(n5996) );
  XOR2X1 U7529 ( .IN1(n4031), .IN2(n5248), .Q(n6713) );
  XOR2X1 U7530 ( .IN1(n6714), .IN2(n4417), .Q(n6712) );
  XOR2X1 U7531 ( .IN1(WX11117), .IN2(n9729), .Q(n6714) );
  NOR2X0 U7532 ( .IN1(n6715), .IN2(n6716), .QN(n6706) );
  NOR2X0 U7533 ( .IN1(n4381), .IN2(n6717), .QN(n6716) );
  NOR2X0 U7534 ( .IN1(DFF_1535_n1), .IN2(n4753), .QN(n6715) );
  NOR2X0 U7535 ( .IN1(n5435), .IN2(WX9536), .QN(WX9597) );
  NOR2X0 U7536 ( .IN1(n5429), .IN2(n6718), .QN(WX9084) );
  XOR2X1 U7537 ( .IN1(n4469), .IN2(DFF_1342_n1), .Q(n6718) );
  NOR2X0 U7538 ( .IN1(n5429), .IN2(n6719), .QN(WX9082) );
  XOR2X1 U7539 ( .IN1(n4470), .IN2(DFF_1341_n1), .Q(n6719) );
  NOR2X0 U7540 ( .IN1(n5429), .IN2(n6720), .QN(WX9080) );
  XOR2X1 U7541 ( .IN1(n4471), .IN2(DFF_1340_n1), .Q(n6720) );
  NOR2X0 U7542 ( .IN1(n5429), .IN2(n6721), .QN(WX9078) );
  XOR2X1 U7543 ( .IN1(n4472), .IN2(DFF_1339_n1), .Q(n6721) );
  NOR2X0 U7544 ( .IN1(n5429), .IN2(n6722), .QN(WX9076) );
  XOR2X1 U7545 ( .IN1(n4473), .IN2(DFF_1338_n1), .Q(n6722) );
  NOR2X0 U7546 ( .IN1(n5429), .IN2(n6723), .QN(WX9074) );
  XNOR2X1 U7547 ( .IN1(DFF_1337_n1), .IN2(test_so74), .Q(n6723) );
  NOR2X0 U7548 ( .IN1(n5429), .IN2(n6724), .QN(WX9072) );
  XOR2X1 U7549 ( .IN1(n4474), .IN2(n4695), .Q(n6724) );
  NOR2X0 U7550 ( .IN1(n5429), .IN2(n6725), .QN(WX9070) );
  XOR2X1 U7551 ( .IN1(n4475), .IN2(DFF_1335_n1), .Q(n6725) );
  NOR2X0 U7552 ( .IN1(n5430), .IN2(n6726), .QN(WX9068) );
  XOR2X1 U7553 ( .IN1(n4476), .IN2(DFF_1334_n1), .Q(n6726) );
  NOR2X0 U7554 ( .IN1(n5430), .IN2(n6727), .QN(WX9066) );
  XOR2X1 U7555 ( .IN1(n4477), .IN2(DFF_1333_n1), .Q(n6727) );
  NOR2X0 U7556 ( .IN1(n5430), .IN2(n6728), .QN(WX9064) );
  XOR2X1 U7557 ( .IN1(n4478), .IN2(DFF_1332_n1), .Q(n6728) );
  NOR2X0 U7558 ( .IN1(n5430), .IN2(n6729), .QN(WX9062) );
  XOR2X1 U7559 ( .IN1(n4479), .IN2(DFF_1331_n1), .Q(n6729) );
  NOR2X0 U7560 ( .IN1(n5430), .IN2(n6730), .QN(WX9060) );
  XOR2X1 U7561 ( .IN1(n4480), .IN2(DFF_1330_n1), .Q(n6730) );
  NOR2X0 U7562 ( .IN1(n5430), .IN2(n6731), .QN(WX9058) );
  XOR2X1 U7563 ( .IN1(n4481), .IN2(DFF_1329_n1), .Q(n6731) );
  NOR2X0 U7564 ( .IN1(n5430), .IN2(n6732), .QN(WX9056) );
  XOR2X1 U7565 ( .IN1(n4482), .IN2(DFF_1328_n1), .Q(n6732) );
  NOR2X0 U7566 ( .IN1(n5430), .IN2(n6733), .QN(WX9054) );
  XNOR2X1 U7567 ( .IN1(DFF_1327_n1), .IN2(n6734), .Q(n6733) );
  XOR2X1 U7568 ( .IN1(n4394), .IN2(DFF_1343_n1), .Q(n6734) );
  NOR2X0 U7569 ( .IN1(n5430), .IN2(n6735), .QN(WX9052) );
  XOR2X1 U7570 ( .IN1(n4483), .IN2(DFF_1326_n1), .Q(n6735) );
  NOR2X0 U7571 ( .IN1(n5430), .IN2(n6736), .QN(WX9050) );
  XOR2X1 U7572 ( .IN1(n4484), .IN2(DFF_1325_n1), .Q(n6736) );
  NOR2X0 U7573 ( .IN1(n5430), .IN2(n6737), .QN(WX9048) );
  XOR2X1 U7574 ( .IN1(n4485), .IN2(DFF_1324_n1), .Q(n6737) );
  NOR2X0 U7575 ( .IN1(n5430), .IN2(n6738), .QN(WX9046) );
  XOR2X1 U7576 ( .IN1(n4486), .IN2(DFF_1323_n1), .Q(n6738) );
  NOR2X0 U7577 ( .IN1(n5430), .IN2(n6739), .QN(WX9044) );
  XNOR2X1 U7578 ( .IN1(DFF_1322_n1), .IN2(n6740), .Q(n6739) );
  XOR2X1 U7579 ( .IN1(n4395), .IN2(DFF_1343_n1), .Q(n6740) );
  NOR2X0 U7580 ( .IN1(n5431), .IN2(n6741), .QN(WX9042) );
  XOR2X1 U7581 ( .IN1(n4487), .IN2(DFF_1321_n1), .Q(n6741) );
  NOR2X0 U7582 ( .IN1(n5431), .IN2(n6742), .QN(WX9040) );
  XNOR2X1 U7583 ( .IN1(DFF_1320_n1), .IN2(test_so75), .Q(n6742) );
  NOR2X0 U7584 ( .IN1(n5431), .IN2(n6743), .QN(WX9038) );
  XOR2X1 U7585 ( .IN1(n4488), .IN2(n4694), .Q(n6743) );
  NOR2X0 U7586 ( .IN1(n5431), .IN2(n6744), .QN(WX9036) );
  XOR2X1 U7587 ( .IN1(n4489), .IN2(DFF_1318_n1), .Q(n6744) );
  NOR2X0 U7588 ( .IN1(n5431), .IN2(n6745), .QN(WX9034) );
  XOR2X1 U7589 ( .IN1(n4490), .IN2(DFF_1317_n1), .Q(n6745) );
  NOR2X0 U7590 ( .IN1(n5431), .IN2(n6746), .QN(WX9032) );
  XOR2X1 U7591 ( .IN1(n4491), .IN2(DFF_1316_n1), .Q(n6746) );
  NOR2X0 U7592 ( .IN1(n5431), .IN2(n6747), .QN(WX9030) );
  XNOR2X1 U7593 ( .IN1(DFF_1315_n1), .IN2(n6748), .Q(n6747) );
  XOR2X1 U7594 ( .IN1(n4396), .IN2(DFF_1343_n1), .Q(n6748) );
  NOR2X0 U7595 ( .IN1(n5431), .IN2(n6749), .QN(WX9028) );
  XOR2X1 U7596 ( .IN1(n4492), .IN2(DFF_1314_n1), .Q(n6749) );
  NOR2X0 U7597 ( .IN1(n5431), .IN2(n6750), .QN(WX9026) );
  XOR2X1 U7598 ( .IN1(n4493), .IN2(DFF_1313_n1), .Q(n6750) );
  NOR2X0 U7599 ( .IN1(n5431), .IN2(n6751), .QN(WX9024) );
  XOR2X1 U7600 ( .IN1(n4494), .IN2(DFF_1312_n1), .Q(n6751) );
  NOR2X0 U7601 ( .IN1(n5431), .IN2(n6752), .QN(WX9022) );
  XOR2X1 U7602 ( .IN1(n4411), .IN2(DFF_1343_n1), .Q(n6752) );
  NOR2X0 U7603 ( .IN1(n9504), .IN2(n5344), .QN(WX8496) );
  NOR2X0 U7604 ( .IN1(n9505), .IN2(n5344), .QN(WX8494) );
  NOR2X0 U7605 ( .IN1(n9506), .IN2(n5344), .QN(WX8492) );
  NOR2X0 U7606 ( .IN1(n9507), .IN2(n5344), .QN(WX8490) );
  NOR2X0 U7607 ( .IN1(n9508), .IN2(n5344), .QN(WX8488) );
  NOR2X0 U7608 ( .IN1(n9509), .IN2(n5344), .QN(WX8486) );
  NOR2X0 U7609 ( .IN1(n9510), .IN2(n5344), .QN(WX8484) );
  NOR2X0 U7610 ( .IN1(n9511), .IN2(n5344), .QN(WX8482) );
  NOR2X0 U7611 ( .IN1(n9512), .IN2(n5345), .QN(WX8480) );
  NOR2X0 U7612 ( .IN1(n9513), .IN2(n5345), .QN(WX8478) );
  NOR2X0 U7613 ( .IN1(n9514), .IN2(n5345), .QN(WX8476) );
  NOR2X0 U7614 ( .IN1(n9515), .IN2(n5345), .QN(WX8474) );
  NOR2X0 U7615 ( .IN1(n9516), .IN2(n5345), .QN(WX8472) );
  NOR2X0 U7616 ( .IN1(n9519), .IN2(n5345), .QN(WX8470) );
  NOR2X0 U7617 ( .IN1(n9520), .IN2(n5345), .QN(WX8468) );
  NOR2X0 U7618 ( .IN1(n9523), .IN2(n5345), .QN(WX8466) );
  NAND2X0 U7619 ( .IN1(n6753), .IN2(n6754), .QN(WX8464) );
  NOR2X0 U7620 ( .IN1(n6755), .IN2(n6756), .QN(n6754) );
  NOR2X0 U7621 ( .IN1(n6757), .IN2(n4721), .QN(n6756) );
  NOR2X0 U7622 ( .IN1(n6393), .IN2(n4772), .QN(n6755) );
  XOR2X1 U7623 ( .IN1(n6758), .IN2(n6759), .Q(n6393) );
  XOR2X1 U7624 ( .IN1(n9453), .IN2(n4410), .Q(n6759) );
  XOR2X1 U7625 ( .IN1(WX9758), .IN2(n4175), .Q(n6758) );
  NOR2X0 U7626 ( .IN1(n6760), .IN2(n6761), .QN(n6753) );
  NOR2X0 U7627 ( .IN1(DFF_1312_n1), .IN2(n4753), .QN(n6761) );
  NOR2X0 U7628 ( .IN1(n4794), .IN2(n6041), .QN(n6760) );
  NAND2X0 U7629 ( .IN1(test_so68), .IN2(n5323), .QN(n6041) );
  NAND2X0 U7630 ( .IN1(n6762), .IN2(n6763), .QN(WX8462) );
  NOR2X0 U7631 ( .IN1(n6764), .IN2(n6765), .QN(n6763) );
  NOR2X0 U7632 ( .IN1(n6766), .IN2(n4721), .QN(n6765) );
  NOR2X0 U7633 ( .IN1(n4785), .IN2(n6403), .QN(n6764) );
  XNOR2X1 U7634 ( .IN1(n6767), .IN2(n6768), .Q(n6403) );
  XOR2X1 U7635 ( .IN1(test_so83), .IN2(n9454), .Q(n6768) );
  XOR2X1 U7636 ( .IN1(WX9756), .IN2(n4468), .Q(n6767) );
  NOR2X0 U7637 ( .IN1(n6769), .IN2(n6770), .QN(n6762) );
  NOR2X0 U7638 ( .IN1(DFF_1313_n1), .IN2(n4753), .QN(n6770) );
  NOR2X0 U7639 ( .IN1(n4794), .IN2(n6042), .QN(n6769) );
  NAND2X0 U7640 ( .IN1(n5285), .IN2(n8381), .QN(n6042) );
  NAND2X0 U7641 ( .IN1(n6771), .IN2(n6772), .QN(WX8460) );
  NOR2X0 U7642 ( .IN1(n6773), .IN2(n6774), .QN(n6772) );
  NOR2X0 U7643 ( .IN1(n6775), .IN2(n4720), .QN(n6774) );
  NOR2X0 U7644 ( .IN1(n6413), .IN2(n4772), .QN(n6773) );
  XOR2X1 U7645 ( .IN1(n6776), .IN2(n6777), .Q(n6413) );
  XOR2X1 U7646 ( .IN1(n9455), .IN2(n4467), .Q(n6777) );
  XOR2X1 U7647 ( .IN1(WX9754), .IN2(n4178), .Q(n6776) );
  NOR2X0 U7648 ( .IN1(n6778), .IN2(n6779), .QN(n6771) );
  NOR2X0 U7649 ( .IN1(DFF_1314_n1), .IN2(n4753), .QN(n6779) );
  NOR2X0 U7650 ( .IN1(n4793), .IN2(n6043), .QN(n6778) );
  NAND2X0 U7651 ( .IN1(n5285), .IN2(n8382), .QN(n6043) );
  NAND2X0 U7652 ( .IN1(n6780), .IN2(n6781), .QN(WX8458) );
  NOR2X0 U7653 ( .IN1(n6782), .IN2(n6783), .QN(n6781) );
  NOR2X0 U7654 ( .IN1(n6784), .IN2(n4720), .QN(n6783) );
  NOR2X0 U7655 ( .IN1(n4786), .IN2(n6422), .QN(n6782) );
  XNOR2X1 U7656 ( .IN1(n6785), .IN2(n6786), .Q(n6422) );
  XOR2X1 U7657 ( .IN1(test_so81), .IN2(n9456), .Q(n6786) );
  XOR2X1 U7658 ( .IN1(WX9880), .IN2(n4466), .Q(n6785) );
  NOR2X0 U7659 ( .IN1(n6787), .IN2(n6788), .QN(n6780) );
  NOR2X0 U7660 ( .IN1(DFF_1315_n1), .IN2(n4753), .QN(n6788) );
  NOR2X0 U7661 ( .IN1(n4793), .IN2(n6044), .QN(n6787) );
  NAND2X0 U7662 ( .IN1(n5285), .IN2(n8383), .QN(n6044) );
  NAND2X0 U7663 ( .IN1(n6789), .IN2(n6790), .QN(WX8456) );
  NOR2X0 U7664 ( .IN1(n6791), .IN2(n6792), .QN(n6790) );
  NOR2X0 U7665 ( .IN1(n6793), .IN2(n4720), .QN(n6792) );
  NOR2X0 U7666 ( .IN1(n6432), .IN2(n4772), .QN(n6791) );
  XOR2X1 U7667 ( .IN1(n6794), .IN2(n6795), .Q(n6432) );
  XOR2X1 U7668 ( .IN1(n9457), .IN2(n4393), .Q(n6795) );
  XOR2X1 U7669 ( .IN1(WX9750), .IN2(n4181), .Q(n6794) );
  NOR2X0 U7670 ( .IN1(n6796), .IN2(n6797), .QN(n6789) );
  NOR2X0 U7671 ( .IN1(DFF_1316_n1), .IN2(n4753), .QN(n6797) );
  NOR2X0 U7672 ( .IN1(n4793), .IN2(n6045), .QN(n6796) );
  NAND2X0 U7673 ( .IN1(n5284), .IN2(n8384), .QN(n6045) );
  NAND2X0 U7674 ( .IN1(n6798), .IN2(n6799), .QN(WX8454) );
  NOR2X0 U7675 ( .IN1(n6800), .IN2(n6801), .QN(n6799) );
  NOR2X0 U7676 ( .IN1(n6802), .IN2(n4720), .QN(n6801) );
  NOR2X0 U7677 ( .IN1(n6441), .IN2(n4772), .QN(n6800) );
  XOR2X1 U7678 ( .IN1(n6803), .IN2(n6804), .Q(n6441) );
  XOR2X1 U7679 ( .IN1(n9458), .IN2(n4465), .Q(n6804) );
  XOR2X1 U7680 ( .IN1(WX9748), .IN2(n4183), .Q(n6803) );
  NOR2X0 U7681 ( .IN1(n6805), .IN2(n6806), .QN(n6798) );
  NOR2X0 U7682 ( .IN1(DFF_1317_n1), .IN2(n4753), .QN(n6806) );
  NOR2X0 U7683 ( .IN1(n4793), .IN2(n6046), .QN(n6805) );
  NAND2X0 U7684 ( .IN1(n5284), .IN2(n8385), .QN(n6046) );
  NAND2X0 U7685 ( .IN1(n6807), .IN2(n6808), .QN(WX8452) );
  NOR2X0 U7686 ( .IN1(n6809), .IN2(n6810), .QN(n6808) );
  NOR2X0 U7687 ( .IN1(n6811), .IN2(n4720), .QN(n6810) );
  NOR2X0 U7688 ( .IN1(n6451), .IN2(n4772), .QN(n6809) );
  XOR2X1 U7689 ( .IN1(n6812), .IN2(n6813), .Q(n6451) );
  XOR2X1 U7690 ( .IN1(n9459), .IN2(n4464), .Q(n6813) );
  XOR2X1 U7691 ( .IN1(WX9746), .IN2(n4185), .Q(n6812) );
  NOR2X0 U7692 ( .IN1(n6814), .IN2(n6815), .QN(n6807) );
  NOR2X0 U7693 ( .IN1(DFF_1318_n1), .IN2(n4752), .QN(n6815) );
  NOR2X0 U7694 ( .IN1(n4793), .IN2(n6047), .QN(n6814) );
  NAND2X0 U7695 ( .IN1(n5284), .IN2(n8386), .QN(n6047) );
  NAND2X0 U7696 ( .IN1(n6816), .IN2(n6817), .QN(WX8450) );
  NOR2X0 U7697 ( .IN1(n6818), .IN2(n6819), .QN(n6817) );
  NOR2X0 U7698 ( .IN1(n6820), .IN2(n4720), .QN(n6819) );
  NOR2X0 U7699 ( .IN1(n6460), .IN2(n4772), .QN(n6818) );
  XOR2X1 U7700 ( .IN1(n6821), .IN2(n6822), .Q(n6460) );
  XOR2X1 U7701 ( .IN1(n9460), .IN2(n4463), .Q(n6822) );
  XOR2X1 U7702 ( .IN1(WX9744), .IN2(n4187), .Q(n6821) );
  NOR2X0 U7703 ( .IN1(n6823), .IN2(n6824), .QN(n6816) );
  NOR2X0 U7704 ( .IN1(n4765), .IN2(n4694), .QN(n6824) );
  NOR2X0 U7705 ( .IN1(n4793), .IN2(n6048), .QN(n6823) );
  NAND2X0 U7706 ( .IN1(n5284), .IN2(n8387), .QN(n6048) );
  NAND2X0 U7707 ( .IN1(n6825), .IN2(n6826), .QN(WX8448) );
  NOR2X0 U7708 ( .IN1(n6827), .IN2(n6828), .QN(n6826) );
  NOR2X0 U7709 ( .IN1(n6829), .IN2(n4720), .QN(n6828) );
  NOR2X0 U7710 ( .IN1(n6470), .IN2(n4772), .QN(n6827) );
  XOR2X1 U7711 ( .IN1(n6830), .IN2(n6831), .Q(n6470) );
  XOR2X1 U7712 ( .IN1(n9461), .IN2(n4462), .Q(n6831) );
  XOR2X1 U7713 ( .IN1(WX9742), .IN2(n4189), .Q(n6830) );
  NOR2X0 U7714 ( .IN1(n6832), .IN2(n6833), .QN(n6825) );
  NOR2X0 U7715 ( .IN1(DFF_1320_n1), .IN2(n4752), .QN(n6833) );
  NOR2X0 U7716 ( .IN1(n4793), .IN2(n6049), .QN(n6832) );
  NAND2X0 U7717 ( .IN1(n5284), .IN2(n8388), .QN(n6049) );
  NAND2X0 U7718 ( .IN1(n6834), .IN2(n6835), .QN(WX8446) );
  NOR2X0 U7719 ( .IN1(n6836), .IN2(n6837), .QN(n6835) );
  NOR2X0 U7720 ( .IN1(n4730), .IN2(n6838), .QN(n6837) );
  NOR2X0 U7721 ( .IN1(n6479), .IN2(n4772), .QN(n6836) );
  XOR2X1 U7722 ( .IN1(n6839), .IN2(n6840), .Q(n6479) );
  XOR2X1 U7723 ( .IN1(n9462), .IN2(n4461), .Q(n6840) );
  XOR2X1 U7724 ( .IN1(WX9740), .IN2(n4191), .Q(n6839) );
  NOR2X0 U7725 ( .IN1(n6841), .IN2(n6842), .QN(n6834) );
  NOR2X0 U7726 ( .IN1(DFF_1321_n1), .IN2(n4752), .QN(n6842) );
  NOR2X0 U7727 ( .IN1(n4793), .IN2(n6050), .QN(n6841) );
  NAND2X0 U7728 ( .IN1(n5284), .IN2(n8389), .QN(n6050) );
  NAND2X0 U7729 ( .IN1(n6843), .IN2(n6844), .QN(WX8444) );
  NOR2X0 U7730 ( .IN1(n6845), .IN2(n6846), .QN(n6844) );
  NOR2X0 U7731 ( .IN1(n6847), .IN2(n4720), .QN(n6846) );
  NOR2X0 U7732 ( .IN1(n6489), .IN2(n4772), .QN(n6845) );
  XOR2X1 U7733 ( .IN1(n6848), .IN2(n6849), .Q(n6489) );
  XOR2X1 U7734 ( .IN1(n9463), .IN2(n4460), .Q(n6849) );
  XOR2X1 U7735 ( .IN1(WX9738), .IN2(n4193), .Q(n6848) );
  NOR2X0 U7736 ( .IN1(n6850), .IN2(n6851), .QN(n6843) );
  NOR2X0 U7737 ( .IN1(DFF_1322_n1), .IN2(n4752), .QN(n6851) );
  NOR2X0 U7738 ( .IN1(n4793), .IN2(n6051), .QN(n6850) );
  NAND2X0 U7739 ( .IN1(n5289), .IN2(n8390), .QN(n6051) );
  NAND2X0 U7740 ( .IN1(n6852), .IN2(n6853), .QN(WX8442) );
  NOR2X0 U7741 ( .IN1(n6854), .IN2(n6855), .QN(n6853) );
  NOR2X0 U7742 ( .IN1(n4729), .IN2(n6856), .QN(n6855) );
  NOR2X0 U7743 ( .IN1(n6499), .IN2(n4772), .QN(n6854) );
  XOR2X1 U7744 ( .IN1(n6857), .IN2(n6858), .Q(n6499) );
  XOR2X1 U7745 ( .IN1(n9464), .IN2(n4392), .Q(n6858) );
  XOR2X1 U7746 ( .IN1(WX9736), .IN2(n4195), .Q(n6857) );
  NOR2X0 U7747 ( .IN1(n6859), .IN2(n6860), .QN(n6852) );
  NOR2X0 U7748 ( .IN1(DFF_1323_n1), .IN2(n4752), .QN(n6860) );
  NOR2X0 U7749 ( .IN1(n4793), .IN2(n6052), .QN(n6859) );
  NAND2X0 U7750 ( .IN1(n5319), .IN2(n8391), .QN(n6052) );
  NAND2X0 U7751 ( .IN1(n6861), .IN2(n6862), .QN(WX8440) );
  NOR2X0 U7752 ( .IN1(n6863), .IN2(n6864), .QN(n6862) );
  NOR2X0 U7753 ( .IN1(n6865), .IN2(n4720), .QN(n6864) );
  NOR2X0 U7754 ( .IN1(n6509), .IN2(n4772), .QN(n6863) );
  XOR2X1 U7755 ( .IN1(n6866), .IN2(n6867), .Q(n6509) );
  XOR2X1 U7756 ( .IN1(n9465), .IN2(n4459), .Q(n6867) );
  XOR2X1 U7757 ( .IN1(WX9734), .IN2(n4197), .Q(n6866) );
  NOR2X0 U7758 ( .IN1(n6868), .IN2(n6869), .QN(n6861) );
  NOR2X0 U7759 ( .IN1(DFF_1324_n1), .IN2(n4752), .QN(n6869) );
  NOR2X0 U7760 ( .IN1(n4793), .IN2(n6053), .QN(n6868) );
  NAND2X0 U7761 ( .IN1(n5322), .IN2(n8392), .QN(n6053) );
  NAND2X0 U7762 ( .IN1(n6870), .IN2(n6871), .QN(WX8438) );
  NOR2X0 U7763 ( .IN1(n6872), .IN2(n6873), .QN(n6871) );
  NOR2X0 U7764 ( .IN1(n4730), .IN2(n6874), .QN(n6873) );
  NOR2X0 U7765 ( .IN1(n6519), .IN2(n4773), .QN(n6872) );
  XOR2X1 U7766 ( .IN1(n6875), .IN2(n6876), .Q(n6519) );
  XOR2X1 U7767 ( .IN1(n9466), .IN2(n4458), .Q(n6876) );
  XOR2X1 U7768 ( .IN1(WX9732), .IN2(n4199), .Q(n6875) );
  NOR2X0 U7769 ( .IN1(n6877), .IN2(n6878), .QN(n6870) );
  NOR2X0 U7770 ( .IN1(DFF_1325_n1), .IN2(n4752), .QN(n6878) );
  NOR2X0 U7771 ( .IN1(n4793), .IN2(n6054), .QN(n6877) );
  NAND2X0 U7772 ( .IN1(n5321), .IN2(n8393), .QN(n6054) );
  NAND2X0 U7773 ( .IN1(n6879), .IN2(n6880), .QN(WX8436) );
  NOR2X0 U7774 ( .IN1(n6881), .IN2(n6882), .QN(n6880) );
  NOR2X0 U7775 ( .IN1(n6883), .IN2(n4720), .QN(n6882) );
  NOR2X0 U7776 ( .IN1(n4786), .IN2(n6529), .QN(n6881) );
  XNOR2X1 U7777 ( .IN1(n6884), .IN2(n6885), .Q(n6529) );
  XOR2X1 U7778 ( .IN1(test_so86), .IN2(n9467), .Q(n6885) );
  XOR2X1 U7779 ( .IN1(WX9730), .IN2(n4201), .Q(n6884) );
  NOR2X0 U7780 ( .IN1(n6886), .IN2(n6887), .QN(n6879) );
  NOR2X0 U7781 ( .IN1(DFF_1326_n1), .IN2(n4752), .QN(n6887) );
  NOR2X0 U7782 ( .IN1(n4793), .IN2(n6055), .QN(n6886) );
  NAND2X0 U7783 ( .IN1(n5321), .IN2(n8394), .QN(n6055) );
  NAND2X0 U7784 ( .IN1(n6888), .IN2(n6889), .QN(WX8434) );
  NOR2X0 U7785 ( .IN1(n6890), .IN2(n6891), .QN(n6889) );
  NOR2X0 U7786 ( .IN1(n4729), .IN2(n6892), .QN(n6891) );
  NOR2X0 U7787 ( .IN1(n6539), .IN2(n4773), .QN(n6890) );
  XOR2X1 U7788 ( .IN1(n6893), .IN2(n6894), .Q(n6539) );
  XOR2X1 U7789 ( .IN1(n9468), .IN2(n4457), .Q(n6894) );
  XOR2X1 U7790 ( .IN1(WX9728), .IN2(n4203), .Q(n6893) );
  NOR2X0 U7791 ( .IN1(n6895), .IN2(n6896), .QN(n6888) );
  NOR2X0 U7792 ( .IN1(DFF_1327_n1), .IN2(n4752), .QN(n6896) );
  NOR2X0 U7793 ( .IN1(n4792), .IN2(n6056), .QN(n6895) );
  NAND2X0 U7794 ( .IN1(n5321), .IN2(n8395), .QN(n6056) );
  NAND2X0 U7795 ( .IN1(n6897), .IN2(n6898), .QN(WX8432) );
  NOR2X0 U7796 ( .IN1(n6899), .IN2(n6900), .QN(n6898) );
  NOR2X0 U7797 ( .IN1(n6901), .IN2(n4720), .QN(n6900) );
  NOR2X0 U7798 ( .IN1(n4786), .IN2(n6549), .QN(n6899) );
  XNOR2X1 U7799 ( .IN1(n6902), .IN2(n6903), .Q(n6549) );
  XOR2X1 U7800 ( .IN1(n4391), .IN2(n5248), .Q(n6903) );
  XOR2X1 U7801 ( .IN1(n6904), .IN2(n9471), .Q(n6902) );
  XOR2X1 U7802 ( .IN1(n9470), .IN2(n9469), .Q(n6904) );
  NOR2X0 U7803 ( .IN1(n6905), .IN2(n6906), .QN(n6897) );
  NOR2X0 U7804 ( .IN1(DFF_1328_n1), .IN2(n4752), .QN(n6906) );
  NOR2X0 U7805 ( .IN1(n4792), .IN2(n6057), .QN(n6905) );
  NAND2X0 U7806 ( .IN1(n5321), .IN2(n8396), .QN(n6057) );
  NAND2X0 U7807 ( .IN1(n6907), .IN2(n6908), .QN(WX8430) );
  NOR2X0 U7808 ( .IN1(n6909), .IN2(n6910), .QN(n6908) );
  NOR2X0 U7809 ( .IN1(n6911), .IN2(n4720), .QN(n6910) );
  NOR2X0 U7810 ( .IN1(n6560), .IN2(n4773), .QN(n6909) );
  XOR2X1 U7811 ( .IN1(n6912), .IN2(n6913), .Q(n6560) );
  XOR2X1 U7812 ( .IN1(n4052), .IN2(n5248), .Q(n6913) );
  XOR2X1 U7813 ( .IN1(n6914), .IN2(n4456), .Q(n6912) );
  XOR2X1 U7814 ( .IN1(WX9852), .IN2(n9472), .Q(n6914) );
  NOR2X0 U7815 ( .IN1(n6915), .IN2(n6916), .QN(n6907) );
  NOR2X0 U7816 ( .IN1(DFF_1329_n1), .IN2(n4752), .QN(n6916) );
  NOR2X0 U7817 ( .IN1(n4792), .IN2(n6058), .QN(n6915) );
  NAND2X0 U7818 ( .IN1(test_so67), .IN2(n5324), .QN(n6058) );
  NAND2X0 U7819 ( .IN1(n6917), .IN2(n6918), .QN(WX8428) );
  NOR2X0 U7820 ( .IN1(n6919), .IN2(n6920), .QN(n6918) );
  NOR2X0 U7821 ( .IN1(n6921), .IN2(n4719), .QN(n6920) );
  NOR2X0 U7822 ( .IN1(n4786), .IN2(n6571), .QN(n6919) );
  XNOR2X1 U7823 ( .IN1(n6922), .IN2(n6923), .Q(n6571) );
  XOR2X1 U7824 ( .IN1(n4455), .IN2(n5248), .Q(n6923) );
  XOR2X1 U7825 ( .IN1(n6924), .IN2(n9475), .Q(n6922) );
  XOR2X1 U7826 ( .IN1(n9474), .IN2(n9473), .Q(n6924) );
  NOR2X0 U7827 ( .IN1(n6925), .IN2(n6926), .QN(n6917) );
  NOR2X0 U7828 ( .IN1(DFF_1330_n1), .IN2(n4752), .QN(n6926) );
  NOR2X0 U7829 ( .IN1(n4792), .IN2(n6315), .QN(n6925) );
  NAND2X0 U7830 ( .IN1(n6927), .IN2(n8399), .QN(n6315) );
  NAND2X0 U7831 ( .IN1(n6928), .IN2(n6929), .QN(WX8426) );
  NOR2X0 U7832 ( .IN1(n6930), .IN2(n6931), .QN(n6929) );
  NOR2X0 U7833 ( .IN1(n6932), .IN2(n4719), .QN(n6931) );
  NOR2X0 U7834 ( .IN1(n6582), .IN2(n4773), .QN(n6930) );
  XOR2X1 U7835 ( .IN1(n6933), .IN2(n6934), .Q(n6582) );
  XOR2X1 U7836 ( .IN1(n4053), .IN2(n5248), .Q(n6934) );
  XOR2X1 U7837 ( .IN1(n6935), .IN2(n4454), .Q(n6933) );
  XOR2X1 U7838 ( .IN1(WX9848), .IN2(n9476), .Q(n6935) );
  NOR2X0 U7839 ( .IN1(n6936), .IN2(n6937), .QN(n6928) );
  NOR2X0 U7840 ( .IN1(DFF_1331_n1), .IN2(n4751), .QN(n6937) );
  NOR2X0 U7841 ( .IN1(n4792), .IN2(n6059), .QN(n6936) );
  NAND2X0 U7842 ( .IN1(n5318), .IN2(n8400), .QN(n6059) );
  NAND2X0 U7843 ( .IN1(n6938), .IN2(n6939), .QN(WX8424) );
  NOR2X0 U7844 ( .IN1(n6940), .IN2(n6941), .QN(n6939) );
  NOR2X0 U7845 ( .IN1(n6942), .IN2(n4719), .QN(n6941) );
  NOR2X0 U7846 ( .IN1(n4786), .IN2(n6592), .QN(n6940) );
  XNOR2X1 U7847 ( .IN1(n6943), .IN2(n6944), .Q(n6592) );
  XOR2X1 U7848 ( .IN1(n4054), .IN2(n5248), .Q(n6944) );
  XOR2X1 U7849 ( .IN1(n6945), .IN2(n4453), .Q(n6943) );
  XOR2X1 U7850 ( .IN1(WX9782), .IN2(test_so80), .Q(n6945) );
  NOR2X0 U7851 ( .IN1(n6946), .IN2(n6947), .QN(n6938) );
  NOR2X0 U7852 ( .IN1(DFF_1332_n1), .IN2(n4751), .QN(n6947) );
  NOR2X0 U7853 ( .IN1(n4796), .IN2(n6060), .QN(n6946) );
  NAND2X0 U7854 ( .IN1(n5320), .IN2(n8401), .QN(n6060) );
  NAND2X0 U7855 ( .IN1(n6948), .IN2(n6949), .QN(WX8422) );
  NOR2X0 U7856 ( .IN1(n6950), .IN2(n6951), .QN(n6949) );
  NOR2X0 U7857 ( .IN1(n6952), .IN2(n4719), .QN(n6951) );
  NOR2X0 U7858 ( .IN1(n6603), .IN2(n4773), .QN(n6950) );
  XOR2X1 U7859 ( .IN1(n6953), .IN2(n6954), .Q(n6603) );
  XOR2X1 U7860 ( .IN1(n4055), .IN2(n5248), .Q(n6954) );
  XOR2X1 U7861 ( .IN1(n6955), .IN2(n4452), .Q(n6953) );
  XOR2X1 U7862 ( .IN1(WX9844), .IN2(n9477), .Q(n6955) );
  NOR2X0 U7863 ( .IN1(n6956), .IN2(n6957), .QN(n6948) );
  NOR2X0 U7864 ( .IN1(DFF_1333_n1), .IN2(n4756), .QN(n6957) );
  NOR2X0 U7865 ( .IN1(n4792), .IN2(n6061), .QN(n6956) );
  NAND2X0 U7866 ( .IN1(n5321), .IN2(n8402), .QN(n6061) );
  NAND2X0 U7867 ( .IN1(n6958), .IN2(n6959), .QN(WX8420) );
  NOR2X0 U7868 ( .IN1(n6960), .IN2(n6961), .QN(n6959) );
  NOR2X0 U7869 ( .IN1(n6962), .IN2(n4719), .QN(n6961) );
  NOR2X0 U7870 ( .IN1(n6613), .IN2(n4773), .QN(n6960) );
  XOR2X1 U7871 ( .IN1(n6963), .IN2(n6964), .Q(n6613) );
  XOR2X1 U7872 ( .IN1(n4056), .IN2(n5248), .Q(n6964) );
  XOR2X1 U7873 ( .IN1(n6965), .IN2(n4451), .Q(n6963) );
  XOR2X1 U7874 ( .IN1(WX9842), .IN2(n9478), .Q(n6965) );
  NOR2X0 U7875 ( .IN1(n6966), .IN2(n6967), .QN(n6958) );
  NOR2X0 U7876 ( .IN1(DFF_1334_n1), .IN2(n4751), .QN(n6967) );
  NOR2X0 U7877 ( .IN1(n4792), .IN2(n6062), .QN(n6966) );
  NAND2X0 U7878 ( .IN1(n5320), .IN2(n8403), .QN(n6062) );
  NAND2X0 U7879 ( .IN1(n6968), .IN2(n6969), .QN(WX8418) );
  NOR2X0 U7880 ( .IN1(n6970), .IN2(n6971), .QN(n6969) );
  NOR2X0 U7881 ( .IN1(n6972), .IN2(n4719), .QN(n6971) );
  NOR2X0 U7882 ( .IN1(n6624), .IN2(n4773), .QN(n6970) );
  XOR2X1 U7883 ( .IN1(n6973), .IN2(n6974), .Q(n6624) );
  XOR2X1 U7884 ( .IN1(n4057), .IN2(n5249), .Q(n6974) );
  XOR2X1 U7885 ( .IN1(n6975), .IN2(n4450), .Q(n6973) );
  XOR2X1 U7886 ( .IN1(WX9840), .IN2(n9479), .Q(n6975) );
  NOR2X0 U7887 ( .IN1(n6976), .IN2(n6977), .QN(n6968) );
  NOR2X0 U7888 ( .IN1(DFF_1335_n1), .IN2(n4751), .QN(n6977) );
  NOR2X0 U7889 ( .IN1(n4792), .IN2(n6063), .QN(n6976) );
  NAND2X0 U7890 ( .IN1(n5321), .IN2(n8404), .QN(n6063) );
  NAND2X0 U7891 ( .IN1(n6978), .IN2(n6979), .QN(WX8416) );
  NOR2X0 U7892 ( .IN1(n6980), .IN2(n6981), .QN(n6979) );
  NOR2X0 U7893 ( .IN1(n6982), .IN2(n4719), .QN(n6981) );
  NOR2X0 U7894 ( .IN1(n6634), .IN2(n4773), .QN(n6980) );
  XOR2X1 U7895 ( .IN1(n6983), .IN2(n6984), .Q(n6634) );
  XOR2X1 U7896 ( .IN1(n4058), .IN2(n5249), .Q(n6984) );
  XOR2X1 U7897 ( .IN1(n6985), .IN2(n4449), .Q(n6983) );
  XOR2X1 U7898 ( .IN1(WX9838), .IN2(n9480), .Q(n6985) );
  NOR2X0 U7899 ( .IN1(n6986), .IN2(n6987), .QN(n6978) );
  NOR2X0 U7900 ( .IN1(n4764), .IN2(n4695), .QN(n6987) );
  NOR2X0 U7901 ( .IN1(n4792), .IN2(n6064), .QN(n6986) );
  NAND2X0 U7902 ( .IN1(n5320), .IN2(n8405), .QN(n6064) );
  NAND2X0 U7903 ( .IN1(n6988), .IN2(n6989), .QN(WX8414) );
  NOR2X0 U7904 ( .IN1(n6990), .IN2(n6991), .QN(n6989) );
  NOR2X0 U7905 ( .IN1(n6992), .IN2(n4719), .QN(n6991) );
  NOR2X0 U7906 ( .IN1(n6645), .IN2(n4773), .QN(n6990) );
  XOR2X1 U7907 ( .IN1(n6993), .IN2(n6994), .Q(n6645) );
  XOR2X1 U7908 ( .IN1(n4059), .IN2(n5249), .Q(n6994) );
  XOR2X1 U7909 ( .IN1(n6995), .IN2(n4448), .Q(n6993) );
  XOR2X1 U7910 ( .IN1(WX9836), .IN2(n9481), .Q(n6995) );
  NOR2X0 U7911 ( .IN1(n6996), .IN2(n6997), .QN(n6988) );
  NOR2X0 U7912 ( .IN1(DFF_1337_n1), .IN2(n4751), .QN(n6997) );
  NOR2X0 U7913 ( .IN1(n4792), .IN2(n6065), .QN(n6996) );
  NAND2X0 U7914 ( .IN1(n5320), .IN2(n8406), .QN(n6065) );
  NAND2X0 U7915 ( .IN1(n6998), .IN2(n6999), .QN(WX8412) );
  NOR2X0 U7916 ( .IN1(n7000), .IN2(n7001), .QN(n6999) );
  NOR2X0 U7917 ( .IN1(n4729), .IN2(n7002), .QN(n7001) );
  NOR2X0 U7918 ( .IN1(n6655), .IN2(n4773), .QN(n7000) );
  XOR2X1 U7919 ( .IN1(n7003), .IN2(n7004), .Q(n6655) );
  XOR2X1 U7920 ( .IN1(n4060), .IN2(n5249), .Q(n7004) );
  XOR2X1 U7921 ( .IN1(n7005), .IN2(n4447), .Q(n7003) );
  XOR2X1 U7922 ( .IN1(WX9834), .IN2(n9482), .Q(n7005) );
  NOR2X0 U7923 ( .IN1(n7006), .IN2(n7007), .QN(n6998) );
  NOR2X0 U7924 ( .IN1(DFF_1338_n1), .IN2(n4751), .QN(n7007) );
  NOR2X0 U7925 ( .IN1(n4792), .IN2(n6066), .QN(n7006) );
  NAND2X0 U7926 ( .IN1(n5318), .IN2(n8407), .QN(n6066) );
  NAND2X0 U7927 ( .IN1(n7008), .IN2(n7009), .QN(WX8410) );
  NOR2X0 U7928 ( .IN1(n7010), .IN2(n7011), .QN(n7009) );
  NOR2X0 U7929 ( .IN1(n7012), .IN2(n4719), .QN(n7011) );
  NOR2X0 U7930 ( .IN1(n6666), .IN2(n4773), .QN(n7010) );
  XOR2X1 U7931 ( .IN1(n7013), .IN2(n7014), .Q(n6666) );
  XOR2X1 U7932 ( .IN1(n4061), .IN2(n5249), .Q(n7014) );
  XOR2X1 U7933 ( .IN1(n7015), .IN2(n4446), .Q(n7013) );
  XOR2X1 U7934 ( .IN1(WX9832), .IN2(n9483), .Q(n7015) );
  NOR2X0 U7935 ( .IN1(n7016), .IN2(n7017), .QN(n7008) );
  NOR2X0 U7936 ( .IN1(DFF_1339_n1), .IN2(n4751), .QN(n7017) );
  NOR2X0 U7937 ( .IN1(n4791), .IN2(n6067), .QN(n7016) );
  NAND2X0 U7938 ( .IN1(n5320), .IN2(n8408), .QN(n6067) );
  NAND2X0 U7939 ( .IN1(n7018), .IN2(n7019), .QN(WX8408) );
  NOR2X0 U7940 ( .IN1(n7020), .IN2(n7021), .QN(n7019) );
  NOR2X0 U7941 ( .IN1(n4730), .IN2(n7022), .QN(n7021) );
  NOR2X0 U7942 ( .IN1(n6677), .IN2(n4773), .QN(n7020) );
  XOR2X1 U7943 ( .IN1(n7023), .IN2(n7024), .Q(n6677) );
  XOR2X1 U7944 ( .IN1(n4062), .IN2(n5249), .Q(n7024) );
  XOR2X1 U7945 ( .IN1(n7025), .IN2(n4445), .Q(n7023) );
  XOR2X1 U7946 ( .IN1(WX9830), .IN2(n9484), .Q(n7025) );
  NOR2X0 U7947 ( .IN1(n7026), .IN2(n7027), .QN(n7018) );
  NOR2X0 U7948 ( .IN1(DFF_1340_n1), .IN2(n4751), .QN(n7027) );
  NOR2X0 U7949 ( .IN1(n4792), .IN2(n6068), .QN(n7026) );
  NAND2X0 U7950 ( .IN1(n5317), .IN2(n8409), .QN(n6068) );
  NAND2X0 U7951 ( .IN1(n7028), .IN2(n7029), .QN(WX8406) );
  NOR2X0 U7952 ( .IN1(n7030), .IN2(n7031), .QN(n7029) );
  NOR2X0 U7953 ( .IN1(n7032), .IN2(n4719), .QN(n7031) );
  NOR2X0 U7954 ( .IN1(n6688), .IN2(n4774), .QN(n7030) );
  XOR2X1 U7955 ( .IN1(n7033), .IN2(n7034), .Q(n6688) );
  XOR2X1 U7956 ( .IN1(n4063), .IN2(n5249), .Q(n7034) );
  XOR2X1 U7957 ( .IN1(n7035), .IN2(n4444), .Q(n7033) );
  XOR2X1 U7958 ( .IN1(WX9828), .IN2(n9485), .Q(n7035) );
  NOR2X0 U7959 ( .IN1(n7036), .IN2(n7037), .QN(n7028) );
  NOR2X0 U7960 ( .IN1(DFF_1341_n1), .IN2(n4751), .QN(n7037) );
  NOR2X0 U7961 ( .IN1(n4791), .IN2(n6069), .QN(n7036) );
  NAND2X0 U7962 ( .IN1(n5319), .IN2(n8410), .QN(n6069) );
  NAND2X0 U7963 ( .IN1(n7038), .IN2(n7039), .QN(WX8404) );
  NOR2X0 U7964 ( .IN1(n7040), .IN2(n7041), .QN(n7039) );
  NOR2X0 U7965 ( .IN1(n4729), .IN2(n7042), .QN(n7041) );
  NOR2X0 U7966 ( .IN1(n6699), .IN2(n4774), .QN(n7040) );
  XOR2X1 U7967 ( .IN1(n7043), .IN2(n7044), .Q(n6699) );
  XOR2X1 U7968 ( .IN1(n4064), .IN2(n5249), .Q(n7044) );
  XOR2X1 U7969 ( .IN1(n7045), .IN2(n4443), .Q(n7043) );
  XOR2X1 U7970 ( .IN1(WX9826), .IN2(n9486), .Q(n7045) );
  NOR2X0 U7971 ( .IN1(n7046), .IN2(n7047), .QN(n7038) );
  NOR2X0 U7972 ( .IN1(DFF_1342_n1), .IN2(n4751), .QN(n7047) );
  NOR2X0 U7973 ( .IN1(n4791), .IN2(n6070), .QN(n7046) );
  NAND2X0 U7974 ( .IN1(n5320), .IN2(n8411), .QN(n6070) );
  NAND2X0 U7975 ( .IN1(n7048), .IN2(n7049), .QN(WX8402) );
  NOR2X0 U7976 ( .IN1(n7050), .IN2(n7051), .QN(n7049) );
  NOR2X0 U7977 ( .IN1(n7052), .IN2(n4719), .QN(n7051) );
  NOR2X0 U7978 ( .IN1(n4786), .IN2(n6710), .QN(n7050) );
  XNOR2X1 U7979 ( .IN1(n7053), .IN2(n7054), .Q(n6710) );
  XOR2X1 U7980 ( .IN1(n4032), .IN2(n5249), .Q(n7054) );
  XOR2X1 U7981 ( .IN1(WX9760), .IN2(n7055), .Q(n7053) );
  XOR2X1 U7982 ( .IN1(test_so85), .IN2(n9487), .Q(n7055) );
  NOR2X0 U7983 ( .IN1(n7056), .IN2(n7057), .QN(n7048) );
  NOR2X0 U7984 ( .IN1(n4382), .IN2(n6717), .QN(n7057) );
  NOR2X0 U7985 ( .IN1(DFF_1343_n1), .IN2(n4751), .QN(n7056) );
  NOR2X0 U7986 ( .IN1(n5431), .IN2(WX8243), .QN(WX8304) );
  NOR2X0 U7987 ( .IN1(n5431), .IN2(n7058), .QN(WX7791) );
  XOR2X1 U7988 ( .IN1(n4495), .IN2(DFF_1150_n1), .Q(n7058) );
  NOR2X0 U7989 ( .IN1(n5432), .IN2(n7059), .QN(WX7789) );
  XOR2X1 U7990 ( .IN1(n4496), .IN2(n4697), .Q(n7059) );
  NOR2X0 U7991 ( .IN1(n5432), .IN2(n7060), .QN(WX7787) );
  XOR2X1 U7992 ( .IN1(n4497), .IN2(DFF_1148_n1), .Q(n7060) );
  NOR2X0 U7993 ( .IN1(n5432), .IN2(n7061), .QN(WX7785) );
  XOR2X1 U7994 ( .IN1(n4498), .IN2(DFF_1147_n1), .Q(n7061) );
  NOR2X0 U7995 ( .IN1(n7062), .IN2(n7063), .QN(WX7783) );
  XOR2X1 U7996 ( .IN1(n4499), .IN2(DFF_1146_n1), .Q(n7063) );
  NOR2X0 U7997 ( .IN1(n5432), .IN2(n7064), .QN(WX7781) );
  XOR2X1 U7998 ( .IN1(n4500), .IN2(DFF_1145_n1), .Q(n7064) );
  NOR2X0 U7999 ( .IN1(n5432), .IN2(n7065), .QN(WX7779) );
  XOR2X1 U8000 ( .IN1(n4501), .IN2(DFF_1144_n1), .Q(n7065) );
  NOR2X0 U8001 ( .IN1(n5432), .IN2(n7066), .QN(WX7777) );
  XOR2X1 U8002 ( .IN1(n4502), .IN2(DFF_1143_n1), .Q(n7066) );
  NOR2X0 U8003 ( .IN1(n5432), .IN2(n7067), .QN(WX7775) );
  XOR2X1 U8004 ( .IN1(n4503), .IN2(DFF_1142_n1), .Q(n7067) );
  NOR2X0 U8005 ( .IN1(n5432), .IN2(n7068), .QN(WX7773) );
  XOR2X1 U8006 ( .IN1(n4504), .IN2(DFF_1141_n1), .Q(n7068) );
  NOR2X0 U8007 ( .IN1(n5432), .IN2(n7069), .QN(WX7771) );
  XNOR2X1 U8008 ( .IN1(DFF_1140_n1), .IN2(test_so63), .Q(n7069) );
  NOR2X0 U8009 ( .IN1(n5432), .IN2(n7070), .QN(WX7769) );
  XOR2X1 U8010 ( .IN1(n4505), .IN2(DFF_1139_n1), .Q(n7070) );
  NOR2X0 U8011 ( .IN1(n5432), .IN2(n7071), .QN(WX7767) );
  XOR2X1 U8012 ( .IN1(n4506), .IN2(DFF_1138_n1), .Q(n7071) );
  NOR2X0 U8013 ( .IN1(n5432), .IN2(n7072), .QN(WX7765) );
  XOR2X1 U8014 ( .IN1(n4507), .IN2(DFF_1137_n1), .Q(n7072) );
  NOR2X0 U8015 ( .IN1(n5432), .IN2(n7073), .QN(WX7763) );
  XOR2X1 U8016 ( .IN1(n4508), .IN2(DFF_1136_n1), .Q(n7073) );
  NOR2X0 U8017 ( .IN1(n5433), .IN2(n7074), .QN(WX7761) );
  XNOR2X1 U8018 ( .IN1(DFF_1135_n1), .IN2(n7075), .Q(n7074) );
  XOR2X1 U8019 ( .IN1(n4397), .IN2(DFF_1151_n1), .Q(n7075) );
  NOR2X0 U8020 ( .IN1(n5433), .IN2(n7076), .QN(WX7759) );
  XOR2X1 U8021 ( .IN1(n4509), .IN2(DFF_1134_n1), .Q(n7076) );
  NOR2X0 U8022 ( .IN1(n5433), .IN2(n7077), .QN(WX7757) );
  XOR2X1 U8023 ( .IN1(n4510), .IN2(DFF_1133_n1), .Q(n7077) );
  NOR2X0 U8024 ( .IN1(n5433), .IN2(n7078), .QN(WX7755) );
  XOR2X1 U8025 ( .IN1(n4511), .IN2(n4696), .Q(n7078) );
  NOR2X0 U8026 ( .IN1(n5433), .IN2(n7079), .QN(WX7753) );
  XOR2X1 U8027 ( .IN1(n4512), .IN2(DFF_1131_n1), .Q(n7079) );
  NOR2X0 U8028 ( .IN1(n5433), .IN2(n7080), .QN(WX7751) );
  XNOR2X1 U8029 ( .IN1(DFF_1130_n1), .IN2(n7081), .Q(n7080) );
  XOR2X1 U8030 ( .IN1(n4398), .IN2(DFF_1151_n1), .Q(n7081) );
  NOR2X0 U8031 ( .IN1(n5433), .IN2(n7082), .QN(WX7749) );
  XOR2X1 U8032 ( .IN1(n4513), .IN2(DFF_1129_n1), .Q(n7082) );
  NOR2X0 U8033 ( .IN1(n5433), .IN2(n7083), .QN(WX7747) );
  XOR2X1 U8034 ( .IN1(n4514), .IN2(DFF_1128_n1), .Q(n7083) );
  NOR2X0 U8035 ( .IN1(n5433), .IN2(n7084), .QN(WX7745) );
  XOR2X1 U8036 ( .IN1(n4515), .IN2(DFF_1127_n1), .Q(n7084) );
  NOR2X0 U8037 ( .IN1(n5433), .IN2(n7085), .QN(WX7743) );
  XOR2X1 U8038 ( .IN1(n4516), .IN2(DFF_1126_n1), .Q(n7085) );
  NOR2X0 U8039 ( .IN1(n5433), .IN2(n7086), .QN(WX7741) );
  XOR2X1 U8040 ( .IN1(n4517), .IN2(DFF_1125_n1), .Q(n7086) );
  NOR2X0 U8041 ( .IN1(n5433), .IN2(n7087), .QN(WX7739) );
  XOR2X1 U8042 ( .IN1(n4518), .IN2(DFF_1124_n1), .Q(n7087) );
  NOR2X0 U8043 ( .IN1(n5433), .IN2(n7088), .QN(WX7737) );
  XOR2X1 U8044 ( .IN1(DFF_1123_n1), .IN2(n7089), .Q(n7088) );
  XOR2X1 U8045 ( .IN1(test_so64), .IN2(DFF_1151_n1), .Q(n7089) );
  NOR2X0 U8046 ( .IN1(n5434), .IN2(n7090), .QN(WX7735) );
  XOR2X1 U8047 ( .IN1(n4519), .IN2(DFF_1122_n1), .Q(n7090) );
  NOR2X0 U8048 ( .IN1(n5434), .IN2(n7091), .QN(WX7733) );
  XOR2X1 U8049 ( .IN1(n4520), .IN2(DFF_1121_n1), .Q(n7091) );
  NOR2X0 U8050 ( .IN1(n5434), .IN2(n7092), .QN(WX7731) );
  XOR2X1 U8051 ( .IN1(n4521), .IN2(DFF_1120_n1), .Q(n7092) );
  NOR2X0 U8052 ( .IN1(n5434), .IN2(n7093), .QN(WX7729) );
  XOR2X1 U8053 ( .IN1(n4412), .IN2(DFF_1151_n1), .Q(n7093) );
  NOR2X0 U8054 ( .IN1(n9540), .IN2(n5345), .QN(WX7203) );
  NOR2X0 U8055 ( .IN1(n9541), .IN2(n5345), .QN(WX7201) );
  NOR2X0 U8056 ( .IN1(n9542), .IN2(n5345), .QN(WX7199) );
  NOR2X0 U8057 ( .IN1(n9543), .IN2(n5345), .QN(WX7197) );
  NOR2X0 U8058 ( .IN1(n9544), .IN2(n5346), .QN(WX7195) );
  NOR2X0 U8059 ( .IN1(n9545), .IN2(n5346), .QN(WX7193) );
  NOR2X0 U8060 ( .IN1(n9546), .IN2(n5346), .QN(WX7191) );
  NOR2X0 U8061 ( .IN1(n9547), .IN2(n5346), .QN(WX7189) );
  NOR2X0 U8062 ( .IN1(n9550), .IN2(n5346), .QN(WX7187) );
  NOR2X0 U8063 ( .IN1(n9551), .IN2(n5346), .QN(WX7185) );
  NOR2X0 U8064 ( .IN1(n9554), .IN2(n5346), .QN(WX7183) );
  NOR2X0 U8065 ( .IN1(n5434), .IN2(n4707), .QN(WX7181) );
  NOR2X0 U8066 ( .IN1(n9555), .IN2(n5346), .QN(WX7179) );
  NOR2X0 U8067 ( .IN1(n9556), .IN2(n5346), .QN(WX7177) );
  NOR2X0 U8068 ( .IN1(n9557), .IN2(n5346), .QN(WX7175) );
  NOR2X0 U8069 ( .IN1(n9558), .IN2(n5346), .QN(WX7173) );
  NAND2X0 U8070 ( .IN1(n7094), .IN2(n7095), .QN(WX7171) );
  NOR2X0 U8071 ( .IN1(n7096), .IN2(n7097), .QN(n7095) );
  NOR2X0 U8072 ( .IN1(n7098), .IN2(n4718), .QN(n7097) );
  NOR2X0 U8073 ( .IN1(n6757), .IN2(n4774), .QN(n7096) );
  XOR2X1 U8074 ( .IN1(n7099), .IN2(n7100), .Q(n6757) );
  XOR2X1 U8075 ( .IN1(n9488), .IN2(n4411), .Q(n7100) );
  XOR2X1 U8076 ( .IN1(WX8465), .IN2(n4205), .Q(n7099) );
  NOR2X0 U8077 ( .IN1(n7101), .IN2(n7102), .QN(n7094) );
  NOR2X0 U8078 ( .IN1(DFF_1120_n1), .IN2(n4750), .QN(n7102) );
  NOR2X0 U8079 ( .IN1(n4791), .IN2(n6071), .QN(n7101) );
  NAND2X0 U8080 ( .IN1(n5319), .IN2(n8438), .QN(n6071) );
  NAND2X0 U8081 ( .IN1(n7103), .IN2(n7104), .QN(WX7169) );
  NOR2X0 U8082 ( .IN1(n7105), .IN2(n7106), .QN(n7104) );
  NOR2X0 U8083 ( .IN1(n7107), .IN2(n4718), .QN(n7106) );
  NOR2X0 U8084 ( .IN1(n6766), .IN2(n4774), .QN(n7105) );
  XOR2X1 U8085 ( .IN1(n7108), .IN2(n7109), .Q(n6766) );
  XOR2X1 U8086 ( .IN1(n9489), .IN2(n4494), .Q(n7109) );
  XOR2X1 U8087 ( .IN1(WX8463), .IN2(n4207), .Q(n7108) );
  NOR2X0 U8088 ( .IN1(n7110), .IN2(n7111), .QN(n7103) );
  NOR2X0 U8089 ( .IN1(DFF_1121_n1), .IN2(n4750), .QN(n7111) );
  NOR2X0 U8090 ( .IN1(n4791), .IN2(n6072), .QN(n7110) );
  NAND2X0 U8091 ( .IN1(n5317), .IN2(n8439), .QN(n6072) );
  NAND2X0 U8092 ( .IN1(n7112), .IN2(n7113), .QN(WX7167) );
  NOR2X0 U8093 ( .IN1(n7114), .IN2(n7115), .QN(n7113) );
  NOR2X0 U8094 ( .IN1(n7116), .IN2(n4718), .QN(n7115) );
  NOR2X0 U8095 ( .IN1(n6775), .IN2(n4774), .QN(n7114) );
  XOR2X1 U8096 ( .IN1(n7117), .IN2(n7118), .Q(n6775) );
  XOR2X1 U8097 ( .IN1(n9490), .IN2(n4493), .Q(n7118) );
  XOR2X1 U8098 ( .IN1(WX8461), .IN2(n4209), .Q(n7117) );
  NOR2X0 U8099 ( .IN1(n7119), .IN2(n7120), .QN(n7112) );
  NOR2X0 U8100 ( .IN1(DFF_1122_n1), .IN2(n4750), .QN(n7120) );
  NOR2X0 U8101 ( .IN1(n4791), .IN2(n6073), .QN(n7119) );
  NAND2X0 U8102 ( .IN1(n5319), .IN2(n8440), .QN(n6073) );
  NAND2X0 U8103 ( .IN1(n7121), .IN2(n7122), .QN(WX7165) );
  NOR2X0 U8104 ( .IN1(n7123), .IN2(n7124), .QN(n7122) );
  NOR2X0 U8105 ( .IN1(n7125), .IN2(n4718), .QN(n7124) );
  NOR2X0 U8106 ( .IN1(n6784), .IN2(n4774), .QN(n7123) );
  XOR2X1 U8107 ( .IN1(n7126), .IN2(n7127), .Q(n6784) );
  XOR2X1 U8108 ( .IN1(n9491), .IN2(n4492), .Q(n7127) );
  XOR2X1 U8109 ( .IN1(WX8459), .IN2(n4211), .Q(n7126) );
  NOR2X0 U8110 ( .IN1(n7128), .IN2(n7129), .QN(n7121) );
  NOR2X0 U8111 ( .IN1(DFF_1123_n1), .IN2(n4750), .QN(n7129) );
  NOR2X0 U8112 ( .IN1(n4791), .IN2(n6074), .QN(n7128) );
  NAND2X0 U8113 ( .IN1(n5319), .IN2(n8441), .QN(n6074) );
  NAND2X0 U8114 ( .IN1(n7130), .IN2(n7131), .QN(WX7163) );
  NOR2X0 U8115 ( .IN1(n7132), .IN2(n7133), .QN(n7131) );
  NOR2X0 U8116 ( .IN1(n4729), .IN2(n7134), .QN(n7133) );
  NOR2X0 U8117 ( .IN1(n6793), .IN2(n4774), .QN(n7132) );
  XOR2X1 U8118 ( .IN1(n7135), .IN2(n7136), .Q(n6793) );
  XOR2X1 U8119 ( .IN1(n9492), .IN2(n4396), .Q(n7136) );
  XOR2X1 U8120 ( .IN1(WX8457), .IN2(n4213), .Q(n7135) );
  NOR2X0 U8121 ( .IN1(n7137), .IN2(n7138), .QN(n7130) );
  NOR2X0 U8122 ( .IN1(DFF_1124_n1), .IN2(n4750), .QN(n7138) );
  NOR2X0 U8123 ( .IN1(n4791), .IN2(n6075), .QN(n7137) );
  NAND2X0 U8124 ( .IN1(n5318), .IN2(n8442), .QN(n6075) );
  NAND2X0 U8125 ( .IN1(n7139), .IN2(n7140), .QN(WX7161) );
  NOR2X0 U8126 ( .IN1(n7141), .IN2(n7142), .QN(n7140) );
  NOR2X0 U8127 ( .IN1(n7143), .IN2(n4718), .QN(n7142) );
  NOR2X0 U8128 ( .IN1(n6802), .IN2(n4774), .QN(n7141) );
  XOR2X1 U8129 ( .IN1(n7144), .IN2(n7145), .Q(n6802) );
  XOR2X1 U8130 ( .IN1(n9493), .IN2(n4491), .Q(n7145) );
  XOR2X1 U8131 ( .IN1(WX8455), .IN2(n4215), .Q(n7144) );
  NOR2X0 U8132 ( .IN1(n7146), .IN2(n7147), .QN(n7139) );
  NOR2X0 U8133 ( .IN1(DFF_1125_n1), .IN2(n4750), .QN(n7147) );
  NOR2X0 U8134 ( .IN1(n4791), .IN2(n6326), .QN(n7146) );
  NAND2X0 U8135 ( .IN1(n6927), .IN2(n8443), .QN(n6326) );
  NAND2X0 U8136 ( .IN1(n7148), .IN2(n7149), .QN(WX7159) );
  NOR2X0 U8137 ( .IN1(n7150), .IN2(n7151), .QN(n7149) );
  NOR2X0 U8138 ( .IN1(n4729), .IN2(n7152), .QN(n7151) );
  NOR2X0 U8139 ( .IN1(n6811), .IN2(n4774), .QN(n7150) );
  XOR2X1 U8140 ( .IN1(n7153), .IN2(n7154), .Q(n6811) );
  XOR2X1 U8141 ( .IN1(n9494), .IN2(n4490), .Q(n7154) );
  XOR2X1 U8142 ( .IN1(WX8453), .IN2(n4217), .Q(n7153) );
  NOR2X0 U8143 ( .IN1(n7155), .IN2(n7156), .QN(n7148) );
  NOR2X0 U8144 ( .IN1(DFF_1126_n1), .IN2(n4750), .QN(n7156) );
  NOR2X0 U8145 ( .IN1(n4791), .IN2(n6076), .QN(n7155) );
  NAND2X0 U8146 ( .IN1(n5319), .IN2(n8444), .QN(n6076) );
  NAND2X0 U8147 ( .IN1(n7157), .IN2(n7158), .QN(WX7157) );
  NOR2X0 U8148 ( .IN1(n7159), .IN2(n7160), .QN(n7158) );
  NOR2X0 U8149 ( .IN1(n7161), .IN2(n4718), .QN(n7160) );
  NOR2X0 U8150 ( .IN1(n6820), .IN2(n4774), .QN(n7159) );
  XOR2X1 U8151 ( .IN1(n7162), .IN2(n7163), .Q(n6820) );
  XOR2X1 U8152 ( .IN1(n9495), .IN2(n4489), .Q(n7163) );
  XOR2X1 U8153 ( .IN1(WX8451), .IN2(n4219), .Q(n7162) );
  NOR2X0 U8154 ( .IN1(n7164), .IN2(n7165), .QN(n7157) );
  NOR2X0 U8155 ( .IN1(DFF_1127_n1), .IN2(n4750), .QN(n7165) );
  NOR2X0 U8156 ( .IN1(n4791), .IN2(n6077), .QN(n7164) );
  NAND2X0 U8157 ( .IN1(n5318), .IN2(n8445), .QN(n6077) );
  NAND2X0 U8158 ( .IN1(n7166), .IN2(n7167), .QN(WX7155) );
  NOR2X0 U8159 ( .IN1(n7168), .IN2(n7169), .QN(n7167) );
  NOR2X0 U8160 ( .IN1(n4730), .IN2(n7170), .QN(n7169) );
  NOR2X0 U8161 ( .IN1(n6829), .IN2(n4774), .QN(n7168) );
  XOR2X1 U8162 ( .IN1(n7171), .IN2(n7172), .Q(n6829) );
  XOR2X1 U8163 ( .IN1(n9496), .IN2(n4488), .Q(n7172) );
  XOR2X1 U8164 ( .IN1(WX8449), .IN2(n4221), .Q(n7171) );
  NOR2X0 U8165 ( .IN1(n7173), .IN2(n7174), .QN(n7166) );
  NOR2X0 U8166 ( .IN1(DFF_1128_n1), .IN2(n4750), .QN(n7174) );
  NOR2X0 U8167 ( .IN1(n4791), .IN2(n6078), .QN(n7173) );
  NAND2X0 U8168 ( .IN1(n5317), .IN2(n8446), .QN(n6078) );
  NAND2X0 U8169 ( .IN1(n7175), .IN2(n7176), .QN(WX7153) );
  NOR2X0 U8170 ( .IN1(n7177), .IN2(n7178), .QN(n7176) );
  NOR2X0 U8171 ( .IN1(n7179), .IN2(n4718), .QN(n7178) );
  NOR2X0 U8172 ( .IN1(n4786), .IN2(n6838), .QN(n7177) );
  XNOR2X1 U8173 ( .IN1(n7180), .IN2(n7181), .Q(n6838) );
  XOR2X1 U8174 ( .IN1(test_so75), .IN2(n9497), .Q(n7181) );
  XOR2X1 U8175 ( .IN1(WX8447), .IN2(n4223), .Q(n7180) );
  NOR2X0 U8176 ( .IN1(n7182), .IN2(n7183), .QN(n7175) );
  NOR2X0 U8177 ( .IN1(DFF_1129_n1), .IN2(n4750), .QN(n7183) );
  NOR2X0 U8178 ( .IN1(n4791), .IN2(n6079), .QN(n7182) );
  NAND2X0 U8179 ( .IN1(n5318), .IN2(n8447), .QN(n6079) );
  NAND2X0 U8180 ( .IN1(n7184), .IN2(n7185), .QN(WX7151) );
  NOR2X0 U8181 ( .IN1(n7186), .IN2(n7187), .QN(n7185) );
  NOR2X0 U8182 ( .IN1(n4729), .IN2(n7188), .QN(n7187) );
  NOR2X0 U8183 ( .IN1(n6847), .IN2(n4774), .QN(n7186) );
  XOR2X1 U8184 ( .IN1(n7189), .IN2(n7190), .Q(n6847) );
  XOR2X1 U8185 ( .IN1(n9498), .IN2(n4487), .Q(n7190) );
  XOR2X1 U8186 ( .IN1(WX8445), .IN2(n4225), .Q(n7189) );
  NOR2X0 U8187 ( .IN1(n7191), .IN2(n7192), .QN(n7184) );
  NOR2X0 U8188 ( .IN1(DFF_1130_n1), .IN2(n4750), .QN(n7192) );
  NOR2X0 U8189 ( .IN1(n4790), .IN2(n6080), .QN(n7191) );
  NAND2X0 U8190 ( .IN1(n5315), .IN2(n8448), .QN(n6080) );
  NAND2X0 U8191 ( .IN1(n7193), .IN2(n7194), .QN(WX7149) );
  NOR2X0 U8192 ( .IN1(n7195), .IN2(n7196), .QN(n7194) );
  NOR2X0 U8193 ( .IN1(n7197), .IN2(n4718), .QN(n7196) );
  NOR2X0 U8194 ( .IN1(n4787), .IN2(n6856), .QN(n7195) );
  XNOR2X1 U8195 ( .IN1(n7198), .IN2(n7199), .Q(n6856) );
  XOR2X1 U8196 ( .IN1(test_so73), .IN2(n9499), .Q(n7199) );
  XOR2X1 U8197 ( .IN1(WX8443), .IN2(n4395), .Q(n7198) );
  NOR2X0 U8198 ( .IN1(n7200), .IN2(n7201), .QN(n7193) );
  NOR2X0 U8199 ( .IN1(DFF_1131_n1), .IN2(n4750), .QN(n7201) );
  NOR2X0 U8200 ( .IN1(n4790), .IN2(n6081), .QN(n7200) );
  NAND2X0 U8201 ( .IN1(n5317), .IN2(n8449), .QN(n6081) );
  NAND2X0 U8202 ( .IN1(n7202), .IN2(n7203), .QN(WX7147) );
  NOR2X0 U8203 ( .IN1(n7204), .IN2(n7205), .QN(n7203) );
  NOR2X0 U8204 ( .IN1(n7206), .IN2(n4718), .QN(n7205) );
  NOR2X0 U8205 ( .IN1(n6865), .IN2(n4775), .QN(n7204) );
  XOR2X1 U8206 ( .IN1(n7207), .IN2(n7208), .Q(n6865) );
  XOR2X1 U8207 ( .IN1(n9500), .IN2(n4486), .Q(n7208) );
  XOR2X1 U8208 ( .IN1(WX8441), .IN2(n4228), .Q(n7207) );
  NOR2X0 U8209 ( .IN1(n7209), .IN2(n7210), .QN(n7202) );
  NOR2X0 U8210 ( .IN1(n4765), .IN2(n4696), .QN(n7210) );
  NOR2X0 U8211 ( .IN1(n4790), .IN2(n6082), .QN(n7209) );
  NAND2X0 U8212 ( .IN1(test_so56), .IN2(n5323), .QN(n6082) );
  NAND2X0 U8213 ( .IN1(n7211), .IN2(n7212), .QN(WX7145) );
  NOR2X0 U8214 ( .IN1(n7213), .IN2(n7214), .QN(n7212) );
  NOR2X0 U8215 ( .IN1(n7215), .IN2(n4718), .QN(n7214) );
  NOR2X0 U8216 ( .IN1(n4787), .IN2(n6874), .QN(n7213) );
  XNOR2X1 U8217 ( .IN1(n7216), .IN2(n7217), .Q(n6874) );
  XOR2X1 U8218 ( .IN1(test_so71), .IN2(n9501), .Q(n7217) );
  XOR2X1 U8219 ( .IN1(WX8439), .IN2(n4485), .Q(n7216) );
  NOR2X0 U8220 ( .IN1(n7218), .IN2(n7219), .QN(n7211) );
  NOR2X0 U8221 ( .IN1(DFF_1133_n1), .IN2(n4749), .QN(n7219) );
  NOR2X0 U8222 ( .IN1(n4790), .IN2(n6083), .QN(n7218) );
  NAND2X0 U8223 ( .IN1(n5318), .IN2(n8452), .QN(n6083) );
  NAND2X0 U8224 ( .IN1(n7220), .IN2(n7221), .QN(WX7143) );
  NOR2X0 U8225 ( .IN1(n7222), .IN2(n7223), .QN(n7221) );
  NOR2X0 U8226 ( .IN1(n7224), .IN2(n4718), .QN(n7223) );
  NOR2X0 U8227 ( .IN1(n6883), .IN2(n4775), .QN(n7222) );
  XOR2X1 U8228 ( .IN1(n7225), .IN2(n7226), .Q(n6883) );
  XOR2X1 U8229 ( .IN1(n9502), .IN2(n4484), .Q(n7226) );
  XOR2X1 U8230 ( .IN1(WX8437), .IN2(n4231), .Q(n7225) );
  NOR2X0 U8231 ( .IN1(n7227), .IN2(n7228), .QN(n7220) );
  NOR2X0 U8232 ( .IN1(DFF_1134_n1), .IN2(n4749), .QN(n7228) );
  NOR2X0 U8233 ( .IN1(n4790), .IN2(n6084), .QN(n7227) );
  NAND2X0 U8234 ( .IN1(n5314), .IN2(n8453), .QN(n6084) );
  NAND2X0 U8235 ( .IN1(n7229), .IN2(n7230), .QN(WX7141) );
  NOR2X0 U8236 ( .IN1(n7231), .IN2(n7232), .QN(n7230) );
  NOR2X0 U8237 ( .IN1(n7233), .IN2(n4718), .QN(n7232) );
  NOR2X0 U8238 ( .IN1(n4787), .IN2(n6892), .QN(n7231) );
  XNOR2X1 U8239 ( .IN1(n7234), .IN2(n7235), .Q(n6892) );
  XOR2X1 U8240 ( .IN1(test_so69), .IN2(n9503), .Q(n7235) );
  XOR2X1 U8241 ( .IN1(WX8563), .IN2(n4483), .Q(n7234) );
  NOR2X0 U8242 ( .IN1(n7236), .IN2(n7237), .QN(n7229) );
  NOR2X0 U8243 ( .IN1(DFF_1135_n1), .IN2(n4749), .QN(n7237) );
  NOR2X0 U8244 ( .IN1(n4790), .IN2(n6085), .QN(n7236) );
  NAND2X0 U8245 ( .IN1(n5317), .IN2(n8454), .QN(n6085) );
  NAND2X0 U8246 ( .IN1(n7238), .IN2(n7239), .QN(WX7139) );
  NOR2X0 U8247 ( .IN1(n7240), .IN2(n7241), .QN(n7239) );
  NOR2X0 U8248 ( .IN1(n7242), .IN2(n4717), .QN(n7241) );
  NOR2X0 U8249 ( .IN1(n6901), .IN2(n4775), .QN(n7240) );
  XOR2X1 U8250 ( .IN1(n7243), .IN2(n7244), .Q(n6901) );
  XOR2X1 U8251 ( .IN1(n4065), .IN2(n5249), .Q(n7244) );
  XOR2X1 U8252 ( .IN1(n7245), .IN2(n4394), .Q(n7243) );
  XOR2X1 U8253 ( .IN1(WX8561), .IN2(n9504), .Q(n7245) );
  NOR2X0 U8254 ( .IN1(n7246), .IN2(n7247), .QN(n7238) );
  NOR2X0 U8255 ( .IN1(DFF_1136_n1), .IN2(n4749), .QN(n7247) );
  NOR2X0 U8256 ( .IN1(n4790), .IN2(n6095), .QN(n7246) );
  NAND2X0 U8257 ( .IN1(n5314), .IN2(n8455), .QN(n6095) );
  NAND2X0 U8258 ( .IN1(n7248), .IN2(n7249), .QN(WX7137) );
  NOR2X0 U8259 ( .IN1(n7250), .IN2(n7251), .QN(n7249) );
  NOR2X0 U8260 ( .IN1(n7252), .IN2(n4717), .QN(n7251) );
  NOR2X0 U8261 ( .IN1(n6911), .IN2(n4775), .QN(n7250) );
  XOR2X1 U8262 ( .IN1(n7253), .IN2(n7254), .Q(n6911) );
  XOR2X1 U8263 ( .IN1(n4066), .IN2(n5249), .Q(n7254) );
  XOR2X1 U8264 ( .IN1(n7255), .IN2(n4482), .Q(n7253) );
  XOR2X1 U8265 ( .IN1(WX8559), .IN2(n9505), .Q(n7255) );
  NOR2X0 U8266 ( .IN1(n7256), .IN2(n7257), .QN(n7248) );
  NOR2X0 U8267 ( .IN1(DFF_1137_n1), .IN2(n4749), .QN(n7257) );
  NOR2X0 U8268 ( .IN1(n4790), .IN2(n6096), .QN(n7256) );
  NAND2X0 U8269 ( .IN1(n5317), .IN2(n8456), .QN(n6096) );
  NAND2X0 U8270 ( .IN1(n7258), .IN2(n7259), .QN(WX7135) );
  NOR2X0 U8271 ( .IN1(n7260), .IN2(n7261), .QN(n7259) );
  NOR2X0 U8272 ( .IN1(n7262), .IN2(n4717), .QN(n7261) );
  NOR2X0 U8273 ( .IN1(n6921), .IN2(n4775), .QN(n7260) );
  XOR2X1 U8274 ( .IN1(n7263), .IN2(n7264), .Q(n6921) );
  XOR2X1 U8275 ( .IN1(n4067), .IN2(n5249), .Q(n7264) );
  XOR2X1 U8276 ( .IN1(n7265), .IN2(n4481), .Q(n7263) );
  XOR2X1 U8277 ( .IN1(WX8557), .IN2(n9506), .Q(n7265) );
  NOR2X0 U8278 ( .IN1(n7266), .IN2(n7267), .QN(n7258) );
  NOR2X0 U8279 ( .IN1(DFF_1138_n1), .IN2(n4749), .QN(n7267) );
  NOR2X0 U8280 ( .IN1(n4790), .IN2(n6097), .QN(n7266) );
  NAND2X0 U8281 ( .IN1(n5316), .IN2(n8457), .QN(n6097) );
  NAND2X0 U8282 ( .IN1(n7268), .IN2(n7269), .QN(WX7133) );
  NOR2X0 U8283 ( .IN1(n7270), .IN2(n7271), .QN(n7269) );
  NOR2X0 U8284 ( .IN1(n7272), .IN2(n4717), .QN(n7271) );
  NOR2X0 U8285 ( .IN1(n6932), .IN2(n4775), .QN(n7270) );
  XOR2X1 U8286 ( .IN1(n7273), .IN2(n7274), .Q(n6932) );
  XOR2X1 U8287 ( .IN1(n4068), .IN2(n5253), .Q(n7274) );
  XOR2X1 U8288 ( .IN1(n7275), .IN2(n4480), .Q(n7273) );
  XOR2X1 U8289 ( .IN1(WX8555), .IN2(n9507), .Q(n7275) );
  NOR2X0 U8290 ( .IN1(n7276), .IN2(n7277), .QN(n7268) );
  NOR2X0 U8291 ( .IN1(DFF_1139_n1), .IN2(n4749), .QN(n7277) );
  NOR2X0 U8292 ( .IN1(n4790), .IN2(n6098), .QN(n7276) );
  NAND2X0 U8293 ( .IN1(n5316), .IN2(n8458), .QN(n6098) );
  NAND2X0 U8294 ( .IN1(n7278), .IN2(n7279), .QN(WX7131) );
  NOR2X0 U8295 ( .IN1(n7280), .IN2(n7281), .QN(n7279) );
  NOR2X0 U8296 ( .IN1(n7282), .IN2(n4717), .QN(n7281) );
  NOR2X0 U8297 ( .IN1(n6942), .IN2(n4775), .QN(n7280) );
  XOR2X1 U8298 ( .IN1(n7283), .IN2(n7284), .Q(n6942) );
  XOR2X1 U8299 ( .IN1(n4069), .IN2(n5250), .Q(n7284) );
  XOR2X1 U8300 ( .IN1(n7285), .IN2(n4479), .Q(n7283) );
  XOR2X1 U8301 ( .IN1(WX8553), .IN2(n9508), .Q(n7285) );
  NOR2X0 U8302 ( .IN1(n7286), .IN2(n7287), .QN(n7278) );
  NOR2X0 U8303 ( .IN1(DFF_1140_n1), .IN2(n4749), .QN(n7287) );
  NOR2X0 U8304 ( .IN1(n4790), .IN2(n6099), .QN(n7286) );
  NAND2X0 U8305 ( .IN1(n5316), .IN2(n8459), .QN(n6099) );
  NAND2X0 U8306 ( .IN1(n7288), .IN2(n7289), .QN(WX7129) );
  NOR2X0 U8307 ( .IN1(n7290), .IN2(n7291), .QN(n7289) );
  NOR2X0 U8308 ( .IN1(n4730), .IN2(n7292), .QN(n7291) );
  NOR2X0 U8309 ( .IN1(n6952), .IN2(n4775), .QN(n7290) );
  XOR2X1 U8310 ( .IN1(n7293), .IN2(n7294), .Q(n6952) );
  XOR2X1 U8311 ( .IN1(n4070), .IN2(n5250), .Q(n7294) );
  XOR2X1 U8312 ( .IN1(n7295), .IN2(n4478), .Q(n7293) );
  XOR2X1 U8313 ( .IN1(WX8551), .IN2(n9509), .Q(n7295) );
  NOR2X0 U8314 ( .IN1(n7296), .IN2(n7297), .QN(n7288) );
  NOR2X0 U8315 ( .IN1(DFF_1141_n1), .IN2(n4749), .QN(n7297) );
  NOR2X0 U8316 ( .IN1(n4790), .IN2(n6100), .QN(n7296) );
  NAND2X0 U8317 ( .IN1(n5316), .IN2(n8460), .QN(n6100) );
  NAND2X0 U8318 ( .IN1(n7298), .IN2(n7299), .QN(WX7127) );
  NOR2X0 U8319 ( .IN1(n7300), .IN2(n7301), .QN(n7299) );
  NOR2X0 U8320 ( .IN1(n7302), .IN2(n4717), .QN(n7301) );
  NOR2X0 U8321 ( .IN1(n6962), .IN2(n4775), .QN(n7300) );
  XOR2X1 U8322 ( .IN1(n7303), .IN2(n7304), .Q(n6962) );
  XOR2X1 U8323 ( .IN1(n4071), .IN2(n5250), .Q(n7304) );
  XOR2X1 U8324 ( .IN1(n7305), .IN2(n4477), .Q(n7303) );
  XOR2X1 U8325 ( .IN1(WX8549), .IN2(n9510), .Q(n7305) );
  NOR2X0 U8326 ( .IN1(n7306), .IN2(n7307), .QN(n7298) );
  NOR2X0 U8327 ( .IN1(DFF_1142_n1), .IN2(n4749), .QN(n7307) );
  NOR2X0 U8328 ( .IN1(n4789), .IN2(n6101), .QN(n7306) );
  NAND2X0 U8329 ( .IN1(n5316), .IN2(n8461), .QN(n6101) );
  NAND2X0 U8330 ( .IN1(n7308), .IN2(n7309), .QN(WX7125) );
  NOR2X0 U8331 ( .IN1(n7310), .IN2(n7311), .QN(n7309) );
  NOR2X0 U8332 ( .IN1(n4729), .IN2(n7312), .QN(n7311) );
  NOR2X0 U8333 ( .IN1(n6972), .IN2(n4775), .QN(n7310) );
  XOR2X1 U8334 ( .IN1(n7313), .IN2(n7314), .Q(n6972) );
  XOR2X1 U8335 ( .IN1(n4072), .IN2(n5250), .Q(n7314) );
  XOR2X1 U8336 ( .IN1(n7315), .IN2(n4476), .Q(n7313) );
  XOR2X1 U8337 ( .IN1(WX8547), .IN2(n9511), .Q(n7315) );
  NOR2X0 U8338 ( .IN1(n7316), .IN2(n7317), .QN(n7308) );
  NOR2X0 U8339 ( .IN1(DFF_1143_n1), .IN2(n4749), .QN(n7317) );
  NOR2X0 U8340 ( .IN1(n4790), .IN2(n6102), .QN(n7316) );
  NAND2X0 U8341 ( .IN1(n5313), .IN2(n8462), .QN(n6102) );
  NAND2X0 U8342 ( .IN1(n7318), .IN2(n7319), .QN(WX7123) );
  NOR2X0 U8343 ( .IN1(n7320), .IN2(n7321), .QN(n7319) );
  NOR2X0 U8344 ( .IN1(n7322), .IN2(n4717), .QN(n7321) );
  NOR2X0 U8345 ( .IN1(n6982), .IN2(n4775), .QN(n7320) );
  XOR2X1 U8346 ( .IN1(n7323), .IN2(n7324), .Q(n6982) );
  XOR2X1 U8347 ( .IN1(n4073), .IN2(n5250), .Q(n7324) );
  XOR2X1 U8348 ( .IN1(n7325), .IN2(n4475), .Q(n7323) );
  XOR2X1 U8349 ( .IN1(WX8545), .IN2(n9512), .Q(n7325) );
  NOR2X0 U8350 ( .IN1(n7326), .IN2(n7327), .QN(n7318) );
  NOR2X0 U8351 ( .IN1(DFF_1144_n1), .IN2(n4749), .QN(n7327) );
  NOR2X0 U8352 ( .IN1(n4789), .IN2(n6103), .QN(n7326) );
  NAND2X0 U8353 ( .IN1(n5316), .IN2(n8463), .QN(n6103) );
  NAND2X0 U8354 ( .IN1(n7328), .IN2(n7329), .QN(WX7121) );
  NOR2X0 U8355 ( .IN1(n7330), .IN2(n7331), .QN(n7329) );
  NOR2X0 U8356 ( .IN1(n4731), .IN2(n7332), .QN(n7331) );
  NOR2X0 U8357 ( .IN1(n6992), .IN2(n4775), .QN(n7330) );
  XOR2X1 U8358 ( .IN1(n7333), .IN2(n7334), .Q(n6992) );
  XOR2X1 U8359 ( .IN1(n4074), .IN2(n5250), .Q(n7334) );
  XOR2X1 U8360 ( .IN1(n7335), .IN2(n4474), .Q(n7333) );
  XOR2X1 U8361 ( .IN1(WX8543), .IN2(n9513), .Q(n7335) );
  NOR2X0 U8362 ( .IN1(n7336), .IN2(n7337), .QN(n7328) );
  NOR2X0 U8363 ( .IN1(DFF_1145_n1), .IN2(n4748), .QN(n7337) );
  NOR2X0 U8364 ( .IN1(n4789), .IN2(n6104), .QN(n7336) );
  NAND2X0 U8365 ( .IN1(n5315), .IN2(n8464), .QN(n6104) );
  NAND2X0 U8366 ( .IN1(n7338), .IN2(n7339), .QN(WX7119) );
  NOR2X0 U8367 ( .IN1(n7340), .IN2(n7341), .QN(n7339) );
  NOR2X0 U8368 ( .IN1(n7342), .IN2(n4717), .QN(n7341) );
  NOR2X0 U8369 ( .IN1(n4787), .IN2(n7002), .QN(n7340) );
  XNOR2X1 U8370 ( .IN1(n7343), .IN2(n7344), .Q(n7002) );
  XOR2X1 U8371 ( .IN1(n4075), .IN2(n5250), .Q(n7344) );
  XOR2X1 U8372 ( .IN1(WX8477), .IN2(n7345), .Q(n7343) );
  XOR2X1 U8373 ( .IN1(test_so74), .IN2(n9514), .Q(n7345) );
  NOR2X0 U8374 ( .IN1(n7346), .IN2(n7347), .QN(n7338) );
  NOR2X0 U8375 ( .IN1(DFF_1146_n1), .IN2(n4748), .QN(n7347) );
  NOR2X0 U8376 ( .IN1(n4789), .IN2(n6105), .QN(n7346) );
  NAND2X0 U8377 ( .IN1(n5315), .IN2(n8465), .QN(n6105) );
  NAND2X0 U8378 ( .IN1(n7348), .IN2(n7349), .QN(WX7117) );
  NOR2X0 U8379 ( .IN1(n7350), .IN2(n7351), .QN(n7349) );
  NOR2X0 U8380 ( .IN1(n4730), .IN2(n7352), .QN(n7351) );
  NOR2X0 U8381 ( .IN1(n7012), .IN2(n4776), .QN(n7350) );
  XOR2X1 U8382 ( .IN1(n7353), .IN2(n7354), .Q(n7012) );
  XOR2X1 U8383 ( .IN1(n4076), .IN2(n5250), .Q(n7354) );
  XOR2X1 U8384 ( .IN1(n7355), .IN2(n4473), .Q(n7353) );
  XOR2X1 U8385 ( .IN1(WX8539), .IN2(n9515), .Q(n7355) );
  NOR2X0 U8386 ( .IN1(n7356), .IN2(n7357), .QN(n7348) );
  NOR2X0 U8387 ( .IN1(DFF_1147_n1), .IN2(n4748), .QN(n7357) );
  NOR2X0 U8388 ( .IN1(n4789), .IN2(n6106), .QN(n7356) );
  NAND2X0 U8389 ( .IN1(n5315), .IN2(n8466), .QN(n6106) );
  NAND2X0 U8390 ( .IN1(n7358), .IN2(n7359), .QN(WX7115) );
  NOR2X0 U8391 ( .IN1(n7360), .IN2(n7361), .QN(n7359) );
  NOR2X0 U8392 ( .IN1(n7362), .IN2(n4717), .QN(n7361) );
  NOR2X0 U8393 ( .IN1(n4787), .IN2(n7022), .QN(n7360) );
  XNOR2X1 U8394 ( .IN1(n7363), .IN2(n7364), .Q(n7022) );
  XOR2X1 U8395 ( .IN1(n4472), .IN2(n5250), .Q(n7364) );
  XOR2X1 U8396 ( .IN1(n7365), .IN2(n9518), .Q(n7363) );
  XOR2X1 U8397 ( .IN1(n9517), .IN2(n9516), .Q(n7365) );
  NOR2X0 U8398 ( .IN1(n7366), .IN2(n7367), .QN(n7358) );
  NOR2X0 U8399 ( .IN1(DFF_1148_n1), .IN2(n4748), .QN(n7367) );
  NOR2X0 U8400 ( .IN1(n4789), .IN2(n6107), .QN(n7366) );
  NAND2X0 U8401 ( .IN1(n5315), .IN2(n8467), .QN(n6107) );
  NAND2X0 U8402 ( .IN1(n7368), .IN2(n7369), .QN(WX7113) );
  NOR2X0 U8403 ( .IN1(n7370), .IN2(n7371), .QN(n7369) );
  NOR2X0 U8404 ( .IN1(n7372), .IN2(n4717), .QN(n7371) );
  NOR2X0 U8405 ( .IN1(n7032), .IN2(n4776), .QN(n7370) );
  XOR2X1 U8406 ( .IN1(n7373), .IN2(n7374), .Q(n7032) );
  XOR2X1 U8407 ( .IN1(n4077), .IN2(n5250), .Q(n7374) );
  XOR2X1 U8408 ( .IN1(n7375), .IN2(n4471), .Q(n7373) );
  XOR2X1 U8409 ( .IN1(WX8535), .IN2(n9519), .Q(n7375) );
  NOR2X0 U8410 ( .IN1(n7376), .IN2(n7377), .QN(n7368) );
  NOR2X0 U8411 ( .IN1(n4764), .IN2(n4697), .QN(n7377) );
  NOR2X0 U8412 ( .IN1(n4789), .IN2(n6108), .QN(n7376) );
  NAND2X0 U8413 ( .IN1(test_so55), .IN2(n5324), .QN(n6108) );
  NAND2X0 U8414 ( .IN1(n7378), .IN2(n7379), .QN(WX7111) );
  NOR2X0 U8415 ( .IN1(n7380), .IN2(n7381), .QN(n7379) );
  NOR2X0 U8416 ( .IN1(n7382), .IN2(n4717), .QN(n7381) );
  NOR2X0 U8417 ( .IN1(n4787), .IN2(n7042), .QN(n7380) );
  XNOR2X1 U8418 ( .IN1(n7383), .IN2(n7384), .Q(n7042) );
  XOR2X1 U8419 ( .IN1(n4470), .IN2(n5250), .Q(n7384) );
  XOR2X1 U8420 ( .IN1(n7385), .IN2(n9522), .Q(n7383) );
  XOR2X1 U8421 ( .IN1(n9521), .IN2(n9520), .Q(n7385) );
  NOR2X0 U8422 ( .IN1(n7386), .IN2(n7387), .QN(n7378) );
  NOR2X0 U8423 ( .IN1(DFF_1150_n1), .IN2(n4748), .QN(n7387) );
  NOR2X0 U8424 ( .IN1(n4789), .IN2(n6109), .QN(n7386) );
  NAND2X0 U8425 ( .IN1(n5315), .IN2(n8470), .QN(n6109) );
  NAND2X0 U8426 ( .IN1(n7388), .IN2(n7389), .QN(WX7109) );
  NOR2X0 U8427 ( .IN1(n7390), .IN2(n7391), .QN(n7389) );
  NOR2X0 U8428 ( .IN1(n7392), .IN2(n4717), .QN(n7391) );
  NOR2X0 U8429 ( .IN1(n7052), .IN2(n4776), .QN(n7390) );
  XOR2X1 U8430 ( .IN1(n7393), .IN2(n7394), .Q(n7052) );
  XOR2X1 U8431 ( .IN1(n4033), .IN2(n5250), .Q(n7394) );
  XOR2X1 U8432 ( .IN1(n7395), .IN2(n4469), .Q(n7393) );
  XOR2X1 U8433 ( .IN1(WX8531), .IN2(n9523), .Q(n7395) );
  NOR2X0 U8434 ( .IN1(n7396), .IN2(n7397), .QN(n7388) );
  NOR2X0 U8435 ( .IN1(n4383), .IN2(n6717), .QN(n7397) );
  NOR2X0 U8436 ( .IN1(DFF_1151_n1), .IN2(n4748), .QN(n7396) );
  NOR2X0 U8437 ( .IN1(n5434), .IN2(WX6950), .QN(WX7011) );
  INVX0 U8438 ( .INP(n7398), .ZN(WX686) );
  NOR2X0 U8439 ( .IN1(n7399), .IN2(n7400), .QN(n7398) );
  NAND2X0 U8440 ( .IN1(n7401), .IN2(n7402), .QN(n7400) );
  NAND2X0 U8441 ( .IN1(n7403), .IN2(n4741), .QN(n7402) );
  NAND2X0 U8442 ( .IN1(n2152), .IN2(CRC_OUT_9_10), .QN(n7401) );
  NAND2X0 U8443 ( .IN1(n7404), .IN2(n7405), .QN(n7399) );
  NAND2X0 U8444 ( .IN1(n7406), .IN2(n2153), .QN(n7405) );
  INVX0 U8445 ( .INP(n7407), .ZN(n7406) );
  NAND2X0 U8446 ( .IN1(WX524), .IN2(n4810), .QN(n7404) );
  NAND2X0 U8447 ( .IN1(n7408), .IN2(n7409), .QN(WX674) );
  NOR2X0 U8448 ( .IN1(n7410), .IN2(n7411), .QN(n7409) );
  NOR2X0 U8449 ( .IN1(n7412), .IN2(n4716), .QN(n7411) );
  NOR2X0 U8450 ( .IN1(n4765), .IN2(DFF_176_n1), .QN(n7410) );
  NOR2X0 U8451 ( .IN1(n7413), .IN2(n7414), .QN(n7408) );
  NOR2X0 U8452 ( .IN1(n4787), .IN2(n7415), .QN(n7414) );
  NOR2X0 U8453 ( .IN1(n7416), .IN2(n6023), .QN(n7413) );
  INVX0 U8454 ( .INP(WX512), .ZN(n7416) );
  NAND2X0 U8455 ( .IN1(n7417), .IN2(n7418), .QN(WX666) );
  NOR2X0 U8456 ( .IN1(n7419), .IN2(n7420), .QN(n7418) );
  NOR2X0 U8457 ( .IN1(n7421), .IN2(n4716), .QN(n7420) );
  NOR2X0 U8458 ( .IN1(n6017), .IN2(DFF_180_n1), .QN(n7419) );
  NOR2X0 U8459 ( .IN1(n7422), .IN2(n7423), .QN(n7417) );
  NOR2X0 U8460 ( .IN1(n4787), .IN2(n7424), .QN(n7423) );
  NOR2X0 U8461 ( .IN1(n7425), .IN2(n6023), .QN(n7422) );
  INVX0 U8462 ( .INP(WX504), .ZN(n7425) );
  NAND2X0 U8463 ( .IN1(n7426), .IN2(n7427), .QN(WX658) );
  NOR2X0 U8464 ( .IN1(n7428), .IN2(n7429), .QN(n7427) );
  NOR2X0 U8465 ( .IN1(n7430), .IN2(n4716), .QN(n7429) );
  NOR2X0 U8466 ( .IN1(n4765), .IN2(DFF_184_n1), .QN(n7428) );
  NOR2X0 U8467 ( .IN1(n7431), .IN2(n7432), .QN(n7426) );
  NOR2X0 U8468 ( .IN1(n4787), .IN2(n7433), .QN(n7432) );
  NOR2X0 U8469 ( .IN1(n7434), .IN2(n6023), .QN(n7431) );
  INVX0 U8470 ( .INP(WX496), .ZN(n7434) );
  NOR2X0 U8471 ( .IN1(n5434), .IN2(n7435), .QN(WX6498) );
  XOR2X1 U8472 ( .IN1(n4522), .IN2(DFF_958_n1), .Q(n7435) );
  NOR2X0 U8473 ( .IN1(n5434), .IN2(n7436), .QN(WX6496) );
  XOR2X1 U8474 ( .IN1(n4523), .IN2(DFF_957_n1), .Q(n7436) );
  NOR2X0 U8475 ( .IN1(n5434), .IN2(n7437), .QN(WX6494) );
  XOR2X1 U8476 ( .IN1(n4524), .IN2(DFF_956_n1), .Q(n7437) );
  NOR2X0 U8477 ( .IN1(n5434), .IN2(n7438), .QN(WX6492) );
  XOR2X1 U8478 ( .IN1(n4525), .IN2(DFF_955_n1), .Q(n7438) );
  NOR2X0 U8479 ( .IN1(n5434), .IN2(n7439), .QN(WX6490) );
  XOR2X1 U8480 ( .IN1(n4526), .IN2(DFF_954_n1), .Q(n7439) );
  NOR2X0 U8481 ( .IN1(n5434), .IN2(n7440), .QN(WX6488) );
  XOR2X1 U8482 ( .IN1(n4527), .IN2(DFF_953_n1), .Q(n7440) );
  NOR2X0 U8483 ( .IN1(n5434), .IN2(n7441), .QN(WX6486) );
  XOR2X1 U8484 ( .IN1(n4528), .IN2(DFF_952_n1), .Q(n7441) );
  NOR2X0 U8485 ( .IN1(n7062), .IN2(n7442), .QN(WX6484) );
  XOR2X1 U8486 ( .IN1(n4529), .IN2(DFF_951_n1), .Q(n7442) );
  INVX0 U8487 ( .INP(n6927), .ZN(n7062) );
  NOR2X0 U8488 ( .IN1(n5435), .IN2(Tj_Trigger), .QN(n6927) );
  NOR2X0 U8489 ( .IN1(n5435), .IN2(n7443), .QN(WX6482) );
  XOR2X1 U8490 ( .IN1(n4530), .IN2(DFF_950_n1), .Q(n7443) );
  NOR2X0 U8491 ( .IN1(n5435), .IN2(n7444), .QN(WX6480) );
  XOR2X1 U8492 ( .IN1(n4531), .IN2(DFF_949_n1), .Q(n7444) );
  NOR2X0 U8493 ( .IN1(n5435), .IN2(n7445), .QN(WX6478) );
  XOR2X1 U8494 ( .IN1(n4532), .IN2(DFF_948_n1), .Q(n7445) );
  NOR2X0 U8495 ( .IN1(n5435), .IN2(n7446), .QN(WX6476) );
  XOR2X1 U8496 ( .IN1(n4533), .IN2(DFF_947_n1), .Q(n7446) );
  NOR2X0 U8497 ( .IN1(n5435), .IN2(n7447), .QN(WX6474) );
  XOR2X1 U8498 ( .IN1(n4534), .IN2(DFF_946_n1), .Q(n7447) );
  NOR2X0 U8499 ( .IN1(n5435), .IN2(n7448), .QN(WX6472) );
  XOR2X1 U8500 ( .IN1(n4535), .IN2(n4699), .Q(n7448) );
  NOR2X0 U8501 ( .IN1(n5435), .IN2(n7449), .QN(WX6470) );
  XOR2X1 U8502 ( .IN1(n4536), .IN2(DFF_944_n1), .Q(n7449) );
  NOR2X0 U8503 ( .IN1(n5435), .IN2(n7450), .QN(WX6468) );
  XOR2X1 U8504 ( .IN1(DFF_943_n1), .IN2(n7451), .Q(n7450) );
  XOR2X1 U8505 ( .IN1(test_so52), .IN2(DFF_959_n1), .Q(n7451) );
  NOR2X0 U8506 ( .IN1(n5435), .IN2(n7452), .QN(WX6466) );
  XOR2X1 U8507 ( .IN1(n4537), .IN2(DFF_942_n1), .Q(n7452) );
  NOR2X0 U8508 ( .IN1(n5435), .IN2(n7453), .QN(WX6464) );
  XOR2X1 U8509 ( .IN1(n4538), .IN2(DFF_941_n1), .Q(n7453) );
  NOR2X0 U8510 ( .IN1(n5435), .IN2(n7454), .QN(WX6462) );
  XOR2X1 U8511 ( .IN1(n4539), .IN2(DFF_940_n1), .Q(n7454) );
  NOR2X0 U8512 ( .IN1(n5436), .IN2(n7455), .QN(WX6460) );
  XOR2X1 U8513 ( .IN1(n4540), .IN2(DFF_939_n1), .Q(n7455) );
  NOR2X0 U8514 ( .IN1(n5436), .IN2(n7456), .QN(WX6458) );
  XNOR2X1 U8515 ( .IN1(DFF_938_n1), .IN2(n7457), .Q(n7456) );
  XOR2X1 U8516 ( .IN1(n4399), .IN2(DFF_959_n1), .Q(n7457) );
  NOR2X0 U8517 ( .IN1(n5436), .IN2(n7458), .QN(WX6456) );
  XOR2X1 U8518 ( .IN1(n4541), .IN2(DFF_937_n1), .Q(n7458) );
  NOR2X0 U8519 ( .IN1(n5436), .IN2(n7459), .QN(WX6454) );
  XOR2X1 U8520 ( .IN1(n4542), .IN2(DFF_936_n1), .Q(n7459) );
  NOR2X0 U8521 ( .IN1(n5436), .IN2(n7460), .QN(WX6452) );
  XOR2X1 U8522 ( .IN1(n4543), .IN2(DFF_935_n1), .Q(n7460) );
  NOR2X0 U8523 ( .IN1(n5436), .IN2(n7461), .QN(WX6450) );
  XOR2X1 U8524 ( .IN1(n4544), .IN2(DFF_934_n1), .Q(n7461) );
  NOR2X0 U8525 ( .IN1(n5436), .IN2(n7462), .QN(WX6448) );
  XOR2X1 U8526 ( .IN1(n4545), .IN2(DFF_933_n1), .Q(n7462) );
  NOR2X0 U8527 ( .IN1(n5436), .IN2(n7463), .QN(WX6446) );
  XOR2X1 U8528 ( .IN1(n4546), .IN2(DFF_932_n1), .Q(n7463) );
  NOR2X0 U8529 ( .IN1(n5436), .IN2(n7464), .QN(WX6444) );
  XNOR2X1 U8530 ( .IN1(DFF_931_n1), .IN2(n7465), .Q(n7464) );
  XOR2X1 U8531 ( .IN1(n4400), .IN2(DFF_959_n1), .Q(n7465) );
  NOR2X0 U8532 ( .IN1(n5436), .IN2(n7466), .QN(WX6442) );
  XOR2X1 U8533 ( .IN1(n4547), .IN2(DFF_930_n1), .Q(n7466) );
  NOR2X0 U8534 ( .IN1(n5436), .IN2(n7467), .QN(WX6440) );
  XOR2X1 U8535 ( .IN1(n4548), .IN2(DFF_929_n1), .Q(n7467) );
  NAND2X0 U8536 ( .IN1(n7468), .IN2(n7469), .QN(WX644) );
  NOR2X0 U8537 ( .IN1(n7470), .IN2(n7471), .QN(n7469) );
  NOR2X0 U8538 ( .IN1(n7472), .IN2(n4716), .QN(n7471) );
  NOR2X0 U8539 ( .IN1(n7473), .IN2(n4776), .QN(n7470) );
  NOR2X0 U8540 ( .IN1(n7474), .IN2(n7475), .QN(n7468) );
  NOR2X0 U8541 ( .IN1(n4379), .IN2(n6717), .QN(n7475) );
  NOR2X0 U8542 ( .IN1(DFF_191_n1), .IN2(n4748), .QN(n7474) );
  NOR2X0 U8543 ( .IN1(n5436), .IN2(n7476), .QN(WX6438) );
  XOR2X1 U8544 ( .IN1(n4549), .IN2(n4698), .Q(n7476) );
  NOR2X0 U8545 ( .IN1(n5436), .IN2(n7477), .QN(WX6436) );
  XOR2X1 U8546 ( .IN1(n4413), .IN2(DFF_959_n1), .Q(n7477) );
  NOR2X0 U8547 ( .IN1(n9575), .IN2(n5346), .QN(WX5910) );
  NOR2X0 U8548 ( .IN1(n9576), .IN2(n5347), .QN(WX5908) );
  NOR2X0 U8549 ( .IN1(n9577), .IN2(n5347), .QN(WX5906) );
  NOR2X0 U8550 ( .IN1(n9580), .IN2(n5347), .QN(WX5904) );
  NOR2X0 U8551 ( .IN1(n9581), .IN2(n5347), .QN(WX5902) );
  NOR2X0 U8552 ( .IN1(n9584), .IN2(n5347), .QN(WX5900) );
  NOR2X0 U8553 ( .IN1(n5437), .IN2(n4708), .QN(WX5898) );
  NOR2X0 U8554 ( .IN1(n9585), .IN2(n5347), .QN(WX5896) );
  NOR2X0 U8555 ( .IN1(n9586), .IN2(n5347), .QN(WX5894) );
  NOR2X0 U8556 ( .IN1(n9587), .IN2(n5347), .QN(WX5892) );
  NOR2X0 U8557 ( .IN1(n9588), .IN2(n5347), .QN(WX5890) );
  NOR2X0 U8558 ( .IN1(n9589), .IN2(n5347), .QN(WX5888) );
  NOR2X0 U8559 ( .IN1(n9590), .IN2(n5347), .QN(WX5886) );
  NOR2X0 U8560 ( .IN1(n9591), .IN2(n5347), .QN(WX5884) );
  NOR2X0 U8561 ( .IN1(n9592), .IN2(n5348), .QN(WX5882) );
  NOR2X0 U8562 ( .IN1(n9593), .IN2(n5412), .QN(WX5880) );
  NAND2X0 U8563 ( .IN1(n7478), .IN2(n7479), .QN(WX5878) );
  NOR2X0 U8564 ( .IN1(n7480), .IN2(n7481), .QN(n7479) );
  NOR2X0 U8565 ( .IN1(n7482), .IN2(n4716), .QN(n7481) );
  NOR2X0 U8566 ( .IN1(n7098), .IN2(n4776), .QN(n7480) );
  XOR2X1 U8567 ( .IN1(n7483), .IN2(n7484), .Q(n7098) );
  XOR2X1 U8568 ( .IN1(n9524), .IN2(n4412), .Q(n7484) );
  XOR2X1 U8569 ( .IN1(WX7172), .IN2(n4234), .Q(n7483) );
  NOR2X0 U8570 ( .IN1(n7485), .IN2(n7486), .QN(n7478) );
  NOR2X0 U8571 ( .IN1(n4764), .IN2(n4698), .QN(n7486) );
  NOR2X0 U8572 ( .IN1(n4789), .IN2(n6129), .QN(n7485) );
  NAND2X0 U8573 ( .IN1(n5312), .IN2(n8496), .QN(n6129) );
  NAND2X0 U8574 ( .IN1(n7487), .IN2(n7488), .QN(WX5876) );
  NOR2X0 U8575 ( .IN1(n7489), .IN2(n7490), .QN(n7488) );
  NOR2X0 U8576 ( .IN1(n4732), .IN2(n7491), .QN(n7490) );
  NOR2X0 U8577 ( .IN1(n7107), .IN2(n4776), .QN(n7489) );
  XOR2X1 U8578 ( .IN1(n7492), .IN2(n7493), .Q(n7107) );
  XOR2X1 U8579 ( .IN1(n9525), .IN2(n4521), .Q(n7493) );
  XOR2X1 U8580 ( .IN1(WX7170), .IN2(n4236), .Q(n7492) );
  NOR2X0 U8581 ( .IN1(n7494), .IN2(n7495), .QN(n7487) );
  NOR2X0 U8582 ( .IN1(DFF_929_n1), .IN2(n4748), .QN(n7495) );
  NOR2X0 U8583 ( .IN1(n4789), .IN2(n6130), .QN(n7494) );
  NAND2X0 U8584 ( .IN1(n5314), .IN2(n8497), .QN(n6130) );
  NAND2X0 U8585 ( .IN1(n7496), .IN2(n7497), .QN(WX5874) );
  NOR2X0 U8586 ( .IN1(n7498), .IN2(n7499), .QN(n7497) );
  NOR2X0 U8587 ( .IN1(n7500), .IN2(n4716), .QN(n7499) );
  NOR2X0 U8588 ( .IN1(n7116), .IN2(n4776), .QN(n7498) );
  XOR2X1 U8589 ( .IN1(n7501), .IN2(n7502), .Q(n7116) );
  XOR2X1 U8590 ( .IN1(n9526), .IN2(n4520), .Q(n7502) );
  XOR2X1 U8591 ( .IN1(WX7168), .IN2(n4238), .Q(n7501) );
  NOR2X0 U8592 ( .IN1(n7503), .IN2(n7504), .QN(n7496) );
  NOR2X0 U8593 ( .IN1(DFF_930_n1), .IN2(n4748), .QN(n7504) );
  NOR2X0 U8594 ( .IN1(n4789), .IN2(n6131), .QN(n7503) );
  NAND2X0 U8595 ( .IN1(n5314), .IN2(n8498), .QN(n6131) );
  NAND2X0 U8596 ( .IN1(n7505), .IN2(n7506), .QN(WX5872) );
  NOR2X0 U8597 ( .IN1(n7507), .IN2(n7508), .QN(n7506) );
  NOR2X0 U8598 ( .IN1(n4731), .IN2(n7509), .QN(n7508) );
  NOR2X0 U8599 ( .IN1(n7125), .IN2(n4776), .QN(n7507) );
  XOR2X1 U8600 ( .IN1(n7510), .IN2(n7511), .Q(n7125) );
  XOR2X1 U8601 ( .IN1(n9527), .IN2(n4519), .Q(n7511) );
  XOR2X1 U8602 ( .IN1(WX7166), .IN2(n4240), .Q(n7510) );
  NOR2X0 U8603 ( .IN1(n7512), .IN2(n7513), .QN(n7505) );
  NOR2X0 U8604 ( .IN1(DFF_931_n1), .IN2(n4748), .QN(n7513) );
  NOR2X0 U8605 ( .IN1(n4789), .IN2(n6132), .QN(n7512) );
  NAND2X0 U8606 ( .IN1(n5314), .IN2(n8499), .QN(n6132) );
  NAND2X0 U8607 ( .IN1(n7514), .IN2(n7515), .QN(WX5870) );
  NOR2X0 U8608 ( .IN1(n7516), .IN2(n7517), .QN(n7515) );
  NOR2X0 U8609 ( .IN1(n7518), .IN2(n4716), .QN(n7517) );
  NOR2X0 U8610 ( .IN1(n4788), .IN2(n7134), .QN(n7516) );
  XNOR2X1 U8611 ( .IN1(n7519), .IN2(n7520), .Q(n7134) );
  XOR2X1 U8612 ( .IN1(test_so64), .IN2(n9528), .Q(n7520) );
  XOR2X1 U8613 ( .IN1(WX7164), .IN2(n4242), .Q(n7519) );
  NOR2X0 U8614 ( .IN1(n7521), .IN2(n7522), .QN(n7514) );
  NOR2X0 U8615 ( .IN1(DFF_932_n1), .IN2(n4748), .QN(n7522) );
  NOR2X0 U8616 ( .IN1(n6023), .IN2(n6133), .QN(n7521) );
  NAND2X0 U8617 ( .IN1(n5314), .IN2(n8500), .QN(n6133) );
  NAND2X0 U8618 ( .IN1(n7523), .IN2(n7524), .QN(WX5868) );
  NOR2X0 U8619 ( .IN1(n7525), .IN2(n7526), .QN(n7524) );
  NOR2X0 U8620 ( .IN1(n4732), .IN2(n7527), .QN(n7526) );
  NOR2X0 U8621 ( .IN1(n7143), .IN2(n4776), .QN(n7525) );
  XOR2X1 U8622 ( .IN1(n7528), .IN2(n7529), .Q(n7143) );
  XOR2X1 U8623 ( .IN1(n9529), .IN2(n4518), .Q(n7529) );
  XOR2X1 U8624 ( .IN1(WX7162), .IN2(n4244), .Q(n7528) );
  NOR2X0 U8625 ( .IN1(n7530), .IN2(n7531), .QN(n7523) );
  NOR2X0 U8626 ( .IN1(DFF_933_n1), .IN2(n4748), .QN(n7531) );
  NOR2X0 U8627 ( .IN1(n4789), .IN2(n6134), .QN(n7530) );
  NAND2X0 U8628 ( .IN1(n5313), .IN2(n8501), .QN(n6134) );
  NAND2X0 U8629 ( .IN1(n7532), .IN2(n7533), .QN(WX5866) );
  NOR2X0 U8630 ( .IN1(n7534), .IN2(n7535), .QN(n7533) );
  NOR2X0 U8631 ( .IN1(n7536), .IN2(n4716), .QN(n7535) );
  NOR2X0 U8632 ( .IN1(n4788), .IN2(n7152), .QN(n7534) );
  XNOR2X1 U8633 ( .IN1(n7537), .IN2(n7538), .Q(n7152) );
  XOR2X1 U8634 ( .IN1(test_so62), .IN2(n9530), .Q(n7538) );
  XOR2X1 U8635 ( .IN1(WX7160), .IN2(n4517), .Q(n7537) );
  NOR2X0 U8636 ( .IN1(n7539), .IN2(n7540), .QN(n7532) );
  NOR2X0 U8637 ( .IN1(DFF_934_n1), .IN2(n4747), .QN(n7540) );
  NOR2X0 U8638 ( .IN1(n6023), .IN2(n6144), .QN(n7539) );
  NAND2X0 U8639 ( .IN1(n5313), .IN2(n8502), .QN(n6144) );
  NAND2X0 U8640 ( .IN1(n7541), .IN2(n7542), .QN(WX5864) );
  NOR2X0 U8641 ( .IN1(n7543), .IN2(n7544), .QN(n7542) );
  NOR2X0 U8642 ( .IN1(n7545), .IN2(n4716), .QN(n7544) );
  NOR2X0 U8643 ( .IN1(n7161), .IN2(n4776), .QN(n7543) );
  XOR2X1 U8644 ( .IN1(n7546), .IN2(n7547), .Q(n7161) );
  XOR2X1 U8645 ( .IN1(n9531), .IN2(n4516), .Q(n7547) );
  XOR2X1 U8646 ( .IN1(WX7158), .IN2(n4247), .Q(n7546) );
  NOR2X0 U8647 ( .IN1(n7548), .IN2(n7549), .QN(n7541) );
  NOR2X0 U8648 ( .IN1(DFF_935_n1), .IN2(n4747), .QN(n7549) );
  NOR2X0 U8649 ( .IN1(n6023), .IN2(n6145), .QN(n7548) );
  NAND2X0 U8650 ( .IN1(test_so45), .IN2(n5323), .QN(n6145) );
  NAND2X0 U8651 ( .IN1(n7550), .IN2(n7551), .QN(WX5862) );
  NOR2X0 U8652 ( .IN1(n7552), .IN2(n7553), .QN(n7551) );
  NOR2X0 U8653 ( .IN1(n7554), .IN2(n4716), .QN(n7553) );
  NOR2X0 U8654 ( .IN1(n4788), .IN2(n7170), .QN(n7552) );
  XNOR2X1 U8655 ( .IN1(n7555), .IN2(n7556), .Q(n7170) );
  XOR2X1 U8656 ( .IN1(test_so60), .IN2(n9532), .Q(n7556) );
  XOR2X1 U8657 ( .IN1(WX7156), .IN2(n4515), .Q(n7555) );
  NOR2X0 U8658 ( .IN1(n7557), .IN2(n7558), .QN(n7550) );
  NOR2X0 U8659 ( .IN1(DFF_936_n1), .IN2(n4747), .QN(n7558) );
  NOR2X0 U8660 ( .IN1(n4798), .IN2(n6146), .QN(n7557) );
  NAND2X0 U8661 ( .IN1(n5313), .IN2(n8505), .QN(n6146) );
  NAND2X0 U8662 ( .IN1(n7559), .IN2(n7560), .QN(WX5860) );
  NOR2X0 U8663 ( .IN1(n7561), .IN2(n7562), .QN(n7560) );
  NOR2X0 U8664 ( .IN1(n7563), .IN2(n4716), .QN(n7562) );
  NOR2X0 U8665 ( .IN1(n7179), .IN2(n4776), .QN(n7561) );
  XOR2X1 U8666 ( .IN1(n7564), .IN2(n7565), .Q(n7179) );
  XOR2X1 U8667 ( .IN1(n9533), .IN2(n4514), .Q(n7565) );
  XOR2X1 U8668 ( .IN1(WX7154), .IN2(n4250), .Q(n7564) );
  NOR2X0 U8669 ( .IN1(n7566), .IN2(n7567), .QN(n7559) );
  NOR2X0 U8670 ( .IN1(DFF_937_n1), .IN2(n4747), .QN(n7567) );
  NOR2X0 U8671 ( .IN1(n6023), .IN2(n6147), .QN(n7566) );
  NAND2X0 U8672 ( .IN1(n5313), .IN2(n8506), .QN(n6147) );
  NAND2X0 U8673 ( .IN1(n7568), .IN2(n7569), .QN(WX5858) );
  NOR2X0 U8674 ( .IN1(n7570), .IN2(n7571), .QN(n7569) );
  NOR2X0 U8675 ( .IN1(n7572), .IN2(n4716), .QN(n7571) );
  NOR2X0 U8676 ( .IN1(n4788), .IN2(n7188), .QN(n7570) );
  XNOR2X1 U8677 ( .IN1(n7573), .IN2(n7574), .Q(n7188) );
  XOR2X1 U8678 ( .IN1(test_so58), .IN2(n9534), .Q(n7574) );
  XOR2X1 U8679 ( .IN1(WX7280), .IN2(n4513), .Q(n7573) );
  NOR2X0 U8680 ( .IN1(n7575), .IN2(n7576), .QN(n7568) );
  NOR2X0 U8681 ( .IN1(DFF_938_n1), .IN2(n4747), .QN(n7576) );
  NOR2X0 U8682 ( .IN1(n4803), .IN2(n6148), .QN(n7575) );
  NAND2X0 U8683 ( .IN1(n5313), .IN2(n8507), .QN(n6148) );
  NAND2X0 U8684 ( .IN1(n7577), .IN2(n7578), .QN(WX5856) );
  NOR2X0 U8685 ( .IN1(n7579), .IN2(n7580), .QN(n7578) );
  NOR2X0 U8686 ( .IN1(n7581), .IN2(n4715), .QN(n7580) );
  NOR2X0 U8687 ( .IN1(n7197), .IN2(n4776), .QN(n7579) );
  XOR2X1 U8688 ( .IN1(n7582), .IN2(n7583), .Q(n7197) );
  XOR2X1 U8689 ( .IN1(n9535), .IN2(n4398), .Q(n7583) );
  XOR2X1 U8690 ( .IN1(WX7150), .IN2(n4253), .Q(n7582) );
  NOR2X0 U8691 ( .IN1(n7584), .IN2(n7585), .QN(n7577) );
  NOR2X0 U8692 ( .IN1(DFF_939_n1), .IN2(n4747), .QN(n7585) );
  NOR2X0 U8693 ( .IN1(n4792), .IN2(n6149), .QN(n7584) );
  NAND2X0 U8694 ( .IN1(n5312), .IN2(n8508), .QN(n6149) );
  NAND2X0 U8695 ( .IN1(n7586), .IN2(n7587), .QN(WX5854) );
  NOR2X0 U8696 ( .IN1(n7588), .IN2(n7589), .QN(n7587) );
  NOR2X0 U8697 ( .IN1(n7590), .IN2(n4715), .QN(n7589) );
  NOR2X0 U8698 ( .IN1(n7206), .IN2(n4777), .QN(n7588) );
  XOR2X1 U8699 ( .IN1(n7591), .IN2(n7592), .Q(n7206) );
  XOR2X1 U8700 ( .IN1(n9536), .IN2(n4512), .Q(n7592) );
  XOR2X1 U8701 ( .IN1(WX7148), .IN2(n4255), .Q(n7591) );
  NOR2X0 U8702 ( .IN1(n7593), .IN2(n7594), .QN(n7586) );
  NOR2X0 U8703 ( .IN1(DFF_940_n1), .IN2(n4747), .QN(n7594) );
  NOR2X0 U8704 ( .IN1(n6023), .IN2(n6150), .QN(n7593) );
  NAND2X0 U8705 ( .IN1(n5312), .IN2(n8509), .QN(n6150) );
  NAND2X0 U8706 ( .IN1(n7595), .IN2(n7596), .QN(WX5852) );
  NOR2X0 U8707 ( .IN1(n7597), .IN2(n7598), .QN(n7596) );
  NOR2X0 U8708 ( .IN1(n7599), .IN2(n4715), .QN(n7598) );
  NOR2X0 U8709 ( .IN1(n7215), .IN2(n4777), .QN(n7597) );
  XOR2X1 U8710 ( .IN1(n7600), .IN2(n7601), .Q(n7215) );
  XOR2X1 U8711 ( .IN1(n9537), .IN2(n4511), .Q(n7601) );
  XOR2X1 U8712 ( .IN1(WX7146), .IN2(n4257), .Q(n7600) );
  NOR2X0 U8713 ( .IN1(n7602), .IN2(n7603), .QN(n7595) );
  NOR2X0 U8714 ( .IN1(DFF_941_n1), .IN2(n4747), .QN(n7603) );
  NOR2X0 U8715 ( .IN1(n6023), .IN2(n6151), .QN(n7602) );
  NAND2X0 U8716 ( .IN1(n5311), .IN2(n8510), .QN(n6151) );
  NAND2X0 U8717 ( .IN1(n7604), .IN2(n7605), .QN(WX5850) );
  NOR2X0 U8718 ( .IN1(n7606), .IN2(n7607), .QN(n7605) );
  NOR2X0 U8719 ( .IN1(n7608), .IN2(n4715), .QN(n7607) );
  NOR2X0 U8720 ( .IN1(n7224), .IN2(n4777), .QN(n7606) );
  XOR2X1 U8721 ( .IN1(n7609), .IN2(n7610), .Q(n7224) );
  XOR2X1 U8722 ( .IN1(n9538), .IN2(n4510), .Q(n7610) );
  XOR2X1 U8723 ( .IN1(WX7144), .IN2(n4259), .Q(n7609) );
  NOR2X0 U8724 ( .IN1(n7611), .IN2(n7612), .QN(n7604) );
  NOR2X0 U8725 ( .IN1(DFF_942_n1), .IN2(n4747), .QN(n7612) );
  NOR2X0 U8726 ( .IN1(n4804), .IN2(n6152), .QN(n7611) );
  NAND2X0 U8727 ( .IN1(n5312), .IN2(n8511), .QN(n6152) );
  NAND2X0 U8728 ( .IN1(n7613), .IN2(n7614), .QN(WX5848) );
  NOR2X0 U8729 ( .IN1(n7615), .IN2(n7616), .QN(n7614) );
  NOR2X0 U8730 ( .IN1(n7617), .IN2(n4715), .QN(n7616) );
  NOR2X0 U8731 ( .IN1(n7233), .IN2(n4777), .QN(n7615) );
  XOR2X1 U8732 ( .IN1(n7618), .IN2(n7619), .Q(n7233) );
  XOR2X1 U8733 ( .IN1(n9539), .IN2(n4509), .Q(n7619) );
  XOR2X1 U8734 ( .IN1(WX7142), .IN2(n4261), .Q(n7618) );
  NOR2X0 U8735 ( .IN1(n7620), .IN2(n7621), .QN(n7613) );
  NOR2X0 U8736 ( .IN1(DFF_943_n1), .IN2(n4747), .QN(n7621) );
  NOR2X0 U8737 ( .IN1(n4804), .IN2(n6153), .QN(n7620) );
  NAND2X0 U8738 ( .IN1(n5312), .IN2(n8512), .QN(n6153) );
  NAND2X0 U8739 ( .IN1(n7622), .IN2(n7623), .QN(WX5846) );
  NOR2X0 U8740 ( .IN1(n7624), .IN2(n7625), .QN(n7623) );
  NOR2X0 U8741 ( .IN1(n4732), .IN2(n7626), .QN(n7625) );
  NOR2X0 U8742 ( .IN1(n7242), .IN2(n4777), .QN(n7624) );
  XOR2X1 U8743 ( .IN1(n7627), .IN2(n7628), .Q(n7242) );
  XOR2X1 U8744 ( .IN1(n4078), .IN2(n5251), .Q(n7628) );
  XOR2X1 U8745 ( .IN1(n7629), .IN2(n4397), .Q(n7627) );
  XOR2X1 U8746 ( .IN1(WX7268), .IN2(n9540), .Q(n7629) );
  NOR2X0 U8747 ( .IN1(n7630), .IN2(n7631), .QN(n7622) );
  NOR2X0 U8748 ( .IN1(DFF_944_n1), .IN2(n4747), .QN(n7631) );
  NOR2X0 U8749 ( .IN1(n4804), .IN2(n6163), .QN(n7630) );
  NAND2X0 U8750 ( .IN1(n5312), .IN2(n8513), .QN(n6163) );
  NAND2X0 U8751 ( .IN1(n7632), .IN2(n7633), .QN(WX5844) );
  NOR2X0 U8752 ( .IN1(n7634), .IN2(n7635), .QN(n7633) );
  NOR2X0 U8753 ( .IN1(n7636), .IN2(n4715), .QN(n7635) );
  NOR2X0 U8754 ( .IN1(n7252), .IN2(n4777), .QN(n7634) );
  XOR2X1 U8755 ( .IN1(n7637), .IN2(n7638), .Q(n7252) );
  XOR2X1 U8756 ( .IN1(n4079), .IN2(n5251), .Q(n7638) );
  XOR2X1 U8757 ( .IN1(n7639), .IN2(n4508), .Q(n7637) );
  XOR2X1 U8758 ( .IN1(WX7266), .IN2(n9541), .Q(n7639) );
  NOR2X0 U8759 ( .IN1(n7640), .IN2(n7641), .QN(n7632) );
  NOR2X0 U8760 ( .IN1(n4765), .IN2(n4699), .QN(n7641) );
  NOR2X0 U8761 ( .IN1(n4804), .IN2(n6164), .QN(n7640) );
  NAND2X0 U8762 ( .IN1(n5311), .IN2(n8514), .QN(n6164) );
  NAND2X0 U8763 ( .IN1(n7642), .IN2(n7643), .QN(WX5842) );
  NOR2X0 U8764 ( .IN1(n7644), .IN2(n7645), .QN(n7643) );
  NOR2X0 U8765 ( .IN1(n4732), .IN2(n7646), .QN(n7645) );
  NOR2X0 U8766 ( .IN1(n7262), .IN2(n4777), .QN(n7644) );
  XOR2X1 U8767 ( .IN1(n7647), .IN2(n7648), .Q(n7262) );
  XOR2X1 U8768 ( .IN1(n4080), .IN2(n5251), .Q(n7648) );
  XOR2X1 U8769 ( .IN1(n7649), .IN2(n4507), .Q(n7647) );
  XOR2X1 U8770 ( .IN1(WX7264), .IN2(n9542), .Q(n7649) );
  NOR2X0 U8771 ( .IN1(n7650), .IN2(n7651), .QN(n7642) );
  NOR2X0 U8772 ( .IN1(DFF_946_n1), .IN2(n4751), .QN(n7651) );
  NOR2X0 U8773 ( .IN1(n4804), .IN2(n6165), .QN(n7650) );
  NAND2X0 U8774 ( .IN1(n5311), .IN2(n8515), .QN(n6165) );
  NAND2X0 U8775 ( .IN1(n7652), .IN2(n7653), .QN(WX5840) );
  NOR2X0 U8776 ( .IN1(n7654), .IN2(n7655), .QN(n7653) );
  NOR2X0 U8777 ( .IN1(n7656), .IN2(n4715), .QN(n7655) );
  NOR2X0 U8778 ( .IN1(n7272), .IN2(n4777), .QN(n7654) );
  XOR2X1 U8779 ( .IN1(n7657), .IN2(n7658), .Q(n7272) );
  XOR2X1 U8780 ( .IN1(n4081), .IN2(n5251), .Q(n7658) );
  XOR2X1 U8781 ( .IN1(n7659), .IN2(n4506), .Q(n7657) );
  XOR2X1 U8782 ( .IN1(WX7262), .IN2(n9543), .Q(n7659) );
  NOR2X0 U8783 ( .IN1(n7660), .IN2(n7661), .QN(n7652) );
  NOR2X0 U8784 ( .IN1(DFF_947_n1), .IN2(n4763), .QN(n7661) );
  NOR2X0 U8785 ( .IN1(n4804), .IN2(n6166), .QN(n7660) );
  NAND2X0 U8786 ( .IN1(n5311), .IN2(n8516), .QN(n6166) );
  NAND2X0 U8787 ( .IN1(n7662), .IN2(n7663), .QN(WX5838) );
  NOR2X0 U8788 ( .IN1(n7664), .IN2(n7665), .QN(n7663) );
  NOR2X0 U8789 ( .IN1(n4732), .IN2(n7666), .QN(n7665) );
  NOR2X0 U8790 ( .IN1(n7282), .IN2(n4777), .QN(n7664) );
  XOR2X1 U8791 ( .IN1(n7667), .IN2(n7668), .Q(n7282) );
  XOR2X1 U8792 ( .IN1(n4082), .IN2(n5251), .Q(n7668) );
  XOR2X1 U8793 ( .IN1(n7669), .IN2(n4505), .Q(n7667) );
  XOR2X1 U8794 ( .IN1(WX7260), .IN2(n9544), .Q(n7669) );
  NOR2X0 U8795 ( .IN1(n7670), .IN2(n7671), .QN(n7662) );
  NOR2X0 U8796 ( .IN1(DFF_948_n1), .IN2(n4764), .QN(n7671) );
  NOR2X0 U8797 ( .IN1(n4804), .IN2(n6167), .QN(n7670) );
  NAND2X0 U8798 ( .IN1(n5311), .IN2(n8517), .QN(n6167) );
  NAND2X0 U8799 ( .IN1(n7672), .IN2(n7673), .QN(WX5836) );
  NOR2X0 U8800 ( .IN1(n7674), .IN2(n7675), .QN(n7673) );
  NOR2X0 U8801 ( .IN1(n7676), .IN2(n4715), .QN(n7675) );
  NOR2X0 U8802 ( .IN1(n4788), .IN2(n7292), .QN(n7674) );
  XNOR2X1 U8803 ( .IN1(n7677), .IN2(n7678), .Q(n7292) );
  XOR2X1 U8804 ( .IN1(n4083), .IN2(n5251), .Q(n7678) );
  XOR2X1 U8805 ( .IN1(WX7194), .IN2(n7679), .Q(n7677) );
  XOR2X1 U8806 ( .IN1(test_so63), .IN2(n9545), .Q(n7679) );
  NOR2X0 U8807 ( .IN1(n7680), .IN2(n7681), .QN(n7672) );
  NOR2X0 U8808 ( .IN1(DFF_949_n1), .IN2(n4764), .QN(n7681) );
  NOR2X0 U8809 ( .IN1(n4804), .IN2(n6168), .QN(n7680) );
  NAND2X0 U8810 ( .IN1(n5310), .IN2(n8518), .QN(n6168) );
  NAND2X0 U8811 ( .IN1(n7682), .IN2(n7683), .QN(WX5834) );
  NOR2X0 U8812 ( .IN1(n7684), .IN2(n7685), .QN(n7683) );
  NOR2X0 U8813 ( .IN1(n4732), .IN2(n7686), .QN(n7685) );
  NOR2X0 U8814 ( .IN1(n7302), .IN2(n4777), .QN(n7684) );
  XOR2X1 U8815 ( .IN1(n7687), .IN2(n7688), .Q(n7302) );
  XOR2X1 U8816 ( .IN1(n4084), .IN2(n5251), .Q(n7688) );
  XOR2X1 U8817 ( .IN1(n7689), .IN2(n4504), .Q(n7687) );
  XOR2X1 U8818 ( .IN1(WX7256), .IN2(n9546), .Q(n7689) );
  NOR2X0 U8819 ( .IN1(n7690), .IN2(n7691), .QN(n7682) );
  NOR2X0 U8820 ( .IN1(DFF_950_n1), .IN2(n4764), .QN(n7691) );
  NOR2X0 U8821 ( .IN1(n4804), .IN2(n6169), .QN(n7690) );
  NAND2X0 U8822 ( .IN1(n5311), .IN2(n8519), .QN(n6169) );
  NAND2X0 U8823 ( .IN1(n7692), .IN2(n7693), .QN(WX5832) );
  NOR2X0 U8824 ( .IN1(n7694), .IN2(n7695), .QN(n7693) );
  NOR2X0 U8825 ( .IN1(n7696), .IN2(n4715), .QN(n7695) );
  NOR2X0 U8826 ( .IN1(n4788), .IN2(n7312), .QN(n7694) );
  XNOR2X1 U8827 ( .IN1(n7697), .IN2(n7698), .Q(n7312) );
  XOR2X1 U8828 ( .IN1(n4503), .IN2(n5251), .Q(n7698) );
  XOR2X1 U8829 ( .IN1(n7699), .IN2(n9549), .Q(n7697) );
  XOR2X1 U8830 ( .IN1(n9548), .IN2(n9547), .Q(n7699) );
  NOR2X0 U8831 ( .IN1(n7700), .IN2(n7701), .QN(n7692) );
  NOR2X0 U8832 ( .IN1(DFF_951_n1), .IN2(n4764), .QN(n7701) );
  NOR2X0 U8833 ( .IN1(n4804), .IN2(n6170), .QN(n7700) );
  NAND2X0 U8834 ( .IN1(n5310), .IN2(n8520), .QN(n6170) );
  NAND2X0 U8835 ( .IN1(n7702), .IN2(n7703), .QN(WX5830) );
  NOR2X0 U8836 ( .IN1(n7704), .IN2(n7705), .QN(n7703) );
  NOR2X0 U8837 ( .IN1(n7706), .IN2(n4715), .QN(n7705) );
  NOR2X0 U8838 ( .IN1(n7322), .IN2(n4777), .QN(n7704) );
  XOR2X1 U8839 ( .IN1(n7707), .IN2(n7708), .Q(n7322) );
  XOR2X1 U8840 ( .IN1(n4085), .IN2(n5251), .Q(n7708) );
  XOR2X1 U8841 ( .IN1(n7709), .IN2(n4502), .Q(n7707) );
  XOR2X1 U8842 ( .IN1(WX7252), .IN2(n9550), .Q(n7709) );
  NOR2X0 U8843 ( .IN1(n7710), .IN2(n7711), .QN(n7702) );
  NOR2X0 U8844 ( .IN1(DFF_952_n1), .IN2(n4763), .QN(n7711) );
  NOR2X0 U8845 ( .IN1(n4804), .IN2(n6171), .QN(n7710) );
  NAND2X0 U8846 ( .IN1(test_so44), .IN2(n5322), .QN(n6171) );
  NAND2X0 U8847 ( .IN1(n7712), .IN2(n7713), .QN(WX5828) );
  NOR2X0 U8848 ( .IN1(n7714), .IN2(n7715), .QN(n7713) );
  NOR2X0 U8849 ( .IN1(n7716), .IN2(n4715), .QN(n7715) );
  NOR2X0 U8850 ( .IN1(n4788), .IN2(n7332), .QN(n7714) );
  XNOR2X1 U8851 ( .IN1(n7717), .IN2(n7718), .Q(n7332) );
  XOR2X1 U8852 ( .IN1(n4501), .IN2(n5251), .Q(n7718) );
  XOR2X1 U8853 ( .IN1(n7719), .IN2(n9553), .Q(n7717) );
  XOR2X1 U8854 ( .IN1(n9552), .IN2(n9551), .Q(n7719) );
  NOR2X0 U8855 ( .IN1(n7720), .IN2(n7721), .QN(n7712) );
  NOR2X0 U8856 ( .IN1(DFF_953_n1), .IN2(n4764), .QN(n7721) );
  NOR2X0 U8857 ( .IN1(n4804), .IN2(n6172), .QN(n7720) );
  NAND2X0 U8858 ( .IN1(n5310), .IN2(n8523), .QN(n6172) );
  NAND2X0 U8859 ( .IN1(n7722), .IN2(n7723), .QN(WX5826) );
  NOR2X0 U8860 ( .IN1(n7724), .IN2(n7725), .QN(n7723) );
  NOR2X0 U8861 ( .IN1(n7726), .IN2(n4719), .QN(n7725) );
  NOR2X0 U8862 ( .IN1(n7342), .IN2(n4777), .QN(n7724) );
  XOR2X1 U8863 ( .IN1(n7727), .IN2(n7728), .Q(n7342) );
  XOR2X1 U8864 ( .IN1(n4086), .IN2(n5251), .Q(n7728) );
  XOR2X1 U8865 ( .IN1(n7729), .IN2(n4500), .Q(n7727) );
  XOR2X1 U8866 ( .IN1(WX7248), .IN2(n9554), .Q(n7729) );
  NOR2X0 U8867 ( .IN1(n7730), .IN2(n7731), .QN(n7722) );
  NOR2X0 U8868 ( .IN1(DFF_954_n1), .IN2(n4763), .QN(n7731) );
  NOR2X0 U8869 ( .IN1(n4804), .IN2(n6183), .QN(n7730) );
  NAND2X0 U8870 ( .IN1(n5310), .IN2(n8524), .QN(n6183) );
  NAND2X0 U8871 ( .IN1(n7732), .IN2(n7733), .QN(WX5824) );
  NOR2X0 U8872 ( .IN1(n7734), .IN2(n7735), .QN(n7733) );
  NOR2X0 U8873 ( .IN1(n7736), .IN2(n4726), .QN(n7735) );
  NOR2X0 U8874 ( .IN1(n4784), .IN2(n7352), .QN(n7734) );
  XNOR2X1 U8875 ( .IN1(n7737), .IN2(n7738), .Q(n7352) );
  XOR2X1 U8876 ( .IN1(n4087), .IN2(n5251), .Q(n7738) );
  XOR2X1 U8877 ( .IN1(n7739), .IN2(n4499), .Q(n7737) );
  XOR2X1 U8878 ( .IN1(WX7182), .IN2(test_so57), .Q(n7739) );
  NOR2X0 U8879 ( .IN1(n7740), .IN2(n7741), .QN(n7732) );
  NOR2X0 U8880 ( .IN1(DFF_955_n1), .IN2(n4762), .QN(n7741) );
  NOR2X0 U8881 ( .IN1(n4803), .IN2(n6184), .QN(n7740) );
  NAND2X0 U8882 ( .IN1(n5310), .IN2(n8525), .QN(n6184) );
  NAND2X0 U8883 ( .IN1(n7742), .IN2(n7743), .QN(WX5822) );
  NOR2X0 U8884 ( .IN1(n7744), .IN2(n7745), .QN(n7743) );
  NOR2X0 U8885 ( .IN1(n7746), .IN2(n4729), .QN(n7745) );
  NOR2X0 U8886 ( .IN1(n7362), .IN2(n4778), .QN(n7744) );
  XOR2X1 U8887 ( .IN1(n7747), .IN2(n7748), .Q(n7362) );
  XOR2X1 U8888 ( .IN1(n4088), .IN2(n5252), .Q(n7748) );
  XOR2X1 U8889 ( .IN1(n7749), .IN2(n4498), .Q(n7747) );
  XOR2X1 U8890 ( .IN1(WX7244), .IN2(n9555), .Q(n7749) );
  NOR2X0 U8891 ( .IN1(n7750), .IN2(n7751), .QN(n7742) );
  NOR2X0 U8892 ( .IN1(DFF_956_n1), .IN2(n4763), .QN(n7751) );
  NOR2X0 U8893 ( .IN1(n4803), .IN2(n6185), .QN(n7750) );
  NAND2X0 U8894 ( .IN1(n5310), .IN2(n8526), .QN(n6185) );
  NAND2X0 U8895 ( .IN1(n7752), .IN2(n7753), .QN(WX5820) );
  NOR2X0 U8896 ( .IN1(n7754), .IN2(n7755), .QN(n7753) );
  NOR2X0 U8897 ( .IN1(n7756), .IN2(n4728), .QN(n7755) );
  NOR2X0 U8898 ( .IN1(n7372), .IN2(n4778), .QN(n7754) );
  XOR2X1 U8899 ( .IN1(n7757), .IN2(n7758), .Q(n7372) );
  XOR2X1 U8900 ( .IN1(n4089), .IN2(n5252), .Q(n7758) );
  XOR2X1 U8901 ( .IN1(n7759), .IN2(n4497), .Q(n7757) );
  XOR2X1 U8902 ( .IN1(WX7242), .IN2(n9556), .Q(n7759) );
  NOR2X0 U8903 ( .IN1(n7760), .IN2(n7761), .QN(n7752) );
  NOR2X0 U8904 ( .IN1(DFF_957_n1), .IN2(n4763), .QN(n7761) );
  NOR2X0 U8905 ( .IN1(n4803), .IN2(n6186), .QN(n7760) );
  NAND2X0 U8906 ( .IN1(n5309), .IN2(n8527), .QN(n6186) );
  NAND2X0 U8907 ( .IN1(n7762), .IN2(n7763), .QN(WX5818) );
  NOR2X0 U8908 ( .IN1(n7764), .IN2(n7765), .QN(n7763) );
  NOR2X0 U8909 ( .IN1(n7766), .IN2(n4727), .QN(n7765) );
  NOR2X0 U8910 ( .IN1(n7382), .IN2(n4778), .QN(n7764) );
  XOR2X1 U8911 ( .IN1(n7767), .IN2(n7768), .Q(n7382) );
  XOR2X1 U8912 ( .IN1(n4090), .IN2(n5252), .Q(n7768) );
  XOR2X1 U8913 ( .IN1(n7769), .IN2(n4496), .Q(n7767) );
  XOR2X1 U8914 ( .IN1(WX7240), .IN2(n9557), .Q(n7769) );
  NOR2X0 U8915 ( .IN1(n7770), .IN2(n7771), .QN(n7762) );
  NOR2X0 U8916 ( .IN1(DFF_958_n1), .IN2(n4763), .QN(n7771) );
  NOR2X0 U8917 ( .IN1(n4803), .IN2(n6187), .QN(n7770) );
  NAND2X0 U8918 ( .IN1(n5309), .IN2(n8528), .QN(n6187) );
  NAND2X0 U8919 ( .IN1(n7772), .IN2(n7773), .QN(WX5816) );
  NOR2X0 U8920 ( .IN1(n7774), .IN2(n7775), .QN(n7773) );
  NOR2X0 U8921 ( .IN1(n7776), .IN2(n4728), .QN(n7775) );
  NOR2X0 U8922 ( .IN1(n7392), .IN2(n4778), .QN(n7774) );
  XOR2X1 U8923 ( .IN1(n7777), .IN2(n7778), .Q(n7392) );
  XOR2X1 U8924 ( .IN1(n4034), .IN2(n5252), .Q(n7778) );
  XOR2X1 U8925 ( .IN1(n7779), .IN2(n4495), .Q(n7777) );
  XOR2X1 U8926 ( .IN1(WX7238), .IN2(n9558), .Q(n7779) );
  NOR2X0 U8927 ( .IN1(n7780), .IN2(n7781), .QN(n7772) );
  NOR2X0 U8928 ( .IN1(n4384), .IN2(n6717), .QN(n7781) );
  NOR2X0 U8929 ( .IN1(DFF_959_n1), .IN2(n4764), .QN(n7780) );
  NOR2X0 U8930 ( .IN1(n5437), .IN2(WX5657), .QN(WX5718) );
  NOR2X0 U8931 ( .IN1(n5437), .IN2(WX485), .QN(WX546) );
  NOR2X0 U8932 ( .IN1(n5437), .IN2(n7782), .QN(WX5205) );
  XOR2X1 U8933 ( .IN1(n4550), .IN2(DFF_766_n1), .Q(n7782) );
  NOR2X0 U8934 ( .IN1(n5437), .IN2(n7783), .QN(WX5203) );
  XOR2X1 U8935 ( .IN1(n4551), .IN2(DFF_765_n1), .Q(n7783) );
  NOR2X0 U8936 ( .IN1(n5437), .IN2(n7784), .QN(WX5201) );
  XOR2X1 U8937 ( .IN1(n4552), .IN2(DFF_764_n1), .Q(n7784) );
  NOR2X0 U8938 ( .IN1(n5437), .IN2(n7785), .QN(WX5199) );
  XNOR2X1 U8939 ( .IN1(DFF_763_n1), .IN2(test_so40), .Q(n7785) );
  NOR2X0 U8940 ( .IN1(n5437), .IN2(n7786), .QN(WX5197) );
  XOR2X1 U8941 ( .IN1(n4553), .IN2(DFF_762_n1), .Q(n7786) );
  NOR2X0 U8942 ( .IN1(n5437), .IN2(n7787), .QN(WX5195) );
  XOR2X1 U8943 ( .IN1(n4554), .IN2(DFF_761_n1), .Q(n7787) );
  NOR2X0 U8944 ( .IN1(n5437), .IN2(n7788), .QN(WX5193) );
  XOR2X1 U8945 ( .IN1(n4555), .IN2(DFF_760_n1), .Q(n7788) );
  NOR2X0 U8946 ( .IN1(n5437), .IN2(n7789), .QN(WX5191) );
  XOR2X1 U8947 ( .IN1(n4556), .IN2(DFF_759_n1), .Q(n7789) );
  NOR2X0 U8948 ( .IN1(n5437), .IN2(n7790), .QN(WX5189) );
  XOR2X1 U8949 ( .IN1(n4557), .IN2(n4701), .Q(n7790) );
  NOR2X0 U8950 ( .IN1(n5437), .IN2(n7791), .QN(WX5187) );
  XOR2X1 U8951 ( .IN1(n4558), .IN2(DFF_757_n1), .Q(n7791) );
  NOR2X0 U8952 ( .IN1(n5438), .IN2(n7792), .QN(WX5185) );
  XOR2X1 U8953 ( .IN1(n4559), .IN2(DFF_756_n1), .Q(n7792) );
  NOR2X0 U8954 ( .IN1(n5438), .IN2(n7793), .QN(WX5183) );
  XOR2X1 U8955 ( .IN1(n4560), .IN2(DFF_755_n1), .Q(n7793) );
  NOR2X0 U8956 ( .IN1(n5438), .IN2(n7794), .QN(WX5181) );
  XOR2X1 U8957 ( .IN1(n4561), .IN2(DFF_754_n1), .Q(n7794) );
  NOR2X0 U8958 ( .IN1(n5438), .IN2(n7795), .QN(WX5179) );
  XOR2X1 U8959 ( .IN1(n4562), .IN2(DFF_753_n1), .Q(n7795) );
  NOR2X0 U8960 ( .IN1(n5438), .IN2(n7796), .QN(WX5177) );
  XOR2X1 U8961 ( .IN1(n4563), .IN2(DFF_752_n1), .Q(n7796) );
  NOR2X0 U8962 ( .IN1(n5438), .IN2(n7797), .QN(WX5175) );
  XNOR2X1 U8963 ( .IN1(DFF_751_n1), .IN2(n7798), .Q(n7797) );
  XOR2X1 U8964 ( .IN1(n4401), .IN2(DFF_767_n1), .Q(n7798) );
  NOR2X0 U8965 ( .IN1(n5438), .IN2(n7799), .QN(WX5173) );
  XOR2X1 U8966 ( .IN1(n4564), .IN2(DFF_750_n1), .Q(n7799) );
  NOR2X0 U8967 ( .IN1(n5438), .IN2(n7800), .QN(WX5171) );
  XOR2X1 U8968 ( .IN1(n4565), .IN2(DFF_749_n1), .Q(n7800) );
  NOR2X0 U8969 ( .IN1(n5438), .IN2(n7801), .QN(WX5169) );
  XOR2X1 U8970 ( .IN1(n4566), .IN2(DFF_748_n1), .Q(n7801) );
  NOR2X0 U8971 ( .IN1(n5438), .IN2(n7802), .QN(WX5167) );
  XOR2X1 U8972 ( .IN1(n4567), .IN2(DFF_747_n1), .Q(n7802) );
  NOR2X0 U8973 ( .IN1(n5438), .IN2(n7803), .QN(WX5165) );
  XOR2X1 U8974 ( .IN1(DFF_746_n1), .IN2(n7804), .Q(n7803) );
  XOR2X1 U8975 ( .IN1(test_so41), .IN2(DFF_767_n1), .Q(n7804) );
  NOR2X0 U8976 ( .IN1(n5438), .IN2(n7805), .QN(WX5163) );
  XOR2X1 U8977 ( .IN1(n4568), .IN2(DFF_745_n1), .Q(n7805) );
  NOR2X0 U8978 ( .IN1(n5438), .IN2(n7806), .QN(WX5161) );
  XOR2X1 U8979 ( .IN1(n4569), .IN2(DFF_744_n1), .Q(n7806) );
  NOR2X0 U8980 ( .IN1(n5439), .IN2(n7807), .QN(WX5159) );
  XOR2X1 U8981 ( .IN1(n4570), .IN2(DFF_743_n1), .Q(n7807) );
  NOR2X0 U8982 ( .IN1(n5439), .IN2(n7808), .QN(WX5157) );
  XOR2X1 U8983 ( .IN1(n4571), .IN2(DFF_742_n1), .Q(n7808) );
  NOR2X0 U8984 ( .IN1(n5439), .IN2(n7809), .QN(WX5155) );
  XOR2X1 U8985 ( .IN1(n4572), .IN2(n4700), .Q(n7809) );
  NOR2X0 U8986 ( .IN1(n5439), .IN2(n7810), .QN(WX5153) );
  XOR2X1 U8987 ( .IN1(n4573), .IN2(DFF_740_n1), .Q(n7810) );
  NOR2X0 U8988 ( .IN1(n5439), .IN2(n7811), .QN(WX5151) );
  XNOR2X1 U8989 ( .IN1(DFF_739_n1), .IN2(n7812), .Q(n7811) );
  XOR2X1 U8990 ( .IN1(n4402), .IN2(DFF_767_n1), .Q(n7812) );
  NOR2X0 U8991 ( .IN1(n5439), .IN2(n7813), .QN(WX5149) );
  XOR2X1 U8992 ( .IN1(n4574), .IN2(DFF_738_n1), .Q(n7813) );
  NOR2X0 U8993 ( .IN1(n5439), .IN2(n7814), .QN(WX5147) );
  XOR2X1 U8994 ( .IN1(n4575), .IN2(DFF_737_n1), .Q(n7814) );
  NOR2X0 U8995 ( .IN1(n5439), .IN2(n7815), .QN(WX5145) );
  XOR2X1 U8996 ( .IN1(n4576), .IN2(DFF_736_n1), .Q(n7815) );
  NOR2X0 U8997 ( .IN1(n5439), .IN2(n7816), .QN(WX5143) );
  XOR2X1 U8998 ( .IN1(n4414), .IN2(DFF_767_n1), .Q(n7816) );
  NOR2X0 U8999 ( .IN1(n9610), .IN2(n5411), .QN(WX4617) );
  NOR2X0 U9000 ( .IN1(n5439), .IN2(n4709), .QN(WX4615) );
  NOR2X0 U9001 ( .IN1(n9611), .IN2(n5410), .QN(WX4613) );
  NOR2X0 U9002 ( .IN1(n9612), .IN2(n5352), .QN(WX4611) );
  NOR2X0 U9003 ( .IN1(n9613), .IN2(n5352), .QN(WX4609) );
  NOR2X0 U9004 ( .IN1(n9614), .IN2(n5352), .QN(WX4607) );
  NOR2X0 U9005 ( .IN1(n9615), .IN2(n5352), .QN(WX4605) );
  NOR2X0 U9006 ( .IN1(n9616), .IN2(n5352), .QN(WX4603) );
  NOR2X0 U9007 ( .IN1(n9617), .IN2(n5352), .QN(WX4601) );
  NOR2X0 U9008 ( .IN1(n9618), .IN2(n5352), .QN(WX4599) );
  NOR2X0 U9009 ( .IN1(n9619), .IN2(n5352), .QN(WX4597) );
  NOR2X0 U9010 ( .IN1(n9620), .IN2(n5352), .QN(WX4595) );
  NOR2X0 U9011 ( .IN1(n9621), .IN2(n5352), .QN(WX4593) );
  NOR2X0 U9012 ( .IN1(n9622), .IN2(n5352), .QN(WX4591) );
  NOR2X0 U9013 ( .IN1(n9623), .IN2(n5352), .QN(WX4589) );
  NOR2X0 U9014 ( .IN1(n9626), .IN2(n5351), .QN(WX4587) );
  NAND2X0 U9015 ( .IN1(n7817), .IN2(n7818), .QN(WX4585) );
  NOR2X0 U9016 ( .IN1(n7819), .IN2(n7820), .QN(n7818) );
  NOR2X0 U9017 ( .IN1(n4732), .IN2(n7821), .QN(n7820) );
  NOR2X0 U9018 ( .IN1(n7482), .IN2(n4778), .QN(n7819) );
  XOR2X1 U9019 ( .IN1(n7822), .IN2(n7823), .Q(n7482) );
  XOR2X1 U9020 ( .IN1(n9559), .IN2(n4413), .Q(n7823) );
  XOR2X1 U9021 ( .IN1(WX5879), .IN2(n4263), .Q(n7822) );
  NOR2X0 U9022 ( .IN1(n7824), .IN2(n7825), .QN(n7817) );
  NOR2X0 U9023 ( .IN1(DFF_736_n1), .IN2(n4763), .QN(n7825) );
  NOR2X0 U9024 ( .IN1(n4803), .IN2(n6206), .QN(n7824) );
  NAND2X0 U9025 ( .IN1(n5309), .IN2(n8554), .QN(n6206) );
  NAND2X0 U9026 ( .IN1(n7826), .IN2(n7827), .QN(WX4583) );
  NOR2X0 U9027 ( .IN1(n7828), .IN2(n7829), .QN(n7827) );
  NOR2X0 U9028 ( .IN1(n7830), .IN2(n4729), .QN(n7829) );
  NOR2X0 U9029 ( .IN1(n4788), .IN2(n7491), .QN(n7828) );
  XNOR2X1 U9030 ( .IN1(n7831), .IN2(n7832), .Q(n7491) );
  XOR2X1 U9031 ( .IN1(test_so51), .IN2(n9560), .Q(n7832) );
  XOR2X1 U9032 ( .IN1(WX5877), .IN2(n4549), .Q(n7831) );
  NOR2X0 U9033 ( .IN1(n7833), .IN2(n7834), .QN(n7826) );
  NOR2X0 U9034 ( .IN1(DFF_737_n1), .IN2(n4764), .QN(n7834) );
  NOR2X0 U9035 ( .IN1(n4803), .IN2(n6207), .QN(n7833) );
  NAND2X0 U9036 ( .IN1(n5309), .IN2(n8555), .QN(n6207) );
  NAND2X0 U9037 ( .IN1(n7835), .IN2(n7836), .QN(WX4581) );
  NOR2X0 U9038 ( .IN1(n7837), .IN2(n7838), .QN(n7836) );
  NOR2X0 U9039 ( .IN1(n7839), .IN2(n4728), .QN(n7838) );
  NOR2X0 U9040 ( .IN1(n7500), .IN2(n4778), .QN(n7837) );
  XOR2X1 U9041 ( .IN1(n7840), .IN2(n7841), .Q(n7500) );
  XOR2X1 U9042 ( .IN1(n9561), .IN2(n4548), .Q(n7841) );
  XOR2X1 U9043 ( .IN1(WX5875), .IN2(n4266), .Q(n7840) );
  NOR2X0 U9044 ( .IN1(n7842), .IN2(n7843), .QN(n7835) );
  NOR2X0 U9045 ( .IN1(DFF_738_n1), .IN2(n4763), .QN(n7843) );
  NOR2X0 U9046 ( .IN1(n4803), .IN2(n6208), .QN(n7842) );
  NAND2X0 U9047 ( .IN1(test_so34), .IN2(n5323), .QN(n6208) );
  NAND2X0 U9048 ( .IN1(n7844), .IN2(n7845), .QN(WX4579) );
  NOR2X0 U9049 ( .IN1(n7846), .IN2(n7847), .QN(n7845) );
  NOR2X0 U9050 ( .IN1(n7848), .IN2(n4727), .QN(n7847) );
  NOR2X0 U9051 ( .IN1(n4788), .IN2(n7509), .QN(n7846) );
  XNOR2X1 U9052 ( .IN1(n7849), .IN2(n7850), .Q(n7509) );
  XOR2X1 U9053 ( .IN1(test_so49), .IN2(n9562), .Q(n7850) );
  XOR2X1 U9054 ( .IN1(WX5873), .IN2(n4547), .Q(n7849) );
  NOR2X0 U9055 ( .IN1(n7851), .IN2(n7852), .QN(n7844) );
  NOR2X0 U9056 ( .IN1(DFF_739_n1), .IN2(n4763), .QN(n7852) );
  NOR2X0 U9057 ( .IN1(n4803), .IN2(n6209), .QN(n7851) );
  NAND2X0 U9058 ( .IN1(n5309), .IN2(n8558), .QN(n6209) );
  NAND2X0 U9059 ( .IN1(n7853), .IN2(n7854), .QN(WX4577) );
  NOR2X0 U9060 ( .IN1(n7855), .IN2(n7856), .QN(n7854) );
  NOR2X0 U9061 ( .IN1(n7857), .IN2(n4728), .QN(n7856) );
  NOR2X0 U9062 ( .IN1(n7518), .IN2(n4779), .QN(n7855) );
  XOR2X1 U9063 ( .IN1(n7858), .IN2(n7859), .Q(n7518) );
  XOR2X1 U9064 ( .IN1(n9563), .IN2(n4400), .Q(n7859) );
  XOR2X1 U9065 ( .IN1(WX5871), .IN2(n4269), .Q(n7858) );
  NOR2X0 U9066 ( .IN1(n7860), .IN2(n7861), .QN(n7853) );
  NOR2X0 U9067 ( .IN1(DFF_740_n1), .IN2(n4763), .QN(n7861) );
  NOR2X0 U9068 ( .IN1(n4803), .IN2(n6210), .QN(n7860) );
  NAND2X0 U9069 ( .IN1(n5308), .IN2(n8559), .QN(n6210) );
  NAND2X0 U9070 ( .IN1(n7862), .IN2(n7863), .QN(WX4575) );
  NOR2X0 U9071 ( .IN1(n7864), .IN2(n7865), .QN(n7863) );
  NOR2X0 U9072 ( .IN1(n7866), .IN2(n4728), .QN(n7865) );
  NOR2X0 U9073 ( .IN1(n4788), .IN2(n7527), .QN(n7864) );
  XNOR2X1 U9074 ( .IN1(n7867), .IN2(n7868), .Q(n7527) );
  XOR2X1 U9075 ( .IN1(test_so47), .IN2(n9564), .Q(n7868) );
  XOR2X1 U9076 ( .IN1(WX5997), .IN2(n4546), .Q(n7867) );
  NOR2X0 U9077 ( .IN1(n7869), .IN2(n7870), .QN(n7862) );
  NOR2X0 U9078 ( .IN1(n4764), .IN2(n4700), .QN(n7870) );
  NOR2X0 U9079 ( .IN1(n4803), .IN2(n6211), .QN(n7869) );
  NAND2X0 U9080 ( .IN1(n5308), .IN2(n8560), .QN(n6211) );
  NAND2X0 U9081 ( .IN1(n7871), .IN2(n7872), .QN(WX4573) );
  NOR2X0 U9082 ( .IN1(n7873), .IN2(n7874), .QN(n7872) );
  NOR2X0 U9083 ( .IN1(n7875), .IN2(n4728), .QN(n7874) );
  NOR2X0 U9084 ( .IN1(n7536), .IN2(n4778), .QN(n7873) );
  XOR2X1 U9085 ( .IN1(n7876), .IN2(n7877), .Q(n7536) );
  XOR2X1 U9086 ( .IN1(n9565), .IN2(n4545), .Q(n7877) );
  XOR2X1 U9087 ( .IN1(WX5867), .IN2(n4272), .Q(n7876) );
  NOR2X0 U9088 ( .IN1(n7878), .IN2(n7879), .QN(n7871) );
  NOR2X0 U9089 ( .IN1(DFF_742_n1), .IN2(n4763), .QN(n7879) );
  NOR2X0 U9090 ( .IN1(n4803), .IN2(n6221), .QN(n7878) );
  NAND2X0 U9091 ( .IN1(n5308), .IN2(n8561), .QN(n6221) );
  NAND2X0 U9092 ( .IN1(n7880), .IN2(n7881), .QN(WX4571) );
  NOR2X0 U9093 ( .IN1(n7882), .IN2(n7883), .QN(n7881) );
  NOR2X0 U9094 ( .IN1(n7884), .IN2(n4728), .QN(n7883) );
  NOR2X0 U9095 ( .IN1(n7545), .IN2(n4778), .QN(n7882) );
  XOR2X1 U9096 ( .IN1(n7885), .IN2(n7886), .Q(n7545) );
  XOR2X1 U9097 ( .IN1(n9566), .IN2(n4544), .Q(n7886) );
  XOR2X1 U9098 ( .IN1(WX5865), .IN2(n4274), .Q(n7885) );
  NOR2X0 U9099 ( .IN1(n7887), .IN2(n7888), .QN(n7880) );
  NOR2X0 U9100 ( .IN1(DFF_743_n1), .IN2(n4762), .QN(n7888) );
  NOR2X0 U9101 ( .IN1(n4803), .IN2(n6222), .QN(n7887) );
  NAND2X0 U9102 ( .IN1(n5308), .IN2(n8562), .QN(n6222) );
  NAND2X0 U9103 ( .IN1(n7889), .IN2(n7890), .QN(WX4569) );
  NOR2X0 U9104 ( .IN1(n7891), .IN2(n7892), .QN(n7890) );
  NOR2X0 U9105 ( .IN1(n7893), .IN2(n4727), .QN(n7892) );
  NOR2X0 U9106 ( .IN1(n7554), .IN2(n4779), .QN(n7891) );
  XOR2X1 U9107 ( .IN1(n7894), .IN2(n7895), .Q(n7554) );
  XOR2X1 U9108 ( .IN1(n9567), .IN2(n4543), .Q(n7895) );
  XOR2X1 U9109 ( .IN1(WX5863), .IN2(n4276), .Q(n7894) );
  NOR2X0 U9110 ( .IN1(n7896), .IN2(n7897), .QN(n7889) );
  NOR2X0 U9111 ( .IN1(DFF_744_n1), .IN2(n4763), .QN(n7897) );
  NOR2X0 U9112 ( .IN1(n4803), .IN2(n6223), .QN(n7896) );
  NAND2X0 U9113 ( .IN1(n5308), .IN2(n8563), .QN(n6223) );
  NAND2X0 U9114 ( .IN1(n7898), .IN2(n7899), .QN(WX4567) );
  NOR2X0 U9115 ( .IN1(n7900), .IN2(n7901), .QN(n7899) );
  NOR2X0 U9116 ( .IN1(n7902), .IN2(n4727), .QN(n7901) );
  NOR2X0 U9117 ( .IN1(n7563), .IN2(n4779), .QN(n7900) );
  XOR2X1 U9118 ( .IN1(n7903), .IN2(n7904), .Q(n7563) );
  XOR2X1 U9119 ( .IN1(n9568), .IN2(n4542), .Q(n7904) );
  XOR2X1 U9120 ( .IN1(WX5861), .IN2(n4278), .Q(n7903) );
  NOR2X0 U9121 ( .IN1(n7905), .IN2(n7906), .QN(n7898) );
  NOR2X0 U9122 ( .IN1(DFF_745_n1), .IN2(n4762), .QN(n7906) );
  NOR2X0 U9123 ( .IN1(n4802), .IN2(n6224), .QN(n7905) );
  NAND2X0 U9124 ( .IN1(n5308), .IN2(n8564), .QN(n6224) );
  NAND2X0 U9125 ( .IN1(n7907), .IN2(n7908), .QN(WX4565) );
  NOR2X0 U9126 ( .IN1(n7909), .IN2(n7910), .QN(n7908) );
  NOR2X0 U9127 ( .IN1(n7911), .IN2(n4728), .QN(n7910) );
  NOR2X0 U9128 ( .IN1(n7572), .IN2(n4779), .QN(n7909) );
  XOR2X1 U9129 ( .IN1(n7912), .IN2(n7913), .Q(n7572) );
  XOR2X1 U9130 ( .IN1(n9569), .IN2(n4541), .Q(n7913) );
  XOR2X1 U9131 ( .IN1(WX5859), .IN2(n4280), .Q(n7912) );
  NOR2X0 U9132 ( .IN1(n7914), .IN2(n7915), .QN(n7907) );
  NOR2X0 U9133 ( .IN1(DFF_746_n1), .IN2(n4762), .QN(n7915) );
  NOR2X0 U9134 ( .IN1(n4802), .IN2(n6225), .QN(n7914) );
  NAND2X0 U9135 ( .IN1(n5307), .IN2(n8565), .QN(n6225) );
  NAND2X0 U9136 ( .IN1(n7916), .IN2(n7917), .QN(WX4563) );
  NOR2X0 U9137 ( .IN1(n7918), .IN2(n7919), .QN(n7917) );
  NOR2X0 U9138 ( .IN1(n4730), .IN2(n7920), .QN(n7919) );
  NOR2X0 U9139 ( .IN1(n7581), .IN2(n4779), .QN(n7918) );
  XOR2X1 U9140 ( .IN1(n7921), .IN2(n7922), .Q(n7581) );
  XOR2X1 U9141 ( .IN1(n9570), .IN2(n4399), .Q(n7922) );
  XOR2X1 U9142 ( .IN1(WX5857), .IN2(n4282), .Q(n7921) );
  NOR2X0 U9143 ( .IN1(n7923), .IN2(n7924), .QN(n7916) );
  NOR2X0 U9144 ( .IN1(DFF_747_n1), .IN2(n4762), .QN(n7924) );
  NOR2X0 U9145 ( .IN1(n4802), .IN2(n6226), .QN(n7923) );
  NAND2X0 U9146 ( .IN1(n5307), .IN2(n8566), .QN(n6226) );
  NAND2X0 U9147 ( .IN1(n7925), .IN2(n7926), .QN(WX4561) );
  NOR2X0 U9148 ( .IN1(n7927), .IN2(n7928), .QN(n7926) );
  NOR2X0 U9149 ( .IN1(n7929), .IN2(n4727), .QN(n7928) );
  NOR2X0 U9150 ( .IN1(n7590), .IN2(n4779), .QN(n7927) );
  XOR2X1 U9151 ( .IN1(n7930), .IN2(n7931), .Q(n7590) );
  XOR2X1 U9152 ( .IN1(n9571), .IN2(n4540), .Q(n7931) );
  XOR2X1 U9153 ( .IN1(WX5855), .IN2(n4284), .Q(n7930) );
  NOR2X0 U9154 ( .IN1(n7932), .IN2(n7933), .QN(n7925) );
  NOR2X0 U9155 ( .IN1(DFF_748_n1), .IN2(n4762), .QN(n7933) );
  NOR2X0 U9156 ( .IN1(n4802), .IN2(n6227), .QN(n7932) );
  NAND2X0 U9157 ( .IN1(n5307), .IN2(n8567), .QN(n6227) );
  NAND2X0 U9158 ( .IN1(n7934), .IN2(n7935), .QN(WX4559) );
  NOR2X0 U9159 ( .IN1(n7936), .IN2(n7937), .QN(n7935) );
  NOR2X0 U9160 ( .IN1(n4730), .IN2(n7938), .QN(n7937) );
  NOR2X0 U9161 ( .IN1(n7599), .IN2(n4779), .QN(n7936) );
  XOR2X1 U9162 ( .IN1(n7939), .IN2(n7940), .Q(n7599) );
  XOR2X1 U9163 ( .IN1(n9572), .IN2(n4539), .Q(n7940) );
  XOR2X1 U9164 ( .IN1(WX5853), .IN2(n4286), .Q(n7939) );
  NOR2X0 U9165 ( .IN1(n7941), .IN2(n7942), .QN(n7934) );
  NOR2X0 U9166 ( .IN1(DFF_749_n1), .IN2(n4762), .QN(n7942) );
  NOR2X0 U9167 ( .IN1(n4802), .IN2(n6228), .QN(n7941) );
  NAND2X0 U9168 ( .IN1(n5307), .IN2(n8568), .QN(n6228) );
  NAND2X0 U9169 ( .IN1(n7943), .IN2(n7944), .QN(WX4557) );
  NOR2X0 U9170 ( .IN1(n7945), .IN2(n7946), .QN(n7944) );
  NOR2X0 U9171 ( .IN1(n7947), .IN2(n4728), .QN(n7946) );
  NOR2X0 U9172 ( .IN1(n7608), .IN2(n4779), .QN(n7945) );
  XOR2X1 U9173 ( .IN1(n7948), .IN2(n7949), .Q(n7608) );
  XOR2X1 U9174 ( .IN1(n9573), .IN2(n4538), .Q(n7949) );
  XOR2X1 U9175 ( .IN1(WX5851), .IN2(n4288), .Q(n7948) );
  NOR2X0 U9176 ( .IN1(n7950), .IN2(n7951), .QN(n7943) );
  NOR2X0 U9177 ( .IN1(DFF_750_n1), .IN2(n4762), .QN(n7951) );
  NOR2X0 U9178 ( .IN1(n4802), .IN2(n6229), .QN(n7950) );
  NAND2X0 U9179 ( .IN1(n5307), .IN2(n8569), .QN(n6229) );
  NAND2X0 U9180 ( .IN1(n7952), .IN2(n7953), .QN(WX4555) );
  NOR2X0 U9181 ( .IN1(n7954), .IN2(n7955), .QN(n7953) );
  NOR2X0 U9182 ( .IN1(n4730), .IN2(n7956), .QN(n7955) );
  NOR2X0 U9183 ( .IN1(n7617), .IN2(n4780), .QN(n7954) );
  XOR2X1 U9184 ( .IN1(n7957), .IN2(n7958), .Q(n7617) );
  XOR2X1 U9185 ( .IN1(n9574), .IN2(n4537), .Q(n7958) );
  XOR2X1 U9186 ( .IN1(WX5849), .IN2(n4290), .Q(n7957) );
  NOR2X0 U9187 ( .IN1(n7959), .IN2(n7960), .QN(n7952) );
  NOR2X0 U9188 ( .IN1(DFF_751_n1), .IN2(n4762), .QN(n7960) );
  NOR2X0 U9189 ( .IN1(n4802), .IN2(n6230), .QN(n7959) );
  NAND2X0 U9190 ( .IN1(n5307), .IN2(n8570), .QN(n6230) );
  NAND2X0 U9191 ( .IN1(n7961), .IN2(n7962), .QN(WX4553) );
  NOR2X0 U9192 ( .IN1(n7963), .IN2(n7964), .QN(n7962) );
  NOR2X0 U9193 ( .IN1(n7965), .IN2(n4726), .QN(n7964) );
  NOR2X0 U9194 ( .IN1(n4788), .IN2(n7626), .QN(n7963) );
  XNOR2X1 U9195 ( .IN1(n7966), .IN2(n7967), .Q(n7626) );
  XOR2X1 U9196 ( .IN1(n4091), .IN2(n5252), .Q(n7967) );
  XOR2X1 U9197 ( .IN1(WX5911), .IN2(n7968), .Q(n7966) );
  XOR2X1 U9198 ( .IN1(test_so52), .IN2(n9575), .Q(n7968) );
  NOR2X0 U9199 ( .IN1(n7969), .IN2(n7970), .QN(n7961) );
  NOR2X0 U9200 ( .IN1(DFF_752_n1), .IN2(n4762), .QN(n7970) );
  NOR2X0 U9201 ( .IN1(n4802), .IN2(n6249), .QN(n7969) );
  NAND2X0 U9202 ( .IN1(n5306), .IN2(n8571), .QN(n6249) );
  NAND2X0 U9203 ( .IN1(n7971), .IN2(n7972), .QN(WX4551) );
  NOR2X0 U9204 ( .IN1(n7973), .IN2(n7974), .QN(n7972) );
  NOR2X0 U9205 ( .IN1(n4731), .IN2(n7975), .QN(n7974) );
  NOR2X0 U9206 ( .IN1(n7636), .IN2(n4779), .QN(n7973) );
  XOR2X1 U9207 ( .IN1(n7976), .IN2(n7977), .Q(n7636) );
  XOR2X1 U9208 ( .IN1(n4092), .IN2(n5252), .Q(n7977) );
  XOR2X1 U9209 ( .IN1(n7978), .IN2(n4536), .Q(n7976) );
  XOR2X1 U9210 ( .IN1(WX5973), .IN2(n9576), .Q(n7978) );
  NOR2X0 U9211 ( .IN1(n7979), .IN2(n7980), .QN(n7971) );
  NOR2X0 U9212 ( .IN1(DFF_753_n1), .IN2(n4762), .QN(n7980) );
  NOR2X0 U9213 ( .IN1(n4802), .IN2(n6250), .QN(n7979) );
  NAND2X0 U9214 ( .IN1(n5306), .IN2(n8572), .QN(n6250) );
  NAND2X0 U9215 ( .IN1(n7981), .IN2(n7982), .QN(WX4549) );
  NOR2X0 U9216 ( .IN1(n7983), .IN2(n7984), .QN(n7982) );
  NOR2X0 U9217 ( .IN1(n7985), .IN2(n4728), .QN(n7984) );
  NOR2X0 U9218 ( .IN1(n4787), .IN2(n7646), .QN(n7983) );
  XNOR2X1 U9219 ( .IN1(n7986), .IN2(n7987), .Q(n7646) );
  XOR2X1 U9220 ( .IN1(n4535), .IN2(n5252), .Q(n7987) );
  XOR2X1 U9221 ( .IN1(n7988), .IN2(n9579), .Q(n7986) );
  XOR2X1 U9222 ( .IN1(n9578), .IN2(n9577), .Q(n7988) );
  NOR2X0 U9223 ( .IN1(n7989), .IN2(n7990), .QN(n7981) );
  NOR2X0 U9224 ( .IN1(DFF_754_n1), .IN2(n4761), .QN(n7990) );
  NOR2X0 U9225 ( .IN1(n4802), .IN2(n6251), .QN(n7989) );
  NAND2X0 U9226 ( .IN1(n5306), .IN2(n8573), .QN(n6251) );
  NAND2X0 U9227 ( .IN1(n7991), .IN2(n7992), .QN(WX4547) );
  NOR2X0 U9228 ( .IN1(n7993), .IN2(n7994), .QN(n7992) );
  NOR2X0 U9229 ( .IN1(n7995), .IN2(n4727), .QN(n7994) );
  NOR2X0 U9230 ( .IN1(n7656), .IN2(n4779), .QN(n7993) );
  XOR2X1 U9231 ( .IN1(n7996), .IN2(n7997), .Q(n7656) );
  XOR2X1 U9232 ( .IN1(n4093), .IN2(n5252), .Q(n7997) );
  XOR2X1 U9233 ( .IN1(n7998), .IN2(n4534), .Q(n7996) );
  XOR2X1 U9234 ( .IN1(WX5969), .IN2(n9580), .Q(n7998) );
  NOR2X0 U9235 ( .IN1(n7999), .IN2(n8000), .QN(n7991) );
  NOR2X0 U9236 ( .IN1(DFF_755_n1), .IN2(n4761), .QN(n8000) );
  NOR2X0 U9237 ( .IN1(n4802), .IN2(n6252), .QN(n7999) );
  NAND2X0 U9238 ( .IN1(test_so33), .IN2(n5322), .QN(n6252) );
  NAND2X0 U9239 ( .IN1(n8001), .IN2(n8002), .QN(WX4545) );
  NOR2X0 U9240 ( .IN1(n8003), .IN2(n8004), .QN(n8002) );
  NOR2X0 U9241 ( .IN1(n8005), .IN2(n4728), .QN(n8004) );
  NOR2X0 U9242 ( .IN1(n4787), .IN2(n7666), .QN(n8003) );
  XNOR2X1 U9243 ( .IN1(n8006), .IN2(n8007), .Q(n7666) );
  XOR2X1 U9244 ( .IN1(n4533), .IN2(n5252), .Q(n8007) );
  XOR2X1 U9245 ( .IN1(n8008), .IN2(n9583), .Q(n8006) );
  XOR2X1 U9246 ( .IN1(n9582), .IN2(n9581), .Q(n8008) );
  NOR2X0 U9247 ( .IN1(n8009), .IN2(n8010), .QN(n8001) );
  NOR2X0 U9248 ( .IN1(DFF_756_n1), .IN2(n4762), .QN(n8010) );
  NOR2X0 U9249 ( .IN1(n4802), .IN2(n6253), .QN(n8009) );
  NAND2X0 U9250 ( .IN1(n5306), .IN2(n8576), .QN(n6253) );
  NAND2X0 U9251 ( .IN1(n8011), .IN2(n8012), .QN(WX4543) );
  NOR2X0 U9252 ( .IN1(n8013), .IN2(n8014), .QN(n8012) );
  NOR2X0 U9253 ( .IN1(n8015), .IN2(n4728), .QN(n8014) );
  NOR2X0 U9254 ( .IN1(n7676), .IN2(n4780), .QN(n8013) );
  XOR2X1 U9255 ( .IN1(n8016), .IN2(n8017), .Q(n7676) );
  XOR2X1 U9256 ( .IN1(n4094), .IN2(n5252), .Q(n8017) );
  XOR2X1 U9257 ( .IN1(n8018), .IN2(n4532), .Q(n8016) );
  XOR2X1 U9258 ( .IN1(WX5965), .IN2(n9584), .Q(n8018) );
  NOR2X0 U9259 ( .IN1(n8019), .IN2(n8020), .QN(n8011) );
  NOR2X0 U9260 ( .IN1(DFF_757_n1), .IN2(n4761), .QN(n8020) );
  NOR2X0 U9261 ( .IN1(n4802), .IN2(n6254), .QN(n8019) );
  NAND2X0 U9262 ( .IN1(n5306), .IN2(n8577), .QN(n6254) );
  NAND2X0 U9263 ( .IN1(n8021), .IN2(n8022), .QN(WX4541) );
  NOR2X0 U9264 ( .IN1(n8023), .IN2(n8024), .QN(n8022) );
  NOR2X0 U9265 ( .IN1(n8025), .IN2(n4727), .QN(n8024) );
  NOR2X0 U9266 ( .IN1(n4787), .IN2(n7686), .QN(n8023) );
  XNOR2X1 U9267 ( .IN1(n8026), .IN2(n8027), .Q(n7686) );
  XOR2X1 U9268 ( .IN1(n4095), .IN2(n5252), .Q(n8027) );
  XOR2X1 U9269 ( .IN1(n8028), .IN2(n4531), .Q(n8026) );
  XOR2X1 U9270 ( .IN1(WX5899), .IN2(test_so46), .Q(n8028) );
  NOR2X0 U9271 ( .IN1(n8029), .IN2(n8030), .QN(n8021) );
  NOR2X0 U9272 ( .IN1(n4764), .IN2(n4701), .QN(n8030) );
  NOR2X0 U9273 ( .IN1(n4801), .IN2(n6255), .QN(n8029) );
  NAND2X0 U9274 ( .IN1(n5306), .IN2(n8578), .QN(n6255) );
  NAND2X0 U9275 ( .IN1(n8031), .IN2(n8032), .QN(WX4539) );
  NOR2X0 U9276 ( .IN1(n8033), .IN2(n8034), .QN(n8032) );
  NOR2X0 U9277 ( .IN1(n8035), .IN2(n4727), .QN(n8034) );
  NOR2X0 U9278 ( .IN1(n7696), .IN2(n4780), .QN(n8033) );
  XOR2X1 U9279 ( .IN1(n8036), .IN2(n8037), .Q(n7696) );
  XOR2X1 U9280 ( .IN1(n4096), .IN2(n5252), .Q(n8037) );
  XOR2X1 U9281 ( .IN1(n8038), .IN2(n4530), .Q(n8036) );
  XOR2X1 U9282 ( .IN1(WX5961), .IN2(n9585), .Q(n8038) );
  NOR2X0 U9283 ( .IN1(n8039), .IN2(n8040), .QN(n8031) );
  NOR2X0 U9284 ( .IN1(DFF_759_n1), .IN2(n4761), .QN(n8040) );
  NOR2X0 U9285 ( .IN1(n4801), .IN2(n6256), .QN(n8039) );
  NAND2X0 U9286 ( .IN1(n5305), .IN2(n8579), .QN(n6256) );
  NAND2X0 U9287 ( .IN1(n8041), .IN2(n8042), .QN(WX4537) );
  NOR2X0 U9288 ( .IN1(n8043), .IN2(n8044), .QN(n8042) );
  NOR2X0 U9289 ( .IN1(n8045), .IN2(n4727), .QN(n8044) );
  NOR2X0 U9290 ( .IN1(n7706), .IN2(n4781), .QN(n8043) );
  XOR2X1 U9291 ( .IN1(n8046), .IN2(n8047), .Q(n7706) );
  XOR2X1 U9292 ( .IN1(n4097), .IN2(n5253), .Q(n8047) );
  XOR2X1 U9293 ( .IN1(n8048), .IN2(n4529), .Q(n8046) );
  XOR2X1 U9294 ( .IN1(WX5959), .IN2(n9586), .Q(n8048) );
  NOR2X0 U9295 ( .IN1(n8049), .IN2(n8050), .QN(n8041) );
  NOR2X0 U9296 ( .IN1(DFF_760_n1), .IN2(n4761), .QN(n8050) );
  NOR2X0 U9297 ( .IN1(n4801), .IN2(n6257), .QN(n8049) );
  NAND2X0 U9298 ( .IN1(n5305), .IN2(n8580), .QN(n6257) );
  NAND2X0 U9299 ( .IN1(n8051), .IN2(n8052), .QN(WX4535) );
  NOR2X0 U9300 ( .IN1(n8053), .IN2(n8054), .QN(n8052) );
  NOR2X0 U9301 ( .IN1(n8055), .IN2(n4727), .QN(n8054) );
  NOR2X0 U9302 ( .IN1(n7716), .IN2(n4781), .QN(n8053) );
  XOR2X1 U9303 ( .IN1(n8056), .IN2(n8057), .Q(n7716) );
  XOR2X1 U9304 ( .IN1(n4098), .IN2(n5253), .Q(n8057) );
  XOR2X1 U9305 ( .IN1(n8058), .IN2(n4528), .Q(n8056) );
  XOR2X1 U9306 ( .IN1(WX5957), .IN2(n9587), .Q(n8058) );
  NOR2X0 U9307 ( .IN1(n8059), .IN2(n8060), .QN(n8051) );
  NOR2X0 U9308 ( .IN1(DFF_761_n1), .IN2(n4761), .QN(n8060) );
  NOR2X0 U9309 ( .IN1(n4801), .IN2(n6258), .QN(n8059) );
  NAND2X0 U9310 ( .IN1(n5305), .IN2(n8581), .QN(n6258) );
  NAND2X0 U9311 ( .IN1(n8061), .IN2(n8062), .QN(WX4533) );
  NOR2X0 U9312 ( .IN1(n8063), .IN2(n8064), .QN(n8062) );
  NOR2X0 U9313 ( .IN1(n8065), .IN2(n4727), .QN(n8064) );
  NOR2X0 U9314 ( .IN1(n7726), .IN2(n4780), .QN(n8063) );
  XOR2X1 U9315 ( .IN1(n8066), .IN2(n8067), .Q(n7726) );
  XOR2X1 U9316 ( .IN1(n4099), .IN2(n5253), .Q(n8067) );
  XOR2X1 U9317 ( .IN1(n8068), .IN2(n4527), .Q(n8066) );
  XOR2X1 U9318 ( .IN1(WX5955), .IN2(n9588), .Q(n8068) );
  NOR2X0 U9319 ( .IN1(n8069), .IN2(n8070), .QN(n8061) );
  NOR2X0 U9320 ( .IN1(DFF_762_n1), .IN2(n4761), .QN(n8070) );
  NOR2X0 U9321 ( .IN1(n4801), .IN2(n6268), .QN(n8069) );
  NAND2X0 U9322 ( .IN1(n5305), .IN2(n8582), .QN(n6268) );
  NAND2X0 U9323 ( .IN1(n8071), .IN2(n8072), .QN(WX4531) );
  NOR2X0 U9324 ( .IN1(n8073), .IN2(n8074), .QN(n8072) );
  NOR2X0 U9325 ( .IN1(n8075), .IN2(n4727), .QN(n8074) );
  NOR2X0 U9326 ( .IN1(n7736), .IN2(n4781), .QN(n8073) );
  XOR2X1 U9327 ( .IN1(n8076), .IN2(n8077), .Q(n7736) );
  XOR2X1 U9328 ( .IN1(n4100), .IN2(n5253), .Q(n8077) );
  XOR2X1 U9329 ( .IN1(n8078), .IN2(n4526), .Q(n8076) );
  XOR2X1 U9330 ( .IN1(WX5953), .IN2(n9589), .Q(n8078) );
  NOR2X0 U9331 ( .IN1(n8079), .IN2(n8080), .QN(n8071) );
  NOR2X0 U9332 ( .IN1(DFF_763_n1), .IN2(n4761), .QN(n8080) );
  NOR2X0 U9333 ( .IN1(n4801), .IN2(n6269), .QN(n8079) );
  NAND2X0 U9334 ( .IN1(n5305), .IN2(n8583), .QN(n6269) );
  NAND2X0 U9335 ( .IN1(n8081), .IN2(n8082), .QN(WX4529) );
  NOR2X0 U9336 ( .IN1(n8083), .IN2(n8084), .QN(n8082) );
  NOR2X0 U9337 ( .IN1(n4731), .IN2(n8085), .QN(n8084) );
  NOR2X0 U9338 ( .IN1(n7746), .IN2(n4781), .QN(n8083) );
  XOR2X1 U9339 ( .IN1(n8086), .IN2(n8087), .Q(n7746) );
  XOR2X1 U9340 ( .IN1(n4101), .IN2(n5253), .Q(n8087) );
  XOR2X1 U9341 ( .IN1(n8088), .IN2(n4525), .Q(n8086) );
  XOR2X1 U9342 ( .IN1(WX5951), .IN2(n9590), .Q(n8088) );
  NOR2X0 U9343 ( .IN1(n8089), .IN2(n8090), .QN(n8081) );
  NOR2X0 U9344 ( .IN1(DFF_764_n1), .IN2(n4761), .QN(n8090) );
  NOR2X0 U9345 ( .IN1(n4801), .IN2(n6270), .QN(n8089) );
  NAND2X0 U9346 ( .IN1(n5305), .IN2(n8584), .QN(n6270) );
  NAND2X0 U9347 ( .IN1(n8091), .IN2(n8092), .QN(WX4527) );
  NOR2X0 U9348 ( .IN1(n8093), .IN2(n8094), .QN(n8092) );
  NOR2X0 U9349 ( .IN1(n8095), .IN2(n4726), .QN(n8094) );
  NOR2X0 U9350 ( .IN1(n7756), .IN2(n4781), .QN(n8093) );
  XOR2X1 U9351 ( .IN1(n8096), .IN2(n8097), .Q(n7756) );
  XOR2X1 U9352 ( .IN1(n4102), .IN2(n5253), .Q(n8097) );
  XOR2X1 U9353 ( .IN1(n8098), .IN2(n4524), .Q(n8096) );
  XOR2X1 U9354 ( .IN1(WX5949), .IN2(n9591), .Q(n8098) );
  NOR2X0 U9355 ( .IN1(n8099), .IN2(n8100), .QN(n8091) );
  NOR2X0 U9356 ( .IN1(DFF_765_n1), .IN2(n4761), .QN(n8100) );
  NOR2X0 U9357 ( .IN1(n4801), .IN2(n6271), .QN(n8099) );
  NAND2X0 U9358 ( .IN1(n5304), .IN2(n8585), .QN(n6271) );
  NAND2X0 U9359 ( .IN1(n8101), .IN2(n8102), .QN(WX4525) );
  NOR2X0 U9360 ( .IN1(n8103), .IN2(n8104), .QN(n8102) );
  NOR2X0 U9361 ( .IN1(n4729), .IN2(n8105), .QN(n8104) );
  NOR2X0 U9362 ( .IN1(n7766), .IN2(n4781), .QN(n8103) );
  XOR2X1 U9363 ( .IN1(n8106), .IN2(n8107), .Q(n7766) );
  XOR2X1 U9364 ( .IN1(n4103), .IN2(n5253), .Q(n8107) );
  XOR2X1 U9365 ( .IN1(n8108), .IN2(n4523), .Q(n8106) );
  XOR2X1 U9366 ( .IN1(WX5947), .IN2(n9592), .Q(n8108) );
  NOR2X0 U9367 ( .IN1(n8109), .IN2(n8110), .QN(n8101) );
  NOR2X0 U9368 ( .IN1(DFF_766_n1), .IN2(n4761), .QN(n8110) );
  NOR2X0 U9369 ( .IN1(n4801), .IN2(n6272), .QN(n8109) );
  NAND2X0 U9370 ( .IN1(n5304), .IN2(n8586), .QN(n6272) );
  NAND2X0 U9371 ( .IN1(n8111), .IN2(n8112), .QN(WX4523) );
  NOR2X0 U9372 ( .IN1(n8113), .IN2(n8114), .QN(n8112) );
  NOR2X0 U9373 ( .IN1(n8115), .IN2(n4726), .QN(n8114) );
  NOR2X0 U9374 ( .IN1(n7776), .IN2(n4781), .QN(n8113) );
  XOR2X1 U9375 ( .IN1(n8116), .IN2(n8117), .Q(n7776) );
  XOR2X1 U9376 ( .IN1(n4035), .IN2(n5253), .Q(n8117) );
  XOR2X1 U9377 ( .IN1(n8118), .IN2(n4522), .Q(n8116) );
  XOR2X1 U9378 ( .IN1(WX5945), .IN2(n9593), .Q(n8118) );
  NOR2X0 U9379 ( .IN1(n8119), .IN2(n8120), .QN(n8111) );
  NOR2X0 U9380 ( .IN1(n4385), .IN2(n6717), .QN(n8120) );
  NOR2X0 U9381 ( .IN1(DFF_767_n1), .IN2(n4761), .QN(n8119) );
  NOR2X0 U9382 ( .IN1(n5439), .IN2(WX4364), .QN(WX4425) );
  NOR2X0 U9383 ( .IN1(n5439), .IN2(n8121), .QN(WX3912) );
  XOR2X1 U9384 ( .IN1(n4577), .IN2(DFF_574_n1), .Q(n8121) );
  NOR2X0 U9385 ( .IN1(n5439), .IN2(n8122), .QN(WX3910) );
  XOR2X1 U9386 ( .IN1(n4578), .IN2(DFF_573_n1), .Q(n8122) );
  NOR2X0 U9387 ( .IN1(n5440), .IN2(n8123), .QN(WX3908) );
  XOR2X1 U9388 ( .IN1(n4579), .IN2(DFF_572_n1), .Q(n8123) );
  NOR2X0 U9389 ( .IN1(n5440), .IN2(n8124), .QN(WX3906) );
  XOR2X1 U9390 ( .IN1(n4580), .IN2(n4702), .Q(n8124) );
  NOR2X0 U9391 ( .IN1(n5440), .IN2(n8125), .QN(WX3904) );
  XOR2X1 U9392 ( .IN1(n4581), .IN2(DFF_570_n1), .Q(n8125) );
  NOR2X0 U9393 ( .IN1(n5440), .IN2(n8126), .QN(WX3902) );
  XOR2X1 U9394 ( .IN1(n4582), .IN2(DFF_569_n1), .Q(n8126) );
  NOR2X0 U9395 ( .IN1(n5440), .IN2(n8127), .QN(WX3900) );
  XOR2X1 U9396 ( .IN1(n4583), .IN2(DFF_568_n1), .Q(n8127) );
  NOR2X0 U9397 ( .IN1(n5440), .IN2(n8128), .QN(WX3898) );
  XOR2X1 U9398 ( .IN1(n4584), .IN2(DFF_567_n1), .Q(n8128) );
  NOR2X0 U9399 ( .IN1(n5440), .IN2(n8129), .QN(WX3896) );
  XNOR2X1 U9400 ( .IN1(DFF_566_n1), .IN2(test_so29), .Q(n8129) );
  NOR2X0 U9401 ( .IN1(n5440), .IN2(n8130), .QN(WX3894) );
  XOR2X1 U9402 ( .IN1(n4585), .IN2(DFF_565_n1), .Q(n8130) );
  NOR2X0 U9403 ( .IN1(n5440), .IN2(n8131), .QN(WX3892) );
  XOR2X1 U9404 ( .IN1(n4586), .IN2(DFF_564_n1), .Q(n8131) );
  NOR2X0 U9405 ( .IN1(n5440), .IN2(n8132), .QN(WX3890) );
  XOR2X1 U9406 ( .IN1(n4587), .IN2(DFF_563_n1), .Q(n8132) );
  NOR2X0 U9407 ( .IN1(n5440), .IN2(n8133), .QN(WX3888) );
  XOR2X1 U9408 ( .IN1(n4588), .IN2(DFF_562_n1), .Q(n8133) );
  NOR2X0 U9409 ( .IN1(n5440), .IN2(n8134), .QN(WX3886) );
  XOR2X1 U9410 ( .IN1(n4589), .IN2(DFF_561_n1), .Q(n8134) );
  NOR2X0 U9411 ( .IN1(n5440), .IN2(n8135), .QN(WX3884) );
  XOR2X1 U9412 ( .IN1(n4590), .IN2(DFF_560_n1), .Q(n8135) );
  NOR2X0 U9413 ( .IN1(n5441), .IN2(n8136), .QN(WX3882) );
  XNOR2X1 U9414 ( .IN1(DFF_559_n1), .IN2(n8137), .Q(n8136) );
  XOR2X1 U9415 ( .IN1(n4403), .IN2(DFF_575_n1), .Q(n8137) );
  NOR2X0 U9416 ( .IN1(n5441), .IN2(n8138), .QN(WX3880) );
  XOR2X1 U9417 ( .IN1(n4591), .IN2(DFF_558_n1), .Q(n8138) );
  NOR2X0 U9418 ( .IN1(n5441), .IN2(n8139), .QN(WX3878) );
  XOR2X1 U9419 ( .IN1(n4592), .IN2(DFF_557_n1), .Q(n8139) );
  NOR2X0 U9420 ( .IN1(n5441), .IN2(n8140), .QN(WX3876) );
  XOR2X1 U9421 ( .IN1(n4593), .IN2(DFF_556_n1), .Q(n8140) );
  NOR2X0 U9422 ( .IN1(n5441), .IN2(n8141), .QN(WX3874) );
  XOR2X1 U9423 ( .IN1(n4594), .IN2(DFF_555_n1), .Q(n8141) );
  NOR2X0 U9424 ( .IN1(n5441), .IN2(n8142), .QN(WX3872) );
  XOR2X1 U9425 ( .IN1(DFF_575_n1), .IN2(n8143), .Q(n8142) );
  XOR2X1 U9426 ( .IN1(test_so31), .IN2(n4404), .Q(n8143) );
  NOR2X0 U9427 ( .IN1(n5441), .IN2(n8144), .QN(WX3870) );
  XOR2X1 U9428 ( .IN1(n4595), .IN2(DFF_553_n1), .Q(n8144) );
  NOR2X0 U9429 ( .IN1(n5441), .IN2(n8145), .QN(WX3868) );
  XOR2X1 U9430 ( .IN1(n4596), .IN2(DFF_552_n1), .Q(n8145) );
  NOR2X0 U9431 ( .IN1(n5441), .IN2(n8146), .QN(WX3866) );
  XOR2X1 U9432 ( .IN1(n4597), .IN2(DFF_551_n1), .Q(n8146) );
  NOR2X0 U9433 ( .IN1(n5441), .IN2(n8147), .QN(WX3864) );
  XOR2X1 U9434 ( .IN1(n4598), .IN2(DFF_550_n1), .Q(n8147) );
  NOR2X0 U9435 ( .IN1(n5441), .IN2(n8148), .QN(WX3862) );
  XNOR2X1 U9436 ( .IN1(DFF_549_n1), .IN2(test_so30), .Q(n8148) );
  NOR2X0 U9437 ( .IN1(n5441), .IN2(n8149), .QN(WX3860) );
  XOR2X1 U9438 ( .IN1(n4599), .IN2(DFF_548_n1), .Q(n8149) );
  NOR2X0 U9439 ( .IN1(n5441), .IN2(n8150), .QN(WX3858) );
  XNOR2X1 U9440 ( .IN1(DFF_547_n1), .IN2(n8151), .Q(n8150) );
  XOR2X1 U9441 ( .IN1(n4405), .IN2(DFF_575_n1), .Q(n8151) );
  NOR2X0 U9442 ( .IN1(n5405), .IN2(n8152), .QN(WX3856) );
  XOR2X1 U9443 ( .IN1(n4600), .IN2(DFF_546_n1), .Q(n8152) );
  NOR2X0 U9444 ( .IN1(n5406), .IN2(n8153), .QN(WX3854) );
  XOR2X1 U9445 ( .IN1(n4601), .IN2(DFF_545_n1), .Q(n8153) );
  NOR2X0 U9446 ( .IN1(n5407), .IN2(n8154), .QN(WX3852) );
  XOR2X1 U9447 ( .IN1(n4602), .IN2(DFF_544_n1), .Q(n8154) );
  NOR2X0 U9448 ( .IN1(n5408), .IN2(n8155), .QN(WX3850) );
  XOR2X1 U9449 ( .IN1(n4415), .IN2(DFF_575_n1), .Q(n8155) );
  NOR2X0 U9450 ( .IN1(n5409), .IN2(n4710), .QN(WX3324) );
  NOR2X0 U9451 ( .IN1(n9661), .IN2(n5351), .QN(WX3322) );
  NOR2X0 U9452 ( .IN1(n9665), .IN2(n5351), .QN(WX3320) );
  NOR2X0 U9453 ( .IN1(n9667), .IN2(n5351), .QN(WX3318) );
  NOR2X0 U9454 ( .IN1(n9669), .IN2(n5351), .QN(WX3316) );
  NOR2X0 U9455 ( .IN1(n9671), .IN2(n5351), .QN(WX3314) );
  NOR2X0 U9456 ( .IN1(n9672), .IN2(n5351), .QN(WX3312) );
  NOR2X0 U9457 ( .IN1(n9674), .IN2(n5351), .QN(WX3310) );
  NOR2X0 U9458 ( .IN1(n9676), .IN2(n5351), .QN(WX3308) );
  NOR2X0 U9459 ( .IN1(n9678), .IN2(n5351), .QN(WX3306) );
  NOR2X0 U9460 ( .IN1(n9680), .IN2(n5351), .QN(WX3304) );
  NOR2X0 U9461 ( .IN1(n9684), .IN2(n5351), .QN(WX3302) );
  NOR2X0 U9462 ( .IN1(n9686), .IN2(n5350), .QN(WX3300) );
  NOR2X0 U9463 ( .IN1(n9688), .IN2(n5350), .QN(WX3298) );
  NOR2X0 U9464 ( .IN1(n9690), .IN2(n5350), .QN(WX3296) );
  NOR2X0 U9465 ( .IN1(n9693), .IN2(n5350), .QN(WX3294) );
  NAND2X0 U9466 ( .IN1(n8156), .IN2(n8157), .QN(WX3292) );
  NOR2X0 U9467 ( .IN1(n8158), .IN2(n8159), .QN(n8157) );
  NOR2X0 U9468 ( .IN1(n8160), .IN2(n4726), .QN(n8159) );
  NOR2X0 U9469 ( .IN1(n4787), .IN2(n7821), .QN(n8158) );
  XNOR2X1 U9470 ( .IN1(n8161), .IN2(n8162), .Q(n7821) );
  XOR2X1 U9471 ( .IN1(test_so36), .IN2(n9594), .Q(n8162) );
  XOR2X1 U9472 ( .IN1(WX4714), .IN2(n4414), .Q(n8161) );
  NOR2X0 U9473 ( .IN1(n8163), .IN2(n8164), .QN(n8156) );
  NOR2X0 U9474 ( .IN1(DFF_544_n1), .IN2(n4760), .QN(n8164) );
  NOR2X0 U9475 ( .IN1(n4801), .IN2(n6291), .QN(n8163) );
  NAND2X0 U9476 ( .IN1(n5304), .IN2(n8612), .QN(n6291) );
  NAND2X0 U9477 ( .IN1(n8165), .IN2(n8166), .QN(WX3290) );
  NOR2X0 U9478 ( .IN1(n8167), .IN2(n8168), .QN(n8166) );
  NOR2X0 U9479 ( .IN1(n8169), .IN2(n4726), .QN(n8168) );
  NOR2X0 U9480 ( .IN1(n7830), .IN2(n4781), .QN(n8167) );
  XOR2X1 U9481 ( .IN1(n8170), .IN2(n8171), .Q(n7830) );
  XOR2X1 U9482 ( .IN1(n9595), .IN2(n4576), .Q(n8171) );
  XOR2X1 U9483 ( .IN1(WX4584), .IN2(n4293), .Q(n8170) );
  NOR2X0 U9484 ( .IN1(n8172), .IN2(n8173), .QN(n8165) );
  NOR2X0 U9485 ( .IN1(DFF_545_n1), .IN2(n4760), .QN(n8173) );
  NOR2X0 U9486 ( .IN1(n4801), .IN2(n6292), .QN(n8172) );
  NAND2X0 U9487 ( .IN1(n5304), .IN2(n8613), .QN(n6292) );
  NAND2X0 U9488 ( .IN1(n8174), .IN2(n8175), .QN(WX3288) );
  NOR2X0 U9489 ( .IN1(n8176), .IN2(n8177), .QN(n8175) );
  NOR2X0 U9490 ( .IN1(n8178), .IN2(n4726), .QN(n8177) );
  NOR2X0 U9491 ( .IN1(n7839), .IN2(n4782), .QN(n8176) );
  XOR2X1 U9492 ( .IN1(n8179), .IN2(n8180), .Q(n7839) );
  XOR2X1 U9493 ( .IN1(n9596), .IN2(n4575), .Q(n8180) );
  XOR2X1 U9494 ( .IN1(WX4582), .IN2(n4295), .Q(n8179) );
  NOR2X0 U9495 ( .IN1(n8181), .IN2(n8182), .QN(n8174) );
  NOR2X0 U9496 ( .IN1(DFF_546_n1), .IN2(n4760), .QN(n8182) );
  NOR2X0 U9497 ( .IN1(n4801), .IN2(n6293), .QN(n8181) );
  NAND2X0 U9498 ( .IN1(test_so23), .IN2(n5324), .QN(n6293) );
  NAND2X0 U9499 ( .IN1(n8183), .IN2(n8184), .QN(WX3286) );
  NOR2X0 U9500 ( .IN1(n8185), .IN2(n8186), .QN(n8184) );
  NOR2X0 U9501 ( .IN1(n8187), .IN2(n4726), .QN(n8186) );
  NOR2X0 U9502 ( .IN1(n7848), .IN2(n4781), .QN(n8185) );
  XOR2X1 U9503 ( .IN1(n8188), .IN2(n8189), .Q(n7848) );
  XOR2X1 U9504 ( .IN1(n9597), .IN2(n4574), .Q(n8189) );
  XOR2X1 U9505 ( .IN1(WX4580), .IN2(n4297), .Q(n8188) );
  NOR2X0 U9506 ( .IN1(n8190), .IN2(n8191), .QN(n8183) );
  NOR2X0 U9507 ( .IN1(DFF_547_n1), .IN2(n4760), .QN(n8191) );
  NOR2X0 U9508 ( .IN1(n4801), .IN2(n6294), .QN(n8190) );
  NAND2X0 U9509 ( .IN1(n5304), .IN2(n8616), .QN(n6294) );
  NAND2X0 U9510 ( .IN1(n8192), .IN2(n8193), .QN(WX3284) );
  NOR2X0 U9511 ( .IN1(n8194), .IN2(n8195), .QN(n8193) );
  NOR2X0 U9512 ( .IN1(n8196), .IN2(n4726), .QN(n8195) );
  NOR2X0 U9513 ( .IN1(n7857), .IN2(n4782), .QN(n8194) );
  XOR2X1 U9514 ( .IN1(n8197), .IN2(n8198), .Q(n7857) );
  XOR2X1 U9515 ( .IN1(n9598), .IN2(n4402), .Q(n8198) );
  XOR2X1 U9516 ( .IN1(WX4578), .IN2(n4299), .Q(n8197) );
  NOR2X0 U9517 ( .IN1(n8199), .IN2(n8200), .QN(n8192) );
  NOR2X0 U9518 ( .IN1(DFF_548_n1), .IN2(n4760), .QN(n8200) );
  NOR2X0 U9519 ( .IN1(n4800), .IN2(n6295), .QN(n8199) );
  NAND2X0 U9520 ( .IN1(n5304), .IN2(n8617), .QN(n6295) );
  NAND2X0 U9521 ( .IN1(n8201), .IN2(n8202), .QN(WX3282) );
  NOR2X0 U9522 ( .IN1(n8203), .IN2(n8204), .QN(n8202) );
  NOR2X0 U9523 ( .IN1(n8205), .IN2(n4726), .QN(n8204) );
  NOR2X0 U9524 ( .IN1(n7866), .IN2(n4781), .QN(n8203) );
  XOR2X1 U9525 ( .IN1(n8206), .IN2(n8207), .Q(n7866) );
  XOR2X1 U9526 ( .IN1(n9599), .IN2(n4573), .Q(n8207) );
  XOR2X1 U9527 ( .IN1(WX4576), .IN2(n4301), .Q(n8206) );
  NOR2X0 U9528 ( .IN1(n8208), .IN2(n8209), .QN(n8201) );
  NOR2X0 U9529 ( .IN1(DFF_549_n1), .IN2(n4760), .QN(n8209) );
  NOR2X0 U9530 ( .IN1(n4800), .IN2(n6296), .QN(n8208) );
  NAND2X0 U9531 ( .IN1(n5303), .IN2(n8618), .QN(n6296) );
  NAND2X0 U9532 ( .IN1(n8210), .IN2(n8211), .QN(WX3280) );
  NOR2X0 U9533 ( .IN1(n8212), .IN2(n8213), .QN(n8211) );
  NOR2X0 U9534 ( .IN1(n4731), .IN2(n8214), .QN(n8213) );
  NOR2X0 U9535 ( .IN1(n7875), .IN2(n4782), .QN(n8212) );
  XOR2X1 U9536 ( .IN1(n8215), .IN2(n8216), .Q(n7875) );
  XOR2X1 U9537 ( .IN1(n9600), .IN2(n4572), .Q(n8216) );
  XOR2X1 U9538 ( .IN1(WX4574), .IN2(n4303), .Q(n8215) );
  NOR2X0 U9539 ( .IN1(n8217), .IN2(n8218), .QN(n8210) );
  NOR2X0 U9540 ( .IN1(DFF_550_n1), .IN2(n4760), .QN(n8218) );
  NOR2X0 U9541 ( .IN1(n4800), .IN2(n6306), .QN(n8217) );
  NAND2X0 U9542 ( .IN1(n5303), .IN2(n8619), .QN(n6306) );
  NAND2X0 U9543 ( .IN1(n8219), .IN2(n8220), .QN(WX3278) );
  NOR2X0 U9544 ( .IN1(n8221), .IN2(n8222), .QN(n8220) );
  NOR2X0 U9545 ( .IN1(n8223), .IN2(n4726), .QN(n8222) );
  NOR2X0 U9546 ( .IN1(n7884), .IN2(n4782), .QN(n8221) );
  XOR2X1 U9547 ( .IN1(n8224), .IN2(n8225), .Q(n7884) );
  XOR2X1 U9548 ( .IN1(n9601), .IN2(n4571), .Q(n8225) );
  XOR2X1 U9549 ( .IN1(WX4572), .IN2(n4305), .Q(n8224) );
  NOR2X0 U9550 ( .IN1(n8226), .IN2(n8227), .QN(n8219) );
  NOR2X0 U9551 ( .IN1(DFF_551_n1), .IN2(n4760), .QN(n8227) );
  NOR2X0 U9552 ( .IN1(n4800), .IN2(n6307), .QN(n8226) );
  NAND2X0 U9553 ( .IN1(n5303), .IN2(n8620), .QN(n6307) );
  NAND2X0 U9554 ( .IN1(n8228), .IN2(n8229), .QN(WX3276) );
  NOR2X0 U9555 ( .IN1(n8230), .IN2(n8231), .QN(n8229) );
  NOR2X0 U9556 ( .IN1(n4729), .IN2(n8232), .QN(n8231) );
  NOR2X0 U9557 ( .IN1(n7893), .IN2(n4782), .QN(n8230) );
  XOR2X1 U9558 ( .IN1(n8233), .IN2(n8234), .Q(n7893) );
  XOR2X1 U9559 ( .IN1(n9602), .IN2(n4570), .Q(n8234) );
  XOR2X1 U9560 ( .IN1(WX4570), .IN2(n4307), .Q(n8233) );
  NOR2X0 U9561 ( .IN1(n8235), .IN2(n8236), .QN(n8228) );
  NOR2X0 U9562 ( .IN1(DFF_552_n1), .IN2(n4760), .QN(n8236) );
  NOR2X0 U9563 ( .IN1(n4800), .IN2(n6308), .QN(n8235) );
  NAND2X0 U9564 ( .IN1(n5303), .IN2(n8621), .QN(n6308) );
  NAND2X0 U9565 ( .IN1(n8237), .IN2(n8238), .QN(WX3274) );
  NOR2X0 U9566 ( .IN1(n8239), .IN2(n8240), .QN(n8238) );
  NOR2X0 U9567 ( .IN1(n8241), .IN2(n4725), .QN(n8240) );
  NOR2X0 U9568 ( .IN1(n7902), .IN2(n4780), .QN(n8239) );
  XOR2X1 U9569 ( .IN1(n8242), .IN2(n8243), .Q(n7902) );
  XOR2X1 U9570 ( .IN1(n9603), .IN2(n4569), .Q(n8243) );
  XOR2X1 U9571 ( .IN1(WX4568), .IN2(n4309), .Q(n8242) );
  NOR2X0 U9572 ( .IN1(n8244), .IN2(n8245), .QN(n8237) );
  NOR2X0 U9573 ( .IN1(DFF_553_n1), .IN2(n4760), .QN(n8245) );
  NOR2X0 U9574 ( .IN1(n4800), .IN2(n6309), .QN(n8244) );
  NAND2X0 U9575 ( .IN1(n5303), .IN2(n8622), .QN(n6309) );
  NAND2X0 U9576 ( .IN1(n8255), .IN2(n8256), .QN(WX3272) );
  NOR2X0 U9577 ( .IN1(n8273), .IN2(n8274), .QN(n8256) );
  NOR2X0 U9578 ( .IN1(n8291), .IN2(n4725), .QN(n8274) );
  NOR2X0 U9579 ( .IN1(n7911), .IN2(n4782), .QN(n8273) );
  XOR2X1 U9580 ( .IN1(n8292), .IN2(n8296), .Q(n7911) );
  XOR2X1 U9581 ( .IN1(n9604), .IN2(n4568), .Q(n8296) );
  XOR2X1 U9582 ( .IN1(WX4566), .IN2(n4311), .Q(n8292) );
  NOR2X0 U9583 ( .IN1(n8297), .IN2(n8298), .QN(n8255) );
  NOR2X0 U9584 ( .IN1(n4765), .IN2(n4705), .QN(n8298) );
  NOR2X0 U9585 ( .IN1(n4800), .IN2(n6310), .QN(n8297) );
  NAND2X0 U9586 ( .IN1(n5303), .IN2(n8623), .QN(n6310) );
  NAND2X0 U9587 ( .IN1(n8299), .IN2(n8300), .QN(WX3270) );
  NOR2X0 U9588 ( .IN1(n8301), .IN2(n8302), .QN(n8300) );
  NOR2X0 U9589 ( .IN1(n8303), .IN2(n4725), .QN(n8302) );
  NOR2X0 U9590 ( .IN1(n4786), .IN2(n7920), .QN(n8301) );
  XNOR2X1 U9591 ( .IN1(n8308), .IN2(n8309), .Q(n7920) );
  XOR2X1 U9592 ( .IN1(test_so41), .IN2(n9605), .Q(n8309) );
  XOR2X1 U9593 ( .IN1(WX4564), .IN2(n4313), .Q(n8308) );
  NOR2X0 U9594 ( .IN1(n8326), .IN2(n8327), .QN(n8299) );
  NOR2X0 U9595 ( .IN1(DFF_555_n1), .IN2(n4760), .QN(n8327) );
  NOR2X0 U9596 ( .IN1(n4800), .IN2(n6311), .QN(n8326) );
  NAND2X0 U9597 ( .IN1(n5302), .IN2(n8624), .QN(n6311) );
  NAND2X0 U9598 ( .IN1(n8344), .IN2(n8345), .QN(WX3268) );
  NOR2X0 U9599 ( .IN1(n8354), .IN2(n8355), .QN(n8345) );
  NOR2X0 U9600 ( .IN1(n4729), .IN2(n8356), .QN(n8355) );
  NOR2X0 U9601 ( .IN1(n7929), .IN2(n4783), .QN(n8354) );
  XOR2X1 U9602 ( .IN1(n8357), .IN2(n8358), .Q(n7929) );
  XOR2X1 U9603 ( .IN1(n9606), .IN2(n4567), .Q(n8358) );
  XOR2X1 U9604 ( .IN1(WX4562), .IN2(n4315), .Q(n8357) );
  NOR2X0 U9605 ( .IN1(n8359), .IN2(n8360), .QN(n8344) );
  NOR2X0 U9606 ( .IN1(DFF_556_n1), .IN2(n4759), .QN(n8360) );
  NOR2X0 U9607 ( .IN1(n4800), .IN2(n6312), .QN(n8359) );
  NAND2X0 U9608 ( .IN1(n5302), .IN2(n8625), .QN(n6312) );
  NAND2X0 U9609 ( .IN1(n8361), .IN2(n8362), .QN(WX3266) );
  NOR2X0 U9610 ( .IN1(n8379), .IN2(n8380), .QN(n8362) );
  NOR2X0 U9611 ( .IN1(n8397), .IN2(n4725), .QN(n8380) );
  NOR2X0 U9612 ( .IN1(n4786), .IN2(n7938), .QN(n8379) );
  XNOR2X1 U9613 ( .IN1(n8398), .IN2(n8412), .Q(n7938) );
  XOR2X1 U9614 ( .IN1(test_so39), .IN2(n9607), .Q(n8412) );
  XOR2X1 U9615 ( .IN1(WX4560), .IN2(n4566), .Q(n8398) );
  NOR2X0 U9616 ( .IN1(n8413), .IN2(n8414), .QN(n8361) );
  NOR2X0 U9617 ( .IN1(DFF_557_n1), .IN2(n4759), .QN(n8414) );
  NOR2X0 U9618 ( .IN1(n4800), .IN2(n6313), .QN(n8413) );
  NAND2X0 U9619 ( .IN1(n5302), .IN2(n8626), .QN(n6313) );
  NAND2X0 U9620 ( .IN1(n8415), .IN2(n8416), .QN(WX3264) );
  NOR2X0 U9621 ( .IN1(n8417), .IN2(n8418), .QN(n8416) );
  NOR2X0 U9622 ( .IN1(n8419), .IN2(n4725), .QN(n8418) );
  NOR2X0 U9623 ( .IN1(n7947), .IN2(n4783), .QN(n8417) );
  XOR2X1 U9624 ( .IN1(n8420), .IN2(n8432), .Q(n7947) );
  XOR2X1 U9625 ( .IN1(n9608), .IN2(n4565), .Q(n8432) );
  XOR2X1 U9626 ( .IN1(WX4558), .IN2(n4318), .Q(n8420) );
  NOR2X0 U9627 ( .IN1(n8433), .IN2(n8450), .QN(n8415) );
  NOR2X0 U9628 ( .IN1(DFF_558_n1), .IN2(n4759), .QN(n8450) );
  NOR2X0 U9629 ( .IN1(n4800), .IN2(n6314), .QN(n8433) );
  NAND2X0 U9630 ( .IN1(n5302), .IN2(n8627), .QN(n6314) );
  NAND2X0 U9631 ( .IN1(n8451), .IN2(n8468), .QN(WX3262) );
  NOR2X0 U9632 ( .IN1(n8469), .IN2(n8471), .QN(n8468) );
  NOR2X0 U9633 ( .IN1(n8472), .IN2(n4725), .QN(n8471) );
  NOR2X0 U9634 ( .IN1(n4786), .IN2(n7956), .QN(n8469) );
  XNOR2X1 U9635 ( .IN1(n8473), .IN2(n8474), .Q(n7956) );
  XOR2X1 U9636 ( .IN1(test_so37), .IN2(n9609), .Q(n8474) );
  XOR2X1 U9637 ( .IN1(WX4556), .IN2(n4564), .Q(n8473) );
  NOR2X0 U9638 ( .IN1(n8475), .IN2(n8476), .QN(n8451) );
  NOR2X0 U9639 ( .IN1(DFF_559_n1), .IN2(n4759), .QN(n8476) );
  NOR2X0 U9640 ( .IN1(n4800), .IN2(n6327), .QN(n8475) );
  NAND2X0 U9641 ( .IN1(n5302), .IN2(n8628), .QN(n6327) );
  NAND2X0 U9642 ( .IN1(n8477), .IN2(n8478), .QN(WX3260) );
  NOR2X0 U9643 ( .IN1(n8485), .IN2(n8486), .QN(n8478) );
  NOR2X0 U9644 ( .IN1(n4730), .IN2(n8503), .QN(n8486) );
  NOR2X0 U9645 ( .IN1(n7965), .IN2(n4782), .QN(n8485) );
  XOR2X1 U9646 ( .IN1(n8504), .IN2(n8521), .Q(n7965) );
  XOR2X1 U9647 ( .IN1(n4104), .IN2(n5253), .Q(n8521) );
  XOR2X1 U9648 ( .IN1(n8522), .IN2(n4401), .Q(n8504) );
  XOR2X1 U9649 ( .IN1(WX4682), .IN2(n9610), .Q(n8522) );
  NOR2X0 U9650 ( .IN1(n8529), .IN2(n8530), .QN(n8477) );
  NOR2X0 U9651 ( .IN1(DFF_560_n1), .IN2(n4759), .QN(n8530) );
  NOR2X0 U9652 ( .IN1(n4799), .IN2(n6328), .QN(n8529) );
  NAND2X0 U9653 ( .IN1(n5302), .IN2(n8629), .QN(n6328) );
  NAND2X0 U9654 ( .IN1(n8531), .IN2(n8532), .QN(WX3258) );
  NOR2X0 U9655 ( .IN1(n8533), .IN2(n8534), .QN(n8532) );
  NOR2X0 U9656 ( .IN1(n8535), .IN2(n4725), .QN(n8534) );
  NOR2X0 U9657 ( .IN1(n4786), .IN2(n7975), .QN(n8533) );
  XNOR2X1 U9658 ( .IN1(n8536), .IN2(n8538), .Q(n7975) );
  XOR2X1 U9659 ( .IN1(n4105), .IN2(n5253), .Q(n8538) );
  XOR2X1 U9660 ( .IN1(n8539), .IN2(n4563), .Q(n8536) );
  XOR2X1 U9661 ( .IN1(WX4616), .IN2(test_so35), .Q(n8539) );
  NOR2X0 U9662 ( .IN1(n8556), .IN2(n8557), .QN(n8531) );
  NOR2X0 U9663 ( .IN1(DFF_561_n1), .IN2(n4759), .QN(n8557) );
  NOR2X0 U9664 ( .IN1(n4799), .IN2(n6329), .QN(n8556) );
  NAND2X0 U9665 ( .IN1(n5301), .IN2(n8630), .QN(n6329) );
  NAND2X0 U9666 ( .IN1(n8574), .IN2(n8575), .QN(WX3256) );
  NOR2X0 U9667 ( .IN1(n8587), .IN2(n8588), .QN(n8575) );
  NOR2X0 U9668 ( .IN1(n8589), .IN2(n4725), .QN(n8588) );
  NOR2X0 U9669 ( .IN1(n7985), .IN2(n4783), .QN(n8587) );
  XOR2X1 U9670 ( .IN1(n8590), .IN2(n8591), .Q(n7985) );
  XOR2X1 U9671 ( .IN1(n4106), .IN2(n5253), .Q(n8591) );
  XOR2X1 U9672 ( .IN1(n8592), .IN2(n4562), .Q(n8590) );
  XOR2X1 U9673 ( .IN1(WX4678), .IN2(n9611), .Q(n8592) );
  NOR2X0 U9674 ( .IN1(n8593), .IN2(n8594), .QN(n8574) );
  NOR2X0 U9675 ( .IN1(DFF_562_n1), .IN2(n4759), .QN(n8594) );
  NOR2X0 U9676 ( .IN1(n4799), .IN2(n6330), .QN(n8593) );
  NAND2X0 U9677 ( .IN1(n5301), .IN2(n8631), .QN(n6330) );
  NAND2X0 U9678 ( .IN1(n8595), .IN2(n8596), .QN(WX3254) );
  NOR2X0 U9679 ( .IN1(n8614), .IN2(n8615), .QN(n8596) );
  NOR2X0 U9680 ( .IN1(n8633), .IN2(n4725), .QN(n8615) );
  NOR2X0 U9681 ( .IN1(n7995), .IN2(n4782), .QN(n8614) );
  XOR2X1 U9682 ( .IN1(n8634), .IN2(n8645), .Q(n7995) );
  XOR2X1 U9683 ( .IN1(n4107), .IN2(n5254), .Q(n8645) );
  XOR2X1 U9684 ( .IN1(n8646), .IN2(n4561), .Q(n8634) );
  XOR2X1 U9685 ( .IN1(WX4676), .IN2(n9612), .Q(n8646) );
  NOR2X0 U9686 ( .IN1(n8647), .IN2(n8648), .QN(n8595) );
  NOR2X0 U9687 ( .IN1(DFF_563_n1), .IN2(n4759), .QN(n8648) );
  NOR2X0 U9688 ( .IN1(n4799), .IN2(n6331), .QN(n8647) );
  NAND2X0 U9689 ( .IN1(n5301), .IN2(n8632), .QN(n6331) );
  NAND2X0 U9690 ( .IN1(n8649), .IN2(n8650), .QN(WX3252) );
  NOR2X0 U9691 ( .IN1(n8651), .IN2(n8652), .QN(n8650) );
  NOR2X0 U9692 ( .IN1(n8659), .IN2(n4725), .QN(n8652) );
  NOR2X0 U9693 ( .IN1(n8005), .IN2(n4783), .QN(n8651) );
  XOR2X1 U9694 ( .IN1(n8660), .IN2(n8678), .Q(n8005) );
  XOR2X1 U9695 ( .IN1(n4108), .IN2(n5254), .Q(n8678) );
  XOR2X1 U9696 ( .IN1(n8679), .IN2(n4560), .Q(n8660) );
  XOR2X1 U9697 ( .IN1(WX4674), .IN2(n9613), .Q(n8679) );
  NOR2X0 U9698 ( .IN1(n8697), .IN2(n8698), .QN(n8649) );
  NOR2X0 U9699 ( .IN1(DFF_564_n1), .IN2(n4759), .QN(n8698) );
  NOR2X0 U9700 ( .IN1(n4799), .IN2(n6332), .QN(n8697) );
  NAND2X0 U9701 ( .IN1(test_so22), .IN2(n5324), .QN(n6332) );
  NAND2X0 U9702 ( .IN1(n8703), .IN2(n8704), .QN(WX3250) );
  NOR2X0 U9703 ( .IN1(n8705), .IN2(n8706), .QN(n8704) );
  NOR2X0 U9704 ( .IN1(n8707), .IN2(n4725), .QN(n8706) );
  NOR2X0 U9705 ( .IN1(n8015), .IN2(n4783), .QN(n8705) );
  XOR2X1 U9706 ( .IN1(n8708), .IN2(n8709), .Q(n8015) );
  XOR2X1 U9707 ( .IN1(n4109), .IN2(n5254), .Q(n8709) );
  XOR2X1 U9708 ( .IN1(n8710), .IN2(n4559), .Q(n8708) );
  XOR2X1 U9709 ( .IN1(WX4672), .IN2(n9614), .Q(n8710) );
  NOR2X0 U9710 ( .IN1(n8711), .IN2(n8712), .QN(n8703) );
  NOR2X0 U9711 ( .IN1(DFF_565_n1), .IN2(n4759), .QN(n8712) );
  NOR2X0 U9712 ( .IN1(n4799), .IN2(n6333), .QN(n8711) );
  NAND2X0 U9713 ( .IN1(n5301), .IN2(n8635), .QN(n6333) );
  NAND2X0 U9714 ( .IN1(n8713), .IN2(n8714), .QN(WX3248) );
  NOR2X0 U9715 ( .IN1(n8715), .IN2(n8716), .QN(n8714) );
  NOR2X0 U9716 ( .IN1(n8717), .IN2(n4725), .QN(n8716) );
  NOR2X0 U9717 ( .IN1(n8025), .IN2(n4782), .QN(n8715) );
  XOR2X1 U9718 ( .IN1(n8718), .IN2(n8719), .Q(n8025) );
  XOR2X1 U9719 ( .IN1(n4110), .IN2(n5254), .Q(n8719) );
  XOR2X1 U9720 ( .IN1(n8720), .IN2(n4558), .Q(n8718) );
  XOR2X1 U9721 ( .IN1(WX4670), .IN2(n9615), .Q(n8720) );
  NOR2X0 U9722 ( .IN1(n8721), .IN2(n8722), .QN(n8713) );
  NOR2X0 U9723 ( .IN1(DFF_566_n1), .IN2(n4759), .QN(n8722) );
  NOR2X0 U9724 ( .IN1(n4799), .IN2(n6334), .QN(n8721) );
  NAND2X0 U9725 ( .IN1(n5301), .IN2(n8636), .QN(n6334) );
  NAND2X0 U9726 ( .IN1(n8723), .IN2(n8724), .QN(WX3246) );
  NOR2X0 U9727 ( .IN1(n8725), .IN2(n8726), .QN(n8724) );
  NOR2X0 U9728 ( .IN1(n4732), .IN2(n8727), .QN(n8726) );
  NOR2X0 U9729 ( .IN1(n8035), .IN2(n4782), .QN(n8725) );
  XOR2X1 U9730 ( .IN1(n8728), .IN2(n8729), .Q(n8035) );
  XOR2X1 U9731 ( .IN1(n4111), .IN2(n5254), .Q(n8729) );
  XOR2X1 U9732 ( .IN1(n8730), .IN2(n4557), .Q(n8728) );
  XOR2X1 U9733 ( .IN1(WX4668), .IN2(n9616), .Q(n8730) );
  NOR2X0 U9734 ( .IN1(n8731), .IN2(n8732), .QN(n8723) );
  NOR2X0 U9735 ( .IN1(DFF_567_n1), .IN2(n4759), .QN(n8732) );
  NOR2X0 U9736 ( .IN1(n4799), .IN2(n6344), .QN(n8731) );
  NAND2X0 U9737 ( .IN1(n5301), .IN2(n8637), .QN(n6344) );
  NAND2X0 U9738 ( .IN1(n8733), .IN2(n8734), .QN(WX3244) );
  NOR2X0 U9739 ( .IN1(n8735), .IN2(n8736), .QN(n8734) );
  NOR2X0 U9740 ( .IN1(n8737), .IN2(n4724), .QN(n8736) );
  NOR2X0 U9741 ( .IN1(n8045), .IN2(n4783), .QN(n8735) );
  XOR2X1 U9742 ( .IN1(n8738), .IN2(n8739), .Q(n8045) );
  XOR2X1 U9743 ( .IN1(n4112), .IN2(n5254), .Q(n8739) );
  XOR2X1 U9744 ( .IN1(n8740), .IN2(n4556), .Q(n8738) );
  XOR2X1 U9745 ( .IN1(WX4666), .IN2(n9617), .Q(n8740) );
  NOR2X0 U9746 ( .IN1(n8741), .IN2(n8742), .QN(n8733) );
  NOR2X0 U9747 ( .IN1(DFF_568_n1), .IN2(n4758), .QN(n8742) );
  NOR2X0 U9748 ( .IN1(n4799), .IN2(n6345), .QN(n8741) );
  NAND2X0 U9749 ( .IN1(n5300), .IN2(n8638), .QN(n6345) );
  NAND2X0 U9750 ( .IN1(n8743), .IN2(n8744), .QN(WX3242) );
  NOR2X0 U9751 ( .IN1(n8745), .IN2(n8746), .QN(n8744) );
  NOR2X0 U9752 ( .IN1(n8747), .IN2(n4724), .QN(n8746) );
  NOR2X0 U9753 ( .IN1(n8055), .IN2(n4783), .QN(n8745) );
  XOR2X1 U9754 ( .IN1(n8748), .IN2(n8749), .Q(n8055) );
  XOR2X1 U9755 ( .IN1(n4113), .IN2(n5254), .Q(n8749) );
  XOR2X1 U9756 ( .IN1(n8750), .IN2(n4555), .Q(n8748) );
  XOR2X1 U9757 ( .IN1(WX4664), .IN2(n9618), .Q(n8750) );
  NOR2X0 U9758 ( .IN1(n8751), .IN2(n8752), .QN(n8743) );
  NOR2X0 U9759 ( .IN1(DFF_569_n1), .IN2(n4758), .QN(n8752) );
  NOR2X0 U9760 ( .IN1(n4799), .IN2(n6346), .QN(n8751) );
  NAND2X0 U9761 ( .IN1(n5300), .IN2(n8639), .QN(n6346) );
  NAND2X0 U9762 ( .IN1(n8753), .IN2(n8754), .QN(WX3240) );
  NOR2X0 U9763 ( .IN1(n8755), .IN2(n8756), .QN(n8754) );
  NOR2X0 U9764 ( .IN1(n4730), .IN2(n8757), .QN(n8756) );
  NOR2X0 U9765 ( .IN1(n8065), .IN2(n4784), .QN(n8755) );
  XOR2X1 U9766 ( .IN1(n8758), .IN2(n8759), .Q(n8065) );
  XOR2X1 U9767 ( .IN1(n4114), .IN2(n5254), .Q(n8759) );
  XOR2X1 U9768 ( .IN1(n8760), .IN2(n4554), .Q(n8758) );
  XOR2X1 U9769 ( .IN1(WX4662), .IN2(n9619), .Q(n8760) );
  NOR2X0 U9770 ( .IN1(n8761), .IN2(n8762), .QN(n8753) );
  NOR2X0 U9771 ( .IN1(DFF_570_n1), .IN2(n4758), .QN(n8762) );
  NOR2X0 U9772 ( .IN1(n4799), .IN2(n6347), .QN(n8761) );
  NAND2X0 U9773 ( .IN1(n5300), .IN2(n8640), .QN(n6347) );
  NAND2X0 U9774 ( .IN1(n8763), .IN2(n8764), .QN(WX3238) );
  NOR2X0 U9775 ( .IN1(n8765), .IN2(n8766), .QN(n8764) );
  NOR2X0 U9776 ( .IN1(n8767), .IN2(n4724), .QN(n8766) );
  NOR2X0 U9777 ( .IN1(n8075), .IN2(n4783), .QN(n8765) );
  XOR2X1 U9778 ( .IN1(n8768), .IN2(n8769), .Q(n8075) );
  XOR2X1 U9779 ( .IN1(n4115), .IN2(n5254), .Q(n8769) );
  XOR2X1 U9780 ( .IN1(n8770), .IN2(n4553), .Q(n8768) );
  XOR2X1 U9781 ( .IN1(WX4660), .IN2(n9620), .Q(n8770) );
  NOR2X0 U9782 ( .IN1(n8771), .IN2(n8772), .QN(n8763) );
  NOR2X0 U9783 ( .IN1(n4765), .IN2(n4702), .QN(n8772) );
  NOR2X0 U9784 ( .IN1(n4799), .IN2(n6348), .QN(n8771) );
  NAND2X0 U9785 ( .IN1(n5300), .IN2(n8641), .QN(n6348) );
  NAND2X0 U9786 ( .IN1(n8773), .IN2(n8774), .QN(WX3236) );
  NOR2X0 U9787 ( .IN1(n8775), .IN2(n8776), .QN(n8774) );
  NOR2X0 U9788 ( .IN1(n8777), .IN2(n4724), .QN(n8776) );
  NOR2X0 U9789 ( .IN1(n4786), .IN2(n8085), .QN(n8775) );
  XNOR2X1 U9790 ( .IN1(n8778), .IN2(n8779), .Q(n8085) );
  XOR2X1 U9791 ( .IN1(n4116), .IN2(n5254), .Q(n8779) );
  XOR2X1 U9792 ( .IN1(WX4594), .IN2(n8780), .Q(n8778) );
  XOR2X1 U9793 ( .IN1(test_so40), .IN2(n9621), .Q(n8780) );
  NOR2X0 U9794 ( .IN1(n8781), .IN2(n8782), .QN(n8773) );
  NOR2X0 U9795 ( .IN1(DFF_572_n1), .IN2(n4758), .QN(n8782) );
  NOR2X0 U9796 ( .IN1(n4799), .IN2(n6349), .QN(n8781) );
  NAND2X0 U9797 ( .IN1(n5300), .IN2(n8642), .QN(n6349) );
  NAND2X0 U9798 ( .IN1(n8783), .IN2(n8784), .QN(WX3234) );
  NOR2X0 U9799 ( .IN1(n8785), .IN2(n8786), .QN(n8784) );
  NOR2X0 U9800 ( .IN1(n8787), .IN2(n4724), .QN(n8786) );
  NOR2X0 U9801 ( .IN1(n8095), .IN2(n4784), .QN(n8785) );
  XOR2X1 U9802 ( .IN1(n8788), .IN2(n8789), .Q(n8095) );
  XOR2X1 U9803 ( .IN1(n4117), .IN2(n5254), .Q(n8789) );
  XOR2X1 U9804 ( .IN1(n8790), .IN2(n4552), .Q(n8788) );
  XOR2X1 U9805 ( .IN1(WX4656), .IN2(n9622), .Q(n8790) );
  NOR2X0 U9806 ( .IN1(n8791), .IN2(n8792), .QN(n8783) );
  NOR2X0 U9807 ( .IN1(DFF_573_n1), .IN2(n4758), .QN(n8792) );
  NOR2X0 U9808 ( .IN1(n4798), .IN2(n6350), .QN(n8791) );
  NAND2X0 U9809 ( .IN1(n5300), .IN2(n8643), .QN(n6350) );
  NAND2X0 U9810 ( .IN1(n8793), .IN2(n8794), .QN(WX3232) );
  NOR2X0 U9811 ( .IN1(n8795), .IN2(n8796), .QN(n8794) );
  NOR2X0 U9812 ( .IN1(n4731), .IN2(n8797), .QN(n8796) );
  NOR2X0 U9813 ( .IN1(n4786), .IN2(n8105), .QN(n8795) );
  XNOR2X1 U9814 ( .IN1(n8798), .IN2(n8799), .Q(n8105) );
  XOR2X1 U9815 ( .IN1(n4551), .IN2(n5254), .Q(n8799) );
  XOR2X1 U9816 ( .IN1(n8800), .IN2(n9625), .Q(n8798) );
  XOR2X1 U9817 ( .IN1(n9624), .IN2(n9623), .Q(n8800) );
  NOR2X0 U9818 ( .IN1(n8801), .IN2(n8802), .QN(n8793) );
  NOR2X0 U9819 ( .IN1(DFF_574_n1), .IN2(n4758), .QN(n8802) );
  NOR2X0 U9820 ( .IN1(n4798), .IN2(n6351), .QN(n8801) );
  NAND2X0 U9821 ( .IN1(n5299), .IN2(n8644), .QN(n6351) );
  NAND2X0 U9822 ( .IN1(n8803), .IN2(n8804), .QN(WX3230) );
  NOR2X0 U9823 ( .IN1(n8805), .IN2(n8806), .QN(n8804) );
  NOR2X0 U9824 ( .IN1(n8807), .IN2(n4724), .QN(n8806) );
  NOR2X0 U9825 ( .IN1(n8115), .IN2(n4784), .QN(n8805) );
  XOR2X1 U9826 ( .IN1(n8808), .IN2(n8809), .Q(n8115) );
  XOR2X1 U9827 ( .IN1(n4036), .IN2(n5255), .Q(n8809) );
  XOR2X1 U9828 ( .IN1(n8810), .IN2(n4550), .Q(n8808) );
  XOR2X1 U9829 ( .IN1(WX4652), .IN2(n9626), .Q(n8810) );
  NOR2X0 U9830 ( .IN1(n8811), .IN2(n8812), .QN(n8803) );
  NOR2X0 U9831 ( .IN1(n4386), .IN2(n6717), .QN(n8812) );
  NOR2X0 U9832 ( .IN1(DFF_575_n1), .IN2(n4758), .QN(n8811) );
  NOR2X0 U9833 ( .IN1(n5420), .IN2(WX3071), .QN(WX3132) );
  NOR2X0 U9834 ( .IN1(n5420), .IN2(n8813), .QN(WX2619) );
  XOR2X1 U9835 ( .IN1(n4603), .IN2(DFF_382_n1), .Q(n8813) );
  NOR2X0 U9836 ( .IN1(n5421), .IN2(n8814), .QN(WX2617) );
  XOR2X1 U9837 ( .IN1(n4604), .IN2(DFF_381_n1), .Q(n8814) );
  NOR2X0 U9838 ( .IN1(n5420), .IN2(n8815), .QN(WX2615) );
  XOR2X1 U9839 ( .IN1(n4605), .IN2(DFF_380_n1), .Q(n8815) );
  NOR2X0 U9840 ( .IN1(n5421), .IN2(n8816), .QN(WX2613) );
  XNOR2X1 U9841 ( .IN1(DFF_379_n1), .IN2(test_so18), .Q(n8816) );
  NOR2X0 U9842 ( .IN1(n5421), .IN2(n8817), .QN(WX2611) );
  XOR2X1 U9843 ( .IN1(n4606), .IN2(DFF_378_n1), .Q(n8817) );
  NOR2X0 U9844 ( .IN1(n5420), .IN2(n8818), .QN(WX2609) );
  XOR2X1 U9845 ( .IN1(n4607), .IN2(n4704), .Q(n8818) );
  NOR2X0 U9846 ( .IN1(n5422), .IN2(n8819), .QN(WX2607) );
  XOR2X1 U9847 ( .IN1(n4608), .IN2(DFF_376_n1), .Q(n8819) );
  NOR2X0 U9848 ( .IN1(n5420), .IN2(n8820), .QN(WX2605) );
  XOR2X1 U9849 ( .IN1(n4609), .IN2(DFF_375_n1), .Q(n8820) );
  NOR2X0 U9850 ( .IN1(n5420), .IN2(n8821), .QN(WX2603) );
  XOR2X1 U9851 ( .IN1(n4610), .IN2(DFF_374_n1), .Q(n8821) );
  NOR2X0 U9852 ( .IN1(n5421), .IN2(n8822), .QN(WX2601) );
  XOR2X1 U9853 ( .IN1(n4611), .IN2(DFF_373_n1), .Q(n8822) );
  NOR2X0 U9854 ( .IN1(n5421), .IN2(n8823), .QN(WX2599) );
  XOR2X1 U9855 ( .IN1(n4612), .IN2(DFF_372_n1), .Q(n8823) );
  NOR2X0 U9856 ( .IN1(n5419), .IN2(n8824), .QN(WX2597) );
  XOR2X1 U9857 ( .IN1(n4613), .IN2(DFF_371_n1), .Q(n8824) );
  NOR2X0 U9858 ( .IN1(n5420), .IN2(n8825), .QN(WX2595) );
  XOR2X1 U9859 ( .IN1(n4614), .IN2(DFF_370_n1), .Q(n8825) );
  NOR2X0 U9860 ( .IN1(n5419), .IN2(n8826), .QN(WX2593) );
  XOR2X1 U9861 ( .IN1(n4615), .IN2(DFF_369_n1), .Q(n8826) );
  NOR2X0 U9862 ( .IN1(n5421), .IN2(n8827), .QN(WX2591) );
  XOR2X1 U9863 ( .IN1(n4616), .IN2(DFF_368_n1), .Q(n8827) );
  NOR2X0 U9864 ( .IN1(n5419), .IN2(n8828), .QN(WX2589) );
  XNOR2X1 U9865 ( .IN1(DFF_367_n1), .IN2(n8829), .Q(n8828) );
  XOR2X1 U9866 ( .IN1(n4406), .IN2(DFF_383_n1), .Q(n8829) );
  NOR2X0 U9867 ( .IN1(n5419), .IN2(n8830), .QN(WX2587) );
  XOR2X1 U9868 ( .IN1(n4617), .IN2(DFF_366_n1), .Q(n8830) );
  NOR2X0 U9869 ( .IN1(n5421), .IN2(n8831), .QN(WX2585) );
  XOR2X1 U9870 ( .IN1(n4618), .IN2(DFF_365_n1), .Q(n8831) );
  NOR2X0 U9871 ( .IN1(n5420), .IN2(n8832), .QN(WX2583) );
  XOR2X1 U9872 ( .IN1(n4619), .IN2(DFF_364_n1), .Q(n8832) );
  NOR2X0 U9873 ( .IN1(n5419), .IN2(n8833), .QN(WX2581) );
  XOR2X1 U9874 ( .IN1(n4620), .IN2(DFF_363_n1), .Q(n8833) );
  NOR2X0 U9875 ( .IN1(n5419), .IN2(n8834), .QN(WX2579) );
  XNOR2X1 U9876 ( .IN1(DFF_362_n1), .IN2(n8835), .Q(n8834) );
  XOR2X1 U9877 ( .IN1(n4407), .IN2(DFF_383_n1), .Q(n8835) );
  NOR2X0 U9878 ( .IN1(n5420), .IN2(n8836), .QN(WX2577) );
  XNOR2X1 U9879 ( .IN1(DFF_361_n1), .IN2(test_so19), .Q(n8836) );
  NOR2X0 U9880 ( .IN1(n5420), .IN2(n8837), .QN(WX2575) );
  XOR2X1 U9881 ( .IN1(n4621), .IN2(DFF_360_n1), .Q(n8837) );
  NOR2X0 U9882 ( .IN1(n5419), .IN2(n8838), .QN(WX2573) );
  XOR2X1 U9883 ( .IN1(n4622), .IN2(n4703), .Q(n8838) );
  NOR2X0 U9884 ( .IN1(n5420), .IN2(n8839), .QN(WX2571) );
  XOR2X1 U9885 ( .IN1(n4623), .IN2(DFF_358_n1), .Q(n8839) );
  NOR2X0 U9886 ( .IN1(n5419), .IN2(n8840), .QN(WX2569) );
  XOR2X1 U9887 ( .IN1(n4624), .IN2(DFF_357_n1), .Q(n8840) );
  NOR2X0 U9888 ( .IN1(n5419), .IN2(n8841), .QN(WX2567) );
  XOR2X1 U9889 ( .IN1(n4625), .IN2(DFF_356_n1), .Q(n8841) );
  NOR2X0 U9890 ( .IN1(n5419), .IN2(n8842), .QN(WX2565) );
  XNOR2X1 U9891 ( .IN1(DFF_355_n1), .IN2(n8843), .Q(n8842) );
  XOR2X1 U9892 ( .IN1(n4408), .IN2(DFF_383_n1), .Q(n8843) );
  NOR2X0 U9893 ( .IN1(n5419), .IN2(n8844), .QN(WX2563) );
  XOR2X1 U9894 ( .IN1(n4626), .IN2(DFF_354_n1), .Q(n8844) );
  NOR2X0 U9895 ( .IN1(n5422), .IN2(n8845), .QN(WX2561) );
  XOR2X1 U9896 ( .IN1(n4627), .IN2(DFF_353_n1), .Q(n8845) );
  NOR2X0 U9897 ( .IN1(n5420), .IN2(n8846), .QN(WX2559) );
  XOR2X1 U9898 ( .IN1(n4628), .IN2(DFF_352_n1), .Q(n8846) );
  NOR2X0 U9899 ( .IN1(n5419), .IN2(n8847), .QN(WX2557) );
  XOR2X1 U9900 ( .IN1(n4416), .IN2(DFF_383_n1), .Q(n8847) );
  NOR2X0 U9901 ( .IN1(n9659), .IN2(n5350), .QN(WX2031) );
  NOR2X0 U9902 ( .IN1(n9660), .IN2(n5350), .QN(WX2029) );
  NOR2X0 U9903 ( .IN1(n9662), .IN2(n5350), .QN(WX2027) );
  NOR2X0 U9904 ( .IN1(n9666), .IN2(n5350), .QN(WX2025) );
  NOR2X0 U9905 ( .IN1(n9668), .IN2(n5350), .QN(WX2023) );
  NOR2X0 U9906 ( .IN1(n9670), .IN2(n5350), .QN(WX2021) );
  NOR2X0 U9907 ( .IN1(n5420), .IN2(n4711), .QN(WX2019) );
  NOR2X0 U9908 ( .IN1(n9673), .IN2(n5350), .QN(WX2017) );
  NOR2X0 U9909 ( .IN1(n9675), .IN2(n5349), .QN(WX2015) );
  NOR2X0 U9910 ( .IN1(n9677), .IN2(n5349), .QN(WX2013) );
  NOR2X0 U9911 ( .IN1(n9679), .IN2(n5349), .QN(WX2011) );
  NOR2X0 U9912 ( .IN1(n9683), .IN2(n5349), .QN(WX2009) );
  NOR2X0 U9913 ( .IN1(n9685), .IN2(n5349), .QN(WX2007) );
  NOR2X0 U9914 ( .IN1(n9687), .IN2(n5349), .QN(WX2005) );
  NOR2X0 U9915 ( .IN1(n9689), .IN2(n5349), .QN(WX2003) );
  NOR2X0 U9916 ( .IN1(n9694), .IN2(n5349), .QN(WX2001) );
  NAND2X0 U9917 ( .IN1(n8848), .IN2(n8849), .QN(WX1999) );
  NOR2X0 U9918 ( .IN1(n8850), .IN2(n8851), .QN(n8849) );
  NOR2X0 U9919 ( .IN1(n8160), .IN2(n4784), .QN(n8851) );
  XOR2X1 U9920 ( .IN1(n8852), .IN2(n8853), .Q(n8160) );
  XOR2X1 U9921 ( .IN1(n9628), .IN2(n4415), .Q(n8853) );
  XOR2X1 U9922 ( .IN1(WX3293), .IN2(n4321), .Q(n8852) );
  NOR2X0 U9923 ( .IN1(n4730), .IN2(n6119), .QN(n8850) );
  XNOR2X1 U9924 ( .IN1(n8854), .IN2(n8855), .Q(n6119) );
  XOR2X1 U9925 ( .IN1(test_so16), .IN2(n9627), .Q(n8855) );
  XOR2X1 U9926 ( .IN1(WX2000), .IN2(n4416), .Q(n8854) );
  NOR2X0 U9927 ( .IN1(n8856), .IN2(n8857), .QN(n8848) );
  NOR2X0 U9928 ( .IN1(DFF_352_n1), .IN2(n4758), .QN(n8857) );
  NOR2X0 U9929 ( .IN1(n4798), .IN2(n5635), .QN(n8856) );
  NAND2X0 U9930 ( .IN1(n5299), .IN2(n8670), .QN(n5635) );
  NAND2X0 U9931 ( .IN1(n8858), .IN2(n8859), .QN(WX1997) );
  NOR2X0 U9932 ( .IN1(n8860), .IN2(n8861), .QN(n8859) );
  NOR2X0 U9933 ( .IN1(n8169), .IN2(n4783), .QN(n8861) );
  XOR2X1 U9934 ( .IN1(n8862), .IN2(n8863), .Q(n8169) );
  XOR2X1 U9935 ( .IN1(n9630), .IN2(n4602), .Q(n8863) );
  XOR2X1 U9936 ( .IN1(WX3291), .IN2(n4323), .Q(n8862) );
  NOR2X0 U9937 ( .IN1(n8864), .IN2(n4724), .QN(n8860) );
  INVX0 U9938 ( .INP(n6128), .ZN(n8864) );
  XNOR2X1 U9939 ( .IN1(n8865), .IN2(n8866), .Q(n6128) );
  XOR2X1 U9940 ( .IN1(n9629), .IN2(n4628), .Q(n8866) );
  XOR2X1 U9941 ( .IN1(WX1998), .IN2(n4352), .Q(n8865) );
  NOR2X0 U9942 ( .IN1(n8867), .IN2(n8868), .QN(n8858) );
  NOR2X0 U9943 ( .IN1(DFF_353_n1), .IN2(n4758), .QN(n8868) );
  NOR2X0 U9944 ( .IN1(n4798), .IN2(n5636), .QN(n8867) );
  NAND2X0 U9945 ( .IN1(n5299), .IN2(n8671), .QN(n5636) );
  NAND2X0 U9946 ( .IN1(n8869), .IN2(n8870), .QN(WX1995) );
  NOR2X0 U9947 ( .IN1(n8871), .IN2(n8872), .QN(n8870) );
  NOR2X0 U9948 ( .IN1(n8178), .IN2(n4784), .QN(n8872) );
  XOR2X1 U9949 ( .IN1(n8873), .IN2(n8874), .Q(n8178) );
  XOR2X1 U9950 ( .IN1(n9632), .IN2(n4601), .Q(n8874) );
  XOR2X1 U9951 ( .IN1(WX3289), .IN2(n4325), .Q(n8873) );
  NOR2X0 U9952 ( .IN1(n6142), .IN2(n4724), .QN(n8871) );
  XOR2X1 U9953 ( .IN1(n8875), .IN2(n8876), .Q(n6142) );
  XOR2X1 U9954 ( .IN1(n9631), .IN2(n4627), .Q(n8876) );
  XOR2X1 U9955 ( .IN1(WX1996), .IN2(n4354), .Q(n8875) );
  NOR2X0 U9956 ( .IN1(n8877), .IN2(n8878), .QN(n8869) );
  NOR2X0 U9957 ( .IN1(DFF_354_n1), .IN2(n4758), .QN(n8878) );
  NOR2X0 U9958 ( .IN1(n4798), .IN2(n5637), .QN(n8877) );
  NAND2X0 U9959 ( .IN1(n5299), .IN2(n8672), .QN(n5637) );
  NAND2X0 U9960 ( .IN1(n8879), .IN2(n8880), .QN(WX1993) );
  NOR2X0 U9961 ( .IN1(n8881), .IN2(n8882), .QN(n8880) );
  NOR2X0 U9962 ( .IN1(n8187), .IN2(n4784), .QN(n8882) );
  XOR2X1 U9963 ( .IN1(n8883), .IN2(n8884), .Q(n8187) );
  XOR2X1 U9964 ( .IN1(n9634), .IN2(n4600), .Q(n8884) );
  XOR2X1 U9965 ( .IN1(WX3287), .IN2(n4327), .Q(n8883) );
  NOR2X0 U9966 ( .IN1(n8885), .IN2(n4724), .QN(n8881) );
  INVX0 U9967 ( .INP(n6162), .ZN(n8885) );
  XNOR2X1 U9968 ( .IN1(n8886), .IN2(n8887), .Q(n6162) );
  XOR2X1 U9969 ( .IN1(n9633), .IN2(n4626), .Q(n8887) );
  XOR2X1 U9970 ( .IN1(WX1994), .IN2(n4356), .Q(n8886) );
  NOR2X0 U9971 ( .IN1(n8888), .IN2(n8889), .QN(n8879) );
  NOR2X0 U9972 ( .IN1(DFF_355_n1), .IN2(n4758), .QN(n8889) );
  NOR2X0 U9973 ( .IN1(n4798), .IN2(n5638), .QN(n8888) );
  NAND2X0 U9974 ( .IN1(n5299), .IN2(n8673), .QN(n5638) );
  NAND2X0 U9975 ( .IN1(n8890), .IN2(n8891), .QN(WX1991) );
  NOR2X0 U9976 ( .IN1(n8892), .IN2(n8893), .QN(n8891) );
  NOR2X0 U9977 ( .IN1(n8196), .IN2(n4781), .QN(n8893) );
  XOR2X1 U9978 ( .IN1(n8894), .IN2(n8895), .Q(n8196) );
  XOR2X1 U9979 ( .IN1(n9636), .IN2(n4405), .Q(n8895) );
  XOR2X1 U9980 ( .IN1(WX3285), .IN2(n4329), .Q(n8894) );
  NOR2X0 U9981 ( .IN1(n4731), .IN2(n6182), .QN(n8892) );
  XNOR2X1 U9982 ( .IN1(n8896), .IN2(n8897), .Q(n6182) );
  XOR2X1 U9983 ( .IN1(test_so14), .IN2(n9635), .Q(n8897) );
  XOR2X1 U9984 ( .IN1(WX2120), .IN2(n4408), .Q(n8896) );
  NOR2X0 U9985 ( .IN1(n8898), .IN2(n8899), .QN(n8890) );
  NOR2X0 U9986 ( .IN1(DFF_356_n1), .IN2(n4758), .QN(n8899) );
  NOR2X0 U9987 ( .IN1(n4798), .IN2(n5639), .QN(n8898) );
  NAND2X0 U9988 ( .IN1(n5299), .IN2(n8674), .QN(n5639) );
  NAND2X0 U9989 ( .IN1(n8900), .IN2(n8901), .QN(WX1989) );
  NOR2X0 U9990 ( .IN1(n8902), .IN2(n8903), .QN(n8901) );
  NOR2X0 U9991 ( .IN1(n8205), .IN2(n4782), .QN(n8903) );
  XOR2X1 U9992 ( .IN1(n8904), .IN2(n8905), .Q(n8205) );
  XOR2X1 U9993 ( .IN1(n9638), .IN2(n4599), .Q(n8905) );
  XOR2X1 U9994 ( .IN1(WX3283), .IN2(n4331), .Q(n8904) );
  NOR2X0 U9995 ( .IN1(n8906), .IN2(n4724), .QN(n8902) );
  INVX0 U9996 ( .INP(n6196), .ZN(n8906) );
  XNOR2X1 U9997 ( .IN1(n8907), .IN2(n8908), .Q(n6196) );
  XOR2X1 U9998 ( .IN1(n9637), .IN2(n4625), .Q(n8908) );
  XOR2X1 U9999 ( .IN1(WX1990), .IN2(n4359), .Q(n8907) );
  NOR2X0 U10000 ( .IN1(n8909), .IN2(n8910), .QN(n8900) );
  NOR2X0 U10001 ( .IN1(DFF_357_n1), .IN2(n4757), .QN(n8910) );
  NOR2X0 U10002 ( .IN1(n4798), .IN2(n5640), .QN(n8909) );
  NAND2X0 U10003 ( .IN1(n5298), .IN2(n8675), .QN(n5640) );
  NAND2X0 U10004 ( .IN1(n8911), .IN2(n8912), .QN(WX1987) );
  NOR2X0 U10005 ( .IN1(n8913), .IN2(n8914), .QN(n8912) );
  NOR2X0 U10006 ( .IN1(n4785), .IN2(n8214), .QN(n8914) );
  XNOR2X1 U10007 ( .IN1(n8915), .IN2(n8916), .Q(n8214) );
  XOR2X1 U10008 ( .IN1(test_so30), .IN2(n9640), .Q(n8916) );
  XOR2X1 U10009 ( .IN1(WX3281), .IN2(n4333), .Q(n8915) );
  NOR2X0 U10010 ( .IN1(n6204), .IN2(n4724), .QN(n8913) );
  XOR2X1 U10011 ( .IN1(n8917), .IN2(n8918), .Q(n6204) );
  XOR2X1 U10012 ( .IN1(n9639), .IN2(n4624), .Q(n8918) );
  XOR2X1 U10013 ( .IN1(WX1988), .IN2(n4361), .Q(n8917) );
  NOR2X0 U10014 ( .IN1(n8919), .IN2(n8920), .QN(n8911) );
  NOR2X0 U10015 ( .IN1(DFF_358_n1), .IN2(n4757), .QN(n8920) );
  NOR2X0 U10016 ( .IN1(n4798), .IN2(n5650), .QN(n8919) );
  NAND2X0 U10017 ( .IN1(n5298), .IN2(n8676), .QN(n5650) );
  NAND2X0 U10018 ( .IN1(n8921), .IN2(n8922), .QN(WX1985) );
  NOR2X0 U10019 ( .IN1(n8923), .IN2(n8924), .QN(n8922) );
  NOR2X0 U10020 ( .IN1(n8223), .IN2(n4784), .QN(n8924) );
  XOR2X1 U10021 ( .IN1(n8925), .IN2(n8926), .Q(n8223) );
  XOR2X1 U10022 ( .IN1(n9642), .IN2(n4598), .Q(n8926) );
  XOR2X1 U10023 ( .IN1(WX3279), .IN2(n4335), .Q(n8925) );
  NOR2X0 U10024 ( .IN1(n8927), .IN2(n4724), .QN(n8923) );
  INVX0 U10025 ( .INP(n6220), .ZN(n8927) );
  XNOR2X1 U10026 ( .IN1(n8928), .IN2(n8929), .Q(n6220) );
  XOR2X1 U10027 ( .IN1(n9641), .IN2(n4623), .Q(n8929) );
  XOR2X1 U10028 ( .IN1(WX1986), .IN2(n4363), .Q(n8928) );
  NOR2X0 U10029 ( .IN1(n8930), .IN2(n8931), .QN(n8921) );
  NOR2X0 U10030 ( .IN1(n4764), .IN2(n4703), .QN(n8931) );
  NOR2X0 U10031 ( .IN1(n4798), .IN2(n5651), .QN(n8930) );
  NAND2X0 U10032 ( .IN1(n5298), .IN2(n8677), .QN(n5651) );
  NAND2X0 U10033 ( .IN1(n8932), .IN2(n8933), .QN(WX1983) );
  NOR2X0 U10034 ( .IN1(n8934), .IN2(n8935), .QN(n8933) );
  NOR2X0 U10035 ( .IN1(n4785), .IN2(n8232), .QN(n8935) );
  XNOR2X1 U10036 ( .IN1(n8936), .IN2(n8937), .Q(n8232) );
  XOR2X1 U10037 ( .IN1(test_so28), .IN2(n9644), .Q(n8937) );
  XOR2X1 U10038 ( .IN1(WX3277), .IN2(n4597), .Q(n8936) );
  NOR2X0 U10039 ( .IN1(n8938), .IN2(n6016), .QN(n8934) );
  INVX0 U10040 ( .INP(n6239), .ZN(n8938) );
  XNOR2X1 U10041 ( .IN1(n8939), .IN2(n8940), .Q(n6239) );
  XOR2X1 U10042 ( .IN1(n9643), .IN2(n4622), .Q(n8940) );
  XOR2X1 U10043 ( .IN1(WX1984), .IN2(n4365), .Q(n8939) );
  NOR2X0 U10044 ( .IN1(n8941), .IN2(n8942), .QN(n8932) );
  NOR2X0 U10045 ( .IN1(DFF_360_n1), .IN2(n4757), .QN(n8942) );
  NOR2X0 U10046 ( .IN1(n4798), .IN2(n5652), .QN(n8941) );
  NAND2X0 U10047 ( .IN1(test_so12), .IN2(n5323), .QN(n5652) );
  NAND2X0 U10048 ( .IN1(n8943), .IN2(n8944), .QN(WX1981) );
  NOR2X0 U10049 ( .IN1(n8945), .IN2(n8946), .QN(n8944) );
  NOR2X0 U10050 ( .IN1(n8241), .IN2(n4783), .QN(n8946) );
  XOR2X1 U10051 ( .IN1(n8947), .IN2(n8948), .Q(n8241) );
  XOR2X1 U10052 ( .IN1(n9646), .IN2(n4596), .Q(n8948) );
  XOR2X1 U10053 ( .IN1(WX3275), .IN2(n4338), .Q(n8947) );
  NOR2X0 U10054 ( .IN1(n8949), .IN2(n6016), .QN(n8945) );
  INVX0 U10055 ( .INP(n6267), .ZN(n8949) );
  XNOR2X1 U10056 ( .IN1(n8950), .IN2(n8951), .Q(n6267) );
  XOR2X1 U10057 ( .IN1(n9645), .IN2(n4621), .Q(n8951) );
  XOR2X1 U10058 ( .IN1(WX1982), .IN2(n4367), .Q(n8950) );
  NOR2X0 U10059 ( .IN1(n8952), .IN2(n8953), .QN(n8943) );
  NOR2X0 U10060 ( .IN1(DFF_361_n1), .IN2(n4757), .QN(n8953) );
  NOR2X0 U10061 ( .IN1(n4798), .IN2(n5653), .QN(n8952) );
  NAND2X0 U10062 ( .IN1(n5298), .IN2(n8680), .QN(n5653) );
  NAND2X0 U10063 ( .IN1(n8954), .IN2(n8955), .QN(WX1979) );
  NOR2X0 U10064 ( .IN1(n8956), .IN2(n8957), .QN(n8955) );
  NOR2X0 U10065 ( .IN1(n8291), .IN2(n4783), .QN(n8957) );
  XOR2X1 U10066 ( .IN1(n8958), .IN2(n8959), .Q(n8291) );
  XOR2X1 U10067 ( .IN1(n9648), .IN2(n4595), .Q(n8959) );
  XOR2X1 U10068 ( .IN1(WX3273), .IN2(n4340), .Q(n8958) );
  NOR2X0 U10069 ( .IN1(n4731), .IN2(n7407), .QN(n8956) );
  XNOR2X1 U10070 ( .IN1(n8960), .IN2(n8961), .Q(n7407) );
  XOR2X1 U10071 ( .IN1(test_so19), .IN2(n9647), .Q(n8961) );
  XOR2X1 U10072 ( .IN1(WX1980), .IN2(n4369), .Q(n8960) );
  NOR2X0 U10073 ( .IN1(n8962), .IN2(n8963), .QN(n8954) );
  NOR2X0 U10074 ( .IN1(DFF_362_n1), .IN2(n4757), .QN(n8963) );
  NOR2X0 U10075 ( .IN1(n4798), .IN2(n5654), .QN(n8962) );
  NAND2X0 U10076 ( .IN1(n5298), .IN2(n8681), .QN(n5654) );
  NAND2X0 U10077 ( .IN1(n8964), .IN2(n8965), .QN(WX1977) );
  NOR2X0 U10078 ( .IN1(n8966), .IN2(n8967), .QN(n8965) );
  NOR2X0 U10079 ( .IN1(n8303), .IN2(n4783), .QN(n8967) );
  XOR2X1 U10080 ( .IN1(n8968), .IN2(n8969), .Q(n8303) );
  XOR2X1 U10081 ( .IN1(n9650), .IN2(n4404), .Q(n8969) );
  XOR2X1 U10082 ( .IN1(WX3271), .IN2(n4342), .Q(n8968) );
  NOR2X0 U10083 ( .IN1(n8970), .IN2(n6016), .QN(n8966) );
  INVX0 U10084 ( .INP(n6281), .ZN(n8970) );
  XNOR2X1 U10085 ( .IN1(n8971), .IN2(n8972), .Q(n6281) );
  XOR2X1 U10086 ( .IN1(n9649), .IN2(n4407), .Q(n8972) );
  XOR2X1 U10087 ( .IN1(WX1978), .IN2(n4371), .Q(n8971) );
  NOR2X0 U10088 ( .IN1(n8973), .IN2(n8974), .QN(n8964) );
  NOR2X0 U10089 ( .IN1(DFF_363_n1), .IN2(n4757), .QN(n8974) );
  NOR2X0 U10090 ( .IN1(n4797), .IN2(n5655), .QN(n8973) );
  NAND2X0 U10091 ( .IN1(n5298), .IN2(n8682), .QN(n5655) );
  NAND2X0 U10092 ( .IN1(n8975), .IN2(n8976), .QN(WX1975) );
  NOR2X0 U10093 ( .IN1(n8977), .IN2(n8978), .QN(n8976) );
  NOR2X0 U10094 ( .IN1(n4785), .IN2(n8356), .QN(n8978) );
  XNOR2X1 U10095 ( .IN1(n8979), .IN2(n8980), .Q(n8356) );
  XOR2X1 U10096 ( .IN1(test_so26), .IN2(n9652), .Q(n8980) );
  XOR2X1 U10097 ( .IN1(WX3269), .IN2(n4594), .Q(n8979) );
  NOR2X0 U10098 ( .IN1(n8981), .IN2(n6016), .QN(n8977) );
  INVX0 U10099 ( .INP(n6290), .ZN(n8981) );
  XNOR2X1 U10100 ( .IN1(n8982), .IN2(n8983), .Q(n6290) );
  XOR2X1 U10101 ( .IN1(n9651), .IN2(n4620), .Q(n8983) );
  XOR2X1 U10102 ( .IN1(WX1976), .IN2(n4373), .Q(n8982) );
  NOR2X0 U10103 ( .IN1(n8984), .IN2(n8985), .QN(n8975) );
  NOR2X0 U10104 ( .IN1(DFF_364_n1), .IN2(n4757), .QN(n8985) );
  NOR2X0 U10105 ( .IN1(n4797), .IN2(n5656), .QN(n8984) );
  NAND2X0 U10106 ( .IN1(n5297), .IN2(n8683), .QN(n5656) );
  NAND2X0 U10107 ( .IN1(n8986), .IN2(n8987), .QN(WX1973) );
  NOR2X0 U10108 ( .IN1(n8988), .IN2(n8989), .QN(n8987) );
  NOR2X0 U10109 ( .IN1(n8397), .IN2(n4782), .QN(n8989) );
  XOR2X1 U10110 ( .IN1(n8990), .IN2(n8991), .Q(n8397) );
  XOR2X1 U10111 ( .IN1(n9654), .IN2(n4593), .Q(n8991) );
  XOR2X1 U10112 ( .IN1(WX3267), .IN2(n4345), .Q(n8990) );
  NOR2X0 U10113 ( .IN1(n8992), .IN2(n6016), .QN(n8988) );
  INVX0 U10114 ( .INP(n6305), .ZN(n8992) );
  XNOR2X1 U10115 ( .IN1(n8993), .IN2(n8994), .Q(n6305) );
  XOR2X1 U10116 ( .IN1(n9653), .IN2(n4619), .Q(n8994) );
  XOR2X1 U10117 ( .IN1(WX1974), .IN2(n4375), .Q(n8993) );
  NOR2X0 U10118 ( .IN1(n8995), .IN2(n8996), .QN(n8986) );
  NOR2X0 U10119 ( .IN1(DFF_365_n1), .IN2(n4757), .QN(n8996) );
  NOR2X0 U10120 ( .IN1(n4797), .IN2(n5657), .QN(n8995) );
  NAND2X0 U10121 ( .IN1(n5297), .IN2(n8684), .QN(n5657) );
  NAND2X0 U10122 ( .IN1(n8997), .IN2(n8998), .QN(WX1971) );
  NOR2X0 U10123 ( .IN1(n8999), .IN2(n9000), .QN(n8998) );
  NOR2X0 U10124 ( .IN1(n8419), .IN2(n4778), .QN(n9000) );
  XOR2X1 U10125 ( .IN1(n9001), .IN2(n9002), .Q(n8419) );
  XOR2X1 U10126 ( .IN1(n9656), .IN2(n4592), .Q(n9002) );
  XOR2X1 U10127 ( .IN1(WX3265), .IN2(n4347), .Q(n9001) );
  NOR2X0 U10128 ( .IN1(n4731), .IN2(n6325), .QN(n8999) );
  XNOR2X1 U10129 ( .IN1(n9003), .IN2(n9004), .Q(n6325) );
  XOR2X1 U10130 ( .IN1(test_so17), .IN2(n9655), .Q(n9004) );
  XOR2X1 U10131 ( .IN1(WX1972), .IN2(n4618), .Q(n9003) );
  NOR2X0 U10132 ( .IN1(n9005), .IN2(n9006), .QN(n8997) );
  NOR2X0 U10133 ( .IN1(DFF_366_n1), .IN2(n4757), .QN(n9006) );
  NOR2X0 U10134 ( .IN1(n4797), .IN2(n5658), .QN(n9005) );
  NAND2X0 U10135 ( .IN1(n5297), .IN2(n8685), .QN(n5658) );
  NAND2X0 U10136 ( .IN1(n9007), .IN2(n9008), .QN(WX1969) );
  NOR2X0 U10137 ( .IN1(n9009), .IN2(n9010), .QN(n9008) );
  NOR2X0 U10138 ( .IN1(n8472), .IN2(n4781), .QN(n9010) );
  XOR2X1 U10139 ( .IN1(n9011), .IN2(n9012), .Q(n8472) );
  XOR2X1 U10140 ( .IN1(n9658), .IN2(n4591), .Q(n9012) );
  XOR2X1 U10141 ( .IN1(WX3263), .IN2(n4349), .Q(n9011) );
  NOR2X0 U10142 ( .IN1(n9013), .IN2(n6016), .QN(n9009) );
  INVX0 U10143 ( .INP(n6343), .ZN(n9013) );
  XNOR2X1 U10144 ( .IN1(n9014), .IN2(n9015), .Q(n6343) );
  XOR2X1 U10145 ( .IN1(n9657), .IN2(n4617), .Q(n9015) );
  XOR2X1 U10146 ( .IN1(WX1970), .IN2(n4378), .Q(n9014) );
  NOR2X0 U10147 ( .IN1(n9016), .IN2(n9017), .QN(n9007) );
  NOR2X0 U10148 ( .IN1(DFF_367_n1), .IN2(n4757), .QN(n9017) );
  NOR2X0 U10149 ( .IN1(n4797), .IN2(n5659), .QN(n9016) );
  NAND2X0 U10150 ( .IN1(n5297), .IN2(n8686), .QN(n5659) );
  NAND2X0 U10151 ( .IN1(n9018), .IN2(n9019), .QN(WX1967) );
  NOR2X0 U10152 ( .IN1(n9020), .IN2(n9021), .QN(n9019) );
  NOR2X0 U10153 ( .IN1(n4784), .IN2(n8503), .QN(n9021) );
  XNOR2X1 U10154 ( .IN1(n9022), .IN2(n9023), .Q(n8503) );
  XOR2X1 U10155 ( .IN1(n4118), .IN2(n5255), .Q(n9023) );
  XOR2X1 U10156 ( .IN1(n9024), .IN2(n4403), .Q(n9022) );
  XOR2X1 U10157 ( .IN1(WX3325), .IN2(test_so24), .Q(n9024) );
  NOR2X0 U10158 ( .IN1(n7415), .IN2(n4726), .QN(n9020) );
  XOR2X1 U10159 ( .IN1(n9025), .IN2(n9026), .Q(n7415) );
  XOR2X1 U10160 ( .IN1(n4131), .IN2(n5255), .Q(n9026) );
  XOR2X1 U10161 ( .IN1(n9027), .IN2(n4406), .Q(n9025) );
  XOR2X1 U10162 ( .IN1(WX2096), .IN2(n9659), .Q(n9027) );
  NOR2X0 U10163 ( .IN1(n9028), .IN2(n9029), .QN(n9018) );
  NOR2X0 U10164 ( .IN1(DFF_368_n1), .IN2(n4757), .QN(n9029) );
  NOR2X0 U10165 ( .IN1(n4797), .IN2(n5669), .QN(n9028) );
  NAND2X0 U10166 ( .IN1(n5297), .IN2(n8687), .QN(n5669) );
  NAND2X0 U10167 ( .IN1(n9030), .IN2(n9031), .QN(WX1965) );
  NOR2X0 U10168 ( .IN1(n9032), .IN2(n9033), .QN(n9031) );
  NOR2X0 U10169 ( .IN1(n8535), .IN2(n4780), .QN(n9033) );
  XOR2X1 U10170 ( .IN1(n9034), .IN2(n9035), .Q(n8535) );
  XOR2X1 U10171 ( .IN1(n4119), .IN2(n5255), .Q(n9035) );
  XOR2X1 U10172 ( .IN1(n9036), .IN2(n4590), .Q(n9034) );
  XOR2X1 U10173 ( .IN1(WX3387), .IN2(n9661), .Q(n9036) );
  NOR2X0 U10174 ( .IN1(n9037), .IN2(n6016), .QN(n9032) );
  INVX0 U10175 ( .INP(n6360), .ZN(n9037) );
  XNOR2X1 U10176 ( .IN1(n9038), .IN2(n9039), .Q(n6360) );
  XOR2X1 U10177 ( .IN1(n4132), .IN2(n5255), .Q(n9039) );
  XOR2X1 U10178 ( .IN1(n9040), .IN2(n4616), .Q(n9038) );
  XOR2X1 U10179 ( .IN1(WX2094), .IN2(n9660), .Q(n9040) );
  NOR2X0 U10180 ( .IN1(n9041), .IN2(n9042), .QN(n9030) );
  NOR2X0 U10181 ( .IN1(DFF_369_n1), .IN2(n4757), .QN(n9042) );
  NOR2X0 U10182 ( .IN1(n4797), .IN2(n5670), .QN(n9041) );
  NAND2X0 U10183 ( .IN1(n5297), .IN2(n8688), .QN(n5670) );
  NAND2X0 U10184 ( .IN1(n9043), .IN2(n9044), .QN(WX1963) );
  NOR2X0 U10185 ( .IN1(n9045), .IN2(n9046), .QN(n9044) );
  NOR2X0 U10186 ( .IN1(n8589), .IN2(n4780), .QN(n9046) );
  XOR2X1 U10187 ( .IN1(n9047), .IN2(n9048), .Q(n8589) );
  XOR2X1 U10188 ( .IN1(n4120), .IN2(n5255), .Q(n9048) );
  XOR2X1 U10189 ( .IN1(n9049), .IN2(n4589), .Q(n9047) );
  XOR2X1 U10190 ( .IN1(WX3385), .IN2(n9665), .Q(n9049) );
  NOR2X0 U10191 ( .IN1(n4732), .IN2(n6370), .QN(n9045) );
  XNOR2X1 U10192 ( .IN1(n9050), .IN2(n9051), .Q(n6370) );
  XOR2X1 U10193 ( .IN1(n4615), .IN2(n5255), .Q(n9051) );
  XOR2X1 U10194 ( .IN1(n9052), .IN2(n9664), .Q(n9050) );
  XOR2X1 U10195 ( .IN1(n9663), .IN2(n9662), .Q(n9052) );
  NOR2X0 U10196 ( .IN1(n9053), .IN2(n9054), .QN(n9043) );
  NOR2X0 U10197 ( .IN1(DFF_370_n1), .IN2(n4756), .QN(n9054) );
  NOR2X0 U10198 ( .IN1(n4797), .IN2(n5671), .QN(n9053) );
  NAND2X0 U10199 ( .IN1(n5296), .IN2(n8689), .QN(n5671) );
  NAND2X0 U10200 ( .IN1(n9055), .IN2(n9056), .QN(WX1961) );
  NOR2X0 U10201 ( .IN1(n9057), .IN2(n9058), .QN(n9056) );
  NOR2X0 U10202 ( .IN1(n8633), .IN2(n4780), .QN(n9058) );
  XOR2X1 U10203 ( .IN1(n9059), .IN2(n9060), .Q(n8633) );
  XOR2X1 U10204 ( .IN1(n4121), .IN2(n5255), .Q(n9060) );
  XOR2X1 U10205 ( .IN1(n9061), .IN2(n4588), .Q(n9059) );
  XOR2X1 U10206 ( .IN1(WX3383), .IN2(n9667), .Q(n9061) );
  NOR2X0 U10207 ( .IN1(n9062), .IN2(n6016), .QN(n9057) );
  INVX0 U10208 ( .INP(n6379), .ZN(n9062) );
  XNOR2X1 U10209 ( .IN1(n9063), .IN2(n9064), .Q(n6379) );
  XOR2X1 U10210 ( .IN1(n4133), .IN2(n5255), .Q(n9064) );
  XOR2X1 U10211 ( .IN1(n9065), .IN2(n4614), .Q(n9063) );
  XOR2X1 U10212 ( .IN1(WX2090), .IN2(n9666), .Q(n9065) );
  NOR2X0 U10213 ( .IN1(n9066), .IN2(n9067), .QN(n9055) );
  NOR2X0 U10214 ( .IN1(DFF_371_n1), .IN2(n4756), .QN(n9067) );
  NOR2X0 U10215 ( .IN1(n4797), .IN2(n5672), .QN(n9066) );
  NAND2X0 U10216 ( .IN1(n5296), .IN2(n8690), .QN(n5672) );
  NAND2X0 U10217 ( .IN1(n9068), .IN2(n9069), .QN(WX1959) );
  NOR2X0 U10218 ( .IN1(n9070), .IN2(n9071), .QN(n9069) );
  NOR2X0 U10219 ( .IN1(n8659), .IN2(n4780), .QN(n9071) );
  XOR2X1 U10220 ( .IN1(n9072), .IN2(n9073), .Q(n8659) );
  XOR2X1 U10221 ( .IN1(n4122), .IN2(n5255), .Q(n9073) );
  XOR2X1 U10222 ( .IN1(n9074), .IN2(n4587), .Q(n9072) );
  XOR2X1 U10223 ( .IN1(WX3381), .IN2(n9669), .Q(n9074) );
  NOR2X0 U10224 ( .IN1(n7424), .IN2(n6016), .QN(n9070) );
  XOR2X1 U10225 ( .IN1(n9075), .IN2(n9076), .Q(n7424) );
  XOR2X1 U10226 ( .IN1(n4134), .IN2(n5255), .Q(n9076) );
  XOR2X1 U10227 ( .IN1(n9077), .IN2(n4613), .Q(n9075) );
  XOR2X1 U10228 ( .IN1(WX2088), .IN2(n9668), .Q(n9077) );
  NOR2X0 U10229 ( .IN1(n9078), .IN2(n9079), .QN(n9068) );
  NOR2X0 U10230 ( .IN1(DFF_372_n1), .IN2(n4756), .QN(n9079) );
  NOR2X0 U10231 ( .IN1(n4797), .IN2(n5673), .QN(n9078) );
  NAND2X0 U10232 ( .IN1(n5296), .IN2(n8691), .QN(n5673) );
  NAND2X0 U10233 ( .IN1(n9080), .IN2(n9081), .QN(WX1957) );
  NOR2X0 U10234 ( .IN1(n9082), .IN2(n9083), .QN(n9081) );
  NOR2X0 U10235 ( .IN1(n8707), .IN2(n4780), .QN(n9083) );
  XOR2X1 U10236 ( .IN1(n9084), .IN2(n9085), .Q(n8707) );
  XOR2X1 U10237 ( .IN1(n4123), .IN2(n5255), .Q(n9085) );
  XOR2X1 U10238 ( .IN1(n9086), .IN2(n4586), .Q(n9084) );
  XOR2X1 U10239 ( .IN1(WX3379), .IN2(n9671), .Q(n9086) );
  NOR2X0 U10240 ( .IN1(n9087), .IN2(n6016), .QN(n9082) );
  INVX0 U10241 ( .INP(n6388), .ZN(n9087) );
  XNOR2X1 U10242 ( .IN1(n9088), .IN2(n9089), .Q(n6388) );
  XOR2X1 U10243 ( .IN1(n4135), .IN2(n5256), .Q(n9089) );
  XOR2X1 U10244 ( .IN1(n9090), .IN2(n4612), .Q(n9088) );
  XOR2X1 U10245 ( .IN1(WX2086), .IN2(n9670), .Q(n9090) );
  NOR2X0 U10246 ( .IN1(n9091), .IN2(n9092), .QN(n9080) );
  NOR2X0 U10247 ( .IN1(DFF_373_n1), .IN2(n4756), .QN(n9092) );
  NOR2X0 U10248 ( .IN1(n4797), .IN2(n5674), .QN(n9091) );
  NAND2X0 U10249 ( .IN1(n5296), .IN2(n8692), .QN(n5674) );
  NAND2X0 U10250 ( .IN1(n9093), .IN2(n9094), .QN(WX1955) );
  NOR2X0 U10251 ( .IN1(n9095), .IN2(n9096), .QN(n9094) );
  NOR2X0 U10252 ( .IN1(n8717), .IN2(n4780), .QN(n9096) );
  XOR2X1 U10253 ( .IN1(n9097), .IN2(n9098), .Q(n8717) );
  XOR2X1 U10254 ( .IN1(n4124), .IN2(n5256), .Q(n9098) );
  XOR2X1 U10255 ( .IN1(n9099), .IN2(n4585), .Q(n9097) );
  XOR2X1 U10256 ( .IN1(WX3377), .IN2(n9672), .Q(n9099) );
  NOR2X0 U10257 ( .IN1(n5634), .IN2(n4732), .QN(n9095) );
  XNOR2X1 U10258 ( .IN1(n9100), .IN2(n9101), .Q(n5634) );
  XOR2X1 U10259 ( .IN1(n4136), .IN2(n5256), .Q(n9101) );
  XOR2X1 U10260 ( .IN1(n9102), .IN2(n4611), .Q(n9100) );
  XOR2X1 U10261 ( .IN1(WX2020), .IN2(test_so13), .Q(n9102) );
  NOR2X0 U10262 ( .IN1(n9103), .IN2(n9104), .QN(n9093) );
  NOR2X0 U10263 ( .IN1(DFF_374_n1), .IN2(n4756), .QN(n9104) );
  NOR2X0 U10264 ( .IN1(n4797), .IN2(n5675), .QN(n9103) );
  NAND2X0 U10265 ( .IN1(n5296), .IN2(n8693), .QN(n5675) );
  NAND2X0 U10266 ( .IN1(n9105), .IN2(n9106), .QN(WX1953) );
  NOR2X0 U10267 ( .IN1(n9107), .IN2(n9108), .QN(n9106) );
  NOR2X0 U10268 ( .IN1(n4785), .IN2(n8727), .QN(n9108) );
  XNOR2X1 U10269 ( .IN1(n9109), .IN2(n9110), .Q(n8727) );
  XOR2X1 U10270 ( .IN1(n4125), .IN2(n5256), .Q(n9110) );
  XOR2X1 U10271 ( .IN1(WX3311), .IN2(n9111), .Q(n9109) );
  XOR2X1 U10272 ( .IN1(test_so29), .IN2(n9674), .Q(n9111) );
  NOR2X0 U10273 ( .IN1(n9112), .IN2(n4723), .QN(n9107) );
  INVX0 U10274 ( .INP(n5649), .ZN(n9112) );
  XNOR2X1 U10275 ( .IN1(n9113), .IN2(n9114), .Q(n5649) );
  XOR2X1 U10276 ( .IN1(n4137), .IN2(n5256), .Q(n9114) );
  XOR2X1 U10277 ( .IN1(n9115), .IN2(n4610), .Q(n9113) );
  XOR2X1 U10278 ( .IN1(WX2082), .IN2(n9673), .Q(n9115) );
  NOR2X0 U10279 ( .IN1(n9116), .IN2(n9117), .QN(n9105) );
  NOR2X0 U10280 ( .IN1(DFF_375_n1), .IN2(n4756), .QN(n9117) );
  NOR2X0 U10281 ( .IN1(n4797), .IN2(n5676), .QN(n9116) );
  NAND2X0 U10282 ( .IN1(n5296), .IN2(n8694), .QN(n5676) );
  NAND2X0 U10283 ( .IN1(n9118), .IN2(n9119), .QN(WX1951) );
  NOR2X0 U10284 ( .IN1(n9120), .IN2(n9121), .QN(n9119) );
  NOR2X0 U10285 ( .IN1(n8737), .IN2(n4780), .QN(n9121) );
  XOR2X1 U10286 ( .IN1(n9122), .IN2(n9123), .Q(n8737) );
  XOR2X1 U10287 ( .IN1(n4126), .IN2(n5256), .Q(n9123) );
  XOR2X1 U10288 ( .IN1(n9124), .IN2(n4584), .Q(n9122) );
  XOR2X1 U10289 ( .IN1(WX3373), .IN2(n9676), .Q(n9124) );
  NOR2X0 U10290 ( .IN1(n7433), .IN2(n4723), .QN(n9120) );
  XOR2X1 U10291 ( .IN1(n9125), .IN2(n9126), .Q(n7433) );
  XOR2X1 U10292 ( .IN1(n4138), .IN2(n5256), .Q(n9126) );
  XOR2X1 U10293 ( .IN1(n9127), .IN2(n4609), .Q(n9125) );
  XOR2X1 U10294 ( .IN1(WX2080), .IN2(n9675), .Q(n9127) );
  NOR2X0 U10295 ( .IN1(n9128), .IN2(n9129), .QN(n9118) );
  NOR2X0 U10296 ( .IN1(DFF_376_n1), .IN2(n4756), .QN(n9129) );
  NOR2X0 U10297 ( .IN1(n4796), .IN2(n5677), .QN(n9128) );
  NAND2X0 U10298 ( .IN1(n5295), .IN2(n8695), .QN(n5677) );
  NAND2X0 U10299 ( .IN1(n9130), .IN2(n9131), .QN(WX1949) );
  NOR2X0 U10300 ( .IN1(n9132), .IN2(n9133), .QN(n9131) );
  NOR2X0 U10301 ( .IN1(n8747), .IN2(n4779), .QN(n9133) );
  XOR2X1 U10302 ( .IN1(n9134), .IN2(n9135), .Q(n8747) );
  XOR2X1 U10303 ( .IN1(n4127), .IN2(n5256), .Q(n9135) );
  XOR2X1 U10304 ( .IN1(n9136), .IN2(n4583), .Q(n9134) );
  XOR2X1 U10305 ( .IN1(WX3371), .IN2(n9678), .Q(n9136) );
  NOR2X0 U10306 ( .IN1(n9137), .IN2(n4723), .QN(n9132) );
  INVX0 U10307 ( .INP(n5668), .ZN(n9137) );
  XNOR2X1 U10308 ( .IN1(n9138), .IN2(n9139), .Q(n5668) );
  XOR2X1 U10309 ( .IN1(n4139), .IN2(n5256), .Q(n9139) );
  XOR2X1 U10310 ( .IN1(n9140), .IN2(n4608), .Q(n9138) );
  XOR2X1 U10311 ( .IN1(WX2078), .IN2(n9677), .Q(n9140) );
  NOR2X0 U10312 ( .IN1(n9141), .IN2(n9142), .QN(n9130) );
  NOR2X0 U10313 ( .IN1(n4765), .IN2(n4704), .QN(n9142) );
  NOR2X0 U10314 ( .IN1(n4796), .IN2(n5678), .QN(n9141) );
  NAND2X0 U10315 ( .IN1(n5295), .IN2(n8696), .QN(n5678) );
  NAND2X0 U10316 ( .IN1(n9143), .IN2(n9144), .QN(WX1947) );
  NOR2X0 U10317 ( .IN1(n9145), .IN2(n9146), .QN(n9144) );
  NOR2X0 U10318 ( .IN1(n4784), .IN2(n8757), .QN(n9146) );
  XNOR2X1 U10319 ( .IN1(n9147), .IN2(n9148), .Q(n8757) );
  XOR2X1 U10320 ( .IN1(n4582), .IN2(n5256), .Q(n9148) );
  XOR2X1 U10321 ( .IN1(n9149), .IN2(n9682), .Q(n9147) );
  XOR2X1 U10322 ( .IN1(n9681), .IN2(n9680), .Q(n9149) );
  NOR2X0 U10323 ( .IN1(n9150), .IN2(n4723), .QN(n9145) );
  INVX0 U10324 ( .INP(n5687), .ZN(n9150) );
  XNOR2X1 U10325 ( .IN1(n9151), .IN2(n9152), .Q(n5687) );
  XOR2X1 U10326 ( .IN1(n4140), .IN2(n5256), .Q(n9152) );
  XOR2X1 U10327 ( .IN1(n9153), .IN2(n4607), .Q(n9151) );
  XOR2X1 U10328 ( .IN1(WX2076), .IN2(n9679), .Q(n9153) );
  NOR2X0 U10329 ( .IN1(n9154), .IN2(n9155), .QN(n9143) );
  NOR2X0 U10330 ( .IN1(DFF_378_n1), .IN2(n4756), .QN(n9155) );
  NOR2X0 U10331 ( .IN1(n4796), .IN2(n5688), .QN(n9154) );
  NAND2X0 U10332 ( .IN1(test_so11), .IN2(n5324), .QN(n5688) );
  NAND2X0 U10333 ( .IN1(n9156), .IN2(n9157), .QN(WX1945) );
  NOR2X0 U10334 ( .IN1(n9158), .IN2(n9159), .QN(n9157) );
  NOR2X0 U10335 ( .IN1(n8767), .IN2(n4779), .QN(n9159) );
  XOR2X1 U10336 ( .IN1(n9160), .IN2(n9161), .Q(n8767) );
  XOR2X1 U10337 ( .IN1(n4128), .IN2(n5257), .Q(n9161) );
  XOR2X1 U10338 ( .IN1(n9162), .IN2(n4581), .Q(n9160) );
  XOR2X1 U10339 ( .IN1(WX3367), .IN2(n9684), .Q(n9162) );
  NOR2X0 U10340 ( .IN1(n9163), .IN2(n4723), .QN(n9158) );
  INVX0 U10341 ( .INP(n5701), .ZN(n9163) );
  XNOR2X1 U10342 ( .IN1(n9164), .IN2(n9165), .Q(n5701) );
  XOR2X1 U10343 ( .IN1(n4141), .IN2(n5257), .Q(n9165) );
  XOR2X1 U10344 ( .IN1(n9166), .IN2(n4606), .Q(n9164) );
  XOR2X1 U10345 ( .IN1(WX2074), .IN2(n9683), .Q(n9166) );
  NOR2X0 U10346 ( .IN1(n9167), .IN2(n9168), .QN(n9156) );
  NOR2X0 U10347 ( .IN1(DFF_379_n1), .IN2(n4756), .QN(n9168) );
  NOR2X0 U10348 ( .IN1(n4796), .IN2(n5689), .QN(n9167) );
  NAND2X0 U10349 ( .IN1(n5295), .IN2(n8699), .QN(n5689) );
  NAND2X0 U10350 ( .IN1(n9169), .IN2(n9170), .QN(WX1943) );
  NOR2X0 U10351 ( .IN1(n9171), .IN2(n9172), .QN(n9170) );
  NOR2X0 U10352 ( .IN1(n8777), .IN2(n4778), .QN(n9172) );
  XOR2X1 U10353 ( .IN1(n9173), .IN2(n9174), .Q(n8777) );
  XOR2X1 U10354 ( .IN1(n4129), .IN2(n5256), .Q(n9174) );
  XOR2X1 U10355 ( .IN1(n9175), .IN2(n4580), .Q(n9173) );
  XOR2X1 U10356 ( .IN1(WX3365), .IN2(n9686), .Q(n9175) );
  NOR2X0 U10357 ( .IN1(n4732), .IN2(n6020), .QN(n9171) );
  XNOR2X1 U10358 ( .IN1(n9176), .IN2(n9177), .Q(n6020) );
  XOR2X1 U10359 ( .IN1(n4142), .IN2(n5257), .Q(n9177) );
  XOR2X1 U10360 ( .IN1(WX2008), .IN2(n9178), .Q(n9176) );
  XOR2X1 U10361 ( .IN1(test_so18), .IN2(n9685), .Q(n9178) );
  NOR2X0 U10362 ( .IN1(n9179), .IN2(n9180), .QN(n9169) );
  NOR2X0 U10363 ( .IN1(DFF_380_n1), .IN2(n4756), .QN(n9180) );
  NOR2X0 U10364 ( .IN1(n4796), .IN2(n5690), .QN(n9179) );
  NAND2X0 U10365 ( .IN1(n5309), .IN2(n8700), .QN(n5690) );
  NAND2X0 U10366 ( .IN1(n9181), .IN2(n9182), .QN(WX1941) );
  NOR2X0 U10367 ( .IN1(n9183), .IN2(n9184), .QN(n9182) );
  NOR2X0 U10368 ( .IN1(n8787), .IN2(n4778), .QN(n9184) );
  XOR2X1 U10369 ( .IN1(n9185), .IN2(n9186), .Q(n8787) );
  XOR2X1 U10370 ( .IN1(n4130), .IN2(n5257), .Q(n9186) );
  XOR2X1 U10371 ( .IN1(n9187), .IN2(n4579), .Q(n9185) );
  XOR2X1 U10372 ( .IN1(WX3363), .IN2(n9688), .Q(n9187) );
  NOR2X0 U10373 ( .IN1(n9188), .IN2(n4723), .QN(n9183) );
  INVX0 U10374 ( .INP(n6094), .ZN(n9188) );
  XNOR2X1 U10375 ( .IN1(n9189), .IN2(n9190), .Q(n6094) );
  XOR2X1 U10376 ( .IN1(n4143), .IN2(n5257), .Q(n9190) );
  XOR2X1 U10377 ( .IN1(n9191), .IN2(n4605), .Q(n9189) );
  XOR2X1 U10378 ( .IN1(WX2070), .IN2(n9687), .Q(n9191) );
  NOR2X0 U10379 ( .IN1(n9192), .IN2(n9193), .QN(n9181) );
  NOR2X0 U10380 ( .IN1(DFF_381_n1), .IN2(n4756), .QN(n9193) );
  NOR2X0 U10381 ( .IN1(n4800), .IN2(n5691), .QN(n9192) );
  NAND2X0 U10382 ( .IN1(n5283), .IN2(n8701), .QN(n5691) );
  NAND2X0 U10383 ( .IN1(n9194), .IN2(n9195), .QN(WX1939) );
  NOR2X0 U10384 ( .IN1(n9196), .IN2(n9197), .QN(n9195) );
  NOR2X0 U10385 ( .IN1(n4785), .IN2(n8797), .QN(n9197) );
  XNOR2X1 U10386 ( .IN1(n9198), .IN2(n9199), .Q(n8797) );
  XOR2X1 U10387 ( .IN1(n4578), .IN2(n5257), .Q(n9199) );
  XOR2X1 U10388 ( .IN1(n9200), .IN2(n9692), .Q(n9198) );
  XOR2X1 U10389 ( .IN1(n9691), .IN2(n9690), .Q(n9200) );
  NOR2X0 U10390 ( .IN1(n9201), .IN2(n6016), .QN(n9196) );
  INVX0 U10391 ( .INP(n6248), .ZN(n9201) );
  XNOR2X1 U10392 ( .IN1(n9202), .IN2(n9203), .Q(n6248) );
  XOR2X1 U10393 ( .IN1(n4144), .IN2(n5257), .Q(n9203) );
  XOR2X1 U10394 ( .IN1(n9204), .IN2(n4604), .Q(n9202) );
  XOR2X1 U10395 ( .IN1(WX2068), .IN2(n9689), .Q(n9204) );
  NOR2X0 U10396 ( .IN1(n9205), .IN2(n9206), .QN(n9194) );
  NOR2X0 U10397 ( .IN1(DFF_382_n1), .IN2(n4760), .QN(n9206) );
  NOR2X0 U10398 ( .IN1(n6023), .IN2(n5692), .QN(n9205) );
  NAND2X0 U10399 ( .IN1(n5295), .IN2(n8702), .QN(n5692) );
  NAND2X0 U10400 ( .IN1(n5259), .IN2(TM0), .QN(n6023) );
  NAND2X0 U10401 ( .IN1(n9207), .IN2(n9208), .QN(WX1937) );
  NOR2X0 U10402 ( .IN1(n9209), .IN2(n9210), .QN(n9208) );
  NOR2X0 U10403 ( .IN1(n7473), .IN2(n4715), .QN(n9210) );
  NAND2X0 U10404 ( .IN1(n9211), .IN2(n5259), .QN(n6016) );
  NOR2X0 U10405 ( .IN1(TM0), .IN2(n5349), .QN(n9211) );
  XOR2X1 U10406 ( .IN1(n9212), .IN2(n9213), .Q(n7473) );
  XOR2X1 U10407 ( .IN1(n4038), .IN2(n5257), .Q(n9213) );
  XOR2X1 U10408 ( .IN1(n9214), .IN2(n4603), .Q(n9212) );
  XOR2X1 U10409 ( .IN1(WX2066), .IN2(n9694), .Q(n9214) );
  NOR2X0 U10410 ( .IN1(n8807), .IN2(n4770), .QN(n9209) );
  INVX0 U10411 ( .INP(n2153), .ZN(n6021) );
  XOR2X1 U10412 ( .IN1(n9215), .IN2(n9216), .Q(n8807) );
  XOR2X1 U10413 ( .IN1(n4037), .IN2(n5257), .Q(n9216) );
  XOR2X1 U10414 ( .IN1(n9217), .IN2(n4577), .Q(n9215) );
  XOR2X1 U10415 ( .IN1(WX3359), .IN2(n9693), .Q(n9217) );
  NOR2X0 U10416 ( .IN1(n9218), .IN2(n9219), .QN(n9207) );
  NOR2X0 U10417 ( .IN1(n4387), .IN2(n6717), .QN(n9219) );
  INVX0 U10418 ( .INP(n2245), .ZN(n6717) );
  NOR2X0 U10419 ( .IN1(DFF_383_n1), .IN2(n4747), .QN(n9218) );
  INVX0 U10420 ( .INP(n2152), .ZN(n6017) );
  NOR2X0 U10421 ( .IN1(n5421), .IN2(WX1778), .QN(WX1839) );
  NOR2X0 U10422 ( .IN1(n5421), .IN2(n9220), .QN(WX1326) );
  XOR2X1 U10423 ( .IN1(n4664), .IN2(DFF_190_n1), .Q(n9220) );
  NOR2X0 U10424 ( .IN1(n5421), .IN2(n9221), .QN(WX1324) );
  XOR2X1 U10425 ( .IN1(n4630), .IN2(DFF_189_n1), .Q(n9221) );
  NOR2X0 U10426 ( .IN1(n5421), .IN2(n9222), .QN(WX1322) );
  XOR2X1 U10427 ( .IN1(n4633), .IN2(DFF_188_n1), .Q(n9222) );
  NOR2X0 U10428 ( .IN1(n5421), .IN2(n9223), .QN(WX1320) );
  XOR2X1 U10429 ( .IN1(n4637), .IN2(DFF_187_n1), .Q(n9223) );
  NOR2X0 U10430 ( .IN1(n5422), .IN2(n9224), .QN(WX1318) );
  XOR2X1 U10431 ( .IN1(n4640), .IN2(DFF_186_n1), .Q(n9224) );
  NOR2X0 U10432 ( .IN1(n5422), .IN2(n9225), .QN(WX1316) );
  XOR2X1 U10433 ( .IN1(n4641), .IN2(DFF_185_n1), .Q(n9225) );
  NOR2X0 U10434 ( .IN1(n5422), .IN2(n9226), .QN(WX1314) );
  XOR2X1 U10435 ( .IN1(n4645), .IN2(DFF_184_n1), .Q(n9226) );
  NOR2X0 U10436 ( .IN1(n5422), .IN2(n9227), .QN(WX1312) );
  XOR2X1 U10437 ( .IN1(n4648), .IN2(DFF_183_n1), .Q(n9227) );
  NOR2X0 U10438 ( .IN1(n5422), .IN2(n9228), .QN(WX1310) );
  XOR2X1 U10439 ( .IN1(n4650), .IN2(DFF_182_n1), .Q(n9228) );
  NOR2X0 U10440 ( .IN1(n5422), .IN2(n9229), .QN(WX1308) );
  XOR2X1 U10441 ( .IN1(n4656), .IN2(DFF_181_n1), .Q(n9229) );
  NOR2X0 U10442 ( .IN1(n5422), .IN2(n9230), .QN(WX1306) );
  XOR2X1 U10443 ( .IN1(n4660), .IN2(DFF_180_n1), .Q(n9230) );
  NOR2X0 U10444 ( .IN1(n5422), .IN2(n9231), .QN(WX1304) );
  XNOR2X1 U10445 ( .IN1(n4662), .IN2(test_so10), .Q(n9231) );
  NOR2X0 U10446 ( .IN1(n5422), .IN2(n9232), .QN(WX1302) );
  XOR2X1 U10447 ( .IN1(n4632), .IN2(DFF_178_n1), .Q(n9232) );
  NOR2X0 U10448 ( .IN1(n5422), .IN2(n9233), .QN(WX1300) );
  XOR2X1 U10449 ( .IN1(n4639), .IN2(DFF_177_n1), .Q(n9233) );
  NOR2X0 U10450 ( .IN1(n5422), .IN2(n9234), .QN(WX1298) );
  XOR2X1 U10451 ( .IN1(n4644), .IN2(DFF_176_n1), .Q(n9234) );
  NOR2X0 U10452 ( .IN1(n5423), .IN2(n9235), .QN(WX1296) );
  XOR2X1 U10453 ( .IN1(DFF_175_n1), .IN2(n9236), .Q(n9235) );
  XOR2X1 U10454 ( .IN1(test_so8), .IN2(DFF_191_n1), .Q(n9236) );
  NOR2X0 U10455 ( .IN1(n5423), .IN2(n9237), .QN(WX1294) );
  XOR2X1 U10456 ( .IN1(n4658), .IN2(DFF_174_n1), .Q(n9237) );
  NOR2X0 U10457 ( .IN1(n5423), .IN2(n9238), .QN(WX1292) );
  XOR2X1 U10458 ( .IN1(n4665), .IN2(DFF_173_n1), .Q(n9238) );
  NOR2X0 U10459 ( .IN1(n5423), .IN2(n9239), .QN(WX1290) );
  XOR2X1 U10460 ( .IN1(n4634), .IN2(DFF_172_n1), .Q(n9239) );
  NOR2X0 U10461 ( .IN1(n5423), .IN2(n9240), .QN(WX1288) );
  XOR2X1 U10462 ( .IN1(n4646), .IN2(DFF_171_n1), .Q(n9240) );
  NOR2X0 U10463 ( .IN1(n5423), .IN2(n9241), .QN(WX1286) );
  XOR2X1 U10464 ( .IN1(CRC_OUT_9_10), .IN2(n9242), .Q(n9241) );
  XOR2X1 U10465 ( .IN1(n4669), .IN2(DFF_191_n1), .Q(n9242) );
  NOR2X0 U10466 ( .IN1(n5423), .IN2(n9243), .QN(WX1284) );
  XOR2X1 U10467 ( .IN1(n4642), .IN2(DFF_169_n1), .Q(n9243) );
  NOR2X0 U10468 ( .IN1(n5423), .IN2(n9244), .QN(WX1282) );
  XOR2X1 U10469 ( .IN1(n4647), .IN2(DFF_168_n1), .Q(n9244) );
  NOR2X0 U10470 ( .IN1(n5423), .IN2(n9245), .QN(WX1280) );
  XOR2X1 U10471 ( .IN1(n4652), .IN2(DFF_167_n1), .Q(n9245) );
  NOR2X0 U10472 ( .IN1(n5423), .IN2(n9246), .QN(WX1278) );
  XOR2X1 U10473 ( .IN1(n4668), .IN2(DFF_166_n1), .Q(n9246) );
  NOR2X0 U10474 ( .IN1(n5423), .IN2(n9247), .QN(WX1276) );
  XOR2X1 U10475 ( .IN1(n4661), .IN2(DFF_165_n1), .Q(n9247) );
  NOR2X0 U10476 ( .IN1(n5423), .IN2(n9248), .QN(WX1274) );
  XOR2X1 U10477 ( .IN1(n4653), .IN2(DFF_164_n1), .Q(n9248) );
  NOR2X0 U10478 ( .IN1(n5423), .IN2(n9249), .QN(WX1272) );
  XOR2X1 U10479 ( .IN1(CRC_OUT_9_3), .IN2(n9250), .Q(n9249) );
  XOR2X1 U10480 ( .IN1(n4654), .IN2(DFF_191_n1), .Q(n9250) );
  NOR2X0 U10481 ( .IN1(n5424), .IN2(n9251), .QN(WX1270) );
  XOR2X1 U10482 ( .IN1(n4631), .IN2(DFF_162_n1), .Q(n9251) );
  NOR2X0 U10483 ( .IN1(n5424), .IN2(n9252), .QN(WX1268) );
  XNOR2X1 U10484 ( .IN1(n4666), .IN2(test_so9), .Q(n9252) );
  NOR2X0 U10485 ( .IN1(n5424), .IN2(n9253), .QN(WX1266) );
  XOR2X1 U10486 ( .IN1(n4635), .IN2(DFF_160_n1), .Q(n9253) );
  NOR2X0 U10487 ( .IN1(n5424), .IN2(n9254), .QN(WX1264) );
  XOR2X1 U10488 ( .IN1(n4671), .IN2(DFF_191_n1), .Q(n9254) );
  NOR2X0 U10489 ( .IN1(n5424), .IN2(n9255), .QN(WX11670) );
  XOR2X1 U10490 ( .IN1(n4417), .IN2(DFF_1726_n1), .Q(n9255) );
  NOR2X0 U10491 ( .IN1(n5424), .IN2(n9256), .QN(WX11668) );
  XOR2X1 U10492 ( .IN1(n4418), .IN2(DFF_1725_n1), .Q(n9256) );
  NOR2X0 U10493 ( .IN1(n5424), .IN2(n9257), .QN(WX11666) );
  XOR2X1 U10494 ( .IN1(n4419), .IN2(DFF_1724_n1), .Q(n9257) );
  NOR2X0 U10495 ( .IN1(n5424), .IN2(n9258), .QN(WX11664) );
  XOR2X1 U10496 ( .IN1(n4420), .IN2(DFF_1723_n1), .Q(n9258) );
  NOR2X0 U10497 ( .IN1(n5424), .IN2(n9259), .QN(WX11662) );
  XOR2X1 U10498 ( .IN1(n4421), .IN2(DFF_1722_n1), .Q(n9259) );
  NOR2X0 U10499 ( .IN1(n5424), .IN2(n9260), .QN(WX11660) );
  XOR2X1 U10500 ( .IN1(n4422), .IN2(DFF_1721_n1), .Q(n9260) );
  NOR2X0 U10501 ( .IN1(n5424), .IN2(n9261), .QN(WX11658) );
  XOR2X1 U10502 ( .IN1(n4423), .IN2(DFF_1720_n1), .Q(n9261) );
  NOR2X0 U10503 ( .IN1(n5424), .IN2(n9262), .QN(WX11656) );
  XOR2X1 U10504 ( .IN1(n4424), .IN2(DFF_1719_n1), .Q(n9262) );
  NOR2X0 U10505 ( .IN1(n5424), .IN2(n9263), .QN(WX11654) );
  XOR2X1 U10506 ( .IN1(n4425), .IN2(DFF_1718_n1), .Q(n9263) );
  NOR2X0 U10507 ( .IN1(n5425), .IN2(n9264), .QN(WX11652) );
  XOR2X1 U10508 ( .IN1(n4426), .IN2(DFF_1717_n1), .Q(n9264) );
  NOR2X0 U10509 ( .IN1(n5425), .IN2(n9265), .QN(WX11650) );
  XOR2X1 U10510 ( .IN1(n4427), .IN2(DFF_1716_n1), .Q(n9265) );
  NOR2X0 U10511 ( .IN1(n5425), .IN2(n9266), .QN(WX11648) );
  XOR2X1 U10512 ( .IN1(n4428), .IN2(DFF_1715_n1), .Q(n9266) );
  NOR2X0 U10513 ( .IN1(n5425), .IN2(n9267), .QN(WX11646) );
  XOR2X1 U10514 ( .IN1(CRC_OUT_1_18), .IN2(test_so97), .Q(n9267) );
  NOR2X0 U10515 ( .IN1(n5425), .IN2(n9268), .QN(WX11644) );
  XOR2X1 U10516 ( .IN1(n4429), .IN2(DFF_1713_n1), .Q(n9268) );
  NOR2X0 U10517 ( .IN1(n5425), .IN2(n9269), .QN(WX11642) );
  XOR2X1 U10518 ( .IN1(n4430), .IN2(DFF_1712_n1), .Q(n9269) );
  NOR2X0 U10519 ( .IN1(n5425), .IN2(n9270), .QN(WX11640) );
  XOR2X1 U10520 ( .IN1(DFF_1711_n1), .IN2(n9271), .Q(n9270) );
  XOR2X1 U10521 ( .IN1(test_so100), .IN2(n4388), .Q(n9271) );
  NOR2X0 U10522 ( .IN1(n5425), .IN2(n9272), .QN(WX11638) );
  XNOR2X1 U10523 ( .IN1(n4431), .IN2(test_so99), .Q(n9272) );
  NOR2X0 U10524 ( .IN1(n5425), .IN2(n9273), .QN(WX11636) );
  XOR2X1 U10525 ( .IN1(n4432), .IN2(DFF_1709_n1), .Q(n9273) );
  NOR2X0 U10526 ( .IN1(n5425), .IN2(n9274), .QN(WX11634) );
  XOR2X1 U10527 ( .IN1(n4433), .IN2(DFF_1708_n1), .Q(n9274) );
  NOR2X0 U10528 ( .IN1(n5425), .IN2(n9275), .QN(WX11632) );
  XOR2X1 U10529 ( .IN1(n4434), .IN2(DFF_1707_n1), .Q(n9275) );
  NOR2X0 U10530 ( .IN1(n5425), .IN2(n9276), .QN(WX11630) );
  XOR2X1 U10531 ( .IN1(DFF_1706_n1), .IN2(n9277), .Q(n9276) );
  XOR2X1 U10532 ( .IN1(test_so100), .IN2(n4389), .Q(n9277) );
  NOR2X0 U10533 ( .IN1(n5425), .IN2(n9278), .QN(WX11628) );
  XOR2X1 U10534 ( .IN1(n4435), .IN2(DFF_1705_n1), .Q(n9278) );
  NOR2X0 U10535 ( .IN1(n5426), .IN2(n9279), .QN(WX11626) );
  XOR2X1 U10536 ( .IN1(n4436), .IN2(DFF_1704_n1), .Q(n9279) );
  NOR2X0 U10537 ( .IN1(n5426), .IN2(n9280), .QN(WX11624) );
  XOR2X1 U10538 ( .IN1(n4437), .IN2(DFF_1703_n1), .Q(n9280) );
  NOR2X0 U10539 ( .IN1(n5426), .IN2(n9281), .QN(WX11622) );
  XOR2X1 U10540 ( .IN1(n4438), .IN2(DFF_1702_n1), .Q(n9281) );
  NOR2X0 U10541 ( .IN1(n5426), .IN2(n9282), .QN(WX11620) );
  XOR2X1 U10542 ( .IN1(n4439), .IN2(DFF_1701_n1), .Q(n9282) );
  NOR2X0 U10543 ( .IN1(n5426), .IN2(n9283), .QN(WX11618) );
  XOR2X1 U10544 ( .IN1(n4440), .IN2(DFF_1700_n1), .Q(n9283) );
  NOR2X0 U10545 ( .IN1(n5426), .IN2(n9284), .QN(WX11616) );
  XOR2X1 U10546 ( .IN1(DFF_1699_n1), .IN2(n9285), .Q(n9284) );
  XOR2X1 U10547 ( .IN1(test_so100), .IN2(n4390), .Q(n9285) );
  NOR2X0 U10548 ( .IN1(n5426), .IN2(n9286), .QN(WX11614) );
  XOR2X1 U10549 ( .IN1(n4441), .IN2(DFF_1698_n1), .Q(n9286) );
  NOR2X0 U10550 ( .IN1(n5426), .IN2(n9287), .QN(WX11612) );
  XOR2X1 U10551 ( .IN1(CRC_OUT_1_1), .IN2(test_so98), .Q(n9287) );
  NOR2X0 U10552 ( .IN1(n5426), .IN2(n9288), .QN(WX11610) );
  XOR2X1 U10553 ( .IN1(n4442), .IN2(DFF_1696_n1), .Q(n9288) );
  NOR2X0 U10554 ( .IN1(n5426), .IN2(n9289), .QN(WX11608) );
  XNOR2X1 U10555 ( .IN1(n4409), .IN2(test_so100), .Q(n9289) );
  NOR2X0 U10556 ( .IN1(n9711), .IN2(n5349), .QN(WX11082) );
  NOR2X0 U10557 ( .IN1(n9712), .IN2(n5349), .QN(WX11080) );
  NOR2X0 U10558 ( .IN1(n9713), .IN2(n5349), .QN(WX11078) );
  NOR2X0 U10559 ( .IN1(n9714), .IN2(n5348), .QN(WX11076) );
  NOR2X0 U10560 ( .IN1(n9715), .IN2(n5348), .QN(WX11074) );
  NOR2X0 U10561 ( .IN1(n9716), .IN2(n5348), .QN(WX11072) );
  NOR2X0 U10562 ( .IN1(n9719), .IN2(n5348), .QN(WX11070) );
  NOR2X0 U10563 ( .IN1(n9720), .IN2(n5348), .QN(WX11068) );
  NOR2X0 U10564 ( .IN1(n9723), .IN2(n5348), .QN(WX11066) );
  NOR2X0 U10565 ( .IN1(n5426), .IN2(n4712), .QN(WX11064) );
  NOR2X0 U10566 ( .IN1(n9724), .IN2(n5348), .QN(WX11062) );
  NOR2X0 U10567 ( .IN1(n9725), .IN2(n5348), .QN(WX11060) );
  NOR2X0 U10568 ( .IN1(n9726), .IN2(n5348), .QN(WX11058) );
  NOR2X0 U10569 ( .IN1(n9727), .IN2(n5348), .QN(WX11056) );
  NOR2X0 U10570 ( .IN1(n9728), .IN2(n5348), .QN(WX11054) );
  NOR2X0 U10571 ( .IN1(n9729), .IN2(n5350), .QN(WX11052) );
  NOR2X0 U10572 ( .IN1(n5426), .IN2(WX10829), .QN(WX10890) );
  NOR2X0 U10573 ( .IN1(n5427), .IN2(n9290), .QN(WX10377) );
  XNOR2X1 U10574 ( .IN1(DFF_1534_n1), .IN2(test_so85), .Q(n9290) );
  NOR2X0 U10575 ( .IN1(n5427), .IN2(n9291), .QN(WX10375) );
  XOR2X1 U10576 ( .IN1(n4443), .IN2(DFF_1533_n1), .Q(n9291) );
  NOR2X0 U10577 ( .IN1(n5427), .IN2(n9292), .QN(WX10373) );
  XOR2X1 U10578 ( .IN1(n4444), .IN2(DFF_1532_n1), .Q(n9292) );
  NOR2X0 U10579 ( .IN1(n5427), .IN2(n9293), .QN(WX10371) );
  XOR2X1 U10580 ( .IN1(n4445), .IN2(DFF_1531_n1), .Q(n9293) );
  NOR2X0 U10581 ( .IN1(n5427), .IN2(n9294), .QN(WX10369) );
  XOR2X1 U10582 ( .IN1(n4446), .IN2(DFF_1530_n1), .Q(n9294) );
  NOR2X0 U10583 ( .IN1(n5427), .IN2(n9295), .QN(WX10367) );
  XOR2X1 U10584 ( .IN1(n4447), .IN2(DFF_1529_n1), .Q(n9295) );
  NOR2X0 U10585 ( .IN1(n5427), .IN2(n9296), .QN(WX10365) );
  XOR2X1 U10586 ( .IN1(n4448), .IN2(DFF_1528_n1), .Q(n9296) );
  NOR2X0 U10587 ( .IN1(n5427), .IN2(n9297), .QN(WX10363) );
  XOR2X1 U10588 ( .IN1(n4449), .IN2(DFF_1527_n1), .Q(n9297) );
  NOR2X0 U10589 ( .IN1(n5427), .IN2(n9298), .QN(WX10361) );
  XOR2X1 U10590 ( .IN1(n4450), .IN2(DFF_1526_n1), .Q(n9298) );
  NOR2X0 U10591 ( .IN1(n5427), .IN2(n9299), .QN(WX10359) );
  XOR2X1 U10592 ( .IN1(n4451), .IN2(DFF_1525_n1), .Q(n9299) );
  NOR2X0 U10593 ( .IN1(n5427), .IN2(n9300), .QN(WX10357) );
  XOR2X1 U10594 ( .IN1(n4452), .IN2(DFF_1524_n1), .Q(n9300) );
  NOR2X0 U10595 ( .IN1(n5427), .IN2(n9301), .QN(WX10355) );
  XNOR2X1 U10596 ( .IN1(n4453), .IN2(test_so88), .Q(n9301) );
  NOR2X0 U10597 ( .IN1(n5427), .IN2(n9302), .QN(WX10353) );
  XOR2X1 U10598 ( .IN1(n4454), .IN2(DFF_1522_n1), .Q(n9302) );
  NOR2X0 U10599 ( .IN1(n5428), .IN2(n9303), .QN(WX10351) );
  XOR2X1 U10600 ( .IN1(n4455), .IN2(DFF_1521_n1), .Q(n9303) );
  NOR2X0 U10601 ( .IN1(n5428), .IN2(n9304), .QN(WX10349) );
  XOR2X1 U10602 ( .IN1(n4456), .IN2(DFF_1520_n1), .Q(n9304) );
  NOR2X0 U10603 ( .IN1(n5428), .IN2(n9305), .QN(WX10347) );
  XNOR2X1 U10604 ( .IN1(DFF_1519_n1), .IN2(n9306), .Q(n9305) );
  XOR2X1 U10605 ( .IN1(n4391), .IN2(DFF_1535_n1), .Q(n9306) );
  NOR2X0 U10606 ( .IN1(n5428), .IN2(n9307), .QN(WX10345) );
  XOR2X1 U10607 ( .IN1(n4457), .IN2(DFF_1518_n1), .Q(n9307) );
  NOR2X0 U10608 ( .IN1(n5428), .IN2(n9308), .QN(WX10343) );
  XNOR2X1 U10609 ( .IN1(DFF_1517_n1), .IN2(test_so86), .Q(n9308) );
  NOR2X0 U10610 ( .IN1(n5428), .IN2(n9309), .QN(WX10341) );
  XOR2X1 U10611 ( .IN1(n4458), .IN2(DFF_1516_n1), .Q(n9309) );
  NOR2X0 U10612 ( .IN1(n5428), .IN2(n9310), .QN(WX10339) );
  XOR2X1 U10613 ( .IN1(n4459), .IN2(DFF_1515_n1), .Q(n9310) );
  NOR2X0 U10614 ( .IN1(n5428), .IN2(n9311), .QN(WX10337) );
  XNOR2X1 U10615 ( .IN1(DFF_1514_n1), .IN2(n9312), .Q(n9311) );
  XOR2X1 U10616 ( .IN1(n4392), .IN2(DFF_1535_n1), .Q(n9312) );
  NOR2X0 U10617 ( .IN1(n5428), .IN2(n9313), .QN(WX10335) );
  XOR2X1 U10618 ( .IN1(n4460), .IN2(DFF_1513_n1), .Q(n9313) );
  NOR2X0 U10619 ( .IN1(n5428), .IN2(n9314), .QN(WX10333) );
  XOR2X1 U10620 ( .IN1(n4461), .IN2(DFF_1512_n1), .Q(n9314) );
  NOR2X0 U10621 ( .IN1(n5428), .IN2(n9315), .QN(WX10331) );
  XOR2X1 U10622 ( .IN1(n4462), .IN2(DFF_1511_n1), .Q(n9315) );
  NOR2X0 U10623 ( .IN1(n5428), .IN2(n9316), .QN(WX10329) );
  XOR2X1 U10624 ( .IN1(n4463), .IN2(DFF_1510_n1), .Q(n9316) );
  NOR2X0 U10625 ( .IN1(n5428), .IN2(n9317), .QN(WX10327) );
  XOR2X1 U10626 ( .IN1(n4464), .IN2(DFF_1509_n1), .Q(n9317) );
  NOR2X0 U10627 ( .IN1(n5429), .IN2(n9318), .QN(WX10325) );
  XOR2X1 U10628 ( .IN1(n4465), .IN2(DFF_1508_n1), .Q(n9318) );
  NOR2X0 U10629 ( .IN1(n5429), .IN2(n9319), .QN(WX10323) );
  XNOR2X1 U10630 ( .IN1(DFF_1507_n1), .IN2(n9320), .Q(n9319) );
  XOR2X1 U10631 ( .IN1(n4393), .IN2(DFF_1535_n1), .Q(n9320) );
  NOR2X0 U10632 ( .IN1(n5429), .IN2(n9321), .QN(WX10321) );
  XNOR2X1 U10633 ( .IN1(n4466), .IN2(test_so87), .Q(n9321) );
  NOR2X0 U10634 ( .IN1(n5429), .IN2(n9322), .QN(WX10319) );
  XOR2X1 U10635 ( .IN1(n4467), .IN2(DFF_1505_n1), .Q(n9322) );
  NOR2X0 U10636 ( .IN1(n5421), .IN2(n9323), .QN(WX10317) );
  XOR2X1 U10637 ( .IN1(n4468), .IN2(DFF_1504_n1), .Q(n9323) );
  NOR2X0 U10638 ( .IN1(n5429), .IN2(n9324), .QN(WX10315) );
  XOR2X1 U10639 ( .IN1(n4410), .IN2(DFF_1535_n1), .Q(n9324) );
  XNOR2X1 U10640 ( .IN1(n9325), .IN2(n6264), .Q(DATA_9_9) );
  XNOR2X1 U10641 ( .IN1(n9326), .IN2(n9327), .Q(n6264) );
  XOR2X1 U10642 ( .IN1(n3485), .IN2(TM0), .Q(n9327) );
  XOR2X1 U10643 ( .IN1(n9328), .IN2(n4647), .Q(n9326) );
  XOR2X1 U10644 ( .IN1(WX753), .IN2(n9730), .Q(n9328) );
  NAND2X0 U10645 ( .IN1(TM0), .IN2(WX529), .QN(n9325) );
  XNOR2X1 U10646 ( .IN1(n9329), .IN2(n6236), .Q(DATA_9_8) );
  XNOR2X1 U10647 ( .IN1(n9330), .IN2(n9331), .Q(n6236) );
  XOR2X1 U10648 ( .IN1(n3483), .IN2(TM0), .Q(n9331) );
  XOR2X1 U10649 ( .IN1(n9332), .IN2(n4652), .Q(n9330) );
  XOR2X1 U10650 ( .IN1(WX819), .IN2(n9731), .Q(n9332) );
  NAND2X0 U10651 ( .IN1(TM0), .IN2(WX531), .QN(n9329) );
  XNOR2X1 U10652 ( .IN1(n9333), .IN2(n6217), .Q(DATA_9_7) );
  XNOR2X1 U10653 ( .IN1(n9334), .IN2(n9335), .Q(n6217) );
  XOR2X1 U10654 ( .IN1(n3481), .IN2(TM0), .Q(n9335) );
  XOR2X1 U10655 ( .IN1(n9336), .IN2(n4667), .Q(n9334) );
  XOR2X1 U10656 ( .IN1(WX821), .IN2(n4668), .Q(n9336) );
  NAND2X0 U10657 ( .IN1(TM0), .IN2(WX533), .QN(n9333) );
  XOR2X1 U10658 ( .IN1(n9337), .IN2(n6201), .Q(DATA_9_6) );
  XNOR2X1 U10659 ( .IN1(n9338), .IN2(n9339), .Q(n6201) );
  XOR2X1 U10660 ( .IN1(n3479), .IN2(TM0), .Q(n9339) );
  XOR2X1 U10661 ( .IN1(n9340), .IN2(n4661), .Q(n9338) );
  XOR2X1 U10662 ( .IN1(WX823), .IN2(test_so5), .Q(n9340) );
  NAND2X0 U10663 ( .IN1(TM0), .IN2(WX535), .QN(n9337) );
  XNOR2X1 U10664 ( .IN1(n9341), .IN2(n6193), .Q(DATA_9_5) );
  XNOR2X1 U10665 ( .IN1(n9342), .IN2(n9343), .Q(n6193) );
  XOR2X1 U10666 ( .IN1(n3477), .IN2(TM0), .Q(n9343) );
  XOR2X1 U10667 ( .IN1(n9344), .IN2(n4653), .Q(n9342) );
  XOR2X1 U10668 ( .IN1(WX825), .IN2(n9732), .Q(n9344) );
  NAND2X0 U10669 ( .IN1(TM0), .IN2(WX537), .QN(n9341) );
  XNOR2X1 U10670 ( .IN1(n9345), .IN2(n6178), .Q(DATA_9_4) );
  XNOR2X1 U10671 ( .IN1(n9346), .IN2(n9347), .Q(n6178) );
  XOR2X1 U10672 ( .IN1(n3475), .IN2(TM0), .Q(n9347) );
  XOR2X1 U10673 ( .IN1(n9348), .IN2(n4654), .Q(n9346) );
  XOR2X1 U10674 ( .IN1(WX827), .IN2(n9733), .Q(n9348) );
  NAND2X0 U10675 ( .IN1(TM0), .IN2(WX539), .QN(n9345) );
  XOR2X1 U10676 ( .IN1(n9349), .IN2(n7472), .Q(DATA_9_31) );
  XOR2X1 U10677 ( .IN1(n9350), .IN2(n9351), .Q(n7472) );
  XOR2X1 U10678 ( .IN1(n3529), .IN2(n5257), .Q(n9351) );
  XOR2X1 U10679 ( .IN1(n9352), .IN2(n4664), .Q(n9350) );
  XOR2X1 U10680 ( .IN1(WX709), .IN2(n9734), .Q(n9352) );
  NAND2X0 U10681 ( .IN1(TM0), .IN2(WX485), .QN(n9349) );
  XNOR2X1 U10682 ( .IN1(n9353), .IN2(n6245), .Q(DATA_9_30) );
  XNOR2X1 U10683 ( .IN1(n9354), .IN2(n9355), .Q(n6245) );
  XOR2X1 U10684 ( .IN1(n3527), .IN2(n5258), .Q(n9355) );
  XOR2X1 U10685 ( .IN1(n9356), .IN2(n4629), .Q(n9354) );
  XOR2X1 U10686 ( .IN1(WX775), .IN2(n4630), .Q(n9356) );
  NAND2X0 U10687 ( .IN1(TM0), .IN2(WX487), .QN(n9353) );
  XNOR2X1 U10688 ( .IN1(n9357), .IN2(n6159), .Q(DATA_9_3) );
  XNOR2X1 U10689 ( .IN1(n9358), .IN2(n9359), .Q(n6159) );
  XOR2X1 U10690 ( .IN1(n3473), .IN2(TM0), .Q(n9359) );
  XOR2X1 U10691 ( .IN1(n9360), .IN2(n4631), .Q(n9358) );
  XOR2X1 U10692 ( .IN1(WX829), .IN2(n9735), .Q(n9360) );
  NAND2X0 U10693 ( .IN1(TM0), .IN2(WX541), .QN(n9357) );
  XNOR2X1 U10694 ( .IN1(n9361), .IN2(n6091), .Q(DATA_9_29) );
  XNOR2X1 U10695 ( .IN1(n9362), .IN2(n9363), .Q(n6091) );
  XOR2X1 U10696 ( .IN1(n3525), .IN2(n5257), .Q(n9363) );
  XOR2X1 U10697 ( .IN1(n9364), .IN2(n4633), .Q(n9362) );
  XOR2X1 U10698 ( .IN1(WX777), .IN2(n9736), .Q(n9364) );
  NAND2X0 U10699 ( .IN1(TM0), .IN2(WX489), .QN(n9361) );
  XOR2X1 U10700 ( .IN1(n9365), .IN2(n6015), .Q(DATA_9_28) );
  XNOR2X1 U10701 ( .IN1(n9366), .IN2(n9367), .Q(n6015) );
  XOR2X1 U10702 ( .IN1(n4637), .IN2(n5258), .Q(n9367) );
  XOR2X1 U10703 ( .IN1(n9368), .IN2(n4638), .Q(n9366) );
  XOR2X1 U10704 ( .IN1(WX779), .IN2(test_so2), .Q(n9368) );
  NAND2X0 U10705 ( .IN1(TM0), .IN2(WX491), .QN(n9365) );
  XNOR2X1 U10706 ( .IN1(n9369), .IN2(n5698), .Q(DATA_9_27) );
  XNOR2X1 U10707 ( .IN1(n9370), .IN2(n9371), .Q(n5698) );
  XOR2X1 U10708 ( .IN1(n3521), .IN2(n5258), .Q(n9371) );
  XOR2X1 U10709 ( .IN1(n9372), .IN2(n4640), .Q(n9370) );
  XOR2X1 U10710 ( .IN1(WX781), .IN2(n9737), .Q(n9372) );
  NAND2X0 U10711 ( .IN1(TM0), .IN2(WX493), .QN(n9369) );
  XNOR2X1 U10712 ( .IN1(n9373), .IN2(n5684), .Q(DATA_9_26) );
  XNOR2X1 U10713 ( .IN1(n9374), .IN2(n9375), .Q(n5684) );
  XOR2X1 U10714 ( .IN1(n3519), .IN2(n5258), .Q(n9375) );
  XOR2X1 U10715 ( .IN1(n9376), .IN2(n4641), .Q(n9374) );
  XOR2X1 U10716 ( .IN1(WX783), .IN2(n9738), .Q(n9376) );
  NAND2X0 U10717 ( .IN1(TM0), .IN2(WX495), .QN(n9373) );
  XNOR2X1 U10718 ( .IN1(n9377), .IN2(n5665), .Q(DATA_9_25) );
  XNOR2X1 U10719 ( .IN1(n9378), .IN2(n9379), .Q(n5665) );
  XOR2X1 U10720 ( .IN1(n3517), .IN2(n5258), .Q(n9379) );
  XOR2X1 U10721 ( .IN1(n9380), .IN2(n4645), .Q(n9378) );
  XOR2X1 U10722 ( .IN1(WX785), .IN2(n9739), .Q(n9380) );
  NAND2X0 U10723 ( .IN1(TM0), .IN2(WX497), .QN(n9377) );
  XOR2X1 U10724 ( .IN1(n9381), .IN2(n7430), .Q(DATA_9_24) );
  XNOR2X1 U10725 ( .IN1(n9382), .IN2(n9383), .Q(n7430) );
  XOR2X1 U10726 ( .IN1(n3515), .IN2(n5258), .Q(n9383) );
  XOR2X1 U10727 ( .IN1(n9384), .IN2(n4648), .Q(n9382) );
  XOR2X1 U10728 ( .IN1(WX787), .IN2(test_so4), .Q(n9384) );
  NAND2X0 U10729 ( .IN1(TM0), .IN2(WX499), .QN(n9381) );
  XNOR2X1 U10730 ( .IN1(n9385), .IN2(n5646), .Q(DATA_9_23) );
  XNOR2X1 U10731 ( .IN1(n9386), .IN2(n9387), .Q(n5646) );
  XOR2X1 U10732 ( .IN1(n3513), .IN2(n5257), .Q(n9387) );
  XOR2X1 U10733 ( .IN1(n9388), .IN2(n4650), .Q(n9386) );
  XOR2X1 U10734 ( .IN1(WX789), .IN2(n9740), .Q(n9388) );
  NAND2X0 U10735 ( .IN1(TM0), .IN2(WX501), .QN(n9385) );
  XNOR2X1 U10736 ( .IN1(n9389), .IN2(n5630), .Q(DATA_9_22) );
  XNOR2X1 U10737 ( .IN1(n9390), .IN2(n9391), .Q(n5630) );
  XOR2X1 U10738 ( .IN1(n3511), .IN2(n5258), .Q(n9391) );
  XOR2X1 U10739 ( .IN1(n9392), .IN2(n4655), .Q(n9390) );
  XOR2X1 U10740 ( .IN1(WX791), .IN2(n4656), .Q(n9392) );
  NAND2X0 U10741 ( .IN1(TM0), .IN2(WX503), .QN(n9389) );
  XNOR2X1 U10742 ( .IN1(n9393), .IN2(n6385), .Q(DATA_9_21) );
  XNOR2X1 U10743 ( .IN1(n9394), .IN2(n9395), .Q(n6385) );
  XOR2X1 U10744 ( .IN1(n3509), .IN2(n5258), .Q(n9395) );
  XOR2X1 U10745 ( .IN1(n9396), .IN2(n4659), .Q(n9394) );
  XOR2X1 U10746 ( .IN1(WX793), .IN2(n4660), .Q(n9396) );
  NAND2X0 U10747 ( .IN1(TM0), .IN2(WX505), .QN(n9393) );
  XOR2X1 U10748 ( .IN1(n9397), .IN2(n7421), .Q(DATA_9_20) );
  XNOR2X1 U10749 ( .IN1(n9398), .IN2(n9399), .Q(n7421) );
  XOR2X1 U10750 ( .IN1(n3507), .IN2(n5258), .Q(n9399) );
  XOR2X1 U10751 ( .IN1(n9400), .IN2(n4662), .Q(n9398) );
  XOR2X1 U10752 ( .IN1(WX731), .IN2(test_so6), .Q(n9400) );
  NAND2X0 U10753 ( .IN1(TM0), .IN2(WX507), .QN(n9397) );
  XOR2X1 U10754 ( .IN1(n9401), .IN2(n6139), .Q(DATA_9_2) );
  XNOR2X1 U10755 ( .IN1(n9402), .IN2(n9403), .Q(n6139) );
  XOR2X1 U10756 ( .IN1(n3471), .IN2(TM0), .Q(n9403) );
  XOR2X1 U10757 ( .IN1(n9404), .IN2(n4666), .Q(n9402) );
  XOR2X1 U10758 ( .IN1(WX767), .IN2(test_so7), .Q(n9404) );
  NAND2X0 U10759 ( .IN1(TM0), .IN2(WX543), .QN(n9401) );
  XNOR2X1 U10760 ( .IN1(n9405), .IN2(n6376), .Q(DATA_9_19) );
  XNOR2X1 U10761 ( .IN1(n9406), .IN2(n9407), .Q(n6376) );
  XOR2X1 U10762 ( .IN1(n3505), .IN2(n5258), .Q(n9407) );
  XOR2X1 U10763 ( .IN1(n9408), .IN2(n4632), .Q(n9406) );
  XOR2X1 U10764 ( .IN1(WX797), .IN2(n9741), .Q(n9408) );
  NAND2X0 U10765 ( .IN1(TM0), .IN2(WX509), .QN(n9405) );
  XNOR2X1 U10766 ( .IN1(n9409), .IN2(n6366), .Q(DATA_9_18) );
  XNOR2X1 U10767 ( .IN1(n9410), .IN2(n9411), .Q(n6366) );
  XOR2X1 U10768 ( .IN1(n3503), .IN2(n5258), .Q(n9411) );
  XOR2X1 U10769 ( .IN1(n9412), .IN2(n4639), .Q(n9410) );
  XOR2X1 U10770 ( .IN1(WX799), .IN2(n9742), .Q(n9412) );
  NAND2X0 U10771 ( .IN1(TM0), .IN2(WX511), .QN(n9409) );
  XNOR2X1 U10772 ( .IN1(n9413), .IN2(n6357), .Q(DATA_9_17) );
  XNOR2X1 U10773 ( .IN1(n9414), .IN2(n9415), .Q(n6357) );
  XOR2X1 U10774 ( .IN1(n3501), .IN2(n5258), .Q(n9415) );
  XOR2X1 U10775 ( .IN1(n9416), .IN2(n4644), .Q(n9414) );
  XOR2X1 U10776 ( .IN1(WX801), .IN2(n9743), .Q(n9416) );
  NAND2X0 U10777 ( .IN1(TM0), .IN2(WX513), .QN(n9413) );
  XOR2X1 U10778 ( .IN1(n9417), .IN2(n7412), .Q(DATA_9_16) );
  XNOR2X1 U10779 ( .IN1(n9418), .IN2(n9419), .Q(n7412) );
  XOR2X1 U10780 ( .IN1(n3499), .IN2(n5247), .Q(n9419) );
  XOR2X1 U10781 ( .IN1(n9420), .IN2(n4651), .Q(n9418) );
  XOR2X1 U10782 ( .IN1(WX739), .IN2(test_so8), .Q(n9420) );
  NAND2X0 U10783 ( .IN1(TM0), .IN2(WX515), .QN(n9417) );
  XNOR2X1 U10784 ( .IN1(n9421), .IN2(n6340), .Q(DATA_9_15) );
  XNOR2X1 U10785 ( .IN1(n9422), .IN2(n9423), .Q(n6340) );
  XOR2X1 U10786 ( .IN1(n3497), .IN2(TM0), .Q(n9423) );
  XOR2X1 U10787 ( .IN1(n9424), .IN2(n4657), .Q(n9422) );
  XOR2X1 U10788 ( .IN1(WX805), .IN2(n4658), .Q(n9424) );
  NAND2X0 U10789 ( .IN1(TM0), .IN2(WX517), .QN(n9421) );
  XNOR2X1 U10790 ( .IN1(n9425), .IN2(n6321), .Q(DATA_9_14) );
  XNOR2X1 U10791 ( .IN1(n9426), .IN2(n9427), .Q(n6321) );
  XOR2X1 U10792 ( .IN1(n3495), .IN2(TM0), .Q(n9427) );
  XOR2X1 U10793 ( .IN1(n9428), .IN2(n4665), .Q(n9426) );
  XOR2X1 U10794 ( .IN1(WX807), .IN2(n9744), .Q(n9428) );
  NAND2X0 U10795 ( .IN1(test_so1), .IN2(TM0), .QN(n9425) );
  XNOR2X1 U10796 ( .IN1(n9429), .IN2(n6302), .Q(DATA_9_13) );
  XNOR2X1 U10797 ( .IN1(n9430), .IN2(n9431), .Q(n6302) );
  XOR2X1 U10798 ( .IN1(n3493), .IN2(TM0), .Q(n9431) );
  XOR2X1 U10799 ( .IN1(n9432), .IN2(n4634), .Q(n9430) );
  XOR2X1 U10800 ( .IN1(WX809), .IN2(n9745), .Q(n9432) );
  NAND2X0 U10801 ( .IN1(TM0), .IN2(WX521), .QN(n9429) );
  XNOR2X1 U10802 ( .IN1(n9433), .IN2(n6287), .Q(DATA_9_12) );
  XNOR2X1 U10803 ( .IN1(n9434), .IN2(n9435), .Q(n6287) );
  XOR2X1 U10804 ( .IN1(n3491), .IN2(TM0), .Q(n9435) );
  XOR2X1 U10805 ( .IN1(n9436), .IN2(n4646), .Q(n9434) );
  XOR2X1 U10806 ( .IN1(WX811), .IN2(n9746), .Q(n9436) );
  NAND2X0 U10807 ( .IN1(TM0), .IN2(WX523), .QN(n9433) );
  XNOR2X1 U10808 ( .IN1(n9437), .IN2(n6278), .Q(DATA_9_11) );
  XNOR2X1 U10809 ( .IN1(n9438), .IN2(n9439), .Q(n6278) );
  XOR2X1 U10810 ( .IN1(n3489), .IN2(TM0), .Q(n9439) );
  XOR2X1 U10811 ( .IN1(n9440), .IN2(n4669), .Q(n9438) );
  XOR2X1 U10812 ( .IN1(WX813), .IN2(n9747), .Q(n9440) );
  NAND2X0 U10813 ( .IN1(TM0), .IN2(WX525), .QN(n9437) );
  XNOR2X1 U10814 ( .IN1(n9441), .IN2(n7403), .Q(DATA_9_10) );
  XOR2X1 U10815 ( .IN1(n9442), .IN2(n9443), .Q(n7403) );
  XOR2X1 U10816 ( .IN1(n4642), .IN2(TM0), .Q(n9443) );
  XOR2X1 U10817 ( .IN1(n9444), .IN2(n4643), .Q(n9442) );
  XOR2X1 U10818 ( .IN1(WX815), .IN2(test_so3), .Q(n9444) );
  NAND2X0 U10819 ( .IN1(TM0), .IN2(WX527), .QN(n9441) );
  XNOR2X1 U10820 ( .IN1(n9445), .IN2(n6125), .Q(DATA_9_1) );
  XNOR2X1 U10821 ( .IN1(n9446), .IN2(n9447), .Q(n6125) );
  XOR2X1 U10822 ( .IN1(n3469), .IN2(TM0), .Q(n9447) );
  XOR2X1 U10823 ( .IN1(n9448), .IN2(n4635), .Q(n9446) );
  XOR2X1 U10824 ( .IN1(WX833), .IN2(n9748), .Q(n9448) );
  NAND2X0 U10825 ( .IN1(TM0), .IN2(WX545), .QN(n9445) );
  XNOR2X1 U10826 ( .IN1(n9449), .IN2(n6115), .Q(DATA_9_0) );
  XNOR2X1 U10827 ( .IN1(n9450), .IN2(n9451), .Q(n6115) );
  XOR2X1 U10828 ( .IN1(n3467), .IN2(TM0), .Q(n9451) );
  XOR2X1 U10829 ( .IN1(n9452), .IN2(n4670), .Q(n9450) );
  XOR2X1 U10830 ( .IN1(WX835), .IN2(n4671), .Q(n9452) );
  NAND2X0 U10831 ( .IN1(TM0), .IN2(WX547), .QN(n9449) );
  NOR2X0 U3558_U2 ( .IN1(n5413), .IN2(U3558_n1), .QN(n2245) );
  INVX0 U3558_U1 ( .INP(n4805), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(n3278), .ZN(U3871_n1) );
  NOR2X0 U3871_U1 ( .IN1(TM0), .IN2(U3871_n1), .QN(n2153) );
  INVX0 U3991_U2 ( .INP(n3278), .ZN(U3991_n1) );
  NOR2X0 U3991_U1 ( .IN1(n583), .IN2(U3991_n1), .QN(n2152) );
  INVX0 U5716_U2 ( .INP(WX547), .ZN(U5716_n1) );
  NOR2X0 U5716_U1 ( .IN1(n5398), .IN2(U5716_n1), .QN(WX544) );
  INVX0 U5717_U2 ( .INP(WX545), .ZN(U5717_n1) );
  NOR2X0 U5717_U1 ( .IN1(n5378), .IN2(U5717_n1), .QN(WX542) );
  INVX0 U5718_U2 ( .INP(WX543), .ZN(U5718_n1) );
  NOR2X0 U5718_U1 ( .IN1(n5393), .IN2(U5718_n1), .QN(WX540) );
  INVX0 U5719_U2 ( .INP(WX541), .ZN(U5719_n1) );
  NOR2X0 U5719_U1 ( .IN1(n5388), .IN2(U5719_n1), .QN(WX538) );
  INVX0 U5720_U2 ( .INP(WX539), .ZN(U5720_n1) );
  NOR2X0 U5720_U1 ( .IN1(n5388), .IN2(U5720_n1), .QN(WX536) );
  INVX0 U5721_U2 ( .INP(WX537), .ZN(U5721_n1) );
  NOR2X0 U5721_U1 ( .IN1(n5388), .IN2(U5721_n1), .QN(WX534) );
  INVX0 U5722_U2 ( .INP(WX535), .ZN(U5722_n1) );
  NOR2X0 U5722_U1 ( .IN1(n5389), .IN2(U5722_n1), .QN(WX532) );
  INVX0 U5723_U2 ( .INP(WX533), .ZN(U5723_n1) );
  NOR2X0 U5723_U1 ( .IN1(n5389), .IN2(U5723_n1), .QN(WX530) );
  INVX0 U5724_U2 ( .INP(WX531), .ZN(U5724_n1) );
  NOR2X0 U5724_U1 ( .IN1(n5389), .IN2(U5724_n1), .QN(WX528) );
  INVX0 U5725_U2 ( .INP(WX529), .ZN(U5725_n1) );
  NOR2X0 U5725_U1 ( .IN1(n5389), .IN2(U5725_n1), .QN(WX526) );
  INVX0 U5726_U2 ( .INP(WX527), .ZN(U5726_n1) );
  NOR2X0 U5726_U1 ( .IN1(n5389), .IN2(U5726_n1), .QN(WX524) );
  INVX0 U5727_U2 ( .INP(WX525), .ZN(U5727_n1) );
  NOR2X0 U5727_U1 ( .IN1(n5389), .IN2(U5727_n1), .QN(WX522) );
  INVX0 U5728_U2 ( .INP(WX523), .ZN(U5728_n1) );
  NOR2X0 U5728_U1 ( .IN1(n5389), .IN2(U5728_n1), .QN(WX520) );
  INVX0 U5729_U2 ( .INP(WX521), .ZN(U5729_n1) );
  NOR2X0 U5729_U1 ( .IN1(n5389), .IN2(U5729_n1), .QN(WX518) );
  INVX0 U5730_U2 ( .INP(test_so1), .ZN(U5730_n1) );
  NOR2X0 U5730_U1 ( .IN1(n5389), .IN2(U5730_n1), .QN(WX516) );
  INVX0 U5731_U2 ( .INP(WX517), .ZN(U5731_n1) );
  NOR2X0 U5731_U1 ( .IN1(n5389), .IN2(U5731_n1), .QN(WX514) );
  INVX0 U5732_U2 ( .INP(WX515), .ZN(U5732_n1) );
  NOR2X0 U5732_U1 ( .IN1(n5389), .IN2(U5732_n1), .QN(WX512) );
  INVX0 U5733_U2 ( .INP(WX513), .ZN(U5733_n1) );
  NOR2X0 U5733_U1 ( .IN1(n5390), .IN2(U5733_n1), .QN(WX510) );
  INVX0 U5734_U2 ( .INP(WX511), .ZN(U5734_n1) );
  NOR2X0 U5734_U1 ( .IN1(n5390), .IN2(U5734_n1), .QN(WX508) );
  INVX0 U5735_U2 ( .INP(WX509), .ZN(U5735_n1) );
  NOR2X0 U5735_U1 ( .IN1(n5390), .IN2(U5735_n1), .QN(WX506) );
  INVX0 U5736_U2 ( .INP(WX507), .ZN(U5736_n1) );
  NOR2X0 U5736_U1 ( .IN1(n5390), .IN2(U5736_n1), .QN(WX504) );
  INVX0 U5737_U2 ( .INP(WX505), .ZN(U5737_n1) );
  NOR2X0 U5737_U1 ( .IN1(n5390), .IN2(U5737_n1), .QN(WX502) );
  INVX0 U5738_U2 ( .INP(WX503), .ZN(U5738_n1) );
  NOR2X0 U5738_U1 ( .IN1(n5390), .IN2(U5738_n1), .QN(WX500) );
  INVX0 U5739_U2 ( .INP(WX501), .ZN(U5739_n1) );
  NOR2X0 U5739_U1 ( .IN1(n5390), .IN2(U5739_n1), .QN(WX498) );
  INVX0 U5740_U2 ( .INP(WX499), .ZN(U5740_n1) );
  NOR2X0 U5740_U1 ( .IN1(n5390), .IN2(U5740_n1), .QN(WX496) );
  INVX0 U5741_U2 ( .INP(WX497), .ZN(U5741_n1) );
  NOR2X0 U5741_U1 ( .IN1(n5390), .IN2(U5741_n1), .QN(WX494) );
  INVX0 U5742_U2 ( .INP(WX495), .ZN(U5742_n1) );
  NOR2X0 U5742_U1 ( .IN1(n5390), .IN2(U5742_n1), .QN(WX492) );
  INVX0 U5743_U2 ( .INP(WX493), .ZN(U5743_n1) );
  NOR2X0 U5743_U1 ( .IN1(n5390), .IN2(U5743_n1), .QN(WX490) );
  INVX0 U5744_U2 ( .INP(WX491), .ZN(U5744_n1) );
  NOR2X0 U5744_U1 ( .IN1(n5391), .IN2(U5744_n1), .QN(WX488) );
  INVX0 U5745_U2 ( .INP(WX489), .ZN(U5745_n1) );
  NOR2X0 U5745_U1 ( .IN1(n5391), .IN2(U5745_n1), .QN(WX486) );
  INVX0 U5746_U2 ( .INP(WX487), .ZN(U5746_n1) );
  NOR2X0 U5746_U1 ( .IN1(n5391), .IN2(U5746_n1), .QN(WX484) );
  INVX0 U5747_U2 ( .INP(WX5939), .ZN(U5747_n1) );
  NOR2X0 U5747_U1 ( .IN1(n5391), .IN2(U5747_n1), .QN(WX6002) );
  INVX0 U5748_U2 ( .INP(test_so49), .ZN(U5748_n1) );
  NOR2X0 U5748_U1 ( .IN1(n5391), .IN2(U5748_n1), .QN(WX6000) );
  INVX0 U5749_U2 ( .INP(WX5935), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n5391), .IN2(U5749_n1), .QN(WX5998) );
  INVX0 U5750_U2 ( .INP(WX5933), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n5391), .IN2(U5750_n1), .QN(WX5996) );
  INVX0 U5751_U2 ( .INP(WX5931), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n5391), .IN2(U5751_n1), .QN(WX5994) );
  INVX0 U5752_U2 ( .INP(WX3269), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n5391), .IN2(U5752_n1), .QN(WX3332) );
  INVX0 U5753_U2 ( .INP(WX3265), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n5391), .IN2(U5753_n1), .QN(WX3328) );
  INVX0 U5754_U2 ( .INP(WX3263), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n5391), .IN2(U5754_n1), .QN(WX3326) );
  INVX0 U5755_U2 ( .INP(WX11179), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n5392), .IN2(U5755_n1), .QN(WX11242) );
  INVX0 U5756_U2 ( .INP(WX11177), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n5392), .IN2(U5756_n1), .QN(WX11240) );
  INVX0 U5757_U2 ( .INP(WX11175), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n5392), .IN2(U5757_n1), .QN(WX11238) );
  INVX0 U5758_U2 ( .INP(WX11173), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n5392), .IN2(U5758_n1), .QN(WX11236) );
  INVX0 U5759_U2 ( .INP(test_so96), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n5392), .IN2(U5759_n1), .QN(WX11234) );
  INVX0 U5760_U2 ( .INP(WX11169), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n5392), .IN2(U5760_n1), .QN(WX11232) );
  INVX0 U5761_U2 ( .INP(WX11167), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n5392), .IN2(U5761_n1), .QN(WX11230) );
  INVX0 U5762_U2 ( .INP(WX11165), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n5392), .IN2(U5762_n1), .QN(WX11228) );
  INVX0 U5763_U2 ( .INP(WX11163), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n5392), .IN2(U5763_n1), .QN(WX11226) );
  INVX0 U5764_U2 ( .INP(WX11161), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n5392), .IN2(U5764_n1), .QN(WX11224) );
  INVX0 U5765_U2 ( .INP(WX11159), .ZN(U5765_n1) );
  NOR2X0 U5765_U1 ( .IN1(n5392), .IN2(U5765_n1), .QN(WX11222) );
  INVX0 U5766_U2 ( .INP(WX11157), .ZN(U5766_n1) );
  NOR2X0 U5766_U1 ( .IN1(n5393), .IN2(U5766_n1), .QN(WX11220) );
  INVX0 U5767_U2 ( .INP(WX11155), .ZN(U5767_n1) );
  NOR2X0 U5767_U1 ( .IN1(n5393), .IN2(U5767_n1), .QN(WX11218) );
  INVX0 U5768_U2 ( .INP(WX11153), .ZN(U5768_n1) );
  NOR2X0 U5768_U1 ( .IN1(n5393), .IN2(U5768_n1), .QN(WX11216) );
  INVX0 U5769_U2 ( .INP(WX11151), .ZN(U5769_n1) );
  NOR2X0 U5769_U1 ( .IN1(n5393), .IN2(U5769_n1), .QN(WX11214) );
  INVX0 U5770_U2 ( .INP(WX11149), .ZN(U5770_n1) );
  NOR2X0 U5770_U1 ( .IN1(n5393), .IN2(U5770_n1), .QN(WX11212) );
  INVX0 U5771_U2 ( .INP(WX11147), .ZN(U5771_n1) );
  NOR2X0 U5771_U1 ( .IN1(n5393), .IN2(U5771_n1), .QN(WX11210) );
  INVX0 U5772_U2 ( .INP(WX11145), .ZN(U5772_n1) );
  NOR2X0 U5772_U1 ( .IN1(n5393), .IN2(U5772_n1), .QN(WX11208) );
  INVX0 U5773_U2 ( .INP(WX11143), .ZN(U5773_n1) );
  NOR2X0 U5773_U1 ( .IN1(n5393), .IN2(U5773_n1), .QN(WX11206) );
  INVX0 U5774_U2 ( .INP(WX11141), .ZN(U5774_n1) );
  NOR2X0 U5774_U1 ( .IN1(n5393), .IN2(U5774_n1), .QN(WX11204) );
  INVX0 U5775_U2 ( .INP(WX11139), .ZN(U5775_n1) );
  NOR2X0 U5775_U1 ( .IN1(n5393), .IN2(U5775_n1), .QN(WX11202) );
  INVX0 U5776_U2 ( .INP(test_so95), .ZN(U5776_n1) );
  NOR2X0 U5776_U1 ( .IN1(n5394), .IN2(U5776_n1), .QN(WX11200) );
  INVX0 U5777_U2 ( .INP(WX11135), .ZN(U5777_n1) );
  NOR2X0 U5777_U1 ( .IN1(n5394), .IN2(U5777_n1), .QN(WX11198) );
  INVX0 U5778_U2 ( .INP(WX11133), .ZN(U5778_n1) );
  NOR2X0 U5778_U1 ( .IN1(n5394), .IN2(U5778_n1), .QN(WX11196) );
  INVX0 U5779_U2 ( .INP(WX11131), .ZN(U5779_n1) );
  NOR2X0 U5779_U1 ( .IN1(n5394), .IN2(U5779_n1), .QN(WX11194) );
  INVX0 U5780_U2 ( .INP(WX11129), .ZN(U5780_n1) );
  NOR2X0 U5780_U1 ( .IN1(n5394), .IN2(U5780_n1), .QN(WX11192) );
  INVX0 U5781_U2 ( .INP(WX11127), .ZN(U5781_n1) );
  NOR2X0 U5781_U1 ( .IN1(n5394), .IN2(U5781_n1), .QN(WX11190) );
  INVX0 U5782_U2 ( .INP(WX11125), .ZN(U5782_n1) );
  NOR2X0 U5782_U1 ( .IN1(n5394), .IN2(U5782_n1), .QN(WX11188) );
  INVX0 U5783_U2 ( .INP(WX11123), .ZN(U5783_n1) );
  NOR2X0 U5783_U1 ( .IN1(n5394), .IN2(U5783_n1), .QN(WX11186) );
  INVX0 U5784_U2 ( .INP(WX11121), .ZN(U5784_n1) );
  NOR2X0 U5784_U1 ( .IN1(n5394), .IN2(U5784_n1), .QN(WX11184) );
  INVX0 U5785_U2 ( .INP(WX11119), .ZN(U5785_n1) );
  NOR2X0 U5785_U1 ( .IN1(n5394), .IN2(U5785_n1), .QN(WX11182) );
  INVX0 U5786_U2 ( .INP(WX11117), .ZN(U5786_n1) );
  NOR2X0 U5786_U1 ( .IN1(n5394), .IN2(U5786_n1), .QN(WX11180) );
  INVX0 U5787_U2 ( .INP(WX11115), .ZN(U5787_n1) );
  NOR2X0 U5787_U1 ( .IN1(n5395), .IN2(U5787_n1), .QN(WX11178) );
  INVX0 U5788_U2 ( .INP(WX11113), .ZN(U5788_n1) );
  NOR2X0 U5788_U1 ( .IN1(n5395), .IN2(U5788_n1), .QN(WX11176) );
  INVX0 U5789_U2 ( .INP(WX11111), .ZN(U5789_n1) );
  NOR2X0 U5789_U1 ( .IN1(n5395), .IN2(U5789_n1), .QN(WX11174) );
  INVX0 U5790_U2 ( .INP(WX11109), .ZN(U5790_n1) );
  NOR2X0 U5790_U1 ( .IN1(n5395), .IN2(U5790_n1), .QN(WX11172) );
  INVX0 U5791_U2 ( .INP(WX11107), .ZN(U5791_n1) );
  NOR2X0 U5791_U1 ( .IN1(n5395), .IN2(U5791_n1), .QN(WX11170) );
  INVX0 U5792_U2 ( .INP(WX11105), .ZN(U5792_n1) );
  NOR2X0 U5792_U1 ( .IN1(n5395), .IN2(U5792_n1), .QN(WX11168) );
  INVX0 U5793_U2 ( .INP(test_so94), .ZN(U5793_n1) );
  NOR2X0 U5793_U1 ( .IN1(n5395), .IN2(U5793_n1), .QN(WX11166) );
  INVX0 U5794_U2 ( .INP(WX11101), .ZN(U5794_n1) );
  NOR2X0 U5794_U1 ( .IN1(n5395), .IN2(U5794_n1), .QN(WX11164) );
  INVX0 U5795_U2 ( .INP(WX11099), .ZN(U5795_n1) );
  NOR2X0 U5795_U1 ( .IN1(n5395), .IN2(U5795_n1), .QN(WX11162) );
  INVX0 U5796_U2 ( .INP(WX11097), .ZN(U5796_n1) );
  NOR2X0 U5796_U1 ( .IN1(n5395), .IN2(U5796_n1), .QN(WX11160) );
  INVX0 U5797_U2 ( .INP(WX11095), .ZN(U5797_n1) );
  NOR2X0 U5797_U1 ( .IN1(n5395), .IN2(U5797_n1), .QN(WX11158) );
  INVX0 U5798_U2 ( .INP(WX11093), .ZN(U5798_n1) );
  NOR2X0 U5798_U1 ( .IN1(n5396), .IN2(U5798_n1), .QN(WX11156) );
  INVX0 U5799_U2 ( .INP(WX11091), .ZN(U5799_n1) );
  NOR2X0 U5799_U1 ( .IN1(n5396), .IN2(U5799_n1), .QN(WX11154) );
  INVX0 U5800_U2 ( .INP(WX11089), .ZN(U5800_n1) );
  NOR2X0 U5800_U1 ( .IN1(n5396), .IN2(U5800_n1), .QN(WX11152) );
  INVX0 U5801_U2 ( .INP(WX11087), .ZN(U5801_n1) );
  NOR2X0 U5801_U1 ( .IN1(n5396), .IN2(U5801_n1), .QN(WX11150) );
  INVX0 U5802_U2 ( .INP(WX11085), .ZN(U5802_n1) );
  NOR2X0 U5802_U1 ( .IN1(n5396), .IN2(U5802_n1), .QN(WX11148) );
  INVX0 U5803_U2 ( .INP(WX11083), .ZN(U5803_n1) );
  NOR2X0 U5803_U1 ( .IN1(n5396), .IN2(U5803_n1), .QN(WX11146) );
  INVX0 U5804_U2 ( .INP(WX11081), .ZN(U5804_n1) );
  NOR2X0 U5804_U1 ( .IN1(n5396), .IN2(U5804_n1), .QN(WX11144) );
  INVX0 U5805_U2 ( .INP(WX11079), .ZN(U5805_n1) );
  NOR2X0 U5805_U1 ( .IN1(n5396), .IN2(U5805_n1), .QN(WX11142) );
  INVX0 U5806_U2 ( .INP(WX11077), .ZN(U5806_n1) );
  NOR2X0 U5806_U1 ( .IN1(n5396), .IN2(U5806_n1), .QN(WX11140) );
  INVX0 U5807_U2 ( .INP(WX11075), .ZN(U5807_n1) );
  NOR2X0 U5807_U1 ( .IN1(n5396), .IN2(U5807_n1), .QN(WX11138) );
  INVX0 U5808_U2 ( .INP(WX11073), .ZN(U5808_n1) );
  NOR2X0 U5808_U1 ( .IN1(n5396), .IN2(U5808_n1), .QN(WX11136) );
  INVX0 U5809_U2 ( .INP(WX11071), .ZN(U5809_n1) );
  NOR2X0 U5809_U1 ( .IN1(n5397), .IN2(U5809_n1), .QN(WX11134) );
  INVX0 U5810_U2 ( .INP(test_so93), .ZN(U5810_n1) );
  NOR2X0 U5810_U1 ( .IN1(n5397), .IN2(U5810_n1), .QN(WX11132) );
  INVX0 U5811_U2 ( .INP(WX11067), .ZN(U5811_n1) );
  NOR2X0 U5811_U1 ( .IN1(n5397), .IN2(U5811_n1), .QN(WX11130) );
  INVX0 U5812_U2 ( .INP(WX11065), .ZN(U5812_n1) );
  NOR2X0 U5812_U1 ( .IN1(n5397), .IN2(U5812_n1), .QN(WX11128) );
  INVX0 U5813_U2 ( .INP(WX11063), .ZN(U5813_n1) );
  NOR2X0 U5813_U1 ( .IN1(n5397), .IN2(U5813_n1), .QN(WX11126) );
  INVX0 U5814_U2 ( .INP(WX11061), .ZN(U5814_n1) );
  NOR2X0 U5814_U1 ( .IN1(n5397), .IN2(U5814_n1), .QN(WX11124) );
  INVX0 U5815_U2 ( .INP(WX11059), .ZN(U5815_n1) );
  NOR2X0 U5815_U1 ( .IN1(n5397), .IN2(U5815_n1), .QN(WX11122) );
  INVX0 U5816_U2 ( .INP(WX11057), .ZN(U5816_n1) );
  NOR2X0 U5816_U1 ( .IN1(n5397), .IN2(U5816_n1), .QN(WX11120) );
  INVX0 U5817_U2 ( .INP(WX11055), .ZN(U5817_n1) );
  NOR2X0 U5817_U1 ( .IN1(n5397), .IN2(U5817_n1), .QN(WX11118) );
  INVX0 U5818_U2 ( .INP(WX11053), .ZN(U5818_n1) );
  NOR2X0 U5818_U1 ( .IN1(n5397), .IN2(U5818_n1), .QN(WX11116) );
  INVX0 U5819_U2 ( .INP(WX11051), .ZN(U5819_n1) );
  NOR2X0 U5819_U1 ( .IN1(n5397), .IN2(U5819_n1), .QN(WX11114) );
  INVX0 U5820_U2 ( .INP(WX11049), .ZN(U5820_n1) );
  NOR2X0 U5820_U1 ( .IN1(n5398), .IN2(U5820_n1), .QN(WX11112) );
  INVX0 U5821_U2 ( .INP(WX11047), .ZN(U5821_n1) );
  NOR2X0 U5821_U1 ( .IN1(n5398), .IN2(U5821_n1), .QN(WX11110) );
  INVX0 U5822_U2 ( .INP(WX11045), .ZN(U5822_n1) );
  NOR2X0 U5822_U1 ( .IN1(n5398), .IN2(U5822_n1), .QN(WX11108) );
  INVX0 U5823_U2 ( .INP(WX11043), .ZN(U5823_n1) );
  NOR2X0 U5823_U1 ( .IN1(n5398), .IN2(U5823_n1), .QN(WX11106) );
  INVX0 U5824_U2 ( .INP(WX11041), .ZN(U5824_n1) );
  NOR2X0 U5824_U1 ( .IN1(n5398), .IN2(U5824_n1), .QN(WX11104) );
  INVX0 U5825_U2 ( .INP(WX11039), .ZN(U5825_n1) );
  NOR2X0 U5825_U1 ( .IN1(n5398), .IN2(U5825_n1), .QN(WX11102) );
  INVX0 U5826_U2 ( .INP(WX11037), .ZN(U5826_n1) );
  NOR2X0 U5826_U1 ( .IN1(n5398), .IN2(U5826_n1), .QN(WX11100) );
  INVX0 U5827_U2 ( .INP(test_so92), .ZN(U5827_n1) );
  NOR2X0 U5827_U1 ( .IN1(n5398), .IN2(U5827_n1), .QN(WX11098) );
  INVX0 U5828_U2 ( .INP(WX11033), .ZN(U5828_n1) );
  NOR2X0 U5828_U1 ( .IN1(n5398), .IN2(U5828_n1), .QN(WX11096) );
  INVX0 U5829_U2 ( .INP(WX11031), .ZN(U5829_n1) );
  NOR2X0 U5829_U1 ( .IN1(n5383), .IN2(U5829_n1), .QN(WX11094) );
  INVX0 U5830_U2 ( .INP(WX11029), .ZN(U5830_n1) );
  NOR2X0 U5830_U1 ( .IN1(n5378), .IN2(U5830_n1), .QN(WX11092) );
  INVX0 U5831_U2 ( .INP(WX11027), .ZN(U5831_n1) );
  NOR2X0 U5831_U1 ( .IN1(n5378), .IN2(U5831_n1), .QN(WX11090) );
  INVX0 U5832_U2 ( .INP(WX11025), .ZN(U5832_n1) );
  NOR2X0 U5832_U1 ( .IN1(n5378), .IN2(U5832_n1), .QN(WX11088) );
  INVX0 U5833_U2 ( .INP(WX11023), .ZN(U5833_n1) );
  NOR2X0 U5833_U1 ( .IN1(n5378), .IN2(U5833_n1), .QN(WX11086) );
  INVX0 U5834_U2 ( .INP(WX11021), .ZN(U5834_n1) );
  NOR2X0 U5834_U1 ( .IN1(n5379), .IN2(U5834_n1), .QN(WX11084) );
  INVX0 U5835_U2 ( .INP(WX9886), .ZN(U5835_n1) );
  NOR2X0 U5835_U1 ( .IN1(n5379), .IN2(U5835_n1), .QN(WX9949) );
  INVX0 U5836_U2 ( .INP(WX9884), .ZN(U5836_n1) );
  NOR2X0 U5836_U1 ( .IN1(n5379), .IN2(U5836_n1), .QN(WX9947) );
  INVX0 U5837_U2 ( .INP(WX9882), .ZN(U5837_n1) );
  NOR2X0 U5837_U1 ( .IN1(n5379), .IN2(U5837_n1), .QN(WX9945) );
  INVX0 U5838_U2 ( .INP(WX9880), .ZN(U5838_n1) );
  NOR2X0 U5838_U1 ( .IN1(n5379), .IN2(U5838_n1), .QN(WX9943) );
  INVX0 U5839_U2 ( .INP(WX9878), .ZN(U5839_n1) );
  NOR2X0 U5839_U1 ( .IN1(n5379), .IN2(U5839_n1), .QN(WX9941) );
  INVX0 U5840_U2 ( .INP(WX9876), .ZN(U5840_n1) );
  NOR2X0 U5840_U1 ( .IN1(n5379), .IN2(U5840_n1), .QN(WX9939) );
  INVX0 U5841_U2 ( .INP(WX9874), .ZN(U5841_n1) );
  NOR2X0 U5841_U1 ( .IN1(n5379), .IN2(U5841_n1), .QN(WX9937) );
  INVX0 U5842_U2 ( .INP(WX9872), .ZN(U5842_n1) );
  NOR2X0 U5842_U1 ( .IN1(n5379), .IN2(U5842_n1), .QN(WX9935) );
  INVX0 U5843_U2 ( .INP(WX9870), .ZN(U5843_n1) );
  NOR2X0 U5843_U1 ( .IN1(n5379), .IN2(U5843_n1), .QN(WX9933) );
  INVX0 U5844_U2 ( .INP(WX9868), .ZN(U5844_n1) );
  NOR2X0 U5844_U1 ( .IN1(n5379), .IN2(U5844_n1), .QN(WX9931) );
  INVX0 U5845_U2 ( .INP(WX9866), .ZN(U5845_n1) );
  NOR2X0 U5845_U1 ( .IN1(n5380), .IN2(U5845_n1), .QN(WX9929) );
  INVX0 U5846_U2 ( .INP(WX9864), .ZN(U5846_n1) );
  NOR2X0 U5846_U1 ( .IN1(n5380), .IN2(U5846_n1), .QN(WX9927) );
  INVX0 U5847_U2 ( .INP(WX9862), .ZN(U5847_n1) );
  NOR2X0 U5847_U1 ( .IN1(n5380), .IN2(U5847_n1), .QN(WX9925) );
  INVX0 U5848_U2 ( .INP(WX9860), .ZN(U5848_n1) );
  NOR2X0 U5848_U1 ( .IN1(n5380), .IN2(U5848_n1), .QN(WX9923) );
  INVX0 U5849_U2 ( .INP(WX9858), .ZN(U5849_n1) );
  NOR2X0 U5849_U1 ( .IN1(n5380), .IN2(U5849_n1), .QN(WX9921) );
  INVX0 U5850_U2 ( .INP(WX9856), .ZN(U5850_n1) );
  NOR2X0 U5850_U1 ( .IN1(n5380), .IN2(U5850_n1), .QN(WX9919) );
  INVX0 U5851_U2 ( .INP(test_so84), .ZN(U5851_n1) );
  NOR2X0 U5851_U1 ( .IN1(n5380), .IN2(U5851_n1), .QN(WX9917) );
  INVX0 U5852_U2 ( .INP(WX9852), .ZN(U5852_n1) );
  NOR2X0 U5852_U1 ( .IN1(n5380), .IN2(U5852_n1), .QN(WX9915) );
  INVX0 U5853_U2 ( .INP(WX9850), .ZN(U5853_n1) );
  NOR2X0 U5853_U1 ( .IN1(n5380), .IN2(U5853_n1), .QN(WX9913) );
  INVX0 U5854_U2 ( .INP(WX9848), .ZN(U5854_n1) );
  NOR2X0 U5854_U1 ( .IN1(n5380), .IN2(U5854_n1), .QN(WX9911) );
  INVX0 U5855_U2 ( .INP(WX9846), .ZN(U5855_n1) );
  NOR2X0 U5855_U1 ( .IN1(n5380), .IN2(U5855_n1), .QN(WX9909) );
  INVX0 U5856_U2 ( .INP(WX9844), .ZN(U5856_n1) );
  NOR2X0 U5856_U1 ( .IN1(n5381), .IN2(U5856_n1), .QN(WX9907) );
  INVX0 U5857_U2 ( .INP(WX9842), .ZN(U5857_n1) );
  NOR2X0 U5857_U1 ( .IN1(n5381), .IN2(U5857_n1), .QN(WX9905) );
  INVX0 U5858_U2 ( .INP(WX9840), .ZN(U5858_n1) );
  NOR2X0 U5858_U1 ( .IN1(n5381), .IN2(U5858_n1), .QN(WX9903) );
  INVX0 U5859_U2 ( .INP(WX9838), .ZN(U5859_n1) );
  NOR2X0 U5859_U1 ( .IN1(n5381), .IN2(U5859_n1), .QN(WX9901) );
  INVX0 U5860_U2 ( .INP(WX9836), .ZN(U5860_n1) );
  NOR2X0 U5860_U1 ( .IN1(n5381), .IN2(U5860_n1), .QN(WX9899) );
  INVX0 U5861_U2 ( .INP(WX9834), .ZN(U5861_n1) );
  NOR2X0 U5861_U1 ( .IN1(n5381), .IN2(U5861_n1), .QN(WX9897) );
  INVX0 U5862_U2 ( .INP(WX9832), .ZN(U5862_n1) );
  NOR2X0 U5862_U1 ( .IN1(n5381), .IN2(U5862_n1), .QN(WX9895) );
  INVX0 U5863_U2 ( .INP(WX9830), .ZN(U5863_n1) );
  NOR2X0 U5863_U1 ( .IN1(n5381), .IN2(U5863_n1), .QN(WX9893) );
  INVX0 U5864_U2 ( .INP(WX9828), .ZN(U5864_n1) );
  NOR2X0 U5864_U1 ( .IN1(n5381), .IN2(U5864_n1), .QN(WX9891) );
  INVX0 U5865_U2 ( .INP(WX9826), .ZN(U5865_n1) );
  NOR2X0 U5865_U1 ( .IN1(n5381), .IN2(U5865_n1), .QN(WX9889) );
  INVX0 U5866_U2 ( .INP(WX9824), .ZN(U5866_n1) );
  NOR2X0 U5866_U1 ( .IN1(n5381), .IN2(U5866_n1), .QN(WX9887) );
  INVX0 U5867_U2 ( .INP(WX9822), .ZN(U5867_n1) );
  NOR2X0 U5867_U1 ( .IN1(n5382), .IN2(U5867_n1), .QN(WX9885) );
  INVX0 U5868_U2 ( .INP(test_so83), .ZN(U5868_n1) );
  NOR2X0 U5868_U1 ( .IN1(n5382), .IN2(U5868_n1), .QN(WX9883) );
  INVX0 U5869_U2 ( .INP(WX9818), .ZN(U5869_n1) );
  NOR2X0 U5869_U1 ( .IN1(n5382), .IN2(U5869_n1), .QN(WX9881) );
  INVX0 U5870_U2 ( .INP(WX9816), .ZN(U5870_n1) );
  NOR2X0 U5870_U1 ( .IN1(n5382), .IN2(U5870_n1), .QN(WX9879) );
  INVX0 U5871_U2 ( .INP(WX9814), .ZN(U5871_n1) );
  NOR2X0 U5871_U1 ( .IN1(n5382), .IN2(U5871_n1), .QN(WX9877) );
  INVX0 U5872_U2 ( .INP(WX9812), .ZN(U5872_n1) );
  NOR2X0 U5872_U1 ( .IN1(n5382), .IN2(U5872_n1), .QN(WX9875) );
  INVX0 U5873_U2 ( .INP(WX9810), .ZN(U5873_n1) );
  NOR2X0 U5873_U1 ( .IN1(n5382), .IN2(U5873_n1), .QN(WX9873) );
  INVX0 U5874_U2 ( .INP(WX9808), .ZN(U5874_n1) );
  NOR2X0 U5874_U1 ( .IN1(n5382), .IN2(U5874_n1), .QN(WX9871) );
  INVX0 U5875_U2 ( .INP(WX9806), .ZN(U5875_n1) );
  NOR2X0 U5875_U1 ( .IN1(n5382), .IN2(U5875_n1), .QN(WX9869) );
  INVX0 U5876_U2 ( .INP(WX9804), .ZN(U5876_n1) );
  NOR2X0 U5876_U1 ( .IN1(n5382), .IN2(U5876_n1), .QN(WX9867) );
  INVX0 U5877_U2 ( .INP(WX9802), .ZN(U5877_n1) );
  NOR2X0 U5877_U1 ( .IN1(n5382), .IN2(U5877_n1), .QN(WX9865) );
  INVX0 U5878_U2 ( .INP(WX9800), .ZN(U5878_n1) );
  NOR2X0 U5878_U1 ( .IN1(n5383), .IN2(U5878_n1), .QN(WX9863) );
  INVX0 U5879_U2 ( .INP(WX9798), .ZN(U5879_n1) );
  NOR2X0 U5879_U1 ( .IN1(n5383), .IN2(U5879_n1), .QN(WX9861) );
  INVX0 U5880_U2 ( .INP(WX9796), .ZN(U5880_n1) );
  NOR2X0 U5880_U1 ( .IN1(n5383), .IN2(U5880_n1), .QN(WX9859) );
  INVX0 U5881_U2 ( .INP(WX9794), .ZN(U5881_n1) );
  NOR2X0 U5881_U1 ( .IN1(n5383), .IN2(U5881_n1), .QN(WX9857) );
  INVX0 U5882_U2 ( .INP(WX9792), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(n5383), .IN2(U5882_n1), .QN(WX9855) );
  INVX0 U5883_U2 ( .INP(WX9790), .ZN(U5883_n1) );
  NOR2X0 U5883_U1 ( .IN1(n5383), .IN2(U5883_n1), .QN(WX9853) );
  INVX0 U5884_U2 ( .INP(WX9788), .ZN(U5884_n1) );
  NOR2X0 U5884_U1 ( .IN1(n5383), .IN2(U5884_n1), .QN(WX9851) );
  INVX0 U5885_U2 ( .INP(test_so82), .ZN(U5885_n1) );
  NOR2X0 U5885_U1 ( .IN1(n5383), .IN2(U5885_n1), .QN(WX9849) );
  INVX0 U5886_U2 ( .INP(WX9784), .ZN(U5886_n1) );
  NOR2X0 U5886_U1 ( .IN1(n5383), .IN2(U5886_n1), .QN(WX9847) );
  INVX0 U5887_U2 ( .INP(WX9782), .ZN(U5887_n1) );
  NOR2X0 U5887_U1 ( .IN1(n5383), .IN2(U5887_n1), .QN(WX9845) );
  INVX0 U5888_U2 ( .INP(WX9780), .ZN(U5888_n1) );
  NOR2X0 U5888_U1 ( .IN1(n5384), .IN2(U5888_n1), .QN(WX9843) );
  INVX0 U5889_U2 ( .INP(WX9778), .ZN(U5889_n1) );
  NOR2X0 U5889_U1 ( .IN1(n5384), .IN2(U5889_n1), .QN(WX9841) );
  INVX0 U5890_U2 ( .INP(WX9776), .ZN(U5890_n1) );
  NOR2X0 U5890_U1 ( .IN1(n5384), .IN2(U5890_n1), .QN(WX9839) );
  INVX0 U5891_U2 ( .INP(WX9774), .ZN(U5891_n1) );
  NOR2X0 U5891_U1 ( .IN1(n5384), .IN2(U5891_n1), .QN(WX9837) );
  INVX0 U5892_U2 ( .INP(WX9772), .ZN(U5892_n1) );
  NOR2X0 U5892_U1 ( .IN1(n5384), .IN2(U5892_n1), .QN(WX9835) );
  INVX0 U5893_U2 ( .INP(WX9770), .ZN(U5893_n1) );
  NOR2X0 U5893_U1 ( .IN1(n5384), .IN2(U5893_n1), .QN(WX9833) );
  INVX0 U5894_U2 ( .INP(WX9768), .ZN(U5894_n1) );
  NOR2X0 U5894_U1 ( .IN1(n5384), .IN2(U5894_n1), .QN(WX9831) );
  INVX0 U5895_U2 ( .INP(WX9766), .ZN(U5895_n1) );
  NOR2X0 U5895_U1 ( .IN1(n5384), .IN2(U5895_n1), .QN(WX9829) );
  INVX0 U5896_U2 ( .INP(WX9764), .ZN(U5896_n1) );
  NOR2X0 U5896_U1 ( .IN1(n5384), .IN2(U5896_n1), .QN(WX9827) );
  INVX0 U5897_U2 ( .INP(WX9762), .ZN(U5897_n1) );
  NOR2X0 U5897_U1 ( .IN1(n5384), .IN2(U5897_n1), .QN(WX9825) );
  INVX0 U5898_U2 ( .INP(WX9760), .ZN(U5898_n1) );
  NOR2X0 U5898_U1 ( .IN1(n5384), .IN2(U5898_n1), .QN(WX9823) );
  INVX0 U5899_U2 ( .INP(WX9758), .ZN(U5899_n1) );
  NOR2X0 U5899_U1 ( .IN1(n5385), .IN2(U5899_n1), .QN(WX9821) );
  INVX0 U5900_U2 ( .INP(WX9756), .ZN(U5900_n1) );
  NOR2X0 U5900_U1 ( .IN1(n5385), .IN2(U5900_n1), .QN(WX9819) );
  INVX0 U5901_U2 ( .INP(WX9754), .ZN(U5901_n1) );
  NOR2X0 U5901_U1 ( .IN1(n5385), .IN2(U5901_n1), .QN(WX9817) );
  INVX0 U5902_U2 ( .INP(test_so81), .ZN(U5902_n1) );
  NOR2X0 U5902_U1 ( .IN1(n5385), .IN2(U5902_n1), .QN(WX9815) );
  INVX0 U5903_U2 ( .INP(WX9750), .ZN(U5903_n1) );
  NOR2X0 U5903_U1 ( .IN1(n5385), .IN2(U5903_n1), .QN(WX9813) );
  INVX0 U5904_U2 ( .INP(WX9748), .ZN(U5904_n1) );
  NOR2X0 U5904_U1 ( .IN1(n5385), .IN2(U5904_n1), .QN(WX9811) );
  INVX0 U5905_U2 ( .INP(WX9746), .ZN(U5905_n1) );
  NOR2X0 U5905_U1 ( .IN1(n5385), .IN2(U5905_n1), .QN(WX9809) );
  INVX0 U5906_U2 ( .INP(WX9744), .ZN(U5906_n1) );
  NOR2X0 U5906_U1 ( .IN1(n5385), .IN2(U5906_n1), .QN(WX9807) );
  INVX0 U5907_U2 ( .INP(WX9742), .ZN(U5907_n1) );
  NOR2X0 U5907_U1 ( .IN1(n5385), .IN2(U5907_n1), .QN(WX9805) );
  INVX0 U5908_U2 ( .INP(WX9740), .ZN(U5908_n1) );
  NOR2X0 U5908_U1 ( .IN1(n5385), .IN2(U5908_n1), .QN(WX9803) );
  INVX0 U5909_U2 ( .INP(WX9738), .ZN(U5909_n1) );
  NOR2X0 U5909_U1 ( .IN1(n5385), .IN2(U5909_n1), .QN(WX9801) );
  INVX0 U5910_U2 ( .INP(WX9736), .ZN(U5910_n1) );
  NOR2X0 U5910_U1 ( .IN1(n5386), .IN2(U5910_n1), .QN(WX9799) );
  INVX0 U5911_U2 ( .INP(WX9734), .ZN(U5911_n1) );
  NOR2X0 U5911_U1 ( .IN1(n5386), .IN2(U5911_n1), .QN(WX9797) );
  INVX0 U5912_U2 ( .INP(WX9732), .ZN(U5912_n1) );
  NOR2X0 U5912_U1 ( .IN1(n5386), .IN2(U5912_n1), .QN(WX9795) );
  INVX0 U5913_U2 ( .INP(WX9730), .ZN(U5913_n1) );
  NOR2X0 U5913_U1 ( .IN1(n5386), .IN2(U5913_n1), .QN(WX9793) );
  INVX0 U5914_U2 ( .INP(WX9728), .ZN(U5914_n1) );
  NOR2X0 U5914_U1 ( .IN1(n5386), .IN2(U5914_n1), .QN(WX9791) );
  INVX0 U5915_U2 ( .INP(WX8593), .ZN(U5915_n1) );
  NOR2X0 U5915_U1 ( .IN1(n5386), .IN2(U5915_n1), .QN(WX8656) );
  INVX0 U5916_U2 ( .INP(WX8591), .ZN(U5916_n1) );
  NOR2X0 U5916_U1 ( .IN1(n5386), .IN2(U5916_n1), .QN(WX8654) );
  INVX0 U5917_U2 ( .INP(WX8589), .ZN(U5917_n1) );
  NOR2X0 U5917_U1 ( .IN1(n5386), .IN2(U5917_n1), .QN(WX8652) );
  INVX0 U5918_U2 ( .INP(WX8587), .ZN(U5918_n1) );
  NOR2X0 U5918_U1 ( .IN1(n5386), .IN2(U5918_n1), .QN(WX8650) );
  INVX0 U5919_U2 ( .INP(WX8585), .ZN(U5919_n1) );
  NOR2X0 U5919_U1 ( .IN1(n5386), .IN2(U5919_n1), .QN(WX8648) );
  INVX0 U5920_U2 ( .INP(WX8583), .ZN(U5920_n1) );
  NOR2X0 U5920_U1 ( .IN1(n5386), .IN2(U5920_n1), .QN(WX8646) );
  INVX0 U5921_U2 ( .INP(WX8581), .ZN(U5921_n1) );
  NOR2X0 U5921_U1 ( .IN1(n5387), .IN2(U5921_n1), .QN(WX8644) );
  INVX0 U5922_U2 ( .INP(WX8579), .ZN(U5922_n1) );
  NOR2X0 U5922_U1 ( .IN1(n5387), .IN2(U5922_n1), .QN(WX8642) );
  INVX0 U5923_U2 ( .INP(WX8577), .ZN(U5923_n1) );
  NOR2X0 U5923_U1 ( .IN1(n5387), .IN2(U5923_n1), .QN(WX8640) );
  INVX0 U5924_U2 ( .INP(WX8575), .ZN(U5924_n1) );
  NOR2X0 U5924_U1 ( .IN1(n5387), .IN2(U5924_n1), .QN(WX8638) );
  INVX0 U5925_U2 ( .INP(WX8573), .ZN(U5925_n1) );
  NOR2X0 U5925_U1 ( .IN1(n5387), .IN2(U5925_n1), .QN(WX8636) );
  INVX0 U5926_U2 ( .INP(test_so73), .ZN(U5926_n1) );
  NOR2X0 U5926_U1 ( .IN1(n5387), .IN2(U5926_n1), .QN(WX8634) );
  INVX0 U5927_U2 ( .INP(WX8569), .ZN(U5927_n1) );
  NOR2X0 U5927_U1 ( .IN1(n5387), .IN2(U5927_n1), .QN(WX8632) );
  INVX0 U5928_U2 ( .INP(WX8567), .ZN(U5928_n1) );
  NOR2X0 U5928_U1 ( .IN1(n5387), .IN2(U5928_n1), .QN(WX8630) );
  INVX0 U5929_U2 ( .INP(WX8565), .ZN(U5929_n1) );
  NOR2X0 U5929_U1 ( .IN1(n5387), .IN2(U5929_n1), .QN(WX8628) );
  INVX0 U5930_U2 ( .INP(WX8563), .ZN(U5930_n1) );
  NOR2X0 U5930_U1 ( .IN1(n5387), .IN2(U5930_n1), .QN(WX8626) );
  INVX0 U5931_U2 ( .INP(WX8561), .ZN(U5931_n1) );
  NOR2X0 U5931_U1 ( .IN1(n5387), .IN2(U5931_n1), .QN(WX8624) );
  INVX0 U5932_U2 ( .INP(WX8559), .ZN(U5932_n1) );
  NOR2X0 U5932_U1 ( .IN1(n5388), .IN2(U5932_n1), .QN(WX8622) );
  INVX0 U5933_U2 ( .INP(WX8557), .ZN(U5933_n1) );
  NOR2X0 U5933_U1 ( .IN1(n5388), .IN2(U5933_n1), .QN(WX8620) );
  INVX0 U5934_U2 ( .INP(WX8555), .ZN(U5934_n1) );
  NOR2X0 U5934_U1 ( .IN1(n5388), .IN2(U5934_n1), .QN(WX8618) );
  INVX0 U5935_U2 ( .INP(WX8553), .ZN(U5935_n1) );
  NOR2X0 U5935_U1 ( .IN1(n5388), .IN2(U5935_n1), .QN(WX8616) );
  INVX0 U5936_U2 ( .INP(WX8551), .ZN(U5936_n1) );
  NOR2X0 U5936_U1 ( .IN1(n5388), .IN2(U5936_n1), .QN(WX8614) );
  INVX0 U5937_U2 ( .INP(WX8549), .ZN(U5937_n1) );
  NOR2X0 U5937_U1 ( .IN1(n5388), .IN2(U5937_n1), .QN(WX8612) );
  INVX0 U5938_U2 ( .INP(WX8547), .ZN(U5938_n1) );
  NOR2X0 U5938_U1 ( .IN1(n5388), .IN2(U5938_n1), .QN(WX8610) );
  INVX0 U5939_U2 ( .INP(WX8545), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n5388), .IN2(U5939_n1), .QN(WX8608) );
  INVX0 U5940_U2 ( .INP(WX8543), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n5411), .IN2(U5940_n1), .QN(WX8606) );
  INVX0 U5941_U2 ( .INP(WX8541), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n5418), .IN2(U5941_n1), .QN(WX8604) );
  INVX0 U5942_U2 ( .INP(WX8539), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n5417), .IN2(U5942_n1), .QN(WX8602) );
  INVX0 U5943_U2 ( .INP(test_so72), .ZN(U5943_n1) );
  NOR2X0 U5943_U1 ( .IN1(n5418), .IN2(U5943_n1), .QN(WX8600) );
  INVX0 U5944_U2 ( .INP(WX8535), .ZN(U5944_n1) );
  NOR2X0 U5944_U1 ( .IN1(n5418), .IN2(U5944_n1), .QN(WX8598) );
  INVX0 U5945_U2 ( .INP(WX8533), .ZN(U5945_n1) );
  NOR2X0 U5945_U1 ( .IN1(n5418), .IN2(U5945_n1), .QN(WX8596) );
  INVX0 U5946_U2 ( .INP(WX8531), .ZN(U5946_n1) );
  NOR2X0 U5946_U1 ( .IN1(n5418), .IN2(U5946_n1), .QN(WX8594) );
  INVX0 U5947_U2 ( .INP(WX8529), .ZN(U5947_n1) );
  NOR2X0 U5947_U1 ( .IN1(n5417), .IN2(U5947_n1), .QN(WX8592) );
  INVX0 U5948_U2 ( .INP(WX8527), .ZN(U5948_n1) );
  NOR2X0 U5948_U1 ( .IN1(n5417), .IN2(U5948_n1), .QN(WX8590) );
  INVX0 U5949_U2 ( .INP(WX8525), .ZN(U5949_n1) );
  NOR2X0 U5949_U1 ( .IN1(n5418), .IN2(U5949_n1), .QN(WX8588) );
  INVX0 U5950_U2 ( .INP(WX8523), .ZN(U5950_n1) );
  NOR2X0 U5950_U1 ( .IN1(n5416), .IN2(U5950_n1), .QN(WX8586) );
  INVX0 U5951_U2 ( .INP(WX8521), .ZN(U5951_n1) );
  NOR2X0 U5951_U1 ( .IN1(n5417), .IN2(U5951_n1), .QN(WX8584) );
  INVX0 U5952_U2 ( .INP(WX8519), .ZN(U5952_n1) );
  NOR2X0 U5952_U1 ( .IN1(n5418), .IN2(U5952_n1), .QN(WX8582) );
  INVX0 U5953_U2 ( .INP(WX8517), .ZN(U5953_n1) );
  NOR2X0 U5953_U1 ( .IN1(n5418), .IN2(U5953_n1), .QN(WX8580) );
  INVX0 U5954_U2 ( .INP(WX8515), .ZN(U5954_n1) );
  NOR2X0 U5954_U1 ( .IN1(n5417), .IN2(U5954_n1), .QN(WX8578) );
  INVX0 U5955_U2 ( .INP(WX8513), .ZN(U5955_n1) );
  NOR2X0 U5955_U1 ( .IN1(n5414), .IN2(U5955_n1), .QN(WX8576) );
  INVX0 U5956_U2 ( .INP(WX8511), .ZN(U5956_n1) );
  NOR2X0 U5956_U1 ( .IN1(n5414), .IN2(U5956_n1), .QN(WX8574) );
  INVX0 U5957_U2 ( .INP(WX8509), .ZN(U5957_n1) );
  NOR2X0 U5957_U1 ( .IN1(n5414), .IN2(U5957_n1), .QN(WX8572) );
  INVX0 U5958_U2 ( .INP(WX8507), .ZN(U5958_n1) );
  NOR2X0 U5958_U1 ( .IN1(n5414), .IN2(U5958_n1), .QN(WX8570) );
  INVX0 U5959_U2 ( .INP(WX8505), .ZN(U5959_n1) );
  NOR2X0 U5959_U1 ( .IN1(n5414), .IN2(U5959_n1), .QN(WX8568) );
  INVX0 U5960_U2 ( .INP(test_so71), .ZN(U5960_n1) );
  NOR2X0 U5960_U1 ( .IN1(n5414), .IN2(U5960_n1), .QN(WX8566) );
  INVX0 U5961_U2 ( .INP(WX8501), .ZN(U5961_n1) );
  NOR2X0 U5961_U1 ( .IN1(n5414), .IN2(U5961_n1), .QN(WX8564) );
  INVX0 U5962_U2 ( .INP(WX8499), .ZN(U5962_n1) );
  NOR2X0 U5962_U1 ( .IN1(n5413), .IN2(U5962_n1), .QN(WX8562) );
  INVX0 U5963_U2 ( .INP(WX8497), .ZN(U5963_n1) );
  NOR2X0 U5963_U1 ( .IN1(n5412), .IN2(U5963_n1), .QN(WX8560) );
  INVX0 U5964_U2 ( .INP(WX8495), .ZN(U5964_n1) );
  NOR2X0 U5964_U1 ( .IN1(n5412), .IN2(U5964_n1), .QN(WX8558) );
  INVX0 U5965_U2 ( .INP(WX8493), .ZN(U5965_n1) );
  NOR2X0 U5965_U1 ( .IN1(n5412), .IN2(U5965_n1), .QN(WX8556) );
  INVX0 U5966_U2 ( .INP(WX8491), .ZN(U5966_n1) );
  NOR2X0 U5966_U1 ( .IN1(n5412), .IN2(U5966_n1), .QN(WX8554) );
  INVX0 U5967_U2 ( .INP(WX8489), .ZN(U5967_n1) );
  NOR2X0 U5967_U1 ( .IN1(n5412), .IN2(U5967_n1), .QN(WX8552) );
  INVX0 U5968_U2 ( .INP(WX8487), .ZN(U5968_n1) );
  NOR2X0 U5968_U1 ( .IN1(n5412), .IN2(U5968_n1), .QN(WX8550) );
  INVX0 U5969_U2 ( .INP(WX8485), .ZN(U5969_n1) );
  NOR2X0 U5969_U1 ( .IN1(n5411), .IN2(U5969_n1), .QN(WX8548) );
  INVX0 U5970_U2 ( .INP(WX8483), .ZN(U5970_n1) );
  NOR2X0 U5970_U1 ( .IN1(n5411), .IN2(U5970_n1), .QN(WX8546) );
  INVX0 U5971_U2 ( .INP(WX8481), .ZN(U5971_n1) );
  NOR2X0 U5971_U1 ( .IN1(n5411), .IN2(U5971_n1), .QN(WX8544) );
  INVX0 U5972_U2 ( .INP(WX8479), .ZN(U5972_n1) );
  NOR2X0 U5972_U1 ( .IN1(n5411), .IN2(U5972_n1), .QN(WX8542) );
  INVX0 U5973_U2 ( .INP(WX8477), .ZN(U5973_n1) );
  NOR2X0 U5973_U1 ( .IN1(n5411), .IN2(U5973_n1), .QN(WX8540) );
  INVX0 U5974_U2 ( .INP(WX8475), .ZN(U5974_n1) );
  NOR2X0 U5974_U1 ( .IN1(n5411), .IN2(U5974_n1), .QN(WX8538) );
  INVX0 U5975_U2 ( .INP(WX8473), .ZN(U5975_n1) );
  NOR2X0 U5975_U1 ( .IN1(n5411), .IN2(U5975_n1), .QN(WX8536) );
  INVX0 U5976_U2 ( .INP(WX8471), .ZN(U5976_n1) );
  NOR2X0 U5976_U1 ( .IN1(n5411), .IN2(U5976_n1), .QN(WX8534) );
  INVX0 U5977_U2 ( .INP(test_so70), .ZN(U5977_n1) );
  NOR2X0 U5977_U1 ( .IN1(n5411), .IN2(U5977_n1), .QN(WX8532) );
  INVX0 U5978_U2 ( .INP(WX8467), .ZN(U5978_n1) );
  NOR2X0 U5978_U1 ( .IN1(n5411), .IN2(U5978_n1), .QN(WX8530) );
  INVX0 U5979_U2 ( .INP(WX8465), .ZN(U5979_n1) );
  NOR2X0 U5979_U1 ( .IN1(n5410), .IN2(U5979_n1), .QN(WX8528) );
  INVX0 U5980_U2 ( .INP(WX8463), .ZN(U5980_n1) );
  NOR2X0 U5980_U1 ( .IN1(n5410), .IN2(U5980_n1), .QN(WX8526) );
  INVX0 U5981_U2 ( .INP(WX8461), .ZN(U5981_n1) );
  NOR2X0 U5981_U1 ( .IN1(n5410), .IN2(U5981_n1), .QN(WX8524) );
  INVX0 U5982_U2 ( .INP(WX8459), .ZN(U5982_n1) );
  NOR2X0 U5982_U1 ( .IN1(n5410), .IN2(U5982_n1), .QN(WX8522) );
  INVX0 U5983_U2 ( .INP(WX8457), .ZN(U5983_n1) );
  NOR2X0 U5983_U1 ( .IN1(n5410), .IN2(U5983_n1), .QN(WX8520) );
  INVX0 U5984_U2 ( .INP(WX8455), .ZN(U5984_n1) );
  NOR2X0 U5984_U1 ( .IN1(n5410), .IN2(U5984_n1), .QN(WX8518) );
  INVX0 U5985_U2 ( .INP(WX8453), .ZN(U5985_n1) );
  NOR2X0 U5985_U1 ( .IN1(n5410), .IN2(U5985_n1), .QN(WX8516) );
  INVX0 U5986_U2 ( .INP(WX8451), .ZN(U5986_n1) );
  NOR2X0 U5986_U1 ( .IN1(n5409), .IN2(U5986_n1), .QN(WX8514) );
  INVX0 U5987_U2 ( .INP(WX8449), .ZN(U5987_n1) );
  NOR2X0 U5987_U1 ( .IN1(n5409), .IN2(U5987_n1), .QN(WX8512) );
  INVX0 U5988_U2 ( .INP(WX8447), .ZN(U5988_n1) );
  NOR2X0 U5988_U1 ( .IN1(n5409), .IN2(U5988_n1), .QN(WX8510) );
  INVX0 U5989_U2 ( .INP(WX8445), .ZN(U5989_n1) );
  NOR2X0 U5989_U1 ( .IN1(n5409), .IN2(U5989_n1), .QN(WX8508) );
  INVX0 U5990_U2 ( .INP(WX8443), .ZN(U5990_n1) );
  NOR2X0 U5990_U1 ( .IN1(n5409), .IN2(U5990_n1), .QN(WX8506) );
  INVX0 U5991_U2 ( .INP(WX8441), .ZN(U5991_n1) );
  NOR2X0 U5991_U1 ( .IN1(n5409), .IN2(U5991_n1), .QN(WX8504) );
  INVX0 U5992_U2 ( .INP(WX8439), .ZN(U5992_n1) );
  NOR2X0 U5992_U1 ( .IN1(n5409), .IN2(U5992_n1), .QN(WX8502) );
  INVX0 U5993_U2 ( .INP(WX8437), .ZN(U5993_n1) );
  NOR2X0 U5993_U1 ( .IN1(n5409), .IN2(U5993_n1), .QN(WX8500) );
  INVX0 U5994_U2 ( .INP(test_so69), .ZN(U5994_n1) );
  NOR2X0 U5994_U1 ( .IN1(n5409), .IN2(U5994_n1), .QN(WX8498) );
  INVX0 U5995_U2 ( .INP(WX7300), .ZN(U5995_n1) );
  NOR2X0 U5995_U1 ( .IN1(n5409), .IN2(U5995_n1), .QN(WX7363) );
  INVX0 U5996_U2 ( .INP(WX7298), .ZN(U5996_n1) );
  NOR2X0 U5996_U1 ( .IN1(n5409), .IN2(U5996_n1), .QN(WX7361) );
  INVX0 U5997_U2 ( .INP(WX7296), .ZN(U5997_n1) );
  NOR2X0 U5997_U1 ( .IN1(n5410), .IN2(U5997_n1), .QN(WX7359) );
  INVX0 U5998_U2 ( .INP(WX7294), .ZN(U5998_n1) );
  NOR2X0 U5998_U1 ( .IN1(n5410), .IN2(U5998_n1), .QN(WX7357) );
  INVX0 U5999_U2 ( .INP(WX7292), .ZN(U5999_n1) );
  NOR2X0 U5999_U1 ( .IN1(n5410), .IN2(U5999_n1), .QN(WX7355) );
  INVX0 U6000_U2 ( .INP(WX7290), .ZN(U6000_n1) );
  NOR2X0 U6000_U1 ( .IN1(n5410), .IN2(U6000_n1), .QN(WX7353) );
  INVX0 U6001_U2 ( .INP(test_so62), .ZN(U6001_n1) );
  NOR2X0 U6001_U1 ( .IN1(n5412), .IN2(U6001_n1), .QN(WX7351) );
  INVX0 U6002_U2 ( .INP(WX7286), .ZN(U6002_n1) );
  NOR2X0 U6002_U1 ( .IN1(n5412), .IN2(U6002_n1), .QN(WX7349) );
  INVX0 U6003_U2 ( .INP(WX7284), .ZN(U6003_n1) );
  NOR2X0 U6003_U1 ( .IN1(n5412), .IN2(U6003_n1), .QN(WX7347) );
  INVX0 U6004_U2 ( .INP(WX7282), .ZN(U6004_n1) );
  NOR2X0 U6004_U1 ( .IN1(n5412), .IN2(U6004_n1), .QN(WX7345) );
  INVX0 U6005_U2 ( .INP(WX7280), .ZN(U6005_n1) );
  NOR2X0 U6005_U1 ( .IN1(n5412), .IN2(U6005_n1), .QN(WX7343) );
  INVX0 U6006_U2 ( .INP(WX7278), .ZN(U6006_n1) );
  NOR2X0 U6006_U1 ( .IN1(n5413), .IN2(U6006_n1), .QN(WX7341) );
  INVX0 U6007_U2 ( .INP(WX7276), .ZN(U6007_n1) );
  NOR2X0 U6007_U1 ( .IN1(n5413), .IN2(U6007_n1), .QN(WX7339) );
  INVX0 U6008_U2 ( .INP(WX7274), .ZN(U6008_n1) );
  NOR2X0 U6008_U1 ( .IN1(n5413), .IN2(U6008_n1), .QN(WX7337) );
  INVX0 U6009_U2 ( .INP(WX7272), .ZN(U6009_n1) );
  NOR2X0 U6009_U1 ( .IN1(n5413), .IN2(U6009_n1), .QN(WX7335) );
  INVX0 U6010_U2 ( .INP(WX7270), .ZN(U6010_n1) );
  NOR2X0 U6010_U1 ( .IN1(n5413), .IN2(U6010_n1), .QN(WX7333) );
  INVX0 U6011_U2 ( .INP(WX7268), .ZN(U6011_n1) );
  NOR2X0 U6011_U1 ( .IN1(n5413), .IN2(U6011_n1), .QN(WX7331) );
  INVX0 U6012_U2 ( .INP(WX7266), .ZN(U6012_n1) );
  NOR2X0 U6012_U1 ( .IN1(n5413), .IN2(U6012_n1), .QN(WX7329) );
  INVX0 U6013_U2 ( .INP(WX7264), .ZN(U6013_n1) );
  NOR2X0 U6013_U1 ( .IN1(n5413), .IN2(U6013_n1), .QN(WX7327) );
  INVX0 U6014_U2 ( .INP(WX7262), .ZN(U6014_n1) );
  NOR2X0 U6014_U1 ( .IN1(n5413), .IN2(U6014_n1), .QN(WX7325) );
  INVX0 U6015_U2 ( .INP(WX7260), .ZN(U6015_n1) );
  NOR2X0 U6015_U1 ( .IN1(n5413), .IN2(U6015_n1), .QN(WX7323) );
  INVX0 U6016_U2 ( .INP(WX7258), .ZN(U6016_n1) );
  NOR2X0 U6016_U1 ( .IN1(n5414), .IN2(U6016_n1), .QN(WX7321) );
  INVX0 U6017_U2 ( .INP(WX7256), .ZN(U6017_n1) );
  NOR2X0 U6017_U1 ( .IN1(n5414), .IN2(U6017_n1), .QN(WX7319) );
  INVX0 U6018_U2 ( .INP(test_so61), .ZN(U6018_n1) );
  NOR2X0 U6018_U1 ( .IN1(n5414), .IN2(U6018_n1), .QN(WX7317) );
  INVX0 U6019_U2 ( .INP(WX7252), .ZN(U6019_n1) );
  NOR2X0 U6019_U1 ( .IN1(n5415), .IN2(U6019_n1), .QN(WX7315) );
  INVX0 U6020_U2 ( .INP(WX7250), .ZN(U6020_n1) );
  NOR2X0 U6020_U1 ( .IN1(n5415), .IN2(U6020_n1), .QN(WX7313) );
  INVX0 U6021_U2 ( .INP(WX7248), .ZN(U6021_n1) );
  NOR2X0 U6021_U1 ( .IN1(n5415), .IN2(U6021_n1), .QN(WX7311) );
  INVX0 U6022_U2 ( .INP(WX7246), .ZN(U6022_n1) );
  NOR2X0 U6022_U1 ( .IN1(n5415), .IN2(U6022_n1), .QN(WX7309) );
  INVX0 U6023_U2 ( .INP(WX7244), .ZN(U6023_n1) );
  NOR2X0 U6023_U1 ( .IN1(n5415), .IN2(U6023_n1), .QN(WX7307) );
  INVX0 U6024_U2 ( .INP(WX7242), .ZN(U6024_n1) );
  NOR2X0 U6024_U1 ( .IN1(n5415), .IN2(U6024_n1), .QN(WX7305) );
  INVX0 U6025_U2 ( .INP(WX7240), .ZN(U6025_n1) );
  NOR2X0 U6025_U1 ( .IN1(n5416), .IN2(U6025_n1), .QN(WX7303) );
  INVX0 U6026_U2 ( .INP(WX7238), .ZN(U6026_n1) );
  NOR2X0 U6026_U1 ( .IN1(n5416), .IN2(U6026_n1), .QN(WX7301) );
  INVX0 U6027_U2 ( .INP(WX7236), .ZN(U6027_n1) );
  NOR2X0 U6027_U1 ( .IN1(n5415), .IN2(U6027_n1), .QN(WX7299) );
  INVX0 U6028_U2 ( .INP(WX7234), .ZN(U6028_n1) );
  NOR2X0 U6028_U1 ( .IN1(n5416), .IN2(U6028_n1), .QN(WX7297) );
  INVX0 U6029_U2 ( .INP(WX7232), .ZN(U6029_n1) );
  NOR2X0 U6029_U1 ( .IN1(n5416), .IN2(U6029_n1), .QN(WX7295) );
  INVX0 U6030_U2 ( .INP(WX7230), .ZN(U6030_n1) );
  NOR2X0 U6030_U1 ( .IN1(n5415), .IN2(U6030_n1), .QN(WX7293) );
  INVX0 U6031_U2 ( .INP(WX7228), .ZN(U6031_n1) );
  NOR2X0 U6031_U1 ( .IN1(n5416), .IN2(U6031_n1), .QN(WX7291) );
  INVX0 U6032_U2 ( .INP(WX7226), .ZN(U6032_n1) );
  NOR2X0 U6032_U1 ( .IN1(n5415), .IN2(U6032_n1), .QN(WX7289) );
  INVX0 U6033_U2 ( .INP(WX7224), .ZN(U6033_n1) );
  NOR2X0 U6033_U1 ( .IN1(n5415), .IN2(U6033_n1), .QN(WX7287) );
  INVX0 U6034_U2 ( .INP(WX7222), .ZN(U6034_n1) );
  NOR2X0 U6034_U1 ( .IN1(n5416), .IN2(U6034_n1), .QN(WX7285) );
  INVX0 U6035_U2 ( .INP(test_so60), .ZN(U6035_n1) );
  NOR2X0 U6035_U1 ( .IN1(n5416), .IN2(U6035_n1), .QN(WX7283) );
  INVX0 U6036_U2 ( .INP(WX7218), .ZN(U6036_n1) );
  NOR2X0 U6036_U1 ( .IN1(n5416), .IN2(U6036_n1), .QN(WX7281) );
  INVX0 U6037_U2 ( .INP(WX7216), .ZN(U6037_n1) );
  NOR2X0 U6037_U1 ( .IN1(n5417), .IN2(U6037_n1), .QN(WX7279) );
  INVX0 U6038_U2 ( .INP(WX7214), .ZN(U6038_n1) );
  NOR2X0 U6038_U1 ( .IN1(n5417), .IN2(U6038_n1), .QN(WX7277) );
  INVX0 U6039_U2 ( .INP(WX7212), .ZN(U6039_n1) );
  NOR2X0 U6039_U1 ( .IN1(n5416), .IN2(U6039_n1), .QN(WX7275) );
  INVX0 U6040_U2 ( .INP(WX7210), .ZN(U6040_n1) );
  NOR2X0 U6040_U1 ( .IN1(n5416), .IN2(U6040_n1), .QN(WX7273) );
  INVX0 U6041_U2 ( .INP(WX7208), .ZN(U6041_n1) );
  NOR2X0 U6041_U1 ( .IN1(n5417), .IN2(U6041_n1), .QN(WX7271) );
  INVX0 U6042_U2 ( .INP(WX7206), .ZN(U6042_n1) );
  NOR2X0 U6042_U1 ( .IN1(n5415), .IN2(U6042_n1), .QN(WX7269) );
  INVX0 U6043_U2 ( .INP(WX7204), .ZN(U6043_n1) );
  NOR2X0 U6043_U1 ( .IN1(n5417), .IN2(U6043_n1), .QN(WX7267) );
  INVX0 U6044_U2 ( .INP(WX7202), .ZN(U6044_n1) );
  NOR2X0 U6044_U1 ( .IN1(n5417), .IN2(U6044_n1), .QN(WX7265) );
  INVX0 U6045_U2 ( .INP(WX7200), .ZN(U6045_n1) );
  NOR2X0 U6045_U1 ( .IN1(n5417), .IN2(U6045_n1), .QN(WX7263) );
  INVX0 U6046_U2 ( .INP(WX7198), .ZN(U6046_n1) );
  NOR2X0 U6046_U1 ( .IN1(n5418), .IN2(U6046_n1), .QN(WX7261) );
  INVX0 U6047_U2 ( .INP(WX7196), .ZN(U6047_n1) );
  NOR2X0 U6047_U1 ( .IN1(n5418), .IN2(U6047_n1), .QN(WX7259) );
  INVX0 U6048_U2 ( .INP(WX7194), .ZN(U6048_n1) );
  NOR2X0 U6048_U1 ( .IN1(n5419), .IN2(U6048_n1), .QN(WX7257) );
  INVX0 U6049_U2 ( .INP(WX7192), .ZN(U6049_n1) );
  NOR2X0 U6049_U1 ( .IN1(n5418), .IN2(U6049_n1), .QN(WX7255) );
  INVX0 U6050_U2 ( .INP(WX7190), .ZN(U6050_n1) );
  NOR2X0 U6050_U1 ( .IN1(n5403), .IN2(U6050_n1), .QN(WX7253) );
  INVX0 U6051_U2 ( .INP(WX7188), .ZN(U6051_n1) );
  NOR2X0 U6051_U1 ( .IN1(n5398), .IN2(U6051_n1), .QN(WX7251) );
  INVX0 U6052_U2 ( .INP(test_so59), .ZN(U6052_n1) );
  NOR2X0 U6052_U1 ( .IN1(n5399), .IN2(U6052_n1), .QN(WX7249) );
  INVX0 U6053_U2 ( .INP(WX7184), .ZN(U6053_n1) );
  NOR2X0 U6053_U1 ( .IN1(n5399), .IN2(U6053_n1), .QN(WX7247) );
  INVX0 U6054_U2 ( .INP(WX7182), .ZN(U6054_n1) );
  NOR2X0 U6054_U1 ( .IN1(n5399), .IN2(U6054_n1), .QN(WX7245) );
  INVX0 U6055_U2 ( .INP(WX7180), .ZN(U6055_n1) );
  NOR2X0 U6055_U1 ( .IN1(n5399), .IN2(U6055_n1), .QN(WX7243) );
  INVX0 U6056_U2 ( .INP(WX7178), .ZN(U6056_n1) );
  NOR2X0 U6056_U1 ( .IN1(n5399), .IN2(U6056_n1), .QN(WX7241) );
  INVX0 U6057_U2 ( .INP(WX7176), .ZN(U6057_n1) );
  NOR2X0 U6057_U1 ( .IN1(n5399), .IN2(U6057_n1), .QN(WX7239) );
  INVX0 U6058_U2 ( .INP(WX7174), .ZN(U6058_n1) );
  NOR2X0 U6058_U1 ( .IN1(n5399), .IN2(U6058_n1), .QN(WX7237) );
  INVX0 U6059_U2 ( .INP(WX7172), .ZN(U6059_n1) );
  NOR2X0 U6059_U1 ( .IN1(n5399), .IN2(U6059_n1), .QN(WX7235) );
  INVX0 U6060_U2 ( .INP(WX7170), .ZN(U6060_n1) );
  NOR2X0 U6060_U1 ( .IN1(n5399), .IN2(U6060_n1), .QN(WX7233) );
  INVX0 U6061_U2 ( .INP(WX7168), .ZN(U6061_n1) );
  NOR2X0 U6061_U1 ( .IN1(n5399), .IN2(U6061_n1), .QN(WX7231) );
  INVX0 U6062_U2 ( .INP(WX7166), .ZN(U6062_n1) );
  NOR2X0 U6062_U1 ( .IN1(n5400), .IN2(U6062_n1), .QN(WX7229) );
  INVX0 U6063_U2 ( .INP(WX7164), .ZN(U6063_n1) );
  NOR2X0 U6063_U1 ( .IN1(n5400), .IN2(U6063_n1), .QN(WX7227) );
  INVX0 U6064_U2 ( .INP(WX7162), .ZN(U6064_n1) );
  NOR2X0 U6064_U1 ( .IN1(n5400), .IN2(U6064_n1), .QN(WX7225) );
  INVX0 U6065_U2 ( .INP(WX7160), .ZN(U6065_n1) );
  NOR2X0 U6065_U1 ( .IN1(n5400), .IN2(U6065_n1), .QN(WX7223) );
  INVX0 U6066_U2 ( .INP(WX7158), .ZN(U6066_n1) );
  NOR2X0 U6066_U1 ( .IN1(n5400), .IN2(U6066_n1), .QN(WX7221) );
  INVX0 U6067_U2 ( .INP(WX7156), .ZN(U6067_n1) );
  NOR2X0 U6067_U1 ( .IN1(n5400), .IN2(U6067_n1), .QN(WX7219) );
  INVX0 U6068_U2 ( .INP(WX7154), .ZN(U6068_n1) );
  NOR2X0 U6068_U1 ( .IN1(n5400), .IN2(U6068_n1), .QN(WX7217) );
  INVX0 U6069_U2 ( .INP(test_so58), .ZN(U6069_n1) );
  NOR2X0 U6069_U1 ( .IN1(n5400), .IN2(U6069_n1), .QN(WX7215) );
  INVX0 U6070_U2 ( .INP(WX7150), .ZN(U6070_n1) );
  NOR2X0 U6070_U1 ( .IN1(n5400), .IN2(U6070_n1), .QN(WX7213) );
  INVX0 U6071_U2 ( .INP(WX7148), .ZN(U6071_n1) );
  NOR2X0 U6071_U1 ( .IN1(n5402), .IN2(U6071_n1), .QN(WX7211) );
  INVX0 U6072_U2 ( .INP(WX7146), .ZN(U6072_n1) );
  NOR2X0 U6072_U1 ( .IN1(n5402), .IN2(U6072_n1), .QN(WX7209) );
  INVX0 U6073_U2 ( .INP(WX7144), .ZN(U6073_n1) );
  NOR2X0 U6073_U1 ( .IN1(n5402), .IN2(U6073_n1), .QN(WX7207) );
  INVX0 U6074_U2 ( .INP(WX7142), .ZN(U6074_n1) );
  NOR2X0 U6074_U1 ( .IN1(n5402), .IN2(U6074_n1), .QN(WX7205) );
  INVX0 U6075_U2 ( .INP(WX6007), .ZN(U6075_n1) );
  NOR2X0 U6075_U1 ( .IN1(n5402), .IN2(U6075_n1), .QN(WX6070) );
  INVX0 U6076_U2 ( .INP(test_so51), .ZN(U6076_n1) );
  NOR2X0 U6076_U1 ( .IN1(n5402), .IN2(U6076_n1), .QN(WX6068) );
  INVX0 U6077_U2 ( .INP(WX6003), .ZN(U6077_n1) );
  NOR2X0 U6077_U1 ( .IN1(n5402), .IN2(U6077_n1), .QN(WX6066) );
  INVX0 U6078_U2 ( .INP(WX6001), .ZN(U6078_n1) );
  NOR2X0 U6078_U1 ( .IN1(n5402), .IN2(U6078_n1), .QN(WX6064) );
  INVX0 U6079_U2 ( .INP(WX5999), .ZN(U6079_n1) );
  NOR2X0 U6079_U1 ( .IN1(n5402), .IN2(U6079_n1), .QN(WX6062) );
  INVX0 U6080_U2 ( .INP(WX5997), .ZN(U6080_n1) );
  NOR2X0 U6080_U1 ( .IN1(n5402), .IN2(U6080_n1), .QN(WX6060) );
  INVX0 U6081_U2 ( .INP(WX5995), .ZN(U6081_n1) );
  NOR2X0 U6081_U1 ( .IN1(n5403), .IN2(U6081_n1), .QN(WX6058) );
  INVX0 U6082_U2 ( .INP(WX5993), .ZN(U6082_n1) );
  NOR2X0 U6082_U1 ( .IN1(n5403), .IN2(U6082_n1), .QN(WX6056) );
  INVX0 U6083_U2 ( .INP(WX5991), .ZN(U6083_n1) );
  NOR2X0 U6083_U1 ( .IN1(n5403), .IN2(U6083_n1), .QN(WX6054) );
  INVX0 U6084_U2 ( .INP(WX5989), .ZN(U6084_n1) );
  NOR2X0 U6084_U1 ( .IN1(n5403), .IN2(U6084_n1), .QN(WX6052) );
  INVX0 U6085_U2 ( .INP(WX5987), .ZN(U6085_n1) );
  NOR2X0 U6085_U1 ( .IN1(n5403), .IN2(U6085_n1), .QN(WX6050) );
  INVX0 U6086_U2 ( .INP(WX5985), .ZN(U6086_n1) );
  NOR2X0 U6086_U1 ( .IN1(n5403), .IN2(U6086_n1), .QN(WX6048) );
  INVX0 U6087_U2 ( .INP(WX5983), .ZN(U6087_n1) );
  NOR2X0 U6087_U1 ( .IN1(n5403), .IN2(U6087_n1), .QN(WX6046) );
  INVX0 U6088_U2 ( .INP(WX5981), .ZN(U6088_n1) );
  NOR2X0 U6088_U1 ( .IN1(n5403), .IN2(U6088_n1), .QN(WX6044) );
  INVX0 U6089_U2 ( .INP(WX5979), .ZN(U6089_n1) );
  NOR2X0 U6089_U1 ( .IN1(n5403), .IN2(U6089_n1), .QN(WX6042) );
  INVX0 U6090_U2 ( .INP(WX5977), .ZN(U6090_n1) );
  NOR2X0 U6090_U1 ( .IN1(n5403), .IN2(U6090_n1), .QN(WX6040) );
  INVX0 U6091_U2 ( .INP(WX5975), .ZN(U6091_n1) );
  NOR2X0 U6091_U1 ( .IN1(n5404), .IN2(U6091_n1), .QN(WX6038) );
  INVX0 U6092_U2 ( .INP(WX5973), .ZN(U6092_n1) );
  NOR2X0 U6092_U1 ( .IN1(n5404), .IN2(U6092_n1), .QN(WX6036) );
  INVX0 U6093_U2 ( .INP(test_so50), .ZN(U6093_n1) );
  NOR2X0 U6093_U1 ( .IN1(n5404), .IN2(U6093_n1), .QN(WX6034) );
  INVX0 U6094_U2 ( .INP(WX5969), .ZN(U6094_n1) );
  NOR2X0 U6094_U1 ( .IN1(n5404), .IN2(U6094_n1), .QN(WX6032) );
  INVX0 U6095_U2 ( .INP(WX5967), .ZN(U6095_n1) );
  NOR2X0 U6095_U1 ( .IN1(n5404), .IN2(U6095_n1), .QN(WX6030) );
  INVX0 U6096_U2 ( .INP(WX5965), .ZN(U6096_n1) );
  NOR2X0 U6096_U1 ( .IN1(n5404), .IN2(U6096_n1), .QN(WX6028) );
  INVX0 U6097_U2 ( .INP(WX5963), .ZN(U6097_n1) );
  NOR2X0 U6097_U1 ( .IN1(n5404), .IN2(U6097_n1), .QN(WX6026) );
  INVX0 U6098_U2 ( .INP(WX5961), .ZN(U6098_n1) );
  NOR2X0 U6098_U1 ( .IN1(n5404), .IN2(U6098_n1), .QN(WX6024) );
  INVX0 U6099_U2 ( .INP(WX5959), .ZN(U6099_n1) );
  NOR2X0 U6099_U1 ( .IN1(n5404), .IN2(U6099_n1), .QN(WX6022) );
  INVX0 U6100_U2 ( .INP(WX5957), .ZN(U6100_n1) );
  NOR2X0 U6100_U1 ( .IN1(n5404), .IN2(U6100_n1), .QN(WX6020) );
  INVX0 U6101_U2 ( .INP(WX5955), .ZN(U6101_n1) );
  NOR2X0 U6101_U1 ( .IN1(n5406), .IN2(U6101_n1), .QN(WX6018) );
  INVX0 U6102_U2 ( .INP(WX5953), .ZN(U6102_n1) );
  NOR2X0 U6102_U1 ( .IN1(n5406), .IN2(U6102_n1), .QN(WX6016) );
  INVX0 U6103_U2 ( .INP(WX5951), .ZN(U6103_n1) );
  NOR2X0 U6103_U1 ( .IN1(n5406), .IN2(U6103_n1), .QN(WX6014) );
  INVX0 U6104_U2 ( .INP(WX5949), .ZN(U6104_n1) );
  NOR2X0 U6104_U1 ( .IN1(n5406), .IN2(U6104_n1), .QN(WX6012) );
  INVX0 U6105_U2 ( .INP(WX5947), .ZN(U6105_n1) );
  NOR2X0 U6105_U1 ( .IN1(n5406), .IN2(U6105_n1), .QN(WX6010) );
  INVX0 U6106_U2 ( .INP(WX5945), .ZN(U6106_n1) );
  NOR2X0 U6106_U1 ( .IN1(n5406), .IN2(U6106_n1), .QN(WX6008) );
  INVX0 U6107_U2 ( .INP(WX5943), .ZN(U6107_n1) );
  NOR2X0 U6107_U1 ( .IN1(n5406), .IN2(U6107_n1), .QN(WX6006) );
  INVX0 U6108_U2 ( .INP(WX5941), .ZN(U6108_n1) );
  NOR2X0 U6108_U1 ( .IN1(n5407), .IN2(U6108_n1), .QN(WX6004) );
  INVX0 U6109_U2 ( .INP(WX5929), .ZN(U6109_n1) );
  NOR2X0 U6109_U1 ( .IN1(n5407), .IN2(U6109_n1), .QN(WX5992) );
  INVX0 U6110_U2 ( .INP(WX5927), .ZN(U6110_n1) );
  NOR2X0 U6110_U1 ( .IN1(n5407), .IN2(U6110_n1), .QN(WX5990) );
  INVX0 U6111_U2 ( .INP(WX5925), .ZN(U6111_n1) );
  NOR2X0 U6111_U1 ( .IN1(n5407), .IN2(U6111_n1), .QN(WX5988) );
  INVX0 U6112_U2 ( .INP(WX5923), .ZN(U6112_n1) );
  NOR2X0 U6112_U1 ( .IN1(n5407), .IN2(U6112_n1), .QN(WX5986) );
  INVX0 U6113_U2 ( .INP(WX5921), .ZN(U6113_n1) );
  NOR2X0 U6113_U1 ( .IN1(n5407), .IN2(U6113_n1), .QN(WX5984) );
  INVX0 U6114_U2 ( .INP(WX5919), .ZN(U6114_n1) );
  NOR2X0 U6114_U1 ( .IN1(n5414), .IN2(U6114_n1), .QN(WX5982) );
  INVX0 U6115_U2 ( .INP(WX5917), .ZN(U6115_n1) );
  NOR2X0 U6115_U1 ( .IN1(n5407), .IN2(U6115_n1), .QN(WX5980) );
  INVX0 U6116_U2 ( .INP(WX5915), .ZN(U6116_n1) );
  NOR2X0 U6116_U1 ( .IN1(n5408), .IN2(U6116_n1), .QN(WX5978) );
  INVX0 U6117_U2 ( .INP(WX5913), .ZN(U6117_n1) );
  NOR2X0 U6117_U1 ( .IN1(n5408), .IN2(U6117_n1), .QN(WX5976) );
  INVX0 U6118_U2 ( .INP(WX5911), .ZN(U6118_n1) );
  NOR2X0 U6118_U1 ( .IN1(n5408), .IN2(U6118_n1), .QN(WX5974) );
  INVX0 U6119_U2 ( .INP(WX5909), .ZN(U6119_n1) );
  NOR2X0 U6119_U1 ( .IN1(n5408), .IN2(U6119_n1), .QN(WX5972) );
  INVX0 U6120_U2 ( .INP(WX5907), .ZN(U6120_n1) );
  NOR2X0 U6120_U1 ( .IN1(n5408), .IN2(U6120_n1), .QN(WX5970) );
  INVX0 U6121_U2 ( .INP(WX5905), .ZN(U6121_n1) );
  NOR2X0 U6121_U1 ( .IN1(n5408), .IN2(U6121_n1), .QN(WX5968) );
  INVX0 U6122_U2 ( .INP(test_so48), .ZN(U6122_n1) );
  NOR2X0 U6122_U1 ( .IN1(n5408), .IN2(U6122_n1), .QN(WX5966) );
  INVX0 U6123_U2 ( .INP(WX5901), .ZN(U6123_n1) );
  NOR2X0 U6123_U1 ( .IN1(n5408), .IN2(U6123_n1), .QN(WX5964) );
  INVX0 U6124_U2 ( .INP(WX5899), .ZN(U6124_n1) );
  NOR2X0 U6124_U1 ( .IN1(n5407), .IN2(U6124_n1), .QN(WX5962) );
  INVX0 U6125_U2 ( .INP(WX5897), .ZN(U6125_n1) );
  NOR2X0 U6125_U1 ( .IN1(n5408), .IN2(U6125_n1), .QN(WX5960) );
  INVX0 U6126_U2 ( .INP(WX5895), .ZN(U6126_n1) );
  NOR2X0 U6126_U1 ( .IN1(n5408), .IN2(U6126_n1), .QN(WX5958) );
  INVX0 U6127_U2 ( .INP(WX5893), .ZN(U6127_n1) );
  NOR2X0 U6127_U1 ( .IN1(n5408), .IN2(U6127_n1), .QN(WX5956) );
  INVX0 U6128_U2 ( .INP(WX5891), .ZN(U6128_n1) );
  NOR2X0 U6128_U1 ( .IN1(n5407), .IN2(U6128_n1), .QN(WX5954) );
  INVX0 U6129_U2 ( .INP(WX5889), .ZN(U6129_n1) );
  NOR2X0 U6129_U1 ( .IN1(n5407), .IN2(U6129_n1), .QN(WX5952) );
  INVX0 U6130_U2 ( .INP(WX5887), .ZN(U6130_n1) );
  NOR2X0 U6130_U1 ( .IN1(n5407), .IN2(U6130_n1), .QN(WX5950) );
  INVX0 U6131_U2 ( .INP(WX5885), .ZN(U6131_n1) );
  NOR2X0 U6131_U1 ( .IN1(n5406), .IN2(U6131_n1), .QN(WX5948) );
  INVX0 U6132_U2 ( .INP(WX5883), .ZN(U6132_n1) );
  NOR2X0 U6132_U1 ( .IN1(n5406), .IN2(U6132_n1), .QN(WX5946) );
  INVX0 U6133_U2 ( .INP(WX5881), .ZN(U6133_n1) );
  NOR2X0 U6133_U1 ( .IN1(n5406), .IN2(U6133_n1), .QN(WX5944) );
  INVX0 U6134_U2 ( .INP(WX5879), .ZN(U6134_n1) );
  NOR2X0 U6134_U1 ( .IN1(n5406), .IN2(U6134_n1), .QN(WX5942) );
  INVX0 U6135_U2 ( .INP(WX5877), .ZN(U6135_n1) );
  NOR2X0 U6135_U1 ( .IN1(n5405), .IN2(U6135_n1), .QN(WX5940) );
  INVX0 U6136_U2 ( .INP(WX5875), .ZN(U6136_n1) );
  NOR2X0 U6136_U1 ( .IN1(n5405), .IN2(U6136_n1), .QN(WX5938) );
  INVX0 U6137_U2 ( .INP(WX5873), .ZN(U6137_n1) );
  NOR2X0 U6137_U1 ( .IN1(n5405), .IN2(U6137_n1), .QN(WX5936) );
  INVX0 U6138_U2 ( .INP(WX5871), .ZN(U6138_n1) );
  NOR2X0 U6138_U1 ( .IN1(n5405), .IN2(U6138_n1), .QN(WX5934) );
  INVX0 U6139_U2 ( .INP(test_so47), .ZN(U6139_n1) );
  NOR2X0 U6139_U1 ( .IN1(n5405), .IN2(U6139_n1), .QN(WX5932) );
  INVX0 U6140_U2 ( .INP(WX5867), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n5405), .IN2(U6140_n1), .QN(WX5930) );
  INVX0 U6141_U2 ( .INP(WX5865), .ZN(U6141_n1) );
  NOR2X0 U6141_U1 ( .IN1(n5405), .IN2(U6141_n1), .QN(WX5928) );
  INVX0 U6142_U2 ( .INP(WX5863), .ZN(U6142_n1) );
  NOR2X0 U6142_U1 ( .IN1(n5405), .IN2(U6142_n1), .QN(WX5926) );
  INVX0 U6143_U2 ( .INP(WX5861), .ZN(U6143_n1) );
  NOR2X0 U6143_U1 ( .IN1(n5405), .IN2(U6143_n1), .QN(WX5924) );
  INVX0 U6144_U2 ( .INP(WX5859), .ZN(U6144_n1) );
  NOR2X0 U6144_U1 ( .IN1(n5405), .IN2(U6144_n1), .QN(WX5922) );
  INVX0 U6145_U2 ( .INP(WX5857), .ZN(U6145_n1) );
  NOR2X0 U6145_U1 ( .IN1(n5405), .IN2(U6145_n1), .QN(WX5920) );
  INVX0 U6146_U2 ( .INP(WX5855), .ZN(U6146_n1) );
  NOR2X0 U6146_U1 ( .IN1(n5404), .IN2(U6146_n1), .QN(WX5918) );
  INVX0 U6147_U2 ( .INP(WX5853), .ZN(U6147_n1) );
  NOR2X0 U6147_U1 ( .IN1(n5402), .IN2(U6147_n1), .QN(WX5916) );
  INVX0 U6148_U2 ( .INP(WX5851), .ZN(U6148_n1) );
  NOR2X0 U6148_U1 ( .IN1(n5401), .IN2(U6148_n1), .QN(WX5914) );
  INVX0 U6149_U2 ( .INP(WX5849), .ZN(U6149_n1) );
  NOR2X0 U6149_U1 ( .IN1(n5401), .IN2(U6149_n1), .QN(WX5912) );
  INVX0 U6150_U2 ( .INP(WX4714), .ZN(U6150_n1) );
  NOR2X0 U6150_U1 ( .IN1(n5401), .IN2(U6150_n1), .QN(WX4777) );
  INVX0 U6151_U2 ( .INP(WX4712), .ZN(U6151_n1) );
  NOR2X0 U6151_U1 ( .IN1(n5401), .IN2(U6151_n1), .QN(WX4775) );
  INVX0 U6152_U2 ( .INP(WX4710), .ZN(U6152_n1) );
  NOR2X0 U6152_U1 ( .IN1(n5401), .IN2(U6152_n1), .QN(WX4773) );
  INVX0 U6153_U2 ( .INP(WX4708), .ZN(U6153_n1) );
  NOR2X0 U6153_U1 ( .IN1(n5401), .IN2(U6153_n1), .QN(WX4771) );
  INVX0 U6154_U2 ( .INP(WX4706), .ZN(U6154_n1) );
  NOR2X0 U6154_U1 ( .IN1(n5401), .IN2(U6154_n1), .QN(WX4769) );
  INVX0 U6155_U2 ( .INP(WX4704), .ZN(U6155_n1) );
  NOR2X0 U6155_U1 ( .IN1(n5401), .IN2(U6155_n1), .QN(WX4767) );
  INVX0 U6156_U2 ( .INP(WX4702), .ZN(U6156_n1) );
  NOR2X0 U6156_U1 ( .IN1(n5401), .IN2(U6156_n1), .QN(WX4765) );
  INVX0 U6157_U2 ( .INP(WX4700), .ZN(U6157_n1) );
  NOR2X0 U6157_U1 ( .IN1(n5401), .IN2(U6157_n1), .QN(WX4763) );
  INVX0 U6158_U2 ( .INP(WX4698), .ZN(U6158_n1) );
  NOR2X0 U6158_U1 ( .IN1(n5401), .IN2(U6158_n1), .QN(WX4761) );
  INVX0 U6159_U2 ( .INP(WX4696), .ZN(U6159_n1) );
  NOR2X0 U6159_U1 ( .IN1(n5400), .IN2(U6159_n1), .QN(WX4759) );
  INVX0 U6160_U2 ( .INP(WX4694), .ZN(U6160_n1) );
  NOR2X0 U6160_U1 ( .IN1(n5400), .IN2(U6160_n1), .QN(WX4757) );
  INVX0 U6161_U2 ( .INP(WX4692), .ZN(U6161_n1) );
  NOR2X0 U6161_U1 ( .IN1(n5399), .IN2(U6161_n1), .QN(WX4755) );
  INVX0 U6162_U2 ( .INP(WX4690), .ZN(U6162_n1) );
  NOR2X0 U6162_U1 ( .IN1(n5363), .IN2(U6162_n1), .QN(WX4753) );
  INVX0 U6163_U2 ( .INP(test_so39), .ZN(U6163_n1) );
  NOR2X0 U6163_U1 ( .IN1(n5363), .IN2(U6163_n1), .QN(WX4751) );
  INVX0 U6164_U2 ( .INP(WX4686), .ZN(U6164_n1) );
  NOR2X0 U6164_U1 ( .IN1(n5363), .IN2(U6164_n1), .QN(WX4749) );
  INVX0 U6165_U2 ( .INP(WX4684), .ZN(U6165_n1) );
  NOR2X0 U6165_U1 ( .IN1(n5363), .IN2(U6165_n1), .QN(WX4747) );
  INVX0 U6166_U2 ( .INP(WX4682), .ZN(U6166_n1) );
  NOR2X0 U6166_U1 ( .IN1(n5363), .IN2(U6166_n1), .QN(WX4745) );
  INVX0 U6167_U2 ( .INP(WX4680), .ZN(U6167_n1) );
  NOR2X0 U6167_U1 ( .IN1(n5363), .IN2(U6167_n1), .QN(WX4743) );
  INVX0 U6168_U2 ( .INP(WX4678), .ZN(U6168_n1) );
  NOR2X0 U6168_U1 ( .IN1(n5363), .IN2(U6168_n1), .QN(WX4741) );
  INVX0 U6169_U2 ( .INP(WX4676), .ZN(U6169_n1) );
  NOR2X0 U6169_U1 ( .IN1(n5363), .IN2(U6169_n1), .QN(WX4739) );
  INVX0 U6170_U2 ( .INP(WX4674), .ZN(U6170_n1) );
  NOR2X0 U6170_U1 ( .IN1(n5363), .IN2(U6170_n1), .QN(WX4737) );
  INVX0 U6171_U2 ( .INP(WX4672), .ZN(U6171_n1) );
  NOR2X0 U6171_U1 ( .IN1(n5363), .IN2(U6171_n1), .QN(WX4735) );
  INVX0 U6172_U2 ( .INP(WX4670), .ZN(U6172_n1) );
  NOR2X0 U6172_U1 ( .IN1(n5363), .IN2(U6172_n1), .QN(WX4733) );
  INVX0 U6173_U2 ( .INP(WX4668), .ZN(U6173_n1) );
  NOR2X0 U6173_U1 ( .IN1(n5362), .IN2(U6173_n1), .QN(WX4731) );
  INVX0 U6174_U2 ( .INP(WX4666), .ZN(U6174_n1) );
  NOR2X0 U6174_U1 ( .IN1(n5362), .IN2(U6174_n1), .QN(WX4729) );
  INVX0 U6175_U2 ( .INP(WX4664), .ZN(U6175_n1) );
  NOR2X0 U6175_U1 ( .IN1(n5362), .IN2(U6175_n1), .QN(WX4727) );
  INVX0 U6176_U2 ( .INP(WX4662), .ZN(U6176_n1) );
  NOR2X0 U6176_U1 ( .IN1(n5362), .IN2(U6176_n1), .QN(WX4725) );
  INVX0 U6177_U2 ( .INP(WX4660), .ZN(U6177_n1) );
  NOR2X0 U6177_U1 ( .IN1(n5362), .IN2(U6177_n1), .QN(WX4723) );
  INVX0 U6178_U2 ( .INP(WX4658), .ZN(U6178_n1) );
  NOR2X0 U6178_U1 ( .IN1(n5362), .IN2(U6178_n1), .QN(WX4721) );
  INVX0 U6179_U2 ( .INP(WX4656), .ZN(U6179_n1) );
  NOR2X0 U6179_U1 ( .IN1(n5362), .IN2(U6179_n1), .QN(WX4719) );
  INVX0 U6180_U2 ( .INP(test_so38), .ZN(U6180_n1) );
  NOR2X0 U6180_U1 ( .IN1(n5362), .IN2(U6180_n1), .QN(WX4717) );
  INVX0 U6181_U2 ( .INP(WX4652), .ZN(U6181_n1) );
  NOR2X0 U6181_U1 ( .IN1(n5362), .IN2(U6181_n1), .QN(WX4715) );
  INVX0 U6182_U2 ( .INP(WX4650), .ZN(U6182_n1) );
  NOR2X0 U6182_U1 ( .IN1(n5362), .IN2(U6182_n1), .QN(WX4713) );
  INVX0 U6183_U2 ( .INP(WX4648), .ZN(U6183_n1) );
  NOR2X0 U6183_U1 ( .IN1(n5362), .IN2(U6183_n1), .QN(WX4711) );
  INVX0 U6184_U2 ( .INP(WX4646), .ZN(U6184_n1) );
  NOR2X0 U6184_U1 ( .IN1(n5361), .IN2(U6184_n1), .QN(WX4709) );
  INVX0 U6185_U2 ( .INP(WX4644), .ZN(U6185_n1) );
  NOR2X0 U6185_U1 ( .IN1(n5361), .IN2(U6185_n1), .QN(WX4707) );
  INVX0 U6186_U2 ( .INP(WX4642), .ZN(U6186_n1) );
  NOR2X0 U6186_U1 ( .IN1(n5361), .IN2(U6186_n1), .QN(WX4705) );
  INVX0 U6187_U2 ( .INP(WX4640), .ZN(U6187_n1) );
  NOR2X0 U6187_U1 ( .IN1(n5361), .IN2(U6187_n1), .QN(WX4703) );
  INVX0 U6188_U2 ( .INP(WX4638), .ZN(U6188_n1) );
  NOR2X0 U6188_U1 ( .IN1(n5361), .IN2(U6188_n1), .QN(WX4701) );
  INVX0 U6189_U2 ( .INP(WX4636), .ZN(U6189_n1) );
  NOR2X0 U6189_U1 ( .IN1(n5361), .IN2(U6189_n1), .QN(WX4699) );
  INVX0 U6190_U2 ( .INP(WX4634), .ZN(U6190_n1) );
  NOR2X0 U6190_U1 ( .IN1(n5361), .IN2(U6190_n1), .QN(WX4697) );
  INVX0 U6191_U2 ( .INP(WX4632), .ZN(U6191_n1) );
  NOR2X0 U6191_U1 ( .IN1(n5361), .IN2(U6191_n1), .QN(WX4695) );
  INVX0 U6192_U2 ( .INP(WX4630), .ZN(U6192_n1) );
  NOR2X0 U6192_U1 ( .IN1(n5361), .IN2(U6192_n1), .QN(WX4693) );
  INVX0 U6193_U2 ( .INP(WX4628), .ZN(U6193_n1) );
  NOR2X0 U6193_U1 ( .IN1(n5361), .IN2(U6193_n1), .QN(WX4691) );
  INVX0 U6194_U2 ( .INP(WX4626), .ZN(U6194_n1) );
  NOR2X0 U6194_U1 ( .IN1(n5361), .IN2(U6194_n1), .QN(WX4689) );
  INVX0 U6195_U2 ( .INP(WX4624), .ZN(U6195_n1) );
  NOR2X0 U6195_U1 ( .IN1(n5360), .IN2(U6195_n1), .QN(WX4687) );
  INVX0 U6196_U2 ( .INP(WX4622), .ZN(U6196_n1) );
  NOR2X0 U6196_U1 ( .IN1(n5360), .IN2(U6196_n1), .QN(WX4685) );
  INVX0 U6197_U2 ( .INP(test_so37), .ZN(U6197_n1) );
  NOR2X0 U6197_U1 ( .IN1(n5360), .IN2(U6197_n1), .QN(WX4683) );
  INVX0 U6198_U2 ( .INP(WX4618), .ZN(U6198_n1) );
  NOR2X0 U6198_U1 ( .IN1(n5360), .IN2(U6198_n1), .QN(WX4681) );
  INVX0 U6199_U2 ( .INP(WX4616), .ZN(U6199_n1) );
  NOR2X0 U6199_U1 ( .IN1(n5360), .IN2(U6199_n1), .QN(WX4679) );
  INVX0 U6200_U2 ( .INP(WX4614), .ZN(U6200_n1) );
  NOR2X0 U6200_U1 ( .IN1(n5360), .IN2(U6200_n1), .QN(WX4677) );
  INVX0 U6201_U2 ( .INP(WX4612), .ZN(U6201_n1) );
  NOR2X0 U6201_U1 ( .IN1(n5360), .IN2(U6201_n1), .QN(WX4675) );
  INVX0 U6202_U2 ( .INP(WX4610), .ZN(U6202_n1) );
  NOR2X0 U6202_U1 ( .IN1(n5360), .IN2(U6202_n1), .QN(WX4673) );
  INVX0 U6203_U2 ( .INP(WX4608), .ZN(U6203_n1) );
  NOR2X0 U6203_U1 ( .IN1(n5360), .IN2(U6203_n1), .QN(WX4671) );
  INVX0 U6204_U2 ( .INP(WX4606), .ZN(U6204_n1) );
  NOR2X0 U6204_U1 ( .IN1(n5360), .IN2(U6204_n1), .QN(WX4669) );
  INVX0 U6205_U2 ( .INP(WX4604), .ZN(U6205_n1) );
  NOR2X0 U6205_U1 ( .IN1(n5360), .IN2(U6205_n1), .QN(WX4667) );
  INVX0 U6206_U2 ( .INP(WX4602), .ZN(U6206_n1) );
  NOR2X0 U6206_U1 ( .IN1(n5359), .IN2(U6206_n1), .QN(WX4665) );
  INVX0 U6207_U2 ( .INP(WX4600), .ZN(U6207_n1) );
  NOR2X0 U6207_U1 ( .IN1(n5359), .IN2(U6207_n1), .QN(WX4663) );
  INVX0 U6208_U2 ( .INP(WX4598), .ZN(U6208_n1) );
  NOR2X0 U6208_U1 ( .IN1(n5359), .IN2(U6208_n1), .QN(WX4661) );
  INVX0 U6209_U2 ( .INP(WX4596), .ZN(U6209_n1) );
  NOR2X0 U6209_U1 ( .IN1(n5359), .IN2(U6209_n1), .QN(WX4659) );
  INVX0 U6210_U2 ( .INP(WX4594), .ZN(U6210_n1) );
  NOR2X0 U6210_U1 ( .IN1(n5359), .IN2(U6210_n1), .QN(WX4657) );
  INVX0 U6211_U2 ( .INP(WX4592), .ZN(U6211_n1) );
  NOR2X0 U6211_U1 ( .IN1(n5359), .IN2(U6211_n1), .QN(WX4655) );
  INVX0 U6212_U2 ( .INP(WX4590), .ZN(U6212_n1) );
  NOR2X0 U6212_U1 ( .IN1(n5359), .IN2(U6212_n1), .QN(WX4653) );
  INVX0 U6213_U2 ( .INP(WX4588), .ZN(U6213_n1) );
  NOR2X0 U6213_U1 ( .IN1(n5359), .IN2(U6213_n1), .QN(WX4651) );
  INVX0 U6214_U2 ( .INP(test_so36), .ZN(U6214_n1) );
  NOR2X0 U6214_U1 ( .IN1(n5359), .IN2(U6214_n1), .QN(WX4649) );
  INVX0 U6215_U2 ( .INP(WX4584), .ZN(U6215_n1) );
  NOR2X0 U6215_U1 ( .IN1(n5359), .IN2(U6215_n1), .QN(WX4647) );
  INVX0 U6216_U2 ( .INP(WX4582), .ZN(U6216_n1) );
  NOR2X0 U6216_U1 ( .IN1(n5359), .IN2(U6216_n1), .QN(WX4645) );
  INVX0 U6217_U2 ( .INP(WX4580), .ZN(U6217_n1) );
  NOR2X0 U6217_U1 ( .IN1(n5358), .IN2(U6217_n1), .QN(WX4643) );
  INVX0 U6218_U2 ( .INP(WX4578), .ZN(U6218_n1) );
  NOR2X0 U6218_U1 ( .IN1(n5358), .IN2(U6218_n1), .QN(WX4641) );
  INVX0 U6219_U2 ( .INP(WX4576), .ZN(U6219_n1) );
  NOR2X0 U6219_U1 ( .IN1(n5358), .IN2(U6219_n1), .QN(WX4639) );
  INVX0 U6220_U2 ( .INP(WX4574), .ZN(U6220_n1) );
  NOR2X0 U6220_U1 ( .IN1(n5358), .IN2(U6220_n1), .QN(WX4637) );
  INVX0 U6221_U2 ( .INP(WX4572), .ZN(U6221_n1) );
  NOR2X0 U6221_U1 ( .IN1(n5358), .IN2(U6221_n1), .QN(WX4635) );
  INVX0 U6222_U2 ( .INP(WX4570), .ZN(U6222_n1) );
  NOR2X0 U6222_U1 ( .IN1(n5358), .IN2(U6222_n1), .QN(WX4633) );
  INVX0 U6223_U2 ( .INP(WX4568), .ZN(U6223_n1) );
  NOR2X0 U6223_U1 ( .IN1(n5358), .IN2(U6223_n1), .QN(WX4631) );
  INVX0 U6224_U2 ( .INP(WX4566), .ZN(U6224_n1) );
  NOR2X0 U6224_U1 ( .IN1(n5358), .IN2(U6224_n1), .QN(WX4629) );
  INVX0 U6225_U2 ( .INP(WX4564), .ZN(U6225_n1) );
  NOR2X0 U6225_U1 ( .IN1(n5358), .IN2(U6225_n1), .QN(WX4627) );
  INVX0 U6226_U2 ( .INP(WX4562), .ZN(U6226_n1) );
  NOR2X0 U6226_U1 ( .IN1(n5358), .IN2(U6226_n1), .QN(WX4625) );
  INVX0 U6227_U2 ( .INP(WX4560), .ZN(U6227_n1) );
  NOR2X0 U6227_U1 ( .IN1(n5358), .IN2(U6227_n1), .QN(WX4623) );
  INVX0 U6228_U2 ( .INP(WX4558), .ZN(U6228_n1) );
  NOR2X0 U6228_U1 ( .IN1(n5357), .IN2(U6228_n1), .QN(WX4621) );
  INVX0 U6229_U2 ( .INP(WX4556), .ZN(U6229_n1) );
  NOR2X0 U6229_U1 ( .IN1(n5357), .IN2(U6229_n1), .QN(WX4619) );
  INVX0 U6230_U2 ( .INP(WX3421), .ZN(U6230_n1) );
  NOR2X0 U6230_U1 ( .IN1(n5357), .IN2(U6230_n1), .QN(WX3484) );
  INVX0 U6231_U2 ( .INP(WX3419), .ZN(U6231_n1) );
  NOR2X0 U6231_U1 ( .IN1(n5357), .IN2(U6231_n1), .QN(WX3482) );
  INVX0 U6232_U2 ( .INP(WX3417), .ZN(U6232_n1) );
  NOR2X0 U6232_U1 ( .IN1(n5357), .IN2(U6232_n1), .QN(WX3480) );
  INVX0 U6233_U2 ( .INP(WX3415), .ZN(U6233_n1) );
  NOR2X0 U6233_U1 ( .IN1(n5357), .IN2(U6233_n1), .QN(WX3478) );
  INVX0 U6234_U2 ( .INP(WX3413), .ZN(U6234_n1) );
  NOR2X0 U6234_U1 ( .IN1(n5357), .IN2(U6234_n1), .QN(WX3476) );
  INVX0 U6235_U2 ( .INP(WX3411), .ZN(U6235_n1) );
  NOR2X0 U6235_U1 ( .IN1(n5357), .IN2(U6235_n1), .QN(WX3474) );
  INVX0 U6236_U2 ( .INP(WX3409), .ZN(U6236_n1) );
  NOR2X0 U6236_U1 ( .IN1(n5357), .IN2(U6236_n1), .QN(WX3472) );
  INVX0 U6237_U2 ( .INP(WX3407), .ZN(U6237_n1) );
  NOR2X0 U6237_U1 ( .IN1(n5357), .IN2(U6237_n1), .QN(WX3470) );
  INVX0 U6238_U2 ( .INP(test_so28), .ZN(U6238_n1) );
  NOR2X0 U6238_U1 ( .IN1(n5357), .IN2(U6238_n1), .QN(WX3468) );
  INVX0 U6239_U2 ( .INP(WX3403), .ZN(U6239_n1) );
  NOR2X0 U6239_U1 ( .IN1(n5356), .IN2(U6239_n1), .QN(WX3466) );
  INVX0 U6240_U2 ( .INP(WX3401), .ZN(U6240_n1) );
  NOR2X0 U6240_U1 ( .IN1(n5356), .IN2(U6240_n1), .QN(WX3464) );
  INVX0 U6241_U2 ( .INP(WX3399), .ZN(U6241_n1) );
  NOR2X0 U6241_U1 ( .IN1(n5356), .IN2(U6241_n1), .QN(WX3462) );
  INVX0 U6242_U2 ( .INP(WX3397), .ZN(U6242_n1) );
  NOR2X0 U6242_U1 ( .IN1(n5356), .IN2(U6242_n1), .QN(WX3460) );
  INVX0 U6243_U2 ( .INP(WX3395), .ZN(U6243_n1) );
  NOR2X0 U6243_U1 ( .IN1(n5377), .IN2(U6243_n1), .QN(WX3458) );
  INVX0 U6244_U2 ( .INP(WX3393), .ZN(U6244_n1) );
  NOR2X0 U6244_U1 ( .IN1(n5414), .IN2(U6244_n1), .QN(WX3456) );
  INVX0 U6245_U2 ( .INP(WX3391), .ZN(U6245_n1) );
  NOR2X0 U6245_U1 ( .IN1(n5415), .IN2(U6245_n1), .QN(WX3454) );
  INVX0 U6246_U2 ( .INP(WX3389), .ZN(U6246_n1) );
  NOR2X0 U6246_U1 ( .IN1(n5416), .IN2(U6246_n1), .QN(WX3452) );
  INVX0 U6247_U2 ( .INP(WX3387), .ZN(U6247_n1) );
  NOR2X0 U6247_U1 ( .IN1(n5417), .IN2(U6247_n1), .QN(WX3450) );
  INVX0 U6248_U2 ( .INP(WX3385), .ZN(U6248_n1) );
  NOR2X0 U6248_U1 ( .IN1(n5418), .IN2(U6248_n1), .QN(WX3448) );
  INVX0 U6249_U2 ( .INP(WX3383), .ZN(U6249_n1) );
  NOR2X0 U6249_U1 ( .IN1(n5403), .IN2(U6249_n1), .QN(WX3446) );
  INVX0 U6250_U2 ( .INP(WX3381), .ZN(U6250_n1) );
  NOR2X0 U6250_U1 ( .IN1(n5404), .IN2(U6250_n1), .QN(WX3444) );
  INVX0 U6251_U2 ( .INP(WX3379), .ZN(U6251_n1) );
  NOR2X0 U6251_U1 ( .IN1(n5353), .IN2(U6251_n1), .QN(WX3442) );
  INVX0 U6252_U2 ( .INP(WX3377), .ZN(U6252_n1) );
  NOR2X0 U6252_U1 ( .IN1(n5353), .IN2(U6252_n1), .QN(WX3440) );
  INVX0 U6253_U2 ( .INP(WX3375), .ZN(U6253_n1) );
  NOR2X0 U6253_U1 ( .IN1(n5353), .IN2(U6253_n1), .QN(WX3438) );
  INVX0 U6254_U2 ( .INP(WX3373), .ZN(U6254_n1) );
  NOR2X0 U6254_U1 ( .IN1(n5353), .IN2(U6254_n1), .QN(WX3436) );
  INVX0 U6255_U2 ( .INP(WX3371), .ZN(U6255_n1) );
  NOR2X0 U6255_U1 ( .IN1(n5353), .IN2(U6255_n1), .QN(WX3434) );
  INVX0 U6256_U2 ( .INP(test_so27), .ZN(U6256_n1) );
  NOR2X0 U6256_U1 ( .IN1(n5353), .IN2(U6256_n1), .QN(WX3432) );
  INVX0 U6257_U2 ( .INP(WX3367), .ZN(U6257_n1) );
  NOR2X0 U6257_U1 ( .IN1(n5353), .IN2(U6257_n1), .QN(WX3430) );
  INVX0 U6258_U2 ( .INP(WX3365), .ZN(U6258_n1) );
  NOR2X0 U6258_U1 ( .IN1(n5353), .IN2(U6258_n1), .QN(WX3428) );
  INVX0 U6259_U2 ( .INP(WX3363), .ZN(U6259_n1) );
  NOR2X0 U6259_U1 ( .IN1(n5353), .IN2(U6259_n1), .QN(WX3426) );
  INVX0 U6260_U2 ( .INP(WX3361), .ZN(U6260_n1) );
  NOR2X0 U6260_U1 ( .IN1(n5353), .IN2(U6260_n1), .QN(WX3424) );
  INVX0 U6261_U2 ( .INP(WX3359), .ZN(U6261_n1) );
  NOR2X0 U6261_U1 ( .IN1(n5353), .IN2(U6261_n1), .QN(WX3422) );
  INVX0 U6262_U2 ( .INP(WX3357), .ZN(U6262_n1) );
  NOR2X0 U6262_U1 ( .IN1(n5360), .IN2(U6262_n1), .QN(WX3420) );
  INVX0 U6263_U2 ( .INP(WX3355), .ZN(U6263_n1) );
  NOR2X0 U6263_U1 ( .IN1(n5361), .IN2(U6263_n1), .QN(WX3418) );
  INVX0 U6264_U2 ( .INP(WX3353), .ZN(U6264_n1) );
  NOR2X0 U6264_U1 ( .IN1(n5362), .IN2(U6264_n1), .QN(WX3416) );
  INVX0 U6265_U2 ( .INP(WX3351), .ZN(U6265_n1) );
  NOR2X0 U6265_U1 ( .IN1(n5363), .IN2(U6265_n1), .QN(WX3414) );
  INVX0 U6266_U2 ( .INP(WX3349), .ZN(U6266_n1) );
  NOR2X0 U6266_U1 ( .IN1(n5389), .IN2(U6266_n1), .QN(WX3412) );
  INVX0 U6267_U2 ( .INP(WX3347), .ZN(U6267_n1) );
  NOR2X0 U6267_U1 ( .IN1(n5390), .IN2(U6267_n1), .QN(WX3410) );
  INVX0 U6268_U2 ( .INP(WX3345), .ZN(U6268_n1) );
  NOR2X0 U6268_U1 ( .IN1(n5391), .IN2(U6268_n1), .QN(WX3408) );
  INVX0 U6269_U2 ( .INP(WX3343), .ZN(U6269_n1) );
  NOR2X0 U6269_U1 ( .IN1(n5392), .IN2(U6269_n1), .QN(WX3406) );
  INVX0 U6270_U2 ( .INP(WX3341), .ZN(U6270_n1) );
  NOR2X0 U6270_U1 ( .IN1(n5384), .IN2(U6270_n1), .QN(WX3404) );
  INVX0 U6271_U2 ( .INP(WX3339), .ZN(U6271_n1) );
  NOR2X0 U6271_U1 ( .IN1(n5385), .IN2(U6271_n1), .QN(WX3402) );
  INVX0 U6272_U2 ( .INP(WX3337), .ZN(U6272_n1) );
  NOR2X0 U6272_U1 ( .IN1(n5386), .IN2(U6272_n1), .QN(WX3400) );
  INVX0 U6273_U2 ( .INP(WX3335), .ZN(U6273_n1) );
  NOR2X0 U6273_U1 ( .IN1(n5387), .IN2(U6273_n1), .QN(WX3398) );
  INVX0 U6274_U2 ( .INP(test_so26), .ZN(U6274_n1) );
  NOR2X0 U6274_U1 ( .IN1(n5388), .IN2(U6274_n1), .QN(WX3396) );
  INVX0 U6275_U2 ( .INP(WX3331), .ZN(U6275_n1) );
  NOR2X0 U6275_U1 ( .IN1(n5393), .IN2(U6275_n1), .QN(WX3394) );
  INVX0 U6276_U2 ( .INP(WX3329), .ZN(U6276_n1) );
  NOR2X0 U6276_U1 ( .IN1(n5394), .IN2(U6276_n1), .QN(WX3392) );
  INVX0 U6277_U2 ( .INP(WX3327), .ZN(U6277_n1) );
  NOR2X0 U6277_U1 ( .IN1(n5395), .IN2(U6277_n1), .QN(WX3390) );
  INVX0 U6278_U2 ( .INP(WX3325), .ZN(U6278_n1) );
  NOR2X0 U6278_U1 ( .IN1(n5396), .IN2(U6278_n1), .QN(WX3388) );
  INVX0 U6279_U2 ( .INP(WX3323), .ZN(U6279_n1) );
  NOR2X0 U6279_U1 ( .IN1(n5397), .IN2(U6279_n1), .QN(WX3386) );
  INVX0 U6280_U2 ( .INP(WX3321), .ZN(U6280_n1) );
  NOR2X0 U6280_U1 ( .IN1(n5374), .IN2(U6280_n1), .QN(WX3384) );
  INVX0 U6281_U2 ( .INP(WX3319), .ZN(U6281_n1) );
  NOR2X0 U6281_U1 ( .IN1(n5375), .IN2(U6281_n1), .QN(WX3382) );
  INVX0 U6282_U2 ( .INP(WX3317), .ZN(U6282_n1) );
  NOR2X0 U6282_U1 ( .IN1(n5376), .IN2(U6282_n1), .QN(WX3380) );
  INVX0 U6283_U2 ( .INP(WX3315), .ZN(U6283_n1) );
  NOR2X0 U6283_U1 ( .IN1(n5378), .IN2(U6283_n1), .QN(WX3378) );
  INVX0 U6284_U2 ( .INP(WX3313), .ZN(U6284_n1) );
  NOR2X0 U6284_U1 ( .IN1(n5379), .IN2(U6284_n1), .QN(WX3376) );
  INVX0 U6285_U2 ( .INP(WX3311), .ZN(U6285_n1) );
  NOR2X0 U6285_U1 ( .IN1(n5380), .IN2(U6285_n1), .QN(WX3374) );
  INVX0 U6286_U2 ( .INP(WX3309), .ZN(U6286_n1) );
  NOR2X0 U6286_U1 ( .IN1(n5381), .IN2(U6286_n1), .QN(WX3372) );
  INVX0 U6287_U2 ( .INP(WX3307), .ZN(U6287_n1) );
  NOR2X0 U6287_U1 ( .IN1(n5382), .IN2(U6287_n1), .QN(WX3370) );
  INVX0 U6288_U2 ( .INP(WX3305), .ZN(U6288_n1) );
  NOR2X0 U6288_U1 ( .IN1(n5383), .IN2(U6288_n1), .QN(WX3368) );
  INVX0 U6289_U2 ( .INP(WX3303), .ZN(U6289_n1) );
  NOR2X0 U6289_U1 ( .IN1(n5398), .IN2(U6289_n1), .QN(WX3366) );
  INVX0 U6290_U2 ( .INP(WX3301), .ZN(U6290_n1) );
  NOR2X0 U6290_U1 ( .IN1(n5399), .IN2(U6290_n1), .QN(WX3364) );
  INVX0 U6291_U2 ( .INP(WX3299), .ZN(U6291_n1) );
  NOR2X0 U6291_U1 ( .IN1(n5400), .IN2(U6291_n1), .QN(WX3362) );
  INVX0 U6292_U2 ( .INP(test_so25), .ZN(U6292_n1) );
  NOR2X0 U6292_U1 ( .IN1(n5401), .IN2(U6292_n1), .QN(WX3360) );
  INVX0 U6293_U2 ( .INP(WX3295), .ZN(U6293_n1) );
  NOR2X0 U6293_U1 ( .IN1(n5402), .IN2(U6293_n1), .QN(WX3358) );
  INVX0 U6294_U2 ( .INP(WX3293), .ZN(U6294_n1) );
  NOR2X0 U6294_U1 ( .IN1(n5354), .IN2(U6294_n1), .QN(WX3356) );
  INVX0 U6295_U2 ( .INP(WX3291), .ZN(U6295_n1) );
  NOR2X0 U6295_U1 ( .IN1(n5354), .IN2(U6295_n1), .QN(WX3354) );
  INVX0 U6296_U2 ( .INP(WX3289), .ZN(U6296_n1) );
  NOR2X0 U6296_U1 ( .IN1(n5354), .IN2(U6296_n1), .QN(WX3352) );
  INVX0 U6297_U2 ( .INP(WX3287), .ZN(U6297_n1) );
  NOR2X0 U6297_U1 ( .IN1(n5354), .IN2(U6297_n1), .QN(WX3350) );
  INVX0 U6298_U2 ( .INP(WX3285), .ZN(U6298_n1) );
  NOR2X0 U6298_U1 ( .IN1(n5354), .IN2(U6298_n1), .QN(WX3348) );
  INVX0 U6299_U2 ( .INP(WX3283), .ZN(U6299_n1) );
  NOR2X0 U6299_U1 ( .IN1(n5354), .IN2(U6299_n1), .QN(WX3346) );
  INVX0 U6300_U2 ( .INP(WX3281), .ZN(U6300_n1) );
  NOR2X0 U6300_U1 ( .IN1(n5354), .IN2(U6300_n1), .QN(WX3344) );
  INVX0 U6301_U2 ( .INP(WX3279), .ZN(U6301_n1) );
  NOR2X0 U6301_U1 ( .IN1(n5354), .IN2(U6301_n1), .QN(WX3342) );
  INVX0 U6302_U2 ( .INP(WX3277), .ZN(U6302_n1) );
  NOR2X0 U6302_U1 ( .IN1(n5354), .IN2(U6302_n1), .QN(WX3340) );
  INVX0 U6303_U2 ( .INP(WX3275), .ZN(U6303_n1) );
  NOR2X0 U6303_U1 ( .IN1(n5354), .IN2(U6303_n1), .QN(WX3338) );
  INVX0 U6304_U2 ( .INP(WX3273), .ZN(U6304_n1) );
  NOR2X0 U6304_U1 ( .IN1(n5354), .IN2(U6304_n1), .QN(WX3336) );
  INVX0 U6305_U2 ( .INP(WX3271), .ZN(U6305_n1) );
  NOR2X0 U6305_U1 ( .IN1(n5355), .IN2(U6305_n1), .QN(WX3334) );
  INVX0 U6306_U2 ( .INP(WX3267), .ZN(U6306_n1) );
  NOR2X0 U6306_U1 ( .IN1(n5355), .IN2(U6306_n1), .QN(WX3330) );
  INVX0 U6307_U2 ( .INP(WX2128), .ZN(U6307_n1) );
  NOR2X0 U6307_U1 ( .IN1(n5355), .IN2(U6307_n1), .QN(WX2191) );
  INVX0 U6308_U2 ( .INP(WX2126), .ZN(U6308_n1) );
  NOR2X0 U6308_U1 ( .IN1(n5355), .IN2(U6308_n1), .QN(WX2189) );
  INVX0 U6309_U2 ( .INP(WX2124), .ZN(U6309_n1) );
  NOR2X0 U6309_U1 ( .IN1(n5355), .IN2(U6309_n1), .QN(WX2187) );
  INVX0 U6310_U2 ( .INP(WX2122), .ZN(U6310_n1) );
  NOR2X0 U6310_U1 ( .IN1(n5355), .IN2(U6310_n1), .QN(WX2185) );
  INVX0 U6311_U2 ( .INP(WX2120), .ZN(U6311_n1) );
  NOR2X0 U6311_U1 ( .IN1(n5355), .IN2(U6311_n1), .QN(WX2183) );
  INVX0 U6312_U2 ( .INP(WX2118), .ZN(U6312_n1) );
  NOR2X0 U6312_U1 ( .IN1(n5355), .IN2(U6312_n1), .QN(WX2181) );
  INVX0 U6313_U2 ( .INP(WX2116), .ZN(U6313_n1) );
  NOR2X0 U6313_U1 ( .IN1(n5355), .IN2(U6313_n1), .QN(WX2179) );
  INVX0 U6314_U2 ( .INP(WX2114), .ZN(U6314_n1) );
  NOR2X0 U6314_U1 ( .IN1(n5355), .IN2(U6314_n1), .QN(WX2177) );
  INVX0 U6315_U2 ( .INP(WX2112), .ZN(U6315_n1) );
  NOR2X0 U6315_U1 ( .IN1(n5355), .IN2(U6315_n1), .QN(WX2175) );
  INVX0 U6316_U2 ( .INP(WX2110), .ZN(U6316_n1) );
  NOR2X0 U6316_U1 ( .IN1(n5356), .IN2(U6316_n1), .QN(WX2173) );
  INVX0 U6317_U2 ( .INP(WX2108), .ZN(U6317_n1) );
  NOR2X0 U6317_U1 ( .IN1(n5356), .IN2(U6317_n1), .QN(WX2171) );
  INVX0 U6318_U2 ( .INP(WX2106), .ZN(U6318_n1) );
  NOR2X0 U6318_U1 ( .IN1(n5356), .IN2(U6318_n1), .QN(WX2169) );
  INVX0 U6319_U2 ( .INP(WX2104), .ZN(U6319_n1) );
  NOR2X0 U6319_U1 ( .IN1(n5356), .IN2(U6319_n1), .QN(WX2167) );
  INVX0 U6320_U2 ( .INP(WX2102), .ZN(U6320_n1) );
  NOR2X0 U6320_U1 ( .IN1(n5356), .IN2(U6320_n1), .QN(WX2165) );
  INVX0 U6321_U2 ( .INP(test_so17), .ZN(U6321_n1) );
  NOR2X0 U6321_U1 ( .IN1(n5356), .IN2(U6321_n1), .QN(WX2163) );
  INVX0 U6322_U2 ( .INP(WX2098), .ZN(U6322_n1) );
  NOR2X0 U6322_U1 ( .IN1(n5356), .IN2(U6322_n1), .QN(WX2161) );
  INVX0 U6323_U2 ( .INP(WX2096), .ZN(U6323_n1) );
  NOR2X0 U6323_U1 ( .IN1(n5378), .IN2(U6323_n1), .QN(WX2159) );
  INVX0 U6324_U2 ( .INP(WX2094), .ZN(U6324_n1) );
  NOR2X0 U6324_U1 ( .IN1(n5378), .IN2(U6324_n1), .QN(WX2157) );
  INVX0 U6325_U2 ( .INP(WX2092), .ZN(U6325_n1) );
  NOR2X0 U6325_U1 ( .IN1(n5378), .IN2(U6325_n1), .QN(WX2155) );
  INVX0 U6326_U2 ( .INP(WX2090), .ZN(U6326_n1) );
  NOR2X0 U6326_U1 ( .IN1(n5378), .IN2(U6326_n1), .QN(WX2153) );
  INVX0 U6327_U2 ( .INP(WX2088), .ZN(U6327_n1) );
  NOR2X0 U6327_U1 ( .IN1(n5378), .IN2(U6327_n1), .QN(WX2151) );
  INVX0 U6328_U2 ( .INP(WX2086), .ZN(U6328_n1) );
  NOR2X0 U6328_U1 ( .IN1(n5378), .IN2(U6328_n1), .QN(WX2149) );
  INVX0 U6329_U2 ( .INP(WX2084), .ZN(U6329_n1) );
  NOR2X0 U6329_U1 ( .IN1(n5377), .IN2(U6329_n1), .QN(WX2147) );
  INVX0 U6330_U2 ( .INP(WX2082), .ZN(U6330_n1) );
  NOR2X0 U6330_U1 ( .IN1(n5377), .IN2(U6330_n1), .QN(WX2145) );
  INVX0 U6331_U2 ( .INP(WX2080), .ZN(U6331_n1) );
  NOR2X0 U6331_U1 ( .IN1(n5377), .IN2(U6331_n1), .QN(WX2143) );
  INVX0 U6332_U2 ( .INP(WX2078), .ZN(U6332_n1) );
  NOR2X0 U6332_U1 ( .IN1(n5377), .IN2(U6332_n1), .QN(WX2141) );
  INVX0 U6333_U2 ( .INP(WX2076), .ZN(U6333_n1) );
  NOR2X0 U6333_U1 ( .IN1(n5377), .IN2(U6333_n1), .QN(WX2139) );
  INVX0 U6334_U2 ( .INP(WX2074), .ZN(U6334_n1) );
  NOR2X0 U6334_U1 ( .IN1(n5377), .IN2(U6334_n1), .QN(WX2137) );
  INVX0 U6335_U2 ( .INP(WX2072), .ZN(U6335_n1) );
  NOR2X0 U6335_U1 ( .IN1(n5377), .IN2(U6335_n1), .QN(WX2135) );
  INVX0 U6336_U2 ( .INP(WX2070), .ZN(U6336_n1) );
  NOR2X0 U6336_U1 ( .IN1(n5377), .IN2(U6336_n1), .QN(WX2133) );
  INVX0 U6337_U2 ( .INP(WX2068), .ZN(U6337_n1) );
  NOR2X0 U6337_U1 ( .IN1(n5377), .IN2(U6337_n1), .QN(WX2131) );
  INVX0 U6338_U2 ( .INP(WX2066), .ZN(U6338_n1) );
  NOR2X0 U6338_U1 ( .IN1(n5377), .IN2(U6338_n1), .QN(WX2129) );
  INVX0 U6339_U2 ( .INP(test_so16), .ZN(U6339_n1) );
  NOR2X0 U6339_U1 ( .IN1(n5377), .IN2(U6339_n1), .QN(WX2127) );
  INVX0 U6340_U2 ( .INP(WX2062), .ZN(U6340_n1) );
  NOR2X0 U6340_U1 ( .IN1(n5376), .IN2(U6340_n1), .QN(WX2125) );
  INVX0 U6341_U2 ( .INP(WX2060), .ZN(U6341_n1) );
  NOR2X0 U6341_U1 ( .IN1(n5376), .IN2(U6341_n1), .QN(WX2123) );
  INVX0 U6342_U2 ( .INP(WX2058), .ZN(U6342_n1) );
  NOR2X0 U6342_U1 ( .IN1(n5376), .IN2(U6342_n1), .QN(WX2121) );
  INVX0 U6343_U2 ( .INP(WX2056), .ZN(U6343_n1) );
  NOR2X0 U6343_U1 ( .IN1(n5376), .IN2(U6343_n1), .QN(WX2119) );
  INVX0 U6344_U2 ( .INP(WX2054), .ZN(U6344_n1) );
  NOR2X0 U6344_U1 ( .IN1(n5376), .IN2(U6344_n1), .QN(WX2117) );
  INVX0 U6345_U2 ( .INP(WX2052), .ZN(U6345_n1) );
  NOR2X0 U6345_U1 ( .IN1(n5376), .IN2(U6345_n1), .QN(WX2115) );
  INVX0 U6346_U2 ( .INP(WX2050), .ZN(U6346_n1) );
  NOR2X0 U6346_U1 ( .IN1(n5376), .IN2(U6346_n1), .QN(WX2113) );
  INVX0 U6347_U2 ( .INP(WX2048), .ZN(U6347_n1) );
  NOR2X0 U6347_U1 ( .IN1(n5376), .IN2(U6347_n1), .QN(WX2111) );
  INVX0 U6348_U2 ( .INP(WX2046), .ZN(U6348_n1) );
  NOR2X0 U6348_U1 ( .IN1(n5376), .IN2(U6348_n1), .QN(WX2109) );
  INVX0 U6349_U2 ( .INP(WX2044), .ZN(U6349_n1) );
  NOR2X0 U6349_U1 ( .IN1(n5376), .IN2(U6349_n1), .QN(WX2107) );
  INVX0 U6350_U2 ( .INP(WX2042), .ZN(U6350_n1) );
  NOR2X0 U6350_U1 ( .IN1(n5376), .IN2(U6350_n1), .QN(WX2105) );
  INVX0 U6351_U2 ( .INP(WX2040), .ZN(U6351_n1) );
  NOR2X0 U6351_U1 ( .IN1(n5375), .IN2(U6351_n1), .QN(WX2103) );
  INVX0 U6352_U2 ( .INP(WX2038), .ZN(U6352_n1) );
  NOR2X0 U6352_U1 ( .IN1(n5375), .IN2(U6352_n1), .QN(WX2101) );
  INVX0 U6353_U2 ( .INP(WX2036), .ZN(U6353_n1) );
  NOR2X0 U6353_U1 ( .IN1(n5375), .IN2(U6353_n1), .QN(WX2099) );
  INVX0 U6354_U2 ( .INP(WX2034), .ZN(U6354_n1) );
  NOR2X0 U6354_U1 ( .IN1(n5375), .IN2(U6354_n1), .QN(WX2097) );
  INVX0 U6355_U2 ( .INP(WX2032), .ZN(U6355_n1) );
  NOR2X0 U6355_U1 ( .IN1(n5375), .IN2(U6355_n1), .QN(WX2095) );
  INVX0 U6356_U2 ( .INP(WX2030), .ZN(U6356_n1) );
  NOR2X0 U6356_U1 ( .IN1(n5375), .IN2(U6356_n1), .QN(WX2093) );
  INVX0 U6357_U2 ( .INP(test_so15), .ZN(U6357_n1) );
  NOR2X0 U6357_U1 ( .IN1(n5375), .IN2(U6357_n1), .QN(WX2091) );
  INVX0 U6358_U2 ( .INP(WX2026), .ZN(U6358_n1) );
  NOR2X0 U6358_U1 ( .IN1(n5375), .IN2(U6358_n1), .QN(WX2089) );
  INVX0 U6359_U2 ( .INP(WX2024), .ZN(U6359_n1) );
  NOR2X0 U6359_U1 ( .IN1(n5375), .IN2(U6359_n1), .QN(WX2087) );
  INVX0 U6360_U2 ( .INP(WX2022), .ZN(U6360_n1) );
  NOR2X0 U6360_U1 ( .IN1(n5375), .IN2(U6360_n1), .QN(WX2085) );
  INVX0 U6361_U2 ( .INP(WX2020), .ZN(U6361_n1) );
  NOR2X0 U6361_U1 ( .IN1(n5375), .IN2(U6361_n1), .QN(WX2083) );
  INVX0 U6362_U2 ( .INP(WX2018), .ZN(U6362_n1) );
  NOR2X0 U6362_U1 ( .IN1(n5374), .IN2(U6362_n1), .QN(WX2081) );
  INVX0 U6363_U2 ( .INP(WX2016), .ZN(U6363_n1) );
  NOR2X0 U6363_U1 ( .IN1(n5374), .IN2(U6363_n1), .QN(WX2079) );
  INVX0 U6364_U2 ( .INP(WX2014), .ZN(U6364_n1) );
  NOR2X0 U6364_U1 ( .IN1(n5374), .IN2(U6364_n1), .QN(WX2077) );
  INVX0 U6365_U2 ( .INP(WX2012), .ZN(U6365_n1) );
  NOR2X0 U6365_U1 ( .IN1(n5374), .IN2(U6365_n1), .QN(WX2075) );
  INVX0 U6366_U2 ( .INP(WX2010), .ZN(U6366_n1) );
  NOR2X0 U6366_U1 ( .IN1(n5374), .IN2(U6366_n1), .QN(WX2073) );
  INVX0 U6367_U2 ( .INP(WX2008), .ZN(U6367_n1) );
  NOR2X0 U6367_U1 ( .IN1(n5374), .IN2(U6367_n1), .QN(WX2071) );
  INVX0 U6368_U2 ( .INP(WX2006), .ZN(U6368_n1) );
  NOR2X0 U6368_U1 ( .IN1(n5374), .IN2(U6368_n1), .QN(WX2069) );
  INVX0 U6369_U2 ( .INP(WX2004), .ZN(U6369_n1) );
  NOR2X0 U6369_U1 ( .IN1(n5374), .IN2(U6369_n1), .QN(WX2067) );
  INVX0 U6370_U2 ( .INP(WX2002), .ZN(U6370_n1) );
  NOR2X0 U6370_U1 ( .IN1(n5374), .IN2(U6370_n1), .QN(WX2065) );
  INVX0 U6371_U2 ( .INP(WX2000), .ZN(U6371_n1) );
  NOR2X0 U6371_U1 ( .IN1(n5374), .IN2(U6371_n1), .QN(WX2063) );
  INVX0 U6372_U2 ( .INP(WX1998), .ZN(U6372_n1) );
  NOR2X0 U6372_U1 ( .IN1(n5374), .IN2(U6372_n1), .QN(WX2061) );
  INVX0 U6373_U2 ( .INP(WX1996), .ZN(U6373_n1) );
  NOR2X0 U6373_U1 ( .IN1(n5373), .IN2(U6373_n1), .QN(WX2059) );
  INVX0 U6374_U2 ( .INP(WX1994), .ZN(U6374_n1) );
  NOR2X0 U6374_U1 ( .IN1(n5373), .IN2(U6374_n1), .QN(WX2057) );
  INVX0 U6375_U2 ( .INP(test_so14), .ZN(U6375_n1) );
  NOR2X0 U6375_U1 ( .IN1(n5373), .IN2(U6375_n1), .QN(WX2055) );
  INVX0 U6376_U2 ( .INP(WX1990), .ZN(U6376_n1) );
  NOR2X0 U6376_U1 ( .IN1(n5373), .IN2(U6376_n1), .QN(WX2053) );
  INVX0 U6377_U2 ( .INP(WX1988), .ZN(U6377_n1) );
  NOR2X0 U6377_U1 ( .IN1(n5373), .IN2(U6377_n1), .QN(WX2051) );
  INVX0 U6378_U2 ( .INP(WX1986), .ZN(U6378_n1) );
  NOR2X0 U6378_U1 ( .IN1(n5373), .IN2(U6378_n1), .QN(WX2049) );
  INVX0 U6379_U2 ( .INP(WX1984), .ZN(U6379_n1) );
  NOR2X0 U6379_U1 ( .IN1(n5373), .IN2(U6379_n1), .QN(WX2047) );
  INVX0 U6380_U2 ( .INP(WX1982), .ZN(U6380_n1) );
  NOR2X0 U6380_U1 ( .IN1(n5373), .IN2(U6380_n1), .QN(WX2045) );
  INVX0 U6381_U2 ( .INP(WX1980), .ZN(U6381_n1) );
  NOR2X0 U6381_U1 ( .IN1(n5373), .IN2(U6381_n1), .QN(WX2043) );
  INVX0 U6382_U2 ( .INP(WX1978), .ZN(U6382_n1) );
  NOR2X0 U6382_U1 ( .IN1(n5373), .IN2(U6382_n1), .QN(WX2041) );
  INVX0 U6383_U2 ( .INP(WX1976), .ZN(U6383_n1) );
  NOR2X0 U6383_U1 ( .IN1(n5373), .IN2(U6383_n1), .QN(WX2039) );
  INVX0 U6384_U2 ( .INP(WX1974), .ZN(U6384_n1) );
  NOR2X0 U6384_U1 ( .IN1(n5372), .IN2(U6384_n1), .QN(WX2037) );
  INVX0 U6385_U2 ( .INP(WX1972), .ZN(U6385_n1) );
  NOR2X0 U6385_U1 ( .IN1(n5372), .IN2(U6385_n1), .QN(WX2035) );
  INVX0 U6386_U2 ( .INP(WX1970), .ZN(U6386_n1) );
  NOR2X0 U6386_U1 ( .IN1(n5372), .IN2(U6386_n1), .QN(WX2033) );
  INVX0 U6387_U2 ( .INP(WX835), .ZN(U6387_n1) );
  NOR2X0 U6387_U1 ( .IN1(n5372), .IN2(U6387_n1), .QN(WX898) );
  INVX0 U6388_U2 ( .INP(WX833), .ZN(U6388_n1) );
  NOR2X0 U6388_U1 ( .IN1(n5372), .IN2(U6388_n1), .QN(WX896) );
  INVX0 U6389_U2 ( .INP(test_so7), .ZN(U6389_n1) );
  NOR2X0 U6389_U1 ( .IN1(n5372), .IN2(U6389_n1), .QN(WX894) );
  INVX0 U6390_U2 ( .INP(WX829), .ZN(U6390_n1) );
  NOR2X0 U6390_U1 ( .IN1(n5372), .IN2(U6390_n1), .QN(WX892) );
  INVX0 U6391_U2 ( .INP(WX827), .ZN(U6391_n1) );
  NOR2X0 U6391_U1 ( .IN1(n5372), .IN2(U6391_n1), .QN(WX890) );
  INVX0 U6392_U2 ( .INP(WX825), .ZN(U6392_n1) );
  NOR2X0 U6392_U1 ( .IN1(n5372), .IN2(U6392_n1), .QN(WX888) );
  INVX0 U6393_U2 ( .INP(WX823), .ZN(U6393_n1) );
  NOR2X0 U6393_U1 ( .IN1(n5372), .IN2(U6393_n1), .QN(WX886) );
  INVX0 U6394_U2 ( .INP(WX821), .ZN(U6394_n1) );
  NOR2X0 U6394_U1 ( .IN1(n5372), .IN2(U6394_n1), .QN(WX884) );
  INVX0 U6395_U2 ( .INP(WX819), .ZN(U6395_n1) );
  NOR2X0 U6395_U1 ( .IN1(n5371), .IN2(U6395_n1), .QN(WX882) );
  INVX0 U6396_U2 ( .INP(WX817), .ZN(U6396_n1) );
  NOR2X0 U6396_U1 ( .IN1(n5371), .IN2(U6396_n1), .QN(WX880) );
  INVX0 U6397_U2 ( .INP(WX815), .ZN(U6397_n1) );
  NOR2X0 U6397_U1 ( .IN1(n5371), .IN2(U6397_n1), .QN(WX878) );
  INVX0 U6398_U2 ( .INP(WX813), .ZN(U6398_n1) );
  NOR2X0 U6398_U1 ( .IN1(n5371), .IN2(U6398_n1), .QN(WX876) );
  INVX0 U6399_U2 ( .INP(WX811), .ZN(U6399_n1) );
  NOR2X0 U6399_U1 ( .IN1(n5371), .IN2(U6399_n1), .QN(WX874) );
  INVX0 U6400_U2 ( .INP(WX809), .ZN(U6400_n1) );
  NOR2X0 U6400_U1 ( .IN1(n5371), .IN2(U6400_n1), .QN(WX872) );
  INVX0 U6401_U2 ( .INP(WX807), .ZN(U6401_n1) );
  NOR2X0 U6401_U1 ( .IN1(n5371), .IN2(U6401_n1), .QN(WX870) );
  INVX0 U6402_U2 ( .INP(WX805), .ZN(U6402_n1) );
  NOR2X0 U6402_U1 ( .IN1(n5371), .IN2(U6402_n1), .QN(WX868) );
  INVX0 U6403_U2 ( .INP(WX803), .ZN(U6403_n1) );
  NOR2X0 U6403_U1 ( .IN1(n5371), .IN2(U6403_n1), .QN(WX866) );
  INVX0 U6404_U2 ( .INP(WX801), .ZN(U6404_n1) );
  NOR2X0 U6404_U1 ( .IN1(n5371), .IN2(U6404_n1), .QN(WX864) );
  INVX0 U6405_U2 ( .INP(WX799), .ZN(U6405_n1) );
  NOR2X0 U6405_U1 ( .IN1(n5370), .IN2(U6405_n1), .QN(WX862) );
  INVX0 U6406_U2 ( .INP(WX797), .ZN(U6406_n1) );
  NOR2X0 U6406_U1 ( .IN1(n5370), .IN2(U6406_n1), .QN(WX860) );
  INVX0 U6407_U2 ( .INP(test_so6), .ZN(U6407_n1) );
  NOR2X0 U6407_U1 ( .IN1(n5370), .IN2(U6407_n1), .QN(WX858) );
  INVX0 U6408_U2 ( .INP(WX793), .ZN(U6408_n1) );
  NOR2X0 U6408_U1 ( .IN1(n5370), .IN2(U6408_n1), .QN(WX856) );
  INVX0 U6409_U2 ( .INP(WX791), .ZN(U6409_n1) );
  NOR2X0 U6409_U1 ( .IN1(n5370), .IN2(U6409_n1), .QN(WX854) );
  INVX0 U6410_U2 ( .INP(WX789), .ZN(U6410_n1) );
  NOR2X0 U6410_U1 ( .IN1(n5370), .IN2(U6410_n1), .QN(WX852) );
  INVX0 U6411_U2 ( .INP(WX787), .ZN(U6411_n1) );
  NOR2X0 U6411_U1 ( .IN1(n5370), .IN2(U6411_n1), .QN(WX850) );
  INVX0 U6412_U2 ( .INP(WX785), .ZN(U6412_n1) );
  NOR2X0 U6412_U1 ( .IN1(n5370), .IN2(U6412_n1), .QN(WX848) );
  INVX0 U6413_U2 ( .INP(WX783), .ZN(U6413_n1) );
  NOR2X0 U6413_U1 ( .IN1(n5370), .IN2(U6413_n1), .QN(WX846) );
  INVX0 U6414_U2 ( .INP(WX781), .ZN(U6414_n1) );
  NOR2X0 U6414_U1 ( .IN1(n5370), .IN2(U6414_n1), .QN(WX844) );
  INVX0 U6415_U2 ( .INP(WX779), .ZN(U6415_n1) );
  NOR2X0 U6415_U1 ( .IN1(n5370), .IN2(U6415_n1), .QN(WX842) );
  INVX0 U6416_U2 ( .INP(WX777), .ZN(U6416_n1) );
  NOR2X0 U6416_U1 ( .IN1(n5369), .IN2(U6416_n1), .QN(WX840) );
  INVX0 U6417_U2 ( .INP(WX775), .ZN(U6417_n1) );
  NOR2X0 U6417_U1 ( .IN1(n5369), .IN2(U6417_n1), .QN(WX838) );
  INVX0 U6418_U2 ( .INP(WX773), .ZN(U6418_n1) );
  NOR2X0 U6418_U1 ( .IN1(n5369), .IN2(U6418_n1), .QN(WX836) );
  INVX0 U6419_U2 ( .INP(WX771), .ZN(U6419_n1) );
  NOR2X0 U6419_U1 ( .IN1(n5369), .IN2(U6419_n1), .QN(WX834) );
  INVX0 U6420_U2 ( .INP(WX769), .ZN(U6420_n1) );
  NOR2X0 U6420_U1 ( .IN1(n5369), .IN2(U6420_n1), .QN(WX832) );
  INVX0 U6421_U2 ( .INP(WX767), .ZN(U6421_n1) );
  NOR2X0 U6421_U1 ( .IN1(n5369), .IN2(U6421_n1), .QN(WX830) );
  INVX0 U6422_U2 ( .INP(WX765), .ZN(U6422_n1) );
  NOR2X0 U6422_U1 ( .IN1(n5369), .IN2(U6422_n1), .QN(WX828) );
  INVX0 U6423_U2 ( .INP(WX763), .ZN(U6423_n1) );
  NOR2X0 U6423_U1 ( .IN1(n5369), .IN2(U6423_n1), .QN(WX826) );
  INVX0 U6424_U2 ( .INP(WX761), .ZN(U6424_n1) );
  NOR2X0 U6424_U1 ( .IN1(n5369), .IN2(U6424_n1), .QN(WX824) );
  INVX0 U6425_U2 ( .INP(test_so5), .ZN(U6425_n1) );
  NOR2X0 U6425_U1 ( .IN1(n5369), .IN2(U6425_n1), .QN(WX822) );
  INVX0 U6426_U2 ( .INP(WX757), .ZN(U6426_n1) );
  NOR2X0 U6426_U1 ( .IN1(n5369), .IN2(U6426_n1), .QN(WX820) );
  INVX0 U6427_U2 ( .INP(WX755), .ZN(U6427_n1) );
  NOR2X0 U6427_U1 ( .IN1(n5368), .IN2(U6427_n1), .QN(WX818) );
  INVX0 U6428_U2 ( .INP(WX753), .ZN(U6428_n1) );
  NOR2X0 U6428_U1 ( .IN1(n5368), .IN2(U6428_n1), .QN(WX816) );
  INVX0 U6429_U2 ( .INP(WX751), .ZN(U6429_n1) );
  NOR2X0 U6429_U1 ( .IN1(n5368), .IN2(U6429_n1), .QN(WX814) );
  INVX0 U6430_U2 ( .INP(WX749), .ZN(U6430_n1) );
  NOR2X0 U6430_U1 ( .IN1(n5368), .IN2(U6430_n1), .QN(WX812) );
  INVX0 U6431_U2 ( .INP(WX747), .ZN(U6431_n1) );
  NOR2X0 U6431_U1 ( .IN1(n5368), .IN2(U6431_n1), .QN(WX810) );
  INVX0 U6432_U2 ( .INP(WX745), .ZN(U6432_n1) );
  NOR2X0 U6432_U1 ( .IN1(n5368), .IN2(U6432_n1), .QN(WX808) );
  INVX0 U6433_U2 ( .INP(WX743), .ZN(U6433_n1) );
  NOR2X0 U6433_U1 ( .IN1(n5368), .IN2(U6433_n1), .QN(WX806) );
  INVX0 U6434_U2 ( .INP(WX741), .ZN(U6434_n1) );
  NOR2X0 U6434_U1 ( .IN1(n5368), .IN2(U6434_n1), .QN(WX804) );
  INVX0 U6435_U2 ( .INP(WX739), .ZN(U6435_n1) );
  NOR2X0 U6435_U1 ( .IN1(n5368), .IN2(U6435_n1), .QN(WX802) );
  INVX0 U6436_U2 ( .INP(WX737), .ZN(U6436_n1) );
  NOR2X0 U6436_U1 ( .IN1(n5368), .IN2(U6436_n1), .QN(WX800) );
  INVX0 U6437_U2 ( .INP(WX735), .ZN(U6437_n1) );
  NOR2X0 U6437_U1 ( .IN1(n5368), .IN2(U6437_n1), .QN(WX798) );
  INVX0 U6438_U2 ( .INP(WX733), .ZN(U6438_n1) );
  NOR2X0 U6438_U1 ( .IN1(n5367), .IN2(U6438_n1), .QN(WX796) );
  INVX0 U6439_U2 ( .INP(WX731), .ZN(U6439_n1) );
  NOR2X0 U6439_U1 ( .IN1(n5367), .IN2(U6439_n1), .QN(WX794) );
  INVX0 U6440_U2 ( .INP(WX729), .ZN(U6440_n1) );
  NOR2X0 U6440_U1 ( .IN1(n5367), .IN2(U6440_n1), .QN(WX792) );
  INVX0 U6441_U2 ( .INP(WX727), .ZN(U6441_n1) );
  NOR2X0 U6441_U1 ( .IN1(n5367), .IN2(U6441_n1), .QN(WX790) );
  INVX0 U6442_U2 ( .INP(WX725), .ZN(U6442_n1) );
  NOR2X0 U6442_U1 ( .IN1(n5367), .IN2(U6442_n1), .QN(WX788) );
  INVX0 U6443_U2 ( .INP(test_so4), .ZN(U6443_n1) );
  NOR2X0 U6443_U1 ( .IN1(n5367), .IN2(U6443_n1), .QN(WX786) );
  INVX0 U6444_U2 ( .INP(WX721), .ZN(U6444_n1) );
  NOR2X0 U6444_U1 ( .IN1(n5367), .IN2(U6444_n1), .QN(WX784) );
  INVX0 U6445_U2 ( .INP(WX719), .ZN(U6445_n1) );
  NOR2X0 U6445_U1 ( .IN1(n5367), .IN2(U6445_n1), .QN(WX782) );
  INVX0 U6446_U2 ( .INP(WX717), .ZN(U6446_n1) );
  NOR2X0 U6446_U1 ( .IN1(n5367), .IN2(U6446_n1), .QN(WX780) );
  INVX0 U6447_U2 ( .INP(WX715), .ZN(U6447_n1) );
  NOR2X0 U6447_U1 ( .IN1(n5367), .IN2(U6447_n1), .QN(WX778) );
  INVX0 U6448_U2 ( .INP(WX713), .ZN(U6448_n1) );
  NOR2X0 U6448_U1 ( .IN1(n5367), .IN2(U6448_n1), .QN(WX776) );
  INVX0 U6449_U2 ( .INP(WX711), .ZN(U6449_n1) );
  NOR2X0 U6449_U1 ( .IN1(n5366), .IN2(U6449_n1), .QN(WX774) );
  INVX0 U6450_U2 ( .INP(WX709), .ZN(U6450_n1) );
  NOR2X0 U6450_U1 ( .IN1(n5366), .IN2(U6450_n1), .QN(WX772) );
  INVX0 U6451_U2 ( .INP(WX707), .ZN(U6451_n1) );
  NOR2X0 U6451_U1 ( .IN1(n5366), .IN2(U6451_n1), .QN(WX770) );
  INVX0 U6452_U2 ( .INP(WX705), .ZN(U6452_n1) );
  NOR2X0 U6452_U1 ( .IN1(n5366), .IN2(U6452_n1), .QN(WX768) );
  INVX0 U6453_U2 ( .INP(WX703), .ZN(U6453_n1) );
  NOR2X0 U6453_U1 ( .IN1(n5366), .IN2(U6453_n1), .QN(WX766) );
  INVX0 U6454_U2 ( .INP(WX701), .ZN(U6454_n1) );
  NOR2X0 U6454_U1 ( .IN1(n5366), .IN2(U6454_n1), .QN(WX764) );
  INVX0 U6455_U2 ( .INP(WX699), .ZN(U6455_n1) );
  NOR2X0 U6455_U1 ( .IN1(n5366), .IN2(U6455_n1), .QN(WX762) );
  INVX0 U6456_U2 ( .INP(WX697), .ZN(U6456_n1) );
  NOR2X0 U6456_U1 ( .IN1(n5366), .IN2(U6456_n1), .QN(WX760) );
  INVX0 U6457_U2 ( .INP(WX695), .ZN(U6457_n1) );
  NOR2X0 U6457_U1 ( .IN1(n5366), .IN2(U6457_n1), .QN(WX758) );
  INVX0 U6458_U2 ( .INP(WX693), .ZN(U6458_n1) );
  NOR2X0 U6458_U1 ( .IN1(n5366), .IN2(U6458_n1), .QN(WX756) );
  INVX0 U6459_U2 ( .INP(WX691), .ZN(U6459_n1) );
  NOR2X0 U6459_U1 ( .IN1(n5366), .IN2(U6459_n1), .QN(WX754) );
  INVX0 U6460_U2 ( .INP(WX689), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(n5365), .IN2(U6460_n1), .QN(WX752) );
  INVX0 U6461_U2 ( .INP(test_so3), .ZN(U6461_n1) );
  NOR2X0 U6461_U1 ( .IN1(n5365), .IN2(U6461_n1), .QN(WX750) );
  INVX0 U6462_U2 ( .INP(WX685), .ZN(U6462_n1) );
  NOR2X0 U6462_U1 ( .IN1(n5365), .IN2(U6462_n1), .QN(WX748) );
  INVX0 U6463_U2 ( .INP(WX683), .ZN(U6463_n1) );
  NOR2X0 U6463_U1 ( .IN1(n5365), .IN2(U6463_n1), .QN(WX746) );
  INVX0 U6464_U2 ( .INP(WX681), .ZN(U6464_n1) );
  NOR2X0 U6464_U1 ( .IN1(n5365), .IN2(U6464_n1), .QN(WX744) );
  INVX0 U6465_U2 ( .INP(WX679), .ZN(U6465_n1) );
  NOR2X0 U6465_U1 ( .IN1(n5365), .IN2(U6465_n1), .QN(WX742) );
  INVX0 U6466_U2 ( .INP(WX677), .ZN(U6466_n1) );
  NOR2X0 U6466_U1 ( .IN1(n5365), .IN2(U6466_n1), .QN(WX740) );
  INVX0 U6467_U2 ( .INP(WX675), .ZN(U6467_n1) );
  NOR2X0 U6467_U1 ( .IN1(n5365), .IN2(U6467_n1), .QN(WX738) );
  INVX0 U6468_U2 ( .INP(WX673), .ZN(U6468_n1) );
  NOR2X0 U6468_U1 ( .IN1(n5365), .IN2(U6468_n1), .QN(WX736) );
  INVX0 U6469_U2 ( .INP(WX671), .ZN(U6469_n1) );
  NOR2X0 U6469_U1 ( .IN1(n5365), .IN2(U6469_n1), .QN(WX734) );
  INVX0 U6470_U2 ( .INP(WX669), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n5365), .IN2(U6470_n1), .QN(WX732) );
  INVX0 U6471_U2 ( .INP(WX667), .ZN(U6471_n1) );
  NOR2X0 U6471_U1 ( .IN1(n5364), .IN2(U6471_n1), .QN(WX730) );
  INVX0 U6472_U2 ( .INP(WX665), .ZN(U6472_n1) );
  NOR2X0 U6472_U1 ( .IN1(n5364), .IN2(U6472_n1), .QN(WX728) );
  INVX0 U6473_U2 ( .INP(WX663), .ZN(U6473_n1) );
  NOR2X0 U6473_U1 ( .IN1(n5364), .IN2(U6473_n1), .QN(WX726) );
  INVX0 U6474_U2 ( .INP(WX661), .ZN(U6474_n1) );
  NOR2X0 U6474_U1 ( .IN1(n5364), .IN2(U6474_n1), .QN(WX724) );
  INVX0 U6475_U2 ( .INP(WX659), .ZN(U6475_n1) );
  NOR2X0 U6475_U1 ( .IN1(n5364), .IN2(U6475_n1), .QN(WX722) );
  INVX0 U6476_U2 ( .INP(WX657), .ZN(U6476_n1) );
  NOR2X0 U6476_U1 ( .IN1(n5364), .IN2(U6476_n1), .QN(WX720) );
  INVX0 U6477_U2 ( .INP(WX655), .ZN(U6477_n1) );
  NOR2X0 U6477_U1 ( .IN1(n5364), .IN2(U6477_n1), .QN(WX718) );
  INVX0 U6478_U2 ( .INP(WX653), .ZN(U6478_n1) );
  NOR2X0 U6478_U1 ( .IN1(n5364), .IN2(U6478_n1), .QN(WX716) );
  INVX0 U6479_U2 ( .INP(test_so2), .ZN(U6479_n1) );
  NOR2X0 U6479_U1 ( .IN1(n5364), .IN2(U6479_n1), .QN(WX714) );
  INVX0 U6480_U2 ( .INP(WX649), .ZN(U6480_n1) );
  NOR2X0 U6480_U1 ( .IN1(n5364), .IN2(U6480_n1), .QN(WX712) );
  INVX0 U6481_U2 ( .INP(WX647), .ZN(U6481_n1) );
  NOR2X0 U6481_U1 ( .IN1(n5364), .IN2(U6481_n1), .QN(WX710) );
  INVX0 U6482_U2 ( .INP(WX645), .ZN(U6482_n1) );
  NOR2X0 U6482_U1 ( .IN1(n5371), .IN2(U6482_n1), .QN(WX708) );
endmodule

