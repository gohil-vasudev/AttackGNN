module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n641_, new_n339_, new_n365_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n691_, new_n456_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n853_, new_n602_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n774_, new_n716_, new_n701_, new_n792_, new_n257_, new_n481_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n634_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n683_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n530_, new_n318_, new_n622_, new_n629_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n498_, new_n492_, new_n496_, new_n650_, new_n708_, new_n750_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n483_, new_n394_, new_n299_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n280_, new_n426_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n267_, new_n473_, new_n790_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n488_, new_n524_, new_n705_, new_n277_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n438_, new_n696_, new_n632_, new_n671_, new_n528_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n384_, new_n410_, new_n851_, new_n543_, new_n775_, new_n371_, new_n509_, new_n454_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n784_, new_n258_, new_n724_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n809_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n749_, new_n310_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n493_, new_n547_, new_n665_, new_n800_, new_n379_, new_n719_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n520_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n825_, new_n557_, new_n260_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n313_, new_n382_, new_n583_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n337_, new_n623_, new_n446_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n519_, new_n563_, new_n662_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n597_, new_n408_, new_n470_, new_n769_, new_n651_, new_n433_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n818_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n643_, new_n474_, new_n467_, new_n404_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n226_, new_n802_, new_n697_, new_n709_, new_n373_, new_n540_, new_n434_, new_n422_, new_n581_, new_n329_, new_n284_, new_n293_, new_n686_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n406_, new_n828_, new_n356_, new_n647_, new_n536_, new_n464_, new_n573_, new_n765_, new_n405_;

nand g000 ( new_n215_, N29, N42, N75 );
not g001 ( N388, new_n215_ );
nand g002 ( new_n217_, N29, N36, N80 );
not g003 ( N389, new_n217_ );
nand g004 ( new_n219_, N29, N36, N42 );
not g005 ( N390, new_n219_ );
nand g006 ( new_n221_, N85, N86 );
not g007 ( N391, new_n221_ );
nand g008 ( new_n223_, N1, N8, N13, N17 );
not g009 ( N418, new_n223_ );
not g010 ( new_n225_, N13 );
not g011 ( new_n226_, N17 );
nand g012 ( new_n227_, N1, N26 );
nor g013 ( new_n228_, new_n227_, new_n225_, new_n226_ );
nand g014 ( N419, new_n228_, new_n219_ );
nand g015 ( N420, N59, N75, N80 );
nand g016 ( N421, N36, N59, N80 );
nand g017 ( N422, N36, N42, N59 );
not g018 ( new_n233_, N90 );
nor g019 ( new_n234_, N87, N88 );
nor g020 ( N423, new_n234_, new_n233_ );
nand g021 ( N446, new_n228_, N390 );
not g022 ( new_n237_, keyIn_0_0 );
nand g023 ( new_n238_, N1, N26, N51 );
nand g024 ( new_n239_, new_n238_, new_n237_ );
nand g025 ( new_n240_, keyIn_0_0, N1, N26, N51 );
nand g026 ( new_n241_, new_n239_, new_n240_ );
not g027 ( N447, new_n241_ );
nand g028 ( new_n243_, N1, N8, N13, N55 );
nand g029 ( new_n244_, N29, N68 );
nor g030 ( N448, new_n243_, new_n244_ );
not g031 ( new_n246_, N74 );
nand g032 ( new_n247_, N59, N68 );
nor g033 ( new_n248_, new_n243_, new_n246_, new_n247_ );
xor g034 ( N449, new_n248_, keyIn_0_10 );
not g035 ( new_n250_, N89 );
nor g036 ( N450, new_n234_, new_n250_ );
not g037 ( new_n252_, N130 );
nor g038 ( new_n253_, N91, N96 );
nand g039 ( new_n254_, N91, N96 );
nand g040 ( new_n255_, new_n254_, keyIn_0_15 );
nor g041 ( new_n256_, new_n255_, new_n253_ );
xor g042 ( new_n257_, N101, N106 );
xnor g043 ( new_n258_, new_n256_, new_n257_ );
xnor g044 ( new_n259_, new_n258_, new_n252_ );
xnor g045 ( new_n260_, N111, N116 );
xnor g046 ( new_n261_, N121, N126 );
xnor g047 ( new_n262_, new_n260_, new_n261_ );
xnor g048 ( new_n263_, new_n262_, N135 );
xnor g049 ( N767, new_n259_, new_n263_ );
xnor g050 ( new_n265_, N159, N165 );
xnor g051 ( new_n266_, N171, N177 );
xnor g052 ( new_n267_, new_n265_, new_n266_ );
xnor g053 ( new_n268_, new_n267_, new_n252_ );
xnor g054 ( new_n269_, N183, N189 );
xnor g055 ( new_n270_, N195, N201 );
xnor g056 ( new_n271_, new_n269_, new_n270_ );
xnor g057 ( new_n272_, new_n271_, N207 );
xnor g058 ( N768, new_n268_, new_n272_ );
not g059 ( new_n274_, keyIn_0_60 );
not g060 ( new_n275_, keyIn_0_38 );
not g061 ( new_n276_, keyIn_0_14 );
nand g062 ( new_n277_, new_n241_, keyIn_0_8 );
not g063 ( new_n278_, keyIn_0_8 );
nand g064 ( new_n279_, new_n239_, new_n278_, new_n240_ );
nand g065 ( new_n280_, new_n277_, new_n279_ );
nand g066 ( new_n281_, new_n280_, new_n276_ );
nand g067 ( new_n282_, new_n277_, keyIn_0_14, new_n279_ );
nand g068 ( new_n283_, new_n281_, new_n282_ );
nand g069 ( new_n284_, N59, N156 );
xnor g070 ( new_n285_, new_n284_, keyIn_0_5 );
nand g071 ( new_n286_, new_n285_, N17 );
not g072 ( new_n287_, new_n286_ );
nand g073 ( new_n288_, new_n283_, keyIn_0_21, new_n287_ );
not g074 ( new_n289_, keyIn_0_21 );
nand g075 ( new_n290_, new_n283_, new_n287_ );
nand g076 ( new_n291_, new_n290_, new_n289_ );
nand g077 ( new_n292_, new_n291_, N1, new_n288_ );
nand g078 ( new_n293_, new_n292_, keyIn_0_25 );
not g079 ( new_n294_, keyIn_0_25 );
nand g080 ( new_n295_, new_n291_, new_n294_, N1, new_n288_ );
nand g081 ( new_n296_, new_n293_, new_n295_ );
nand g082 ( new_n297_, new_n296_, N153 );
nand g083 ( new_n298_, new_n297_, new_n275_ );
nand g084 ( new_n299_, new_n296_, keyIn_0_38, N153 );
nand g085 ( new_n300_, new_n298_, new_n299_ );
not g086 ( new_n301_, keyIn_0_13 );
nand g087 ( new_n302_, N17, N42 );
nand g088 ( new_n303_, new_n302_, keyIn_0_7 );
not g089 ( new_n304_, N42 );
nand g090 ( new_n305_, new_n226_, new_n304_ );
nand g091 ( new_n306_, new_n305_, keyIn_0_6 );
nor g092 ( new_n307_, keyIn_0_6, N17, N42 );
nor g093 ( new_n308_, new_n302_, keyIn_0_7 );
nor g094 ( new_n309_, new_n308_, new_n307_ );
nand g095 ( new_n310_, new_n309_, new_n301_, new_n303_, new_n306_ );
not g096 ( new_n311_, keyIn_0_6 );
nand g097 ( new_n312_, new_n311_, new_n226_, new_n304_ );
not g098 ( new_n313_, keyIn_0_7 );
nand g099 ( new_n314_, new_n313_, N17, N42 );
nand g100 ( new_n315_, new_n306_, new_n303_, new_n312_, new_n314_ );
nand g101 ( new_n316_, new_n315_, keyIn_0_13 );
nand g102 ( new_n317_, new_n316_, new_n310_, N59, N156 );
not g103 ( new_n318_, new_n317_ );
nand g104 ( new_n319_, new_n318_, new_n283_ );
nand g105 ( new_n320_, new_n319_, keyIn_0_20 );
not g106 ( new_n321_, keyIn_0_20 );
nand g107 ( new_n322_, new_n318_, new_n283_, new_n321_ );
not g108 ( new_n323_, keyIn_0_16 );
not g109 ( new_n324_, keyIn_0_1 );
nand g110 ( new_n325_, N1, N8, N17, N51 );
xnor g111 ( new_n326_, new_n325_, new_n324_ );
nand g112 ( new_n327_, new_n326_, keyIn_0_9 );
not g113 ( new_n328_, keyIn_0_9 );
xnor g114 ( new_n329_, new_n325_, keyIn_0_1 );
nand g115 ( new_n330_, new_n329_, new_n328_ );
nand g116 ( new_n331_, new_n327_, new_n330_ );
nand g117 ( new_n332_, N42, N59, N75 );
xnor g118 ( new_n333_, new_n332_, keyIn_0_3 );
xnor g119 ( new_n334_, new_n333_, keyIn_0_11 );
nand g120 ( new_n335_, new_n334_, new_n331_ );
nand g121 ( new_n336_, new_n335_, new_n323_ );
nand g122 ( new_n337_, new_n334_, new_n331_, keyIn_0_16 );
nand g123 ( new_n338_, new_n336_, new_n337_ );
nand g124 ( new_n339_, new_n338_, new_n320_, keyIn_0_22, new_n322_ );
not g125 ( new_n340_, keyIn_0_22 );
nand g126 ( new_n341_, new_n338_, new_n320_, new_n322_ );
nand g127 ( new_n342_, new_n341_, new_n340_ );
nand g128 ( new_n343_, new_n342_, N126, new_n339_ );
nand g129 ( new_n344_, new_n343_, keyIn_0_39 );
not g130 ( new_n345_, keyIn_0_39 );
nand g131 ( new_n346_, new_n342_, new_n345_, N126, new_n339_ );
nand g132 ( new_n347_, new_n344_, new_n346_ );
nand g133 ( new_n348_, new_n300_, new_n347_ );
nand g134 ( new_n349_, new_n348_, keyIn_0_45 );
not g135 ( new_n350_, keyIn_0_45 );
nand g136 ( new_n351_, new_n300_, new_n350_, new_n347_ );
nand g137 ( new_n352_, new_n349_, new_n351_ );
nand g138 ( new_n353_, N29, N75, N80 );
xor g139 ( new_n354_, new_n353_, keyIn_0_2 );
nand g140 ( new_n355_, new_n283_, new_n354_ );
not g141 ( new_n356_, new_n355_ );
nand g142 ( new_n357_, new_n356_, N55 );
xnor g143 ( new_n358_, new_n357_, keyIn_0_19 );
xnor g144 ( new_n359_, keyIn_0_4, N268 );
xor g145 ( new_n360_, new_n359_, keyIn_0_12 );
nand g146 ( new_n361_, new_n358_, new_n360_ );
xnor g147 ( new_n362_, new_n361_, keyIn_0_29 );
nand g148 ( new_n363_, new_n352_, new_n362_ );
nand g149 ( new_n364_, new_n363_, keyIn_0_50 );
not g150 ( new_n365_, keyIn_0_50 );
nand g151 ( new_n366_, new_n352_, new_n365_, new_n362_ );
nand g152 ( new_n367_, new_n364_, new_n366_ );
nand g153 ( new_n368_, new_n367_, N201 );
nand g154 ( new_n369_, new_n368_, new_n274_ );
nand g155 ( new_n370_, new_n367_, keyIn_0_60, N201 );
nand g156 ( new_n371_, new_n369_, new_n370_ );
not g157 ( new_n372_, new_n371_ );
not g158 ( new_n373_, N201 );
nand g159 ( new_n374_, new_n364_, new_n373_, new_n366_ );
nand g160 ( new_n375_, new_n374_, keyIn_0_61 );
not g161 ( new_n376_, keyIn_0_61 );
nand g162 ( new_n377_, new_n364_, new_n376_, new_n373_, new_n366_ );
nand g163 ( new_n378_, new_n375_, new_n377_ );
nand g164 ( new_n379_, new_n372_, new_n378_ );
not g165 ( new_n380_, new_n379_ );
nand g166 ( new_n381_, new_n380_, N261 );
not g167 ( new_n382_, N261 );
nand g168 ( new_n383_, new_n379_, new_n382_ );
nand g169 ( new_n384_, new_n381_, N219, new_n383_ );
nand g170 ( new_n385_, new_n371_, keyIn_0_67 );
not g171 ( new_n386_, keyIn_0_67 );
nand g172 ( new_n387_, new_n369_, new_n386_, new_n370_ );
nand g173 ( new_n388_, new_n385_, new_n387_ );
nand g174 ( new_n389_, new_n388_, N237 );
nand g175 ( new_n390_, new_n380_, N228 );
nand g176 ( new_n391_, new_n367_, N246 );
nand g177 ( new_n392_, N42, N72, N73 );
nor g178 ( new_n393_, new_n243_, new_n392_, new_n247_ );
nand g179 ( new_n394_, new_n393_, N201 );
nand g180 ( new_n395_, N121, N210 );
nand g181 ( new_n396_, N255, N267 );
nand g182 ( new_n397_, new_n391_, new_n394_, new_n395_, new_n396_ );
not g183 ( new_n398_, new_n397_ );
nand g184 ( N850, new_n384_, new_n389_, new_n390_, new_n398_ );
not g185 ( new_n400_, keyIn_0_80 );
not g186 ( new_n401_, keyIn_0_77 );
xnor g187 ( new_n402_, new_n341_, keyIn_0_22 );
nand g188 ( new_n403_, new_n402_, N111 );
xor g189 ( new_n404_, new_n403_, keyIn_0_33 );
nand g190 ( new_n405_, new_n296_, N143 );
xnor g191 ( new_n406_, new_n405_, keyIn_0_32 );
nand g192 ( new_n407_, new_n404_, new_n406_ );
xnor g193 ( new_n408_, new_n407_, keyIn_0_42 );
xor g194 ( new_n409_, new_n361_, keyIn_0_26 );
nand g195 ( new_n410_, new_n408_, new_n409_ );
xor g196 ( new_n411_, new_n410_, keyIn_0_47 );
nand g197 ( new_n412_, new_n411_, N183 );
xnor g198 ( new_n413_, new_n412_, keyIn_0_54 );
not g199 ( new_n414_, N183 );
not g200 ( new_n415_, new_n411_ );
nand g201 ( new_n416_, new_n415_, new_n414_ );
xor g202 ( new_n417_, new_n416_, keyIn_0_55 );
nand g203 ( new_n418_, new_n417_, new_n413_ );
not g204 ( new_n419_, new_n418_ );
not g205 ( new_n420_, keyIn_0_75 );
not g206 ( new_n421_, N195 );
not g207 ( new_n422_, keyIn_0_49 );
nand g208 ( new_n423_, new_n296_, N149 );
nand g209 ( new_n424_, new_n423_, keyIn_0_36 );
not g210 ( new_n425_, keyIn_0_36 );
nand g211 ( new_n426_, new_n296_, new_n425_, N149 );
nand g212 ( new_n427_, new_n424_, new_n426_ );
nand g213 ( new_n428_, new_n342_, N121, new_n339_ );
nand g214 ( new_n429_, new_n428_, keyIn_0_37 );
not g215 ( new_n430_, keyIn_0_37 );
nand g216 ( new_n431_, new_n342_, new_n430_, N121, new_n339_ );
nand g217 ( new_n432_, new_n429_, new_n431_ );
nand g218 ( new_n433_, new_n427_, keyIn_0_44, new_n432_ );
xor g219 ( new_n434_, new_n361_, keyIn_0_28 );
not g220 ( new_n435_, keyIn_0_44 );
nand g221 ( new_n436_, new_n427_, new_n432_ );
nand g222 ( new_n437_, new_n436_, new_n435_ );
nand g223 ( new_n438_, new_n437_, new_n433_, new_n434_ );
nand g224 ( new_n439_, new_n438_, new_n422_ );
nand g225 ( new_n440_, new_n437_, keyIn_0_49, new_n433_, new_n434_ );
nand g226 ( new_n441_, new_n439_, new_n440_ );
nand g227 ( new_n442_, new_n441_, new_n421_ );
nand g228 ( new_n443_, new_n442_, keyIn_0_59 );
not g229 ( new_n444_, keyIn_0_59 );
nand g230 ( new_n445_, new_n441_, new_n444_, new_n421_ );
nand g231 ( new_n446_, new_n443_, new_n445_ );
not g232 ( new_n447_, N189 );
not g233 ( new_n448_, keyIn_0_43 );
not g234 ( new_n449_, keyIn_0_35 );
nand g235 ( new_n450_, new_n342_, N116, new_n339_ );
nand g236 ( new_n451_, new_n450_, new_n449_ );
nand g237 ( new_n452_, new_n342_, keyIn_0_35, N116, new_n339_ );
nand g238 ( new_n453_, new_n451_, new_n452_ );
nand g239 ( new_n454_, new_n296_, N146 );
nand g240 ( new_n455_, new_n454_, keyIn_0_34 );
not g241 ( new_n456_, keyIn_0_34 );
nand g242 ( new_n457_, new_n296_, new_n456_, N146 );
nand g243 ( new_n458_, new_n453_, new_n448_, new_n455_, new_n457_ );
xnor g244 ( new_n459_, new_n361_, keyIn_0_27 );
nand g245 ( new_n460_, new_n453_, new_n455_, new_n457_ );
nand g246 ( new_n461_, new_n460_, keyIn_0_43 );
nand g247 ( new_n462_, new_n461_, new_n458_, new_n459_ );
nand g248 ( new_n463_, new_n462_, keyIn_0_48 );
not g249 ( new_n464_, keyIn_0_48 );
nand g250 ( new_n465_, new_n461_, new_n458_, new_n464_, new_n459_ );
nand g251 ( new_n466_, new_n463_, new_n447_, new_n465_ );
xnor g252 ( new_n467_, new_n466_, keyIn_0_57 );
nand g253 ( new_n468_, new_n446_, new_n467_ );
not g254 ( new_n469_, new_n468_ );
nand g255 ( new_n470_, new_n388_, new_n469_ );
nand g256 ( new_n471_, new_n470_, keyIn_0_73 );
not g257 ( new_n472_, keyIn_0_73 );
nand g258 ( new_n473_, new_n388_, new_n472_, new_n469_ );
nand g259 ( new_n474_, new_n471_, new_n473_ );
nand g260 ( new_n475_, new_n439_, N195, new_n440_ );
xnor g261 ( new_n476_, new_n475_, keyIn_0_58 );
xnor g262 ( new_n477_, new_n476_, keyIn_0_66 );
nand g263 ( new_n478_, new_n477_, new_n467_ );
nand g264 ( new_n479_, new_n478_, keyIn_0_72 );
not g265 ( new_n480_, keyIn_0_72 );
nand g266 ( new_n481_, new_n477_, new_n480_, new_n467_ );
nand g267 ( new_n482_, new_n479_, new_n481_ );
nand g268 ( new_n483_, new_n378_, new_n446_, new_n467_, N261 );
xnor g269 ( new_n484_, new_n483_, keyIn_0_68 );
not g270 ( new_n485_, keyIn_0_65 );
nand g271 ( new_n486_, new_n463_, new_n465_ );
nand g272 ( new_n487_, new_n486_, N189 );
nand g273 ( new_n488_, new_n487_, keyIn_0_56 );
not g274 ( new_n489_, keyIn_0_56 );
nand g275 ( new_n490_, new_n486_, new_n489_, N189 );
nand g276 ( new_n491_, new_n488_, new_n490_ );
nand g277 ( new_n492_, new_n491_, new_n485_ );
nand g278 ( new_n493_, new_n488_, keyIn_0_65, new_n490_ );
nand g279 ( new_n494_, new_n492_, new_n493_ );
nand g280 ( new_n495_, new_n494_, keyIn_0_71 );
not g281 ( new_n496_, keyIn_0_71 );
nand g282 ( new_n497_, new_n492_, new_n496_, new_n493_ );
nand g283 ( new_n498_, new_n495_, new_n497_ );
nor g284 ( new_n499_, new_n484_, new_n498_ );
nand g285 ( new_n500_, new_n474_, new_n482_, new_n499_ );
nand g286 ( new_n501_, new_n500_, new_n420_ );
nand g287 ( new_n502_, new_n474_, new_n499_, new_n482_, keyIn_0_75 );
nand g288 ( new_n503_, new_n501_, new_n502_ );
not g289 ( new_n504_, new_n503_ );
nand g290 ( new_n505_, new_n504_, new_n419_ );
nand g291 ( new_n506_, new_n505_, new_n401_ );
nand g292 ( new_n507_, new_n503_, keyIn_0_76, new_n418_ );
not g293 ( new_n508_, keyIn_0_76 );
nand g294 ( new_n509_, new_n503_, new_n418_ );
nand g295 ( new_n510_, new_n509_, new_n508_ );
nand g296 ( new_n511_, new_n504_, keyIn_0_77, new_n419_ );
nand g297 ( new_n512_, new_n506_, new_n507_, new_n510_, new_n511_ );
not g298 ( new_n513_, new_n512_ );
nand g299 ( new_n514_, new_n513_, new_n400_ );
nand g300 ( new_n515_, new_n512_, keyIn_0_80 );
nand g301 ( new_n516_, new_n514_, keyIn_0_83, N219, new_n515_ );
nand g302 ( new_n517_, N106, N210 );
not g303 ( new_n518_, keyIn_0_83 );
nand g304 ( new_n519_, new_n514_, N219, new_n515_ );
nand g305 ( new_n520_, new_n519_, new_n518_ );
nand g306 ( new_n521_, new_n520_, new_n516_, new_n517_ );
xor g307 ( new_n522_, new_n521_, keyIn_0_92 );
xor g308 ( new_n523_, new_n413_, keyIn_0_64 );
not g309 ( new_n524_, new_n523_ );
nand g310 ( new_n525_, new_n524_, N237 );
nand g311 ( new_n526_, new_n419_, N228 );
nand g312 ( new_n527_, new_n393_, N183 );
nand g313 ( new_n528_, new_n411_, N246 );
nand g314 ( new_n529_, new_n526_, new_n527_, new_n528_ );
not g315 ( new_n530_, new_n529_ );
nand g316 ( new_n531_, new_n522_, new_n525_, new_n530_ );
xor g317 ( new_n532_, new_n531_, keyIn_0_100 );
xnor g318 ( new_n533_, new_n532_, keyIn_0_106 );
xnor g319 ( N863, new_n533_, keyIn_0_112 );
not g320 ( new_n535_, new_n491_ );
nand g321 ( new_n536_, new_n535_, new_n467_ );
not g322 ( new_n537_, new_n536_ );
not g323 ( new_n538_, new_n477_ );
not g324 ( new_n539_, new_n388_ );
nand g325 ( new_n540_, new_n378_, N261 );
nand g326 ( new_n541_, new_n539_, new_n540_ );
nand g327 ( new_n542_, new_n541_, new_n446_ );
nand g328 ( new_n543_, new_n542_, new_n538_ );
nand g329 ( new_n544_, new_n543_, new_n537_ );
nand g330 ( new_n545_, new_n542_, new_n538_, new_n536_ );
nand g331 ( new_n546_, new_n544_, N219, new_n545_ );
nand g332 ( new_n547_, new_n492_, N237, new_n493_ );
nand g333 ( new_n548_, new_n537_, N228 );
nand g334 ( new_n549_, new_n486_, N246 );
nand g335 ( new_n550_, new_n393_, N189 );
nand g336 ( new_n551_, N111, N210 );
nand g337 ( new_n552_, N255, N259 );
nand g338 ( new_n553_, new_n549_, new_n550_, new_n551_, new_n552_ );
not g339 ( new_n554_, new_n553_ );
nand g340 ( N864, new_n546_, new_n547_, new_n548_, new_n554_ );
nand g341 ( new_n556_, new_n446_, new_n476_ );
not g342 ( new_n557_, new_n556_ );
nand g343 ( new_n558_, new_n541_, new_n557_ );
nand g344 ( new_n559_, new_n539_, new_n540_, new_n556_ );
nand g345 ( new_n560_, new_n558_, keyIn_0_84, N219, new_n559_ );
not g346 ( new_n561_, keyIn_0_84 );
nand g347 ( new_n562_, new_n558_, N219, new_n559_ );
nand g348 ( new_n563_, new_n562_, new_n561_ );
nand g349 ( new_n564_, new_n477_, N237 );
nand g350 ( new_n565_, new_n557_, N228 );
nand g351 ( new_n566_, new_n439_, N246, new_n440_ );
nand g352 ( new_n567_, new_n393_, N195 );
nand g353 ( new_n568_, N255, N260 );
nand g354 ( new_n569_, N116, N210 );
nand g355 ( new_n570_, new_n568_, new_n569_ );
not g356 ( new_n571_, new_n570_ );
nand g357 ( new_n572_, new_n565_, new_n566_, new_n567_, new_n571_ );
not g358 ( new_n573_, new_n572_ );
nand g359 ( N865, new_n563_, new_n560_, new_n564_, new_n573_ );
not g360 ( new_n575_, keyIn_0_88 );
not g361 ( new_n576_, keyIn_0_87 );
nand g362 ( new_n577_, new_n402_, N96 );
not g363 ( new_n578_, new_n359_ );
nand g364 ( new_n579_, new_n356_, keyIn_0_18, N17 );
not g365 ( new_n580_, keyIn_0_18 );
nand g366 ( new_n581_, new_n356_, N17 );
nand g367 ( new_n582_, new_n581_, new_n580_ );
nand g368 ( new_n583_, new_n582_, new_n578_, new_n579_ );
nand g369 ( new_n584_, new_n283_, N55, new_n285_ );
xor g370 ( new_n585_, new_n584_, keyIn_0_17 );
nand g371 ( new_n586_, new_n585_, N146 );
nand g372 ( new_n587_, N51, N138 );
nand g373 ( new_n588_, new_n577_, new_n583_, new_n586_, new_n587_ );
nor g374 ( new_n589_, new_n588_, N165 );
not g375 ( new_n590_, new_n589_ );
nand g376 ( new_n591_, new_n402_, N101 );
nand g377 ( new_n592_, new_n585_, N149 );
nand g378 ( new_n593_, N17, N138 );
nand g379 ( new_n594_, new_n591_, new_n583_, new_n592_, new_n593_ );
nor g380 ( new_n595_, new_n594_, N171 );
not g381 ( new_n596_, new_n595_ );
nand g382 ( new_n597_, new_n590_, new_n596_ );
not g383 ( new_n598_, new_n597_ );
not g384 ( new_n599_, N177 );
nand g385 ( new_n600_, new_n402_, keyIn_0_30, N106 );
not g386 ( new_n601_, keyIn_0_30 );
nand g387 ( new_n602_, new_n402_, N106 );
nand g388 ( new_n603_, new_n602_, new_n601_ );
nand g389 ( new_n604_, N138, N152 );
nand g390 ( new_n605_, new_n603_, new_n600_, new_n604_ );
xor g391 ( new_n606_, new_n605_, keyIn_0_41 );
nand g392 ( new_n607_, new_n585_, N153 );
xnor g393 ( new_n608_, new_n607_, keyIn_0_23 );
xnor g394 ( new_n609_, new_n583_, keyIn_0_24 );
nand g395 ( new_n610_, new_n608_, new_n609_ );
xor g396 ( new_n611_, new_n610_, keyIn_0_31 );
nand g397 ( new_n612_, new_n606_, new_n611_ );
xor g398 ( new_n613_, new_n612_, keyIn_0_46 );
nand g399 ( new_n614_, new_n613_, new_n599_ );
xor g400 ( new_n615_, new_n614_, keyIn_0_53 );
not g401 ( new_n616_, keyIn_0_78 );
nand g402 ( new_n617_, new_n501_, new_n417_, new_n502_ );
nand g403 ( new_n618_, new_n617_, new_n616_ );
nand g404 ( new_n619_, new_n501_, keyIn_0_78, new_n417_, new_n502_ );
nand g405 ( new_n620_, new_n618_, new_n619_ );
not g406 ( new_n621_, keyIn_0_70 );
xnor g407 ( new_n622_, new_n523_, new_n621_ );
nand g408 ( new_n623_, new_n620_, new_n622_ );
xnor g409 ( new_n624_, new_n623_, keyIn_0_79 );
nand g410 ( new_n625_, new_n624_, new_n576_, new_n598_, new_n615_ );
not g411 ( new_n626_, keyIn_0_79 );
nand g412 ( new_n627_, new_n623_, new_n626_ );
nand g413 ( new_n628_, new_n620_, keyIn_0_79, new_n622_ );
nand g414 ( new_n629_, new_n627_, new_n598_, new_n615_, new_n628_ );
nand g415 ( new_n630_, new_n629_, keyIn_0_87 );
not g416 ( new_n631_, new_n613_ );
nand g417 ( new_n632_, new_n631_, N177 );
xnor g418 ( new_n633_, new_n632_, keyIn_0_52 );
xor g419 ( new_n634_, new_n633_, keyIn_0_63 );
not g420 ( new_n635_, new_n634_ );
nand g421 ( new_n636_, new_n635_, keyIn_0_74, new_n598_ );
not g422 ( new_n637_, keyIn_0_74 );
nand g423 ( new_n638_, new_n635_, new_n598_ );
nand g424 ( new_n639_, new_n638_, new_n637_ );
nand g425 ( new_n640_, new_n594_, N171 );
not g426 ( new_n641_, new_n640_ );
nand g427 ( new_n642_, new_n590_, new_n641_ );
nand g428 ( new_n643_, new_n588_, N165 );
nand g429 ( new_n644_, new_n639_, new_n636_, new_n642_, new_n643_ );
not g430 ( new_n645_, new_n644_ );
nand g431 ( new_n646_, new_n625_, new_n630_, new_n645_ );
nand g432 ( new_n647_, new_n646_, new_n575_ );
nand g433 ( new_n648_, new_n625_, keyIn_0_88, new_n630_, new_n645_ );
nand g434 ( new_n649_, new_n647_, new_n648_ );
not g435 ( new_n650_, N159 );
nand g436 ( new_n651_, new_n402_, N91 );
nand g437 ( new_n652_, N8, N138 );
nand g438 ( new_n653_, new_n651_, keyIn_0_40, new_n652_ );
not g439 ( new_n654_, keyIn_0_40 );
nand g440 ( new_n655_, new_n651_, new_n652_ );
nand g441 ( new_n656_, new_n655_, new_n654_ );
nand g442 ( new_n657_, new_n585_, N143 );
nand g443 ( new_n658_, new_n657_, new_n583_ );
not g444 ( new_n659_, new_n658_ );
nand g445 ( new_n660_, new_n656_, new_n650_, new_n653_, new_n659_ );
nand g446 ( new_n661_, new_n649_, keyIn_0_101, new_n660_ );
not g447 ( new_n662_, keyIn_0_101 );
nand g448 ( new_n663_, new_n649_, new_n660_ );
nand g449 ( new_n664_, new_n663_, new_n662_ );
nand g450 ( new_n665_, new_n656_, new_n653_, new_n659_ );
nand g451 ( new_n666_, new_n665_, N159 );
xor g452 ( new_n667_, new_n666_, keyIn_0_51 );
nand g453 ( new_n668_, new_n664_, new_n661_, new_n667_ );
xor g454 ( new_n669_, new_n668_, keyIn_0_107 );
xnor g455 ( N866, new_n669_, keyIn_0_113 );
not g456 ( new_n671_, keyIn_0_91 );
nand g457 ( new_n672_, new_n627_, new_n628_ );
nand g458 ( new_n673_, new_n633_, new_n615_ );
nand g459 ( new_n674_, new_n672_, new_n673_ );
xnor g460 ( new_n675_, new_n674_, keyIn_0_81 );
not g461 ( new_n676_, keyIn_0_82 );
not g462 ( new_n677_, new_n673_ );
nand g463 ( new_n678_, new_n624_, new_n677_ );
xnor g464 ( new_n679_, new_n678_, new_n676_ );
nand g465 ( new_n680_, new_n679_, new_n675_ );
nand g466 ( new_n681_, new_n680_, new_n671_ );
nand g467 ( new_n682_, new_n679_, keyIn_0_91, new_n675_ );
nand g468 ( new_n683_, new_n681_, keyIn_0_99, N219, new_n682_ );
nand g469 ( new_n684_, N101, N210 );
not g470 ( new_n685_, keyIn_0_99 );
nand g471 ( new_n686_, new_n681_, N219, new_n682_ );
nand g472 ( new_n687_, new_n686_, new_n685_ );
nand g473 ( new_n688_, new_n687_, new_n683_, new_n684_ );
xnor g474 ( new_n689_, new_n688_, keyIn_0_105 );
not g475 ( new_n690_, keyIn_0_69 );
nand g476 ( new_n691_, new_n635_, new_n690_, N237 );
nand g477 ( new_n692_, new_n635_, N237 );
nand g478 ( new_n693_, new_n692_, keyIn_0_69 );
nand g479 ( new_n694_, new_n677_, N228 );
nand g480 ( new_n695_, new_n631_, N246 );
nand g481 ( new_n696_, new_n393_, N177 );
nand g482 ( new_n697_, new_n694_, new_n695_, new_n696_ );
not g483 ( new_n698_, new_n697_ );
nand g484 ( new_n699_, new_n689_, new_n691_, new_n693_, new_n698_ );
xor g485 ( new_n700_, new_n699_, keyIn_0_111 );
xnor g486 ( new_n701_, new_n700_, keyIn_0_117 );
xnor g487 ( N874, new_n701_, keyIn_0_121 );
not g488 ( new_n703_, keyIn_0_118 );
not g489 ( new_n704_, keyIn_0_102 );
nand g490 ( new_n705_, new_n667_, new_n660_ );
xnor g491 ( new_n706_, new_n705_, keyIn_0_62 );
not g492 ( new_n707_, new_n706_ );
nand g493 ( new_n708_, new_n649_, new_n707_ );
nand g494 ( new_n709_, new_n708_, keyIn_0_94 );
not g495 ( new_n710_, keyIn_0_94 );
nand g496 ( new_n711_, new_n649_, new_n710_, new_n707_ );
nand g497 ( new_n712_, new_n709_, new_n711_ );
nand g498 ( new_n713_, new_n647_, new_n648_, new_n706_ );
xnor g499 ( new_n714_, new_n713_, keyIn_0_93 );
nand g500 ( new_n715_, new_n712_, new_n714_ );
nand g501 ( new_n716_, new_n715_, new_n704_ );
nand g502 ( new_n717_, new_n712_, new_n714_, keyIn_0_102 );
nand g503 ( new_n718_, new_n716_, keyIn_0_108, N219, new_n717_ );
not g504 ( new_n719_, new_n360_ );
nand g505 ( new_n720_, new_n719_, N210 );
not g506 ( new_n721_, keyIn_0_108 );
nand g507 ( new_n722_, new_n716_, N219, new_n717_ );
nand g508 ( new_n723_, new_n722_, new_n721_ );
nand g509 ( new_n724_, new_n723_, new_n718_, new_n720_ );
nand g510 ( new_n725_, new_n724_, keyIn_0_114 );
not g511 ( new_n726_, keyIn_0_114 );
nand g512 ( new_n727_, new_n723_, new_n726_, new_n718_, new_n720_ );
nand g513 ( new_n728_, new_n725_, new_n727_ );
nand g514 ( new_n729_, new_n707_, N228 );
not g515 ( new_n730_, new_n667_ );
nand g516 ( new_n731_, new_n730_, N237 );
nand g517 ( new_n732_, new_n393_, N159 );
nand g518 ( new_n733_, new_n665_, N246 );
nand g519 ( new_n734_, new_n729_, new_n731_, new_n732_, new_n733_ );
not g520 ( new_n735_, new_n734_ );
nand g521 ( new_n736_, new_n728_, new_n735_ );
nand g522 ( new_n737_, new_n736_, new_n703_ );
nand g523 ( new_n738_, new_n728_, keyIn_0_118, new_n735_ );
nand g524 ( new_n739_, new_n737_, new_n738_ );
nand g525 ( new_n740_, new_n739_, keyIn_0_122 );
not g526 ( new_n741_, keyIn_0_122 );
nand g527 ( new_n742_, new_n737_, new_n741_, new_n738_ );
nand g528 ( new_n743_, new_n740_, new_n742_ );
nand g529 ( new_n744_, new_n743_, keyIn_0_125 );
not g530 ( new_n745_, keyIn_0_125 );
nand g531 ( new_n746_, new_n740_, new_n745_, new_n742_ );
nand g532 ( N878, new_n744_, new_n746_ );
not g533 ( new_n748_, keyIn_0_119 );
not g534 ( new_n749_, keyIn_0_115 );
not g535 ( new_n750_, keyIn_0_103 );
not g536 ( new_n751_, new_n643_ );
nor g537 ( new_n752_, new_n751_, new_n589_ );
not g538 ( new_n753_, new_n752_ );
not g539 ( new_n754_, keyIn_0_89 );
not g540 ( new_n755_, keyIn_0_86 );
nand g541 ( new_n756_, new_n624_, new_n755_, new_n596_, new_n615_ );
nand g542 ( new_n757_, new_n627_, new_n596_, new_n615_, new_n628_ );
nand g543 ( new_n758_, new_n757_, keyIn_0_86 );
nand g544 ( new_n759_, new_n635_, new_n596_ );
nand g545 ( new_n760_, new_n759_, new_n640_ );
not g546 ( new_n761_, new_n760_ );
nand g547 ( new_n762_, new_n756_, new_n758_, new_n761_ );
nand g548 ( new_n763_, new_n762_, new_n754_ );
nand g549 ( new_n764_, new_n756_, keyIn_0_89, new_n758_, new_n761_ );
nand g550 ( new_n765_, new_n763_, new_n764_ );
nand g551 ( new_n766_, new_n765_, new_n753_ );
nand g552 ( new_n767_, new_n766_, keyIn_0_95 );
not g553 ( new_n768_, keyIn_0_95 );
nand g554 ( new_n769_, new_n765_, new_n768_, new_n753_ );
nand g555 ( new_n770_, new_n767_, new_n769_ );
not g556 ( new_n771_, keyIn_0_96 );
nand g557 ( new_n772_, new_n763_, new_n752_, new_n764_ );
xnor g558 ( new_n773_, new_n772_, new_n771_ );
nand g559 ( new_n774_, new_n770_, new_n773_ );
nand g560 ( new_n775_, new_n774_, new_n750_ );
nand g561 ( new_n776_, new_n770_, new_n773_, keyIn_0_103 );
nand g562 ( new_n777_, new_n775_, new_n776_ );
nand g563 ( new_n778_, new_n777_, keyIn_0_109, N219 );
nand g564 ( new_n779_, N91, N210 );
not g565 ( new_n780_, keyIn_0_109 );
nand g566 ( new_n781_, new_n777_, N219 );
nand g567 ( new_n782_, new_n781_, new_n780_ );
nand g568 ( new_n783_, new_n782_, new_n749_, new_n778_, new_n779_ );
nand g569 ( new_n784_, new_n782_, new_n778_, new_n779_ );
nand g570 ( new_n785_, new_n784_, keyIn_0_115 );
nand g571 ( new_n786_, new_n752_, N228 );
not g572 ( new_n787_, new_n786_ );
nand g573 ( new_n788_, new_n751_, N237 );
nand g574 ( new_n789_, new_n393_, N165 );
nand g575 ( new_n790_, new_n588_, N246 );
nand g576 ( new_n791_, new_n788_, new_n789_, new_n790_ );
nor g577 ( new_n792_, new_n787_, new_n791_ );
nand g578 ( new_n793_, new_n785_, new_n783_, new_n792_ );
nand g579 ( new_n794_, new_n793_, new_n748_ );
nand g580 ( new_n795_, new_n785_, keyIn_0_119, new_n783_, new_n792_ );
nand g581 ( new_n796_, new_n794_, new_n795_ );
nand g582 ( new_n797_, new_n796_, keyIn_0_123 );
not g583 ( new_n798_, keyIn_0_123 );
nand g584 ( new_n799_, new_n794_, new_n798_, new_n795_ );
nand g585 ( new_n800_, new_n797_, new_n799_ );
nand g586 ( new_n801_, new_n800_, keyIn_0_126 );
not g587 ( new_n802_, keyIn_0_126 );
nand g588 ( new_n803_, new_n797_, new_n802_, new_n799_ );
nand g589 ( N879, new_n801_, new_n803_ );
not g590 ( new_n805_, keyIn_0_120 );
not g591 ( new_n806_, keyIn_0_110 );
not g592 ( new_n807_, keyIn_0_104 );
nor g593 ( new_n808_, new_n641_, new_n595_ );
nand g594 ( new_n809_, new_n624_, keyIn_0_85, new_n615_ );
not g595 ( new_n810_, keyIn_0_85 );
nand g596 ( new_n811_, new_n624_, new_n615_ );
nand g597 ( new_n812_, new_n811_, new_n810_ );
nand g598 ( new_n813_, new_n812_, new_n634_, new_n809_ );
nand g599 ( new_n814_, new_n813_, keyIn_0_90 );
not g600 ( new_n815_, keyIn_0_90 );
nand g601 ( new_n816_, new_n812_, new_n815_, new_n634_, new_n809_ );
nand g602 ( new_n817_, new_n814_, new_n808_, new_n816_ );
nand g603 ( new_n818_, new_n817_, keyIn_0_98 );
not g604 ( new_n819_, keyIn_0_97 );
not g605 ( new_n820_, new_n808_ );
nand g606 ( new_n821_, new_n814_, new_n816_ );
nand g607 ( new_n822_, new_n821_, new_n819_, new_n820_ );
nand g608 ( new_n823_, new_n818_, new_n822_ );
not g609 ( new_n824_, new_n823_ );
not g610 ( new_n825_, keyIn_0_98 );
nand g611 ( new_n826_, new_n814_, new_n825_, new_n808_, new_n816_ );
nand g612 ( new_n827_, new_n821_, new_n820_ );
nand g613 ( new_n828_, new_n827_, keyIn_0_97 );
nand g614 ( new_n829_, new_n824_, new_n807_, new_n826_, new_n828_ );
nand g615 ( new_n830_, new_n828_, new_n826_, new_n818_, new_n822_ );
nand g616 ( new_n831_, new_n830_, keyIn_0_104 );
nand g617 ( new_n832_, new_n829_, new_n831_, new_n806_, N219 );
nand g618 ( new_n833_, N96, N210 );
nand g619 ( new_n834_, new_n829_, new_n831_, N219 );
nand g620 ( new_n835_, new_n834_, keyIn_0_110 );
nand g621 ( new_n836_, new_n835_, keyIn_0_116, new_n832_, new_n833_ );
not g622 ( new_n837_, keyIn_0_116 );
nand g623 ( new_n838_, new_n835_, new_n832_, new_n833_ );
nand g624 ( new_n839_, new_n838_, new_n837_ );
nand g625 ( new_n840_, new_n808_, N228 );
not g626 ( new_n841_, new_n840_ );
nand g627 ( new_n842_, new_n641_, N237 );
nand g628 ( new_n843_, new_n393_, N171 );
nand g629 ( new_n844_, new_n594_, N246 );
nand g630 ( new_n845_, new_n842_, new_n843_, new_n844_ );
nor g631 ( new_n846_, new_n841_, new_n845_ );
nand g632 ( new_n847_, new_n839_, new_n836_, new_n846_ );
nand g633 ( new_n848_, new_n847_, new_n805_ );
nand g634 ( new_n849_, new_n839_, keyIn_0_120, new_n836_, new_n846_ );
nand g635 ( new_n850_, new_n848_, new_n849_ );
nand g636 ( new_n851_, new_n850_, keyIn_0_124 );
not g637 ( new_n852_, keyIn_0_124 );
nand g638 ( new_n853_, new_n848_, new_n852_, new_n849_ );
nand g639 ( new_n854_, new_n851_, new_n853_ );
nand g640 ( new_n855_, new_n854_, keyIn_0_127 );
not g641 ( new_n856_, keyIn_0_127 );
nand g642 ( new_n857_, new_n851_, new_n856_, new_n853_ );
nand g643 ( N880, new_n855_, new_n857_ );
endmodule