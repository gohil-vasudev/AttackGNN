module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, WX1266, WX1268, WX1270, DFF_163_n1, WX1272,
         WX1274, WX1276, WX1278, WX1280, WX1282, WX1284, DFF_170_n1, WX1286,
         WX1288, WX1290, WX1292, WX1294, WX1296, WX1298, WX1300, WX1302,
         WX1304, WX1306, WX1308, WX1310, WX1312, WX1314, WX1316, WX1318,
         WX1320, WX1322, WX1324, WX1326, DFF_191_n1, WX1778, n8702, n4033,
         n8701, n4032, n8700, n4031, n8699, n4030, n4029, n8696, n4028, n8695,
         n4027, n8694, n4026, n8693, n4025, n8692, n4024, n8691, n4023, n8690,
         n4022, n8689, n4021, n8688, n4020, n8687, n4019, n8686, n4018, n8685,
         n4017, n8684, n4016, n8683, n4015, n8682, n4014, n8681, n4013, n8680,
         n4012, n4011, n8677, n4010, n8676, n4009, n8675, n4008, n8674, n4007,
         n8673, n4006, n8672, n4005, n8671, n4004, WX1839, n8670, n4003,
         WX1937, n8669, WX1939, n8668, WX1941, n8667, WX1943, n8666, WX1945,
         n8665, WX1947, n8664, WX1949, n8663, WX1951, n8662, WX1953, n8661,
         WX1955, WX1957, n8658, WX1959, n8657, WX1961, n8656, WX1963, n8655,
         WX1965, n8654, WX1967, n8653, WX1969, WX1970, WX1971, WX1972, WX1973,
         WX1974, WX1975, WX1976, WX1977, WX1978, WX1979, WX1980, WX1981,
         WX1982, WX1983, WX1984, WX1985, WX1986, WX1987, WX1988, WX1989,
         WX1990, WX1991, WX1993, WX1994, WX1995, WX1996, WX1997, WX1998,
         WX1999, WX2000, WX2001, WX2002, WX2003, WX2004, WX2005, WX2006,
         WX2007, WX2008, WX2009, WX2010, WX2011, WX2012, WX2013, WX2014,
         WX2015, WX2016, WX2017, WX2018, WX2019, WX2020, WX2021, WX2022,
         WX2023, WX2024, WX2025, WX2026, WX2027, WX2029, WX2030, WX2031,
         WX2032, WX2033, WX2034, WX2035, WX2036, WX2037, WX2038, WX2039,
         WX2040, WX2041, WX2042, WX2043, WX2044, WX2045, WX2046, WX2047,
         WX2048, WX2049, WX2050, WX2051, WX2052, WX2053, WX2054, WX2055,
         WX2056, WX2057, WX2058, WX2059, WX2060, WX2061, WX2062, WX2063,
         WX2065, WX2066, WX2067, WX2068, WX2069, WX2070, WX2071, WX2072,
         WX2073, WX2074, WX2075, WX2076, WX2077, WX2078, WX2079, WX2080,
         WX2081, WX2082, WX2083, WX2084, WX2085, WX2086, WX2087, WX2088,
         WX2089, WX2090, WX2091, WX2092, WX2093, WX2094, WX2095, WX2096,
         WX2097, WX2098, WX2099, WX2101, WX2102, WX2103, WX2104, WX2105,
         WX2106, WX2107, WX2108, WX2109, WX2110, WX2111, WX2112, WX2113,
         WX2114, WX2115, WX2116, WX2117, WX2118, WX2119, WX2120, WX2121,
         WX2122, WX2123, WX2124, WX2125, WX2126, WX2127, WX2128, WX2129,
         WX2130, WX2131, WX2132, WX2133, WX2134, WX2135, WX2137, WX2138,
         WX2139, WX2140, WX2141, WX2142, WX2143, WX2144, WX2145, WX2146,
         WX2147, WX2148, WX2149, WX2150, WX2151, WX2152, WX2153, WX2154,
         WX2155, WX2156, WX2157, WX2158, WX2159, WX2160, WX2161, WX2162,
         WX2163, WX2164, WX2165, WX2166, WX2167, WX2168, WX2169, WX2170,
         WX2171, WX2173, WX2174, WX2175, WX2176, WX2177, WX2178, WX2179,
         WX2180, WX2181, WX2182, WX2183, WX2184, WX2185, WX2186, WX2187,
         WX2188, WX2189, WX2190, WX2191, WX2192, WX2557, WX2559, WX2561,
         WX2563, DFF_355_n1, WX2565, WX2567, WX2569, WX2571, WX2573, WX2575,
         DFF_361_n1, WX2577, DFF_362_n1, WX2579, WX2581, WX2583, WX2585,
         WX2587, DFF_367_n1, WX2589, WX2591, WX2593, WX2595, WX2597, WX2599,
         WX2601, WX2603, WX2605, WX2607, WX2609, WX2611, DFF_379_n1, WX2613,
         WX2615, WX2617, WX2619, DFF_383_n1, WX3071, n8644, n4002, n8643,
         n4001, n8642, n4000, n8641, n3999, n8640, n3998, n8639, n3997, n8638,
         n3996, n8637, n3995, n8636, n3994, n8635, n3993, n3992, n8632, n3991,
         n8631, n3990, n8630, n3989, n8629, n3988, n8628, n3987, n8627, n3986,
         n8626, n3985, n8625, n3984, n8624, n3983, n8623, n3982, n8622, n3981,
         n8621, n3980, n8620, n3979, n8619, n3978, n8618, n3977, n8617, n3976,
         n8616, n3975, n3974, n8613, n3973, WX3132, n8612, n3972, WX3230,
         n8611, WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238, n8607,
         WX3240, n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603, WX3248,
         n8602, WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256, n8598,
         WX3258, n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266, WX3267,
         WX3268, WX3269, WX3270, WX3271, WX3272, WX3273, WX3274, WX3275,
         WX3276, WX3277, WX3278, WX3279, WX3280, WX3281, WX3282, WX3283,
         WX3284, WX3285, WX3286, WX3287, WX3288, WX3289, WX3290, WX3291,
         WX3292, WX3293, WX3294, WX3295, WX3296, WX3298, WX3299, WX3300,
         WX3301, WX3302, WX3303, WX3304, WX3305, WX3306, WX3307, WX3308,
         WX3309, WX3310, WX3311, WX3312, WX3313, WX3314, WX3315, WX3316,
         WX3317, WX3318, WX3319, WX3320, WX3321, WX3322, WX3323, WX3324,
         WX3325, WX3326, WX3327, WX3328, WX3329, WX3330, WX3331, WX3332,
         WX3334, WX3335, WX3336, WX3337, WX3338, WX3339, WX3340, WX3341,
         WX3342, WX3343, WX3344, WX3345, WX3346, WX3347, WX3348, WX3349,
         WX3350, WX3351, WX3352, WX3353, WX3354, WX3355, WX3356, WX3357,
         WX3358, WX3359, WX3360, WX3361, WX3362, WX3363, WX3364, WX3365,
         WX3366, WX3367, WX3368, WX3370, WX3371, WX3372, WX3373, WX3374,
         WX3375, WX3376, WX3377, WX3378, WX3379, WX3380, WX3381, WX3382,
         WX3383, WX3384, WX3385, WX3386, WX3387, WX3388, WX3389, WX3390,
         WX3391, WX3392, WX3393, WX3394, WX3395, WX3396, WX3397, WX3398,
         WX3399, WX3400, WX3401, WX3402, WX3403, WX3404, WX3406, WX3407,
         WX3408, WX3409, WX3410, WX3411, WX3412, WX3413, WX3414, WX3415,
         WX3416, WX3417, WX3418, WX3419, WX3420, WX3421, WX3422, WX3423,
         WX3424, WX3425, WX3426, WX3427, WX3428, WX3429, WX3430, WX3431,
         WX3432, WX3433, WX3434, WX3435, WX3436, WX3437, WX3438, WX3440,
         WX3441, WX3442, WX3443, WX3444, WX3445, WX3446, WX3447, WX3448,
         WX3449, WX3450, WX3451, WX3452, WX3453, WX3454, WX3455, WX3456,
         WX3457, WX3458, WX3459, WX3460, WX3461, WX3462, WX3463, WX3464,
         WX3465, WX3466, WX3467, WX3468, WX3469, WX3470, WX3471, WX3472,
         WX3474, WX3475, WX3476, WX3477, WX3478, WX3479, WX3480, WX3481,
         WX3482, WX3483, WX3484, WX3485, WX3850, WX3852, WX3854, WX3856,
         DFF_547_n1, WX3858, WX3860, DFF_549_n1, WX3862, WX3864, WX3866,
         WX3868, WX3870, WX3872, WX3874, WX3876, WX3878, WX3880, DFF_559_n1,
         WX3882, WX3884, WX3886, WX3888, WX3890, WX3892, WX3894, DFF_566_n1,
         WX3896, WX3898, WX3900, WX3902, WX3904, WX3906, WX3908, WX3910,
         WX3912, DFF_575_n1, WX4364, n8586, n3971, n8585, n3970, n8584, n3969,
         n8583, n3968, n8582, n3967, n8581, n3966, n8580, n3965, n8579, n3964,
         n8578, n3963, n8577, n3962, n8576, n3961, n3960, n8573, n3959, n8572,
         n3958, n8571, n3957, n8570, n3956, n8569, n3955, n8568, n3954, n8567,
         n3953, n8566, n3952, n8565, n3951, n8564, n3950, n8563, n3949, n8562,
         n3948, n8561, n3947, n8560, n3946, n8559, n3945, n8558, n3944, n3943,
         n8555, n3942, WX4425, n8554, n3941, WX4523, n8553, WX4525, n8552,
         WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533, n8548, WX4535,
         n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544, WX4543, n8543,
         WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551, WX4553, n8537,
         WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561, WX4562,
         WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569, WX4570,
         WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577, WX4578,
         WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585, WX4587,
         WX4588, WX4589, WX4590, WX4591, WX4592, WX4593, WX4594, WX4595,
         WX4596, WX4597, WX4598, WX4599, WX4600, WX4601, WX4602, WX4603,
         WX4604, WX4605, WX4606, WX4607, WX4608, WX4609, WX4610, WX4611,
         WX4612, WX4613, WX4614, WX4615, WX4616, WX4617, WX4618, WX4619,
         WX4621, WX4622, WX4623, WX4624, WX4625, WX4626, WX4627, WX4628,
         WX4629, WX4630, WX4631, WX4632, WX4633, WX4634, WX4635, WX4636,
         WX4637, WX4638, WX4639, WX4640, WX4641, WX4642, WX4643, WX4644,
         WX4645, WX4646, WX4647, WX4648, WX4649, WX4650, WX4651, WX4652,
         WX4653, WX4655, WX4656, WX4657, WX4658, WX4659, WX4660, WX4661,
         WX4662, WX4663, WX4664, WX4665, WX4666, WX4667, WX4668, WX4669,
         WX4670, WX4671, WX4672, WX4673, WX4674, WX4675, WX4676, WX4677,
         WX4678, WX4679, WX4680, WX4681, WX4682, WX4683, WX4684, WX4685,
         WX4686, WX4687, WX4689, WX4690, WX4691, WX4692, WX4693, WX4694,
         WX4695, WX4696, WX4697, WX4698, WX4699, WX4700, WX4701, WX4702,
         WX4703, WX4704, WX4705, WX4706, WX4707, WX4708, WX4709, WX4710,
         WX4711, WX4712, WX4713, WX4714, WX4715, WX4716, WX4717, WX4718,
         WX4719, WX4720, WX4721, WX4723, WX4724, WX4725, WX4726, WX4727,
         WX4728, WX4729, WX4730, WX4731, WX4732, WX4733, WX4734, WX4735,
         WX4736, WX4737, WX4738, WX4739, WX4740, WX4741, WX4742, WX4743,
         WX4744, WX4745, WX4746, WX4747, WX4748, WX4749, WX4750, WX4751,
         WX4752, WX4753, WX4754, WX4755, WX4757, WX4758, WX4759, WX4760,
         WX4761, WX4762, WX4763, WX4764, WX4765, WX4766, WX4767, WX4768,
         WX4769, WX4770, WX4771, WX4772, WX4773, WX4774, WX4775, WX4776,
         WX4777, WX4778, WX5143, WX5145, WX5147, WX5149, DFF_739_n1, WX5151,
         WX5153, WX5155, WX5157, WX5159, WX5161, WX5163, WX5165, WX5167,
         WX5169, WX5171, WX5173, DFF_751_n1, WX5175, WX5177, WX5179, WX5181,
         WX5183, WX5185, WX5187, WX5189, WX5191, WX5193, WX5195, WX5197,
         DFF_763_n1, WX5199, WX5201, WX5203, WX5205, DFF_767_n1, WX5657, n8528,
         n3940, n8527, n3939, n8526, n3938, n8525, n3937, n8524, n3936, n8523,
         n3935, n3934, n8520, n3933, n8519, n3932, n8518, n3931, n8517, n3930,
         n8516, n3929, n8515, n3928, n8514, n3927, n8513, n3926, n8512, n3925,
         n8511, n3924, n8510, n3923, n8509, n3922, n8508, n3921, n8507, n3920,
         n8506, n3919, n8505, n3918, n3917, n8502, n3916, n8501, n3915, n8500,
         n3914, n8499, n3913, n8498, n3912, n8497, n3911, WX5718, n8496, n3910,
         WX5816, n8495, WX5818, n8494, WX5820, n8493, WX5822, n8492, WX5824,
         n8491, WX5826, n8490, WX5828, n8489, WX5830, n8488, WX5832, n8487,
         WX5834, WX5836, n8484, WX5838, n8483, WX5840, n8482, WX5842, n8481,
         WX5844, n8480, WX5846, n8479, WX5848, WX5849, WX5850, WX5851, WX5852,
         WX5853, WX5854, WX5855, WX5856, WX5857, WX5858, WX5859, WX5860,
         WX5861, WX5862, WX5863, WX5864, WX5865, WX5866, WX5867, WX5868,
         WX5870, WX5871, WX5872, WX5873, WX5874, WX5875, WX5876, WX5877,
         WX5878, WX5879, WX5880, WX5881, WX5882, WX5883, WX5884, WX5885,
         WX5886, WX5887, WX5888, WX5889, WX5890, WX5891, WX5892, WX5893,
         WX5894, WX5895, WX5896, WX5897, WX5898, WX5899, WX5900, WX5901,
         WX5902, WX5904, WX5905, WX5906, WX5907, WX5908, WX5909, WX5910,
         WX5911, WX5912, WX5913, WX5914, WX5915, WX5916, WX5917, WX5918,
         WX5919, WX5920, WX5921, WX5922, WX5923, WX5924, WX5925, WX5926,
         WX5927, WX5928, WX5929, WX5930, WX5931, WX5932, WX5933, WX5934,
         WX5935, WX5936, WX5938, WX5939, WX5940, WX5941, WX5942, WX5943,
         WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950, WX5951,
         WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958, WX5959,
         WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966, WX5967,
         WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975, WX5976,
         WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983, WX5984,
         WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991, WX5992,
         WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999, WX6000,
         WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008, WX6009,
         WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016, WX6017,
         WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024, WX6025,
         WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032, WX6033,
         WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041, WX6042,
         WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049, WX6050,
         WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057, WX6058,
         WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065, WX6066,
         WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438, WX6440,
         WX6442, DFF_931_n1, WX6444, WX6446, WX6448, WX6450, WX6452, WX6454,
         WX6456, DFF_938_n1, WX6458, WX6460, WX6462, WX6464, WX6466, WX6468,
         WX6470, WX6472, WX6474, WX6476, WX6478, WX6480, WX6482, WX6484,
         WX6486, WX6488, WX6490, WX6492, WX6494, WX6496, WX6498, DFF_959_n1,
         WX6950, n8470, n3909, n3908, n8467, n3907, n8466, n3906, n8465, n3905,
         n8464, n3904, n8463, n3903, n8462, n3902, n8461, n3901, n8460, n3900,
         n8459, n3899, n8458, n3898, n8457, n3897, n8456, n3896, n8455, n3895,
         n8454, n3894, n8453, n3893, n8452, n3892, n3891, n8449, n3890, n8448,
         n3889, n8447, n3888, n8446, n3887, n8445, n3886, WX6999, n8444, n3885,
         n8443, n8442, n3883, n8441, n3882, n8440, n3881, n8439, n3880, WX7011,
         n8438, n3879, WX7109, n8437, WX7111, n8436, WX7113, n8435, WX7115,
         n8434, WX7117, WX7119, n8431, WX7121, n8430, WX7123, n8429, WX7125,
         n8428, WX7127, n8427, WX7129, n8426, WX7131, n8425, WX7133, n8424,
         WX7135, n8423, WX7137, n8422, WX7139, n8421, WX7141, WX7142, WX7143,
         WX7144, WX7145, WX7146, WX7147, WX7148, WX7149, WX7150, WX7151,
         WX7153, WX7154, WX7155, WX7156, WX7157, WX7158, WX7159, WX7160,
         WX7161, WX7162, WX7163, WX7164, WX7165, WX7166, WX7167, WX7168,
         WX7169, WX7170, WX7171, WX7172, WX7173, WX7174, WX7175, WX7176,
         WX7177, WX7178, WX7179, WX7180, WX7181, WX7182, WX7183, WX7184,
         WX7185, WX7187, WX7188, WX7189, WX7190, WX7191, WX7192, WX7193,
         WX7194, WX7195, WX7196, WX7197, WX7198, WX7199, WX7200, WX7201,
         WX7202, WX7203, WX7204, WX7205, WX7206, WX7207, WX7208, WX7209,
         WX7210, WX7211, WX7212, WX7213, WX7214, WX7215, WX7216, WX7217,
         WX7218, WX7219, WX7221, WX7222, WX7223, WX7224, WX7225, WX7226,
         WX7227, WX7228, WX7229, WX7230, WX7231, WX7232, WX7233, WX7234,
         WX7235, WX7236, WX7237, WX7238, WX7239, WX7240, WX7241, WX7242,
         WX7243, WX7244, WX7245, WX7246, WX7247, WX7248, WX7249, WX7250,
         WX7251, WX7252, WX7253, WX7255, WX7256, WX7257, WX7258, WX7259,
         WX7260, WX7261, WX7262, WX7263, WX7264, WX7265, WX7266, WX7267,
         WX7268, WX7269, WX7270, WX7271, WX7272, WX7273, WX7274, WX7275,
         WX7276, WX7277, WX7278, WX7279, WX7280, WX7281, WX7282, WX7283,
         WX7284, WX7285, WX7286, WX7287, WX7289, WX7290, WX7291, WX7292,
         WX7293, WX7294, WX7295, WX7296, WX7297, WX7298, WX7299, WX7300,
         WX7301, WX7302, WX7303, WX7304, WX7305, WX7306, WX7307, WX7308,
         WX7309, WX7310, WX7311, WX7312, WX7313, WX7314, WX7315, WX7316,
         WX7317, WX7318, WX7319, WX7320, WX7321, WX7323, WX7324, WX7325,
         WX7326, WX7327, WX7328, WX7329, WX7330, WX7331, WX7332, WX7333,
         WX7334, WX7335, WX7336, WX7337, WX7338, WX7339, WX7340, WX7341,
         WX7342, WX7343, WX7344, WX7345, WX7346, WX7347, WX7348, WX7349,
         WX7350, WX7351, WX7352, WX7353, WX7354, WX7355, WX7357, WX7358,
         WX7359, WX7360, WX7361, WX7362, WX7363, WX7364, WX7729, WX7731,
         WX7733, WX7735, WX7737, WX7739, WX7741, WX7743, WX7745, WX7747,
         WX7749, DFF_1130_n1, WX7751, WX7753, WX7755, WX7757, WX7759,
         DFF_1135_n1, WX7761, WX7763, WX7765, WX7767, WX7769, DFF_1140_n1,
         WX7771, WX7773, WX7775, WX7777, WX7779, WX7781, WX7783, WX7785,
         WX7787, WX7789, WX7791, DFF_1151_n1, WX8243, n8411, n3878, n8410,
         n3877, n8409, n3876, n8408, n3875, n8407, n3874, n8406, n3873, n8405,
         n3872, n8404, n3871, n8403, n3870, n8402, n3869, n8401, n3868, WX8266,
         n8400, n3867, n8399, n3865, n8396, n3864, n8395, n3863, n8394, n3862,
         n8393, n3861, n8392, n3860, n8391, n3859, n8390, n3858, n8389, n3857,
         n8388, n3856, n8387, n3855, n8386, n3854, n8385, n3853, n8384, n3852,
         n8383, n3851, n8382, n3850, n8381, n3849, WX8304, n3848, WX8402,
         n8378, WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410, n8374,
         WX8412, n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370, WX8420,
         n8369, WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428, n8365,
         WX8430, n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438, WX8439,
         WX8440, WX8441, WX8442, WX8443, WX8444, WX8445, WX8446, WX8447,
         WX8448, WX8449, WX8450, WX8451, WX8452, WX8453, WX8454, WX8455,
         WX8456, WX8457, WX8458, WX8459, WX8460, WX8461, WX8462, WX8463,
         WX8464, WX8465, WX8466, WX8467, WX8468, WX8470, WX8471, WX8472,
         WX8473, WX8474, WX8475, WX8476, WX8477, WX8478, WX8479, WX8480,
         WX8481, WX8482, WX8483, WX8484, WX8485, WX8486, WX8487, WX8488,
         WX8489, WX8490, WX8491, WX8492, WX8493, WX8494, WX8495, WX8496,
         WX8497, WX8498, WX8499, WX8500, WX8501, WX8502, WX8504, WX8505,
         WX8506, WX8507, WX8508, WX8509, WX8510, WX8511, WX8512, WX8513,
         WX8514, WX8515, WX8516, WX8517, WX8518, WX8519, WX8520, WX8521,
         WX8522, WX8523, WX8524, WX8525, WX8526, WX8527, WX8528, WX8529,
         WX8530, WX8531, WX8532, WX8533, WX8534, WX8535, WX8536, WX8538,
         WX8539, WX8540, WX8541, WX8542, WX8543, WX8544, WX8545, WX8546,
         WX8547, WX8548, WX8549, WX8550, WX8551, WX8552, WX8553, WX8554,
         WX8555, WX8556, WX8557, WX8558, WX8559, WX8560, WX8561, WX8562,
         WX8563, WX8564, WX8565, WX8566, WX8567, WX8568, WX8569, WX8570,
         WX8572, WX8573, WX8574, WX8575, WX8576, WX8577, WX8578, WX8579,
         WX8580, WX8581, WX8582, WX8583, WX8584, WX8585, WX8586, WX8587,
         WX8588, WX8589, WX8590, WX8591, WX8592, WX8593, WX8594, WX8595,
         WX8596, WX8597, WX8598, WX8599, WX8600, WX8601, WX8602, WX8603,
         WX8604, WX8606, WX8607, WX8608, WX8609, WX8610, WX8611, WX8612,
         WX8613, WX8614, WX8615, WX8616, WX8617, WX8618, WX8619, WX8620,
         WX8621, WX8622, WX8623, WX8624, WX8625, WX8626, WX8627, WX8628,
         WX8629, WX8630, WX8631, WX8632, WX8633, WX8634, WX8635, WX8636,
         WX8637, WX8638, WX8640, WX8641, WX8642, WX8643, WX8644, WX8645,
         WX8646, WX8647, WX8648, WX8649, WX8650, WX8651, WX8652, WX8653,
         WX8654, WX8655, WX8656, WX8657, WX9022, WX9024, WX9026, WX9028,
         DFF_1315_n1, WX9030, WX9032, WX9034, WX9036, WX9038, DFF_1320_n1,
         WX9040, WX9042, DFF_1322_n1, WX9044, WX9046, WX9048, WX9050, WX9052,
         DFF_1327_n1, WX9054, WX9056, WX9058, WX9060, WX9062, WX9064, WX9066,
         WX9068, WX9070, WX9072, DFF_1337_n1, WX9074, WX9076, WX9078, WX9080,
         WX9082, WX9084, DFF_1343_n1, WX9536, n8353, n3847, n8352, n3846,
         n8351, n3845, n8350, n3844, n8349, n3843, n8348, n3842, n8347, n3841,
         n8346, n3840, n3839, n8343, n3838, n8342, n3837, n8341, n3836, n8340,
         n3835, n8339, n3834, n8338, n3833, n8337, n3832, n8336, n3831, n8335,
         n3830, n8334, n3829, n8333, n3828, n8332, n3827, n8331, n3826, n8330,
         n3825, n8329, n3824, n8328, n3823, n3822, n8325, n3821, n8324, n3820,
         n8323, n3819, n8322, n3818, WX9597, n8321, n3817, WX9695, n8320,
         WX9697, n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705,
         n8315, WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311,
         WX9715, n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305,
         WX9725, n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733,
         WX9734, WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741,
         WX9742, WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749,
         WX9750, WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758,
         WX9759, WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766,
         WX9767, WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774,
         WX9775, WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782,
         WX9783, WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791,
         WX9792, WX9793, WX9794, WX9795, WX9796, WX9797, WX9798, WX9799,
         WX9800, WX9801, WX9802, WX9803, WX9804, WX9805, WX9806, WX9807,
         WX9808, WX9809, WX9810, WX9811, WX9812, WX9813, WX9814, WX9815,
         WX9816, WX9817, WX9818, WX9819, WX9821, WX9822, WX9823, WX9824,
         WX9825, WX9826, WX9827, WX9828, WX9829, WX9830, WX9831, WX9832,
         WX9833, WX9834, WX9835, WX9836, WX9837, WX9838, WX9839, WX9840,
         WX9841, WX9842, WX9843, WX9844, WX9845, WX9846, WX9847, WX9848,
         WX9849, WX9850, WX9851, WX9852, WX9853, WX9855, WX9856, WX9857,
         WX9858, WX9859, WX9860, WX9861, WX9862, WX9863, WX9864, WX9865,
         WX9866, WX9867, WX9868, WX9869, WX9870, WX9871, WX9872, WX9873,
         WX9874, WX9875, WX9876, WX9877, WX9878, WX9879, WX9880, WX9881,
         WX9882, WX9883, WX9884, WX9885, WX9886, WX9887, WX9889, WX9890,
         WX9891, WX9892, WX9893, WX9894, WX9895, WX9896, WX9897, WX9898,
         WX9899, WX9900, WX9901, WX9902, WX9903, WX9904, WX9905, WX9906,
         WX9907, WX9908, WX9909, WX9910, WX9911, WX9912, WX9913, WX9914,
         WX9915, WX9916, WX9917, WX9918, WX9919, WX9920, WX9921, WX9923,
         WX9924, WX9925, WX9926, WX9927, WX9928, WX9929, WX9930, WX9931,
         WX9932, WX9933, WX9934, WX9935, WX9936, WX9937, WX9938, WX9939,
         WX9940, WX9941, WX9942, WX9943, WX9944, WX9945, WX9946, WX9947,
         WX9948, WX9949, WX9950, WX10315, WX10317, WX10319, WX10321,
         DFF_1507_n1, WX10323, WX10325, WX10327, WX10329, WX10331, WX10333,
         WX10335, DFF_1514_n1, WX10337, WX10339, WX10341, DFF_1517_n1, WX10343,
         WX10345, DFF_1519_n1, WX10347, WX10349, WX10351, WX10353, WX10355,
         WX10357, WX10359, WX10361, WX10363, WX10365, WX10367, WX10369,
         WX10371, WX10373, WX10375, DFF_1534_n1, WX10377, DFF_1535_n1, WX10829,
         n8295, n3816, n8294, n3815, n8293, n3814, n3813, n8290, n3812, n8289,
         n3811, n8288, n3810, n8287, n3809, n8286, n3808, n8285, n3807, n8284,
         n3806, n8283, n3805, n8282, n3804, n8281, n3803, n8280, n3802, n8279,
         n3801, n8278, n3800, n8277, n3799, n8276, n3798, n8275, n3797, n3796,
         n8272, n3795, n8271, n3794, n8270, n3793, n8269, n3792, n8268, n3791,
         n8267, n3790, n8266, n3789, n8265, n3788, n8264, n3787, WX10890,
         n8263, n3786, WX10988, n8262, WX10990, n8261, WX10992, n8260, WX10994,
         n8259, WX10996, n8258, WX10998, n8257, WX11000, WX11002, n8254,
         WX11004, n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250,
         WX11012, n8249, WX11014, n8248, WX11016, n8247, WX11018, n8246,
         WX11020, WX11021, WX11022, WX11023, WX11024, WX11025, WX11026,
         WX11027, WX11028, WX11029, WX11030, WX11031, WX11032, WX11033,
         WX11034, WX11036, WX11037, WX11038, WX11039, WX11040, WX11041,
         WX11042, WX11043, WX11044, WX11045, WX11046, WX11047, WX11048,
         WX11049, WX11050, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, WX11086, WX11087, WX11088, WX11089, WX11090, WX11091,
         WX11092, WX11093, WX11094, WX11095, WX11096, WX11097, WX11098,
         WX11099, WX11100, WX11101, WX11102, WX11104, WX11105, WX11106,
         WX11107, WX11108, WX11109, WX11110, WX11111, WX11112, WX11113,
         WX11114, WX11115, WX11116, WX11117, WX11118, WX11119, WX11120,
         WX11121, WX11122, WX11123, WX11124, WX11125, WX11126, WX11127,
         WX11128, WX11129, WX11130, WX11131, WX11132, WX11133, WX11134,
         WX11135, WX11136, WX11138, WX11139, WX11140, WX11141, WX11142,
         WX11143, WX11144, WX11145, WX11146, WX11147, WX11148, WX11149,
         WX11150, WX11151, WX11152, WX11153, WX11154, WX11155, WX11156,
         WX11157, WX11158, WX11159, WX11160, WX11161, WX11162, WX11163,
         WX11164, WX11165, WX11166, WX11167, WX11168, WX11169, WX11170,
         WX11172, WX11173, WX11174, WX11175, WX11176, WX11177, WX11178,
         WX11179, WX11180, WX11181, WX11182, WX11183, WX11184, WX11185,
         WX11186, WX11187, WX11188, WX11189, WX11190, WX11191, WX11192,
         WX11193, WX11194, WX11195, WX11196, WX11197, WX11198, WX11199,
         WX11200, WX11201, WX11202, WX11203, WX11204, WX11206, WX11207,
         WX11208, WX11209, WX11210, WX11211, WX11212, WX11213, WX11214,
         WX11215, WX11216, WX11217, WX11218, WX11219, WX11220, WX11221,
         WX11222, WX11223, WX11224, WX11225, WX11226, WX11227, WX11228,
         WX11229, WX11230, WX11231, WX11232, WX11233, WX11234, WX11235,
         WX11236, WX11237, WX11238, WX11240, WX11241, WX11242, WX11243,
         WX11608, WX11610, DFF_1697_n1, WX11612, WX11614, WX11616, WX11618,
         WX11620, WX11622, WX11624, WX11626, WX11628, WX11630, WX11632,
         WX11634, WX11636, WX11638, WX11640, WX11642, WX11644, DFF_1714_n1,
         WX11646, WX11648, WX11650, WX11652, WX11654, WX11656, WX11658,
         WX11660, WX11662, WX11664, WX11666, WX11668, WX11670, n2245, n2153,
         n3278, n2152, n2148, Tj_Trigger, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4,
         Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n308, n309, n310, n311, n312, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n530,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4280, n4282, n4284, n4286, n4289, n4292,
         n4295, n4297, n4299, n4301, n4303, n4305, n4307, n4309, n4312, n4315,
         n4317, n4319, n4321, n4323, n4325, n4327, n4329, n4331, n4333, n4335,
         n4337, n4339, n4341, n4343, n4345, n4347, n4349, n4351, n4353, n4355,
         n4357, n4359, n4362, n4365, n4368, n4370, n4372, n4374, n4376, n4378,
         n4381, n4384, n4387, n4389, n4391, n4393, n4395, n4397, n4400, n4403,
         n4406, n4408, n4410, n4412, n4414, n4416, n4418, n4420, n4422, n4424,
         n4427, n4429, n4431, n4433, n4435, n4437, n4439, n4441, n4443, n4445,
         n4447, n4449, n4452, n4455, n4457, n4459, n4461, n4463, n4465, n4467,
         n4469, n4472, n4474, n4476, n4479, n4481, n4483, n4486, n4488, n4490,
         n4493, n4495, n4497, n4499, n4501, n4503, n4505, n4507, n4509, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8255, n8256,
         n8273, n8274, n8291, n8292, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8308, n8309, n8326, n8327, n8344, n8345, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8379, n8380, n8397,
         n8398, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8432, n8433, n8450, n8451, n8468, n8469, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8485, n8486, n8503, n8504, n8521, n8522,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8538, n8539,
         n8556, n8557, n8574, n8575, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8614, n8615, n8633, n8634, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8659, n8660, n8678, n8679,
         n8697, n8698, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1,
         U5718_n1, U5719_n1, U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1,
         U5725_n1, U5726_n1, U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1,
         U5732_n1, U5733_n1, U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1,
         U5739_n1, U5740_n1, U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1,
         U5746_n1, U5747_n1, U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1,
         U5753_n1, U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1,
         U5760_n1, U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1,
         U5767_n1, U5768_n1, U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1,
         U5774_n1, U5775_n1, U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1,
         U5781_n1, U5782_n1, U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1,
         U5788_n1, U5789_n1, U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1,
         U5795_n1, U5796_n1, U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1,
         U5802_n1, U5803_n1, U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1,
         U5809_n1, U5810_n1, U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1,
         U5816_n1, U5817_n1, U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1,
         U5823_n1, U5824_n1, U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1,
         U5830_n1, U5831_n1, U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1,
         U5837_n1, U5838_n1, U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1,
         U5844_n1, U5845_n1, U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1,
         U5851_n1, U5852_n1, U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1,
         U5858_n1, U5859_n1, U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1,
         U5865_n1, U5866_n1, U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1,
         U5872_n1, U5873_n1, U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1,
         U5879_n1, U5880_n1, U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1,
         U5886_n1, U5887_n1, U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1,
         U5893_n1, U5894_n1, U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1,
         U5900_n1, U5901_n1, U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1,
         U5907_n1, U5908_n1, U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1,
         U5914_n1, U5915_n1, U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1,
         U5921_n1, U5922_n1, U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1,
         U5928_n1, U5929_n1, U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1,
         U5935_n1, U5936_n1, U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1,
         U5942_n1, U5943_n1, U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1,
         U5949_n1, U5950_n1, U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1,
         U5956_n1, U5957_n1, U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1,
         U5963_n1, U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1,
         U5970_n1, U5971_n1, U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1,
         U5977_n1, U5978_n1, U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1,
         U5984_n1, U5985_n1, U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1,
         U5991_n1, U5992_n1, U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1,
         U5998_n1, U5999_n1, U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1,
         U6005_n1, U6006_n1, U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1,
         U6012_n1, U6013_n1, U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1,
         U6019_n1, U6020_n1, U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1,
         U6026_n1, U6027_n1, U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1,
         U6033_n1, U6034_n1, U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1,
         U6040_n1, U6041_n1, U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1,
         U6047_n1, U6048_n1, U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1,
         U6054_n1, U6055_n1, U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1,
         U6061_n1, U6062_n1, U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1,
         U6068_n1, U6069_n1, U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1,
         U6075_n1, U6076_n1, U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1,
         U6082_n1, U6083_n1, U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1,
         U6089_n1, U6090_n1, U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1,
         U6096_n1, U6097_n1, U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1,
         U6103_n1, U6104_n1, U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1,
         U6110_n1, U6111_n1, U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1,
         U6117_n1, U6118_n1, U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1,
         U6124_n1, U6125_n1, U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1,
         U6131_n1, U6132_n1, U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1,
         U6138_n1, U6139_n1, U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1,
         U6145_n1, U6146_n1, U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1,
         U6152_n1, U6153_n1, U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1,
         U6159_n1, U6160_n1, U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1,
         U6166_n1, U6167_n1, U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1,
         U6173_n1, U6174_n1, U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1,
         U6180_n1, U6181_n1, U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1,
         U6187_n1, U6188_n1, U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1,
         U6194_n1, U6195_n1, U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1,
         U6201_n1, U6202_n1, U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1,
         U6208_n1, U6209_n1, U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1,
         U6215_n1, U6216_n1, U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1,
         U6222_n1, U6223_n1, U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1,
         U6229_n1, U6230_n1, U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1,
         U6236_n1, U6237_n1, U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1,
         U6243_n1, U6244_n1, U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1,
         U6250_n1, U6251_n1, U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1,
         U6257_n1, U6258_n1, U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1,
         U6264_n1, U6265_n1, U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1,
         U6271_n1, U6272_n1, U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1,
         U6278_n1, U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1,
         U6285_n1, U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1,
         U6292_n1, U6293_n1, U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1,
         U6299_n1, U6300_n1, U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1,
         U6306_n1, U6307_n1, U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1,
         U6313_n1, U6314_n1, U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1,
         U6320_n1, U6321_n1, U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1,
         U6327_n1, U6328_n1, U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1,
         U6334_n1, U6335_n1, U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1,
         U6341_n1, U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1,
         U6348_n1, U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1,
         U6355_n1, U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1,
         U6362_n1, U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1,
         U6369_n1, U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1,
         U6376_n1, U6377_n1, U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1,
         U6383_n1, U6384_n1, U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1,
         U6390_n1, U6391_n1, U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1,
         U6397_n1, U6398_n1, U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1,
         U6404_n1, U6405_n1, U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1,
         U6411_n1, U6412_n1, U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1,
         U6418_n1, U6419_n1, U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1,
         U6425_n1, U6426_n1, U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1,
         U6432_n1, U6433_n1, U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1,
         U6439_n1, U6440_n1, U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1,
         U6446_n1, U6447_n1, U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1,
         U6453_n1, U6454_n1, U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1,
         U6460_n1, U6461_n1, U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1,
         U6467_n1, U6468_n1, U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1,
         U6474_n1, U6475_n1, U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1,
         U6481_n1, U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n5232), .CLK(n5542), .Q(
        WX485), .QN(n4827) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n5227), .CLK(n5544), .Q(
        WX487) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n5227), .CLK(n5544), .Q(
        WX489) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n5228), .CLK(n5544), .Q(
        WX491) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n5228), .CLK(n5544), .Q(
        WX493) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n5228), .CLK(n5544), .Q(
        WX495) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n5228), .CLK(n5544), .Q(
        WX497) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n5228), .CLK(n5544), .Q(
        WX499) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n5228), .CLK(n5544), .Q(
        WX501) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n5229), .CLK(n5543), .Q(
        WX503) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n5229), .CLK(n5543), .Q(
        WX505) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n5229), .CLK(n5543), .Q(
        WX507) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n5229), .CLK(n5543), .Q(
        WX509) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n5229), .CLK(n5543), .Q(
        WX511) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n5229), .CLK(n5543), .Q(
        WX513) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n5230), .CLK(n5543), .Q(
        WX515) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n5230), .CLK(n5543), .Q(
        WX517) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n5230), .CLK(n5543), .Q(
        test_so1) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n5230), .CLK(n5543), .Q(
        WX521) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n5230), .CLK(n5543), .Q(
        WX523) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n5230), .CLK(n5543), .Q(
        WX525) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n5231), .CLK(n5542), .Q(
        WX527) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n5231), .CLK(n5542), .Q(
        WX529) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n5231), .CLK(n5542), .Q(
        WX531) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n5231), .CLK(n5542), .Q(
        WX533) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n5231), .CLK(n5542), .Q(
        WX535) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n5231), .CLK(n5542), .Q(
        WX537) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n5232), .CLK(n5542), .Q(
        WX539) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n5232), .CLK(n5542), .Q(
        WX541) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n5232), .CLK(n5542), .Q(
        WX543) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n5232), .CLK(n5542), .Q(
        WX545) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n5232), .CLK(n5542), .Q(
        WX547) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n5227), .CLK(n5544), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n5227), .CLK(n5544), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n5227), .CLK(n5544), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n5227), .CLK(n5544), .Q(
        test_so2) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n5226), .CLK(n5545), .Q(
        WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n5226), .CLK(n5545), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n5226), .CLK(n5545), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n5225), .CLK(n5545), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n5225), .CLK(n5545), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n5225), .CLK(n5545), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n5224), .CLK(n5546), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n5224), .CLK(n5546), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n5224), .CLK(n5546), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n5223), .CLK(n5546), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n5223), .CLK(n5546), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n5222), .CLK(n5547), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n5222), .CLK(n5547), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n5221), .CLK(n5547), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n5220), .CLK(n5548), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n5220), .CLK(n5548), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n5219), .CLK(n5548), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n5218), .CLK(n5549), .Q(
        test_so3) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n4945), .CLK(n5685), .Q(
        WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n5217), .CLK(n5549), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n5216), .CLK(n5550), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n5216), .CLK(n5550), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n5215), .CLK(n5550), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n5214), .CLK(n5551), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n5214), .CLK(n5551), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n5213), .CLK(n5551), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n5212), .CLK(n5552), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n5212), .CLK(n5552), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n5211), .CLK(n5552), .Q(
        WX709) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n5211), .CLK(n5552), .Q(
        WX711), .QN(n4754) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n5210), .CLK(n5553), .Q(
        WX713), .QN(n9771) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n5226), .CLK(n5545), .Q(
        WX715), .QN(n4763) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n5226), .CLK(n5545), .Q(
        WX717), .QN(n9772) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n5226), .CLK(n5545), .Q(
        WX719), .QN(n9773) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n5225), .CLK(n5545), .Q(
        WX721), .QN(n9774) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n5225), .CLK(n5545), .Q(
        test_so4) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n5225), .CLK(n5545), .Q(
        WX725), .QN(n9775) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n5224), .CLK(n5546), .Q(
        WX727), .QN(n4780) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n5224), .CLK(n5546), .Q(
        WX729), .QN(n4784) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n5224), .CLK(n5546), .Q(
        WX731) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n5223), .CLK(n5546), .Q(
        WX733), .QN(n9776) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n5223), .CLK(n5546), .Q(
        WX735), .QN(n9777) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n5222), .CLK(n5547), .Q(
        WX737), .QN(n9778) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n5222), .CLK(n5547), .Q(
        WX739) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n5221), .CLK(n5547), .Q(
        WX741), .QN(n4782) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n5221), .CLK(n5547), .Q(
        WX743), .QN(n9779) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n5220), .CLK(n5548), .Q(
        WX745), .QN(n9780) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n5219), .CLK(n5548), .Q(
        WX747), .QN(n9781) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n5219), .CLK(n5548), .Q(
        WX749), .QN(n9782) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n5218), .CLK(n5549), .Q(
        WX751), .QN(n4768) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n5218), .CLK(n5549), .Q(
        WX753) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n5217), .CLK(n5549), .Q(
        WX755), .QN(n9766) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n5216), .CLK(n5550), .Q(
        WX757), .QN(n4792) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n5216), .CLK(n5550), .Q(
        test_so5) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n5215), .CLK(n5550), .Q(
        WX761), .QN(n9767) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n5214), .CLK(n5551), .Q(
        WX763), .QN(n9768) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n5214), .CLK(n5551), .Q(
        WX765), .QN(n9770) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n5213), .CLK(n5551), .Q(
        WX767) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n5212), .CLK(n5552), .Q(
        WX769), .QN(n9783) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n5212), .CLK(n5552), .Q(
        WX771), .QN(n4795) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n5211), .CLK(n5552), .Q(
        WX773), .QN(n9769) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n5210), .CLK(n5553), .Q(
        WX775) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n5210), .CLK(n5553), .Q(
        WX777) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n5210), .CLK(n5553), .Q(
        WX779) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n5209), .CLK(n5553), .Q(
        WX781) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n5209), .CLK(n5553), .Q(
        WX783) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n5209), .CLK(n5553), .Q(
        WX785) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n5208), .CLK(n5554), .Q(
        WX787) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n5208), .CLK(n5554), .Q(
        WX789) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n5208), .CLK(n5554), .Q(
        WX791) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n5207), .CLK(n5554), .Q(
        WX793) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n5207), .CLK(n5554), .Q(
        test_so6) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n5223), .CLK(n5546), 
        .Q(WX797) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n5223), .CLK(n5546), .Q(
        WX799) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n5222), .CLK(n5547), .Q(
        WX801) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n5222), .CLK(n5547), .Q(
        WX803), .QN(n4776) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n5221), .CLK(n5547), .Q(
        WX805) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n5221), .CLK(n5547), .Q(
        WX807) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n5220), .CLK(n5548), .Q(
        WX809) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n5219), .CLK(n5548), .Q(
        WX811) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n5219), .CLK(n5548), .Q(
        WX813) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n5218), .CLK(n5549), .Q(
        WX815) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n5217), .CLK(n5549), .Q(
        WX817), .QN(n9765) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n5217), .CLK(n5549), .Q(
        WX819) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n5216), .CLK(n5550), .Q(
        WX821) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n5215), .CLK(n5550), .Q(
        WX823) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n5215), .CLK(n5550), .Q(
        WX825) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n5214), .CLK(n5551), .Q(
        WX827) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n5213), .CLK(n5551), .Q(
        WX829) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n5213), .CLK(n5551), .Q(
        test_so7) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n5212), .CLK(n5552), 
        .Q(WX833) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n5211), .CLK(n5552), .Q(
        WX835) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n5211), .CLK(n5552), .Q(
        WX837), .QN(n4789) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n5210), .CLK(n5553), .Q(
        WX839), .QN(n4755) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n5210), .CLK(n5553), .Q(
        WX841), .QN(n4758) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n5209), .CLK(n5553), .Q(
        WX843), .QN(n4762) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n5209), .CLK(n5553), .Q(
        WX845), .QN(n4765) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n5209), .CLK(n5553), .Q(
        WX847), .QN(n4766) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n5208), .CLK(n5554), .Q(
        WX849), .QN(n4770) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n5208), .CLK(n5554), .Q(
        WX851), .QN(n4773) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n5208), .CLK(n5554), .Q(
        WX853), .QN(n4775) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n5207), .CLK(n5554), .Q(
        WX855), .QN(n4781) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n5207), .CLK(n5554), .Q(
        WX857), .QN(n4785) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n5207), .CLK(n5554), .Q(
        WX859), .QN(n4787) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n5207), .CLK(n5554), .Q(
        WX861), .QN(n4757) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n5206), .CLK(n5555), .Q(
        WX863), .QN(n4764) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n5206), .CLK(n5555), .Q(
        WX865), .QN(n4769) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n5206), .CLK(n5555), .Q(
        test_so8) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n5221), .CLK(n5547), 
        .Q(WX869), .QN(n4783) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n5220), .CLK(n5548), .Q(
        WX871), .QN(n4790) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n5220), .CLK(n5548), .Q(
        WX873), .QN(n4759) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n5219), .CLK(n5548), .Q(
        WX875), .QN(n4771) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n5218), .CLK(n5549), .Q(
        WX877), .QN(n4794) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n5218), .CLK(n5549), .Q(
        WX879), .QN(n4767) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n5217), .CLK(n5549), .Q(
        WX881), .QN(n4772) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n5217), .CLK(n5549), .Q(
        WX883), .QN(n4777) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n5216), .CLK(n5550), .Q(
        WX885), .QN(n4793) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n5215), .CLK(n5550), .Q(
        WX887), .QN(n4786) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n5215), .CLK(n5550), .Q(
        WX889), .QN(n4778) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n5214), .CLK(n5551), .Q(
        WX891), .QN(n4779) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n5213), .CLK(n5551), .Q(
        WX893), .QN(n4756) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n5213), .CLK(n5551), .Q(
        WX895), .QN(n4791) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n5212), .CLK(n5552), .Q(
        WX897), .QN(n4760) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n5211), .CLK(n5552), .Q(
        WX899), .QN(n4796) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n4948), .CLK(n5684), .Q(
        CRC_OUT_9_0) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n4948), .CLK(n5684), 
        .Q(test_so9) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n4948), .CLK(n5684), 
        .Q(CRC_OUT_9_2) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_4) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_5) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_6) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_7) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n4947), .CLK(n5684), 
        .Q(CRC_OUT_9_8) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n4946), .CLK(n5685), 
        .Q(CRC_OUT_9_9) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n4946), .CLK(n5685), 
        .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n4946), .CLK(n5685), .Q(CRC_OUT_9_11) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n4946), .CLK(n5685), .Q(CRC_OUT_9_12) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n4946), .CLK(n5685), .Q(CRC_OUT_9_13) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n4946), .CLK(n5685), .Q(CRC_OUT_9_14) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n4945), .CLK(n5685), .Q(CRC_OUT_9_15) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n4945), .CLK(n5685), .Q(CRC_OUT_9_16) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n4945), .CLK(n5685), .Q(CRC_OUT_9_17) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n4945), .CLK(n5685), .Q(CRC_OUT_9_18) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n4945), .CLK(n5685), .Q(test_so10) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n5206), .CLK(n5555), 
        .Q(CRC_OUT_9_20) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n5206), .CLK(n5555), .Q(CRC_OUT_9_21) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n5206), .CLK(n5555), .Q(CRC_OUT_9_22) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_23) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_24) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_25) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_26) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_27) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n5205), .CLK(n5555), .Q(CRC_OUT_9_28) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n5204), .CLK(n5556), .Q(CRC_OUT_9_29) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n5204), .CLK(n5556), .Q(CRC_OUT_9_30) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n5204), .CLK(n5556), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n33), .SI(CRC_OUT_9_31), .SE(n5204), .CLK(n5556), 
        .Q(WX1778), .QN(n4819) );
  SDFFX1 DFF_193_Q_reg ( .D(n34), .SI(WX1778), .SE(n5199), .CLK(n5558), .Q(
        n8702), .QN(n4033) );
  SDFFX1 DFF_194_Q_reg ( .D(n35), .SI(n8702), .SE(n5199), .CLK(n5558), .Q(
        n8701), .QN(n4032) );
  SDFFX1 DFF_195_Q_reg ( .D(n36), .SI(n8701), .SE(n5199), .CLK(n5558), .Q(
        n8700), .QN(n4031) );
  SDFFX1 DFF_196_Q_reg ( .D(n37), .SI(n8700), .SE(n5199), .CLK(n5558), .Q(
        n8699), .QN(n4030) );
  SDFFX1 DFF_197_Q_reg ( .D(n38), .SI(n8699), .SE(n5199), .CLK(n5558), .Q(
        test_so11), .QN(n4029) );
  SDFFX1 DFF_198_Q_reg ( .D(n39), .SI(test_si12), .SE(n5200), .CLK(n5558), .Q(
        n8696), .QN(n4028) );
  SDFFX1 DFF_199_Q_reg ( .D(n40), .SI(n8696), .SE(n5200), .CLK(n5558), .Q(
        n8695), .QN(n4027) );
  SDFFX1 DFF_200_Q_reg ( .D(n41), .SI(n8695), .SE(n5200), .CLK(n5558), .Q(
        n8694), .QN(n4026) );
  SDFFX1 DFF_201_Q_reg ( .D(n42), .SI(n8694), .SE(n5200), .CLK(n5558), .Q(
        n8693), .QN(n4025) );
  SDFFX1 DFF_202_Q_reg ( .D(n43), .SI(n8693), .SE(n5200), .CLK(n5558), .Q(
        n8692), .QN(n4024) );
  SDFFX1 DFF_203_Q_reg ( .D(n44), .SI(n8692), .SE(n5200), .CLK(n5558), .Q(
        n8691), .QN(n4023) );
  SDFFX1 DFF_204_Q_reg ( .D(n45), .SI(n8691), .SE(n5201), .CLK(n5557), .Q(
        n8690), .QN(n4022) );
  SDFFX1 DFF_205_Q_reg ( .D(n46), .SI(n8690), .SE(n5201), .CLK(n5557), .Q(
        n8689), .QN(n4021) );
  SDFFX1 DFF_206_Q_reg ( .D(n47), .SI(n8689), .SE(n5201), .CLK(n5557), .Q(
        n8688), .QN(n4020) );
  SDFFX1 DFF_207_Q_reg ( .D(n48), .SI(n8688), .SE(n5201), .CLK(n5557), .Q(
        n8687), .QN(n4019) );
  SDFFX1 DFF_208_Q_reg ( .D(n49), .SI(n8687), .SE(n5201), .CLK(n5557), .Q(
        n8686), .QN(n4018) );
  SDFFX1 DFF_209_Q_reg ( .D(n50), .SI(n8686), .SE(n5201), .CLK(n5557), .Q(
        n8685), .QN(n4017) );
  SDFFX1 DFF_210_Q_reg ( .D(n51), .SI(n8685), .SE(n5202), .CLK(n5557), .Q(
        n8684), .QN(n4016) );
  SDFFX1 DFF_211_Q_reg ( .D(n52), .SI(n8684), .SE(n5202), .CLK(n5557), .Q(
        n8683), .QN(n4015) );
  SDFFX1 DFF_212_Q_reg ( .D(n53), .SI(n8683), .SE(n5202), .CLK(n5557), .Q(
        n8682), .QN(n4014) );
  SDFFX1 DFF_213_Q_reg ( .D(n54), .SI(n8682), .SE(n5202), .CLK(n5557), .Q(
        n8681), .QN(n4013) );
  SDFFX1 DFF_214_Q_reg ( .D(n55), .SI(n8681), .SE(n5202), .CLK(n5557), .Q(
        n8680), .QN(n4012) );
  SDFFX1 DFF_215_Q_reg ( .D(n56), .SI(n8680), .SE(n5202), .CLK(n5557), .Q(
        test_so12), .QN(n4011) );
  SDFFX1 DFF_216_Q_reg ( .D(n57), .SI(test_si13), .SE(n5203), .CLK(n5556), .Q(
        n8677), .QN(n4010) );
  SDFFX1 DFF_217_Q_reg ( .D(n58), .SI(n8677), .SE(n5203), .CLK(n5556), .Q(
        n8676), .QN(n4009) );
  SDFFX1 DFF_218_Q_reg ( .D(n59), .SI(n8676), .SE(n5203), .CLK(n5556), .Q(
        n8675), .QN(n4008) );
  SDFFX1 DFF_219_Q_reg ( .D(n60), .SI(n8675), .SE(n5203), .CLK(n5556), .Q(
        n8674), .QN(n4007) );
  SDFFX1 DFF_220_Q_reg ( .D(n61), .SI(n8674), .SE(n5203), .CLK(n5556), .Q(
        n8673), .QN(n4006) );
  SDFFX1 DFF_221_Q_reg ( .D(n62), .SI(n8673), .SE(n5203), .CLK(n5556), .Q(
        n8672), .QN(n4005) );
  SDFFX1 DFF_222_Q_reg ( .D(n63), .SI(n8672), .SE(n5204), .CLK(n5556), .Q(
        n8671), .QN(n4004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n5204), .CLK(n5556), .Q(
        n8670), .QN(n4003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n4948), .CLK(n5684), .Q(
        n8669) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n5199), .CLK(n5558), .Q(
        n8668) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n5198), .CLK(n5559), .Q(
        n8667) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n5198), .CLK(n5559), .Q(
        n8666) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n5197), .CLK(n5559), .Q(
        n8665) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n5197), .CLK(n5559), .Q(
        n8664) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n5197), .CLK(n5559), .Q(
        n8663) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n5197), .CLK(n5559), .Q(
        n8662) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n5196), .CLK(n5560), .Q(
        n8661) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n5196), .CLK(n5560), .Q(
        test_so13) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n5195), .CLK(n5560), 
        .Q(n8658) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n5195), .CLK(n5560), .Q(
        n8657) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n5195), .CLK(n5560), .Q(
        n8656) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n5195), .CLK(n5560), .Q(
        n8655) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n4956), .CLK(n5680), .Q(
        n8654) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n4948), .CLK(n5684), .Q(
        n8653) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n5194), .CLK(n5561), .Q(
        WX1970) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n5193), .CLK(n5561), .Q(
        WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n5193), .CLK(n5561), .Q(
        WX1974) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n5193), .CLK(n5561), .Q(
        WX1976) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n5193), .CLK(n5561), .Q(
        WX1978) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n5193), .CLK(n5561), .Q(
        WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n5193), .CLK(n5561), .Q(
        WX1982) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n5192), .CLK(n5562), .Q(
        WX1984) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n5192), .CLK(n5562), .Q(
        WX1986) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n5192), .CLK(n5562), .Q(
        WX1988) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n5192), .CLK(n5562), .Q(
        WX1990) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n5192), .CLK(n5562), .Q(
        test_so14) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n5191), .CLK(n5562), 
        .Q(WX1994) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n5191), .CLK(n5562), .Q(
        WX1996) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n5191), .CLK(n5562), .Q(
        WX1998) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n5190), .CLK(n5563), .Q(
        WX2000) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n5190), .CLK(n5563), .Q(
        WX2002), .QN(n4172) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n5198), .CLK(n5559), .Q(
        WX2004), .QN(n4278) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n5198), .CLK(n5559), .Q(
        WX2006), .QN(n4277) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n5198), .CLK(n5559), .Q(
        WX2008) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n5198), .CLK(n5559), .Q(
        WX2010), .QN(n4275) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n5197), .CLK(n5559), .Q(
        WX2012), .QN(n4274) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n5197), .CLK(n5559), .Q(
        WX2014), .QN(n4273) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n5196), .CLK(n5560), .Q(
        WX2016), .QN(n4272) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n5196), .CLK(n5560), .Q(
        WX2018), .QN(n4271) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n5196), .CLK(n5560), .Q(
        WX2020) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n5196), .CLK(n5560), .Q(
        WX2022), .QN(n4269) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n5195), .CLK(n5560), .Q(
        WX2024), .QN(n4268) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n5195), .CLK(n5560), .Q(
        WX2026), .QN(n4267) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n5194), .CLK(n5561), .Q(
        test_so15), .QN(n9725) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n4956), .CLK(n5680), 
        .Q(WX2030), .QN(n4266) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n4956), .CLK(n5680), .Q(
        WX2032), .QN(n4265) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n4956), .CLK(n5680), .Q(
        WX2034), .QN(n9722) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n4956), .CLK(n5680), .Q(
        WX2036), .QN(n9720) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n4955), .CLK(n5680), .Q(
        WX2038), .QN(n9718) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n4955), .CLK(n5680), .Q(
        WX2040), .QN(n9716) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n4954), .CLK(n5681), .Q(
        WX2042), .QN(n9714) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n4954), .CLK(n5681), .Q(
        WX2044), .QN(n9712) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n4953), .CLK(n5681), .Q(
        WX2046), .QN(n9710) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n4953), .CLK(n5681), .Q(
        WX2048), .QN(n9708) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n4952), .CLK(n5682), .Q(
        WX2050), .QN(n9706) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n4952), .CLK(n5682), .Q(
        WX2052), .QN(n9704) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n4951), .CLK(n5682), .Q(
        WX2054), .QN(n9702) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n5192), .CLK(n5562), .Q(
        WX2056), .QN(n9700) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n5191), .CLK(n5562), .Q(
        WX2058), .QN(n9698) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n5191), .CLK(n5562), .Q(
        WX2060), .QN(n9696) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n5191), .CLK(n5562), .Q(
        WX2062), .QN(n9694) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n5190), .CLK(n5563), .Q(
        test_so16) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n5190), .CLK(n5563), 
        .Q(WX2066) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n5190), .CLK(n5563), .Q(
        WX2068) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n5190), .CLK(n5563), .Q(
        WX2070) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n5189), .CLK(n5563), .Q(
        WX2072), .QN(n4276) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n5189), .CLK(n5563), .Q(
        WX2074) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n5189), .CLK(n5563), .Q(
        WX2076) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n5189), .CLK(n5563), .Q(
        WX2078) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n5188), .CLK(n5564), .Q(
        WX2080) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n5188), .CLK(n5564), .Q(
        WX2082) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n5188), .CLK(n5564), .Q(
        WX2084), .QN(n4270) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n5187), .CLK(n5564), .Q(
        WX2086) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n5187), .CLK(n5564), .Q(
        WX2088) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n5187), .CLK(n5564), .Q(
        WX2090) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n5194), .CLK(n5561), .Q(
        WX2092), .QN(n9726) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n5194), .CLK(n5561), .Q(
        WX2094) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n5194), .CLK(n5561), .Q(
        WX2096) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n5194), .CLK(n5561), .Q(
        WX2098), .QN(n4512) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n4956), .CLK(n5680), .Q(
        test_so17) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n4955), .CLK(n5680), 
        .Q(WX2102), .QN(n4509) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n4955), .CLK(n5680), .Q(
        WX2104), .QN(n4507) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n4954), .CLK(n5681), .Q(
        WX2106), .QN(n4505) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n4954), .CLK(n5681), .Q(
        WX2108), .QN(n4503) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n4953), .CLK(n5681), .Q(
        WX2110), .QN(n4501) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n4953), .CLK(n5681), .Q(
        WX2112), .QN(n4499) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n4952), .CLK(n5682), .Q(
        WX2114), .QN(n4497) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n4952), .CLK(n5682), .Q(
        WX2116), .QN(n4495) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n4951), .CLK(n5682), .Q(
        WX2118), .QN(n4493) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n4951), .CLK(n5682), .Q(
        WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n4950), .CLK(n5683), .Q(
        WX2122), .QN(n4490) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n4950), .CLK(n5683), .Q(
        WX2124), .QN(n4488) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n4950), .CLK(n5683), .Q(
        WX2126), .QN(n4486) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n4949), .CLK(n5683), .Q(
        WX2128), .QN(n9692) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n4949), .CLK(n5683), .Q(
        WX2130), .QN(n4728) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n4949), .CLK(n5683), .Q(
        WX2132), .QN(n4729) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n4949), .CLK(n5683), .Q(
        WX2134), .QN(n4730) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n4949), .CLK(n5683), .Q(
        test_so18) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n5189), .CLK(n5563), 
        .Q(WX2138), .QN(n4731) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n5189), .CLK(n5563), .Q(
        WX2140), .QN(n4732) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n5188), .CLK(n5564), .Q(
        WX2142), .QN(n4733) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n5188), .CLK(n5564), .Q(
        WX2144), .QN(n4734) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n5188), .CLK(n5564), .Q(
        WX2146), .QN(n4735) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n5187), .CLK(n5564), .Q(
        WX2148), .QN(n4736) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n5187), .CLK(n5564), .Q(
        WX2150), .QN(n4737) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n5187), .CLK(n5564), .Q(
        WX2152), .QN(n4738) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n5186), .CLK(n5565), .Q(
        WX2154), .QN(n4739) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n5186), .CLK(n5565), .Q(
        WX2156), .QN(n4740) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n5186), .CLK(n5565), .Q(
        WX2158), .QN(n4741) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n5186), .CLK(n5565), .Q(
        WX2160), .QN(n4531) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n5186), .CLK(n5565), .Q(
        WX2162), .QN(n4742) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n4955), .CLK(n5680), .Q(
        WX2164), .QN(n4743) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n4955), .CLK(n5680), .Q(
        WX2166), .QN(n4744) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n4954), .CLK(n5681), .Q(
        WX2168), .QN(n4745) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n4954), .CLK(n5681), .Q(
        WX2170), .QN(n4532) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n4953), .CLK(n5681), .Q(
        test_so19) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n4953), .CLK(n5681), 
        .Q(WX2174), .QN(n4746) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n4952), .CLK(n5682), .Q(
        WX2176), .QN(n4747) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n4952), .CLK(n5682), .Q(
        WX2178), .QN(n4748) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n4951), .CLK(n5682), .Q(
        WX2180), .QN(n4749) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n4951), .CLK(n5682), .Q(
        WX2182), .QN(n4750) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n4951), .CLK(n5682), .Q(
        WX2184), .QN(n4533) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n4950), .CLK(n5683), .Q(
        WX2186), .QN(n4751) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n4950), .CLK(n5683), .Q(
        WX2188), .QN(n4752) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n4950), .CLK(n5683), .Q(
        WX2190), .QN(n4753) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n4949), .CLK(n5683), .Q(
        WX2192), .QN(n4541) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n4959), .CLK(n5678), .Q(
        CRC_OUT_8_0) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n4959), .CLK(n5678), 
        .Q(CRC_OUT_8_1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n4959), .CLK(n5678), 
        .Q(CRC_OUT_8_2) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n4959), .CLK(n5678), 
        .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n4959), .CLK(n5678), 
        .Q(CRC_OUT_8_4) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n4959), .CLK(n5678), 
        .Q(CRC_OUT_8_5) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n4958), .CLK(n5679), 
        .Q(CRC_OUT_8_6) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n4958), .CLK(n5679), 
        .Q(test_so20) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n4958), .CLK(n5679), 
        .Q(CRC_OUT_8_8) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n4958), .CLK(n5679), 
        .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n4958), .CLK(n5679), 
        .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n4958), .CLK(n5679), .Q(CRC_OUT_8_11) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_12) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_13) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_14) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_16) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n4957), .CLK(n5679), .Q(CRC_OUT_8_17) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n4948), .CLK(n5684), .Q(CRC_OUT_8_18) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n5186), .CLK(n5565), .Q(CRC_OUT_8_19) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n5185), .CLK(n5565), .Q(CRC_OUT_8_20) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n5185), .CLK(n5565), .Q(CRC_OUT_8_21) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n5185), .CLK(n5565), .Q(CRC_OUT_8_22) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n5185), .CLK(n5565), .Q(CRC_OUT_8_23) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n5185), .CLK(n5565), .Q(CRC_OUT_8_24) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n5185), .CLK(n5565), .Q(test_so21) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n5184), .CLK(n5566), 
        .Q(CRC_OUT_8_26) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n5184), .CLK(n5566), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n5184), .CLK(n5566), .Q(CRC_OUT_8_28) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n5184), .CLK(n5566), .Q(CRC_OUT_8_29) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n5184), .CLK(n5566), .Q(CRC_OUT_8_30) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n5184), .CLK(n5566), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n95), .SI(CRC_OUT_8_31), .SE(n5183), .CLK(n5566), 
        .Q(WX3071), .QN(n4820) );
  SDFFX1 DFF_385_Q_reg ( .D(n96), .SI(WX3071), .SE(n5178), .CLK(n5569), .Q(
        n8644), .QN(n4002) );
  SDFFX1 DFF_386_Q_reg ( .D(n97), .SI(n8644), .SE(n5178), .CLK(n5569), .Q(
        n8643), .QN(n4001) );
  SDFFX1 DFF_387_Q_reg ( .D(n98), .SI(n8643), .SE(n5179), .CLK(n5568), .Q(
        n8642), .QN(n4000) );
  SDFFX1 DFF_388_Q_reg ( .D(n99), .SI(n8642), .SE(n5179), .CLK(n5568), .Q(
        n8641), .QN(n3999) );
  SDFFX1 DFF_389_Q_reg ( .D(n100), .SI(n8641), .SE(n5179), .CLK(n5568), .Q(
        n8640), .QN(n3998) );
  SDFFX1 DFF_390_Q_reg ( .D(n101), .SI(n8640), .SE(n5179), .CLK(n5568), .Q(
        n8639), .QN(n3997) );
  SDFFX1 DFF_391_Q_reg ( .D(n102), .SI(n8639), .SE(n5179), .CLK(n5568), .Q(
        n8638), .QN(n3996) );
  SDFFX1 DFF_392_Q_reg ( .D(n103), .SI(n8638), .SE(n5179), .CLK(n5568), .Q(
        n8637), .QN(n3995) );
  SDFFX1 DFF_393_Q_reg ( .D(n104), .SI(n8637), .SE(n5180), .CLK(n5568), .Q(
        n8636), .QN(n3994) );
  SDFFX1 DFF_394_Q_reg ( .D(n105), .SI(n8636), .SE(n5180), .CLK(n5568), .Q(
        n8635), .QN(n3993) );
  SDFFX1 DFF_395_Q_reg ( .D(n106), .SI(n8635), .SE(n5180), .CLK(n5568), .Q(
        test_so22), .QN(n3992) );
  SDFFX1 DFF_396_Q_reg ( .D(n107), .SI(test_si23), .SE(n5180), .CLK(n5568), 
        .Q(n8632), .QN(n3991) );
  SDFFX1 DFF_397_Q_reg ( .D(n108), .SI(n8632), .SE(n5180), .CLK(n5568), .Q(
        n8631), .QN(n3990) );
  SDFFX1 DFF_398_Q_reg ( .D(n109), .SI(n8631), .SE(n5180), .CLK(n5568), .Q(
        n8630), .QN(n3989) );
  SDFFX1 DFF_399_Q_reg ( .D(n110), .SI(n8630), .SE(n5181), .CLK(n5567), .Q(
        n8629), .QN(n3988) );
  SDFFX1 DFF_400_Q_reg ( .D(n112), .SI(n8629), .SE(n5181), .CLK(n5567), .Q(
        n8628), .QN(n3987) );
  SDFFX1 DFF_401_Q_reg ( .D(n113), .SI(n8628), .SE(n5181), .CLK(n5567), .Q(
        n8627), .QN(n3986) );
  SDFFX1 DFF_402_Q_reg ( .D(n114), .SI(n8627), .SE(n5181), .CLK(n5567), .Q(
        n8626), .QN(n3985) );
  SDFFX1 DFF_403_Q_reg ( .D(n115), .SI(n8626), .SE(n5181), .CLK(n5567), .Q(
        n8625), .QN(n3984) );
  SDFFX1 DFF_404_Q_reg ( .D(n116), .SI(n8625), .SE(n5181), .CLK(n5567), .Q(
        n8624), .QN(n3983) );
  SDFFX1 DFF_405_Q_reg ( .D(n117), .SI(n8624), .SE(n5182), .CLK(n5567), .Q(
        n8623), .QN(n3982) );
  SDFFX1 DFF_406_Q_reg ( .D(n118), .SI(n8623), .SE(n5182), .CLK(n5567), .Q(
        n8622), .QN(n3981) );
  SDFFX1 DFF_407_Q_reg ( .D(n119), .SI(n8622), .SE(n5182), .CLK(n5567), .Q(
        n8621), .QN(n3980) );
  SDFFX1 DFF_408_Q_reg ( .D(n120), .SI(n8621), .SE(n5182), .CLK(n5567), .Q(
        n8620), .QN(n3979) );
  SDFFX1 DFF_409_Q_reg ( .D(n121), .SI(n8620), .SE(n5182), .CLK(n5567), .Q(
        n8619), .QN(n3978) );
  SDFFX1 DFF_410_Q_reg ( .D(n122), .SI(n8619), .SE(n5182), .CLK(n5567), .Q(
        n8618), .QN(n3977) );
  SDFFX1 DFF_411_Q_reg ( .D(n123), .SI(n8618), .SE(n5183), .CLK(n5566), .Q(
        n8617), .QN(n3976) );
  SDFFX1 DFF_412_Q_reg ( .D(n124), .SI(n8617), .SE(n5183), .CLK(n5566), .Q(
        n8616), .QN(n3975) );
  SDFFX1 DFF_413_Q_reg ( .D(n125), .SI(n8616), .SE(n5183), .CLK(n5566), .Q(
        test_so23), .QN(n3974) );
  SDFFX1 DFF_414_Q_reg ( .D(n126), .SI(test_si24), .SE(n5183), .CLK(n5566), 
        .Q(n8613), .QN(n3973) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n5183), .CLK(n5566), .Q(
        n8612), .QN(n3972) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n5073), .CLK(n5621), .Q(
        n8611), .QN(n9744) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n5073), .CLK(n5621), .Q(
        n8610), .QN(n9741) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n5052), .CLK(n5632), .Q(
        n8609), .QN(n9740) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n4962), .CLK(n5677), .Q(
        n8608), .QN(n9739) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n4960), .CLK(n5678), .Q(
        n8607), .QN(n9738) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n5071), .CLK(n5622), .Q(
        n8606), .QN(n9735) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n5070), .CLK(n5623), .Q(
        n8605), .QN(n9734) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n5070), .CLK(n5623), .Q(
        n8604), .QN(n9733) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n5048), .CLK(n5634), .Q(
        n8603), .QN(n9732) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n5068), .CLK(n5624), .Q(
        n8602), .QN(n9731) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n5068), .CLK(n5624), .Q(
        n8601), .QN(n9730) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n5067), .CLK(n5624), .Q(
        n8600), .QN(n9729) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n5067), .CLK(n5624), .Q(
        n8599), .QN(n9728) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n4960), .CLK(n5678), .Q(
        n8598), .QN(n9727) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n5082), .CLK(n5617), .Q(
        n8597), .QN(n9724) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n4960), .CLK(n5678), .Q(
        test_so24) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n5081), .CLK(n5617), 
        .Q(WX3263) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n5081), .CLK(n5617), .Q(
        WX3265) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n5081), .CLK(n5617), .Q(
        WX3267) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n5080), .CLK(n5618), .Q(
        WX3269) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n5080), .CLK(n5618), .Q(
        WX3271) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n5080), .CLK(n5618), .Q(
        WX3273) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n5079), .CLK(n5618), .Q(
        WX3275) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n5079), .CLK(n5618), .Q(
        WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n5079), .CLK(n5618), .Q(
        WX3279) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n5078), .CLK(n5619), .Q(
        WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n5078), .CLK(n5619), .Q(
        WX3283) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n5077), .CLK(n5619), .Q(
        WX3285) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n5076), .CLK(n5620), .Q(
        WX3287) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n5076), .CLK(n5620), .Q(
        WX3289) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n5075), .CLK(n5620), .Q(
        WX3291) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n5074), .CLK(n5621), .Q(
        WX3293) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n5074), .CLK(n5621), .Q(
        WX3295), .QN(n4171) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n5073), .CLK(n5621), .Q(
        test_so25), .QN(n9742) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n5052), .CLK(n5632), 
        .Q(WX3299), .QN(n4264) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n4962), .CLK(n5677), .Q(
        WX3301), .QN(n4263) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n4960), .CLK(n5678), .Q(
        WX3303), .QN(n4262) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n5071), .CLK(n5622), .Q(
        WX3305), .QN(n9737) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n5071), .CLK(n5622), .Q(
        WX3307), .QN(n4261) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n5070), .CLK(n5623), .Q(
        WX3309), .QN(n4260) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n5069), .CLK(n5623), .Q(
        WX3311) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n5069), .CLK(n5623), .Q(
        WX3313), .QN(n4258) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n5068), .CLK(n5624), .Q(
        WX3315), .QN(n4257) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n5067), .CLK(n5624), .Q(
        WX3317), .QN(n4256) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n5067), .CLK(n5624), .Q(
        WX3319), .QN(n4255) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n5066), .CLK(n5625), .Q(
        WX3321), .QN(n4254) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n5082), .CLK(n5617), .Q(
        WX3323), .QN(n4253) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n5081), .CLK(n5617), .Q(
        WX3325) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n5081), .CLK(n5617), .Q(
        WX3327), .QN(n9723) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n5081), .CLK(n5617), .Q(
        WX3329), .QN(n9721) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n5080), .CLK(n5618), .Q(
        WX3331), .QN(n9719) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n5080), .CLK(n5618), .Q(
        test_so26) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n5080), .CLK(n5618), 
        .Q(WX3335), .QN(n9715) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n5079), .CLK(n5618), .Q(
        WX3337), .QN(n9713) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n5079), .CLK(n5618), .Q(
        WX3339), .QN(n9711) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n5079), .CLK(n5618), .Q(
        WX3341), .QN(n9709) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n5078), .CLK(n5619), .Q(
        WX3343), .QN(n9707) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n5078), .CLK(n5619), .Q(
        WX3345), .QN(n9705) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n5077), .CLK(n5619), .Q(
        WX3347), .QN(n9703) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n5077), .CLK(n5619), .Q(
        WX3349), .QN(n9701) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n5076), .CLK(n5620), .Q(
        WX3351), .QN(n9699) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n5075), .CLK(n5620), .Q(
        WX3353), .QN(n9697) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n5075), .CLK(n5620), .Q(
        WX3355), .QN(n9695) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n5074), .CLK(n5621), .Q(
        WX3357), .QN(n9693) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n5073), .CLK(n5621), .Q(
        WX3359) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n5073), .CLK(n5621), .Q(
        WX3361), .QN(n9743) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n5072), .CLK(n5622), .Q(
        WX3363) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n5072), .CLK(n5622), .Q(
        WX3365) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n5072), .CLK(n5622), .Q(
        WX3367) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n5071), .CLK(n5622), .Q(
        test_so27), .QN(n9736) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n5070), .CLK(n5623), 
        .Q(WX3371) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n5070), .CLK(n5623), .Q(
        WX3373) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n5069), .CLK(n5623), .Q(
        WX3375), .QN(n4259) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n5069), .CLK(n5623), .Q(
        WX3377) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n5068), .CLK(n5624), .Q(
        WX3379) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n5067), .CLK(n5624), .Q(
        WX3381) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n5066), .CLK(n5625), .Q(
        WX3383) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n5066), .CLK(n5625), .Q(
        WX3385) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n5066), .CLK(n5625), .Q(
        WX3387) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n5065), .CLK(n5625), .Q(
        WX3389), .QN(n4252) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n5065), .CLK(n5625), .Q(
        WX3391), .QN(n4483) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n5065), .CLK(n5625), .Q(
        WX3393), .QN(n4481) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n5064), .CLK(n5626), .Q(
        WX3395), .QN(n4479) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n5064), .CLK(n5626), .Q(
        WX3397), .QN(n9717) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n5064), .CLK(n5626), .Q(
        WX3399), .QN(n4476) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n5063), .CLK(n5626), .Q(
        WX3401), .QN(n4474) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n5063), .CLK(n5626), .Q(
        WX3403), .QN(n4472) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n5063), .CLK(n5626), .Q(
        test_so28) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n5078), .CLK(n5619), 
        .Q(WX3407), .QN(n4469) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n5078), .CLK(n5619), .Q(
        WX3409), .QN(n4467) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n5077), .CLK(n5619), .Q(
        WX3411), .QN(n4465) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n5077), .CLK(n5619), .Q(
        WX3413), .QN(n4463) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n5076), .CLK(n5620), .Q(
        WX3415), .QN(n4461) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n5075), .CLK(n5620), .Q(
        WX3417), .QN(n4459) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n5075), .CLK(n5620), .Q(
        WX3419), .QN(n4457) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n5074), .CLK(n5621), .Q(
        WX3421), .QN(n4455) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n5073), .CLK(n5621), .Q(
        WX3423), .QN(n4702) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n5072), .CLK(n5622), .Q(
        WX3425), .QN(n4703) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n5072), .CLK(n5622), .Q(
        WX3427), .QN(n4704) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n5072), .CLK(n5622), .Q(
        WX3429), .QN(n4705) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n5071), .CLK(n5622), .Q(
        WX3431), .QN(n4706) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n5071), .CLK(n5622), .Q(
        WX3433), .QN(n4707) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n5070), .CLK(n5623), .Q(
        WX3435), .QN(n4708) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n5069), .CLK(n5623), .Q(
        WX3437), .QN(n4709) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n5069), .CLK(n5623), .Q(
        test_so29) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n5068), .CLK(n5624), 
        .Q(WX3441), .QN(n4710) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n5068), .CLK(n5624), .Q(
        WX3443), .QN(n4711) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n5067), .CLK(n5624), .Q(
        WX3445), .QN(n4712) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n5066), .CLK(n5625), .Q(
        WX3447), .QN(n4713) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n5066), .CLK(n5625), .Q(
        WX3449), .QN(n4714) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n5065), .CLK(n5625), .Q(
        WX3451), .QN(n4715) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n5065), .CLK(n5625), .Q(
        WX3453), .QN(n4528) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n5065), .CLK(n5625), .Q(
        WX3455), .QN(n4716) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n5064), .CLK(n5626), .Q(
        WX3457), .QN(n4717) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n5064), .CLK(n5626), .Q(
        WX3459), .QN(n4718) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n5064), .CLK(n5626), .Q(
        WX3461), .QN(n4719) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n5063), .CLK(n5626), .Q(
        WX3463), .QN(n4529) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n5063), .CLK(n5626), .Q(
        WX3465), .QN(n4720) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n5063), .CLK(n5626), .Q(
        WX3467), .QN(n4721) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n5062), .CLK(n5627), .Q(
        WX3469), .QN(n4722) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n5062), .CLK(n5627), .Q(
        WX3471), .QN(n4723) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n5062), .CLK(n5627), .Q(
        test_so30) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n5077), .CLK(n5619), 
        .Q(WX3475), .QN(n4724) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n5076), .CLK(n5620), .Q(
        WX3477), .QN(n4530) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n5076), .CLK(n5620), .Q(
        WX3479), .QN(n4725) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n5075), .CLK(n5620), .Q(
        WX3481), .QN(n4726) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n5074), .CLK(n5621), .Q(
        WX3483), .QN(n4727) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n5074), .CLK(n5621), .Q(
        WX3485), .QN(n4540) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n4962), .CLK(n5677), .Q(
        CRC_OUT_7_0) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_2) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_4) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n4961), .CLK(n5677), 
        .Q(CRC_OUT_7_6) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n4960), .CLK(n5678), 
        .Q(CRC_OUT_7_7) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n5062), .CLK(n5627), 
        .Q(CRC_OUT_7_8) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n5062), .CLK(n5627), 
        .Q(CRC_OUT_7_9) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n5062), .CLK(n5627), 
        .Q(test_so31) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n5061), .CLK(n5627), 
        .Q(CRC_OUT_7_11) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n5061), .CLK(n5627), .Q(CRC_OUT_7_12) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n5061), .CLK(n5627), .Q(CRC_OUT_7_13) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n5061), .CLK(n5627), .Q(CRC_OUT_7_14) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n5061), .CLK(n5627), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n5061), .CLK(n5627), .Q(CRC_OUT_7_16) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_17) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_18) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_19) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_20) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_21) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n5060), .CLK(n5628), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n5059), .CLK(n5628), .Q(CRC_OUT_7_23) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n5059), .CLK(n5628), .Q(CRC_OUT_7_24) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n5059), .CLK(n5628), .Q(CRC_OUT_7_25) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n5059), .CLK(n5628), .Q(CRC_OUT_7_26) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n5059), .CLK(n5628), .Q(test_so32) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n5059), .CLK(n5628), 
        .Q(CRC_OUT_7_28) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n5058), .CLK(n5629), .Q(CRC_OUT_7_29) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n5058), .CLK(n5629), .Q(CRC_OUT_7_30) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n5058), .CLK(n5629), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n158), .SI(CRC_OUT_7_31), .SE(n5058), .CLK(n5629), 
        .Q(WX4364), .QN(n4821) );
  SDFFX1 DFF_577_Q_reg ( .D(n159), .SI(WX4364), .SE(n5053), .CLK(n5631), .Q(
        n8586), .QN(n3971) );
  SDFFX1 DFF_578_Q_reg ( .D(n160), .SI(n8586), .SE(n5053), .CLK(n5631), .Q(
        n8585), .QN(n3970) );
  SDFFX1 DFF_579_Q_reg ( .D(n161), .SI(n8585), .SE(n5053), .CLK(n5631), .Q(
        n8584), .QN(n3969) );
  SDFFX1 DFF_580_Q_reg ( .D(n162), .SI(n8584), .SE(n5053), .CLK(n5631), .Q(
        n8583), .QN(n3968) );
  SDFFX1 DFF_581_Q_reg ( .D(n163), .SI(n8583), .SE(n5053), .CLK(n5631), .Q(
        n8582), .QN(n3967) );
  SDFFX1 DFF_582_Q_reg ( .D(n164), .SI(n8582), .SE(n5054), .CLK(n5631), .Q(
        n8581), .QN(n3966) );
  SDFFX1 DFF_583_Q_reg ( .D(n165), .SI(n8581), .SE(n5054), .CLK(n5631), .Q(
        n8580), .QN(n3965) );
  SDFFX1 DFF_584_Q_reg ( .D(n166), .SI(n8580), .SE(n5054), .CLK(n5631), .Q(
        n8579), .QN(n3964) );
  SDFFX1 DFF_585_Q_reg ( .D(n167), .SI(n8579), .SE(n5054), .CLK(n5631), .Q(
        n8578), .QN(n3963) );
  SDFFX1 DFF_586_Q_reg ( .D(n168), .SI(n8578), .SE(n5054), .CLK(n5631), .Q(
        n8577), .QN(n3962) );
  SDFFX1 DFF_587_Q_reg ( .D(n169), .SI(n8577), .SE(n5054), .CLK(n5631), .Q(
        n8576), .QN(n3961) );
  SDFFX1 DFF_588_Q_reg ( .D(n170), .SI(n8576), .SE(n5055), .CLK(n5630), .Q(
        test_so33), .QN(n3960) );
  SDFFX1 DFF_589_Q_reg ( .D(n171), .SI(test_si34), .SE(n5055), .CLK(n5630), 
        .Q(n8573), .QN(n3959) );
  SDFFX1 DFF_590_Q_reg ( .D(n172), .SI(n8573), .SE(n5055), .CLK(n5630), .Q(
        n8572), .QN(n3958) );
  SDFFX1 DFF_591_Q_reg ( .D(n173), .SI(n8572), .SE(n5055), .CLK(n5630), .Q(
        n8571), .QN(n3957) );
  SDFFX1 DFF_592_Q_reg ( .D(n174), .SI(n8571), .SE(n5055), .CLK(n5630), .Q(
        n8570), .QN(n3956) );
  SDFFX1 DFF_593_Q_reg ( .D(n175), .SI(n8570), .SE(n5055), .CLK(n5630), .Q(
        n8569), .QN(n3955) );
  SDFFX1 DFF_594_Q_reg ( .D(n176), .SI(n8569), .SE(n5056), .CLK(n5630), .Q(
        n8568), .QN(n3954) );
  SDFFX1 DFF_595_Q_reg ( .D(n177), .SI(n8568), .SE(n5056), .CLK(n5630), .Q(
        n8567), .QN(n3953) );
  SDFFX1 DFF_596_Q_reg ( .D(n178), .SI(n8567), .SE(n5056), .CLK(n5630), .Q(
        n8566), .QN(n3952) );
  SDFFX1 DFF_597_Q_reg ( .D(n179), .SI(n8566), .SE(n5056), .CLK(n5630), .Q(
        n8565), .QN(n3951) );
  SDFFX1 DFF_598_Q_reg ( .D(n180), .SI(n8565), .SE(n5056), .CLK(n5630), .Q(
        n8564), .QN(n3950) );
  SDFFX1 DFF_599_Q_reg ( .D(n181), .SI(n8564), .SE(n5056), .CLK(n5630), .Q(
        n8563), .QN(n3949) );
  SDFFX1 DFF_600_Q_reg ( .D(n182), .SI(n8563), .SE(n5057), .CLK(n5629), .Q(
        n8562), .QN(n3948) );
  SDFFX1 DFF_601_Q_reg ( .D(n183), .SI(n8562), .SE(n5057), .CLK(n5629), .Q(
        n8561), .QN(n3947) );
  SDFFX1 DFF_602_Q_reg ( .D(n184), .SI(n8561), .SE(n5057), .CLK(n5629), .Q(
        n8560), .QN(n3946) );
  SDFFX1 DFF_603_Q_reg ( .D(n185), .SI(n8560), .SE(n5057), .CLK(n5629), .Q(
        n8559), .QN(n3945) );
  SDFFX1 DFF_604_Q_reg ( .D(n186), .SI(n8559), .SE(n5057), .CLK(n5629), .Q(
        n8558), .QN(n3944) );
  SDFFX1 DFF_605_Q_reg ( .D(n187), .SI(n8558), .SE(n5057), .CLK(n5629), .Q(
        test_so34), .QN(n3943) );
  SDFFX1 DFF_606_Q_reg ( .D(n188), .SI(test_si35), .SE(n5058), .CLK(n5629), 
        .Q(n8555), .QN(n3942) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n5058), .CLK(n5629), .Q(
        n8554), .QN(n3941) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n4967), .CLK(n5674), .Q(
        n8553), .QN(n9691) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n5053), .CLK(n5631), .Q(
        n8552), .QN(n9688) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n5052), .CLK(n5632), .Q(
        n8551), .QN(n9687) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n5051), .CLK(n5632), .Q(
        n8550), .QN(n9686) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n5050), .CLK(n5633), .Q(
        n8549), .QN(n9685) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n5050), .CLK(n5633), .Q(
        n8548), .QN(n9684) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n5049), .CLK(n5633), .Q(
        n8547), .QN(n9683) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n5049), .CLK(n5633), .Q(
        n8546), .QN(n9682) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n5048), .CLK(n5634), .Q(
        n8545), .QN(n9681) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n5047), .CLK(n5634), .Q(
        n8544), .QN(n9680) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n5046), .CLK(n5635), .Q(
        n8543), .QN(n9679) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n5046), .CLK(n5635), .Q(
        n8542), .QN(n9678) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n5045), .CLK(n5635), .Q(
        n8541), .QN(n9677) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n5045), .CLK(n5635), .Q(
        n8540), .QN(n9676) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n5082), .CLK(n5617), .Q(
        test_so35) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n5043), .CLK(n5636), 
        .Q(n8537), .QN(n9675) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n5043), .CLK(n5636), .Q(
        WX4556) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n5042), .CLK(n5637), .Q(
        WX4558) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n5042), .CLK(n5637), .Q(
        WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n5041), .CLK(n5637), .Q(
        WX4562) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n5040), .CLK(n5638), .Q(
        WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n5040), .CLK(n5638), .Q(
        WX4566) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n5039), .CLK(n5638), .Q(
        WX4568) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n5038), .CLK(n5639), .Q(
        WX4570) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n5038), .CLK(n5639), .Q(
        WX4572) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n5037), .CLK(n5639), .Q(
        WX4574) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n5036), .CLK(n5640), .Q(
        WX4576) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n5036), .CLK(n5640), .Q(
        WX4578) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n5035), .CLK(n5640), .Q(
        WX4580) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n5034), .CLK(n5641), .Q(
        WX4582) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n5034), .CLK(n5641), .Q(
        WX4584) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n5033), .CLK(n5641), .Q(
        test_so36) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n4967), .CLK(n5674), 
        .Q(WX4588), .QN(n4170) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n5052), .CLK(n5632), .Q(
        WX4590), .QN(n9690) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n5052), .CLK(n5632), .Q(
        WX4592), .QN(n4251) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n5051), .CLK(n5632), .Q(
        WX4594) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n5051), .CLK(n5632), .Q(
        WX4596), .QN(n4249) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n5050), .CLK(n5633), .Q(
        WX4598), .QN(n4248) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n5050), .CLK(n5633), .Q(
        WX4600), .QN(n4247) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n5049), .CLK(n5633), .Q(
        WX4602), .QN(n4246) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n5048), .CLK(n5634), .Q(
        WX4604), .QN(n4245) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n5047), .CLK(n5634), .Q(
        WX4606), .QN(n4244) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n5047), .CLK(n5634), .Q(
        WX4608), .QN(n4243) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n5046), .CLK(n5635), .Q(
        WX4610), .QN(n4242) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n5045), .CLK(n5635), .Q(
        WX4612), .QN(n4241) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n5045), .CLK(n5635), .Q(
        WX4614), .QN(n4240) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n5044), .CLK(n5636), .Q(
        WX4616) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n5044), .CLK(n5636), .Q(
        WX4618), .QN(n4238) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n5043), .CLK(n5636), .Q(
        test_so37) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n5042), .CLK(n5637), 
        .Q(WX4622), .QN(n9673) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n5041), .CLK(n5637), .Q(
        WX4624), .QN(n9672) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n5041), .CLK(n5637), .Q(
        WX4626), .QN(n9671) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n5040), .CLK(n5638), .Q(
        WX4628), .QN(n9670) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n5039), .CLK(n5638), .Q(
        WX4630), .QN(n9669) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n5039), .CLK(n5638), .Q(
        WX4632), .QN(n9668) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n5038), .CLK(n5639), .Q(
        WX4634), .QN(n9667) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n5037), .CLK(n5639), .Q(
        WX4636), .QN(n9666) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n5037), .CLK(n5639), .Q(
        WX4638), .QN(n9665) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n5036), .CLK(n5640), .Q(
        WX4640), .QN(n9664) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n5035), .CLK(n5640), .Q(
        WX4642), .QN(n9663) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n5035), .CLK(n5640), .Q(
        WX4644), .QN(n9662) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n5034), .CLK(n5641), .Q(
        WX4646), .QN(n9661) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n5033), .CLK(n5641), .Q(
        WX4648), .QN(n9660) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n5033), .CLK(n5641), .Q(
        WX4650), .QN(n9659) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n5032), .CLK(n5642), .Q(
        WX4652) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n5032), .CLK(n5642), .Q(
        test_so38), .QN(n9689) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n5052), .CLK(n5632), 
        .Q(WX4656) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n5051), .CLK(n5632), .Q(
        WX4658), .QN(n4250) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n5051), .CLK(n5632), .Q(
        WX4660) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n5050), .CLK(n5633), .Q(
        WX4662) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n5049), .CLK(n5633), .Q(
        WX4664) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n5049), .CLK(n5633), .Q(
        WX4666) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n5048), .CLK(n5634), .Q(
        WX4668) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n5047), .CLK(n5634), .Q(
        WX4670) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n5047), .CLK(n5634), .Q(
        WX4672) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n5046), .CLK(n5635), .Q(
        WX4674) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n5045), .CLK(n5635), .Q(
        WX4676) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n5044), .CLK(n5636), .Q(
        WX4678) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n5044), .CLK(n5636), .Q(
        WX4680), .QN(n4239) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n5043), .CLK(n5636), .Q(
        WX4682) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n5043), .CLK(n5636), .Q(
        WX4684), .QN(n9674) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n5042), .CLK(n5637), .Q(
        WX4686), .QN(n4452) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n5041), .CLK(n5637), .Q(
        test_so39) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n5041), .CLK(n5637), 
        .Q(WX4690), .QN(n4449) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n5040), .CLK(n5638), .Q(
        WX4692), .QN(n4447) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n5039), .CLK(n5638), .Q(
        WX4694), .QN(n4445) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n5039), .CLK(n5638), .Q(
        WX4696), .QN(n4443) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n5038), .CLK(n5639), .Q(
        WX4698), .QN(n4441) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n5037), .CLK(n5639), .Q(
        WX4700), .QN(n4439) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n5037), .CLK(n5639), .Q(
        WX4702), .QN(n4437) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n5036), .CLK(n5640), .Q(
        WX4704), .QN(n4435) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n5035), .CLK(n5640), .Q(
        WX4706), .QN(n4433) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n5035), .CLK(n5640), .Q(
        WX4708), .QN(n4431) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n5034), .CLK(n5641), .Q(
        WX4710), .QN(n4429) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n5033), .CLK(n5641), .Q(
        WX4712), .QN(n4427) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n5033), .CLK(n5641), .Q(
        WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n5032), .CLK(n5642), .Q(
        WX4716), .QN(n4675) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n5032), .CLK(n5642), .Q(
        WX4718), .QN(n4676) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n5032), .CLK(n5642), .Q(
        WX4720), .QN(n4677) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n5031), .CLK(n5642), .Q(
        test_so40) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n5051), .CLK(n5632), 
        .Q(WX4724), .QN(n4678) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n5050), .CLK(n5633), .Q(
        WX4726), .QN(n4679) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n5049), .CLK(n5633), .Q(
        WX4728), .QN(n4680) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n5048), .CLK(n5634), .Q(
        WX4730), .QN(n4681) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n5048), .CLK(n5634), .Q(
        WX4732), .QN(n4682) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n5047), .CLK(n5634), .Q(
        WX4734), .QN(n4683) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n5046), .CLK(n5635), .Q(
        WX4736), .QN(n4684) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n5046), .CLK(n5635), .Q(
        WX4738), .QN(n4685) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n5045), .CLK(n5635), .Q(
        WX4740), .QN(n4686) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n5044), .CLK(n5636), .Q(
        WX4742), .QN(n4687) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n5044), .CLK(n5636), .Q(
        WX4744), .QN(n4688) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n5043), .CLK(n5636), .Q(
        WX4746), .QN(n4526) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n5042), .CLK(n5637), .Q(
        WX4748), .QN(n4689) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n5042), .CLK(n5637), .Q(
        WX4750), .QN(n4690) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n5041), .CLK(n5637), .Q(
        WX4752), .QN(n4691) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n5040), .CLK(n5638), .Q(
        WX4754), .QN(n4692) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n5040), .CLK(n5638), .Q(
        test_so41) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n5039), .CLK(n5638), 
        .Q(WX4758), .QN(n4693) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n5038), .CLK(n5639), .Q(
        WX4760), .QN(n4694) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n5038), .CLK(n5639), .Q(
        WX4762), .QN(n4695) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n5037), .CLK(n5639), .Q(
        WX4764), .QN(n4696) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n5036), .CLK(n5640), .Q(
        WX4766), .QN(n4697) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n5036), .CLK(n5640), .Q(
        WX4768), .QN(n4698) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n5035), .CLK(n5640), .Q(
        WX4770), .QN(n4527) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n5034), .CLK(n5641), .Q(
        WX4772), .QN(n4699) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n5034), .CLK(n5641), .Q(
        WX4774), .QN(n4700) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n5033), .CLK(n5641), .Q(
        WX4776), .QN(n4701) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n5032), .CLK(n5642), .Q(
        WX4778), .QN(n4539) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n4967), .CLK(n5674), .Q(
        CRC_OUT_6_0) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n4967), .CLK(n5674), 
        .Q(CRC_OUT_6_1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n4967), .CLK(n5674), 
        .Q(CRC_OUT_6_2) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n4966), .CLK(n5675), 
        .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n4966), .CLK(n5675), 
        .Q(CRC_OUT_6_4) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n4966), .CLK(n5675), 
        .Q(test_so42) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n4966), .CLK(n5675), 
        .Q(CRC_OUT_6_6) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n4966), .CLK(n5675), 
        .Q(CRC_OUT_6_7) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n4966), .CLK(n5675), 
        .Q(CRC_OUT_6_8) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n4965), .CLK(n5675), 
        .Q(CRC_OUT_6_9) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n4965), .CLK(n5675), 
        .Q(CRC_OUT_6_10) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n4965), .CLK(n5675), .Q(CRC_OUT_6_11) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n4965), .CLK(n5675), .Q(CRC_OUT_6_12) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n4965), .CLK(n5675), .Q(CRC_OUT_6_13) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n4965), .CLK(n5675), .Q(CRC_OUT_6_14) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_16) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_17) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_18) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_19) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n4964), .CLK(n5676), .Q(CRC_OUT_6_20) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n4963), .CLK(n5676), .Q(CRC_OUT_6_21) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n4963), .CLK(n5676), .Q(test_so43) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n4963), .CLK(n5676), 
        .Q(CRC_OUT_6_23) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n4963), .CLK(n5676), .Q(CRC_OUT_6_24) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n4963), .CLK(n5676), .Q(CRC_OUT_6_25) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n4963), .CLK(n5676), .Q(CRC_OUT_6_26) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n4962), .CLK(n5677), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n4962), .CLK(n5677), .Q(CRC_OUT_6_28) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n4962), .CLK(n5677), .Q(CRC_OUT_6_29) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n5031), .CLK(n5642), .Q(CRC_OUT_6_30) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n5031), .CLK(n5642), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n220), .SI(CRC_OUT_6_31), .SE(n5031), .CLK(n5642), 
        .Q(WX5657), .QN(n4822) );
  SDFFX1 DFF_769_Q_reg ( .D(n221), .SI(WX5657), .SE(n5026), .CLK(n5645), .Q(
        n8528), .QN(n3940) );
  SDFFX1 DFF_770_Q_reg ( .D(n222), .SI(n8528), .SE(n5026), .CLK(n5645), .Q(
        n8527), .QN(n3939) );
  SDFFX1 DFF_771_Q_reg ( .D(n223), .SI(n8527), .SE(n5026), .CLK(n5645), .Q(
        n8526), .QN(n3938) );
  SDFFX1 DFF_772_Q_reg ( .D(n224), .SI(n8526), .SE(n5026), .CLK(n5645), .Q(
        n8525), .QN(n3937) );
  SDFFX1 DFF_773_Q_reg ( .D(n225), .SI(n8525), .SE(n5026), .CLK(n5645), .Q(
        n8524), .QN(n3936) );
  SDFFX1 DFF_774_Q_reg ( .D(n226), .SI(n8524), .SE(n5027), .CLK(n5644), .Q(
        n8523), .QN(n3935) );
  SDFFX1 DFF_775_Q_reg ( .D(n227), .SI(n8523), .SE(n5027), .CLK(n5644), .Q(
        test_so44), .QN(n3934) );
  SDFFX1 DFF_776_Q_reg ( .D(n228), .SI(test_si45), .SE(n5027), .CLK(n5644), 
        .Q(n8520), .QN(n3933) );
  SDFFX1 DFF_777_Q_reg ( .D(n229), .SI(n8520), .SE(n5027), .CLK(n5644), .Q(
        n8519), .QN(n3932) );
  SDFFX1 DFF_778_Q_reg ( .D(n230), .SI(n8519), .SE(n5027), .CLK(n5644), .Q(
        n8518), .QN(n3931) );
  SDFFX1 DFF_779_Q_reg ( .D(n231), .SI(n8518), .SE(n5027), .CLK(n5644), .Q(
        n8517), .QN(n3930) );
  SDFFX1 DFF_780_Q_reg ( .D(n232), .SI(n8517), .SE(n5028), .CLK(n5644), .Q(
        n8516), .QN(n3929) );
  SDFFX1 DFF_781_Q_reg ( .D(n233), .SI(n8516), .SE(n5028), .CLK(n5644), .Q(
        n8515), .QN(n3928) );
  SDFFX1 DFF_782_Q_reg ( .D(n234), .SI(n8515), .SE(n5028), .CLK(n5644), .Q(
        n8514), .QN(n3927) );
  SDFFX1 DFF_783_Q_reg ( .D(n235), .SI(n8514), .SE(n5028), .CLK(n5644), .Q(
        n8513), .QN(n3926) );
  SDFFX1 DFF_784_Q_reg ( .D(n236), .SI(n8513), .SE(n5028), .CLK(n5644), .Q(
        n8512), .QN(n3925) );
  SDFFX1 DFF_785_Q_reg ( .D(n237), .SI(n8512), .SE(n5028), .CLK(n5644), .Q(
        n8511), .QN(n3924) );
  SDFFX1 DFF_786_Q_reg ( .D(n238), .SI(n8511), .SE(n5029), .CLK(n5643), .Q(
        n8510), .QN(n3923) );
  SDFFX1 DFF_787_Q_reg ( .D(n239), .SI(n8510), .SE(n5029), .CLK(n5643), .Q(
        n8509), .QN(n3922) );
  SDFFX1 DFF_788_Q_reg ( .D(n240), .SI(n8509), .SE(n5029), .CLK(n5643), .Q(
        n8508), .QN(n3921) );
  SDFFX1 DFF_789_Q_reg ( .D(n241), .SI(n8508), .SE(n5029), .CLK(n5643), .Q(
        n8507), .QN(n3920) );
  SDFFX1 DFF_790_Q_reg ( .D(n242), .SI(n8507), .SE(n5029), .CLK(n5643), .Q(
        n8506), .QN(n3919) );
  SDFFX1 DFF_791_Q_reg ( .D(n243), .SI(n8506), .SE(n5029), .CLK(n5643), .Q(
        n8505), .QN(n3918) );
  SDFFX1 DFF_792_Q_reg ( .D(n244), .SI(n8505), .SE(n5030), .CLK(n5643), .Q(
        test_so45), .QN(n3917) );
  SDFFX1 DFF_793_Q_reg ( .D(n245), .SI(test_si46), .SE(n5030), .CLK(n5643), 
        .Q(n8502), .QN(n3916) );
  SDFFX1 DFF_794_Q_reg ( .D(n246), .SI(n8502), .SE(n5030), .CLK(n5643), .Q(
        n8501), .QN(n3915) );
  SDFFX1 DFF_795_Q_reg ( .D(n247), .SI(n8501), .SE(n5030), .CLK(n5643), .Q(
        n8500), .QN(n3914) );
  SDFFX1 DFF_796_Q_reg ( .D(n248), .SI(n8500), .SE(n5030), .CLK(n5643), .Q(
        n8499), .QN(n3913) );
  SDFFX1 DFF_797_Q_reg ( .D(n249), .SI(n8499), .SE(n5030), .CLK(n5643), .Q(
        n8498), .QN(n3912) );
  SDFFX1 DFF_798_Q_reg ( .D(n250), .SI(n8498), .SE(n5031), .CLK(n5642), .Q(
        n8497), .QN(n3911) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n5031), .CLK(n5642), .Q(
        n8496), .QN(n3910) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n4967), .CLK(n5674), .Q(
        n8495), .QN(n9658) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n5026), .CLK(n5645), .Q(
        n8494), .QN(n9657) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n5025), .CLK(n5645), .Q(
        n8493), .QN(n9656) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n5025), .CLK(n5645), .Q(
        n8492), .QN(n9655) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n5024), .CLK(n5646), .Q(
        n8491), .QN(n9654) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n5024), .CLK(n5646), .Q(
        n8490), .QN(n9653) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n5024), .CLK(n5646), .Q(
        n8489), .QN(n9652) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n5024), .CLK(n5646), .Q(
        n8488), .QN(n9651) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n5023), .CLK(n5646), .Q(
        n8487), .QN(n9650) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n5023), .CLK(n5646), .Q(
        test_so46) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n5022), .CLK(n5647), 
        .Q(n8484), .QN(n9649) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n5022), .CLK(n5647), .Q(
        n8483), .QN(n9646) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n4968), .CLK(n5674), .Q(
        n8482), .QN(n9645) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n5021), .CLK(n5647), .Q(
        n8481), .QN(n9642) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n5082), .CLK(n5617), .Q(
        n8480), .QN(n9641) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n4969), .CLK(n5673), .Q(
        n8479), .QN(n9640) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n5020), .CLK(n5648), .Q(
        WX5849) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n5020), .CLK(n5648), .Q(
        WX5851) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n5019), .CLK(n5648), .Q(
        WX5853) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n5018), .CLK(n5649), .Q(
        WX5855) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n5018), .CLK(n5649), .Q(
        WX5857) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n5017), .CLK(n5649), .Q(
        WX5859) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n5016), .CLK(n5650), .Q(
        WX5861) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n5016), .CLK(n5650), .Q(
        WX5863) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n5015), .CLK(n5650), .Q(
        WX5865) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n5014), .CLK(n5651), .Q(
        WX5867) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n5014), .CLK(n5651), .Q(
        test_so47) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n5013), .CLK(n5651), 
        .Q(WX5871) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n5012), .CLK(n5652), .Q(
        WX5873) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n5012), .CLK(n5652), .Q(
        WX5875) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n5011), .CLK(n5652), .Q(
        WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n5010), .CLK(n5653), .Q(
        WX5879) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n5010), .CLK(n5653), .Q(
        WX5881), .QN(n4169) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n5025), .CLK(n5645), .Q(
        WX5883), .QN(n4237) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n5025), .CLK(n5645), .Q(
        WX5885), .QN(n4236) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n5025), .CLK(n5645), .Q(
        WX5887), .QN(n4235) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n5025), .CLK(n5645), .Q(
        WX5889), .QN(n4234) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n5024), .CLK(n5646), .Q(
        WX5891), .QN(n4233) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n5024), .CLK(n5646), .Q(
        WX5893), .QN(n4232) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n5023), .CLK(n5646), .Q(
        WX5895), .QN(n4231) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n5023), .CLK(n5646), .Q(
        WX5897), .QN(n4230) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n5023), .CLK(n5646), .Q(
        WX5899) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n5023), .CLK(n5646), .Q(
        WX5901), .QN(n4228) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n5022), .CLK(n5647), .Q(
        test_so48), .QN(n9647) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n4968), .CLK(n5674), 
        .Q(WX5905), .QN(n4227) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n5021), .CLK(n5647), .Q(
        WX5907), .QN(n9644) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n5021), .CLK(n5647), .Q(
        WX5909), .QN(n4226) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n5021), .CLK(n5647), .Q(
        WX5911) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n5020), .CLK(n5648), .Q(
        WX5913), .QN(n9639) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n5020), .CLK(n5648), .Q(
        WX5915), .QN(n9638) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n5019), .CLK(n5648), .Q(
        WX5917), .QN(n9637) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n5018), .CLK(n5649), .Q(
        WX5919), .QN(n9636) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n5018), .CLK(n5649), .Q(
        WX5921), .QN(n9635) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n5017), .CLK(n5649), .Q(
        WX5923), .QN(n9634) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n5016), .CLK(n5650), .Q(
        WX5925), .QN(n9633) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n5016), .CLK(n5650), .Q(
        WX5927), .QN(n9632) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n5015), .CLK(n5650), .Q(
        WX5929), .QN(n9631) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n5014), .CLK(n5651), .Q(
        WX5931), .QN(n9630) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n5014), .CLK(n5651), .Q(
        WX5933), .QN(n9629) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n5013), .CLK(n5651), .Q(
        WX5935), .QN(n9628) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n5012), .CLK(n5652), .Q(
        test_so49) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n5012), .CLK(n5652), 
        .Q(WX5939), .QN(n9626) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n5011), .CLK(n5652), .Q(
        WX5941), .QN(n9625) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n5010), .CLK(n5653), .Q(
        WX5943), .QN(n9624) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n5010), .CLK(n5653), .Q(
        WX5945) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n5009), .CLK(n5653), .Q(
        WX5947) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n5009), .CLK(n5653), .Q(
        WX5949) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n5009), .CLK(n5653), .Q(
        WX5951) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n5008), .CLK(n5654), .Q(
        WX5953) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n5008), .CLK(n5654), .Q(
        WX5955) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n5008), .CLK(n5654), .Q(
        WX5957) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n5007), .CLK(n5654), .Q(
        WX5959) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n5007), .CLK(n5654), .Q(
        WX5961) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n5007), .CLK(n5654), .Q(
        WX5963), .QN(n4229) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n5006), .CLK(n5655), .Q(
        WX5965) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n5022), .CLK(n5647), .Q(
        WX5967), .QN(n9648) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n5022), .CLK(n5647), .Q(
        WX5969) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n5022), .CLK(n5647), .Q(
        test_so50), .QN(n9643) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n5021), .CLK(n5647), 
        .Q(WX5973) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n5021), .CLK(n5647), .Q(
        WX5975), .QN(n4225) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n5020), .CLK(n5648), .Q(
        WX5977), .QN(n4424) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n5019), .CLK(n5648), .Q(
        WX5979), .QN(n4422) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n5019), .CLK(n5648), .Q(
        WX5981), .QN(n4420) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n5018), .CLK(n5649), .Q(
        WX5983), .QN(n4418) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n5017), .CLK(n5649), .Q(
        WX5985), .QN(n4416) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n5017), .CLK(n5649), .Q(
        WX5987), .QN(n4414) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n5016), .CLK(n5650), .Q(
        WX5989), .QN(n4412) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n5015), .CLK(n5650), .Q(
        WX5991), .QN(n4410) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n5015), .CLK(n5650), .Q(
        WX5993), .QN(n4408) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n5014), .CLK(n5651), .Q(
        WX5995), .QN(n4406) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n5013), .CLK(n5651), .Q(
        WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n5013), .CLK(n5651), .Q(
        WX5999), .QN(n4403) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n5012), .CLK(n5652), .Q(
        WX6001), .QN(n9627) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n5011), .CLK(n5652), .Q(
        WX6003), .QN(n4400) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n5011), .CLK(n5652), .Q(
        test_so51) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n5010), .CLK(n5653), 
        .Q(WX6007), .QN(n4397) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n5009), .CLK(n5653), .Q(
        WX6009), .QN(n4647) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n5009), .CLK(n5653), .Q(
        WX6011), .QN(n4648) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n5009), .CLK(n5653), .Q(
        WX6013), .QN(n4649) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n5008), .CLK(n5654), .Q(
        WX6015), .QN(n4650) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n5008), .CLK(n5654), .Q(
        WX6017), .QN(n4651) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n5008), .CLK(n5654), .Q(
        WX6019), .QN(n4652) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n5007), .CLK(n5654), .Q(
        WX6021), .QN(n4653) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n5007), .CLK(n5654), .Q(
        WX6023), .QN(n4654) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n5007), .CLK(n5654), .Q(
        WX6025), .QN(n4655) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n5006), .CLK(n5655), .Q(
        WX6027), .QN(n4656) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n5006), .CLK(n5655), .Q(
        WX6029), .QN(n4657) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n5006), .CLK(n5655), .Q(
        WX6031), .QN(n4658) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n5006), .CLK(n5655), .Q(
        WX6033), .QN(n4659) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n5006), .CLK(n5655), .Q(
        WX6035), .QN(n4660) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n5005), .CLK(n5655), .Q(
        WX6037), .QN(n4661) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n5005), .CLK(n5655), .Q(
        test_so52) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n5020), .CLK(n5648), 
        .Q(WX6041), .QN(n4662) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n5019), .CLK(n5648), .Q(
        WX6043), .QN(n4663) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n5019), .CLK(n5648), .Q(
        WX6045), .QN(n4664) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n5018), .CLK(n5649), .Q(
        WX6047), .QN(n4665) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n5017), .CLK(n5649), .Q(
        WX6049), .QN(n4524) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n5017), .CLK(n5649), .Q(
        WX6051), .QN(n4666) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n5016), .CLK(n5650), .Q(
        WX6053), .QN(n4667) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n5015), .CLK(n5650), .Q(
        WX6055), .QN(n4668) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n5015), .CLK(n5650), .Q(
        WX6057), .QN(n4669) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n5014), .CLK(n5651), .Q(
        WX6059), .QN(n4670) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n5013), .CLK(n5651), .Q(
        WX6061), .QN(n4671) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n5013), .CLK(n5651), .Q(
        WX6063), .QN(n4525) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n5012), .CLK(n5652), .Q(
        WX6065), .QN(n4672) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n5011), .CLK(n5652), .Q(
        WX6067), .QN(n4673) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n5011), .CLK(n5652), .Q(
        WX6069), .QN(n4674) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n5010), .CLK(n5653), .Q(
        WX6071), .QN(n4538) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n4971), .CLK(n5672), .Q(
        test_so53) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n4971), .CLK(n5672), 
        .Q(CRC_OUT_5_1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n4971), .CLK(n5672), 
        .Q(CRC_OUT_5_2) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n4971), .CLK(n5672), 
        .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n4971), .CLK(n5672), 
        .Q(CRC_OUT_5_4) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n4971), .CLK(n5672), 
        .Q(CRC_OUT_5_5) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n4970), .CLK(n5673), 
        .Q(CRC_OUT_5_6) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n4970), .CLK(n5673), 
        .Q(CRC_OUT_5_7) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n4970), .CLK(n5673), 
        .Q(CRC_OUT_5_8) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n4970), .CLK(n5673), 
        .Q(CRC_OUT_5_9) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n4970), .CLK(n5673), 
        .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n4970), .CLK(n5673), .Q(CRC_OUT_5_11) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n4969), .CLK(n5673), .Q(CRC_OUT_5_12) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n4969), .CLK(n5673), .Q(CRC_OUT_5_13) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n4969), .CLK(n5673), .Q(CRC_OUT_5_14) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n4969), .CLK(n5673), .Q(CRC_OUT_5_15) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n4969), .CLK(n5673), .Q(CRC_OUT_5_16) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n4968), .CLK(n5674), .Q(test_so54) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n4968), .CLK(n5674), 
        .Q(CRC_OUT_5_18) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n4968), .CLK(n5674), .Q(CRC_OUT_5_19) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n4968), .CLK(n5674), .Q(CRC_OUT_5_20) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n5005), .CLK(n5655), .Q(CRC_OUT_5_21) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n5005), .CLK(n5655), .Q(CRC_OUT_5_22) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n5005), .CLK(n5655), .Q(CRC_OUT_5_23) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n5005), .CLK(n5655), .Q(CRC_OUT_5_24) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_25) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_26) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_27) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_28) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_29) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n5004), .CLK(n5656), .Q(CRC_OUT_5_30) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n5003), .CLK(n5656), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n282), .SI(CRC_OUT_5_31), .SE(n5003), .CLK(n5656), 
        .Q(WX6950), .QN(n4823) );
  SDFFX1 DFF_961_Q_reg ( .D(n283), .SI(WX6950), .SE(n4998), .CLK(n5659), .Q(
        n8470), .QN(n3909) );
  SDFFX1 DFF_962_Q_reg ( .D(n284), .SI(n8470), .SE(n4998), .CLK(n5659), .Q(
        test_so55), .QN(n3908) );
  SDFFX1 DFF_963_Q_reg ( .D(n285), .SI(test_si56), .SE(n4998), .CLK(n5659), 
        .Q(n8467), .QN(n3907) );
  SDFFX1 DFF_964_Q_reg ( .D(n286), .SI(n8467), .SE(n4999), .CLK(n5658), .Q(
        n8466), .QN(n3906) );
  SDFFX1 DFF_965_Q_reg ( .D(n287), .SI(n8466), .SE(n4999), .CLK(n5658), .Q(
        n8465), .QN(n3905) );
  SDFFX1 DFF_966_Q_reg ( .D(n288), .SI(n8465), .SE(n4999), .CLK(n5658), .Q(
        n8464), .QN(n3904) );
  SDFFX1 DFF_967_Q_reg ( .D(n289), .SI(n8464), .SE(n4999), .CLK(n5658), .Q(
        n8463), .QN(n3903) );
  SDFFX1 DFF_968_Q_reg ( .D(n290), .SI(n8463), .SE(n4999), .CLK(n5658), .Q(
        n8462), .QN(n3902) );
  SDFFX1 DFF_969_Q_reg ( .D(n291), .SI(n8462), .SE(n4999), .CLK(n5658), .Q(
        n8461), .QN(n3901) );
  SDFFX1 DFF_970_Q_reg ( .D(n292), .SI(n8461), .SE(n5000), .CLK(n5658), .Q(
        n8460), .QN(n3900) );
  SDFFX1 DFF_971_Q_reg ( .D(n293), .SI(n8460), .SE(n5000), .CLK(n5658), .Q(
        n8459), .QN(n3899) );
  SDFFX1 DFF_972_Q_reg ( .D(n294), .SI(n8459), .SE(n5000), .CLK(n5658), .Q(
        n8458), .QN(n3898) );
  SDFFX1 DFF_973_Q_reg ( .D(n295), .SI(n8458), .SE(n5000), .CLK(n5658), .Q(
        n8457), .QN(n3897) );
  SDFFX1 DFF_974_Q_reg ( .D(n296), .SI(n8457), .SE(n5000), .CLK(n5658), .Q(
        n8456), .QN(n3896) );
  SDFFX1 DFF_975_Q_reg ( .D(n297), .SI(n8456), .SE(n5000), .CLK(n5658), .Q(
        n8455), .QN(n3895) );
  SDFFX1 DFF_976_Q_reg ( .D(n298), .SI(n8455), .SE(n5001), .CLK(n5657), .Q(
        n8454), .QN(n3894) );
  SDFFX1 DFF_977_Q_reg ( .D(n299), .SI(n8454), .SE(n5001), .CLK(n5657), .Q(
        n8453), .QN(n3893) );
  SDFFX1 DFF_978_Q_reg ( .D(n300), .SI(n8453), .SE(n5001), .CLK(n5657), .Q(
        n8452), .QN(n3892) );
  SDFFX1 DFF_979_Q_reg ( .D(n301), .SI(n8452), .SE(n5001), .CLK(n5657), .Q(
        test_so56), .QN(n3891) );
  SDFFX1 DFF_980_Q_reg ( .D(n302), .SI(test_si57), .SE(n5001), .CLK(n5657), 
        .Q(n8449), .QN(n3890) );
  SDFFX1 DFF_981_Q_reg ( .D(n303), .SI(n8449), .SE(n5001), .CLK(n5657), .Q(
        n8448), .QN(n3889) );
  SDFFX1 DFF_982_Q_reg ( .D(n304), .SI(n8448), .SE(n5002), .CLK(n5657), .Q(
        n8447), .QN(n3888) );
  SDFFX1 DFF_983_Q_reg ( .D(n305), .SI(n8447), .SE(n5002), .CLK(n5657), .Q(
        n8446), .QN(n3887) );
  SDFFX1 DFF_984_Q_reg ( .D(n306), .SI(n8446), .SE(n5002), .CLK(n5657), .Q(
        n8445), .QN(n3886) );
  SDFFX1 DFF_985_Q_reg ( .D(WX6999), .SI(n8445), .SE(n5002), .CLK(n5657), .Q(
        n8444), .QN(n3885) );
  SDFFX1 DFF_986_Q_reg ( .D(n308), .SI(n8444), .SE(n5002), .CLK(n5657), .Q(
        n8443) );
  SDFFX1 DFF_987_Q_reg ( .D(n309), .SI(n8443), .SE(n5002), .CLK(n5657), .Q(
        n8442), .QN(n3883) );
  SDFFX1 DFF_988_Q_reg ( .D(n310), .SI(n8442), .SE(n5003), .CLK(n5656), .Q(
        n8441), .QN(n3882) );
  SDFFX1 DFF_989_Q_reg ( .D(n311), .SI(n8441), .SE(n5003), .CLK(n5656), .Q(
        n8440), .QN(n3881) );
  SDFFX1 DFF_990_Q_reg ( .D(n312), .SI(n8440), .SE(n5003), .CLK(n5656), .Q(
        n8439), .QN(n3880) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n5003), .CLK(n5656), .Q(
        n8438), .QN(n3879) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n4972), .CLK(n5672), .Q(
        n8437), .QN(n9623) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n4998), .CLK(n5659), .Q(
        n8436), .QN(n9622) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n4997), .CLK(n5659), .Q(
        n8435), .QN(n9621) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n4997), .CLK(n5659), .Q(
        n8434), .QN(n9620) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n4972), .CLK(n5672), .Q(
        test_so57) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n4997), .CLK(n5659), 
        .Q(n8431), .QN(n9619) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n4996), .CLK(n5660), .Q(
        n8430), .QN(n9616) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n4972), .CLK(n5672), .Q(
        n8429), .QN(n9615) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n4996), .CLK(n5660), .Q(
        n8428), .QN(n9612) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n4995), .CLK(n5660), .Q(
        n8427), .QN(n9611) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n4995), .CLK(n5660), .Q(
        n8426), .QN(n9610) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n4994), .CLK(n5661), .Q(
        n8425), .QN(n9609) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n4994), .CLK(n5661), .Q(
        n8424), .QN(n9608) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n4972), .CLK(n5672), .Q(
        n8423), .QN(n9607) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n5082), .CLK(n5617), .Q(
        n8422), .QN(n9606) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n4991), .CLK(n5662), .Q(
        n8421), .QN(n9605) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n4991), .CLK(n5662), .Q(
        WX7142) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n4991), .CLK(n5662), 
        .Q(WX7144) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n4990), .CLK(n5663), 
        .Q(WX7146) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n4989), .CLK(n5663), 
        .Q(WX7148) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n4989), .CLK(n5663), 
        .Q(WX7150) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n4988), .CLK(n5664), 
        .Q(test_so58) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n4987), .CLK(n5664), 
        .Q(WX7154) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n4987), .CLK(n5664), 
        .Q(WX7156) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n4986), .CLK(n5665), 
        .Q(WX7158) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n4985), .CLK(n5665), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n4985), .CLK(n5665), 
        .Q(WX7162) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n4984), .CLK(n5666), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n4983), .CLK(n5666), 
        .Q(WX7166) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n4983), .CLK(n5666), 
        .Q(WX7168) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n4982), .CLK(n5667), 
        .Q(WX7170) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n4981), .CLK(n5667), 
        .Q(WX7172) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n4981), .CLK(n5667), 
        .Q(WX7174), .QN(n4168) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n4998), .CLK(n5659), 
        .Q(WX7176), .QN(n4224) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n4998), .CLK(n5659), 
        .Q(WX7178), .QN(n4223) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n4997), .CLK(n5659), 
        .Q(WX7180), .QN(n4222) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n4997), .CLK(n5659), 
        .Q(WX7182) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n4997), .CLK(n5659), 
        .Q(WX7184), .QN(n4220) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n4996), .CLK(n5660), 
        .Q(test_so59), .QN(n9617) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n4972), .CLK(n5672), 
        .Q(WX7188), .QN(n4219) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n4995), .CLK(n5660), 
        .Q(WX7190), .QN(n9614) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n4995), .CLK(n5660), 
        .Q(WX7192), .QN(n4218) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n4995), .CLK(n5660), 
        .Q(WX7194) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n4994), .CLK(n5661), 
        .Q(WX7196), .QN(n4216) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n4993), .CLK(n5661), 
        .Q(WX7198), .QN(n4215) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n4993), .CLK(n5661), 
        .Q(WX7200), .QN(n4214) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n4992), .CLK(n5662), 
        .Q(WX7202), .QN(n4213) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n4992), .CLK(n5662), 
        .Q(WX7204), .QN(n4212) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n4991), .CLK(n5662), 
        .Q(WX7206), .QN(n9604) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n4990), .CLK(n5663), 
        .Q(WX7208), .QN(n9603) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n4990), .CLK(n5663), 
        .Q(WX7210), .QN(n9602) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n4989), .CLK(n5663), 
        .Q(WX7212), .QN(n9601) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n4988), .CLK(n5664), 
        .Q(WX7214), .QN(n9600) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n4988), .CLK(n5664), 
        .Q(WX7216), .QN(n9599) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n4987), .CLK(n5664), 
        .Q(WX7218), .QN(n9598) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n4986), .CLK(n5665), 
        .Q(test_so60) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n4986), .CLK(n5665), 
        .Q(WX7222), .QN(n9596) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n4985), .CLK(n5665), 
        .Q(WX7224), .QN(n9595) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n4984), .CLK(n5666), 
        .Q(WX7226), .QN(n9594) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n4984), .CLK(n5666), 
        .Q(WX7228), .QN(n9593) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n4983), .CLK(n5666), 
        .Q(WX7230), .QN(n9592) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n4982), .CLK(n5667), 
        .Q(WX7232), .QN(n9591) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n4982), .CLK(n5667), 
        .Q(WX7234), .QN(n9590) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n4981), .CLK(n5667), 
        .Q(WX7236), .QN(n9589) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n4980), .CLK(n5668), 
        .Q(WX7238) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n4980), .CLK(n5668), 
        .Q(WX7240) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n4980), .CLK(n5668), 
        .Q(WX7242) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n4979), .CLK(n5668), 
        .Q(WX7244) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n4979), .CLK(n5668), 
        .Q(WX7246), .QN(n4221) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n4979), .CLK(n5668), 
        .Q(WX7248) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n4996), .CLK(n5660), 
        .Q(WX7250), .QN(n9618) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n4996), .CLK(n5660), 
        .Q(WX7252) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n4996), .CLK(n5660), 
        .Q(test_so61), .QN(n9613) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n4995), .CLK(n5660), 
        .Q(WX7256) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n4994), .CLK(n5661), 
        .Q(WX7258), .QN(n4217) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n4994), .CLK(n5661), 
        .Q(WX7260) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n4993), .CLK(n5661), 
        .Q(WX7262) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n4993), .CLK(n5661), 
        .Q(WX7264) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n4992), .CLK(n5662), 
        .Q(WX7266) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n4992), .CLK(n5662), 
        .Q(WX7268) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n4991), .CLK(n5662), 
        .Q(WX7270), .QN(n4395) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n4990), .CLK(n5663), 
        .Q(WX7272), .QN(n4393) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n4990), .CLK(n5663), 
        .Q(WX7274), .QN(n4391) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n4989), .CLK(n5663), 
        .Q(WX7276), .QN(n4389) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n4988), .CLK(n5664), 
        .Q(WX7278), .QN(n4387) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n4988), .CLK(n5664), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n4987), .CLK(n5664), 
        .Q(WX7282), .QN(n4384) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n4986), .CLK(n5665), 
        .Q(WX7284), .QN(n9597) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n4986), .CLK(n5665), 
        .Q(WX7286), .QN(n4381) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n4985), .CLK(n5665), 
        .Q(test_so62) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n4984), .CLK(n5666), 
        .Q(WX7290), .QN(n4378) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n4984), .CLK(n5666), 
        .Q(WX7292), .QN(n4376) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n4983), .CLK(n5666), 
        .Q(WX7294), .QN(n4374) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n4982), .CLK(n5667), 
        .Q(WX7296), .QN(n4372) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n4982), .CLK(n5667), 
        .Q(WX7298), .QN(n4370) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n4981), .CLK(n5667), 
        .Q(WX7300), .QN(n4368) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n4980), .CLK(n5668), 
        .Q(WX7302), .QN(n4620) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n4980), .CLK(n5668), 
        .Q(WX7304), .QN(n4621) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n4980), .CLK(n5668), 
        .Q(WX7306), .QN(n4622) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n4979), .CLK(n5668), 
        .Q(WX7308), .QN(n4623) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n4979), .CLK(n5668), 
        .Q(WX7310), .QN(n4624) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n4979), .CLK(n5668), 
        .Q(WX7312), .QN(n4625) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n4978), .CLK(n5669), 
        .Q(WX7314), .QN(n4626) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n4978), .CLK(n5669), 
        .Q(WX7316), .QN(n4627) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n4978), .CLK(n5669), 
        .Q(WX7318), .QN(n4628) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n4978), .CLK(n5669), 
        .Q(WX7320), .QN(n4629) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n4978), .CLK(n5669), 
        .Q(test_so63) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n4994), .CLK(n5661), 
        .Q(WX7324), .QN(n4630) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n4993), .CLK(n5661), 
        .Q(WX7326), .QN(n4631) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n4993), .CLK(n5661), 
        .Q(WX7328), .QN(n4632) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n4992), .CLK(n5662), 
        .Q(WX7330), .QN(n4633) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n4992), .CLK(n5662), 
        .Q(WX7332), .QN(n4522) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n4991), .CLK(n5662), 
        .Q(WX7334), .QN(n4634) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n4990), .CLK(n5663), 
        .Q(WX7336), .QN(n4635) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n4989), .CLK(n5663), 
        .Q(WX7338), .QN(n4636) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n4989), .CLK(n5663), 
        .Q(WX7340), .QN(n4637) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n4988), .CLK(n5664), 
        .Q(WX7342), .QN(n4523) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n4987), .CLK(n5664), 
        .Q(WX7344), .QN(n4638) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n4987), .CLK(n5664), 
        .Q(WX7346), .QN(n4639) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n4986), .CLK(n5665), 
        .Q(WX7348), .QN(n4640) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n4985), .CLK(n5665), 
        .Q(WX7350), .QN(n4641) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n4985), .CLK(n5665), 
        .Q(WX7352), .QN(n4642) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n4984), .CLK(n5666), 
        .Q(WX7354), .QN(n4643) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n4983), .CLK(n5666), 
        .Q(test_so64) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n4983), .CLK(n5666), 
        .Q(WX7358), .QN(n4644) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n4982), .CLK(n5667), 
        .Q(WX7360), .QN(n4645) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n4981), .CLK(n5667), 
        .Q(WX7362), .QN(n4646) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n4981), .CLK(n5667), 
        .Q(WX7364), .QN(n4537) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n4977), .CLK(n5669), 
        .Q(CRC_OUT_4_0) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_2) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_3) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_4) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_5) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n4976), .CLK(n5670), .Q(CRC_OUT_4_6) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n4975), .CLK(n5670), .Q(CRC_OUT_4_7) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n4975), .CLK(n5670), .Q(CRC_OUT_4_8) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n4975), .CLK(n5670), .Q(CRC_OUT_4_9) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n4975), .CLK(n5670), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n4975), .CLK(
        n5670), .Q(CRC_OUT_4_11) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n4975), .CLK(
        n5670), .Q(test_so65) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n4974), .CLK(n5671), 
        .Q(CRC_OUT_4_13) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n4974), .CLK(
        n5671), .Q(CRC_OUT_4_14) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n4974), .CLK(
        n5671), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n4974), .CLK(
        n5671), .Q(CRC_OUT_4_16) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n4974), .CLK(
        n5671), .Q(CRC_OUT_4_17) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n4974), .CLK(
        n5671), .Q(CRC_OUT_4_18) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_19) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_21) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_22) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_23) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n4973), .CLK(
        n5671), .Q(CRC_OUT_4_24) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n4972), .CLK(
        n5672), .Q(CRC_OUT_4_25) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n4978), .CLK(
        n5669), .Q(CRC_OUT_4_26) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n4977), .CLK(
        n5669), .Q(CRC_OUT_4_27) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n4977), .CLK(
        n5669), .Q(CRC_OUT_4_28) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n4977), .CLK(
        n5669), .Q(test_so66) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n4977), .CLK(n5669), 
        .Q(CRC_OUT_4_30) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n4977), .CLK(
        n5669), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n344), .SI(CRC_OUT_4_31), .SE(n5176), .CLK(n5570), 
        .Q(WX8243), .QN(n4824) );
  SDFFX1 DFF_1153_Q_reg ( .D(n345), .SI(WX8243), .SE(n5176), .CLK(n5570), .Q(
        n8411), .QN(n3878) );
  SDFFX1 DFF_1154_Q_reg ( .D(n346), .SI(n8411), .SE(n5176), .CLK(n5570), .Q(
        n8410), .QN(n3877) );
  SDFFX1 DFF_1155_Q_reg ( .D(n347), .SI(n8410), .SE(n5177), .CLK(n5569), .Q(
        n8409), .QN(n3876) );
  SDFFX1 DFF_1156_Q_reg ( .D(n348), .SI(n8409), .SE(n5177), .CLK(n5569), .Q(
        n8408), .QN(n3875) );
  SDFFX1 DFF_1157_Q_reg ( .D(n349), .SI(n8408), .SE(n5177), .CLK(n5569), .Q(
        n8407), .QN(n3874) );
  SDFFX1 DFF_1158_Q_reg ( .D(n350), .SI(n8407), .SE(n5177), .CLK(n5569), .Q(
        n8406), .QN(n3873) );
  SDFFX1 DFF_1159_Q_reg ( .D(n351), .SI(n8406), .SE(n5177), .CLK(n5569), .Q(
        n8405), .QN(n3872) );
  SDFFX1 DFF_1160_Q_reg ( .D(n352), .SI(n8405), .SE(n5177), .CLK(n5569), .Q(
        n8404), .QN(n3871) );
  SDFFX1 DFF_1161_Q_reg ( .D(n353), .SI(n8404), .SE(n5178), .CLK(n5569), .Q(
        n8403), .QN(n3870) );
  SDFFX1 DFF_1162_Q_reg ( .D(n354), .SI(n8403), .SE(n5178), .CLK(n5569), .Q(
        n8402), .QN(n3869) );
  SDFFX1 DFF_1163_Q_reg ( .D(n355), .SI(n8402), .SE(n5178), .CLK(n5569), .Q(
        n8401), .QN(n3868) );
  SDFFX1 DFF_1164_Q_reg ( .D(WX8266), .SI(n8401), .SE(n5178), .CLK(n5569), .Q(
        n8400), .QN(n3867) );
  SDFFX1 DFF_1165_Q_reg ( .D(n357), .SI(n8400), .SE(n4960), .CLK(n5678), .Q(
        n8399) );
  SDFFX1 DFF_1166_Q_reg ( .D(n358), .SI(n8399), .SE(n5173), .CLK(n5571), .Q(
        test_so67), .QN(n3865) );
  SDFFX1 DFF_1167_Q_reg ( .D(n359), .SI(test_si68), .SE(n5173), .CLK(n5571), 
        .Q(n8396), .QN(n3864) );
  SDFFX1 DFF_1168_Q_reg ( .D(n360), .SI(n8396), .SE(n5173), .CLK(n5571), .Q(
        n8395), .QN(n3863) );
  SDFFX1 DFF_1169_Q_reg ( .D(n361), .SI(n8395), .SE(n5174), .CLK(n5571), .Q(
        n8394), .QN(n3862) );
  SDFFX1 DFF_1170_Q_reg ( .D(n362), .SI(n8394), .SE(n5174), .CLK(n5571), .Q(
        n8393), .QN(n3861) );
  SDFFX1 DFF_1171_Q_reg ( .D(n363), .SI(n8393), .SE(n5174), .CLK(n5571), .Q(
        n8392), .QN(n3860) );
  SDFFX1 DFF_1172_Q_reg ( .D(n364), .SI(n8392), .SE(n5174), .CLK(n5571), .Q(
        n8391), .QN(n3859) );
  SDFFX1 DFF_1173_Q_reg ( .D(n365), .SI(n8391), .SE(n5174), .CLK(n5571), .Q(
        n8390), .QN(n3858) );
  SDFFX1 DFF_1174_Q_reg ( .D(n366), .SI(n8390), .SE(n5174), .CLK(n5571), .Q(
        n8389), .QN(n3857) );
  SDFFX1 DFF_1175_Q_reg ( .D(n367), .SI(n8389), .SE(n5175), .CLK(n5570), .Q(
        n8388), .QN(n3856) );
  SDFFX1 DFF_1176_Q_reg ( .D(n368), .SI(n8388), .SE(n5175), .CLK(n5570), .Q(
        n8387), .QN(n3855) );
  SDFFX1 DFF_1177_Q_reg ( .D(n369), .SI(n8387), .SE(n5175), .CLK(n5570), .Q(
        n8386), .QN(n3854) );
  SDFFX1 DFF_1178_Q_reg ( .D(n370), .SI(n8386), .SE(n5175), .CLK(n5570), .Q(
        n8385), .QN(n3853) );
  SDFFX1 DFF_1179_Q_reg ( .D(n371), .SI(n8385), .SE(n5175), .CLK(n5570), .Q(
        n8384), .QN(n3852) );
  SDFFX1 DFF_1180_Q_reg ( .D(n372), .SI(n8384), .SE(n5175), .CLK(n5570), .Q(
        n8383), .QN(n3851) );
  SDFFX1 DFF_1181_Q_reg ( .D(n373), .SI(n8383), .SE(n5176), .CLK(n5570), .Q(
        n8382), .QN(n3850) );
  SDFFX1 DFF_1182_Q_reg ( .D(n374), .SI(n8382), .SE(n5176), .CLK(n5570), .Q(
        n8381), .QN(n3849) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n5176), .CLK(n5570), .Q(
        test_so68), .QN(n3848) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n5163), .CLK(n5576), 
        .Q(n8378), .QN(n9588) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n5163), .CLK(n5576), .Q(
        n8377), .QN(n9585) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n5143), .CLK(n5586), .Q(
        n8376), .QN(n9584) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n5162), .CLK(n5577), .Q(
        n8375), .QN(n9581) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n5161), .CLK(n5577), .Q(
        n8374), .QN(n9580) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n5161), .CLK(n5577), .Q(
        n8373), .QN(n9579) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n5159), .CLK(n5578), .Q(
        n8372), .QN(n9578) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n5159), .CLK(n5578), .Q(
        n8371), .QN(n9577) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n5158), .CLK(n5579), .Q(
        n8370), .QN(n9576) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n5158), .CLK(n5579), .Q(
        n8369), .QN(n9575) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n5157), .CLK(n5579), .Q(
        n8368), .QN(n9574) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n5157), .CLK(n5579), .Q(
        n8367), .QN(n9573) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n5155), .CLK(n5580), .Q(
        n8366), .QN(n9572) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n5155), .CLK(n5580), .Q(
        n8365), .QN(n9571) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n5173), .CLK(n5571), .Q(
        n8364), .QN(n9570) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n5172), .CLK(n5572), .Q(
        n8363), .QN(n9569) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n5172), .CLK(n5572), .Q(
        test_so69) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n5172), .CLK(n5572), 
        .Q(WX8437) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n5172), .CLK(n5572), 
        .Q(WX8439) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n5171), .CLK(n5572), 
        .Q(WX8441) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n5171), .CLK(n5572), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n5171), .CLK(n5572), 
        .Q(WX8445) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n5170), .CLK(n5573), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n5170), .CLK(n5573), 
        .Q(WX8449) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n5169), .CLK(n5573), 
        .Q(WX8451) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n5168), .CLK(n5574), 
        .Q(WX8453) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n5168), .CLK(n5574), 
        .Q(WX8455) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n5167), .CLK(n5574), 
        .Q(WX8457) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n5166), .CLK(n5575), 
        .Q(WX8459) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n5166), .CLK(n5575), 
        .Q(WX8461) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n5165), .CLK(n5575), 
        .Q(WX8463) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n5164), .CLK(n5576), 
        .Q(WX8465) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n5164), .CLK(n5576), 
        .Q(WX8467), .QN(n4167) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n5163), .CLK(n5576), 
        .Q(test_so70), .QN(n9586) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n5142), .CLK(n5587), 
        .Q(WX8471), .QN(n4211) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n5161), .CLK(n5577), 
        .Q(WX8473), .QN(n9583) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n5161), .CLK(n5577), 
        .Q(WX8475), .QN(n4210) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n5160), .CLK(n5578), 
        .Q(WX8477) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n5160), .CLK(n5578), 
        .Q(WX8479), .QN(n4208) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n5159), .CLK(n5578), 
        .Q(WX8481), .QN(n4207) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n5159), .CLK(n5578), 
        .Q(WX8483), .QN(n4206) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n5158), .CLK(n5579), 
        .Q(WX8485), .QN(n4205) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n5157), .CLK(n5579), 
        .Q(WX8487), .QN(n4204) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n5156), .CLK(n5580), 
        .Q(WX8489), .QN(n4203) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n5156), .CLK(n5580), 
        .Q(WX8491), .QN(n4202) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n5155), .CLK(n5580), 
        .Q(WX8493), .QN(n4201) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n5173), .CLK(n5571), 
        .Q(WX8495), .QN(n4200) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n5173), .CLK(n5571), 
        .Q(WX8497), .QN(n4199) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n5172), .CLK(n5572), 
        .Q(WX8499), .QN(n9568) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n5172), .CLK(n5572), 
        .Q(WX8501), .QN(n9567) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n5171), .CLK(n5572), 
        .Q(test_so71) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n5171), .CLK(n5572), 
        .Q(WX8505), .QN(n9565) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n5171), .CLK(n5572), 
        .Q(WX8507), .QN(n9564) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n5170), .CLK(n5573), 
        .Q(WX8509), .QN(n9563) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n5170), .CLK(n5573), 
        .Q(WX8511), .QN(n9562) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n5169), .CLK(n5573), 
        .Q(WX8513), .QN(n9561) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n5169), .CLK(n5573), 
        .Q(WX8515), .QN(n9560) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n5168), .CLK(n5574), 
        .Q(WX8517), .QN(n9559) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n5167), .CLK(n5574), 
        .Q(WX8519), .QN(n9558) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n5167), .CLK(n5574), 
        .Q(WX8521), .QN(n9557) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n5166), .CLK(n5575), 
        .Q(WX8523), .QN(n9556) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n5165), .CLK(n5575), 
        .Q(WX8525), .QN(n9555) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n5165), .CLK(n5575), 
        .Q(WX8527), .QN(n9554) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n5164), .CLK(n5576), 
        .Q(WX8529), .QN(n9553) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n5163), .CLK(n5576), 
        .Q(WX8531) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n5163), .CLK(n5576), 
        .Q(WX8533), .QN(n9587) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n5162), .CLK(n5577), 
        .Q(WX8535) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n5162), .CLK(n5577), 
        .Q(test_so72), .QN(n9582) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n5161), .CLK(n5577), 
        .Q(WX8539) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n5160), .CLK(n5578), 
        .Q(WX8541), .QN(n4209) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n5160), .CLK(n5578), 
        .Q(WX8543) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n5159), .CLK(n5578), 
        .Q(WX8545) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n5158), .CLK(n5579), 
        .Q(WX8547) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n5158), .CLK(n5579), 
        .Q(WX8549) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n5157), .CLK(n5579), 
        .Q(WX8551) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n5156), .CLK(n5580), 
        .Q(WX8553) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n5156), .CLK(n5580), 
        .Q(WX8555) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n5155), .CLK(n5580), 
        .Q(WX8557) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n5155), .CLK(n5580), 
        .Q(WX8559) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n5154), .CLK(n5581), 
        .Q(WX8561) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n5154), .CLK(n5581), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n5154), .CLK(n5581), 
        .Q(WX8565), .QN(n4365) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n5153), .CLK(n5581), 
        .Q(WX8567), .QN(n9566) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n5153), .CLK(n5581), 
        .Q(WX8569), .QN(n4362) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n5153), .CLK(n5581), 
        .Q(test_so73) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n5170), .CLK(n5573), 
        .Q(WX8573), .QN(n4359) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n5170), .CLK(n5573), 
        .Q(WX8575), .QN(n4357) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n5169), .CLK(n5573), 
        .Q(WX8577), .QN(n4355) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n5169), .CLK(n5573), 
        .Q(WX8579), .QN(n4353) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n5168), .CLK(n5574), 
        .Q(WX8581), .QN(n4351) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n5167), .CLK(n5574), 
        .Q(WX8583), .QN(n4349) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n5167), .CLK(n5574), 
        .Q(WX8585), .QN(n4347) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n5166), .CLK(n5575), 
        .Q(WX8587), .QN(n4345) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n5165), .CLK(n5575), 
        .Q(WX8589), .QN(n4343) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n5165), .CLK(n5575), 
        .Q(WX8591), .QN(n4341) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n5164), .CLK(n5576), 
        .Q(WX8593), .QN(n4339) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n5163), .CLK(n5576), 
        .Q(WX8595), .QN(n4594) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n5162), .CLK(n5577), 
        .Q(WX8597), .QN(n4595) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n5162), .CLK(n5577), 
        .Q(WX8599), .QN(n4596) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n5162), .CLK(n5577), 
        .Q(WX8601), .QN(n4597) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n5161), .CLK(n5577), 
        .Q(WX8603), .QN(n4598) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n5160), .CLK(n5578), 
        .Q(test_so74) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n5160), .CLK(n5578), 
        .Q(WX8607), .QN(n4599) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n5159), .CLK(n5578), 
        .Q(WX8609), .QN(n4600) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n5158), .CLK(n5579), 
        .Q(WX8611), .QN(n4601) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n5157), .CLK(n5579), 
        .Q(WX8613), .QN(n4602) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n5157), .CLK(n5579), 
        .Q(WX8615), .QN(n4603) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n5156), .CLK(n5580), 
        .Q(WX8617), .QN(n4604) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n5156), .CLK(n5580), 
        .Q(WX8619), .QN(n4605) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n5155), .CLK(n5580), 
        .Q(WX8621), .QN(n4606) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n5154), .CLK(n5581), 
        .Q(WX8623), .QN(n4607) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n5154), .CLK(n5581), 
        .Q(WX8625), .QN(n4519) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n5154), .CLK(n5581), 
        .Q(WX8627), .QN(n4608) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n5153), .CLK(n5581), 
        .Q(WX8629), .QN(n4609) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n5153), .CLK(n5581), 
        .Q(WX8631), .QN(n4610) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n5153), .CLK(n5581), 
        .Q(WX8633), .QN(n4611) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n5152), .CLK(n5582), 
        .Q(WX8635), .QN(n4520) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n5152), .CLK(n5582), 
        .Q(WX8637), .QN(n4612) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n5152), .CLK(n5582), 
        .Q(test_so75) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n5169), .CLK(n5573), 
        .Q(WX8641), .QN(n4613) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n5168), .CLK(n5574), 
        .Q(WX8643), .QN(n4614) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n5168), .CLK(n5574), 
        .Q(WX8645), .QN(n4615) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n5167), .CLK(n5574), 
        .Q(WX8647), .QN(n4616) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n5166), .CLK(n5575), 
        .Q(WX8649), .QN(n4521) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n5166), .CLK(n5575), 
        .Q(WX8651), .QN(n4617) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n5165), .CLK(n5575), 
        .Q(WX8653), .QN(n4618) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n5164), .CLK(n5576), 
        .Q(WX8655), .QN(n4619) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n5164), .CLK(n5576), 
        .Q(WX8657), .QN(n4536) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n5084), .CLK(n5616), 
        .Q(CRC_OUT_3_0) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n5084), .CLK(n5616), .Q(CRC_OUT_3_1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n5084), .CLK(n5616), .Q(CRC_OUT_3_2) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n5084), .CLK(n5616), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n5083), .CLK(n5616), .Q(CRC_OUT_3_4) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n5083), .CLK(n5616), .Q(CRC_OUT_3_5) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n5083), .CLK(n5616), .Q(CRC_OUT_3_6) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n5083), .CLK(n5616), .Q(test_so76) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n5083), .CLK(n5616), 
        .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n5083), .CLK(n5616), .Q(CRC_OUT_3_9) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n5082), .CLK(n5617), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n5152), .CLK(
        n5582), .Q(CRC_OUT_3_11) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n5152), .CLK(
        n5582), .Q(CRC_OUT_3_12) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n5152), .CLK(
        n5582), .Q(CRC_OUT_3_13) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_14) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_16) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_17) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_18) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n5151), .CLK(
        n5582), .Q(CRC_OUT_3_19) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n5150), .CLK(
        n5583), .Q(CRC_OUT_3_20) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n5150), .CLK(
        n5583), .Q(CRC_OUT_3_21) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n5150), .CLK(
        n5583), .Q(CRC_OUT_3_22) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n5150), .CLK(
        n5583), .Q(CRC_OUT_3_23) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n5150), .CLK(
        n5583), .Q(test_so77) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n5150), .CLK(n5583), 
        .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_26) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_27) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_28) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_29) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_30) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n5149), .CLK(
        n5583), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n406), .SI(CRC_OUT_3_31), .SE(n5148), .CLK(n5584), 
        .Q(WX9536), .QN(n4825) );
  SDFFX1 DFF_1345_Q_reg ( .D(n407), .SI(WX9536), .SE(n5143), .CLK(n5586), .Q(
        n8353), .QN(n3847) );
  SDFFX1 DFF_1346_Q_reg ( .D(n408), .SI(n8353), .SE(n5143), .CLK(n5586), .Q(
        n8352), .QN(n3846) );
  SDFFX1 DFF_1347_Q_reg ( .D(n409), .SI(n8352), .SE(n5144), .CLK(n5586), .Q(
        n8351), .QN(n3845) );
  SDFFX1 DFF_1348_Q_reg ( .D(n410), .SI(n8351), .SE(n5144), .CLK(n5586), .Q(
        n8350), .QN(n3844) );
  SDFFX1 DFF_1349_Q_reg ( .D(n411), .SI(n8350), .SE(n5144), .CLK(n5586), .Q(
        n8349), .QN(n3843) );
  SDFFX1 DFF_1350_Q_reg ( .D(n412), .SI(n8349), .SE(n5144), .CLK(n5586), .Q(
        n8348), .QN(n3842) );
  SDFFX1 DFF_1351_Q_reg ( .D(n413), .SI(n8348), .SE(n5144), .CLK(n5586), .Q(
        n8347), .QN(n3841) );
  SDFFX1 DFF_1352_Q_reg ( .D(n414), .SI(n8347), .SE(n5144), .CLK(n5586), .Q(
        n8346), .QN(n3840) );
  SDFFX1 DFF_1353_Q_reg ( .D(n415), .SI(n8346), .SE(n5145), .CLK(n5585), .Q(
        test_so78), .QN(n3839) );
  SDFFX1 DFF_1354_Q_reg ( .D(n416), .SI(test_si79), .SE(n5145), .CLK(n5585), 
        .Q(n8343), .QN(n3838) );
  SDFFX1 DFF_1355_Q_reg ( .D(n417), .SI(n8343), .SE(n5145), .CLK(n5585), .Q(
        n8342), .QN(n3837) );
  SDFFX1 DFF_1356_Q_reg ( .D(n418), .SI(n8342), .SE(n5145), .CLK(n5585), .Q(
        n8341), .QN(n3836) );
  SDFFX1 DFF_1357_Q_reg ( .D(n419), .SI(n8341), .SE(n5145), .CLK(n5585), .Q(
        n8340), .QN(n3835) );
  SDFFX1 DFF_1358_Q_reg ( .D(n420), .SI(n8340), .SE(n5145), .CLK(n5585), .Q(
        n8339), .QN(n3834) );
  SDFFX1 DFF_1359_Q_reg ( .D(n421), .SI(n8339), .SE(n5146), .CLK(n5585), .Q(
        n8338), .QN(n3833) );
  SDFFX1 DFF_1360_Q_reg ( .D(n422), .SI(n8338), .SE(n5146), .CLK(n5585), .Q(
        n8337), .QN(n3832) );
  SDFFX1 DFF_1361_Q_reg ( .D(n423), .SI(n8337), .SE(n5146), .CLK(n5585), .Q(
        n8336), .QN(n3831) );
  SDFFX1 DFF_1362_Q_reg ( .D(n424), .SI(n8336), .SE(n5146), .CLK(n5585), .Q(
        n8335), .QN(n3830) );
  SDFFX1 DFF_1363_Q_reg ( .D(n425), .SI(n8335), .SE(n5146), .CLK(n5585), .Q(
        n8334), .QN(n3829) );
  SDFFX1 DFF_1364_Q_reg ( .D(n426), .SI(n8334), .SE(n5146), .CLK(n5585), .Q(
        n8333), .QN(n3828) );
  SDFFX1 DFF_1365_Q_reg ( .D(n427), .SI(n8333), .SE(n5147), .CLK(n5584), .Q(
        n8332), .QN(n3827) );
  SDFFX1 DFF_1366_Q_reg ( .D(n428), .SI(n8332), .SE(n5147), .CLK(n5584), .Q(
        n8331), .QN(n3826) );
  SDFFX1 DFF_1367_Q_reg ( .D(n429), .SI(n8331), .SE(n5147), .CLK(n5584), .Q(
        n8330), .QN(n3825) );
  SDFFX1 DFF_1368_Q_reg ( .D(n430), .SI(n8330), .SE(n5147), .CLK(n5584), .Q(
        n8329), .QN(n3824) );
  SDFFX1 DFF_1369_Q_reg ( .D(n431), .SI(n8329), .SE(n5147), .CLK(n5584), .Q(
        n8328), .QN(n3823) );
  SDFFX1 DFF_1370_Q_reg ( .D(n432), .SI(n8328), .SE(n5147), .CLK(n5584), .Q(
        test_so79), .QN(n3822) );
  SDFFX1 DFF_1371_Q_reg ( .D(n433), .SI(test_si80), .SE(n5148), .CLK(n5584), 
        .Q(n8325), .QN(n3821) );
  SDFFX1 DFF_1372_Q_reg ( .D(n434), .SI(n8325), .SE(n5148), .CLK(n5584), .Q(
        n8324), .QN(n3820) );
  SDFFX1 DFF_1373_Q_reg ( .D(n435), .SI(n8324), .SE(n5148), .CLK(n5584), .Q(
        n8323), .QN(n3819) );
  SDFFX1 DFF_1374_Q_reg ( .D(n436), .SI(n8323), .SE(n5148), .CLK(n5584), .Q(
        n8322), .QN(n3818) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n5148), .CLK(n5584), .Q(
        n8321), .QN(n3817) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n5084), .CLK(n5616), .Q(
        n8320), .QN(n9552) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n5143), .CLK(n5586), .Q(
        n8319), .QN(n9551) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n5142), .CLK(n5587), .Q(
        n8318), .QN(n9550) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n5142), .CLK(n5587), .Q(
        n8317), .QN(n9549) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n5142), .CLK(n5587), .Q(
        n8316), .QN(n9548) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n5141), .CLK(n5587), .Q(
        n8315), .QN(n9547) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n5141), .CLK(n5587), .Q(
        n8314), .QN(n9546) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n5141), .CLK(n5587), .Q(
        n8313), .QN(n9545) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n5140), .CLK(n5588), .Q(
        n8312), .QN(n9544) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n5140), .CLK(n5588), .Q(
        n8311), .QN(n9543) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n5140), .CLK(n5588), .Q(
        n8310), .QN(n9542) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n5139), .CLK(n5588), .Q(
        test_so80) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n5139), .CLK(n5588), 
        .Q(n8307), .QN(n9541) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n5139), .CLK(n5588), .Q(
        n8306), .QN(n9538) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n5085), .CLK(n5615), .Q(
        n8305), .QN(n9537) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n5138), .CLK(n5589), .Q(
        n8304), .QN(n9534) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n5137), .CLK(n5589), .Q(
        WX9728) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n5137), .CLK(n5589), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n5137), .CLK(n5589), 
        .Q(WX9732) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n5136), .CLK(n5590), 
        .Q(WX9734) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n5135), .CLK(n5590), 
        .Q(WX9736) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n5135), .CLK(n5590), 
        .Q(WX9738) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n5134), .CLK(n5591), 
        .Q(WX9740) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n5133), .CLK(n5591), 
        .Q(WX9742) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n5133), .CLK(n5591), 
        .Q(WX9744) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n5132), .CLK(n5592), 
        .Q(WX9746) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n5131), .CLK(n5592), 
        .Q(WX9748) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n5131), .CLK(n5592), 
        .Q(WX9750) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n5130), .CLK(n5593), 
        .Q(test_so81) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n5129), .CLK(n5593), 
        .Q(WX9754) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n5129), .CLK(n5593), 
        .Q(WX9756) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n5128), .CLK(n5594), 
        .Q(WX9758) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n5127), .CLK(n5594), 
        .Q(WX9760) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n5143), .CLK(n5586), 
        .Q(WX9762), .QN(n4198) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n5143), .CLK(n5586), 
        .Q(WX9764), .QN(n4197) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n5142), .CLK(n5587), 
        .Q(WX9766), .QN(n4196) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n5142), .CLK(n5587), 
        .Q(WX9768), .QN(n4195) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n5141), .CLK(n5587), 
        .Q(WX9770), .QN(n4194) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n5141), .CLK(n5587), 
        .Q(WX9772), .QN(n4193) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n5141), .CLK(n5587), 
        .Q(WX9774), .QN(n4192) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n5140), .CLK(n5588), 
        .Q(WX9776), .QN(n4191) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n5140), .CLK(n5588), 
        .Q(WX9778), .QN(n4190) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n5140), .CLK(n5588), 
        .Q(WX9780), .QN(n4189) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n5139), .CLK(n5588), 
        .Q(WX9782) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n5139), .CLK(n5588), 
        .Q(WX9784), .QN(n4187) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n5139), .CLK(n5588), 
        .Q(test_so82), .QN(n9539) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n5084), .CLK(n5616), 
        .Q(WX9788), .QN(n4186) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n5138), .CLK(n5589), 
        .Q(WX9790), .QN(n9536) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n5138), .CLK(n5589), 
        .Q(WX9792), .QN(n9533) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n5137), .CLK(n5589), 
        .Q(WX9794), .QN(n9532) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n5136), .CLK(n5590), 
        .Q(WX9796), .QN(n9531) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n5136), .CLK(n5590), 
        .Q(WX9798), .QN(n9530) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n5135), .CLK(n5590), 
        .Q(WX9800), .QN(n9529) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n5134), .CLK(n5591), 
        .Q(WX9802), .QN(n9528) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n5134), .CLK(n5591), 
        .Q(WX9804), .QN(n9527) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n5133), .CLK(n5591), 
        .Q(WX9806), .QN(n9526) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n5132), .CLK(n5592), 
        .Q(WX9808), .QN(n9525) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n5132), .CLK(n5592), 
        .Q(WX9810), .QN(n9524) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n5131), .CLK(n5592), 
        .Q(WX9812), .QN(n9523) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n5130), .CLK(n5593), 
        .Q(WX9814), .QN(n9522) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n5130), .CLK(n5593), 
        .Q(WX9816), .QN(n9521) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n5129), .CLK(n5593), 
        .Q(WX9818), .QN(n9520) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n5128), .CLK(n5594), 
        .Q(test_so83) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n5128), .CLK(n5594), 
        .Q(WX9822), .QN(n9518) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n5127), .CLK(n5594), 
        .Q(WX9824), .QN(n4166) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n5127), .CLK(n5594), 
        .Q(WX9826) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n5126), .CLK(n5595), 
        .Q(WX9828) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n5126), .CLK(n5595), 
        .Q(WX9830) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n5126), .CLK(n5595), 
        .Q(WX9832) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n5125), .CLK(n5595), 
        .Q(WX9834) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n5125), .CLK(n5595), 
        .Q(WX9836) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n5125), .CLK(n5595), 
        .Q(WX9838) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n5124), .CLK(n5596), 
        .Q(WX9840) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n5124), .CLK(n5596), 
        .Q(WX9842) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n5124), .CLK(n5596), 
        .Q(WX9844) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n5123), .CLK(n5596), 
        .Q(WX9846), .QN(n4188) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n5123), .CLK(n5596), 
        .Q(WX9848) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n5138), .CLK(n5589), 
        .Q(WX9850), .QN(n9540) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n5138), .CLK(n5589), 
        .Q(WX9852) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n5138), .CLK(n5589), 
        .Q(test_so84), .QN(n9535) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n5137), .CLK(n5589), 
        .Q(WX9856), .QN(n4337) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n5137), .CLK(n5589), 
        .Q(WX9858), .QN(n4335) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n5136), .CLK(n5590), 
        .Q(WX9860), .QN(n4333) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n5136), .CLK(n5590), 
        .Q(WX9862), .QN(n4331) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n5135), .CLK(n5590), 
        .Q(WX9864), .QN(n4329) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n5134), .CLK(n5591), 
        .Q(WX9866), .QN(n4327) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n5134), .CLK(n5591), 
        .Q(WX9868), .QN(n4325) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n5133), .CLK(n5591), 
        .Q(WX9870), .QN(n4323) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n5132), .CLK(n5592), 
        .Q(WX9872), .QN(n4321) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n5132), .CLK(n5592), 
        .Q(WX9874), .QN(n4319) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n5131), .CLK(n5592), 
        .Q(WX9876), .QN(n4317) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n5130), .CLK(n5593), 
        .Q(WX9878), .QN(n4315) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n5130), .CLK(n5593), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n5129), .CLK(n5593), 
        .Q(WX9882), .QN(n4312) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n5128), .CLK(n5594), 
        .Q(WX9884), .QN(n9519) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n5128), .CLK(n5594), 
        .Q(WX9886), .QN(n4309) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n5127), .CLK(n5594), 
        .Q(test_so85) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n5127), .CLK(n5594), 
        .Q(WX9890), .QN(n4568) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n5126), .CLK(n5595), 
        .Q(WX9892), .QN(n4569) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n5126), .CLK(n5595), 
        .Q(WX9894), .QN(n4570) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n5126), .CLK(n5595), 
        .Q(WX9896), .QN(n4571) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n5125), .CLK(n5595), 
        .Q(WX9898), .QN(n4572) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n5125), .CLK(n5595), 
        .Q(WX9900), .QN(n4573) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n5125), .CLK(n5595), 
        .Q(WX9902), .QN(n4574) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n5124), .CLK(n5596), 
        .Q(WX9904), .QN(n4575) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n5124), .CLK(n5596), 
        .Q(WX9906), .QN(n4576) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n5124), .CLK(n5596), 
        .Q(WX9908), .QN(n4577) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n5123), .CLK(n5596), 
        .Q(WX9910), .QN(n4578) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n5123), .CLK(n5596), 
        .Q(WX9912), .QN(n4579) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n5123), .CLK(n5596), 
        .Q(WX9914), .QN(n4580) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n5123), .CLK(n5596), 
        .Q(WX9916), .QN(n4581) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n5122), .CLK(n5597), 
        .Q(WX9918), .QN(n4516) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n5122), .CLK(n5597), 
        .Q(WX9920), .QN(n4582) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n5122), .CLK(n5597), 
        .Q(test_so86) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n5136), .CLK(n5590), 
        .Q(WX9924), .QN(n4583) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n5135), .CLK(n5590), 
        .Q(WX9926), .QN(n4584) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n5135), .CLK(n5590), 
        .Q(WX9928), .QN(n4517) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n5134), .CLK(n5591), 
        .Q(WX9930), .QN(n4585) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n5133), .CLK(n5591), 
        .Q(WX9932), .QN(n4586) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n5133), .CLK(n5591), 
        .Q(WX9934), .QN(n4587) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n5132), .CLK(n5592), 
        .Q(WX9936), .QN(n4588) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n5131), .CLK(n5592), 
        .Q(WX9938), .QN(n4589) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n5131), .CLK(n5592), 
        .Q(WX9940), .QN(n4590) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n5130), .CLK(n5593), 
        .Q(WX9942), .QN(n4518) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n5129), .CLK(n5593), 
        .Q(WX9944), .QN(n4591) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n5129), .CLK(n5593), 
        .Q(WX9946), .QN(n4592) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n5128), .CLK(n5594), 
        .Q(WX9948), .QN(n4593) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n5127), .CLK(n5594), 
        .Q(WX9950), .QN(n4535) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n5088), .CLK(n5614), 
        .Q(CRC_OUT_2_0) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n5088), .CLK(
        n5614), .Q(CRC_OUT_2_1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n5087), .CLK(
        n5614), .Q(test_so87) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n5087), .CLK(n5614), 
        .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n5087), .CLK(
        n5614), .Q(CRC_OUT_2_4) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n5087), .CLK(
        n5614), .Q(CRC_OUT_2_5) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n5087), .CLK(
        n5614), .Q(CRC_OUT_2_6) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n5087), .CLK(
        n5614), .Q(CRC_OUT_2_7) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_8) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_9) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_11) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_12) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n5086), .CLK(
        n5615), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n5085), .CLK(
        n5615), .Q(CRC_OUT_2_14) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n5085), .CLK(
        n5615), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n5085), .CLK(
        n5615), .Q(CRC_OUT_2_16) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n5085), .CLK(
        n5615), .Q(CRC_OUT_2_17) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n5085), .CLK(
        n5615), .Q(CRC_OUT_2_18) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n5122), .CLK(
        n5597), .Q(test_so88) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n5122), .CLK(n5597), 
        .Q(CRC_OUT_2_20) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n5122), .CLK(
        n5597), .Q(CRC_OUT_2_21) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_22) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_23) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_24) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_25) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_26) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n5121), .CLK(
        n5597), .Q(CRC_OUT_2_27) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n5120), .CLK(
        n5598), .Q(CRC_OUT_2_28) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n5120), .CLK(
        n5598), .Q(CRC_OUT_2_29) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n5120), .CLK(
        n5598), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n5120), .CLK(
        n5598), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n468), .SI(CRC_OUT_2_31), .SE(n5120), .CLK(n5598), 
        .Q(WX10829), .QN(n4826) );
  SDFFX1 DFF_1537_Q_reg ( .D(n469), .SI(WX10829), .SE(n5115), .CLK(n5600), .Q(
        n8295), .QN(n3816) );
  SDFFX1 DFF_1538_Q_reg ( .D(n470), .SI(n8295), .SE(n5115), .CLK(n5600), .Q(
        n8294), .QN(n3815) );
  SDFFX1 DFF_1539_Q_reg ( .D(n471), .SI(n8294), .SE(n5115), .CLK(n5600), .Q(
        n8293), .QN(n3814) );
  SDFFX1 DFF_1540_Q_reg ( .D(n472), .SI(n8293), .SE(n5115), .CLK(n5600), .Q(
        test_so89), .QN(n3813) );
  SDFFX1 DFF_1541_Q_reg ( .D(n473), .SI(test_si90), .SE(n5115), .CLK(n5600), 
        .Q(n8290), .QN(n3812) );
  SDFFX1 DFF_1542_Q_reg ( .D(n474), .SI(n8290), .SE(n5115), .CLK(n5600), .Q(
        n8289), .QN(n3811) );
  SDFFX1 DFF_1543_Q_reg ( .D(n475), .SI(n8289), .SE(n5116), .CLK(n5600), .Q(
        n8288), .QN(n3810) );
  SDFFX1 DFF_1544_Q_reg ( .D(n476), .SI(n8288), .SE(n5116), .CLK(n5600), .Q(
        n8287), .QN(n3809) );
  SDFFX1 DFF_1545_Q_reg ( .D(n477), .SI(n8287), .SE(n5116), .CLK(n5600), .Q(
        n8286), .QN(n3808) );
  SDFFX1 DFF_1546_Q_reg ( .D(n478), .SI(n8286), .SE(n5116), .CLK(n5600), .Q(
        n8285), .QN(n3807) );
  SDFFX1 DFF_1547_Q_reg ( .D(n479), .SI(n8285), .SE(n5116), .CLK(n5600), .Q(
        n8284), .QN(n3806) );
  SDFFX1 DFF_1548_Q_reg ( .D(n480), .SI(n8284), .SE(n5116), .CLK(n5600), .Q(
        n8283), .QN(n3805) );
  SDFFX1 DFF_1549_Q_reg ( .D(n481), .SI(n8283), .SE(n5117), .CLK(n5599), .Q(
        n8282), .QN(n3804) );
  SDFFX1 DFF_1550_Q_reg ( .D(n482), .SI(n8282), .SE(n5117), .CLK(n5599), .Q(
        n8281), .QN(n3803) );
  SDFFX1 DFF_1551_Q_reg ( .D(n483), .SI(n8281), .SE(n5117), .CLK(n5599), .Q(
        n8280), .QN(n3802) );
  SDFFX1 DFF_1552_Q_reg ( .D(n484), .SI(n8280), .SE(n5117), .CLK(n5599), .Q(
        n8279), .QN(n3801) );
  SDFFX1 DFF_1553_Q_reg ( .D(n485), .SI(n8279), .SE(n5117), .CLK(n5599), .Q(
        n8278), .QN(n3800) );
  SDFFX1 DFF_1554_Q_reg ( .D(n486), .SI(n8278), .SE(n5117), .CLK(n5599), .Q(
        n8277), .QN(n3799) );
  SDFFX1 DFF_1555_Q_reg ( .D(n487), .SI(n8277), .SE(n5118), .CLK(n5599), .Q(
        n8276), .QN(n3798) );
  SDFFX1 DFF_1556_Q_reg ( .D(n488), .SI(n8276), .SE(n5118), .CLK(n5599), .Q(
        n8275), .QN(n3797) );
  SDFFX1 DFF_1557_Q_reg ( .D(n489), .SI(n8275), .SE(n5118), .CLK(n5599), .Q(
        test_so90), .QN(n3796) );
  SDFFX1 DFF_1558_Q_reg ( .D(n490), .SI(test_si91), .SE(n5118), .CLK(n5599), 
        .Q(n8272), .QN(n3795) );
  SDFFX1 DFF_1559_Q_reg ( .D(n491), .SI(n8272), .SE(n5118), .CLK(n5599), .Q(
        n8271), .QN(n3794) );
  SDFFX1 DFF_1560_Q_reg ( .D(n492), .SI(n8271), .SE(n5118), .CLK(n5599), .Q(
        n8270), .QN(n3793) );
  SDFFX1 DFF_1561_Q_reg ( .D(n493), .SI(n8270), .SE(n5119), .CLK(n5598), .Q(
        n8269), .QN(n3792) );
  SDFFX1 DFF_1562_Q_reg ( .D(n494), .SI(n8269), .SE(n5119), .CLK(n5598), .Q(
        n8268), .QN(n3791) );
  SDFFX1 DFF_1563_Q_reg ( .D(n495), .SI(n8268), .SE(n5119), .CLK(n5598), .Q(
        n8267), .QN(n3790) );
  SDFFX1 DFF_1564_Q_reg ( .D(n496), .SI(n8267), .SE(n5119), .CLK(n5598), .Q(
        n8266), .QN(n3789) );
  SDFFX1 DFF_1565_Q_reg ( .D(n497), .SI(n8266), .SE(n5119), .CLK(n5598), .Q(
        n8265), .QN(n3788) );
  SDFFX1 DFF_1566_Q_reg ( .D(n498), .SI(n8265), .SE(n5119), .CLK(n5598), .Q(
        n8264), .QN(n3787) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n5120), .CLK(n5598), 
        .Q(n8263), .QN(n3786) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n5088), .CLK(n5614), 
        .Q(n8262) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n5114), .CLK(n5601), 
        .Q(n8261) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n5114), .CLK(n5601), 
        .Q(n8260) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n5114), .CLK(n5601), 
        .Q(n8259) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n5113), .CLK(n5601), 
        .Q(n8258) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n5113), .CLK(n5601), 
        .Q(n8257) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n5088), .CLK(n5614), 
        .Q(test_so91) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n5112), .CLK(n5602), 
        .Q(n8254) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n5112), .CLK(n5602), 
        .Q(n8253) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n5089), .CLK(n5613), 
        .Q(n8252) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n5111), .CLK(n5602), 
        .Q(n8251) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n5111), .CLK(n5602), 
        .Q(n8250) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n5111), .CLK(n5602), 
        .Q(n8249) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n5110), .CLK(n5603), 
        .Q(n8248) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n5109), .CLK(n5603), 
        .Q(n8247) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n5108), .CLK(n5604), 
        .Q(n8246) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n5108), .CLK(n5604), 
        .Q(WX11021) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n5107), .CLK(n5604), 
        .Q(WX11023) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n5107), .CLK(n5604), 
        .Q(WX11025) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n5106), .CLK(n5605), 
        .Q(WX11027) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n5105), .CLK(n5605), 
        .Q(WX11029) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n5105), .CLK(n5605), 
        .Q(WX11031) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n5104), .CLK(n5606), 
        .Q(WX11033) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n5103), .CLK(n5606), 
        .Q(test_so92) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n5102), .CLK(n5607), 
        .Q(WX11037) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n5102), .CLK(n5607), 
        .Q(WX11039) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n5101), .CLK(n5607), 
        .Q(WX11041) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n5101), .CLK(n5607), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n5100), .CLK(n5608), 
        .Q(WX11045) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n5099), .CLK(n5608), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n5099), .CLK(n5608), 
        .Q(WX11049) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n5098), .CLK(n5609), 
        .Q(WX11051) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n5097), .CLK(n5609), 
        .Q(WX11053), .QN(n4165) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n5114), .CLK(n5601), 
        .Q(WX11055), .QN(n4185) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n5114), .CLK(n5601), 
        .Q(WX11057), .QN(n4184) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n5114), .CLK(n5601), 
        .Q(WX11059), .QN(n4183) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n5113), .CLK(n5601), 
        .Q(WX11061), .QN(n4182) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n5113), .CLK(n5601), 
        .Q(WX11063), .QN(n4181) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n5113), .CLK(n5601), 
        .Q(WX11065) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n5113), .CLK(n5601), 
        .Q(WX11067), .QN(n4179) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n5112), .CLK(n5602), 
        .Q(test_so93), .QN(n9763) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n5088), .CLK(n5614), 
        .Q(WX11071), .QN(n4178) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n5111), .CLK(n5602), 
        .Q(WX11073), .QN(n9762) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n5111), .CLK(n5602), 
        .Q(WX11075), .QN(n4177) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n5110), .CLK(n5603), 
        .Q(WX11077) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n5110), .CLK(n5603), 
        .Q(WX11079), .QN(n4175) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n5109), .CLK(n5603), 
        .Q(WX11081), .QN(n4174) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n5109), .CLK(n5603), 
        .Q(WX11083), .QN(n4173) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n5108), .CLK(n5604), 
        .Q(WX11085), .QN(n9760) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n5107), .CLK(n5604), 
        .Q(WX11087), .QN(n9759) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n5107), .CLK(n5604), 
        .Q(WX11089), .QN(n9758) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n5106), .CLK(n5605), 
        .Q(WX11091), .QN(n9757) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n5105), .CLK(n5605), 
        .Q(WX11093), .QN(n9756) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n5105), .CLK(n5605), 
        .Q(WX11095), .QN(n9755) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n5104), .CLK(n5606), 
        .Q(WX11097), .QN(n9754) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n5103), .CLK(n5606), 
        .Q(WX11099), .QN(n9753) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n5103), .CLK(n5606), 
        .Q(WX11101), .QN(n9752) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n5102), .CLK(n5607), 
        .Q(test_so94) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n5101), .CLK(n5607), 
        .Q(WX11105), .QN(n9750) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n5101), .CLK(n5607), 
        .Q(WX11107), .QN(n9749) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n5100), .CLK(n5608), 
        .Q(WX11109), .QN(n9748) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n5099), .CLK(n5608), 
        .Q(WX11111), .QN(n9747) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n5099), .CLK(n5608), 
        .Q(WX11113), .QN(n9746) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n5098), .CLK(n5609), 
        .Q(WX11115), .QN(n9745) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n5097), .CLK(n5609), 
        .Q(WX11117) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n5097), .CLK(n5609), 
        .Q(WX11119) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n5097), .CLK(n5609), 
        .Q(WX11121) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n5096), .CLK(n5610), 
        .Q(WX11123) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n5096), .CLK(n5610), 
        .Q(WX11125) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n5096), .CLK(n5610), 
        .Q(WX11127) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n5095), .CLK(n5610), 
        .Q(WX11129), .QN(n4180) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n5095), .CLK(n5610), 
        .Q(WX11131) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n5112), .CLK(n5602), 
        .Q(WX11133), .QN(n9764) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n5112), .CLK(n5602), 
        .Q(WX11135) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n5112), .CLK(n5602), 
        .Q(test_so95), .QN(n9761) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n5111), .CLK(n5602), 
        .Q(WX11139) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n5110), .CLK(n5603), 
        .Q(WX11141), .QN(n4176) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n5110), .CLK(n5603), 
        .Q(WX11143) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n5109), .CLK(n5603), 
        .Q(WX11145) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n5109), .CLK(n5603), 
        .Q(WX11147) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n5108), .CLK(n5604), 
        .Q(WX11149), .QN(n4307) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n5107), .CLK(n5604), 
        .Q(WX11151), .QN(n4305) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n5106), .CLK(n5605), 
        .Q(WX11153), .QN(n4303) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n5106), .CLK(n5605), 
        .Q(WX11155), .QN(n4301) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155), .SE(n5105), .CLK(n5605), 
        .Q(WX11157), .QN(n4299) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(n5104), .CLK(n5606), 
        .Q(WX11159), .QN(n4297) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(n5104), .CLK(n5606), 
        .Q(WX11161), .QN(n4295) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(n5103), .CLK(n5606), 
        .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(n5103), .CLK(n5606), 
        .Q(WX11165), .QN(n4292) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(n5102), .CLK(n5607), 
        .Q(WX11167), .QN(n9751) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(n5101), .CLK(n5607), 
        .Q(WX11169), .QN(n4289) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(n5100), .CLK(n5608), 
        .Q(test_so96) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n5100), .CLK(n5608), 
        .Q(WX11173), .QN(n4286) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n5099), .CLK(n5608), 
        .Q(WX11175), .QN(n4284) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n5098), .CLK(n5609), 
        .Q(WX11177), .QN(n4282) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n5098), .CLK(n5609), 
        .Q(WX11179), .QN(n4280) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n5097), .CLK(n5609), 
        .Q(WX11181), .QN(n4542) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n5097), .CLK(n5609), 
        .Q(WX11183), .QN(n4543) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n5096), .CLK(n5610), 
        .Q(WX11185), .QN(n4544) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n5096), .CLK(n5610), 
        .Q(WX11187), .QN(n4545) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n5096), .CLK(n5610), 
        .Q(WX11189), .QN(n4546) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n5095), .CLK(n5610), 
        .Q(WX11191), .QN(n4547) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n5095), .CLK(n5610), 
        .Q(WX11193), .QN(n4548) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n5095), .CLK(n5610), 
        .Q(WX11195), .QN(n4549) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n5095), .CLK(n5610), 
        .Q(WX11197), .QN(n4550) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n5094), .CLK(n5611), 
        .Q(WX11199), .QN(n4551) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n5094), .CLK(n5611), 
        .Q(WX11201), .QN(n4552) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n5094), .CLK(n5611), 
        .Q(WX11203), .QN(n4553) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n5094), .CLK(n5611), 
        .Q(test_so97) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n5110), .CLK(n5603), 
        .Q(WX11207), .QN(n4554) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n5109), .CLK(n5603), 
        .Q(WX11209), .QN(n4555) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n5108), .CLK(n5604), 
        .Q(WX11211), .QN(n4513) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n5108), .CLK(n5604), 
        .Q(WX11213), .QN(n4556) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n5107), .CLK(n5604), 
        .Q(WX11215), .QN(n4557) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n5106), .CLK(n5605), 
        .Q(WX11217), .QN(n4558) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n5106), .CLK(n5605), 
        .Q(WX11219), .QN(n4559) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n5105), .CLK(n5605), 
        .Q(WX11221), .QN(n4514) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n5104), .CLK(n5606), 
        .Q(WX11223), .QN(n4560) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n5104), .CLK(n5606), 
        .Q(WX11225), .QN(n4561) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n5103), .CLK(n5606), 
        .Q(WX11227), .QN(n4562) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n5102), .CLK(n5607), 
        .Q(WX11229), .QN(n4563) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n5102), .CLK(n5607), 
        .Q(WX11231), .QN(n4564) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n5101), .CLK(n5607), 
        .Q(WX11233), .QN(n4565) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n5100), .CLK(n5608), 
        .Q(WX11235), .QN(n4515) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n5100), .CLK(n5608), 
        .Q(WX11237), .QN(n4566) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n5099), .CLK(n5608), 
        .Q(test_so98) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n5098), .CLK(n5609), 
        .Q(WX11241), .QN(n4567) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n5098), .CLK(n5609), 
        .Q(WX11243), .QN(n4534) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n5092), .CLK(n5612), 
        .Q(CRC_OUT_1_0) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n5092), .CLK(
        n5612), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n5092), .CLK(
        n5612), .Q(CRC_OUT_1_2) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n5092), .CLK(
        n5612), .Q(CRC_OUT_1_3) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n5092), .CLK(
        n5612), .Q(CRC_OUT_1_4) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n5092), .CLK(
        n5612), .Q(CRC_OUT_1_5) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_6) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_7) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_8) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_9) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_10) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n5091), .CLK(
        n5612), .Q(CRC_OUT_1_11) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n5090), .CLK(
        n5613), .Q(CRC_OUT_1_12) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n5090), .CLK(
        n5613), .Q(CRC_OUT_1_13) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n5090), .CLK(
        n5613), .Q(test_so99) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n5090), .CLK(n5613), .Q(CRC_OUT_1_15) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n5090), .CLK(
        n5613), .Q(CRC_OUT_1_16) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n5090), .CLK(
        n5613), .Q(CRC_OUT_1_17) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n5089), .CLK(
        n5613), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n5089), .CLK(
        n5613), .Q(CRC_OUT_1_19) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n5089), .CLK(
        n5613), .Q(CRC_OUT_1_20) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n5089), .CLK(
        n5613), .Q(CRC_OUT_1_21) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n5089), .CLK(
        n5613), .Q(CRC_OUT_1_22) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n5088), .CLK(
        n5614), .Q(CRC_OUT_1_23) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n5094), .CLK(
        n5611), .Q(CRC_OUT_1_24) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n5094), .CLK(
        n5611), .Q(CRC_OUT_1_25) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n5093), .CLK(
        n5611), .Q(CRC_OUT_1_26) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n5093), .CLK(
        n5611), .Q(CRC_OUT_1_27) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n5093), .CLK(
        n5611), .Q(CRC_OUT_1_28) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n5093), .CLK(
        n5611), .Q(CRC_OUT_1_29) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n5093), .CLK(
        n5611), .Q(CRC_OUT_1_30) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n5093), .CLK(
        n5611), .Q(test_so100) );
  NOR2X0 Trojan1 ( .IN1(WX3442), .IN2(WX5974), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(WX806), .IN2(WX782), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(WX11632), .IN2(n112), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(WX5964), .IN2(WX3324), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(WX8634), .IN2(WX3330), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n124), .IN2(n116), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(WX862), .IN2(WX7227), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(WX11616), .IN2(n485), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  INVX0 TrojanINVtest_se ( .INP(n5362), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  NBUFFX2 U4632 ( .INP(n4914), .Z(n4888) );
  NBUFFX2 U4633 ( .INP(n4914), .Z(n4889) );
  NBUFFX2 U4634 ( .INP(n4912), .Z(n4897) );
  NBUFFX2 U4635 ( .INP(n4912), .Z(n4899) );
  NBUFFX2 U4636 ( .INP(n4911), .Z(n4900) );
  NBUFFX2 U4637 ( .INP(n4911), .Z(n4901) );
  NBUFFX2 U4638 ( .INP(n4911), .Z(n4902) );
  NBUFFX2 U4639 ( .INP(n4911), .Z(n4903) );
  NBUFFX2 U4640 ( .INP(n4911), .Z(n4904) );
  NBUFFX2 U4641 ( .INP(n4910), .Z(n4908) );
  NBUFFX2 U4642 ( .INP(n4913), .Z(n4890) );
  NBUFFX2 U4643 ( .INP(n4913), .Z(n4891) );
  NBUFFX2 U4644 ( .INP(n4913), .Z(n4892) );
  NBUFFX2 U4645 ( .INP(n4912), .Z(n4898) );
  NBUFFX2 U4646 ( .INP(n4913), .Z(n4893) );
  NBUFFX2 U4647 ( .INP(n4913), .Z(n4894) );
  NBUFFX2 U4648 ( .INP(n4912), .Z(n4895) );
  NBUFFX2 U4649 ( .INP(n4912), .Z(n4896) );
  NBUFFX2 U4650 ( .INP(n4910), .Z(n4905) );
  NBUFFX2 U4651 ( .INP(n4910), .Z(n4906) );
  NBUFFX2 U4652 ( .INP(n4910), .Z(n4907) );
  NBUFFX2 U4653 ( .INP(n4914), .Z(n4887) );
  NBUFFX2 U4654 ( .INP(n5714), .Z(n5545) );
  NBUFFX2 U4655 ( .INP(n5714), .Z(n5543) );
  NBUFFX2 U4656 ( .INP(n5714), .Z(n5544) );
  NBUFFX2 U4657 ( .INP(n5714), .Z(n5542) );
  NBUFFX2 U4658 ( .INP(n5700), .Z(n5612) );
  NBUFFX2 U4659 ( .INP(n5700), .Z(n5611) );
  NBUFFX2 U4660 ( .INP(n5701), .Z(n5610) );
  NBUFFX2 U4661 ( .INP(n5701), .Z(n5609) );
  NBUFFX2 U4662 ( .INP(n5701), .Z(n5608) );
  NBUFFX2 U4663 ( .INP(n5701), .Z(n5607) );
  NBUFFX2 U4664 ( .INP(n5701), .Z(n5606) );
  NBUFFX2 U4665 ( .INP(n5702), .Z(n5605) );
  NBUFFX2 U4666 ( .INP(n5702), .Z(n5604) );
  NBUFFX2 U4667 ( .INP(n5702), .Z(n5603) );
  NBUFFX2 U4668 ( .INP(n5700), .Z(n5613) );
  NBUFFX2 U4669 ( .INP(n5702), .Z(n5602) );
  NBUFFX2 U4670 ( .INP(n5702), .Z(n5601) );
  NBUFFX2 U4671 ( .INP(n5703), .Z(n5599) );
  NBUFFX2 U4672 ( .INP(n5703), .Z(n5600) );
  NBUFFX2 U4673 ( .INP(n5703), .Z(n5598) );
  NBUFFX2 U4674 ( .INP(n5700), .Z(n5614) );
  NBUFFX2 U4675 ( .INP(n5703), .Z(n5597) );
  NBUFFX2 U4676 ( .INP(n5703), .Z(n5596) );
  NBUFFX2 U4677 ( .INP(n5704), .Z(n5595) );
  NBUFFX2 U4678 ( .INP(n5704), .Z(n5594) );
  NBUFFX2 U4679 ( .INP(n5704), .Z(n5593) );
  NBUFFX2 U4680 ( .INP(n5704), .Z(n5592) );
  NBUFFX2 U4681 ( .INP(n5704), .Z(n5591) );
  NBUFFX2 U4682 ( .INP(n5705), .Z(n5590) );
  NBUFFX2 U4683 ( .INP(n5705), .Z(n5589) );
  NBUFFX2 U4684 ( .INP(n5700), .Z(n5615) );
  NBUFFX2 U4685 ( .INP(n5705), .Z(n5588) );
  NBUFFX2 U4686 ( .INP(n5706), .Z(n5585) );
  NBUFFX2 U4687 ( .INP(n5706), .Z(n5584) );
  NBUFFX2 U4688 ( .INP(n5706), .Z(n5583) );
  NBUFFX2 U4689 ( .INP(n5699), .Z(n5616) );
  NBUFFX2 U4690 ( .INP(n5706), .Z(n5582) );
  NBUFFX2 U4691 ( .INP(n5706), .Z(n5581) );
  NBUFFX2 U4692 ( .INP(n5705), .Z(n5587) );
  NBUFFX2 U4693 ( .INP(n5708), .Z(n5575) );
  NBUFFX2 U4694 ( .INP(n5708), .Z(n5574) );
  NBUFFX2 U4695 ( .INP(n5708), .Z(n5573) );
  NBUFFX2 U4696 ( .INP(n5708), .Z(n5572) );
  NBUFFX2 U4697 ( .INP(n5707), .Z(n5580) );
  NBUFFX2 U4698 ( .INP(n5707), .Z(n5579) );
  NBUFFX2 U4699 ( .INP(n5707), .Z(n5578) );
  NBUFFX2 U4700 ( .INP(n5707), .Z(n5577) );
  NBUFFX2 U4701 ( .INP(n5705), .Z(n5586) );
  NBUFFX2 U4702 ( .INP(n5707), .Z(n5576) );
  NBUFFX2 U4703 ( .INP(n5708), .Z(n5571) );
  NBUFFX2 U4704 ( .INP(n5709), .Z(n5570) );
  NBUFFX2 U4705 ( .INP(n5688), .Z(n5671) );
  NBUFFX2 U4706 ( .INP(n5689), .Z(n5670) );
  NBUFFX2 U4707 ( .INP(n5689), .Z(n5669) );
  NBUFFX2 U4708 ( .INP(n5689), .Z(n5668) );
  NBUFFX2 U4709 ( .INP(n5689), .Z(n5667) );
  NBUFFX2 U4710 ( .INP(n5689), .Z(n5666) );
  NBUFFX2 U4711 ( .INP(n5690), .Z(n5665) );
  NBUFFX2 U4712 ( .INP(n5690), .Z(n5664) );
  NBUFFX2 U4713 ( .INP(n5690), .Z(n5663) );
  NBUFFX2 U4714 ( .INP(n5690), .Z(n5662) );
  NBUFFX2 U4715 ( .INP(n5690), .Z(n5661) );
  NBUFFX2 U4716 ( .INP(n5691), .Z(n5660) );
  NBUFFX2 U4717 ( .INP(n5691), .Z(n5657) );
  NBUFFX2 U4718 ( .INP(n5691), .Z(n5658) );
  NBUFFX2 U4719 ( .INP(n5691), .Z(n5659) );
  NBUFFX2 U4720 ( .INP(n5691), .Z(n5656) );
  NBUFFX2 U4721 ( .INP(n5688), .Z(n5672) );
  NBUFFX2 U4722 ( .INP(n5692), .Z(n5655) );
  NBUFFX2 U4723 ( .INP(n5692), .Z(n5654) );
  NBUFFX2 U4724 ( .INP(n5692), .Z(n5653) );
  NBUFFX2 U4725 ( .INP(n5692), .Z(n5652) );
  NBUFFX2 U4726 ( .INP(n5692), .Z(n5651) );
  NBUFFX2 U4727 ( .INP(n5693), .Z(n5650) );
  NBUFFX2 U4728 ( .INP(n5693), .Z(n5649) );
  NBUFFX2 U4729 ( .INP(n5693), .Z(n5648) );
  NBUFFX2 U4730 ( .INP(n5688), .Z(n5673) );
  NBUFFX2 U4731 ( .INP(n5693), .Z(n5647) );
  NBUFFX2 U4732 ( .INP(n5693), .Z(n5646) );
  NBUFFX2 U4733 ( .INP(n5694), .Z(n5643) );
  NBUFFX2 U4734 ( .INP(n5694), .Z(n5644) );
  NBUFFX2 U4735 ( .INP(n5694), .Z(n5645) );
  NBUFFX2 U4736 ( .INP(n5687), .Z(n5676) );
  NBUFFX2 U4737 ( .INP(n5688), .Z(n5675) );
  NBUFFX2 U4738 ( .INP(n5694), .Z(n5642) );
  NBUFFX2 U4739 ( .INP(n5694), .Z(n5641) );
  NBUFFX2 U4740 ( .INP(n5695), .Z(n5640) );
  NBUFFX2 U4741 ( .INP(n5695), .Z(n5639) );
  NBUFFX2 U4742 ( .INP(n5695), .Z(n5638) );
  NBUFFX2 U4743 ( .INP(n5695), .Z(n5637) );
  NBUFFX2 U4744 ( .INP(n5695), .Z(n5636) );
  NBUFFX2 U4745 ( .INP(n5696), .Z(n5635) );
  NBUFFX2 U4746 ( .INP(n5696), .Z(n5633) );
  NBUFFX2 U4747 ( .INP(n5688), .Z(n5674) );
  NBUFFX2 U4748 ( .INP(n5697), .Z(n5630) );
  NBUFFX2 U4749 ( .INP(n5696), .Z(n5631) );
  NBUFFX2 U4750 ( .INP(n5697), .Z(n5629) );
  NBUFFX2 U4751 ( .INP(n5697), .Z(n5628) );
  NBUFFX2 U4752 ( .INP(n5697), .Z(n5627) );
  NBUFFX2 U4753 ( .INP(n5697), .Z(n5626) );
  NBUFFX2 U4754 ( .INP(n5698), .Z(n5625) );
  NBUFFX2 U4755 ( .INP(n5699), .Z(n5620) );
  NBUFFX2 U4756 ( .INP(n5699), .Z(n5619) );
  NBUFFX2 U4757 ( .INP(n5699), .Z(n5618) );
  NBUFFX2 U4758 ( .INP(n5699), .Z(n5617) );
  NBUFFX2 U4759 ( .INP(n5698), .Z(n5624) );
  NBUFFX2 U4760 ( .INP(n5696), .Z(n5634) );
  NBUFFX2 U4761 ( .INP(n5698), .Z(n5623) );
  NBUFFX2 U4762 ( .INP(n5698), .Z(n5622) );
  NBUFFX2 U4763 ( .INP(n5687), .Z(n5677) );
  NBUFFX2 U4764 ( .INP(n5696), .Z(n5632) );
  NBUFFX2 U4765 ( .INP(n5698), .Z(n5621) );
  NBUFFX2 U4766 ( .INP(n5709), .Z(n5567) );
  NBUFFX2 U4767 ( .INP(n5709), .Z(n5568) );
  NBUFFX2 U4768 ( .INP(n5709), .Z(n5569) );
  NBUFFX2 U4769 ( .INP(n5709), .Z(n5566) );
  NBUFFX2 U4770 ( .INP(n5687), .Z(n5679) );
  NBUFFX2 U4771 ( .INP(n5687), .Z(n5678) );
  NBUFFX2 U4772 ( .INP(n5710), .Z(n5565) );
  NBUFFX2 U4773 ( .INP(n5686), .Z(n5683) );
  NBUFFX2 U4774 ( .INP(n5710), .Z(n5564) );
  NBUFFX2 U4775 ( .INP(n5686), .Z(n5682) );
  NBUFFX2 U4776 ( .INP(n5686), .Z(n5681) );
  NBUFFX2 U4777 ( .INP(n5710), .Z(n5563) );
  NBUFFX2 U4778 ( .INP(n5710), .Z(n5562) );
  NBUFFX2 U4779 ( .INP(n5710), .Z(n5561) );
  NBUFFX2 U4780 ( .INP(n5687), .Z(n5680) );
  NBUFFX2 U4781 ( .INP(n5711), .Z(n5560) );
  NBUFFX2 U4782 ( .INP(n5711), .Z(n5559) );
  NBUFFX2 U4783 ( .INP(n5711), .Z(n5557) );
  NBUFFX2 U4784 ( .INP(n5711), .Z(n5558) );
  NBUFFX2 U4785 ( .INP(n5711), .Z(n5556) );
  NBUFFX2 U4786 ( .INP(n5686), .Z(n5684) );
  NBUFFX2 U4787 ( .INP(n5712), .Z(n5555) );
  NBUFFX2 U4788 ( .INP(n5712), .Z(n5554) );
  NBUFFX2 U4789 ( .INP(n5712), .Z(n5553) );
  NBUFFX2 U4790 ( .INP(n5712), .Z(n5552) );
  NBUFFX2 U4791 ( .INP(n5712), .Z(n5551) );
  NBUFFX2 U4792 ( .INP(n5713), .Z(n5550) );
  NBUFFX2 U4793 ( .INP(n5686), .Z(n5685) );
  NBUFFX2 U4794 ( .INP(n5713), .Z(n5549) );
  NBUFFX2 U4795 ( .INP(n5713), .Z(n5548) );
  NBUFFX2 U4796 ( .INP(n5713), .Z(n5547) );
  NBUFFX2 U4797 ( .INP(n5713), .Z(n5546) );
  NBUFFX2 U4798 ( .INP(n4910), .Z(n4909) );
  NBUFFX2 U4799 ( .INP(n4943), .Z(n4924) );
  NBUFFX2 U4800 ( .INP(n4829), .Z(n4838) );
  NBUFFX2 U4801 ( .INP(n4832), .Z(n4854) );
  NBUFFX2 U4802 ( .INP(n4832), .Z(n4853) );
  NBUFFX2 U4803 ( .INP(n4941), .Z(n4931) );
  NBUFFX2 U4804 ( .INP(n4941), .Z(n4932) );
  NBUFFX2 U4805 ( .INP(n4941), .Z(n4933) );
  NBUFFX2 U4806 ( .INP(n4941), .Z(n4934) );
  NBUFFX2 U4807 ( .INP(n4940), .Z(n4938) );
  NBUFFX2 U4808 ( .INP(n4942), .Z(n4926) );
  NBUFFX2 U4809 ( .INP(n4942), .Z(n4927) );
  NBUFFX2 U4810 ( .INP(n4942), .Z(n4928) );
  NBUFFX2 U4811 ( .INP(n4942), .Z(n4925) );
  NBUFFX2 U4812 ( .INP(n4941), .Z(n4930) );
  NBUFFX2 U4813 ( .INP(n4942), .Z(n4929) );
  NBUFFX2 U4814 ( .INP(n4940), .Z(n4935) );
  NBUFFX2 U4815 ( .INP(n4940), .Z(n4936) );
  NBUFFX2 U4816 ( .INP(n4940), .Z(n4937) );
  NBUFFX2 U4817 ( .INP(n4830), .Z(n4846) );
  NBUFFX2 U4818 ( .INP(n4830), .Z(n4845) );
  NBUFFX2 U4819 ( .INP(n4830), .Z(n4844) );
  NBUFFX2 U4820 ( .INP(n4830), .Z(n4843) );
  NBUFFX2 U4821 ( .INP(n4829), .Z(n4842) );
  NBUFFX2 U4822 ( .INP(n4831), .Z(n4852) );
  NBUFFX2 U4823 ( .INP(n4831), .Z(n4851) );
  NBUFFX2 U4824 ( .INP(n4831), .Z(n4850) );
  NBUFFX2 U4825 ( .INP(n4831), .Z(n4849) );
  NBUFFX2 U4826 ( .INP(n4831), .Z(n4848) );
  NBUFFX2 U4827 ( .INP(n4830), .Z(n4847) );
  NBUFFX2 U4828 ( .INP(n4829), .Z(n4839) );
  NBUFFX2 U4829 ( .INP(n4829), .Z(n4840) );
  NBUFFX2 U4830 ( .INP(n4829), .Z(n4841) );
  NBUFFX2 U4831 ( .INP(n4944), .Z(n4917) );
  NBUFFX2 U4832 ( .INP(n4944), .Z(n4919) );
  NBUFFX2 U4833 ( .INP(n4944), .Z(n4918) );
  NBUFFX2 U4834 ( .INP(n4943), .Z(n4923) );
  NBUFFX2 U4835 ( .INP(n4943), .Z(n4922) );
  NBUFFX2 U4836 ( .INP(n4943), .Z(n4920) );
  NBUFFX2 U4837 ( .INP(n4943), .Z(n4921) );
  NBUFFX2 U4838 ( .INP(n4828), .Z(n4837) );
  NBUFFX2 U4839 ( .INP(n4828), .Z(n4836) );
  NBUFFX2 U4840 ( .INP(n4828), .Z(n4835) );
  NBUFFX2 U4841 ( .INP(n4828), .Z(n4834) );
  NBUFFX2 U4842 ( .INP(n4828), .Z(n4833) );
  NBUFFX2 U4843 ( .INP(n4940), .Z(n4939) );
  NBUFFX2 U4844 ( .INP(n4832), .Z(n4855) );
  NBUFFX2 U4845 ( .INP(n4860), .Z(n4883) );
  NBUFFX2 U4846 ( .INP(n4860), .Z(n4882) );
  NBUFFX2 U4847 ( .INP(n4860), .Z(n4881) );
  NBUFFX2 U4848 ( .INP(n4856), .Z(n4862) );
  NBUFFX2 U4849 ( .INP(n4856), .Z(n4861) );
  NBUFFX2 U4850 ( .INP(n4859), .Z(n4880) );
  NBUFFX2 U4851 ( .INP(n4859), .Z(n4879) );
  NBUFFX2 U4852 ( .INP(n4859), .Z(n4878) );
  NBUFFX2 U4853 ( .INP(n4859), .Z(n4877) );
  NBUFFX2 U4854 ( .INP(n4858), .Z(n4872) );
  NBUFFX2 U4855 ( .INP(n4858), .Z(n4871) );
  NBUFFX2 U4856 ( .INP(n4857), .Z(n4870) );
  NBUFFX2 U4857 ( .INP(n4857), .Z(n4869) );
  NBUFFX2 U4858 ( .INP(n4857), .Z(n4868) );
  NBUFFX2 U4859 ( .INP(n4857), .Z(n4867) );
  NBUFFX2 U4860 ( .INP(n4857), .Z(n4866) );
  NBUFFX2 U4861 ( .INP(n4856), .Z(n4865) );
  NBUFFX2 U4862 ( .INP(n4856), .Z(n4864) );
  NBUFFX2 U4863 ( .INP(n4856), .Z(n4863) );
  NBUFFX2 U4864 ( .INP(n4859), .Z(n4876) );
  NBUFFX2 U4865 ( .INP(n4858), .Z(n4875) );
  NBUFFX2 U4866 ( .INP(n4858), .Z(n4874) );
  NBUFFX2 U4867 ( .INP(n4858), .Z(n4873) );
  NBUFFX2 U4868 ( .INP(n4860), .Z(n4884) );
  NBUFFX2 U4869 ( .INP(n5748), .Z(n4828) );
  NBUFFX2 U4870 ( .INP(n5748), .Z(n4829) );
  NBUFFX2 U4871 ( .INP(n5748), .Z(n4830) );
  NBUFFX2 U4872 ( .INP(n5748), .Z(n4831) );
  NBUFFX2 U4873 ( .INP(n5748), .Z(n4832) );
  NBUFFX2 U4874 ( .INP(n2148), .Z(n4856) );
  NBUFFX2 U4875 ( .INP(n2148), .Z(n4857) );
  NBUFFX2 U4876 ( .INP(n2148), .Z(n4858) );
  NBUFFX2 U4877 ( .INP(n2148), .Z(n4859) );
  NBUFFX2 U4878 ( .INP(n2148), .Z(n4860) );
  NBUFFX2 U4879 ( .INP(n2152), .Z(n4885) );
  NBUFFX2 U4880 ( .INP(n2152), .Z(n4886) );
  NBUFFX2 U4881 ( .INP(n4885), .Z(n4910) );
  NBUFFX2 U4882 ( .INP(n4885), .Z(n4911) );
  NBUFFX2 U4883 ( .INP(n4885), .Z(n4912) );
  NBUFFX2 U4884 ( .INP(n4886), .Z(n4913) );
  NBUFFX2 U4885 ( .INP(n4886), .Z(n4914) );
  NBUFFX2 U4886 ( .INP(n2153), .Z(n4915) );
  NBUFFX2 U4887 ( .INP(n2153), .Z(n4916) );
  NBUFFX2 U4888 ( .INP(n4915), .Z(n4940) );
  NBUFFX2 U4889 ( .INP(n4915), .Z(n4941) );
  NBUFFX2 U4890 ( .INP(n4915), .Z(n4942) );
  NBUFFX2 U4891 ( .INP(n4916), .Z(n4943) );
  NBUFFX2 U4892 ( .INP(n4916), .Z(n4944) );
  NBUFFX2 U4893 ( .INP(n5329), .Z(n4945) );
  NBUFFX2 U4894 ( .INP(n5328), .Z(n4946) );
  NBUFFX2 U4895 ( .INP(n5328), .Z(n4947) );
  NBUFFX2 U4896 ( .INP(n5328), .Z(n4948) );
  NBUFFX2 U4897 ( .INP(n5327), .Z(n4949) );
  NBUFFX2 U4898 ( .INP(n5327), .Z(n4950) );
  NBUFFX2 U4899 ( .INP(n5327), .Z(n4951) );
  NBUFFX2 U4900 ( .INP(n5326), .Z(n4952) );
  NBUFFX2 U4901 ( .INP(n5326), .Z(n4953) );
  NBUFFX2 U4902 ( .INP(n5326), .Z(n4954) );
  NBUFFX2 U4903 ( .INP(n5325), .Z(n4955) );
  NBUFFX2 U4904 ( .INP(n5325), .Z(n4956) );
  NBUFFX2 U4905 ( .INP(n5325), .Z(n4957) );
  NBUFFX2 U4906 ( .INP(n5324), .Z(n4958) );
  NBUFFX2 U4907 ( .INP(n5324), .Z(n4959) );
  NBUFFX2 U4908 ( .INP(n5324), .Z(n4960) );
  NBUFFX2 U4909 ( .INP(n5323), .Z(n4961) );
  NBUFFX2 U4910 ( .INP(n5323), .Z(n4962) );
  NBUFFX2 U4911 ( .INP(n5323), .Z(n4963) );
  NBUFFX2 U4912 ( .INP(n5322), .Z(n4964) );
  NBUFFX2 U4913 ( .INP(n5322), .Z(n4965) );
  NBUFFX2 U4914 ( .INP(n5322), .Z(n4966) );
  NBUFFX2 U4915 ( .INP(n5321), .Z(n4967) );
  NBUFFX2 U4916 ( .INP(n5321), .Z(n4968) );
  NBUFFX2 U4917 ( .INP(n5321), .Z(n4969) );
  NBUFFX2 U4918 ( .INP(n5320), .Z(n4970) );
  NBUFFX2 U4919 ( .INP(n5320), .Z(n4971) );
  NBUFFX2 U4920 ( .INP(n5320), .Z(n4972) );
  NBUFFX2 U4921 ( .INP(n5319), .Z(n4973) );
  NBUFFX2 U4922 ( .INP(n5319), .Z(n4974) );
  NBUFFX2 U4923 ( .INP(n5319), .Z(n4975) );
  NBUFFX2 U4924 ( .INP(n5318), .Z(n4976) );
  NBUFFX2 U4925 ( .INP(n5318), .Z(n4977) );
  NBUFFX2 U4926 ( .INP(n5318), .Z(n4978) );
  NBUFFX2 U4927 ( .INP(n5317), .Z(n4979) );
  NBUFFX2 U4928 ( .INP(n5317), .Z(n4980) );
  NBUFFX2 U4929 ( .INP(n5317), .Z(n4981) );
  NBUFFX2 U4930 ( .INP(n5316), .Z(n4982) );
  NBUFFX2 U4931 ( .INP(n5316), .Z(n4983) );
  NBUFFX2 U4932 ( .INP(n5316), .Z(n4984) );
  NBUFFX2 U4933 ( .INP(n5315), .Z(n4985) );
  NBUFFX2 U4934 ( .INP(n5315), .Z(n4986) );
  NBUFFX2 U4935 ( .INP(n5315), .Z(n4987) );
  NBUFFX2 U4936 ( .INP(n5314), .Z(n4988) );
  NBUFFX2 U4937 ( .INP(n5314), .Z(n4989) );
  NBUFFX2 U4938 ( .INP(n5314), .Z(n4990) );
  NBUFFX2 U4939 ( .INP(n5313), .Z(n4991) );
  NBUFFX2 U4940 ( .INP(n5313), .Z(n4992) );
  NBUFFX2 U4941 ( .INP(n5313), .Z(n4993) );
  NBUFFX2 U4942 ( .INP(n5312), .Z(n4994) );
  NBUFFX2 U4943 ( .INP(n5312), .Z(n4995) );
  NBUFFX2 U4944 ( .INP(n5312), .Z(n4996) );
  NBUFFX2 U4945 ( .INP(n5311), .Z(n4997) );
  NBUFFX2 U4946 ( .INP(n5311), .Z(n4998) );
  NBUFFX2 U4947 ( .INP(n5311), .Z(n4999) );
  NBUFFX2 U4948 ( .INP(n5310), .Z(n5000) );
  NBUFFX2 U4949 ( .INP(n5310), .Z(n5001) );
  NBUFFX2 U4950 ( .INP(n5310), .Z(n5002) );
  NBUFFX2 U4951 ( .INP(n5309), .Z(n5003) );
  NBUFFX2 U4952 ( .INP(n5309), .Z(n5004) );
  NBUFFX2 U4953 ( .INP(n5309), .Z(n5005) );
  NBUFFX2 U4954 ( .INP(n5308), .Z(n5006) );
  NBUFFX2 U4955 ( .INP(n5308), .Z(n5007) );
  NBUFFX2 U4956 ( .INP(n5308), .Z(n5008) );
  NBUFFX2 U4957 ( .INP(n5307), .Z(n5009) );
  NBUFFX2 U4958 ( .INP(n5307), .Z(n5010) );
  NBUFFX2 U4959 ( .INP(n5307), .Z(n5011) );
  NBUFFX2 U4960 ( .INP(n5306), .Z(n5012) );
  NBUFFX2 U4961 ( .INP(n5306), .Z(n5013) );
  NBUFFX2 U4962 ( .INP(n5306), .Z(n5014) );
  NBUFFX2 U4963 ( .INP(n5305), .Z(n5015) );
  NBUFFX2 U4964 ( .INP(n5305), .Z(n5016) );
  NBUFFX2 U4965 ( .INP(n5305), .Z(n5017) );
  NBUFFX2 U4966 ( .INP(n5304), .Z(n5018) );
  NBUFFX2 U4967 ( .INP(n5304), .Z(n5019) );
  NBUFFX2 U4968 ( .INP(n5304), .Z(n5020) );
  NBUFFX2 U4969 ( .INP(n5303), .Z(n5021) );
  NBUFFX2 U4970 ( .INP(n5303), .Z(n5022) );
  NBUFFX2 U4971 ( .INP(n5303), .Z(n5023) );
  NBUFFX2 U4972 ( .INP(n5302), .Z(n5024) );
  NBUFFX2 U4973 ( .INP(n5302), .Z(n5025) );
  NBUFFX2 U4974 ( .INP(n5302), .Z(n5026) );
  NBUFFX2 U4975 ( .INP(n5301), .Z(n5027) );
  NBUFFX2 U4976 ( .INP(n5301), .Z(n5028) );
  NBUFFX2 U4977 ( .INP(n5301), .Z(n5029) );
  NBUFFX2 U4978 ( .INP(n5300), .Z(n5030) );
  NBUFFX2 U4979 ( .INP(n5300), .Z(n5031) );
  NBUFFX2 U4980 ( .INP(n5300), .Z(n5032) );
  NBUFFX2 U4981 ( .INP(n5299), .Z(n5033) );
  NBUFFX2 U4982 ( .INP(n5299), .Z(n5034) );
  NBUFFX2 U4983 ( .INP(n5299), .Z(n5035) );
  NBUFFX2 U4984 ( .INP(n5298), .Z(n5036) );
  NBUFFX2 U4985 ( .INP(n5298), .Z(n5037) );
  NBUFFX2 U4986 ( .INP(n5298), .Z(n5038) );
  NBUFFX2 U4987 ( .INP(n5297), .Z(n5039) );
  NBUFFX2 U4988 ( .INP(n5297), .Z(n5040) );
  NBUFFX2 U4989 ( .INP(n5297), .Z(n5041) );
  NBUFFX2 U4990 ( .INP(n5296), .Z(n5042) );
  NBUFFX2 U4991 ( .INP(n5296), .Z(n5043) );
  NBUFFX2 U4992 ( .INP(n5296), .Z(n5044) );
  NBUFFX2 U4993 ( .INP(n5295), .Z(n5045) );
  NBUFFX2 U4994 ( .INP(n5295), .Z(n5046) );
  NBUFFX2 U4995 ( .INP(n5295), .Z(n5047) );
  NBUFFX2 U4996 ( .INP(n5294), .Z(n5048) );
  NBUFFX2 U4997 ( .INP(n5294), .Z(n5049) );
  NBUFFX2 U4998 ( .INP(n5294), .Z(n5050) );
  NBUFFX2 U4999 ( .INP(n5293), .Z(n5051) );
  NBUFFX2 U5000 ( .INP(n5293), .Z(n5052) );
  NBUFFX2 U5001 ( .INP(n5293), .Z(n5053) );
  NBUFFX2 U5002 ( .INP(n5292), .Z(n5054) );
  NBUFFX2 U5003 ( .INP(n5292), .Z(n5055) );
  NBUFFX2 U5004 ( .INP(n5292), .Z(n5056) );
  NBUFFX2 U5005 ( .INP(n5291), .Z(n5057) );
  NBUFFX2 U5006 ( .INP(n5291), .Z(n5058) );
  NBUFFX2 U5007 ( .INP(n5291), .Z(n5059) );
  NBUFFX2 U5008 ( .INP(n5290), .Z(n5060) );
  NBUFFX2 U5009 ( .INP(n5290), .Z(n5061) );
  NBUFFX2 U5010 ( .INP(n5290), .Z(n5062) );
  NBUFFX2 U5011 ( .INP(n5289), .Z(n5063) );
  NBUFFX2 U5012 ( .INP(n5289), .Z(n5064) );
  NBUFFX2 U5013 ( .INP(n5289), .Z(n5065) );
  NBUFFX2 U5014 ( .INP(n5288), .Z(n5066) );
  NBUFFX2 U5015 ( .INP(n5288), .Z(n5067) );
  NBUFFX2 U5016 ( .INP(n5288), .Z(n5068) );
  NBUFFX2 U5017 ( .INP(n5287), .Z(n5069) );
  NBUFFX2 U5018 ( .INP(n5287), .Z(n5070) );
  NBUFFX2 U5019 ( .INP(n5287), .Z(n5071) );
  NBUFFX2 U5020 ( .INP(n5286), .Z(n5072) );
  NBUFFX2 U5021 ( .INP(n5286), .Z(n5073) );
  NBUFFX2 U5022 ( .INP(n5286), .Z(n5074) );
  NBUFFX2 U5023 ( .INP(n5285), .Z(n5075) );
  NBUFFX2 U5024 ( .INP(n5285), .Z(n5076) );
  NBUFFX2 U5025 ( .INP(n5285), .Z(n5077) );
  NBUFFX2 U5026 ( .INP(n5284), .Z(n5078) );
  NBUFFX2 U5027 ( .INP(n5284), .Z(n5079) );
  NBUFFX2 U5028 ( .INP(n5284), .Z(n5080) );
  NBUFFX2 U5029 ( .INP(n5283), .Z(n5081) );
  NBUFFX2 U5030 ( .INP(n5283), .Z(n5082) );
  NBUFFX2 U5031 ( .INP(n5283), .Z(n5083) );
  NBUFFX2 U5032 ( .INP(n5282), .Z(n5084) );
  NBUFFX2 U5033 ( .INP(n5282), .Z(n5085) );
  NBUFFX2 U5034 ( .INP(n5282), .Z(n5086) );
  NBUFFX2 U5035 ( .INP(n5281), .Z(n5087) );
  NBUFFX2 U5036 ( .INP(n5281), .Z(n5088) );
  NBUFFX2 U5037 ( .INP(n5281), .Z(n5089) );
  NBUFFX2 U5038 ( .INP(n5280), .Z(n5090) );
  NBUFFX2 U5039 ( .INP(n5280), .Z(n5091) );
  NBUFFX2 U5040 ( .INP(n5280), .Z(n5092) );
  NBUFFX2 U5041 ( .INP(n5279), .Z(n5093) );
  NBUFFX2 U5042 ( .INP(n5279), .Z(n5094) );
  NBUFFX2 U5043 ( .INP(n5279), .Z(n5095) );
  NBUFFX2 U5044 ( .INP(n5278), .Z(n5096) );
  NBUFFX2 U5045 ( .INP(n5278), .Z(n5097) );
  NBUFFX2 U5046 ( .INP(n5278), .Z(n5098) );
  NBUFFX2 U5047 ( .INP(n5277), .Z(n5099) );
  NBUFFX2 U5048 ( .INP(n5277), .Z(n5100) );
  NBUFFX2 U5049 ( .INP(n5277), .Z(n5101) );
  NBUFFX2 U5050 ( .INP(n5276), .Z(n5102) );
  NBUFFX2 U5051 ( .INP(n5276), .Z(n5103) );
  NBUFFX2 U5052 ( .INP(n5276), .Z(n5104) );
  NBUFFX2 U5053 ( .INP(n5275), .Z(n5105) );
  NBUFFX2 U5054 ( .INP(n5275), .Z(n5106) );
  NBUFFX2 U5055 ( .INP(n5275), .Z(n5107) );
  NBUFFX2 U5056 ( .INP(n5274), .Z(n5108) );
  NBUFFX2 U5057 ( .INP(n5274), .Z(n5109) );
  NBUFFX2 U5058 ( .INP(n5274), .Z(n5110) );
  NBUFFX2 U5059 ( .INP(n5273), .Z(n5111) );
  NBUFFX2 U5060 ( .INP(n5273), .Z(n5112) );
  NBUFFX2 U5061 ( .INP(n5273), .Z(n5113) );
  NBUFFX2 U5062 ( .INP(n5272), .Z(n5114) );
  NBUFFX2 U5063 ( .INP(n5272), .Z(n5115) );
  NBUFFX2 U5064 ( .INP(n5272), .Z(n5116) );
  NBUFFX2 U5065 ( .INP(n5271), .Z(n5117) );
  NBUFFX2 U5066 ( .INP(n5271), .Z(n5118) );
  NBUFFX2 U5067 ( .INP(n5271), .Z(n5119) );
  NBUFFX2 U5068 ( .INP(n5270), .Z(n5120) );
  NBUFFX2 U5069 ( .INP(n5270), .Z(n5121) );
  NBUFFX2 U5070 ( .INP(n5270), .Z(n5122) );
  NBUFFX2 U5071 ( .INP(n5269), .Z(n5123) );
  NBUFFX2 U5072 ( .INP(n5269), .Z(n5124) );
  NBUFFX2 U5073 ( .INP(n5269), .Z(n5125) );
  NBUFFX2 U5074 ( .INP(n5268), .Z(n5126) );
  NBUFFX2 U5075 ( .INP(n5268), .Z(n5127) );
  NBUFFX2 U5076 ( .INP(n5268), .Z(n5128) );
  NBUFFX2 U5077 ( .INP(n5267), .Z(n5129) );
  NBUFFX2 U5078 ( .INP(n5267), .Z(n5130) );
  NBUFFX2 U5079 ( .INP(n5267), .Z(n5131) );
  NBUFFX2 U5080 ( .INP(n5266), .Z(n5132) );
  NBUFFX2 U5081 ( .INP(n5266), .Z(n5133) );
  NBUFFX2 U5082 ( .INP(n5266), .Z(n5134) );
  NBUFFX2 U5083 ( .INP(n5265), .Z(n5135) );
  NBUFFX2 U5084 ( .INP(n5265), .Z(n5136) );
  NBUFFX2 U5085 ( .INP(n5265), .Z(n5137) );
  NBUFFX2 U5086 ( .INP(n5264), .Z(n5138) );
  NBUFFX2 U5087 ( .INP(n5264), .Z(n5139) );
  NBUFFX2 U5088 ( .INP(n5264), .Z(n5140) );
  NBUFFX2 U5089 ( .INP(n5263), .Z(n5141) );
  NBUFFX2 U5090 ( .INP(n5263), .Z(n5142) );
  NBUFFX2 U5091 ( .INP(n5263), .Z(n5143) );
  NBUFFX2 U5092 ( .INP(n5262), .Z(n5144) );
  NBUFFX2 U5093 ( .INP(n5262), .Z(n5145) );
  NBUFFX2 U5094 ( .INP(n5262), .Z(n5146) );
  NBUFFX2 U5095 ( .INP(n5261), .Z(n5147) );
  NBUFFX2 U5096 ( .INP(n5261), .Z(n5148) );
  NBUFFX2 U5097 ( .INP(n5261), .Z(n5149) );
  NBUFFX2 U5098 ( .INP(n5260), .Z(n5150) );
  NBUFFX2 U5099 ( .INP(n5260), .Z(n5151) );
  NBUFFX2 U5100 ( .INP(n5260), .Z(n5152) );
  NBUFFX2 U5101 ( .INP(n5259), .Z(n5153) );
  NBUFFX2 U5102 ( .INP(n5259), .Z(n5154) );
  NBUFFX2 U5103 ( .INP(n5259), .Z(n5155) );
  NBUFFX2 U5104 ( .INP(n5258), .Z(n5156) );
  NBUFFX2 U5105 ( .INP(n5258), .Z(n5157) );
  NBUFFX2 U5106 ( .INP(n5258), .Z(n5158) );
  NBUFFX2 U5107 ( .INP(n5257), .Z(n5159) );
  NBUFFX2 U5108 ( .INP(n5257), .Z(n5160) );
  NBUFFX2 U5109 ( .INP(n5257), .Z(n5161) );
  NBUFFX2 U5110 ( .INP(n5256), .Z(n5162) );
  NBUFFX2 U5111 ( .INP(n5256), .Z(n5163) );
  NBUFFX2 U5112 ( .INP(n5256), .Z(n5164) );
  NBUFFX2 U5113 ( .INP(n5255), .Z(n5165) );
  NBUFFX2 U5114 ( .INP(n5255), .Z(n5166) );
  NBUFFX2 U5115 ( .INP(n5255), .Z(n5167) );
  NBUFFX2 U5116 ( .INP(n5254), .Z(n5168) );
  NBUFFX2 U5117 ( .INP(n5254), .Z(n5169) );
  NBUFFX2 U5118 ( .INP(n5254), .Z(n5170) );
  NBUFFX2 U5119 ( .INP(n5253), .Z(n5171) );
  NBUFFX2 U5120 ( .INP(n5253), .Z(n5172) );
  NBUFFX2 U5121 ( .INP(n5253), .Z(n5173) );
  NBUFFX2 U5122 ( .INP(n5252), .Z(n5174) );
  NBUFFX2 U5123 ( .INP(n5252), .Z(n5175) );
  NBUFFX2 U5124 ( .INP(n5252), .Z(n5176) );
  NBUFFX2 U5125 ( .INP(n5251), .Z(n5177) );
  NBUFFX2 U5126 ( .INP(n5251), .Z(n5178) );
  NBUFFX2 U5127 ( .INP(n5251), .Z(n5179) );
  NBUFFX2 U5128 ( .INP(n5250), .Z(n5180) );
  NBUFFX2 U5129 ( .INP(n5250), .Z(n5181) );
  NBUFFX2 U5130 ( .INP(n5250), .Z(n5182) );
  NBUFFX2 U5131 ( .INP(n5249), .Z(n5183) );
  NBUFFX2 U5132 ( .INP(n5249), .Z(n5184) );
  NBUFFX2 U5133 ( .INP(n5249), .Z(n5185) );
  NBUFFX2 U5134 ( .INP(n5248), .Z(n5186) );
  NBUFFX2 U5135 ( .INP(n5248), .Z(n5187) );
  NBUFFX2 U5136 ( .INP(n5248), .Z(n5188) );
  NBUFFX2 U5137 ( .INP(n5247), .Z(n5189) );
  NBUFFX2 U5138 ( .INP(n5247), .Z(n5190) );
  NBUFFX2 U5139 ( .INP(n5247), .Z(n5191) );
  NBUFFX2 U5140 ( .INP(n5246), .Z(n5192) );
  NBUFFX2 U5141 ( .INP(n5246), .Z(n5193) );
  NBUFFX2 U5142 ( .INP(n5246), .Z(n5194) );
  NBUFFX2 U5143 ( .INP(n5245), .Z(n5195) );
  NBUFFX2 U5144 ( .INP(n5245), .Z(n5196) );
  NBUFFX2 U5145 ( .INP(n5245), .Z(n5197) );
  NBUFFX2 U5146 ( .INP(n5244), .Z(n5198) );
  NBUFFX2 U5147 ( .INP(n5244), .Z(n5199) );
  NBUFFX2 U5148 ( .INP(n5244), .Z(n5200) );
  NBUFFX2 U5149 ( .INP(n5243), .Z(n5201) );
  NBUFFX2 U5150 ( .INP(n5243), .Z(n5202) );
  NBUFFX2 U5151 ( .INP(n5243), .Z(n5203) );
  NBUFFX2 U5152 ( .INP(n5242), .Z(n5204) );
  NBUFFX2 U5153 ( .INP(n5242), .Z(n5205) );
  NBUFFX2 U5154 ( .INP(n5242), .Z(n5206) );
  NBUFFX2 U5155 ( .INP(n5241), .Z(n5207) );
  NBUFFX2 U5156 ( .INP(n5241), .Z(n5208) );
  NBUFFX2 U5157 ( .INP(n5241), .Z(n5209) );
  NBUFFX2 U5158 ( .INP(n5240), .Z(n5210) );
  NBUFFX2 U5159 ( .INP(n5240), .Z(n5211) );
  NBUFFX2 U5160 ( .INP(n5240), .Z(n5212) );
  NBUFFX2 U5161 ( .INP(n5239), .Z(n5213) );
  NBUFFX2 U5162 ( .INP(n5239), .Z(n5214) );
  NBUFFX2 U5163 ( .INP(n5239), .Z(n5215) );
  NBUFFX2 U5164 ( .INP(n5238), .Z(n5216) );
  NBUFFX2 U5165 ( .INP(n5238), .Z(n5217) );
  NBUFFX2 U5166 ( .INP(n5238), .Z(n5218) );
  NBUFFX2 U5167 ( .INP(n5237), .Z(n5219) );
  NBUFFX2 U5168 ( .INP(n5237), .Z(n5220) );
  NBUFFX2 U5169 ( .INP(n5237), .Z(n5221) );
  NBUFFX2 U5170 ( .INP(n5236), .Z(n5222) );
  NBUFFX2 U5171 ( .INP(n5236), .Z(n5223) );
  NBUFFX2 U5172 ( .INP(n5236), .Z(n5224) );
  NBUFFX2 U5173 ( .INP(n5235), .Z(n5225) );
  NBUFFX2 U5174 ( .INP(n5235), .Z(n5226) );
  NBUFFX2 U5175 ( .INP(n5235), .Z(n5227) );
  NBUFFX2 U5176 ( .INP(n5234), .Z(n5228) );
  NBUFFX2 U5177 ( .INP(n5234), .Z(n5229) );
  NBUFFX2 U5178 ( .INP(n5234), .Z(n5230) );
  NBUFFX2 U5179 ( .INP(n5233), .Z(n5231) );
  NBUFFX2 U5180 ( .INP(n5233), .Z(n5232) );
  NBUFFX2 U5181 ( .INP(n5362), .Z(n5233) );
  NBUFFX2 U5182 ( .INP(n5361), .Z(n5234) );
  NBUFFX2 U5183 ( .INP(n5361), .Z(n5235) );
  NBUFFX2 U5184 ( .INP(n5361), .Z(n5236) );
  NBUFFX2 U5185 ( .INP(n5360), .Z(n5237) );
  NBUFFX2 U5186 ( .INP(n5360), .Z(n5238) );
  NBUFFX2 U5187 ( .INP(n5360), .Z(n5239) );
  NBUFFX2 U5188 ( .INP(n5359), .Z(n5240) );
  NBUFFX2 U5189 ( .INP(n5359), .Z(n5241) );
  NBUFFX2 U5190 ( .INP(n5359), .Z(n5242) );
  NBUFFX2 U5191 ( .INP(n5358), .Z(n5243) );
  NBUFFX2 U5192 ( .INP(n5358), .Z(n5244) );
  NBUFFX2 U5193 ( .INP(n5358), .Z(n5245) );
  NBUFFX2 U5194 ( .INP(n5357), .Z(n5246) );
  NBUFFX2 U5195 ( .INP(n5357), .Z(n5247) );
  NBUFFX2 U5196 ( .INP(n5357), .Z(n5248) );
  NBUFFX2 U5197 ( .INP(n5356), .Z(n5249) );
  NBUFFX2 U5198 ( .INP(n5356), .Z(n5250) );
  NBUFFX2 U5199 ( .INP(n5356), .Z(n5251) );
  NBUFFX2 U5200 ( .INP(n5355), .Z(n5252) );
  NBUFFX2 U5201 ( .INP(n5355), .Z(n5253) );
  NBUFFX2 U5202 ( .INP(n5355), .Z(n5254) );
  NBUFFX2 U5203 ( .INP(n5354), .Z(n5255) );
  NBUFFX2 U5204 ( .INP(n5354), .Z(n5256) );
  NBUFFX2 U5205 ( .INP(n5354), .Z(n5257) );
  NBUFFX2 U5206 ( .INP(n5353), .Z(n5258) );
  NBUFFX2 U5207 ( .INP(n5353), .Z(n5259) );
  NBUFFX2 U5208 ( .INP(n5353), .Z(n5260) );
  NBUFFX2 U5209 ( .INP(n5352), .Z(n5261) );
  NBUFFX2 U5210 ( .INP(n5352), .Z(n5262) );
  NBUFFX2 U5211 ( .INP(n5352), .Z(n5263) );
  NBUFFX2 U5212 ( .INP(n5351), .Z(n5264) );
  NBUFFX2 U5213 ( .INP(n5351), .Z(n5265) );
  NBUFFX2 U5214 ( .INP(n5351), .Z(n5266) );
  NBUFFX2 U5215 ( .INP(n5350), .Z(n5267) );
  NBUFFX2 U5216 ( .INP(n5350), .Z(n5268) );
  NBUFFX2 U5217 ( .INP(n5350), .Z(n5269) );
  NBUFFX2 U5218 ( .INP(n5349), .Z(n5270) );
  NBUFFX2 U5219 ( .INP(n5349), .Z(n5271) );
  NBUFFX2 U5220 ( .INP(n5349), .Z(n5272) );
  NBUFFX2 U5221 ( .INP(n5348), .Z(n5273) );
  NBUFFX2 U5222 ( .INP(n5348), .Z(n5274) );
  NBUFFX2 U5223 ( .INP(n5348), .Z(n5275) );
  NBUFFX2 U5224 ( .INP(n5347), .Z(n5276) );
  NBUFFX2 U5225 ( .INP(n5347), .Z(n5277) );
  NBUFFX2 U5226 ( .INP(n5347), .Z(n5278) );
  NBUFFX2 U5227 ( .INP(n5346), .Z(n5279) );
  NBUFFX2 U5228 ( .INP(n5346), .Z(n5280) );
  NBUFFX2 U5229 ( .INP(n5346), .Z(n5281) );
  NBUFFX2 U5230 ( .INP(n5345), .Z(n5282) );
  NBUFFX2 U5231 ( .INP(n5345), .Z(n5283) );
  NBUFFX2 U5232 ( .INP(n5345), .Z(n5284) );
  NBUFFX2 U5233 ( .INP(n5344), .Z(n5285) );
  NBUFFX2 U5234 ( .INP(n5344), .Z(n5286) );
  NBUFFX2 U5235 ( .INP(n5344), .Z(n5287) );
  NBUFFX2 U5236 ( .INP(n5343), .Z(n5288) );
  NBUFFX2 U5237 ( .INP(n5343), .Z(n5289) );
  NBUFFX2 U5238 ( .INP(n5343), .Z(n5290) );
  NBUFFX2 U5239 ( .INP(n5342), .Z(n5291) );
  NBUFFX2 U5240 ( .INP(n5342), .Z(n5292) );
  NBUFFX2 U5241 ( .INP(n5342), .Z(n5293) );
  NBUFFX2 U5242 ( .INP(n5341), .Z(n5294) );
  NBUFFX2 U5243 ( .INP(n5341), .Z(n5295) );
  NBUFFX2 U5244 ( .INP(n5341), .Z(n5296) );
  NBUFFX2 U5245 ( .INP(n5340), .Z(n5297) );
  NBUFFX2 U5246 ( .INP(n5340), .Z(n5298) );
  NBUFFX2 U5247 ( .INP(n5340), .Z(n5299) );
  NBUFFX2 U5248 ( .INP(n5339), .Z(n5300) );
  NBUFFX2 U5249 ( .INP(n5339), .Z(n5301) );
  NBUFFX2 U5250 ( .INP(n5339), .Z(n5302) );
  NBUFFX2 U5251 ( .INP(n5338), .Z(n5303) );
  NBUFFX2 U5252 ( .INP(n5338), .Z(n5304) );
  NBUFFX2 U5253 ( .INP(n5338), .Z(n5305) );
  NBUFFX2 U5254 ( .INP(n5337), .Z(n5306) );
  NBUFFX2 U5255 ( .INP(n5337), .Z(n5307) );
  NBUFFX2 U5256 ( .INP(n5337), .Z(n5308) );
  NBUFFX2 U5257 ( .INP(n5336), .Z(n5309) );
  NBUFFX2 U5258 ( .INP(n5336), .Z(n5310) );
  NBUFFX2 U5259 ( .INP(n5336), .Z(n5311) );
  NBUFFX2 U5260 ( .INP(n5335), .Z(n5312) );
  NBUFFX2 U5261 ( .INP(n5335), .Z(n5313) );
  NBUFFX2 U5262 ( .INP(n5335), .Z(n5314) );
  NBUFFX2 U5263 ( .INP(n5334), .Z(n5315) );
  NBUFFX2 U5264 ( .INP(n5334), .Z(n5316) );
  NBUFFX2 U5265 ( .INP(n5334), .Z(n5317) );
  NBUFFX2 U5266 ( .INP(n5333), .Z(n5318) );
  NBUFFX2 U5267 ( .INP(n5333), .Z(n5319) );
  NBUFFX2 U5268 ( .INP(n5333), .Z(n5320) );
  NBUFFX2 U5269 ( .INP(n5332), .Z(n5321) );
  NBUFFX2 U5270 ( .INP(n5332), .Z(n5322) );
  NBUFFX2 U5271 ( .INP(n5332), .Z(n5323) );
  NBUFFX2 U5272 ( .INP(n5331), .Z(n5324) );
  NBUFFX2 U5273 ( .INP(n5331), .Z(n5325) );
  NBUFFX2 U5274 ( .INP(n5331), .Z(n5326) );
  NBUFFX2 U5275 ( .INP(n5330), .Z(n5327) );
  NBUFFX2 U5276 ( .INP(n5330), .Z(n5328) );
  NBUFFX2 U5277 ( .INP(n5330), .Z(n5329) );
  NBUFFX2 U5278 ( .INP(n5373), .Z(n5330) );
  NBUFFX2 U5279 ( .INP(n5373), .Z(n5331) );
  NBUFFX2 U5280 ( .INP(n5373), .Z(n5332) );
  NBUFFX2 U5281 ( .INP(n5372), .Z(n5333) );
  NBUFFX2 U5282 ( .INP(n5372), .Z(n5334) );
  NBUFFX2 U5283 ( .INP(n5372), .Z(n5335) );
  NBUFFX2 U5284 ( .INP(n5371), .Z(n5336) );
  NBUFFX2 U5285 ( .INP(n5371), .Z(n5337) );
  NBUFFX2 U5286 ( .INP(n5371), .Z(n5338) );
  NBUFFX2 U5287 ( .INP(n5370), .Z(n5339) );
  NBUFFX2 U5288 ( .INP(n5370), .Z(n5340) );
  NBUFFX2 U5289 ( .INP(n5370), .Z(n5341) );
  NBUFFX2 U5290 ( .INP(n5369), .Z(n5342) );
  NBUFFX2 U5291 ( .INP(n5369), .Z(n5343) );
  NBUFFX2 U5292 ( .INP(n5369), .Z(n5344) );
  NBUFFX2 U5293 ( .INP(n5368), .Z(n5345) );
  NBUFFX2 U5294 ( .INP(n5368), .Z(n5346) );
  NBUFFX2 U5295 ( .INP(n5368), .Z(n5347) );
  NBUFFX2 U5296 ( .INP(n5367), .Z(n5348) );
  NBUFFX2 U5297 ( .INP(n5367), .Z(n5349) );
  NBUFFX2 U5298 ( .INP(n5367), .Z(n5350) );
  NBUFFX2 U5299 ( .INP(n5366), .Z(n5351) );
  NBUFFX2 U5300 ( .INP(n5366), .Z(n5352) );
  NBUFFX2 U5301 ( .INP(n5366), .Z(n5353) );
  NBUFFX2 U5302 ( .INP(n5365), .Z(n5354) );
  NBUFFX2 U5303 ( .INP(n5365), .Z(n5355) );
  NBUFFX2 U5304 ( .INP(n5365), .Z(n5356) );
  NBUFFX2 U5305 ( .INP(n5364), .Z(n5357) );
  NBUFFX2 U5306 ( .INP(n5364), .Z(n5358) );
  NBUFFX2 U5307 ( .INP(n5364), .Z(n5359) );
  NBUFFX2 U5308 ( .INP(n5363), .Z(n5360) );
  NBUFFX2 U5309 ( .INP(n5363), .Z(n5361) );
  NBUFFX2 U5310 ( .INP(n5363), .Z(n5362) );
  NBUFFX2 U5311 ( .INP(n5377), .Z(n5363) );
  NBUFFX2 U5312 ( .INP(n5377), .Z(n5364) );
  NBUFFX2 U5313 ( .INP(n5376), .Z(n5365) );
  NBUFFX2 U5314 ( .INP(n5376), .Z(n5366) );
  NBUFFX2 U5315 ( .INP(n5376), .Z(n5367) );
  NBUFFX2 U5316 ( .INP(n5375), .Z(n5368) );
  NBUFFX2 U5317 ( .INP(n5375), .Z(n5369) );
  NBUFFX2 U5318 ( .INP(n5375), .Z(n5370) );
  NBUFFX2 U5319 ( .INP(n5374), .Z(n5371) );
  NBUFFX2 U5320 ( .INP(n5374), .Z(n5372) );
  NBUFFX2 U5321 ( .INP(n5374), .Z(n5373) );
  NBUFFX2 U5322 ( .INP(test_se), .Z(n5374) );
  NBUFFX2 U5323 ( .INP(test_se), .Z(n5375) );
  NBUFFX2 U5324 ( .INP(test_se), .Z(n5376) );
  NBUFFX2 U5325 ( .INP(test_se), .Z(n5377) );
  INVX0 U5326 ( .INP(n5390), .ZN(n5378) );
  INVX0 U5327 ( .INP(n5390), .ZN(n5379) );
  INVX0 U5328 ( .INP(n5390), .ZN(n5380) );
  INVX0 U5329 ( .INP(n5390), .ZN(n5381) );
  INVX0 U5330 ( .INP(n5390), .ZN(n5382) );
  INVX0 U5331 ( .INP(n5390), .ZN(n5383) );
  INVX0 U5332 ( .INP(n5390), .ZN(n5384) );
  INVX0 U5333 ( .INP(n5390), .ZN(n5385) );
  INVX0 U5334 ( .INP(n5390), .ZN(n5386) );
  INVX0 U5335 ( .INP(n5390), .ZN(n5387) );
  INVX0 U5336 ( .INP(n5390), .ZN(n5388) );
  INVX0 U5337 ( .INP(n5390), .ZN(n5389) );
  INVX0 U5338 ( .INP(TM1), .ZN(n5390) );
  NBUFFX2 U5339 ( .INP(n5454), .Z(n5391) );
  NBUFFX2 U5340 ( .INP(n5454), .Z(n5392) );
  NBUFFX2 U5341 ( .INP(n5454), .Z(n5393) );
  NBUFFX2 U5342 ( .INP(n5453), .Z(n5394) );
  NBUFFX2 U5343 ( .INP(n5453), .Z(n5395) );
  NBUFFX2 U5344 ( .INP(n5453), .Z(n5396) );
  NBUFFX2 U5345 ( .INP(n5452), .Z(n5397) );
  NBUFFX2 U5346 ( .INP(n5452), .Z(n5398) );
  NBUFFX2 U5347 ( .INP(n5452), .Z(n5399) );
  NBUFFX2 U5348 ( .INP(n5451), .Z(n5400) );
  NBUFFX2 U5349 ( .INP(n5451), .Z(n5401) );
  NBUFFX2 U5350 ( .INP(n5451), .Z(n5402) );
  NBUFFX2 U5351 ( .INP(n5450), .Z(n5403) );
  NBUFFX2 U5352 ( .INP(n5450), .Z(n5404) );
  NBUFFX2 U5353 ( .INP(n5450), .Z(n5405) );
  NBUFFX2 U5354 ( .INP(n5449), .Z(n5406) );
  NBUFFX2 U5355 ( .INP(n5449), .Z(n5407) );
  NBUFFX2 U5356 ( .INP(n5449), .Z(n5408) );
  NBUFFX2 U5357 ( .INP(n5448), .Z(n5409) );
  NBUFFX2 U5358 ( .INP(n5448), .Z(n5410) );
  NBUFFX2 U5359 ( .INP(n5448), .Z(n5411) );
  NBUFFX2 U5360 ( .INP(n5447), .Z(n5412) );
  NBUFFX2 U5361 ( .INP(n5447), .Z(n5413) );
  NBUFFX2 U5362 ( .INP(n5447), .Z(n5414) );
  NBUFFX2 U5363 ( .INP(n5446), .Z(n5415) );
  NBUFFX2 U5364 ( .INP(n5446), .Z(n5416) );
  NBUFFX2 U5365 ( .INP(n5446), .Z(n5417) );
  NBUFFX2 U5366 ( .INP(n5445), .Z(n5418) );
  NBUFFX2 U5367 ( .INP(n5445), .Z(n5419) );
  NBUFFX2 U5368 ( .INP(n5445), .Z(n5420) );
  NBUFFX2 U5369 ( .INP(n5444), .Z(n5421) );
  NBUFFX2 U5370 ( .INP(n5444), .Z(n5422) );
  NBUFFX2 U5371 ( .INP(n5444), .Z(n5423) );
  NBUFFX2 U5372 ( .INP(n5443), .Z(n5424) );
  NBUFFX2 U5373 ( .INP(n5443), .Z(n5425) );
  NBUFFX2 U5374 ( .INP(n5443), .Z(n5426) );
  NBUFFX2 U5375 ( .INP(n5442), .Z(n5427) );
  NBUFFX2 U5376 ( .INP(n5442), .Z(n5428) );
  NBUFFX2 U5377 ( .INP(n5442), .Z(n5429) );
  NBUFFX2 U5378 ( .INP(n5441), .Z(n5430) );
  NBUFFX2 U5379 ( .INP(n5441), .Z(n5431) );
  NBUFFX2 U5380 ( .INP(n5441), .Z(n5432) );
  NBUFFX2 U5381 ( .INP(n5440), .Z(n5433) );
  NBUFFX2 U5382 ( .INP(n5440), .Z(n5434) );
  NBUFFX2 U5383 ( .INP(n5440), .Z(n5435) );
  NBUFFX2 U5384 ( .INP(n5439), .Z(n5436) );
  NBUFFX2 U5385 ( .INP(n5439), .Z(n5437) );
  NBUFFX2 U5386 ( .INP(n5439), .Z(n5438) );
  NBUFFX2 U5387 ( .INP(n5460), .Z(n5439) );
  NBUFFX2 U5388 ( .INP(n5459), .Z(n5440) );
  NBUFFX2 U5389 ( .INP(n5459), .Z(n5441) );
  NBUFFX2 U5390 ( .INP(n5459), .Z(n5442) );
  NBUFFX2 U5391 ( .INP(n5458), .Z(n5443) );
  NBUFFX2 U5392 ( .INP(n5458), .Z(n5444) );
  NBUFFX2 U5393 ( .INP(n5458), .Z(n5445) );
  NBUFFX2 U5394 ( .INP(n5457), .Z(n5446) );
  NBUFFX2 U5395 ( .INP(n5457), .Z(n5447) );
  NBUFFX2 U5396 ( .INP(n5457), .Z(n5448) );
  NBUFFX2 U5397 ( .INP(n5456), .Z(n5449) );
  NBUFFX2 U5398 ( .INP(n5456), .Z(n5450) );
  NBUFFX2 U5399 ( .INP(n5456), .Z(n5451) );
  NBUFFX2 U5400 ( .INP(n5455), .Z(n5452) );
  NBUFFX2 U5401 ( .INP(n5455), .Z(n5453) );
  NBUFFX2 U5402 ( .INP(n5455), .Z(n5454) );
  NBUFFX2 U5403 ( .INP(RESET), .Z(n5455) );
  NBUFFX2 U5404 ( .INP(RESET), .Z(n5456) );
  NBUFFX2 U5405 ( .INP(RESET), .Z(n5457) );
  NBUFFX2 U5406 ( .INP(RESET), .Z(n5458) );
  NBUFFX2 U5407 ( .INP(RESET), .Z(n5459) );
  NBUFFX2 U5408 ( .INP(RESET), .Z(n5460) );
  INVX0 U5409 ( .INP(n5391), .ZN(n5461) );
  INVX0 U5410 ( .INP(n5391), .ZN(n5462) );
  INVX0 U5411 ( .INP(n5391), .ZN(n5463) );
  INVX0 U5412 ( .INP(n5391), .ZN(n5464) );
  INVX0 U5413 ( .INP(n5391), .ZN(n5465) );
  INVX0 U5414 ( .INP(n5391), .ZN(n5466) );
  INVX0 U5415 ( .INP(n5391), .ZN(n5467) );
  INVX0 U5416 ( .INP(n5391), .ZN(n5468) );
  INVX0 U5417 ( .INP(n5392), .ZN(n5469) );
  INVX0 U5418 ( .INP(n5392), .ZN(n5470) );
  INVX0 U5419 ( .INP(n5392), .ZN(n5471) );
  INVX0 U5420 ( .INP(n5392), .ZN(n5472) );
  INVX0 U5421 ( .INP(n5392), .ZN(n5473) );
  INVX0 U5422 ( .INP(n5392), .ZN(n5474) );
  INVX0 U5423 ( .INP(n5392), .ZN(n5475) );
  INVX0 U5424 ( .INP(n5392), .ZN(n5476) );
  INVX0 U5425 ( .INP(n5393), .ZN(n5477) );
  INVX0 U5426 ( .INP(n5393), .ZN(n5478) );
  INVX0 U5427 ( .INP(n5393), .ZN(n5479) );
  INVX0 U5428 ( .INP(n5393), .ZN(n5480) );
  INVX0 U5429 ( .INP(n5393), .ZN(n5481) );
  INVX0 U5430 ( .INP(n5393), .ZN(n5482) );
  INVX0 U5431 ( .INP(n5393), .ZN(n5483) );
  INVX0 U5432 ( .INP(n5393), .ZN(n5484) );
  INVX0 U5433 ( .INP(n5394), .ZN(n5485) );
  INVX0 U5434 ( .INP(n5394), .ZN(n5486) );
  INVX0 U5435 ( .INP(n5394), .ZN(n5487) );
  INVX0 U5436 ( .INP(n5394), .ZN(n5488) );
  INVX0 U5437 ( .INP(n5394), .ZN(n5489) );
  INVX0 U5438 ( .INP(n5394), .ZN(n5490) );
  INVX0 U5439 ( .INP(n5394), .ZN(n5491) );
  INVX0 U5440 ( .INP(n5394), .ZN(n5492) );
  INVX0 U5441 ( .INP(n5395), .ZN(n5493) );
  INVX0 U5442 ( .INP(n5395), .ZN(n5494) );
  INVX0 U5443 ( .INP(n5395), .ZN(n5495) );
  INVX0 U5444 ( .INP(n5395), .ZN(n5496) );
  INVX0 U5445 ( .INP(n5395), .ZN(n5497) );
  INVX0 U5446 ( .INP(n5395), .ZN(n5498) );
  INVX0 U5447 ( .INP(n5395), .ZN(n5499) );
  INVX0 U5448 ( .INP(n5395), .ZN(n5500) );
  INVX0 U5449 ( .INP(n5396), .ZN(n5501) );
  INVX0 U5450 ( .INP(n5396), .ZN(n5502) );
  INVX0 U5451 ( .INP(n5396), .ZN(n5503) );
  INVX0 U5452 ( .INP(n5396), .ZN(n5504) );
  INVX0 U5453 ( .INP(n5396), .ZN(n5505) );
  INVX0 U5454 ( .INP(n5396), .ZN(n5506) );
  INVX0 U5455 ( .INP(n5396), .ZN(n5507) );
  INVX0 U5456 ( .INP(n5397), .ZN(n5508) );
  INVX0 U5457 ( .INP(n5397), .ZN(n5509) );
  INVX0 U5458 ( .INP(n5397), .ZN(n5510) );
  INVX0 U5459 ( .INP(n5397), .ZN(n5511) );
  INVX0 U5460 ( .INP(n5397), .ZN(n5512) );
  INVX0 U5461 ( .INP(n5397), .ZN(n5513) );
  INVX0 U5462 ( .INP(n5397), .ZN(n5514) );
  INVX0 U5463 ( .INP(n5397), .ZN(n5515) );
  INVX0 U5464 ( .INP(n5398), .ZN(n5516) );
  INVX0 U5465 ( .INP(n5398), .ZN(n5517) );
  INVX0 U5466 ( .INP(n5398), .ZN(n5518) );
  INVX0 U5467 ( .INP(n5398), .ZN(n5519) );
  INVX0 U5468 ( .INP(n5398), .ZN(n5520) );
  INVX0 U5469 ( .INP(n5398), .ZN(n5521) );
  INVX0 U5470 ( .INP(n5398), .ZN(n5522) );
  INVX0 U5471 ( .INP(n5398), .ZN(n5523) );
  INVX0 U5472 ( .INP(n5399), .ZN(n5524) );
  INVX0 U5473 ( .INP(n5399), .ZN(n5525) );
  INVX0 U5474 ( .INP(n5399), .ZN(n5526) );
  INVX0 U5475 ( .INP(n5399), .ZN(n5527) );
  INVX0 U5476 ( .INP(n5399), .ZN(n5528) );
  INVX0 U5477 ( .INP(n5399), .ZN(n5529) );
  INVX0 U5478 ( .INP(n5399), .ZN(n5530) );
  INVX0 U5479 ( .INP(n5399), .ZN(n5531) );
  INVX0 U5480 ( .INP(n5400), .ZN(n5532) );
  INVX0 U5481 ( .INP(n5400), .ZN(n5533) );
  INVX0 U5482 ( .INP(n5400), .ZN(n5534) );
  INVX0 U5483 ( .INP(n5400), .ZN(n5535) );
  INVX0 U5484 ( .INP(n5400), .ZN(n5536) );
  INVX0 U5485 ( .INP(n5400), .ZN(n5537) );
  INVX0 U5486 ( .INP(n5400), .ZN(n5538) );
  INVX0 U5487 ( .INP(n5400), .ZN(n5539) );
  INVX0 U5488 ( .INP(n5401), .ZN(n5540) );
  INVX0 U5489 ( .INP(n5396), .ZN(n5541) );
  NBUFFX2 U5490 ( .INP(n5724), .Z(n5686) );
  NBUFFX2 U5491 ( .INP(n5724), .Z(n5687) );
  NBUFFX2 U5492 ( .INP(n5723), .Z(n5688) );
  NBUFFX2 U5493 ( .INP(n5723), .Z(n5689) );
  NBUFFX2 U5494 ( .INP(n5723), .Z(n5690) );
  NBUFFX2 U5495 ( .INP(n5722), .Z(n5691) );
  NBUFFX2 U5496 ( .INP(n5722), .Z(n5692) );
  NBUFFX2 U5497 ( .INP(n5722), .Z(n5693) );
  NBUFFX2 U5498 ( .INP(n5721), .Z(n5694) );
  NBUFFX2 U5499 ( .INP(n5721), .Z(n5695) );
  NBUFFX2 U5500 ( .INP(n5721), .Z(n5696) );
  NBUFFX2 U5501 ( .INP(n5720), .Z(n5697) );
  NBUFFX2 U5502 ( .INP(n5720), .Z(n5698) );
  NBUFFX2 U5503 ( .INP(n5720), .Z(n5699) );
  NBUFFX2 U5504 ( .INP(n5719), .Z(n5700) );
  NBUFFX2 U5505 ( .INP(n5719), .Z(n5701) );
  NBUFFX2 U5506 ( .INP(n5719), .Z(n5702) );
  NBUFFX2 U5507 ( .INP(n5718), .Z(n5703) );
  NBUFFX2 U5508 ( .INP(n5718), .Z(n5704) );
  NBUFFX2 U5509 ( .INP(n5718), .Z(n5705) );
  NBUFFX2 U5510 ( .INP(n5717), .Z(n5706) );
  NBUFFX2 U5511 ( .INP(n5717), .Z(n5707) );
  NBUFFX2 U5512 ( .INP(n5717), .Z(n5708) );
  NBUFFX2 U5513 ( .INP(n5716), .Z(n5709) );
  NBUFFX2 U5514 ( .INP(n5716), .Z(n5710) );
  NBUFFX2 U5515 ( .INP(n5716), .Z(n5711) );
  NBUFFX2 U5516 ( .INP(n5715), .Z(n5712) );
  NBUFFX2 U5517 ( .INP(n5715), .Z(n5713) );
  NBUFFX2 U5518 ( .INP(n5715), .Z(n5714) );
  NBUFFX2 U5519 ( .INP(CK), .Z(n5715) );
  NBUFFX2 U5520 ( .INP(CK), .Z(n5716) );
  NBUFFX2 U5521 ( .INP(n5724), .Z(n5717) );
  NBUFFX2 U5522 ( .INP(CK), .Z(n5718) );
  NBUFFX2 U5523 ( .INP(n5720), .Z(n5719) );
  NBUFFX2 U5524 ( .INP(CK), .Z(n5720) );
  NBUFFX2 U5525 ( .INP(n5715), .Z(n5721) );
  NBUFFX2 U5526 ( .INP(n5716), .Z(n5722) );
  NBUFFX2 U5527 ( .INP(n5718), .Z(n5723) );
  NBUFFX2 U5528 ( .INP(n5555), .Z(n5724) );
  AND2X1 U5529 ( .IN1(n5435), .IN2(n5390), .Q(n3278) );
  INVX0 U5530 ( .INP(n5725), .ZN(WX9789) );
  OR2X1 U5531 ( .IN1(n5461), .IN2(n9534), .Q(n5725) );
  INVX0 U5532 ( .INP(n5726), .ZN(WX9787) );
  OR2X1 U5533 ( .IN1(n5473), .IN2(n9537), .Q(n5726) );
  INVX0 U5534 ( .INP(n5727), .ZN(WX9785) );
  OR2X1 U5535 ( .IN1(n5473), .IN2(n9538), .Q(n5727) );
  INVX0 U5536 ( .INP(n5728), .ZN(WX9783) );
  OR2X1 U5537 ( .IN1(n5473), .IN2(n9541), .Q(n5728) );
  AND2X1 U5538 ( .IN1(test_so80), .IN2(n5415), .Q(WX9781) );
  INVX0 U5539 ( .INP(n5729), .ZN(WX9779) );
  OR2X1 U5540 ( .IN1(n5473), .IN2(n9542), .Q(n5729) );
  INVX0 U5541 ( .INP(n5730), .ZN(WX9777) );
  OR2X1 U5542 ( .IN1(n5473), .IN2(n9543), .Q(n5730) );
  INVX0 U5543 ( .INP(n5731), .ZN(WX9775) );
  OR2X1 U5544 ( .IN1(n5473), .IN2(n9544), .Q(n5731) );
  INVX0 U5545 ( .INP(n5732), .ZN(WX9773) );
  OR2X1 U5546 ( .IN1(n5473), .IN2(n9545), .Q(n5732) );
  INVX0 U5547 ( .INP(n5733), .ZN(WX9771) );
  OR2X1 U5548 ( .IN1(n5473), .IN2(n9546), .Q(n5733) );
  INVX0 U5549 ( .INP(n5734), .ZN(WX9769) );
  OR2X1 U5550 ( .IN1(n5473), .IN2(n9547), .Q(n5734) );
  INVX0 U5551 ( .INP(n5735), .ZN(WX9767) );
  OR2X1 U5552 ( .IN1(n5473), .IN2(n9548), .Q(n5735) );
  INVX0 U5553 ( .INP(n5736), .ZN(WX9765) );
  OR2X1 U5554 ( .IN1(n5473), .IN2(n9549), .Q(n5736) );
  INVX0 U5555 ( .INP(n5737), .ZN(WX9763) );
  OR2X1 U5556 ( .IN1(n5473), .IN2(n9550), .Q(n5737) );
  INVX0 U5557 ( .INP(n5738), .ZN(WX9761) );
  OR2X1 U5558 ( .IN1(n5473), .IN2(n9551), .Q(n5738) );
  INVX0 U5559 ( .INP(n5739), .ZN(WX9759) );
  OR2X1 U5560 ( .IN1(n5472), .IN2(n9552), .Q(n5739) );
  OR2X1 U5561 ( .IN1(n5740), .IN2(n5741), .Q(WX9757) );
  OR2X1 U5562 ( .IN1(n5742), .IN2(n5743), .Q(n5741) );
  AND2X1 U5563 ( .IN1(n4889), .IN2(CRC_OUT_2_0), .Q(n5743) );
  AND2X1 U5564 ( .IN1(n436), .IN2(n4884), .Q(n5742) );
  INVX0 U5565 ( .INP(n5744), .ZN(n436) );
  OR2X1 U5566 ( .IN1(n5472), .IN2(n3817), .Q(n5744) );
  OR2X1 U5567 ( .IN1(n5745), .IN2(n5746), .Q(n5740) );
  AND2X1 U5568 ( .IN1(n4926), .IN2(n5747), .Q(n5746) );
  AND2X1 U5569 ( .IN1(n4845), .IN2(n5749), .Q(n5745) );
  OR2X1 U5570 ( .IN1(n5750), .IN2(n5751), .Q(WX9755) );
  OR2X1 U5571 ( .IN1(n5752), .IN2(n5753), .Q(n5751) );
  AND2X1 U5572 ( .IN1(n4903), .IN2(CRC_OUT_2_1), .Q(n5753) );
  AND2X1 U5573 ( .IN1(n435), .IN2(n4884), .Q(n5752) );
  INVX0 U5574 ( .INP(n5754), .ZN(n435) );
  OR2X1 U5575 ( .IN1(n5472), .IN2(n3818), .Q(n5754) );
  OR2X1 U5576 ( .IN1(n5755), .IN2(n5756), .Q(n5750) );
  AND2X1 U5577 ( .IN1(n4934), .IN2(n5757), .Q(n5756) );
  AND2X1 U5578 ( .IN1(n5758), .IN2(n4833), .Q(n5755) );
  OR2X1 U5579 ( .IN1(n5759), .IN2(n5760), .Q(WX9753) );
  OR2X1 U5580 ( .IN1(n5761), .IN2(n5762), .Q(n5760) );
  AND2X1 U5581 ( .IN1(test_so87), .IN2(n4887), .Q(n5762) );
  AND2X1 U5582 ( .IN1(n434), .IN2(n4884), .Q(n5761) );
  INVX0 U5583 ( .INP(n5763), .ZN(n434) );
  OR2X1 U5584 ( .IN1(n5472), .IN2(n3819), .Q(n5763) );
  OR2X1 U5585 ( .IN1(n5764), .IN2(n5765), .Q(n5759) );
  AND2X1 U5586 ( .IN1(n5766), .IN2(n4921), .Q(n5765) );
  AND2X1 U5587 ( .IN1(n4845), .IN2(n5767), .Q(n5764) );
  OR2X1 U5588 ( .IN1(n5768), .IN2(n5769), .Q(WX9751) );
  OR2X1 U5589 ( .IN1(n5770), .IN2(n5771), .Q(n5769) );
  AND2X1 U5590 ( .IN1(n4898), .IN2(CRC_OUT_2_3), .Q(n5771) );
  AND2X1 U5591 ( .IN1(n433), .IN2(n4883), .Q(n5770) );
  INVX0 U5592 ( .INP(n5772), .ZN(n433) );
  OR2X1 U5593 ( .IN1(n5472), .IN2(n3820), .Q(n5772) );
  OR2X1 U5594 ( .IN1(n5773), .IN2(n5774), .Q(n5768) );
  AND2X1 U5595 ( .IN1(n4930), .IN2(n5775), .Q(n5774) );
  AND2X1 U5596 ( .IN1(n5776), .IN2(n4833), .Q(n5773) );
  OR2X1 U5597 ( .IN1(n5777), .IN2(n5778), .Q(WX9749) );
  OR2X1 U5598 ( .IN1(n5779), .IN2(n5780), .Q(n5778) );
  AND2X1 U5599 ( .IN1(n4898), .IN2(CRC_OUT_2_4), .Q(n5780) );
  AND2X1 U5600 ( .IN1(n432), .IN2(n4883), .Q(n5779) );
  INVX0 U5601 ( .INP(n5781), .ZN(n432) );
  OR2X1 U5602 ( .IN1(n5472), .IN2(n3821), .Q(n5781) );
  OR2X1 U5603 ( .IN1(n5782), .IN2(n5783), .Q(n5777) );
  AND2X1 U5604 ( .IN1(n5784), .IN2(n4921), .Q(n5783) );
  AND2X1 U5605 ( .IN1(n4845), .IN2(n5785), .Q(n5782) );
  OR2X1 U5606 ( .IN1(n5786), .IN2(n5787), .Q(WX9747) );
  OR2X1 U5607 ( .IN1(n5788), .IN2(n5789), .Q(n5787) );
  AND2X1 U5608 ( .IN1(n4898), .IN2(CRC_OUT_2_5), .Q(n5789) );
  AND2X1 U5609 ( .IN1(n431), .IN2(n4883), .Q(n5788) );
  INVX0 U5610 ( .INP(n5790), .ZN(n431) );
  OR2X1 U5611 ( .IN1(n5472), .IN2(n3822), .Q(n5790) );
  OR2X1 U5612 ( .IN1(n5791), .IN2(n5792), .Q(n5786) );
  AND2X1 U5613 ( .IN1(n4930), .IN2(n5793), .Q(n5792) );
  AND2X1 U5614 ( .IN1(n4845), .IN2(n5794), .Q(n5791) );
  OR2X1 U5615 ( .IN1(n5795), .IN2(n5796), .Q(WX9745) );
  OR2X1 U5616 ( .IN1(n5797), .IN2(n5798), .Q(n5796) );
  AND2X1 U5617 ( .IN1(n4898), .IN2(CRC_OUT_2_6), .Q(n5798) );
  AND2X1 U5618 ( .IN1(n430), .IN2(n4883), .Q(n5797) );
  INVX0 U5619 ( .INP(n5799), .ZN(n430) );
  OR2X1 U5620 ( .IN1(n5472), .IN2(n3823), .Q(n5799) );
  OR2X1 U5621 ( .IN1(n5800), .IN2(n5801), .Q(n5795) );
  AND2X1 U5622 ( .IN1(n5802), .IN2(n4922), .Q(n5801) );
  AND2X1 U5623 ( .IN1(n4845), .IN2(n5803), .Q(n5800) );
  OR2X1 U5624 ( .IN1(n5804), .IN2(n5805), .Q(WX9743) );
  OR2X1 U5625 ( .IN1(n5806), .IN2(n5807), .Q(n5805) );
  AND2X1 U5626 ( .IN1(n4898), .IN2(CRC_OUT_2_7), .Q(n5807) );
  AND2X1 U5627 ( .IN1(n429), .IN2(n4883), .Q(n5806) );
  INVX0 U5628 ( .INP(n5808), .ZN(n429) );
  OR2X1 U5629 ( .IN1(n5472), .IN2(n3824), .Q(n5808) );
  OR2X1 U5630 ( .IN1(n5809), .IN2(n5810), .Q(n5804) );
  AND2X1 U5631 ( .IN1(n4930), .IN2(n5811), .Q(n5810) );
  AND2X1 U5632 ( .IN1(n4845), .IN2(n5812), .Q(n5809) );
  OR2X1 U5633 ( .IN1(n5813), .IN2(n5814), .Q(WX9741) );
  OR2X1 U5634 ( .IN1(n5815), .IN2(n5816), .Q(n5814) );
  AND2X1 U5635 ( .IN1(n4899), .IN2(CRC_OUT_2_8), .Q(n5816) );
  AND2X1 U5636 ( .IN1(n428), .IN2(n4883), .Q(n5815) );
  INVX0 U5637 ( .INP(n5817), .ZN(n428) );
  OR2X1 U5638 ( .IN1(n5472), .IN2(n3825), .Q(n5817) );
  OR2X1 U5639 ( .IN1(n5818), .IN2(n5819), .Q(n5813) );
  AND2X1 U5640 ( .IN1(n5820), .IN2(n4922), .Q(n5819) );
  AND2X1 U5641 ( .IN1(n4845), .IN2(n5821), .Q(n5818) );
  OR2X1 U5642 ( .IN1(n5822), .IN2(n5823), .Q(WX9739) );
  OR2X1 U5643 ( .IN1(n5824), .IN2(n5825), .Q(n5823) );
  AND2X1 U5644 ( .IN1(n4899), .IN2(CRC_OUT_2_9), .Q(n5825) );
  AND2X1 U5645 ( .IN1(n427), .IN2(n4883), .Q(n5824) );
  INVX0 U5646 ( .INP(n5826), .ZN(n427) );
  OR2X1 U5647 ( .IN1(n5472), .IN2(n3826), .Q(n5826) );
  OR2X1 U5648 ( .IN1(n5827), .IN2(n5828), .Q(n5822) );
  AND2X1 U5649 ( .IN1(n4930), .IN2(n5829), .Q(n5828) );
  AND2X1 U5650 ( .IN1(n4845), .IN2(n5830), .Q(n5827) );
  OR2X1 U5651 ( .IN1(n5831), .IN2(n5832), .Q(WX9737) );
  OR2X1 U5652 ( .IN1(n5833), .IN2(n5834), .Q(n5832) );
  AND2X1 U5653 ( .IN1(n4899), .IN2(CRC_OUT_2_10), .Q(n5834) );
  AND2X1 U5654 ( .IN1(n426), .IN2(n4883), .Q(n5833) );
  INVX0 U5655 ( .INP(n5835), .ZN(n426) );
  OR2X1 U5656 ( .IN1(n5472), .IN2(n3827), .Q(n5835) );
  OR2X1 U5657 ( .IN1(n5836), .IN2(n5837), .Q(n5831) );
  AND2X1 U5658 ( .IN1(n4930), .IN2(n5838), .Q(n5837) );
  AND2X1 U5659 ( .IN1(n4845), .IN2(n5839), .Q(n5836) );
  OR2X1 U5660 ( .IN1(n5840), .IN2(n5841), .Q(WX9735) );
  OR2X1 U5661 ( .IN1(n5842), .IN2(n5843), .Q(n5841) );
  AND2X1 U5662 ( .IN1(n4899), .IN2(CRC_OUT_2_11), .Q(n5843) );
  AND2X1 U5663 ( .IN1(n425), .IN2(n4883), .Q(n5842) );
  INVX0 U5664 ( .INP(n5844), .ZN(n425) );
  OR2X1 U5665 ( .IN1(n5472), .IN2(n3828), .Q(n5844) );
  OR2X1 U5666 ( .IN1(n5845), .IN2(n5846), .Q(n5840) );
  AND2X1 U5667 ( .IN1(n4930), .IN2(n5847), .Q(n5846) );
  AND2X1 U5668 ( .IN1(n4845), .IN2(n5848), .Q(n5845) );
  OR2X1 U5669 ( .IN1(n5849), .IN2(n5850), .Q(WX9733) );
  OR2X1 U5670 ( .IN1(n5851), .IN2(n5852), .Q(n5850) );
  AND2X1 U5671 ( .IN1(n4899), .IN2(CRC_OUT_2_12), .Q(n5852) );
  AND2X1 U5672 ( .IN1(n424), .IN2(n4883), .Q(n5851) );
  INVX0 U5673 ( .INP(n5853), .ZN(n424) );
  OR2X1 U5674 ( .IN1(n5471), .IN2(n3829), .Q(n5853) );
  OR2X1 U5675 ( .IN1(n5854), .IN2(n5855), .Q(n5849) );
  AND2X1 U5676 ( .IN1(n4930), .IN2(n5856), .Q(n5855) );
  AND2X1 U5677 ( .IN1(n4845), .IN2(n5857), .Q(n5854) );
  OR2X1 U5678 ( .IN1(n5858), .IN2(n5859), .Q(WX9731) );
  OR2X1 U5679 ( .IN1(n5860), .IN2(n5861), .Q(n5859) );
  AND2X1 U5680 ( .IN1(n4899), .IN2(CRC_OUT_2_13), .Q(n5861) );
  AND2X1 U5681 ( .IN1(n423), .IN2(n4883), .Q(n5860) );
  INVX0 U5682 ( .INP(n5862), .ZN(n423) );
  OR2X1 U5683 ( .IN1(n5471), .IN2(n3830), .Q(n5862) );
  OR2X1 U5684 ( .IN1(n5863), .IN2(n5864), .Q(n5858) );
  AND2X1 U5685 ( .IN1(n4930), .IN2(n5865), .Q(n5864) );
  AND2X1 U5686 ( .IN1(n4845), .IN2(n5866), .Q(n5863) );
  OR2X1 U5687 ( .IN1(n5867), .IN2(n5868), .Q(WX9729) );
  OR2X1 U5688 ( .IN1(n5869), .IN2(n5870), .Q(n5868) );
  AND2X1 U5689 ( .IN1(n4899), .IN2(CRC_OUT_2_14), .Q(n5870) );
  AND2X1 U5690 ( .IN1(n422), .IN2(n4883), .Q(n5869) );
  INVX0 U5691 ( .INP(n5871), .ZN(n422) );
  OR2X1 U5692 ( .IN1(n5471), .IN2(n3831), .Q(n5871) );
  OR2X1 U5693 ( .IN1(n5872), .IN2(n5873), .Q(n5867) );
  AND2X1 U5694 ( .IN1(n4930), .IN2(n5874), .Q(n5873) );
  AND2X1 U5695 ( .IN1(n5875), .IN2(n4834), .Q(n5872) );
  OR2X1 U5696 ( .IN1(n5876), .IN2(n5877), .Q(WX9727) );
  OR2X1 U5697 ( .IN1(n5878), .IN2(n5879), .Q(n5877) );
  AND2X1 U5698 ( .IN1(n4899), .IN2(CRC_OUT_2_15), .Q(n5879) );
  AND2X1 U5699 ( .IN1(n421), .IN2(n4882), .Q(n5878) );
  INVX0 U5700 ( .INP(n5880), .ZN(n421) );
  OR2X1 U5701 ( .IN1(n5471), .IN2(n3832), .Q(n5880) );
  OR2X1 U5702 ( .IN1(n5881), .IN2(n5882), .Q(n5876) );
  AND2X1 U5703 ( .IN1(n4930), .IN2(n5883), .Q(n5882) );
  AND2X1 U5704 ( .IN1(n4844), .IN2(n5884), .Q(n5881) );
  OR2X1 U5705 ( .IN1(n5885), .IN2(n5886), .Q(WX9725) );
  OR2X1 U5706 ( .IN1(n5887), .IN2(n5888), .Q(n5886) );
  AND2X1 U5707 ( .IN1(n4899), .IN2(CRC_OUT_2_16), .Q(n5888) );
  AND2X1 U5708 ( .IN1(n420), .IN2(n4882), .Q(n5887) );
  INVX0 U5709 ( .INP(n5889), .ZN(n420) );
  OR2X1 U5710 ( .IN1(n5471), .IN2(n3833), .Q(n5889) );
  OR2X1 U5711 ( .IN1(n5890), .IN2(n5891), .Q(n5885) );
  AND2X1 U5712 ( .IN1(n4930), .IN2(n5892), .Q(n5891) );
  AND2X1 U5713 ( .IN1(n5893), .IN2(n4834), .Q(n5890) );
  OR2X1 U5714 ( .IN1(n5894), .IN2(n5895), .Q(WX9723) );
  OR2X1 U5715 ( .IN1(n5896), .IN2(n5897), .Q(n5895) );
  AND2X1 U6483 ( .IN1(n4899), .IN2(CRC_OUT_2_17), .Q(n5897) );
  AND2X1 U6484 ( .IN1(n419), .IN2(n4882), .Q(n5896) );
  INVX0 U6485 ( .INP(n5898), .ZN(n419) );
  OR2X1 U6486 ( .IN1(n5471), .IN2(n3834), .Q(n5898) );
  OR2X1 U6487 ( .IN1(n5899), .IN2(n5900), .Q(n5894) );
  AND2X1 U6488 ( .IN1(n4931), .IN2(n5901), .Q(n5900) );
  AND2X1 U6489 ( .IN1(n4844), .IN2(n5902), .Q(n5899) );
  OR2X1 U6490 ( .IN1(n5903), .IN2(n5904), .Q(WX9721) );
  OR2X1 U6491 ( .IN1(n5905), .IN2(n5906), .Q(n5904) );
  AND2X1 U6492 ( .IN1(n4899), .IN2(CRC_OUT_2_18), .Q(n5906) );
  AND2X1 U6493 ( .IN1(n418), .IN2(n4882), .Q(n5905) );
  INVX0 U6494 ( .INP(n5907), .ZN(n418) );
  OR2X1 U6495 ( .IN1(n5471), .IN2(n3835), .Q(n5907) );
  OR2X1 U6496 ( .IN1(n5908), .IN2(n5909), .Q(n5903) );
  AND2X1 U6497 ( .IN1(n4931), .IN2(n5910), .Q(n5909) );
  AND2X1 U6498 ( .IN1(n5911), .IN2(n4834), .Q(n5908) );
  OR2X1 U6499 ( .IN1(n5912), .IN2(n5913), .Q(WX9719) );
  OR2X1 U6500 ( .IN1(n5914), .IN2(n5915), .Q(n5913) );
  AND2X1 U6501 ( .IN1(test_so88), .IN2(n4887), .Q(n5915) );
  AND2X1 U6502 ( .IN1(n417), .IN2(n4882), .Q(n5914) );
  INVX0 U6503 ( .INP(n5916), .ZN(n417) );
  OR2X1 U6504 ( .IN1(n5471), .IN2(n3836), .Q(n5916) );
  OR2X1 U6505 ( .IN1(n5917), .IN2(n5918), .Q(n5912) );
  AND2X1 U6506 ( .IN1(n5919), .IN2(n4924), .Q(n5918) );
  AND2X1 U6507 ( .IN1(n4844), .IN2(n5920), .Q(n5917) );
  OR2X1 U6508 ( .IN1(n5921), .IN2(n5922), .Q(WX9717) );
  OR2X1 U6509 ( .IN1(n5923), .IN2(n5924), .Q(n5922) );
  AND2X1 U6510 ( .IN1(n4899), .IN2(CRC_OUT_2_20), .Q(n5924) );
  AND2X1 U6511 ( .IN1(n416), .IN2(n4882), .Q(n5923) );
  INVX0 U6512 ( .INP(n5925), .ZN(n416) );
  OR2X1 U6513 ( .IN1(n5471), .IN2(n3837), .Q(n5925) );
  OR2X1 U6514 ( .IN1(n5926), .IN2(n5927), .Q(n5921) );
  AND2X1 U6515 ( .IN1(n4931), .IN2(n5928), .Q(n5927) );
  AND2X1 U6516 ( .IN1(n5929), .IN2(n4834), .Q(n5926) );
  OR2X1 U6517 ( .IN1(n5930), .IN2(n5931), .Q(WX9715) );
  OR2X1 U6518 ( .IN1(n5932), .IN2(n5933), .Q(n5931) );
  AND2X1 U6519 ( .IN1(n4899), .IN2(CRC_OUT_2_21), .Q(n5933) );
  AND2X1 U6520 ( .IN1(n415), .IN2(n4882), .Q(n5932) );
  INVX0 U6521 ( .INP(n5934), .ZN(n415) );
  OR2X1 U6522 ( .IN1(n5471), .IN2(n3838), .Q(n5934) );
  OR2X1 U6523 ( .IN1(n5935), .IN2(n5936), .Q(n5930) );
  AND2X1 U6524 ( .IN1(n5937), .IN2(n4923), .Q(n5936) );
  AND2X1 U6525 ( .IN1(n4844), .IN2(n5938), .Q(n5935) );
  OR2X1 U6526 ( .IN1(n5939), .IN2(n5940), .Q(WX9713) );
  OR2X1 U6527 ( .IN1(n5941), .IN2(n5942), .Q(n5940) );
  AND2X1 U6528 ( .IN1(n4900), .IN2(CRC_OUT_2_22), .Q(n5942) );
  AND2X1 U6529 ( .IN1(n414), .IN2(n4882), .Q(n5941) );
  INVX0 U6530 ( .INP(n5943), .ZN(n414) );
  OR2X1 U6531 ( .IN1(n5471), .IN2(n3839), .Q(n5943) );
  OR2X1 U6532 ( .IN1(n5944), .IN2(n5945), .Q(n5939) );
  AND2X1 U6533 ( .IN1(n4931), .IN2(n5946), .Q(n5945) );
  AND2X1 U6534 ( .IN1(n4844), .IN2(n5947), .Q(n5944) );
  OR2X1 U6535 ( .IN1(n5948), .IN2(n5949), .Q(WX9711) );
  OR2X1 U6536 ( .IN1(n5950), .IN2(n5951), .Q(n5949) );
  AND2X1 U6537 ( .IN1(n4900), .IN2(CRC_OUT_2_23), .Q(n5951) );
  AND2X1 U6538 ( .IN1(n413), .IN2(n4882), .Q(n5950) );
  INVX0 U6539 ( .INP(n5952), .ZN(n413) );
  OR2X1 U6540 ( .IN1(n5471), .IN2(n3840), .Q(n5952) );
  OR2X1 U6541 ( .IN1(n5953), .IN2(n5954), .Q(n5948) );
  AND2X1 U6542 ( .IN1(n5955), .IN2(n4924), .Q(n5954) );
  AND2X1 U6543 ( .IN1(n4844), .IN2(n5956), .Q(n5953) );
  OR2X1 U6544 ( .IN1(n5957), .IN2(n5958), .Q(WX9709) );
  OR2X1 U6545 ( .IN1(n5959), .IN2(n5960), .Q(n5958) );
  AND2X1 U6546 ( .IN1(n4900), .IN2(CRC_OUT_2_24), .Q(n5960) );
  AND2X1 U6547 ( .IN1(n412), .IN2(n4882), .Q(n5959) );
  INVX0 U6548 ( .INP(n5961), .ZN(n412) );
  OR2X1 U6549 ( .IN1(n5471), .IN2(n3841), .Q(n5961) );
  OR2X1 U6550 ( .IN1(n5962), .IN2(n5963), .Q(n5957) );
  AND2X1 U6551 ( .IN1(n4931), .IN2(n5964), .Q(n5963) );
  AND2X1 U6552 ( .IN1(n4844), .IN2(n5965), .Q(n5962) );
  OR2X1 U6553 ( .IN1(n5966), .IN2(n5967), .Q(WX9707) );
  OR2X1 U6554 ( .IN1(n5968), .IN2(n5969), .Q(n5967) );
  AND2X1 U6555 ( .IN1(n4900), .IN2(CRC_OUT_2_25), .Q(n5969) );
  AND2X1 U6556 ( .IN1(n411), .IN2(n4882), .Q(n5968) );
  INVX0 U6557 ( .INP(n5970), .ZN(n411) );
  OR2X1 U6558 ( .IN1(n5470), .IN2(n3842), .Q(n5970) );
  OR2X1 U6559 ( .IN1(n5971), .IN2(n5972), .Q(n5966) );
  AND2X1 U6560 ( .IN1(n5973), .IN2(n4923), .Q(n5972) );
  AND2X1 U6561 ( .IN1(n4844), .IN2(n5974), .Q(n5971) );
  OR2X1 U6562 ( .IN1(n5975), .IN2(n5976), .Q(WX9705) );
  OR2X1 U6563 ( .IN1(n5977), .IN2(n5978), .Q(n5976) );
  AND2X1 U6564 ( .IN1(n4900), .IN2(CRC_OUT_2_26), .Q(n5978) );
  AND2X1 U6565 ( .IN1(n410), .IN2(n4882), .Q(n5977) );
  INVX0 U6566 ( .INP(n5979), .ZN(n410) );
  OR2X1 U6567 ( .IN1(n5470), .IN2(n3843), .Q(n5979) );
  OR2X1 U6568 ( .IN1(n5980), .IN2(n5981), .Q(n5975) );
  AND2X1 U6569 ( .IN1(n4931), .IN2(n5982), .Q(n5981) );
  AND2X1 U6570 ( .IN1(n4844), .IN2(n5983), .Q(n5980) );
  OR2X1 U6571 ( .IN1(n5984), .IN2(n5985), .Q(WX9703) );
  OR2X1 U6572 ( .IN1(n5986), .IN2(n5987), .Q(n5985) );
  AND2X1 U6573 ( .IN1(n4900), .IN2(CRC_OUT_2_27), .Q(n5987) );
  AND2X1 U6574 ( .IN1(n409), .IN2(n4881), .Q(n5986) );
  INVX0 U6575 ( .INP(n5988), .ZN(n409) );
  OR2X1 U6576 ( .IN1(n5470), .IN2(n3844), .Q(n5988) );
  OR2X1 U6577 ( .IN1(n5989), .IN2(n5990), .Q(n5984) );
  AND2X1 U6578 ( .IN1(n4931), .IN2(n5991), .Q(n5990) );
  AND2X1 U6579 ( .IN1(n4844), .IN2(n5992), .Q(n5989) );
  OR2X1 U6580 ( .IN1(n5993), .IN2(n5994), .Q(WX9701) );
  OR2X1 U6581 ( .IN1(n5995), .IN2(n5996), .Q(n5994) );
  AND2X1 U6582 ( .IN1(n4900), .IN2(CRC_OUT_2_28), .Q(n5996) );
  AND2X1 U6583 ( .IN1(n408), .IN2(n4881), .Q(n5995) );
  INVX0 U6584 ( .INP(n5997), .ZN(n408) );
  OR2X1 U6585 ( .IN1(n5470), .IN2(n3845), .Q(n5997) );
  OR2X1 U6586 ( .IN1(n5998), .IN2(n5999), .Q(n5993) );
  AND2X1 U6587 ( .IN1(n4931), .IN2(n6000), .Q(n5999) );
  AND2X1 U6588 ( .IN1(n4844), .IN2(n6001), .Q(n5998) );
  OR2X1 U6589 ( .IN1(n6002), .IN2(n6003), .Q(WX9699) );
  OR2X1 U6590 ( .IN1(n6004), .IN2(n6005), .Q(n6003) );
  AND2X1 U6591 ( .IN1(n4900), .IN2(CRC_OUT_2_29), .Q(n6005) );
  AND2X1 U6592 ( .IN1(n407), .IN2(n4881), .Q(n6004) );
  INVX0 U6593 ( .INP(n6006), .ZN(n407) );
  OR2X1 U6594 ( .IN1(n5470), .IN2(n3846), .Q(n6006) );
  OR2X1 U6595 ( .IN1(n6007), .IN2(n6008), .Q(n6002) );
  AND2X1 U6596 ( .IN1(n4931), .IN2(n6009), .Q(n6008) );
  AND2X1 U6597 ( .IN1(n4844), .IN2(n6010), .Q(n6007) );
  OR2X1 U6598 ( .IN1(n6011), .IN2(n6012), .Q(WX9697) );
  OR2X1 U6599 ( .IN1(n6013), .IN2(n6014), .Q(n6012) );
  AND2X1 U6600 ( .IN1(n4900), .IN2(CRC_OUT_2_30), .Q(n6014) );
  AND2X1 U6601 ( .IN1(n406), .IN2(n4881), .Q(n6013) );
  INVX0 U6602 ( .INP(n6015), .ZN(n406) );
  OR2X1 U6603 ( .IN1(n5470), .IN2(n3847), .Q(n6015) );
  OR2X1 U6604 ( .IN1(n6016), .IN2(n6017), .Q(n6011) );
  AND2X1 U6605 ( .IN1(n4931), .IN2(n6018), .Q(n6017) );
  AND2X1 U6606 ( .IN1(n4844), .IN2(n6019), .Q(n6016) );
  OR2X1 U6607 ( .IN1(n6020), .IN2(n6021), .Q(WX9695) );
  OR2X1 U6608 ( .IN1(n6022), .IN2(n6023), .Q(n6021) );
  AND2X1 U6609 ( .IN1(n2245), .IN2(WX9536), .Q(n6023) );
  AND2X1 U6610 ( .IN1(n4900), .IN2(CRC_OUT_2_31), .Q(n6022) );
  OR2X1 U6611 ( .IN1(n6024), .IN2(n6025), .Q(n6020) );
  AND2X1 U6612 ( .IN1(n4931), .IN2(n6026), .Q(n6025) );
  AND2X1 U6613 ( .IN1(n6027), .IN2(n4836), .Q(n6024) );
  AND2X1 U6614 ( .IN1(n4825), .IN2(n5414), .Q(WX9597) );
  AND2X1 U6615 ( .IN1(n6028), .IN2(n5414), .Q(WX9084) );
  XOR2X1 U6616 ( .IN1(CRC_OUT_3_30), .IN2(n4594), .Q(n6028) );
  AND2X1 U6617 ( .IN1(n6029), .IN2(n5414), .Q(WX9082) );
  XOR2X1 U6618 ( .IN1(CRC_OUT_3_29), .IN2(n4595), .Q(n6029) );
  AND2X1 U6619 ( .IN1(n6030), .IN2(n5414), .Q(WX9080) );
  XOR2X1 U6620 ( .IN1(CRC_OUT_3_28), .IN2(n4596), .Q(n6030) );
  AND2X1 U6621 ( .IN1(n6031), .IN2(n5414), .Q(WX9078) );
  XOR2X1 U6622 ( .IN1(CRC_OUT_3_27), .IN2(n4597), .Q(n6031) );
  AND2X1 U6623 ( .IN1(n6032), .IN2(n5414), .Q(WX9076) );
  XOR2X1 U6624 ( .IN1(CRC_OUT_3_26), .IN2(n4598), .Q(n6032) );
  AND2X1 U6625 ( .IN1(n6033), .IN2(n5414), .Q(WX9074) );
  XOR2X1 U6626 ( .IN1(test_so74), .IN2(DFF_1337_n1), .Q(n6033) );
  AND2X1 U6627 ( .IN1(n6034), .IN2(n5414), .Q(WX9072) );
  XOR2X1 U6628 ( .IN1(test_so77), .IN2(n4599), .Q(n6034) );
  AND2X1 U6629 ( .IN1(n6035), .IN2(n5414), .Q(WX9070) );
  XOR2X1 U6630 ( .IN1(CRC_OUT_3_23), .IN2(n4600), .Q(n6035) );
  AND2X1 U6631 ( .IN1(n6036), .IN2(n5413), .Q(WX9068) );
  XOR2X1 U6632 ( .IN1(CRC_OUT_3_22), .IN2(n4601), .Q(n6036) );
  AND2X1 U6633 ( .IN1(n6037), .IN2(n5413), .Q(WX9066) );
  XOR2X1 U6634 ( .IN1(CRC_OUT_3_21), .IN2(n4602), .Q(n6037) );
  AND2X1 U6635 ( .IN1(n6038), .IN2(n5413), .Q(WX9064) );
  XOR2X1 U6636 ( .IN1(CRC_OUT_3_20), .IN2(n4603), .Q(n6038) );
  AND2X1 U6637 ( .IN1(n6039), .IN2(n5413), .Q(WX9062) );
  XOR2X1 U6638 ( .IN1(CRC_OUT_3_19), .IN2(n4604), .Q(n6039) );
  AND2X1 U6639 ( .IN1(n6040), .IN2(n5413), .Q(WX9060) );
  XOR2X1 U6640 ( .IN1(CRC_OUT_3_18), .IN2(n4605), .Q(n6040) );
  AND2X1 U6641 ( .IN1(n6041), .IN2(n5413), .Q(WX9058) );
  XOR2X1 U6642 ( .IN1(CRC_OUT_3_17), .IN2(n4606), .Q(n6041) );
  AND2X1 U6643 ( .IN1(n6042), .IN2(n5413), .Q(WX9056) );
  XOR2X1 U6644 ( .IN1(CRC_OUT_3_16), .IN2(n4607), .Q(n6042) );
  AND2X1 U6645 ( .IN1(n6043), .IN2(n5413), .Q(WX9054) );
  XOR2X1 U6646 ( .IN1(DFF_1327_n1), .IN2(n6044), .Q(n6043) );
  XOR2X1 U6647 ( .IN1(n4519), .IN2(DFF_1343_n1), .Q(n6044) );
  AND2X1 U6648 ( .IN1(n6045), .IN2(n5413), .Q(WX9052) );
  XOR2X1 U6649 ( .IN1(CRC_OUT_3_14), .IN2(n4608), .Q(n6045) );
  AND2X1 U6650 ( .IN1(n6046), .IN2(n5412), .Q(WX9050) );
  XOR2X1 U6651 ( .IN1(CRC_OUT_3_13), .IN2(n4609), .Q(n6046) );
  AND2X1 U6652 ( .IN1(n6047), .IN2(n5412), .Q(WX9048) );
  XOR2X1 U6653 ( .IN1(CRC_OUT_3_12), .IN2(n4610), .Q(n6047) );
  AND2X1 U6654 ( .IN1(n6048), .IN2(n5412), .Q(WX9046) );
  XOR2X1 U6655 ( .IN1(CRC_OUT_3_11), .IN2(n4611), .Q(n6048) );
  AND2X1 U6656 ( .IN1(n6049), .IN2(n5412), .Q(WX9044) );
  XOR2X1 U6657 ( .IN1(DFF_1322_n1), .IN2(n6050), .Q(n6049) );
  XOR2X1 U6658 ( .IN1(n4520), .IN2(DFF_1343_n1), .Q(n6050) );
  AND2X1 U6659 ( .IN1(n6051), .IN2(n5412), .Q(WX9042) );
  XOR2X1 U6660 ( .IN1(CRC_OUT_3_9), .IN2(n4612), .Q(n6051) );
  AND2X1 U6661 ( .IN1(n6052), .IN2(n5412), .Q(WX9040) );
  XOR2X1 U6662 ( .IN1(test_so75), .IN2(DFF_1320_n1), .Q(n6052) );
  AND2X1 U6663 ( .IN1(n6053), .IN2(n5412), .Q(WX9038) );
  XOR2X1 U6664 ( .IN1(test_so76), .IN2(n4613), .Q(n6053) );
  AND2X1 U6665 ( .IN1(n6054), .IN2(n5412), .Q(WX9036) );
  XOR2X1 U6666 ( .IN1(CRC_OUT_3_6), .IN2(n4614), .Q(n6054) );
  AND2X1 U6667 ( .IN1(n6055), .IN2(n5412), .Q(WX9034) );
  XOR2X1 U6668 ( .IN1(CRC_OUT_3_5), .IN2(n4615), .Q(n6055) );
  AND2X1 U6669 ( .IN1(n6056), .IN2(n5411), .Q(WX9032) );
  XOR2X1 U6670 ( .IN1(CRC_OUT_3_4), .IN2(n4616), .Q(n6056) );
  AND2X1 U6671 ( .IN1(n6057), .IN2(n5411), .Q(WX9030) );
  XOR2X1 U6672 ( .IN1(DFF_1315_n1), .IN2(n6058), .Q(n6057) );
  XOR2X1 U6673 ( .IN1(n4521), .IN2(DFF_1343_n1), .Q(n6058) );
  AND2X1 U6674 ( .IN1(n6059), .IN2(n5411), .Q(WX9028) );
  XOR2X1 U6675 ( .IN1(CRC_OUT_3_2), .IN2(n4617), .Q(n6059) );
  AND2X1 U6676 ( .IN1(n6060), .IN2(n5411), .Q(WX9026) );
  XOR2X1 U6677 ( .IN1(CRC_OUT_3_1), .IN2(n4618), .Q(n6060) );
  AND2X1 U6678 ( .IN1(n6061), .IN2(n5411), .Q(WX9024) );
  XOR2X1 U6679 ( .IN1(CRC_OUT_3_0), .IN2(n4619), .Q(n6061) );
  AND2X1 U6680 ( .IN1(n6062), .IN2(n5411), .Q(WX9022) );
  XOR2X1 U6681 ( .IN1(n4536), .IN2(CRC_OUT_3_31), .Q(n6062) );
  INVX0 U6682 ( .INP(n6063), .ZN(WX8496) );
  OR2X1 U6683 ( .IN1(n5470), .IN2(n9569), .Q(n6063) );
  INVX0 U6684 ( .INP(n6064), .ZN(WX8494) );
  OR2X1 U6685 ( .IN1(n5470), .IN2(n9570), .Q(n6064) );
  INVX0 U6686 ( .INP(n6065), .ZN(WX8492) );
  OR2X1 U6687 ( .IN1(n5470), .IN2(n9571), .Q(n6065) );
  INVX0 U6688 ( .INP(n6066), .ZN(WX8490) );
  OR2X1 U6689 ( .IN1(n5470), .IN2(n9572), .Q(n6066) );
  INVX0 U6690 ( .INP(n6067), .ZN(WX8488) );
  OR2X1 U6691 ( .IN1(n5470), .IN2(n9573), .Q(n6067) );
  INVX0 U6692 ( .INP(n6068), .ZN(WX8486) );
  OR2X1 U6693 ( .IN1(n5470), .IN2(n9574), .Q(n6068) );
  INVX0 U6694 ( .INP(n6069), .ZN(WX8484) );
  OR2X1 U6695 ( .IN1(n5470), .IN2(n9575), .Q(n6069) );
  INVX0 U6696 ( .INP(n6070), .ZN(WX8482) );
  OR2X1 U6697 ( .IN1(n5469), .IN2(n9576), .Q(n6070) );
  INVX0 U6698 ( .INP(n6071), .ZN(WX8480) );
  OR2X1 U6699 ( .IN1(n5469), .IN2(n9577), .Q(n6071) );
  INVX0 U6700 ( .INP(n6072), .ZN(WX8478) );
  OR2X1 U6701 ( .IN1(n5469), .IN2(n9578), .Q(n6072) );
  INVX0 U6702 ( .INP(n6073), .ZN(WX8476) );
  OR2X1 U6703 ( .IN1(n5469), .IN2(n9579), .Q(n6073) );
  INVX0 U6704 ( .INP(n6074), .ZN(WX8474) );
  OR2X1 U6705 ( .IN1(n5469), .IN2(n9580), .Q(n6074) );
  INVX0 U6706 ( .INP(n6075), .ZN(WX8472) );
  OR2X1 U6707 ( .IN1(n5469), .IN2(n9581), .Q(n6075) );
  INVX0 U6708 ( .INP(n6076), .ZN(WX8470) );
  OR2X1 U6709 ( .IN1(n5469), .IN2(n9584), .Q(n6076) );
  INVX0 U6710 ( .INP(n6077), .ZN(WX8468) );
  OR2X1 U6711 ( .IN1(n5469), .IN2(n9585), .Q(n6077) );
  INVX0 U6712 ( .INP(n6078), .ZN(WX8466) );
  OR2X1 U6713 ( .IN1(n5469), .IN2(n9588), .Q(n6078) );
  OR2X1 U6714 ( .IN1(n6079), .IN2(n6080), .Q(WX8464) );
  OR2X1 U6715 ( .IN1(n6081), .IN2(n6082), .Q(n6080) );
  AND2X1 U6716 ( .IN1(n4900), .IN2(CRC_OUT_3_0), .Q(n6082) );
  AND2X1 U6717 ( .IN1(n374), .IN2(n4881), .Q(n6081) );
  INVX0 U6718 ( .INP(n6083), .ZN(n374) );
  OR2X1 U6719 ( .IN1(n5469), .IN2(n3848), .Q(n6083) );
  OR2X1 U6720 ( .IN1(n6084), .IN2(n6085), .Q(n6079) );
  AND2X1 U6721 ( .IN1(n4843), .IN2(n6086), .Q(n6085) );
  AND2X1 U6722 ( .IN1(n4931), .IN2(n5749), .Q(n6084) );
  XNOR2X1 U6723 ( .IN1(n6087), .IN2(n6088), .Q(n5749) );
  XOR2X1 U6724 ( .IN1(n9518), .IN2(n4535), .Q(n6088) );
  XOR2X1 U6725 ( .IN1(WX9758), .IN2(n4309), .Q(n6087) );
  OR2X1 U6726 ( .IN1(n6089), .IN2(n6090), .Q(WX8462) );
  OR2X1 U6727 ( .IN1(n6091), .IN2(n6092), .Q(n6090) );
  AND2X1 U6728 ( .IN1(n4900), .IN2(CRC_OUT_3_1), .Q(n6092) );
  AND2X1 U6729 ( .IN1(n373), .IN2(n4881), .Q(n6091) );
  INVX0 U6730 ( .INP(n6093), .ZN(n373) );
  OR2X1 U6731 ( .IN1(n5469), .IN2(n3849), .Q(n6093) );
  OR2X1 U6732 ( .IN1(n6094), .IN2(n6095), .Q(n6089) );
  AND2X1 U6733 ( .IN1(n4843), .IN2(n6096), .Q(n6095) );
  AND2X1 U6734 ( .IN1(n5758), .IN2(n4922), .Q(n6094) );
  XOR2X1 U6735 ( .IN1(n6097), .IN2(n6098), .Q(n5758) );
  XOR2X1 U6736 ( .IN1(test_so83), .IN2(n9519), .Q(n6098) );
  XOR2X1 U6737 ( .IN1(WX9756), .IN2(n4593), .Q(n6097) );
  OR2X1 U6738 ( .IN1(n6099), .IN2(n6100), .Q(WX8460) );
  OR2X1 U6739 ( .IN1(n6101), .IN2(n6102), .Q(n6100) );
  AND2X1 U6740 ( .IN1(n4900), .IN2(CRC_OUT_3_2), .Q(n6102) );
  AND2X1 U6741 ( .IN1(n372), .IN2(n4881), .Q(n6101) );
  INVX0 U6742 ( .INP(n6103), .ZN(n372) );
  OR2X1 U6743 ( .IN1(n5469), .IN2(n3850), .Q(n6103) );
  OR2X1 U6744 ( .IN1(n6104), .IN2(n6105), .Q(n6099) );
  AND2X1 U6745 ( .IN1(n4843), .IN2(n6106), .Q(n6105) );
  AND2X1 U6746 ( .IN1(n4931), .IN2(n5767), .Q(n6104) );
  XNOR2X1 U6747 ( .IN1(n6107), .IN2(n6108), .Q(n5767) );
  XOR2X1 U6748 ( .IN1(n9520), .IN2(n4592), .Q(n6108) );
  XOR2X1 U6749 ( .IN1(WX9754), .IN2(n4312), .Q(n6107) );
  OR2X1 U6750 ( .IN1(n6109), .IN2(n6110), .Q(WX8458) );
  OR2X1 U6751 ( .IN1(n6111), .IN2(n6112), .Q(n6110) );
  AND2X1 U6752 ( .IN1(n4901), .IN2(CRC_OUT_3_3), .Q(n6112) );
  AND2X1 U6753 ( .IN1(n371), .IN2(n4881), .Q(n6111) );
  INVX0 U6754 ( .INP(n6113), .ZN(n371) );
  OR2X1 U6755 ( .IN1(n5469), .IN2(n3851), .Q(n6113) );
  OR2X1 U6756 ( .IN1(n6114), .IN2(n6115), .Q(n6109) );
  AND2X1 U6757 ( .IN1(n4843), .IN2(n6116), .Q(n6115) );
  AND2X1 U6758 ( .IN1(n5776), .IN2(n4921), .Q(n6114) );
  XOR2X1 U6759 ( .IN1(n6117), .IN2(n6118), .Q(n5776) );
  XOR2X1 U6760 ( .IN1(test_so81), .IN2(n9521), .Q(n6118) );
  XOR2X1 U6761 ( .IN1(WX9880), .IN2(n4591), .Q(n6117) );
  OR2X1 U6762 ( .IN1(n6119), .IN2(n6120), .Q(WX8456) );
  OR2X1 U6763 ( .IN1(n6121), .IN2(n6122), .Q(n6120) );
  AND2X1 U6764 ( .IN1(n4901), .IN2(CRC_OUT_3_4), .Q(n6122) );
  AND2X1 U6765 ( .IN1(n370), .IN2(n4881), .Q(n6121) );
  INVX0 U6766 ( .INP(n6123), .ZN(n370) );
  OR2X1 U6767 ( .IN1(n5468), .IN2(n3852), .Q(n6123) );
  OR2X1 U6768 ( .IN1(n6124), .IN2(n6125), .Q(n6119) );
  AND2X1 U6769 ( .IN1(n4843), .IN2(n6126), .Q(n6125) );
  AND2X1 U6770 ( .IN1(n4932), .IN2(n5785), .Q(n6124) );
  XNOR2X1 U6771 ( .IN1(n6127), .IN2(n6128), .Q(n5785) );
  XOR2X1 U6772 ( .IN1(n9522), .IN2(n4518), .Q(n6128) );
  XOR2X1 U6773 ( .IN1(WX9750), .IN2(n4315), .Q(n6127) );
  OR2X1 U6774 ( .IN1(n6129), .IN2(n6130), .Q(WX8454) );
  OR2X1 U6775 ( .IN1(n6131), .IN2(n6132), .Q(n6130) );
  AND2X1 U6776 ( .IN1(n4901), .IN2(CRC_OUT_3_5), .Q(n6132) );
  AND2X1 U6777 ( .IN1(n369), .IN2(n4881), .Q(n6131) );
  INVX0 U6778 ( .INP(n6133), .ZN(n369) );
  OR2X1 U6779 ( .IN1(n5468), .IN2(n3853), .Q(n6133) );
  OR2X1 U6780 ( .IN1(n6134), .IN2(n6135), .Q(n6129) );
  AND2X1 U6781 ( .IN1(n4843), .IN2(n6136), .Q(n6135) );
  AND2X1 U6782 ( .IN1(n4932), .IN2(n5794), .Q(n6134) );
  XNOR2X1 U6783 ( .IN1(n6137), .IN2(n6138), .Q(n5794) );
  XOR2X1 U6784 ( .IN1(n9523), .IN2(n4590), .Q(n6138) );
  XOR2X1 U6785 ( .IN1(WX9748), .IN2(n4317), .Q(n6137) );
  OR2X1 U6786 ( .IN1(n6139), .IN2(n6140), .Q(WX8452) );
  OR2X1 U6787 ( .IN1(n6141), .IN2(n6142), .Q(n6140) );
  AND2X1 U6788 ( .IN1(n4901), .IN2(CRC_OUT_3_6), .Q(n6142) );
  AND2X1 U6789 ( .IN1(n368), .IN2(n4881), .Q(n6141) );
  INVX0 U6790 ( .INP(n6143), .ZN(n368) );
  OR2X1 U6791 ( .IN1(n5468), .IN2(n3854), .Q(n6143) );
  OR2X1 U6792 ( .IN1(n6144), .IN2(n6145), .Q(n6139) );
  AND2X1 U6793 ( .IN1(n4843), .IN2(n6146), .Q(n6145) );
  AND2X1 U6794 ( .IN1(n4932), .IN2(n5803), .Q(n6144) );
  XNOR2X1 U6795 ( .IN1(n6147), .IN2(n6148), .Q(n5803) );
  XOR2X1 U6796 ( .IN1(n9524), .IN2(n4589), .Q(n6148) );
  XOR2X1 U6797 ( .IN1(WX9746), .IN2(n4319), .Q(n6147) );
  OR2X1 U6798 ( .IN1(n6149), .IN2(n6150), .Q(WX8450) );
  OR2X1 U6799 ( .IN1(n6151), .IN2(n6152), .Q(n6150) );
  AND2X1 U6800 ( .IN1(test_so76), .IN2(n4888), .Q(n6152) );
  AND2X1 U6801 ( .IN1(n367), .IN2(n4881), .Q(n6151) );
  INVX0 U6802 ( .INP(n6153), .ZN(n367) );
  OR2X1 U6803 ( .IN1(n5468), .IN2(n3855), .Q(n6153) );
  OR2X1 U6804 ( .IN1(n6154), .IN2(n6155), .Q(n6149) );
  AND2X1 U6805 ( .IN1(n4843), .IN2(n6156), .Q(n6155) );
  AND2X1 U6806 ( .IN1(n4932), .IN2(n5812), .Q(n6154) );
  XNOR2X1 U6807 ( .IN1(n6157), .IN2(n6158), .Q(n5812) );
  XOR2X1 U6808 ( .IN1(n9525), .IN2(n4588), .Q(n6158) );
  XOR2X1 U6809 ( .IN1(WX9744), .IN2(n4321), .Q(n6157) );
  OR2X1 U6810 ( .IN1(n6159), .IN2(n6160), .Q(WX8448) );
  OR2X1 U6811 ( .IN1(n6161), .IN2(n6162), .Q(n6160) );
  AND2X1 U6812 ( .IN1(n4901), .IN2(CRC_OUT_3_8), .Q(n6162) );
  AND2X1 U6813 ( .IN1(n366), .IN2(n4880), .Q(n6161) );
  INVX0 U6814 ( .INP(n6163), .ZN(n366) );
  OR2X1 U6815 ( .IN1(n5468), .IN2(n3856), .Q(n6163) );
  OR2X1 U6816 ( .IN1(n6164), .IN2(n6165), .Q(n6159) );
  AND2X1 U6817 ( .IN1(n4843), .IN2(n6166), .Q(n6165) );
  AND2X1 U6818 ( .IN1(n4932), .IN2(n5821), .Q(n6164) );
  XNOR2X1 U6819 ( .IN1(n6167), .IN2(n6168), .Q(n5821) );
  XOR2X1 U6820 ( .IN1(n9526), .IN2(n4587), .Q(n6168) );
  XOR2X1 U6821 ( .IN1(WX9742), .IN2(n4323), .Q(n6167) );
  OR2X1 U6822 ( .IN1(n6169), .IN2(n6170), .Q(WX8446) );
  OR2X1 U6823 ( .IN1(n6171), .IN2(n6172), .Q(n6170) );
  AND2X1 U6824 ( .IN1(n4901), .IN2(CRC_OUT_3_9), .Q(n6172) );
  AND2X1 U6825 ( .IN1(n365), .IN2(n4880), .Q(n6171) );
  INVX0 U6826 ( .INP(n6173), .ZN(n365) );
  OR2X1 U6827 ( .IN1(n5468), .IN2(n3857), .Q(n6173) );
  OR2X1 U6828 ( .IN1(n6174), .IN2(n6175), .Q(n6169) );
  AND2X1 U6829 ( .IN1(n6176), .IN2(n4837), .Q(n6175) );
  AND2X1 U6830 ( .IN1(n4932), .IN2(n5830), .Q(n6174) );
  XNOR2X1 U6831 ( .IN1(n6177), .IN2(n6178), .Q(n5830) );
  XOR2X1 U6832 ( .IN1(n9527), .IN2(n4586), .Q(n6178) );
  XOR2X1 U6833 ( .IN1(WX9740), .IN2(n4325), .Q(n6177) );
  OR2X1 U6834 ( .IN1(n6179), .IN2(n6180), .Q(WX8444) );
  OR2X1 U6835 ( .IN1(n6181), .IN2(n6182), .Q(n6180) );
  AND2X1 U6836 ( .IN1(n4901), .IN2(CRC_OUT_3_10), .Q(n6182) );
  AND2X1 U6837 ( .IN1(n364), .IN2(n4880), .Q(n6181) );
  INVX0 U6838 ( .INP(n6183), .ZN(n364) );
  OR2X1 U6839 ( .IN1(n5468), .IN2(n3858), .Q(n6183) );
  OR2X1 U6840 ( .IN1(n6184), .IN2(n6185), .Q(n6179) );
  AND2X1 U6841 ( .IN1(n4843), .IN2(n6186), .Q(n6185) );
  AND2X1 U6842 ( .IN1(n4932), .IN2(n5839), .Q(n6184) );
  XNOR2X1 U6843 ( .IN1(n6187), .IN2(n6188), .Q(n5839) );
  XOR2X1 U6844 ( .IN1(n9528), .IN2(n4585), .Q(n6188) );
  XOR2X1 U6845 ( .IN1(WX9738), .IN2(n4327), .Q(n6187) );
  OR2X1 U6846 ( .IN1(n6189), .IN2(n6190), .Q(WX8442) );
  OR2X1 U6847 ( .IN1(n6191), .IN2(n6192), .Q(n6190) );
  AND2X1 U6848 ( .IN1(n4901), .IN2(CRC_OUT_3_11), .Q(n6192) );
  AND2X1 U6849 ( .IN1(n363), .IN2(n4880), .Q(n6191) );
  INVX0 U6850 ( .INP(n6193), .ZN(n363) );
  OR2X1 U6851 ( .IN1(n5468), .IN2(n3859), .Q(n6193) );
  OR2X1 U6852 ( .IN1(n6194), .IN2(n6195), .Q(n6189) );
  AND2X1 U6853 ( .IN1(n6196), .IN2(n4837), .Q(n6195) );
  AND2X1 U6854 ( .IN1(n4932), .IN2(n5848), .Q(n6194) );
  XNOR2X1 U6855 ( .IN1(n6197), .IN2(n6198), .Q(n5848) );
  XOR2X1 U6856 ( .IN1(n9529), .IN2(n4517), .Q(n6198) );
  XOR2X1 U6857 ( .IN1(WX9736), .IN2(n4329), .Q(n6197) );
  OR2X1 U6858 ( .IN1(n6199), .IN2(n6200), .Q(WX8440) );
  OR2X1 U6859 ( .IN1(n6201), .IN2(n6202), .Q(n6200) );
  AND2X1 U6860 ( .IN1(n4901), .IN2(CRC_OUT_3_12), .Q(n6202) );
  AND2X1 U6861 ( .IN1(n362), .IN2(n4880), .Q(n6201) );
  INVX0 U6862 ( .INP(n6203), .ZN(n362) );
  OR2X1 U6863 ( .IN1(n5468), .IN2(n3860), .Q(n6203) );
  OR2X1 U6864 ( .IN1(n6204), .IN2(n6205), .Q(n6199) );
  AND2X1 U6865 ( .IN1(n4843), .IN2(n6206), .Q(n6205) );
  AND2X1 U6866 ( .IN1(n4932), .IN2(n5857), .Q(n6204) );
  XNOR2X1 U6867 ( .IN1(n6207), .IN2(n6208), .Q(n5857) );
  XOR2X1 U6868 ( .IN1(n9530), .IN2(n4584), .Q(n6208) );
  XOR2X1 U6869 ( .IN1(WX9734), .IN2(n4331), .Q(n6207) );
  OR2X1 U6870 ( .IN1(n6209), .IN2(n6210), .Q(WX8438) );
  OR2X1 U6871 ( .IN1(n6211), .IN2(n6212), .Q(n6210) );
  AND2X1 U6872 ( .IN1(n4901), .IN2(CRC_OUT_3_13), .Q(n6212) );
  AND2X1 U6873 ( .IN1(n361), .IN2(n4880), .Q(n6211) );
  INVX0 U6874 ( .INP(n6213), .ZN(n361) );
  OR2X1 U6875 ( .IN1(n5468), .IN2(n3861), .Q(n6213) );
  OR2X1 U6876 ( .IN1(n6214), .IN2(n6215), .Q(n6209) );
  AND2X1 U6877 ( .IN1(n6216), .IN2(n4837), .Q(n6215) );
  AND2X1 U6878 ( .IN1(n4932), .IN2(n5866), .Q(n6214) );
  XNOR2X1 U6879 ( .IN1(n6217), .IN2(n6218), .Q(n5866) );
  XOR2X1 U6880 ( .IN1(n9531), .IN2(n4583), .Q(n6218) );
  XOR2X1 U6881 ( .IN1(WX9732), .IN2(n4333), .Q(n6217) );
  OR2X1 U6882 ( .IN1(n6219), .IN2(n6220), .Q(WX8436) );
  OR2X1 U6883 ( .IN1(n6221), .IN2(n6222), .Q(n6220) );
  AND2X1 U6884 ( .IN1(n4901), .IN2(CRC_OUT_3_14), .Q(n6222) );
  AND2X1 U6885 ( .IN1(n360), .IN2(n4880), .Q(n6221) );
  INVX0 U6886 ( .INP(n6223), .ZN(n360) );
  OR2X1 U6887 ( .IN1(n5468), .IN2(n3862), .Q(n6223) );
  OR2X1 U6888 ( .IN1(n6224), .IN2(n6225), .Q(n6219) );
  AND2X1 U6889 ( .IN1(n4843), .IN2(n6226), .Q(n6225) );
  AND2X1 U6890 ( .IN1(n5875), .IN2(n4921), .Q(n6224) );
  XOR2X1 U6891 ( .IN1(n6227), .IN2(n6228), .Q(n5875) );
  XOR2X1 U6892 ( .IN1(test_so86), .IN2(n9532), .Q(n6228) );
  XOR2X1 U6893 ( .IN1(WX9730), .IN2(n4335), .Q(n6227) );
  OR2X1 U6894 ( .IN1(n6229), .IN2(n6230), .Q(WX8434) );
  OR2X1 U6895 ( .IN1(n6231), .IN2(n6232), .Q(n6230) );
  AND2X1 U6896 ( .IN1(n4901), .IN2(CRC_OUT_3_15), .Q(n6232) );
  AND2X1 U6897 ( .IN1(n359), .IN2(n4880), .Q(n6231) );
  INVX0 U6898 ( .INP(n6233), .ZN(n359) );
  OR2X1 U6899 ( .IN1(n5468), .IN2(n3863), .Q(n6233) );
  OR2X1 U6900 ( .IN1(n6234), .IN2(n6235), .Q(n6229) );
  AND2X1 U6901 ( .IN1(n6236), .IN2(n4836), .Q(n6235) );
  AND2X1 U6902 ( .IN1(n4932), .IN2(n5884), .Q(n6234) );
  XNOR2X1 U6903 ( .IN1(n6237), .IN2(n6238), .Q(n5884) );
  XOR2X1 U6904 ( .IN1(n9533), .IN2(n4582), .Q(n6238) );
  XOR2X1 U6905 ( .IN1(WX9728), .IN2(n4337), .Q(n6237) );
  OR2X1 U6906 ( .IN1(n6239), .IN2(n6240), .Q(WX8432) );
  OR2X1 U6907 ( .IN1(n6241), .IN2(n6242), .Q(n6240) );
  AND2X1 U6908 ( .IN1(n4901), .IN2(CRC_OUT_3_16), .Q(n6242) );
  AND2X1 U6909 ( .IN1(n358), .IN2(n4880), .Q(n6241) );
  INVX0 U6910 ( .INP(n6243), .ZN(n358) );
  OR2X1 U6911 ( .IN1(n5468), .IN2(n3864), .Q(n6243) );
  OR2X1 U6912 ( .IN1(n6244), .IN2(n6245), .Q(n6239) );
  AND2X1 U6913 ( .IN1(n4843), .IN2(n6246), .Q(n6245) );
  AND2X1 U6914 ( .IN1(n5893), .IN2(n4920), .Q(n6244) );
  XOR2X1 U6915 ( .IN1(n6247), .IN2(n6248), .Q(n5893) );
  XOR2X1 U6916 ( .IN1(n4516), .IN2(n5378), .Q(n6248) );
  XOR2X1 U6917 ( .IN1(n6249), .IN2(n9536), .Q(n6247) );
  XOR2X1 U6918 ( .IN1(n9535), .IN2(n9534), .Q(n6249) );
  OR2X1 U6919 ( .IN1(n6250), .IN2(n6251), .Q(WX8430) );
  OR2X1 U6920 ( .IN1(n6252), .IN2(n6253), .Q(n6251) );
  AND2X1 U6921 ( .IN1(n4902), .IN2(CRC_OUT_3_17), .Q(n6253) );
  AND2X1 U6922 ( .IN1(n357), .IN2(n4880), .Q(n6252) );
  INVX0 U6923 ( .INP(n6254), .ZN(n357) );
  OR2X1 U6924 ( .IN1(n5467), .IN2(n3865), .Q(n6254) );
  OR2X1 U6925 ( .IN1(n6255), .IN2(n6256), .Q(n6250) );
  AND2X1 U6926 ( .IN1(n4842), .IN2(n6257), .Q(n6256) );
  AND2X1 U6927 ( .IN1(n4932), .IN2(n5902), .Q(n6255) );
  XNOR2X1 U6928 ( .IN1(n6258), .IN2(n6259), .Q(n5902) );
  XOR2X1 U6929 ( .IN1(n4186), .IN2(n5389), .Q(n6259) );
  XOR2X1 U6930 ( .IN1(n6260), .IN2(n4581), .Q(n6258) );
  XOR2X1 U6931 ( .IN1(WX9852), .IN2(n9537), .Q(n6260) );
  OR2X1 U6932 ( .IN1(n6261), .IN2(n6262), .Q(WX8428) );
  OR2X1 U6933 ( .IN1(n6263), .IN2(n6264), .Q(n6262) );
  AND2X1 U6934 ( .IN1(n4902), .IN2(CRC_OUT_3_18), .Q(n6264) );
  AND2X1 U6935 ( .IN1(WX8266), .IN2(n4880), .Q(n6263) );
  OR2X1 U6936 ( .IN1(n6265), .IN2(n6266), .Q(n6261) );
  AND2X1 U6937 ( .IN1(n4842), .IN2(n6267), .Q(n6266) );
  AND2X1 U6938 ( .IN1(n5911), .IN2(n4920), .Q(n6265) );
  XOR2X1 U6939 ( .IN1(n6268), .IN2(n6269), .Q(n5911) );
  XOR2X1 U6940 ( .IN1(n4580), .IN2(n5389), .Q(n6269) );
  XOR2X1 U6941 ( .IN1(n6270), .IN2(n9540), .Q(n6268) );
  XOR2X1 U6942 ( .IN1(n9539), .IN2(n9538), .Q(n6270) );
  OR2X1 U6943 ( .IN1(n6271), .IN2(n6272), .Q(WX8426) );
  OR2X1 U6944 ( .IN1(n6273), .IN2(n6274), .Q(n6272) );
  AND2X1 U6945 ( .IN1(n4902), .IN2(CRC_OUT_3_19), .Q(n6274) );
  AND2X1 U6946 ( .IN1(n355), .IN2(n4880), .Q(n6273) );
  INVX0 U6947 ( .INP(n6275), .ZN(n355) );
  OR2X1 U6948 ( .IN1(n5467), .IN2(n3867), .Q(n6275) );
  OR2X1 U6949 ( .IN1(n6276), .IN2(n6277), .Q(n6271) );
  AND2X1 U6950 ( .IN1(n4842), .IN2(n6278), .Q(n6277) );
  AND2X1 U6951 ( .IN1(n4932), .IN2(n5920), .Q(n6276) );
  XNOR2X1 U6952 ( .IN1(n6279), .IN2(n6280), .Q(n5920) );
  XOR2X1 U6953 ( .IN1(n4187), .IN2(n5389), .Q(n6280) );
  XOR2X1 U6954 ( .IN1(n6281), .IN2(n4579), .Q(n6279) );
  XOR2X1 U6955 ( .IN1(WX9848), .IN2(n9541), .Q(n6281) );
  OR2X1 U6956 ( .IN1(n6282), .IN2(n6283), .Q(WX8424) );
  OR2X1 U6957 ( .IN1(n6284), .IN2(n6285), .Q(n6283) );
  AND2X1 U6958 ( .IN1(n4902), .IN2(CRC_OUT_3_20), .Q(n6285) );
  AND2X1 U6959 ( .IN1(n354), .IN2(n4879), .Q(n6284) );
  INVX0 U6960 ( .INP(n6286), .ZN(n354) );
  OR2X1 U6961 ( .IN1(n5467), .IN2(n3868), .Q(n6286) );
  OR2X1 U6962 ( .IN1(n6287), .IN2(n6288), .Q(n6282) );
  AND2X1 U6963 ( .IN1(n4842), .IN2(n6289), .Q(n6288) );
  AND2X1 U6964 ( .IN1(n5929), .IN2(n4920), .Q(n6287) );
  XOR2X1 U6965 ( .IN1(n6290), .IN2(n6291), .Q(n5929) );
  XOR2X1 U6966 ( .IN1(n4188), .IN2(n5389), .Q(n6291) );
  XOR2X1 U6967 ( .IN1(n6292), .IN2(n4578), .Q(n6290) );
  XOR2X1 U6968 ( .IN1(WX9782), .IN2(test_so80), .Q(n6292) );
  OR2X1 U6969 ( .IN1(n6293), .IN2(n6294), .Q(WX8422) );
  OR2X1 U6970 ( .IN1(n6295), .IN2(n6296), .Q(n6294) );
  AND2X1 U6971 ( .IN1(n4902), .IN2(CRC_OUT_3_21), .Q(n6296) );
  AND2X1 U6972 ( .IN1(n353), .IN2(n4879), .Q(n6295) );
  INVX0 U6973 ( .INP(n6297), .ZN(n353) );
  OR2X1 U6974 ( .IN1(n5467), .IN2(n3869), .Q(n6297) );
  OR2X1 U6975 ( .IN1(n6298), .IN2(n6299), .Q(n6293) );
  AND2X1 U6976 ( .IN1(n4842), .IN2(n6300), .Q(n6299) );
  AND2X1 U6977 ( .IN1(n4933), .IN2(n5938), .Q(n6298) );
  XNOR2X1 U6978 ( .IN1(n6301), .IN2(n6302), .Q(n5938) );
  XOR2X1 U6979 ( .IN1(n4189), .IN2(n5389), .Q(n6302) );
  XOR2X1 U6980 ( .IN1(n6303), .IN2(n4577), .Q(n6301) );
  XOR2X1 U6981 ( .IN1(WX9844), .IN2(n9542), .Q(n6303) );
  OR2X1 U6982 ( .IN1(n6304), .IN2(n6305), .Q(WX8420) );
  OR2X1 U6983 ( .IN1(n6306), .IN2(n6307), .Q(n6305) );
  AND2X1 U6984 ( .IN1(n4902), .IN2(CRC_OUT_3_22), .Q(n6307) );
  AND2X1 U6985 ( .IN1(n352), .IN2(n4879), .Q(n6306) );
  INVX0 U6986 ( .INP(n6308), .ZN(n352) );
  OR2X1 U6987 ( .IN1(n5467), .IN2(n3870), .Q(n6308) );
  OR2X1 U6988 ( .IN1(n6309), .IN2(n6310), .Q(n6304) );
  AND2X1 U6989 ( .IN1(n4842), .IN2(n6311), .Q(n6310) );
  AND2X1 U6990 ( .IN1(n4933), .IN2(n5947), .Q(n6309) );
  XNOR2X1 U6991 ( .IN1(n6312), .IN2(n6313), .Q(n5947) );
  XOR2X1 U6992 ( .IN1(n4190), .IN2(n5389), .Q(n6313) );
  XOR2X1 U6993 ( .IN1(n6314), .IN2(n4576), .Q(n6312) );
  XOR2X1 U6994 ( .IN1(WX9842), .IN2(n9543), .Q(n6314) );
  OR2X1 U6995 ( .IN1(n6315), .IN2(n6316), .Q(WX8418) );
  OR2X1 U6996 ( .IN1(n6317), .IN2(n6318), .Q(n6316) );
  AND2X1 U6997 ( .IN1(n4902), .IN2(CRC_OUT_3_23), .Q(n6318) );
  AND2X1 U6998 ( .IN1(n351), .IN2(n4879), .Q(n6317) );
  INVX0 U6999 ( .INP(n6319), .ZN(n351) );
  OR2X1 U7000 ( .IN1(n5467), .IN2(n3871), .Q(n6319) );
  OR2X1 U7001 ( .IN1(n6320), .IN2(n6321), .Q(n6315) );
  AND2X1 U7002 ( .IN1(n4842), .IN2(n6322), .Q(n6321) );
  AND2X1 U7003 ( .IN1(n4933), .IN2(n5956), .Q(n6320) );
  XNOR2X1 U7004 ( .IN1(n6323), .IN2(n6324), .Q(n5956) );
  XOR2X1 U7005 ( .IN1(n4191), .IN2(n5389), .Q(n6324) );
  XOR2X1 U7006 ( .IN1(n6325), .IN2(n4575), .Q(n6323) );
  XOR2X1 U7007 ( .IN1(WX9840), .IN2(n9544), .Q(n6325) );
  OR2X1 U7008 ( .IN1(n6326), .IN2(n6327), .Q(WX8416) );
  OR2X1 U7009 ( .IN1(n6328), .IN2(n6329), .Q(n6327) );
  AND2X1 U7010 ( .IN1(test_so77), .IN2(n4887), .Q(n6329) );
  AND2X1 U7011 ( .IN1(n350), .IN2(n4879), .Q(n6328) );
  INVX0 U7012 ( .INP(n6330), .ZN(n350) );
  OR2X1 U7013 ( .IN1(n5467), .IN2(n3872), .Q(n6330) );
  OR2X1 U7014 ( .IN1(n6331), .IN2(n6332), .Q(n6326) );
  AND2X1 U7015 ( .IN1(n4842), .IN2(n6333), .Q(n6332) );
  AND2X1 U7016 ( .IN1(n4933), .IN2(n5965), .Q(n6331) );
  XNOR2X1 U7017 ( .IN1(n6334), .IN2(n6335), .Q(n5965) );
  XOR2X1 U7018 ( .IN1(n4192), .IN2(n5389), .Q(n6335) );
  XOR2X1 U7019 ( .IN1(n6336), .IN2(n4574), .Q(n6334) );
  XOR2X1 U7020 ( .IN1(WX9838), .IN2(n9545), .Q(n6336) );
  OR2X1 U7021 ( .IN1(n6337), .IN2(n6338), .Q(WX8414) );
  OR2X1 U7022 ( .IN1(n6339), .IN2(n6340), .Q(n6338) );
  AND2X1 U7023 ( .IN1(n4902), .IN2(CRC_OUT_3_25), .Q(n6340) );
  AND2X1 U7024 ( .IN1(n349), .IN2(n4879), .Q(n6339) );
  INVX0 U7025 ( .INP(n6341), .ZN(n349) );
  OR2X1 U7026 ( .IN1(n5467), .IN2(n3873), .Q(n6341) );
  OR2X1 U7027 ( .IN1(n6342), .IN2(n6343), .Q(n6337) );
  AND2X1 U7028 ( .IN1(n4842), .IN2(n6344), .Q(n6343) );
  AND2X1 U7029 ( .IN1(n4933), .IN2(n5974), .Q(n6342) );
  XNOR2X1 U7030 ( .IN1(n6345), .IN2(n6346), .Q(n5974) );
  XOR2X1 U7031 ( .IN1(n4193), .IN2(n5389), .Q(n6346) );
  XOR2X1 U7032 ( .IN1(n6347), .IN2(n4573), .Q(n6345) );
  XOR2X1 U7033 ( .IN1(WX9836), .IN2(n9546), .Q(n6347) );
  OR2X1 U7034 ( .IN1(n6348), .IN2(n6349), .Q(WX8412) );
  OR2X1 U7035 ( .IN1(n6350), .IN2(n6351), .Q(n6349) );
  AND2X1 U7036 ( .IN1(n4902), .IN2(CRC_OUT_3_26), .Q(n6351) );
  AND2X1 U7037 ( .IN1(n348), .IN2(n4879), .Q(n6350) );
  INVX0 U7038 ( .INP(n6352), .ZN(n348) );
  OR2X1 U7039 ( .IN1(n5467), .IN2(n3874), .Q(n6352) );
  OR2X1 U7040 ( .IN1(n6353), .IN2(n6354), .Q(n6348) );
  AND2X1 U7041 ( .IN1(n6355), .IN2(n4837), .Q(n6354) );
  AND2X1 U7042 ( .IN1(n4933), .IN2(n5983), .Q(n6353) );
  XNOR2X1 U7043 ( .IN1(n6356), .IN2(n6357), .Q(n5983) );
  XOR2X1 U7044 ( .IN1(n4194), .IN2(n5389), .Q(n6357) );
  XOR2X1 U7045 ( .IN1(n6358), .IN2(n4572), .Q(n6356) );
  XOR2X1 U7046 ( .IN1(WX9834), .IN2(n9547), .Q(n6358) );
  OR2X1 U7047 ( .IN1(n6359), .IN2(n6360), .Q(WX8410) );
  OR2X1 U7048 ( .IN1(n6361), .IN2(n6362), .Q(n6360) );
  AND2X1 U7049 ( .IN1(n4902), .IN2(CRC_OUT_3_27), .Q(n6362) );
  AND2X1 U7050 ( .IN1(n347), .IN2(n4879), .Q(n6361) );
  INVX0 U7051 ( .INP(n6363), .ZN(n347) );
  OR2X1 U7052 ( .IN1(n5467), .IN2(n3875), .Q(n6363) );
  OR2X1 U7053 ( .IN1(n6364), .IN2(n6365), .Q(n6359) );
  AND2X1 U7054 ( .IN1(n4842), .IN2(n6366), .Q(n6365) );
  AND2X1 U7055 ( .IN1(n4933), .IN2(n5992), .Q(n6364) );
  XNOR2X1 U7056 ( .IN1(n6367), .IN2(n6368), .Q(n5992) );
  XOR2X1 U7057 ( .IN1(n4195), .IN2(n5389), .Q(n6368) );
  XOR2X1 U7058 ( .IN1(n6369), .IN2(n4571), .Q(n6367) );
  XOR2X1 U7059 ( .IN1(WX9832), .IN2(n9548), .Q(n6369) );
  OR2X1 U7060 ( .IN1(n6370), .IN2(n6371), .Q(WX8408) );
  OR2X1 U7061 ( .IN1(n6372), .IN2(n6373), .Q(n6371) );
  AND2X1 U7062 ( .IN1(n4902), .IN2(CRC_OUT_3_28), .Q(n6373) );
  AND2X1 U7063 ( .IN1(n346), .IN2(n4879), .Q(n6372) );
  INVX0 U7064 ( .INP(n6374), .ZN(n346) );
  OR2X1 U7065 ( .IN1(n5467), .IN2(n3876), .Q(n6374) );
  OR2X1 U7066 ( .IN1(n6375), .IN2(n6376), .Q(n6370) );
  AND2X1 U7067 ( .IN1(n6377), .IN2(n4838), .Q(n6376) );
  AND2X1 U7068 ( .IN1(n4933), .IN2(n6001), .Q(n6375) );
  XNOR2X1 U7069 ( .IN1(n6378), .IN2(n6379), .Q(n6001) );
  XOR2X1 U7070 ( .IN1(n4196), .IN2(n5389), .Q(n6379) );
  XOR2X1 U7071 ( .IN1(n6380), .IN2(n4570), .Q(n6378) );
  XOR2X1 U7072 ( .IN1(WX9830), .IN2(n9549), .Q(n6380) );
  OR2X1 U7073 ( .IN1(n6381), .IN2(n6382), .Q(WX8406) );
  OR2X1 U7074 ( .IN1(n6383), .IN2(n6384), .Q(n6382) );
  AND2X1 U7075 ( .IN1(n4902), .IN2(CRC_OUT_3_29), .Q(n6384) );
  AND2X1 U7076 ( .IN1(n345), .IN2(n4879), .Q(n6383) );
  INVX0 U7077 ( .INP(n6385), .ZN(n345) );
  OR2X1 U7078 ( .IN1(n5467), .IN2(n3877), .Q(n6385) );
  OR2X1 U7079 ( .IN1(n6386), .IN2(n6387), .Q(n6381) );
  AND2X1 U7080 ( .IN1(n4842), .IN2(n6388), .Q(n6387) );
  AND2X1 U7081 ( .IN1(n4933), .IN2(n6010), .Q(n6386) );
  XNOR2X1 U7082 ( .IN1(n6389), .IN2(n6390), .Q(n6010) );
  XOR2X1 U7083 ( .IN1(n4197), .IN2(n5388), .Q(n6390) );
  XOR2X1 U7084 ( .IN1(n6391), .IN2(n4569), .Q(n6389) );
  XOR2X1 U7085 ( .IN1(WX9828), .IN2(n9550), .Q(n6391) );
  OR2X1 U7086 ( .IN1(n6392), .IN2(n6393), .Q(WX8404) );
  OR2X1 U7087 ( .IN1(n6394), .IN2(n6395), .Q(n6393) );
  AND2X1 U7088 ( .IN1(n4902), .IN2(CRC_OUT_3_30), .Q(n6395) );
  AND2X1 U7089 ( .IN1(n344), .IN2(n4879), .Q(n6394) );
  INVX0 U7090 ( .INP(n6396), .ZN(n344) );
  OR2X1 U7091 ( .IN1(n5466), .IN2(n3878), .Q(n6396) );
  OR2X1 U7092 ( .IN1(n6397), .IN2(n6398), .Q(n6392) );
  AND2X1 U7093 ( .IN1(n6399), .IN2(n4837), .Q(n6398) );
  AND2X1 U7094 ( .IN1(n4933), .IN2(n6019), .Q(n6397) );
  XNOR2X1 U7095 ( .IN1(n6400), .IN2(n6401), .Q(n6019) );
  XOR2X1 U7096 ( .IN1(n4198), .IN2(n5388), .Q(n6401) );
  XOR2X1 U7097 ( .IN1(n6402), .IN2(n4568), .Q(n6400) );
  XOR2X1 U7098 ( .IN1(WX9826), .IN2(n9551), .Q(n6402) );
  OR2X1 U7099 ( .IN1(n6403), .IN2(n6404), .Q(WX8402) );
  OR2X1 U7100 ( .IN1(n6405), .IN2(n6406), .Q(n6404) );
  AND2X1 U7101 ( .IN1(n2245), .IN2(WX8243), .Q(n6406) );
  AND2X1 U7102 ( .IN1(n4903), .IN2(CRC_OUT_3_31), .Q(n6405) );
  OR2X1 U7103 ( .IN1(n6407), .IN2(n6408), .Q(n6403) );
  AND2X1 U7104 ( .IN1(n4842), .IN2(n6409), .Q(n6408) );
  AND2X1 U7105 ( .IN1(n6027), .IN2(n4920), .Q(n6407) );
  XOR2X1 U7106 ( .IN1(n6410), .IN2(n6411), .Q(n6027) );
  XOR2X1 U7107 ( .IN1(n4166), .IN2(n5388), .Q(n6411) );
  XOR2X1 U7108 ( .IN1(WX9760), .IN2(n6412), .Q(n6410) );
  XOR2X1 U7109 ( .IN1(test_so85), .IN2(n9552), .Q(n6412) );
  AND2X1 U7110 ( .IN1(n4824), .IN2(n5411), .Q(WX8304) );
  AND2X1 U7111 ( .IN1(n6413), .IN2(n8399), .Q(WX8266) );
  AND2X1 U7112 ( .IN1(n6414), .IN2(n5411), .Q(WX7791) );
  XOR2X1 U7113 ( .IN1(CRC_OUT_4_30), .IN2(n4620), .Q(n6414) );
  AND2X1 U7114 ( .IN1(n6415), .IN2(n5411), .Q(WX7789) );
  XOR2X1 U7115 ( .IN1(test_so66), .IN2(n4621), .Q(n6415) );
  AND2X1 U7116 ( .IN1(n6416), .IN2(n5410), .Q(WX7787) );
  XOR2X1 U7117 ( .IN1(CRC_OUT_4_28), .IN2(n4622), .Q(n6416) );
  AND2X1 U7118 ( .IN1(n6417), .IN2(n5410), .Q(WX7785) );
  XOR2X1 U7119 ( .IN1(CRC_OUT_4_27), .IN2(n4623), .Q(n6417) );
  AND2X1 U7120 ( .IN1(n6418), .IN2(n6413), .Q(WX7783) );
  XOR2X1 U7121 ( .IN1(CRC_OUT_4_26), .IN2(n4624), .Q(n6418) );
  AND2X1 U7122 ( .IN1(n6419), .IN2(n5410), .Q(WX7781) );
  XOR2X1 U7123 ( .IN1(CRC_OUT_4_25), .IN2(n4625), .Q(n6419) );
  AND2X1 U7124 ( .IN1(n6420), .IN2(n5410), .Q(WX7779) );
  XOR2X1 U7125 ( .IN1(CRC_OUT_4_24), .IN2(n4626), .Q(n6420) );
  AND2X1 U7126 ( .IN1(n6421), .IN2(n5410), .Q(WX7777) );
  XOR2X1 U7127 ( .IN1(CRC_OUT_4_23), .IN2(n4627), .Q(n6421) );
  AND2X1 U7128 ( .IN1(n6422), .IN2(n5410), .Q(WX7775) );
  XOR2X1 U7129 ( .IN1(CRC_OUT_4_22), .IN2(n4628), .Q(n6422) );
  AND2X1 U7130 ( .IN1(n6423), .IN2(n5410), .Q(WX7773) );
  XOR2X1 U7131 ( .IN1(CRC_OUT_4_21), .IN2(n4629), .Q(n6423) );
  AND2X1 U7132 ( .IN1(n6424), .IN2(n5410), .Q(WX7771) );
  XOR2X1 U7133 ( .IN1(test_so63), .IN2(DFF_1140_n1), .Q(n6424) );
  AND2X1 U7134 ( .IN1(n6425), .IN2(n5410), .Q(WX7769) );
  XOR2X1 U7135 ( .IN1(CRC_OUT_4_19), .IN2(n4630), .Q(n6425) );
  AND2X1 U7136 ( .IN1(n6426), .IN2(n5409), .Q(WX7767) );
  XOR2X1 U7137 ( .IN1(CRC_OUT_4_18), .IN2(n4631), .Q(n6426) );
  AND2X1 U7138 ( .IN1(n6427), .IN2(n5409), .Q(WX7765) );
  XOR2X1 U7139 ( .IN1(CRC_OUT_4_17), .IN2(n4632), .Q(n6427) );
  AND2X1 U7140 ( .IN1(n6428), .IN2(n5409), .Q(WX7763) );
  XOR2X1 U7141 ( .IN1(CRC_OUT_4_16), .IN2(n4633), .Q(n6428) );
  AND2X1 U7142 ( .IN1(n6429), .IN2(n5409), .Q(WX7761) );
  XOR2X1 U7143 ( .IN1(DFF_1135_n1), .IN2(n6430), .Q(n6429) );
  XOR2X1 U7144 ( .IN1(n4522), .IN2(DFF_1151_n1), .Q(n6430) );
  AND2X1 U7145 ( .IN1(n6431), .IN2(n5409), .Q(WX7759) );
  XOR2X1 U7146 ( .IN1(CRC_OUT_4_14), .IN2(n4634), .Q(n6431) );
  AND2X1 U7147 ( .IN1(n6432), .IN2(n5409), .Q(WX7757) );
  XOR2X1 U7148 ( .IN1(CRC_OUT_4_13), .IN2(n4635), .Q(n6432) );
  AND2X1 U7149 ( .IN1(n6433), .IN2(n5409), .Q(WX7755) );
  XOR2X1 U7150 ( .IN1(test_so65), .IN2(n4636), .Q(n6433) );
  AND2X1 U7151 ( .IN1(n6434), .IN2(n5409), .Q(WX7753) );
  XOR2X1 U7152 ( .IN1(CRC_OUT_4_11), .IN2(n4637), .Q(n6434) );
  AND2X1 U7153 ( .IN1(n6435), .IN2(n5409), .Q(WX7751) );
  XOR2X1 U7154 ( .IN1(DFF_1130_n1), .IN2(n6436), .Q(n6435) );
  XOR2X1 U7155 ( .IN1(n4523), .IN2(DFF_1151_n1), .Q(n6436) );
  AND2X1 U7156 ( .IN1(n6437), .IN2(n5408), .Q(WX7749) );
  XOR2X1 U7157 ( .IN1(CRC_OUT_4_9), .IN2(n4638), .Q(n6437) );
  AND2X1 U7158 ( .IN1(n6438), .IN2(n5408), .Q(WX7747) );
  XOR2X1 U7159 ( .IN1(CRC_OUT_4_8), .IN2(n4639), .Q(n6438) );
  AND2X1 U7160 ( .IN1(n6439), .IN2(n5408), .Q(WX7745) );
  XOR2X1 U7161 ( .IN1(CRC_OUT_4_7), .IN2(n4640), .Q(n6439) );
  AND2X1 U7162 ( .IN1(n6440), .IN2(n5408), .Q(WX7743) );
  XOR2X1 U7163 ( .IN1(CRC_OUT_4_6), .IN2(n4641), .Q(n6440) );
  AND2X1 U7164 ( .IN1(n6441), .IN2(n5408), .Q(WX7741) );
  XOR2X1 U7165 ( .IN1(CRC_OUT_4_5), .IN2(n4642), .Q(n6441) );
  AND2X1 U7166 ( .IN1(n6442), .IN2(n5408), .Q(WX7739) );
  XOR2X1 U7167 ( .IN1(CRC_OUT_4_4), .IN2(n4643), .Q(n6442) );
  AND2X1 U7168 ( .IN1(n6443), .IN2(n5408), .Q(WX7737) );
  XOR2X1 U7169 ( .IN1(CRC_OUT_4_3), .IN2(n6444), .Q(n6443) );
  XOR2X1 U7170 ( .IN1(test_so64), .IN2(DFF_1151_n1), .Q(n6444) );
  AND2X1 U7171 ( .IN1(n6445), .IN2(n5404), .Q(WX7735) );
  XOR2X1 U7172 ( .IN1(CRC_OUT_4_2), .IN2(n4644), .Q(n6445) );
  AND2X1 U7173 ( .IN1(n6446), .IN2(n5401), .Q(WX7733) );
  XOR2X1 U7174 ( .IN1(CRC_OUT_4_1), .IN2(n4645), .Q(n6446) );
  AND2X1 U7175 ( .IN1(n6447), .IN2(n5401), .Q(WX7731) );
  XOR2X1 U7176 ( .IN1(CRC_OUT_4_0), .IN2(n4646), .Q(n6447) );
  AND2X1 U7177 ( .IN1(n6448), .IN2(n5401), .Q(WX7729) );
  XOR2X1 U7178 ( .IN1(n4537), .IN2(CRC_OUT_4_31), .Q(n6448) );
  INVX0 U7179 ( .INP(n6449), .ZN(WX7203) );
  OR2X1 U7180 ( .IN1(n5466), .IN2(n9605), .Q(n6449) );
  INVX0 U7181 ( .INP(n6450), .ZN(WX7201) );
  OR2X1 U7182 ( .IN1(n5466), .IN2(n9606), .Q(n6450) );
  INVX0 U7183 ( .INP(n6451), .ZN(WX7199) );
  OR2X1 U7184 ( .IN1(n5466), .IN2(n9607), .Q(n6451) );
  INVX0 U7185 ( .INP(n6452), .ZN(WX7197) );
  OR2X1 U7186 ( .IN1(n5466), .IN2(n9608), .Q(n6452) );
  INVX0 U7187 ( .INP(n6453), .ZN(WX7195) );
  OR2X1 U7188 ( .IN1(n5466), .IN2(n9609), .Q(n6453) );
  INVX0 U7189 ( .INP(n6454), .ZN(WX7193) );
  OR2X1 U7190 ( .IN1(n5466), .IN2(n9610), .Q(n6454) );
  INVX0 U7191 ( .INP(n6455), .ZN(WX7191) );
  OR2X1 U7192 ( .IN1(n5466), .IN2(n9611), .Q(n6455) );
  INVX0 U7193 ( .INP(n6456), .ZN(WX7189) );
  OR2X1 U7194 ( .IN1(n5466), .IN2(n9612), .Q(n6456) );
  INVX0 U7195 ( .INP(n6457), .ZN(WX7187) );
  OR2X1 U7196 ( .IN1(n5466), .IN2(n9615), .Q(n6457) );
  INVX0 U7197 ( .INP(n6458), .ZN(WX7185) );
  OR2X1 U7198 ( .IN1(n5466), .IN2(n9616), .Q(n6458) );
  INVX0 U7199 ( .INP(n6459), .ZN(WX7183) );
  OR2X1 U7200 ( .IN1(n5466), .IN2(n9619), .Q(n6459) );
  AND2X1 U7201 ( .IN1(test_so57), .IN2(n5401), .Q(WX7181) );
  INVX0 U7202 ( .INP(n6460), .ZN(WX7179) );
  OR2X1 U7203 ( .IN1(n5466), .IN2(n9620), .Q(n6460) );
  INVX0 U7204 ( .INP(n6461), .ZN(WX7177) );
  OR2X1 U7205 ( .IN1(n5465), .IN2(n9621), .Q(n6461) );
  INVX0 U7206 ( .INP(n6462), .ZN(WX7175) );
  OR2X1 U7207 ( .IN1(n5465), .IN2(n9622), .Q(n6462) );
  INVX0 U7208 ( .INP(n6463), .ZN(WX7173) );
  OR2X1 U7209 ( .IN1(n5465), .IN2(n9623), .Q(n6463) );
  OR2X1 U7210 ( .IN1(n6464), .IN2(n6465), .Q(WX7171) );
  OR2X1 U7211 ( .IN1(n6466), .IN2(n6467), .Q(n6465) );
  AND2X1 U7212 ( .IN1(n4903), .IN2(CRC_OUT_4_0), .Q(n6467) );
  AND2X1 U7213 ( .IN1(n312), .IN2(n4879), .Q(n6466) );
  INVX0 U7214 ( .INP(n6468), .ZN(n312) );
  OR2X1 U7215 ( .IN1(n5465), .IN2(n3879), .Q(n6468) );
  OR2X1 U7216 ( .IN1(n6469), .IN2(n6470), .Q(n6464) );
  AND2X1 U7217 ( .IN1(n4842), .IN2(n6471), .Q(n6470) );
  AND2X1 U7218 ( .IN1(n4933), .IN2(n6086), .Q(n6469) );
  XNOR2X1 U7219 ( .IN1(n6472), .IN2(n6473), .Q(n6086) );
  XOR2X1 U7220 ( .IN1(n9553), .IN2(n4536), .Q(n6473) );
  XOR2X1 U7221 ( .IN1(WX8465), .IN2(n4339), .Q(n6472) );
  OR2X1 U7222 ( .IN1(n6474), .IN2(n6475), .Q(WX7169) );
  OR2X1 U7223 ( .IN1(n6476), .IN2(n6477), .Q(n6475) );
  AND2X1 U7224 ( .IN1(n4903), .IN2(CRC_OUT_4_1), .Q(n6477) );
  AND2X1 U7225 ( .IN1(n311), .IN2(n4878), .Q(n6476) );
  INVX0 U7226 ( .INP(n6478), .ZN(n311) );
  OR2X1 U7227 ( .IN1(n5465), .IN2(n3880), .Q(n6478) );
  OR2X1 U7228 ( .IN1(n6479), .IN2(n6480), .Q(n6474) );
  AND2X1 U7229 ( .IN1(n4841), .IN2(n6481), .Q(n6480) );
  AND2X1 U7230 ( .IN1(n4933), .IN2(n6096), .Q(n6479) );
  XNOR2X1 U7231 ( .IN1(n6482), .IN2(n6483), .Q(n6096) );
  XOR2X1 U7232 ( .IN1(n9554), .IN2(n4619), .Q(n6483) );
  XOR2X1 U7233 ( .IN1(WX8463), .IN2(n4341), .Q(n6482) );
  OR2X1 U7234 ( .IN1(n6484), .IN2(n6485), .Q(WX7167) );
  OR2X1 U7235 ( .IN1(n6486), .IN2(n6487), .Q(n6485) );
  AND2X1 U7236 ( .IN1(n4903), .IN2(CRC_OUT_4_2), .Q(n6487) );
  AND2X1 U7237 ( .IN1(n310), .IN2(n4878), .Q(n6486) );
  INVX0 U7238 ( .INP(n6488), .ZN(n310) );
  OR2X1 U7239 ( .IN1(n5465), .IN2(n3881), .Q(n6488) );
  OR2X1 U7240 ( .IN1(n6489), .IN2(n6490), .Q(n6484) );
  AND2X1 U7241 ( .IN1(n4841), .IN2(n6491), .Q(n6490) );
  AND2X1 U7242 ( .IN1(n4933), .IN2(n6106), .Q(n6489) );
  XNOR2X1 U7243 ( .IN1(n6492), .IN2(n6493), .Q(n6106) );
  XOR2X1 U7244 ( .IN1(n9555), .IN2(n4618), .Q(n6493) );
  XOR2X1 U7245 ( .IN1(WX8461), .IN2(n4343), .Q(n6492) );
  OR2X1 U7246 ( .IN1(n6494), .IN2(n6495), .Q(WX7165) );
  OR2X1 U7247 ( .IN1(n6496), .IN2(n6497), .Q(n6495) );
  AND2X1 U7248 ( .IN1(n4903), .IN2(CRC_OUT_4_3), .Q(n6497) );
  AND2X1 U7249 ( .IN1(n309), .IN2(n4878), .Q(n6496) );
  INVX0 U7250 ( .INP(n6498), .ZN(n309) );
  OR2X1 U7251 ( .IN1(n5465), .IN2(n3882), .Q(n6498) );
  OR2X1 U7252 ( .IN1(n6499), .IN2(n6500), .Q(n6494) );
  AND2X1 U7253 ( .IN1(n4841), .IN2(n6501), .Q(n6500) );
  AND2X1 U7254 ( .IN1(n4934), .IN2(n6116), .Q(n6499) );
  XNOR2X1 U7255 ( .IN1(n6502), .IN2(n6503), .Q(n6116) );
  XOR2X1 U7256 ( .IN1(n9556), .IN2(n4617), .Q(n6503) );
  XOR2X1 U7257 ( .IN1(WX8459), .IN2(n4345), .Q(n6502) );
  OR2X1 U7258 ( .IN1(n6504), .IN2(n6505), .Q(WX7163) );
  OR2X1 U7259 ( .IN1(n6506), .IN2(n6507), .Q(n6505) );
  AND2X1 U7260 ( .IN1(n4903), .IN2(CRC_OUT_4_4), .Q(n6507) );
  AND2X1 U7261 ( .IN1(n308), .IN2(n4878), .Q(n6506) );
  INVX0 U7262 ( .INP(n6508), .ZN(n308) );
  OR2X1 U7263 ( .IN1(n5465), .IN2(n3883), .Q(n6508) );
  OR2X1 U7264 ( .IN1(n6509), .IN2(n6510), .Q(n6504) );
  AND2X1 U7265 ( .IN1(n6511), .IN2(n4835), .Q(n6510) );
  AND2X1 U7266 ( .IN1(n4934), .IN2(n6126), .Q(n6509) );
  XNOR2X1 U7267 ( .IN1(n6512), .IN2(n6513), .Q(n6126) );
  XOR2X1 U7268 ( .IN1(n9557), .IN2(n4521), .Q(n6513) );
  XOR2X1 U7269 ( .IN1(WX8457), .IN2(n4347), .Q(n6512) );
  OR2X1 U7270 ( .IN1(n6514), .IN2(n6515), .Q(WX7161) );
  OR2X1 U7271 ( .IN1(n6516), .IN2(n6517), .Q(n6515) );
  AND2X1 U7272 ( .IN1(n4903), .IN2(CRC_OUT_4_5), .Q(n6517) );
  AND2X1 U7273 ( .IN1(WX6999), .IN2(n4878), .Q(n6516) );
  OR2X1 U7274 ( .IN1(n6518), .IN2(n6519), .Q(n6514) );
  AND2X1 U7275 ( .IN1(n4841), .IN2(n6520), .Q(n6519) );
  AND2X1 U7276 ( .IN1(n4934), .IN2(n6136), .Q(n6518) );
  XNOR2X1 U7277 ( .IN1(n6521), .IN2(n6522), .Q(n6136) );
  XOR2X1 U7278 ( .IN1(n9558), .IN2(n4616), .Q(n6522) );
  XOR2X1 U7279 ( .IN1(WX8455), .IN2(n4349), .Q(n6521) );
  OR2X1 U7280 ( .IN1(n6523), .IN2(n6524), .Q(WX7159) );
  OR2X1 U7281 ( .IN1(n6525), .IN2(n6526), .Q(n6524) );
  AND2X1 U7282 ( .IN1(n4903), .IN2(CRC_OUT_4_6), .Q(n6526) );
  AND2X1 U7283 ( .IN1(n306), .IN2(n4878), .Q(n6525) );
  INVX0 U7284 ( .INP(n6527), .ZN(n306) );
  OR2X1 U7285 ( .IN1(n5465), .IN2(n3885), .Q(n6527) );
  OR2X1 U7286 ( .IN1(n6528), .IN2(n6529), .Q(n6523) );
  AND2X1 U7287 ( .IN1(n6530), .IN2(n4835), .Q(n6529) );
  AND2X1 U7288 ( .IN1(n4934), .IN2(n6146), .Q(n6528) );
  XNOR2X1 U7289 ( .IN1(n6531), .IN2(n6532), .Q(n6146) );
  XOR2X1 U7290 ( .IN1(n9559), .IN2(n4615), .Q(n6532) );
  XOR2X1 U7291 ( .IN1(WX8453), .IN2(n4351), .Q(n6531) );
  OR2X1 U7292 ( .IN1(n6533), .IN2(n6534), .Q(WX7157) );
  OR2X1 U7293 ( .IN1(n6535), .IN2(n6536), .Q(n6534) );
  AND2X1 U7294 ( .IN1(n4903), .IN2(CRC_OUT_4_7), .Q(n6536) );
  AND2X1 U7295 ( .IN1(n305), .IN2(n4878), .Q(n6535) );
  INVX0 U7296 ( .INP(n6537), .ZN(n305) );
  OR2X1 U7297 ( .IN1(n5465), .IN2(n3886), .Q(n6537) );
  OR2X1 U7298 ( .IN1(n6538), .IN2(n6539), .Q(n6533) );
  AND2X1 U7299 ( .IN1(n4841), .IN2(n6540), .Q(n6539) );
  AND2X1 U7300 ( .IN1(n4934), .IN2(n6156), .Q(n6538) );
  XNOR2X1 U7301 ( .IN1(n6541), .IN2(n6542), .Q(n6156) );
  XOR2X1 U7302 ( .IN1(n9560), .IN2(n4614), .Q(n6542) );
  XOR2X1 U7303 ( .IN1(WX8451), .IN2(n4353), .Q(n6541) );
  OR2X1 U7304 ( .IN1(n6543), .IN2(n6544), .Q(WX7155) );
  OR2X1 U7305 ( .IN1(n6545), .IN2(n6546), .Q(n6544) );
  AND2X1 U7306 ( .IN1(n4903), .IN2(CRC_OUT_4_8), .Q(n6546) );
  AND2X1 U7307 ( .IN1(n304), .IN2(n4878), .Q(n6545) );
  INVX0 U7308 ( .INP(n6547), .ZN(n304) );
  OR2X1 U7309 ( .IN1(n5465), .IN2(n3887), .Q(n6547) );
  OR2X1 U7310 ( .IN1(n6548), .IN2(n6549), .Q(n6543) );
  AND2X1 U7311 ( .IN1(n6550), .IN2(n4834), .Q(n6549) );
  AND2X1 U7312 ( .IN1(n4934), .IN2(n6166), .Q(n6548) );
  XNOR2X1 U7313 ( .IN1(n6551), .IN2(n6552), .Q(n6166) );
  XOR2X1 U7314 ( .IN1(n9561), .IN2(n4613), .Q(n6552) );
  XOR2X1 U7315 ( .IN1(WX8449), .IN2(n4355), .Q(n6551) );
  OR2X1 U7316 ( .IN1(n6553), .IN2(n6554), .Q(WX7153) );
  OR2X1 U7317 ( .IN1(n6555), .IN2(n6556), .Q(n6554) );
  AND2X1 U7318 ( .IN1(n4903), .IN2(CRC_OUT_4_9), .Q(n6556) );
  AND2X1 U7319 ( .IN1(n303), .IN2(n4878), .Q(n6555) );
  INVX0 U7320 ( .INP(n6557), .ZN(n303) );
  OR2X1 U7321 ( .IN1(n5465), .IN2(n3888), .Q(n6557) );
  OR2X1 U7322 ( .IN1(n6558), .IN2(n6559), .Q(n6553) );
  AND2X1 U7323 ( .IN1(n4841), .IN2(n6560), .Q(n6559) );
  AND2X1 U7324 ( .IN1(n6176), .IN2(n4919), .Q(n6558) );
  XOR2X1 U7325 ( .IN1(n6561), .IN2(n6562), .Q(n6176) );
  XOR2X1 U7326 ( .IN1(test_so75), .IN2(n9562), .Q(n6562) );
  XOR2X1 U7327 ( .IN1(WX8447), .IN2(n4357), .Q(n6561) );
  OR2X1 U7328 ( .IN1(n6563), .IN2(n6564), .Q(WX7151) );
  OR2X1 U7329 ( .IN1(n6565), .IN2(n6566), .Q(n6564) );
  AND2X1 U7330 ( .IN1(n4903), .IN2(CRC_OUT_4_10), .Q(n6566) );
  AND2X1 U7331 ( .IN1(n302), .IN2(n4878), .Q(n6565) );
  INVX0 U7332 ( .INP(n6567), .ZN(n302) );
  OR2X1 U7333 ( .IN1(n5465), .IN2(n3889), .Q(n6567) );
  OR2X1 U7334 ( .IN1(n6568), .IN2(n6569), .Q(n6563) );
  AND2X1 U7335 ( .IN1(n6570), .IN2(n4834), .Q(n6569) );
  AND2X1 U7336 ( .IN1(n4934), .IN2(n6186), .Q(n6568) );
  XNOR2X1 U7337 ( .IN1(n6571), .IN2(n6572), .Q(n6186) );
  XOR2X1 U7338 ( .IN1(n9563), .IN2(n4612), .Q(n6572) );
  XOR2X1 U7339 ( .IN1(WX8445), .IN2(n4359), .Q(n6571) );
  OR2X1 U7340 ( .IN1(n6573), .IN2(n6574), .Q(WX7149) );
  OR2X1 U7341 ( .IN1(n6575), .IN2(n6576), .Q(n6574) );
  AND2X1 U7342 ( .IN1(n4904), .IN2(CRC_OUT_4_11), .Q(n6576) );
  AND2X1 U7343 ( .IN1(n301), .IN2(n4878), .Q(n6575) );
  INVX0 U7344 ( .INP(n6577), .ZN(n301) );
  OR2X1 U7345 ( .IN1(n5464), .IN2(n3890), .Q(n6577) );
  OR2X1 U7346 ( .IN1(n6578), .IN2(n6579), .Q(n6573) );
  AND2X1 U7347 ( .IN1(n4841), .IN2(n6580), .Q(n6579) );
  AND2X1 U7348 ( .IN1(n6196), .IN2(n4919), .Q(n6578) );
  XOR2X1 U7349 ( .IN1(n6581), .IN2(n6582), .Q(n6196) );
  XOR2X1 U7350 ( .IN1(test_so73), .IN2(n9564), .Q(n6582) );
  XOR2X1 U7351 ( .IN1(WX8443), .IN2(n4520), .Q(n6581) );
  OR2X1 U7352 ( .IN1(n6583), .IN2(n6584), .Q(WX7147) );
  OR2X1 U7353 ( .IN1(n6585), .IN2(n6586), .Q(n6584) );
  AND2X1 U7354 ( .IN1(test_so65), .IN2(n4887), .Q(n6586) );
  AND2X1 U7355 ( .IN1(n300), .IN2(n4878), .Q(n6585) );
  INVX0 U7356 ( .INP(n6587), .ZN(n300) );
  OR2X1 U7357 ( .IN1(n5464), .IN2(n3891), .Q(n6587) );
  OR2X1 U7358 ( .IN1(n6588), .IN2(n6589), .Q(n6583) );
  AND2X1 U7359 ( .IN1(n4841), .IN2(n6590), .Q(n6589) );
  AND2X1 U7360 ( .IN1(n4934), .IN2(n6206), .Q(n6588) );
  XNOR2X1 U7361 ( .IN1(n6591), .IN2(n6592), .Q(n6206) );
  XOR2X1 U7362 ( .IN1(n9565), .IN2(n4611), .Q(n6592) );
  XOR2X1 U7363 ( .IN1(WX8441), .IN2(n4362), .Q(n6591) );
  OR2X1 U7364 ( .IN1(n6593), .IN2(n6594), .Q(WX7145) );
  OR2X1 U7365 ( .IN1(n6595), .IN2(n6596), .Q(n6594) );
  AND2X1 U7366 ( .IN1(n4904), .IN2(CRC_OUT_4_13), .Q(n6596) );
  AND2X1 U7367 ( .IN1(n299), .IN2(n4877), .Q(n6595) );
  INVX0 U7368 ( .INP(n6597), .ZN(n299) );
  OR2X1 U7369 ( .IN1(n5464), .IN2(n3892), .Q(n6597) );
  OR2X1 U7370 ( .IN1(n6598), .IN2(n6599), .Q(n6593) );
  AND2X1 U7371 ( .IN1(n4841), .IN2(n6600), .Q(n6599) );
  AND2X1 U7372 ( .IN1(n6216), .IN2(n4919), .Q(n6598) );
  XOR2X1 U7373 ( .IN1(n6601), .IN2(n6602), .Q(n6216) );
  XOR2X1 U7374 ( .IN1(test_so71), .IN2(n9566), .Q(n6602) );
  XOR2X1 U7375 ( .IN1(WX8439), .IN2(n4610), .Q(n6601) );
  OR2X1 U7376 ( .IN1(n6603), .IN2(n6604), .Q(WX7143) );
  OR2X1 U7377 ( .IN1(n6605), .IN2(n6606), .Q(n6604) );
  AND2X1 U7378 ( .IN1(n4904), .IN2(CRC_OUT_4_14), .Q(n6606) );
  AND2X1 U7379 ( .IN1(n298), .IN2(n4877), .Q(n6605) );
  INVX0 U7380 ( .INP(n6607), .ZN(n298) );
  OR2X1 U7381 ( .IN1(n5464), .IN2(n3893), .Q(n6607) );
  OR2X1 U7382 ( .IN1(n6608), .IN2(n6609), .Q(n6603) );
  AND2X1 U7383 ( .IN1(n4838), .IN2(n6610), .Q(n6609) );
  AND2X1 U7384 ( .IN1(n4934), .IN2(n6226), .Q(n6608) );
  XNOR2X1 U7385 ( .IN1(n6611), .IN2(n6612), .Q(n6226) );
  XOR2X1 U7386 ( .IN1(n9567), .IN2(n4609), .Q(n6612) );
  XOR2X1 U7387 ( .IN1(WX8437), .IN2(n4365), .Q(n6611) );
  OR2X1 U7388 ( .IN1(n6613), .IN2(n6614), .Q(WX7141) );
  OR2X1 U7389 ( .IN1(n6615), .IN2(n6616), .Q(n6614) );
  AND2X1 U7390 ( .IN1(n4904), .IN2(CRC_OUT_4_15), .Q(n6616) );
  AND2X1 U7391 ( .IN1(n297), .IN2(n4877), .Q(n6615) );
  INVX0 U7392 ( .INP(n6617), .ZN(n297) );
  OR2X1 U7393 ( .IN1(n5464), .IN2(n3894), .Q(n6617) );
  OR2X1 U7394 ( .IN1(n6618), .IN2(n6619), .Q(n6613) );
  AND2X1 U7395 ( .IN1(n4838), .IN2(n6620), .Q(n6619) );
  AND2X1 U7396 ( .IN1(n6236), .IN2(n4919), .Q(n6618) );
  XOR2X1 U7397 ( .IN1(n6621), .IN2(n6622), .Q(n6236) );
  XOR2X1 U7398 ( .IN1(test_so69), .IN2(n9568), .Q(n6622) );
  XOR2X1 U7399 ( .IN1(WX8563), .IN2(n4608), .Q(n6621) );
  OR2X1 U7400 ( .IN1(n6623), .IN2(n6624), .Q(WX7139) );
  OR2X1 U7401 ( .IN1(n6625), .IN2(n6626), .Q(n6624) );
  AND2X1 U7402 ( .IN1(n4904), .IN2(CRC_OUT_4_16), .Q(n6626) );
  AND2X1 U7403 ( .IN1(n296), .IN2(n4877), .Q(n6625) );
  INVX0 U7404 ( .INP(n6627), .ZN(n296) );
  OR2X1 U7405 ( .IN1(n5464), .IN2(n3895), .Q(n6627) );
  OR2X1 U7406 ( .IN1(n6628), .IN2(n6629), .Q(n6623) );
  AND2X1 U7407 ( .IN1(n4838), .IN2(n6630), .Q(n6629) );
  AND2X1 U7408 ( .IN1(n4934), .IN2(n6246), .Q(n6628) );
  XNOR2X1 U7409 ( .IN1(n6631), .IN2(n6632), .Q(n6246) );
  XOR2X1 U7410 ( .IN1(n4199), .IN2(n5388), .Q(n6632) );
  XOR2X1 U7411 ( .IN1(n6633), .IN2(n4519), .Q(n6631) );
  XOR2X1 U7412 ( .IN1(WX8561), .IN2(n9569), .Q(n6633) );
  OR2X1 U7413 ( .IN1(n6634), .IN2(n6635), .Q(WX7137) );
  OR2X1 U7414 ( .IN1(n6636), .IN2(n6637), .Q(n6635) );
  AND2X1 U7415 ( .IN1(n4904), .IN2(CRC_OUT_4_17), .Q(n6637) );
  AND2X1 U7416 ( .IN1(n295), .IN2(n4877), .Q(n6636) );
  INVX0 U7417 ( .INP(n6638), .ZN(n295) );
  OR2X1 U7418 ( .IN1(n5464), .IN2(n3896), .Q(n6638) );
  OR2X1 U7419 ( .IN1(n6639), .IN2(n6640), .Q(n6634) );
  AND2X1 U7420 ( .IN1(n4838), .IN2(n6641), .Q(n6640) );
  AND2X1 U7421 ( .IN1(n4934), .IN2(n6257), .Q(n6639) );
  XNOR2X1 U7422 ( .IN1(n6642), .IN2(n6643), .Q(n6257) );
  XOR2X1 U7423 ( .IN1(n4200), .IN2(n5388), .Q(n6643) );
  XOR2X1 U7424 ( .IN1(n6644), .IN2(n4607), .Q(n6642) );
  XOR2X1 U7425 ( .IN1(WX8559), .IN2(n9570), .Q(n6644) );
  OR2X1 U7426 ( .IN1(n6645), .IN2(n6646), .Q(WX7135) );
  OR2X1 U7427 ( .IN1(n6647), .IN2(n6648), .Q(n6646) );
  AND2X1 U7428 ( .IN1(n4904), .IN2(CRC_OUT_4_18), .Q(n6648) );
  AND2X1 U7429 ( .IN1(n294), .IN2(n4877), .Q(n6647) );
  INVX0 U7430 ( .INP(n6649), .ZN(n294) );
  OR2X1 U7431 ( .IN1(n5464), .IN2(n3897), .Q(n6649) );
  OR2X1 U7432 ( .IN1(n6650), .IN2(n6651), .Q(n6645) );
  AND2X1 U7433 ( .IN1(n4838), .IN2(n6652), .Q(n6651) );
  AND2X1 U7434 ( .IN1(n4934), .IN2(n6267), .Q(n6650) );
  XNOR2X1 U7435 ( .IN1(n6653), .IN2(n6654), .Q(n6267) );
  XOR2X1 U7436 ( .IN1(n4201), .IN2(n5388), .Q(n6654) );
  XOR2X1 U7437 ( .IN1(n6655), .IN2(n4606), .Q(n6653) );
  XOR2X1 U7438 ( .IN1(WX8557), .IN2(n9571), .Q(n6655) );
  OR2X1 U7439 ( .IN1(n6656), .IN2(n6657), .Q(WX7133) );
  OR2X1 U7440 ( .IN1(n6658), .IN2(n6659), .Q(n6657) );
  AND2X1 U7441 ( .IN1(n4904), .IN2(CRC_OUT_4_19), .Q(n6659) );
  AND2X1 U7442 ( .IN1(n293), .IN2(n4877), .Q(n6658) );
  INVX0 U7443 ( .INP(n6660), .ZN(n293) );
  OR2X1 U7444 ( .IN1(n5464), .IN2(n3898), .Q(n6660) );
  OR2X1 U7445 ( .IN1(n6661), .IN2(n6662), .Q(n6656) );
  AND2X1 U7446 ( .IN1(n4839), .IN2(n6663), .Q(n6662) );
  AND2X1 U7447 ( .IN1(n4935), .IN2(n6278), .Q(n6661) );
  XNOR2X1 U7448 ( .IN1(n6664), .IN2(n6665), .Q(n6278) );
  XOR2X1 U7449 ( .IN1(n4202), .IN2(n5388), .Q(n6665) );
  XOR2X1 U7450 ( .IN1(n6666), .IN2(n4605), .Q(n6664) );
  XOR2X1 U7451 ( .IN1(WX8555), .IN2(n9572), .Q(n6666) );
  OR2X1 U7452 ( .IN1(n6667), .IN2(n6668), .Q(WX7131) );
  OR2X1 U7453 ( .IN1(n6669), .IN2(n6670), .Q(n6668) );
  AND2X1 U7454 ( .IN1(n4904), .IN2(CRC_OUT_4_20), .Q(n6670) );
  AND2X1 U7455 ( .IN1(n292), .IN2(n4877), .Q(n6669) );
  INVX0 U7456 ( .INP(n6671), .ZN(n292) );
  OR2X1 U7457 ( .IN1(n5464), .IN2(n3899), .Q(n6671) );
  OR2X1 U7458 ( .IN1(n6672), .IN2(n6673), .Q(n6667) );
  AND2X1 U7459 ( .IN1(n4838), .IN2(n6674), .Q(n6673) );
  AND2X1 U7460 ( .IN1(n4935), .IN2(n6289), .Q(n6672) );
  XNOR2X1 U7461 ( .IN1(n6675), .IN2(n6676), .Q(n6289) );
  XOR2X1 U7462 ( .IN1(n4203), .IN2(n5388), .Q(n6676) );
  XOR2X1 U7463 ( .IN1(n6677), .IN2(n4604), .Q(n6675) );
  XOR2X1 U7464 ( .IN1(WX8553), .IN2(n9573), .Q(n6677) );
  OR2X1 U7465 ( .IN1(n6678), .IN2(n6679), .Q(WX7129) );
  OR2X1 U7466 ( .IN1(n6680), .IN2(n6681), .Q(n6679) );
  AND2X1 U7467 ( .IN1(n4904), .IN2(CRC_OUT_4_21), .Q(n6681) );
  AND2X1 U7468 ( .IN1(n291), .IN2(n4877), .Q(n6680) );
  INVX0 U7469 ( .INP(n6682), .ZN(n291) );
  OR2X1 U7470 ( .IN1(n5464), .IN2(n3900), .Q(n6682) );
  OR2X1 U7471 ( .IN1(n6683), .IN2(n6684), .Q(n6678) );
  AND2X1 U7472 ( .IN1(n6685), .IN2(n4836), .Q(n6684) );
  AND2X1 U7473 ( .IN1(n4935), .IN2(n6300), .Q(n6683) );
  XNOR2X1 U7474 ( .IN1(n6686), .IN2(n6687), .Q(n6300) );
  XOR2X1 U7475 ( .IN1(n4204), .IN2(n5388), .Q(n6687) );
  XOR2X1 U7476 ( .IN1(n6688), .IN2(n4603), .Q(n6686) );
  XOR2X1 U7477 ( .IN1(WX8551), .IN2(n9574), .Q(n6688) );
  OR2X1 U7478 ( .IN1(n6689), .IN2(n6690), .Q(WX7127) );
  OR2X1 U7479 ( .IN1(n6691), .IN2(n6692), .Q(n6690) );
  AND2X1 U7480 ( .IN1(n4904), .IN2(CRC_OUT_4_22), .Q(n6692) );
  AND2X1 U7481 ( .IN1(n290), .IN2(n4877), .Q(n6691) );
  INVX0 U7482 ( .INP(n6693), .ZN(n290) );
  OR2X1 U7483 ( .IN1(n5464), .IN2(n3901), .Q(n6693) );
  OR2X1 U7484 ( .IN1(n6694), .IN2(n6695), .Q(n6689) );
  AND2X1 U7485 ( .IN1(n4838), .IN2(n6696), .Q(n6695) );
  AND2X1 U7486 ( .IN1(n4935), .IN2(n6311), .Q(n6694) );
  XNOR2X1 U7487 ( .IN1(n6697), .IN2(n6698), .Q(n6311) );
  XOR2X1 U7488 ( .IN1(n4205), .IN2(n5388), .Q(n6698) );
  XOR2X1 U7489 ( .IN1(n6699), .IN2(n4602), .Q(n6697) );
  XOR2X1 U7490 ( .IN1(WX8549), .IN2(n9575), .Q(n6699) );
  OR2X1 U7491 ( .IN1(n6700), .IN2(n6701), .Q(WX7125) );
  OR2X1 U7492 ( .IN1(n6702), .IN2(n6703), .Q(n6701) );
  AND2X1 U7493 ( .IN1(n4904), .IN2(CRC_OUT_4_23), .Q(n6703) );
  AND2X1 U7494 ( .IN1(n289), .IN2(n4877), .Q(n6702) );
  INVX0 U7495 ( .INP(n6704), .ZN(n289) );
  OR2X1 U7496 ( .IN1(n5464), .IN2(n3902), .Q(n6704) );
  OR2X1 U7497 ( .IN1(n6705), .IN2(n6706), .Q(n6700) );
  AND2X1 U7498 ( .IN1(n6707), .IN2(n4837), .Q(n6706) );
  AND2X1 U7499 ( .IN1(n4935), .IN2(n6322), .Q(n6705) );
  XNOR2X1 U7500 ( .IN1(n6708), .IN2(n6709), .Q(n6322) );
  XOR2X1 U7501 ( .IN1(n4206), .IN2(n5388), .Q(n6709) );
  XOR2X1 U7502 ( .IN1(n6710), .IN2(n4601), .Q(n6708) );
  XOR2X1 U7503 ( .IN1(WX8547), .IN2(n9576), .Q(n6710) );
  OR2X1 U7504 ( .IN1(n6711), .IN2(n6712), .Q(WX7123) );
  OR2X1 U7505 ( .IN1(n6713), .IN2(n6714), .Q(n6712) );
  AND2X1 U7506 ( .IN1(n4904), .IN2(CRC_OUT_4_24), .Q(n6714) );
  AND2X1 U7507 ( .IN1(n288), .IN2(n4877), .Q(n6713) );
  INVX0 U7508 ( .INP(n6715), .ZN(n288) );
  OR2X1 U7509 ( .IN1(n5463), .IN2(n3903), .Q(n6715) );
  OR2X1 U7510 ( .IN1(n6716), .IN2(n6717), .Q(n6711) );
  AND2X1 U7511 ( .IN1(n4838), .IN2(n6718), .Q(n6717) );
  AND2X1 U7512 ( .IN1(n4935), .IN2(n6333), .Q(n6716) );
  XNOR2X1 U7513 ( .IN1(n6719), .IN2(n6720), .Q(n6333) );
  XOR2X1 U7514 ( .IN1(n4207), .IN2(n5388), .Q(n6720) );
  XOR2X1 U7515 ( .IN1(n6721), .IN2(n4600), .Q(n6719) );
  XOR2X1 U7516 ( .IN1(WX8545), .IN2(n9577), .Q(n6721) );
  OR2X1 U7517 ( .IN1(n6722), .IN2(n6723), .Q(WX7121) );
  OR2X1 U7518 ( .IN1(n6724), .IN2(n6725), .Q(n6723) );
  AND2X1 U7519 ( .IN1(n4905), .IN2(CRC_OUT_4_25), .Q(n6725) );
  AND2X1 U7520 ( .IN1(n287), .IN2(n4876), .Q(n6724) );
  INVX0 U7521 ( .INP(n6726), .ZN(n287) );
  OR2X1 U7522 ( .IN1(n5463), .IN2(n3904), .Q(n6726) );
  OR2X1 U7523 ( .IN1(n6727), .IN2(n6728), .Q(n6722) );
  AND2X1 U7524 ( .IN1(n6729), .IN2(n4837), .Q(n6728) );
  AND2X1 U7525 ( .IN1(n4935), .IN2(n6344), .Q(n6727) );
  XNOR2X1 U7526 ( .IN1(n6730), .IN2(n6731), .Q(n6344) );
  XOR2X1 U7527 ( .IN1(n4208), .IN2(n5387), .Q(n6731) );
  XOR2X1 U7528 ( .IN1(n6732), .IN2(n4599), .Q(n6730) );
  XOR2X1 U7529 ( .IN1(WX8543), .IN2(n9578), .Q(n6732) );
  OR2X1 U7530 ( .IN1(n6733), .IN2(n6734), .Q(WX7119) );
  OR2X1 U7531 ( .IN1(n6735), .IN2(n6736), .Q(n6734) );
  AND2X1 U7532 ( .IN1(n4905), .IN2(CRC_OUT_4_26), .Q(n6736) );
  AND2X1 U7533 ( .IN1(n286), .IN2(n4876), .Q(n6735) );
  INVX0 U7534 ( .INP(n6737), .ZN(n286) );
  OR2X1 U7535 ( .IN1(n5463), .IN2(n3905), .Q(n6737) );
  OR2X1 U7536 ( .IN1(n6738), .IN2(n6739), .Q(n6733) );
  AND2X1 U7537 ( .IN1(n4839), .IN2(n6740), .Q(n6739) );
  AND2X1 U7538 ( .IN1(n6355), .IN2(n4919), .Q(n6738) );
  XOR2X1 U7539 ( .IN1(n6741), .IN2(n6742), .Q(n6355) );
  XOR2X1 U7540 ( .IN1(n4209), .IN2(n5387), .Q(n6742) );
  XOR2X1 U7541 ( .IN1(WX8477), .IN2(n6743), .Q(n6741) );
  XOR2X1 U7542 ( .IN1(test_so74), .IN2(n9579), .Q(n6743) );
  OR2X1 U7543 ( .IN1(n6744), .IN2(n6745), .Q(WX7117) );
  OR2X1 U7544 ( .IN1(n6746), .IN2(n6747), .Q(n6745) );
  AND2X1 U7545 ( .IN1(n4905), .IN2(CRC_OUT_4_27), .Q(n6747) );
  AND2X1 U7546 ( .IN1(n285), .IN2(n4876), .Q(n6746) );
  INVX0 U7547 ( .INP(n6748), .ZN(n285) );
  OR2X1 U7548 ( .IN1(n5463), .IN2(n3906), .Q(n6748) );
  OR2X1 U7549 ( .IN1(n6749), .IN2(n6750), .Q(n6744) );
  AND2X1 U7550 ( .IN1(n6751), .IN2(n4838), .Q(n6750) );
  AND2X1 U7551 ( .IN1(n4935), .IN2(n6366), .Q(n6749) );
  XNOR2X1 U7552 ( .IN1(n6752), .IN2(n6753), .Q(n6366) );
  XOR2X1 U7553 ( .IN1(n4210), .IN2(n5387), .Q(n6753) );
  XOR2X1 U7554 ( .IN1(n6754), .IN2(n4598), .Q(n6752) );
  XOR2X1 U7555 ( .IN1(WX8539), .IN2(n9580), .Q(n6754) );
  OR2X1 U7556 ( .IN1(n6755), .IN2(n6756), .Q(WX7115) );
  OR2X1 U7557 ( .IN1(n6757), .IN2(n6758), .Q(n6756) );
  AND2X1 U7558 ( .IN1(n4905), .IN2(CRC_OUT_4_28), .Q(n6758) );
  AND2X1 U7559 ( .IN1(n284), .IN2(n4876), .Q(n6757) );
  INVX0 U7560 ( .INP(n6759), .ZN(n284) );
  OR2X1 U7561 ( .IN1(n5463), .IN2(n3907), .Q(n6759) );
  OR2X1 U7562 ( .IN1(n6760), .IN2(n6761), .Q(n6755) );
  AND2X1 U7563 ( .IN1(n4839), .IN2(n6762), .Q(n6761) );
  AND2X1 U7564 ( .IN1(n6377), .IN2(n4919), .Q(n6760) );
  XOR2X1 U7565 ( .IN1(n6763), .IN2(n6764), .Q(n6377) );
  XOR2X1 U7566 ( .IN1(n4597), .IN2(n5387), .Q(n6764) );
  XOR2X1 U7567 ( .IN1(n6765), .IN2(n9583), .Q(n6763) );
  XOR2X1 U7568 ( .IN1(n9582), .IN2(n9581), .Q(n6765) );
  OR2X1 U7569 ( .IN1(n6766), .IN2(n6767), .Q(WX7113) );
  OR2X1 U7570 ( .IN1(n6768), .IN2(n6769), .Q(n6767) );
  AND2X1 U7571 ( .IN1(test_so66), .IN2(n4887), .Q(n6769) );
  AND2X1 U7572 ( .IN1(n283), .IN2(n4876), .Q(n6768) );
  INVX0 U7573 ( .INP(n6770), .ZN(n283) );
  OR2X1 U7574 ( .IN1(n5463), .IN2(n3908), .Q(n6770) );
  OR2X1 U7575 ( .IN1(n6771), .IN2(n6772), .Q(n6766) );
  AND2X1 U7576 ( .IN1(n4839), .IN2(n6773), .Q(n6772) );
  AND2X1 U7577 ( .IN1(n4935), .IN2(n6388), .Q(n6771) );
  XNOR2X1 U7578 ( .IN1(n6774), .IN2(n6775), .Q(n6388) );
  XOR2X1 U7579 ( .IN1(n4211), .IN2(n5387), .Q(n6775) );
  XOR2X1 U7580 ( .IN1(n6776), .IN2(n4596), .Q(n6774) );
  XOR2X1 U7581 ( .IN1(WX8535), .IN2(n9584), .Q(n6776) );
  OR2X1 U7582 ( .IN1(n6777), .IN2(n6778), .Q(WX7111) );
  OR2X1 U7583 ( .IN1(n6779), .IN2(n6780), .Q(n6778) );
  AND2X1 U7584 ( .IN1(n4905), .IN2(CRC_OUT_4_30), .Q(n6780) );
  AND2X1 U7585 ( .IN1(n282), .IN2(n4876), .Q(n6779) );
  INVX0 U7586 ( .INP(n6781), .ZN(n282) );
  OR2X1 U7587 ( .IN1(n5463), .IN2(n3909), .Q(n6781) );
  OR2X1 U7588 ( .IN1(n6782), .IN2(n6783), .Q(n6777) );
  AND2X1 U7589 ( .IN1(n4839), .IN2(n6784), .Q(n6783) );
  AND2X1 U7590 ( .IN1(n6399), .IN2(n4919), .Q(n6782) );
  XOR2X1 U7591 ( .IN1(n6785), .IN2(n6786), .Q(n6399) );
  XOR2X1 U7592 ( .IN1(n4595), .IN2(n5387), .Q(n6786) );
  XOR2X1 U7593 ( .IN1(n6787), .IN2(n9587), .Q(n6785) );
  XOR2X1 U7594 ( .IN1(n9586), .IN2(n9585), .Q(n6787) );
  OR2X1 U7595 ( .IN1(n6788), .IN2(n6789), .Q(WX7109) );
  OR2X1 U7596 ( .IN1(n6790), .IN2(n6791), .Q(n6789) );
  AND2X1 U7597 ( .IN1(n2245), .IN2(WX6950), .Q(n6791) );
  AND2X1 U7598 ( .IN1(n4905), .IN2(CRC_OUT_4_31), .Q(n6790) );
  OR2X1 U7599 ( .IN1(n6792), .IN2(n6793), .Q(n6788) );
  AND2X1 U7600 ( .IN1(n4839), .IN2(n6794), .Q(n6793) );
  AND2X1 U7601 ( .IN1(n4935), .IN2(n6409), .Q(n6792) );
  XNOR2X1 U7602 ( .IN1(n6795), .IN2(n6796), .Q(n6409) );
  XOR2X1 U7603 ( .IN1(n4167), .IN2(n5387), .Q(n6796) );
  XOR2X1 U7604 ( .IN1(n6797), .IN2(n4594), .Q(n6795) );
  XOR2X1 U7605 ( .IN1(WX8531), .IN2(n9588), .Q(n6797) );
  OR2X1 U7606 ( .IN1(n6798), .IN2(n6799), .Q(WX706) );
  OR2X1 U7607 ( .IN1(n6800), .IN2(n6801), .Q(n6799) );
  AND2X1 U7608 ( .IN1(n4905), .IN2(CRC_OUT_9_0), .Q(n6801) );
  AND2X1 U7609 ( .IN1(WX544), .IN2(n4876), .Q(n6800) );
  OR2X1 U7610 ( .IN1(n6802), .IN2(n6803), .Q(n6798) );
  AND2X1 U7611 ( .IN1(n4839), .IN2(n6804), .Q(n6803) );
  AND2X1 U7612 ( .IN1(n6805), .IN2(n4919), .Q(n6802) );
  OR2X1 U7613 ( .IN1(n6806), .IN2(n6807), .Q(WX704) );
  OR2X1 U7614 ( .IN1(n6808), .IN2(n6809), .Q(n6807) );
  AND2X1 U7615 ( .IN1(test_so9), .IN2(n4888), .Q(n6809) );
  AND2X1 U7616 ( .IN1(WX542), .IN2(n4876), .Q(n6808) );
  OR2X1 U7617 ( .IN1(n6810), .IN2(n6811), .Q(n6806) );
  AND2X1 U7618 ( .IN1(n4839), .IN2(n6812), .Q(n6811) );
  AND2X1 U7619 ( .IN1(n4935), .IN2(n6813), .Q(n6810) );
  OR2X1 U7620 ( .IN1(n6814), .IN2(n6815), .Q(WX702) );
  OR2X1 U7621 ( .IN1(n6816), .IN2(n6817), .Q(n6815) );
  AND2X1 U7622 ( .IN1(n4905), .IN2(CRC_OUT_9_2), .Q(n6817) );
  AND2X1 U7623 ( .IN1(WX540), .IN2(n4876), .Q(n6816) );
  OR2X1 U7624 ( .IN1(n6818), .IN2(n6819), .Q(n6814) );
  AND2X1 U7625 ( .IN1(n6820), .IN2(n4836), .Q(n6819) );
  AND2X1 U7626 ( .IN1(n4935), .IN2(n6821), .Q(n6818) );
  AND2X1 U7627 ( .IN1(n4823), .IN2(n5401), .Q(WX7011) );
  OR2X1 U7628 ( .IN1(n6822), .IN2(n6823), .Q(WX700) );
  OR2X1 U7629 ( .IN1(n6824), .IN2(n6825), .Q(n6823) );
  AND2X1 U7630 ( .IN1(n4905), .IN2(CRC_OUT_9_3), .Q(n6825) );
  AND2X1 U7631 ( .IN1(WX538), .IN2(n4876), .Q(n6824) );
  OR2X1 U7632 ( .IN1(n6826), .IN2(n6827), .Q(n6822) );
  AND2X1 U7633 ( .IN1(n4839), .IN2(n6828), .Q(n6827) );
  AND2X1 U7634 ( .IN1(n4935), .IN2(n6829), .Q(n6826) );
  AND2X1 U7635 ( .IN1(n6413), .IN2(n8443), .Q(WX6999) );
  OR2X1 U7636 ( .IN1(n6830), .IN2(n6831), .Q(WX698) );
  OR2X1 U7637 ( .IN1(n6832), .IN2(n6833), .Q(n6831) );
  AND2X1 U7638 ( .IN1(n4905), .IN2(CRC_OUT_9_4), .Q(n6833) );
  AND2X1 U7639 ( .IN1(WX536), .IN2(n4876), .Q(n6832) );
  OR2X1 U7640 ( .IN1(n6834), .IN2(n6835), .Q(n6830) );
  AND2X1 U7641 ( .IN1(n4839), .IN2(n6836), .Q(n6835) );
  AND2X1 U7642 ( .IN1(n6837), .IN2(n4919), .Q(n6834) );
  OR2X1 U7643 ( .IN1(n6838), .IN2(n6839), .Q(WX696) );
  OR2X1 U7644 ( .IN1(n6840), .IN2(n6841), .Q(n6839) );
  AND2X1 U7645 ( .IN1(n4905), .IN2(CRC_OUT_9_5), .Q(n6841) );
  AND2X1 U7646 ( .IN1(WX534), .IN2(n4876), .Q(n6840) );
  OR2X1 U7647 ( .IN1(n6842), .IN2(n6843), .Q(n6838) );
  AND2X1 U7648 ( .IN1(n4839), .IN2(n6844), .Q(n6843) );
  AND2X1 U7649 ( .IN1(n4936), .IN2(n6845), .Q(n6842) );
  OR2X1 U7650 ( .IN1(n6846), .IN2(n6847), .Q(WX694) );
  OR2X1 U7651 ( .IN1(n6848), .IN2(n6849), .Q(n6847) );
  AND2X1 U7652 ( .IN1(n4905), .IN2(CRC_OUT_9_6), .Q(n6849) );
  AND2X1 U7653 ( .IN1(WX532), .IN2(n4875), .Q(n6848) );
  OR2X1 U7654 ( .IN1(n6850), .IN2(n6851), .Q(n6846) );
  AND2X1 U7655 ( .IN1(n6852), .IN2(n4836), .Q(n6851) );
  AND2X1 U7656 ( .IN1(n4936), .IN2(n6853), .Q(n6850) );
  OR2X1 U7657 ( .IN1(n6854), .IN2(n6855), .Q(WX692) );
  OR2X1 U7658 ( .IN1(n6856), .IN2(n6857), .Q(n6855) );
  AND2X1 U7659 ( .IN1(n4905), .IN2(CRC_OUT_9_7), .Q(n6857) );
  AND2X1 U7660 ( .IN1(WX530), .IN2(n4875), .Q(n6856) );
  OR2X1 U7661 ( .IN1(n6858), .IN2(n6859), .Q(n6854) );
  AND2X1 U7662 ( .IN1(n4839), .IN2(n6860), .Q(n6859) );
  AND2X1 U7663 ( .IN1(n4936), .IN2(n6861), .Q(n6858) );
  OR2X1 U7664 ( .IN1(n6862), .IN2(n6863), .Q(WX690) );
  OR2X1 U7665 ( .IN1(n6864), .IN2(n6865), .Q(n6863) );
  AND2X1 U7666 ( .IN1(n4906), .IN2(CRC_OUT_9_8), .Q(n6865) );
  AND2X1 U7667 ( .IN1(WX528), .IN2(n4875), .Q(n6864) );
  OR2X1 U7668 ( .IN1(n6866), .IN2(n6867), .Q(n6862) );
  AND2X1 U7669 ( .IN1(n4840), .IN2(n6868), .Q(n6867) );
  AND2X1 U7670 ( .IN1(n4936), .IN2(n6869), .Q(n6866) );
  OR2X1 U7671 ( .IN1(n6870), .IN2(n6871), .Q(WX688) );
  OR2X1 U7672 ( .IN1(n6872), .IN2(n6873), .Q(n6871) );
  AND2X1 U7673 ( .IN1(n4906), .IN2(CRC_OUT_9_9), .Q(n6873) );
  AND2X1 U7674 ( .IN1(WX526), .IN2(n4875), .Q(n6872) );
  OR2X1 U7675 ( .IN1(n6874), .IN2(n6875), .Q(n6870) );
  AND2X1 U7676 ( .IN1(n4840), .IN2(n6876), .Q(n6875) );
  AND2X1 U7677 ( .IN1(n4936), .IN2(n6877), .Q(n6874) );
  OR2X1 U7678 ( .IN1(n6878), .IN2(n6879), .Q(WX686) );
  OR2X1 U7679 ( .IN1(n6880), .IN2(n6881), .Q(n6879) );
  AND2X1 U7680 ( .IN1(n4906), .IN2(CRC_OUT_9_10), .Q(n6881) );
  AND2X1 U7681 ( .IN1(WX524), .IN2(n4875), .Q(n6880) );
  OR2X1 U7682 ( .IN1(n6882), .IN2(n6883), .Q(n6878) );
  AND2X1 U7683 ( .IN1(n6884), .IN2(n4835), .Q(n6883) );
  AND2X1 U7684 ( .IN1(n6885), .IN2(n4918), .Q(n6882) );
  OR2X1 U7685 ( .IN1(n6886), .IN2(n6887), .Q(WX684) );
  OR2X1 U7686 ( .IN1(n6888), .IN2(n6889), .Q(n6887) );
  AND2X1 U7687 ( .IN1(n4906), .IN2(CRC_OUT_9_11), .Q(n6889) );
  AND2X1 U7688 ( .IN1(WX522), .IN2(n4875), .Q(n6888) );
  OR2X1 U7689 ( .IN1(n6890), .IN2(n6891), .Q(n6886) );
  AND2X1 U7690 ( .IN1(n4840), .IN2(n6892), .Q(n6891) );
  AND2X1 U7691 ( .IN1(n4936), .IN2(n6893), .Q(n6890) );
  OR2X1 U7692 ( .IN1(n6894), .IN2(n6895), .Q(WX682) );
  OR2X1 U7693 ( .IN1(n6896), .IN2(n6897), .Q(n6895) );
  AND2X1 U7694 ( .IN1(n4906), .IN2(CRC_OUT_9_12), .Q(n6897) );
  AND2X1 U7695 ( .IN1(WX520), .IN2(n4875), .Q(n6896) );
  OR2X1 U7696 ( .IN1(n6898), .IN2(n6899), .Q(n6894) );
  AND2X1 U7697 ( .IN1(n4840), .IN2(n6900), .Q(n6899) );
  AND2X1 U7698 ( .IN1(n4936), .IN2(n6901), .Q(n6898) );
  OR2X1 U7699 ( .IN1(n6902), .IN2(n6903), .Q(WX680) );
  OR2X1 U7700 ( .IN1(n6904), .IN2(n6905), .Q(n6903) );
  AND2X1 U7701 ( .IN1(n4906), .IN2(CRC_OUT_9_13), .Q(n6905) );
  AND2X1 U7702 ( .IN1(WX518), .IN2(n4875), .Q(n6904) );
  OR2X1 U7703 ( .IN1(n6906), .IN2(n6907), .Q(n6902) );
  AND2X1 U7704 ( .IN1(n4840), .IN2(n6908), .Q(n6907) );
  AND2X1 U7705 ( .IN1(n4936), .IN2(n6909), .Q(n6906) );
  OR2X1 U7706 ( .IN1(n6910), .IN2(n6911), .Q(WX678) );
  OR2X1 U7707 ( .IN1(n6912), .IN2(n6913), .Q(n6911) );
  AND2X1 U7708 ( .IN1(n4906), .IN2(CRC_OUT_9_14), .Q(n6913) );
  AND2X1 U7709 ( .IN1(WX516), .IN2(n4875), .Q(n6912) );
  OR2X1 U7710 ( .IN1(n6914), .IN2(n6915), .Q(n6910) );
  AND2X1 U7711 ( .IN1(n4840), .IN2(n6916), .Q(n6915) );
  AND2X1 U7712 ( .IN1(n6917), .IN2(n4918), .Q(n6914) );
  OR2X1 U7713 ( .IN1(n6918), .IN2(n6919), .Q(WX676) );
  OR2X1 U7714 ( .IN1(n6920), .IN2(n6921), .Q(n6919) );
  AND2X1 U7715 ( .IN1(n4906), .IN2(CRC_OUT_9_15), .Q(n6921) );
  AND2X1 U7716 ( .IN1(WX514), .IN2(n4875), .Q(n6920) );
  OR2X1 U7717 ( .IN1(n6922), .IN2(n6923), .Q(n6918) );
  AND2X1 U7718 ( .IN1(n4840), .IN2(n6924), .Q(n6923) );
  AND2X1 U7719 ( .IN1(n4936), .IN2(n6925), .Q(n6922) );
  OR2X1 U7720 ( .IN1(n6926), .IN2(n6927), .Q(WX674) );
  OR2X1 U7721 ( .IN1(n6928), .IN2(n6929), .Q(n6927) );
  AND2X1 U7722 ( .IN1(n4906), .IN2(CRC_OUT_9_16), .Q(n6929) );
  AND2X1 U7723 ( .IN1(WX512), .IN2(n4875), .Q(n6928) );
  OR2X1 U7724 ( .IN1(n6930), .IN2(n6931), .Q(n6926) );
  AND2X1 U7725 ( .IN1(n6932), .IN2(n4835), .Q(n6931) );
  AND2X1 U7726 ( .IN1(n4936), .IN2(n6933), .Q(n6930) );
  OR2X1 U7727 ( .IN1(n6934), .IN2(n6935), .Q(WX672) );
  OR2X1 U7728 ( .IN1(n6936), .IN2(n6937), .Q(n6935) );
  AND2X1 U7729 ( .IN1(n4906), .IN2(CRC_OUT_9_17), .Q(n6937) );
  AND2X1 U7730 ( .IN1(WX510), .IN2(n4875), .Q(n6936) );
  OR2X1 U7731 ( .IN1(n6938), .IN2(n6939), .Q(n6934) );
  AND2X1 U7732 ( .IN1(n4840), .IN2(n6940), .Q(n6939) );
  AND2X1 U7733 ( .IN1(n4936), .IN2(n6941), .Q(n6938) );
  OR2X1 U7734 ( .IN1(n6942), .IN2(n6943), .Q(WX670) );
  OR2X1 U7735 ( .IN1(n6944), .IN2(n6945), .Q(n6943) );
  AND2X1 U7736 ( .IN1(n4906), .IN2(CRC_OUT_9_18), .Q(n6945) );
  AND2X1 U7737 ( .IN1(WX508), .IN2(n4874), .Q(n6944) );
  OR2X1 U7738 ( .IN1(n6946), .IN2(n6947), .Q(n6942) );
  AND2X1 U7739 ( .IN1(n4840), .IN2(n6948), .Q(n6947) );
  AND2X1 U7740 ( .IN1(n6949), .IN2(n4918), .Q(n6946) );
  OR2X1 U7741 ( .IN1(n6950), .IN2(n6951), .Q(WX668) );
  OR2X1 U7742 ( .IN1(n6952), .IN2(n6953), .Q(n6951) );
  AND2X1 U7743 ( .IN1(test_so10), .IN2(n4887), .Q(n6953) );
  AND2X1 U7744 ( .IN1(WX506), .IN2(n4874), .Q(n6952) );
  OR2X1 U7745 ( .IN1(n6954), .IN2(n6955), .Q(n6950) );
  AND2X1 U7746 ( .IN1(n4840), .IN2(n6956), .Q(n6955) );
  AND2X1 U7747 ( .IN1(n4936), .IN2(n6957), .Q(n6954) );
  OR2X1 U7748 ( .IN1(n6958), .IN2(n6959), .Q(WX666) );
  OR2X1 U7749 ( .IN1(n6960), .IN2(n6961), .Q(n6959) );
  AND2X1 U7750 ( .IN1(n4906), .IN2(CRC_OUT_9_20), .Q(n6961) );
  AND2X1 U7751 ( .IN1(WX504), .IN2(n4874), .Q(n6960) );
  OR2X1 U7752 ( .IN1(n6962), .IN2(n6963), .Q(n6958) );
  AND2X1 U7753 ( .IN1(n6964), .IN2(n4834), .Q(n6963) );
  AND2X1 U7754 ( .IN1(n4936), .IN2(n6965), .Q(n6962) );
  OR2X1 U7755 ( .IN1(n6966), .IN2(n6967), .Q(WX664) );
  OR2X1 U7756 ( .IN1(n6968), .IN2(n6969), .Q(n6967) );
  AND2X1 U7757 ( .IN1(n4906), .IN2(CRC_OUT_9_21), .Q(n6969) );
  AND2X1 U7758 ( .IN1(WX502), .IN2(n4874), .Q(n6968) );
  OR2X1 U7759 ( .IN1(n6970), .IN2(n6971), .Q(n6966) );
  AND2X1 U7760 ( .IN1(n4840), .IN2(n6972), .Q(n6971) );
  AND2X1 U7761 ( .IN1(n4937), .IN2(n6973), .Q(n6970) );
  OR2X1 U7762 ( .IN1(n6974), .IN2(n6975), .Q(WX662) );
  OR2X1 U7763 ( .IN1(n6976), .IN2(n6977), .Q(n6975) );
  AND2X1 U7764 ( .IN1(n4907), .IN2(CRC_OUT_9_22), .Q(n6977) );
  AND2X1 U7765 ( .IN1(WX500), .IN2(n4874), .Q(n6976) );
  OR2X1 U7766 ( .IN1(n6978), .IN2(n6979), .Q(n6974) );
  AND2X1 U7767 ( .IN1(n4840), .IN2(n6980), .Q(n6979) );
  AND2X1 U7768 ( .IN1(n6981), .IN2(n4918), .Q(n6978) );
  OR2X1 U7769 ( .IN1(n6982), .IN2(n6983), .Q(WX660) );
  OR2X1 U7770 ( .IN1(n6984), .IN2(n6985), .Q(n6983) );
  AND2X1 U7771 ( .IN1(n4907), .IN2(CRC_OUT_9_23), .Q(n6985) );
  AND2X1 U7772 ( .IN1(WX498), .IN2(n4874), .Q(n6984) );
  OR2X1 U7773 ( .IN1(n6986), .IN2(n6987), .Q(n6982) );
  AND2X1 U7774 ( .IN1(n4840), .IN2(n6988), .Q(n6987) );
  AND2X1 U7775 ( .IN1(n4937), .IN2(n6989), .Q(n6986) );
  OR2X1 U7776 ( .IN1(n6990), .IN2(n6991), .Q(WX658) );
  OR2X1 U7777 ( .IN1(n6992), .IN2(n6993), .Q(n6991) );
  AND2X1 U7778 ( .IN1(n4907), .IN2(CRC_OUT_9_24), .Q(n6993) );
  AND2X1 U7779 ( .IN1(WX496), .IN2(n4874), .Q(n6992) );
  OR2X1 U7780 ( .IN1(n6994), .IN2(n6995), .Q(n6990) );
  AND2X1 U7781 ( .IN1(n6996), .IN2(n4834), .Q(n6995) );
  AND2X1 U7782 ( .IN1(n4937), .IN2(n6997), .Q(n6994) );
  OR2X1 U7783 ( .IN1(n6998), .IN2(n6999), .Q(WX656) );
  OR2X1 U7784 ( .IN1(n7000), .IN2(n7001), .Q(n6999) );
  AND2X1 U7785 ( .IN1(n4907), .IN2(CRC_OUT_9_25), .Q(n7001) );
  AND2X1 U7786 ( .IN1(WX494), .IN2(n4874), .Q(n7000) );
  OR2X1 U7787 ( .IN1(n7002), .IN2(n7003), .Q(n6998) );
  AND2X1 U7788 ( .IN1(n4841), .IN2(n7004), .Q(n7003) );
  AND2X1 U7789 ( .IN1(n4937), .IN2(n7005), .Q(n7002) );
  OR2X1 U7790 ( .IN1(n7006), .IN2(n7007), .Q(WX654) );
  OR2X1 U7791 ( .IN1(n7008), .IN2(n7009), .Q(n7007) );
  AND2X1 U7792 ( .IN1(n4907), .IN2(CRC_OUT_9_26), .Q(n7009) );
  AND2X1 U7793 ( .IN1(WX492), .IN2(n4874), .Q(n7008) );
  OR2X1 U7794 ( .IN1(n7010), .IN2(n7011), .Q(n7006) );
  AND2X1 U7795 ( .IN1(n4841), .IN2(n7012), .Q(n7011) );
  AND2X1 U7796 ( .IN1(n4937), .IN2(n7013), .Q(n7010) );
  OR2X1 U7797 ( .IN1(n7014), .IN2(n7015), .Q(WX652) );
  OR2X1 U7798 ( .IN1(n7016), .IN2(n7017), .Q(n7015) );
  AND2X1 U7799 ( .IN1(n4907), .IN2(CRC_OUT_9_27), .Q(n7017) );
  AND2X1 U7800 ( .IN1(WX490), .IN2(n4874), .Q(n7016) );
  OR2X1 U7801 ( .IN1(n7018), .IN2(n7019), .Q(n7014) );
  AND2X1 U7802 ( .IN1(n4841), .IN2(n7020), .Q(n7019) );
  AND2X1 U7803 ( .IN1(n4937), .IN2(n7021), .Q(n7018) );
  OR2X1 U7804 ( .IN1(n7022), .IN2(n7023), .Q(WX650) );
  OR2X1 U7805 ( .IN1(n7024), .IN2(n7025), .Q(n7023) );
  AND2X1 U7806 ( .IN1(n4907), .IN2(CRC_OUT_9_28), .Q(n7025) );
  AND2X1 U7807 ( .IN1(WX488), .IN2(n4874), .Q(n7024) );
  OR2X1 U7808 ( .IN1(n7026), .IN2(n7027), .Q(n7022) );
  AND2X1 U7809 ( .IN1(n7028), .IN2(n4833), .Q(n7027) );
  AND2X1 U7810 ( .IN1(n7029), .IN2(n4918), .Q(n7026) );
  AND2X1 U7811 ( .IN1(n7030), .IN2(n5401), .Q(WX6498) );
  XOR2X1 U7812 ( .IN1(CRC_OUT_5_30), .IN2(n4647), .Q(n7030) );
  AND2X1 U7813 ( .IN1(n7031), .IN2(n5401), .Q(WX6496) );
  XOR2X1 U7814 ( .IN1(CRC_OUT_5_29), .IN2(n4648), .Q(n7031) );
  AND2X1 U7815 ( .IN1(n7032), .IN2(n5402), .Q(WX6494) );
  XOR2X1 U7816 ( .IN1(CRC_OUT_5_28), .IN2(n4649), .Q(n7032) );
  AND2X1 U7817 ( .IN1(n7033), .IN2(n5402), .Q(WX6492) );
  XOR2X1 U7818 ( .IN1(CRC_OUT_5_27), .IN2(n4650), .Q(n7033) );
  AND2X1 U7819 ( .IN1(n7034), .IN2(n5402), .Q(WX6490) );
  XOR2X1 U7820 ( .IN1(CRC_OUT_5_26), .IN2(n4651), .Q(n7034) );
  AND2X1 U7821 ( .IN1(n7035), .IN2(n5402), .Q(WX6488) );
  XOR2X1 U7822 ( .IN1(CRC_OUT_5_25), .IN2(n4652), .Q(n7035) );
  AND2X1 U7823 ( .IN1(n7036), .IN2(n5402), .Q(WX6486) );
  XOR2X1 U7824 ( .IN1(CRC_OUT_5_24), .IN2(n4653), .Q(n7036) );
  AND2X1 U7825 ( .IN1(n7037), .IN2(n6413), .Q(WX6484) );
  INVX0 U7826 ( .INP(n7038), .ZN(n6413) );
  OR2X1 U7827 ( .IN1(Tj_Trigger), .IN2(n5461), .Q(n7038) );
  XOR2X1 U7828 ( .IN1(CRC_OUT_5_23), .IN2(n4654), .Q(n7037) );
  AND2X1 U7829 ( .IN1(n7039), .IN2(n5402), .Q(WX6482) );
  XOR2X1 U7830 ( .IN1(CRC_OUT_5_22), .IN2(n4655), .Q(n7039) );
  AND2X1 U7831 ( .IN1(n7040), .IN2(n5402), .Q(WX6480) );
  XOR2X1 U7832 ( .IN1(CRC_OUT_5_21), .IN2(n4656), .Q(n7040) );
  OR2X1 U7833 ( .IN1(n7041), .IN2(n7042), .Q(WX648) );
  OR2X1 U7834 ( .IN1(n7043), .IN2(n7044), .Q(n7042) );
  AND2X1 U7835 ( .IN1(n4907), .IN2(CRC_OUT_9_29), .Q(n7044) );
  AND2X1 U7836 ( .IN1(WX486), .IN2(n4874), .Q(n7043) );
  OR2X1 U7837 ( .IN1(n7045), .IN2(n7046), .Q(n7041) );
  AND2X1 U7838 ( .IN1(n4841), .IN2(n7047), .Q(n7046) );
  AND2X1 U7839 ( .IN1(n4937), .IN2(n7048), .Q(n7045) );
  AND2X1 U7840 ( .IN1(n7049), .IN2(n5402), .Q(WX6478) );
  XOR2X1 U7841 ( .IN1(CRC_OUT_5_20), .IN2(n4657), .Q(n7049) );
  AND2X1 U7842 ( .IN1(n7050), .IN2(n5402), .Q(WX6476) );
  XOR2X1 U7843 ( .IN1(CRC_OUT_5_19), .IN2(n4658), .Q(n7050) );
  AND2X1 U7844 ( .IN1(n7051), .IN2(n5403), .Q(WX6474) );
  XOR2X1 U7845 ( .IN1(CRC_OUT_5_18), .IN2(n4659), .Q(n7051) );
  AND2X1 U7846 ( .IN1(n7052), .IN2(n5403), .Q(WX6472) );
  XOR2X1 U7847 ( .IN1(test_so54), .IN2(n4660), .Q(n7052) );
  AND2X1 U7848 ( .IN1(n7053), .IN2(n5403), .Q(WX6470) );
  XOR2X1 U7849 ( .IN1(CRC_OUT_5_16), .IN2(n4661), .Q(n7053) );
  AND2X1 U7850 ( .IN1(n7054), .IN2(n5403), .Q(WX6468) );
  XOR2X1 U7851 ( .IN1(CRC_OUT_5_15), .IN2(n7055), .Q(n7054) );
  XOR2X1 U7852 ( .IN1(test_so52), .IN2(DFF_959_n1), .Q(n7055) );
  AND2X1 U7853 ( .IN1(n7056), .IN2(n5403), .Q(WX6466) );
  XOR2X1 U7854 ( .IN1(CRC_OUT_5_14), .IN2(n4662), .Q(n7056) );
  AND2X1 U7855 ( .IN1(n7057), .IN2(n5403), .Q(WX6464) );
  XOR2X1 U7856 ( .IN1(CRC_OUT_5_13), .IN2(n4663), .Q(n7057) );
  AND2X1 U7857 ( .IN1(n7058), .IN2(n5403), .Q(WX6462) );
  XOR2X1 U7858 ( .IN1(CRC_OUT_5_12), .IN2(n4664), .Q(n7058) );
  AND2X1 U7859 ( .IN1(n7059), .IN2(n5403), .Q(WX6460) );
  XOR2X1 U7860 ( .IN1(CRC_OUT_5_11), .IN2(n4665), .Q(n7059) );
  OR2X1 U7861 ( .IN1(n7060), .IN2(n7061), .Q(WX646) );
  OR2X1 U7862 ( .IN1(n7062), .IN2(n7063), .Q(n7061) );
  AND2X1 U7863 ( .IN1(n4907), .IN2(CRC_OUT_9_30), .Q(n7063) );
  AND2X1 U7864 ( .IN1(WX484), .IN2(n4873), .Q(n7062) );
  OR2X1 U7865 ( .IN1(n7064), .IN2(n7065), .Q(n7060) );
  AND2X1 U7866 ( .IN1(n4855), .IN2(n7066), .Q(n7065) );
  AND2X1 U7867 ( .IN1(n4937), .IN2(n7067), .Q(n7064) );
  AND2X1 U7868 ( .IN1(n7068), .IN2(n5403), .Q(WX6458) );
  XOR2X1 U7869 ( .IN1(DFF_938_n1), .IN2(n7069), .Q(n7068) );
  XOR2X1 U7870 ( .IN1(n4524), .IN2(DFF_959_n1), .Q(n7069) );
  AND2X1 U7871 ( .IN1(n7070), .IN2(n5404), .Q(WX6456) );
  XOR2X1 U7872 ( .IN1(CRC_OUT_5_9), .IN2(n4666), .Q(n7070) );
  AND2X1 U7873 ( .IN1(n7071), .IN2(n5404), .Q(WX6454) );
  XOR2X1 U7874 ( .IN1(CRC_OUT_5_8), .IN2(n4667), .Q(n7071) );
  AND2X1 U7875 ( .IN1(n7072), .IN2(n5404), .Q(WX6452) );
  XOR2X1 U7876 ( .IN1(CRC_OUT_5_7), .IN2(n4668), .Q(n7072) );
  AND2X1 U7877 ( .IN1(n7073), .IN2(n5404), .Q(WX6450) );
  XOR2X1 U7878 ( .IN1(CRC_OUT_5_6), .IN2(n4669), .Q(n7073) );
  AND2X1 U7879 ( .IN1(n7074), .IN2(n5404), .Q(WX6448) );
  XOR2X1 U7880 ( .IN1(CRC_OUT_5_5), .IN2(n4670), .Q(n7074) );
  AND2X1 U7881 ( .IN1(n7075), .IN2(n5404), .Q(WX6446) );
  XOR2X1 U7882 ( .IN1(CRC_OUT_5_4), .IN2(n4671), .Q(n7075) );
  AND2X1 U7883 ( .IN1(n7076), .IN2(n5404), .Q(WX6444) );
  XOR2X1 U7884 ( .IN1(DFF_931_n1), .IN2(n7077), .Q(n7076) );
  XOR2X1 U7885 ( .IN1(n4525), .IN2(DFF_959_n1), .Q(n7077) );
  AND2X1 U7886 ( .IN1(n7078), .IN2(n5404), .Q(WX6442) );
  XOR2X1 U7887 ( .IN1(CRC_OUT_5_2), .IN2(n4672), .Q(n7078) );
  AND2X1 U7888 ( .IN1(n7079), .IN2(n5405), .Q(WX6440) );
  XOR2X1 U7889 ( .IN1(CRC_OUT_5_1), .IN2(n4673), .Q(n7079) );
  OR2X1 U7890 ( .IN1(n7080), .IN2(n7081), .Q(WX644) );
  OR2X1 U7891 ( .IN1(n7082), .IN2(n7083), .Q(n7081) );
  AND2X1 U7892 ( .IN1(n2245), .IN2(WX485), .Q(n7083) );
  AND2X1 U7893 ( .IN1(n4907), .IN2(CRC_OUT_9_31), .Q(n7082) );
  OR2X1 U7894 ( .IN1(n7084), .IN2(n7085), .Q(n7080) );
  AND2X1 U7895 ( .IN1(n4855), .IN2(n7086), .Q(n7085) );
  AND2X1 U7896 ( .IN1(n4937), .IN2(n7087), .Q(n7084) );
  AND2X1 U7897 ( .IN1(n7088), .IN2(n5405), .Q(WX6438) );
  XOR2X1 U7898 ( .IN1(test_so53), .IN2(n4674), .Q(n7088) );
  AND2X1 U7899 ( .IN1(n7089), .IN2(n5405), .Q(WX6436) );
  XOR2X1 U7900 ( .IN1(n4538), .IN2(CRC_OUT_5_31), .Q(n7089) );
  INVX0 U7901 ( .INP(n7090), .ZN(WX5910) );
  OR2X1 U7902 ( .IN1(n5463), .IN2(n9640), .Q(n7090) );
  INVX0 U7903 ( .INP(n7091), .ZN(WX5908) );
  OR2X1 U7904 ( .IN1(n5463), .IN2(n9641), .Q(n7091) );
  INVX0 U7905 ( .INP(n7092), .ZN(WX5906) );
  OR2X1 U7906 ( .IN1(n5463), .IN2(n9642), .Q(n7092) );
  INVX0 U7907 ( .INP(n7093), .ZN(WX5904) );
  OR2X1 U7908 ( .IN1(n5463), .IN2(n9645), .Q(n7093) );
  INVX0 U7909 ( .INP(n7094), .ZN(WX5902) );
  OR2X1 U7910 ( .IN1(n5463), .IN2(n9646), .Q(n7094) );
  INVX0 U7911 ( .INP(n7095), .ZN(WX5900) );
  OR2X1 U7912 ( .IN1(n5463), .IN2(n9649), .Q(n7095) );
  AND2X1 U7913 ( .IN1(test_so46), .IN2(n5405), .Q(WX5898) );
  INVX0 U7914 ( .INP(n7096), .ZN(WX5896) );
  OR2X1 U7915 ( .IN1(n5462), .IN2(n9650), .Q(n7096) );
  INVX0 U7916 ( .INP(n7097), .ZN(WX5894) );
  OR2X1 U7917 ( .IN1(n5462), .IN2(n9651), .Q(n7097) );
  INVX0 U7918 ( .INP(n7098), .ZN(WX5892) );
  OR2X1 U7919 ( .IN1(n5462), .IN2(n9652), .Q(n7098) );
  INVX0 U7920 ( .INP(n7099), .ZN(WX5890) );
  OR2X1 U7921 ( .IN1(n5462), .IN2(n9653), .Q(n7099) );
  INVX0 U7922 ( .INP(n7100), .ZN(WX5888) );
  OR2X1 U7923 ( .IN1(n5462), .IN2(n9654), .Q(n7100) );
  INVX0 U7924 ( .INP(n7101), .ZN(WX5886) );
  OR2X1 U7925 ( .IN1(n5462), .IN2(n9655), .Q(n7101) );
  INVX0 U7926 ( .INP(n7102), .ZN(WX5884) );
  OR2X1 U7927 ( .IN1(n5462), .IN2(n9656), .Q(n7102) );
  INVX0 U7928 ( .INP(n7103), .ZN(WX5882) );
  OR2X1 U7929 ( .IN1(n5462), .IN2(n9657), .Q(n7103) );
  INVX0 U7930 ( .INP(n7104), .ZN(WX5880) );
  OR2X1 U7931 ( .IN1(n5462), .IN2(n9658), .Q(n7104) );
  OR2X1 U7932 ( .IN1(n7105), .IN2(n7106), .Q(WX5878) );
  OR2X1 U7933 ( .IN1(n7107), .IN2(n7108), .Q(n7106) );
  AND2X1 U7934 ( .IN1(test_so53), .IN2(n4888), .Q(n7108) );
  AND2X1 U7935 ( .IN1(n250), .IN2(n4873), .Q(n7107) );
  INVX0 U7936 ( .INP(n7109), .ZN(n250) );
  OR2X1 U7937 ( .IN1(n5462), .IN2(n3910), .Q(n7109) );
  OR2X1 U7938 ( .IN1(n7110), .IN2(n7111), .Q(n7105) );
  AND2X1 U7939 ( .IN1(n4855), .IN2(n7112), .Q(n7111) );
  AND2X1 U7940 ( .IN1(n4937), .IN2(n6471), .Q(n7110) );
  XNOR2X1 U7941 ( .IN1(n7113), .IN2(n7114), .Q(n6471) );
  XOR2X1 U7942 ( .IN1(n9589), .IN2(n4537), .Q(n7114) );
  XOR2X1 U7943 ( .IN1(WX7172), .IN2(n4368), .Q(n7113) );
  OR2X1 U7944 ( .IN1(n7115), .IN2(n7116), .Q(WX5876) );
  OR2X1 U7945 ( .IN1(n7117), .IN2(n7118), .Q(n7116) );
  AND2X1 U7946 ( .IN1(n4907), .IN2(CRC_OUT_5_1), .Q(n7118) );
  AND2X1 U7947 ( .IN1(n249), .IN2(n4873), .Q(n7117) );
  INVX0 U7948 ( .INP(n7119), .ZN(n249) );
  OR2X1 U7949 ( .IN1(n5462), .IN2(n3911), .Q(n7119) );
  OR2X1 U7950 ( .IN1(n7120), .IN2(n7121), .Q(n7115) );
  AND2X1 U7951 ( .IN1(n7122), .IN2(n4833), .Q(n7121) );
  AND2X1 U7952 ( .IN1(n4937), .IN2(n6481), .Q(n7120) );
  XNOR2X1 U7953 ( .IN1(n7123), .IN2(n7124), .Q(n6481) );
  XOR2X1 U7954 ( .IN1(n9590), .IN2(n4646), .Q(n7124) );
  XOR2X1 U7955 ( .IN1(WX7170), .IN2(n4370), .Q(n7123) );
  OR2X1 U7956 ( .IN1(n7125), .IN2(n7126), .Q(WX5874) );
  OR2X1 U7957 ( .IN1(n7127), .IN2(n7128), .Q(n7126) );
  AND2X1 U7958 ( .IN1(n4907), .IN2(CRC_OUT_5_2), .Q(n7128) );
  AND2X1 U7959 ( .IN1(n248), .IN2(n4873), .Q(n7127) );
  INVX0 U7960 ( .INP(n7129), .ZN(n248) );
  OR2X1 U7961 ( .IN1(n5462), .IN2(n3912), .Q(n7129) );
  OR2X1 U7962 ( .IN1(n7130), .IN2(n7131), .Q(n7125) );
  AND2X1 U7963 ( .IN1(n4855), .IN2(n7132), .Q(n7131) );
  AND2X1 U7964 ( .IN1(n4937), .IN2(n6491), .Q(n7130) );
  XNOR2X1 U7965 ( .IN1(n7133), .IN2(n7134), .Q(n6491) );
  XOR2X1 U7966 ( .IN1(n9591), .IN2(n4645), .Q(n7134) );
  XOR2X1 U7967 ( .IN1(WX7168), .IN2(n4372), .Q(n7133) );
  OR2X1 U7968 ( .IN1(n7135), .IN2(n7136), .Q(WX5872) );
  OR2X1 U7969 ( .IN1(n7137), .IN2(n7138), .Q(n7136) );
  AND2X1 U7970 ( .IN1(n4907), .IN2(CRC_OUT_5_3), .Q(n7138) );
  AND2X1 U7971 ( .IN1(n247), .IN2(n4873), .Q(n7137) );
  INVX0 U7972 ( .INP(n7139), .ZN(n247) );
  OR2X1 U7973 ( .IN1(n5462), .IN2(n3913), .Q(n7139) );
  OR2X1 U7974 ( .IN1(n7140), .IN2(n7141), .Q(n7135) );
  AND2X1 U7975 ( .IN1(n7142), .IN2(n4833), .Q(n7141) );
  AND2X1 U7976 ( .IN1(n4937), .IN2(n6501), .Q(n7140) );
  XNOR2X1 U7977 ( .IN1(n7143), .IN2(n7144), .Q(n6501) );
  XOR2X1 U7978 ( .IN1(n9592), .IN2(n4644), .Q(n7144) );
  XOR2X1 U7979 ( .IN1(WX7166), .IN2(n4374), .Q(n7143) );
  OR2X1 U7980 ( .IN1(n7145), .IN2(n7146), .Q(WX5870) );
  OR2X1 U7981 ( .IN1(n7147), .IN2(n7148), .Q(n7146) );
  AND2X1 U7982 ( .IN1(n4908), .IN2(CRC_OUT_5_4), .Q(n7148) );
  AND2X1 U7983 ( .IN1(n246), .IN2(n4873), .Q(n7147) );
  INVX0 U7984 ( .INP(n7149), .ZN(n246) );
  OR2X1 U7985 ( .IN1(n5461), .IN2(n3914), .Q(n7149) );
  OR2X1 U7986 ( .IN1(n7150), .IN2(n7151), .Q(n7145) );
  AND2X1 U7987 ( .IN1(n4855), .IN2(n7152), .Q(n7151) );
  AND2X1 U7988 ( .IN1(n6511), .IN2(n4918), .Q(n7150) );
  XOR2X1 U7989 ( .IN1(n7153), .IN2(n7154), .Q(n6511) );
  XOR2X1 U7990 ( .IN1(test_so64), .IN2(n9593), .Q(n7154) );
  XOR2X1 U7991 ( .IN1(WX7164), .IN2(n4376), .Q(n7153) );
  OR2X1 U7992 ( .IN1(n7155), .IN2(n7156), .Q(WX5868) );
  OR2X1 U7993 ( .IN1(n7157), .IN2(n7158), .Q(n7156) );
  AND2X1 U7994 ( .IN1(n4908), .IN2(CRC_OUT_5_5), .Q(n7158) );
  AND2X1 U7995 ( .IN1(n245), .IN2(n4873), .Q(n7157) );
  INVX0 U7996 ( .INP(n7159), .ZN(n245) );
  OR2X1 U7997 ( .IN1(n5461), .IN2(n3915), .Q(n7159) );
  OR2X1 U7998 ( .IN1(n7160), .IN2(n7161), .Q(n7155) );
  AND2X1 U7999 ( .IN1(n7162), .IN2(n4833), .Q(n7161) );
  AND2X1 U8000 ( .IN1(n4938), .IN2(n6520), .Q(n7160) );
  XNOR2X1 U8001 ( .IN1(n7163), .IN2(n7164), .Q(n6520) );
  XOR2X1 U8002 ( .IN1(n9594), .IN2(n4643), .Q(n7164) );
  XOR2X1 U8003 ( .IN1(WX7162), .IN2(n4378), .Q(n7163) );
  OR2X1 U8004 ( .IN1(n7165), .IN2(n7166), .Q(WX5866) );
  OR2X1 U8005 ( .IN1(n7167), .IN2(n7168), .Q(n7166) );
  AND2X1 U8006 ( .IN1(n4908), .IN2(CRC_OUT_5_6), .Q(n7168) );
  AND2X1 U8007 ( .IN1(n244), .IN2(n4873), .Q(n7167) );
  INVX0 U8008 ( .INP(n7169), .ZN(n244) );
  OR2X1 U8009 ( .IN1(n5461), .IN2(n3916), .Q(n7169) );
  OR2X1 U8010 ( .IN1(n7170), .IN2(n7171), .Q(n7165) );
  AND2X1 U8011 ( .IN1(n4855), .IN2(n7172), .Q(n7171) );
  AND2X1 U8012 ( .IN1(n6530), .IN2(n4918), .Q(n7170) );
  XOR2X1 U8013 ( .IN1(n7173), .IN2(n7174), .Q(n6530) );
  XOR2X1 U8014 ( .IN1(test_so62), .IN2(n9595), .Q(n7174) );
  XOR2X1 U8015 ( .IN1(WX7160), .IN2(n4642), .Q(n7173) );
  OR2X1 U8016 ( .IN1(n7175), .IN2(n7176), .Q(WX5864) );
  OR2X1 U8017 ( .IN1(n7177), .IN2(n7178), .Q(n7176) );
  AND2X1 U8018 ( .IN1(n4908), .IN2(CRC_OUT_5_7), .Q(n7178) );
  AND2X1 U8019 ( .IN1(n243), .IN2(n4873), .Q(n7177) );
  INVX0 U8020 ( .INP(n7179), .ZN(n243) );
  OR2X1 U8021 ( .IN1(n5461), .IN2(n3917), .Q(n7179) );
  OR2X1 U8022 ( .IN1(n7180), .IN2(n7181), .Q(n7175) );
  AND2X1 U8023 ( .IN1(n4855), .IN2(n7182), .Q(n7181) );
  AND2X1 U8024 ( .IN1(n4938), .IN2(n6540), .Q(n7180) );
  XNOR2X1 U8025 ( .IN1(n7183), .IN2(n7184), .Q(n6540) );
  XOR2X1 U8026 ( .IN1(n9596), .IN2(n4641), .Q(n7184) );
  XOR2X1 U8027 ( .IN1(WX7158), .IN2(n4381), .Q(n7183) );
  OR2X1 U8028 ( .IN1(n7185), .IN2(n7186), .Q(WX5862) );
  OR2X1 U8029 ( .IN1(n7187), .IN2(n7188), .Q(n7186) );
  AND2X1 U8030 ( .IN1(n4908), .IN2(CRC_OUT_5_8), .Q(n7188) );
  AND2X1 U8031 ( .IN1(n242), .IN2(n4873), .Q(n7187) );
  INVX0 U8032 ( .INP(n7189), .ZN(n242) );
  OR2X1 U8033 ( .IN1(n5461), .IN2(n3918), .Q(n7189) );
  OR2X1 U8034 ( .IN1(n7190), .IN2(n7191), .Q(n7185) );
  AND2X1 U8035 ( .IN1(n4854), .IN2(n7192), .Q(n7191) );
  AND2X1 U8036 ( .IN1(n6550), .IN2(n4917), .Q(n7190) );
  XOR2X1 U8037 ( .IN1(n7193), .IN2(n7194), .Q(n6550) );
  XOR2X1 U8038 ( .IN1(test_so60), .IN2(n9597), .Q(n7194) );
  XOR2X1 U8039 ( .IN1(WX7156), .IN2(n4640), .Q(n7193) );
  OR2X1 U8040 ( .IN1(n7195), .IN2(n7196), .Q(WX5860) );
  OR2X1 U8041 ( .IN1(n7197), .IN2(n7198), .Q(n7196) );
  AND2X1 U8042 ( .IN1(n4908), .IN2(CRC_OUT_5_9), .Q(n7198) );
  AND2X1 U8043 ( .IN1(n241), .IN2(n4873), .Q(n7197) );
  INVX0 U8044 ( .INP(n7199), .ZN(n241) );
  OR2X1 U8045 ( .IN1(n5461), .IN2(n3919), .Q(n7199) );
  OR2X1 U8046 ( .IN1(n7200), .IN2(n7201), .Q(n7195) );
  AND2X1 U8047 ( .IN1(n4854), .IN2(n7202), .Q(n7201) );
  AND2X1 U8048 ( .IN1(n4938), .IN2(n6560), .Q(n7200) );
  XNOR2X1 U8049 ( .IN1(n7203), .IN2(n7204), .Q(n6560) );
  XOR2X1 U8050 ( .IN1(n9598), .IN2(n4639), .Q(n7204) );
  XOR2X1 U8051 ( .IN1(WX7154), .IN2(n4384), .Q(n7203) );
  OR2X1 U8052 ( .IN1(n7205), .IN2(n7206), .Q(WX5858) );
  OR2X1 U8053 ( .IN1(n7207), .IN2(n7208), .Q(n7206) );
  AND2X1 U8054 ( .IN1(n4908), .IN2(CRC_OUT_5_10), .Q(n7208) );
  AND2X1 U8055 ( .IN1(n240), .IN2(n4873), .Q(n7207) );
  INVX0 U8056 ( .INP(n7209), .ZN(n240) );
  OR2X1 U8057 ( .IN1(n5461), .IN2(n3920), .Q(n7209) );
  OR2X1 U8058 ( .IN1(n7210), .IN2(n7211), .Q(n7205) );
  AND2X1 U8059 ( .IN1(n4854), .IN2(n7212), .Q(n7211) );
  AND2X1 U8060 ( .IN1(n6570), .IN2(n4917), .Q(n7210) );
  XOR2X1 U8061 ( .IN1(n7213), .IN2(n7214), .Q(n6570) );
  XOR2X1 U8062 ( .IN1(test_so58), .IN2(n9599), .Q(n7214) );
  XOR2X1 U8063 ( .IN1(WX7280), .IN2(n4638), .Q(n7213) );
  OR2X1 U8064 ( .IN1(n7215), .IN2(n7216), .Q(WX5856) );
  OR2X1 U8065 ( .IN1(n7217), .IN2(n7218), .Q(n7216) );
  AND2X1 U8066 ( .IN1(n4908), .IN2(CRC_OUT_5_11), .Q(n7218) );
  AND2X1 U8067 ( .IN1(n239), .IN2(n4872), .Q(n7217) );
  INVX0 U8068 ( .INP(n7219), .ZN(n239) );
  OR2X1 U8069 ( .IN1(n5461), .IN2(n3921), .Q(n7219) );
  OR2X1 U8070 ( .IN1(n7220), .IN2(n7221), .Q(n7215) );
  AND2X1 U8071 ( .IN1(n4854), .IN2(n7222), .Q(n7221) );
  AND2X1 U8072 ( .IN1(n4938), .IN2(n6580), .Q(n7220) );
  XNOR2X1 U8073 ( .IN1(n7223), .IN2(n7224), .Q(n6580) );
  XOR2X1 U8074 ( .IN1(n9600), .IN2(n4523), .Q(n7224) );
  XOR2X1 U8075 ( .IN1(WX7150), .IN2(n4387), .Q(n7223) );
  OR2X1 U8076 ( .IN1(n7225), .IN2(n7226), .Q(WX5854) );
  OR2X1 U8077 ( .IN1(n7227), .IN2(n7228), .Q(n7226) );
  AND2X1 U8078 ( .IN1(n4908), .IN2(CRC_OUT_5_12), .Q(n7228) );
  AND2X1 U8079 ( .IN1(n238), .IN2(n4872), .Q(n7227) );
  INVX0 U8080 ( .INP(n7229), .ZN(n238) );
  OR2X1 U8081 ( .IN1(n5461), .IN2(n3922), .Q(n7229) );
  OR2X1 U8082 ( .IN1(n7230), .IN2(n7231), .Q(n7225) );
  AND2X1 U8083 ( .IN1(n4854), .IN2(n7232), .Q(n7231) );
  AND2X1 U8084 ( .IN1(n4938), .IN2(n6590), .Q(n7230) );
  XNOR2X1 U8085 ( .IN1(n7233), .IN2(n7234), .Q(n6590) );
  XOR2X1 U8086 ( .IN1(n9601), .IN2(n4637), .Q(n7234) );
  XOR2X1 U8087 ( .IN1(WX7148), .IN2(n4389), .Q(n7233) );
  OR2X1 U8088 ( .IN1(n7235), .IN2(n7236), .Q(WX5852) );
  OR2X1 U8089 ( .IN1(n7237), .IN2(n7238), .Q(n7236) );
  AND2X1 U8090 ( .IN1(n4908), .IN2(CRC_OUT_5_13), .Q(n7238) );
  AND2X1 U8091 ( .IN1(n237), .IN2(n4872), .Q(n7237) );
  INVX0 U8092 ( .INP(n7239), .ZN(n237) );
  OR2X1 U8093 ( .IN1(n5461), .IN2(n3923), .Q(n7239) );
  OR2X1 U8094 ( .IN1(n7240), .IN2(n7241), .Q(n7235) );
  AND2X1 U8095 ( .IN1(n4854), .IN2(n7242), .Q(n7241) );
  AND2X1 U8096 ( .IN1(n4938), .IN2(n6600), .Q(n7240) );
  XNOR2X1 U8097 ( .IN1(n7243), .IN2(n7244), .Q(n6600) );
  XOR2X1 U8098 ( .IN1(n9602), .IN2(n4636), .Q(n7244) );
  XOR2X1 U8099 ( .IN1(WX7146), .IN2(n4391), .Q(n7243) );
  OR2X1 U8100 ( .IN1(n7245), .IN2(n7246), .Q(WX5850) );
  OR2X1 U8101 ( .IN1(n7247), .IN2(n7248), .Q(n7246) );
  AND2X1 U8102 ( .IN1(n4908), .IN2(CRC_OUT_5_14), .Q(n7248) );
  AND2X1 U8103 ( .IN1(n236), .IN2(n4872), .Q(n7247) );
  INVX0 U8104 ( .INP(n7249), .ZN(n236) );
  OR2X1 U8105 ( .IN1(n5461), .IN2(n3924), .Q(n7249) );
  OR2X1 U8106 ( .IN1(n7250), .IN2(n7251), .Q(n7245) );
  AND2X1 U8107 ( .IN1(n4854), .IN2(n7252), .Q(n7251) );
  AND2X1 U8108 ( .IN1(n4938), .IN2(n6610), .Q(n7250) );
  XNOR2X1 U8109 ( .IN1(n7253), .IN2(n7254), .Q(n6610) );
  XOR2X1 U8110 ( .IN1(n9603), .IN2(n4635), .Q(n7254) );
  XOR2X1 U8111 ( .IN1(WX7144), .IN2(n4393), .Q(n7253) );
  OR2X1 U8112 ( .IN1(n7255), .IN2(n7256), .Q(WX5848) );
  OR2X1 U8113 ( .IN1(n7257), .IN2(n7258), .Q(n7256) );
  AND2X1 U8114 ( .IN1(n4908), .IN2(CRC_OUT_5_15), .Q(n7258) );
  AND2X1 U8115 ( .IN1(n235), .IN2(n4872), .Q(n7257) );
  INVX0 U8116 ( .INP(n7259), .ZN(n235) );
  OR2X1 U8117 ( .IN1(n5467), .IN2(n3925), .Q(n7259) );
  OR2X1 U8118 ( .IN1(n7260), .IN2(n7261), .Q(n7255) );
  AND2X1 U8119 ( .IN1(n4854), .IN2(n7262), .Q(n7261) );
  AND2X1 U8120 ( .IN1(n4938), .IN2(n6620), .Q(n7260) );
  XNOR2X1 U8121 ( .IN1(n7263), .IN2(n7264), .Q(n6620) );
  XOR2X1 U8122 ( .IN1(n9604), .IN2(n4634), .Q(n7264) );
  XOR2X1 U8123 ( .IN1(WX7142), .IN2(n4395), .Q(n7263) );
  OR2X1 U8124 ( .IN1(n7265), .IN2(n7266), .Q(WX5846) );
  OR2X1 U8125 ( .IN1(n7267), .IN2(n7268), .Q(n7266) );
  AND2X1 U8126 ( .IN1(n4908), .IN2(CRC_OUT_5_16), .Q(n7268) );
  AND2X1 U8127 ( .IN1(n234), .IN2(n4872), .Q(n7267) );
  INVX0 U8128 ( .INP(n7269), .ZN(n234) );
  OR2X1 U8129 ( .IN1(n5480), .IN2(n3926), .Q(n7269) );
  OR2X1 U8130 ( .IN1(n7270), .IN2(n7271), .Q(n7265) );
  AND2X1 U8131 ( .IN1(n7272), .IN2(n4835), .Q(n7271) );
  AND2X1 U8132 ( .IN1(n4938), .IN2(n6630), .Q(n7270) );
  XNOR2X1 U8133 ( .IN1(n7273), .IN2(n7274), .Q(n6630) );
  XOR2X1 U8134 ( .IN1(n4212), .IN2(n5387), .Q(n7274) );
  XOR2X1 U8135 ( .IN1(n7275), .IN2(n4522), .Q(n7273) );
  XOR2X1 U8136 ( .IN1(WX7268), .IN2(n9605), .Q(n7275) );
  OR2X1 U8137 ( .IN1(n7276), .IN2(n7277), .Q(WX5844) );
  OR2X1 U8138 ( .IN1(n7278), .IN2(n7279), .Q(n7277) );
  AND2X1 U8139 ( .IN1(test_so54), .IN2(n4887), .Q(n7279) );
  AND2X1 U8140 ( .IN1(n233), .IN2(n4872), .Q(n7278) );
  INVX0 U8141 ( .INP(n7280), .ZN(n233) );
  OR2X1 U8142 ( .IN1(n5480), .IN2(n3927), .Q(n7280) );
  OR2X1 U8143 ( .IN1(n7281), .IN2(n7282), .Q(n7276) );
  AND2X1 U8144 ( .IN1(n4854), .IN2(n7283), .Q(n7282) );
  AND2X1 U8145 ( .IN1(n4938), .IN2(n6641), .Q(n7281) );
  XNOR2X1 U8146 ( .IN1(n7284), .IN2(n7285), .Q(n6641) );
  XOR2X1 U8147 ( .IN1(n4213), .IN2(n5387), .Q(n7285) );
  XOR2X1 U8148 ( .IN1(n7286), .IN2(n4633), .Q(n7284) );
  XOR2X1 U8149 ( .IN1(WX7266), .IN2(n9606), .Q(n7286) );
  OR2X1 U8150 ( .IN1(n7287), .IN2(n7288), .Q(WX5842) );
  OR2X1 U8151 ( .IN1(n7289), .IN2(n7290), .Q(n7288) );
  AND2X1 U8152 ( .IN1(n4909), .IN2(CRC_OUT_5_18), .Q(n7290) );
  AND2X1 U8153 ( .IN1(n232), .IN2(n4872), .Q(n7289) );
  INVX0 U8154 ( .INP(n7291), .ZN(n232) );
  OR2X1 U8155 ( .IN1(n5480), .IN2(n3928), .Q(n7291) );
  OR2X1 U8156 ( .IN1(n7292), .IN2(n7293), .Q(n7287) );
  AND2X1 U8157 ( .IN1(n7294), .IN2(n4835), .Q(n7293) );
  AND2X1 U8158 ( .IN1(n4938), .IN2(n6652), .Q(n7292) );
  XNOR2X1 U8159 ( .IN1(n7295), .IN2(n7296), .Q(n6652) );
  XOR2X1 U8160 ( .IN1(n4214), .IN2(n5387), .Q(n7296) );
  XOR2X1 U8161 ( .IN1(n7297), .IN2(n4632), .Q(n7295) );
  XOR2X1 U8162 ( .IN1(WX7264), .IN2(n9607), .Q(n7297) );
  OR2X1 U8163 ( .IN1(n7298), .IN2(n7299), .Q(WX5840) );
  OR2X1 U8164 ( .IN1(n7300), .IN2(n7301), .Q(n7299) );
  AND2X1 U8165 ( .IN1(n4909), .IN2(CRC_OUT_5_19), .Q(n7301) );
  AND2X1 U8166 ( .IN1(n231), .IN2(n4872), .Q(n7300) );
  INVX0 U8167 ( .INP(n7302), .ZN(n231) );
  OR2X1 U8168 ( .IN1(n5480), .IN2(n3929), .Q(n7302) );
  OR2X1 U8169 ( .IN1(n7303), .IN2(n7304), .Q(n7298) );
  AND2X1 U8170 ( .IN1(n4854), .IN2(n7305), .Q(n7304) );
  AND2X1 U8171 ( .IN1(n4938), .IN2(n6663), .Q(n7303) );
  XNOR2X1 U8172 ( .IN1(n7306), .IN2(n7307), .Q(n6663) );
  XOR2X1 U8173 ( .IN1(n4215), .IN2(n5387), .Q(n7307) );
  XOR2X1 U8174 ( .IN1(n7308), .IN2(n4631), .Q(n7306) );
  XOR2X1 U8175 ( .IN1(WX7262), .IN2(n9608), .Q(n7308) );
  OR2X1 U8176 ( .IN1(n7309), .IN2(n7310), .Q(WX5838) );
  OR2X1 U8177 ( .IN1(n7311), .IN2(n7312), .Q(n7310) );
  AND2X1 U8178 ( .IN1(n4909), .IN2(CRC_OUT_5_20), .Q(n7312) );
  AND2X1 U8179 ( .IN1(n230), .IN2(n4872), .Q(n7311) );
  INVX0 U8180 ( .INP(n7313), .ZN(n230) );
  OR2X1 U8181 ( .IN1(n5480), .IN2(n3930), .Q(n7313) );
  OR2X1 U8182 ( .IN1(n7314), .IN2(n7315), .Q(n7309) );
  AND2X1 U8183 ( .IN1(n7316), .IN2(n4835), .Q(n7315) );
  AND2X1 U8184 ( .IN1(n4938), .IN2(n6674), .Q(n7314) );
  XNOR2X1 U8185 ( .IN1(n7317), .IN2(n7318), .Q(n6674) );
  XOR2X1 U8186 ( .IN1(n4216), .IN2(n5387), .Q(n7318) );
  XOR2X1 U8187 ( .IN1(n7319), .IN2(n4630), .Q(n7317) );
  XOR2X1 U8188 ( .IN1(WX7260), .IN2(n9609), .Q(n7319) );
  OR2X1 U8189 ( .IN1(n7320), .IN2(n7321), .Q(WX5836) );
  OR2X1 U8190 ( .IN1(n7322), .IN2(n7323), .Q(n7321) );
  AND2X1 U8191 ( .IN1(n4893), .IN2(CRC_OUT_5_21), .Q(n7323) );
  AND2X1 U8192 ( .IN1(n229), .IN2(n4872), .Q(n7322) );
  INVX0 U8193 ( .INP(n7324), .ZN(n229) );
  OR2X1 U8194 ( .IN1(n5480), .IN2(n3931), .Q(n7324) );
  OR2X1 U8195 ( .IN1(n7325), .IN2(n7326), .Q(n7320) );
  AND2X1 U8196 ( .IN1(n4854), .IN2(n7327), .Q(n7326) );
  AND2X1 U8197 ( .IN1(n6685), .IN2(n4917), .Q(n7325) );
  XOR2X1 U8198 ( .IN1(n7328), .IN2(n7329), .Q(n6685) );
  XOR2X1 U8199 ( .IN1(n4217), .IN2(n5386), .Q(n7329) );
  XOR2X1 U8200 ( .IN1(WX7194), .IN2(n7330), .Q(n7328) );
  XOR2X1 U8201 ( .IN1(test_so63), .IN2(n9610), .Q(n7330) );
  OR2X1 U8202 ( .IN1(n7331), .IN2(n7332), .Q(WX5834) );
  OR2X1 U8203 ( .IN1(n7333), .IN2(n7334), .Q(n7332) );
  AND2X1 U8204 ( .IN1(n4888), .IN2(CRC_OUT_5_22), .Q(n7334) );
  AND2X1 U8205 ( .IN1(n228), .IN2(n4872), .Q(n7333) );
  INVX0 U8206 ( .INP(n7335), .ZN(n228) );
  OR2X1 U8207 ( .IN1(n5480), .IN2(n3932), .Q(n7335) );
  OR2X1 U8208 ( .IN1(n7336), .IN2(n7337), .Q(n7331) );
  AND2X1 U8209 ( .IN1(n7338), .IN2(n4835), .Q(n7337) );
  AND2X1 U8210 ( .IN1(n4939), .IN2(n6696), .Q(n7336) );
  XNOR2X1 U8211 ( .IN1(n7339), .IN2(n7340), .Q(n6696) );
  XOR2X1 U8212 ( .IN1(n4218), .IN2(n5386), .Q(n7340) );
  XOR2X1 U8213 ( .IN1(n7341), .IN2(n4629), .Q(n7339) );
  XOR2X1 U8214 ( .IN1(WX7256), .IN2(n9611), .Q(n7341) );
  OR2X1 U8215 ( .IN1(n7342), .IN2(n7343), .Q(WX5832) );
  OR2X1 U8216 ( .IN1(n7344), .IN2(n7345), .Q(n7343) );
  AND2X1 U8217 ( .IN1(n4890), .IN2(CRC_OUT_5_23), .Q(n7345) );
  AND2X1 U8218 ( .IN1(n227), .IN2(n4871), .Q(n7344) );
  INVX0 U8219 ( .INP(n7346), .ZN(n227) );
  OR2X1 U8220 ( .IN1(n5481), .IN2(n3933), .Q(n7346) );
  OR2X1 U8221 ( .IN1(n7347), .IN2(n7348), .Q(n7342) );
  AND2X1 U8222 ( .IN1(n4854), .IN2(n7349), .Q(n7348) );
  AND2X1 U8223 ( .IN1(n6707), .IN2(n4917), .Q(n7347) );
  XOR2X1 U8224 ( .IN1(n7350), .IN2(n7351), .Q(n6707) );
  XOR2X1 U8225 ( .IN1(n4628), .IN2(n5386), .Q(n7351) );
  XOR2X1 U8226 ( .IN1(n7352), .IN2(n9614), .Q(n7350) );
  XOR2X1 U8227 ( .IN1(n9613), .IN2(n9612), .Q(n7352) );
  OR2X1 U8228 ( .IN1(n7353), .IN2(n7354), .Q(WX5830) );
  OR2X1 U8229 ( .IN1(n7355), .IN2(n7356), .Q(n7354) );
  AND2X1 U8230 ( .IN1(n4888), .IN2(CRC_OUT_5_24), .Q(n7356) );
  AND2X1 U8231 ( .IN1(n226), .IN2(n4871), .Q(n7355) );
  INVX0 U8232 ( .INP(n7357), .ZN(n226) );
  OR2X1 U8233 ( .IN1(n5481), .IN2(n3934), .Q(n7357) );
  OR2X1 U8234 ( .IN1(n7358), .IN2(n7359), .Q(n7353) );
  AND2X1 U8235 ( .IN1(n4854), .IN2(n7360), .Q(n7359) );
  AND2X1 U8236 ( .IN1(n4939), .IN2(n6718), .Q(n7358) );
  XNOR2X1 U8237 ( .IN1(n7361), .IN2(n7362), .Q(n6718) );
  XOR2X1 U8238 ( .IN1(n4219), .IN2(n5386), .Q(n7362) );
  XOR2X1 U8239 ( .IN1(n7363), .IN2(n4627), .Q(n7361) );
  XOR2X1 U8240 ( .IN1(WX7252), .IN2(n9615), .Q(n7363) );
  OR2X1 U8241 ( .IN1(n7364), .IN2(n7365), .Q(WX5828) );
  OR2X1 U8242 ( .IN1(n7366), .IN2(n7367), .Q(n7365) );
  AND2X1 U8243 ( .IN1(n4889), .IN2(CRC_OUT_5_25), .Q(n7367) );
  AND2X1 U8244 ( .IN1(n225), .IN2(n4871), .Q(n7366) );
  INVX0 U8245 ( .INP(n7368), .ZN(n225) );
  OR2X1 U8246 ( .IN1(n5481), .IN2(n3935), .Q(n7368) );
  OR2X1 U8247 ( .IN1(n7369), .IN2(n7370), .Q(n7364) );
  AND2X1 U8248 ( .IN1(n4853), .IN2(n7371), .Q(n7370) );
  AND2X1 U8249 ( .IN1(n6729), .IN2(n4917), .Q(n7369) );
  XOR2X1 U8250 ( .IN1(n7372), .IN2(n7373), .Q(n6729) );
  XOR2X1 U8251 ( .IN1(n4626), .IN2(n5386), .Q(n7373) );
  XOR2X1 U8252 ( .IN1(n7374), .IN2(n9618), .Q(n7372) );
  XOR2X1 U8253 ( .IN1(n9617), .IN2(n9616), .Q(n7374) );
  OR2X1 U8254 ( .IN1(n7375), .IN2(n7376), .Q(WX5826) );
  OR2X1 U8255 ( .IN1(n7377), .IN2(n7378), .Q(n7376) );
  AND2X1 U8256 ( .IN1(n4888), .IN2(CRC_OUT_5_26), .Q(n7378) );
  AND2X1 U8257 ( .IN1(n224), .IN2(n4871), .Q(n7377) );
  INVX0 U8258 ( .INP(n7379), .ZN(n224) );
  OR2X1 U8259 ( .IN1(n5481), .IN2(n3936), .Q(n7379) );
  OR2X1 U8260 ( .IN1(n7380), .IN2(n7381), .Q(n7375) );
  AND2X1 U8261 ( .IN1(n4853), .IN2(n7382), .Q(n7381) );
  AND2X1 U8262 ( .IN1(n4939), .IN2(n6740), .Q(n7380) );
  XNOR2X1 U8263 ( .IN1(n7383), .IN2(n7384), .Q(n6740) );
  XOR2X1 U8264 ( .IN1(n4220), .IN2(n5386), .Q(n7384) );
  XOR2X1 U8265 ( .IN1(n7385), .IN2(n4625), .Q(n7383) );
  XOR2X1 U8266 ( .IN1(WX7248), .IN2(n9619), .Q(n7385) );
  OR2X1 U8267 ( .IN1(n7386), .IN2(n7387), .Q(WX5824) );
  OR2X1 U8268 ( .IN1(n7388), .IN2(n7389), .Q(n7387) );
  AND2X1 U8269 ( .IN1(n4889), .IN2(CRC_OUT_5_27), .Q(n7389) );
  AND2X1 U8270 ( .IN1(n223), .IN2(n4871), .Q(n7388) );
  INVX0 U8271 ( .INP(n7390), .ZN(n223) );
  OR2X1 U8272 ( .IN1(n5481), .IN2(n3937), .Q(n7390) );
  OR2X1 U8273 ( .IN1(n7391), .IN2(n7392), .Q(n7386) );
  AND2X1 U8274 ( .IN1(n4853), .IN2(n7393), .Q(n7392) );
  AND2X1 U8275 ( .IN1(n6751), .IN2(n4917), .Q(n7391) );
  XOR2X1 U8276 ( .IN1(n7394), .IN2(n7395), .Q(n6751) );
  XOR2X1 U8277 ( .IN1(n4221), .IN2(n5386), .Q(n7395) );
  XOR2X1 U8278 ( .IN1(n7396), .IN2(n4624), .Q(n7394) );
  XOR2X1 U8279 ( .IN1(WX7182), .IN2(test_so57), .Q(n7396) );
  OR2X1 U8280 ( .IN1(n7397), .IN2(n7398), .Q(WX5822) );
  OR2X1 U8281 ( .IN1(n7399), .IN2(n7400), .Q(n7398) );
  AND2X1 U8282 ( .IN1(n4888), .IN2(CRC_OUT_5_28), .Q(n7400) );
  AND2X1 U8283 ( .IN1(n222), .IN2(n4871), .Q(n7399) );
  INVX0 U8284 ( .INP(n7401), .ZN(n222) );
  OR2X1 U8285 ( .IN1(n5481), .IN2(n3938), .Q(n7401) );
  OR2X1 U8286 ( .IN1(n7402), .IN2(n7403), .Q(n7397) );
  AND2X1 U8287 ( .IN1(n4853), .IN2(n7404), .Q(n7403) );
  AND2X1 U8288 ( .IN1(n4939), .IN2(n6762), .Q(n7402) );
  XNOR2X1 U8289 ( .IN1(n7405), .IN2(n7406), .Q(n6762) );
  XOR2X1 U8290 ( .IN1(n4222), .IN2(n5386), .Q(n7406) );
  XOR2X1 U8291 ( .IN1(n7407), .IN2(n4623), .Q(n7405) );
  XOR2X1 U8292 ( .IN1(WX7244), .IN2(n9620), .Q(n7407) );
  OR2X1 U8293 ( .IN1(n7408), .IN2(n7409), .Q(WX5820) );
  OR2X1 U8294 ( .IN1(n7410), .IN2(n7411), .Q(n7409) );
  AND2X1 U8295 ( .IN1(n4889), .IN2(CRC_OUT_5_29), .Q(n7411) );
  AND2X1 U8296 ( .IN1(n221), .IN2(n4871), .Q(n7410) );
  INVX0 U8297 ( .INP(n7412), .ZN(n221) );
  OR2X1 U8298 ( .IN1(n5481), .IN2(n3939), .Q(n7412) );
  OR2X1 U8299 ( .IN1(n7413), .IN2(n7414), .Q(n7408) );
  AND2X1 U8300 ( .IN1(n4853), .IN2(n7415), .Q(n7414) );
  AND2X1 U8301 ( .IN1(n4939), .IN2(n6773), .Q(n7413) );
  XNOR2X1 U8302 ( .IN1(n7416), .IN2(n7417), .Q(n6773) );
  XOR2X1 U8303 ( .IN1(n4223), .IN2(n5386), .Q(n7417) );
  XOR2X1 U8304 ( .IN1(n7418), .IN2(n4622), .Q(n7416) );
  XOR2X1 U8305 ( .IN1(WX7242), .IN2(n9621), .Q(n7418) );
  OR2X1 U8306 ( .IN1(n7419), .IN2(n7420), .Q(WX5818) );
  OR2X1 U8307 ( .IN1(n7421), .IN2(n7422), .Q(n7420) );
  AND2X1 U8308 ( .IN1(n4888), .IN2(CRC_OUT_5_30), .Q(n7422) );
  AND2X1 U8309 ( .IN1(n220), .IN2(n4871), .Q(n7421) );
  INVX0 U8310 ( .INP(n7423), .ZN(n220) );
  OR2X1 U8311 ( .IN1(n5481), .IN2(n3940), .Q(n7423) );
  OR2X1 U8312 ( .IN1(n7424), .IN2(n7425), .Q(n7419) );
  AND2X1 U8313 ( .IN1(n4853), .IN2(n7426), .Q(n7425) );
  AND2X1 U8314 ( .IN1(n4939), .IN2(n6784), .Q(n7424) );
  XNOR2X1 U8315 ( .IN1(n7427), .IN2(n7428), .Q(n6784) );
  XOR2X1 U8316 ( .IN1(n4224), .IN2(n5386), .Q(n7428) );
  XOR2X1 U8317 ( .IN1(n7429), .IN2(n4621), .Q(n7427) );
  XOR2X1 U8318 ( .IN1(WX7240), .IN2(n9622), .Q(n7429) );
  OR2X1 U8319 ( .IN1(n7430), .IN2(n7431), .Q(WX5816) );
  OR2X1 U8320 ( .IN1(n7432), .IN2(n7433), .Q(n7431) );
  AND2X1 U8321 ( .IN1(n2245), .IN2(WX5657), .Q(n7433) );
  AND2X1 U8322 ( .IN1(n4890), .IN2(CRC_OUT_5_31), .Q(n7432) );
  OR2X1 U8323 ( .IN1(n7434), .IN2(n7435), .Q(n7430) );
  AND2X1 U8324 ( .IN1(n4853), .IN2(n7436), .Q(n7435) );
  AND2X1 U8325 ( .IN1(n4939), .IN2(n6794), .Q(n7434) );
  XNOR2X1 U8326 ( .IN1(n7437), .IN2(n7438), .Q(n6794) );
  XOR2X1 U8327 ( .IN1(n4168), .IN2(n5386), .Q(n7438) );
  XOR2X1 U8328 ( .IN1(n7439), .IN2(n4620), .Q(n7437) );
  XOR2X1 U8329 ( .IN1(WX7238), .IN2(n9623), .Q(n7439) );
  AND2X1 U8330 ( .IN1(n4822), .IN2(n5405), .Q(WX5718) );
  AND2X1 U8331 ( .IN1(n4827), .IN2(n5405), .Q(WX546) );
  AND2X1 U8332 ( .IN1(n7440), .IN2(n5405), .Q(WX5205) );
  XOR2X1 U8333 ( .IN1(CRC_OUT_6_30), .IN2(n4675), .Q(n7440) );
  AND2X1 U8334 ( .IN1(n7441), .IN2(n5405), .Q(WX5203) );
  XOR2X1 U8335 ( .IN1(CRC_OUT_6_29), .IN2(n4676), .Q(n7441) );
  AND2X1 U8336 ( .IN1(n7442), .IN2(n5405), .Q(WX5201) );
  XOR2X1 U8337 ( .IN1(CRC_OUT_6_28), .IN2(n4677), .Q(n7442) );
  AND2X1 U8338 ( .IN1(n7443), .IN2(n5406), .Q(WX5199) );
  XOR2X1 U8339 ( .IN1(test_so40), .IN2(DFF_763_n1), .Q(n7443) );
  AND2X1 U8340 ( .IN1(n7444), .IN2(n5406), .Q(WX5197) );
  XOR2X1 U8341 ( .IN1(CRC_OUT_6_26), .IN2(n4678), .Q(n7444) );
  AND2X1 U8342 ( .IN1(n7445), .IN2(n5406), .Q(WX5195) );
  XOR2X1 U8343 ( .IN1(CRC_OUT_6_25), .IN2(n4679), .Q(n7445) );
  AND2X1 U8344 ( .IN1(n7446), .IN2(n5406), .Q(WX5193) );
  XOR2X1 U8345 ( .IN1(CRC_OUT_6_24), .IN2(n4680), .Q(n7446) );
  AND2X1 U8346 ( .IN1(n7447), .IN2(n5406), .Q(WX5191) );
  XOR2X1 U8347 ( .IN1(CRC_OUT_6_23), .IN2(n4681), .Q(n7447) );
  AND2X1 U8348 ( .IN1(n7448), .IN2(n5406), .Q(WX5189) );
  XOR2X1 U8349 ( .IN1(test_so43), .IN2(n4682), .Q(n7448) );
  AND2X1 U8350 ( .IN1(n7449), .IN2(n5406), .Q(WX5187) );
  XOR2X1 U8351 ( .IN1(CRC_OUT_6_21), .IN2(n4683), .Q(n7449) );
  AND2X1 U8352 ( .IN1(n7450), .IN2(n5406), .Q(WX5185) );
  XOR2X1 U8353 ( .IN1(CRC_OUT_6_20), .IN2(n4684), .Q(n7450) );
  AND2X1 U8354 ( .IN1(n7451), .IN2(n5406), .Q(WX5183) );
  XOR2X1 U8355 ( .IN1(CRC_OUT_6_19), .IN2(n4685), .Q(n7451) );
  AND2X1 U8356 ( .IN1(n7452), .IN2(n5407), .Q(WX5181) );
  XOR2X1 U8357 ( .IN1(CRC_OUT_6_18), .IN2(n4686), .Q(n7452) );
  AND2X1 U8358 ( .IN1(n7453), .IN2(n5407), .Q(WX5179) );
  XOR2X1 U8359 ( .IN1(CRC_OUT_6_17), .IN2(n4687), .Q(n7453) );
  AND2X1 U8360 ( .IN1(n7454), .IN2(n5407), .Q(WX5177) );
  XOR2X1 U8361 ( .IN1(CRC_OUT_6_16), .IN2(n4688), .Q(n7454) );
  AND2X1 U8362 ( .IN1(n7455), .IN2(n5407), .Q(WX5175) );
  XOR2X1 U8363 ( .IN1(DFF_751_n1), .IN2(n7456), .Q(n7455) );
  XOR2X1 U8364 ( .IN1(n4526), .IN2(DFF_767_n1), .Q(n7456) );
  AND2X1 U8365 ( .IN1(n7457), .IN2(n5407), .Q(WX5173) );
  XOR2X1 U8366 ( .IN1(CRC_OUT_6_14), .IN2(n4689), .Q(n7457) );
  AND2X1 U8367 ( .IN1(n7458), .IN2(n5407), .Q(WX5171) );
  XOR2X1 U8368 ( .IN1(CRC_OUT_6_13), .IN2(n4690), .Q(n7458) );
  AND2X1 U8369 ( .IN1(n7459), .IN2(n5407), .Q(WX5169) );
  XOR2X1 U8370 ( .IN1(CRC_OUT_6_12), .IN2(n4691), .Q(n7459) );
  AND2X1 U8371 ( .IN1(n7460), .IN2(n5407), .Q(WX5167) );
  XOR2X1 U8372 ( .IN1(CRC_OUT_6_11), .IN2(n4692), .Q(n7460) );
  AND2X1 U8373 ( .IN1(n7461), .IN2(n5407), .Q(WX5165) );
  XOR2X1 U8374 ( .IN1(CRC_OUT_6_10), .IN2(n7462), .Q(n7461) );
  XOR2X1 U8375 ( .IN1(test_so41), .IN2(DFF_767_n1), .Q(n7462) );
  AND2X1 U8376 ( .IN1(n7463), .IN2(n5408), .Q(WX5163) );
  XOR2X1 U8377 ( .IN1(CRC_OUT_6_9), .IN2(n4693), .Q(n7463) );
  AND2X1 U8378 ( .IN1(n7464), .IN2(n5408), .Q(WX5161) );
  XOR2X1 U8379 ( .IN1(CRC_OUT_6_8), .IN2(n4694), .Q(n7464) );
  AND2X1 U8380 ( .IN1(n7465), .IN2(n5431), .Q(WX5159) );
  XOR2X1 U8381 ( .IN1(CRC_OUT_6_7), .IN2(n4695), .Q(n7465) );
  AND2X1 U8382 ( .IN1(n7466), .IN2(n5425), .Q(WX5157) );
  XOR2X1 U8383 ( .IN1(CRC_OUT_6_6), .IN2(n4696), .Q(n7466) );
  AND2X1 U8384 ( .IN1(n7467), .IN2(n5426), .Q(WX5155) );
  XOR2X1 U8385 ( .IN1(test_so42), .IN2(n4697), .Q(n7467) );
  AND2X1 U8386 ( .IN1(n7468), .IN2(n5426), .Q(WX5153) );
  XOR2X1 U8387 ( .IN1(CRC_OUT_6_4), .IN2(n4698), .Q(n7468) );
  AND2X1 U8388 ( .IN1(n7469), .IN2(n5426), .Q(WX5151) );
  XOR2X1 U8389 ( .IN1(DFF_739_n1), .IN2(n7470), .Q(n7469) );
  XOR2X1 U8390 ( .IN1(n4527), .IN2(DFF_767_n1), .Q(n7470) );
  AND2X1 U8391 ( .IN1(n7471), .IN2(n5426), .Q(WX5149) );
  XOR2X1 U8392 ( .IN1(CRC_OUT_6_2), .IN2(n4699), .Q(n7471) );
  AND2X1 U8393 ( .IN1(n7472), .IN2(n5426), .Q(WX5147) );
  XOR2X1 U8394 ( .IN1(CRC_OUT_6_1), .IN2(n4700), .Q(n7472) );
  AND2X1 U8395 ( .IN1(n7473), .IN2(n5426), .Q(WX5145) );
  XOR2X1 U8396 ( .IN1(CRC_OUT_6_0), .IN2(n4701), .Q(n7473) );
  AND2X1 U8397 ( .IN1(n7474), .IN2(n5426), .Q(WX5143) );
  XOR2X1 U8398 ( .IN1(n4539), .IN2(CRC_OUT_6_31), .Q(n7474) );
  INVX0 U8399 ( .INP(n7475), .ZN(WX4617) );
  OR2X1 U8400 ( .IN1(n5481), .IN2(n9675), .Q(n7475) );
  AND2X1 U8401 ( .IN1(test_so35), .IN2(n5426), .Q(WX4615) );
  INVX0 U8402 ( .INP(n7476), .ZN(WX4613) );
  OR2X1 U8403 ( .IN1(n5481), .IN2(n9676), .Q(n7476) );
  INVX0 U8404 ( .INP(n7477), .ZN(WX4611) );
  OR2X1 U8405 ( .IN1(n5481), .IN2(n9677), .Q(n7477) );
  INVX0 U8406 ( .INP(n7478), .ZN(WX4609) );
  OR2X1 U8407 ( .IN1(n5481), .IN2(n9678), .Q(n7478) );
  INVX0 U8408 ( .INP(n7479), .ZN(WX4607) );
  OR2X1 U8409 ( .IN1(n5481), .IN2(n9679), .Q(n7479) );
  INVX0 U8410 ( .INP(n7480), .ZN(WX4605) );
  OR2X1 U8411 ( .IN1(n5482), .IN2(n9680), .Q(n7480) );
  INVX0 U8412 ( .INP(n7481), .ZN(WX4603) );
  OR2X1 U8413 ( .IN1(n5482), .IN2(n9681), .Q(n7481) );
  INVX0 U8414 ( .INP(n7482), .ZN(WX4601) );
  OR2X1 U8415 ( .IN1(n5482), .IN2(n9682), .Q(n7482) );
  INVX0 U8416 ( .INP(n7483), .ZN(WX4599) );
  OR2X1 U8417 ( .IN1(n5482), .IN2(n9683), .Q(n7483) );
  INVX0 U8418 ( .INP(n7484), .ZN(WX4597) );
  OR2X1 U8419 ( .IN1(n5482), .IN2(n9684), .Q(n7484) );
  INVX0 U8420 ( .INP(n7485), .ZN(WX4595) );
  OR2X1 U8421 ( .IN1(n5482), .IN2(n9685), .Q(n7485) );
  INVX0 U8422 ( .INP(n7486), .ZN(WX4593) );
  OR2X1 U8423 ( .IN1(n5482), .IN2(n9686), .Q(n7486) );
  INVX0 U8424 ( .INP(n7487), .ZN(WX4591) );
  OR2X1 U8425 ( .IN1(n5482), .IN2(n9687), .Q(n7487) );
  INVX0 U8426 ( .INP(n7488), .ZN(WX4589) );
  OR2X1 U8427 ( .IN1(n5482), .IN2(n9688), .Q(n7488) );
  INVX0 U8428 ( .INP(n7489), .ZN(WX4587) );
  OR2X1 U8429 ( .IN1(n5482), .IN2(n9691), .Q(n7489) );
  OR2X1 U8430 ( .IN1(n7490), .IN2(n7491), .Q(WX4585) );
  OR2X1 U8431 ( .IN1(n7492), .IN2(n7493), .Q(n7491) );
  AND2X1 U8432 ( .IN1(n4888), .IN2(CRC_OUT_6_0), .Q(n7493) );
  AND2X1 U8433 ( .IN1(n188), .IN2(n4871), .Q(n7492) );
  INVX0 U8434 ( .INP(n7494), .ZN(n188) );
  OR2X1 U8435 ( .IN1(n5482), .IN2(n3941), .Q(n7494) );
  OR2X1 U8436 ( .IN1(n7495), .IN2(n7496), .Q(n7490) );
  AND2X1 U8437 ( .IN1(n7497), .IN2(n4836), .Q(n7496) );
  AND2X1 U8438 ( .IN1(n4939), .IN2(n7112), .Q(n7495) );
  XNOR2X1 U8439 ( .IN1(n7498), .IN2(n7499), .Q(n7112) );
  XOR2X1 U8440 ( .IN1(n9624), .IN2(n4538), .Q(n7499) );
  XOR2X1 U8441 ( .IN1(WX5879), .IN2(n4397), .Q(n7498) );
  OR2X1 U8442 ( .IN1(n7500), .IN2(n7501), .Q(WX4583) );
  OR2X1 U8443 ( .IN1(n7502), .IN2(n7503), .Q(n7501) );
  AND2X1 U8444 ( .IN1(n4889), .IN2(CRC_OUT_6_1), .Q(n7503) );
  AND2X1 U8445 ( .IN1(n187), .IN2(n4871), .Q(n7502) );
  INVX0 U8446 ( .INP(n7504), .ZN(n187) );
  OR2X1 U8447 ( .IN1(n5482), .IN2(n3942), .Q(n7504) );
  OR2X1 U8448 ( .IN1(n7505), .IN2(n7506), .Q(n7500) );
  AND2X1 U8449 ( .IN1(n4853), .IN2(n7507), .Q(n7506) );
  AND2X1 U8450 ( .IN1(n7122), .IN2(n4917), .Q(n7505) );
  XOR2X1 U8451 ( .IN1(n7508), .IN2(n7509), .Q(n7122) );
  XOR2X1 U8452 ( .IN1(test_so51), .IN2(n9625), .Q(n7509) );
  XOR2X1 U8453 ( .IN1(WX5877), .IN2(n4674), .Q(n7508) );
  OR2X1 U8454 ( .IN1(n7510), .IN2(n7511), .Q(WX4581) );
  OR2X1 U8455 ( .IN1(n7512), .IN2(n7513), .Q(n7511) );
  AND2X1 U8456 ( .IN1(n4888), .IN2(CRC_OUT_6_2), .Q(n7513) );
  AND2X1 U8457 ( .IN1(n186), .IN2(n4871), .Q(n7512) );
  INVX0 U8458 ( .INP(n7514), .ZN(n186) );
  OR2X1 U8459 ( .IN1(n5482), .IN2(n3943), .Q(n7514) );
  OR2X1 U8460 ( .IN1(n7515), .IN2(n7516), .Q(n7510) );
  AND2X1 U8461 ( .IN1(n4853), .IN2(n7517), .Q(n7516) );
  AND2X1 U8462 ( .IN1(n4939), .IN2(n7132), .Q(n7515) );
  XNOR2X1 U8463 ( .IN1(n7518), .IN2(n7519), .Q(n7132) );
  XOR2X1 U8464 ( .IN1(n9626), .IN2(n4673), .Q(n7519) );
  XOR2X1 U8465 ( .IN1(WX5875), .IN2(n4400), .Q(n7518) );
  OR2X1 U8466 ( .IN1(n7520), .IN2(n7521), .Q(WX4579) );
  OR2X1 U8467 ( .IN1(n7522), .IN2(n7523), .Q(n7521) );
  AND2X1 U8468 ( .IN1(n4889), .IN2(CRC_OUT_6_3), .Q(n7523) );
  AND2X1 U8469 ( .IN1(n185), .IN2(n4871), .Q(n7522) );
  INVX0 U8470 ( .INP(n7524), .ZN(n185) );
  OR2X1 U8471 ( .IN1(n5483), .IN2(n3944), .Q(n7524) );
  OR2X1 U8472 ( .IN1(n7525), .IN2(n7526), .Q(n7520) );
  AND2X1 U8473 ( .IN1(n4853), .IN2(n7527), .Q(n7526) );
  AND2X1 U8474 ( .IN1(n7142), .IN2(n4917), .Q(n7525) );
  XOR2X1 U8475 ( .IN1(n7528), .IN2(n7529), .Q(n7142) );
  XOR2X1 U8476 ( .IN1(test_so49), .IN2(n9627), .Q(n7529) );
  XOR2X1 U8477 ( .IN1(WX5873), .IN2(n4672), .Q(n7528) );
  OR2X1 U8478 ( .IN1(n7530), .IN2(n7531), .Q(WX4577) );
  OR2X1 U8479 ( .IN1(n7532), .IN2(n7533), .Q(n7531) );
  AND2X1 U8480 ( .IN1(n4889), .IN2(CRC_OUT_6_4), .Q(n7533) );
  AND2X1 U8481 ( .IN1(n184), .IN2(n4870), .Q(n7532) );
  INVX0 U8482 ( .INP(n7534), .ZN(n184) );
  OR2X1 U8483 ( .IN1(n5483), .IN2(n3945), .Q(n7534) );
  OR2X1 U8484 ( .IN1(n7535), .IN2(n7536), .Q(n7530) );
  AND2X1 U8485 ( .IN1(n4853), .IN2(n7537), .Q(n7536) );
  AND2X1 U8486 ( .IN1(n4924), .IN2(n7152), .Q(n7535) );
  XNOR2X1 U8487 ( .IN1(n7538), .IN2(n7539), .Q(n7152) );
  XOR2X1 U8488 ( .IN1(n9628), .IN2(n4525), .Q(n7539) );
  XOR2X1 U8489 ( .IN1(WX5871), .IN2(n4403), .Q(n7538) );
  OR2X1 U8490 ( .IN1(n7540), .IN2(n7541), .Q(WX4575) );
  OR2X1 U8491 ( .IN1(n7542), .IN2(n7543), .Q(n7541) );
  AND2X1 U8492 ( .IN1(test_so42), .IN2(n4887), .Q(n7543) );
  AND2X1 U8493 ( .IN1(n183), .IN2(n4870), .Q(n7542) );
  INVX0 U8494 ( .INP(n7544), .ZN(n183) );
  OR2X1 U8495 ( .IN1(n5483), .IN2(n3946), .Q(n7544) );
  OR2X1 U8496 ( .IN1(n7545), .IN2(n7546), .Q(n7540) );
  AND2X1 U8497 ( .IN1(n4853), .IN2(n7547), .Q(n7546) );
  AND2X1 U8498 ( .IN1(n7162), .IN2(n4917), .Q(n7545) );
  XOR2X1 U8499 ( .IN1(n7548), .IN2(n7549), .Q(n7162) );
  XOR2X1 U8500 ( .IN1(test_so47), .IN2(n9629), .Q(n7549) );
  XOR2X1 U8501 ( .IN1(WX5997), .IN2(n4671), .Q(n7548) );
  OR2X1 U8502 ( .IN1(n7550), .IN2(n7551), .Q(WX4573) );
  OR2X1 U8503 ( .IN1(n7552), .IN2(n7553), .Q(n7551) );
  AND2X1 U8504 ( .IN1(n4889), .IN2(CRC_OUT_6_6), .Q(n7553) );
  AND2X1 U8505 ( .IN1(n182), .IN2(n4870), .Q(n7552) );
  INVX0 U8506 ( .INP(n7554), .ZN(n182) );
  OR2X1 U8507 ( .IN1(n5483), .IN2(n3947), .Q(n7554) );
  OR2X1 U8508 ( .IN1(n7555), .IN2(n7556), .Q(n7550) );
  AND2X1 U8509 ( .IN1(n4853), .IN2(n7557), .Q(n7556) );
  AND2X1 U8510 ( .IN1(n4926), .IN2(n7172), .Q(n7555) );
  XNOR2X1 U8511 ( .IN1(n7558), .IN2(n7559), .Q(n7172) );
  XOR2X1 U8512 ( .IN1(n9630), .IN2(n4670), .Q(n7559) );
  XOR2X1 U8513 ( .IN1(WX5867), .IN2(n4406), .Q(n7558) );
  OR2X1 U8514 ( .IN1(n7560), .IN2(n7561), .Q(WX4571) );
  OR2X1 U8515 ( .IN1(n7562), .IN2(n7563), .Q(n7561) );
  AND2X1 U8516 ( .IN1(n4889), .IN2(CRC_OUT_6_7), .Q(n7563) );
  AND2X1 U8517 ( .IN1(n181), .IN2(n4870), .Q(n7562) );
  INVX0 U8518 ( .INP(n7564), .ZN(n181) );
  OR2X1 U8519 ( .IN1(n5483), .IN2(n3948), .Q(n7564) );
  OR2X1 U8520 ( .IN1(n7565), .IN2(n7566), .Q(n7560) );
  AND2X1 U8521 ( .IN1(n4852), .IN2(n7567), .Q(n7566) );
  AND2X1 U8522 ( .IN1(n4924), .IN2(n7182), .Q(n7565) );
  XNOR2X1 U8523 ( .IN1(n7568), .IN2(n7569), .Q(n7182) );
  XOR2X1 U8524 ( .IN1(n9631), .IN2(n4669), .Q(n7569) );
  XOR2X1 U8525 ( .IN1(WX5865), .IN2(n4408), .Q(n7568) );
  OR2X1 U8526 ( .IN1(n7570), .IN2(n7571), .Q(WX4569) );
  OR2X1 U8527 ( .IN1(n7572), .IN2(n7573), .Q(n7571) );
  AND2X1 U8528 ( .IN1(n4891), .IN2(CRC_OUT_6_8), .Q(n7573) );
  AND2X1 U8529 ( .IN1(n180), .IN2(n4870), .Q(n7572) );
  INVX0 U8530 ( .INP(n7574), .ZN(n180) );
  OR2X1 U8531 ( .IN1(n5483), .IN2(n3949), .Q(n7574) );
  OR2X1 U8532 ( .IN1(n7575), .IN2(n7576), .Q(n7570) );
  AND2X1 U8533 ( .IN1(n4852), .IN2(n7577), .Q(n7576) );
  AND2X1 U8534 ( .IN1(n4924), .IN2(n7192), .Q(n7575) );
  XNOR2X1 U8535 ( .IN1(n7578), .IN2(n7579), .Q(n7192) );
  XOR2X1 U8536 ( .IN1(n9632), .IN2(n4668), .Q(n7579) );
  XOR2X1 U8537 ( .IN1(WX5863), .IN2(n4410), .Q(n7578) );
  OR2X1 U8538 ( .IN1(n7580), .IN2(n7581), .Q(WX4567) );
  OR2X1 U8539 ( .IN1(n7582), .IN2(n7583), .Q(n7581) );
  AND2X1 U8540 ( .IN1(n4889), .IN2(CRC_OUT_6_9), .Q(n7583) );
  AND2X1 U8541 ( .IN1(n179), .IN2(n4870), .Q(n7582) );
  INVX0 U8542 ( .INP(n7584), .ZN(n179) );
  OR2X1 U8543 ( .IN1(n5483), .IN2(n3950), .Q(n7584) );
  OR2X1 U8544 ( .IN1(n7585), .IN2(n7586), .Q(n7580) );
  AND2X1 U8545 ( .IN1(n4852), .IN2(n7587), .Q(n7586) );
  AND2X1 U8546 ( .IN1(n4925), .IN2(n7202), .Q(n7585) );
  XNOR2X1 U8547 ( .IN1(n7588), .IN2(n7589), .Q(n7202) );
  XOR2X1 U8548 ( .IN1(n9633), .IN2(n4667), .Q(n7589) );
  XOR2X1 U8549 ( .IN1(WX5861), .IN2(n4412), .Q(n7588) );
  OR2X1 U8550 ( .IN1(n7590), .IN2(n7591), .Q(WX4565) );
  OR2X1 U8551 ( .IN1(n7592), .IN2(n7593), .Q(n7591) );
  AND2X1 U8552 ( .IN1(n4890), .IN2(CRC_OUT_6_10), .Q(n7593) );
  AND2X1 U8553 ( .IN1(n178), .IN2(n4870), .Q(n7592) );
  INVX0 U8554 ( .INP(n7594), .ZN(n178) );
  OR2X1 U8555 ( .IN1(n5483), .IN2(n3951), .Q(n7594) );
  OR2X1 U8556 ( .IN1(n7595), .IN2(n7596), .Q(n7590) );
  AND2X1 U8557 ( .IN1(n4852), .IN2(n7597), .Q(n7596) );
  AND2X1 U8558 ( .IN1(n4925), .IN2(n7212), .Q(n7595) );
  XNOR2X1 U8559 ( .IN1(n7598), .IN2(n7599), .Q(n7212) );
  XOR2X1 U8560 ( .IN1(n9634), .IN2(n4666), .Q(n7599) );
  XOR2X1 U8561 ( .IN1(WX5859), .IN2(n4414), .Q(n7598) );
  OR2X1 U8562 ( .IN1(n7600), .IN2(n7601), .Q(WX4563) );
  OR2X1 U8563 ( .IN1(n7602), .IN2(n7603), .Q(n7601) );
  AND2X1 U8564 ( .IN1(n4889), .IN2(CRC_OUT_6_11), .Q(n7603) );
  AND2X1 U8565 ( .IN1(n177), .IN2(n4870), .Q(n7602) );
  INVX0 U8566 ( .INP(n7604), .ZN(n177) );
  OR2X1 U8567 ( .IN1(n5483), .IN2(n3952), .Q(n7604) );
  OR2X1 U8568 ( .IN1(n7605), .IN2(n7606), .Q(n7600) );
  AND2X1 U8569 ( .IN1(n7607), .IN2(n4838), .Q(n7606) );
  AND2X1 U8570 ( .IN1(n4924), .IN2(n7222), .Q(n7605) );
  XNOR2X1 U8571 ( .IN1(n7608), .IN2(n7609), .Q(n7222) );
  XOR2X1 U8572 ( .IN1(n9635), .IN2(n4524), .Q(n7609) );
  XOR2X1 U8573 ( .IN1(WX5857), .IN2(n4416), .Q(n7608) );
  OR2X1 U8574 ( .IN1(n7610), .IN2(n7611), .Q(WX4561) );
  OR2X1 U8575 ( .IN1(n7612), .IN2(n7613), .Q(n7611) );
  AND2X1 U8576 ( .IN1(n4890), .IN2(CRC_OUT_6_12), .Q(n7613) );
  AND2X1 U8577 ( .IN1(n176), .IN2(n4870), .Q(n7612) );
  INVX0 U8578 ( .INP(n7614), .ZN(n176) );
  OR2X1 U8579 ( .IN1(n5483), .IN2(n3953), .Q(n7614) );
  OR2X1 U8580 ( .IN1(n7615), .IN2(n7616), .Q(n7610) );
  AND2X1 U8581 ( .IN1(n4852), .IN2(n7617), .Q(n7616) );
  AND2X1 U8582 ( .IN1(n4925), .IN2(n7232), .Q(n7615) );
  XNOR2X1 U8583 ( .IN1(n7618), .IN2(n7619), .Q(n7232) );
  XOR2X1 U8584 ( .IN1(n9636), .IN2(n4665), .Q(n7619) );
  XOR2X1 U8585 ( .IN1(WX5855), .IN2(n4418), .Q(n7618) );
  OR2X1 U8586 ( .IN1(n7620), .IN2(n7621), .Q(WX4559) );
  OR2X1 U8587 ( .IN1(n7622), .IN2(n7623), .Q(n7621) );
  AND2X1 U8588 ( .IN1(n4889), .IN2(CRC_OUT_6_13), .Q(n7623) );
  AND2X1 U8589 ( .IN1(n175), .IN2(n4870), .Q(n7622) );
  INVX0 U8590 ( .INP(n7624), .ZN(n175) );
  OR2X1 U8591 ( .IN1(n5483), .IN2(n3954), .Q(n7624) );
  OR2X1 U8592 ( .IN1(n7625), .IN2(n7626), .Q(n7620) );
  AND2X1 U8593 ( .IN1(n7627), .IN2(n4838), .Q(n7626) );
  AND2X1 U8594 ( .IN1(n4925), .IN2(n7242), .Q(n7625) );
  XNOR2X1 U8595 ( .IN1(n7628), .IN2(n7629), .Q(n7242) );
  XOR2X1 U8596 ( .IN1(n9637), .IN2(n4664), .Q(n7629) );
  XOR2X1 U8597 ( .IN1(WX5853), .IN2(n4420), .Q(n7628) );
  OR2X1 U8598 ( .IN1(n7630), .IN2(n7631), .Q(WX4557) );
  OR2X1 U8599 ( .IN1(n7632), .IN2(n7633), .Q(n7631) );
  AND2X1 U8600 ( .IN1(n4891), .IN2(CRC_OUT_6_14), .Q(n7633) );
  AND2X1 U8601 ( .IN1(n174), .IN2(n4870), .Q(n7632) );
  INVX0 U8602 ( .INP(n7634), .ZN(n174) );
  OR2X1 U8603 ( .IN1(n5483), .IN2(n3955), .Q(n7634) );
  OR2X1 U8604 ( .IN1(n7635), .IN2(n7636), .Q(n7630) );
  AND2X1 U8605 ( .IN1(n4852), .IN2(n7637), .Q(n7636) );
  AND2X1 U8606 ( .IN1(n4924), .IN2(n7252), .Q(n7635) );
  XNOR2X1 U8607 ( .IN1(n7638), .IN2(n7639), .Q(n7252) );
  XOR2X1 U8608 ( .IN1(n9638), .IN2(n4663), .Q(n7639) );
  XOR2X1 U8609 ( .IN1(WX5851), .IN2(n4422), .Q(n7638) );
  OR2X1 U8610 ( .IN1(n7640), .IN2(n7641), .Q(WX4555) );
  OR2X1 U8611 ( .IN1(n7642), .IN2(n7643), .Q(n7641) );
  AND2X1 U8612 ( .IN1(n4889), .IN2(CRC_OUT_6_15), .Q(n7643) );
  AND2X1 U8613 ( .IN1(n173), .IN2(n4870), .Q(n7642) );
  INVX0 U8614 ( .INP(n7644), .ZN(n173) );
  OR2X1 U8615 ( .IN1(n5484), .IN2(n3956), .Q(n7644) );
  OR2X1 U8616 ( .IN1(n7645), .IN2(n7646), .Q(n7640) );
  AND2X1 U8617 ( .IN1(n7647), .IN2(n4836), .Q(n7646) );
  AND2X1 U8618 ( .IN1(n4925), .IN2(n7262), .Q(n7645) );
  XNOR2X1 U8619 ( .IN1(n7648), .IN2(n7649), .Q(n7262) );
  XOR2X1 U8620 ( .IN1(n9639), .IN2(n4662), .Q(n7649) );
  XOR2X1 U8621 ( .IN1(WX5849), .IN2(n4424), .Q(n7648) );
  OR2X1 U8622 ( .IN1(n7650), .IN2(n7651), .Q(WX4553) );
  OR2X1 U8623 ( .IN1(n7652), .IN2(n7653), .Q(n7651) );
  AND2X1 U8624 ( .IN1(n4890), .IN2(CRC_OUT_6_16), .Q(n7653) );
  AND2X1 U8625 ( .IN1(n172), .IN2(n4869), .Q(n7652) );
  INVX0 U8626 ( .INP(n7654), .ZN(n172) );
  OR2X1 U8627 ( .IN1(n5484), .IN2(n3957), .Q(n7654) );
  OR2X1 U8628 ( .IN1(n7655), .IN2(n7656), .Q(n7650) );
  AND2X1 U8629 ( .IN1(n4852), .IN2(n7657), .Q(n7656) );
  AND2X1 U8630 ( .IN1(n7272), .IN2(n4917), .Q(n7655) );
  XOR2X1 U8631 ( .IN1(n7658), .IN2(n7659), .Q(n7272) );
  XOR2X1 U8632 ( .IN1(n4225), .IN2(n5386), .Q(n7659) );
  XOR2X1 U8633 ( .IN1(WX5911), .IN2(n7660), .Q(n7658) );
  XOR2X1 U8634 ( .IN1(test_so52), .IN2(n9640), .Q(n7660) );
  OR2X1 U8635 ( .IN1(n7661), .IN2(n7662), .Q(WX4551) );
  OR2X1 U8636 ( .IN1(n7663), .IN2(n7664), .Q(n7662) );
  AND2X1 U8637 ( .IN1(n4890), .IN2(CRC_OUT_6_17), .Q(n7664) );
  AND2X1 U8638 ( .IN1(n171), .IN2(n4869), .Q(n7663) );
  INVX0 U8639 ( .INP(n7665), .ZN(n171) );
  OR2X1 U8640 ( .IN1(n5484), .IN2(n3958), .Q(n7665) );
  OR2X1 U8641 ( .IN1(n7666), .IN2(n7667), .Q(n7661) );
  AND2X1 U8642 ( .IN1(n7668), .IN2(n4836), .Q(n7667) );
  AND2X1 U8643 ( .IN1(n4924), .IN2(n7283), .Q(n7666) );
  XNOR2X1 U8644 ( .IN1(n7669), .IN2(n7670), .Q(n7283) );
  XOR2X1 U8645 ( .IN1(n4226), .IN2(n5385), .Q(n7670) );
  XOR2X1 U8646 ( .IN1(n7671), .IN2(n4661), .Q(n7669) );
  XOR2X1 U8647 ( .IN1(WX5973), .IN2(n9641), .Q(n7671) );
  OR2X1 U8648 ( .IN1(n7672), .IN2(n7673), .Q(WX4549) );
  OR2X1 U8649 ( .IN1(n7674), .IN2(n7675), .Q(n7673) );
  AND2X1 U8650 ( .IN1(n4890), .IN2(CRC_OUT_6_18), .Q(n7675) );
  AND2X1 U8651 ( .IN1(n170), .IN2(n4869), .Q(n7674) );
  INVX0 U8652 ( .INP(n7676), .ZN(n170) );
  OR2X1 U8653 ( .IN1(n5484), .IN2(n3959), .Q(n7676) );
  OR2X1 U8654 ( .IN1(n7677), .IN2(n7678), .Q(n7672) );
  AND2X1 U8655 ( .IN1(n4852), .IN2(n7679), .Q(n7678) );
  AND2X1 U8656 ( .IN1(n7294), .IN2(n4920), .Q(n7677) );
  XOR2X1 U8657 ( .IN1(n7680), .IN2(n7681), .Q(n7294) );
  XOR2X1 U8658 ( .IN1(n4660), .IN2(n5385), .Q(n7681) );
  XOR2X1 U8659 ( .IN1(n7682), .IN2(n9644), .Q(n7680) );
  XOR2X1 U8660 ( .IN1(n9643), .IN2(n9642), .Q(n7682) );
  OR2X1 U8661 ( .IN1(n7683), .IN2(n7684), .Q(WX4547) );
  OR2X1 U8662 ( .IN1(n7685), .IN2(n7686), .Q(n7684) );
  AND2X1 U8663 ( .IN1(n4890), .IN2(CRC_OUT_6_19), .Q(n7686) );
  AND2X1 U8664 ( .IN1(n169), .IN2(n4869), .Q(n7685) );
  INVX0 U8665 ( .INP(n7687), .ZN(n169) );
  OR2X1 U8666 ( .IN1(n5484), .IN2(n3960), .Q(n7687) );
  OR2X1 U8667 ( .IN1(n7688), .IN2(n7689), .Q(n7683) );
  AND2X1 U8668 ( .IN1(n4852), .IN2(n7690), .Q(n7689) );
  AND2X1 U8669 ( .IN1(n4924), .IN2(n7305), .Q(n7688) );
  XNOR2X1 U8670 ( .IN1(n7691), .IN2(n7692), .Q(n7305) );
  XOR2X1 U8671 ( .IN1(n4227), .IN2(n5385), .Q(n7692) );
  XOR2X1 U8672 ( .IN1(n7693), .IN2(n4659), .Q(n7691) );
  XOR2X1 U8673 ( .IN1(WX5969), .IN2(n9645), .Q(n7693) );
  OR2X1 U8674 ( .IN1(n7694), .IN2(n7695), .Q(WX4545) );
  OR2X1 U8675 ( .IN1(n7696), .IN2(n7697), .Q(n7695) );
  AND2X1 U8676 ( .IN1(n4890), .IN2(CRC_OUT_6_20), .Q(n7697) );
  AND2X1 U8677 ( .IN1(n168), .IN2(n4869), .Q(n7696) );
  INVX0 U8678 ( .INP(n7698), .ZN(n168) );
  OR2X1 U8679 ( .IN1(n5484), .IN2(n3961), .Q(n7698) );
  OR2X1 U8680 ( .IN1(n7699), .IN2(n7700), .Q(n7694) );
  AND2X1 U8681 ( .IN1(n4852), .IN2(n7701), .Q(n7700) );
  AND2X1 U8682 ( .IN1(n7316), .IN2(n4917), .Q(n7699) );
  XOR2X1 U8683 ( .IN1(n7702), .IN2(n7703), .Q(n7316) );
  XOR2X1 U8684 ( .IN1(n4658), .IN2(n5385), .Q(n7703) );
  XOR2X1 U8685 ( .IN1(n7704), .IN2(n9648), .Q(n7702) );
  XOR2X1 U8686 ( .IN1(n9647), .IN2(n9646), .Q(n7704) );
  OR2X1 U8687 ( .IN1(n7705), .IN2(n7706), .Q(WX4543) );
  OR2X1 U8688 ( .IN1(n7707), .IN2(n7708), .Q(n7706) );
  AND2X1 U8689 ( .IN1(n4890), .IN2(CRC_OUT_6_21), .Q(n7708) );
  AND2X1 U8690 ( .IN1(n167), .IN2(n4869), .Q(n7707) );
  INVX0 U8691 ( .INP(n7709), .ZN(n167) );
  OR2X1 U8692 ( .IN1(n5484), .IN2(n3962), .Q(n7709) );
  OR2X1 U8693 ( .IN1(n7710), .IN2(n7711), .Q(n7705) );
  AND2X1 U8694 ( .IN1(n4852), .IN2(n7712), .Q(n7711) );
  AND2X1 U8695 ( .IN1(n4925), .IN2(n7327), .Q(n7710) );
  XNOR2X1 U8696 ( .IN1(n7713), .IN2(n7714), .Q(n7327) );
  XOR2X1 U8697 ( .IN1(n4228), .IN2(n5385), .Q(n7714) );
  XOR2X1 U8698 ( .IN1(n7715), .IN2(n4657), .Q(n7713) );
  XOR2X1 U8699 ( .IN1(WX5965), .IN2(n9649), .Q(n7715) );
  OR2X1 U8700 ( .IN1(n7716), .IN2(n7717), .Q(WX4541) );
  OR2X1 U8701 ( .IN1(n7718), .IN2(n7719), .Q(n7717) );
  AND2X1 U8702 ( .IN1(test_so43), .IN2(n4887), .Q(n7719) );
  AND2X1 U8703 ( .IN1(n166), .IN2(n4869), .Q(n7718) );
  INVX0 U8704 ( .INP(n7720), .ZN(n166) );
  OR2X1 U8705 ( .IN1(n5484), .IN2(n3963), .Q(n7720) );
  OR2X1 U8706 ( .IN1(n7721), .IN2(n7722), .Q(n7716) );
  AND2X1 U8707 ( .IN1(n4852), .IN2(n7723), .Q(n7722) );
  AND2X1 U8708 ( .IN1(n7338), .IN2(n4917), .Q(n7721) );
  XOR2X1 U8709 ( .IN1(n7724), .IN2(n7725), .Q(n7338) );
  XOR2X1 U8710 ( .IN1(n4229), .IN2(n5385), .Q(n7725) );
  XOR2X1 U8711 ( .IN1(n7726), .IN2(n4656), .Q(n7724) );
  XOR2X1 U8712 ( .IN1(WX5899), .IN2(test_so46), .Q(n7726) );
  OR2X1 U8713 ( .IN1(n7727), .IN2(n7728), .Q(WX4539) );
  OR2X1 U8714 ( .IN1(n7729), .IN2(n7730), .Q(n7728) );
  AND2X1 U8715 ( .IN1(n4891), .IN2(CRC_OUT_6_23), .Q(n7730) );
  AND2X1 U8716 ( .IN1(n165), .IN2(n4869), .Q(n7729) );
  INVX0 U8717 ( .INP(n7731), .ZN(n165) );
  OR2X1 U8718 ( .IN1(n5484), .IN2(n3964), .Q(n7731) );
  OR2X1 U8719 ( .IN1(n7732), .IN2(n7733), .Q(n7727) );
  AND2X1 U8720 ( .IN1(n4852), .IN2(n7734), .Q(n7733) );
  AND2X1 U8721 ( .IN1(n4925), .IN2(n7349), .Q(n7732) );
  XNOR2X1 U8722 ( .IN1(n7735), .IN2(n7736), .Q(n7349) );
  XOR2X1 U8723 ( .IN1(n4230), .IN2(n5385), .Q(n7736) );
  XOR2X1 U8724 ( .IN1(n7737), .IN2(n4655), .Q(n7735) );
  XOR2X1 U8725 ( .IN1(WX5961), .IN2(n9650), .Q(n7737) );
  OR2X1 U8726 ( .IN1(n7738), .IN2(n7739), .Q(WX4537) );
  OR2X1 U8727 ( .IN1(n7740), .IN2(n7741), .Q(n7739) );
  AND2X1 U8728 ( .IN1(n4890), .IN2(CRC_OUT_6_24), .Q(n7741) );
  AND2X1 U8729 ( .IN1(n164), .IN2(n4869), .Q(n7740) );
  INVX0 U8730 ( .INP(n7742), .ZN(n164) );
  OR2X1 U8731 ( .IN1(n5484), .IN2(n3965), .Q(n7742) );
  OR2X1 U8732 ( .IN1(n7743), .IN2(n7744), .Q(n7738) );
  AND2X1 U8733 ( .IN1(n4851), .IN2(n7745), .Q(n7744) );
  AND2X1 U8734 ( .IN1(n4925), .IN2(n7360), .Q(n7743) );
  XNOR2X1 U8735 ( .IN1(n7746), .IN2(n7747), .Q(n7360) );
  XOR2X1 U8736 ( .IN1(n4231), .IN2(n5385), .Q(n7747) );
  XOR2X1 U8737 ( .IN1(n7748), .IN2(n4654), .Q(n7746) );
  XOR2X1 U8738 ( .IN1(WX5959), .IN2(n9651), .Q(n7748) );
  OR2X1 U8739 ( .IN1(n7749), .IN2(n7750), .Q(WX4535) );
  OR2X1 U8740 ( .IN1(n7751), .IN2(n7752), .Q(n7750) );
  AND2X1 U8741 ( .IN1(n4891), .IN2(CRC_OUT_6_25), .Q(n7752) );
  AND2X1 U8742 ( .IN1(n163), .IN2(n4869), .Q(n7751) );
  INVX0 U8743 ( .INP(n7753), .ZN(n163) );
  OR2X1 U8744 ( .IN1(n5484), .IN2(n3966), .Q(n7753) );
  OR2X1 U8745 ( .IN1(n7754), .IN2(n7755), .Q(n7749) );
  AND2X1 U8746 ( .IN1(n4851), .IN2(n7756), .Q(n7755) );
  AND2X1 U8747 ( .IN1(n4925), .IN2(n7371), .Q(n7754) );
  XNOR2X1 U8748 ( .IN1(n7757), .IN2(n7758), .Q(n7371) );
  XOR2X1 U8749 ( .IN1(n4232), .IN2(n5385), .Q(n7758) );
  XOR2X1 U8750 ( .IN1(n7759), .IN2(n4653), .Q(n7757) );
  XOR2X1 U8751 ( .IN1(WX5957), .IN2(n9652), .Q(n7759) );
  OR2X1 U8752 ( .IN1(n7760), .IN2(n7761), .Q(WX4533) );
  OR2X1 U8753 ( .IN1(n7762), .IN2(n7763), .Q(n7761) );
  AND2X1 U8754 ( .IN1(n4890), .IN2(CRC_OUT_6_26), .Q(n7763) );
  AND2X1 U8755 ( .IN1(n162), .IN2(n4869), .Q(n7762) );
  INVX0 U8756 ( .INP(n7764), .ZN(n162) );
  OR2X1 U8757 ( .IN1(n5484), .IN2(n3967), .Q(n7764) );
  OR2X1 U8758 ( .IN1(n7765), .IN2(n7766), .Q(n7760) );
  AND2X1 U8759 ( .IN1(n4851), .IN2(n7767), .Q(n7766) );
  AND2X1 U8760 ( .IN1(n4925), .IN2(n7382), .Q(n7765) );
  XNOR2X1 U8761 ( .IN1(n7768), .IN2(n7769), .Q(n7382) );
  XOR2X1 U8762 ( .IN1(n4233), .IN2(n5385), .Q(n7769) );
  XOR2X1 U8763 ( .IN1(n7770), .IN2(n4652), .Q(n7768) );
  XOR2X1 U8764 ( .IN1(WX5955), .IN2(n9653), .Q(n7770) );
  OR2X1 U8765 ( .IN1(n7771), .IN2(n7772), .Q(WX4531) );
  OR2X1 U8766 ( .IN1(n7773), .IN2(n7774), .Q(n7772) );
  AND2X1 U8767 ( .IN1(n4891), .IN2(CRC_OUT_6_27), .Q(n7774) );
  AND2X1 U8768 ( .IN1(n161), .IN2(n4869), .Q(n7773) );
  INVX0 U8769 ( .INP(n7775), .ZN(n161) );
  OR2X1 U8770 ( .IN1(n5484), .IN2(n3968), .Q(n7775) );
  OR2X1 U8771 ( .IN1(n7776), .IN2(n7777), .Q(n7771) );
  AND2X1 U8772 ( .IN1(n4851), .IN2(n7778), .Q(n7777) );
  AND2X1 U8773 ( .IN1(n4925), .IN2(n7393), .Q(n7776) );
  XNOR2X1 U8774 ( .IN1(n7779), .IN2(n7780), .Q(n7393) );
  XOR2X1 U8775 ( .IN1(n4234), .IN2(n5385), .Q(n7780) );
  XOR2X1 U8776 ( .IN1(n7781), .IN2(n4651), .Q(n7779) );
  XOR2X1 U8777 ( .IN1(WX5953), .IN2(n9654), .Q(n7781) );
  OR2X1 U8778 ( .IN1(n7782), .IN2(n7783), .Q(WX4529) );
  OR2X1 U8779 ( .IN1(n7784), .IN2(n7785), .Q(n7783) );
  AND2X1 U8780 ( .IN1(n4890), .IN2(CRC_OUT_6_28), .Q(n7785) );
  AND2X1 U8781 ( .IN1(n160), .IN2(n4868), .Q(n7784) );
  INVX0 U8782 ( .INP(n7786), .ZN(n160) );
  OR2X1 U8783 ( .IN1(n5485), .IN2(n3969), .Q(n7786) );
  OR2X1 U8784 ( .IN1(n7787), .IN2(n7788), .Q(n7782) );
  AND2X1 U8785 ( .IN1(n7789), .IN2(n4833), .Q(n7788) );
  AND2X1 U8786 ( .IN1(n4926), .IN2(n7404), .Q(n7787) );
  XNOR2X1 U8787 ( .IN1(n7790), .IN2(n7791), .Q(n7404) );
  XOR2X1 U8788 ( .IN1(n4235), .IN2(n5385), .Q(n7791) );
  XOR2X1 U8789 ( .IN1(n7792), .IN2(n4650), .Q(n7790) );
  XOR2X1 U8790 ( .IN1(WX5951), .IN2(n9655), .Q(n7792) );
  OR2X1 U8791 ( .IN1(n7793), .IN2(n7794), .Q(WX4527) );
  OR2X1 U8792 ( .IN1(n7795), .IN2(n7796), .Q(n7794) );
  AND2X1 U8793 ( .IN1(n4892), .IN2(CRC_OUT_6_29), .Q(n7796) );
  AND2X1 U8794 ( .IN1(n159), .IN2(n4868), .Q(n7795) );
  INVX0 U8795 ( .INP(n7797), .ZN(n159) );
  OR2X1 U8796 ( .IN1(n5485), .IN2(n3970), .Q(n7797) );
  OR2X1 U8797 ( .IN1(n7798), .IN2(n7799), .Q(n7793) );
  AND2X1 U8798 ( .IN1(n4851), .IN2(n7800), .Q(n7799) );
  AND2X1 U8799 ( .IN1(n4925), .IN2(n7415), .Q(n7798) );
  XNOR2X1 U8800 ( .IN1(n7801), .IN2(n7802), .Q(n7415) );
  XOR2X1 U8801 ( .IN1(n4236), .IN2(n5384), .Q(n7802) );
  XOR2X1 U8802 ( .IN1(n7803), .IN2(n4649), .Q(n7801) );
  XOR2X1 U8803 ( .IN1(WX5949), .IN2(n9656), .Q(n7803) );
  OR2X1 U8804 ( .IN1(n7804), .IN2(n7805), .Q(WX4525) );
  OR2X1 U8805 ( .IN1(n7806), .IN2(n7807), .Q(n7805) );
  AND2X1 U8806 ( .IN1(n4891), .IN2(CRC_OUT_6_30), .Q(n7807) );
  AND2X1 U8807 ( .IN1(n158), .IN2(n4868), .Q(n7806) );
  INVX0 U8808 ( .INP(n7808), .ZN(n158) );
  OR2X1 U8809 ( .IN1(n5485), .IN2(n3971), .Q(n7808) );
  OR2X1 U8810 ( .IN1(n7809), .IN2(n7810), .Q(n7804) );
  AND2X1 U8811 ( .IN1(n7811), .IN2(n4833), .Q(n7810) );
  AND2X1 U8812 ( .IN1(n4926), .IN2(n7426), .Q(n7809) );
  XNOR2X1 U8813 ( .IN1(n7812), .IN2(n7813), .Q(n7426) );
  XOR2X1 U8814 ( .IN1(n4237), .IN2(n5384), .Q(n7813) );
  XOR2X1 U8815 ( .IN1(n7814), .IN2(n4648), .Q(n7812) );
  XOR2X1 U8816 ( .IN1(WX5947), .IN2(n9657), .Q(n7814) );
  OR2X1 U8817 ( .IN1(n7815), .IN2(n7816), .Q(WX4523) );
  OR2X1 U8818 ( .IN1(n7817), .IN2(n7818), .Q(n7816) );
  AND2X1 U8819 ( .IN1(n2245), .IN2(WX4364), .Q(n7818) );
  AND2X1 U8820 ( .IN1(n4891), .IN2(CRC_OUT_6_31), .Q(n7817) );
  OR2X1 U8821 ( .IN1(n7819), .IN2(n7820), .Q(n7815) );
  AND2X1 U8822 ( .IN1(n4851), .IN2(n7821), .Q(n7820) );
  AND2X1 U8823 ( .IN1(n4926), .IN2(n7436), .Q(n7819) );
  XNOR2X1 U8824 ( .IN1(n7822), .IN2(n7823), .Q(n7436) );
  XOR2X1 U8825 ( .IN1(n4169), .IN2(n5384), .Q(n7823) );
  XOR2X1 U8826 ( .IN1(n7824), .IN2(n4647), .Q(n7822) );
  XOR2X1 U8827 ( .IN1(WX5945), .IN2(n9658), .Q(n7824) );
  AND2X1 U8828 ( .IN1(n4821), .IN2(n5426), .Q(WX4425) );
  AND2X1 U8829 ( .IN1(n7825), .IN2(n5427), .Q(WX3912) );
  XOR2X1 U8830 ( .IN1(CRC_OUT_7_30), .IN2(n4702), .Q(n7825) );
  AND2X1 U8831 ( .IN1(n7826), .IN2(n5427), .Q(WX3910) );
  XOR2X1 U8832 ( .IN1(CRC_OUT_7_29), .IN2(n4703), .Q(n7826) );
  AND2X1 U8833 ( .IN1(n7827), .IN2(n5427), .Q(WX3908) );
  XOR2X1 U8834 ( .IN1(CRC_OUT_7_28), .IN2(n4704), .Q(n7827) );
  AND2X1 U8835 ( .IN1(n7828), .IN2(n5427), .Q(WX3906) );
  XOR2X1 U8836 ( .IN1(test_so32), .IN2(n4705), .Q(n7828) );
  AND2X1 U8837 ( .IN1(n7829), .IN2(n5427), .Q(WX3904) );
  XOR2X1 U8838 ( .IN1(CRC_OUT_7_26), .IN2(n4706), .Q(n7829) );
  AND2X1 U8839 ( .IN1(n7830), .IN2(n5427), .Q(WX3902) );
  XOR2X1 U8840 ( .IN1(CRC_OUT_7_25), .IN2(n4707), .Q(n7830) );
  AND2X1 U8841 ( .IN1(n7831), .IN2(n5427), .Q(WX3900) );
  XOR2X1 U8842 ( .IN1(CRC_OUT_7_24), .IN2(n4708), .Q(n7831) );
  AND2X1 U8843 ( .IN1(n7832), .IN2(n5427), .Q(WX3898) );
  XOR2X1 U8844 ( .IN1(CRC_OUT_7_23), .IN2(n4709), .Q(n7832) );
  AND2X1 U8845 ( .IN1(n7833), .IN2(n5427), .Q(WX3896) );
  XOR2X1 U8846 ( .IN1(test_so29), .IN2(DFF_566_n1), .Q(n7833) );
  AND2X1 U8847 ( .IN1(n7834), .IN2(n5428), .Q(WX3894) );
  XOR2X1 U8848 ( .IN1(CRC_OUT_7_21), .IN2(n4710), .Q(n7834) );
  AND2X1 U8849 ( .IN1(n7835), .IN2(n5428), .Q(WX3892) );
  XOR2X1 U8850 ( .IN1(CRC_OUT_7_20), .IN2(n4711), .Q(n7835) );
  AND2X1 U8851 ( .IN1(n7836), .IN2(n5428), .Q(WX3890) );
  XOR2X1 U8852 ( .IN1(CRC_OUT_7_19), .IN2(n4712), .Q(n7836) );
  AND2X1 U8853 ( .IN1(n7837), .IN2(n5428), .Q(WX3888) );
  XOR2X1 U8854 ( .IN1(CRC_OUT_7_18), .IN2(n4713), .Q(n7837) );
  AND2X1 U8855 ( .IN1(n7838), .IN2(n5428), .Q(WX3886) );
  XOR2X1 U8856 ( .IN1(CRC_OUT_7_17), .IN2(n4714), .Q(n7838) );
  AND2X1 U8857 ( .IN1(n7839), .IN2(n5428), .Q(WX3884) );
  XOR2X1 U8858 ( .IN1(CRC_OUT_7_16), .IN2(n4715), .Q(n7839) );
  AND2X1 U8859 ( .IN1(n7840), .IN2(n5428), .Q(WX3882) );
  XOR2X1 U8860 ( .IN1(DFF_559_n1), .IN2(n7841), .Q(n7840) );
  XOR2X1 U8861 ( .IN1(n4528), .IN2(DFF_575_n1), .Q(n7841) );
  AND2X1 U8862 ( .IN1(n7842), .IN2(n5428), .Q(WX3880) );
  XOR2X1 U8863 ( .IN1(CRC_OUT_7_14), .IN2(n4716), .Q(n7842) );
  AND2X1 U8864 ( .IN1(n7843), .IN2(n5428), .Q(WX3878) );
  XOR2X1 U8865 ( .IN1(CRC_OUT_7_13), .IN2(n4717), .Q(n7843) );
  AND2X1 U8866 ( .IN1(n7844), .IN2(n5429), .Q(WX3876) );
  XOR2X1 U8867 ( .IN1(CRC_OUT_7_12), .IN2(n4718), .Q(n7844) );
  AND2X1 U8868 ( .IN1(n7845), .IN2(n5429), .Q(WX3874) );
  XOR2X1 U8869 ( .IN1(CRC_OUT_7_11), .IN2(n4719), .Q(n7845) );
  AND2X1 U8870 ( .IN1(n7846), .IN2(n5429), .Q(WX3872) );
  XOR2X1 U8871 ( .IN1(CRC_OUT_7_31), .IN2(n7847), .Q(n7846) );
  XOR2X1 U8872 ( .IN1(test_so31), .IN2(n4529), .Q(n7847) );
  AND2X1 U8873 ( .IN1(n7848), .IN2(n5429), .Q(WX3870) );
  XOR2X1 U8874 ( .IN1(CRC_OUT_7_9), .IN2(n4720), .Q(n7848) );
  AND2X1 U8875 ( .IN1(n7849), .IN2(n5429), .Q(WX3868) );
  XOR2X1 U8876 ( .IN1(CRC_OUT_7_8), .IN2(n4721), .Q(n7849) );
  AND2X1 U8877 ( .IN1(n7850), .IN2(n5429), .Q(WX3866) );
  XOR2X1 U8878 ( .IN1(CRC_OUT_7_7), .IN2(n4722), .Q(n7850) );
  AND2X1 U8879 ( .IN1(n7851), .IN2(n5429), .Q(WX3864) );
  XOR2X1 U8880 ( .IN1(CRC_OUT_7_6), .IN2(n4723), .Q(n7851) );
  AND2X1 U8881 ( .IN1(n7852), .IN2(n5429), .Q(WX3862) );
  XOR2X1 U8882 ( .IN1(test_so30), .IN2(DFF_549_n1), .Q(n7852) );
  AND2X1 U8883 ( .IN1(n7853), .IN2(n5429), .Q(WX3860) );
  XOR2X1 U8884 ( .IN1(CRC_OUT_7_4), .IN2(n4724), .Q(n7853) );
  AND2X1 U8885 ( .IN1(n7854), .IN2(n5430), .Q(WX3858) );
  XOR2X1 U8886 ( .IN1(DFF_547_n1), .IN2(n7855), .Q(n7854) );
  XOR2X1 U8887 ( .IN1(n4530), .IN2(DFF_575_n1), .Q(n7855) );
  AND2X1 U8888 ( .IN1(n7856), .IN2(n5430), .Q(WX3856) );
  XOR2X1 U8889 ( .IN1(CRC_OUT_7_2), .IN2(n4725), .Q(n7856) );
  AND2X1 U8890 ( .IN1(n7857), .IN2(n5430), .Q(WX3854) );
  XOR2X1 U8891 ( .IN1(CRC_OUT_7_1), .IN2(n4726), .Q(n7857) );
  AND2X1 U8892 ( .IN1(n7858), .IN2(n5430), .Q(WX3852) );
  XOR2X1 U8893 ( .IN1(CRC_OUT_7_0), .IN2(n4727), .Q(n7858) );
  AND2X1 U8894 ( .IN1(n7859), .IN2(n5430), .Q(WX3850) );
  XOR2X1 U8895 ( .IN1(n4540), .IN2(CRC_OUT_7_31), .Q(n7859) );
  AND2X1 U8896 ( .IN1(test_so24), .IN2(n5430), .Q(WX3324) );
  INVX0 U8897 ( .INP(n7860), .ZN(WX3322) );
  OR2X1 U8898 ( .IN1(n5485), .IN2(n9724), .Q(n7860) );
  INVX0 U8899 ( .INP(n7861), .ZN(WX3320) );
  OR2X1 U8900 ( .IN1(n5485), .IN2(n9727), .Q(n7861) );
  INVX0 U8901 ( .INP(n7862), .ZN(WX3318) );
  OR2X1 U8902 ( .IN1(n5485), .IN2(n9728), .Q(n7862) );
  INVX0 U8903 ( .INP(n7863), .ZN(WX3316) );
  OR2X1 U8904 ( .IN1(n5485), .IN2(n9729), .Q(n7863) );
  INVX0 U8905 ( .INP(n7864), .ZN(WX3314) );
  OR2X1 U8906 ( .IN1(n5485), .IN2(n9730), .Q(n7864) );
  INVX0 U8907 ( .INP(n7865), .ZN(WX3312) );
  OR2X1 U8908 ( .IN1(n5485), .IN2(n9731), .Q(n7865) );
  INVX0 U8909 ( .INP(n7866), .ZN(WX3310) );
  OR2X1 U8910 ( .IN1(n5485), .IN2(n9732), .Q(n7866) );
  INVX0 U8911 ( .INP(n7867), .ZN(WX3308) );
  OR2X1 U8912 ( .IN1(n5485), .IN2(n9733), .Q(n7867) );
  INVX0 U8913 ( .INP(n7868), .ZN(WX3306) );
  OR2X1 U8914 ( .IN1(n5485), .IN2(n9734), .Q(n7868) );
  INVX0 U8915 ( .INP(n7869), .ZN(WX3304) );
  OR2X1 U8916 ( .IN1(n5485), .IN2(n9735), .Q(n7869) );
  INVX0 U8917 ( .INP(n7870), .ZN(WX3302) );
  OR2X1 U8918 ( .IN1(n5486), .IN2(n9738), .Q(n7870) );
  INVX0 U8919 ( .INP(n7871), .ZN(WX3300) );
  OR2X1 U8920 ( .IN1(n5486), .IN2(n9739), .Q(n7871) );
  INVX0 U8921 ( .INP(n7872), .ZN(WX3298) );
  OR2X1 U8922 ( .IN1(n5486), .IN2(n9740), .Q(n7872) );
  INVX0 U8923 ( .INP(n7873), .ZN(WX3296) );
  OR2X1 U8924 ( .IN1(n5486), .IN2(n9741), .Q(n7873) );
  INVX0 U8925 ( .INP(n7874), .ZN(WX3294) );
  OR2X1 U8926 ( .IN1(n5486), .IN2(n9744), .Q(n7874) );
  OR2X1 U8927 ( .IN1(n7875), .IN2(n7876), .Q(WX3292) );
  OR2X1 U8928 ( .IN1(n7877), .IN2(n7878), .Q(n7876) );
  AND2X1 U8929 ( .IN1(n4891), .IN2(CRC_OUT_7_0), .Q(n7878) );
  AND2X1 U8930 ( .IN1(n126), .IN2(n4868), .Q(n7877) );
  INVX0 U8931 ( .INP(n7879), .ZN(n126) );
  OR2X1 U8932 ( .IN1(n5486), .IN2(n3972), .Q(n7879) );
  OR2X1 U8933 ( .IN1(n7880), .IN2(n7881), .Q(n7875) );
  AND2X1 U8934 ( .IN1(n4851), .IN2(n7882), .Q(n7881) );
  AND2X1 U8935 ( .IN1(n7497), .IN2(n4918), .Q(n7880) );
  XOR2X1 U8936 ( .IN1(n7883), .IN2(n7884), .Q(n7497) );
  XOR2X1 U8937 ( .IN1(test_so36), .IN2(n9659), .Q(n7884) );
  XOR2X1 U8938 ( .IN1(WX4714), .IN2(n4539), .Q(n7883) );
  OR2X1 U8939 ( .IN1(n7885), .IN2(n7886), .Q(WX3290) );
  OR2X1 U8940 ( .IN1(n7887), .IN2(n7888), .Q(n7886) );
  AND2X1 U8941 ( .IN1(n4891), .IN2(CRC_OUT_7_1), .Q(n7888) );
  AND2X1 U8942 ( .IN1(n125), .IN2(n4868), .Q(n7887) );
  INVX0 U8943 ( .INP(n7889), .ZN(n125) );
  OR2X1 U8944 ( .IN1(n5486), .IN2(n3973), .Q(n7889) );
  OR2X1 U8945 ( .IN1(n7890), .IN2(n7891), .Q(n7885) );
  AND2X1 U8946 ( .IN1(n4851), .IN2(n7892), .Q(n7891) );
  AND2X1 U8947 ( .IN1(n4926), .IN2(n7507), .Q(n7890) );
  XNOR2X1 U8948 ( .IN1(n7893), .IN2(n7894), .Q(n7507) );
  XOR2X1 U8949 ( .IN1(n9660), .IN2(n4701), .Q(n7894) );
  XOR2X1 U8950 ( .IN1(WX4584), .IN2(n4427), .Q(n7893) );
  OR2X1 U8951 ( .IN1(n7895), .IN2(n7896), .Q(WX3288) );
  OR2X1 U8952 ( .IN1(n7897), .IN2(n7898), .Q(n7896) );
  AND2X1 U8953 ( .IN1(n4891), .IN2(CRC_OUT_7_2), .Q(n7898) );
  AND2X1 U8954 ( .IN1(n124), .IN2(n4868), .Q(n7897) );
  INVX0 U8955 ( .INP(n7899), .ZN(n124) );
  OR2X1 U8956 ( .IN1(n5486), .IN2(n3974), .Q(n7899) );
  OR2X1 U8957 ( .IN1(n7900), .IN2(n7901), .Q(n7895) );
  AND2X1 U8958 ( .IN1(n4851), .IN2(n7902), .Q(n7901) );
  AND2X1 U8959 ( .IN1(n4926), .IN2(n7517), .Q(n7900) );
  XNOR2X1 U8960 ( .IN1(n7903), .IN2(n7904), .Q(n7517) );
  XOR2X1 U8961 ( .IN1(n9661), .IN2(n4700), .Q(n7904) );
  XOR2X1 U8962 ( .IN1(WX4582), .IN2(n4429), .Q(n7903) );
  OR2X1 U8963 ( .IN1(n7905), .IN2(n7906), .Q(WX3286) );
  OR2X1 U8964 ( .IN1(n7907), .IN2(n7908), .Q(n7906) );
  AND2X1 U8965 ( .IN1(n4892), .IN2(CRC_OUT_7_3), .Q(n7908) );
  AND2X1 U8966 ( .IN1(n123), .IN2(n4868), .Q(n7907) );
  INVX0 U8967 ( .INP(n7909), .ZN(n123) );
  OR2X1 U8968 ( .IN1(n5486), .IN2(n3975), .Q(n7909) );
  OR2X1 U8969 ( .IN1(n7910), .IN2(n7911), .Q(n7905) );
  AND2X1 U8970 ( .IN1(n4851), .IN2(n7912), .Q(n7911) );
  AND2X1 U8971 ( .IN1(n4926), .IN2(n7527), .Q(n7910) );
  XNOR2X1 U8972 ( .IN1(n7913), .IN2(n7914), .Q(n7527) );
  XOR2X1 U8973 ( .IN1(n9662), .IN2(n4699), .Q(n7914) );
  XOR2X1 U8974 ( .IN1(WX4580), .IN2(n4431), .Q(n7913) );
  OR2X1 U8975 ( .IN1(n7915), .IN2(n7916), .Q(WX3284) );
  OR2X1 U8976 ( .IN1(n7917), .IN2(n7918), .Q(n7916) );
  AND2X1 U8977 ( .IN1(n4891), .IN2(CRC_OUT_7_4), .Q(n7918) );
  AND2X1 U8978 ( .IN1(n122), .IN2(n4868), .Q(n7917) );
  INVX0 U8979 ( .INP(n7919), .ZN(n122) );
  OR2X1 U8980 ( .IN1(n5486), .IN2(n3976), .Q(n7919) );
  OR2X1 U8981 ( .IN1(n7920), .IN2(n7921), .Q(n7915) );
  AND2X1 U8982 ( .IN1(n4851), .IN2(n7922), .Q(n7921) );
  AND2X1 U8983 ( .IN1(n4926), .IN2(n7537), .Q(n7920) );
  XNOR2X1 U8984 ( .IN1(n7923), .IN2(n7924), .Q(n7537) );
  XOR2X1 U8985 ( .IN1(n9663), .IN2(n4527), .Q(n7924) );
  XOR2X1 U8986 ( .IN1(WX4578), .IN2(n4433), .Q(n7923) );
  OR2X1 U8987 ( .IN1(n7925), .IN2(n7926), .Q(WX3282) );
  OR2X1 U8988 ( .IN1(n7927), .IN2(n7928), .Q(n7926) );
  AND2X1 U8989 ( .IN1(n4892), .IN2(CRC_OUT_7_5), .Q(n7928) );
  AND2X1 U8990 ( .IN1(n121), .IN2(n4868), .Q(n7927) );
  INVX0 U8991 ( .INP(n7929), .ZN(n121) );
  OR2X1 U8992 ( .IN1(n5486), .IN2(n3977), .Q(n7929) );
  OR2X1 U8993 ( .IN1(n7930), .IN2(n7931), .Q(n7925) );
  AND2X1 U8994 ( .IN1(n4851), .IN2(n7932), .Q(n7931) );
  AND2X1 U8995 ( .IN1(n4926), .IN2(n7547), .Q(n7930) );
  XNOR2X1 U8996 ( .IN1(n7933), .IN2(n7934), .Q(n7547) );
  XOR2X1 U8997 ( .IN1(n9664), .IN2(n4698), .Q(n7934) );
  XOR2X1 U8998 ( .IN1(WX4576), .IN2(n4435), .Q(n7933) );
  OR2X1 U8999 ( .IN1(n7935), .IN2(n7936), .Q(WX3280) );
  OR2X1 U9000 ( .IN1(n7937), .IN2(n7938), .Q(n7936) );
  AND2X1 U9001 ( .IN1(n4891), .IN2(CRC_OUT_7_6), .Q(n7938) );
  AND2X1 U9002 ( .IN1(n120), .IN2(n4868), .Q(n7937) );
  INVX0 U9003 ( .INP(n7939), .ZN(n120) );
  OR2X1 U9004 ( .IN1(n5486), .IN2(n3978), .Q(n7939) );
  OR2X1 U9005 ( .IN1(n7940), .IN2(n7941), .Q(n7935) );
  AND2X1 U9006 ( .IN1(n7942), .IN2(n4835), .Q(n7941) );
  AND2X1 U9007 ( .IN1(n4926), .IN2(n7557), .Q(n7940) );
  XNOR2X1 U9008 ( .IN1(n7943), .IN2(n7944), .Q(n7557) );
  XOR2X1 U9009 ( .IN1(n9665), .IN2(n4697), .Q(n7944) );
  XOR2X1 U9010 ( .IN1(WX4574), .IN2(n4437), .Q(n7943) );
  OR2X1 U9011 ( .IN1(n7945), .IN2(n7946), .Q(WX3278) );
  OR2X1 U9012 ( .IN1(n7947), .IN2(n7948), .Q(n7946) );
  AND2X1 U9013 ( .IN1(n4891), .IN2(CRC_OUT_7_7), .Q(n7948) );
  AND2X1 U9014 ( .IN1(n119), .IN2(n4868), .Q(n7947) );
  INVX0 U9015 ( .INP(n7949), .ZN(n119) );
  OR2X1 U9016 ( .IN1(n5486), .IN2(n3979), .Q(n7949) );
  OR2X1 U9017 ( .IN1(n7950), .IN2(n7951), .Q(n7945) );
  AND2X1 U9018 ( .IN1(n4851), .IN2(n7952), .Q(n7951) );
  AND2X1 U9019 ( .IN1(n4926), .IN2(n7567), .Q(n7950) );
  XNOR2X1 U9020 ( .IN1(n7953), .IN2(n7954), .Q(n7567) );
  XOR2X1 U9021 ( .IN1(n9666), .IN2(n4696), .Q(n7954) );
  XOR2X1 U9022 ( .IN1(WX4572), .IN2(n4439), .Q(n7953) );
  OR2X1 U9023 ( .IN1(n7955), .IN2(n7956), .Q(WX3276) );
  OR2X1 U9024 ( .IN1(n7957), .IN2(n7958), .Q(n7956) );
  AND2X1 U9025 ( .IN1(n4892), .IN2(CRC_OUT_7_8), .Q(n7958) );
  AND2X1 U9026 ( .IN1(n118), .IN2(n4868), .Q(n7957) );
  INVX0 U9027 ( .INP(n7959), .ZN(n118) );
  OR2X1 U9028 ( .IN1(n5480), .IN2(n3980), .Q(n7959) );
  OR2X1 U9029 ( .IN1(n7960), .IN2(n7961), .Q(n7955) );
  AND2X1 U9030 ( .IN1(n7962), .IN2(n4836), .Q(n7961) );
  AND2X1 U9031 ( .IN1(n4926), .IN2(n7577), .Q(n7960) );
  XNOR2X1 U9032 ( .IN1(n7963), .IN2(n7964), .Q(n7577) );
  XOR2X1 U9033 ( .IN1(n9667), .IN2(n4695), .Q(n7964) );
  XOR2X1 U9034 ( .IN1(WX4570), .IN2(n4441), .Q(n7963) );
  OR2X1 U9035 ( .IN1(n7965), .IN2(n7966), .Q(WX3274) );
  OR2X1 U9036 ( .IN1(n7967), .IN2(n7968), .Q(n7966) );
  AND2X1 U9037 ( .IN1(n4892), .IN2(CRC_OUT_7_9), .Q(n7968) );
  AND2X1 U9038 ( .IN1(n117), .IN2(n4867), .Q(n7967) );
  INVX0 U9039 ( .INP(n7969), .ZN(n117) );
  OR2X1 U9040 ( .IN1(n5480), .IN2(n3981), .Q(n7969) );
  OR2X1 U9041 ( .IN1(n7970), .IN2(n7971), .Q(n7965) );
  AND2X1 U9042 ( .IN1(n4850), .IN2(n7972), .Q(n7971) );
  AND2X1 U9043 ( .IN1(n4927), .IN2(n7587), .Q(n7970) );
  XNOR2X1 U9044 ( .IN1(n7973), .IN2(n7974), .Q(n7587) );
  XOR2X1 U9045 ( .IN1(n9668), .IN2(n4694), .Q(n7974) );
  XOR2X1 U9046 ( .IN1(WX4568), .IN2(n4443), .Q(n7973) );
  OR2X1 U9047 ( .IN1(n7975), .IN2(n7976), .Q(WX3272) );
  OR2X1 U9048 ( .IN1(n7977), .IN2(n7978), .Q(n7976) );
  AND2X1 U9049 ( .IN1(test_so31), .IN2(n4888), .Q(n7978) );
  AND2X1 U9050 ( .IN1(n116), .IN2(n4867), .Q(n7977) );
  INVX0 U9051 ( .INP(n7979), .ZN(n116) );
  OR2X1 U9052 ( .IN1(n5480), .IN2(n3982), .Q(n7979) );
  OR2X1 U9053 ( .IN1(n7980), .IN2(n7981), .Q(n7975) );
  AND2X1 U9054 ( .IN1(n4850), .IN2(n7982), .Q(n7981) );
  AND2X1 U9055 ( .IN1(n4927), .IN2(n7597), .Q(n7980) );
  XNOR2X1 U9056 ( .IN1(n7983), .IN2(n7984), .Q(n7597) );
  XOR2X1 U9057 ( .IN1(n9669), .IN2(n4693), .Q(n7984) );
  XOR2X1 U9058 ( .IN1(WX4566), .IN2(n4445), .Q(n7983) );
  OR2X1 U9059 ( .IN1(n7985), .IN2(n7986), .Q(WX3270) );
  OR2X1 U9060 ( .IN1(n7987), .IN2(n7988), .Q(n7986) );
  AND2X1 U9061 ( .IN1(n4892), .IN2(CRC_OUT_7_11), .Q(n7988) );
  AND2X1 U9062 ( .IN1(n115), .IN2(n4867), .Q(n7987) );
  INVX0 U9063 ( .INP(n7989), .ZN(n115) );
  OR2X1 U9064 ( .IN1(n5480), .IN2(n3983), .Q(n7989) );
  OR2X1 U9065 ( .IN1(n7990), .IN2(n7991), .Q(n7985) );
  AND2X1 U9066 ( .IN1(n4850), .IN2(n7992), .Q(n7991) );
  AND2X1 U9067 ( .IN1(n7607), .IN2(n4918), .Q(n7990) );
  XOR2X1 U9068 ( .IN1(n7993), .IN2(n7994), .Q(n7607) );
  XOR2X1 U9069 ( .IN1(test_so41), .IN2(n9670), .Q(n7994) );
  XOR2X1 U9070 ( .IN1(WX4564), .IN2(n4447), .Q(n7993) );
  OR2X1 U9071 ( .IN1(n7995), .IN2(n7996), .Q(WX3268) );
  OR2X1 U9072 ( .IN1(n7997), .IN2(n7998), .Q(n7996) );
  AND2X1 U9073 ( .IN1(n4892), .IN2(CRC_OUT_7_12), .Q(n7998) );
  AND2X1 U9074 ( .IN1(n114), .IN2(n4867), .Q(n7997) );
  INVX0 U9075 ( .INP(n7999), .ZN(n114) );
  OR2X1 U9076 ( .IN1(n5480), .IN2(n3984), .Q(n7999) );
  OR2X1 U9077 ( .IN1(n8000), .IN2(n8001), .Q(n7995) );
  AND2X1 U9078 ( .IN1(n8002), .IN2(n4836), .Q(n8001) );
  AND2X1 U9079 ( .IN1(n4927), .IN2(n7617), .Q(n8000) );
  XNOR2X1 U9080 ( .IN1(n8003), .IN2(n8004), .Q(n7617) );
  XOR2X1 U9081 ( .IN1(n9671), .IN2(n4692), .Q(n8004) );
  XOR2X1 U9082 ( .IN1(WX4562), .IN2(n4449), .Q(n8003) );
  OR2X1 U9083 ( .IN1(n8005), .IN2(n8006), .Q(WX3266) );
  OR2X1 U9084 ( .IN1(n8007), .IN2(n8008), .Q(n8006) );
  AND2X1 U9085 ( .IN1(n4892), .IN2(CRC_OUT_7_13), .Q(n8008) );
  AND2X1 U9086 ( .IN1(n113), .IN2(n4867), .Q(n8007) );
  INVX0 U9087 ( .INP(n8009), .ZN(n113) );
  OR2X1 U9088 ( .IN1(n5480), .IN2(n3985), .Q(n8009) );
  OR2X1 U9089 ( .IN1(n8010), .IN2(n8011), .Q(n8005) );
  AND2X1 U9090 ( .IN1(n4850), .IN2(n8012), .Q(n8011) );
  AND2X1 U9091 ( .IN1(n7627), .IN2(n4918), .Q(n8010) );
  XOR2X1 U9092 ( .IN1(n8013), .IN2(n8014), .Q(n7627) );
  XOR2X1 U9093 ( .IN1(test_so39), .IN2(n9672), .Q(n8014) );
  XOR2X1 U9094 ( .IN1(WX4560), .IN2(n4691), .Q(n8013) );
  OR2X1 U9095 ( .IN1(n8015), .IN2(n8016), .Q(WX3264) );
  OR2X1 U9096 ( .IN1(n8017), .IN2(n8018), .Q(n8016) );
  AND2X1 U9097 ( .IN1(n4892), .IN2(CRC_OUT_7_14), .Q(n8018) );
  AND2X1 U9098 ( .IN1(n112), .IN2(n4867), .Q(n8017) );
  INVX0 U9099 ( .INP(n8019), .ZN(n112) );
  OR2X1 U9100 ( .IN1(n5479), .IN2(n3986), .Q(n8019) );
  OR2X1 U9101 ( .IN1(n8020), .IN2(n8021), .Q(n8015) );
  AND2X1 U9102 ( .IN1(n4850), .IN2(n8022), .Q(n8021) );
  AND2X1 U9103 ( .IN1(n4927), .IN2(n7637), .Q(n8020) );
  XNOR2X1 U9104 ( .IN1(n8023), .IN2(n8024), .Q(n7637) );
  XOR2X1 U9105 ( .IN1(n9673), .IN2(n4690), .Q(n8024) );
  XOR2X1 U9106 ( .IN1(WX4558), .IN2(n4452), .Q(n8023) );
  OR2X1 U9107 ( .IN1(n8025), .IN2(n8026), .Q(WX3262) );
  OR2X1 U9108 ( .IN1(n8027), .IN2(n8028), .Q(n8026) );
  AND2X1 U9109 ( .IN1(n4892), .IN2(CRC_OUT_7_15), .Q(n8028) );
  AND2X1 U9110 ( .IN1(n110), .IN2(n4867), .Q(n8027) );
  INVX0 U9111 ( .INP(n8029), .ZN(n110) );
  OR2X1 U9112 ( .IN1(n5479), .IN2(n3987), .Q(n8029) );
  OR2X1 U9113 ( .IN1(n8030), .IN2(n8031), .Q(n8025) );
  AND2X1 U9114 ( .IN1(n4850), .IN2(n8032), .Q(n8031) );
  AND2X1 U9115 ( .IN1(n7647), .IN2(n4918), .Q(n8030) );
  XOR2X1 U9116 ( .IN1(n8033), .IN2(n8034), .Q(n7647) );
  XOR2X1 U9117 ( .IN1(test_so37), .IN2(n9674), .Q(n8034) );
  XOR2X1 U9118 ( .IN1(WX4556), .IN2(n4689), .Q(n8033) );
  OR2X1 U9119 ( .IN1(n8035), .IN2(n8036), .Q(WX3260) );
  OR2X1 U9120 ( .IN1(n8037), .IN2(n8038), .Q(n8036) );
  AND2X1 U9121 ( .IN1(n4892), .IN2(CRC_OUT_7_16), .Q(n8038) );
  AND2X1 U9122 ( .IN1(n109), .IN2(n4867), .Q(n8037) );
  INVX0 U9123 ( .INP(n8039), .ZN(n109) );
  OR2X1 U9124 ( .IN1(n5479), .IN2(n3988), .Q(n8039) );
  OR2X1 U9125 ( .IN1(n8040), .IN2(n8041), .Q(n8035) );
  AND2X1 U9126 ( .IN1(n8042), .IN2(n4837), .Q(n8041) );
  AND2X1 U9127 ( .IN1(n4927), .IN2(n7657), .Q(n8040) );
  XNOR2X1 U9128 ( .IN1(n8043), .IN2(n8044), .Q(n7657) );
  XOR2X1 U9129 ( .IN1(n4238), .IN2(n5384), .Q(n8044) );
  XOR2X1 U9130 ( .IN1(n8045), .IN2(n4526), .Q(n8043) );
  XOR2X1 U9131 ( .IN1(WX4682), .IN2(n9675), .Q(n8045) );
  OR2X1 U9132 ( .IN1(n8046), .IN2(n8047), .Q(WX3258) );
  OR2X1 U9133 ( .IN1(n8048), .IN2(n8049), .Q(n8047) );
  AND2X1 U9134 ( .IN1(n4892), .IN2(CRC_OUT_7_17), .Q(n8049) );
  AND2X1 U9135 ( .IN1(n108), .IN2(n4867), .Q(n8048) );
  INVX0 U9136 ( .INP(n8050), .ZN(n108) );
  OR2X1 U9137 ( .IN1(n5479), .IN2(n3989), .Q(n8050) );
  OR2X1 U9138 ( .IN1(n8051), .IN2(n8052), .Q(n8046) );
  AND2X1 U9139 ( .IN1(n4850), .IN2(n8053), .Q(n8052) );
  AND2X1 U9140 ( .IN1(n7668), .IN2(n4918), .Q(n8051) );
  XOR2X1 U9141 ( .IN1(n8054), .IN2(n8055), .Q(n7668) );
  XOR2X1 U9142 ( .IN1(n4239), .IN2(n5384), .Q(n8055) );
  XOR2X1 U9143 ( .IN1(n8056), .IN2(n4688), .Q(n8054) );
  XOR2X1 U9144 ( .IN1(WX4616), .IN2(test_so35), .Q(n8056) );
  OR2X1 U9145 ( .IN1(n8057), .IN2(n8058), .Q(WX3256) );
  OR2X1 U9146 ( .IN1(n8059), .IN2(n8060), .Q(n8058) );
  AND2X1 U9147 ( .IN1(n4893), .IN2(CRC_OUT_7_18), .Q(n8060) );
  AND2X1 U9148 ( .IN1(n107), .IN2(n4867), .Q(n8059) );
  INVX0 U9149 ( .INP(n8061), .ZN(n107) );
  OR2X1 U9150 ( .IN1(n5479), .IN2(n3990), .Q(n8061) );
  OR2X1 U9151 ( .IN1(n8062), .IN2(n8063), .Q(n8057) );
  AND2X1 U9152 ( .IN1(n4850), .IN2(n8064), .Q(n8063) );
  AND2X1 U9153 ( .IN1(n4927), .IN2(n7679), .Q(n8062) );
  XNOR2X1 U9154 ( .IN1(n8065), .IN2(n8066), .Q(n7679) );
  XOR2X1 U9155 ( .IN1(n4240), .IN2(n5384), .Q(n8066) );
  XOR2X1 U9156 ( .IN1(n8067), .IN2(n4687), .Q(n8065) );
  XOR2X1 U9157 ( .IN1(WX4678), .IN2(n9676), .Q(n8067) );
  OR2X1 U9158 ( .IN1(n8068), .IN2(n8069), .Q(WX3254) );
  OR2X1 U9159 ( .IN1(n8070), .IN2(n8071), .Q(n8069) );
  AND2X1 U9160 ( .IN1(n4892), .IN2(CRC_OUT_7_19), .Q(n8071) );
  AND2X1 U9161 ( .IN1(n106), .IN2(n4867), .Q(n8070) );
  INVX0 U9162 ( .INP(n8072), .ZN(n106) );
  OR2X1 U9163 ( .IN1(n5479), .IN2(n3991), .Q(n8072) );
  OR2X1 U9164 ( .IN1(n8073), .IN2(n8074), .Q(n8068) );
  AND2X1 U9165 ( .IN1(n4850), .IN2(n8075), .Q(n8074) );
  AND2X1 U9166 ( .IN1(n4927), .IN2(n7690), .Q(n8073) );
  XNOR2X1 U9167 ( .IN1(n8076), .IN2(n8077), .Q(n7690) );
  XOR2X1 U9168 ( .IN1(n4241), .IN2(n5384), .Q(n8077) );
  XOR2X1 U9169 ( .IN1(n8078), .IN2(n4686), .Q(n8076) );
  XOR2X1 U9170 ( .IN1(WX4676), .IN2(n9677), .Q(n8078) );
  OR2X1 U9171 ( .IN1(n8079), .IN2(n8080), .Q(WX3252) );
  OR2X1 U9172 ( .IN1(n8081), .IN2(n8082), .Q(n8080) );
  AND2X1 U9173 ( .IN1(n4893), .IN2(CRC_OUT_7_20), .Q(n8082) );
  AND2X1 U9174 ( .IN1(n105), .IN2(n4867), .Q(n8081) );
  INVX0 U9175 ( .INP(n8083), .ZN(n105) );
  OR2X1 U9176 ( .IN1(n5479), .IN2(n3992), .Q(n8083) );
  OR2X1 U9177 ( .IN1(n8084), .IN2(n8085), .Q(n8079) );
  AND2X1 U9178 ( .IN1(n4850), .IN2(n8086), .Q(n8085) );
  AND2X1 U9179 ( .IN1(n4927), .IN2(n7701), .Q(n8084) );
  XNOR2X1 U9180 ( .IN1(n8087), .IN2(n8088), .Q(n7701) );
  XOR2X1 U9181 ( .IN1(n4242), .IN2(n5384), .Q(n8088) );
  XOR2X1 U9182 ( .IN1(n8089), .IN2(n4685), .Q(n8087) );
  XOR2X1 U9183 ( .IN1(WX4674), .IN2(n9678), .Q(n8089) );
  OR2X1 U9184 ( .IN1(n8090), .IN2(n8091), .Q(WX3250) );
  OR2X1 U9185 ( .IN1(n8092), .IN2(n8093), .Q(n8091) );
  AND2X1 U9186 ( .IN1(n4893), .IN2(CRC_OUT_7_21), .Q(n8093) );
  AND2X1 U9187 ( .IN1(n104), .IN2(n4866), .Q(n8092) );
  INVX0 U9188 ( .INP(n8094), .ZN(n104) );
  OR2X1 U9189 ( .IN1(n5479), .IN2(n3993), .Q(n8094) );
  OR2X1 U9190 ( .IN1(n8095), .IN2(n8096), .Q(n8090) );
  AND2X1 U9191 ( .IN1(n4850), .IN2(n8097), .Q(n8096) );
  AND2X1 U9192 ( .IN1(n4927), .IN2(n7712), .Q(n8095) );
  XNOR2X1 U9193 ( .IN1(n8098), .IN2(n8099), .Q(n7712) );
  XOR2X1 U9194 ( .IN1(n4243), .IN2(n5384), .Q(n8099) );
  XOR2X1 U9195 ( .IN1(n8100), .IN2(n4684), .Q(n8098) );
  XOR2X1 U9196 ( .IN1(WX4672), .IN2(n9679), .Q(n8100) );
  OR2X1 U9197 ( .IN1(n8101), .IN2(n8102), .Q(WX3248) );
  OR2X1 U9198 ( .IN1(n8103), .IN2(n8104), .Q(n8102) );
  AND2X1 U9199 ( .IN1(n4893), .IN2(CRC_OUT_7_22), .Q(n8104) );
  AND2X1 U9200 ( .IN1(n103), .IN2(n4866), .Q(n8103) );
  INVX0 U9201 ( .INP(n8105), .ZN(n103) );
  OR2X1 U9202 ( .IN1(n5479), .IN2(n3994), .Q(n8105) );
  OR2X1 U9203 ( .IN1(n8106), .IN2(n8107), .Q(n8101) );
  AND2X1 U9204 ( .IN1(n4850), .IN2(n8108), .Q(n8107) );
  AND2X1 U9205 ( .IN1(n4927), .IN2(n7723), .Q(n8106) );
  XNOR2X1 U9206 ( .IN1(n8109), .IN2(n8110), .Q(n7723) );
  XOR2X1 U9207 ( .IN1(n4244), .IN2(n5384), .Q(n8110) );
  XOR2X1 U9208 ( .IN1(n8111), .IN2(n4683), .Q(n8109) );
  XOR2X1 U9209 ( .IN1(WX4670), .IN2(n9680), .Q(n8111) );
  OR2X1 U9210 ( .IN1(n8112), .IN2(n8113), .Q(WX3246) );
  OR2X1 U9211 ( .IN1(n8114), .IN2(n8115), .Q(n8113) );
  AND2X1 U9212 ( .IN1(n4898), .IN2(CRC_OUT_7_23), .Q(n8115) );
  AND2X1 U9213 ( .IN1(n102), .IN2(n4866), .Q(n8114) );
  INVX0 U9214 ( .INP(n8116), .ZN(n102) );
  OR2X1 U9215 ( .IN1(n5479), .IN2(n3995), .Q(n8116) );
  OR2X1 U9216 ( .IN1(n8117), .IN2(n8118), .Q(n8112) );
  AND2X1 U9217 ( .IN1(n8119), .IN2(n4838), .Q(n8118) );
  AND2X1 U9218 ( .IN1(n4930), .IN2(n7734), .Q(n8117) );
  XNOR2X1 U9219 ( .IN1(n8120), .IN2(n8121), .Q(n7734) );
  XOR2X1 U9220 ( .IN1(n4245), .IN2(n5384), .Q(n8121) );
  XOR2X1 U9221 ( .IN1(n8122), .IN2(n4682), .Q(n8120) );
  XOR2X1 U9222 ( .IN1(WX4668), .IN2(n9681), .Q(n8122) );
  OR2X1 U9223 ( .IN1(n8123), .IN2(n8124), .Q(WX3244) );
  OR2X1 U9224 ( .IN1(n8125), .IN2(n8126), .Q(n8124) );
  AND2X1 U9225 ( .IN1(n4893), .IN2(CRC_OUT_7_24), .Q(n8126) );
  AND2X1 U9226 ( .IN1(n101), .IN2(n4866), .Q(n8125) );
  INVX0 U9227 ( .INP(n8127), .ZN(n101) );
  OR2X1 U9228 ( .IN1(n5479), .IN2(n3996), .Q(n8127) );
  OR2X1 U9229 ( .IN1(n8128), .IN2(n8129), .Q(n8123) );
  AND2X1 U9230 ( .IN1(n4849), .IN2(n8130), .Q(n8129) );
  AND2X1 U9231 ( .IN1(n4927), .IN2(n7745), .Q(n8128) );
  XNOR2X1 U9232 ( .IN1(n8131), .IN2(n8132), .Q(n7745) );
  XOR2X1 U9233 ( .IN1(n4246), .IN2(n5383), .Q(n8132) );
  XOR2X1 U9234 ( .IN1(n8133), .IN2(n4681), .Q(n8131) );
  XOR2X1 U9235 ( .IN1(WX4666), .IN2(n9682), .Q(n8133) );
  OR2X1 U9236 ( .IN1(n8134), .IN2(n8135), .Q(WX3242) );
  OR2X1 U9237 ( .IN1(n8136), .IN2(n8137), .Q(n8135) );
  AND2X1 U9238 ( .IN1(n4893), .IN2(CRC_OUT_7_25), .Q(n8137) );
  AND2X1 U9239 ( .IN1(n100), .IN2(n4866), .Q(n8136) );
  INVX0 U9240 ( .INP(n8138), .ZN(n100) );
  OR2X1 U9241 ( .IN1(n5479), .IN2(n3997), .Q(n8138) );
  OR2X1 U9242 ( .IN1(n8139), .IN2(n8140), .Q(n8134) );
  AND2X1 U9243 ( .IN1(n4849), .IN2(n8141), .Q(n8140) );
  AND2X1 U9244 ( .IN1(n4927), .IN2(n7756), .Q(n8139) );
  XNOR2X1 U9245 ( .IN1(n8142), .IN2(n8143), .Q(n7756) );
  XOR2X1 U9246 ( .IN1(n4247), .IN2(n5383), .Q(n8143) );
  XOR2X1 U9247 ( .IN1(n8144), .IN2(n4680), .Q(n8142) );
  XOR2X1 U9248 ( .IN1(WX4664), .IN2(n9683), .Q(n8144) );
  OR2X1 U9249 ( .IN1(n8145), .IN2(n8146), .Q(WX3240) );
  OR2X1 U9250 ( .IN1(n8147), .IN2(n8148), .Q(n8146) );
  AND2X1 U9251 ( .IN1(n4893), .IN2(CRC_OUT_7_26), .Q(n8148) );
  AND2X1 U9252 ( .IN1(n99), .IN2(n4866), .Q(n8147) );
  INVX0 U9253 ( .INP(n8149), .ZN(n99) );
  OR2X1 U9254 ( .IN1(n5479), .IN2(n3998), .Q(n8149) );
  OR2X1 U9255 ( .IN1(n8150), .IN2(n8151), .Q(n8145) );
  AND2X1 U9256 ( .IN1(n8152), .IN2(n4837), .Q(n8151) );
  AND2X1 U9257 ( .IN1(n4927), .IN2(n7767), .Q(n8150) );
  XNOR2X1 U9258 ( .IN1(n8153), .IN2(n8154), .Q(n7767) );
  XOR2X1 U9259 ( .IN1(n4248), .IN2(n5383), .Q(n8154) );
  XOR2X1 U9260 ( .IN1(n8155), .IN2(n4679), .Q(n8153) );
  XOR2X1 U9261 ( .IN1(WX4662), .IN2(n9684), .Q(n8155) );
  OR2X1 U9262 ( .IN1(n8156), .IN2(n8157), .Q(WX3238) );
  OR2X1 U9263 ( .IN1(n8158), .IN2(n8159), .Q(n8157) );
  AND2X1 U9264 ( .IN1(test_so32), .IN2(n4887), .Q(n8159) );
  AND2X1 U9265 ( .IN1(n98), .IN2(n4866), .Q(n8158) );
  INVX0 U9266 ( .INP(n8160), .ZN(n98) );
  OR2X1 U9267 ( .IN1(n5478), .IN2(n3999), .Q(n8160) );
  OR2X1 U9268 ( .IN1(n8161), .IN2(n8162), .Q(n8156) );
  AND2X1 U9269 ( .IN1(n4849), .IN2(n8163), .Q(n8162) );
  AND2X1 U9270 ( .IN1(n4928), .IN2(n7778), .Q(n8161) );
  XNOR2X1 U9271 ( .IN1(n8164), .IN2(n8165), .Q(n7778) );
  XOR2X1 U9272 ( .IN1(n4249), .IN2(n5383), .Q(n8165) );
  XOR2X1 U9273 ( .IN1(n8166), .IN2(n4678), .Q(n8164) );
  XOR2X1 U9274 ( .IN1(WX4660), .IN2(n9685), .Q(n8166) );
  OR2X1 U9275 ( .IN1(n8167), .IN2(n8168), .Q(WX3236) );
  OR2X1 U9276 ( .IN1(n8169), .IN2(n8170), .Q(n8168) );
  AND2X1 U9277 ( .IN1(n4893), .IN2(CRC_OUT_7_28), .Q(n8170) );
  AND2X1 U9278 ( .IN1(n97), .IN2(n4866), .Q(n8169) );
  INVX0 U9279 ( .INP(n8171), .ZN(n97) );
  OR2X1 U9280 ( .IN1(n5478), .IN2(n4000), .Q(n8171) );
  OR2X1 U9281 ( .IN1(n8172), .IN2(n8173), .Q(n8167) );
  AND2X1 U9282 ( .IN1(n4849), .IN2(n8174), .Q(n8173) );
  AND2X1 U9283 ( .IN1(n7789), .IN2(n4919), .Q(n8172) );
  XOR2X1 U9284 ( .IN1(n8175), .IN2(n8176), .Q(n7789) );
  XOR2X1 U9285 ( .IN1(n4250), .IN2(n5383), .Q(n8176) );
  XOR2X1 U9286 ( .IN1(WX4594), .IN2(n8177), .Q(n8175) );
  XOR2X1 U9287 ( .IN1(test_so40), .IN2(n9686), .Q(n8177) );
  OR2X1 U9288 ( .IN1(n8178), .IN2(n8179), .Q(WX3234) );
  OR2X1 U9289 ( .IN1(n8180), .IN2(n8181), .Q(n8179) );
  AND2X1 U9290 ( .IN1(n4893), .IN2(CRC_OUT_7_29), .Q(n8181) );
  AND2X1 U9291 ( .IN1(n96), .IN2(n4866), .Q(n8180) );
  INVX0 U9292 ( .INP(n8182), .ZN(n96) );
  OR2X1 U9293 ( .IN1(n5478), .IN2(n4001), .Q(n8182) );
  OR2X1 U9294 ( .IN1(n8183), .IN2(n8184), .Q(n8178) );
  AND2X1 U9295 ( .IN1(n4849), .IN2(n8185), .Q(n8184) );
  AND2X1 U9296 ( .IN1(n4928), .IN2(n7800), .Q(n8183) );
  XNOR2X1 U9297 ( .IN1(n8186), .IN2(n8187), .Q(n7800) );
  XOR2X1 U9298 ( .IN1(n4251), .IN2(n5383), .Q(n8187) );
  XOR2X1 U9299 ( .IN1(n8188), .IN2(n4677), .Q(n8186) );
  XOR2X1 U9300 ( .IN1(WX4656), .IN2(n9687), .Q(n8188) );
  OR2X1 U9301 ( .IN1(n8189), .IN2(n8190), .Q(WX3232) );
  OR2X1 U9302 ( .IN1(n8191), .IN2(n8192), .Q(n8190) );
  AND2X1 U9303 ( .IN1(n4893), .IN2(CRC_OUT_7_30), .Q(n8192) );
  AND2X1 U9304 ( .IN1(n95), .IN2(n4866), .Q(n8191) );
  INVX0 U9305 ( .INP(n8193), .ZN(n95) );
  OR2X1 U9306 ( .IN1(n5478), .IN2(n4002), .Q(n8193) );
  OR2X1 U9307 ( .IN1(n8194), .IN2(n8195), .Q(n8189) );
  AND2X1 U9308 ( .IN1(n8196), .IN2(n4837), .Q(n8195) );
  AND2X1 U9309 ( .IN1(n7811), .IN2(n4919), .Q(n8194) );
  XOR2X1 U9310 ( .IN1(n8197), .IN2(n8198), .Q(n7811) );
  XOR2X1 U9311 ( .IN1(n4676), .IN2(n5383), .Q(n8198) );
  XOR2X1 U9312 ( .IN1(n8199), .IN2(n9690), .Q(n8197) );
  XOR2X1 U9313 ( .IN1(n9689), .IN2(n9688), .Q(n8199) );
  OR2X1 U9314 ( .IN1(n8200), .IN2(n8201), .Q(WX3230) );
  OR2X1 U9315 ( .IN1(n8202), .IN2(n8203), .Q(n8201) );
  AND2X1 U9316 ( .IN1(n2245), .IN2(WX3071), .Q(n8203) );
  AND2X1 U9317 ( .IN1(n4893), .IN2(CRC_OUT_7_31), .Q(n8202) );
  OR2X1 U9318 ( .IN1(n8204), .IN2(n8205), .Q(n8200) );
  AND2X1 U9319 ( .IN1(n4849), .IN2(n8206), .Q(n8205) );
  AND2X1 U9320 ( .IN1(n4928), .IN2(n7821), .Q(n8204) );
  XNOR2X1 U9321 ( .IN1(n8207), .IN2(n8208), .Q(n7821) );
  XOR2X1 U9322 ( .IN1(n4170), .IN2(n5383), .Q(n8208) );
  XOR2X1 U9323 ( .IN1(n8209), .IN2(n4675), .Q(n8207) );
  XOR2X1 U9324 ( .IN1(WX4652), .IN2(n9691), .Q(n8209) );
  AND2X1 U9325 ( .IN1(n4820), .IN2(n5430), .Q(WX3132) );
  AND2X1 U9326 ( .IN1(n8210), .IN2(n5430), .Q(WX2619) );
  XOR2X1 U9327 ( .IN1(CRC_OUT_8_30), .IN2(n4728), .Q(n8210) );
  AND2X1 U9328 ( .IN1(n8211), .IN2(n5430), .Q(WX2617) );
  XOR2X1 U9329 ( .IN1(CRC_OUT_8_29), .IN2(n4729), .Q(n8211) );
  AND2X1 U9330 ( .IN1(n8212), .IN2(n5431), .Q(WX2615) );
  XOR2X1 U9331 ( .IN1(CRC_OUT_8_28), .IN2(n4730), .Q(n8212) );
  AND2X1 U9332 ( .IN1(n8213), .IN2(n5431), .Q(WX2613) );
  XOR2X1 U9333 ( .IN1(test_so18), .IN2(DFF_379_n1), .Q(n8213) );
  AND2X1 U9334 ( .IN1(n8214), .IN2(n5431), .Q(WX2611) );
  XOR2X1 U9335 ( .IN1(CRC_OUT_8_26), .IN2(n4731), .Q(n8214) );
  AND2X1 U9336 ( .IN1(n8215), .IN2(n5431), .Q(WX2609) );
  XOR2X1 U9337 ( .IN1(test_so21), .IN2(n4732), .Q(n8215) );
  AND2X1 U9338 ( .IN1(n8216), .IN2(n5431), .Q(WX2607) );
  XOR2X1 U9339 ( .IN1(CRC_OUT_8_24), .IN2(n4733), .Q(n8216) );
  AND2X1 U9340 ( .IN1(n8217), .IN2(n5431), .Q(WX2605) );
  XOR2X1 U9341 ( .IN1(CRC_OUT_8_23), .IN2(n4734), .Q(n8217) );
  AND2X1 U9342 ( .IN1(n8218), .IN2(n5431), .Q(WX2603) );
  XOR2X1 U9343 ( .IN1(CRC_OUT_8_22), .IN2(n4735), .Q(n8218) );
  AND2X1 U9344 ( .IN1(n8219), .IN2(n5431), .Q(WX2601) );
  XOR2X1 U9345 ( .IN1(CRC_OUT_8_21), .IN2(n4736), .Q(n8219) );
  AND2X1 U9346 ( .IN1(n8220), .IN2(n5432), .Q(WX2599) );
  XOR2X1 U9347 ( .IN1(CRC_OUT_8_20), .IN2(n4737), .Q(n8220) );
  AND2X1 U9348 ( .IN1(n8221), .IN2(n5432), .Q(WX2597) );
  XOR2X1 U9349 ( .IN1(CRC_OUT_8_19), .IN2(n4738), .Q(n8221) );
  AND2X1 U9350 ( .IN1(n8222), .IN2(n5432), .Q(WX2595) );
  XOR2X1 U9351 ( .IN1(CRC_OUT_8_18), .IN2(n4739), .Q(n8222) );
  AND2X1 U9352 ( .IN1(n8223), .IN2(n5432), .Q(WX2593) );
  XOR2X1 U9353 ( .IN1(CRC_OUT_8_17), .IN2(n4740), .Q(n8223) );
  AND2X1 U9354 ( .IN1(n8224), .IN2(n5432), .Q(WX2591) );
  XOR2X1 U9355 ( .IN1(CRC_OUT_8_16), .IN2(n4741), .Q(n8224) );
  AND2X1 U9356 ( .IN1(n8225), .IN2(n5432), .Q(WX2589) );
  XOR2X1 U9357 ( .IN1(DFF_367_n1), .IN2(n8226), .Q(n8225) );
  XOR2X1 U9358 ( .IN1(n4531), .IN2(DFF_383_n1), .Q(n8226) );
  AND2X1 U9359 ( .IN1(n8227), .IN2(n5432), .Q(WX2587) );
  XOR2X1 U9360 ( .IN1(CRC_OUT_8_14), .IN2(n4742), .Q(n8227) );
  AND2X1 U9361 ( .IN1(n8228), .IN2(n5432), .Q(WX2585) );
  XOR2X1 U9362 ( .IN1(CRC_OUT_8_13), .IN2(n4743), .Q(n8228) );
  AND2X1 U9363 ( .IN1(n8229), .IN2(n5433), .Q(WX2583) );
  XOR2X1 U9364 ( .IN1(CRC_OUT_8_12), .IN2(n4744), .Q(n8229) );
  AND2X1 U9365 ( .IN1(n8230), .IN2(n5434), .Q(WX2581) );
  XOR2X1 U9366 ( .IN1(CRC_OUT_8_11), .IN2(n4745), .Q(n8230) );
  AND2X1 U9367 ( .IN1(n8231), .IN2(n5433), .Q(WX2579) );
  XOR2X1 U9368 ( .IN1(DFF_362_n1), .IN2(n8232), .Q(n8231) );
  XOR2X1 U9369 ( .IN1(n4532), .IN2(DFF_383_n1), .Q(n8232) );
  AND2X1 U9370 ( .IN1(n8233), .IN2(n5433), .Q(WX2577) );
  XOR2X1 U9371 ( .IN1(test_so19), .IN2(DFF_361_n1), .Q(n8233) );
  AND2X1 U9372 ( .IN1(n8234), .IN2(n5434), .Q(WX2575) );
  XOR2X1 U9373 ( .IN1(CRC_OUT_8_8), .IN2(n4746), .Q(n8234) );
  AND2X1 U9374 ( .IN1(n8235), .IN2(n5433), .Q(WX2573) );
  XOR2X1 U9375 ( .IN1(test_so20), .IN2(n4747), .Q(n8235) );
  AND2X1 U9376 ( .IN1(n8236), .IN2(n5432), .Q(WX2571) );
  XOR2X1 U9377 ( .IN1(CRC_OUT_8_6), .IN2(n4748), .Q(n8236) );
  AND2X1 U9378 ( .IN1(n8237), .IN2(n5433), .Q(WX2569) );
  XOR2X1 U9379 ( .IN1(CRC_OUT_8_5), .IN2(n4749), .Q(n8237) );
  AND2X1 U9380 ( .IN1(n8238), .IN2(n5434), .Q(WX2567) );
  XOR2X1 U9381 ( .IN1(CRC_OUT_8_4), .IN2(n4750), .Q(n8238) );
  AND2X1 U9382 ( .IN1(n8239), .IN2(n5433), .Q(WX2565) );
  XOR2X1 U9383 ( .IN1(DFF_355_n1), .IN2(n8240), .Q(n8239) );
  XOR2X1 U9384 ( .IN1(n4533), .IN2(DFF_383_n1), .Q(n8240) );
  AND2X1 U9385 ( .IN1(n8241), .IN2(n5434), .Q(WX2563) );
  XOR2X1 U9386 ( .IN1(CRC_OUT_8_2), .IN2(n4751), .Q(n8241) );
  AND2X1 U9387 ( .IN1(n8242), .IN2(n5433), .Q(WX2561) );
  XOR2X1 U9388 ( .IN1(CRC_OUT_8_1), .IN2(n4752), .Q(n8242) );
  AND2X1 U9389 ( .IN1(n8243), .IN2(n5434), .Q(WX2559) );
  XOR2X1 U9390 ( .IN1(CRC_OUT_8_0), .IN2(n4753), .Q(n8243) );
  AND2X1 U9391 ( .IN1(n8244), .IN2(n5433), .Q(WX2557) );
  XOR2X1 U9392 ( .IN1(n4541), .IN2(CRC_OUT_8_31), .Q(n8244) );
  AND2X1 U9393 ( .IN1(n5436), .IN2(n8653), .Q(WX2031) );
  AND2X1 U9394 ( .IN1(n5436), .IN2(n8654), .Q(WX2029) );
  AND2X1 U9395 ( .IN1(n5436), .IN2(n8655), .Q(WX2027) );
  AND2X1 U9396 ( .IN1(n5436), .IN2(n8656), .Q(WX2025) );
  AND2X1 U9397 ( .IN1(n5436), .IN2(n8657), .Q(WX2023) );
  AND2X1 U9398 ( .IN1(n5438), .IN2(n8658), .Q(WX2021) );
  AND2X1 U9399 ( .IN1(test_so13), .IN2(n5434), .Q(WX2019) );
  AND2X1 U9400 ( .IN1(n5437), .IN2(n8661), .Q(WX2017) );
  AND2X1 U9401 ( .IN1(n5437), .IN2(n8662), .Q(WX2015) );
  AND2X1 U9402 ( .IN1(n5437), .IN2(n8663), .Q(WX2013) );
  AND2X1 U9403 ( .IN1(n5437), .IN2(n8664), .Q(WX2011) );
  AND2X1 U9404 ( .IN1(n5437), .IN2(n8665), .Q(WX2009) );
  AND2X1 U9405 ( .IN1(n5437), .IN2(n8666), .Q(WX2007) );
  AND2X1 U9406 ( .IN1(n5437), .IN2(n8667), .Q(WX2005) );
  AND2X1 U9407 ( .IN1(n5437), .IN2(n8668), .Q(WX2003) );
  AND2X1 U9408 ( .IN1(n5438), .IN2(n8669), .Q(WX2001) );
  OR2X1 U9409 ( .IN1(n8245), .IN2(n8255), .Q(WX1999) );
  OR2X1 U9410 ( .IN1(n8256), .IN2(n8273), .Q(n8255) );
  AND2X1 U9411 ( .IN1(n4893), .IN2(CRC_OUT_8_0), .Q(n8273) );
  AND2X1 U9412 ( .IN1(n63), .IN2(n4866), .Q(n8256) );
  INVX0 U9413 ( .INP(n8274), .ZN(n63) );
  OR2X1 U9414 ( .IN1(n5478), .IN2(n4003), .Q(n8274) );
  OR2X1 U9415 ( .IN1(n8291), .IN2(n8292), .Q(n8245) );
  AND2X1 U9416 ( .IN1(n4928), .IN2(n7882), .Q(n8292) );
  XNOR2X1 U9417 ( .IN1(n8296), .IN2(n8297), .Q(n7882) );
  XOR2X1 U9418 ( .IN1(n9693), .IN2(n4540), .Q(n8297) );
  XOR2X1 U9419 ( .IN1(WX3293), .IN2(n4455), .Q(n8296) );
  AND2X1 U9420 ( .IN1(n6805), .IN2(n4837), .Q(n8291) );
  XOR2X1 U9421 ( .IN1(n8298), .IN2(n8299), .Q(n6805) );
  XOR2X1 U9422 ( .IN1(test_so16), .IN2(n9692), .Q(n8299) );
  XOR2X1 U9423 ( .IN1(WX2000), .IN2(n4541), .Q(n8298) );
  OR2X1 U9424 ( .IN1(n8300), .IN2(n8301), .Q(WX1997) );
  OR2X1 U9425 ( .IN1(n8302), .IN2(n8303), .Q(n8301) );
  AND2X1 U9426 ( .IN1(n4894), .IN2(CRC_OUT_8_1), .Q(n8303) );
  AND2X1 U9427 ( .IN1(n62), .IN2(n4866), .Q(n8302) );
  INVX0 U9428 ( .INP(n8308), .ZN(n62) );
  OR2X1 U9429 ( .IN1(n5478), .IN2(n4004), .Q(n8308) );
  OR2X1 U9430 ( .IN1(n8309), .IN2(n8326), .Q(n8300) );
  AND2X1 U9431 ( .IN1(n4928), .IN2(n7892), .Q(n8326) );
  XNOR2X1 U9432 ( .IN1(n8327), .IN2(n8344), .Q(n7892) );
  XOR2X1 U9433 ( .IN1(n9695), .IN2(n4727), .Q(n8344) );
  XOR2X1 U9434 ( .IN1(WX3291), .IN2(n4457), .Q(n8327) );
  AND2X1 U9435 ( .IN1(n4849), .IN2(n6813), .Q(n8309) );
  XNOR2X1 U9436 ( .IN1(n8345), .IN2(n8354), .Q(n6813) );
  XOR2X1 U9437 ( .IN1(n9694), .IN2(n4753), .Q(n8354) );
  XOR2X1 U9438 ( .IN1(WX1998), .IN2(n4486), .Q(n8345) );
  OR2X1 U9439 ( .IN1(n8355), .IN2(n8356), .Q(WX1995) );
  OR2X1 U9440 ( .IN1(n8357), .IN2(n8358), .Q(n8356) );
  AND2X1 U9441 ( .IN1(n4894), .IN2(CRC_OUT_8_2), .Q(n8358) );
  AND2X1 U9442 ( .IN1(n61), .IN2(n4865), .Q(n8357) );
  INVX0 U9443 ( .INP(n8359), .ZN(n61) );
  OR2X1 U9444 ( .IN1(n5478), .IN2(n4005), .Q(n8359) );
  OR2X1 U9445 ( .IN1(n8360), .IN2(n8361), .Q(n8355) );
  AND2X1 U9446 ( .IN1(n4928), .IN2(n7902), .Q(n8361) );
  XNOR2X1 U9447 ( .IN1(n8362), .IN2(n8379), .Q(n7902) );
  XOR2X1 U9448 ( .IN1(n9697), .IN2(n4726), .Q(n8379) );
  XOR2X1 U9449 ( .IN1(WX3289), .IN2(n4459), .Q(n8362) );
  AND2X1 U9450 ( .IN1(n4849), .IN2(n6821), .Q(n8360) );
  XNOR2X1 U9451 ( .IN1(n8380), .IN2(n8397), .Q(n6821) );
  XOR2X1 U9452 ( .IN1(n9696), .IN2(n4752), .Q(n8397) );
  XOR2X1 U9453 ( .IN1(WX1996), .IN2(n4488), .Q(n8380) );
  OR2X1 U9454 ( .IN1(n8398), .IN2(n8412), .Q(WX1993) );
  OR2X1 U9455 ( .IN1(n8413), .IN2(n8414), .Q(n8412) );
  AND2X1 U9456 ( .IN1(n4894), .IN2(CRC_OUT_8_3), .Q(n8414) );
  AND2X1 U9457 ( .IN1(n60), .IN2(n4865), .Q(n8413) );
  INVX0 U9458 ( .INP(n8415), .ZN(n60) );
  OR2X1 U9459 ( .IN1(n5478), .IN2(n4006), .Q(n8415) );
  OR2X1 U9460 ( .IN1(n8416), .IN2(n8417), .Q(n8398) );
  AND2X1 U9461 ( .IN1(n4928), .IN2(n7912), .Q(n8417) );
  XNOR2X1 U9462 ( .IN1(n8418), .IN2(n8419), .Q(n7912) );
  XOR2X1 U9463 ( .IN1(n9699), .IN2(n4725), .Q(n8419) );
  XOR2X1 U9464 ( .IN1(WX3287), .IN2(n4461), .Q(n8418) );
  AND2X1 U9465 ( .IN1(n4849), .IN2(n6829), .Q(n8416) );
  XNOR2X1 U9466 ( .IN1(n8420), .IN2(n8432), .Q(n6829) );
  XOR2X1 U9467 ( .IN1(n9698), .IN2(n4751), .Q(n8432) );
  XOR2X1 U9468 ( .IN1(WX1994), .IN2(n4490), .Q(n8420) );
  OR2X1 U9469 ( .IN1(n8433), .IN2(n8450), .Q(WX1991) );
  OR2X1 U9470 ( .IN1(n8451), .IN2(n8468), .Q(n8450) );
  AND2X1 U9471 ( .IN1(n4894), .IN2(CRC_OUT_8_4), .Q(n8468) );
  AND2X1 U9472 ( .IN1(n59), .IN2(n4865), .Q(n8451) );
  INVX0 U9473 ( .INP(n8469), .ZN(n59) );
  OR2X1 U9474 ( .IN1(n5478), .IN2(n4007), .Q(n8469) );
  OR2X1 U9475 ( .IN1(n8471), .IN2(n8472), .Q(n8433) );
  AND2X1 U9476 ( .IN1(n4928), .IN2(n7922), .Q(n8472) );
  XNOR2X1 U9477 ( .IN1(n8473), .IN2(n8474), .Q(n7922) );
  XOR2X1 U9478 ( .IN1(n9701), .IN2(n4530), .Q(n8474) );
  XOR2X1 U9479 ( .IN1(WX3285), .IN2(n4463), .Q(n8473) );
  AND2X1 U9480 ( .IN1(n6837), .IN2(n4837), .Q(n8471) );
  XOR2X1 U9481 ( .IN1(n8475), .IN2(n8476), .Q(n6837) );
  XOR2X1 U9482 ( .IN1(test_so14), .IN2(n9700), .Q(n8476) );
  XOR2X1 U9483 ( .IN1(WX2120), .IN2(n4533), .Q(n8475) );
  OR2X1 U9484 ( .IN1(n8477), .IN2(n8478), .Q(WX1989) );
  OR2X1 U9485 ( .IN1(n8485), .IN2(n8486), .Q(n8478) );
  AND2X1 U9486 ( .IN1(n4894), .IN2(CRC_OUT_8_5), .Q(n8486) );
  AND2X1 U9487 ( .IN1(n58), .IN2(n4865), .Q(n8485) );
  INVX0 U9488 ( .INP(n8503), .ZN(n58) );
  OR2X1 U9489 ( .IN1(n5478), .IN2(n4008), .Q(n8503) );
  OR2X1 U9490 ( .IN1(n8504), .IN2(n8521), .Q(n8477) );
  AND2X1 U9491 ( .IN1(n4928), .IN2(n7932), .Q(n8521) );
  XNOR2X1 U9492 ( .IN1(n8522), .IN2(n8529), .Q(n7932) );
  XOR2X1 U9493 ( .IN1(n9703), .IN2(n4724), .Q(n8529) );
  XOR2X1 U9494 ( .IN1(WX3283), .IN2(n4465), .Q(n8522) );
  AND2X1 U9495 ( .IN1(n4849), .IN2(n6845), .Q(n8504) );
  XNOR2X1 U9496 ( .IN1(n8530), .IN2(n8531), .Q(n6845) );
  XOR2X1 U9497 ( .IN1(n9702), .IN2(n4750), .Q(n8531) );
  XOR2X1 U9498 ( .IN1(WX1990), .IN2(n4493), .Q(n8530) );
  OR2X1 U9499 ( .IN1(n8532), .IN2(n8533), .Q(WX1987) );
  OR2X1 U9500 ( .IN1(n8534), .IN2(n8535), .Q(n8533) );
  AND2X1 U9501 ( .IN1(n4894), .IN2(CRC_OUT_8_6), .Q(n8535) );
  AND2X1 U9502 ( .IN1(n57), .IN2(n4865), .Q(n8534) );
  INVX0 U9503 ( .INP(n8536), .ZN(n57) );
  OR2X1 U9504 ( .IN1(n5478), .IN2(n4009), .Q(n8536) );
  OR2X1 U9505 ( .IN1(n8538), .IN2(n8539), .Q(n8532) );
  AND2X1 U9506 ( .IN1(n7942), .IN2(n4920), .Q(n8539) );
  XOR2X1 U9507 ( .IN1(n8556), .IN2(n8557), .Q(n7942) );
  XOR2X1 U9508 ( .IN1(test_so30), .IN2(n9705), .Q(n8557) );
  XOR2X1 U9509 ( .IN1(WX3281), .IN2(n4467), .Q(n8556) );
  AND2X1 U9510 ( .IN1(n4849), .IN2(n6853), .Q(n8538) );
  XNOR2X1 U9511 ( .IN1(n8574), .IN2(n8575), .Q(n6853) );
  XOR2X1 U9512 ( .IN1(n9704), .IN2(n4749), .Q(n8575) );
  XOR2X1 U9513 ( .IN1(WX1988), .IN2(n4495), .Q(n8574) );
  OR2X1 U9514 ( .IN1(n8587), .IN2(n8588), .Q(WX1985) );
  OR2X1 U9515 ( .IN1(n8589), .IN2(n8590), .Q(n8588) );
  AND2X1 U9516 ( .IN1(test_so20), .IN2(n4887), .Q(n8590) );
  AND2X1 U9517 ( .IN1(n56), .IN2(n4865), .Q(n8589) );
  INVX0 U9518 ( .INP(n8591), .ZN(n56) );
  OR2X1 U9519 ( .IN1(n5478), .IN2(n4010), .Q(n8591) );
  OR2X1 U9520 ( .IN1(n8592), .IN2(n8593), .Q(n8587) );
  AND2X1 U9521 ( .IN1(n4928), .IN2(n7952), .Q(n8593) );
  XNOR2X1 U9522 ( .IN1(n8594), .IN2(n8595), .Q(n7952) );
  XOR2X1 U9523 ( .IN1(n9707), .IN2(n4723), .Q(n8595) );
  XOR2X1 U9524 ( .IN1(WX3279), .IN2(n4469), .Q(n8594) );
  AND2X1 U9525 ( .IN1(n4849), .IN2(n6861), .Q(n8592) );
  XNOR2X1 U9526 ( .IN1(n8596), .IN2(n8614), .Q(n6861) );
  XOR2X1 U9527 ( .IN1(n9706), .IN2(n4748), .Q(n8614) );
  XOR2X1 U9528 ( .IN1(WX1986), .IN2(n4497), .Q(n8596) );
  OR2X1 U9529 ( .IN1(n8615), .IN2(n8633), .Q(WX1983) );
  OR2X1 U9530 ( .IN1(n8634), .IN2(n8645), .Q(n8633) );
  AND2X1 U9531 ( .IN1(n4894), .IN2(CRC_OUT_8_8), .Q(n8645) );
  AND2X1 U9532 ( .IN1(n55), .IN2(n4865), .Q(n8634) );
  INVX0 U9533 ( .INP(n8646), .ZN(n55) );
  OR2X1 U9534 ( .IN1(n5478), .IN2(n4011), .Q(n8646) );
  OR2X1 U9535 ( .IN1(n8647), .IN2(n8648), .Q(n8615) );
  AND2X1 U9536 ( .IN1(n7962), .IN2(n4920), .Q(n8648) );
  XOR2X1 U9537 ( .IN1(n8649), .IN2(n8650), .Q(n7962) );
  XOR2X1 U9538 ( .IN1(test_so28), .IN2(n9709), .Q(n8650) );
  XOR2X1 U9539 ( .IN1(WX3277), .IN2(n4722), .Q(n8649) );
  AND2X1 U9540 ( .IN1(n4849), .IN2(n6869), .Q(n8647) );
  XNOR2X1 U9541 ( .IN1(n8651), .IN2(n8652), .Q(n6869) );
  XOR2X1 U9542 ( .IN1(n9708), .IN2(n4747), .Q(n8652) );
  XOR2X1 U9543 ( .IN1(WX1984), .IN2(n4499), .Q(n8651) );
  OR2X1 U9544 ( .IN1(n8659), .IN2(n8660), .Q(WX1981) );
  OR2X1 U9545 ( .IN1(n8678), .IN2(n8679), .Q(n8660) );
  AND2X1 U9546 ( .IN1(n4894), .IN2(CRC_OUT_8_9), .Q(n8679) );
  AND2X1 U9547 ( .IN1(n54), .IN2(n4865), .Q(n8678) );
  INVX0 U9548 ( .INP(n8697), .ZN(n54) );
  OR2X1 U9549 ( .IN1(n5477), .IN2(n4012), .Q(n8697) );
  OR2X1 U9550 ( .IN1(n8698), .IN2(n8703), .Q(n8659) );
  AND2X1 U9551 ( .IN1(n4928), .IN2(n7972), .Q(n8703) );
  XNOR2X1 U9552 ( .IN1(n8704), .IN2(n8705), .Q(n7972) );
  XOR2X1 U9553 ( .IN1(n9711), .IN2(n4721), .Q(n8705) );
  XOR2X1 U9554 ( .IN1(WX3275), .IN2(n4472), .Q(n8704) );
  AND2X1 U9555 ( .IN1(n4848), .IN2(n6877), .Q(n8698) );
  XNOR2X1 U9556 ( .IN1(n8706), .IN2(n8707), .Q(n6877) );
  XOR2X1 U9557 ( .IN1(n9710), .IN2(n4746), .Q(n8707) );
  XOR2X1 U9558 ( .IN1(WX1982), .IN2(n4501), .Q(n8706) );
  OR2X1 U9559 ( .IN1(n8708), .IN2(n8709), .Q(WX1979) );
  OR2X1 U9560 ( .IN1(n8710), .IN2(n8711), .Q(n8709) );
  AND2X1 U9561 ( .IN1(n4894), .IN2(CRC_OUT_8_10), .Q(n8711) );
  AND2X1 U9562 ( .IN1(n53), .IN2(n4865), .Q(n8710) );
  INVX0 U9563 ( .INP(n8712), .ZN(n53) );
  OR2X1 U9564 ( .IN1(n5477), .IN2(n4013), .Q(n8712) );
  OR2X1 U9565 ( .IN1(n8713), .IN2(n8714), .Q(n8708) );
  AND2X1 U9566 ( .IN1(n4928), .IN2(n7982), .Q(n8714) );
  XNOR2X1 U9567 ( .IN1(n8715), .IN2(n8716), .Q(n7982) );
  XOR2X1 U9568 ( .IN1(n9713), .IN2(n4720), .Q(n8716) );
  XOR2X1 U9569 ( .IN1(WX3273), .IN2(n4474), .Q(n8715) );
  AND2X1 U9570 ( .IN1(n6885), .IN2(n4836), .Q(n8713) );
  XOR2X1 U9571 ( .IN1(n8717), .IN2(n8718), .Q(n6885) );
  XOR2X1 U9572 ( .IN1(test_so19), .IN2(n9712), .Q(n8718) );
  XOR2X1 U9573 ( .IN1(WX1980), .IN2(n4503), .Q(n8717) );
  OR2X1 U9574 ( .IN1(n8719), .IN2(n8720), .Q(WX1977) );
  OR2X1 U9575 ( .IN1(n8721), .IN2(n8722), .Q(n8720) );
  AND2X1 U9576 ( .IN1(n4894), .IN2(CRC_OUT_8_11), .Q(n8722) );
  AND2X1 U9577 ( .IN1(n52), .IN2(n4865), .Q(n8721) );
  INVX0 U9578 ( .INP(n8723), .ZN(n52) );
  OR2X1 U9579 ( .IN1(n5477), .IN2(n4014), .Q(n8723) );
  OR2X1 U9580 ( .IN1(n8724), .IN2(n8725), .Q(n8719) );
  AND2X1 U9581 ( .IN1(n4928), .IN2(n7992), .Q(n8725) );
  XNOR2X1 U9582 ( .IN1(n8726), .IN2(n8727), .Q(n7992) );
  XOR2X1 U9583 ( .IN1(n9715), .IN2(n4529), .Q(n8727) );
  XOR2X1 U9584 ( .IN1(WX3271), .IN2(n4476), .Q(n8726) );
  AND2X1 U9585 ( .IN1(n4848), .IN2(n6893), .Q(n8724) );
  XNOR2X1 U9586 ( .IN1(n8728), .IN2(n8729), .Q(n6893) );
  XOR2X1 U9587 ( .IN1(n9714), .IN2(n4532), .Q(n8729) );
  XOR2X1 U9588 ( .IN1(WX1978), .IN2(n4505), .Q(n8728) );
  OR2X1 U9589 ( .IN1(n8730), .IN2(n8731), .Q(WX1975) );
  OR2X1 U9590 ( .IN1(n8732), .IN2(n8733), .Q(n8731) );
  AND2X1 U9591 ( .IN1(n4894), .IN2(CRC_OUT_8_12), .Q(n8733) );
  AND2X1 U9592 ( .IN1(n51), .IN2(n4865), .Q(n8732) );
  INVX0 U9593 ( .INP(n8734), .ZN(n51) );
  OR2X1 U9594 ( .IN1(n5477), .IN2(n4015), .Q(n8734) );
  OR2X1 U9595 ( .IN1(n8735), .IN2(n8736), .Q(n8730) );
  AND2X1 U9596 ( .IN1(n8002), .IN2(n4920), .Q(n8736) );
  XOR2X1 U9597 ( .IN1(n8737), .IN2(n8738), .Q(n8002) );
  XOR2X1 U9598 ( .IN1(test_so26), .IN2(n9717), .Q(n8738) );
  XOR2X1 U9599 ( .IN1(WX3269), .IN2(n4719), .Q(n8737) );
  AND2X1 U9600 ( .IN1(n4848), .IN2(n6901), .Q(n8735) );
  XNOR2X1 U9601 ( .IN1(n8739), .IN2(n8740), .Q(n6901) );
  XOR2X1 U9602 ( .IN1(n9716), .IN2(n4745), .Q(n8740) );
  XOR2X1 U9603 ( .IN1(WX1976), .IN2(n4507), .Q(n8739) );
  OR2X1 U9604 ( .IN1(n8741), .IN2(n8742), .Q(WX1973) );
  OR2X1 U9605 ( .IN1(n8743), .IN2(n8744), .Q(n8742) );
  AND2X1 U9606 ( .IN1(n4894), .IN2(CRC_OUT_8_13), .Q(n8744) );
  AND2X1 U9607 ( .IN1(n50), .IN2(n4865), .Q(n8743) );
  INVX0 U9608 ( .INP(n8745), .ZN(n50) );
  OR2X1 U9609 ( .IN1(n5477), .IN2(n4016), .Q(n8745) );
  OR2X1 U9610 ( .IN1(n8746), .IN2(n8747), .Q(n8741) );
  AND2X1 U9611 ( .IN1(n4929), .IN2(n8012), .Q(n8747) );
  XNOR2X1 U9612 ( .IN1(n8748), .IN2(n8749), .Q(n8012) );
  XOR2X1 U9613 ( .IN1(n9719), .IN2(n4718), .Q(n8749) );
  XOR2X1 U9614 ( .IN1(WX3267), .IN2(n4479), .Q(n8748) );
  AND2X1 U9615 ( .IN1(n4848), .IN2(n6909), .Q(n8746) );
  XNOR2X1 U9616 ( .IN1(n8750), .IN2(n8751), .Q(n6909) );
  XOR2X1 U9617 ( .IN1(n9718), .IN2(n4744), .Q(n8751) );
  XOR2X1 U9618 ( .IN1(WX1974), .IN2(n4509), .Q(n8750) );
  OR2X1 U9619 ( .IN1(n8752), .IN2(n8753), .Q(WX1971) );
  OR2X1 U9620 ( .IN1(n8754), .IN2(n8755), .Q(n8753) );
  AND2X1 U9621 ( .IN1(n4894), .IN2(CRC_OUT_8_14), .Q(n8755) );
  AND2X1 U9622 ( .IN1(n49), .IN2(n4864), .Q(n8754) );
  INVX0 U9623 ( .INP(n8756), .ZN(n49) );
  OR2X1 U9624 ( .IN1(n5477), .IN2(n4017), .Q(n8756) );
  OR2X1 U9625 ( .IN1(n8757), .IN2(n8758), .Q(n8752) );
  AND2X1 U9626 ( .IN1(n4929), .IN2(n8022), .Q(n8758) );
  XNOR2X1 U9627 ( .IN1(n8759), .IN2(n8760), .Q(n8022) );
  XOR2X1 U9628 ( .IN1(n9721), .IN2(n4717), .Q(n8760) );
  XOR2X1 U9629 ( .IN1(WX3265), .IN2(n4481), .Q(n8759) );
  AND2X1 U9630 ( .IN1(n6917), .IN2(n4835), .Q(n8757) );
  XOR2X1 U9631 ( .IN1(n8761), .IN2(n8762), .Q(n6917) );
  XOR2X1 U9632 ( .IN1(test_so17), .IN2(n9720), .Q(n8762) );
  XOR2X1 U9633 ( .IN1(WX1972), .IN2(n4743), .Q(n8761) );
  OR2X1 U9634 ( .IN1(n8763), .IN2(n8764), .Q(WX1969) );
  OR2X1 U9635 ( .IN1(n8765), .IN2(n8766), .Q(n8764) );
  AND2X1 U9636 ( .IN1(n4895), .IN2(CRC_OUT_8_15), .Q(n8766) );
  AND2X1 U9637 ( .IN1(n48), .IN2(n4864), .Q(n8765) );
  INVX0 U9638 ( .INP(n8767), .ZN(n48) );
  OR2X1 U9639 ( .IN1(n5477), .IN2(n4018), .Q(n8767) );
  OR2X1 U9640 ( .IN1(n8768), .IN2(n8769), .Q(n8763) );
  AND2X1 U9641 ( .IN1(n4929), .IN2(n8032), .Q(n8769) );
  XNOR2X1 U9642 ( .IN1(n8770), .IN2(n8771), .Q(n8032) );
  XOR2X1 U9643 ( .IN1(n9723), .IN2(n4716), .Q(n8771) );
  XOR2X1 U9644 ( .IN1(WX3263), .IN2(n4483), .Q(n8770) );
  AND2X1 U9645 ( .IN1(n4848), .IN2(n6925), .Q(n8768) );
  XNOR2X1 U9646 ( .IN1(n8772), .IN2(n8773), .Q(n6925) );
  XOR2X1 U9647 ( .IN1(n9722), .IN2(n4742), .Q(n8773) );
  XOR2X1 U9648 ( .IN1(WX1970), .IN2(n4512), .Q(n8772) );
  OR2X1 U9649 ( .IN1(n8774), .IN2(n8775), .Q(WX1967) );
  OR2X1 U9650 ( .IN1(n8776), .IN2(n8777), .Q(n8775) );
  AND2X1 U9651 ( .IN1(n4895), .IN2(CRC_OUT_8_16), .Q(n8777) );
  AND2X1 U9652 ( .IN1(n47), .IN2(n4864), .Q(n8776) );
  INVX0 U9653 ( .INP(n8778), .ZN(n47) );
  OR2X1 U9654 ( .IN1(n5477), .IN2(n4019), .Q(n8778) );
  OR2X1 U9655 ( .IN1(n8779), .IN2(n8780), .Q(n8774) );
  AND2X1 U9656 ( .IN1(n8042), .IN2(n4920), .Q(n8780) );
  XOR2X1 U9657 ( .IN1(n8781), .IN2(n8782), .Q(n8042) );
  XOR2X1 U9658 ( .IN1(n4252), .IN2(n5383), .Q(n8782) );
  XOR2X1 U9659 ( .IN1(n8783), .IN2(n4528), .Q(n8781) );
  XOR2X1 U9660 ( .IN1(WX3325), .IN2(test_so24), .Q(n8783) );
  AND2X1 U9661 ( .IN1(n4848), .IN2(n6933), .Q(n8779) );
  XNOR2X1 U9662 ( .IN1(n8784), .IN2(n8785), .Q(n6933) );
  XOR2X1 U9663 ( .IN1(n4265), .IN2(n5383), .Q(n8785) );
  XOR2X1 U9664 ( .IN1(n8786), .IN2(n4531), .Q(n8784) );
  XNOR2X1 U9665 ( .IN1(WX2096), .IN2(n8653), .Q(n8786) );
  OR2X1 U9666 ( .IN1(n8787), .IN2(n8788), .Q(WX1965) );
  OR2X1 U9667 ( .IN1(n8789), .IN2(n8790), .Q(n8788) );
  AND2X1 U9668 ( .IN1(n4895), .IN2(CRC_OUT_8_17), .Q(n8790) );
  AND2X1 U9669 ( .IN1(n46), .IN2(n4864), .Q(n8789) );
  INVX0 U9670 ( .INP(n8791), .ZN(n46) );
  OR2X1 U9671 ( .IN1(n5477), .IN2(n4020), .Q(n8791) );
  OR2X1 U9672 ( .IN1(n8792), .IN2(n8793), .Q(n8787) );
  AND2X1 U9673 ( .IN1(n4929), .IN2(n8053), .Q(n8793) );
  XNOR2X1 U9674 ( .IN1(n8794), .IN2(n8795), .Q(n8053) );
  XOR2X1 U9675 ( .IN1(n4253), .IN2(n5383), .Q(n8795) );
  XOR2X1 U9676 ( .IN1(n8796), .IN2(n4715), .Q(n8794) );
  XOR2X1 U9677 ( .IN1(WX3387), .IN2(n9724), .Q(n8796) );
  AND2X1 U9678 ( .IN1(n4848), .IN2(n6941), .Q(n8792) );
  XNOR2X1 U9679 ( .IN1(n8797), .IN2(n8798), .Q(n6941) );
  XOR2X1 U9680 ( .IN1(n4266), .IN2(n5383), .Q(n8798) );
  XOR2X1 U9681 ( .IN1(n8799), .IN2(n4741), .Q(n8797) );
  XNOR2X1 U9682 ( .IN1(WX2094), .IN2(n8654), .Q(n8799) );
  OR2X1 U9683 ( .IN1(n8800), .IN2(n8801), .Q(WX1963) );
  OR2X1 U9684 ( .IN1(n8802), .IN2(n8803), .Q(n8801) );
  AND2X1 U9685 ( .IN1(n4895), .IN2(CRC_OUT_8_18), .Q(n8803) );
  AND2X1 U9686 ( .IN1(n45), .IN2(n4864), .Q(n8802) );
  INVX0 U9687 ( .INP(n8804), .ZN(n45) );
  OR2X1 U9688 ( .IN1(n5477), .IN2(n4021), .Q(n8804) );
  OR2X1 U9689 ( .IN1(n8805), .IN2(n8806), .Q(n8800) );
  AND2X1 U9690 ( .IN1(n4929), .IN2(n8064), .Q(n8806) );
  XNOR2X1 U9691 ( .IN1(n8807), .IN2(n8808), .Q(n8064) );
  XOR2X1 U9692 ( .IN1(n4254), .IN2(n5382), .Q(n8808) );
  XOR2X1 U9693 ( .IN1(n8809), .IN2(n4714), .Q(n8807) );
  XOR2X1 U9694 ( .IN1(WX3385), .IN2(n9727), .Q(n8809) );
  AND2X1 U9695 ( .IN1(n6949), .IN2(n4836), .Q(n8805) );
  XOR2X1 U9696 ( .IN1(n8810), .IN2(n8811), .Q(n6949) );
  XOR2X1 U9697 ( .IN1(n4740), .IN2(n5382), .Q(n8811) );
  XOR2X1 U9698 ( .IN1(n8812), .IN2(n9726), .Q(n8810) );
  XNOR2X1 U9699 ( .IN1(n9725), .IN2(n8655), .Q(n8812) );
  OR2X1 U9700 ( .IN1(n8813), .IN2(n8814), .Q(WX1961) );
  OR2X1 U9701 ( .IN1(n8815), .IN2(n8816), .Q(n8814) );
  AND2X1 U9702 ( .IN1(n4895), .IN2(CRC_OUT_8_19), .Q(n8816) );
  AND2X1 U9703 ( .IN1(n44), .IN2(n4864), .Q(n8815) );
  INVX0 U9704 ( .INP(n8817), .ZN(n44) );
  OR2X1 U9705 ( .IN1(n5477), .IN2(n4022), .Q(n8817) );
  OR2X1 U9706 ( .IN1(n8818), .IN2(n8819), .Q(n8813) );
  AND2X1 U9707 ( .IN1(n4929), .IN2(n8075), .Q(n8819) );
  XNOR2X1 U9708 ( .IN1(n8820), .IN2(n8821), .Q(n8075) );
  XOR2X1 U9709 ( .IN1(n4255), .IN2(n5382), .Q(n8821) );
  XOR2X1 U9710 ( .IN1(n8822), .IN2(n4713), .Q(n8820) );
  XOR2X1 U9711 ( .IN1(WX3383), .IN2(n9728), .Q(n8822) );
  AND2X1 U9712 ( .IN1(n4848), .IN2(n6957), .Q(n8818) );
  XNOR2X1 U9713 ( .IN1(n8823), .IN2(n8824), .Q(n6957) );
  XOR2X1 U9714 ( .IN1(n4267), .IN2(n5382), .Q(n8824) );
  XOR2X1 U9715 ( .IN1(n8825), .IN2(n4739), .Q(n8823) );
  XNOR2X1 U9716 ( .IN1(WX2090), .IN2(n8656), .Q(n8825) );
  OR2X1 U9717 ( .IN1(n8826), .IN2(n8827), .Q(WX1959) );
  OR2X1 U9718 ( .IN1(n8828), .IN2(n8829), .Q(n8827) );
  AND2X1 U9719 ( .IN1(n4895), .IN2(CRC_OUT_8_20), .Q(n8829) );
  AND2X1 U9720 ( .IN1(n43), .IN2(n4864), .Q(n8828) );
  INVX0 U9721 ( .INP(n8830), .ZN(n43) );
  OR2X1 U9722 ( .IN1(n5477), .IN2(n4023), .Q(n8830) );
  OR2X1 U9723 ( .IN1(n8831), .IN2(n8832), .Q(n8826) );
  AND2X1 U9724 ( .IN1(n4929), .IN2(n8086), .Q(n8832) );
  XNOR2X1 U9725 ( .IN1(n8833), .IN2(n8834), .Q(n8086) );
  XOR2X1 U9726 ( .IN1(n4256), .IN2(n5382), .Q(n8834) );
  XOR2X1 U9727 ( .IN1(n8835), .IN2(n4712), .Q(n8833) );
  XOR2X1 U9728 ( .IN1(WX3381), .IN2(n9729), .Q(n8835) );
  AND2X1 U9729 ( .IN1(n4848), .IN2(n6965), .Q(n8831) );
  XNOR2X1 U9730 ( .IN1(n8836), .IN2(n8837), .Q(n6965) );
  XOR2X1 U9731 ( .IN1(n4268), .IN2(n5382), .Q(n8837) );
  XOR2X1 U9732 ( .IN1(n8838), .IN2(n4738), .Q(n8836) );
  XNOR2X1 U9733 ( .IN1(WX2088), .IN2(n8657), .Q(n8838) );
  OR2X1 U9734 ( .IN1(n8839), .IN2(n8840), .Q(WX1957) );
  OR2X1 U9735 ( .IN1(n8841), .IN2(n8842), .Q(n8840) );
  AND2X1 U9736 ( .IN1(n4895), .IN2(CRC_OUT_8_21), .Q(n8842) );
  AND2X1 U9737 ( .IN1(n42), .IN2(n4864), .Q(n8841) );
  INVX0 U9738 ( .INP(n8843), .ZN(n42) );
  OR2X1 U9739 ( .IN1(n5477), .IN2(n4024), .Q(n8843) );
  OR2X1 U9740 ( .IN1(n8844), .IN2(n8845), .Q(n8839) );
  AND2X1 U9741 ( .IN1(n4929), .IN2(n8097), .Q(n8845) );
  XNOR2X1 U9742 ( .IN1(n8846), .IN2(n8847), .Q(n8097) );
  XOR2X1 U9743 ( .IN1(n4257), .IN2(n5382), .Q(n8847) );
  XOR2X1 U9744 ( .IN1(n8848), .IN2(n4711), .Q(n8846) );
  XOR2X1 U9745 ( .IN1(WX3379), .IN2(n9730), .Q(n8848) );
  AND2X1 U9746 ( .IN1(n4848), .IN2(n6973), .Q(n8844) );
  XNOR2X1 U9747 ( .IN1(n8849), .IN2(n8850), .Q(n6973) );
  XOR2X1 U9748 ( .IN1(n4269), .IN2(n5382), .Q(n8850) );
  XOR2X1 U9749 ( .IN1(n8851), .IN2(n4737), .Q(n8849) );
  XNOR2X1 U9750 ( .IN1(WX2086), .IN2(n8658), .Q(n8851) );
  OR2X1 U9751 ( .IN1(n8852), .IN2(n8853), .Q(WX1955) );
  OR2X1 U9752 ( .IN1(n8854), .IN2(n8855), .Q(n8853) );
  AND2X1 U9753 ( .IN1(n4895), .IN2(CRC_OUT_8_22), .Q(n8855) );
  AND2X1 U9754 ( .IN1(n41), .IN2(n4864), .Q(n8854) );
  INVX0 U9755 ( .INP(n8856), .ZN(n41) );
  OR2X1 U9756 ( .IN1(n5476), .IN2(n4025), .Q(n8856) );
  OR2X1 U9757 ( .IN1(n8857), .IN2(n8858), .Q(n8852) );
  AND2X1 U9758 ( .IN1(n4929), .IN2(n8108), .Q(n8858) );
  XNOR2X1 U9759 ( .IN1(n8859), .IN2(n8860), .Q(n8108) );
  XOR2X1 U9760 ( .IN1(n4258), .IN2(n5382), .Q(n8860) );
  XOR2X1 U9761 ( .IN1(n8861), .IN2(n4710), .Q(n8859) );
  XOR2X1 U9762 ( .IN1(WX3377), .IN2(n9731), .Q(n8861) );
  AND2X1 U9763 ( .IN1(n6981), .IN2(n4835), .Q(n8857) );
  XOR2X1 U9764 ( .IN1(n8862), .IN2(n8863), .Q(n6981) );
  XOR2X1 U9765 ( .IN1(n4270), .IN2(n5382), .Q(n8863) );
  XOR2X1 U9766 ( .IN1(n8864), .IN2(n4736), .Q(n8862) );
  XOR2X1 U9767 ( .IN1(WX2020), .IN2(test_so13), .Q(n8864) );
  OR2X1 U9768 ( .IN1(n8865), .IN2(n8866), .Q(WX1953) );
  OR2X1 U9769 ( .IN1(n8867), .IN2(n8868), .Q(n8866) );
  AND2X1 U9770 ( .IN1(n4895), .IN2(CRC_OUT_8_23), .Q(n8868) );
  AND2X1 U9771 ( .IN1(n40), .IN2(n4864), .Q(n8867) );
  INVX0 U9772 ( .INP(n8869), .ZN(n40) );
  OR2X1 U9773 ( .IN1(n5476), .IN2(n4026), .Q(n8869) );
  OR2X1 U9774 ( .IN1(n8870), .IN2(n8871), .Q(n8865) );
  AND2X1 U9775 ( .IN1(n8119), .IN2(n4920), .Q(n8871) );
  XOR2X1 U9776 ( .IN1(n8872), .IN2(n8873), .Q(n8119) );
  XOR2X1 U9777 ( .IN1(n4259), .IN2(n5382), .Q(n8873) );
  XOR2X1 U9778 ( .IN1(WX3311), .IN2(n8874), .Q(n8872) );
  XOR2X1 U9779 ( .IN1(test_so29), .IN2(n9732), .Q(n8874) );
  AND2X1 U9780 ( .IN1(n4848), .IN2(n6989), .Q(n8870) );
  XNOR2X1 U9781 ( .IN1(n8875), .IN2(n8876), .Q(n6989) );
  XOR2X1 U9782 ( .IN1(n4271), .IN2(n5382), .Q(n8876) );
  XOR2X1 U9783 ( .IN1(n8877), .IN2(n4735), .Q(n8875) );
  XNOR2X1 U9784 ( .IN1(WX2082), .IN2(n8661), .Q(n8877) );
  OR2X1 U9785 ( .IN1(n8878), .IN2(n8879), .Q(WX1951) );
  OR2X1 U9786 ( .IN1(n8880), .IN2(n8881), .Q(n8879) );
  AND2X1 U9787 ( .IN1(n4895), .IN2(CRC_OUT_8_24), .Q(n8881) );
  AND2X1 U9788 ( .IN1(n39), .IN2(n4864), .Q(n8880) );
  INVX0 U9789 ( .INP(n8882), .ZN(n39) );
  OR2X1 U9790 ( .IN1(n5476), .IN2(n4027), .Q(n8882) );
  OR2X1 U9791 ( .IN1(n8883), .IN2(n8884), .Q(n8878) );
  AND2X1 U9792 ( .IN1(n4929), .IN2(n8130), .Q(n8884) );
  XNOR2X1 U9793 ( .IN1(n8885), .IN2(n8886), .Q(n8130) );
  XOR2X1 U9794 ( .IN1(n4260), .IN2(n5381), .Q(n8886) );
  XOR2X1 U9795 ( .IN1(n8887), .IN2(n4709), .Q(n8885) );
  XOR2X1 U9796 ( .IN1(WX3373), .IN2(n9733), .Q(n8887) );
  AND2X1 U9797 ( .IN1(n4848), .IN2(n6997), .Q(n8883) );
  XNOR2X1 U9798 ( .IN1(n8888), .IN2(n8889), .Q(n6997) );
  XOR2X1 U9799 ( .IN1(n4272), .IN2(n5381), .Q(n8889) );
  XOR2X1 U9800 ( .IN1(n8890), .IN2(n4734), .Q(n8888) );
  XNOR2X1 U9801 ( .IN1(WX2080), .IN2(n8662), .Q(n8890) );
  OR2X1 U9802 ( .IN1(n8891), .IN2(n8892), .Q(WX1949) );
  OR2X1 U9803 ( .IN1(n8893), .IN2(n8894), .Q(n8892) );
  AND2X1 U9804 ( .IN1(test_so21), .IN2(n4888), .Q(n8894) );
  AND2X1 U9805 ( .IN1(n38), .IN2(n4864), .Q(n8893) );
  INVX0 U9806 ( .INP(n8895), .ZN(n38) );
  OR2X1 U9807 ( .IN1(n5476), .IN2(n4028), .Q(n8895) );
  OR2X1 U9808 ( .IN1(n8896), .IN2(n8897), .Q(n8891) );
  AND2X1 U9809 ( .IN1(n4929), .IN2(n8141), .Q(n8897) );
  XNOR2X1 U9810 ( .IN1(n8898), .IN2(n8899), .Q(n8141) );
  XOR2X1 U9811 ( .IN1(n4261), .IN2(n5381), .Q(n8899) );
  XOR2X1 U9812 ( .IN1(n8900), .IN2(n4708), .Q(n8898) );
  XOR2X1 U9813 ( .IN1(WX3371), .IN2(n9734), .Q(n8900) );
  AND2X1 U9814 ( .IN1(n4848), .IN2(n7005), .Q(n8896) );
  XNOR2X1 U9815 ( .IN1(n8901), .IN2(n8902), .Q(n7005) );
  XOR2X1 U9816 ( .IN1(n4273), .IN2(n5381), .Q(n8902) );
  XOR2X1 U9817 ( .IN1(n8903), .IN2(n4733), .Q(n8901) );
  XNOR2X1 U9818 ( .IN1(WX2078), .IN2(n8663), .Q(n8903) );
  OR2X1 U9819 ( .IN1(n8904), .IN2(n8905), .Q(WX1947) );
  OR2X1 U9820 ( .IN1(n8906), .IN2(n8907), .Q(n8905) );
  AND2X1 U9821 ( .IN1(n4895), .IN2(CRC_OUT_8_26), .Q(n8907) );
  AND2X1 U9822 ( .IN1(n37), .IN2(n4863), .Q(n8906) );
  INVX0 U9823 ( .INP(n8908), .ZN(n37) );
  OR2X1 U9824 ( .IN1(n5476), .IN2(n4029), .Q(n8908) );
  OR2X1 U9825 ( .IN1(n8909), .IN2(n8910), .Q(n8904) );
  AND2X1 U9826 ( .IN1(n8152), .IN2(n4920), .Q(n8910) );
  XOR2X1 U9827 ( .IN1(n8911), .IN2(n8912), .Q(n8152) );
  XOR2X1 U9828 ( .IN1(n4707), .IN2(n5381), .Q(n8912) );
  XOR2X1 U9829 ( .IN1(n8913), .IN2(n9737), .Q(n8911) );
  XOR2X1 U9830 ( .IN1(n9736), .IN2(n9735), .Q(n8913) );
  AND2X1 U9831 ( .IN1(n4847), .IN2(n7013), .Q(n8909) );
  XNOR2X1 U9832 ( .IN1(n8914), .IN2(n8915), .Q(n7013) );
  XOR2X1 U9833 ( .IN1(n4274), .IN2(n5381), .Q(n8915) );
  XOR2X1 U9834 ( .IN1(n8916), .IN2(n4732), .Q(n8914) );
  XNOR2X1 U9835 ( .IN1(WX2076), .IN2(n8664), .Q(n8916) );
  OR2X1 U9836 ( .IN1(n8917), .IN2(n8918), .Q(WX1945) );
  OR2X1 U9837 ( .IN1(n8919), .IN2(n8920), .Q(n8918) );
  AND2X1 U9838 ( .IN1(n4895), .IN2(CRC_OUT_8_27), .Q(n8920) );
  AND2X1 U9839 ( .IN1(n36), .IN2(n4863), .Q(n8919) );
  INVX0 U9840 ( .INP(n8921), .ZN(n36) );
  OR2X1 U9841 ( .IN1(n5476), .IN2(n4030), .Q(n8921) );
  OR2X1 U9842 ( .IN1(n8922), .IN2(n8923), .Q(n8917) );
  AND2X1 U9843 ( .IN1(n4925), .IN2(n8163), .Q(n8923) );
  XNOR2X1 U9844 ( .IN1(n8924), .IN2(n8925), .Q(n8163) );
  XOR2X1 U9845 ( .IN1(n4262), .IN2(n5381), .Q(n8925) );
  XOR2X1 U9846 ( .IN1(n8926), .IN2(n4706), .Q(n8924) );
  XOR2X1 U9847 ( .IN1(WX3367), .IN2(n9738), .Q(n8926) );
  AND2X1 U9848 ( .IN1(n4847), .IN2(n7021), .Q(n8922) );
  XNOR2X1 U9849 ( .IN1(n8927), .IN2(n8928), .Q(n7021) );
  XOR2X1 U9850 ( .IN1(n4275), .IN2(n5381), .Q(n8928) );
  XOR2X1 U9851 ( .IN1(n8929), .IN2(n4731), .Q(n8927) );
  XNOR2X1 U9852 ( .IN1(WX2074), .IN2(n8665), .Q(n8929) );
  OR2X1 U9853 ( .IN1(n8930), .IN2(n8931), .Q(WX1943) );
  OR2X1 U9854 ( .IN1(n8932), .IN2(n8933), .Q(n8931) );
  AND2X1 U9855 ( .IN1(n4895), .IN2(CRC_OUT_8_28), .Q(n8933) );
  AND2X1 U9856 ( .IN1(n35), .IN2(n4863), .Q(n8932) );
  INVX0 U9857 ( .INP(n8934), .ZN(n35) );
  OR2X1 U9858 ( .IN1(n5476), .IN2(n4031), .Q(n8934) );
  OR2X1 U9859 ( .IN1(n8935), .IN2(n8936), .Q(n8930) );
  AND2X1 U9860 ( .IN1(n4930), .IN2(n8174), .Q(n8936) );
  XNOR2X1 U9861 ( .IN1(n8937), .IN2(n8938), .Q(n8174) );
  XOR2X1 U9862 ( .IN1(n4263), .IN2(n5381), .Q(n8938) );
  XOR2X1 U9863 ( .IN1(n8939), .IN2(n4705), .Q(n8937) );
  XOR2X1 U9864 ( .IN1(WX3365), .IN2(n9739), .Q(n8939) );
  AND2X1 U9865 ( .IN1(n7029), .IN2(n4835), .Q(n8935) );
  XOR2X1 U9866 ( .IN1(n8940), .IN2(n8941), .Q(n7029) );
  XOR2X1 U9867 ( .IN1(n4276), .IN2(n5381), .Q(n8941) );
  XOR2X1 U9868 ( .IN1(WX2008), .IN2(n8942), .Q(n8940) );
  XNOR2X1 U9869 ( .IN1(test_so18), .IN2(n8666), .Q(n8942) );
  OR2X1 U9870 ( .IN1(n8943), .IN2(n8944), .Q(WX1941) );
  OR2X1 U9871 ( .IN1(n8945), .IN2(n8946), .Q(n8944) );
  AND2X1 U9872 ( .IN1(n4896), .IN2(CRC_OUT_8_29), .Q(n8946) );
  AND2X1 U9873 ( .IN1(n34), .IN2(n4863), .Q(n8945) );
  INVX0 U9874 ( .INP(n8947), .ZN(n34) );
  OR2X1 U9875 ( .IN1(n5476), .IN2(n4032), .Q(n8947) );
  OR2X1 U9876 ( .IN1(n8948), .IN2(n8949), .Q(n8943) );
  AND2X1 U9877 ( .IN1(n4929), .IN2(n8185), .Q(n8949) );
  XNOR2X1 U9878 ( .IN1(n8950), .IN2(n8951), .Q(n8185) );
  XOR2X1 U9879 ( .IN1(n4264), .IN2(n5381), .Q(n8951) );
  XOR2X1 U9880 ( .IN1(n8952), .IN2(n4704), .Q(n8950) );
  XOR2X1 U9881 ( .IN1(WX3363), .IN2(n9740), .Q(n8952) );
  AND2X1 U9882 ( .IN1(n4847), .IN2(n7048), .Q(n8948) );
  XNOR2X1 U9883 ( .IN1(n8953), .IN2(n8954), .Q(n7048) );
  XOR2X1 U9884 ( .IN1(n4277), .IN2(n5381), .Q(n8954) );
  XOR2X1 U9885 ( .IN1(n8955), .IN2(n4730), .Q(n8953) );
  XNOR2X1 U9886 ( .IN1(WX2070), .IN2(n8667), .Q(n8955) );
  OR2X1 U9887 ( .IN1(n8956), .IN2(n8957), .Q(WX1939) );
  OR2X1 U9888 ( .IN1(n8958), .IN2(n8959), .Q(n8957) );
  AND2X1 U9889 ( .IN1(n4896), .IN2(CRC_OUT_8_30), .Q(n8959) );
  AND2X1 U9890 ( .IN1(n33), .IN2(n4863), .Q(n8958) );
  INVX0 U9891 ( .INP(n8960), .ZN(n33) );
  OR2X1 U9892 ( .IN1(n5476), .IN2(n4033), .Q(n8960) );
  OR2X1 U9893 ( .IN1(n8961), .IN2(n8962), .Q(n8956) );
  AND2X1 U9894 ( .IN1(n8196), .IN2(n4921), .Q(n8962) );
  XOR2X1 U9895 ( .IN1(n8963), .IN2(n8964), .Q(n8196) );
  XOR2X1 U9896 ( .IN1(n4703), .IN2(n5380), .Q(n8964) );
  XOR2X1 U9897 ( .IN1(n8965), .IN2(n9743), .Q(n8963) );
  XOR2X1 U9898 ( .IN1(n9742), .IN2(n9741), .Q(n8965) );
  AND2X1 U9899 ( .IN1(n4847), .IN2(n7067), .Q(n8961) );
  XNOR2X1 U9900 ( .IN1(n8966), .IN2(n8967), .Q(n7067) );
  XOR2X1 U9901 ( .IN1(n4278), .IN2(n5380), .Q(n8967) );
  XOR2X1 U9902 ( .IN1(n8968), .IN2(n4729), .Q(n8966) );
  XNOR2X1 U9903 ( .IN1(WX2068), .IN2(n8668), .Q(n8968) );
  OR2X1 U9904 ( .IN1(n8969), .IN2(n8970), .Q(WX1937) );
  OR2X1 U9905 ( .IN1(n8971), .IN2(n8972), .Q(n8970) );
  AND2X1 U9906 ( .IN1(n2245), .IN2(WX1778), .Q(n8972) );
  AND2X1 U9907 ( .IN1(n4896), .IN2(CRC_OUT_8_31), .Q(n8971) );
  OR2X1 U9908 ( .IN1(n8973), .IN2(n8974), .Q(n8969) );
  AND2X1 U9909 ( .IN1(n4847), .IN2(n7087), .Q(n8974) );
  XNOR2X1 U9910 ( .IN1(n8975), .IN2(n8976), .Q(n7087) );
  XOR2X1 U9911 ( .IN1(n4172), .IN2(n5380), .Q(n8976) );
  XOR2X1 U9912 ( .IN1(n8977), .IN2(n4728), .Q(n8975) );
  XNOR2X1 U9913 ( .IN1(WX2066), .IN2(n8669), .Q(n8977) );
  AND2X1 U9914 ( .IN1(n4929), .IN2(n8206), .Q(n8973) );
  XNOR2X1 U9915 ( .IN1(n8978), .IN2(n8979), .Q(n8206) );
  XOR2X1 U9916 ( .IN1(n4171), .IN2(n5380), .Q(n8979) );
  XOR2X1 U9917 ( .IN1(n8980), .IN2(n4702), .Q(n8978) );
  XOR2X1 U9918 ( .IN1(WX3359), .IN2(n9744), .Q(n8980) );
  AND2X1 U9919 ( .IN1(n4819), .IN2(n5434), .Q(WX1839) );
  AND2X1 U9920 ( .IN1(n8981), .IN2(n5433), .Q(WX1326) );
  XOR2X1 U9921 ( .IN1(CRC_OUT_9_30), .IN2(n4789), .Q(n8981) );
  AND2X1 U9922 ( .IN1(n8982), .IN2(n5425), .Q(WX1324) );
  XOR2X1 U9923 ( .IN1(CRC_OUT_9_29), .IN2(n4755), .Q(n8982) );
  AND2X1 U9924 ( .IN1(n8983), .IN2(n5425), .Q(WX1322) );
  XOR2X1 U9925 ( .IN1(CRC_OUT_9_28), .IN2(n4758), .Q(n8983) );
  AND2X1 U9926 ( .IN1(n8984), .IN2(n5425), .Q(WX1320) );
  XOR2X1 U9927 ( .IN1(CRC_OUT_9_27), .IN2(n4762), .Q(n8984) );
  AND2X1 U9928 ( .IN1(n8985), .IN2(n5425), .Q(WX1318) );
  XOR2X1 U9929 ( .IN1(CRC_OUT_9_26), .IN2(n4765), .Q(n8985) );
  AND2X1 U9930 ( .IN1(n8986), .IN2(n5425), .Q(WX1316) );
  XOR2X1 U9931 ( .IN1(CRC_OUT_9_25), .IN2(n4766), .Q(n8986) );
  AND2X1 U9932 ( .IN1(n8987), .IN2(n5425), .Q(WX1314) );
  XOR2X1 U9933 ( .IN1(CRC_OUT_9_24), .IN2(n4770), .Q(n8987) );
  AND2X1 U9934 ( .IN1(n8988), .IN2(n5425), .Q(WX1312) );
  XOR2X1 U9935 ( .IN1(CRC_OUT_9_23), .IN2(n4773), .Q(n8988) );
  AND2X1 U9936 ( .IN1(n8989), .IN2(n5424), .Q(WX1310) );
  XOR2X1 U9937 ( .IN1(CRC_OUT_9_22), .IN2(n4775), .Q(n8989) );
  AND2X1 U9938 ( .IN1(n8990), .IN2(n5424), .Q(WX1308) );
  XOR2X1 U9939 ( .IN1(CRC_OUT_9_21), .IN2(n4781), .Q(n8990) );
  AND2X1 U9940 ( .IN1(n8991), .IN2(n5424), .Q(WX1306) );
  XOR2X1 U9941 ( .IN1(CRC_OUT_9_20), .IN2(n4785), .Q(n8991) );
  AND2X1 U9942 ( .IN1(n8992), .IN2(n5424), .Q(WX1304) );
  XOR2X1 U9943 ( .IN1(test_so10), .IN2(n4787), .Q(n8992) );
  AND2X1 U9944 ( .IN1(n8993), .IN2(n5424), .Q(WX1302) );
  XOR2X1 U9945 ( .IN1(CRC_OUT_9_18), .IN2(n4757), .Q(n8993) );
  AND2X1 U9946 ( .IN1(n8994), .IN2(n5424), .Q(WX1300) );
  XOR2X1 U9947 ( .IN1(CRC_OUT_9_17), .IN2(n4764), .Q(n8994) );
  AND2X1 U9948 ( .IN1(n8995), .IN2(n5424), .Q(WX1298) );
  XOR2X1 U9949 ( .IN1(CRC_OUT_9_16), .IN2(n4769), .Q(n8995) );
  AND2X1 U9950 ( .IN1(n8996), .IN2(n5424), .Q(WX1296) );
  XOR2X1 U9951 ( .IN1(CRC_OUT_9_15), .IN2(n8997), .Q(n8996) );
  XOR2X1 U9952 ( .IN1(test_so8), .IN2(DFF_191_n1), .Q(n8997) );
  AND2X1 U9953 ( .IN1(n8998), .IN2(n5424), .Q(WX1294) );
  XOR2X1 U9954 ( .IN1(CRC_OUT_9_14), .IN2(n4783), .Q(n8998) );
  AND2X1 U9955 ( .IN1(n8999), .IN2(n5423), .Q(WX1292) );
  XOR2X1 U9956 ( .IN1(CRC_OUT_9_13), .IN2(n4790), .Q(n8999) );
  AND2X1 U9957 ( .IN1(n9000), .IN2(n5423), .Q(WX1290) );
  XOR2X1 U9958 ( .IN1(CRC_OUT_9_12), .IN2(n4759), .Q(n9000) );
  AND2X1 U9959 ( .IN1(n9001), .IN2(n5423), .Q(WX1288) );
  XOR2X1 U9960 ( .IN1(CRC_OUT_9_11), .IN2(n4771), .Q(n9001) );
  AND2X1 U9961 ( .IN1(n9002), .IN2(n5423), .Q(WX1286) );
  XOR2X1 U9962 ( .IN1(DFF_170_n1), .IN2(n9003), .Q(n9002) );
  XOR2X1 U9963 ( .IN1(n4794), .IN2(DFF_191_n1), .Q(n9003) );
  AND2X1 U9964 ( .IN1(n9004), .IN2(n5423), .Q(WX1284) );
  XOR2X1 U9965 ( .IN1(CRC_OUT_9_9), .IN2(n4767), .Q(n9004) );
  AND2X1 U9966 ( .IN1(n9005), .IN2(n5423), .Q(WX1282) );
  XOR2X1 U9967 ( .IN1(CRC_OUT_9_8), .IN2(n4772), .Q(n9005) );
  AND2X1 U9968 ( .IN1(n9006), .IN2(n5423), .Q(WX1280) );
  XOR2X1 U9969 ( .IN1(CRC_OUT_9_7), .IN2(n4777), .Q(n9006) );
  AND2X1 U9970 ( .IN1(n9007), .IN2(n5423), .Q(WX1278) );
  XOR2X1 U9971 ( .IN1(CRC_OUT_9_6), .IN2(n4793), .Q(n9007) );
  AND2X1 U9972 ( .IN1(n9008), .IN2(n5423), .Q(WX1276) );
  XOR2X1 U9973 ( .IN1(CRC_OUT_9_5), .IN2(n4786), .Q(n9008) );
  AND2X1 U9974 ( .IN1(n9009), .IN2(n5422), .Q(WX1274) );
  XOR2X1 U9975 ( .IN1(CRC_OUT_9_4), .IN2(n4778), .Q(n9009) );
  AND2X1 U9976 ( .IN1(n9010), .IN2(n5422), .Q(WX1272) );
  XOR2X1 U9977 ( .IN1(DFF_163_n1), .IN2(n9011), .Q(n9010) );
  XOR2X1 U9978 ( .IN1(n4779), .IN2(DFF_191_n1), .Q(n9011) );
  AND2X1 U9979 ( .IN1(n9012), .IN2(n5422), .Q(WX1270) );
  XOR2X1 U9980 ( .IN1(CRC_OUT_9_2), .IN2(n4756), .Q(n9012) );
  AND2X1 U9981 ( .IN1(n9013), .IN2(n5422), .Q(WX1268) );
  XOR2X1 U9982 ( .IN1(test_so9), .IN2(n4791), .Q(n9013) );
  AND2X1 U9983 ( .IN1(n9014), .IN2(n5422), .Q(WX1266) );
  XOR2X1 U9984 ( .IN1(CRC_OUT_9_0), .IN2(n4760), .Q(n9014) );
  AND2X1 U9985 ( .IN1(n9015), .IN2(n5422), .Q(WX1264) );
  XOR2X1 U9986 ( .IN1(n4796), .IN2(CRC_OUT_9_31), .Q(n9015) );
  AND2X1 U9987 ( .IN1(n9016), .IN2(n5422), .Q(WX11670) );
  XOR2X1 U9988 ( .IN1(CRC_OUT_1_30), .IN2(n4542), .Q(n9016) );
  AND2X1 U9989 ( .IN1(n9017), .IN2(n5422), .Q(WX11668) );
  XOR2X1 U9990 ( .IN1(CRC_OUT_1_29), .IN2(n4543), .Q(n9017) );
  AND2X1 U9991 ( .IN1(n9018), .IN2(n5422), .Q(WX11666) );
  XOR2X1 U9992 ( .IN1(CRC_OUT_1_28), .IN2(n4544), .Q(n9018) );
  AND2X1 U9993 ( .IN1(n9019), .IN2(n5421), .Q(WX11664) );
  XOR2X1 U9994 ( .IN1(CRC_OUT_1_27), .IN2(n4545), .Q(n9019) );
  AND2X1 U9995 ( .IN1(n9020), .IN2(n5421), .Q(WX11662) );
  XOR2X1 U9996 ( .IN1(CRC_OUT_1_26), .IN2(n4546), .Q(n9020) );
  AND2X1 U9997 ( .IN1(n9021), .IN2(n5421), .Q(WX11660) );
  XOR2X1 U9998 ( .IN1(CRC_OUT_1_25), .IN2(n4547), .Q(n9021) );
  AND2X1 U9999 ( .IN1(n9022), .IN2(n5421), .Q(WX11658) );
  XOR2X1 U10000 ( .IN1(CRC_OUT_1_24), .IN2(n4548), .Q(n9022) );
  AND2X1 U10001 ( .IN1(n9023), .IN2(n5421), .Q(WX11656) );
  XOR2X1 U10002 ( .IN1(CRC_OUT_1_23), .IN2(n4549), .Q(n9023) );
  AND2X1 U10003 ( .IN1(n9024), .IN2(n5421), .Q(WX11654) );
  XOR2X1 U10004 ( .IN1(CRC_OUT_1_22), .IN2(n4550), .Q(n9024) );
  AND2X1 U10005 ( .IN1(n9025), .IN2(n5421), .Q(WX11652) );
  XOR2X1 U10006 ( .IN1(CRC_OUT_1_21), .IN2(n4551), .Q(n9025) );
  AND2X1 U10007 ( .IN1(n9026), .IN2(n5421), .Q(WX11650) );
  XOR2X1 U10008 ( .IN1(CRC_OUT_1_20), .IN2(n4552), .Q(n9026) );
  AND2X1 U10009 ( .IN1(n9027), .IN2(n5421), .Q(WX11648) );
  XOR2X1 U10010 ( .IN1(CRC_OUT_1_19), .IN2(n4553), .Q(n9027) );
  AND2X1 U10011 ( .IN1(n9028), .IN2(n5420), .Q(WX11646) );
  XOR2X1 U10012 ( .IN1(test_so97), .IN2(DFF_1714_n1), .Q(n9028) );
  AND2X1 U10013 ( .IN1(n9029), .IN2(n5420), .Q(WX11644) );
  XOR2X1 U10014 ( .IN1(CRC_OUT_1_17), .IN2(n4554), .Q(n9029) );
  AND2X1 U10015 ( .IN1(n9030), .IN2(n5420), .Q(WX11642) );
  XOR2X1 U10016 ( .IN1(CRC_OUT_1_16), .IN2(n4555), .Q(n9030) );
  AND2X1 U10017 ( .IN1(n9031), .IN2(n5420), .Q(WX11640) );
  XOR2X1 U10018 ( .IN1(CRC_OUT_1_15), .IN2(n9032), .Q(n9031) );
  XOR2X1 U10019 ( .IN1(test_so100), .IN2(n4513), .Q(n9032) );
  AND2X1 U10020 ( .IN1(n9033), .IN2(n5420), .Q(WX11638) );
  XOR2X1 U10021 ( .IN1(test_so99), .IN2(n4556), .Q(n9033) );
  AND2X1 U10022 ( .IN1(n9034), .IN2(n5420), .Q(WX11636) );
  XOR2X1 U10023 ( .IN1(CRC_OUT_1_13), .IN2(n4557), .Q(n9034) );
  AND2X1 U10024 ( .IN1(n9035), .IN2(n5420), .Q(WX11634) );
  XOR2X1 U10025 ( .IN1(CRC_OUT_1_12), .IN2(n4558), .Q(n9035) );
  AND2X1 U10026 ( .IN1(n9036), .IN2(n5420), .Q(WX11632) );
  XOR2X1 U10027 ( .IN1(CRC_OUT_1_11), .IN2(n4559), .Q(n9036) );
  AND2X1 U10028 ( .IN1(n9037), .IN2(n5420), .Q(WX11630) );
  XOR2X1 U10029 ( .IN1(CRC_OUT_1_10), .IN2(n9038), .Q(n9037) );
  XOR2X1 U10030 ( .IN1(test_so100), .IN2(n4514), .Q(n9038) );
  AND2X1 U10031 ( .IN1(n9039), .IN2(n5419), .Q(WX11628) );
  XOR2X1 U10032 ( .IN1(CRC_OUT_1_9), .IN2(n4560), .Q(n9039) );
  AND2X1 U10033 ( .IN1(n9040), .IN2(n5419), .Q(WX11626) );
  XOR2X1 U10034 ( .IN1(CRC_OUT_1_8), .IN2(n4561), .Q(n9040) );
  AND2X1 U10035 ( .IN1(n9041), .IN2(n5419), .Q(WX11624) );
  XOR2X1 U10036 ( .IN1(CRC_OUT_1_7), .IN2(n4562), .Q(n9041) );
  AND2X1 U10037 ( .IN1(n9042), .IN2(n5419), .Q(WX11622) );
  XOR2X1 U10038 ( .IN1(CRC_OUT_1_6), .IN2(n4563), .Q(n9042) );
  AND2X1 U10039 ( .IN1(n9043), .IN2(n5419), .Q(WX11620) );
  XOR2X1 U10040 ( .IN1(CRC_OUT_1_5), .IN2(n4564), .Q(n9043) );
  AND2X1 U10041 ( .IN1(n9044), .IN2(n5419), .Q(WX11618) );
  XOR2X1 U10042 ( .IN1(CRC_OUT_1_4), .IN2(n4565), .Q(n9044) );
  AND2X1 U10043 ( .IN1(n9045), .IN2(n5419), .Q(WX11616) );
  XOR2X1 U10044 ( .IN1(CRC_OUT_1_3), .IN2(n9046), .Q(n9045) );
  XOR2X1 U10045 ( .IN1(test_so100), .IN2(n4515), .Q(n9046) );
  AND2X1 U10046 ( .IN1(n9047), .IN2(n5419), .Q(WX11614) );
  XOR2X1 U10047 ( .IN1(CRC_OUT_1_2), .IN2(n4566), .Q(n9047) );
  AND2X1 U10048 ( .IN1(n9048), .IN2(n5419), .Q(WX11612) );
  XOR2X1 U10049 ( .IN1(test_so98), .IN2(DFF_1697_n1), .Q(n9048) );
  AND2X1 U10050 ( .IN1(n9049), .IN2(n5418), .Q(WX11610) );
  XOR2X1 U10051 ( .IN1(CRC_OUT_1_0), .IN2(n4567), .Q(n9049) );
  AND2X1 U10052 ( .IN1(n9050), .IN2(n5418), .Q(WX11608) );
  XOR2X1 U10053 ( .IN1(test_so100), .IN2(n4534), .Q(n9050) );
  AND2X1 U10054 ( .IN1(n5434), .IN2(n8246), .Q(WX11082) );
  AND2X1 U10055 ( .IN1(n5435), .IN2(n8247), .Q(WX11080) );
  AND2X1 U10056 ( .IN1(n5436), .IN2(n8248), .Q(WX11078) );
  AND2X1 U10057 ( .IN1(n5435), .IN2(n8249), .Q(WX11076) );
  AND2X1 U10058 ( .IN1(n5434), .IN2(n8250), .Q(WX11074) );
  AND2X1 U10059 ( .IN1(n5435), .IN2(n8251), .Q(WX11072) );
  AND2X1 U10060 ( .IN1(n5435), .IN2(n8252), .Q(WX11070) );
  AND2X1 U10061 ( .IN1(n5435), .IN2(n8253), .Q(WX11068) );
  AND2X1 U10062 ( .IN1(n5435), .IN2(n8254), .Q(WX11066) );
  AND2X1 U10063 ( .IN1(test_so91), .IN2(n5418), .Q(WX11064) );
  AND2X1 U10064 ( .IN1(n5435), .IN2(n8257), .Q(WX11062) );
  AND2X1 U10065 ( .IN1(n5437), .IN2(n8258), .Q(WX11060) );
  AND2X1 U10066 ( .IN1(n5436), .IN2(n8259), .Q(WX11058) );
  AND2X1 U10067 ( .IN1(n5436), .IN2(n8260), .Q(WX11056) );
  AND2X1 U10068 ( .IN1(n5435), .IN2(n8261), .Q(WX11054) );
  AND2X1 U10069 ( .IN1(n5436), .IN2(n8262), .Q(WX11052) );
  OR2X1 U10070 ( .IN1(n9051), .IN2(n9052), .Q(WX11050) );
  OR2X1 U10071 ( .IN1(n9053), .IN2(n9054), .Q(n9052) );
  AND2X1 U10072 ( .IN1(n4896), .IN2(CRC_OUT_1_0), .Q(n9054) );
  AND2X1 U10073 ( .IN1(DATA_0_0), .IN2(n4920), .Q(n9053) );
  OR2X1 U10074 ( .IN1(n9055), .IN2(n9056), .Q(n9051) );
  AND2X1 U10075 ( .IN1(n498), .IN2(n4863), .Q(n9056) );
  INVX0 U10076 ( .INP(n9057), .ZN(n498) );
  OR2X1 U10077 ( .IN1(n5476), .IN2(n3786), .Q(n9057) );
  AND2X1 U10078 ( .IN1(n4847), .IN2(n5747), .Q(n9055) );
  XNOR2X1 U10079 ( .IN1(n9058), .IN2(n9059), .Q(n5747) );
  XOR2X1 U10080 ( .IN1(n9745), .IN2(n4534), .Q(n9059) );
  XOR2X1 U10081 ( .IN1(WX11051), .IN2(n4280), .Q(n9058) );
  OR2X1 U10082 ( .IN1(n9060), .IN2(n9061), .Q(WX11048) );
  OR2X1 U10083 ( .IN1(n9062), .IN2(n9063), .Q(n9061) );
  AND2X1 U10084 ( .IN1(n4896), .IN2(CRC_OUT_1_1), .Q(n9063) );
  AND2X1 U10085 ( .IN1(DATA_0_1), .IN2(n4921), .Q(n9062) );
  OR2X1 U10086 ( .IN1(n9064), .IN2(n9065), .Q(n9060) );
  AND2X1 U10087 ( .IN1(n497), .IN2(n4863), .Q(n9065) );
  INVX0 U10088 ( .INP(n9066), .ZN(n497) );
  OR2X1 U10089 ( .IN1(n5476), .IN2(n3787), .Q(n9066) );
  AND2X1 U10090 ( .IN1(n4847), .IN2(n5757), .Q(n9064) );
  XNOR2X1 U10091 ( .IN1(n9067), .IN2(n9068), .Q(n5757) );
  XOR2X1 U10092 ( .IN1(n9746), .IN2(n4567), .Q(n9068) );
  XOR2X1 U10093 ( .IN1(WX11049), .IN2(n4282), .Q(n9067) );
  OR2X1 U10094 ( .IN1(n9069), .IN2(n9070), .Q(WX11046) );
  OR2X1 U10095 ( .IN1(n9071), .IN2(n9072), .Q(n9070) );
  AND2X1 U10096 ( .IN1(n4896), .IN2(CRC_OUT_1_2), .Q(n9072) );
  AND2X1 U10097 ( .IN1(DATA_0_2), .IN2(n4922), .Q(n9071) );
  OR2X1 U10098 ( .IN1(n9073), .IN2(n9074), .Q(n9069) );
  AND2X1 U10099 ( .IN1(n496), .IN2(n4863), .Q(n9074) );
  INVX0 U10100 ( .INP(n9075), .ZN(n496) );
  OR2X1 U10101 ( .IN1(n5476), .IN2(n3788), .Q(n9075) );
  AND2X1 U10102 ( .IN1(n5766), .IN2(n4834), .Q(n9073) );
  XOR2X1 U10103 ( .IN1(n9076), .IN2(n9077), .Q(n5766) );
  XOR2X1 U10104 ( .IN1(test_so98), .IN2(n9747), .Q(n9077) );
  XOR2X1 U10105 ( .IN1(WX11047), .IN2(n4284), .Q(n9076) );
  OR2X1 U10106 ( .IN1(n9078), .IN2(n9079), .Q(WX11044) );
  OR2X1 U10107 ( .IN1(n9080), .IN2(n9081), .Q(n9079) );
  AND2X1 U10108 ( .IN1(n4896), .IN2(CRC_OUT_1_3), .Q(n9081) );
  AND2X1 U10109 ( .IN1(DATA_0_3), .IN2(n4922), .Q(n9080) );
  OR2X1 U10110 ( .IN1(n9082), .IN2(n9083), .Q(n9078) );
  AND2X1 U10111 ( .IN1(n495), .IN2(n4863), .Q(n9083) );
  INVX0 U10112 ( .INP(n9084), .ZN(n495) );
  OR2X1 U10113 ( .IN1(n5476), .IN2(n3789), .Q(n9084) );
  AND2X1 U10114 ( .IN1(n4847), .IN2(n5775), .Q(n9082) );
  XNOR2X1 U10115 ( .IN1(n9085), .IN2(n9086), .Q(n5775) );
  XOR2X1 U10116 ( .IN1(n9748), .IN2(n4566), .Q(n9086) );
  XOR2X1 U10117 ( .IN1(WX11045), .IN2(n4286), .Q(n9085) );
  OR2X1 U10118 ( .IN1(n9087), .IN2(n9088), .Q(WX11042) );
  OR2X1 U10119 ( .IN1(n9089), .IN2(n9090), .Q(n9088) );
  AND2X1 U10120 ( .IN1(n4896), .IN2(CRC_OUT_1_4), .Q(n9090) );
  AND2X1 U10121 ( .IN1(DATA_0_4), .IN2(n4922), .Q(n9089) );
  OR2X1 U10122 ( .IN1(n9091), .IN2(n9092), .Q(n9087) );
  AND2X1 U10123 ( .IN1(n494), .IN2(n4863), .Q(n9092) );
  INVX0 U10124 ( .INP(n9093), .ZN(n494) );
  OR2X1 U10125 ( .IN1(n5475), .IN2(n3790), .Q(n9093) );
  AND2X1 U10126 ( .IN1(n5784), .IN2(n4834), .Q(n9091) );
  XOR2X1 U10127 ( .IN1(n9094), .IN2(n9095), .Q(n5784) );
  XOR2X1 U10128 ( .IN1(test_so96), .IN2(n9749), .Q(n9095) );
  XOR2X1 U10129 ( .IN1(WX11043), .IN2(n4515), .Q(n9094) );
  OR2X1 U10130 ( .IN1(n9096), .IN2(n9097), .Q(WX11040) );
  OR2X1 U10131 ( .IN1(n9098), .IN2(n9099), .Q(n9097) );
  AND2X1 U10132 ( .IN1(n4896), .IN2(CRC_OUT_1_5), .Q(n9099) );
  AND2X1 U10133 ( .IN1(DATA_0_5), .IN2(n4922), .Q(n9098) );
  OR2X1 U10134 ( .IN1(n9100), .IN2(n9101), .Q(n9096) );
  AND2X1 U10135 ( .IN1(n493), .IN2(n4863), .Q(n9101) );
  INVX0 U10136 ( .INP(n9102), .ZN(n493) );
  OR2X1 U10137 ( .IN1(n5475), .IN2(n3791), .Q(n9102) );
  AND2X1 U10138 ( .IN1(n4847), .IN2(n5793), .Q(n9100) );
  XNOR2X1 U10139 ( .IN1(n9103), .IN2(n9104), .Q(n5793) );
  XOR2X1 U10140 ( .IN1(n9750), .IN2(n4565), .Q(n9104) );
  XOR2X1 U10141 ( .IN1(WX11041), .IN2(n4289), .Q(n9103) );
  OR2X1 U10142 ( .IN1(n9105), .IN2(n9106), .Q(WX11038) );
  OR2X1 U10143 ( .IN1(n9107), .IN2(n9108), .Q(n9106) );
  AND2X1 U10144 ( .IN1(n4896), .IN2(CRC_OUT_1_6), .Q(n9108) );
  AND2X1 U10145 ( .IN1(DATA_0_6), .IN2(n4922), .Q(n9107) );
  OR2X1 U10146 ( .IN1(n9109), .IN2(n9110), .Q(n9105) );
  AND2X1 U10147 ( .IN1(n492), .IN2(n4863), .Q(n9110) );
  INVX0 U10148 ( .INP(n9111), .ZN(n492) );
  OR2X1 U10149 ( .IN1(n5475), .IN2(n3792), .Q(n9111) );
  AND2X1 U10150 ( .IN1(n5802), .IN2(n4834), .Q(n9109) );
  XOR2X1 U10151 ( .IN1(n9112), .IN2(n9113), .Q(n5802) );
  XOR2X1 U10152 ( .IN1(test_so94), .IN2(n9751), .Q(n9113) );
  XOR2X1 U10153 ( .IN1(WX11039), .IN2(n4564), .Q(n9112) );
  OR2X1 U10154 ( .IN1(n9114), .IN2(n9115), .Q(WX11036) );
  OR2X1 U10155 ( .IN1(n9116), .IN2(n9117), .Q(n9115) );
  AND2X1 U10156 ( .IN1(n4896), .IN2(CRC_OUT_1_7), .Q(n9117) );
  AND2X1 U10157 ( .IN1(DATA_0_7), .IN2(n4923), .Q(n9116) );
  OR2X1 U10158 ( .IN1(n9118), .IN2(n9119), .Q(n9114) );
  AND2X1 U10159 ( .IN1(n491), .IN2(n4862), .Q(n9119) );
  INVX0 U10160 ( .INP(n9120), .ZN(n491) );
  OR2X1 U10161 ( .IN1(n5475), .IN2(n3793), .Q(n9120) );
  AND2X1 U10162 ( .IN1(n4847), .IN2(n5811), .Q(n9118) );
  XNOR2X1 U10163 ( .IN1(n9121), .IN2(n9122), .Q(n5811) );
  XOR2X1 U10164 ( .IN1(n9752), .IN2(n4563), .Q(n9122) );
  XOR2X1 U10165 ( .IN1(WX11037), .IN2(n4292), .Q(n9121) );
  OR2X1 U10166 ( .IN1(n9123), .IN2(n9124), .Q(WX11034) );
  OR2X1 U10167 ( .IN1(n9125), .IN2(n9126), .Q(n9124) );
  AND2X1 U10168 ( .IN1(n4896), .IN2(CRC_OUT_1_8), .Q(n9126) );
  AND2X1 U10169 ( .IN1(DATA_0_8), .IN2(n4923), .Q(n9125) );
  OR2X1 U10170 ( .IN1(n9127), .IN2(n9128), .Q(n9123) );
  AND2X1 U10171 ( .IN1(n490), .IN2(n4862), .Q(n9128) );
  INVX0 U10172 ( .INP(n9129), .ZN(n490) );
  OR2X1 U10173 ( .IN1(n5475), .IN2(n3794), .Q(n9129) );
  AND2X1 U10174 ( .IN1(n5820), .IN2(n4834), .Q(n9127) );
  XOR2X1 U10175 ( .IN1(n9130), .IN2(n9131), .Q(n5820) );
  XOR2X1 U10176 ( .IN1(test_so92), .IN2(n9753), .Q(n9131) );
  XOR2X1 U10177 ( .IN1(WX11163), .IN2(n4562), .Q(n9130) );
  OR2X1 U10178 ( .IN1(n9132), .IN2(n9133), .Q(WX11032) );
  OR2X1 U10179 ( .IN1(n9134), .IN2(n9135), .Q(n9133) );
  AND2X1 U10180 ( .IN1(n4896), .IN2(CRC_OUT_1_9), .Q(n9135) );
  AND2X1 U10181 ( .IN1(DATA_0_9), .IN2(n4923), .Q(n9134) );
  OR2X1 U10182 ( .IN1(n9136), .IN2(n9137), .Q(n9132) );
  AND2X1 U10183 ( .IN1(n489), .IN2(n4862), .Q(n9137) );
  INVX0 U10184 ( .INP(n9138), .ZN(n489) );
  OR2X1 U10185 ( .IN1(n5475), .IN2(n3795), .Q(n9138) );
  AND2X1 U10186 ( .IN1(n4847), .IN2(n5829), .Q(n9136) );
  XNOR2X1 U10187 ( .IN1(n9139), .IN2(n9140), .Q(n5829) );
  XOR2X1 U10188 ( .IN1(n9754), .IN2(n4561), .Q(n9140) );
  XOR2X1 U10189 ( .IN1(WX11033), .IN2(n4295), .Q(n9139) );
  OR2X1 U10190 ( .IN1(n9141), .IN2(n9142), .Q(WX11030) );
  OR2X1 U10191 ( .IN1(n9143), .IN2(n9144), .Q(n9142) );
  AND2X1 U10192 ( .IN1(n4897), .IN2(CRC_OUT_1_10), .Q(n9144) );
  AND2X1 U10193 ( .IN1(DATA_0_10), .IN2(n4923), .Q(n9143) );
  OR2X1 U10194 ( .IN1(n9145), .IN2(n9146), .Q(n9141) );
  AND2X1 U10195 ( .IN1(n488), .IN2(n4862), .Q(n9146) );
  INVX0 U10196 ( .INP(n9147), .ZN(n488) );
  OR2X1 U10197 ( .IN1(n5475), .IN2(n3796), .Q(n9147) );
  AND2X1 U10198 ( .IN1(n4847), .IN2(n5838), .Q(n9145) );
  XNOR2X1 U10199 ( .IN1(n9148), .IN2(n9149), .Q(n5838) );
  XOR2X1 U10200 ( .IN1(n9755), .IN2(n4560), .Q(n9149) );
  XOR2X1 U10201 ( .IN1(WX11031), .IN2(n4297), .Q(n9148) );
  OR2X1 U10202 ( .IN1(n9150), .IN2(n9151), .Q(WX11028) );
  OR2X1 U10203 ( .IN1(n9152), .IN2(n9153), .Q(n9151) );
  AND2X1 U10204 ( .IN1(n4897), .IN2(CRC_OUT_1_11), .Q(n9153) );
  AND2X1 U10205 ( .IN1(DATA_0_11), .IN2(n4921), .Q(n9152) );
  OR2X1 U10206 ( .IN1(n9154), .IN2(n9155), .Q(n9150) );
  AND2X1 U10207 ( .IN1(n487), .IN2(n4862), .Q(n9155) );
  INVX0 U10208 ( .INP(n9156), .ZN(n487) );
  OR2X1 U10209 ( .IN1(n5475), .IN2(n3797), .Q(n9156) );
  AND2X1 U10210 ( .IN1(n4847), .IN2(n5847), .Q(n9154) );
  XNOR2X1 U10211 ( .IN1(n9157), .IN2(n9158), .Q(n5847) );
  XOR2X1 U10212 ( .IN1(n9756), .IN2(n4514), .Q(n9158) );
  XOR2X1 U10213 ( .IN1(WX11029), .IN2(n4299), .Q(n9157) );
  OR2X1 U10214 ( .IN1(n9159), .IN2(n9160), .Q(WX11026) );
  OR2X1 U10215 ( .IN1(n9161), .IN2(n9162), .Q(n9160) );
  AND2X1 U10216 ( .IN1(n4897), .IN2(CRC_OUT_1_12), .Q(n9162) );
  AND2X1 U10217 ( .IN1(DATA_0_12), .IN2(n4923), .Q(n9161) );
  OR2X1 U10218 ( .IN1(n9163), .IN2(n9164), .Q(n9159) );
  AND2X1 U10219 ( .IN1(n486), .IN2(n4862), .Q(n9164) );
  INVX0 U10220 ( .INP(n9165), .ZN(n486) );
  OR2X1 U10221 ( .IN1(n5475), .IN2(n3798), .Q(n9165) );
  AND2X1 U10222 ( .IN1(n4846), .IN2(n5856), .Q(n9163) );
  XNOR2X1 U10223 ( .IN1(n9166), .IN2(n9167), .Q(n5856) );
  XOR2X1 U10224 ( .IN1(n9757), .IN2(n4559), .Q(n9167) );
  XOR2X1 U10225 ( .IN1(WX11027), .IN2(n4301), .Q(n9166) );
  OR2X1 U10226 ( .IN1(n9168), .IN2(n9169), .Q(WX11024) );
  OR2X1 U10227 ( .IN1(n9170), .IN2(n9171), .Q(n9169) );
  AND2X1 U10228 ( .IN1(n4897), .IN2(CRC_OUT_1_13), .Q(n9171) );
  AND2X1 U10229 ( .IN1(DATA_0_13), .IN2(n4923), .Q(n9170) );
  OR2X1 U10230 ( .IN1(n9172), .IN2(n9173), .Q(n9168) );
  AND2X1 U10231 ( .IN1(n485), .IN2(n4862), .Q(n9173) );
  INVX0 U10232 ( .INP(n9174), .ZN(n485) );
  OR2X1 U10233 ( .IN1(n5475), .IN2(n3799), .Q(n9174) );
  AND2X1 U10234 ( .IN1(n4846), .IN2(n5865), .Q(n9172) );
  XNOR2X1 U10235 ( .IN1(n9175), .IN2(n9176), .Q(n5865) );
  XOR2X1 U10236 ( .IN1(n9758), .IN2(n4558), .Q(n9176) );
  XOR2X1 U10237 ( .IN1(WX11025), .IN2(n4303), .Q(n9175) );
  OR2X1 U10238 ( .IN1(n9177), .IN2(n9178), .Q(WX11022) );
  OR2X1 U10239 ( .IN1(n9179), .IN2(n9180), .Q(n9178) );
  AND2X1 U10240 ( .IN1(test_so99), .IN2(n4887), .Q(n9180) );
  AND2X1 U10241 ( .IN1(DATA_0_14), .IN2(n4924), .Q(n9179) );
  OR2X1 U10242 ( .IN1(n9181), .IN2(n9182), .Q(n9177) );
  AND2X1 U10243 ( .IN1(n484), .IN2(n4862), .Q(n9182) );
  INVX0 U10244 ( .INP(n9183), .ZN(n484) );
  OR2X1 U10245 ( .IN1(n5475), .IN2(n3800), .Q(n9183) );
  AND2X1 U10246 ( .IN1(n4846), .IN2(n5874), .Q(n9181) );
  XNOR2X1 U10247 ( .IN1(n9184), .IN2(n9185), .Q(n5874) );
  XOR2X1 U10248 ( .IN1(n9759), .IN2(n4557), .Q(n9185) );
  XOR2X1 U10249 ( .IN1(WX11023), .IN2(n4305), .Q(n9184) );
  OR2X1 U10250 ( .IN1(n9186), .IN2(n9187), .Q(WX11020) );
  OR2X1 U10251 ( .IN1(n9188), .IN2(n9189), .Q(n9187) );
  AND2X1 U10252 ( .IN1(n4897), .IN2(CRC_OUT_1_15), .Q(n9189) );
  AND2X1 U10253 ( .IN1(DATA_0_15), .IN2(n4924), .Q(n9188) );
  OR2X1 U10254 ( .IN1(n9190), .IN2(n9191), .Q(n9186) );
  AND2X1 U10255 ( .IN1(n483), .IN2(n4862), .Q(n9191) );
  INVX0 U10256 ( .INP(n9192), .ZN(n483) );
  OR2X1 U10257 ( .IN1(n5475), .IN2(n3801), .Q(n9192) );
  AND2X1 U10258 ( .IN1(n4846), .IN2(n5883), .Q(n9190) );
  XNOR2X1 U10259 ( .IN1(n9193), .IN2(n9194), .Q(n5883) );
  XOR2X1 U10260 ( .IN1(n9760), .IN2(n4556), .Q(n9194) );
  XOR2X1 U10261 ( .IN1(WX11021), .IN2(n4307), .Q(n9193) );
  OR2X1 U10262 ( .IN1(n9195), .IN2(n9196), .Q(WX11018) );
  OR2X1 U10263 ( .IN1(n9197), .IN2(n9198), .Q(n9196) );
  AND2X1 U10264 ( .IN1(n4897), .IN2(CRC_OUT_1_16), .Q(n9198) );
  AND2X1 U10265 ( .IN1(DATA_0_16), .IN2(n4923), .Q(n9197) );
  OR2X1 U10266 ( .IN1(n9199), .IN2(n9200), .Q(n9195) );
  AND2X1 U10267 ( .IN1(n482), .IN2(n4862), .Q(n9200) );
  INVX0 U10268 ( .INP(n9201), .ZN(n482) );
  OR2X1 U10269 ( .IN1(n5475), .IN2(n3802), .Q(n9201) );
  AND2X1 U10270 ( .IN1(n4846), .IN2(n5892), .Q(n9199) );
  XNOR2X1 U10271 ( .IN1(n9202), .IN2(n9203), .Q(n5892) );
  XOR2X1 U10272 ( .IN1(n4173), .IN2(n5380), .Q(n9203) );
  XOR2X1 U10273 ( .IN1(n9204), .IN2(n4513), .Q(n9202) );
  XNOR2X1 U10274 ( .IN1(WX11147), .IN2(n8246), .Q(n9204) );
  OR2X1 U10275 ( .IN1(n9205), .IN2(n9206), .Q(WX11016) );
  OR2X1 U10276 ( .IN1(n9207), .IN2(n9208), .Q(n9206) );
  AND2X1 U10277 ( .IN1(n4897), .IN2(CRC_OUT_1_17), .Q(n9208) );
  AND2X1 U10278 ( .IN1(DATA_0_17), .IN2(n4924), .Q(n9207) );
  OR2X1 U10279 ( .IN1(n9209), .IN2(n9210), .Q(n9205) );
  AND2X1 U10280 ( .IN1(n481), .IN2(n4862), .Q(n9210) );
  INVX0 U10281 ( .INP(n9211), .ZN(n481) );
  OR2X1 U10282 ( .IN1(n5474), .IN2(n3803), .Q(n9211) );
  AND2X1 U10283 ( .IN1(n4846), .IN2(n5901), .Q(n9209) );
  XNOR2X1 U10284 ( .IN1(n9212), .IN2(n9213), .Q(n5901) );
  XOR2X1 U10285 ( .IN1(n4174), .IN2(n5380), .Q(n9213) );
  XOR2X1 U10286 ( .IN1(n9214), .IN2(n4555), .Q(n9212) );
  XNOR2X1 U10287 ( .IN1(WX11145), .IN2(n8247), .Q(n9214) );
  OR2X1 U10288 ( .IN1(n9215), .IN2(n9216), .Q(WX11014) );
  OR2X1 U10289 ( .IN1(n9217), .IN2(n9218), .Q(n9216) );
  AND2X1 U10290 ( .IN1(n4897), .IN2(CRC_OUT_1_18), .Q(n9218) );
  AND2X1 U10291 ( .IN1(DATA_0_18), .IN2(n4922), .Q(n9217) );
  OR2X1 U10292 ( .IN1(n9219), .IN2(n9220), .Q(n9215) );
  AND2X1 U10293 ( .IN1(n480), .IN2(n4862), .Q(n9220) );
  INVX0 U10294 ( .INP(n9221), .ZN(n480) );
  OR2X1 U10295 ( .IN1(n5474), .IN2(n3804), .Q(n9221) );
  AND2X1 U10296 ( .IN1(n4846), .IN2(n5910), .Q(n9219) );
  XNOR2X1 U10297 ( .IN1(n9222), .IN2(n9223), .Q(n5910) );
  XOR2X1 U10298 ( .IN1(n4175), .IN2(n5380), .Q(n9223) );
  XOR2X1 U10299 ( .IN1(n9224), .IN2(n4554), .Q(n9222) );
  XNOR2X1 U10300 ( .IN1(WX11143), .IN2(n8248), .Q(n9224) );
  OR2X1 U10301 ( .IN1(n9225), .IN2(n9226), .Q(WX11012) );
  OR2X1 U10302 ( .IN1(n9227), .IN2(n9228), .Q(n9226) );
  AND2X1 U10303 ( .IN1(n4897), .IN2(CRC_OUT_1_19), .Q(n9228) );
  AND2X1 U10304 ( .IN1(DATA_0_19), .IN2(n4921), .Q(n9227) );
  OR2X1 U10305 ( .IN1(n9229), .IN2(n9230), .Q(n9225) );
  AND2X1 U10306 ( .IN1(n479), .IN2(n4861), .Q(n9230) );
  INVX0 U10307 ( .INP(n9231), .ZN(n479) );
  OR2X1 U10308 ( .IN1(n5474), .IN2(n3805), .Q(n9231) );
  AND2X1 U10309 ( .IN1(n5919), .IN2(n4833), .Q(n9229) );
  XOR2X1 U10310 ( .IN1(n9232), .IN2(n9233), .Q(n5919) );
  XOR2X1 U10311 ( .IN1(n4176), .IN2(n5380), .Q(n9233) );
  XOR2X1 U10312 ( .IN1(WX11077), .IN2(n9234), .Q(n9232) );
  XNOR2X1 U10313 ( .IN1(test_so97), .IN2(n8249), .Q(n9234) );
  OR2X1 U10314 ( .IN1(n9235), .IN2(n9236), .Q(WX11010) );
  OR2X1 U10315 ( .IN1(n9237), .IN2(n9238), .Q(n9236) );
  AND2X1 U10316 ( .IN1(n4897), .IN2(CRC_OUT_1_20), .Q(n9238) );
  AND2X1 U10317 ( .IN1(DATA_0_20), .IN2(n4924), .Q(n9237) );
  OR2X1 U10318 ( .IN1(n9239), .IN2(n9240), .Q(n9235) );
  AND2X1 U10319 ( .IN1(n478), .IN2(n4861), .Q(n9240) );
  INVX0 U10320 ( .INP(n9241), .ZN(n478) );
  OR2X1 U10321 ( .IN1(n5474), .IN2(n3806), .Q(n9241) );
  AND2X1 U10322 ( .IN1(n4846), .IN2(n5928), .Q(n9239) );
  XNOR2X1 U10323 ( .IN1(n9242), .IN2(n9243), .Q(n5928) );
  XOR2X1 U10324 ( .IN1(n4177), .IN2(n5380), .Q(n9243) );
  XOR2X1 U10325 ( .IN1(n9244), .IN2(n4553), .Q(n9242) );
  XNOR2X1 U10326 ( .IN1(WX11139), .IN2(n8250), .Q(n9244) );
  OR2X1 U10327 ( .IN1(n9245), .IN2(n9246), .Q(WX11008) );
  OR2X1 U10328 ( .IN1(n9247), .IN2(n9248), .Q(n9246) );
  AND2X1 U10329 ( .IN1(n4897), .IN2(CRC_OUT_1_21), .Q(n9248) );
  AND2X1 U10330 ( .IN1(DATA_0_21), .IN2(n4922), .Q(n9247) );
  OR2X1 U10331 ( .IN1(n9249), .IN2(n9250), .Q(n9245) );
  AND2X1 U10332 ( .IN1(n477), .IN2(n4861), .Q(n9250) );
  INVX0 U10333 ( .INP(n9251), .ZN(n477) );
  OR2X1 U10334 ( .IN1(n5474), .IN2(n3807), .Q(n9251) );
  AND2X1 U10335 ( .IN1(n5937), .IN2(n4833), .Q(n9249) );
  XOR2X1 U10336 ( .IN1(n9252), .IN2(n9253), .Q(n5937) );
  XOR2X1 U10337 ( .IN1(n4552), .IN2(n5380), .Q(n9253) );
  XOR2X1 U10338 ( .IN1(n9254), .IN2(n9762), .Q(n9252) );
  XNOR2X1 U10339 ( .IN1(n9761), .IN2(n8251), .Q(n9254) );
  OR2X1 U10340 ( .IN1(n9255), .IN2(n9256), .Q(WX11006) );
  OR2X1 U10341 ( .IN1(n9257), .IN2(n9258), .Q(n9256) );
  AND2X1 U10342 ( .IN1(n4897), .IN2(CRC_OUT_1_22), .Q(n9258) );
  AND2X1 U10343 ( .IN1(DATA_0_22), .IN2(n4923), .Q(n9257) );
  OR2X1 U10344 ( .IN1(n9259), .IN2(n9260), .Q(n9255) );
  AND2X1 U10345 ( .IN1(n476), .IN2(n4861), .Q(n9260) );
  INVX0 U10346 ( .INP(n9261), .ZN(n476) );
  OR2X1 U10347 ( .IN1(n5474), .IN2(n3808), .Q(n9261) );
  AND2X1 U10348 ( .IN1(n4846), .IN2(n5946), .Q(n9259) );
  XNOR2X1 U10349 ( .IN1(n9262), .IN2(n9263), .Q(n5946) );
  XOR2X1 U10350 ( .IN1(n4178), .IN2(n5380), .Q(n9263) );
  XOR2X1 U10351 ( .IN1(n9264), .IN2(n4551), .Q(n9262) );
  XNOR2X1 U10352 ( .IN1(WX11135), .IN2(n8252), .Q(n9264) );
  OR2X1 U10353 ( .IN1(n9265), .IN2(n9266), .Q(WX11004) );
  OR2X1 U10354 ( .IN1(n9267), .IN2(n9268), .Q(n9266) );
  AND2X1 U10355 ( .IN1(n4897), .IN2(CRC_OUT_1_23), .Q(n9268) );
  AND2X1 U10356 ( .IN1(DATA_0_23), .IN2(n4921), .Q(n9267) );
  OR2X1 U10357 ( .IN1(n9269), .IN2(n9270), .Q(n9265) );
  AND2X1 U10358 ( .IN1(n475), .IN2(n4861), .Q(n9270) );
  INVX0 U10359 ( .INP(n9271), .ZN(n475) );
  OR2X1 U10360 ( .IN1(n5474), .IN2(n3809), .Q(n9271) );
  AND2X1 U10361 ( .IN1(n5955), .IN2(n4833), .Q(n9269) );
  XOR2X1 U10362 ( .IN1(n9272), .IN2(n9273), .Q(n5955) );
  XOR2X1 U10363 ( .IN1(n4550), .IN2(n5380), .Q(n9273) );
  XOR2X1 U10364 ( .IN1(n9274), .IN2(n9764), .Q(n9272) );
  XNOR2X1 U10365 ( .IN1(n9763), .IN2(n8253), .Q(n9274) );
  OR2X1 U10366 ( .IN1(n9275), .IN2(n9276), .Q(WX11002) );
  OR2X1 U10367 ( .IN1(n9277), .IN2(n9278), .Q(n9276) );
  AND2X1 U10368 ( .IN1(n4898), .IN2(CRC_OUT_1_24), .Q(n9278) );
  AND2X1 U10369 ( .IN1(DATA_0_24), .IN2(n4922), .Q(n9277) );
  OR2X1 U10370 ( .IN1(n9279), .IN2(n9280), .Q(n9275) );
  AND2X1 U10371 ( .IN1(n474), .IN2(n4861), .Q(n9280) );
  INVX0 U10372 ( .INP(n9281), .ZN(n474) );
  OR2X1 U10373 ( .IN1(n5474), .IN2(n3810), .Q(n9281) );
  AND2X1 U10374 ( .IN1(n4846), .IN2(n5964), .Q(n9279) );
  XNOR2X1 U10375 ( .IN1(n9282), .IN2(n9283), .Q(n5964) );
  XOR2X1 U10376 ( .IN1(n4179), .IN2(n5379), .Q(n9283) );
  XOR2X1 U10377 ( .IN1(n9284), .IN2(n4549), .Q(n9282) );
  XNOR2X1 U10378 ( .IN1(WX11131), .IN2(n8254), .Q(n9284) );
  OR2X1 U10379 ( .IN1(n9285), .IN2(n9286), .Q(WX11000) );
  OR2X1 U10380 ( .IN1(n9287), .IN2(n9288), .Q(n9286) );
  AND2X1 U10381 ( .IN1(n4898), .IN2(CRC_OUT_1_25), .Q(n9288) );
  AND2X1 U10382 ( .IN1(DATA_0_25), .IN2(n4923), .Q(n9287) );
  OR2X1 U10383 ( .IN1(n9289), .IN2(n9290), .Q(n9285) );
  AND2X1 U10384 ( .IN1(n473), .IN2(n4861), .Q(n9290) );
  INVX0 U10385 ( .INP(n9291), .ZN(n473) );
  OR2X1 U10386 ( .IN1(n5474), .IN2(n3811), .Q(n9291) );
  AND2X1 U10387 ( .IN1(n5973), .IN2(n4833), .Q(n9289) );
  XOR2X1 U10388 ( .IN1(n9292), .IN2(n9293), .Q(n5973) );
  XOR2X1 U10389 ( .IN1(n4180), .IN2(n5379), .Q(n9293) );
  XOR2X1 U10390 ( .IN1(n9294), .IN2(n4548), .Q(n9292) );
  XOR2X1 U10391 ( .IN1(WX11065), .IN2(test_so91), .Q(n9294) );
  OR2X1 U10392 ( .IN1(n9295), .IN2(n9296), .Q(WX10998) );
  OR2X1 U10393 ( .IN1(n9297), .IN2(n9298), .Q(n9296) );
  AND2X1 U10394 ( .IN1(n4898), .IN2(CRC_OUT_1_26), .Q(n9298) );
  AND2X1 U10395 ( .IN1(DATA_0_26), .IN2(n4923), .Q(n9297) );
  OR2X1 U10396 ( .IN1(n9299), .IN2(n9300), .Q(n9295) );
  AND2X1 U10397 ( .IN1(n472), .IN2(n4861), .Q(n9300) );
  INVX0 U10398 ( .INP(n9301), .ZN(n472) );
  OR2X1 U10399 ( .IN1(n5474), .IN2(n3812), .Q(n9301) );
  AND2X1 U10400 ( .IN1(n4846), .IN2(n5982), .Q(n9299) );
  XNOR2X1 U10401 ( .IN1(n9302), .IN2(n9303), .Q(n5982) );
  XOR2X1 U10402 ( .IN1(n4181), .IN2(n5379), .Q(n9303) );
  XOR2X1 U10403 ( .IN1(n9304), .IN2(n4547), .Q(n9302) );
  XNOR2X1 U10404 ( .IN1(WX11127), .IN2(n8257), .Q(n9304) );
  OR2X1 U10405 ( .IN1(n9305), .IN2(n9306), .Q(WX10996) );
  OR2X1 U10406 ( .IN1(n9307), .IN2(n9308), .Q(n9306) );
  AND2X1 U10407 ( .IN1(n4898), .IN2(CRC_OUT_1_27), .Q(n9308) );
  AND2X1 U10408 ( .IN1(DATA_0_27), .IN2(n4922), .Q(n9307) );
  OR2X1 U10409 ( .IN1(n9309), .IN2(n9310), .Q(n9305) );
  AND2X1 U10410 ( .IN1(n471), .IN2(n4861), .Q(n9310) );
  INVX0 U10411 ( .INP(n9311), .ZN(n471) );
  OR2X1 U10412 ( .IN1(n5474), .IN2(n3813), .Q(n9311) );
  AND2X1 U10413 ( .IN1(n4846), .IN2(n5991), .Q(n9309) );
  XNOR2X1 U10414 ( .IN1(n9312), .IN2(n9313), .Q(n5991) );
  XOR2X1 U10415 ( .IN1(n4182), .IN2(n5379), .Q(n9313) );
  XOR2X1 U10416 ( .IN1(n9314), .IN2(n4546), .Q(n9312) );
  XNOR2X1 U10417 ( .IN1(WX11125), .IN2(n8258), .Q(n9314) );
  OR2X1 U10418 ( .IN1(n9315), .IN2(n9316), .Q(WX10994) );
  OR2X1 U10419 ( .IN1(n9317), .IN2(n9318), .Q(n9316) );
  AND2X1 U10420 ( .IN1(n4898), .IN2(CRC_OUT_1_28), .Q(n9318) );
  AND2X1 U10421 ( .IN1(DATA_0_28), .IN2(n4921), .Q(n9317) );
  OR2X1 U10422 ( .IN1(n9319), .IN2(n9320), .Q(n9315) );
  AND2X1 U10423 ( .IN1(n470), .IN2(n4861), .Q(n9320) );
  INVX0 U10424 ( .INP(n9321), .ZN(n470) );
  OR2X1 U10425 ( .IN1(n5474), .IN2(n3814), .Q(n9321) );
  AND2X1 U10426 ( .IN1(n4846), .IN2(n6000), .Q(n9319) );
  XNOR2X1 U10427 ( .IN1(n9322), .IN2(n9323), .Q(n6000) );
  XOR2X1 U10428 ( .IN1(n4183), .IN2(n5379), .Q(n9323) );
  XOR2X1 U10429 ( .IN1(n9324), .IN2(n4545), .Q(n9322) );
  XNOR2X1 U10430 ( .IN1(WX11123), .IN2(n8259), .Q(n9324) );
  OR2X1 U10431 ( .IN1(n9325), .IN2(n9326), .Q(WX10992) );
  OR2X1 U10432 ( .IN1(n9327), .IN2(n9328), .Q(n9326) );
  AND2X1 U10433 ( .IN1(n4898), .IN2(CRC_OUT_1_29), .Q(n9328) );
  AND2X1 U10434 ( .IN1(DATA_0_29), .IN2(n4921), .Q(n9327) );
  OR2X1 U10435 ( .IN1(n9329), .IN2(n9330), .Q(n9325) );
  AND2X1 U10436 ( .IN1(n469), .IN2(n4861), .Q(n9330) );
  INVX0 U10437 ( .INP(n9331), .ZN(n469) );
  OR2X1 U10438 ( .IN1(n5474), .IN2(n3815), .Q(n9331) );
  AND2X1 U10439 ( .IN1(n4845), .IN2(n6009), .Q(n9329) );
  XNOR2X1 U10440 ( .IN1(n9332), .IN2(n9333), .Q(n6009) );
  XOR2X1 U10441 ( .IN1(n4184), .IN2(n5379), .Q(n9333) );
  XOR2X1 U10442 ( .IN1(n9334), .IN2(n4544), .Q(n9332) );
  XNOR2X1 U10443 ( .IN1(WX11121), .IN2(n8260), .Q(n9334) );
  OR2X1 U10444 ( .IN1(n9335), .IN2(n9336), .Q(WX10990) );
  OR2X1 U10445 ( .IN1(n9337), .IN2(n9338), .Q(n9336) );
  AND2X1 U10446 ( .IN1(n4898), .IN2(CRC_OUT_1_30), .Q(n9338) );
  AND2X1 U10447 ( .IN1(DATA_0_30), .IN2(n4921), .Q(n9337) );
  OR2X1 U10448 ( .IN1(n9339), .IN2(n9340), .Q(n9335) );
  AND2X1 U10449 ( .IN1(n468), .IN2(n4861), .Q(n9340) );
  AND2X1 U10450 ( .IN1(TM0), .IN2(TM1), .Q(n2148) );
  INVX0 U10451 ( .INP(n9341), .ZN(n468) );
  OR2X1 U10452 ( .IN1(n5483), .IN2(n3816), .Q(n9341) );
  AND2X1 U10453 ( .IN1(n4850), .IN2(n6018), .Q(n9339) );
  XNOR2X1 U10454 ( .IN1(n9342), .IN2(n9343), .Q(n6018) );
  XOR2X1 U10455 ( .IN1(n4185), .IN2(n5379), .Q(n9343) );
  XOR2X1 U10456 ( .IN1(n9344), .IN2(n4543), .Q(n9342) );
  XNOR2X1 U10457 ( .IN1(WX11119), .IN2(n8261), .Q(n9344) );
  OR2X1 U10458 ( .IN1(n9345), .IN2(n9346), .Q(WX10988) );
  OR2X1 U10459 ( .IN1(n9347), .IN2(n9348), .Q(n9346) );
  AND2X1 U10460 ( .IN1(n2245), .IN2(WX10829), .Q(n9348) );
  AND2X1 U10461 ( .IN1(test_so100), .IN2(n4888), .Q(n9347) );
  OR2X1 U10462 ( .IN1(n9349), .IN2(n9350), .Q(n9345) );
  AND2X1 U10463 ( .IN1(DATA_0_31), .IN2(n4919), .Q(n9350) );
  AND2X1 U10464 ( .IN1(n4839), .IN2(n6026), .Q(n9349) );
  XNOR2X1 U10465 ( .IN1(n9351), .IN2(n9352), .Q(n6026) );
  XOR2X1 U10466 ( .IN1(n4165), .IN2(n5379), .Q(n9352) );
  XOR2X1 U10467 ( .IN1(n9353), .IN2(n4542), .Q(n9351) );
  XNOR2X1 U10468 ( .IN1(WX11117), .IN2(n8262), .Q(n9353) );
  AND2X1 U10469 ( .IN1(TM1), .IN2(n9354), .Q(n5748) );
  AND2X1 U10470 ( .IN1(n530), .IN2(n5418), .Q(n9354) );
  INVX0 U10471 ( .INP(TM0), .ZN(n530) );
  AND2X1 U10472 ( .IN1(n4826), .IN2(n5418), .Q(WX10890) );
  AND2X1 U10473 ( .IN1(n9355), .IN2(n5418), .Q(WX10377) );
  XOR2X1 U10474 ( .IN1(test_so85), .IN2(DFF_1534_n1), .Q(n9355) );
  AND2X1 U10475 ( .IN1(n9356), .IN2(n5418), .Q(WX10375) );
  XOR2X1 U10476 ( .IN1(CRC_OUT_2_29), .IN2(n4568), .Q(n9356) );
  AND2X1 U10477 ( .IN1(n9357), .IN2(n5418), .Q(WX10373) );
  XOR2X1 U10478 ( .IN1(CRC_OUT_2_28), .IN2(n4569), .Q(n9357) );
  AND2X1 U10479 ( .IN1(n9358), .IN2(n5418), .Q(WX10371) );
  XOR2X1 U10480 ( .IN1(CRC_OUT_2_27), .IN2(n4570), .Q(n9358) );
  AND2X1 U10481 ( .IN1(n9359), .IN2(n5417), .Q(WX10369) );
  XOR2X1 U10482 ( .IN1(CRC_OUT_2_26), .IN2(n4571), .Q(n9359) );
  AND2X1 U10483 ( .IN1(n9360), .IN2(n5417), .Q(WX10367) );
  XOR2X1 U10484 ( .IN1(CRC_OUT_2_25), .IN2(n4572), .Q(n9360) );
  AND2X1 U10485 ( .IN1(n9361), .IN2(n5417), .Q(WX10365) );
  XOR2X1 U10486 ( .IN1(CRC_OUT_2_24), .IN2(n4573), .Q(n9361) );
  AND2X1 U10487 ( .IN1(n9362), .IN2(n5417), .Q(WX10363) );
  XOR2X1 U10488 ( .IN1(CRC_OUT_2_23), .IN2(n4574), .Q(n9362) );
  AND2X1 U10489 ( .IN1(n9363), .IN2(n5417), .Q(WX10361) );
  XOR2X1 U10490 ( .IN1(CRC_OUT_2_22), .IN2(n4575), .Q(n9363) );
  AND2X1 U10491 ( .IN1(n9364), .IN2(n5417), .Q(WX10359) );
  XOR2X1 U10492 ( .IN1(CRC_OUT_2_21), .IN2(n4576), .Q(n9364) );
  AND2X1 U10493 ( .IN1(n9365), .IN2(n5417), .Q(WX10357) );
  XOR2X1 U10494 ( .IN1(CRC_OUT_2_20), .IN2(n4577), .Q(n9365) );
  AND2X1 U10495 ( .IN1(n9366), .IN2(n5417), .Q(WX10355) );
  XOR2X1 U10496 ( .IN1(test_so88), .IN2(n4578), .Q(n9366) );
  AND2X1 U10497 ( .IN1(n9367), .IN2(n5417), .Q(WX10353) );
  XOR2X1 U10498 ( .IN1(CRC_OUT_2_18), .IN2(n4579), .Q(n9367) );
  AND2X1 U10499 ( .IN1(n9368), .IN2(n5416), .Q(WX10351) );
  XOR2X1 U10500 ( .IN1(CRC_OUT_2_17), .IN2(n4580), .Q(n9368) );
  AND2X1 U10501 ( .IN1(n9369), .IN2(n5416), .Q(WX10349) );
  XOR2X1 U10502 ( .IN1(CRC_OUT_2_16), .IN2(n4581), .Q(n9369) );
  AND2X1 U10503 ( .IN1(n9370), .IN2(n5416), .Q(WX10347) );
  XOR2X1 U10504 ( .IN1(DFF_1519_n1), .IN2(n9371), .Q(n9370) );
  XOR2X1 U10505 ( .IN1(n4516), .IN2(DFF_1535_n1), .Q(n9371) );
  AND2X1 U10506 ( .IN1(n9372), .IN2(n5416), .Q(WX10345) );
  XOR2X1 U10507 ( .IN1(CRC_OUT_2_14), .IN2(n4582), .Q(n9372) );
  AND2X1 U10508 ( .IN1(n9373), .IN2(n5416), .Q(WX10343) );
  XOR2X1 U10509 ( .IN1(test_so86), .IN2(DFF_1517_n1), .Q(n9373) );
  AND2X1 U10510 ( .IN1(n9374), .IN2(n5416), .Q(WX10341) );
  XOR2X1 U10511 ( .IN1(CRC_OUT_2_12), .IN2(n4583), .Q(n9374) );
  AND2X1 U10512 ( .IN1(n9375), .IN2(n5416), .Q(WX10339) );
  XOR2X1 U10513 ( .IN1(CRC_OUT_2_11), .IN2(n4584), .Q(n9375) );
  AND2X1 U10514 ( .IN1(n9376), .IN2(n5416), .Q(WX10337) );
  XOR2X1 U10515 ( .IN1(DFF_1514_n1), .IN2(n9377), .Q(n9376) );
  XOR2X1 U10516 ( .IN1(n4517), .IN2(DFF_1535_n1), .Q(n9377) );
  AND2X1 U10517 ( .IN1(n9378), .IN2(n5416), .Q(WX10335) );
  XOR2X1 U10518 ( .IN1(CRC_OUT_2_9), .IN2(n4585), .Q(n9378) );
  AND2X1 U10519 ( .IN1(n9379), .IN2(n5415), .Q(WX10333) );
  XOR2X1 U10520 ( .IN1(CRC_OUT_2_8), .IN2(n4586), .Q(n9379) );
  AND2X1 U10521 ( .IN1(n9380), .IN2(n5415), .Q(WX10331) );
  XOR2X1 U10522 ( .IN1(CRC_OUT_2_7), .IN2(n4587), .Q(n9380) );
  AND2X1 U10523 ( .IN1(n9381), .IN2(n5415), .Q(WX10329) );
  XOR2X1 U10524 ( .IN1(CRC_OUT_2_6), .IN2(n4588), .Q(n9381) );
  AND2X1 U10525 ( .IN1(n9382), .IN2(n5415), .Q(WX10327) );
  XOR2X1 U10526 ( .IN1(CRC_OUT_2_5), .IN2(n4589), .Q(n9382) );
  AND2X1 U10527 ( .IN1(n9383), .IN2(n5415), .Q(WX10325) );
  XOR2X1 U10528 ( .IN1(CRC_OUT_2_4), .IN2(n4590), .Q(n9383) );
  AND2X1 U10529 ( .IN1(n9384), .IN2(n5415), .Q(WX10323) );
  XOR2X1 U10530 ( .IN1(DFF_1507_n1), .IN2(n9385), .Q(n9384) );
  XOR2X1 U10531 ( .IN1(n4518), .IN2(DFF_1535_n1), .Q(n9385) );
  AND2X1 U10532 ( .IN1(n9386), .IN2(n5415), .Q(WX10321) );
  XOR2X1 U10533 ( .IN1(test_so87), .IN2(n4591), .Q(n9386) );
  AND2X1 U10534 ( .IN1(n9387), .IN2(n5425), .Q(WX10319) );
  XOR2X1 U10535 ( .IN1(CRC_OUT_2_1), .IN2(n4592), .Q(n9387) );
  AND2X1 U10536 ( .IN1(n9388), .IN2(n5401), .Q(WX10317) );
  XOR2X1 U10537 ( .IN1(CRC_OUT_2_0), .IN2(n4593), .Q(n9388) );
  AND2X1 U10538 ( .IN1(n9389), .IN2(n5415), .Q(WX10315) );
  XOR2X1 U10539 ( .IN1(n4535), .IN2(CRC_OUT_2_31), .Q(n9389) );
  XOR2X1 U10540 ( .IN1(n9390), .IN2(n6876), .Q(DATA_9_9) );
  XNOR2X1 U10541 ( .IN1(n9391), .IN2(n9392), .Q(n6876) );
  XOR2X1 U10542 ( .IN1(n3485), .IN2(TM0), .Q(n9392) );
  XOR2X1 U10543 ( .IN1(n9393), .IN2(n4772), .Q(n9391) );
  XOR2X1 U10544 ( .IN1(WX753), .IN2(n9765), .Q(n9393) );
  AND2X1 U10545 ( .IN1(TM0), .IN2(WX529), .Q(n9390) );
  XOR2X1 U10546 ( .IN1(n9394), .IN2(n6868), .Q(DATA_9_8) );
  XNOR2X1 U10547 ( .IN1(n9395), .IN2(n9396), .Q(n6868) );
  XOR2X1 U10548 ( .IN1(n3483), .IN2(TM0), .Q(n9396) );
  XOR2X1 U10549 ( .IN1(n9397), .IN2(n4777), .Q(n9395) );
  XOR2X1 U10550 ( .IN1(WX819), .IN2(n9766), .Q(n9397) );
  AND2X1 U10551 ( .IN1(TM0), .IN2(WX531), .Q(n9394) );
  XOR2X1 U10552 ( .IN1(n9398), .IN2(n6860), .Q(DATA_9_7) );
  XNOR2X1 U10553 ( .IN1(n9399), .IN2(n9400), .Q(n6860) );
  XOR2X1 U10554 ( .IN1(n3481), .IN2(TM0), .Q(n9400) );
  XOR2X1 U10555 ( .IN1(n9401), .IN2(n4792), .Q(n9399) );
  XOR2X1 U10556 ( .IN1(WX821), .IN2(n4793), .Q(n9401) );
  AND2X1 U10557 ( .IN1(TM0), .IN2(WX533), .Q(n9398) );
  XOR2X1 U10558 ( .IN1(n6852), .IN2(n9402), .Q(DATA_9_6) );
  AND2X1 U10559 ( .IN1(TM0), .IN2(WX535), .Q(n9402) );
  XOR2X1 U10560 ( .IN1(n9403), .IN2(n9404), .Q(n6852) );
  XOR2X1 U10561 ( .IN1(n3479), .IN2(TM0), .Q(n9404) );
  XOR2X1 U10562 ( .IN1(n9405), .IN2(n4786), .Q(n9403) );
  XOR2X1 U10563 ( .IN1(WX823), .IN2(test_so5), .Q(n9405) );
  XOR2X1 U10564 ( .IN1(n9406), .IN2(n6844), .Q(DATA_9_5) );
  XNOR2X1 U10565 ( .IN1(n9407), .IN2(n9408), .Q(n6844) );
  XOR2X1 U10566 ( .IN1(n3477), .IN2(TM0), .Q(n9408) );
  XOR2X1 U10567 ( .IN1(n9409), .IN2(n4778), .Q(n9407) );
  XOR2X1 U10568 ( .IN1(WX825), .IN2(n9767), .Q(n9409) );
  AND2X1 U10569 ( .IN1(TM0), .IN2(WX537), .Q(n9406) );
  XOR2X1 U10570 ( .IN1(n9410), .IN2(n6836), .Q(DATA_9_4) );
  XNOR2X1 U10571 ( .IN1(n9411), .IN2(n9412), .Q(n6836) );
  XOR2X1 U10572 ( .IN1(n3475), .IN2(TM0), .Q(n9412) );
  XOR2X1 U10573 ( .IN1(n9413), .IN2(n4779), .Q(n9411) );
  XOR2X1 U10574 ( .IN1(WX827), .IN2(n9768), .Q(n9413) );
  AND2X1 U10575 ( .IN1(TM0), .IN2(WX539), .Q(n9410) );
  XOR2X1 U10576 ( .IN1(n9414), .IN2(n7086), .Q(DATA_9_31) );
  XNOR2X1 U10577 ( .IN1(n9415), .IN2(n9416), .Q(n7086) );
  XOR2X1 U10578 ( .IN1(n3529), .IN2(n5379), .Q(n9416) );
  XOR2X1 U10579 ( .IN1(n9417), .IN2(n4789), .Q(n9415) );
  XOR2X1 U10580 ( .IN1(WX709), .IN2(n9769), .Q(n9417) );
  AND2X1 U10581 ( .IN1(TM0), .IN2(WX485), .Q(n9414) );
  XOR2X1 U10582 ( .IN1(n9418), .IN2(n7066), .Q(DATA_9_30) );
  XNOR2X1 U10583 ( .IN1(n9419), .IN2(n9420), .Q(n7066) );
  XOR2X1 U10584 ( .IN1(n3527), .IN2(n5379), .Q(n9420) );
  XOR2X1 U10585 ( .IN1(n9421), .IN2(n4754), .Q(n9419) );
  XOR2X1 U10586 ( .IN1(WX775), .IN2(n4755), .Q(n9421) );
  AND2X1 U10587 ( .IN1(TM0), .IN2(WX487), .Q(n9418) );
  XOR2X1 U10588 ( .IN1(n9422), .IN2(n6828), .Q(DATA_9_3) );
  XNOR2X1 U10589 ( .IN1(n9423), .IN2(n9424), .Q(n6828) );
  XOR2X1 U10590 ( .IN1(n3473), .IN2(TM0), .Q(n9424) );
  XOR2X1 U10591 ( .IN1(n9425), .IN2(n4756), .Q(n9423) );
  XOR2X1 U10592 ( .IN1(WX829), .IN2(n9770), .Q(n9425) );
  AND2X1 U10593 ( .IN1(TM0), .IN2(WX541), .Q(n9422) );
  XOR2X1 U10594 ( .IN1(n9426), .IN2(n7047), .Q(DATA_9_29) );
  XNOR2X1 U10595 ( .IN1(n9427), .IN2(n9428), .Q(n7047) );
  XOR2X1 U10596 ( .IN1(n3525), .IN2(n5379), .Q(n9428) );
  XOR2X1 U10597 ( .IN1(n9429), .IN2(n4758), .Q(n9427) );
  XOR2X1 U10598 ( .IN1(WX777), .IN2(n9771), .Q(n9429) );
  AND2X1 U10599 ( .IN1(TM0), .IN2(WX489), .Q(n9426) );
  XOR2X1 U10600 ( .IN1(n7028), .IN2(n9430), .Q(DATA_9_28) );
  AND2X1 U10601 ( .IN1(TM0), .IN2(WX491), .Q(n9430) );
  XOR2X1 U10602 ( .IN1(n9431), .IN2(n9432), .Q(n7028) );
  XOR2X1 U10603 ( .IN1(n4762), .IN2(n5379), .Q(n9432) );
  XOR2X1 U10604 ( .IN1(n9433), .IN2(n4763), .Q(n9431) );
  XOR2X1 U10605 ( .IN1(WX779), .IN2(test_so2), .Q(n9433) );
  XOR2X1 U10606 ( .IN1(n9434), .IN2(n7020), .Q(DATA_9_27) );
  XNOR2X1 U10607 ( .IN1(n9435), .IN2(n9436), .Q(n7020) );
  XOR2X1 U10608 ( .IN1(n3521), .IN2(n5378), .Q(n9436) );
  XOR2X1 U10609 ( .IN1(n9437), .IN2(n4765), .Q(n9435) );
  XOR2X1 U10610 ( .IN1(WX781), .IN2(n9772), .Q(n9437) );
  AND2X1 U10611 ( .IN1(TM0), .IN2(WX493), .Q(n9434) );
  XOR2X1 U10612 ( .IN1(n9438), .IN2(n7012), .Q(DATA_9_26) );
  XNOR2X1 U10613 ( .IN1(n9439), .IN2(n9440), .Q(n7012) );
  XOR2X1 U10614 ( .IN1(n3519), .IN2(n5378), .Q(n9440) );
  XOR2X1 U10615 ( .IN1(n9441), .IN2(n4766), .Q(n9439) );
  XOR2X1 U10616 ( .IN1(WX783), .IN2(n9773), .Q(n9441) );
  AND2X1 U10617 ( .IN1(TM0), .IN2(WX495), .Q(n9438) );
  XOR2X1 U10618 ( .IN1(n9442), .IN2(n7004), .Q(DATA_9_25) );
  XNOR2X1 U10619 ( .IN1(n9443), .IN2(n9444), .Q(n7004) );
  XOR2X1 U10620 ( .IN1(n3517), .IN2(n5378), .Q(n9444) );
  XOR2X1 U10621 ( .IN1(n9445), .IN2(n4770), .Q(n9443) );
  XOR2X1 U10622 ( .IN1(WX785), .IN2(n9774), .Q(n9445) );
  AND2X1 U10623 ( .IN1(TM0), .IN2(WX497), .Q(n9442) );
  XOR2X1 U10624 ( .IN1(n6996), .IN2(n9446), .Q(DATA_9_24) );
  AND2X1 U10625 ( .IN1(TM0), .IN2(WX499), .Q(n9446) );
  XOR2X1 U10626 ( .IN1(n9447), .IN2(n9448), .Q(n6996) );
  XOR2X1 U10627 ( .IN1(n3515), .IN2(n5378), .Q(n9448) );
  XOR2X1 U10628 ( .IN1(n9449), .IN2(n4773), .Q(n9447) );
  XOR2X1 U10629 ( .IN1(WX787), .IN2(test_so4), .Q(n9449) );
  XOR2X1 U10630 ( .IN1(n9450), .IN2(n6988), .Q(DATA_9_23) );
  XNOR2X1 U10631 ( .IN1(n9451), .IN2(n9452), .Q(n6988) );
  XOR2X1 U10632 ( .IN1(n3513), .IN2(n5378), .Q(n9452) );
  XOR2X1 U10633 ( .IN1(n9453), .IN2(n4775), .Q(n9451) );
  XOR2X1 U10634 ( .IN1(WX789), .IN2(n9775), .Q(n9453) );
  AND2X1 U10635 ( .IN1(TM0), .IN2(WX501), .Q(n9450) );
  XOR2X1 U10636 ( .IN1(n9454), .IN2(n6980), .Q(DATA_9_22) );
  XNOR2X1 U10637 ( .IN1(n9455), .IN2(n9456), .Q(n6980) );
  XOR2X1 U10638 ( .IN1(n3511), .IN2(n5378), .Q(n9456) );
  XOR2X1 U10639 ( .IN1(n9457), .IN2(n4780), .Q(n9455) );
  XOR2X1 U10640 ( .IN1(WX791), .IN2(n4781), .Q(n9457) );
  AND2X1 U10641 ( .IN1(TM0), .IN2(WX503), .Q(n9454) );
  XOR2X1 U10642 ( .IN1(n9458), .IN2(n6972), .Q(DATA_9_21) );
  XNOR2X1 U10643 ( .IN1(n9459), .IN2(n9460), .Q(n6972) );
  XOR2X1 U10644 ( .IN1(n3509), .IN2(n5378), .Q(n9460) );
  XOR2X1 U10645 ( .IN1(n9461), .IN2(n4784), .Q(n9459) );
  XOR2X1 U10646 ( .IN1(WX793), .IN2(n4785), .Q(n9461) );
  AND2X1 U10647 ( .IN1(TM0), .IN2(WX505), .Q(n9458) );
  XOR2X1 U10648 ( .IN1(n6964), .IN2(n9462), .Q(DATA_9_20) );
  AND2X1 U10649 ( .IN1(TM0), .IN2(WX507), .Q(n9462) );
  XOR2X1 U10650 ( .IN1(n9463), .IN2(n9464), .Q(n6964) );
  XOR2X1 U10651 ( .IN1(n3507), .IN2(n5378), .Q(n9464) );
  XOR2X1 U10652 ( .IN1(n9465), .IN2(n4787), .Q(n9463) );
  XOR2X1 U10653 ( .IN1(WX731), .IN2(test_so6), .Q(n9465) );
  XOR2X1 U10654 ( .IN1(n6820), .IN2(n9466), .Q(DATA_9_2) );
  AND2X1 U10655 ( .IN1(TM0), .IN2(WX543), .Q(n9466) );
  XOR2X1 U10656 ( .IN1(n9467), .IN2(n9468), .Q(n6820) );
  XOR2X1 U10657 ( .IN1(n3471), .IN2(TM0), .Q(n9468) );
  XOR2X1 U10658 ( .IN1(n9469), .IN2(n4791), .Q(n9467) );
  XOR2X1 U10659 ( .IN1(WX767), .IN2(test_so7), .Q(n9469) );
  XOR2X1 U10660 ( .IN1(n9470), .IN2(n6956), .Q(DATA_9_19) );
  XNOR2X1 U10661 ( .IN1(n9471), .IN2(n9472), .Q(n6956) );
  XOR2X1 U10662 ( .IN1(n3505), .IN2(n5378), .Q(n9472) );
  XOR2X1 U10663 ( .IN1(n9473), .IN2(n4757), .Q(n9471) );
  XOR2X1 U10664 ( .IN1(WX797), .IN2(n9776), .Q(n9473) );
  AND2X1 U10665 ( .IN1(TM0), .IN2(WX509), .Q(n9470) );
  XOR2X1 U10666 ( .IN1(n9474), .IN2(n6948), .Q(DATA_9_18) );
  XNOR2X1 U10667 ( .IN1(n9475), .IN2(n9476), .Q(n6948) );
  XOR2X1 U10668 ( .IN1(n3503), .IN2(n5378), .Q(n9476) );
  XOR2X1 U10669 ( .IN1(n9477), .IN2(n4764), .Q(n9475) );
  XOR2X1 U10670 ( .IN1(WX799), .IN2(n9777), .Q(n9477) );
  AND2X1 U10671 ( .IN1(TM0), .IN2(WX511), .Q(n9474) );
  XOR2X1 U10672 ( .IN1(n9478), .IN2(n6940), .Q(DATA_9_17) );
  XNOR2X1 U10673 ( .IN1(n9479), .IN2(n9480), .Q(n6940) );
  XOR2X1 U10674 ( .IN1(n3501), .IN2(n5378), .Q(n9480) );
  XOR2X1 U10675 ( .IN1(n9481), .IN2(n4769), .Q(n9479) );
  XOR2X1 U10676 ( .IN1(WX801), .IN2(n9778), .Q(n9481) );
  AND2X1 U10677 ( .IN1(TM0), .IN2(WX513), .Q(n9478) );
  XOR2X1 U10678 ( .IN1(n6932), .IN2(n9482), .Q(DATA_9_16) );
  AND2X1 U10679 ( .IN1(TM0), .IN2(WX515), .Q(n9482) );
  XOR2X1 U10680 ( .IN1(n9483), .IN2(n9484), .Q(n6932) );
  XOR2X1 U10681 ( .IN1(n3499), .IN2(n5384), .Q(n9484) );
  XOR2X1 U10682 ( .IN1(n9485), .IN2(n4776), .Q(n9483) );
  XOR2X1 U10683 ( .IN1(WX739), .IN2(test_so8), .Q(n9485) );
  XOR2X1 U10684 ( .IN1(n9486), .IN2(n6924), .Q(DATA_9_15) );
  XNOR2X1 U10685 ( .IN1(n9487), .IN2(n9488), .Q(n6924) );
  XOR2X1 U10686 ( .IN1(n3497), .IN2(TM0), .Q(n9488) );
  XOR2X1 U10687 ( .IN1(n9489), .IN2(n4782), .Q(n9487) );
  XOR2X1 U10688 ( .IN1(WX805), .IN2(n4783), .Q(n9489) );
  AND2X1 U10689 ( .IN1(TM0), .IN2(WX517), .Q(n9486) );
  XOR2X1 U10690 ( .IN1(n9490), .IN2(n6916), .Q(DATA_9_14) );
  XNOR2X1 U10691 ( .IN1(n9491), .IN2(n9492), .Q(n6916) );
  XOR2X1 U10692 ( .IN1(n3495), .IN2(TM0), .Q(n9492) );
  XOR2X1 U10693 ( .IN1(n9493), .IN2(n4790), .Q(n9491) );
  XOR2X1 U10694 ( .IN1(WX807), .IN2(n9779), .Q(n9493) );
  AND2X1 U10695 ( .IN1(test_so1), .IN2(TM0), .Q(n9490) );
  XOR2X1 U10696 ( .IN1(n9494), .IN2(n6908), .Q(DATA_9_13) );
  XNOR2X1 U10697 ( .IN1(n9495), .IN2(n9496), .Q(n6908) );
  XOR2X1 U10698 ( .IN1(n3493), .IN2(TM0), .Q(n9496) );
  XOR2X1 U10699 ( .IN1(n9497), .IN2(n4759), .Q(n9495) );
  XOR2X1 U10700 ( .IN1(WX809), .IN2(n9780), .Q(n9497) );
  AND2X1 U10701 ( .IN1(TM0), .IN2(WX521), .Q(n9494) );
  XOR2X1 U10702 ( .IN1(n9498), .IN2(n6900), .Q(DATA_9_12) );
  XNOR2X1 U10703 ( .IN1(n9499), .IN2(n9500), .Q(n6900) );
  XOR2X1 U10704 ( .IN1(n3491), .IN2(TM0), .Q(n9500) );
  XOR2X1 U10705 ( .IN1(n9501), .IN2(n4771), .Q(n9499) );
  XOR2X1 U10706 ( .IN1(WX811), .IN2(n9781), .Q(n9501) );
  AND2X1 U10707 ( .IN1(TM0), .IN2(WX523), .Q(n9498) );
  XOR2X1 U10708 ( .IN1(n9502), .IN2(n6892), .Q(DATA_9_11) );
  XNOR2X1 U10709 ( .IN1(n9503), .IN2(n9504), .Q(n6892) );
  XOR2X1 U10710 ( .IN1(n3489), .IN2(TM0), .Q(n9504) );
  XOR2X1 U10711 ( .IN1(n9505), .IN2(n4794), .Q(n9503) );
  XOR2X1 U10712 ( .IN1(WX813), .IN2(n9782), .Q(n9505) );
  AND2X1 U10713 ( .IN1(TM0), .IN2(WX525), .Q(n9502) );
  XOR2X1 U10714 ( .IN1(n6884), .IN2(n9506), .Q(DATA_9_10) );
  AND2X1 U10715 ( .IN1(TM0), .IN2(WX527), .Q(n9506) );
  XOR2X1 U10716 ( .IN1(n9507), .IN2(n9508), .Q(n6884) );
  XOR2X1 U10717 ( .IN1(n4767), .IN2(TM0), .Q(n9508) );
  XOR2X1 U10718 ( .IN1(n9509), .IN2(n4768), .Q(n9507) );
  XOR2X1 U10719 ( .IN1(WX815), .IN2(test_so3), .Q(n9509) );
  XOR2X1 U10720 ( .IN1(n9510), .IN2(n6812), .Q(DATA_9_1) );
  XNOR2X1 U10721 ( .IN1(n9511), .IN2(n9512), .Q(n6812) );
  XOR2X1 U10722 ( .IN1(n3469), .IN2(TM0), .Q(n9512) );
  XOR2X1 U10723 ( .IN1(n9513), .IN2(n4760), .Q(n9511) );
  XOR2X1 U10724 ( .IN1(WX833), .IN2(n9783), .Q(n9513) );
  AND2X1 U10725 ( .IN1(TM0), .IN2(WX545), .Q(n9510) );
  XOR2X1 U10726 ( .IN1(n9514), .IN2(n6804), .Q(DATA_9_0) );
  XNOR2X1 U10727 ( .IN1(n9515), .IN2(n9516), .Q(n6804) );
  XOR2X1 U10728 ( .IN1(n3467), .IN2(TM0), .Q(n9516) );
  XOR2X1 U10729 ( .IN1(n9517), .IN2(n4795), .Q(n9515) );
  XOR2X1 U10730 ( .IN1(WX835), .IN2(n4796), .Q(n9517) );
  AND2X1 U10731 ( .IN1(TM0), .IN2(WX547), .Q(n9514) );
  AND2X1 U3558_U2 ( .IN1(n4884), .IN2(U3558_n1), .Q(n2245) );
  INVX0 U3558_U1 ( .INP(n5498), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(TM0), .ZN(U3871_n1) );
  AND2X1 U3871_U1 ( .IN1(n3278), .IN2(U3871_n1), .Q(n2153) );
  INVX0 U3991_U2 ( .INP(n530), .ZN(U3991_n1) );
  AND2X1 U3991_U1 ( .IN1(n3278), .IN2(U3991_n1), .Q(n2152) );
  AND2X1 U5716_U2 ( .IN1(WX547), .IN2(U5716_n1), .Q(WX544) );
  INVX0 U5716_U1 ( .INP(n5502), .ZN(U5716_n1) );
  AND2X1 U5717_U2 ( .IN1(WX545), .IN2(U5717_n1), .Q(WX542) );
  INVX0 U5717_U1 ( .INP(n5487), .ZN(U5717_n1) );
  AND2X1 U5718_U2 ( .IN1(WX543), .IN2(U5718_n1), .Q(WX540) );
  INVX0 U5718_U1 ( .INP(n5522), .ZN(U5718_n1) );
  AND2X1 U5719_U2 ( .IN1(WX541), .IN2(U5719_n1), .Q(WX538) );
  INVX0 U5719_U1 ( .INP(n5517), .ZN(U5719_n1) );
  AND2X1 U5720_U2 ( .IN1(WX539), .IN2(U5720_n1), .Q(WX536) );
  INVX0 U5720_U1 ( .INP(n5512), .ZN(U5720_n1) );
  AND2X1 U5721_U2 ( .IN1(WX537), .IN2(U5721_n1), .Q(WX534) );
  INVX0 U5721_U1 ( .INP(n5512), .ZN(U5721_n1) );
  AND2X1 U5722_U2 ( .IN1(WX535), .IN2(U5722_n1), .Q(WX532) );
  INVX0 U5722_U1 ( .INP(n5512), .ZN(U5722_n1) );
  AND2X1 U5723_U2 ( .IN1(WX533), .IN2(U5723_n1), .Q(WX530) );
  INVX0 U5723_U1 ( .INP(n5512), .ZN(U5723_n1) );
  AND2X1 U5724_U2 ( .IN1(WX531), .IN2(U5724_n1), .Q(WX528) );
  INVX0 U5724_U1 ( .INP(n5512), .ZN(U5724_n1) );
  AND2X1 U5725_U2 ( .IN1(WX529), .IN2(U5725_n1), .Q(WX526) );
  INVX0 U5725_U1 ( .INP(n5512), .ZN(U5725_n1) );
  AND2X1 U5726_U2 ( .IN1(WX527), .IN2(U5726_n1), .Q(WX524) );
  INVX0 U5726_U1 ( .INP(n5512), .ZN(U5726_n1) );
  AND2X1 U5727_U2 ( .IN1(WX525), .IN2(U5727_n1), .Q(WX522) );
  INVX0 U5727_U1 ( .INP(n5512), .ZN(U5727_n1) );
  AND2X1 U5728_U2 ( .IN1(WX523), .IN2(U5728_n1), .Q(WX520) );
  INVX0 U5728_U1 ( .INP(n5512), .ZN(U5728_n1) );
  AND2X1 U5729_U2 ( .IN1(WX521), .IN2(U5729_n1), .Q(WX518) );
  INVX0 U5729_U1 ( .INP(n5512), .ZN(U5729_n1) );
  AND2X1 U5730_U2 ( .IN1(test_so1), .IN2(U5730_n1), .Q(WX516) );
  INVX0 U5730_U1 ( .INP(n5513), .ZN(U5730_n1) );
  AND2X1 U5731_U2 ( .IN1(WX517), .IN2(U5731_n1), .Q(WX514) );
  INVX0 U5731_U1 ( .INP(n5513), .ZN(U5731_n1) );
  AND2X1 U5732_U2 ( .IN1(WX515), .IN2(U5732_n1), .Q(WX512) );
  INVX0 U5732_U1 ( .INP(n5513), .ZN(U5732_n1) );
  AND2X1 U5733_U2 ( .IN1(WX513), .IN2(U5733_n1), .Q(WX510) );
  INVX0 U5733_U1 ( .INP(n5513), .ZN(U5733_n1) );
  AND2X1 U5734_U2 ( .IN1(WX511), .IN2(U5734_n1), .Q(WX508) );
  INVX0 U5734_U1 ( .INP(n5513), .ZN(U5734_n1) );
  AND2X1 U5735_U2 ( .IN1(WX509), .IN2(U5735_n1), .Q(WX506) );
  INVX0 U5735_U1 ( .INP(n5513), .ZN(U5735_n1) );
  AND2X1 U5736_U2 ( .IN1(WX507), .IN2(U5736_n1), .Q(WX504) );
  INVX0 U5736_U1 ( .INP(n5513), .ZN(U5736_n1) );
  AND2X1 U5737_U2 ( .IN1(WX505), .IN2(U5737_n1), .Q(WX502) );
  INVX0 U5737_U1 ( .INP(n5513), .ZN(U5737_n1) );
  AND2X1 U5738_U2 ( .IN1(WX503), .IN2(U5738_n1), .Q(WX500) );
  INVX0 U5738_U1 ( .INP(n5513), .ZN(U5738_n1) );
  AND2X1 U5739_U2 ( .IN1(WX501), .IN2(U5739_n1), .Q(WX498) );
  INVX0 U5739_U1 ( .INP(n5513), .ZN(U5739_n1) );
  AND2X1 U5740_U2 ( .IN1(WX499), .IN2(U5740_n1), .Q(WX496) );
  INVX0 U5740_U1 ( .INP(n5513), .ZN(U5740_n1) );
  AND2X1 U5741_U2 ( .IN1(WX497), .IN2(U5741_n1), .Q(WX494) );
  INVX0 U5741_U1 ( .INP(n5513), .ZN(U5741_n1) );
  AND2X1 U5742_U2 ( .IN1(WX495), .IN2(U5742_n1), .Q(WX492) );
  INVX0 U5742_U1 ( .INP(n5513), .ZN(U5742_n1) );
  AND2X1 U5743_U2 ( .IN1(WX493), .IN2(U5743_n1), .Q(WX490) );
  INVX0 U5743_U1 ( .INP(n5513), .ZN(U5743_n1) );
  AND2X1 U5744_U2 ( .IN1(WX491), .IN2(U5744_n1), .Q(WX488) );
  INVX0 U5744_U1 ( .INP(n5514), .ZN(U5744_n1) );
  AND2X1 U5745_U2 ( .IN1(WX489), .IN2(U5745_n1), .Q(WX486) );
  INVX0 U5745_U1 ( .INP(n5514), .ZN(U5745_n1) );
  AND2X1 U5746_U2 ( .IN1(WX487), .IN2(U5746_n1), .Q(WX484) );
  INVX0 U5746_U1 ( .INP(n5514), .ZN(U5746_n1) );
  AND2X1 U5747_U2 ( .IN1(WX5939), .IN2(U5747_n1), .Q(WX6002) );
  INVX0 U5747_U1 ( .INP(n5514), .ZN(U5747_n1) );
  AND2X1 U5748_U2 ( .IN1(test_so49), .IN2(U5748_n1), .Q(WX6000) );
  INVX0 U5748_U1 ( .INP(n5514), .ZN(U5748_n1) );
  AND2X1 U5749_U2 ( .IN1(WX5935), .IN2(U5749_n1), .Q(WX5998) );
  INVX0 U5749_U1 ( .INP(n5514), .ZN(U5749_n1) );
  AND2X1 U5750_U2 ( .IN1(WX5933), .IN2(U5750_n1), .Q(WX5996) );
  INVX0 U5750_U1 ( .INP(n5514), .ZN(U5750_n1) );
  AND2X1 U5751_U2 ( .IN1(WX5931), .IN2(U5751_n1), .Q(WX5994) );
  INVX0 U5751_U1 ( .INP(n5514), .ZN(U5751_n1) );
  AND2X1 U5752_U2 ( .IN1(WX3269), .IN2(U5752_n1), .Q(WX3332) );
  INVX0 U5752_U1 ( .INP(n5514), .ZN(U5752_n1) );
  AND2X1 U5753_U2 ( .IN1(WX3265), .IN2(U5753_n1), .Q(WX3328) );
  INVX0 U5753_U1 ( .INP(n5514), .ZN(U5753_n1) );
  AND2X1 U5754_U2 ( .IN1(WX3263), .IN2(U5754_n1), .Q(WX3326) );
  INVX0 U5754_U1 ( .INP(n5514), .ZN(U5754_n1) );
  AND2X1 U5755_U2 ( .IN1(WX11179), .IN2(U5755_n1), .Q(WX11242) );
  INVX0 U5755_U1 ( .INP(n5514), .ZN(U5755_n1) );
  AND2X1 U5756_U2 ( .IN1(WX11177), .IN2(U5756_n1), .Q(WX11240) );
  INVX0 U5756_U1 ( .INP(n5514), .ZN(U5756_n1) );
  AND2X1 U5757_U2 ( .IN1(WX11175), .IN2(U5757_n1), .Q(WX11238) );
  INVX0 U5757_U1 ( .INP(n5514), .ZN(U5757_n1) );
  AND2X1 U5758_U2 ( .IN1(WX11173), .IN2(U5758_n1), .Q(WX11236) );
  INVX0 U5758_U1 ( .INP(n5515), .ZN(U5758_n1) );
  AND2X1 U5759_U2 ( .IN1(test_so96), .IN2(U5759_n1), .Q(WX11234) );
  INVX0 U5759_U1 ( .INP(n5515), .ZN(U5759_n1) );
  AND2X1 U5760_U2 ( .IN1(WX11169), .IN2(U5760_n1), .Q(WX11232) );
  INVX0 U5760_U1 ( .INP(n5515), .ZN(U5760_n1) );
  AND2X1 U5761_U2 ( .IN1(WX11167), .IN2(U5761_n1), .Q(WX11230) );
  INVX0 U5761_U1 ( .INP(n5515), .ZN(U5761_n1) );
  AND2X1 U5762_U2 ( .IN1(WX11165), .IN2(U5762_n1), .Q(WX11228) );
  INVX0 U5762_U1 ( .INP(n5515), .ZN(U5762_n1) );
  AND2X1 U5763_U2 ( .IN1(WX11163), .IN2(U5763_n1), .Q(WX11226) );
  INVX0 U5763_U1 ( .INP(n5515), .ZN(U5763_n1) );
  AND2X1 U5764_U2 ( .IN1(WX11161), .IN2(U5764_n1), .Q(WX11224) );
  INVX0 U5764_U1 ( .INP(n5515), .ZN(U5764_n1) );
  AND2X1 U5765_U2 ( .IN1(WX11159), .IN2(U5765_n1), .Q(WX11222) );
  INVX0 U5765_U1 ( .INP(n5515), .ZN(U5765_n1) );
  AND2X1 U5766_U2 ( .IN1(WX11157), .IN2(U5766_n1), .Q(WX11220) );
  INVX0 U5766_U1 ( .INP(n5515), .ZN(U5766_n1) );
  AND2X1 U5767_U2 ( .IN1(WX11155), .IN2(U5767_n1), .Q(WX11218) );
  INVX0 U5767_U1 ( .INP(n5515), .ZN(U5767_n1) );
  AND2X1 U5768_U2 ( .IN1(WX11153), .IN2(U5768_n1), .Q(WX11216) );
  INVX0 U5768_U1 ( .INP(n5515), .ZN(U5768_n1) );
  AND2X1 U5769_U2 ( .IN1(WX11151), .IN2(U5769_n1), .Q(WX11214) );
  INVX0 U5769_U1 ( .INP(n5515), .ZN(U5769_n1) );
  AND2X1 U5770_U2 ( .IN1(WX11149), .IN2(U5770_n1), .Q(WX11212) );
  INVX0 U5770_U1 ( .INP(n5515), .ZN(U5770_n1) );
  AND2X1 U5771_U2 ( .IN1(WX11147), .IN2(U5771_n1), .Q(WX11210) );
  INVX0 U5771_U1 ( .INP(n5515), .ZN(U5771_n1) );
  AND2X1 U5772_U2 ( .IN1(WX11145), .IN2(U5772_n1), .Q(WX11208) );
  INVX0 U5772_U1 ( .INP(n5516), .ZN(U5772_n1) );
  AND2X1 U5773_U2 ( .IN1(WX11143), .IN2(U5773_n1), .Q(WX11206) );
  INVX0 U5773_U1 ( .INP(n5516), .ZN(U5773_n1) );
  AND2X1 U5774_U2 ( .IN1(WX11141), .IN2(U5774_n1), .Q(WX11204) );
  INVX0 U5774_U1 ( .INP(n5516), .ZN(U5774_n1) );
  AND2X1 U5775_U2 ( .IN1(WX11139), .IN2(U5775_n1), .Q(WX11202) );
  INVX0 U5775_U1 ( .INP(n5516), .ZN(U5775_n1) );
  AND2X1 U5776_U2 ( .IN1(test_so95), .IN2(U5776_n1), .Q(WX11200) );
  INVX0 U5776_U1 ( .INP(n5516), .ZN(U5776_n1) );
  AND2X1 U5777_U2 ( .IN1(WX11135), .IN2(U5777_n1), .Q(WX11198) );
  INVX0 U5777_U1 ( .INP(n5516), .ZN(U5777_n1) );
  AND2X1 U5778_U2 ( .IN1(WX11133), .IN2(U5778_n1), .Q(WX11196) );
  INVX0 U5778_U1 ( .INP(n5516), .ZN(U5778_n1) );
  AND2X1 U5779_U2 ( .IN1(WX11131), .IN2(U5779_n1), .Q(WX11194) );
  INVX0 U5779_U1 ( .INP(n5516), .ZN(U5779_n1) );
  AND2X1 U5780_U2 ( .IN1(WX11129), .IN2(U5780_n1), .Q(WX11192) );
  INVX0 U5780_U1 ( .INP(n5516), .ZN(U5780_n1) );
  AND2X1 U5781_U2 ( .IN1(WX11127), .IN2(U5781_n1), .Q(WX11190) );
  INVX0 U5781_U1 ( .INP(n5516), .ZN(U5781_n1) );
  AND2X1 U5782_U2 ( .IN1(WX11125), .IN2(U5782_n1), .Q(WX11188) );
  INVX0 U5782_U1 ( .INP(n5516), .ZN(U5782_n1) );
  AND2X1 U5783_U2 ( .IN1(WX11123), .IN2(U5783_n1), .Q(WX11186) );
  INVX0 U5783_U1 ( .INP(n5516), .ZN(U5783_n1) );
  AND2X1 U5784_U2 ( .IN1(WX11121), .IN2(U5784_n1), .Q(WX11184) );
  INVX0 U5784_U1 ( .INP(n5516), .ZN(U5784_n1) );
  AND2X1 U5785_U2 ( .IN1(WX11119), .IN2(U5785_n1), .Q(WX11182) );
  INVX0 U5785_U1 ( .INP(n5516), .ZN(U5785_n1) );
  AND2X1 U5786_U2 ( .IN1(WX11117), .IN2(U5786_n1), .Q(WX11180) );
  INVX0 U5786_U1 ( .INP(n5517), .ZN(U5786_n1) );
  AND2X1 U5787_U2 ( .IN1(WX11115), .IN2(U5787_n1), .Q(WX11178) );
  INVX0 U5787_U1 ( .INP(n5517), .ZN(U5787_n1) );
  AND2X1 U5788_U2 ( .IN1(WX11113), .IN2(U5788_n1), .Q(WX11176) );
  INVX0 U5788_U1 ( .INP(n5517), .ZN(U5788_n1) );
  AND2X1 U5789_U2 ( .IN1(WX11111), .IN2(U5789_n1), .Q(WX11174) );
  INVX0 U5789_U1 ( .INP(n5517), .ZN(U5789_n1) );
  AND2X1 U5790_U2 ( .IN1(WX11109), .IN2(U5790_n1), .Q(WX11172) );
  INVX0 U5790_U1 ( .INP(n5517), .ZN(U5790_n1) );
  AND2X1 U5791_U2 ( .IN1(WX11107), .IN2(U5791_n1), .Q(WX11170) );
  INVX0 U5791_U1 ( .INP(n5517), .ZN(U5791_n1) );
  AND2X1 U5792_U2 ( .IN1(WX11105), .IN2(U5792_n1), .Q(WX11168) );
  INVX0 U5792_U1 ( .INP(n5517), .ZN(U5792_n1) );
  AND2X1 U5793_U2 ( .IN1(test_so94), .IN2(U5793_n1), .Q(WX11166) );
  INVX0 U5793_U1 ( .INP(n5517), .ZN(U5793_n1) );
  AND2X1 U5794_U2 ( .IN1(WX11101), .IN2(U5794_n1), .Q(WX11164) );
  INVX0 U5794_U1 ( .INP(n5517), .ZN(U5794_n1) );
  AND2X1 U5795_U2 ( .IN1(WX11099), .IN2(U5795_n1), .Q(WX11162) );
  INVX0 U5795_U1 ( .INP(n5517), .ZN(U5795_n1) );
  AND2X1 U5796_U2 ( .IN1(WX11097), .IN2(U5796_n1), .Q(WX11160) );
  INVX0 U5796_U1 ( .INP(n5517), .ZN(U5796_n1) );
  AND2X1 U5797_U2 ( .IN1(WX11095), .IN2(U5797_n1), .Q(WX11158) );
  INVX0 U5797_U1 ( .INP(n5517), .ZN(U5797_n1) );
  AND2X1 U5798_U2 ( .IN1(WX11093), .IN2(U5798_n1), .Q(WX11156) );
  INVX0 U5798_U1 ( .INP(n5517), .ZN(U5798_n1) );
  AND2X1 U5799_U2 ( .IN1(WX11091), .IN2(U5799_n1), .Q(WX11154) );
  INVX0 U5799_U1 ( .INP(n5518), .ZN(U5799_n1) );
  AND2X1 U5800_U2 ( .IN1(WX11089), .IN2(U5800_n1), .Q(WX11152) );
  INVX0 U5800_U1 ( .INP(n5518), .ZN(U5800_n1) );
  AND2X1 U5801_U2 ( .IN1(WX11087), .IN2(U5801_n1), .Q(WX11150) );
  INVX0 U5801_U1 ( .INP(n5518), .ZN(U5801_n1) );
  AND2X1 U5802_U2 ( .IN1(WX11085), .IN2(U5802_n1), .Q(WX11148) );
  INVX0 U5802_U1 ( .INP(n5518), .ZN(U5802_n1) );
  AND2X1 U5803_U2 ( .IN1(WX11083), .IN2(U5803_n1), .Q(WX11146) );
  INVX0 U5803_U1 ( .INP(n5518), .ZN(U5803_n1) );
  AND2X1 U5804_U2 ( .IN1(WX11081), .IN2(U5804_n1), .Q(WX11144) );
  INVX0 U5804_U1 ( .INP(n5518), .ZN(U5804_n1) );
  AND2X1 U5805_U2 ( .IN1(WX11079), .IN2(U5805_n1), .Q(WX11142) );
  INVX0 U5805_U1 ( .INP(n5518), .ZN(U5805_n1) );
  AND2X1 U5806_U2 ( .IN1(WX11077), .IN2(U5806_n1), .Q(WX11140) );
  INVX0 U5806_U1 ( .INP(n5518), .ZN(U5806_n1) );
  AND2X1 U5807_U2 ( .IN1(WX11075), .IN2(U5807_n1), .Q(WX11138) );
  INVX0 U5807_U1 ( .INP(n5518), .ZN(U5807_n1) );
  AND2X1 U5808_U2 ( .IN1(WX11073), .IN2(U5808_n1), .Q(WX11136) );
  INVX0 U5808_U1 ( .INP(n5518), .ZN(U5808_n1) );
  AND2X1 U5809_U2 ( .IN1(WX11071), .IN2(U5809_n1), .Q(WX11134) );
  INVX0 U5809_U1 ( .INP(n5518), .ZN(U5809_n1) );
  AND2X1 U5810_U2 ( .IN1(test_so93), .IN2(U5810_n1), .Q(WX11132) );
  INVX0 U5810_U1 ( .INP(n5518), .ZN(U5810_n1) );
  AND2X1 U5811_U2 ( .IN1(WX11067), .IN2(U5811_n1), .Q(WX11130) );
  INVX0 U5811_U1 ( .INP(n5518), .ZN(U5811_n1) );
  AND2X1 U5812_U2 ( .IN1(WX11065), .IN2(U5812_n1), .Q(WX11128) );
  INVX0 U5812_U1 ( .INP(n5518), .ZN(U5812_n1) );
  AND2X1 U5813_U2 ( .IN1(WX11063), .IN2(U5813_n1), .Q(WX11126) );
  INVX0 U5813_U1 ( .INP(n5519), .ZN(U5813_n1) );
  AND2X1 U5814_U2 ( .IN1(WX11061), .IN2(U5814_n1), .Q(WX11124) );
  INVX0 U5814_U1 ( .INP(n5519), .ZN(U5814_n1) );
  AND2X1 U5815_U2 ( .IN1(WX11059), .IN2(U5815_n1), .Q(WX11122) );
  INVX0 U5815_U1 ( .INP(n5519), .ZN(U5815_n1) );
  AND2X1 U5816_U2 ( .IN1(WX11057), .IN2(U5816_n1), .Q(WX11120) );
  INVX0 U5816_U1 ( .INP(n5519), .ZN(U5816_n1) );
  AND2X1 U5817_U2 ( .IN1(WX11055), .IN2(U5817_n1), .Q(WX11118) );
  INVX0 U5817_U1 ( .INP(n5519), .ZN(U5817_n1) );
  AND2X1 U5818_U2 ( .IN1(WX11053), .IN2(U5818_n1), .Q(WX11116) );
  INVX0 U5818_U1 ( .INP(n5519), .ZN(U5818_n1) );
  AND2X1 U5819_U2 ( .IN1(WX11051), .IN2(U5819_n1), .Q(WX11114) );
  INVX0 U5819_U1 ( .INP(n5519), .ZN(U5819_n1) );
  AND2X1 U5820_U2 ( .IN1(WX11049), .IN2(U5820_n1), .Q(WX11112) );
  INVX0 U5820_U1 ( .INP(n5519), .ZN(U5820_n1) );
  AND2X1 U5821_U2 ( .IN1(WX11047), .IN2(U5821_n1), .Q(WX11110) );
  INVX0 U5821_U1 ( .INP(n5519), .ZN(U5821_n1) );
  AND2X1 U5822_U2 ( .IN1(WX11045), .IN2(U5822_n1), .Q(WX11108) );
  INVX0 U5822_U1 ( .INP(n5519), .ZN(U5822_n1) );
  AND2X1 U5823_U2 ( .IN1(WX11043), .IN2(U5823_n1), .Q(WX11106) );
  INVX0 U5823_U1 ( .INP(n5519), .ZN(U5823_n1) );
  AND2X1 U5824_U2 ( .IN1(WX11041), .IN2(U5824_n1), .Q(WX11104) );
  INVX0 U5824_U1 ( .INP(n5519), .ZN(U5824_n1) );
  AND2X1 U5825_U2 ( .IN1(WX11039), .IN2(U5825_n1), .Q(WX11102) );
  INVX0 U5825_U1 ( .INP(n5519), .ZN(U5825_n1) );
  AND2X1 U5826_U2 ( .IN1(WX11037), .IN2(U5826_n1), .Q(WX11100) );
  INVX0 U5826_U1 ( .INP(n5519), .ZN(U5826_n1) );
  AND2X1 U5827_U2 ( .IN1(test_so92), .IN2(U5827_n1), .Q(WX11098) );
  INVX0 U5827_U1 ( .INP(n5520), .ZN(U5827_n1) );
  AND2X1 U5828_U2 ( .IN1(WX11033), .IN2(U5828_n1), .Q(WX11096) );
  INVX0 U5828_U1 ( .INP(n5520), .ZN(U5828_n1) );
  AND2X1 U5829_U2 ( .IN1(WX11031), .IN2(U5829_n1), .Q(WX11094) );
  INVX0 U5829_U1 ( .INP(n5520), .ZN(U5829_n1) );
  AND2X1 U5830_U2 ( .IN1(WX11029), .IN2(U5830_n1), .Q(WX11092) );
  INVX0 U5830_U1 ( .INP(n5520), .ZN(U5830_n1) );
  AND2X1 U5831_U2 ( .IN1(WX11027), .IN2(U5831_n1), .Q(WX11090) );
  INVX0 U5831_U1 ( .INP(n5520), .ZN(U5831_n1) );
  AND2X1 U5832_U2 ( .IN1(WX11025), .IN2(U5832_n1), .Q(WX11088) );
  INVX0 U5832_U1 ( .INP(n5520), .ZN(U5832_n1) );
  AND2X1 U5833_U2 ( .IN1(WX11023), .IN2(U5833_n1), .Q(WX11086) );
  INVX0 U5833_U1 ( .INP(n5520), .ZN(U5833_n1) );
  AND2X1 U5834_U2 ( .IN1(WX11021), .IN2(U5834_n1), .Q(WX11084) );
  INVX0 U5834_U1 ( .INP(n5520), .ZN(U5834_n1) );
  AND2X1 U5835_U2 ( .IN1(WX9886), .IN2(U5835_n1), .Q(WX9949) );
  INVX0 U5835_U1 ( .INP(n5520), .ZN(U5835_n1) );
  AND2X1 U5836_U2 ( .IN1(WX9884), .IN2(U5836_n1), .Q(WX9947) );
  INVX0 U5836_U1 ( .INP(n5520), .ZN(U5836_n1) );
  AND2X1 U5837_U2 ( .IN1(WX9882), .IN2(U5837_n1), .Q(WX9945) );
  INVX0 U5837_U1 ( .INP(n5520), .ZN(U5837_n1) );
  AND2X1 U5838_U2 ( .IN1(WX9880), .IN2(U5838_n1), .Q(WX9943) );
  INVX0 U5838_U1 ( .INP(n5520), .ZN(U5838_n1) );
  AND2X1 U5839_U2 ( .IN1(WX9878), .IN2(U5839_n1), .Q(WX9941) );
  INVX0 U5839_U1 ( .INP(n5520), .ZN(U5839_n1) );
  AND2X1 U5840_U2 ( .IN1(WX9876), .IN2(U5840_n1), .Q(WX9939) );
  INVX0 U5840_U1 ( .INP(n5520), .ZN(U5840_n1) );
  AND2X1 U5841_U2 ( .IN1(WX9874), .IN2(U5841_n1), .Q(WX9937) );
  INVX0 U5841_U1 ( .INP(n5521), .ZN(U5841_n1) );
  AND2X1 U5842_U2 ( .IN1(WX9872), .IN2(U5842_n1), .Q(WX9935) );
  INVX0 U5842_U1 ( .INP(n5521), .ZN(U5842_n1) );
  AND2X1 U5843_U2 ( .IN1(WX9870), .IN2(U5843_n1), .Q(WX9933) );
  INVX0 U5843_U1 ( .INP(n5521), .ZN(U5843_n1) );
  AND2X1 U5844_U2 ( .IN1(WX9868), .IN2(U5844_n1), .Q(WX9931) );
  INVX0 U5844_U1 ( .INP(n5521), .ZN(U5844_n1) );
  AND2X1 U5845_U2 ( .IN1(WX9866), .IN2(U5845_n1), .Q(WX9929) );
  INVX0 U5845_U1 ( .INP(n5521), .ZN(U5845_n1) );
  AND2X1 U5846_U2 ( .IN1(WX9864), .IN2(U5846_n1), .Q(WX9927) );
  INVX0 U5846_U1 ( .INP(n5521), .ZN(U5846_n1) );
  AND2X1 U5847_U2 ( .IN1(WX9862), .IN2(U5847_n1), .Q(WX9925) );
  INVX0 U5847_U1 ( .INP(n5521), .ZN(U5847_n1) );
  AND2X1 U5848_U2 ( .IN1(WX9860), .IN2(U5848_n1), .Q(WX9923) );
  INVX0 U5848_U1 ( .INP(n5521), .ZN(U5848_n1) );
  AND2X1 U5849_U2 ( .IN1(WX9858), .IN2(U5849_n1), .Q(WX9921) );
  INVX0 U5849_U1 ( .INP(n5521), .ZN(U5849_n1) );
  AND2X1 U5850_U2 ( .IN1(WX9856), .IN2(U5850_n1), .Q(WX9919) );
  INVX0 U5850_U1 ( .INP(n5521), .ZN(U5850_n1) );
  AND2X1 U5851_U2 ( .IN1(test_so84), .IN2(U5851_n1), .Q(WX9917) );
  INVX0 U5851_U1 ( .INP(n5521), .ZN(U5851_n1) );
  AND2X1 U5852_U2 ( .IN1(WX9852), .IN2(U5852_n1), .Q(WX9915) );
  INVX0 U5852_U1 ( .INP(n5521), .ZN(U5852_n1) );
  AND2X1 U5853_U2 ( .IN1(WX9850), .IN2(U5853_n1), .Q(WX9913) );
  INVX0 U5853_U1 ( .INP(n5521), .ZN(U5853_n1) );
  AND2X1 U5854_U2 ( .IN1(WX9848), .IN2(U5854_n1), .Q(WX9911) );
  INVX0 U5854_U1 ( .INP(n5521), .ZN(U5854_n1) );
  AND2X1 U5855_U2 ( .IN1(WX9846), .IN2(U5855_n1), .Q(WX9909) );
  INVX0 U5855_U1 ( .INP(n5522), .ZN(U5855_n1) );
  AND2X1 U5856_U2 ( .IN1(WX9844), .IN2(U5856_n1), .Q(WX9907) );
  INVX0 U5856_U1 ( .INP(n5507), .ZN(U5856_n1) );
  AND2X1 U5857_U2 ( .IN1(WX9842), .IN2(U5857_n1), .Q(WX9905) );
  INVX0 U5857_U1 ( .INP(n5502), .ZN(U5857_n1) );
  AND2X1 U5858_U2 ( .IN1(WX9840), .IN2(U5858_n1), .Q(WX9903) );
  INVX0 U5858_U1 ( .INP(n5502), .ZN(U5858_n1) );
  AND2X1 U5859_U2 ( .IN1(WX9838), .IN2(U5859_n1), .Q(WX9901) );
  INVX0 U5859_U1 ( .INP(n5502), .ZN(U5859_n1) );
  AND2X1 U5860_U2 ( .IN1(WX9836), .IN2(U5860_n1), .Q(WX9899) );
  INVX0 U5860_U1 ( .INP(n5502), .ZN(U5860_n1) );
  AND2X1 U5861_U2 ( .IN1(WX9834), .IN2(U5861_n1), .Q(WX9897) );
  INVX0 U5861_U1 ( .INP(n5502), .ZN(U5861_n1) );
  AND2X1 U5862_U2 ( .IN1(WX9832), .IN2(U5862_n1), .Q(WX9895) );
  INVX0 U5862_U1 ( .INP(n5502), .ZN(U5862_n1) );
  AND2X1 U5863_U2 ( .IN1(WX9830), .IN2(U5863_n1), .Q(WX9893) );
  INVX0 U5863_U1 ( .INP(n5502), .ZN(U5863_n1) );
  AND2X1 U5864_U2 ( .IN1(WX9828), .IN2(U5864_n1), .Q(WX9891) );
  INVX0 U5864_U1 ( .INP(n5502), .ZN(U5864_n1) );
  AND2X1 U5865_U2 ( .IN1(WX9826), .IN2(U5865_n1), .Q(WX9889) );
  INVX0 U5865_U1 ( .INP(n5503), .ZN(U5865_n1) );
  AND2X1 U5866_U2 ( .IN1(WX9824), .IN2(U5866_n1), .Q(WX9887) );
  INVX0 U5866_U1 ( .INP(n5503), .ZN(U5866_n1) );
  AND2X1 U5867_U2 ( .IN1(WX9822), .IN2(U5867_n1), .Q(WX9885) );
  INVX0 U5867_U1 ( .INP(n5503), .ZN(U5867_n1) );
  AND2X1 U5868_U2 ( .IN1(test_so83), .IN2(U5868_n1), .Q(WX9883) );
  INVX0 U5868_U1 ( .INP(n5503), .ZN(U5868_n1) );
  AND2X1 U5869_U2 ( .IN1(WX9818), .IN2(U5869_n1), .Q(WX9881) );
  INVX0 U5869_U1 ( .INP(n5503), .ZN(U5869_n1) );
  AND2X1 U5870_U2 ( .IN1(WX9816), .IN2(U5870_n1), .Q(WX9879) );
  INVX0 U5870_U1 ( .INP(n5503), .ZN(U5870_n1) );
  AND2X1 U5871_U2 ( .IN1(WX9814), .IN2(U5871_n1), .Q(WX9877) );
  INVX0 U5871_U1 ( .INP(n5503), .ZN(U5871_n1) );
  AND2X1 U5872_U2 ( .IN1(WX9812), .IN2(U5872_n1), .Q(WX9875) );
  INVX0 U5872_U1 ( .INP(n5503), .ZN(U5872_n1) );
  AND2X1 U5873_U2 ( .IN1(WX9810), .IN2(U5873_n1), .Q(WX9873) );
  INVX0 U5873_U1 ( .INP(n5503), .ZN(U5873_n1) );
  AND2X1 U5874_U2 ( .IN1(WX9808), .IN2(U5874_n1), .Q(WX9871) );
  INVX0 U5874_U1 ( .INP(n5503), .ZN(U5874_n1) );
  AND2X1 U5875_U2 ( .IN1(WX9806), .IN2(U5875_n1), .Q(WX9869) );
  INVX0 U5875_U1 ( .INP(n5503), .ZN(U5875_n1) );
  AND2X1 U5876_U2 ( .IN1(WX9804), .IN2(U5876_n1), .Q(WX9867) );
  INVX0 U5876_U1 ( .INP(n5503), .ZN(U5876_n1) );
  AND2X1 U5877_U2 ( .IN1(WX9802), .IN2(U5877_n1), .Q(WX9865) );
  INVX0 U5877_U1 ( .INP(n5503), .ZN(U5877_n1) );
  AND2X1 U5878_U2 ( .IN1(WX9800), .IN2(U5878_n1), .Q(WX9863) );
  INVX0 U5878_U1 ( .INP(n5503), .ZN(U5878_n1) );
  AND2X1 U5879_U2 ( .IN1(WX9798), .IN2(U5879_n1), .Q(WX9861) );
  INVX0 U5879_U1 ( .INP(n5504), .ZN(U5879_n1) );
  AND2X1 U5880_U2 ( .IN1(WX9796), .IN2(U5880_n1), .Q(WX9859) );
  INVX0 U5880_U1 ( .INP(n5504), .ZN(U5880_n1) );
  AND2X1 U5881_U2 ( .IN1(WX9794), .IN2(U5881_n1), .Q(WX9857) );
  INVX0 U5881_U1 ( .INP(n5504), .ZN(U5881_n1) );
  AND2X1 U5882_U2 ( .IN1(WX9792), .IN2(U5882_n1), .Q(WX9855) );
  INVX0 U5882_U1 ( .INP(n5504), .ZN(U5882_n1) );
  AND2X1 U5883_U2 ( .IN1(WX9790), .IN2(U5883_n1), .Q(WX9853) );
  INVX0 U5883_U1 ( .INP(n5504), .ZN(U5883_n1) );
  AND2X1 U5884_U2 ( .IN1(WX9788), .IN2(U5884_n1), .Q(WX9851) );
  INVX0 U5884_U1 ( .INP(n5504), .ZN(U5884_n1) );
  AND2X1 U5885_U2 ( .IN1(test_so82), .IN2(U5885_n1), .Q(WX9849) );
  INVX0 U5885_U1 ( .INP(n5504), .ZN(U5885_n1) );
  AND2X1 U5886_U2 ( .IN1(WX9784), .IN2(U5886_n1), .Q(WX9847) );
  INVX0 U5886_U1 ( .INP(n5504), .ZN(U5886_n1) );
  AND2X1 U5887_U2 ( .IN1(WX9782), .IN2(U5887_n1), .Q(WX9845) );
  INVX0 U5887_U1 ( .INP(n5504), .ZN(U5887_n1) );
  AND2X1 U5888_U2 ( .IN1(WX9780), .IN2(U5888_n1), .Q(WX9843) );
  INVX0 U5888_U1 ( .INP(n5504), .ZN(U5888_n1) );
  AND2X1 U5889_U2 ( .IN1(WX9778), .IN2(U5889_n1), .Q(WX9841) );
  INVX0 U5889_U1 ( .INP(n5504), .ZN(U5889_n1) );
  AND2X1 U5890_U2 ( .IN1(WX9776), .IN2(U5890_n1), .Q(WX9839) );
  INVX0 U5890_U1 ( .INP(n5504), .ZN(U5890_n1) );
  AND2X1 U5891_U2 ( .IN1(WX9774), .IN2(U5891_n1), .Q(WX9837) );
  INVX0 U5891_U1 ( .INP(n5504), .ZN(U5891_n1) );
  AND2X1 U5892_U2 ( .IN1(WX9772), .IN2(U5892_n1), .Q(WX9835) );
  INVX0 U5892_U1 ( .INP(n5504), .ZN(U5892_n1) );
  AND2X1 U5893_U2 ( .IN1(WX9770), .IN2(U5893_n1), .Q(WX9833) );
  INVX0 U5893_U1 ( .INP(n5505), .ZN(U5893_n1) );
  AND2X1 U5894_U2 ( .IN1(WX9768), .IN2(U5894_n1), .Q(WX9831) );
  INVX0 U5894_U1 ( .INP(n5505), .ZN(U5894_n1) );
  AND2X1 U5895_U2 ( .IN1(WX9766), .IN2(U5895_n1), .Q(WX9829) );
  INVX0 U5895_U1 ( .INP(n5505), .ZN(U5895_n1) );
  AND2X1 U5896_U2 ( .IN1(WX9764), .IN2(U5896_n1), .Q(WX9827) );
  INVX0 U5896_U1 ( .INP(n5505), .ZN(U5896_n1) );
  AND2X1 U5897_U2 ( .IN1(WX9762), .IN2(U5897_n1), .Q(WX9825) );
  INVX0 U5897_U1 ( .INP(n5505), .ZN(U5897_n1) );
  AND2X1 U5898_U2 ( .IN1(WX9760), .IN2(U5898_n1), .Q(WX9823) );
  INVX0 U5898_U1 ( .INP(n5505), .ZN(U5898_n1) );
  AND2X1 U5899_U2 ( .IN1(WX9758), .IN2(U5899_n1), .Q(WX9821) );
  INVX0 U5899_U1 ( .INP(n5505), .ZN(U5899_n1) );
  AND2X1 U5900_U2 ( .IN1(WX9756), .IN2(U5900_n1), .Q(WX9819) );
  INVX0 U5900_U1 ( .INP(n5505), .ZN(U5900_n1) );
  AND2X1 U5901_U2 ( .IN1(WX9754), .IN2(U5901_n1), .Q(WX9817) );
  INVX0 U5901_U1 ( .INP(n5505), .ZN(U5901_n1) );
  AND2X1 U5902_U2 ( .IN1(test_so81), .IN2(U5902_n1), .Q(WX9815) );
  INVX0 U5902_U1 ( .INP(n5505), .ZN(U5902_n1) );
  AND2X1 U5903_U2 ( .IN1(WX9750), .IN2(U5903_n1), .Q(WX9813) );
  INVX0 U5903_U1 ( .INP(n5505), .ZN(U5903_n1) );
  AND2X1 U5904_U2 ( .IN1(WX9748), .IN2(U5904_n1), .Q(WX9811) );
  INVX0 U5904_U1 ( .INP(n5505), .ZN(U5904_n1) );
  AND2X1 U5905_U2 ( .IN1(WX9746), .IN2(U5905_n1), .Q(WX9809) );
  INVX0 U5905_U1 ( .INP(n5505), .ZN(U5905_n1) );
  AND2X1 U5906_U2 ( .IN1(WX9744), .IN2(U5906_n1), .Q(WX9807) );
  INVX0 U5906_U1 ( .INP(n5505), .ZN(U5906_n1) );
  AND2X1 U5907_U2 ( .IN1(WX9742), .IN2(U5907_n1), .Q(WX9805) );
  INVX0 U5907_U1 ( .INP(n5506), .ZN(U5907_n1) );
  AND2X1 U5908_U2 ( .IN1(WX9740), .IN2(U5908_n1), .Q(WX9803) );
  INVX0 U5908_U1 ( .INP(n5506), .ZN(U5908_n1) );
  AND2X1 U5909_U2 ( .IN1(WX9738), .IN2(U5909_n1), .Q(WX9801) );
  INVX0 U5909_U1 ( .INP(n5506), .ZN(U5909_n1) );
  AND2X1 U5910_U2 ( .IN1(WX9736), .IN2(U5910_n1), .Q(WX9799) );
  INVX0 U5910_U1 ( .INP(n5506), .ZN(U5910_n1) );
  AND2X1 U5911_U2 ( .IN1(WX9734), .IN2(U5911_n1), .Q(WX9797) );
  INVX0 U5911_U1 ( .INP(n5506), .ZN(U5911_n1) );
  AND2X1 U5912_U2 ( .IN1(WX9732), .IN2(U5912_n1), .Q(WX9795) );
  INVX0 U5912_U1 ( .INP(n5506), .ZN(U5912_n1) );
  AND2X1 U5913_U2 ( .IN1(WX9730), .IN2(U5913_n1), .Q(WX9793) );
  INVX0 U5913_U1 ( .INP(n5506), .ZN(U5913_n1) );
  AND2X1 U5914_U2 ( .IN1(WX9728), .IN2(U5914_n1), .Q(WX9791) );
  INVX0 U5914_U1 ( .INP(n5506), .ZN(U5914_n1) );
  AND2X1 U5915_U2 ( .IN1(WX8593), .IN2(U5915_n1), .Q(WX8656) );
  INVX0 U5915_U1 ( .INP(n5506), .ZN(U5915_n1) );
  AND2X1 U5916_U2 ( .IN1(WX8591), .IN2(U5916_n1), .Q(WX8654) );
  INVX0 U5916_U1 ( .INP(n5506), .ZN(U5916_n1) );
  AND2X1 U5917_U2 ( .IN1(WX8589), .IN2(U5917_n1), .Q(WX8652) );
  INVX0 U5917_U1 ( .INP(n5506), .ZN(U5917_n1) );
  AND2X1 U5918_U2 ( .IN1(WX8587), .IN2(U5918_n1), .Q(WX8650) );
  INVX0 U5918_U1 ( .INP(n5506), .ZN(U5918_n1) );
  AND2X1 U5919_U2 ( .IN1(WX8585), .IN2(U5919_n1), .Q(WX8648) );
  INVX0 U5919_U1 ( .INP(n5506), .ZN(U5919_n1) );
  AND2X1 U5920_U2 ( .IN1(WX8583), .IN2(U5920_n1), .Q(WX8646) );
  INVX0 U5920_U1 ( .INP(n5506), .ZN(U5920_n1) );
  AND2X1 U5921_U2 ( .IN1(WX8581), .IN2(U5921_n1), .Q(WX8644) );
  INVX0 U5921_U1 ( .INP(n5507), .ZN(U5921_n1) );
  AND2X1 U5922_U2 ( .IN1(WX8579), .IN2(U5922_n1), .Q(WX8642) );
  INVX0 U5922_U1 ( .INP(n5507), .ZN(U5922_n1) );
  AND2X1 U5923_U2 ( .IN1(WX8577), .IN2(U5923_n1), .Q(WX8640) );
  INVX0 U5923_U1 ( .INP(n5507), .ZN(U5923_n1) );
  AND2X1 U5924_U2 ( .IN1(WX8575), .IN2(U5924_n1), .Q(WX8638) );
  INVX0 U5924_U1 ( .INP(n5507), .ZN(U5924_n1) );
  AND2X1 U5925_U2 ( .IN1(WX8573), .IN2(U5925_n1), .Q(WX8636) );
  INVX0 U5925_U1 ( .INP(n5507), .ZN(U5925_n1) );
  AND2X1 U5926_U2 ( .IN1(test_so73), .IN2(U5926_n1), .Q(WX8634) );
  INVX0 U5926_U1 ( .INP(n5507), .ZN(U5926_n1) );
  AND2X1 U5927_U2 ( .IN1(WX8569), .IN2(U5927_n1), .Q(WX8632) );
  INVX0 U5927_U1 ( .INP(n5507), .ZN(U5927_n1) );
  AND2X1 U5928_U2 ( .IN1(WX8567), .IN2(U5928_n1), .Q(WX8630) );
  INVX0 U5928_U1 ( .INP(n5507), .ZN(U5928_n1) );
  AND2X1 U5929_U2 ( .IN1(WX8565), .IN2(U5929_n1), .Q(WX8628) );
  INVX0 U5929_U1 ( .INP(n5507), .ZN(U5929_n1) );
  AND2X1 U5930_U2 ( .IN1(WX8563), .IN2(U5930_n1), .Q(WX8626) );
  INVX0 U5930_U1 ( .INP(n5507), .ZN(U5930_n1) );
  AND2X1 U5931_U2 ( .IN1(WX8561), .IN2(U5931_n1), .Q(WX8624) );
  INVX0 U5931_U1 ( .INP(n5507), .ZN(U5931_n1) );
  AND2X1 U5932_U2 ( .IN1(WX8559), .IN2(U5932_n1), .Q(WX8622) );
  INVX0 U5932_U1 ( .INP(n5507), .ZN(U5932_n1) );
  AND2X1 U5933_U2 ( .IN1(WX8557), .IN2(U5933_n1), .Q(WX8620) );
  INVX0 U5933_U1 ( .INP(n5507), .ZN(U5933_n1) );
  AND2X1 U5934_U2 ( .IN1(WX8555), .IN2(U5934_n1), .Q(WX8618) );
  INVX0 U5934_U1 ( .INP(n5508), .ZN(U5934_n1) );
  AND2X1 U5935_U2 ( .IN1(WX8553), .IN2(U5935_n1), .Q(WX8616) );
  INVX0 U5935_U1 ( .INP(n5508), .ZN(U5935_n1) );
  AND2X1 U5936_U2 ( .IN1(WX8551), .IN2(U5936_n1), .Q(WX8614) );
  INVX0 U5936_U1 ( .INP(n5508), .ZN(U5936_n1) );
  AND2X1 U5937_U2 ( .IN1(WX8549), .IN2(U5937_n1), .Q(WX8612) );
  INVX0 U5937_U1 ( .INP(n5508), .ZN(U5937_n1) );
  AND2X1 U5938_U2 ( .IN1(WX8547), .IN2(U5938_n1), .Q(WX8610) );
  INVX0 U5938_U1 ( .INP(n5508), .ZN(U5938_n1) );
  AND2X1 U5939_U2 ( .IN1(WX8545), .IN2(U5939_n1), .Q(WX8608) );
  INVX0 U5939_U1 ( .INP(n5508), .ZN(U5939_n1) );
  AND2X1 U5940_U2 ( .IN1(WX8543), .IN2(U5940_n1), .Q(WX8606) );
  INVX0 U5940_U1 ( .INP(n5508), .ZN(U5940_n1) );
  AND2X1 U5941_U2 ( .IN1(WX8541), .IN2(U5941_n1), .Q(WX8604) );
  INVX0 U5941_U1 ( .INP(n5508), .ZN(U5941_n1) );
  AND2X1 U5942_U2 ( .IN1(WX8539), .IN2(U5942_n1), .Q(WX8602) );
  INVX0 U5942_U1 ( .INP(n5508), .ZN(U5942_n1) );
  AND2X1 U5943_U2 ( .IN1(test_so72), .IN2(U5943_n1), .Q(WX8600) );
  INVX0 U5943_U1 ( .INP(n5508), .ZN(U5943_n1) );
  AND2X1 U5944_U2 ( .IN1(WX8535), .IN2(U5944_n1), .Q(WX8598) );
  INVX0 U5944_U1 ( .INP(n5508), .ZN(U5944_n1) );
  AND2X1 U5945_U2 ( .IN1(WX8533), .IN2(U5945_n1), .Q(WX8596) );
  INVX0 U5945_U1 ( .INP(n5508), .ZN(U5945_n1) );
  AND2X1 U5946_U2 ( .IN1(WX8531), .IN2(U5946_n1), .Q(WX8594) );
  INVX0 U5946_U1 ( .INP(n5508), .ZN(U5946_n1) );
  AND2X1 U5947_U2 ( .IN1(WX8529), .IN2(U5947_n1), .Q(WX8592) );
  INVX0 U5947_U1 ( .INP(n5508), .ZN(U5947_n1) );
  AND2X1 U5948_U2 ( .IN1(WX8527), .IN2(U5948_n1), .Q(WX8590) );
  INVX0 U5948_U1 ( .INP(n5509), .ZN(U5948_n1) );
  AND2X1 U5949_U2 ( .IN1(WX8525), .IN2(U5949_n1), .Q(WX8588) );
  INVX0 U5949_U1 ( .INP(n5509), .ZN(U5949_n1) );
  AND2X1 U5950_U2 ( .IN1(WX8523), .IN2(U5950_n1), .Q(WX8586) );
  INVX0 U5950_U1 ( .INP(n5509), .ZN(U5950_n1) );
  AND2X1 U5951_U2 ( .IN1(WX8521), .IN2(U5951_n1), .Q(WX8584) );
  INVX0 U5951_U1 ( .INP(n5509), .ZN(U5951_n1) );
  AND2X1 U5952_U2 ( .IN1(WX8519), .IN2(U5952_n1), .Q(WX8582) );
  INVX0 U5952_U1 ( .INP(n5509), .ZN(U5952_n1) );
  AND2X1 U5953_U2 ( .IN1(WX8517), .IN2(U5953_n1), .Q(WX8580) );
  INVX0 U5953_U1 ( .INP(n5509), .ZN(U5953_n1) );
  AND2X1 U5954_U2 ( .IN1(WX8515), .IN2(U5954_n1), .Q(WX8578) );
  INVX0 U5954_U1 ( .INP(n5509), .ZN(U5954_n1) );
  AND2X1 U5955_U2 ( .IN1(WX8513), .IN2(U5955_n1), .Q(WX8576) );
  INVX0 U5955_U1 ( .INP(n5509), .ZN(U5955_n1) );
  AND2X1 U5956_U2 ( .IN1(WX8511), .IN2(U5956_n1), .Q(WX8574) );
  INVX0 U5956_U1 ( .INP(n5509), .ZN(U5956_n1) );
  AND2X1 U5957_U2 ( .IN1(WX8509), .IN2(U5957_n1), .Q(WX8572) );
  INVX0 U5957_U1 ( .INP(n5509), .ZN(U5957_n1) );
  AND2X1 U5958_U2 ( .IN1(WX8507), .IN2(U5958_n1), .Q(WX8570) );
  INVX0 U5958_U1 ( .INP(n5509), .ZN(U5958_n1) );
  AND2X1 U5959_U2 ( .IN1(WX8505), .IN2(U5959_n1), .Q(WX8568) );
  INVX0 U5959_U1 ( .INP(n5509), .ZN(U5959_n1) );
  AND2X1 U5960_U2 ( .IN1(test_so71), .IN2(U5960_n1), .Q(WX8566) );
  INVX0 U5960_U1 ( .INP(n5509), .ZN(U5960_n1) );
  AND2X1 U5961_U2 ( .IN1(WX8501), .IN2(U5961_n1), .Q(WX8564) );
  INVX0 U5961_U1 ( .INP(n5509), .ZN(U5961_n1) );
  AND2X1 U5962_U2 ( .IN1(WX8499), .IN2(U5962_n1), .Q(WX8562) );
  INVX0 U5962_U1 ( .INP(n5510), .ZN(U5962_n1) );
  AND2X1 U5963_U2 ( .IN1(WX8497), .IN2(U5963_n1), .Q(WX8560) );
  INVX0 U5963_U1 ( .INP(n5510), .ZN(U5963_n1) );
  AND2X1 U5964_U2 ( .IN1(WX8495), .IN2(U5964_n1), .Q(WX8558) );
  INVX0 U5964_U1 ( .INP(n5510), .ZN(U5964_n1) );
  AND2X1 U5965_U2 ( .IN1(WX8493), .IN2(U5965_n1), .Q(WX8556) );
  INVX0 U5965_U1 ( .INP(n5510), .ZN(U5965_n1) );
  AND2X1 U5966_U2 ( .IN1(WX8491), .IN2(U5966_n1), .Q(WX8554) );
  INVX0 U5966_U1 ( .INP(n5510), .ZN(U5966_n1) );
  AND2X1 U5967_U2 ( .IN1(WX8489), .IN2(U5967_n1), .Q(WX8552) );
  INVX0 U5967_U1 ( .INP(n5510), .ZN(U5967_n1) );
  AND2X1 U5968_U2 ( .IN1(WX8487), .IN2(U5968_n1), .Q(WX8550) );
  INVX0 U5968_U1 ( .INP(n5510), .ZN(U5968_n1) );
  AND2X1 U5969_U2 ( .IN1(WX8485), .IN2(U5969_n1), .Q(WX8548) );
  INVX0 U5969_U1 ( .INP(n5510), .ZN(U5969_n1) );
  AND2X1 U5970_U2 ( .IN1(WX8483), .IN2(U5970_n1), .Q(WX8546) );
  INVX0 U5970_U1 ( .INP(n5510), .ZN(U5970_n1) );
  AND2X1 U5971_U2 ( .IN1(WX8481), .IN2(U5971_n1), .Q(WX8544) );
  INVX0 U5971_U1 ( .INP(n5510), .ZN(U5971_n1) );
  AND2X1 U5972_U2 ( .IN1(WX8479), .IN2(U5972_n1), .Q(WX8542) );
  INVX0 U5972_U1 ( .INP(n5510), .ZN(U5972_n1) );
  AND2X1 U5973_U2 ( .IN1(WX8477), .IN2(U5973_n1), .Q(WX8540) );
  INVX0 U5973_U1 ( .INP(n5510), .ZN(U5973_n1) );
  AND2X1 U5974_U2 ( .IN1(WX8475), .IN2(U5974_n1), .Q(WX8538) );
  INVX0 U5974_U1 ( .INP(n5510), .ZN(U5974_n1) );
  AND2X1 U5975_U2 ( .IN1(WX8473), .IN2(U5975_n1), .Q(WX8536) );
  INVX0 U5975_U1 ( .INP(n5510), .ZN(U5975_n1) );
  AND2X1 U5976_U2 ( .IN1(WX8471), .IN2(U5976_n1), .Q(WX8534) );
  INVX0 U5976_U1 ( .INP(n5511), .ZN(U5976_n1) );
  AND2X1 U5977_U2 ( .IN1(test_so70), .IN2(U5977_n1), .Q(WX8532) );
  INVX0 U5977_U1 ( .INP(n5511), .ZN(U5977_n1) );
  AND2X1 U5978_U2 ( .IN1(WX8467), .IN2(U5978_n1), .Q(WX8530) );
  INVX0 U5978_U1 ( .INP(n5511), .ZN(U5978_n1) );
  AND2X1 U5979_U2 ( .IN1(WX8465), .IN2(U5979_n1), .Q(WX8528) );
  INVX0 U5979_U1 ( .INP(n5511), .ZN(U5979_n1) );
  AND2X1 U5980_U2 ( .IN1(WX8463), .IN2(U5980_n1), .Q(WX8526) );
  INVX0 U5980_U1 ( .INP(n5511), .ZN(U5980_n1) );
  AND2X1 U5981_U2 ( .IN1(WX8461), .IN2(U5981_n1), .Q(WX8524) );
  INVX0 U5981_U1 ( .INP(n5511), .ZN(U5981_n1) );
  AND2X1 U5982_U2 ( .IN1(WX8459), .IN2(U5982_n1), .Q(WX8522) );
  INVX0 U5982_U1 ( .INP(n5511), .ZN(U5982_n1) );
  AND2X1 U5983_U2 ( .IN1(WX8457), .IN2(U5983_n1), .Q(WX8520) );
  INVX0 U5983_U1 ( .INP(n5511), .ZN(U5983_n1) );
  AND2X1 U5984_U2 ( .IN1(WX8455), .IN2(U5984_n1), .Q(WX8518) );
  INVX0 U5984_U1 ( .INP(n5511), .ZN(U5984_n1) );
  AND2X1 U5985_U2 ( .IN1(WX8453), .IN2(U5985_n1), .Q(WX8516) );
  INVX0 U5985_U1 ( .INP(n5511), .ZN(U5985_n1) );
  AND2X1 U5986_U2 ( .IN1(WX8451), .IN2(U5986_n1), .Q(WX8514) );
  INVX0 U5986_U1 ( .INP(n5511), .ZN(U5986_n1) );
  AND2X1 U5987_U2 ( .IN1(WX8449), .IN2(U5987_n1), .Q(WX8512) );
  INVX0 U5987_U1 ( .INP(n5511), .ZN(U5987_n1) );
  AND2X1 U5988_U2 ( .IN1(WX8447), .IN2(U5988_n1), .Q(WX8510) );
  INVX0 U5988_U1 ( .INP(n5511), .ZN(U5988_n1) );
  AND2X1 U5989_U2 ( .IN1(WX8445), .IN2(U5989_n1), .Q(WX8508) );
  INVX0 U5989_U1 ( .INP(n5511), .ZN(U5989_n1) );
  AND2X1 U5990_U2 ( .IN1(WX8443), .IN2(U5990_n1), .Q(WX8506) );
  INVX0 U5990_U1 ( .INP(n5512), .ZN(U5990_n1) );
  AND2X1 U5991_U2 ( .IN1(WX8441), .IN2(U5991_n1), .Q(WX8504) );
  INVX0 U5991_U1 ( .INP(n5512), .ZN(U5991_n1) );
  AND2X1 U5992_U2 ( .IN1(WX8439), .IN2(U5992_n1), .Q(WX8502) );
  INVX0 U5992_U1 ( .INP(n5512), .ZN(U5992_n1) );
  AND2X1 U5993_U2 ( .IN1(WX8437), .IN2(U5993_n1), .Q(WX8500) );
  INVX0 U5993_U1 ( .INP(n5512), .ZN(U5993_n1) );
  AND2X1 U5994_U2 ( .IN1(test_so69), .IN2(U5994_n1), .Q(WX8498) );
  INVX0 U5994_U1 ( .INP(n5536), .ZN(U5994_n1) );
  AND2X1 U5995_U2 ( .IN1(WX7300), .IN2(U5995_n1), .Q(WX7363) );
  INVX0 U5995_U1 ( .INP(n5532), .ZN(U5995_n1) );
  AND2X1 U5996_U2 ( .IN1(WX7298), .IN2(U5996_n1), .Q(WX7361) );
  INVX0 U5996_U1 ( .INP(n5532), .ZN(U5996_n1) );
  AND2X1 U5997_U2 ( .IN1(WX7296), .IN2(U5997_n1), .Q(WX7359) );
  INVX0 U5997_U1 ( .INP(n5532), .ZN(U5997_n1) );
  AND2X1 U5998_U2 ( .IN1(WX7294), .IN2(U5998_n1), .Q(WX7357) );
  INVX0 U5998_U1 ( .INP(n5532), .ZN(U5998_n1) );
  AND2X1 U5999_U2 ( .IN1(WX7292), .IN2(U5999_n1), .Q(WX7355) );
  INVX0 U5999_U1 ( .INP(n5532), .ZN(U5999_n1) );
  AND2X1 U6000_U2 ( .IN1(WX7290), .IN2(U6000_n1), .Q(WX7353) );
  INVX0 U6000_U1 ( .INP(n5532), .ZN(U6000_n1) );
  AND2X1 U6001_U2 ( .IN1(test_so62), .IN2(U6001_n1), .Q(WX7351) );
  INVX0 U6001_U1 ( .INP(n5532), .ZN(U6001_n1) );
  AND2X1 U6002_U2 ( .IN1(WX7286), .IN2(U6002_n1), .Q(WX7349) );
  INVX0 U6002_U1 ( .INP(n5532), .ZN(U6002_n1) );
  AND2X1 U6003_U2 ( .IN1(WX7284), .IN2(U6003_n1), .Q(WX7347) );
  INVX0 U6003_U1 ( .INP(n5532), .ZN(U6003_n1) );
  AND2X1 U6004_U2 ( .IN1(WX7282), .IN2(U6004_n1), .Q(WX7345) );
  INVX0 U6004_U1 ( .INP(n5532), .ZN(U6004_n1) );
  AND2X1 U6005_U2 ( .IN1(WX7280), .IN2(U6005_n1), .Q(WX7343) );
  INVX0 U6005_U1 ( .INP(n5532), .ZN(U6005_n1) );
  AND2X1 U6006_U2 ( .IN1(WX7278), .IN2(U6006_n1), .Q(WX7341) );
  INVX0 U6006_U1 ( .INP(n5532), .ZN(U6006_n1) );
  AND2X1 U6007_U2 ( .IN1(WX7276), .IN2(U6007_n1), .Q(WX7339) );
  INVX0 U6007_U1 ( .INP(n5532), .ZN(U6007_n1) );
  AND2X1 U6008_U2 ( .IN1(WX7274), .IN2(U6008_n1), .Q(WX7337) );
  INVX0 U6008_U1 ( .INP(n5532), .ZN(U6008_n1) );
  AND2X1 U6009_U2 ( .IN1(WX7272), .IN2(U6009_n1), .Q(WX7335) );
  INVX0 U6009_U1 ( .INP(n5533), .ZN(U6009_n1) );
  AND2X1 U6010_U2 ( .IN1(WX7270), .IN2(U6010_n1), .Q(WX7333) );
  INVX0 U6010_U1 ( .INP(n5533), .ZN(U6010_n1) );
  AND2X1 U6011_U2 ( .IN1(WX7268), .IN2(U6011_n1), .Q(WX7331) );
  INVX0 U6011_U1 ( .INP(n5533), .ZN(U6011_n1) );
  AND2X1 U6012_U2 ( .IN1(WX7266), .IN2(U6012_n1), .Q(WX7329) );
  INVX0 U6012_U1 ( .INP(n5533), .ZN(U6012_n1) );
  AND2X1 U6013_U2 ( .IN1(WX7264), .IN2(U6013_n1), .Q(WX7327) );
  INVX0 U6013_U1 ( .INP(n5533), .ZN(U6013_n1) );
  AND2X1 U6014_U2 ( .IN1(WX7262), .IN2(U6014_n1), .Q(WX7325) );
  INVX0 U6014_U1 ( .INP(n5533), .ZN(U6014_n1) );
  AND2X1 U6015_U2 ( .IN1(WX7260), .IN2(U6015_n1), .Q(WX7323) );
  INVX0 U6015_U1 ( .INP(n5533), .ZN(U6015_n1) );
  AND2X1 U6016_U2 ( .IN1(WX7258), .IN2(U6016_n1), .Q(WX7321) );
  INVX0 U6016_U1 ( .INP(n5533), .ZN(U6016_n1) );
  AND2X1 U6017_U2 ( .IN1(WX7256), .IN2(U6017_n1), .Q(WX7319) );
  INVX0 U6017_U1 ( .INP(n5533), .ZN(U6017_n1) );
  AND2X1 U6018_U2 ( .IN1(test_so61), .IN2(U6018_n1), .Q(WX7317) );
  INVX0 U6018_U1 ( .INP(n5533), .ZN(U6018_n1) );
  AND2X1 U6019_U2 ( .IN1(WX7252), .IN2(U6019_n1), .Q(WX7315) );
  INVX0 U6019_U1 ( .INP(n5533), .ZN(U6019_n1) );
  AND2X1 U6020_U2 ( .IN1(WX7250), .IN2(U6020_n1), .Q(WX7313) );
  INVX0 U6020_U1 ( .INP(n5533), .ZN(U6020_n1) );
  AND2X1 U6021_U2 ( .IN1(WX7248), .IN2(U6021_n1), .Q(WX7311) );
  INVX0 U6021_U1 ( .INP(n5533), .ZN(U6021_n1) );
  AND2X1 U6022_U2 ( .IN1(WX7246), .IN2(U6022_n1), .Q(WX7309) );
  INVX0 U6022_U1 ( .INP(n5533), .ZN(U6022_n1) );
  AND2X1 U6023_U2 ( .IN1(WX7244), .IN2(U6023_n1), .Q(WX7307) );
  INVX0 U6023_U1 ( .INP(n5534), .ZN(U6023_n1) );
  AND2X1 U6024_U2 ( .IN1(WX7242), .IN2(U6024_n1), .Q(WX7305) );
  INVX0 U6024_U1 ( .INP(n5534), .ZN(U6024_n1) );
  AND2X1 U6025_U2 ( .IN1(WX7240), .IN2(U6025_n1), .Q(WX7303) );
  INVX0 U6025_U1 ( .INP(n5534), .ZN(U6025_n1) );
  AND2X1 U6026_U2 ( .IN1(WX7238), .IN2(U6026_n1), .Q(WX7301) );
  INVX0 U6026_U1 ( .INP(n5534), .ZN(U6026_n1) );
  AND2X1 U6027_U2 ( .IN1(WX7236), .IN2(U6027_n1), .Q(WX7299) );
  INVX0 U6027_U1 ( .INP(n5534), .ZN(U6027_n1) );
  AND2X1 U6028_U2 ( .IN1(WX7234), .IN2(U6028_n1), .Q(WX7297) );
  INVX0 U6028_U1 ( .INP(n5534), .ZN(U6028_n1) );
  AND2X1 U6029_U2 ( .IN1(WX7232), .IN2(U6029_n1), .Q(WX7295) );
  INVX0 U6029_U1 ( .INP(n5534), .ZN(U6029_n1) );
  AND2X1 U6030_U2 ( .IN1(WX7230), .IN2(U6030_n1), .Q(WX7293) );
  INVX0 U6030_U1 ( .INP(n5534), .ZN(U6030_n1) );
  AND2X1 U6031_U2 ( .IN1(WX7228), .IN2(U6031_n1), .Q(WX7291) );
  INVX0 U6031_U1 ( .INP(n5534), .ZN(U6031_n1) );
  AND2X1 U6032_U2 ( .IN1(WX7226), .IN2(U6032_n1), .Q(WX7289) );
  INVX0 U6032_U1 ( .INP(n5534), .ZN(U6032_n1) );
  AND2X1 U6033_U2 ( .IN1(WX7224), .IN2(U6033_n1), .Q(WX7287) );
  INVX0 U6033_U1 ( .INP(n5534), .ZN(U6033_n1) );
  AND2X1 U6034_U2 ( .IN1(WX7222), .IN2(U6034_n1), .Q(WX7285) );
  INVX0 U6034_U1 ( .INP(n5534), .ZN(U6034_n1) );
  AND2X1 U6035_U2 ( .IN1(test_so60), .IN2(U6035_n1), .Q(WX7283) );
  INVX0 U6035_U1 ( .INP(n5534), .ZN(U6035_n1) );
  AND2X1 U6036_U2 ( .IN1(WX7218), .IN2(U6036_n1), .Q(WX7281) );
  INVX0 U6036_U1 ( .INP(n5534), .ZN(U6036_n1) );
  AND2X1 U6037_U2 ( .IN1(WX7216), .IN2(U6037_n1), .Q(WX7279) );
  INVX0 U6037_U1 ( .INP(n5535), .ZN(U6037_n1) );
  AND2X1 U6038_U2 ( .IN1(WX7214), .IN2(U6038_n1), .Q(WX7277) );
  INVX0 U6038_U1 ( .INP(n5535), .ZN(U6038_n1) );
  AND2X1 U6039_U2 ( .IN1(WX7212), .IN2(U6039_n1), .Q(WX7275) );
  INVX0 U6039_U1 ( .INP(n5535), .ZN(U6039_n1) );
  AND2X1 U6040_U2 ( .IN1(WX7210), .IN2(U6040_n1), .Q(WX7273) );
  INVX0 U6040_U1 ( .INP(n5535), .ZN(U6040_n1) );
  AND2X1 U6041_U2 ( .IN1(WX7208), .IN2(U6041_n1), .Q(WX7271) );
  INVX0 U6041_U1 ( .INP(n5535), .ZN(U6041_n1) );
  AND2X1 U6042_U2 ( .IN1(WX7206), .IN2(U6042_n1), .Q(WX7269) );
  INVX0 U6042_U1 ( .INP(n5535), .ZN(U6042_n1) );
  AND2X1 U6043_U2 ( .IN1(WX7204), .IN2(U6043_n1), .Q(WX7267) );
  INVX0 U6043_U1 ( .INP(n5535), .ZN(U6043_n1) );
  AND2X1 U6044_U2 ( .IN1(WX7202), .IN2(U6044_n1), .Q(WX7265) );
  INVX0 U6044_U1 ( .INP(n5535), .ZN(U6044_n1) );
  AND2X1 U6045_U2 ( .IN1(WX7200), .IN2(U6045_n1), .Q(WX7263) );
  INVX0 U6045_U1 ( .INP(n5535), .ZN(U6045_n1) );
  AND2X1 U6046_U2 ( .IN1(WX7198), .IN2(U6046_n1), .Q(WX7261) );
  INVX0 U6046_U1 ( .INP(n5535), .ZN(U6046_n1) );
  AND2X1 U6047_U2 ( .IN1(WX7196), .IN2(U6047_n1), .Q(WX7259) );
  INVX0 U6047_U1 ( .INP(n5535), .ZN(U6047_n1) );
  AND2X1 U6048_U2 ( .IN1(WX7194), .IN2(U6048_n1), .Q(WX7257) );
  INVX0 U6048_U1 ( .INP(n5535), .ZN(U6048_n1) );
  AND2X1 U6049_U2 ( .IN1(WX7192), .IN2(U6049_n1), .Q(WX7255) );
  INVX0 U6049_U1 ( .INP(n5535), .ZN(U6049_n1) );
  AND2X1 U6050_U2 ( .IN1(WX7190), .IN2(U6050_n1), .Q(WX7253) );
  INVX0 U6050_U1 ( .INP(n5535), .ZN(U6050_n1) );
  AND2X1 U6051_U2 ( .IN1(WX7188), .IN2(U6051_n1), .Q(WX7251) );
  INVX0 U6051_U1 ( .INP(n5536), .ZN(U6051_n1) );
  AND2X1 U6052_U2 ( .IN1(test_so59), .IN2(U6052_n1), .Q(WX7249) );
  INVX0 U6052_U1 ( .INP(n5536), .ZN(U6052_n1) );
  AND2X1 U6053_U2 ( .IN1(WX7184), .IN2(U6053_n1), .Q(WX7247) );
  INVX0 U6053_U1 ( .INP(n5536), .ZN(U6053_n1) );
  AND2X1 U6054_U2 ( .IN1(WX7182), .IN2(U6054_n1), .Q(WX7245) );
  INVX0 U6054_U1 ( .INP(n5536), .ZN(U6054_n1) );
  AND2X1 U6055_U2 ( .IN1(WX7180), .IN2(U6055_n1), .Q(WX7243) );
  INVX0 U6055_U1 ( .INP(n5536), .ZN(U6055_n1) );
  AND2X1 U6056_U2 ( .IN1(WX7178), .IN2(U6056_n1), .Q(WX7241) );
  INVX0 U6056_U1 ( .INP(n5536), .ZN(U6056_n1) );
  AND2X1 U6057_U2 ( .IN1(WX7176), .IN2(U6057_n1), .Q(WX7239) );
  INVX0 U6057_U1 ( .INP(n5536), .ZN(U6057_n1) );
  AND2X1 U6058_U2 ( .IN1(WX7174), .IN2(U6058_n1), .Q(WX7237) );
  INVX0 U6058_U1 ( .INP(n5536), .ZN(U6058_n1) );
  AND2X1 U6059_U2 ( .IN1(WX7172), .IN2(U6059_n1), .Q(WX7235) );
  INVX0 U6059_U1 ( .INP(n5536), .ZN(U6059_n1) );
  AND2X1 U6060_U2 ( .IN1(WX7170), .IN2(U6060_n1), .Q(WX7233) );
  INVX0 U6060_U1 ( .INP(n5536), .ZN(U6060_n1) );
  AND2X1 U6061_U2 ( .IN1(WX7168), .IN2(U6061_n1), .Q(WX7231) );
  INVX0 U6061_U1 ( .INP(n5536), .ZN(U6061_n1) );
  AND2X1 U6062_U2 ( .IN1(WX7166), .IN2(U6062_n1), .Q(WX7229) );
  INVX0 U6062_U1 ( .INP(n5536), .ZN(U6062_n1) );
  AND2X1 U6063_U2 ( .IN1(WX7164), .IN2(U6063_n1), .Q(WX7227) );
  INVX0 U6063_U1 ( .INP(n5536), .ZN(U6063_n1) );
  AND2X1 U6064_U2 ( .IN1(WX7162), .IN2(U6064_n1), .Q(WX7225) );
  INVX0 U6064_U1 ( .INP(n5537), .ZN(U6064_n1) );
  AND2X1 U6065_U2 ( .IN1(WX7160), .IN2(U6065_n1), .Q(WX7223) );
  INVX0 U6065_U1 ( .INP(n5537), .ZN(U6065_n1) );
  AND2X1 U6066_U2 ( .IN1(WX7158), .IN2(U6066_n1), .Q(WX7221) );
  INVX0 U6066_U1 ( .INP(n5537), .ZN(U6066_n1) );
  AND2X1 U6067_U2 ( .IN1(WX7156), .IN2(U6067_n1), .Q(WX7219) );
  INVX0 U6067_U1 ( .INP(n5537), .ZN(U6067_n1) );
  AND2X1 U6068_U2 ( .IN1(WX7154), .IN2(U6068_n1), .Q(WX7217) );
  INVX0 U6068_U1 ( .INP(n5537), .ZN(U6068_n1) );
  AND2X1 U6069_U2 ( .IN1(test_so58), .IN2(U6069_n1), .Q(WX7215) );
  INVX0 U6069_U1 ( .INP(n5537), .ZN(U6069_n1) );
  AND2X1 U6070_U2 ( .IN1(WX7150), .IN2(U6070_n1), .Q(WX7213) );
  INVX0 U6070_U1 ( .INP(n5537), .ZN(U6070_n1) );
  AND2X1 U6071_U2 ( .IN1(WX7148), .IN2(U6071_n1), .Q(WX7211) );
  INVX0 U6071_U1 ( .INP(n5537), .ZN(U6071_n1) );
  AND2X1 U6072_U2 ( .IN1(WX7146), .IN2(U6072_n1), .Q(WX7209) );
  INVX0 U6072_U1 ( .INP(n5537), .ZN(U6072_n1) );
  AND2X1 U6073_U2 ( .IN1(WX7144), .IN2(U6073_n1), .Q(WX7207) );
  INVX0 U6073_U1 ( .INP(n5537), .ZN(U6073_n1) );
  AND2X1 U6074_U2 ( .IN1(WX7142), .IN2(U6074_n1), .Q(WX7205) );
  INVX0 U6074_U1 ( .INP(n5537), .ZN(U6074_n1) );
  AND2X1 U6075_U2 ( .IN1(WX6007), .IN2(U6075_n1), .Q(WX6070) );
  INVX0 U6075_U1 ( .INP(n5537), .ZN(U6075_n1) );
  AND2X1 U6076_U2 ( .IN1(test_so51), .IN2(U6076_n1), .Q(WX6068) );
  INVX0 U6076_U1 ( .INP(n5537), .ZN(U6076_n1) );
  AND2X1 U6077_U2 ( .IN1(WX6003), .IN2(U6077_n1), .Q(WX6066) );
  INVX0 U6077_U1 ( .INP(n5537), .ZN(U6077_n1) );
  AND2X1 U6078_U2 ( .IN1(WX6001), .IN2(U6078_n1), .Q(WX6064) );
  INVX0 U6078_U1 ( .INP(n5538), .ZN(U6078_n1) );
  AND2X1 U6079_U2 ( .IN1(WX5999), .IN2(U6079_n1), .Q(WX6062) );
  INVX0 U6079_U1 ( .INP(n5538), .ZN(U6079_n1) );
  AND2X1 U6080_U2 ( .IN1(WX5997), .IN2(U6080_n1), .Q(WX6060) );
  INVX0 U6080_U1 ( .INP(n5538), .ZN(U6080_n1) );
  AND2X1 U6081_U2 ( .IN1(WX5995), .IN2(U6081_n1), .Q(WX6058) );
  INVX0 U6081_U1 ( .INP(n5538), .ZN(U6081_n1) );
  AND2X1 U6082_U2 ( .IN1(WX5993), .IN2(U6082_n1), .Q(WX6056) );
  INVX0 U6082_U1 ( .INP(n5538), .ZN(U6082_n1) );
  AND2X1 U6083_U2 ( .IN1(WX5991), .IN2(U6083_n1), .Q(WX6054) );
  INVX0 U6083_U1 ( .INP(n5538), .ZN(U6083_n1) );
  AND2X1 U6084_U2 ( .IN1(WX5989), .IN2(U6084_n1), .Q(WX6052) );
  INVX0 U6084_U1 ( .INP(n5538), .ZN(U6084_n1) );
  AND2X1 U6085_U2 ( .IN1(WX5987), .IN2(U6085_n1), .Q(WX6050) );
  INVX0 U6085_U1 ( .INP(n5538), .ZN(U6085_n1) );
  AND2X1 U6086_U2 ( .IN1(WX5985), .IN2(U6086_n1), .Q(WX6048) );
  INVX0 U6086_U1 ( .INP(n5538), .ZN(U6086_n1) );
  AND2X1 U6087_U2 ( .IN1(WX5983), .IN2(U6087_n1), .Q(WX6046) );
  INVX0 U6087_U1 ( .INP(n5538), .ZN(U6087_n1) );
  AND2X1 U6088_U2 ( .IN1(WX5981), .IN2(U6088_n1), .Q(WX6044) );
  INVX0 U6088_U1 ( .INP(n5538), .ZN(U6088_n1) );
  AND2X1 U6089_U2 ( .IN1(WX5979), .IN2(U6089_n1), .Q(WX6042) );
  INVX0 U6089_U1 ( .INP(n5538), .ZN(U6089_n1) );
  AND2X1 U6090_U2 ( .IN1(WX5977), .IN2(U6090_n1), .Q(WX6040) );
  INVX0 U6090_U1 ( .INP(n5538), .ZN(U6090_n1) );
  AND2X1 U6091_U2 ( .IN1(WX5975), .IN2(U6091_n1), .Q(WX6038) );
  INVX0 U6091_U1 ( .INP(n5538), .ZN(U6091_n1) );
  AND2X1 U6092_U2 ( .IN1(WX5973), .IN2(U6092_n1), .Q(WX6036) );
  INVX0 U6092_U1 ( .INP(n5539), .ZN(U6092_n1) );
  AND2X1 U6093_U2 ( .IN1(test_so50), .IN2(U6093_n1), .Q(WX6034) );
  INVX0 U6093_U1 ( .INP(n5539), .ZN(U6093_n1) );
  AND2X1 U6094_U2 ( .IN1(WX5969), .IN2(U6094_n1), .Q(WX6032) );
  INVX0 U6094_U1 ( .INP(n5539), .ZN(U6094_n1) );
  AND2X1 U6095_U2 ( .IN1(WX5967), .IN2(U6095_n1), .Q(WX6030) );
  INVX0 U6095_U1 ( .INP(n5539), .ZN(U6095_n1) );
  AND2X1 U6096_U2 ( .IN1(WX5965), .IN2(U6096_n1), .Q(WX6028) );
  INVX0 U6096_U1 ( .INP(n5539), .ZN(U6096_n1) );
  AND2X1 U6097_U2 ( .IN1(WX5963), .IN2(U6097_n1), .Q(WX6026) );
  INVX0 U6097_U1 ( .INP(n5539), .ZN(U6097_n1) );
  AND2X1 U6098_U2 ( .IN1(WX5961), .IN2(U6098_n1), .Q(WX6024) );
  INVX0 U6098_U1 ( .INP(n5539), .ZN(U6098_n1) );
  AND2X1 U6099_U2 ( .IN1(WX5959), .IN2(U6099_n1), .Q(WX6022) );
  INVX0 U6099_U1 ( .INP(n5539), .ZN(U6099_n1) );
  AND2X1 U6100_U2 ( .IN1(WX5957), .IN2(U6100_n1), .Q(WX6020) );
  INVX0 U6100_U1 ( .INP(n5539), .ZN(U6100_n1) );
  AND2X1 U6101_U2 ( .IN1(WX5955), .IN2(U6101_n1), .Q(WX6018) );
  INVX0 U6101_U1 ( .INP(n5539), .ZN(U6101_n1) );
  AND2X1 U6102_U2 ( .IN1(WX5953), .IN2(U6102_n1), .Q(WX6016) );
  INVX0 U6102_U1 ( .INP(n5539), .ZN(U6102_n1) );
  AND2X1 U6103_U2 ( .IN1(WX5951), .IN2(U6103_n1), .Q(WX6014) );
  INVX0 U6103_U1 ( .INP(n5539), .ZN(U6103_n1) );
  AND2X1 U6104_U2 ( .IN1(WX5949), .IN2(U6104_n1), .Q(WX6012) );
  INVX0 U6104_U1 ( .INP(n5539), .ZN(U6104_n1) );
  AND2X1 U6105_U2 ( .IN1(WX5947), .IN2(U6105_n1), .Q(WX6010) );
  INVX0 U6105_U1 ( .INP(n5539), .ZN(U6105_n1) );
  AND2X1 U6106_U2 ( .IN1(WX5945), .IN2(U6106_n1), .Q(WX6008) );
  INVX0 U6106_U1 ( .INP(n5540), .ZN(U6106_n1) );
  AND2X1 U6107_U2 ( .IN1(WX5943), .IN2(U6107_n1), .Q(WX6006) );
  INVX0 U6107_U1 ( .INP(n5540), .ZN(U6107_n1) );
  AND2X1 U6108_U2 ( .IN1(WX5941), .IN2(U6108_n1), .Q(WX6004) );
  INVX0 U6108_U1 ( .INP(n5540), .ZN(U6108_n1) );
  AND2X1 U6109_U2 ( .IN1(WX5929), .IN2(U6109_n1), .Q(WX5992) );
  INVX0 U6109_U1 ( .INP(n5540), .ZN(U6109_n1) );
  AND2X1 U6110_U2 ( .IN1(WX5927), .IN2(U6110_n1), .Q(WX5990) );
  INVX0 U6110_U1 ( .INP(n5540), .ZN(U6110_n1) );
  AND2X1 U6111_U2 ( .IN1(WX5925), .IN2(U6111_n1), .Q(WX5988) );
  INVX0 U6111_U1 ( .INP(n5540), .ZN(U6111_n1) );
  AND2X1 U6112_U2 ( .IN1(WX5923), .IN2(U6112_n1), .Q(WX5986) );
  INVX0 U6112_U1 ( .INP(n5540), .ZN(U6112_n1) );
  AND2X1 U6113_U2 ( .IN1(WX5921), .IN2(U6113_n1), .Q(WX5984) );
  INVX0 U6113_U1 ( .INP(n5540), .ZN(U6113_n1) );
  AND2X1 U6114_U2 ( .IN1(WX5919), .IN2(U6114_n1), .Q(WX5982) );
  INVX0 U6114_U1 ( .INP(n5540), .ZN(U6114_n1) );
  AND2X1 U6115_U2 ( .IN1(WX5917), .IN2(U6115_n1), .Q(WX5980) );
  INVX0 U6115_U1 ( .INP(n5540), .ZN(U6115_n1) );
  AND2X1 U6116_U2 ( .IN1(WX5915), .IN2(U6116_n1), .Q(WX5978) );
  INVX0 U6116_U1 ( .INP(n5540), .ZN(U6116_n1) );
  AND2X1 U6117_U2 ( .IN1(WX5913), .IN2(U6117_n1), .Q(WX5976) );
  INVX0 U6117_U1 ( .INP(n5540), .ZN(U6117_n1) );
  AND2X1 U6118_U2 ( .IN1(WX5911), .IN2(U6118_n1), .Q(WX5974) );
  INVX0 U6118_U1 ( .INP(n5540), .ZN(U6118_n1) );
  AND2X1 U6119_U2 ( .IN1(WX5909), .IN2(U6119_n1), .Q(WX5972) );
  INVX0 U6119_U1 ( .INP(n5540), .ZN(U6119_n1) );
  AND2X1 U6120_U2 ( .IN1(WX5907), .IN2(U6120_n1), .Q(WX5970) );
  INVX0 U6120_U1 ( .INP(n5541), .ZN(U6120_n1) );
  AND2X1 U6121_U2 ( .IN1(WX5905), .IN2(U6121_n1), .Q(WX5968) );
  INVX0 U6121_U1 ( .INP(n5541), .ZN(U6121_n1) );
  AND2X1 U6122_U2 ( .IN1(test_so48), .IN2(U6122_n1), .Q(WX5966) );
  INVX0 U6122_U1 ( .INP(n5541), .ZN(U6122_n1) );
  AND2X1 U6123_U2 ( .IN1(WX5901), .IN2(U6123_n1), .Q(WX5964) );
  INVX0 U6123_U1 ( .INP(n5541), .ZN(U6123_n1) );
  AND2X1 U6124_U2 ( .IN1(WX5899), .IN2(U6124_n1), .Q(WX5962) );
  INVX0 U6124_U1 ( .INP(n5541), .ZN(U6124_n1) );
  AND2X1 U6125_U2 ( .IN1(WX5897), .IN2(U6125_n1), .Q(WX5960) );
  INVX0 U6125_U1 ( .INP(n5541), .ZN(U6125_n1) );
  AND2X1 U6126_U2 ( .IN1(WX5895), .IN2(U6126_n1), .Q(WX5958) );
  INVX0 U6126_U1 ( .INP(n5541), .ZN(U6126_n1) );
  AND2X1 U6127_U2 ( .IN1(WX5893), .IN2(U6127_n1), .Q(WX5956) );
  INVX0 U6127_U1 ( .INP(n5541), .ZN(U6127_n1) );
  AND2X1 U6128_U2 ( .IN1(WX5891), .IN2(U6128_n1), .Q(WX5954) );
  INVX0 U6128_U1 ( .INP(n5541), .ZN(U6128_n1) );
  AND2X1 U6129_U2 ( .IN1(WX5889), .IN2(U6129_n1), .Q(WX5952) );
  INVX0 U6129_U1 ( .INP(n5541), .ZN(U6129_n1) );
  AND2X1 U6130_U2 ( .IN1(WX5887), .IN2(U6130_n1), .Q(WX5950) );
  INVX0 U6130_U1 ( .INP(n5541), .ZN(U6130_n1) );
  AND2X1 U6131_U2 ( .IN1(WX5885), .IN2(U6131_n1), .Q(WX5948) );
  INVX0 U6131_U1 ( .INP(n5541), .ZN(U6131_n1) );
  AND2X1 U6132_U2 ( .IN1(WX5883), .IN2(U6132_n1), .Q(WX5946) );
  INVX0 U6132_U1 ( .INP(n5527), .ZN(U6132_n1) );
  AND2X1 U6133_U2 ( .IN1(WX5881), .IN2(U6133_n1), .Q(WX5944) );
  INVX0 U6133_U1 ( .INP(n5522), .ZN(U6133_n1) );
  AND2X1 U6134_U2 ( .IN1(WX5879), .IN2(U6134_n1), .Q(WX5942) );
  INVX0 U6134_U1 ( .INP(n5522), .ZN(U6134_n1) );
  AND2X1 U6135_U2 ( .IN1(WX5877), .IN2(U6135_n1), .Q(WX5940) );
  INVX0 U6135_U1 ( .INP(n5522), .ZN(U6135_n1) );
  AND2X1 U6136_U2 ( .IN1(WX5875), .IN2(U6136_n1), .Q(WX5938) );
  INVX0 U6136_U1 ( .INP(n5522), .ZN(U6136_n1) );
  AND2X1 U6137_U2 ( .IN1(WX5873), .IN2(U6137_n1), .Q(WX5936) );
  INVX0 U6137_U1 ( .INP(n5522), .ZN(U6137_n1) );
  AND2X1 U6138_U2 ( .IN1(WX5871), .IN2(U6138_n1), .Q(WX5934) );
  INVX0 U6138_U1 ( .INP(n5522), .ZN(U6138_n1) );
  AND2X1 U6139_U2 ( .IN1(test_so47), .IN2(U6139_n1), .Q(WX5932) );
  INVX0 U6139_U1 ( .INP(n5522), .ZN(U6139_n1) );
  AND2X1 U6140_U2 ( .IN1(WX5867), .IN2(U6140_n1), .Q(WX5930) );
  INVX0 U6140_U1 ( .INP(n5522), .ZN(U6140_n1) );
  AND2X1 U6141_U2 ( .IN1(WX5865), .IN2(U6141_n1), .Q(WX5928) );
  INVX0 U6141_U1 ( .INP(n5522), .ZN(U6141_n1) );
  AND2X1 U6142_U2 ( .IN1(WX5863), .IN2(U6142_n1), .Q(WX5926) );
  INVX0 U6142_U1 ( .INP(n5522), .ZN(U6142_n1) );
  AND2X1 U6143_U2 ( .IN1(WX5861), .IN2(U6143_n1), .Q(WX5924) );
  INVX0 U6143_U1 ( .INP(n5522), .ZN(U6143_n1) );
  AND2X1 U6144_U2 ( .IN1(WX5859), .IN2(U6144_n1), .Q(WX5922) );
  INVX0 U6144_U1 ( .INP(n5522), .ZN(U6144_n1) );
  AND2X1 U6145_U2 ( .IN1(WX5857), .IN2(U6145_n1), .Q(WX5920) );
  INVX0 U6145_U1 ( .INP(n5523), .ZN(U6145_n1) );
  AND2X1 U6146_U2 ( .IN1(WX5855), .IN2(U6146_n1), .Q(WX5918) );
  INVX0 U6146_U1 ( .INP(n5523), .ZN(U6146_n1) );
  AND2X1 U6147_U2 ( .IN1(WX5853), .IN2(U6147_n1), .Q(WX5916) );
  INVX0 U6147_U1 ( .INP(n5523), .ZN(U6147_n1) );
  AND2X1 U6148_U2 ( .IN1(WX5851), .IN2(U6148_n1), .Q(WX5914) );
  INVX0 U6148_U1 ( .INP(n5523), .ZN(U6148_n1) );
  AND2X1 U6149_U2 ( .IN1(WX5849), .IN2(U6149_n1), .Q(WX5912) );
  INVX0 U6149_U1 ( .INP(n5523), .ZN(U6149_n1) );
  AND2X1 U6150_U2 ( .IN1(WX4714), .IN2(U6150_n1), .Q(WX4777) );
  INVX0 U6150_U1 ( .INP(n5523), .ZN(U6150_n1) );
  AND2X1 U6151_U2 ( .IN1(WX4712), .IN2(U6151_n1), .Q(WX4775) );
  INVX0 U6151_U1 ( .INP(n5523), .ZN(U6151_n1) );
  AND2X1 U6152_U2 ( .IN1(WX4710), .IN2(U6152_n1), .Q(WX4773) );
  INVX0 U6152_U1 ( .INP(n5523), .ZN(U6152_n1) );
  AND2X1 U6153_U2 ( .IN1(WX4708), .IN2(U6153_n1), .Q(WX4771) );
  INVX0 U6153_U1 ( .INP(n5523), .ZN(U6153_n1) );
  AND2X1 U6154_U2 ( .IN1(WX4706), .IN2(U6154_n1), .Q(WX4769) );
  INVX0 U6154_U1 ( .INP(n5523), .ZN(U6154_n1) );
  AND2X1 U6155_U2 ( .IN1(WX4704), .IN2(U6155_n1), .Q(WX4767) );
  INVX0 U6155_U1 ( .INP(n5523), .ZN(U6155_n1) );
  AND2X1 U6156_U2 ( .IN1(WX4702), .IN2(U6156_n1), .Q(WX4765) );
  INVX0 U6156_U1 ( .INP(n5523), .ZN(U6156_n1) );
  AND2X1 U6157_U2 ( .IN1(WX4700), .IN2(U6157_n1), .Q(WX4763) );
  INVX0 U6157_U1 ( .INP(n5523), .ZN(U6157_n1) );
  AND2X1 U6158_U2 ( .IN1(WX4698), .IN2(U6158_n1), .Q(WX4761) );
  INVX0 U6158_U1 ( .INP(n5523), .ZN(U6158_n1) );
  AND2X1 U6159_U2 ( .IN1(WX4696), .IN2(U6159_n1), .Q(WX4759) );
  INVX0 U6159_U1 ( .INP(n5524), .ZN(U6159_n1) );
  AND2X1 U6160_U2 ( .IN1(WX4694), .IN2(U6160_n1), .Q(WX4757) );
  INVX0 U6160_U1 ( .INP(n5524), .ZN(U6160_n1) );
  AND2X1 U6161_U2 ( .IN1(WX4692), .IN2(U6161_n1), .Q(WX4755) );
  INVX0 U6161_U1 ( .INP(n5524), .ZN(U6161_n1) );
  AND2X1 U6162_U2 ( .IN1(WX4690), .IN2(U6162_n1), .Q(WX4753) );
  INVX0 U6162_U1 ( .INP(n5524), .ZN(U6162_n1) );
  AND2X1 U6163_U2 ( .IN1(test_so39), .IN2(U6163_n1), .Q(WX4751) );
  INVX0 U6163_U1 ( .INP(n5524), .ZN(U6163_n1) );
  AND2X1 U6164_U2 ( .IN1(WX4686), .IN2(U6164_n1), .Q(WX4749) );
  INVX0 U6164_U1 ( .INP(n5524), .ZN(U6164_n1) );
  AND2X1 U6165_U2 ( .IN1(WX4684), .IN2(U6165_n1), .Q(WX4747) );
  INVX0 U6165_U1 ( .INP(n5524), .ZN(U6165_n1) );
  AND2X1 U6166_U2 ( .IN1(WX4682), .IN2(U6166_n1), .Q(WX4745) );
  INVX0 U6166_U1 ( .INP(n5524), .ZN(U6166_n1) );
  AND2X1 U6167_U2 ( .IN1(WX4680), .IN2(U6167_n1), .Q(WX4743) );
  INVX0 U6167_U1 ( .INP(n5524), .ZN(U6167_n1) );
  AND2X1 U6168_U2 ( .IN1(WX4678), .IN2(U6168_n1), .Q(WX4741) );
  INVX0 U6168_U1 ( .INP(n5524), .ZN(U6168_n1) );
  AND2X1 U6169_U2 ( .IN1(WX4676), .IN2(U6169_n1), .Q(WX4739) );
  INVX0 U6169_U1 ( .INP(n5524), .ZN(U6169_n1) );
  AND2X1 U6170_U2 ( .IN1(WX4674), .IN2(U6170_n1), .Q(WX4737) );
  INVX0 U6170_U1 ( .INP(n5524), .ZN(U6170_n1) );
  AND2X1 U6171_U2 ( .IN1(WX4672), .IN2(U6171_n1), .Q(WX4735) );
  INVX0 U6171_U1 ( .INP(n5524), .ZN(U6171_n1) );
  AND2X1 U6172_U2 ( .IN1(WX4670), .IN2(U6172_n1), .Q(WX4733) );
  INVX0 U6172_U1 ( .INP(n5524), .ZN(U6172_n1) );
  AND2X1 U6173_U2 ( .IN1(WX4668), .IN2(U6173_n1), .Q(WX4731) );
  INVX0 U6173_U1 ( .INP(n5525), .ZN(U6173_n1) );
  AND2X1 U6174_U2 ( .IN1(WX4666), .IN2(U6174_n1), .Q(WX4729) );
  INVX0 U6174_U1 ( .INP(n5525), .ZN(U6174_n1) );
  AND2X1 U6175_U2 ( .IN1(WX4664), .IN2(U6175_n1), .Q(WX4727) );
  INVX0 U6175_U1 ( .INP(n5525), .ZN(U6175_n1) );
  AND2X1 U6176_U2 ( .IN1(WX4662), .IN2(U6176_n1), .Q(WX4725) );
  INVX0 U6176_U1 ( .INP(n5525), .ZN(U6176_n1) );
  AND2X1 U6177_U2 ( .IN1(WX4660), .IN2(U6177_n1), .Q(WX4723) );
  INVX0 U6177_U1 ( .INP(n5525), .ZN(U6177_n1) );
  AND2X1 U6178_U2 ( .IN1(WX4658), .IN2(U6178_n1), .Q(WX4721) );
  INVX0 U6178_U1 ( .INP(n5525), .ZN(U6178_n1) );
  AND2X1 U6179_U2 ( .IN1(WX4656), .IN2(U6179_n1), .Q(WX4719) );
  INVX0 U6179_U1 ( .INP(n5525), .ZN(U6179_n1) );
  AND2X1 U6180_U2 ( .IN1(test_so38), .IN2(U6180_n1), .Q(WX4717) );
  INVX0 U6180_U1 ( .INP(n5525), .ZN(U6180_n1) );
  AND2X1 U6181_U2 ( .IN1(WX4652), .IN2(U6181_n1), .Q(WX4715) );
  INVX0 U6181_U1 ( .INP(n5525), .ZN(U6181_n1) );
  AND2X1 U6182_U2 ( .IN1(WX4650), .IN2(U6182_n1), .Q(WX4713) );
  INVX0 U6182_U1 ( .INP(n5525), .ZN(U6182_n1) );
  AND2X1 U6183_U2 ( .IN1(WX4648), .IN2(U6183_n1), .Q(WX4711) );
  INVX0 U6183_U1 ( .INP(n5525), .ZN(U6183_n1) );
  AND2X1 U6184_U2 ( .IN1(WX4646), .IN2(U6184_n1), .Q(WX4709) );
  INVX0 U6184_U1 ( .INP(n5525), .ZN(U6184_n1) );
  AND2X1 U6185_U2 ( .IN1(WX4644), .IN2(U6185_n1), .Q(WX4707) );
  INVX0 U6185_U1 ( .INP(n5525), .ZN(U6185_n1) );
  AND2X1 U6186_U2 ( .IN1(WX4642), .IN2(U6186_n1), .Q(WX4705) );
  INVX0 U6186_U1 ( .INP(n5525), .ZN(U6186_n1) );
  AND2X1 U6187_U2 ( .IN1(WX4640), .IN2(U6187_n1), .Q(WX4703) );
  INVX0 U6187_U1 ( .INP(n5526), .ZN(U6187_n1) );
  AND2X1 U6188_U2 ( .IN1(WX4638), .IN2(U6188_n1), .Q(WX4701) );
  INVX0 U6188_U1 ( .INP(n5526), .ZN(U6188_n1) );
  AND2X1 U6189_U2 ( .IN1(WX4636), .IN2(U6189_n1), .Q(WX4699) );
  INVX0 U6189_U1 ( .INP(n5526), .ZN(U6189_n1) );
  AND2X1 U6190_U2 ( .IN1(WX4634), .IN2(U6190_n1), .Q(WX4697) );
  INVX0 U6190_U1 ( .INP(n5526), .ZN(U6190_n1) );
  AND2X1 U6191_U2 ( .IN1(WX4632), .IN2(U6191_n1), .Q(WX4695) );
  INVX0 U6191_U1 ( .INP(n5526), .ZN(U6191_n1) );
  AND2X1 U6192_U2 ( .IN1(WX4630), .IN2(U6192_n1), .Q(WX4693) );
  INVX0 U6192_U1 ( .INP(n5526), .ZN(U6192_n1) );
  AND2X1 U6193_U2 ( .IN1(WX4628), .IN2(U6193_n1), .Q(WX4691) );
  INVX0 U6193_U1 ( .INP(n5526), .ZN(U6193_n1) );
  AND2X1 U6194_U2 ( .IN1(WX4626), .IN2(U6194_n1), .Q(WX4689) );
  INVX0 U6194_U1 ( .INP(n5526), .ZN(U6194_n1) );
  AND2X1 U6195_U2 ( .IN1(WX4624), .IN2(U6195_n1), .Q(WX4687) );
  INVX0 U6195_U1 ( .INP(n5526), .ZN(U6195_n1) );
  AND2X1 U6196_U2 ( .IN1(WX4622), .IN2(U6196_n1), .Q(WX4685) );
  INVX0 U6196_U1 ( .INP(n5526), .ZN(U6196_n1) );
  AND2X1 U6197_U2 ( .IN1(test_so37), .IN2(U6197_n1), .Q(WX4683) );
  INVX0 U6197_U1 ( .INP(n5526), .ZN(U6197_n1) );
  AND2X1 U6198_U2 ( .IN1(WX4618), .IN2(U6198_n1), .Q(WX4681) );
  INVX0 U6198_U1 ( .INP(n5526), .ZN(U6198_n1) );
  AND2X1 U6199_U2 ( .IN1(WX4616), .IN2(U6199_n1), .Q(WX4679) );
  INVX0 U6199_U1 ( .INP(n5526), .ZN(U6199_n1) );
  AND2X1 U6200_U2 ( .IN1(WX4614), .IN2(U6200_n1), .Q(WX4677) );
  INVX0 U6200_U1 ( .INP(n5526), .ZN(U6200_n1) );
  AND2X1 U6201_U2 ( .IN1(WX4612), .IN2(U6201_n1), .Q(WX4675) );
  INVX0 U6201_U1 ( .INP(n5527), .ZN(U6201_n1) );
  AND2X1 U6202_U2 ( .IN1(WX4610), .IN2(U6202_n1), .Q(WX4673) );
  INVX0 U6202_U1 ( .INP(n5527), .ZN(U6202_n1) );
  AND2X1 U6203_U2 ( .IN1(WX4608), .IN2(U6203_n1), .Q(WX4671) );
  INVX0 U6203_U1 ( .INP(n5527), .ZN(U6203_n1) );
  AND2X1 U6204_U2 ( .IN1(WX4606), .IN2(U6204_n1), .Q(WX4669) );
  INVX0 U6204_U1 ( .INP(n5527), .ZN(U6204_n1) );
  AND2X1 U6205_U2 ( .IN1(WX4604), .IN2(U6205_n1), .Q(WX4667) );
  INVX0 U6205_U1 ( .INP(n5527), .ZN(U6205_n1) );
  AND2X1 U6206_U2 ( .IN1(WX4602), .IN2(U6206_n1), .Q(WX4665) );
  INVX0 U6206_U1 ( .INP(n5527), .ZN(U6206_n1) );
  AND2X1 U6207_U2 ( .IN1(WX4600), .IN2(U6207_n1), .Q(WX4663) );
  INVX0 U6207_U1 ( .INP(n5527), .ZN(U6207_n1) );
  AND2X1 U6208_U2 ( .IN1(WX4598), .IN2(U6208_n1), .Q(WX4661) );
  INVX0 U6208_U1 ( .INP(n5527), .ZN(U6208_n1) );
  AND2X1 U6209_U2 ( .IN1(WX4596), .IN2(U6209_n1), .Q(WX4659) );
  INVX0 U6209_U1 ( .INP(n5527), .ZN(U6209_n1) );
  AND2X1 U6210_U2 ( .IN1(WX4594), .IN2(U6210_n1), .Q(WX4657) );
  INVX0 U6210_U1 ( .INP(n5527), .ZN(U6210_n1) );
  AND2X1 U6211_U2 ( .IN1(WX4592), .IN2(U6211_n1), .Q(WX4655) );
  INVX0 U6211_U1 ( .INP(n5527), .ZN(U6211_n1) );
  AND2X1 U6212_U2 ( .IN1(WX4590), .IN2(U6212_n1), .Q(WX4653) );
  INVX0 U6212_U1 ( .INP(n5527), .ZN(U6212_n1) );
  AND2X1 U6213_U2 ( .IN1(WX4588), .IN2(U6213_n1), .Q(WX4651) );
  INVX0 U6213_U1 ( .INP(n5527), .ZN(U6213_n1) );
  AND2X1 U6214_U2 ( .IN1(test_so36), .IN2(U6214_n1), .Q(WX4649) );
  INVX0 U6214_U1 ( .INP(n5528), .ZN(U6214_n1) );
  AND2X1 U6215_U2 ( .IN1(WX4584), .IN2(U6215_n1), .Q(WX4647) );
  INVX0 U6215_U1 ( .INP(n5528), .ZN(U6215_n1) );
  AND2X1 U6216_U2 ( .IN1(WX4582), .IN2(U6216_n1), .Q(WX4645) );
  INVX0 U6216_U1 ( .INP(n5528), .ZN(U6216_n1) );
  AND2X1 U6217_U2 ( .IN1(WX4580), .IN2(U6217_n1), .Q(WX4643) );
  INVX0 U6217_U1 ( .INP(n5528), .ZN(U6217_n1) );
  AND2X1 U6218_U2 ( .IN1(WX4578), .IN2(U6218_n1), .Q(WX4641) );
  INVX0 U6218_U1 ( .INP(n5528), .ZN(U6218_n1) );
  AND2X1 U6219_U2 ( .IN1(WX4576), .IN2(U6219_n1), .Q(WX4639) );
  INVX0 U6219_U1 ( .INP(n5528), .ZN(U6219_n1) );
  AND2X1 U6220_U2 ( .IN1(WX4574), .IN2(U6220_n1), .Q(WX4637) );
  INVX0 U6220_U1 ( .INP(n5528), .ZN(U6220_n1) );
  AND2X1 U6221_U2 ( .IN1(WX4572), .IN2(U6221_n1), .Q(WX4635) );
  INVX0 U6221_U1 ( .INP(n5528), .ZN(U6221_n1) );
  AND2X1 U6222_U2 ( .IN1(WX4570), .IN2(U6222_n1), .Q(WX4633) );
  INVX0 U6222_U1 ( .INP(n5528), .ZN(U6222_n1) );
  AND2X1 U6223_U2 ( .IN1(WX4568), .IN2(U6223_n1), .Q(WX4631) );
  INVX0 U6223_U1 ( .INP(n5528), .ZN(U6223_n1) );
  AND2X1 U6224_U2 ( .IN1(WX4566), .IN2(U6224_n1), .Q(WX4629) );
  INVX0 U6224_U1 ( .INP(n5528), .ZN(U6224_n1) );
  AND2X1 U6225_U2 ( .IN1(WX4564), .IN2(U6225_n1), .Q(WX4627) );
  INVX0 U6225_U1 ( .INP(n5528), .ZN(U6225_n1) );
  AND2X1 U6226_U2 ( .IN1(WX4562), .IN2(U6226_n1), .Q(WX4625) );
  INVX0 U6226_U1 ( .INP(n5528), .ZN(U6226_n1) );
  AND2X1 U6227_U2 ( .IN1(WX4560), .IN2(U6227_n1), .Q(WX4623) );
  INVX0 U6227_U1 ( .INP(n5528), .ZN(U6227_n1) );
  AND2X1 U6228_U2 ( .IN1(WX4558), .IN2(U6228_n1), .Q(WX4621) );
  INVX0 U6228_U1 ( .INP(n5529), .ZN(U6228_n1) );
  AND2X1 U6229_U2 ( .IN1(WX4556), .IN2(U6229_n1), .Q(WX4619) );
  INVX0 U6229_U1 ( .INP(n5529), .ZN(U6229_n1) );
  AND2X1 U6230_U2 ( .IN1(WX3421), .IN2(U6230_n1), .Q(WX3484) );
  INVX0 U6230_U1 ( .INP(n5529), .ZN(U6230_n1) );
  AND2X1 U6231_U2 ( .IN1(WX3419), .IN2(U6231_n1), .Q(WX3482) );
  INVX0 U6231_U1 ( .INP(n5529), .ZN(U6231_n1) );
  AND2X1 U6232_U2 ( .IN1(WX3417), .IN2(U6232_n1), .Q(WX3480) );
  INVX0 U6232_U1 ( .INP(n5529), .ZN(U6232_n1) );
  AND2X1 U6233_U2 ( .IN1(WX3415), .IN2(U6233_n1), .Q(WX3478) );
  INVX0 U6233_U1 ( .INP(n5529), .ZN(U6233_n1) );
  AND2X1 U6234_U2 ( .IN1(WX3413), .IN2(U6234_n1), .Q(WX3476) );
  INVX0 U6234_U1 ( .INP(n5529), .ZN(U6234_n1) );
  AND2X1 U6235_U2 ( .IN1(WX3411), .IN2(U6235_n1), .Q(WX3474) );
  INVX0 U6235_U1 ( .INP(n5529), .ZN(U6235_n1) );
  AND2X1 U6236_U2 ( .IN1(WX3409), .IN2(U6236_n1), .Q(WX3472) );
  INVX0 U6236_U1 ( .INP(n5529), .ZN(U6236_n1) );
  AND2X1 U6237_U2 ( .IN1(WX3407), .IN2(U6237_n1), .Q(WX3470) );
  INVX0 U6237_U1 ( .INP(n5529), .ZN(U6237_n1) );
  AND2X1 U6238_U2 ( .IN1(test_so28), .IN2(U6238_n1), .Q(WX3468) );
  INVX0 U6238_U1 ( .INP(n5529), .ZN(U6238_n1) );
  AND2X1 U6239_U2 ( .IN1(WX3403), .IN2(U6239_n1), .Q(WX3466) );
  INVX0 U6239_U1 ( .INP(n5529), .ZN(U6239_n1) );
  AND2X1 U6240_U2 ( .IN1(WX3401), .IN2(U6240_n1), .Q(WX3464) );
  INVX0 U6240_U1 ( .INP(n5529), .ZN(U6240_n1) );
  AND2X1 U6241_U2 ( .IN1(WX3399), .IN2(U6241_n1), .Q(WX3462) );
  INVX0 U6241_U1 ( .INP(n5529), .ZN(U6241_n1) );
  AND2X1 U6242_U2 ( .IN1(WX3397), .IN2(U6242_n1), .Q(WX3460) );
  INVX0 U6242_U1 ( .INP(n5530), .ZN(U6242_n1) );
  AND2X1 U6243_U2 ( .IN1(WX3395), .IN2(U6243_n1), .Q(WX3458) );
  INVX0 U6243_U1 ( .INP(n5530), .ZN(U6243_n1) );
  AND2X1 U6244_U2 ( .IN1(WX3393), .IN2(U6244_n1), .Q(WX3456) );
  INVX0 U6244_U1 ( .INP(n5530), .ZN(U6244_n1) );
  AND2X1 U6245_U2 ( .IN1(WX3391), .IN2(U6245_n1), .Q(WX3454) );
  INVX0 U6245_U1 ( .INP(n5530), .ZN(U6245_n1) );
  AND2X1 U6246_U2 ( .IN1(WX3389), .IN2(U6246_n1), .Q(WX3452) );
  INVX0 U6246_U1 ( .INP(n5530), .ZN(U6246_n1) );
  AND2X1 U6247_U2 ( .IN1(WX3387), .IN2(U6247_n1), .Q(WX3450) );
  INVX0 U6247_U1 ( .INP(n5530), .ZN(U6247_n1) );
  AND2X1 U6248_U2 ( .IN1(WX3385), .IN2(U6248_n1), .Q(WX3448) );
  INVX0 U6248_U1 ( .INP(n5530), .ZN(U6248_n1) );
  AND2X1 U6249_U2 ( .IN1(WX3383), .IN2(U6249_n1), .Q(WX3446) );
  INVX0 U6249_U1 ( .INP(n5530), .ZN(U6249_n1) );
  AND2X1 U6250_U2 ( .IN1(WX3381), .IN2(U6250_n1), .Q(WX3444) );
  INVX0 U6250_U1 ( .INP(n5530), .ZN(U6250_n1) );
  AND2X1 U6251_U2 ( .IN1(WX3379), .IN2(U6251_n1), .Q(WX3442) );
  INVX0 U6251_U1 ( .INP(n5530), .ZN(U6251_n1) );
  AND2X1 U6252_U2 ( .IN1(WX3377), .IN2(U6252_n1), .Q(WX3440) );
  INVX0 U6252_U1 ( .INP(n5530), .ZN(U6252_n1) );
  AND2X1 U6253_U2 ( .IN1(WX3375), .IN2(U6253_n1), .Q(WX3438) );
  INVX0 U6253_U1 ( .INP(n5530), .ZN(U6253_n1) );
  AND2X1 U6254_U2 ( .IN1(WX3373), .IN2(U6254_n1), .Q(WX3436) );
  INVX0 U6254_U1 ( .INP(n5530), .ZN(U6254_n1) );
  AND2X1 U6255_U2 ( .IN1(WX3371), .IN2(U6255_n1), .Q(WX3434) );
  INVX0 U6255_U1 ( .INP(n5530), .ZN(U6255_n1) );
  AND2X1 U6256_U2 ( .IN1(test_so27), .IN2(U6256_n1), .Q(WX3432) );
  INVX0 U6256_U1 ( .INP(n5531), .ZN(U6256_n1) );
  AND2X1 U6257_U2 ( .IN1(WX3367), .IN2(U6257_n1), .Q(WX3430) );
  INVX0 U6257_U1 ( .INP(n5531), .ZN(U6257_n1) );
  AND2X1 U6258_U2 ( .IN1(WX3365), .IN2(U6258_n1), .Q(WX3428) );
  INVX0 U6258_U1 ( .INP(n5531), .ZN(U6258_n1) );
  AND2X1 U6259_U2 ( .IN1(WX3363), .IN2(U6259_n1), .Q(WX3426) );
  INVX0 U6259_U1 ( .INP(n5531), .ZN(U6259_n1) );
  AND2X1 U6260_U2 ( .IN1(WX3361), .IN2(U6260_n1), .Q(WX3424) );
  INVX0 U6260_U1 ( .INP(n5531), .ZN(U6260_n1) );
  AND2X1 U6261_U2 ( .IN1(WX3359), .IN2(U6261_n1), .Q(WX3422) );
  INVX0 U6261_U1 ( .INP(n5531), .ZN(U6261_n1) );
  AND2X1 U6262_U2 ( .IN1(WX3357), .IN2(U6262_n1), .Q(WX3420) );
  INVX0 U6262_U1 ( .INP(n5531), .ZN(U6262_n1) );
  AND2X1 U6263_U2 ( .IN1(WX3355), .IN2(U6263_n1), .Q(WX3418) );
  INVX0 U6263_U1 ( .INP(n5531), .ZN(U6263_n1) );
  AND2X1 U6264_U2 ( .IN1(WX3353), .IN2(U6264_n1), .Q(WX3416) );
  INVX0 U6264_U1 ( .INP(n5531), .ZN(U6264_n1) );
  AND2X1 U6265_U2 ( .IN1(WX3351), .IN2(U6265_n1), .Q(WX3414) );
  INVX0 U6265_U1 ( .INP(n5531), .ZN(U6265_n1) );
  AND2X1 U6266_U2 ( .IN1(WX3349), .IN2(U6266_n1), .Q(WX3412) );
  INVX0 U6266_U1 ( .INP(n5531), .ZN(U6266_n1) );
  AND2X1 U6267_U2 ( .IN1(WX3347), .IN2(U6267_n1), .Q(WX3410) );
  INVX0 U6267_U1 ( .INP(n5531), .ZN(U6267_n1) );
  AND2X1 U6268_U2 ( .IN1(WX3345), .IN2(U6268_n1), .Q(WX3408) );
  INVX0 U6268_U1 ( .INP(n5531), .ZN(U6268_n1) );
  AND2X1 U6269_U2 ( .IN1(WX3343), .IN2(U6269_n1), .Q(WX3406) );
  INVX0 U6269_U1 ( .INP(n5531), .ZN(U6269_n1) );
  AND2X1 U6270_U2 ( .IN1(WX3341), .IN2(U6270_n1), .Q(WX3404) );
  INVX0 U6270_U1 ( .INP(n5494), .ZN(U6270_n1) );
  AND2X1 U6271_U2 ( .IN1(WX3339), .IN2(U6271_n1), .Q(WX3402) );
  INVX0 U6271_U1 ( .INP(n5494), .ZN(U6271_n1) );
  AND2X1 U6272_U2 ( .IN1(WX3337), .IN2(U6272_n1), .Q(WX3400) );
  INVX0 U6272_U1 ( .INP(n5494), .ZN(U6272_n1) );
  AND2X1 U6273_U2 ( .IN1(WX3335), .IN2(U6273_n1), .Q(WX3398) );
  INVX0 U6273_U1 ( .INP(n5494), .ZN(U6273_n1) );
  AND2X1 U6274_U2 ( .IN1(test_so26), .IN2(U6274_n1), .Q(WX3396) );
  INVX0 U6274_U1 ( .INP(n5494), .ZN(U6274_n1) );
  AND2X1 U6275_U2 ( .IN1(WX3331), .IN2(U6275_n1), .Q(WX3394) );
  INVX0 U6275_U1 ( .INP(n5494), .ZN(U6275_n1) );
  AND2X1 U6276_U2 ( .IN1(WX3329), .IN2(U6276_n1), .Q(WX3392) );
  INVX0 U6276_U1 ( .INP(n5494), .ZN(U6276_n1) );
  AND2X1 U6277_U2 ( .IN1(WX3327), .IN2(U6277_n1), .Q(WX3390) );
  INVX0 U6277_U1 ( .INP(n5494), .ZN(U6277_n1) );
  AND2X1 U6278_U2 ( .IN1(WX3325), .IN2(U6278_n1), .Q(WX3388) );
  INVX0 U6278_U1 ( .INP(n5494), .ZN(U6278_n1) );
  AND2X1 U6279_U2 ( .IN1(WX3323), .IN2(U6279_n1), .Q(WX3386) );
  INVX0 U6279_U1 ( .INP(n5494), .ZN(U6279_n1) );
  AND2X1 U6280_U2 ( .IN1(WX3321), .IN2(U6280_n1), .Q(WX3384) );
  INVX0 U6280_U1 ( .INP(n5493), .ZN(U6280_n1) );
  AND2X1 U6281_U2 ( .IN1(WX3319), .IN2(U6281_n1), .Q(WX3382) );
  INVX0 U6281_U1 ( .INP(n5493), .ZN(U6281_n1) );
  AND2X1 U6282_U2 ( .IN1(WX3317), .IN2(U6282_n1), .Q(WX3380) );
  INVX0 U6282_U1 ( .INP(n5493), .ZN(U6282_n1) );
  AND2X1 U6283_U2 ( .IN1(WX3315), .IN2(U6283_n1), .Q(WX3378) );
  INVX0 U6283_U1 ( .INP(n5493), .ZN(U6283_n1) );
  AND2X1 U6284_U2 ( .IN1(WX3313), .IN2(U6284_n1), .Q(WX3376) );
  INVX0 U6284_U1 ( .INP(n5493), .ZN(U6284_n1) );
  AND2X1 U6285_U2 ( .IN1(WX3311), .IN2(U6285_n1), .Q(WX3374) );
  INVX0 U6285_U1 ( .INP(n5493), .ZN(U6285_n1) );
  AND2X1 U6286_U2 ( .IN1(WX3309), .IN2(U6286_n1), .Q(WX3372) );
  INVX0 U6286_U1 ( .INP(n5493), .ZN(U6286_n1) );
  AND2X1 U6287_U2 ( .IN1(WX3307), .IN2(U6287_n1), .Q(WX3370) );
  INVX0 U6287_U1 ( .INP(n5493), .ZN(U6287_n1) );
  AND2X1 U6288_U2 ( .IN1(WX3305), .IN2(U6288_n1), .Q(WX3368) );
  INVX0 U6288_U1 ( .INP(n5493), .ZN(U6288_n1) );
  AND2X1 U6289_U2 ( .IN1(WX3303), .IN2(U6289_n1), .Q(WX3366) );
  INVX0 U6289_U1 ( .INP(n5493), .ZN(U6289_n1) );
  AND2X1 U6290_U2 ( .IN1(WX3301), .IN2(U6290_n1), .Q(WX3364) );
  INVX0 U6290_U1 ( .INP(n5493), .ZN(U6290_n1) );
  AND2X1 U6291_U2 ( .IN1(WX3299), .IN2(U6291_n1), .Q(WX3362) );
  INVX0 U6291_U1 ( .INP(n5493), .ZN(U6291_n1) );
  AND2X1 U6292_U2 ( .IN1(test_so25), .IN2(U6292_n1), .Q(WX3360) );
  INVX0 U6292_U1 ( .INP(n5493), .ZN(U6292_n1) );
  AND2X1 U6293_U2 ( .IN1(WX3295), .IN2(U6293_n1), .Q(WX3358) );
  INVX0 U6293_U1 ( .INP(n5493), .ZN(U6293_n1) );
  AND2X1 U6294_U2 ( .IN1(WX3293), .IN2(U6294_n1), .Q(WX3356) );
  INVX0 U6294_U1 ( .INP(n5492), .ZN(U6294_n1) );
  AND2X1 U6295_U2 ( .IN1(WX3291), .IN2(U6295_n1), .Q(WX3354) );
  INVX0 U6295_U1 ( .INP(n5492), .ZN(U6295_n1) );
  AND2X1 U6296_U2 ( .IN1(WX3289), .IN2(U6296_n1), .Q(WX3352) );
  INVX0 U6296_U1 ( .INP(n5492), .ZN(U6296_n1) );
  AND2X1 U6297_U2 ( .IN1(WX3287), .IN2(U6297_n1), .Q(WX3350) );
  INVX0 U6297_U1 ( .INP(n5492), .ZN(U6297_n1) );
  AND2X1 U6298_U2 ( .IN1(WX3285), .IN2(U6298_n1), .Q(WX3348) );
  INVX0 U6298_U1 ( .INP(n5492), .ZN(U6298_n1) );
  AND2X1 U6299_U2 ( .IN1(WX3283), .IN2(U6299_n1), .Q(WX3346) );
  INVX0 U6299_U1 ( .INP(n5492), .ZN(U6299_n1) );
  AND2X1 U6300_U2 ( .IN1(WX3281), .IN2(U6300_n1), .Q(WX3344) );
  INVX0 U6300_U1 ( .INP(n5492), .ZN(U6300_n1) );
  AND2X1 U6301_U2 ( .IN1(WX3279), .IN2(U6301_n1), .Q(WX3342) );
  INVX0 U6301_U1 ( .INP(n5492), .ZN(U6301_n1) );
  AND2X1 U6302_U2 ( .IN1(WX3277), .IN2(U6302_n1), .Q(WX3340) );
  INVX0 U6302_U1 ( .INP(n5492), .ZN(U6302_n1) );
  AND2X1 U6303_U2 ( .IN1(WX3275), .IN2(U6303_n1), .Q(WX3338) );
  INVX0 U6303_U1 ( .INP(n5492), .ZN(U6303_n1) );
  AND2X1 U6304_U2 ( .IN1(WX3273), .IN2(U6304_n1), .Q(WX3336) );
  INVX0 U6304_U1 ( .INP(n5492), .ZN(U6304_n1) );
  AND2X1 U6305_U2 ( .IN1(WX3271), .IN2(U6305_n1), .Q(WX3334) );
  INVX0 U6305_U1 ( .INP(n5492), .ZN(U6305_n1) );
  AND2X1 U6306_U2 ( .IN1(WX3267), .IN2(U6306_n1), .Q(WX3330) );
  INVX0 U6306_U1 ( .INP(n5492), .ZN(U6306_n1) );
  AND2X1 U6307_U2 ( .IN1(WX2128), .IN2(U6307_n1), .Q(WX2191) );
  INVX0 U6307_U1 ( .INP(n5492), .ZN(U6307_n1) );
  AND2X1 U6308_U2 ( .IN1(WX2126), .IN2(U6308_n1), .Q(WX2189) );
  INVX0 U6308_U1 ( .INP(n5491), .ZN(U6308_n1) );
  AND2X1 U6309_U2 ( .IN1(WX2124), .IN2(U6309_n1), .Q(WX2187) );
  INVX0 U6309_U1 ( .INP(n5491), .ZN(U6309_n1) );
  AND2X1 U6310_U2 ( .IN1(WX2122), .IN2(U6310_n1), .Q(WX2185) );
  INVX0 U6310_U1 ( .INP(n5491), .ZN(U6310_n1) );
  AND2X1 U6311_U2 ( .IN1(WX2120), .IN2(U6311_n1), .Q(WX2183) );
  INVX0 U6311_U1 ( .INP(n5491), .ZN(U6311_n1) );
  AND2X1 U6312_U2 ( .IN1(WX2118), .IN2(U6312_n1), .Q(WX2181) );
  INVX0 U6312_U1 ( .INP(n5491), .ZN(U6312_n1) );
  AND2X1 U6313_U2 ( .IN1(WX2116), .IN2(U6313_n1), .Q(WX2179) );
  INVX0 U6313_U1 ( .INP(n5491), .ZN(U6313_n1) );
  AND2X1 U6314_U2 ( .IN1(WX2114), .IN2(U6314_n1), .Q(WX2177) );
  INVX0 U6314_U1 ( .INP(n5491), .ZN(U6314_n1) );
  AND2X1 U6315_U2 ( .IN1(WX2112), .IN2(U6315_n1), .Q(WX2175) );
  INVX0 U6315_U1 ( .INP(n5491), .ZN(U6315_n1) );
  AND2X1 U6316_U2 ( .IN1(WX2110), .IN2(U6316_n1), .Q(WX2173) );
  INVX0 U6316_U1 ( .INP(n5491), .ZN(U6316_n1) );
  AND2X1 U6317_U2 ( .IN1(WX2108), .IN2(U6317_n1), .Q(WX2171) );
  INVX0 U6317_U1 ( .INP(n5491), .ZN(U6317_n1) );
  AND2X1 U6318_U2 ( .IN1(WX2106), .IN2(U6318_n1), .Q(WX2169) );
  INVX0 U6318_U1 ( .INP(n5491), .ZN(U6318_n1) );
  AND2X1 U6319_U2 ( .IN1(WX2104), .IN2(U6319_n1), .Q(WX2167) );
  INVX0 U6319_U1 ( .INP(n5491), .ZN(U6319_n1) );
  AND2X1 U6320_U2 ( .IN1(WX2102), .IN2(U6320_n1), .Q(WX2165) );
  INVX0 U6320_U1 ( .INP(n5491), .ZN(U6320_n1) );
  AND2X1 U6321_U2 ( .IN1(test_so17), .IN2(U6321_n1), .Q(WX2163) );
  INVX0 U6321_U1 ( .INP(n5491), .ZN(U6321_n1) );
  AND2X1 U6322_U2 ( .IN1(WX2098), .IN2(U6322_n1), .Q(WX2161) );
  INVX0 U6322_U1 ( .INP(n5490), .ZN(U6322_n1) );
  AND2X1 U6323_U2 ( .IN1(WX2096), .IN2(U6323_n1), .Q(WX2159) );
  INVX0 U6323_U1 ( .INP(n5490), .ZN(U6323_n1) );
  AND2X1 U6324_U2 ( .IN1(WX2094), .IN2(U6324_n1), .Q(WX2157) );
  INVX0 U6324_U1 ( .INP(n5490), .ZN(U6324_n1) );
  AND2X1 U6325_U2 ( .IN1(WX2092), .IN2(U6325_n1), .Q(WX2155) );
  INVX0 U6325_U1 ( .INP(n5490), .ZN(U6325_n1) );
  AND2X1 U6326_U2 ( .IN1(WX2090), .IN2(U6326_n1), .Q(WX2153) );
  INVX0 U6326_U1 ( .INP(n5490), .ZN(U6326_n1) );
  AND2X1 U6327_U2 ( .IN1(WX2088), .IN2(U6327_n1), .Q(WX2151) );
  INVX0 U6327_U1 ( .INP(n5490), .ZN(U6327_n1) );
  AND2X1 U6328_U2 ( .IN1(WX2086), .IN2(U6328_n1), .Q(WX2149) );
  INVX0 U6328_U1 ( .INP(n5490), .ZN(U6328_n1) );
  AND2X1 U6329_U2 ( .IN1(WX2084), .IN2(U6329_n1), .Q(WX2147) );
  INVX0 U6329_U1 ( .INP(n5490), .ZN(U6329_n1) );
  AND2X1 U6330_U2 ( .IN1(WX2082), .IN2(U6330_n1), .Q(WX2145) );
  INVX0 U6330_U1 ( .INP(n5490), .ZN(U6330_n1) );
  AND2X1 U6331_U2 ( .IN1(WX2080), .IN2(U6331_n1), .Q(WX2143) );
  INVX0 U6331_U1 ( .INP(n5490), .ZN(U6331_n1) );
  AND2X1 U6332_U2 ( .IN1(WX2078), .IN2(U6332_n1), .Q(WX2141) );
  INVX0 U6332_U1 ( .INP(n5490), .ZN(U6332_n1) );
  AND2X1 U6333_U2 ( .IN1(WX2076), .IN2(U6333_n1), .Q(WX2139) );
  INVX0 U6333_U1 ( .INP(n5490), .ZN(U6333_n1) );
  AND2X1 U6334_U2 ( .IN1(WX2074), .IN2(U6334_n1), .Q(WX2137) );
  INVX0 U6334_U1 ( .INP(n5490), .ZN(U6334_n1) );
  AND2X1 U6335_U2 ( .IN1(WX2072), .IN2(U6335_n1), .Q(WX2135) );
  INVX0 U6335_U1 ( .INP(n5489), .ZN(U6335_n1) );
  AND2X1 U6336_U2 ( .IN1(WX2070), .IN2(U6336_n1), .Q(WX2133) );
  INVX0 U6336_U1 ( .INP(n5489), .ZN(U6336_n1) );
  AND2X1 U6337_U2 ( .IN1(WX2068), .IN2(U6337_n1), .Q(WX2131) );
  INVX0 U6337_U1 ( .INP(n5489), .ZN(U6337_n1) );
  AND2X1 U6338_U2 ( .IN1(WX2066), .IN2(U6338_n1), .Q(WX2129) );
  INVX0 U6338_U1 ( .INP(n5489), .ZN(U6338_n1) );
  AND2X1 U6339_U2 ( .IN1(test_so16), .IN2(U6339_n1), .Q(WX2127) );
  INVX0 U6339_U1 ( .INP(n5489), .ZN(U6339_n1) );
  AND2X1 U6340_U2 ( .IN1(WX2062), .IN2(U6340_n1), .Q(WX2125) );
  INVX0 U6340_U1 ( .INP(n5489), .ZN(U6340_n1) );
  AND2X1 U6341_U2 ( .IN1(WX2060), .IN2(U6341_n1), .Q(WX2123) );
  INVX0 U6341_U1 ( .INP(n5489), .ZN(U6341_n1) );
  AND2X1 U6342_U2 ( .IN1(WX2058), .IN2(U6342_n1), .Q(WX2121) );
  INVX0 U6342_U1 ( .INP(n5489), .ZN(U6342_n1) );
  AND2X1 U6343_U2 ( .IN1(WX2056), .IN2(U6343_n1), .Q(WX2119) );
  INVX0 U6343_U1 ( .INP(n5489), .ZN(U6343_n1) );
  AND2X1 U6344_U2 ( .IN1(WX2054), .IN2(U6344_n1), .Q(WX2117) );
  INVX0 U6344_U1 ( .INP(n5489), .ZN(U6344_n1) );
  AND2X1 U6345_U2 ( .IN1(WX2052), .IN2(U6345_n1), .Q(WX2115) );
  INVX0 U6345_U1 ( .INP(n5489), .ZN(U6345_n1) );
  AND2X1 U6346_U2 ( .IN1(WX2050), .IN2(U6346_n1), .Q(WX2113) );
  INVX0 U6346_U1 ( .INP(n5489), .ZN(U6346_n1) );
  AND2X1 U6347_U2 ( .IN1(WX2048), .IN2(U6347_n1), .Q(WX2111) );
  INVX0 U6347_U1 ( .INP(n5489), .ZN(U6347_n1) );
  AND2X1 U6348_U2 ( .IN1(WX2046), .IN2(U6348_n1), .Q(WX2109) );
  INVX0 U6348_U1 ( .INP(n5489), .ZN(U6348_n1) );
  AND2X1 U6349_U2 ( .IN1(WX2044), .IN2(U6349_n1), .Q(WX2107) );
  INVX0 U6349_U1 ( .INP(n5488), .ZN(U6349_n1) );
  AND2X1 U6350_U2 ( .IN1(WX2042), .IN2(U6350_n1), .Q(WX2105) );
  INVX0 U6350_U1 ( .INP(n5488), .ZN(U6350_n1) );
  AND2X1 U6351_U2 ( .IN1(WX2040), .IN2(U6351_n1), .Q(WX2103) );
  INVX0 U6351_U1 ( .INP(n5488), .ZN(U6351_n1) );
  AND2X1 U6352_U2 ( .IN1(WX2038), .IN2(U6352_n1), .Q(WX2101) );
  INVX0 U6352_U1 ( .INP(n5488), .ZN(U6352_n1) );
  AND2X1 U6353_U2 ( .IN1(WX2036), .IN2(U6353_n1), .Q(WX2099) );
  INVX0 U6353_U1 ( .INP(n5488), .ZN(U6353_n1) );
  AND2X1 U6354_U2 ( .IN1(WX2034), .IN2(U6354_n1), .Q(WX2097) );
  INVX0 U6354_U1 ( .INP(n5488), .ZN(U6354_n1) );
  AND2X1 U6355_U2 ( .IN1(WX2032), .IN2(U6355_n1), .Q(WX2095) );
  INVX0 U6355_U1 ( .INP(n5488), .ZN(U6355_n1) );
  AND2X1 U6356_U2 ( .IN1(WX2030), .IN2(U6356_n1), .Q(WX2093) );
  INVX0 U6356_U1 ( .INP(n5488), .ZN(U6356_n1) );
  AND2X1 U6357_U2 ( .IN1(test_so15), .IN2(U6357_n1), .Q(WX2091) );
  INVX0 U6357_U1 ( .INP(n5488), .ZN(U6357_n1) );
  AND2X1 U6358_U2 ( .IN1(WX2026), .IN2(U6358_n1), .Q(WX2089) );
  INVX0 U6358_U1 ( .INP(n5488), .ZN(U6358_n1) );
  AND2X1 U6359_U2 ( .IN1(WX2024), .IN2(U6359_n1), .Q(WX2087) );
  INVX0 U6359_U1 ( .INP(n5488), .ZN(U6359_n1) );
  AND2X1 U6360_U2 ( .IN1(WX2022), .IN2(U6360_n1), .Q(WX2085) );
  INVX0 U6360_U1 ( .INP(n5488), .ZN(U6360_n1) );
  AND2X1 U6361_U2 ( .IN1(WX2020), .IN2(U6361_n1), .Q(WX2083) );
  INVX0 U6361_U1 ( .INP(n5488), .ZN(U6361_n1) );
  AND2X1 U6362_U2 ( .IN1(WX2018), .IN2(U6362_n1), .Q(WX2081) );
  INVX0 U6362_U1 ( .INP(n5488), .ZN(U6362_n1) );
  AND2X1 U6363_U2 ( .IN1(WX2016), .IN2(U6363_n1), .Q(WX2079) );
  INVX0 U6363_U1 ( .INP(n5487), .ZN(U6363_n1) );
  AND2X1 U6364_U2 ( .IN1(WX2014), .IN2(U6364_n1), .Q(WX2077) );
  INVX0 U6364_U1 ( .INP(n5487), .ZN(U6364_n1) );
  AND2X1 U6365_U2 ( .IN1(WX2012), .IN2(U6365_n1), .Q(WX2075) );
  INVX0 U6365_U1 ( .INP(n5487), .ZN(U6365_n1) );
  AND2X1 U6366_U2 ( .IN1(WX2010), .IN2(U6366_n1), .Q(WX2073) );
  INVX0 U6366_U1 ( .INP(n5487), .ZN(U6366_n1) );
  AND2X1 U6367_U2 ( .IN1(WX2008), .IN2(U6367_n1), .Q(WX2071) );
  INVX0 U6367_U1 ( .INP(n5487), .ZN(U6367_n1) );
  AND2X1 U6368_U2 ( .IN1(WX2006), .IN2(U6368_n1), .Q(WX2069) );
  INVX0 U6368_U1 ( .INP(n5487), .ZN(U6368_n1) );
  AND2X1 U6369_U2 ( .IN1(WX2004), .IN2(U6369_n1), .Q(WX2067) );
  INVX0 U6369_U1 ( .INP(n5487), .ZN(U6369_n1) );
  AND2X1 U6370_U2 ( .IN1(WX2002), .IN2(U6370_n1), .Q(WX2065) );
  INVX0 U6370_U1 ( .INP(n5487), .ZN(U6370_n1) );
  AND2X1 U6371_U2 ( .IN1(WX2000), .IN2(U6371_n1), .Q(WX2063) );
  INVX0 U6371_U1 ( .INP(n5487), .ZN(U6371_n1) );
  AND2X1 U6372_U2 ( .IN1(WX1998), .IN2(U6372_n1), .Q(WX2061) );
  INVX0 U6372_U1 ( .INP(n5487), .ZN(U6372_n1) );
  AND2X1 U6373_U2 ( .IN1(WX1996), .IN2(U6373_n1), .Q(WX2059) );
  INVX0 U6373_U1 ( .INP(n5487), .ZN(U6373_n1) );
  AND2X1 U6374_U2 ( .IN1(WX1994), .IN2(U6374_n1), .Q(WX2057) );
  INVX0 U6374_U1 ( .INP(n5487), .ZN(U6374_n1) );
  AND2X1 U6375_U2 ( .IN1(test_so14), .IN2(U6375_n1), .Q(WX2055) );
  INVX0 U6375_U1 ( .INP(n5487), .ZN(U6375_n1) );
  AND2X1 U6376_U2 ( .IN1(WX1990), .IN2(U6376_n1), .Q(WX2053) );
  INVX0 U6376_U1 ( .INP(n5490), .ZN(U6376_n1) );
  AND2X1 U6377_U2 ( .IN1(WX1988), .IN2(U6377_n1), .Q(WX2051) );
  INVX0 U6377_U1 ( .INP(n5502), .ZN(U6377_n1) );
  AND2X1 U6378_U2 ( .IN1(WX1986), .IN2(U6378_n1), .Q(WX2049) );
  INVX0 U6378_U1 ( .INP(n5502), .ZN(U6378_n1) );
  AND2X1 U6379_U2 ( .IN1(WX1984), .IN2(U6379_n1), .Q(WX2047) );
  INVX0 U6379_U1 ( .INP(n5502), .ZN(U6379_n1) );
  AND2X1 U6380_U2 ( .IN1(WX1982), .IN2(U6380_n1), .Q(WX2045) );
  INVX0 U6380_U1 ( .INP(n5502), .ZN(U6380_n1) );
  AND2X1 U6381_U2 ( .IN1(WX1980), .IN2(U6381_n1), .Q(WX2043) );
  INVX0 U6381_U1 ( .INP(n5502), .ZN(U6381_n1) );
  AND2X1 U6382_U2 ( .IN1(WX1978), .IN2(U6382_n1), .Q(WX2041) );
  INVX0 U6382_U1 ( .INP(n5501), .ZN(U6382_n1) );
  AND2X1 U6383_U2 ( .IN1(WX1976), .IN2(U6383_n1), .Q(WX2039) );
  INVX0 U6383_U1 ( .INP(n5501), .ZN(U6383_n1) );
  AND2X1 U6384_U2 ( .IN1(WX1974), .IN2(U6384_n1), .Q(WX2037) );
  INVX0 U6384_U1 ( .INP(n5501), .ZN(U6384_n1) );
  AND2X1 U6385_U2 ( .IN1(WX1972), .IN2(U6385_n1), .Q(WX2035) );
  INVX0 U6385_U1 ( .INP(n5501), .ZN(U6385_n1) );
  AND2X1 U6386_U2 ( .IN1(WX1970), .IN2(U6386_n1), .Q(WX2033) );
  INVX0 U6386_U1 ( .INP(n5501), .ZN(U6386_n1) );
  AND2X1 U6387_U2 ( .IN1(WX835), .IN2(U6387_n1), .Q(WX898) );
  INVX0 U6387_U1 ( .INP(n5501), .ZN(U6387_n1) );
  AND2X1 U6388_U2 ( .IN1(WX833), .IN2(U6388_n1), .Q(WX896) );
  INVX0 U6388_U1 ( .INP(n5501), .ZN(U6388_n1) );
  AND2X1 U6389_U2 ( .IN1(test_so7), .IN2(U6389_n1), .Q(WX894) );
  INVX0 U6389_U1 ( .INP(n5501), .ZN(U6389_n1) );
  AND2X1 U6390_U2 ( .IN1(WX829), .IN2(U6390_n1), .Q(WX892) );
  INVX0 U6390_U1 ( .INP(n5501), .ZN(U6390_n1) );
  AND2X1 U6391_U2 ( .IN1(WX827), .IN2(U6391_n1), .Q(WX890) );
  INVX0 U6391_U1 ( .INP(n5501), .ZN(U6391_n1) );
  AND2X1 U6392_U2 ( .IN1(WX825), .IN2(U6392_n1), .Q(WX888) );
  INVX0 U6392_U1 ( .INP(n5501), .ZN(U6392_n1) );
  AND2X1 U6393_U2 ( .IN1(WX823), .IN2(U6393_n1), .Q(WX886) );
  INVX0 U6393_U1 ( .INP(n5501), .ZN(U6393_n1) );
  AND2X1 U6394_U2 ( .IN1(WX821), .IN2(U6394_n1), .Q(WX884) );
  INVX0 U6394_U1 ( .INP(n5501), .ZN(U6394_n1) );
  AND2X1 U6395_U2 ( .IN1(WX819), .IN2(U6395_n1), .Q(WX882) );
  INVX0 U6395_U1 ( .INP(n5501), .ZN(U6395_n1) );
  AND2X1 U6396_U2 ( .IN1(WX817), .IN2(U6396_n1), .Q(WX880) );
  INVX0 U6396_U1 ( .INP(n5500), .ZN(U6396_n1) );
  AND2X1 U6397_U2 ( .IN1(WX815), .IN2(U6397_n1), .Q(WX878) );
  INVX0 U6397_U1 ( .INP(n5500), .ZN(U6397_n1) );
  AND2X1 U6398_U2 ( .IN1(WX813), .IN2(U6398_n1), .Q(WX876) );
  INVX0 U6398_U1 ( .INP(n5500), .ZN(U6398_n1) );
  AND2X1 U6399_U2 ( .IN1(WX811), .IN2(U6399_n1), .Q(WX874) );
  INVX0 U6399_U1 ( .INP(n5500), .ZN(U6399_n1) );
  AND2X1 U6400_U2 ( .IN1(WX809), .IN2(U6400_n1), .Q(WX872) );
  INVX0 U6400_U1 ( .INP(n5500), .ZN(U6400_n1) );
  AND2X1 U6401_U2 ( .IN1(WX807), .IN2(U6401_n1), .Q(WX870) );
  INVX0 U6401_U1 ( .INP(n5500), .ZN(U6401_n1) );
  AND2X1 U6402_U2 ( .IN1(WX805), .IN2(U6402_n1), .Q(WX868) );
  INVX0 U6402_U1 ( .INP(n5500), .ZN(U6402_n1) );
  AND2X1 U6403_U2 ( .IN1(WX803), .IN2(U6403_n1), .Q(WX866) );
  INVX0 U6403_U1 ( .INP(n5500), .ZN(U6403_n1) );
  AND2X1 U6404_U2 ( .IN1(WX801), .IN2(U6404_n1), .Q(WX864) );
  INVX0 U6404_U1 ( .INP(n5500), .ZN(U6404_n1) );
  AND2X1 U6405_U2 ( .IN1(WX799), .IN2(U6405_n1), .Q(WX862) );
  INVX0 U6405_U1 ( .INP(n5500), .ZN(U6405_n1) );
  AND2X1 U6406_U2 ( .IN1(WX797), .IN2(U6406_n1), .Q(WX860) );
  INVX0 U6406_U1 ( .INP(n5500), .ZN(U6406_n1) );
  AND2X1 U6407_U2 ( .IN1(test_so6), .IN2(U6407_n1), .Q(WX858) );
  INVX0 U6407_U1 ( .INP(n5500), .ZN(U6407_n1) );
  AND2X1 U6408_U2 ( .IN1(WX793), .IN2(U6408_n1), .Q(WX856) );
  INVX0 U6408_U1 ( .INP(n5500), .ZN(U6408_n1) );
  AND2X1 U6409_U2 ( .IN1(WX791), .IN2(U6409_n1), .Q(WX854) );
  INVX0 U6409_U1 ( .INP(n5500), .ZN(U6409_n1) );
  AND2X1 U6410_U2 ( .IN1(WX789), .IN2(U6410_n1), .Q(WX852) );
  INVX0 U6410_U1 ( .INP(n5499), .ZN(U6410_n1) );
  AND2X1 U6411_U2 ( .IN1(WX787), .IN2(U6411_n1), .Q(WX850) );
  INVX0 U6411_U1 ( .INP(n5499), .ZN(U6411_n1) );
  AND2X1 U6412_U2 ( .IN1(WX785), .IN2(U6412_n1), .Q(WX848) );
  INVX0 U6412_U1 ( .INP(n5499), .ZN(U6412_n1) );
  AND2X1 U6413_U2 ( .IN1(WX783), .IN2(U6413_n1), .Q(WX846) );
  INVX0 U6413_U1 ( .INP(n5499), .ZN(U6413_n1) );
  AND2X1 U6414_U2 ( .IN1(WX781), .IN2(U6414_n1), .Q(WX844) );
  INVX0 U6414_U1 ( .INP(n5499), .ZN(U6414_n1) );
  AND2X1 U6415_U2 ( .IN1(WX779), .IN2(U6415_n1), .Q(WX842) );
  INVX0 U6415_U1 ( .INP(n5499), .ZN(U6415_n1) );
  AND2X1 U6416_U2 ( .IN1(WX777), .IN2(U6416_n1), .Q(WX840) );
  INVX0 U6416_U1 ( .INP(n5499), .ZN(U6416_n1) );
  AND2X1 U6417_U2 ( .IN1(WX775), .IN2(U6417_n1), .Q(WX838) );
  INVX0 U6417_U1 ( .INP(n5499), .ZN(U6417_n1) );
  AND2X1 U6418_U2 ( .IN1(WX773), .IN2(U6418_n1), .Q(WX836) );
  INVX0 U6418_U1 ( .INP(n5499), .ZN(U6418_n1) );
  AND2X1 U6419_U2 ( .IN1(WX771), .IN2(U6419_n1), .Q(WX834) );
  INVX0 U6419_U1 ( .INP(n5499), .ZN(U6419_n1) );
  AND2X1 U6420_U2 ( .IN1(WX769), .IN2(U6420_n1), .Q(WX832) );
  INVX0 U6420_U1 ( .INP(n5499), .ZN(U6420_n1) );
  AND2X1 U6421_U2 ( .IN1(WX767), .IN2(U6421_n1), .Q(WX830) );
  INVX0 U6421_U1 ( .INP(n5499), .ZN(U6421_n1) );
  AND2X1 U6422_U2 ( .IN1(WX765), .IN2(U6422_n1), .Q(WX828) );
  INVX0 U6422_U1 ( .INP(n5499), .ZN(U6422_n1) );
  AND2X1 U6423_U2 ( .IN1(WX763), .IN2(U6423_n1), .Q(WX826) );
  INVX0 U6423_U1 ( .INP(n5499), .ZN(U6423_n1) );
  AND2X1 U6424_U2 ( .IN1(WX761), .IN2(U6424_n1), .Q(WX824) );
  INVX0 U6424_U1 ( .INP(n5498), .ZN(U6424_n1) );
  AND2X1 U6425_U2 ( .IN1(test_so5), .IN2(U6425_n1), .Q(WX822) );
  INVX0 U6425_U1 ( .INP(n5498), .ZN(U6425_n1) );
  AND2X1 U6426_U2 ( .IN1(WX757), .IN2(U6426_n1), .Q(WX820) );
  INVX0 U6426_U1 ( .INP(n5498), .ZN(U6426_n1) );
  AND2X1 U6427_U2 ( .IN1(WX755), .IN2(U6427_n1), .Q(WX818) );
  INVX0 U6427_U1 ( .INP(n5498), .ZN(U6427_n1) );
  AND2X1 U6428_U2 ( .IN1(WX753), .IN2(U6428_n1), .Q(WX816) );
  INVX0 U6428_U1 ( .INP(n5498), .ZN(U6428_n1) );
  AND2X1 U6429_U2 ( .IN1(WX751), .IN2(U6429_n1), .Q(WX814) );
  INVX0 U6429_U1 ( .INP(n5498), .ZN(U6429_n1) );
  AND2X1 U6430_U2 ( .IN1(WX749), .IN2(U6430_n1), .Q(WX812) );
  INVX0 U6430_U1 ( .INP(n5498), .ZN(U6430_n1) );
  AND2X1 U6431_U2 ( .IN1(WX747), .IN2(U6431_n1), .Q(WX810) );
  INVX0 U6431_U1 ( .INP(n5498), .ZN(U6431_n1) );
  AND2X1 U6432_U2 ( .IN1(WX745), .IN2(U6432_n1), .Q(WX808) );
  INVX0 U6432_U1 ( .INP(n5498), .ZN(U6432_n1) );
  AND2X1 U6433_U2 ( .IN1(WX743), .IN2(U6433_n1), .Q(WX806) );
  INVX0 U6433_U1 ( .INP(n5498), .ZN(U6433_n1) );
  AND2X1 U6434_U2 ( .IN1(WX741), .IN2(U6434_n1), .Q(WX804) );
  INVX0 U6434_U1 ( .INP(n5498), .ZN(U6434_n1) );
  AND2X1 U6435_U2 ( .IN1(WX739), .IN2(U6435_n1), .Q(WX802) );
  INVX0 U6435_U1 ( .INP(n5498), .ZN(U6435_n1) );
  AND2X1 U6436_U2 ( .IN1(WX737), .IN2(U6436_n1), .Q(WX800) );
  INVX0 U6436_U1 ( .INP(n5498), .ZN(U6436_n1) );
  AND2X1 U6437_U2 ( .IN1(WX735), .IN2(U6437_n1), .Q(WX798) );
  INVX0 U6437_U1 ( .INP(n5497), .ZN(U6437_n1) );
  AND2X1 U6438_U2 ( .IN1(WX733), .IN2(U6438_n1), .Q(WX796) );
  INVX0 U6438_U1 ( .INP(n5497), .ZN(U6438_n1) );
  AND2X1 U6439_U2 ( .IN1(WX731), .IN2(U6439_n1), .Q(WX794) );
  INVX0 U6439_U1 ( .INP(n5497), .ZN(U6439_n1) );
  AND2X1 U6440_U2 ( .IN1(WX729), .IN2(U6440_n1), .Q(WX792) );
  INVX0 U6440_U1 ( .INP(n5497), .ZN(U6440_n1) );
  AND2X1 U6441_U2 ( .IN1(WX727), .IN2(U6441_n1), .Q(WX790) );
  INVX0 U6441_U1 ( .INP(n5497), .ZN(U6441_n1) );
  AND2X1 U6442_U2 ( .IN1(WX725), .IN2(U6442_n1), .Q(WX788) );
  INVX0 U6442_U1 ( .INP(n5497), .ZN(U6442_n1) );
  AND2X1 U6443_U2 ( .IN1(test_so4), .IN2(U6443_n1), .Q(WX786) );
  INVX0 U6443_U1 ( .INP(n5497), .ZN(U6443_n1) );
  AND2X1 U6444_U2 ( .IN1(WX721), .IN2(U6444_n1), .Q(WX784) );
  INVX0 U6444_U1 ( .INP(n5497), .ZN(U6444_n1) );
  AND2X1 U6445_U2 ( .IN1(WX719), .IN2(U6445_n1), .Q(WX782) );
  INVX0 U6445_U1 ( .INP(n5497), .ZN(U6445_n1) );
  AND2X1 U6446_U2 ( .IN1(WX717), .IN2(U6446_n1), .Q(WX780) );
  INVX0 U6446_U1 ( .INP(n5497), .ZN(U6446_n1) );
  AND2X1 U6447_U2 ( .IN1(WX715), .IN2(U6447_n1), .Q(WX778) );
  INVX0 U6447_U1 ( .INP(n5497), .ZN(U6447_n1) );
  AND2X1 U6448_U2 ( .IN1(WX713), .IN2(U6448_n1), .Q(WX776) );
  INVX0 U6448_U1 ( .INP(n5497), .ZN(U6448_n1) );
  AND2X1 U6449_U2 ( .IN1(WX711), .IN2(U6449_n1), .Q(WX774) );
  INVX0 U6449_U1 ( .INP(n5497), .ZN(U6449_n1) );
  AND2X1 U6450_U2 ( .IN1(WX709), .IN2(U6450_n1), .Q(WX772) );
  INVX0 U6450_U1 ( .INP(n5497), .ZN(U6450_n1) );
  AND2X1 U6451_U2 ( .IN1(WX707), .IN2(U6451_n1), .Q(WX770) );
  INVX0 U6451_U1 ( .INP(n5496), .ZN(U6451_n1) );
  AND2X1 U6452_U2 ( .IN1(WX705), .IN2(U6452_n1), .Q(WX768) );
  INVX0 U6452_U1 ( .INP(n5496), .ZN(U6452_n1) );
  AND2X1 U6453_U2 ( .IN1(WX703), .IN2(U6453_n1), .Q(WX766) );
  INVX0 U6453_U1 ( .INP(n5496), .ZN(U6453_n1) );
  AND2X1 U6454_U2 ( .IN1(WX701), .IN2(U6454_n1), .Q(WX764) );
  INVX0 U6454_U1 ( .INP(n5496), .ZN(U6454_n1) );
  AND2X1 U6455_U2 ( .IN1(WX699), .IN2(U6455_n1), .Q(WX762) );
  INVX0 U6455_U1 ( .INP(n5496), .ZN(U6455_n1) );
  AND2X1 U6456_U2 ( .IN1(WX697), .IN2(U6456_n1), .Q(WX760) );
  INVX0 U6456_U1 ( .INP(n5496), .ZN(U6456_n1) );
  AND2X1 U6457_U2 ( .IN1(WX695), .IN2(U6457_n1), .Q(WX758) );
  INVX0 U6457_U1 ( .INP(n5496), .ZN(U6457_n1) );
  AND2X1 U6458_U2 ( .IN1(WX693), .IN2(U6458_n1), .Q(WX756) );
  INVX0 U6458_U1 ( .INP(n5496), .ZN(U6458_n1) );
  AND2X1 U6459_U2 ( .IN1(WX691), .IN2(U6459_n1), .Q(WX754) );
  INVX0 U6459_U1 ( .INP(n5496), .ZN(U6459_n1) );
  AND2X1 U6460_U2 ( .IN1(WX689), .IN2(U6460_n1), .Q(WX752) );
  INVX0 U6460_U1 ( .INP(n5496), .ZN(U6460_n1) );
  AND2X1 U6461_U2 ( .IN1(test_so3), .IN2(U6461_n1), .Q(WX750) );
  INVX0 U6461_U1 ( .INP(n5496), .ZN(U6461_n1) );
  AND2X1 U6462_U2 ( .IN1(WX685), .IN2(U6462_n1), .Q(WX748) );
  INVX0 U6462_U1 ( .INP(n5496), .ZN(U6462_n1) );
  AND2X1 U6463_U2 ( .IN1(WX683), .IN2(U6463_n1), .Q(WX746) );
  INVX0 U6463_U1 ( .INP(n5496), .ZN(U6463_n1) );
  AND2X1 U6464_U2 ( .IN1(WX681), .IN2(U6464_n1), .Q(WX744) );
  INVX0 U6464_U1 ( .INP(n5496), .ZN(U6464_n1) );
  AND2X1 U6465_U2 ( .IN1(WX679), .IN2(U6465_n1), .Q(WX742) );
  INVX0 U6465_U1 ( .INP(n5495), .ZN(U6465_n1) );
  AND2X1 U6466_U2 ( .IN1(WX677), .IN2(U6466_n1), .Q(WX740) );
  INVX0 U6466_U1 ( .INP(n5495), .ZN(U6466_n1) );
  AND2X1 U6467_U2 ( .IN1(WX675), .IN2(U6467_n1), .Q(WX738) );
  INVX0 U6467_U1 ( .INP(n5495), .ZN(U6467_n1) );
  AND2X1 U6468_U2 ( .IN1(WX673), .IN2(U6468_n1), .Q(WX736) );
  INVX0 U6468_U1 ( .INP(n5495), .ZN(U6468_n1) );
  AND2X1 U6469_U2 ( .IN1(WX671), .IN2(U6469_n1), .Q(WX734) );
  INVX0 U6469_U1 ( .INP(n5495), .ZN(U6469_n1) );
  AND2X1 U6470_U2 ( .IN1(WX669), .IN2(U6470_n1), .Q(WX732) );
  INVX0 U6470_U1 ( .INP(n5495), .ZN(U6470_n1) );
  AND2X1 U6471_U2 ( .IN1(WX667), .IN2(U6471_n1), .Q(WX730) );
  INVX0 U6471_U1 ( .INP(n5495), .ZN(U6471_n1) );
  AND2X1 U6472_U2 ( .IN1(WX665), .IN2(U6472_n1), .Q(WX728) );
  INVX0 U6472_U1 ( .INP(n5495), .ZN(U6472_n1) );
  AND2X1 U6473_U2 ( .IN1(WX663), .IN2(U6473_n1), .Q(WX726) );
  INVX0 U6473_U1 ( .INP(n5495), .ZN(U6473_n1) );
  AND2X1 U6474_U2 ( .IN1(WX661), .IN2(U6474_n1), .Q(WX724) );
  INVX0 U6474_U1 ( .INP(n5495), .ZN(U6474_n1) );
  AND2X1 U6475_U2 ( .IN1(WX659), .IN2(U6475_n1), .Q(WX722) );
  INVX0 U6475_U1 ( .INP(n5495), .ZN(U6475_n1) );
  AND2X1 U6476_U2 ( .IN1(WX657), .IN2(U6476_n1), .Q(WX720) );
  INVX0 U6476_U1 ( .INP(n5495), .ZN(U6476_n1) );
  AND2X1 U6477_U2 ( .IN1(WX655), .IN2(U6477_n1), .Q(WX718) );
  INVX0 U6477_U1 ( .INP(n5495), .ZN(U6477_n1) );
  AND2X1 U6478_U2 ( .IN1(WX653), .IN2(U6478_n1), .Q(WX716) );
  INVX0 U6478_U1 ( .INP(n5495), .ZN(U6478_n1) );
  AND2X1 U6479_U2 ( .IN1(test_so2), .IN2(U6479_n1), .Q(WX714) );
  INVX0 U6479_U1 ( .INP(n5494), .ZN(U6479_n1) );
  AND2X1 U6480_U2 ( .IN1(WX649), .IN2(U6480_n1), .Q(WX712) );
  INVX0 U6480_U1 ( .INP(n5494), .ZN(U6480_n1) );
  AND2X1 U6481_U2 ( .IN1(WX647), .IN2(U6481_n1), .Q(WX710) );
  INVX0 U6481_U1 ( .INP(n5494), .ZN(U6481_n1) );
  AND2X1 U6482_U2 ( .IN1(WX645), .IN2(U6482_n1), .Q(WX708) );
  INVX0 U6482_U1 ( .INP(n5494), .ZN(U6482_n1) );
endmodule

