module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, 
        CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, 
        CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, 
        CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, 
        CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, 
        CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, 
        CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, 
        CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, 
        CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, 
        CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, 
        CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, 
        CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, 
        CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, 
        CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, 
        CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, 
        CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, 
        CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, 
        CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, 
        CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, 
        CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, 
        CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, 
        CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, 
        CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, 
        CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, 
        CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, 
        CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, 
        CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, 
        CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, 
        CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, 
        CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, 
        CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, 
        CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, 
        CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, 
        CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, 
        CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, 
        CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, 
        CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, 
        CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, 
        CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, 
        CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, 
        CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, 
        CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, 
        CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, 
        CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, 
        CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, 
        CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, 
        CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, 
        CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, 
        CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, 
        CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, 
        CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, 
        CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, 
        CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, 
        CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, 
        CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, 
        CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, 
        CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, 
        CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_0_0, DATA_0_1, 
        DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, DATA_0_14, DATA_0_15, 
        DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, DATA_0_2, DATA_0_20, 
        DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, DATA_0_25, DATA_0_26, 
        DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, DATA_0_30, DATA_0_31, 
        DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, DATA_0_9, DATA_9_0, 
        DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, 
        DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, 
        DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, 
        DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, 
        DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, 
        RESET, TM0, TM1, test_se, test_si1, test_so1, test_si2, test_so2, 
        test_si3, test_so3, test_si4, test_so4, test_si5, test_so5, test_si6, 
        test_so6, test_si7, test_so7, test_si8, test_so8, test_si9, test_so9, 
        test_si10, test_so10, test_si11, test_so11, test_si12, test_so12, 
        test_si13, test_so13, test_si14, test_so14, test_si15, test_so15, 
        test_si16, test_so16, test_si17, test_so17, test_si18, test_so18, 
        test_si19, test_so19, test_si20, test_so20, test_si21, test_so21, 
        test_si22, test_so22, test_si23, test_so23, test_si24, test_so24, 
        test_si25, test_so25, test_si26, test_so26, test_si27, test_so27, 
        test_si28, test_so28, test_si29, test_so29, test_si30, test_so30, 
        test_si31, test_so31, test_si32, test_so32, test_si33, test_so33, 
        test_si34, test_so34, test_si35, test_so35, test_si36, test_so36, 
        test_si37, test_so37, test_si38, test_so38, test_si39, test_so39, 
        test_si40, test_so40, test_si41, test_so41, test_si42, test_so42, 
        test_si43, test_so43, test_si44, test_so44, test_si45, test_so45, 
        test_si46, test_so46, test_si47, test_so47, test_si48, test_so48, 
        test_si49, test_so49, test_si50, test_so50, test_si51, test_so51, 
        test_si52, test_so52, test_si53, test_so53, test_si54, test_so54, 
        test_si55, test_so55, test_si56, test_so56, test_si57, test_so57, 
        test_si58, test_so58, test_si59, test_so59, test_si60, test_so60, 
        test_si61, test_so61, test_si62, test_so62, test_si63, test_so63, 
        test_si64, test_so64, test_si65, test_so65, test_si66, test_so66, 
        test_si67, test_so67, test_si68, test_so68, test_si69, test_so69, 
        test_si70, test_so70, test_si71, test_so71, test_si72, test_so72, 
        test_si73, test_so73, test_si74, test_so74, test_si75, test_so75, 
        test_si76, test_so76, test_si77, test_so77, test_si78, test_so78, 
        test_si79, test_so79, test_si80, test_so80, test_si81, test_so81, 
        test_si82, test_so82, test_si83, test_so83, test_si84, test_so84, 
        test_si85, test_so85, test_si86, test_so86, test_si87, test_so87, 
        test_si88, test_so88, test_si89, test_so89, test_si90, test_so90, 
        test_si91, test_so91, test_si92, test_so92, test_si93, test_so93, 
        test_si94, test_so94, test_si95, test_so95, test_si96, test_so96, 
        test_si97, test_so97, test_si98, test_so98, test_si99, test_so99, 
        test_si100, test_so100 );
  input CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13,
         DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19,
         DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24,
         DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3,
         DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7,
         DATA_0_8, DATA_0_9, RESET, TM0, TM1, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10, test_si11, test_si12, test_si13, test_si14, test_si15,
         test_si16, test_si17, test_si18, test_si19, test_si20, test_si21,
         test_si22, test_si23, test_si24, test_si25, test_si26, test_si27,
         test_si28, test_si29, test_si30, test_si31, test_si32, test_si33,
         test_si34, test_si35, test_si36, test_si37, test_si38, test_si39,
         test_si40, test_si41, test_si42, test_si43, test_si44, test_si45,
         test_si46, test_si47, test_si48, test_si49, test_si50, test_si51,
         test_si52, test_si53, test_si54, test_si55, test_si56, test_si57,
         test_si58, test_si59, test_si60, test_si61, test_si62, test_si63,
         test_si64, test_si65, test_si66, test_si67, test_si68, test_si69,
         test_si70, test_si71, test_si72, test_si73, test_si74, test_si75,
         test_si76, test_si77, test_si78, test_si79, test_si80, test_si81,
         test_si82, test_si83, test_si84, test_si85, test_si86, test_si87,
         test_si88, test_si89, test_si90, test_si91, test_si92, test_si93,
         test_si94, test_si95, test_si96, test_si97, test_si98, test_si99,
         test_si100;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9, test_so1, test_so2,
         test_so3, test_so4, test_so5, test_so6, test_so7, test_so8, test_so9,
         test_so10, test_so11, test_so12, test_so13, test_so14, test_so15,
         test_so16, test_so17, test_so18, test_so19, test_so20, test_so21,
         test_so22, test_so23, test_so24, test_so25, test_so26, test_so27,
         test_so28, test_so29, test_so30, test_so31, test_so32, test_so33,
         test_so34, test_so35, test_so36, test_so37, test_so38, test_so39,
         test_so40, test_so41, test_so42, test_so43, test_so44, test_so45,
         test_so46, test_so47, test_so48, test_so49, test_so50, test_so51,
         test_so52, test_so53, test_so54, test_so55, test_so56, test_so57,
         test_so58, test_so59, test_so60, test_so61, test_so62, test_so63,
         test_so64, test_so65, test_so66, test_so67, test_so68, test_so69,
         test_so70, test_so71, test_so72, test_so73, test_so74, test_so75,
         test_so76, test_so77, test_so78, test_so79, test_so80, test_so81,
         test_so82, test_so83, test_so84, test_so85, test_so86, test_so87,
         test_so88, test_so89, test_so90, test_so91, test_so92, test_so93,
         test_so94, test_so95, test_so96, test_so97, test_so98, test_so99,
         test_so100;
  wire   test_so9, test_so10, test_so20, test_so21, test_so31, test_so32,
         test_so42, test_so43, test_so53, test_so54, test_so65, test_so66,
         test_so76, test_so77, test_so87, test_so88, test_so99, test_so100,
         WX484, WX485, WX486, WX487, WX488, WX489, WX490, WX491, WX492, WX493,
         WX494, WX495, WX496, WX497, WX498, WX499, WX500, WX501, WX502, WX503,
         WX504, WX505, WX506, WX507, WX508, WX509, WX510, WX511, WX512, WX513,
         WX514, WX515, WX516, WX517, WX518, WX520, WX521, WX522, WX523, WX524,
         WX525, WX526, WX527, WX528, WX529, WX530, WX531, WX532, WX533, WX534,
         WX535, WX536, WX537, WX538, WX539, WX540, WX541, WX542, WX543, WX544,
         WX545, WX546, WX547, WX644, WX645, n3529, WX646, WX647, n3527, WX648,
         WX649, n3525, WX650, WX652, WX653, n3521, WX654, WX655, n3519, WX656,
         WX657, n3517, WX658, WX659, n3515, WX660, WX661, n3513, WX662, WX663,
         n3511, WX664, WX665, n3509, WX666, WX667, n3507, WX668, WX669, n3505,
         WX670, WX671, n3503, WX672, WX673, n3501, WX674, WX675, n3499, WX676,
         WX677, n3497, WX678, WX679, n3495, WX680, WX681, n3493, WX682, WX683,
         n3491, WX684, WX685, n3489, WX686, WX688, WX689, n3485, WX690, WX691,
         n3483, WX692, WX693, n3481, WX694, WX695, n3479, WX696, WX697, n3477,
         WX698, WX699, n3475, WX700, WX701, n3473, WX702, WX703, n3471, WX704,
         WX705, n3469, WX706, WX707, n3467, WX708, WX709, WX710, WX711, WX712,
         WX713, WX714, WX715, WX716, WX717, WX718, WX719, WX720, WX721, WX722,
         WX724, WX725, WX726, WX727, WX728, WX729, WX730, WX731, WX732, WX733,
         WX734, WX735, WX736, WX737, WX738, WX739, WX740, WX741, WX742, WX743,
         WX744, WX745, WX746, WX747, WX748, WX749, WX750, WX751, WX752, WX753,
         WX754, WX755, WX756, WX757, WX758, WX760, WX761, WX762, WX763, WX764,
         WX765, WX766, WX767, WX768, WX769, WX770, WX771, WX772, WX773, WX774,
         WX775, WX776, WX777, WX778, WX779, WX780, WX781, WX782, WX783, WX784,
         WX785, WX786, WX787, WX788, WX789, WX790, WX791, WX792, WX793, WX794,
         WX796, WX797, WX798, WX799, WX800, WX801, WX802, WX803, WX804, WX805,
         WX806, WX807, WX808, WX809, WX810, WX811, WX812, WX813, WX814, WX815,
         WX816, WX817, WX818, WX819, WX820, WX821, WX822, WX823, WX824, WX825,
         WX826, WX827, WX828, WX829, WX830, WX832, WX833, WX834, WX835, WX836,
         WX837, WX838, WX839, WX840, WX841, WX842, WX843, WX844, WX845, WX846,
         WX847, WX848, WX849, WX850, WX851, WX852, WX853, WX854, WX855, WX856,
         WX857, WX858, WX859, WX860, WX861, WX862, WX863, WX864, WX865, WX866,
         WX868, WX869, WX870, WX871, WX872, WX873, WX874, WX875, WX876, WX877,
         WX878, WX879, WX880, WX881, WX882, WX883, WX884, WX885, WX886, WX887,
         WX888, WX889, WX890, WX891, WX892, WX893, WX894, WX895, WX896, WX897,
         WX898, WX899, WX1264, WX1266, WX1268, DFF_162_n1, WX1270, DFF_163_n1,
         WX1272, DFF_164_n1, WX1274, DFF_165_n1, WX1276, DFF_166_n1, WX1278,
         DFF_167_n1, WX1280, DFF_168_n1, WX1282, DFF_169_n1, WX1284,
         DFF_170_n1, WX1286, DFF_171_n1, WX1288, DFF_172_n1, WX1290,
         DFF_173_n1, WX1292, DFF_174_n1, WX1294, DFF_175_n1, WX1296,
         DFF_176_n1, WX1298, DFF_177_n1, WX1300, DFF_178_n1, WX1302, WX1304,
         DFF_180_n1, WX1306, DFF_181_n1, WX1308, DFF_182_n1, WX1310,
         DFF_183_n1, WX1312, DFF_184_n1, WX1314, DFF_185_n1, WX1316,
         DFF_186_n1, WX1318, DFF_187_n1, WX1320, DFF_188_n1, WX1322,
         DFF_189_n1, WX1324, DFF_190_n1, WX1326, DFF_191_n1, WX1778, n8702,
         n4033, n8701, n4032, n8700, n4031, n8699, n4030, n4029, n8696, n4028,
         n8695, n4027, n8694, n4026, n8693, n4025, n8692, n4024, n8691, n4023,
         n8690, n4022, n8689, n4021, n8688, n4020, n8687, n4019, n8686, n4018,
         n8685, n4017, n8684, n4016, n8683, n4015, n8682, n4014, n8681, n4013,
         n8680, n4012, n4011, n8677, n4010, n8676, n4009, n8675, n4008, n8674,
         n4007, n8673, n4006, n8672, n4005, n8671, n4004, WX1839, n8670, n4003,
         WX1937, n8669, WX1939, n8668, WX1941, n8667, WX1943, n8666, WX1945,
         n8665, WX1947, n8664, WX1949, n8663, WX1951, n8662, WX1953, n8661,
         WX1955, WX1957, n8658, WX1959, n8657, WX1961, n8656, WX1963, n8655,
         WX1965, n8654, WX1967, n8653, WX1969, WX1970, WX1971, WX1972, WX1973,
         WX1974, WX1975, WX1976, WX1977, WX1978, WX1979, WX1980, WX1981,
         WX1982, WX1983, WX1984, WX1985, WX1986, WX1987, WX1988, WX1989,
         WX1990, WX1991, WX1993, WX1994, WX1995, WX1996, WX1997, WX1998,
         WX1999, WX2000, WX2001, WX2002, WX2003, WX2004, WX2005, WX2006,
         WX2007, WX2008, WX2009, WX2010, WX2011, WX2012, WX2013, WX2014,
         WX2015, WX2016, WX2017, WX2018, WX2019, WX2020, WX2021, WX2022,
         WX2023, WX2024, WX2025, WX2026, WX2027, WX2029, WX2030, WX2031,
         WX2032, WX2033, WX2034, n3785, WX2035, WX2036, n3783, WX2037, WX2038,
         n3781, WX2039, WX2040, n3779, WX2041, WX2042, n3777, WX2043, WX2044,
         n3775, WX2045, WX2046, n3773, WX2047, WX2048, n3771, WX2049, WX2050,
         n3769, WX2051, WX2052, n3767, WX2053, WX2054, n3765, WX2055, WX2056,
         n3763, WX2057, WX2058, n3761, WX2059, WX2060, n3759, WX2061, WX2062,
         n3757, WX2063, WX2065, WX2066, WX2067, WX2068, WX2069, WX2070, WX2071,
         WX2072, WX2073, WX2074, WX2075, WX2076, WX2077, WX2078, WX2079,
         WX2080, WX2081, WX2082, WX2083, WX2084, WX2085, WX2086, WX2087,
         WX2088, WX2089, WX2090, WX2091, WX2092, WX2093, WX2094, WX2095,
         WX2096, WX2097, WX2098, WX2099, WX2101, WX2102, WX2103, WX2104,
         WX2105, WX2106, WX2107, WX2108, WX2109, WX2110, WX2111, WX2112,
         WX2113, WX2114, WX2115, WX2116, WX2117, WX2118, WX2119, WX2120,
         WX2121, WX2122, WX2123, WX2124, WX2125, WX2126, WX2127, WX2128,
         WX2129, WX2130, WX2131, WX2132, WX2133, WX2134, WX2135, WX2137,
         WX2138, WX2139, WX2140, WX2141, WX2142, WX2143, WX2144, WX2145,
         WX2146, WX2147, WX2148, WX2149, WX2150, WX2151, WX2152, WX2153,
         WX2154, WX2155, WX2156, WX2157, WX2158, WX2159, WX2160, WX2161,
         WX2162, WX2163, WX2164, WX2165, WX2166, WX2167, WX2168, WX2169,
         WX2170, WX2171, WX2173, WX2174, WX2175, WX2176, WX2177, WX2178,
         WX2179, WX2180, WX2181, WX2182, WX2183, WX2184, WX2185, WX2186,
         WX2187, WX2188, WX2189, WX2190, WX2191, WX2192, WX2557, DFF_352_n1,
         WX2559, DFF_353_n1, WX2561, DFF_354_n1, WX2563, DFF_355_n1, WX2565,
         DFF_356_n1, WX2567, DFF_357_n1, WX2569, DFF_358_n1, WX2571, WX2573,
         DFF_360_n1, WX2575, DFF_361_n1, WX2577, DFF_362_n1, WX2579,
         DFF_363_n1, WX2581, DFF_364_n1, WX2583, DFF_365_n1, WX2585,
         DFF_366_n1, WX2587, DFF_367_n1, WX2589, DFF_368_n1, WX2591,
         DFF_369_n1, WX2593, DFF_370_n1, WX2595, DFF_371_n1, WX2597,
         DFF_372_n1, WX2599, DFF_373_n1, WX2601, DFF_374_n1, WX2603,
         DFF_375_n1, WX2605, DFF_376_n1, WX2607, WX2609, DFF_378_n1, WX2611,
         DFF_379_n1, WX2613, DFF_380_n1, WX2615, DFF_381_n1, WX2617,
         DFF_382_n1, WX2619, DFF_383_n1, WX3071, n8644, n4002, n8643, n4001,
         n8642, n4000, n8641, n3999, n8640, n3998, n8639, n3997, n8638, n3996,
         n8637, n3995, n8636, n3994, n8635, n3993, n3992, n8632, n3991, n8631,
         n3990, n8630, n3989, n8629, n3988, n8628, n3987, n8627, n3986, n8626,
         n3985, n8625, n3984, n8624, n3983, n8623, n3982, n8622, n3981, n8621,
         n3980, n8620, n3979, n8619, n3978, n8618, n3977, n8617, n3976, n8616,
         n3975, n3974, n8613, n3973, WX3132, n8612, n3972, WX3230, n8611,
         WX3232, n8610, WX3234, n8609, WX3236, n8608, WX3238, n8607, WX3240,
         n8606, WX3242, n8605, WX3244, n8604, WX3246, n8603, WX3248, n8602,
         WX3250, n8601, WX3252, n8600, WX3254, n8599, WX3256, n8598, WX3258,
         n8597, WX3260, WX3262, WX3263, WX3264, WX3265, WX3266, WX3267, WX3268,
         WX3269, WX3270, WX3271, WX3272, WX3273, WX3274, WX3275, WX3276,
         WX3277, WX3278, WX3279, WX3280, WX3281, WX3282, WX3283, WX3284,
         WX3285, WX3286, WX3287, WX3288, WX3289, WX3290, WX3291, WX3292,
         WX3293, WX3294, WX3295, WX3296, WX3298, WX3299, WX3300, WX3301,
         WX3302, WX3303, WX3304, WX3305, WX3306, WX3307, WX3308, WX3309,
         WX3310, WX3311, WX3312, WX3313, WX3314, WX3315, WX3316, WX3317,
         WX3318, WX3319, WX3320, WX3321, WX3322, WX3323, WX3324, WX3325,
         WX3326, WX3327, n3753, WX3328, WX3329, n3751, WX3330, WX3331, n3749,
         WX3332, WX3334, WX3335, n3745, WX3336, WX3337, n3743, WX3338, WX3339,
         n3741, WX3340, WX3341, n3739, WX3342, WX3343, n3737, WX3344, WX3345,
         n3735, WX3346, WX3347, n3733, WX3348, WX3349, n3731, WX3350, WX3351,
         n3729, WX3352, WX3353, n3727, WX3354, WX3355, n3725, WX3356, WX3357,
         n3723, WX3358, WX3359, WX3360, WX3361, WX3362, WX3363, WX3364, WX3365,
         WX3366, WX3367, WX3368, WX3370, WX3371, WX3372, WX3373, WX3374,
         WX3375, WX3376, WX3377, WX3378, WX3379, WX3380, WX3381, WX3382,
         WX3383, WX3384, WX3385, WX3386, WX3387, WX3388, WX3389, WX3390,
         WX3391, WX3392, WX3393, WX3394, WX3395, WX3396, WX3397, WX3398,
         WX3399, WX3400, WX3401, WX3402, WX3403, WX3404, WX3406, WX3407,
         WX3408, WX3409, WX3410, WX3411, WX3412, WX3413, WX3414, WX3415,
         WX3416, WX3417, WX3418, WX3419, WX3420, WX3421, WX3422, WX3423,
         WX3424, WX3425, WX3426, WX3427, WX3428, WX3429, WX3430, WX3431,
         WX3432, WX3433, WX3434, WX3435, WX3436, WX3437, WX3438, WX3440,
         WX3441, WX3442, WX3443, WX3444, WX3445, WX3446, WX3447, WX3448,
         WX3449, WX3450, WX3451, WX3452, WX3453, WX3454, WX3455, WX3456,
         WX3457, WX3458, WX3459, WX3460, WX3461, WX3462, WX3463, WX3464,
         WX3465, WX3466, WX3467, WX3468, WX3469, WX3470, WX3471, WX3472,
         WX3474, WX3475, WX3476, WX3477, WX3478, WX3479, WX3480, WX3481,
         WX3482, WX3483, WX3484, WX3485, WX3850, DFF_544_n1, WX3852,
         DFF_545_n1, WX3854, DFF_546_n1, WX3856, DFF_547_n1, WX3858,
         DFF_548_n1, WX3860, DFF_549_n1, WX3862, DFF_550_n1, WX3864,
         DFF_551_n1, WX3866, DFF_552_n1, WX3868, DFF_553_n1, WX3870, WX3872,
         DFF_555_n1, WX3874, DFF_556_n1, WX3876, DFF_557_n1, WX3878,
         DFF_558_n1, WX3880, DFF_559_n1, WX3882, DFF_560_n1, WX3884,
         DFF_561_n1, WX3886, DFF_562_n1, WX3888, DFF_563_n1, WX3890,
         DFF_564_n1, WX3892, DFF_565_n1, WX3894, DFF_566_n1, WX3896,
         DFF_567_n1, WX3898, DFF_568_n1, WX3900, DFF_569_n1, WX3902,
         DFF_570_n1, WX3904, WX3906, DFF_572_n1, WX3908, DFF_573_n1, WX3910,
         DFF_574_n1, WX3912, DFF_575_n1, WX4364, n8586, n3971, n8585, n3970,
         n8584, n3969, n8583, n3968, n8582, n3967, n8581, n3966, n8580, n3965,
         n8579, n3964, n8578, n3963, n8577, n3962, n8576, n3961, n3960, n8573,
         n3959, n8572, n3958, n8571, n3957, n8570, n3956, n8569, n3955, n8568,
         n3954, n8567, n3953, n8566, n3952, n8565, n3951, n8564, n3950, n8563,
         n3949, n8562, n3948, n8561, n3947, n8560, n3946, n8559, n3945, n8558,
         n3944, n3943, n8555, n3942, WX4425, n8554, n3941, WX4523, n8553,
         WX4525, n8552, WX4527, n8551, WX4529, n8550, WX4531, n8549, WX4533,
         n8548, WX4535, n8547, WX4537, n8546, WX4539, n8545, WX4541, n8544,
         WX4543, n8543, WX4545, n8542, WX4547, n8541, WX4549, n8540, WX4551,
         WX4553, n8537, WX4555, WX4556, WX4557, WX4558, WX4559, WX4560, WX4561,
         WX4562, WX4563, WX4564, WX4565, WX4566, WX4567, WX4568, WX4569,
         WX4570, WX4571, WX4572, WX4573, WX4574, WX4575, WX4576, WX4577,
         WX4578, WX4579, WX4580, WX4581, WX4582, WX4583, WX4584, WX4585,
         WX4587, WX4588, WX4589, WX4590, WX4591, WX4592, WX4593, WX4594,
         WX4595, WX4596, WX4597, WX4598, WX4599, WX4600, WX4601, WX4602,
         WX4603, WX4604, WX4605, WX4606, WX4607, WX4608, WX4609, WX4610,
         WX4611, WX4612, WX4613, WX4614, WX4615, WX4616, WX4617, WX4618,
         WX4619, WX4621, WX4622, n3719, WX4623, WX4624, n3717, WX4625, WX4626,
         n3715, WX4627, WX4628, n3713, WX4629, WX4630, n3711, WX4631, WX4632,
         n3709, WX4633, WX4634, n3707, WX4635, WX4636, n3705, WX4637, WX4638,
         n3703, WX4639, WX4640, n3701, WX4641, WX4642, n3699, WX4643, WX4644,
         n3697, WX4645, WX4646, n3695, WX4647, WX4648, n3693, WX4649, WX4650,
         n3691, WX4651, WX4652, WX4653, WX4655, WX4656, WX4657, WX4658, WX4659,
         WX4660, WX4661, WX4662, WX4663, WX4664, WX4665, WX4666, WX4667,
         WX4668, WX4669, WX4670, WX4671, WX4672, WX4673, WX4674, WX4675,
         WX4676, WX4677, WX4678, WX4679, WX4680, WX4681, WX4682, WX4683,
         WX4684, WX4685, WX4686, WX4687, WX4689, WX4690, WX4691, WX4692,
         WX4693, WX4694, WX4695, WX4696, WX4697, WX4698, WX4699, WX4700,
         WX4701, WX4702, WX4703, WX4704, WX4705, WX4706, WX4707, WX4708,
         WX4709, WX4710, WX4711, WX4712, WX4713, WX4714, WX4715, WX4716,
         WX4717, WX4718, WX4719, WX4720, WX4721, WX4723, WX4724, WX4725,
         WX4726, WX4727, WX4728, WX4729, WX4730, WX4731, WX4732, WX4733,
         WX4734, WX4735, WX4736, WX4737, WX4738, WX4739, WX4740, WX4741,
         WX4742, WX4743, WX4744, WX4745, WX4746, WX4747, WX4748, WX4749,
         WX4750, WX4751, WX4752, WX4753, WX4754, WX4755, WX4757, WX4758,
         WX4759, WX4760, WX4761, WX4762, WX4763, WX4764, WX4765, WX4766,
         WX4767, WX4768, WX4769, WX4770, WX4771, WX4772, WX4773, WX4774,
         WX4775, WX4776, WX4777, WX4778, WX5143, DFF_736_n1, WX5145,
         DFF_737_n1, WX5147, DFF_738_n1, WX5149, DFF_739_n1, WX5151,
         DFF_740_n1, WX5153, WX5155, DFF_742_n1, WX5157, DFF_743_n1, WX5159,
         DFF_744_n1, WX5161, DFF_745_n1, WX5163, DFF_746_n1, WX5165,
         DFF_747_n1, WX5167, DFF_748_n1, WX5169, DFF_749_n1, WX5171,
         DFF_750_n1, WX5173, DFF_751_n1, WX5175, DFF_752_n1, WX5177,
         DFF_753_n1, WX5179, DFF_754_n1, WX5181, DFF_755_n1, WX5183,
         DFF_756_n1, WX5185, DFF_757_n1, WX5187, WX5189, DFF_759_n1, WX5191,
         DFF_760_n1, WX5193, DFF_761_n1, WX5195, DFF_762_n1, WX5197,
         DFF_763_n1, WX5199, DFF_764_n1, WX5201, DFF_765_n1, WX5203,
         DFF_766_n1, WX5205, DFF_767_n1, WX5657, n8528, n3940, n8527, n3939,
         n8526, n3938, n8525, n3937, n8524, n3936, n8523, n3935, n3934, n8520,
         n3933, n8519, n3932, n8518, n3931, n8517, n3930, n8516, n3929, n8515,
         n3928, n8514, n3927, n8513, n3926, n8512, n3925, n8511, n3924, n8510,
         n3923, n8509, n3922, n8508, n3921, n8507, n3920, n8506, n3919, n8505,
         n3918, n3917, n8502, n3916, n8501, n3915, n8500, n3914, n8499, n3913,
         n8498, n3912, n8497, n3911, WX5718, n8496, n3910, WX5816, n8495,
         WX5818, n8494, WX5820, n8493, WX5822, n8492, WX5824, n8491, WX5826,
         n8490, WX5828, n8489, WX5830, n8488, WX5832, n8487, WX5834, WX5836,
         n8484, WX5838, n8483, WX5840, n8482, WX5842, n8481, WX5844, n8480,
         WX5846, n8479, WX5848, WX5849, WX5850, WX5851, WX5852, WX5853, WX5854,
         WX5855, WX5856, WX5857, WX5858, WX5859, WX5860, WX5861, WX5862,
         WX5863, WX5864, WX5865, WX5866, WX5867, WX5868, WX5870, WX5871,
         WX5872, WX5873, WX5874, WX5875, WX5876, WX5877, WX5878, WX5879,
         WX5880, WX5881, WX5882, WX5883, WX5884, WX5885, WX5886, WX5887,
         WX5888, WX5889, WX5890, WX5891, WX5892, WX5893, WX5894, WX5895,
         WX5896, WX5897, WX5898, WX5899, WX5900, WX5901, WX5902, WX5904,
         WX5905, WX5906, WX5907, WX5908, WX5909, WX5910, WX5911, WX5912,
         WX5913, n3689, WX5914, WX5915, n3687, WX5916, WX5917, n3685, WX5918,
         WX5919, n3683, WX5920, WX5921, n3681, WX5922, WX5923, n3679, WX5924,
         WX5925, n3677, WX5926, WX5927, n3675, WX5928, WX5929, n3673, WX5930,
         WX5931, n3671, WX5932, WX5933, n3669, WX5934, WX5935, n3667, WX5936,
         WX5938, WX5939, n3663, WX5940, WX5941, n3661, WX5942, WX5943, n3659,
         WX5944, WX5945, WX5946, WX5947, WX5948, WX5949, WX5950, WX5951,
         WX5952, WX5953, WX5954, WX5955, WX5956, WX5957, WX5958, WX5959,
         WX5960, WX5961, WX5962, WX5963, WX5964, WX5965, WX5966, WX5967,
         WX5968, WX5969, WX5970, WX5972, WX5973, WX5974, WX5975, WX5976,
         WX5977, WX5978, WX5979, WX5980, WX5981, WX5982, WX5983, WX5984,
         WX5985, WX5986, WX5987, WX5988, WX5989, WX5990, WX5991, WX5992,
         WX5993, WX5994, WX5995, WX5996, WX5997, WX5998, WX5999, WX6000,
         WX6001, WX6002, WX6003, WX6004, WX6006, WX6007, WX6008, WX6009,
         WX6010, WX6011, WX6012, WX6013, WX6014, WX6015, WX6016, WX6017,
         WX6018, WX6019, WX6020, WX6021, WX6022, WX6023, WX6024, WX6025,
         WX6026, WX6027, WX6028, WX6029, WX6030, WX6031, WX6032, WX6033,
         WX6034, WX6035, WX6036, WX6037, WX6038, WX6040, WX6041, WX6042,
         WX6043, WX6044, WX6045, WX6046, WX6047, WX6048, WX6049, WX6050,
         WX6051, WX6052, WX6053, WX6054, WX6055, WX6056, WX6057, WX6058,
         WX6059, WX6060, WX6061, WX6062, WX6063, WX6064, WX6065, WX6066,
         WX6067, WX6068, WX6069, WX6070, WX6071, WX6436, WX6438, DFF_929_n1,
         WX6440, DFF_930_n1, WX6442, DFF_931_n1, WX6444, DFF_932_n1, WX6446,
         DFF_933_n1, WX6448, DFF_934_n1, WX6450, DFF_935_n1, WX6452,
         DFF_936_n1, WX6454, DFF_937_n1, WX6456, DFF_938_n1, WX6458,
         DFF_939_n1, WX6460, DFF_940_n1, WX6462, DFF_941_n1, WX6464,
         DFF_942_n1, WX6466, DFF_943_n1, WX6468, DFF_944_n1, WX6470, WX6472,
         DFF_946_n1, WX6474, DFF_947_n1, WX6476, DFF_948_n1, WX6478,
         DFF_949_n1, WX6480, DFF_950_n1, WX6482, DFF_951_n1, WX6484,
         DFF_952_n1, WX6486, DFF_953_n1, WX6488, DFF_954_n1, WX6490,
         DFF_955_n1, WX6492, DFF_956_n1, WX6494, DFF_957_n1, WX6496,
         DFF_958_n1, WX6498, DFF_959_n1, WX6950, n8470, n3909, n3908, n8467,
         n3907, n8466, n3906, n8465, n3905, n8464, n3904, n8463, n3903, n8462,
         n3902, n8461, n3901, n8460, n3900, n8459, n3899, n8458, n3898, n8457,
         n3897, n8456, n3896, n8455, n3895, n8454, n3894, n8453, n3893, n8452,
         n3892, n3891, n8449, n3890, n8448, n3889, n8447, n3888, n8446, n3887,
         n8445, n3886, n8444, n3885, n8443, n3884, n8442, n3883, n8441, n3882,
         n8440, n3881, n8439, n3880, WX7011, n8438, n3879, WX7109, n8437,
         WX7111, n8436, WX7113, n8435, WX7115, n8434, WX7117, WX7119, n8431,
         WX7121, n8430, WX7123, n8429, WX7125, n8428, WX7127, n8427, WX7129,
         n8426, WX7131, n8425, WX7133, n8424, WX7135, n8423, WX7137, n8422,
         WX7139, n8421, WX7141, WX7142, WX7143, WX7144, WX7145, WX7146, WX7147,
         WX7148, WX7149, WX7150, WX7151, WX7153, WX7154, WX7155, WX7156,
         WX7157, WX7158, WX7159, WX7160, WX7161, WX7162, WX7163, WX7164,
         WX7165, WX7166, WX7167, WX7168, WX7169, WX7170, WX7171, WX7172,
         WX7173, WX7174, WX7175, WX7176, WX7177, WX7178, WX7179, WX7180,
         WX7181, WX7182, WX7183, WX7184, WX7185, WX7187, WX7188, WX7189,
         WX7190, WX7191, WX7192, WX7193, WX7194, WX7195, WX7196, WX7197,
         WX7198, WX7199, WX7200, WX7201, WX7202, WX7203, WX7204, WX7205,
         WX7206, n3657, WX7207, WX7208, n3655, WX7209, WX7210, n3653, WX7211,
         WX7212, n3651, WX7213, WX7214, n3649, WX7215, WX7216, n3647, WX7217,
         WX7218, n3645, WX7219, WX7221, WX7222, n3641, WX7223, WX7224, n3639,
         WX7225, WX7226, n3637, WX7227, WX7228, n3635, WX7229, WX7230, n3633,
         WX7231, WX7232, n3631, WX7233, WX7234, n3629, WX7235, WX7236, n3627,
         WX7237, WX7238, WX7239, WX7240, WX7241, WX7242, WX7243, WX7244,
         WX7245, WX7246, WX7247, WX7248, WX7249, WX7250, WX7251, WX7252,
         WX7253, WX7255, WX7256, WX7257, WX7258, WX7259, WX7260, WX7261,
         WX7262, WX7263, WX7264, WX7265, WX7266, WX7267, WX7268, WX7269,
         WX7270, WX7271, WX7272, WX7273, WX7274, WX7275, WX7276, WX7277,
         WX7278, WX7279, WX7280, WX7281, WX7282, WX7283, WX7284, WX7285,
         WX7286, WX7287, WX7289, WX7290, WX7291, WX7292, WX7293, WX7294,
         WX7295, WX7296, WX7297, WX7298, WX7299, WX7300, WX7301, WX7302,
         WX7303, WX7304, WX7305, WX7306, WX7307, WX7308, WX7309, WX7310,
         WX7311, WX7312, WX7313, WX7314, WX7315, WX7316, WX7317, WX7318,
         WX7319, WX7320, WX7321, WX7323, WX7324, WX7325, WX7326, WX7327,
         WX7328, WX7329, WX7330, WX7331, WX7332, WX7333, WX7334, WX7335,
         WX7336, WX7337, WX7338, WX7339, WX7340, WX7341, WX7342, WX7343,
         WX7344, WX7345, WX7346, WX7347, WX7348, WX7349, WX7350, WX7351,
         WX7352, WX7353, WX7354, WX7355, WX7357, WX7358, WX7359, WX7360,
         WX7361, WX7362, WX7363, WX7364, WX7729, DFF_1120_n1, WX7731,
         DFF_1121_n1, WX7733, DFF_1122_n1, WX7735, DFF_1123_n1, WX7737,
         DFF_1124_n1, WX7739, DFF_1125_n1, WX7741, DFF_1126_n1, WX7743,
         DFF_1127_n1, WX7745, DFF_1128_n1, WX7747, DFF_1129_n1, WX7749,
         DFF_1130_n1, WX7751, DFF_1131_n1, WX7753, WX7755, DFF_1133_n1, WX7757,
         DFF_1134_n1, WX7759, DFF_1135_n1, WX7761, DFF_1136_n1, WX7763,
         DFF_1137_n1, WX7765, DFF_1138_n1, WX7767, DFF_1139_n1, WX7769,
         DFF_1140_n1, WX7771, DFF_1141_n1, WX7773, DFF_1142_n1, WX7775,
         DFF_1143_n1, WX7777, DFF_1144_n1, WX7779, DFF_1145_n1, WX7781,
         DFF_1146_n1, WX7783, DFF_1147_n1, WX7785, DFF_1148_n1, WX7787, WX7789,
         DFF_1150_n1, WX7791, DFF_1151_n1, WX8243, n8411, n3878, n8410, n3877,
         n8409, n3876, n8408, n3875, n8407, n3874, n8406, n3873, n8405, n3872,
         n8404, n3871, n8403, n3870, n8402, n3869, n8401, n3868, n8400, n3867,
         n8399, n3866, n3865, n8396, n3864, n8395, n3863, n8394, n3862, n8393,
         n3861, n8392, n3860, n8391, n3859, n8390, n3858, n8389, n3857, n8388,
         n3856, n8387, n3855, n8386, n3854, n8385, n3853, n8384, n3852, n8383,
         n3851, n8382, n3850, n8381, n3849, WX8304, n3848, WX8402, n8378,
         WX8404, n8377, WX8406, n8376, WX8408, n8375, WX8410, n8374, WX8412,
         n8373, WX8414, n8372, WX8416, n8371, WX8418, n8370, WX8420, n8369,
         WX8422, n8368, WX8424, n8367, WX8426, n8366, WX8428, n8365, WX8430,
         n8364, WX8432, n8363, WX8434, WX8436, WX8437, WX8438, WX8439, WX8440,
         WX8441, WX8442, WX8443, WX8444, WX8445, WX8446, WX8447, WX8448,
         WX8449, WX8450, WX8451, WX8452, WX8453, WX8454, WX8455, WX8456,
         WX8457, WX8458, WX8459, WX8460, WX8461, WX8462, WX8463, WX8464,
         WX8465, WX8466, WX8467, WX8468, WX8470, WX8471, WX8472, WX8473,
         WX8474, WX8475, WX8476, WX8477, WX8478, WX8479, WX8480, WX8481,
         WX8482, WX8483, WX8484, WX8485, WX8486, WX8487, WX8488, WX8489,
         WX8490, WX8491, WX8492, WX8493, WX8494, WX8495, WX8496, WX8497,
         WX8498, WX8499, n3625, WX8500, WX8501, n3623, WX8502, WX8504, WX8505,
         n3619, WX8506, WX8507, n3617, WX8508, WX8509, n3615, WX8510, WX8511,
         n3613, WX8512, WX8513, n3611, WX8514, WX8515, n3609, WX8516, WX8517,
         n3607, WX8518, WX8519, n3605, WX8520, WX8521, n3603, WX8522, WX8523,
         n3601, WX8524, WX8525, n3599, WX8526, WX8527, n3597, WX8528, WX8529,
         n3595, WX8530, WX8531, WX8532, WX8533, WX8534, WX8535, WX8536, WX8538,
         WX8539, WX8540, WX8541, WX8542, WX8543, WX8544, WX8545, WX8546,
         WX8547, WX8548, WX8549, WX8550, WX8551, WX8552, WX8553, WX8554,
         WX8555, WX8556, WX8557, WX8558, WX8559, WX8560, WX8561, WX8562,
         WX8563, WX8564, WX8565, WX8566, WX8567, WX8568, WX8569, WX8570,
         WX8572, WX8573, WX8574, WX8575, WX8576, WX8577, WX8578, WX8579,
         WX8580, WX8581, WX8582, WX8583, WX8584, WX8585, WX8586, WX8587,
         WX8588, WX8589, WX8590, WX8591, WX8592, WX8593, WX8594, WX8595,
         WX8596, WX8597, WX8598, WX8599, WX8600, WX8601, WX8602, WX8603,
         WX8604, WX8606, WX8607, WX8608, WX8609, WX8610, WX8611, WX8612,
         WX8613, WX8614, WX8615, WX8616, WX8617, WX8618, WX8619, WX8620,
         WX8621, WX8622, WX8623, WX8624, WX8625, WX8626, WX8627, WX8628,
         WX8629, WX8630, WX8631, WX8632, WX8633, WX8634, WX8635, WX8636,
         WX8637, WX8638, WX8640, WX8641, WX8642, WX8643, WX8644, WX8645,
         WX8646, WX8647, WX8648, WX8649, WX8650, WX8651, WX8652, WX8653,
         WX8654, WX8655, WX8656, WX8657, WX9022, DFF_1312_n1, WX9024,
         DFF_1313_n1, WX9026, DFF_1314_n1, WX9028, DFF_1315_n1, WX9030,
         DFF_1316_n1, WX9032, DFF_1317_n1, WX9034, DFF_1318_n1, WX9036, WX9038,
         DFF_1320_n1, WX9040, DFF_1321_n1, WX9042, DFF_1322_n1, WX9044,
         DFF_1323_n1, WX9046, DFF_1324_n1, WX9048, DFF_1325_n1, WX9050,
         DFF_1326_n1, WX9052, DFF_1327_n1, WX9054, DFF_1328_n1, WX9056,
         DFF_1329_n1, WX9058, DFF_1330_n1, WX9060, DFF_1331_n1, WX9062,
         DFF_1332_n1, WX9064, DFF_1333_n1, WX9066, DFF_1334_n1, WX9068,
         DFF_1335_n1, WX9070, WX9072, DFF_1337_n1, WX9074, DFF_1338_n1, WX9076,
         DFF_1339_n1, WX9078, DFF_1340_n1, WX9080, DFF_1341_n1, WX9082,
         DFF_1342_n1, WX9084, DFF_1343_n1, WX9536, n8353, n3847, n8352, n3846,
         n8351, n3845, n8350, n3844, n8349, n3843, n8348, n3842, n8347, n3841,
         n8346, n3840, n3839, n8343, n3838, n8342, n3837, n8341, n3836, n8340,
         n3835, n8339, n3834, n8338, n3833, n8337, n3832, n8336, n3831, n8335,
         n3830, n8334, n3829, n8333, n3828, n8332, n3827, n8331, n3826, n8330,
         n3825, n8329, n3824, n8328, n3823, n3822, n8325, n3821, n8324, n3820,
         n8323, n3819, n8322, n3818, WX9597, n8321, n3817, WX9695, n8320,
         WX9697, n8319, WX9699, n8318, WX9701, n8317, WX9703, n8316, WX9705,
         n8315, WX9707, n8314, WX9709, n8313, WX9711, n8312, WX9713, n8311,
         WX9715, n8310, WX9717, WX9719, n8307, WX9721, n8306, WX9723, n8305,
         WX9725, n8304, WX9727, WX9728, WX9729, WX9730, WX9731, WX9732, WX9733,
         WX9734, WX9735, WX9736, WX9737, WX9738, WX9739, WX9740, WX9741,
         WX9742, WX9743, WX9744, WX9745, WX9746, WX9747, WX9748, WX9749,
         WX9750, WX9751, WX9753, WX9754, WX9755, WX9756, WX9757, WX9758,
         WX9759, WX9760, WX9761, WX9762, WX9763, WX9764, WX9765, WX9766,
         WX9767, WX9768, WX9769, WX9770, WX9771, WX9772, WX9773, WX9774,
         WX9775, WX9776, WX9777, WX9778, WX9779, WX9780, WX9781, WX9782,
         WX9783, WX9784, WX9785, WX9787, WX9788, WX9789, WX9790, WX9791,
         WX9792, n3593, WX9793, WX9794, n3591, WX9795, WX9796, n3589, WX9797,
         WX9798, n3587, WX9799, WX9800, n3585, WX9801, WX9802, n3583, WX9803,
         WX9804, n3581, WX9805, WX9806, n3579, WX9807, WX9808, n3577, WX9809,
         WX9810, n3575, WX9811, WX9812, n3573, WX9813, WX9814, n3571, WX9815,
         WX9816, n3569, WX9817, WX9818, n3567, WX9819, WX9821, WX9822, n3563,
         WX9823, WX9824, WX9825, WX9826, WX9827, WX9828, WX9829, WX9830,
         WX9831, WX9832, WX9833, WX9834, WX9835, WX9836, WX9837, WX9838,
         WX9839, WX9840, WX9841, WX9842, WX9843, WX9844, WX9845, WX9846,
         WX9847, WX9848, WX9849, WX9850, WX9851, WX9852, WX9853, WX9855,
         WX9856, WX9857, WX9858, WX9859, WX9860, WX9861, WX9862, WX9863,
         WX9864, WX9865, WX9866, WX9867, WX9868, WX9869, WX9870, WX9871,
         WX9872, WX9873, WX9874, WX9875, WX9876, WX9877, WX9878, WX9879,
         WX9880, WX9881, WX9882, WX9883, WX9884, WX9885, WX9886, WX9887,
         WX9889, WX9890, WX9891, WX9892, WX9893, WX9894, WX9895, WX9896,
         WX9897, WX9898, WX9899, WX9900, WX9901, WX9902, WX9903, WX9904,
         WX9905, WX9906, WX9907, WX9908, WX9909, WX9910, WX9911, WX9912,
         WX9913, WX9914, WX9915, WX9916, WX9917, WX9918, WX9919, WX9920,
         WX9921, WX9923, WX9924, WX9925, WX9926, WX9927, WX9928, WX9929,
         WX9930, WX9931, WX9932, WX9933, WX9934, WX9935, WX9936, WX9937,
         WX9938, WX9939, WX9940, WX9941, WX9942, WX9943, WX9944, WX9945,
         WX9946, WX9947, WX9948, WX9949, WX9950, WX10315, DFF_1504_n1, WX10317,
         DFF_1505_n1, WX10319, WX10321, DFF_1507_n1, WX10323, DFF_1508_n1,
         WX10325, DFF_1509_n1, WX10327, DFF_1510_n1, WX10329, DFF_1511_n1,
         WX10331, DFF_1512_n1, WX10333, DFF_1513_n1, WX10335, DFF_1514_n1,
         WX10337, DFF_1515_n1, WX10339, DFF_1516_n1, WX10341, DFF_1517_n1,
         WX10343, DFF_1518_n1, WX10345, DFF_1519_n1, WX10347, DFF_1520_n1,
         WX10349, DFF_1521_n1, WX10351, DFF_1522_n1, WX10353, WX10355,
         DFF_1524_n1, WX10357, DFF_1525_n1, WX10359, DFF_1526_n1, WX10361,
         DFF_1527_n1, WX10363, DFF_1528_n1, WX10365, DFF_1529_n1, WX10367,
         DFF_1530_n1, WX10369, DFF_1531_n1, WX10371, DFF_1532_n1, WX10373,
         DFF_1533_n1, WX10375, DFF_1534_n1, WX10377, DFF_1535_n1, WX10829,
         n8295, n3816, n8294, n3815, n8293, n3814, n3813, n8290, n3812, n8289,
         n3811, n8288, n3810, n8287, n3809, n8286, n3808, n8285, n3807, n8284,
         n3806, n8283, n3805, n8282, n3804, n8281, n3803, n8280, n3802, n8279,
         n3801, n8278, n3800, n8277, n3799, n8276, n3798, n8275, n3797, n3796,
         n8272, n3795, n8271, n3794, n8270, n3793, n8269, n3792, n8268, n3791,
         n8267, n3790, n8266, n3789, n8265, n3788, n8264, n3787, WX10890,
         n8263, n3786, WX10988, n8262, WX10990, n8261, WX10992, n8260, WX10994,
         n8259, WX10996, n8258, WX10998, n8257, WX11000, WX11002, n8254,
         WX11004, n8253, WX11006, n8252, WX11008, n8251, WX11010, n8250,
         WX11012, n8249, WX11014, n8248, WX11016, n8247, WX11018, n8246,
         WX11020, WX11021, WX11022, WX11023, WX11024, WX11025, WX11026,
         WX11027, WX11028, WX11029, WX11030, WX11031, WX11032, WX11033,
         WX11034, WX11036, WX11037, WX11038, WX11039, WX11040, WX11041,
         WX11042, WX11043, WX11044, WX11045, WX11046, WX11047, WX11048,
         WX11049, WX11050, WX11051, WX11052, WX11053, WX11054, WX11055,
         WX11056, WX11057, WX11058, WX11059, WX11060, WX11061, WX11062,
         WX11063, WX11064, WX11065, WX11066, WX11067, WX11068, WX11070,
         WX11071, WX11072, WX11073, WX11074, WX11075, WX11076, WX11077,
         WX11078, WX11079, WX11080, WX11081, WX11082, WX11083, WX11084,
         WX11085, n3561, WX11086, WX11087, n3559, WX11088, WX11089, n3557,
         WX11090, WX11091, n3555, WX11092, WX11093, n3553, WX11094, WX11095,
         n3551, WX11096, WX11097, n3549, WX11098, WX11099, n3547, WX11100,
         WX11101, n3545, WX11102, WX11104, WX11105, n3541, WX11106, WX11107,
         n3539, WX11108, WX11109, n3537, WX11110, WX11111, n3535, WX11112,
         WX11113, n3533, WX11114, WX11115, n3531, WX11116, WX11117, WX11118,
         WX11119, WX11120, WX11121, WX11122, WX11123, WX11124, WX11125,
         WX11126, WX11127, WX11128, WX11129, WX11130, WX11131, WX11132,
         WX11133, WX11134, WX11135, WX11136, WX11138, WX11139, WX11140,
         WX11141, WX11142, WX11143, WX11144, WX11145, WX11146, WX11147,
         WX11148, WX11149, WX11150, WX11151, WX11152, WX11153, WX11154,
         WX11155, WX11156, WX11155_Tj_Payload, test_se_Trojan, WX11157,
         WX11158, WX11159, WX11160, WX11161, WX11162, WX11163, WX11164,
         WX11165, WX11166, WX11167, WX11168, WX11169, WX11170, WX11172,
         WX11173, WX11174, WX11175, WX11176, WX11177, WX11178, WX11179,
         WX11180, WX11181, WX11182, WX11183, WX11184, WX11185, WX11186,
         WX11187, WX11188, WX11189, WX11190, WX11191, WX11192, WX11193,
         WX11194, WX11195, WX11196, WX11197, WX11198, WX11199, WX11200,
         WX11201, WX11202, WX11203, WX11204, WX11206, WX11207, WX11208,
         WX11209, WX11210, WX11211, WX11212, WX11213, WX11214, WX11215,
         WX11216, WX11217, WX11218, WX11219, WX11220, WX11221, WX11222,
         WX11223, WX11224, WX11225, WX11226, WX11227, WX11228, WX11229,
         WX11230, WX11231, WX11232, WX11233, WX11234, WX11235, WX11236,
         WX11237, WX11238, WX11240, WX11241, WX11242, WX11243, WX11608,
         DFF_1696_n1, WX11610, DFF_1697_n1, WX11612, DFF_1698_n1, WX11614,
         DFF_1699_n1, WX11616, DFF_1700_n1, WX11618, DFF_1701_n1, WX11620,
         DFF_1702_n1, WX11622, DFF_1703_n1, WX11624, DFF_1704_n1, WX11626,
         DFF_1705_n1, WX11628, DFF_1706_n1, WX11630, DFF_1707_n1, WX11632,
         DFF_1708_n1, WX11634, DFF_1709_n1, WX11636, WX11638, DFF_1711_n1,
         WX11640, DFF_1712_n1, WX11642, DFF_1713_n1, WX11644, DFF_1714_n1,
         WX11646, DFF_1715_n1, WX11648, DFF_1716_n1, WX11650, DFF_1717_n1,
         WX11652, DFF_1718_n1, WX11654, DFF_1719_n1, WX11656, DFF_1720_n1,
         WX11658, DFF_1721_n1, WX11660, DFF_1722_n1, WX11662, DFF_1723_n1,
         WX11664, DFF_1724_n1, WX11666, DFF_1725_n1, WX11668, DFF_1726_n1,
         WX11670, n2245, n2153, n3278, n2152, n2148, Tj_OUT1, Tj_OUT2, Tj_OUT3,
         Tj_OUT4, Tj_OUT1234, Tj_OUT5, Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678,
         test_se_NOT, Tj_Trigger, Trojan_SE, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n2182, n9028, n9029, n9030, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9275, n9276, n9277, n9279, n9280, n9281, n9283, n9284,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9304, n9305, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9350, n9351, n9352, n9354, n9355, n9356, n9358, n9359, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9370, n9371, n9372, n9374,
         n9375, n9376, n9378, n9379, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9394, n9395, n9396, n9398,
         n9399, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9443, n9444, n9445, n9447, n9448, n9449, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9464,
         n9465, n9466, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9484, n9485, n9486, n9487,
         n9488, n9489, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, U3558_n1, U3871_n1, U3991_n1, U5716_n1, U5717_n1, U5718_n1,
         U5719_n1, U5720_n1, U5721_n1, U5722_n1, U5723_n1, U5724_n1, U5725_n1,
         U5726_n1, U5727_n1, U5728_n1, U5729_n1, U5730_n1, U5731_n1, U5732_n1,
         U5733_n1, U5734_n1, U5735_n1, U5736_n1, U5737_n1, U5738_n1, U5739_n1,
         U5740_n1, U5741_n1, U5742_n1, U5743_n1, U5744_n1, U5745_n1, U5746_n1,
         U5747_n1, U5748_n1, U5749_n1, U5750_n1, U5751_n1, U5752_n1, U5753_n1,
         U5754_n1, U5755_n1, U5756_n1, U5757_n1, U5758_n1, U5759_n1, U5760_n1,
         U5761_n1, U5762_n1, U5763_n1, U5764_n1, U5765_n1, U5766_n1, U5767_n1,
         U5768_n1, U5769_n1, U5770_n1, U5771_n1, U5772_n1, U5773_n1, U5774_n1,
         U5775_n1, U5776_n1, U5777_n1, U5778_n1, U5779_n1, U5780_n1, U5781_n1,
         U5782_n1, U5783_n1, U5784_n1, U5785_n1, U5786_n1, U5787_n1, U5788_n1,
         U5789_n1, U5790_n1, U5791_n1, U5792_n1, U5793_n1, U5794_n1, U5795_n1,
         U5796_n1, U5797_n1, U5798_n1, U5799_n1, U5800_n1, U5801_n1, U5802_n1,
         U5803_n1, U5804_n1, U5805_n1, U5806_n1, U5807_n1, U5808_n1, U5809_n1,
         U5810_n1, U5811_n1, U5812_n1, U5813_n1, U5814_n1, U5815_n1, U5816_n1,
         U5817_n1, U5818_n1, U5819_n1, U5820_n1, U5821_n1, U5822_n1, U5823_n1,
         U5824_n1, U5825_n1, U5826_n1, U5827_n1, U5828_n1, U5829_n1, U5830_n1,
         U5831_n1, U5832_n1, U5833_n1, U5834_n1, U5835_n1, U5836_n1, U5837_n1,
         U5838_n1, U5839_n1, U5840_n1, U5841_n1, U5842_n1, U5843_n1, U5844_n1,
         U5845_n1, U5846_n1, U5847_n1, U5848_n1, U5849_n1, U5850_n1, U5851_n1,
         U5852_n1, U5853_n1, U5854_n1, U5855_n1, U5856_n1, U5857_n1, U5858_n1,
         U5859_n1, U5860_n1, U5861_n1, U5862_n1, U5863_n1, U5864_n1, U5865_n1,
         U5866_n1, U5867_n1, U5868_n1, U5869_n1, U5870_n1, U5871_n1, U5872_n1,
         U5873_n1, U5874_n1, U5875_n1, U5876_n1, U5877_n1, U5878_n1, U5879_n1,
         U5880_n1, U5881_n1, U5882_n1, U5883_n1, U5884_n1, U5885_n1, U5886_n1,
         U5887_n1, U5888_n1, U5889_n1, U5890_n1, U5891_n1, U5892_n1, U5893_n1,
         U5894_n1, U5895_n1, U5896_n1, U5897_n1, U5898_n1, U5899_n1, U5900_n1,
         U5901_n1, U5902_n1, U5903_n1, U5904_n1, U5905_n1, U5906_n1, U5907_n1,
         U5908_n1, U5909_n1, U5910_n1, U5911_n1, U5912_n1, U5913_n1, U5914_n1,
         U5915_n1, U5916_n1, U5917_n1, U5918_n1, U5919_n1, U5920_n1, U5921_n1,
         U5922_n1, U5923_n1, U5924_n1, U5925_n1, U5926_n1, U5927_n1, U5928_n1,
         U5929_n1, U5930_n1, U5931_n1, U5932_n1, U5933_n1, U5934_n1, U5935_n1,
         U5936_n1, U5937_n1, U5938_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1,
         U5943_n1, U5944_n1, U5945_n1, U5946_n1, U5947_n1, U5948_n1, U5949_n1,
         U5950_n1, U5951_n1, U5952_n1, U5953_n1, U5954_n1, U5955_n1, U5956_n1,
         U5957_n1, U5958_n1, U5959_n1, U5960_n1, U5961_n1, U5962_n1, U5963_n1,
         U5964_n1, U5965_n1, U5966_n1, U5967_n1, U5968_n1, U5969_n1, U5970_n1,
         U5971_n1, U5972_n1, U5973_n1, U5974_n1, U5975_n1, U5976_n1, U5977_n1,
         U5978_n1, U5979_n1, U5980_n1, U5981_n1, U5982_n1, U5983_n1, U5984_n1,
         U5985_n1, U5986_n1, U5987_n1, U5988_n1, U5989_n1, U5990_n1, U5991_n1,
         U5992_n1, U5993_n1, U5994_n1, U5995_n1, U5996_n1, U5997_n1, U5998_n1,
         U5999_n1, U6000_n1, U6001_n1, U6002_n1, U6003_n1, U6004_n1, U6005_n1,
         U6006_n1, U6007_n1, U6008_n1, U6009_n1, U6010_n1, U6011_n1, U6012_n1,
         U6013_n1, U6014_n1, U6015_n1, U6016_n1, U6017_n1, U6018_n1, U6019_n1,
         U6020_n1, U6021_n1, U6022_n1, U6023_n1, U6024_n1, U6025_n1, U6026_n1,
         U6027_n1, U6028_n1, U6029_n1, U6030_n1, U6031_n1, U6032_n1, U6033_n1,
         U6034_n1, U6035_n1, U6036_n1, U6037_n1, U6038_n1, U6039_n1, U6040_n1,
         U6041_n1, U6042_n1, U6043_n1, U6044_n1, U6045_n1, U6046_n1, U6047_n1,
         U6048_n1, U6049_n1, U6050_n1, U6051_n1, U6052_n1, U6053_n1, U6054_n1,
         U6055_n1, U6056_n1, U6057_n1, U6058_n1, U6059_n1, U6060_n1, U6061_n1,
         U6062_n1, U6063_n1, U6064_n1, U6065_n1, U6066_n1, U6067_n1, U6068_n1,
         U6069_n1, U6070_n1, U6071_n1, U6072_n1, U6073_n1, U6074_n1, U6075_n1,
         U6076_n1, U6077_n1, U6078_n1, U6079_n1, U6080_n1, U6081_n1, U6082_n1,
         U6083_n1, U6084_n1, U6085_n1, U6086_n1, U6087_n1, U6088_n1, U6089_n1,
         U6090_n1, U6091_n1, U6092_n1, U6093_n1, U6094_n1, U6095_n1, U6096_n1,
         U6097_n1, U6098_n1, U6099_n1, U6100_n1, U6101_n1, U6102_n1, U6103_n1,
         U6104_n1, U6105_n1, U6106_n1, U6107_n1, U6108_n1, U6109_n1, U6110_n1,
         U6111_n1, U6112_n1, U6113_n1, U6114_n1, U6115_n1, U6116_n1, U6117_n1,
         U6118_n1, U6119_n1, U6120_n1, U6121_n1, U6122_n1, U6123_n1, U6124_n1,
         U6125_n1, U6126_n1, U6127_n1, U6128_n1, U6129_n1, U6130_n1, U6131_n1,
         U6132_n1, U6133_n1, U6134_n1, U6135_n1, U6136_n1, U6137_n1, U6138_n1,
         U6139_n1, U6140_n1, U6141_n1, U6142_n1, U6143_n1, U6144_n1, U6145_n1,
         U6146_n1, U6147_n1, U6148_n1, U6149_n1, U6150_n1, U6151_n1, U6152_n1,
         U6153_n1, U6154_n1, U6155_n1, U6156_n1, U6157_n1, U6158_n1, U6159_n1,
         U6160_n1, U6161_n1, U6162_n1, U6163_n1, U6164_n1, U6165_n1, U6166_n1,
         U6167_n1, U6168_n1, U6169_n1, U6170_n1, U6171_n1, U6172_n1, U6173_n1,
         U6174_n1, U6175_n1, U6176_n1, U6177_n1, U6178_n1, U6179_n1, U6180_n1,
         U6181_n1, U6182_n1, U6183_n1, U6184_n1, U6185_n1, U6186_n1, U6187_n1,
         U6188_n1, U6189_n1, U6190_n1, U6191_n1, U6192_n1, U6193_n1, U6194_n1,
         U6195_n1, U6196_n1, U6197_n1, U6198_n1, U6199_n1, U6200_n1, U6201_n1,
         U6202_n1, U6203_n1, U6204_n1, U6205_n1, U6206_n1, U6207_n1, U6208_n1,
         U6209_n1, U6210_n1, U6211_n1, U6212_n1, U6213_n1, U6214_n1, U6215_n1,
         U6216_n1, U6217_n1, U6218_n1, U6219_n1, U6220_n1, U6221_n1, U6222_n1,
         U6223_n1, U6224_n1, U6225_n1, U6226_n1, U6227_n1, U6228_n1, U6229_n1,
         U6230_n1, U6231_n1, U6232_n1, U6233_n1, U6234_n1, U6235_n1, U6236_n1,
         U6237_n1, U6238_n1, U6239_n1, U6240_n1, U6241_n1, U6242_n1, U6243_n1,
         U6244_n1, U6245_n1, U6246_n1, U6247_n1, U6248_n1, U6249_n1, U6250_n1,
         U6251_n1, U6252_n1, U6253_n1, U6254_n1, U6255_n1, U6256_n1, U6257_n1,
         U6258_n1, U6259_n1, U6260_n1, U6261_n1, U6262_n1, U6263_n1, U6264_n1,
         U6265_n1, U6266_n1, U6267_n1, U6268_n1, U6269_n1, U6270_n1, U6271_n1,
         U6272_n1, U6273_n1, U6274_n1, U6275_n1, U6276_n1, U6277_n1, U6278_n1,
         U6279_n1, U6280_n1, U6281_n1, U6282_n1, U6283_n1, U6284_n1, U6285_n1,
         U6286_n1, U6287_n1, U6288_n1, U6289_n1, U6290_n1, U6291_n1, U6292_n1,
         U6293_n1, U6294_n1, U6295_n1, U6296_n1, U6297_n1, U6298_n1, U6299_n1,
         U6300_n1, U6301_n1, U6302_n1, U6303_n1, U6304_n1, U6305_n1, U6306_n1,
         U6307_n1, U6308_n1, U6309_n1, U6310_n1, U6311_n1, U6312_n1, U6313_n1,
         U6314_n1, U6315_n1, U6316_n1, U6317_n1, U6318_n1, U6319_n1, U6320_n1,
         U6321_n1, U6322_n1, U6323_n1, U6324_n1, U6325_n1, U6326_n1, U6327_n1,
         U6328_n1, U6329_n1, U6330_n1, U6331_n1, U6332_n1, U6333_n1, U6334_n1,
         U6335_n1, U6336_n1, U6337_n1, U6338_n1, U6339_n1, U6340_n1, U6341_n1,
         U6342_n1, U6343_n1, U6344_n1, U6345_n1, U6346_n1, U6347_n1, U6348_n1,
         U6349_n1, U6350_n1, U6351_n1, U6352_n1, U6353_n1, U6354_n1, U6355_n1,
         U6356_n1, U6357_n1, U6358_n1, U6359_n1, U6360_n1, U6361_n1, U6362_n1,
         U6363_n1, U6364_n1, U6365_n1, U6366_n1, U6367_n1, U6368_n1, U6369_n1,
         U6370_n1, U6371_n1, U6372_n1, U6373_n1, U6374_n1, U6375_n1, U6376_n1,
         U6377_n1, U6378_n1, U6379_n1, U6380_n1, U6381_n1, U6382_n1, U6383_n1,
         U6384_n1, U6385_n1, U6386_n1, U6387_n1, U6388_n1, U6389_n1, U6390_n1,
         U6391_n1, U6392_n1, U6393_n1, U6394_n1, U6395_n1, U6396_n1, U6397_n1,
         U6398_n1, U6399_n1, U6400_n1, U6401_n1, U6402_n1, U6403_n1, U6404_n1,
         U6405_n1, U6406_n1, U6407_n1, U6408_n1, U6409_n1, U6410_n1, U6411_n1,
         U6412_n1, U6413_n1, U6414_n1, U6415_n1, U6416_n1, U6417_n1, U6418_n1,
         U6419_n1, U6420_n1, U6421_n1, U6422_n1, U6423_n1, U6424_n1, U6425_n1,
         U6426_n1, U6427_n1, U6428_n1, U6429_n1, U6430_n1, U6431_n1, U6432_n1,
         U6433_n1, U6434_n1, U6435_n1, U6436_n1, U6437_n1, U6438_n1, U6439_n1,
         U6440_n1, U6441_n1, U6442_n1, U6443_n1, U6444_n1, U6445_n1, U6446_n1,
         U6447_n1, U6448_n1, U6449_n1, U6450_n1, U6451_n1, U6452_n1, U6453_n1,
         U6454_n1, U6455_n1, U6456_n1, U6457_n1, U6458_n1, U6459_n1, U6460_n1,
         U6461_n1, U6462_n1, U6463_n1, U6464_n1, U6465_n1, U6466_n1, U6467_n1,
         U6468_n1, U6469_n1, U6470_n1, U6471_n1, U6472_n1, U6473_n1, U6474_n1,
         U6475_n1, U6476_n1, U6477_n1, U6478_n1, U6479_n1, U6480_n1, U6481_n1,
         U6482_n1;
  assign CRC_OUT_9_1 = test_so9;
  assign CRC_OUT_9_19 = test_so10;
  assign CRC_OUT_8_7 = test_so20;
  assign CRC_OUT_8_25 = test_so21;
  assign CRC_OUT_7_10 = test_so31;
  assign CRC_OUT_7_27 = test_so32;
  assign CRC_OUT_6_5 = test_so42;
  assign CRC_OUT_6_22 = test_so43;
  assign CRC_OUT_5_0 = test_so53;
  assign CRC_OUT_5_17 = test_so54;
  assign CRC_OUT_4_12 = test_so65;
  assign CRC_OUT_4_29 = test_so66;
  assign CRC_OUT_3_7 = test_so76;
  assign CRC_OUT_3_24 = test_so77;
  assign CRC_OUT_2_2 = test_so87;
  assign CRC_OUT_2_19 = test_so88;
  assign CRC_OUT_1_14 = test_so99;
  assign CRC_OUT_1_31 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(WX484), .SI(test_si1), .SE(n10370), .CLK(n10705), 
        .Q(WX485), .QN(n9877) );
  SDFFX1 DFF_1_Q_reg ( .D(WX486), .SI(WX485), .SE(n10365), .CLK(n10707), .Q(
        WX487), .QN(n9876) );
  SDFFX1 DFF_2_Q_reg ( .D(WX488), .SI(WX487), .SE(n10365), .CLK(n10707), .Q(
        WX489), .QN(n9874) );
  SDFFX1 DFF_3_Q_reg ( .D(WX490), .SI(WX489), .SE(n10365), .CLK(n10707), .Q(
        WX491), .QN(n9873) );
  SDFFX1 DFF_4_Q_reg ( .D(WX492), .SI(WX491), .SE(n10365), .CLK(n10707), .Q(
        WX493), .QN(n9872) );
  SDFFX1 DFF_5_Q_reg ( .D(WX494), .SI(WX493), .SE(n10366), .CLK(n10707), .Q(
        WX495), .QN(n9871) );
  SDFFX1 DFF_6_Q_reg ( .D(WX496), .SI(WX495), .SE(n10366), .CLK(n10707), .Q(
        WX497), .QN(n9870) );
  SDFFX1 DFF_7_Q_reg ( .D(WX498), .SI(WX497), .SE(n10366), .CLK(n10707), .Q(
        WX499), .QN(n9869) );
  SDFFX1 DFF_8_Q_reg ( .D(WX500), .SI(WX499), .SE(n10366), .CLK(n10707), .Q(
        WX501), .QN(n9868) );
  SDFFX1 DFF_9_Q_reg ( .D(WX502), .SI(WX501), .SE(n10366), .CLK(n10706), .Q(
        WX503), .QN(n9867) );
  SDFFX1 DFF_10_Q_reg ( .D(WX504), .SI(WX503), .SE(n10366), .CLK(n10706), .Q(
        WX505), .QN(n9866) );
  SDFFX1 DFF_11_Q_reg ( .D(WX506), .SI(WX505), .SE(n10367), .CLK(n10706), .Q(
        WX507), .QN(n9865) );
  SDFFX1 DFF_12_Q_reg ( .D(WX508), .SI(WX507), .SE(n10367), .CLK(n10706), .Q(
        WX509), .QN(n9863) );
  SDFFX1 DFF_13_Q_reg ( .D(WX510), .SI(WX509), .SE(n10367), .CLK(n10706), .Q(
        WX511), .QN(n9862) );
  SDFFX1 DFF_14_Q_reg ( .D(WX512), .SI(WX511), .SE(n10367), .CLK(n10706), .Q(
        WX513), .QN(n9861) );
  SDFFX1 DFF_15_Q_reg ( .D(WX514), .SI(WX513), .SE(n10367), .CLK(n10706), .Q(
        WX515), .QN(n9860) );
  SDFFX1 DFF_16_Q_reg ( .D(WX516), .SI(WX515), .SE(n10367), .CLK(n10706), .Q(
        WX517), .QN(n9859) );
  SDFFX1 DFF_17_Q_reg ( .D(WX518), .SI(WX517), .SE(n10368), .CLK(n10706), .Q(
        test_so1), .QN(n9858) );
  SDFFX1 DFF_18_Q_reg ( .D(WX520), .SI(test_si2), .SE(n10368), .CLK(n10706), 
        .Q(WX521), .QN(n9857) );
  SDFFX1 DFF_19_Q_reg ( .D(WX522), .SI(WX521), .SE(n10368), .CLK(n10706), .Q(
        WX523), .QN(n9856) );
  SDFFX1 DFF_20_Q_reg ( .D(WX524), .SI(WX523), .SE(n10368), .CLK(n10706), .Q(
        WX525), .QN(n9855) );
  SDFFX1 DFF_21_Q_reg ( .D(WX526), .SI(WX525), .SE(n10368), .CLK(n10705), .Q(
        WX527), .QN(n9854) );
  SDFFX1 DFF_22_Q_reg ( .D(WX528), .SI(WX527), .SE(n10368), .CLK(n10705), .Q(
        WX529), .QN(n9883) );
  SDFFX1 DFF_23_Q_reg ( .D(WX530), .SI(WX529), .SE(n10369), .CLK(n10705), .Q(
        WX531), .QN(n9882) );
  SDFFX1 DFF_24_Q_reg ( .D(WX532), .SI(WX531), .SE(n10369), .CLK(n10705), .Q(
        WX533), .QN(n9881) );
  SDFFX1 DFF_25_Q_reg ( .D(WX534), .SI(WX533), .SE(n10369), .CLK(n10705), .Q(
        WX535), .QN(n9880) );
  SDFFX1 DFF_26_Q_reg ( .D(WX536), .SI(WX535), .SE(n10369), .CLK(n10705), .Q(
        WX537), .QN(n9879) );
  SDFFX1 DFF_27_Q_reg ( .D(WX538), .SI(WX537), .SE(n10369), .CLK(n10705), .Q(
        WX539), .QN(n9878) );
  SDFFX1 DFF_28_Q_reg ( .D(WX540), .SI(WX539), .SE(n10369), .CLK(n10705), .Q(
        WX541), .QN(n9875) );
  SDFFX1 DFF_29_Q_reg ( .D(WX542), .SI(WX541), .SE(n10370), .CLK(n10705), .Q(
        WX543), .QN(n9864) );
  SDFFX1 DFF_30_Q_reg ( .D(WX544), .SI(WX543), .SE(n10370), .CLK(n10705), .Q(
        WX545), .QN(n9853) );
  SDFFX1 DFF_31_Q_reg ( .D(WX546), .SI(WX545), .SE(n10370), .CLK(n10705), .Q(
        WX547), .QN(n9852) );
  SDFFX1 DFF_32_Q_reg ( .D(WX644), .SI(WX547), .SE(n10365), .CLK(n10707), .Q(
        WX645), .QN(n3529) );
  SDFFX1 DFF_33_Q_reg ( .D(WX646), .SI(WX645), .SE(n10365), .CLK(n10707), .Q(
        WX647), .QN(n3527) );
  SDFFX1 DFF_34_Q_reg ( .D(WX648), .SI(WX647), .SE(n10364), .CLK(n10707), .Q(
        WX649), .QN(n3525) );
  SDFFX1 DFF_35_Q_reg ( .D(WX650), .SI(WX649), .SE(n10364), .CLK(n10707), .Q(
        test_so2), .QN(n9898) );
  SDFFX1 DFF_36_Q_reg ( .D(WX652), .SI(test_si3), .SE(n10364), .CLK(n10708), 
        .Q(WX653), .QN(n3521) );
  SDFFX1 DFF_37_Q_reg ( .D(WX654), .SI(WX653), .SE(n10364), .CLK(n10708), .Q(
        WX655), .QN(n3519) );
  SDFFX1 DFF_38_Q_reg ( .D(WX656), .SI(WX655), .SE(n10363), .CLK(n10708), .Q(
        WX657), .QN(n3517) );
  SDFFX1 DFF_39_Q_reg ( .D(WX658), .SI(WX657), .SE(n10363), .CLK(n10708), .Q(
        WX659), .QN(n3515) );
  SDFFX1 DFF_40_Q_reg ( .D(WX660), .SI(WX659), .SE(n10363), .CLK(n10708), .Q(
        WX661), .QN(n3513) );
  SDFFX1 DFF_41_Q_reg ( .D(WX662), .SI(WX661), .SE(n10362), .CLK(n10708), .Q(
        WX663), .QN(n3511) );
  SDFFX1 DFF_42_Q_reg ( .D(WX664), .SI(WX663), .SE(n10362), .CLK(n10709), .Q(
        WX665), .QN(n3509) );
  SDFFX1 DFF_43_Q_reg ( .D(WX666), .SI(WX665), .SE(n10362), .CLK(n10709), .Q(
        WX667), .QN(n3507) );
  SDFFX1 DFF_44_Q_reg ( .D(WX668), .SI(WX667), .SE(n10361), .CLK(n10709), .Q(
        WX669), .QN(n3505) );
  SDFFX1 DFF_45_Q_reg ( .D(WX670), .SI(WX669), .SE(n10361), .CLK(n10709), .Q(
        WX671), .QN(n3503) );
  SDFFX1 DFF_46_Q_reg ( .D(WX672), .SI(WX671), .SE(n10360), .CLK(n10709), .Q(
        WX673), .QN(n3501) );
  SDFFX1 DFF_47_Q_reg ( .D(WX674), .SI(WX673), .SE(n10360), .CLK(n10710), .Q(
        WX675), .QN(n3499) );
  SDFFX1 DFF_48_Q_reg ( .D(WX676), .SI(WX675), .SE(n10359), .CLK(n10710), .Q(
        WX677), .QN(n3497) );
  SDFFX1 DFF_49_Q_reg ( .D(WX678), .SI(WX677), .SE(n10359), .CLK(n10710), .Q(
        WX679), .QN(n3495) );
  SDFFX1 DFF_50_Q_reg ( .D(WX680), .SI(WX679), .SE(n10358), .CLK(n10711), .Q(
        WX681), .QN(n3493) );
  SDFFX1 DFF_51_Q_reg ( .D(WX682), .SI(WX681), .SE(n10357), .CLK(n10711), .Q(
        WX683), .QN(n3491) );
  SDFFX1 DFF_52_Q_reg ( .D(WX684), .SI(WX683), .SE(n10357), .CLK(n10711), .Q(
        WX685), .QN(n3489) );
  SDFFX1 DFF_53_Q_reg ( .D(WX686), .SI(WX685), .SE(n10356), .CLK(n10712), .Q(
        test_so3), .QN(n9902) );
  SDFFX1 DFF_54_Q_reg ( .D(WX688), .SI(test_si4), .SE(n10355), .CLK(n10712), 
        .Q(WX689), .QN(n3485) );
  SDFFX1 DFF_55_Q_reg ( .D(WX690), .SI(WX689), .SE(n10355), .CLK(n10712), .Q(
        WX691), .QN(n3483) );
  SDFFX1 DFF_56_Q_reg ( .D(WX692), .SI(WX691), .SE(n10354), .CLK(n10713), .Q(
        WX693), .QN(n3481) );
  SDFFX1 DFF_57_Q_reg ( .D(WX694), .SI(WX693), .SE(n10353), .CLK(n10713), .Q(
        WX695), .QN(n3479) );
  SDFFX1 DFF_58_Q_reg ( .D(WX696), .SI(WX695), .SE(n10353), .CLK(n10713), .Q(
        WX697), .QN(n3477) );
  SDFFX1 DFF_59_Q_reg ( .D(WX698), .SI(WX697), .SE(n10352), .CLK(n10714), .Q(
        WX699), .QN(n3475) );
  SDFFX1 DFF_60_Q_reg ( .D(WX700), .SI(WX699), .SE(n10351), .CLK(n10714), .Q(
        WX701), .QN(n3473) );
  SDFFX1 DFF_61_Q_reg ( .D(WX702), .SI(WX701), .SE(n10351), .CLK(n10714), .Q(
        WX703), .QN(n3471) );
  SDFFX1 DFF_62_Q_reg ( .D(WX704), .SI(WX703), .SE(n10350), .CLK(n10715), .Q(
        WX705), .QN(n3469) );
  SDFFX1 DFF_63_Q_reg ( .D(WX706), .SI(WX705), .SE(n10349), .CLK(n10715), .Q(
        WX707), .QN(n3467) );
  SDFFX1 DFF_64_Q_reg ( .D(WX708), .SI(WX707), .SE(n10349), .CLK(n10715), .Q(
        WX709), .QN(n9827) );
  SDFFX1 DFF_65_Q_reg ( .D(WX710), .SI(WX709), .SE(n10348), .CLK(n10716), .Q(
        WX711), .QN(n9753) );
  SDFFX1 DFF_66_Q_reg ( .D(WX712), .SI(WX711), .SE(n10348), .CLK(n10716), .Q(
        WX713), .QN(n9764) );
  SDFFX1 DFF_67_Q_reg ( .D(WX714), .SI(WX713), .SE(n10364), .CLK(n10708), .Q(
        WX715), .QN(n9773) );
  SDFFX1 DFF_68_Q_reg ( .D(WX716), .SI(WX715), .SE(n10364), .CLK(n10708), .Q(
        WX717), .QN(n9779) );
  SDFFX1 DFF_69_Q_reg ( .D(WX718), .SI(WX717), .SE(n10363), .CLK(n10708), .Q(
        WX719), .QN(n9782) );
  SDFFX1 DFF_70_Q_reg ( .D(WX720), .SI(WX719), .SE(n10363), .CLK(n10708), .Q(
        WX721), .QN(n9791) );
  SDFFX1 DFF_71_Q_reg ( .D(WX722), .SI(WX721), .SE(n10363), .CLK(n10708), .Q(
        test_so4), .QN(n9899) );
  SDFFX1 DFF_72_Q_reg ( .D(WX724), .SI(test_si5), .SE(n10362), .CLK(n10708), 
        .Q(WX725), .QN(n9802) );
  SDFFX1 DFF_73_Q_reg ( .D(WX726), .SI(WX725), .SE(n10362), .CLK(n10709), .Q(
        WX727), .QN(n9814) );
  SDFFX1 DFF_74_Q_reg ( .D(WX728), .SI(WX727), .SE(n10362), .CLK(n10709), .Q(
        WX729), .QN(n9820) );
  SDFFX1 DFF_75_Q_reg ( .D(WX730), .SI(WX729), .SE(n10361), .CLK(n10709), .Q(
        WX731), .QN(n9826) );
  SDFFX1 DFF_76_Q_reg ( .D(WX732), .SI(WX731), .SE(n10361), .CLK(n10709), .Q(
        WX733), .QN(n9761) );
  SDFFX1 DFF_77_Q_reg ( .D(WX734), .SI(WX733), .SE(n10361), .CLK(n10709), .Q(
        WX735), .QN(n9776) );
  SDFFX1 DFF_78_Q_reg ( .D(WX736), .SI(WX735), .SE(n10360), .CLK(n10710), .Q(
        WX737), .QN(n9788) );
  SDFFX1 DFF_79_Q_reg ( .D(WX738), .SI(WX737), .SE(n10360), .CLK(n10710), .Q(
        WX739), .QN(n9803) );
  SDFFX1 DFF_80_Q_reg ( .D(WX740), .SI(WX739), .SE(n10359), .CLK(n10710), .Q(
        WX741), .QN(n9817) );
  SDFFX1 DFF_81_Q_reg ( .D(WX742), .SI(WX741), .SE(n10358), .CLK(n10710), .Q(
        WX743), .QN(n9832) );
  SDFFX1 DFF_82_Q_reg ( .D(WX744), .SI(WX743), .SE(n10358), .CLK(n10711), .Q(
        WX745), .QN(n9767) );
  SDFFX1 DFF_83_Q_reg ( .D(WX746), .SI(WX745), .SE(n10357), .CLK(n10711), .Q(
        WX747), .QN(n9794) );
  SDFFX1 DFF_84_Q_reg ( .D(WX748), .SI(WX747), .SE(n10356), .CLK(n10711), .Q(
        WX749), .QN(n9840) );
  SDFFX1 DFF_85_Q_reg ( .D(WX750), .SI(WX749), .SE(n10356), .CLK(n10712), .Q(
        WX751), .QN(n9785) );
  SDFFX1 DFF_86_Q_reg ( .D(WX752), .SI(WX751), .SE(n10355), .CLK(n10712), .Q(
        WX753), .QN(n9795) );
  SDFFX1 DFF_87_Q_reg ( .D(WX754), .SI(WX753), .SE(n10354), .CLK(n10712), .Q(
        WX755), .QN(n9807) );
  SDFFX1 DFF_88_Q_reg ( .D(WX756), .SI(WX755), .SE(n10354), .CLK(n10713), .Q(
        WX757), .QN(n9835) );
  SDFFX1 DFF_89_Q_reg ( .D(WX758), .SI(WX757), .SE(n10353), .CLK(n10713), .Q(
        test_so5), .QN(n9897) );
  SDFFX1 DFF_90_Q_reg ( .D(WX760), .SI(test_si6), .SE(n10352), .CLK(n10713), 
        .Q(WX761), .QN(n9810) );
  SDFFX1 DFF_91_Q_reg ( .D(WX762), .SI(WX761), .SE(n10352), .CLK(n10714), .Q(
        WX763), .QN(n9813) );
  SDFFX1 DFF_92_Q_reg ( .D(WX764), .SI(WX763), .SE(n10351), .CLK(n10714), .Q(
        WX765), .QN(n9758) );
  SDFFX1 DFF_93_Q_reg ( .D(WX766), .SI(WX765), .SE(n10350), .CLK(n10714), .Q(
        WX767), .QN(n9833) );
  SDFFX1 DFF_94_Q_reg ( .D(WX768), .SI(WX767), .SE(n10350), .CLK(n10715), .Q(
        WX769) );
  SDFFX1 DFF_95_Q_reg ( .D(WX770), .SI(WX769), .SE(n10349), .CLK(n10715), .Q(
        WX771), .QN(n9841) );
  SDFFX1 DFF_96_Q_reg ( .D(WX772), .SI(WX771), .SE(n10348), .CLK(n10715), .Q(
        WX773), .QN(n9828) );
  SDFFX1 DFF_97_Q_reg ( .D(WX774), .SI(WX773), .SE(n10348), .CLK(n10716), .Q(
        WX775), .QN(n9754) );
  SDFFX1 DFF_98_Q_reg ( .D(WX776), .SI(WX775), .SE(n10347), .CLK(n10716), .Q(
        WX777), .QN(n9762) );
  SDFFX1 DFF_99_Q_reg ( .D(WX778), .SI(WX777), .SE(n10347), .CLK(n10716), .Q(
        WX779), .QN(n9771) );
  SDFFX1 DFF_100_Q_reg ( .D(WX780), .SI(WX779), .SE(n10347), .CLK(n10716), .Q(
        WX781), .QN(n9777) );
  SDFFX1 DFF_101_Q_reg ( .D(WX782), .SI(WX781), .SE(n10346), .CLK(n10716), .Q(
        WX783), .QN(n9780) );
  SDFFX1 DFF_102_Q_reg ( .D(WX784), .SI(WX783), .SE(n10346), .CLK(n10717), .Q(
        WX785), .QN(n9789) );
  SDFFX1 DFF_103_Q_reg ( .D(WX786), .SI(WX785), .SE(n10346), .CLK(n10717), .Q(
        WX787), .QN(n9798) );
  SDFFX1 DFF_104_Q_reg ( .D(WX788), .SI(WX787), .SE(n10345), .CLK(n10717), .Q(
        WX789), .QN(n9800) );
  SDFFX1 DFF_105_Q_reg ( .D(WX790), .SI(WX789), .SE(n10345), .CLK(n10717), .Q(
        WX791), .QN(n9815) );
  SDFFX1 DFF_106_Q_reg ( .D(WX792), .SI(WX791), .SE(n10345), .CLK(n10717), .Q(
        WX793), .QN(n9821) );
  SDFFX1 DFF_107_Q_reg ( .D(WX794), .SI(WX793), .SE(n10344), .CLK(n10717), .Q(
        test_so6), .QN(n9900) );
  SDFFX1 DFF_108_Q_reg ( .D(WX796), .SI(test_si7), .SE(n10361), .CLK(n10709), 
        .Q(WX797), .QN(n9759) );
  SDFFX1 DFF_109_Q_reg ( .D(WX798), .SI(WX797), .SE(n10360), .CLK(n10709), .Q(
        WX799), .QN(n9774) );
  SDFFX1 DFF_110_Q_reg ( .D(WX800), .SI(WX799), .SE(n10360), .CLK(n10710), .Q(
        WX801), .QN(n9786) );
  SDFFX1 DFF_111_Q_reg ( .D(WX802), .SI(WX801), .SE(n10359), .CLK(n10710), .Q(
        WX803), .QN(n9804) );
  SDFFX1 DFF_112_Q_reg ( .D(WX804), .SI(WX803), .SE(n10359), .CLK(n10710), .Q(
        WX805), .QN(n9818) );
  SDFFX1 DFF_113_Q_reg ( .D(WX806), .SI(WX805), .SE(n10358), .CLK(n10710), .Q(
        WX807), .QN(n9830) );
  SDFFX1 DFF_114_Q_reg ( .D(WX808), .SI(WX807), .SE(n10358), .CLK(n10711), .Q(
        WX809), .QN(n9765) );
  SDFFX1 DFF_115_Q_reg ( .D(WX810), .SI(WX809), .SE(n10357), .CLK(n10711), .Q(
        WX811), .QN(n9792) );
  SDFFX1 DFF_116_Q_reg ( .D(WX812), .SI(WX811), .SE(n10356), .CLK(n10711), .Q(
        WX813), .QN(n9838) );
  SDFFX1 DFF_117_Q_reg ( .D(WX814), .SI(WX813), .SE(n10356), .CLK(n10712), .Q(
        WX815), .QN(n9783) );
  SDFFX1 DFF_118_Q_reg ( .D(WX816), .SI(WX815), .SE(n10355), .CLK(n10712), .Q(
        WX817), .QN(n9796) );
  SDFFX1 DFF_119_Q_reg ( .D(WX818), .SI(WX817), .SE(n10354), .CLK(n10712), .Q(
        WX819), .QN(n9805) );
  SDFFX1 DFF_120_Q_reg ( .D(WX820), .SI(WX819), .SE(n10354), .CLK(n10713), .Q(
        WX821), .QN(n9836) );
  SDFFX1 DFF_121_Q_reg ( .D(WX822), .SI(WX821), .SE(n10353), .CLK(n10713), .Q(
        WX823), .QN(n9823) );
  SDFFX1 DFF_122_Q_reg ( .D(WX824), .SI(WX823), .SE(n10352), .CLK(n10713), .Q(
        WX825), .QN(n9808) );
  SDFFX1 DFF_123_Q_reg ( .D(WX826), .SI(WX825), .SE(n10352), .CLK(n10714), .Q(
        WX827), .QN(n9811) );
  SDFFX1 DFF_124_Q_reg ( .D(WX828), .SI(WX827), .SE(n10351), .CLK(n10714), .Q(
        WX829), .QN(n9756) );
  SDFFX1 DFF_125_Q_reg ( .D(WX830), .SI(WX829), .SE(n10350), .CLK(n10714), .Q(
        test_so7), .QN(n9901) );
  SDFFX1 DFF_126_Q_reg ( .D(WX832), .SI(test_si8), .SE(n10350), .CLK(n10715), 
        .Q(WX833), .QN(n9770) );
  SDFFX1 DFF_127_Q_reg ( .D(WX834), .SI(WX833), .SE(n10349), .CLK(n10715), .Q(
        WX835), .QN(n9842) );
  SDFFX1 DFF_128_Q_reg ( .D(WX836), .SI(WX835), .SE(n10348), .CLK(n10715), .Q(
        WX837), .QN(n9829) );
  SDFFX1 DFF_129_Q_reg ( .D(WX838), .SI(WX837), .SE(n10348), .CLK(n10716), .Q(
        WX839), .QN(n9755) );
  SDFFX1 DFF_130_Q_reg ( .D(WX840), .SI(WX839), .SE(n10347), .CLK(n10716), .Q(
        WX841), .QN(n9763) );
  SDFFX1 DFF_131_Q_reg ( .D(WX842), .SI(WX841), .SE(n10347), .CLK(n10716), .Q(
        WX843), .QN(n9772) );
  SDFFX1 DFF_132_Q_reg ( .D(WX844), .SI(WX843), .SE(n10347), .CLK(n10716), .Q(
        WX845), .QN(n9778) );
  SDFFX1 DFF_133_Q_reg ( .D(WX846), .SI(WX845), .SE(n10346), .CLK(n10716), .Q(
        WX847), .QN(n9781) );
  SDFFX1 DFF_134_Q_reg ( .D(WX848), .SI(WX847), .SE(n10346), .CLK(n10717), .Q(
        WX849), .QN(n9790) );
  SDFFX1 DFF_135_Q_reg ( .D(WX850), .SI(WX849), .SE(n10346), .CLK(n10717), .Q(
        WX851), .QN(n9799) );
  SDFFX1 DFF_136_Q_reg ( .D(WX852), .SI(WX851), .SE(n10345), .CLK(n10717), .Q(
        WX853), .QN(n9801) );
  SDFFX1 DFF_137_Q_reg ( .D(WX854), .SI(WX853), .SE(n10345), .CLK(n10717), .Q(
        WX855), .QN(n9816) );
  SDFFX1 DFF_138_Q_reg ( .D(WX856), .SI(WX855), .SE(n10345), .CLK(n10717), .Q(
        WX857), .QN(n9822) );
  SDFFX1 DFF_139_Q_reg ( .D(WX858), .SI(WX857), .SE(n10344), .CLK(n10717), .Q(
        WX859), .QN(n9825) );
  SDFFX1 DFF_140_Q_reg ( .D(WX860), .SI(WX859), .SE(n10344), .CLK(n10718), .Q(
        WX861), .QN(n9760) );
  SDFFX1 DFF_141_Q_reg ( .D(WX862), .SI(WX861), .SE(n10344), .CLK(n10718), .Q(
        WX863), .QN(n9775) );
  SDFFX1 DFF_142_Q_reg ( .D(WX864), .SI(WX863), .SE(n10344), .CLK(n10718), .Q(
        WX865), .QN(n9787) );
  SDFFX1 DFF_143_Q_reg ( .D(WX866), .SI(WX865), .SE(n10344), .CLK(n10718), .Q(
        test_so8), .QN(n9885) );
  SDFFX1 DFF_144_Q_reg ( .D(WX868), .SI(test_si9), .SE(n10359), .CLK(n10710), 
        .Q(WX869), .QN(n9819) );
  SDFFX1 DFF_145_Q_reg ( .D(WX870), .SI(WX869), .SE(n10358), .CLK(n10711), .Q(
        WX871), .QN(n9831) );
  SDFFX1 DFF_146_Q_reg ( .D(WX872), .SI(WX871), .SE(n10357), .CLK(n10711), .Q(
        WX873), .QN(n9766) );
  SDFFX1 DFF_147_Q_reg ( .D(WX874), .SI(WX873), .SE(n10357), .CLK(n10711), .Q(
        WX875), .QN(n9793) );
  SDFFX1 DFF_148_Q_reg ( .D(WX876), .SI(WX875), .SE(n10356), .CLK(n10712), .Q(
        WX877), .QN(n9839) );
  SDFFX1 DFF_149_Q_reg ( .D(WX878), .SI(WX877), .SE(n10355), .CLK(n10712), .Q(
        WX879), .QN(n9784) );
  SDFFX1 DFF_150_Q_reg ( .D(WX880), .SI(WX879), .SE(n10355), .CLK(n10712), .Q(
        WX881), .QN(n9797) );
  SDFFX1 DFF_151_Q_reg ( .D(WX882), .SI(WX881), .SE(n10354), .CLK(n10713), .Q(
        WX883), .QN(n9806) );
  SDFFX1 DFF_152_Q_reg ( .D(WX884), .SI(WX883), .SE(n10353), .CLK(n10713), .Q(
        WX885), .QN(n9837) );
  SDFFX1 DFF_153_Q_reg ( .D(WX886), .SI(WX885), .SE(n10353), .CLK(n10713), .Q(
        WX887), .QN(n9824) );
  SDFFX1 DFF_154_Q_reg ( .D(WX888), .SI(WX887), .SE(n10352), .CLK(n10714), .Q(
        WX889), .QN(n9809) );
  SDFFX1 DFF_155_Q_reg ( .D(WX890), .SI(WX889), .SE(n10351), .CLK(n10714), .Q(
        WX891), .QN(n9812) );
  SDFFX1 DFF_156_Q_reg ( .D(WX892), .SI(WX891), .SE(n10351), .CLK(n10714), .Q(
        WX893), .QN(n9757) );
  SDFFX1 DFF_157_Q_reg ( .D(WX894), .SI(WX893), .SE(n10350), .CLK(n10715), .Q(
        WX895), .QN(n9834) );
  SDFFX1 DFF_158_Q_reg ( .D(WX896), .SI(WX895), .SE(n10349), .CLK(n10715), .Q(
        WX897), .QN(n9768) );
  SDFFX1 DFF_159_Q_reg ( .D(WX898), .SI(WX897), .SE(n10349), .CLK(n10715), .Q(
        WX899), .QN(n9843) );
  SDFFX1 DFF_160_Q_reg ( .D(WX1264), .SI(WX899), .SE(n10087), .CLK(n10847), 
        .Q(CRC_OUT_9_0) );
  SDFFX1 DFF_161_Q_reg ( .D(WX1266), .SI(CRC_OUT_9_0), .SE(n10087), .CLK(
        n10847), .Q(test_so9), .QN(n9949) );
  SDFFX1 DFF_162_Q_reg ( .D(WX1268), .SI(test_si10), .SE(n10086), .CLK(n10847), 
        .Q(CRC_OUT_9_2), .QN(DFF_162_n1) );
  SDFFX1 DFF_163_Q_reg ( .D(WX1270), .SI(CRC_OUT_9_2), .SE(n10086), .CLK(
        n10847), .Q(CRC_OUT_9_3), .QN(DFF_163_n1) );
  SDFFX1 DFF_164_Q_reg ( .D(WX1272), .SI(CRC_OUT_9_3), .SE(n10086), .CLK(
        n10847), .Q(CRC_OUT_9_4), .QN(DFF_164_n1) );
  SDFFX1 DFF_165_Q_reg ( .D(WX1274), .SI(CRC_OUT_9_4), .SE(n10086), .CLK(
        n10847), .Q(CRC_OUT_9_5), .QN(DFF_165_n1) );
  SDFFX1 DFF_166_Q_reg ( .D(WX1276), .SI(CRC_OUT_9_5), .SE(n10086), .CLK(
        n10847), .Q(CRC_OUT_9_6), .QN(DFF_166_n1) );
  SDFFX1 DFF_167_Q_reg ( .D(WX1278), .SI(CRC_OUT_9_6), .SE(n10086), .CLK(
        n10847), .Q(CRC_OUT_9_7), .QN(DFF_167_n1) );
  SDFFX1 DFF_168_Q_reg ( .D(WX1280), .SI(CRC_OUT_9_7), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_8), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(WX1282), .SI(CRC_OUT_9_8), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_9), .QN(DFF_169_n1) );
  SDFFX1 DFF_170_Q_reg ( .D(WX1284), .SI(CRC_OUT_9_9), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_10), .QN(DFF_170_n1) );
  SDFFX1 DFF_171_Q_reg ( .D(WX1286), .SI(CRC_OUT_9_10), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_11), .QN(DFF_171_n1) );
  SDFFX1 DFF_172_Q_reg ( .D(WX1288), .SI(CRC_OUT_9_11), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_12), .QN(DFF_172_n1) );
  SDFFX1 DFF_173_Q_reg ( .D(WX1290), .SI(CRC_OUT_9_12), .SE(n10085), .CLK(
        n10848), .Q(CRC_OUT_9_13), .QN(DFF_173_n1) );
  SDFFX1 DFF_174_Q_reg ( .D(WX1292), .SI(CRC_OUT_9_13), .SE(n10084), .CLK(
        n10848), .Q(CRC_OUT_9_14), .QN(DFF_174_n1) );
  SDFFX1 DFF_175_Q_reg ( .D(WX1294), .SI(CRC_OUT_9_14), .SE(n10084), .CLK(
        n10848), .Q(CRC_OUT_9_15), .QN(DFF_175_n1) );
  SDFFX1 DFF_176_Q_reg ( .D(WX1296), .SI(CRC_OUT_9_15), .SE(n10084), .CLK(
        n10848), .Q(CRC_OUT_9_16), .QN(DFF_176_n1) );
  SDFFX1 DFF_177_Q_reg ( .D(WX1298), .SI(CRC_OUT_9_16), .SE(n10084), .CLK(
        n10848), .Q(CRC_OUT_9_17), .QN(DFF_177_n1) );
  SDFFX1 DFF_178_Q_reg ( .D(WX1300), .SI(CRC_OUT_9_17), .SE(n10084), .CLK(
        n10848), .Q(CRC_OUT_9_18), .QN(DFF_178_n1) );
  SDFFX1 DFF_179_Q_reg ( .D(WX1302), .SI(CRC_OUT_9_18), .SE(n10084), .CLK(
        n10848), .Q(test_so10), .QN(n9948) );
  SDFFX1 DFF_180_Q_reg ( .D(WX1304), .SI(test_si11), .SE(n10343), .CLK(n10718), 
        .Q(CRC_OUT_9_20), .QN(DFF_180_n1) );
  SDFFX1 DFF_181_Q_reg ( .D(WX1306), .SI(CRC_OUT_9_20), .SE(n10343), .CLK(
        n10718), .Q(CRC_OUT_9_21), .QN(DFF_181_n1) );
  SDFFX1 DFF_182_Q_reg ( .D(WX1308), .SI(CRC_OUT_9_21), .SE(n10343), .CLK(
        n10718), .Q(CRC_OUT_9_22), .QN(DFF_182_n1) );
  SDFFX1 DFF_183_Q_reg ( .D(WX1310), .SI(CRC_OUT_9_22), .SE(n10343), .CLK(
        n10718), .Q(CRC_OUT_9_23), .QN(DFF_183_n1) );
  SDFFX1 DFF_184_Q_reg ( .D(WX1312), .SI(CRC_OUT_9_23), .SE(n10343), .CLK(
        n10718), .Q(CRC_OUT_9_24), .QN(DFF_184_n1) );
  SDFFX1 DFF_185_Q_reg ( .D(WX1314), .SI(CRC_OUT_9_24), .SE(n10343), .CLK(
        n10718), .Q(CRC_OUT_9_25), .QN(DFF_185_n1) );
  SDFFX1 DFF_186_Q_reg ( .D(WX1316), .SI(CRC_OUT_9_25), .SE(n10342), .CLK(
        n10718), .Q(CRC_OUT_9_26), .QN(DFF_186_n1) );
  SDFFX1 DFF_187_Q_reg ( .D(WX1318), .SI(CRC_OUT_9_26), .SE(n10342), .CLK(
        n10718), .Q(CRC_OUT_9_27), .QN(DFF_187_n1) );
  SDFFX1 DFF_188_Q_reg ( .D(WX1320), .SI(CRC_OUT_9_27), .SE(n10342), .CLK(
        n10719), .Q(CRC_OUT_9_28), .QN(DFF_188_n1) );
  SDFFX1 DFF_189_Q_reg ( .D(WX1322), .SI(CRC_OUT_9_28), .SE(n10342), .CLK(
        n10719), .Q(CRC_OUT_9_29), .QN(DFF_189_n1) );
  SDFFX1 DFF_190_Q_reg ( .D(WX1324), .SI(CRC_OUT_9_29), .SE(n10342), .CLK(
        n10719), .Q(CRC_OUT_9_30), .QN(DFF_190_n1) );
  SDFFX1 DFF_191_Q_reg ( .D(WX1326), .SI(CRC_OUT_9_30), .SE(n10342), .CLK(
        n10719), .Q(CRC_OUT_9_31), .QN(DFF_191_n1) );
  SDFFX1 DFF_192_Q_reg ( .D(n250), .SI(CRC_OUT_9_31), .SE(n10341), .CLK(n10719), .Q(WX1778), .QN(n9844) );
  SDFFX1 DFF_193_Q_reg ( .D(n251), .SI(WX1778), .SE(n10336), .CLK(n10721), .Q(
        n8702), .QN(n4033) );
  SDFFX1 DFF_194_Q_reg ( .D(n252), .SI(n8702), .SE(n10336), .CLK(n10721), .Q(
        n8701), .QN(n4032) );
  SDFFX1 DFF_195_Q_reg ( .D(n253), .SI(n8701), .SE(n10337), .CLK(n10721), .Q(
        n8700), .QN(n4031) );
  SDFFX1 DFF_196_Q_reg ( .D(n254), .SI(n8700), .SE(n10337), .CLK(n10721), .Q(
        n8699), .QN(n4030) );
  SDFFX1 DFF_197_Q_reg ( .D(n255), .SI(n8699), .SE(n10337), .CLK(n10721), .Q(
        test_so11), .QN(n4029) );
  SDFFX1 DFF_198_Q_reg ( .D(n256), .SI(test_si12), .SE(n10337), .CLK(n10721), 
        .Q(n8696), .QN(n4028) );
  SDFFX1 DFF_199_Q_reg ( .D(n257), .SI(n8696), .SE(n10337), .CLK(n10721), .Q(
        n8695), .QN(n4027) );
  SDFFX1 DFF_200_Q_reg ( .D(n258), .SI(n8695), .SE(n10337), .CLK(n10721), .Q(
        n8694), .QN(n4026) );
  SDFFX1 DFF_201_Q_reg ( .D(n259), .SI(n8694), .SE(n10338), .CLK(n10721), .Q(
        n8693), .QN(n4025) );
  SDFFX1 DFF_202_Q_reg ( .D(n260), .SI(n8693), .SE(n10338), .CLK(n10721), .Q(
        n8692), .QN(n4024) );
  SDFFX1 DFF_203_Q_reg ( .D(n261), .SI(n8692), .SE(n10338), .CLK(n10721), .Q(
        n8691), .QN(n4023) );
  SDFFX1 DFF_204_Q_reg ( .D(n262), .SI(n8691), .SE(n10338), .CLK(n10721), .Q(
        n8690), .QN(n4022) );
  SDFFX1 DFF_205_Q_reg ( .D(n263), .SI(n8690), .SE(n10338), .CLK(n10720), .Q(
        n8689), .QN(n4021) );
  SDFFX1 DFF_206_Q_reg ( .D(n264), .SI(n8689), .SE(n10338), .CLK(n10720), .Q(
        n8688), .QN(n4020) );
  SDFFX1 DFF_207_Q_reg ( .D(n265), .SI(n8688), .SE(n10339), .CLK(n10720), .Q(
        n8687), .QN(n4019) );
  SDFFX1 DFF_208_Q_reg ( .D(n266), .SI(n8687), .SE(n10339), .CLK(n10720), .Q(
        n8686), .QN(n4018) );
  SDFFX1 DFF_209_Q_reg ( .D(n267), .SI(n8686), .SE(n10339), .CLK(n10720), .Q(
        n8685), .QN(n4017) );
  SDFFX1 DFF_210_Q_reg ( .D(n268), .SI(n8685), .SE(n10339), .CLK(n10720), .Q(
        n8684), .QN(n4016) );
  SDFFX1 DFF_211_Q_reg ( .D(n269), .SI(n8684), .SE(n10339), .CLK(n10720), .Q(
        n8683), .QN(n4015) );
  SDFFX1 DFF_212_Q_reg ( .D(n270), .SI(n8683), .SE(n10339), .CLK(n10720), .Q(
        n8682), .QN(n4014) );
  SDFFX1 DFF_213_Q_reg ( .D(n271), .SI(n8682), .SE(n10340), .CLK(n10720), .Q(
        n8681), .QN(n4013) );
  SDFFX1 DFF_214_Q_reg ( .D(n272), .SI(n8681), .SE(n10340), .CLK(n10720), .Q(
        n8680), .QN(n4012) );
  SDFFX1 DFF_215_Q_reg ( .D(n273), .SI(n8680), .SE(n10340), .CLK(n10720), .Q(
        test_so12), .QN(n4011) );
  SDFFX1 DFF_216_Q_reg ( .D(n274), .SI(test_si13), .SE(n10340), .CLK(n10720), 
        .Q(n8677), .QN(n4010) );
  SDFFX1 DFF_217_Q_reg ( .D(n275), .SI(n8677), .SE(n10340), .CLK(n10719), .Q(
        n8676), .QN(n4009) );
  SDFFX1 DFF_218_Q_reg ( .D(n276), .SI(n8676), .SE(n10340), .CLK(n10719), .Q(
        n8675), .QN(n4008) );
  SDFFX1 DFF_219_Q_reg ( .D(n277), .SI(n8675), .SE(n10341), .CLK(n10719), .Q(
        n8674), .QN(n4007) );
  SDFFX1 DFF_220_Q_reg ( .D(n278), .SI(n8674), .SE(n10341), .CLK(n10719), .Q(
        n8673), .QN(n4006) );
  SDFFX1 DFF_221_Q_reg ( .D(n279), .SI(n8673), .SE(n10341), .CLK(n10719), .Q(
        n8672), .QN(n4005) );
  SDFFX1 DFF_222_Q_reg ( .D(n280), .SI(n8672), .SE(n10341), .CLK(n10719), .Q(
        n8671), .QN(n4004) );
  SDFFX1 DFF_223_Q_reg ( .D(WX1839), .SI(n8671), .SE(n10341), .CLK(n10719), 
        .Q(n8670), .QN(n4003) );
  SDFFX1 DFF_224_Q_reg ( .D(WX1937), .SI(n8670), .SE(n10332), .CLK(n10724), 
        .Q(n8669), .QN(n17986) );
  SDFFX1 DFF_225_Q_reg ( .D(WX1939), .SI(n8669), .SE(n10332), .CLK(n10724), 
        .Q(n8668), .QN(n17983) );
  SDFFX1 DFF_226_Q_reg ( .D(WX1941), .SI(n8668), .SE(n10331), .CLK(n10724), 
        .Q(n8667), .QN(n17981) );
  SDFFX1 DFF_227_Q_reg ( .D(WX1943), .SI(n8667), .SE(n10331), .CLK(n10724), 
        .Q(n8666), .QN(n17979) );
  SDFFX1 DFF_228_Q_reg ( .D(WX1945), .SI(n8666), .SE(n10330), .CLK(n10725), 
        .Q(n8665), .QN(n17977) );
  SDFFX1 DFF_229_Q_reg ( .D(WX1947), .SI(n8665), .SE(n10329), .CLK(n10725), 
        .Q(n8664), .QN(n17975) );
  SDFFX1 DFF_230_Q_reg ( .D(WX1949), .SI(n8664), .SE(n10328), .CLK(n10726), 
        .Q(n8663), .QN(n17973) );
  SDFFX1 DFF_231_Q_reg ( .D(WX1951), .SI(n8663), .SE(n10328), .CLK(n10726), 
        .Q(n8662), .QN(n17971) );
  SDFFX1 DFF_232_Q_reg ( .D(WX1953), .SI(n8662), .SE(n10327), .CLK(n10726), 
        .Q(n8661), .QN(n17969) );
  SDFFX1 DFF_233_Q_reg ( .D(WX1955), .SI(n8661), .SE(n10327), .CLK(n10726), 
        .Q(test_so13), .QN(n9895) );
  SDFFX1 DFF_234_Q_reg ( .D(WX1957), .SI(test_si14), .SE(n10326), .CLK(n10727), 
        .Q(n8658), .QN(n17966) );
  SDFFX1 DFF_235_Q_reg ( .D(WX1959), .SI(n8658), .SE(n10325), .CLK(n10727), 
        .Q(n8657), .QN(n17964) );
  SDFFX1 DFF_236_Q_reg ( .D(WX1961), .SI(n8657), .SE(n10324), .CLK(n10728), 
        .Q(n8656), .QN(n17962) );
  SDFFX1 DFF_237_Q_reg ( .D(WX1963), .SI(n8656), .SE(n10324), .CLK(n10728), 
        .Q(n8655), .QN(n17960) );
  SDFFX1 DFF_238_Q_reg ( .D(WX1965), .SI(n8655), .SE(n10323), .CLK(n10728), 
        .Q(n8654), .QN(n17958) );
  SDFFX1 DFF_239_Q_reg ( .D(WX1967), .SI(n8654), .SE(n10322), .CLK(n10729), 
        .Q(n8653), .QN(n17957) );
  SDFFX1 DFF_240_Q_reg ( .D(WX1969), .SI(n8653), .SE(n10322), .CLK(n10729), 
        .Q(WX1970), .QN(n9510) );
  SDFFX1 DFF_241_Q_reg ( .D(WX1971), .SI(WX1970), .SE(n10321), .CLK(n10729), 
        .Q(WX1972) );
  SDFFX1 DFF_242_Q_reg ( .D(WX1973), .SI(WX1972), .SE(n10321), .CLK(n10729), 
        .Q(WX1974), .QN(n9507) );
  SDFFX1 DFF_243_Q_reg ( .D(WX1975), .SI(WX1974), .SE(n10320), .CLK(n10730), 
        .Q(WX1976), .QN(n9505) );
  SDFFX1 DFF_244_Q_reg ( .D(WX1977), .SI(WX1976), .SE(n10335), .CLK(n10722), 
        .Q(WX1978), .QN(n9503) );
  SDFFX1 DFF_245_Q_reg ( .D(WX1979), .SI(WX1978), .SE(n10335), .CLK(n10722), 
        .Q(WX1980) );
  SDFFX1 DFF_246_Q_reg ( .D(WX1981), .SI(WX1980), .SE(n10335), .CLK(n10722), 
        .Q(WX1982), .QN(n9499) );
  SDFFX1 DFF_247_Q_reg ( .D(WX1983), .SI(WX1982), .SE(n10334), .CLK(n10722), 
        .Q(WX1984), .QN(n9497) );
  SDFFX1 DFF_248_Q_reg ( .D(WX1985), .SI(WX1984), .SE(n10334), .CLK(n10723), 
        .Q(WX1986), .QN(n9495) );
  SDFFX1 DFF_249_Q_reg ( .D(WX1987), .SI(WX1986), .SE(n10334), .CLK(n10723), 
        .Q(WX1988), .QN(n9493) );
  SDFFX1 DFF_250_Q_reg ( .D(WX1989), .SI(WX1988), .SE(n10334), .CLK(n10723), 
        .Q(WX1990), .QN(n9491) );
  SDFFX1 DFF_251_Q_reg ( .D(WX1991), .SI(WX1990), .SE(n10334), .CLK(n10723), 
        .Q(test_so14), .QN(n9930) );
  SDFFX1 DFF_252_Q_reg ( .D(WX1993), .SI(test_si15), .SE(n10333), .CLK(n10723), 
        .Q(WX1994), .QN(n9488) );
  SDFFX1 DFF_253_Q_reg ( .D(WX1995), .SI(WX1994), .SE(n10333), .CLK(n10723), 
        .Q(WX1996), .QN(n9486) );
  SDFFX1 DFF_254_Q_reg ( .D(WX1997), .SI(WX1996), .SE(n10333), .CLK(n10723), 
        .Q(WX1998), .QN(n9484) );
  SDFFX1 DFF_255_Q_reg ( .D(WX1999), .SI(WX1998), .SE(n10332), .CLK(n10723), 
        .Q(WX2000), .QN(n9482) );
  SDFFX1 DFF_256_Q_reg ( .D(WX2001), .SI(WX2000), .SE(n10332), .CLK(n10724), 
        .Q(WX2002), .QN(n9042) );
  SDFFX1 DFF_257_Q_reg ( .D(WX2003), .SI(WX2002), .SE(n10331), .CLK(n10724), 
        .Q(WX2004), .QN(n9268) );
  SDFFX1 DFF_258_Q_reg ( .D(WX2005), .SI(WX2004), .SE(n10331), .CLK(n10724), 
        .Q(WX2006), .QN(n9266) );
  SDFFX1 DFF_259_Q_reg ( .D(WX2007), .SI(WX2006), .SE(n10330), .CLK(n10724), 
        .Q(WX2008), .QN(n9264) );
  SDFFX1 DFF_260_Q_reg ( .D(WX2009), .SI(WX2008), .SE(n10330), .CLK(n10725), 
        .Q(WX2010), .QN(n9262) );
  SDFFX1 DFF_261_Q_reg ( .D(WX2011), .SI(WX2010), .SE(n10329), .CLK(n10725), 
        .Q(WX2012), .QN(n9260) );
  SDFFX1 DFF_262_Q_reg ( .D(WX2013), .SI(WX2012), .SE(n10329), .CLK(n10725), 
        .Q(WX2014), .QN(n9258) );
  SDFFX1 DFF_263_Q_reg ( .D(WX2015), .SI(WX2014), .SE(n10328), .CLK(n10726), 
        .Q(WX2016), .QN(n9256) );
  SDFFX1 DFF_264_Q_reg ( .D(WX2017), .SI(WX2016), .SE(n10327), .CLK(n10726), 
        .Q(WX2018), .QN(n9254) );
  SDFFX1 DFF_265_Q_reg ( .D(WX2019), .SI(WX2018), .SE(n10327), .CLK(n10726), 
        .Q(WX2020), .QN(n9252) );
  SDFFX1 DFF_266_Q_reg ( .D(WX2021), .SI(WX2020), .SE(n10326), .CLK(n10727), 
        .Q(WX2022), .QN(n9250) );
  SDFFX1 DFF_267_Q_reg ( .D(WX2023), .SI(WX2022), .SE(n10325), .CLK(n10727), 
        .Q(WX2024), .QN(n9248) );
  SDFFX1 DFF_268_Q_reg ( .D(WX2025), .SI(WX2024), .SE(n10325), .CLK(n10727), 
        .Q(WX2026), .QN(n9246) );
  SDFFX1 DFF_269_Q_reg ( .D(WX2027), .SI(WX2026), .SE(n10324), .CLK(n10728), 
        .Q(test_so15), .QN(n9962) );
  SDFFX1 DFF_270_Q_reg ( .D(WX2029), .SI(test_si16), .SE(n10323), .CLK(n10728), 
        .Q(WX2030), .QN(n9243) );
  SDFFX1 DFF_271_Q_reg ( .D(WX2031), .SI(WX2030), .SE(n10323), .CLK(n10728), 
        .Q(WX2032), .QN(n9241) );
  SDFFX1 DFF_272_Q_reg ( .D(WX2033), .SI(WX2032), .SE(n10322), .CLK(n10729), 
        .Q(WX2034), .QN(n3785) );
  SDFFX1 DFF_273_Q_reg ( .D(WX2035), .SI(WX2034), .SE(n10321), .CLK(n10729), 
        .Q(WX2036), .QN(n3783) );
  SDFFX1 DFF_274_Q_reg ( .D(WX2037), .SI(WX2036), .SE(n10321), .CLK(n10729), 
        .Q(WX2038), .QN(n3781) );
  SDFFX1 DFF_275_Q_reg ( .D(WX2039), .SI(WX2038), .SE(n10320), .CLK(n10730), 
        .Q(WX2040), .QN(n3779) );
  SDFFX1 DFF_276_Q_reg ( .D(WX2041), .SI(WX2040), .SE(n10319), .CLK(n10730), 
        .Q(WX2042), .QN(n3777) );
  SDFFX1 DFF_277_Q_reg ( .D(WX2043), .SI(WX2042), .SE(n10319), .CLK(n10730), 
        .Q(WX2044), .QN(n3775) );
  SDFFX1 DFF_278_Q_reg ( .D(WX2045), .SI(WX2044), .SE(n10318), .CLK(n10730), 
        .Q(WX2046), .QN(n3773) );
  SDFFX1 DFF_279_Q_reg ( .D(WX2047), .SI(WX2046), .SE(n10318), .CLK(n10731), 
        .Q(WX2048), .QN(n3771) );
  SDFFX1 DFF_280_Q_reg ( .D(WX2049), .SI(WX2048), .SE(n10317), .CLK(n10731), 
        .Q(WX2050), .QN(n3769) );
  SDFFX1 DFF_281_Q_reg ( .D(WX2051), .SI(WX2050), .SE(n10317), .CLK(n10731), 
        .Q(WX2052), .QN(n3767) );
  SDFFX1 DFF_282_Q_reg ( .D(WX2053), .SI(WX2052), .SE(n10316), .CLK(n10731), 
        .Q(WX2054), .QN(n3765) );
  SDFFX1 DFF_283_Q_reg ( .D(WX2055), .SI(WX2054), .SE(n10334), .CLK(n10723), 
        .Q(WX2056), .QN(n3763) );
  SDFFX1 DFF_284_Q_reg ( .D(WX2057), .SI(WX2056), .SE(n10333), .CLK(n10723), 
        .Q(WX2058), .QN(n3761) );
  SDFFX1 DFF_285_Q_reg ( .D(WX2059), .SI(WX2058), .SE(n10333), .CLK(n10723), 
        .Q(WX2060), .QN(n3759) );
  SDFFX1 DFF_286_Q_reg ( .D(WX2061), .SI(WX2060), .SE(n10333), .CLK(n10723), 
        .Q(WX2062), .QN(n3757) );
  SDFFX1 DFF_287_Q_reg ( .D(WX2063), .SI(WX2062), .SE(n10332), .CLK(n10724), 
        .Q(test_so16), .QN(n9929) );
  SDFFX1 DFF_288_Q_reg ( .D(WX2065), .SI(test_si17), .SE(n10332), .CLK(n10724), 
        .Q(WX2066), .QN(n9043) );
  SDFFX1 DFF_289_Q_reg ( .D(WX2067), .SI(WX2066), .SE(n10331), .CLK(n10724), 
        .Q(WX2068), .QN(n9269) );
  SDFFX1 DFF_290_Q_reg ( .D(WX2069), .SI(WX2068), .SE(n10331), .CLK(n10724), 
        .Q(WX2070), .QN(n9267) );
  SDFFX1 DFF_291_Q_reg ( .D(WX2071), .SI(WX2070), .SE(n10330), .CLK(n10725), 
        .Q(WX2072) );
  SDFFX1 DFF_292_Q_reg ( .D(WX2073), .SI(WX2072), .SE(n10330), .CLK(n10725), 
        .Q(WX2074), .QN(n9263) );
  SDFFX1 DFF_293_Q_reg ( .D(WX2075), .SI(WX2074), .SE(n10329), .CLK(n10725), 
        .Q(WX2076), .QN(n9261) );
  SDFFX1 DFF_294_Q_reg ( .D(WX2077), .SI(WX2076), .SE(n10329), .CLK(n10725), 
        .Q(WX2078), .QN(n9259) );
  SDFFX1 DFF_295_Q_reg ( .D(WX2079), .SI(WX2078), .SE(n10328), .CLK(n10726), 
        .Q(WX2080), .QN(n9257) );
  SDFFX1 DFF_296_Q_reg ( .D(WX2081), .SI(WX2080), .SE(n10327), .CLK(n10726), 
        .Q(WX2082), .QN(n9255) );
  SDFFX1 DFF_297_Q_reg ( .D(WX2083), .SI(WX2082), .SE(n10326), .CLK(n10726), 
        .Q(WX2084), .QN(n9253) );
  SDFFX1 DFF_298_Q_reg ( .D(WX2085), .SI(WX2084), .SE(n10326), .CLK(n10727), 
        .Q(WX2086), .QN(n9251) );
  SDFFX1 DFF_299_Q_reg ( .D(WX2087), .SI(WX2086), .SE(n10325), .CLK(n10727), 
        .Q(WX2088), .QN(n9249) );
  SDFFX1 DFF_300_Q_reg ( .D(WX2089), .SI(WX2088), .SE(n10325), .CLK(n10727), 
        .Q(WX2090), .QN(n9247) );
  SDFFX1 DFF_301_Q_reg ( .D(WX2091), .SI(WX2090), .SE(n10324), .CLK(n10728), 
        .Q(WX2092), .QN(n9245) );
  SDFFX1 DFF_302_Q_reg ( .D(WX2093), .SI(WX2092), .SE(n10323), .CLK(n10728), 
        .Q(WX2094), .QN(n9244) );
  SDFFX1 DFF_303_Q_reg ( .D(WX2095), .SI(WX2094), .SE(n10323), .CLK(n10728), 
        .Q(WX2096), .QN(n9242) );
  SDFFX1 DFF_304_Q_reg ( .D(WX2097), .SI(WX2096), .SE(n10322), .CLK(n10729), 
        .Q(WX2098), .QN(n9511) );
  SDFFX1 DFF_305_Q_reg ( .D(WX2099), .SI(WX2098), .SE(n10321), .CLK(n10729), 
        .Q(test_so17), .QN(n9933) );
  SDFFX1 DFF_306_Q_reg ( .D(WX2101), .SI(test_si18), .SE(n10320), .CLK(n10729), 
        .Q(WX2102), .QN(n9508) );
  SDFFX1 DFF_307_Q_reg ( .D(WX2103), .SI(WX2102), .SE(n10320), .CLK(n10730), 
        .Q(WX2104), .QN(n9506) );
  SDFFX1 DFF_308_Q_reg ( .D(WX2105), .SI(WX2104), .SE(n10319), .CLK(n10730), 
        .Q(WX2106), .QN(n9504) );
  SDFFX1 DFF_309_Q_reg ( .D(WX2107), .SI(WX2106), .SE(n10319), .CLK(n10730), 
        .Q(WX2108), .QN(n9502) );
  SDFFX1 DFF_310_Q_reg ( .D(WX2109), .SI(WX2108), .SE(n10318), .CLK(n10731), 
        .Q(WX2110), .QN(n9500) );
  SDFFX1 DFF_311_Q_reg ( .D(WX2111), .SI(WX2110), .SE(n10318), .CLK(n10731), 
        .Q(WX2112), .QN(n9498) );
  SDFFX1 DFF_312_Q_reg ( .D(WX2113), .SI(WX2112), .SE(n10317), .CLK(n10731), 
        .Q(WX2114), .QN(n9496) );
  SDFFX1 DFF_313_Q_reg ( .D(WX2115), .SI(WX2114), .SE(n10317), .CLK(n10731), 
        .Q(WX2116), .QN(n9494) );
  SDFFX1 DFF_314_Q_reg ( .D(WX2117), .SI(WX2116), .SE(n10316), .CLK(n10732), 
        .Q(WX2118), .QN(n9492) );
  SDFFX1 DFF_315_Q_reg ( .D(WX2119), .SI(WX2118), .SE(n10316), .CLK(n10732), 
        .Q(WX2120) );
  SDFFX1 DFF_316_Q_reg ( .D(WX2121), .SI(WX2120), .SE(n10316), .CLK(n10732), 
        .Q(WX2122), .QN(n9489) );
  SDFFX1 DFF_317_Q_reg ( .D(WX2123), .SI(WX2122), .SE(n10315), .CLK(n10732), 
        .Q(WX2124), .QN(n9487) );
  SDFFX1 DFF_318_Q_reg ( .D(WX2125), .SI(WX2124), .SE(n10315), .CLK(n10732), 
        .Q(WX2126), .QN(n9485) );
  SDFFX1 DFF_319_Q_reg ( .D(WX2127), .SI(WX2126), .SE(n10315), .CLK(n10732), 
        .Q(WX2128) );
  SDFFX1 DFF_320_Q_reg ( .D(WX2129), .SI(WX2128), .SE(n10314), .CLK(n10733), 
        .Q(WX2130), .QN(n9727) );
  SDFFX1 DFF_321_Q_reg ( .D(WX2131), .SI(WX2130), .SE(n10314), .CLK(n10733), 
        .Q(WX2132), .QN(n9728) );
  SDFFX1 DFF_322_Q_reg ( .D(WX2133), .SI(WX2132), .SE(n10314), .CLK(n10733), 
        .Q(WX2134), .QN(n9729) );
  SDFFX1 DFF_323_Q_reg ( .D(WX2135), .SI(WX2134), .SE(n10314), .CLK(n10733), 
        .Q(test_so18), .QN(n9912) );
  SDFFX1 DFF_324_Q_reg ( .D(WX2137), .SI(test_si19), .SE(n10330), .CLK(n10725), 
        .Q(WX2138), .QN(n9730) );
  SDFFX1 DFF_325_Q_reg ( .D(WX2139), .SI(WX2138), .SE(n10329), .CLK(n10725), 
        .Q(WX2140), .QN(n9731) );
  SDFFX1 DFF_326_Q_reg ( .D(WX2141), .SI(WX2140), .SE(n10328), .CLK(n10725), 
        .Q(WX2142), .QN(n9732) );
  SDFFX1 DFF_327_Q_reg ( .D(WX2143), .SI(WX2142), .SE(n10328), .CLK(n10726), 
        .Q(WX2144), .QN(n9733) );
  SDFFX1 DFF_328_Q_reg ( .D(WX2145), .SI(WX2144), .SE(n10327), .CLK(n10726), 
        .Q(WX2146), .QN(n9734) );
  SDFFX1 DFF_329_Q_reg ( .D(WX2147), .SI(WX2146), .SE(n10326), .CLK(n10727), 
        .Q(WX2148), .QN(n9735) );
  SDFFX1 DFF_330_Q_reg ( .D(WX2149), .SI(WX2148), .SE(n10326), .CLK(n10727), 
        .Q(WX2150), .QN(n9736) );
  SDFFX1 DFF_331_Q_reg ( .D(WX2151), .SI(WX2150), .SE(n10325), .CLK(n10727), 
        .Q(WX2152), .QN(n9737) );
  SDFFX1 DFF_332_Q_reg ( .D(WX2153), .SI(WX2152), .SE(n10324), .CLK(n10727), 
        .Q(WX2154), .QN(n9738) );
  SDFFX1 DFF_333_Q_reg ( .D(WX2155), .SI(WX2154), .SE(n10324), .CLK(n10728), 
        .Q(WX2156), .QN(n9739) );
  SDFFX1 DFF_334_Q_reg ( .D(WX2157), .SI(WX2156), .SE(n10323), .CLK(n10728), 
        .Q(WX2158), .QN(n9740) );
  SDFFX1 DFF_335_Q_reg ( .D(WX2159), .SI(WX2158), .SE(n10322), .CLK(n10728), 
        .Q(WX2160), .QN(n9530) );
  SDFFX1 DFF_336_Q_reg ( .D(WX2161), .SI(WX2160), .SE(n10322), .CLK(n10729), 
        .Q(WX2162), .QN(n9741) );
  SDFFX1 DFF_337_Q_reg ( .D(WX2163), .SI(WX2162), .SE(n10321), .CLK(n10729), 
        .Q(WX2164), .QN(n9742) );
  SDFFX1 DFF_338_Q_reg ( .D(WX2165), .SI(WX2164), .SE(n10320), .CLK(n10730), 
        .Q(WX2166), .QN(n9743) );
  SDFFX1 DFF_339_Q_reg ( .D(WX2167), .SI(WX2166), .SE(n10320), .CLK(n10730), 
        .Q(WX2168), .QN(n9744) );
  SDFFX1 DFF_340_Q_reg ( .D(WX2169), .SI(WX2168), .SE(n10319), .CLK(n10730), 
        .Q(WX2170), .QN(n9531) );
  SDFFX1 DFF_341_Q_reg ( .D(WX2171), .SI(WX2170), .SE(n10319), .CLK(n10730), 
        .Q(test_so19), .QN(n9905) );
  SDFFX1 DFF_342_Q_reg ( .D(WX2173), .SI(test_si20), .SE(n10318), .CLK(n10731), 
        .Q(WX2174), .QN(n9745) );
  SDFFX1 DFF_343_Q_reg ( .D(WX2175), .SI(WX2174), .SE(n10318), .CLK(n10731), 
        .Q(WX2176), .QN(n9746) );
  SDFFX1 DFF_344_Q_reg ( .D(WX2177), .SI(WX2176), .SE(n10317), .CLK(n10731), 
        .Q(WX2178), .QN(n9747) );
  SDFFX1 DFF_345_Q_reg ( .D(WX2179), .SI(WX2178), .SE(n10317), .CLK(n10731), 
        .Q(WX2180), .QN(n9748) );
  SDFFX1 DFF_346_Q_reg ( .D(WX2181), .SI(WX2180), .SE(n10316), .CLK(n10732), 
        .Q(WX2182), .QN(n9749) );
  SDFFX1 DFF_347_Q_reg ( .D(WX2183), .SI(WX2182), .SE(n10316), .CLK(n10732), 
        .Q(WX2184), .QN(n9532) );
  SDFFX1 DFF_348_Q_reg ( .D(WX2185), .SI(WX2184), .SE(n10315), .CLK(n10732), 
        .Q(WX2186), .QN(n9750) );
  SDFFX1 DFF_349_Q_reg ( .D(WX2187), .SI(WX2186), .SE(n10315), .CLK(n10732), 
        .Q(WX2188), .QN(n9751) );
  SDFFX1 DFF_350_Q_reg ( .D(WX2189), .SI(WX2188), .SE(n10315), .CLK(n10732), 
        .Q(WX2190), .QN(n9752) );
  SDFFX1 DFF_351_Q_reg ( .D(WX2191), .SI(WX2190), .SE(n10314), .CLK(n10732), 
        .Q(WX2192), .QN(n9540) );
  SDFFX1 DFF_352_Q_reg ( .D(WX2557), .SI(WX2192), .SE(n10092), .CLK(n10844), 
        .Q(CRC_OUT_8_0), .QN(DFF_352_n1) );
  SDFFX1 DFF_353_Q_reg ( .D(WX2559), .SI(CRC_OUT_8_0), .SE(n10092), .CLK(
        n10844), .Q(CRC_OUT_8_1), .QN(DFF_353_n1) );
  SDFFX1 DFF_354_Q_reg ( .D(WX2561), .SI(CRC_OUT_8_1), .SE(n10092), .CLK(
        n10844), .Q(CRC_OUT_8_2), .QN(DFF_354_n1) );
  SDFFX1 DFF_355_Q_reg ( .D(WX2563), .SI(CRC_OUT_8_2), .SE(n10091), .CLK(
        n10845), .Q(CRC_OUT_8_3), .QN(DFF_355_n1) );
  SDFFX1 DFF_356_Q_reg ( .D(WX2565), .SI(CRC_OUT_8_3), .SE(n10091), .CLK(
        n10845), .Q(CRC_OUT_8_4), .QN(DFF_356_n1) );
  SDFFX1 DFF_357_Q_reg ( .D(WX2567), .SI(CRC_OUT_8_4), .SE(n10091), .CLK(
        n10845), .Q(CRC_OUT_8_5), .QN(DFF_357_n1) );
  SDFFX1 DFF_358_Q_reg ( .D(WX2569), .SI(CRC_OUT_8_5), .SE(n10091), .CLK(
        n10845), .Q(CRC_OUT_8_6), .QN(DFF_358_n1) );
  SDFFX1 DFF_359_Q_reg ( .D(WX2571), .SI(CRC_OUT_8_6), .SE(n10091), .CLK(
        n10845), .Q(test_so20), .QN(n9947) );
  SDFFX1 DFF_360_Q_reg ( .D(WX2573), .SI(test_si21), .SE(n10091), .CLK(n10845), 
        .Q(CRC_OUT_8_8), .QN(DFF_360_n1) );
  SDFFX1 DFF_361_Q_reg ( .D(WX2575), .SI(CRC_OUT_8_8), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_9), .QN(DFF_361_n1) );
  SDFFX1 DFF_362_Q_reg ( .D(WX2577), .SI(CRC_OUT_8_9), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_10), .QN(DFF_362_n1) );
  SDFFX1 DFF_363_Q_reg ( .D(WX2579), .SI(CRC_OUT_8_10), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_11), .QN(DFF_363_n1) );
  SDFFX1 DFF_364_Q_reg ( .D(WX2581), .SI(CRC_OUT_8_11), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_12), .QN(DFF_364_n1) );
  SDFFX1 DFF_365_Q_reg ( .D(WX2583), .SI(CRC_OUT_8_12), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_13), .QN(DFF_365_n1) );
  SDFFX1 DFF_366_Q_reg ( .D(WX2585), .SI(CRC_OUT_8_13), .SE(n10090), .CLK(
        n10845), .Q(CRC_OUT_8_14), .QN(DFF_366_n1) );
  SDFFX1 DFF_367_Q_reg ( .D(WX2587), .SI(CRC_OUT_8_14), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_15), .QN(DFF_367_n1) );
  SDFFX1 DFF_368_Q_reg ( .D(WX2589), .SI(CRC_OUT_8_15), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_16), .QN(DFF_368_n1) );
  SDFFX1 DFF_369_Q_reg ( .D(WX2591), .SI(CRC_OUT_8_16), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_17), .QN(DFF_369_n1) );
  SDFFX1 DFF_370_Q_reg ( .D(WX2593), .SI(CRC_OUT_8_17), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_18), .QN(DFF_370_n1) );
  SDFFX1 DFF_371_Q_reg ( .D(WX2595), .SI(CRC_OUT_8_18), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_19), .QN(DFF_371_n1) );
  SDFFX1 DFF_372_Q_reg ( .D(WX2597), .SI(CRC_OUT_8_19), .SE(n10089), .CLK(
        n10846), .Q(CRC_OUT_8_20), .QN(DFF_372_n1) );
  SDFFX1 DFF_373_Q_reg ( .D(WX2599), .SI(CRC_OUT_8_20), .SE(n10088), .CLK(
        n10846), .Q(CRC_OUT_8_21), .QN(DFF_373_n1) );
  SDFFX1 DFF_374_Q_reg ( .D(WX2601), .SI(CRC_OUT_8_21), .SE(n10088), .CLK(
        n10846), .Q(CRC_OUT_8_22), .QN(DFF_374_n1) );
  SDFFX1 DFF_375_Q_reg ( .D(WX2603), .SI(CRC_OUT_8_22), .SE(n10088), .CLK(
        n10846), .Q(CRC_OUT_8_23), .QN(DFF_375_n1) );
  SDFFX1 DFF_376_Q_reg ( .D(WX2605), .SI(CRC_OUT_8_23), .SE(n10088), .CLK(
        n10846), .Q(CRC_OUT_8_24), .QN(DFF_376_n1) );
  SDFFX1 DFF_377_Q_reg ( .D(WX2607), .SI(CRC_OUT_8_24), .SE(n10088), .CLK(
        n10846), .Q(test_so21), .QN(n9946) );
  SDFFX1 DFF_378_Q_reg ( .D(WX2609), .SI(test_si22), .SE(n10088), .CLK(n10846), 
        .Q(CRC_OUT_8_26), .QN(DFF_378_n1) );
  SDFFX1 DFF_379_Q_reg ( .D(WX2611), .SI(CRC_OUT_8_26), .SE(n10087), .CLK(
        n10847), .Q(CRC_OUT_8_27), .QN(DFF_379_n1) );
  SDFFX1 DFF_380_Q_reg ( .D(WX2613), .SI(CRC_OUT_8_27), .SE(n10087), .CLK(
        n10847), .Q(CRC_OUT_8_28), .QN(DFF_380_n1) );
  SDFFX1 DFF_381_Q_reg ( .D(WX2615), .SI(CRC_OUT_8_28), .SE(n10087), .CLK(
        n10847), .Q(CRC_OUT_8_29), .QN(DFF_381_n1) );
  SDFFX1 DFF_382_Q_reg ( .D(WX2617), .SI(CRC_OUT_8_29), .SE(n10087), .CLK(
        n10847), .Q(CRC_OUT_8_30), .QN(DFF_382_n1) );
  SDFFX1 DFF_383_Q_reg ( .D(WX2619), .SI(CRC_OUT_8_30), .SE(n10314), .CLK(
        n10733), .Q(CRC_OUT_8_31), .QN(DFF_383_n1) );
  SDFFX1 DFF_384_Q_reg ( .D(n491), .SI(CRC_OUT_8_31), .SE(n10313), .CLK(n10733), .Q(WX3071), .QN(n9845) );
  SDFFX1 DFF_385_Q_reg ( .D(n492), .SI(WX3071), .SE(n10308), .CLK(n10736), .Q(
        n8644), .QN(n4002) );
  SDFFX1 DFF_386_Q_reg ( .D(n493), .SI(n8644), .SE(n10308), .CLK(n10735), .Q(
        n8643), .QN(n4001) );
  SDFFX1 DFF_387_Q_reg ( .D(n494), .SI(n8643), .SE(n10309), .CLK(n10735), .Q(
        n8642), .QN(n4000) );
  SDFFX1 DFF_388_Q_reg ( .D(n495), .SI(n8642), .SE(n10309), .CLK(n10735), .Q(
        n8641), .QN(n3999) );
  SDFFX1 DFF_389_Q_reg ( .D(n496), .SI(n8641), .SE(n10309), .CLK(n10735), .Q(
        n8640), .QN(n3998) );
  SDFFX1 DFF_390_Q_reg ( .D(n497), .SI(n8640), .SE(n10309), .CLK(n10735), .Q(
        n8639), .QN(n3997) );
  SDFFX1 DFF_391_Q_reg ( .D(n498), .SI(n8639), .SE(n10309), .CLK(n10735), .Q(
        n8638), .QN(n3996) );
  SDFFX1 DFF_392_Q_reg ( .D(n499), .SI(n8638), .SE(n10309), .CLK(n10735), .Q(
        n8637), .QN(n3995) );
  SDFFX1 DFF_393_Q_reg ( .D(n500), .SI(n8637), .SE(n10310), .CLK(n10735), .Q(
        n8636), .QN(n3994) );
  SDFFX1 DFF_394_Q_reg ( .D(n501), .SI(n8636), .SE(n10310), .CLK(n10735), .Q(
        n8635), .QN(n3993) );
  SDFFX1 DFF_395_Q_reg ( .D(n502), .SI(n8635), .SE(n10310), .CLK(n10735), .Q(
        test_so22), .QN(n3992) );
  SDFFX1 DFF_396_Q_reg ( .D(n503), .SI(test_si23), .SE(n10310), .CLK(n10735), 
        .Q(n8632), .QN(n3991) );
  SDFFX1 DFF_397_Q_reg ( .D(n504), .SI(n8632), .SE(n10310), .CLK(n10735), .Q(
        n8631), .QN(n3990) );
  SDFFX1 DFF_398_Q_reg ( .D(n505), .SI(n8631), .SE(n10310), .CLK(n10734), .Q(
        n8630), .QN(n3989) );
  SDFFX1 DFF_399_Q_reg ( .D(n506), .SI(n8630), .SE(n10311), .CLK(n10734), .Q(
        n8629), .QN(n3988) );
  SDFFX1 DFF_400_Q_reg ( .D(n507), .SI(n8629), .SE(n10311), .CLK(n10734), .Q(
        n8628), .QN(n3987) );
  SDFFX1 DFF_401_Q_reg ( .D(n508), .SI(n8628), .SE(n10311), .CLK(n10734), .Q(
        n8627), .QN(n3986) );
  SDFFX1 DFF_402_Q_reg ( .D(n509), .SI(n8627), .SE(n10311), .CLK(n10734), .Q(
        n8626), .QN(n3985) );
  SDFFX1 DFF_403_Q_reg ( .D(n510), .SI(n8626), .SE(n10311), .CLK(n10734), .Q(
        n8625), .QN(n3984) );
  SDFFX1 DFF_404_Q_reg ( .D(n511), .SI(n8625), .SE(n10311), .CLK(n10734), .Q(
        n8624), .QN(n3983) );
  SDFFX1 DFF_405_Q_reg ( .D(n512), .SI(n8624), .SE(n10312), .CLK(n10734), .Q(
        n8623), .QN(n3982) );
  SDFFX1 DFF_406_Q_reg ( .D(n513), .SI(n8623), .SE(n10312), .CLK(n10734), .Q(
        n8622), .QN(n3981) );
  SDFFX1 DFF_407_Q_reg ( .D(n514), .SI(n8622), .SE(n10312), .CLK(n10734), .Q(
        n8621), .QN(n3980) );
  SDFFX1 DFF_408_Q_reg ( .D(n515), .SI(n8621), .SE(n10312), .CLK(n10734), .Q(
        n8620), .QN(n3979) );
  SDFFX1 DFF_409_Q_reg ( .D(n516), .SI(n8620), .SE(n10312), .CLK(n10734), .Q(
        n8619), .QN(n3978) );
  SDFFX1 DFF_410_Q_reg ( .D(n517), .SI(n8619), .SE(n10312), .CLK(n10733), .Q(
        n8618), .QN(n3977) );
  SDFFX1 DFF_411_Q_reg ( .D(n518), .SI(n8618), .SE(n10313), .CLK(n10733), .Q(
        n8617), .QN(n3976) );
  SDFFX1 DFF_412_Q_reg ( .D(n519), .SI(n8617), .SE(n10313), .CLK(n10733), .Q(
        n8616), .QN(n3975) );
  SDFFX1 DFF_413_Q_reg ( .D(n520), .SI(n8616), .SE(n10313), .CLK(n10733), .Q(
        test_so23), .QN(n3974) );
  SDFFX1 DFF_414_Q_reg ( .D(n521), .SI(test_si24), .SE(n10313), .CLK(n10733), 
        .Q(n8613), .QN(n3973) );
  SDFFX1 DFF_415_Q_reg ( .D(WX3132), .SI(n8613), .SE(n10313), .CLK(n10733), 
        .Q(n8612), .QN(n3972) );
  SDFFX1 DFF_416_Q_reg ( .D(WX3230), .SI(n8612), .SE(n10092), .CLK(n10844), 
        .Q(n8611), .QN(n17985) );
  SDFFX1 DFF_417_Q_reg ( .D(WX3232), .SI(n8611), .SE(n10308), .CLK(n10736), 
        .Q(n8610), .QN(n17984) );
  SDFFX1 DFF_418_Q_reg ( .D(WX3234), .SI(n8610), .SE(n10307), .CLK(n10736), 
        .Q(n8609), .QN(n17982) );
  SDFFX1 DFF_419_Q_reg ( .D(WX3236), .SI(n8609), .SE(n10307), .CLK(n10736), 
        .Q(n8608), .QN(n17980) );
  SDFFX1 DFF_420_Q_reg ( .D(WX3238), .SI(n8608), .SE(n10307), .CLK(n10736), 
        .Q(n8607), .QN(n17978) );
  SDFFX1 DFF_421_Q_reg ( .D(WX3240), .SI(n8607), .SE(n10306), .CLK(n10737), 
        .Q(n8606), .QN(n17976) );
  SDFFX1 DFF_422_Q_reg ( .D(WX3242), .SI(n8606), .SE(n10306), .CLK(n10737), 
        .Q(n8605), .QN(n17974) );
  SDFFX1 DFF_423_Q_reg ( .D(WX3244), .SI(n8605), .SE(n10305), .CLK(n10737), 
        .Q(n8604), .QN(n17972) );
  SDFFX1 DFF_424_Q_reg ( .D(WX3246), .SI(n8604), .SE(n10305), .CLK(n10737), 
        .Q(n8603), .QN(n17970) );
  SDFFX1 DFF_425_Q_reg ( .D(WX3248), .SI(n8603), .SE(n10304), .CLK(n10738), 
        .Q(n8602), .QN(n17968) );
  SDFFX1 DFF_426_Q_reg ( .D(WX3250), .SI(n8602), .SE(n10303), .CLK(n10738), 
        .Q(n8601), .QN(n17967) );
  SDFFX1 DFF_427_Q_reg ( .D(WX3252), .SI(n8601), .SE(n10302), .CLK(n10739), 
        .Q(n8600), .QN(n17965) );
  SDFFX1 DFF_428_Q_reg ( .D(WX3254), .SI(n8600), .SE(n10302), .CLK(n10739), 
        .Q(n8599), .QN(n17963) );
  SDFFX1 DFF_429_Q_reg ( .D(WX3256), .SI(n8599), .SE(n10301), .CLK(n10739), 
        .Q(n8598), .QN(n17961) );
  SDFFX1 DFF_430_Q_reg ( .D(WX3258), .SI(n8598), .SE(n10301), .CLK(n10739), 
        .Q(n8597), .QN(n17959) );
  SDFFX1 DFF_431_Q_reg ( .D(WX3260), .SI(n8597), .SE(n10092), .CLK(n10844), 
        .Q(test_so24), .QN(n9894) );
  SDFFX1 DFF_432_Q_reg ( .D(WX3262), .SI(test_si25), .SE(n10299), .CLK(n10740), 
        .Q(WX3263), .QN(n9480) );
  SDFFX1 DFF_433_Q_reg ( .D(WX3264), .SI(WX3263), .SE(n10299), .CLK(n10740), 
        .Q(WX3265), .QN(n9478) );
  SDFFX1 DFF_434_Q_reg ( .D(WX3266), .SI(WX3265), .SE(n10298), .CLK(n10741), 
        .Q(WX3267), .QN(n9476) );
  SDFFX1 DFF_435_Q_reg ( .D(WX3268), .SI(WX3267), .SE(n10298), .CLK(n10741), 
        .Q(WX3269), .QN(n9474) );
  SDFFX1 DFF_436_Q_reg ( .D(WX3270), .SI(WX3269), .SE(n10335), .CLK(n10722), 
        .Q(WX3271), .QN(n9472) );
  SDFFX1 DFF_437_Q_reg ( .D(WX3272), .SI(WX3271), .SE(n10296), .CLK(n10742), 
        .Q(WX3273), .QN(n9470) );
  SDFFX1 DFF_438_Q_reg ( .D(WX3274), .SI(WX3273), .SE(n10296), .CLK(n10742), 
        .Q(WX3275), .QN(n9468) );
  SDFFX1 DFF_439_Q_reg ( .D(WX3276), .SI(WX3275), .SE(n10295), .CLK(n10742), 
        .Q(WX3277) );
  SDFFX1 DFF_440_Q_reg ( .D(WX3278), .SI(WX3277), .SE(n10295), .CLK(n10742), 
        .Q(WX3279), .QN(n9465) );
  SDFFX1 DFF_441_Q_reg ( .D(WX3280), .SI(WX3279), .SE(n10294), .CLK(n10743), 
        .Q(WX3281) );
  SDFFX1 DFF_442_Q_reg ( .D(WX3282), .SI(WX3281), .SE(n10293), .CLK(n10743), 
        .Q(WX3283), .QN(n9461) );
  SDFFX1 DFF_443_Q_reg ( .D(WX3284), .SI(WX3283), .SE(n10293), .CLK(n10743), 
        .Q(WX3285), .QN(n9459) );
  SDFFX1 DFF_444_Q_reg ( .D(WX3286), .SI(WX3285), .SE(n10292), .CLK(n10744), 
        .Q(WX3287), .QN(n9457) );
  SDFFX1 DFF_445_Q_reg ( .D(WX3288), .SI(WX3287), .SE(n10291), .CLK(n10744), 
        .Q(WX3289), .QN(n9455) );
  SDFFX1 DFF_446_Q_reg ( .D(WX3290), .SI(WX3289), .SE(n10291), .CLK(n10744), 
        .Q(WX3291), .QN(n9453) );
  SDFFX1 DFF_447_Q_reg ( .D(WX3292), .SI(WX3291), .SE(n10290), .CLK(n10745), 
        .Q(WX3293), .QN(n9451) );
  SDFFX1 DFF_448_Q_reg ( .D(WX3294), .SI(WX3293), .SE(n10289), .CLK(n10745), 
        .Q(WX3295), .QN(n9040) );
  SDFFX1 DFF_449_Q_reg ( .D(WX3296), .SI(WX3295), .SE(n10308), .CLK(n10736), 
        .Q(test_so25), .QN(n9964) );
  SDFFX1 DFF_450_Q_reg ( .D(WX3298), .SI(test_si26), .SE(n10307), .CLK(n10736), 
        .Q(WX3299), .QN(n9238) );
  SDFFX1 DFF_451_Q_reg ( .D(WX3300), .SI(WX3299), .SE(n10307), .CLK(n10736), 
        .Q(WX3301), .QN(n9236) );
  SDFFX1 DFF_452_Q_reg ( .D(WX3302), .SI(WX3301), .SE(n10306), .CLK(n10736), 
        .Q(WX3303), .QN(n9234) );
  SDFFX1 DFF_453_Q_reg ( .D(WX3304), .SI(WX3303), .SE(n10306), .CLK(n10737), 
        .Q(WX3305), .QN(n9233) );
  SDFFX1 DFF_454_Q_reg ( .D(WX3306), .SI(WX3305), .SE(n10305), .CLK(n10737), 
        .Q(WX3307), .QN(n9231) );
  SDFFX1 DFF_455_Q_reg ( .D(WX3308), .SI(WX3307), .SE(n10305), .CLK(n10737), 
        .Q(WX3309), .QN(n9229) );
  SDFFX1 DFF_456_Q_reg ( .D(WX3310), .SI(WX3309), .SE(n10304), .CLK(n10737), 
        .Q(WX3311), .QN(n9227) );
  SDFFX1 DFF_457_Q_reg ( .D(WX3312), .SI(WX3311), .SE(n10304), .CLK(n10738), 
        .Q(WX3313), .QN(n9225) );
  SDFFX1 DFF_458_Q_reg ( .D(WX3314), .SI(WX3313), .SE(n10303), .CLK(n10738), 
        .Q(WX3315), .QN(n9223) );
  SDFFX1 DFF_459_Q_reg ( .D(WX3316), .SI(WX3315), .SE(n10303), .CLK(n10738), 
        .Q(WX3317), .QN(n9221) );
  SDFFX1 DFF_460_Q_reg ( .D(WX3318), .SI(WX3317), .SE(n10302), .CLK(n10739), 
        .Q(WX3319), .QN(n9219) );
  SDFFX1 DFF_461_Q_reg ( .D(WX3320), .SI(WX3319), .SE(n10301), .CLK(n10739), 
        .Q(WX3321), .QN(n9217) );
  SDFFX1 DFF_462_Q_reg ( .D(WX3322), .SI(WX3321), .SE(n10301), .CLK(n10739), 
        .Q(WX3323), .QN(n9215) );
  SDFFX1 DFF_463_Q_reg ( .D(WX3324), .SI(WX3323), .SE(n10300), .CLK(n10740), 
        .Q(WX3325), .QN(n9213) );
  SDFFX1 DFF_464_Q_reg ( .D(WX3326), .SI(WX3325), .SE(n10300), .CLK(n10740), 
        .Q(WX3327), .QN(n3753) );
  SDFFX1 DFF_465_Q_reg ( .D(WX3328), .SI(WX3327), .SE(n10299), .CLK(n10740), 
        .Q(WX3329), .QN(n3751) );
  SDFFX1 DFF_466_Q_reg ( .D(WX3330), .SI(WX3329), .SE(n10298), .CLK(n10741), 
        .Q(WX3331), .QN(n3749) );
  SDFFX1 DFF_467_Q_reg ( .D(WX3332), .SI(WX3331), .SE(n10297), .CLK(n10741), 
        .Q(test_so26), .QN(n9932) );
  SDFFX1 DFF_468_Q_reg ( .D(WX3334), .SI(test_si27), .SE(n10335), .CLK(n10722), 
        .Q(WX3335), .QN(n3745) );
  SDFFX1 DFF_469_Q_reg ( .D(WX3336), .SI(WX3335), .SE(n10296), .CLK(n10742), 
        .Q(WX3337), .QN(n3743) );
  SDFFX1 DFF_470_Q_reg ( .D(WX3338), .SI(WX3337), .SE(n10296), .CLK(n10742), 
        .Q(WX3339), .QN(n3741) );
  SDFFX1 DFF_471_Q_reg ( .D(WX3340), .SI(WX3339), .SE(n10295), .CLK(n10742), 
        .Q(WX3341), .QN(n3739) );
  SDFFX1 DFF_472_Q_reg ( .D(WX3342), .SI(WX3341), .SE(n10294), .CLK(n10742), 
        .Q(WX3343), .QN(n3737) );
  SDFFX1 DFF_473_Q_reg ( .D(WX3344), .SI(WX3343), .SE(n10294), .CLK(n10743), 
        .Q(WX3345), .QN(n3735) );
  SDFFX1 DFF_474_Q_reg ( .D(WX3346), .SI(WX3345), .SE(n10293), .CLK(n10743), 
        .Q(WX3347), .QN(n3733) );
  SDFFX1 DFF_475_Q_reg ( .D(WX3348), .SI(WX3347), .SE(n10292), .CLK(n10743), 
        .Q(WX3349), .QN(n3731) );
  SDFFX1 DFF_476_Q_reg ( .D(WX3350), .SI(WX3349), .SE(n10292), .CLK(n10744), 
        .Q(WX3351), .QN(n3729) );
  SDFFX1 DFF_477_Q_reg ( .D(WX3352), .SI(WX3351), .SE(n10291), .CLK(n10744), 
        .Q(WX3353), .QN(n3727) );
  SDFFX1 DFF_478_Q_reg ( .D(WX3354), .SI(WX3353), .SE(n10290), .CLK(n10744), 
        .Q(WX3355), .QN(n3725) );
  SDFFX1 DFF_479_Q_reg ( .D(WX3356), .SI(WX3355), .SE(n10290), .CLK(n10745), 
        .Q(WX3357), .QN(n3723) );
  SDFFX1 DFF_480_Q_reg ( .D(WX3358), .SI(WX3357), .SE(n10289), .CLK(n10745), 
        .Q(WX3359), .QN(n9041) );
  SDFFX1 DFF_481_Q_reg ( .D(WX3360), .SI(WX3359), .SE(n10308), .CLK(n10736), 
        .Q(WX3361), .QN(n9240) );
  SDFFX1 DFF_482_Q_reg ( .D(WX3362), .SI(WX3361), .SE(n10308), .CLK(n10736), 
        .Q(WX3363), .QN(n9239) );
  SDFFX1 DFF_483_Q_reg ( .D(WX3364), .SI(WX3363), .SE(n10307), .CLK(n10736), 
        .Q(WX3365), .QN(n9237) );
  SDFFX1 DFF_484_Q_reg ( .D(WX3366), .SI(WX3365), .SE(n10306), .CLK(n10737), 
        .Q(WX3367), .QN(n9235) );
  SDFFX1 DFF_485_Q_reg ( .D(WX3368), .SI(WX3367), .SE(n10306), .CLK(n10737), 
        .Q(test_so27), .QN(n9963) );
  SDFFX1 DFF_486_Q_reg ( .D(WX3370), .SI(test_si28), .SE(n10305), .CLK(n10737), 
        .Q(WX3371), .QN(n9232) );
  SDFFX1 DFF_487_Q_reg ( .D(WX3372), .SI(WX3371), .SE(n10305), .CLK(n10737), 
        .Q(WX3373), .QN(n9230) );
  SDFFX1 DFF_488_Q_reg ( .D(WX3374), .SI(WX3373), .SE(n10304), .CLK(n10738), 
        .Q(WX3375) );
  SDFFX1 DFF_489_Q_reg ( .D(WX3376), .SI(WX3375), .SE(n10304), .CLK(n10738), 
        .Q(WX3377), .QN(n9226) );
  SDFFX1 DFF_490_Q_reg ( .D(WX3378), .SI(WX3377), .SE(n10303), .CLK(n10738), 
        .Q(WX3379), .QN(n9224) );
  SDFFX1 DFF_491_Q_reg ( .D(WX3380), .SI(WX3379), .SE(n10303), .CLK(n10738), 
        .Q(WX3381), .QN(n9222) );
  SDFFX1 DFF_492_Q_reg ( .D(WX3382), .SI(WX3381), .SE(n10302), .CLK(n10739), 
        .Q(WX3383), .QN(n9220) );
  SDFFX1 DFF_493_Q_reg ( .D(WX3384), .SI(WX3383), .SE(n10301), .CLK(n10739), 
        .Q(WX3385), .QN(n9218) );
  SDFFX1 DFF_494_Q_reg ( .D(WX3386), .SI(WX3385), .SE(n10300), .CLK(n10739), 
        .Q(WX3387), .QN(n9216) );
  SDFFX1 DFF_495_Q_reg ( .D(WX3388), .SI(WX3387), .SE(n10300), .CLK(n10740), 
        .Q(WX3389), .QN(n9214) );
  SDFFX1 DFF_496_Q_reg ( .D(WX3390), .SI(WX3389), .SE(n10299), .CLK(n10740), 
        .Q(WX3391), .QN(n9481) );
  SDFFX1 DFF_497_Q_reg ( .D(WX3392), .SI(WX3391), .SE(n10299), .CLK(n10740), 
        .Q(WX3393), .QN(n9479) );
  SDFFX1 DFF_498_Q_reg ( .D(WX3394), .SI(WX3393), .SE(n10298), .CLK(n10741), 
        .Q(WX3395), .QN(n9477) );
  SDFFX1 DFF_499_Q_reg ( .D(WX3396), .SI(WX3395), .SE(n10297), .CLK(n10741), 
        .Q(WX3397) );
  SDFFX1 DFF_500_Q_reg ( .D(WX3398), .SI(WX3397), .SE(n10297), .CLK(n10741), 
        .Q(WX3399), .QN(n9473) );
  SDFFX1 DFF_501_Q_reg ( .D(WX3400), .SI(WX3399), .SE(n10297), .CLK(n10741), 
        .Q(WX3401), .QN(n9471) );
  SDFFX1 DFF_502_Q_reg ( .D(WX3402), .SI(WX3401), .SE(n10296), .CLK(n10742), 
        .Q(WX3403), .QN(n9469) );
  SDFFX1 DFF_503_Q_reg ( .D(WX3404), .SI(WX3403), .SE(n10295), .CLK(n10742), 
        .Q(test_so28), .QN(n9931) );
  SDFFX1 DFF_504_Q_reg ( .D(WX3406), .SI(test_si29), .SE(n10294), .CLK(n10743), 
        .Q(WX3407), .QN(n9466) );
  SDFFX1 DFF_505_Q_reg ( .D(WX3408), .SI(WX3407), .SE(n10294), .CLK(n10743), 
        .Q(WX3409), .QN(n9464) );
  SDFFX1 DFF_506_Q_reg ( .D(WX3410), .SI(WX3409), .SE(n10293), .CLK(n10743), 
        .Q(WX3411), .QN(n9462) );
  SDFFX1 DFF_507_Q_reg ( .D(WX3412), .SI(WX3411), .SE(n10292), .CLK(n10744), 
        .Q(WX3413), .QN(n9460) );
  SDFFX1 DFF_508_Q_reg ( .D(WX3414), .SI(WX3413), .SE(n10292), .CLK(n10744), 
        .Q(WX3415), .QN(n9458) );
  SDFFX1 DFF_509_Q_reg ( .D(WX3416), .SI(WX3415), .SE(n10291), .CLK(n10744), 
        .Q(WX3417), .QN(n9456) );
  SDFFX1 DFF_510_Q_reg ( .D(WX3418), .SI(WX3417), .SE(n10290), .CLK(n10745), 
        .Q(WX3419), .QN(n9454) );
  SDFFX1 DFF_511_Q_reg ( .D(WX3420), .SI(WX3419), .SE(n10290), .CLK(n10745), 
        .Q(WX3421), .QN(n9452) );
  SDFFX1 DFF_512_Q_reg ( .D(WX3422), .SI(WX3421), .SE(n10289), .CLK(n10745), 
        .Q(WX3423), .QN(n9701) );
  SDFFX1 DFF_513_Q_reg ( .D(WX3424), .SI(WX3423), .SE(n10289), .CLK(n10745), 
        .Q(WX3425), .QN(n9702) );
  SDFFX1 DFF_514_Q_reg ( .D(WX3426), .SI(WX3425), .SE(n10289), .CLK(n10745), 
        .Q(WX3427), .QN(n9703) );
  SDFFX1 DFF_515_Q_reg ( .D(WX3428), .SI(WX3427), .SE(n10288), .CLK(n10745), 
        .Q(WX3429), .QN(n9704) );
  SDFFX1 DFF_516_Q_reg ( .D(WX3430), .SI(WX3429), .SE(n10288), .CLK(n10746), 
        .Q(WX3431), .QN(n9705) );
  SDFFX1 DFF_517_Q_reg ( .D(WX3432), .SI(WX3431), .SE(n10288), .CLK(n10746), 
        .Q(WX3433), .QN(n9706) );
  SDFFX1 DFF_518_Q_reg ( .D(WX3434), .SI(WX3433), .SE(n10288), .CLK(n10746), 
        .Q(WX3435), .QN(n9707) );
  SDFFX1 DFF_519_Q_reg ( .D(WX3436), .SI(WX3435), .SE(n10288), .CLK(n10746), 
        .Q(WX3437), .QN(n9708) );
  SDFFX1 DFF_520_Q_reg ( .D(WX3438), .SI(WX3437), .SE(n10288), .CLK(n10746), 
        .Q(test_so29), .QN(n9911) );
  SDFFX1 DFF_521_Q_reg ( .D(WX3440), .SI(test_si30), .SE(n10304), .CLK(n10738), 
        .Q(WX3441), .QN(n9709) );
  SDFFX1 DFF_522_Q_reg ( .D(WX3442), .SI(WX3441), .SE(n10303), .CLK(n10738), 
        .Q(WX3443), .QN(n9710) );
  SDFFX1 DFF_523_Q_reg ( .D(WX3444), .SI(WX3443), .SE(n10302), .CLK(n10738), 
        .Q(WX3445), .QN(n9711) );
  SDFFX1 DFF_524_Q_reg ( .D(WX3446), .SI(WX3445), .SE(n10302), .CLK(n10739), 
        .Q(WX3447), .QN(n9712) );
  SDFFX1 DFF_525_Q_reg ( .D(WX3448), .SI(WX3447), .SE(n10301), .CLK(n10739), 
        .Q(WX3449), .QN(n9713) );
  SDFFX1 DFF_526_Q_reg ( .D(WX3450), .SI(WX3449), .SE(n10300), .CLK(n10740), 
        .Q(WX3451), .QN(n9714) );
  SDFFX1 DFF_527_Q_reg ( .D(WX3452), .SI(WX3451), .SE(n10300), .CLK(n10740), 
        .Q(WX3453), .QN(n9527) );
  SDFFX1 DFF_528_Q_reg ( .D(WX3454), .SI(WX3453), .SE(n10299), .CLK(n10740), 
        .Q(WX3455), .QN(n9715) );
  SDFFX1 DFF_529_Q_reg ( .D(WX3456), .SI(WX3455), .SE(n10298), .CLK(n10740), 
        .Q(WX3457), .QN(n9716) );
  SDFFX1 DFF_530_Q_reg ( .D(WX3458), .SI(WX3457), .SE(n10298), .CLK(n10741), 
        .Q(WX3459), .QN(n9717) );
  SDFFX1 DFF_531_Q_reg ( .D(WX3460), .SI(WX3459), .SE(n10297), .CLK(n10741), 
        .Q(WX3461), .QN(n9718) );
  SDFFX1 DFF_532_Q_reg ( .D(WX3462), .SI(WX3461), .SE(n10297), .CLK(n10741), 
        .Q(WX3463), .QN(n9528) );
  SDFFX1 DFF_533_Q_reg ( .D(WX3464), .SI(WX3463), .SE(n10296), .CLK(n10741), 
        .Q(WX3465), .QN(n9719) );
  SDFFX1 DFF_534_Q_reg ( .D(WX3466), .SI(WX3465), .SE(n10295), .CLK(n10742), 
        .Q(WX3467), .QN(n9720) );
  SDFFX1 DFF_535_Q_reg ( .D(WX3468), .SI(WX3467), .SE(n10295), .CLK(n10742), 
        .Q(WX3469), .QN(n9721) );
  SDFFX1 DFF_536_Q_reg ( .D(WX3470), .SI(WX3469), .SE(n10294), .CLK(n10743), 
        .Q(WX3471), .QN(n9722) );
  SDFFX1 DFF_537_Q_reg ( .D(WX3472), .SI(WX3471), .SE(n10293), .CLK(n10743), 
        .Q(test_so30), .QN(n9904) );
  SDFFX1 DFF_538_Q_reg ( .D(WX3474), .SI(test_si31), .SE(n10293), .CLK(n10743), 
        .Q(WX3475), .QN(n9723) );
  SDFFX1 DFF_539_Q_reg ( .D(WX3476), .SI(WX3475), .SE(n10292), .CLK(n10744), 
        .Q(WX3477), .QN(n9529) );
  SDFFX1 DFF_540_Q_reg ( .D(WX3478), .SI(WX3477), .SE(n10291), .CLK(n10744), 
        .Q(WX3479), .QN(n9724) );
  SDFFX1 DFF_541_Q_reg ( .D(WX3480), .SI(WX3479), .SE(n10291), .CLK(n10744), 
        .Q(WX3481), .QN(n9725) );
  SDFFX1 DFF_542_Q_reg ( .D(WX3482), .SI(WX3481), .SE(n10290), .CLK(n10745), 
        .Q(WX3483), .QN(n9726) );
  SDFFX1 DFF_543_Q_reg ( .D(WX3484), .SI(WX3483), .SE(n10289), .CLK(n10745), 
        .Q(WX3485), .QN(n9539) );
  SDFFX1 DFF_544_Q_reg ( .D(WX3850), .SI(WX3485), .SE(n10097), .CLK(n10842), 
        .Q(CRC_OUT_7_0), .QN(DFF_544_n1) );
  SDFFX1 DFF_545_Q_reg ( .D(WX3852), .SI(CRC_OUT_7_0), .SE(n10097), .CLK(
        n10842), .Q(CRC_OUT_7_1), .QN(DFF_545_n1) );
  SDFFX1 DFF_546_Q_reg ( .D(WX3854), .SI(CRC_OUT_7_1), .SE(n10097), .CLK(
        n10842), .Q(CRC_OUT_7_2), .QN(DFF_546_n1) );
  SDFFX1 DFF_547_Q_reg ( .D(WX3856), .SI(CRC_OUT_7_2), .SE(n10097), .CLK(
        n10842), .Q(CRC_OUT_7_3), .QN(DFF_547_n1) );
  SDFFX1 DFF_548_Q_reg ( .D(WX3858), .SI(CRC_OUT_7_3), .SE(n10097), .CLK(
        n10842), .Q(CRC_OUT_7_4), .QN(DFF_548_n1) );
  SDFFX1 DFF_549_Q_reg ( .D(WX3860), .SI(CRC_OUT_7_4), .SE(n10097), .CLK(
        n10842), .Q(CRC_OUT_7_5), .QN(DFF_549_n1) );
  SDFFX1 DFF_550_Q_reg ( .D(WX3862), .SI(CRC_OUT_7_5), .SE(n10096), .CLK(
        n10842), .Q(CRC_OUT_7_6), .QN(DFF_550_n1) );
  SDFFX1 DFF_551_Q_reg ( .D(WX3864), .SI(CRC_OUT_7_6), .SE(n10096), .CLK(
        n10842), .Q(CRC_OUT_7_7), .QN(DFF_551_n1) );
  SDFFX1 DFF_552_Q_reg ( .D(WX3866), .SI(CRC_OUT_7_7), .SE(n10096), .CLK(
        n10842), .Q(CRC_OUT_7_8), .QN(DFF_552_n1) );
  SDFFX1 DFF_553_Q_reg ( .D(WX3868), .SI(CRC_OUT_7_8), .SE(n10096), .CLK(
        n10842), .Q(CRC_OUT_7_9), .QN(DFF_553_n1) );
  SDFFX1 DFF_554_Q_reg ( .D(WX3870), .SI(CRC_OUT_7_9), .SE(n10096), .CLK(
        n10842), .Q(test_so31), .QN(n9889) );
  SDFFX1 DFF_555_Q_reg ( .D(WX3872), .SI(test_si32), .SE(n10096), .CLK(n10842), 
        .Q(CRC_OUT_7_11), .QN(DFF_555_n1) );
  SDFFX1 DFF_556_Q_reg ( .D(WX3874), .SI(CRC_OUT_7_11), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_12), .QN(DFF_556_n1) );
  SDFFX1 DFF_557_Q_reg ( .D(WX3876), .SI(CRC_OUT_7_12), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_13), .QN(DFF_557_n1) );
  SDFFX1 DFF_558_Q_reg ( .D(WX3878), .SI(CRC_OUT_7_13), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_14), .QN(DFF_558_n1) );
  SDFFX1 DFF_559_Q_reg ( .D(WX3880), .SI(CRC_OUT_7_14), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_15), .QN(DFF_559_n1) );
  SDFFX1 DFF_560_Q_reg ( .D(WX3882), .SI(CRC_OUT_7_15), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_16), .QN(DFF_560_n1) );
  SDFFX1 DFF_561_Q_reg ( .D(WX3884), .SI(CRC_OUT_7_16), .SE(n10095), .CLK(
        n10843), .Q(CRC_OUT_7_17), .QN(DFF_561_n1) );
  SDFFX1 DFF_562_Q_reg ( .D(WX3886), .SI(CRC_OUT_7_17), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_18), .QN(DFF_562_n1) );
  SDFFX1 DFF_563_Q_reg ( .D(WX3888), .SI(CRC_OUT_7_18), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_19), .QN(DFF_563_n1) );
  SDFFX1 DFF_564_Q_reg ( .D(WX3890), .SI(CRC_OUT_7_19), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_20), .QN(DFF_564_n1) );
  SDFFX1 DFF_565_Q_reg ( .D(WX3892), .SI(CRC_OUT_7_20), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_21), .QN(DFF_565_n1) );
  SDFFX1 DFF_566_Q_reg ( .D(WX3894), .SI(CRC_OUT_7_21), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_22), .QN(DFF_566_n1) );
  SDFFX1 DFF_567_Q_reg ( .D(WX3896), .SI(CRC_OUT_7_22), .SE(n10094), .CLK(
        n10843), .Q(CRC_OUT_7_23), .QN(DFF_567_n1) );
  SDFFX1 DFF_568_Q_reg ( .D(WX3898), .SI(CRC_OUT_7_23), .SE(n10093), .CLK(
        n10844), .Q(CRC_OUT_7_24), .QN(DFF_568_n1) );
  SDFFX1 DFF_569_Q_reg ( .D(WX3900), .SI(CRC_OUT_7_24), .SE(n10093), .CLK(
        n10844), .Q(CRC_OUT_7_25), .QN(DFF_569_n1) );
  SDFFX1 DFF_570_Q_reg ( .D(WX3902), .SI(CRC_OUT_7_25), .SE(n10093), .CLK(
        n10844), .Q(CRC_OUT_7_26), .QN(DFF_570_n1) );
  SDFFX1 DFF_571_Q_reg ( .D(WX3904), .SI(CRC_OUT_7_26), .SE(n10093), .CLK(
        n10844), .Q(test_so32), .QN(n9945) );
  SDFFX1 DFF_572_Q_reg ( .D(WX3906), .SI(test_si33), .SE(n10093), .CLK(n10844), 
        .Q(CRC_OUT_7_28), .QN(DFF_572_n1) );
  SDFFX1 DFF_573_Q_reg ( .D(WX3908), .SI(CRC_OUT_7_28), .SE(n10093), .CLK(
        n10844), .Q(CRC_OUT_7_29), .QN(DFF_573_n1) );
  SDFFX1 DFF_574_Q_reg ( .D(WX3910), .SI(CRC_OUT_7_29), .SE(n10092), .CLK(
        n10844), .Q(CRC_OUT_7_30), .QN(DFF_574_n1) );
  SDFFX1 DFF_575_Q_reg ( .D(WX3912), .SI(CRC_OUT_7_30), .SE(n10287), .CLK(
        n10746), .Q(CRC_OUT_7_31), .QN(DFF_575_n1) );
  SDFFX1 DFF_576_Q_reg ( .D(n732), .SI(CRC_OUT_7_31), .SE(n10287), .CLK(n10746), .Q(WX4364), .QN(n9846) );
  SDFFX1 DFF_577_Q_reg ( .D(n733), .SI(WX4364), .SE(n10282), .CLK(n10749), .Q(
        n8586), .QN(n3971) );
  SDFFX1 DFF_578_Q_reg ( .D(n734), .SI(n8586), .SE(n10282), .CLK(n10749), .Q(
        n8585), .QN(n3970) );
  SDFFX1 DFF_579_Q_reg ( .D(n735), .SI(n8585), .SE(n10282), .CLK(n10748), .Q(
        n8584), .QN(n3969) );
  SDFFX1 DFF_580_Q_reg ( .D(n736), .SI(n8584), .SE(n10283), .CLK(n10748), .Q(
        n8583), .QN(n3968) );
  SDFFX1 DFF_581_Q_reg ( .D(n737), .SI(n8583), .SE(n10283), .CLK(n10748), .Q(
        n8582), .QN(n3967) );
  SDFFX1 DFF_582_Q_reg ( .D(n738), .SI(n8582), .SE(n10283), .CLK(n10748), .Q(
        n8581), .QN(n3966) );
  SDFFX1 DFF_583_Q_reg ( .D(n739), .SI(n8581), .SE(n10283), .CLK(n10748), .Q(
        n8580), .QN(n3965) );
  SDFFX1 DFF_584_Q_reg ( .D(n740), .SI(n8580), .SE(n10283), .CLK(n10748), .Q(
        n8579), .QN(n3964) );
  SDFFX1 DFF_585_Q_reg ( .D(n741), .SI(n8579), .SE(n10283), .CLK(n10748), .Q(
        n8578), .QN(n3963) );
  SDFFX1 DFF_586_Q_reg ( .D(n742), .SI(n8578), .SE(n10284), .CLK(n10748), .Q(
        n8577), .QN(n3962) );
  SDFFX1 DFF_587_Q_reg ( .D(n743), .SI(n8577), .SE(n10284), .CLK(n10748), .Q(
        n8576), .QN(n3961) );
  SDFFX1 DFF_588_Q_reg ( .D(n744), .SI(n8576), .SE(n10284), .CLK(n10748), .Q(
        test_so33), .QN(n3960) );
  SDFFX1 DFF_589_Q_reg ( .D(n745), .SI(test_si34), .SE(n10284), .CLK(n10748), 
        .Q(n8573), .QN(n3959) );
  SDFFX1 DFF_590_Q_reg ( .D(n746), .SI(n8573), .SE(n10284), .CLK(n10748), .Q(
        n8572), .QN(n3958) );
  SDFFX1 DFF_591_Q_reg ( .D(n747), .SI(n8572), .SE(n10284), .CLK(n10747), .Q(
        n8571), .QN(n3957) );
  SDFFX1 DFF_592_Q_reg ( .D(n748), .SI(n8571), .SE(n10285), .CLK(n10747), .Q(
        n8570), .QN(n3956) );
  SDFFX1 DFF_593_Q_reg ( .D(n749), .SI(n8570), .SE(n10285), .CLK(n10747), .Q(
        n8569), .QN(n3955) );
  SDFFX1 DFF_594_Q_reg ( .D(n750), .SI(n8569), .SE(n10285), .CLK(n10747), .Q(
        n8568), .QN(n3954) );
  SDFFX1 DFF_595_Q_reg ( .D(n751), .SI(n8568), .SE(n10285), .CLK(n10747), .Q(
        n8567), .QN(n3953) );
  SDFFX1 DFF_596_Q_reg ( .D(n752), .SI(n8567), .SE(n10285), .CLK(n10747), .Q(
        n8566), .QN(n3952) );
  SDFFX1 DFF_597_Q_reg ( .D(n753), .SI(n8566), .SE(n10285), .CLK(n10747), .Q(
        n8565), .QN(n3951) );
  SDFFX1 DFF_598_Q_reg ( .D(n754), .SI(n8565), .SE(n10286), .CLK(n10747), .Q(
        n8564), .QN(n3950) );
  SDFFX1 DFF_599_Q_reg ( .D(n755), .SI(n8564), .SE(n10286), .CLK(n10747), .Q(
        n8563), .QN(n3949) );
  SDFFX1 DFF_600_Q_reg ( .D(n756), .SI(n8563), .SE(n10286), .CLK(n10747), .Q(
        n8562), .QN(n3948) );
  SDFFX1 DFF_601_Q_reg ( .D(n757), .SI(n8562), .SE(n10286), .CLK(n10747), .Q(
        n8561), .QN(n3947) );
  SDFFX1 DFF_602_Q_reg ( .D(n758), .SI(n8561), .SE(n10286), .CLK(n10747), .Q(
        n8560), .QN(n3946) );
  SDFFX1 DFF_603_Q_reg ( .D(n759), .SI(n8560), .SE(n10286), .CLK(n10746), .Q(
        n8559), .QN(n3945) );
  SDFFX1 DFF_604_Q_reg ( .D(n760), .SI(n8559), .SE(n10287), .CLK(n10746), .Q(
        n8558), .QN(n3944) );
  SDFFX1 DFF_605_Q_reg ( .D(n761), .SI(n8558), .SE(n10287), .CLK(n10746), .Q(
        test_so34), .QN(n3943) );
  SDFFX1 DFF_606_Q_reg ( .D(n762), .SI(test_si35), .SE(n10287), .CLK(n10746), 
        .Q(n8555), .QN(n3942) );
  SDFFX1 DFF_607_Q_reg ( .D(WX4425), .SI(n8555), .SE(n10287), .CLK(n10746), 
        .Q(n8554), .QN(n3941) );
  SDFFX1 DFF_608_Q_reg ( .D(WX4523), .SI(n8554), .SE(n10098), .CLK(n10841), 
        .Q(n8553), .QN(n17956) );
  SDFFX1 DFF_609_Q_reg ( .D(WX4525), .SI(n8553), .SE(n10282), .CLK(n10749), 
        .Q(n8552), .QN(n17955) );
  SDFFX1 DFF_610_Q_reg ( .D(WX4527), .SI(n8552), .SE(n10281), .CLK(n10749), 
        .Q(n8551), .QN(n17954) );
  SDFFX1 DFF_611_Q_reg ( .D(WX4529), .SI(n8551), .SE(n10281), .CLK(n10749), 
        .Q(n8550), .QN(n17953) );
  SDFFX1 DFF_612_Q_reg ( .D(WX4531), .SI(n8550), .SE(n10280), .CLK(n10750), 
        .Q(n8549), .QN(n17952) );
  SDFFX1 DFF_613_Q_reg ( .D(WX4533), .SI(n8549), .SE(n10280), .CLK(n10750), 
        .Q(n8548), .QN(n17951) );
  SDFFX1 DFF_614_Q_reg ( .D(WX4535), .SI(n8548), .SE(n10279), .CLK(n10750), 
        .Q(n8547), .QN(n17950) );
  SDFFX1 DFF_615_Q_reg ( .D(WX4537), .SI(n8547), .SE(n10279), .CLK(n10750), 
        .Q(n8546), .QN(n17949) );
  SDFFX1 DFF_616_Q_reg ( .D(WX4539), .SI(n8546), .SE(n10277), .CLK(n10751), 
        .Q(n8545), .QN(n17948) );
  SDFFX1 DFF_617_Q_reg ( .D(WX4541), .SI(n8545), .SE(n10277), .CLK(n10751), 
        .Q(n8544), .QN(n17947) );
  SDFFX1 DFF_618_Q_reg ( .D(WX4543), .SI(n8544), .SE(n10276), .CLK(n10752), 
        .Q(n8543), .QN(n17946) );
  SDFFX1 DFF_619_Q_reg ( .D(WX4545), .SI(n8543), .SE(n10276), .CLK(n10752), 
        .Q(n8542), .QN(n17945) );
  SDFFX1 DFF_620_Q_reg ( .D(WX4547), .SI(n8542), .SE(n10275), .CLK(n10752), 
        .Q(n8541), .QN(n17944) );
  SDFFX1 DFF_621_Q_reg ( .D(WX4549), .SI(n8541), .SE(n10275), .CLK(n10752), 
        .Q(n8540), .QN(n17943) );
  SDFFX1 DFF_622_Q_reg ( .D(WX4551), .SI(n8540), .SE(n10098), .CLK(n10841), 
        .Q(test_so35), .QN(n9893) );
  SDFFX1 DFF_623_Q_reg ( .D(WX4553), .SI(test_si36), .SE(n10273), .CLK(n10753), 
        .Q(n8537), .QN(n17942) );
  SDFFX1 DFF_624_Q_reg ( .D(WX4555), .SI(n8537), .SE(n10273), .CLK(n10753), 
        .Q(WX4556), .QN(n9449) );
  SDFFX1 DFF_625_Q_reg ( .D(WX4557), .SI(WX4556), .SE(n10272), .CLK(n10754), 
        .Q(WX4558), .QN(n9447) );
  SDFFX1 DFF_626_Q_reg ( .D(WX4559), .SI(WX4558), .SE(n10271), .CLK(n10754), 
        .Q(WX4560) );
  SDFFX1 DFF_627_Q_reg ( .D(WX4561), .SI(WX4560), .SE(n10271), .CLK(n10754), 
        .Q(WX4562), .QN(n9444) );
  SDFFX1 DFF_628_Q_reg ( .D(WX4563), .SI(WX4562), .SE(n10335), .CLK(n10722), 
        .Q(WX4564) );
  SDFFX1 DFF_629_Q_reg ( .D(WX4565), .SI(WX4564), .SE(n10269), .CLK(n10755), 
        .Q(WX4566), .QN(n9440) );
  SDFFX1 DFF_630_Q_reg ( .D(WX4567), .SI(WX4566), .SE(n10269), .CLK(n10755), 
        .Q(WX4568), .QN(n9438) );
  SDFFX1 DFF_631_Q_reg ( .D(WX4569), .SI(WX4568), .SE(n10268), .CLK(n10756), 
        .Q(WX4570), .QN(n9436) );
  SDFFX1 DFF_632_Q_reg ( .D(WX4571), .SI(WX4570), .SE(n10268), .CLK(n10756), 
        .Q(WX4572), .QN(n9434) );
  SDFFX1 DFF_633_Q_reg ( .D(WX4573), .SI(WX4572), .SE(n10267), .CLK(n10756), 
        .Q(WX4574), .QN(n9432) );
  SDFFX1 DFF_634_Q_reg ( .D(WX4575), .SI(WX4574), .SE(n10266), .CLK(n10757), 
        .Q(WX4576), .QN(n9430) );
  SDFFX1 DFF_635_Q_reg ( .D(WX4577), .SI(WX4576), .SE(n10266), .CLK(n10757), 
        .Q(WX4578), .QN(n9428) );
  SDFFX1 DFF_636_Q_reg ( .D(WX4579), .SI(WX4578), .SE(n10265), .CLK(n10757), 
        .Q(WX4580), .QN(n9426) );
  SDFFX1 DFF_637_Q_reg ( .D(WX4581), .SI(WX4580), .SE(n10264), .CLK(n10758), 
        .Q(WX4582), .QN(n9424) );
  SDFFX1 DFF_638_Q_reg ( .D(WX4583), .SI(WX4582), .SE(n10264), .CLK(n10758), 
        .Q(WX4584), .QN(n9422) );
  SDFFX1 DFF_639_Q_reg ( .D(WX4585), .SI(WX4584), .SE(n10263), .CLK(n10758), 
        .Q(test_so36), .QN(n9926) );
  SDFFX1 DFF_640_Q_reg ( .D(WX4587), .SI(test_si37), .SE(n10098), .CLK(n10841), 
        .Q(WX4588), .QN(n9038) );
  SDFFX1 DFF_641_Q_reg ( .D(WX4589), .SI(WX4588), .SE(n10282), .CLK(n10749), 
        .Q(WX4590), .QN(n9212) );
  SDFFX1 DFF_642_Q_reg ( .D(WX4591), .SI(WX4590), .SE(n10282), .CLK(n10749), 
        .Q(WX4592), .QN(n9210) );
  SDFFX1 DFF_643_Q_reg ( .D(WX4593), .SI(WX4592), .SE(n10281), .CLK(n10749), 
        .Q(WX4594), .QN(n9208) );
  SDFFX1 DFF_644_Q_reg ( .D(WX4595), .SI(WX4594), .SE(n10281), .CLK(n10749), 
        .Q(WX4596), .QN(n9206) );
  SDFFX1 DFF_645_Q_reg ( .D(WX4597), .SI(WX4596), .SE(n10280), .CLK(n10750), 
        .Q(WX4598), .QN(n9204) );
  SDFFX1 DFF_646_Q_reg ( .D(WX4599), .SI(WX4598), .SE(n10279), .CLK(n10750), 
        .Q(WX4600), .QN(n9202) );
  SDFFX1 DFF_647_Q_reg ( .D(WX4601), .SI(WX4600), .SE(n10278), .CLK(n10750), 
        .Q(WX4602), .QN(n9200) );
  SDFFX1 DFF_648_Q_reg ( .D(WX4603), .SI(WX4602), .SE(n10278), .CLK(n10751), 
        .Q(WX4604), .QN(n9198) );
  SDFFX1 DFF_649_Q_reg ( .D(WX4605), .SI(WX4604), .SE(n10277), .CLK(n10751), 
        .Q(WX4606), .QN(n9196) );
  SDFFX1 DFF_650_Q_reg ( .D(WX4607), .SI(WX4606), .SE(n10277), .CLK(n10751), 
        .Q(WX4608), .QN(n9194) );
  SDFFX1 DFF_651_Q_reg ( .D(WX4609), .SI(WX4608), .SE(n10276), .CLK(n10752), 
        .Q(WX4610), .QN(n9192) );
  SDFFX1 DFF_652_Q_reg ( .D(WX4611), .SI(WX4610), .SE(n10275), .CLK(n10752), 
        .Q(WX4612), .QN(n9190) );
  SDFFX1 DFF_653_Q_reg ( .D(WX4613), .SI(WX4612), .SE(n10274), .CLK(n10752), 
        .Q(WX4614), .QN(n9188) );
  SDFFX1 DFF_654_Q_reg ( .D(WX4615), .SI(WX4614), .SE(n10274), .CLK(n10753), 
        .Q(WX4616), .QN(n9186) );
  SDFFX1 DFF_655_Q_reg ( .D(WX4617), .SI(WX4616), .SE(n10273), .CLK(n10753), 
        .Q(WX4618), .QN(n9184) );
  SDFFX1 DFF_656_Q_reg ( .D(WX4619), .SI(WX4618), .SE(n10273), .CLK(n10753), 
        .Q(test_so37), .QN(n9928) );
  SDFFX1 DFF_657_Q_reg ( .D(WX4621), .SI(test_si38), .SE(n10272), .CLK(n10754), 
        .Q(WX4622), .QN(n3719) );
  SDFFX1 DFF_658_Q_reg ( .D(WX4623), .SI(WX4622), .SE(n10271), .CLK(n10754), 
        .Q(WX4624), .QN(n3717) );
  SDFFX1 DFF_659_Q_reg ( .D(WX4625), .SI(WX4624), .SE(n10271), .CLK(n10754), 
        .Q(WX4626), .QN(n3715) );
  SDFFX1 DFF_660_Q_reg ( .D(WX4627), .SI(WX4626), .SE(n10270), .CLK(n10755), 
        .Q(WX4628), .QN(n3713) );
  SDFFX1 DFF_661_Q_reg ( .D(WX4629), .SI(WX4628), .SE(n10270), .CLK(n10755), 
        .Q(WX4630), .QN(n3711) );
  SDFFX1 DFF_662_Q_reg ( .D(WX4631), .SI(WX4630), .SE(n10269), .CLK(n10755), 
        .Q(WX4632), .QN(n3709) );
  SDFFX1 DFF_663_Q_reg ( .D(WX4633), .SI(WX4632), .SE(n10268), .CLK(n10756), 
        .Q(WX4634), .QN(n3707) );
  SDFFX1 DFF_664_Q_reg ( .D(WX4635), .SI(WX4634), .SE(n10267), .CLK(n10756), 
        .Q(WX4636), .QN(n3705) );
  SDFFX1 DFF_665_Q_reg ( .D(WX4637), .SI(WX4636), .SE(n10267), .CLK(n10756), 
        .Q(WX4638), .QN(n3703) );
  SDFFX1 DFF_666_Q_reg ( .D(WX4639), .SI(WX4638), .SE(n10266), .CLK(n10757), 
        .Q(WX4640), .QN(n3701) );
  SDFFX1 DFF_667_Q_reg ( .D(WX4641), .SI(WX4640), .SE(n10265), .CLK(n10757), 
        .Q(WX4642), .QN(n3699) );
  SDFFX1 DFF_668_Q_reg ( .D(WX4643), .SI(WX4642), .SE(n10265), .CLK(n10757), 
        .Q(WX4644), .QN(n3697) );
  SDFFX1 DFF_669_Q_reg ( .D(WX4645), .SI(WX4644), .SE(n10264), .CLK(n10758), 
        .Q(WX4646), .QN(n3695) );
  SDFFX1 DFF_670_Q_reg ( .D(WX4647), .SI(WX4646), .SE(n10263), .CLK(n10758), 
        .Q(WX4648), .QN(n3693) );
  SDFFX1 DFF_671_Q_reg ( .D(WX4649), .SI(WX4648), .SE(n10263), .CLK(n10758), 
        .Q(WX4650), .QN(n3691) );
  SDFFX1 DFF_672_Q_reg ( .D(WX4651), .SI(WX4650), .SE(n10262), .CLK(n10759), 
        .Q(WX4652), .QN(n9039) );
  SDFFX1 DFF_673_Q_reg ( .D(WX4653), .SI(WX4652), .SE(n10262), .CLK(n10759), 
        .Q(test_so38), .QN(n9961) );
  SDFFX1 DFF_674_Q_reg ( .D(WX4655), .SI(test_si39), .SE(n10281), .CLK(n10749), 
        .Q(WX4656), .QN(n9211) );
  SDFFX1 DFF_675_Q_reg ( .D(WX4657), .SI(WX4656), .SE(n10281), .CLK(n10749), 
        .Q(WX4658) );
  SDFFX1 DFF_676_Q_reg ( .D(WX4659), .SI(WX4658), .SE(n10280), .CLK(n10749), 
        .Q(WX4660), .QN(n9207) );
  SDFFX1 DFF_677_Q_reg ( .D(WX4661), .SI(WX4660), .SE(n10280), .CLK(n10750), 
        .Q(WX4662), .QN(n9205) );
  SDFFX1 DFF_678_Q_reg ( .D(WX4663), .SI(WX4662), .SE(n10279), .CLK(n10750), 
        .Q(WX4664), .QN(n9203) );
  SDFFX1 DFF_679_Q_reg ( .D(WX4665), .SI(WX4664), .SE(n10278), .CLK(n10751), 
        .Q(WX4666), .QN(n9201) );
  SDFFX1 DFF_680_Q_reg ( .D(WX4667), .SI(WX4666), .SE(n10278), .CLK(n10751), 
        .Q(WX4668), .QN(n9199) );
  SDFFX1 DFF_681_Q_reg ( .D(WX4669), .SI(WX4668), .SE(n10277), .CLK(n10751), 
        .Q(WX4670), .QN(n9197) );
  SDFFX1 DFF_682_Q_reg ( .D(WX4671), .SI(WX4670), .SE(n10276), .CLK(n10751), 
        .Q(WX4672), .QN(n9195) );
  SDFFX1 DFF_683_Q_reg ( .D(WX4673), .SI(WX4672), .SE(n10276), .CLK(n10752), 
        .Q(WX4674), .QN(n9193) );
  SDFFX1 DFF_684_Q_reg ( .D(WX4675), .SI(WX4674), .SE(n10275), .CLK(n10752), 
        .Q(WX4676), .QN(n9191) );
  SDFFX1 DFF_685_Q_reg ( .D(WX4677), .SI(WX4676), .SE(n10274), .CLK(n10753), 
        .Q(WX4678), .QN(n9189) );
  SDFFX1 DFF_686_Q_reg ( .D(WX4679), .SI(WX4678), .SE(n10274), .CLK(n10753), 
        .Q(WX4680), .QN(n9187) );
  SDFFX1 DFF_687_Q_reg ( .D(WX4681), .SI(WX4680), .SE(n10273), .CLK(n10753), 
        .Q(WX4682), .QN(n9185) );
  SDFFX1 DFF_688_Q_reg ( .D(WX4683), .SI(WX4682), .SE(n10272), .CLK(n10753), 
        .Q(WX4684) );
  SDFFX1 DFF_689_Q_reg ( .D(WX4685), .SI(WX4684), .SE(n10272), .CLK(n10754), 
        .Q(WX4686), .QN(n9448) );
  SDFFX1 DFF_690_Q_reg ( .D(WX4687), .SI(WX4686), .SE(n10271), .CLK(n10754), 
        .Q(test_so39), .QN(n9927) );
  SDFFX1 DFF_691_Q_reg ( .D(WX4689), .SI(test_si40), .SE(n10270), .CLK(n10754), 
        .Q(WX4690), .QN(n9445) );
  SDFFX1 DFF_692_Q_reg ( .D(WX4691), .SI(WX4690), .SE(n10270), .CLK(n10755), 
        .Q(WX4692), .QN(n9443) );
  SDFFX1 DFF_693_Q_reg ( .D(WX4693), .SI(WX4692), .SE(n10269), .CLK(n10755), 
        .Q(WX4694), .QN(n9441) );
  SDFFX1 DFF_694_Q_reg ( .D(WX4695), .SI(WX4694), .SE(n10269), .CLK(n10755), 
        .Q(WX4696), .QN(n9439) );
  SDFFX1 DFF_695_Q_reg ( .D(WX4697), .SI(WX4696), .SE(n10268), .CLK(n10756), 
        .Q(WX4698), .QN(n9437) );
  SDFFX1 DFF_696_Q_reg ( .D(WX4699), .SI(WX4698), .SE(n10267), .CLK(n10756), 
        .Q(WX4700), .QN(n9435) );
  SDFFX1 DFF_697_Q_reg ( .D(WX4701), .SI(WX4700), .SE(n10267), .CLK(n10756), 
        .Q(WX4702), .QN(n9433) );
  SDFFX1 DFF_698_Q_reg ( .D(WX4703), .SI(WX4702), .SE(n10266), .CLK(n10757), 
        .Q(WX4704), .QN(n9431) );
  SDFFX1 DFF_699_Q_reg ( .D(WX4705), .SI(WX4704), .SE(n10265), .CLK(n10757), 
        .Q(WX4706), .QN(n9429) );
  SDFFX1 DFF_700_Q_reg ( .D(WX4707), .SI(WX4706), .SE(n10265), .CLK(n10757), 
        .Q(WX4708), .QN(n9427) );
  SDFFX1 DFF_701_Q_reg ( .D(WX4709), .SI(WX4708), .SE(n10264), .CLK(n10758), 
        .Q(WX4710), .QN(n9425) );
  SDFFX1 DFF_702_Q_reg ( .D(WX4711), .SI(WX4710), .SE(n10263), .CLK(n10758), 
        .Q(WX4712), .QN(n9423) );
  SDFFX1 DFF_703_Q_reg ( .D(WX4713), .SI(WX4712), .SE(n10263), .CLK(n10758), 
        .Q(WX4714) );
  SDFFX1 DFF_704_Q_reg ( .D(WX4715), .SI(WX4714), .SE(n10262), .CLK(n10759), 
        .Q(WX4716), .QN(n9674) );
  SDFFX1 DFF_705_Q_reg ( .D(WX4717), .SI(WX4716), .SE(n10262), .CLK(n10759), 
        .Q(WX4718), .QN(n9675) );
  SDFFX1 DFF_706_Q_reg ( .D(WX4719), .SI(WX4718), .SE(n10262), .CLK(n10759), 
        .Q(WX4720), .QN(n9676) );
  SDFFX1 DFF_707_Q_reg ( .D(WX4721), .SI(WX4720), .SE(n10261), .CLK(n10759), 
        .Q(test_so40), .QN(n9910) );
  SDFFX1 DFF_708_Q_reg ( .D(WX4723), .SI(test_si41), .SE(n10280), .CLK(n10750), 
        .Q(WX4724), .QN(n9677) );
  SDFFX1 DFF_709_Q_reg ( .D(WX4725), .SI(WX4724), .SE(n10279), .CLK(n10750), 
        .Q(WX4726), .QN(n9678) );
  SDFFX1 DFF_710_Q_reg ( .D(WX4727), .SI(WX4726), .SE(n10279), .CLK(n10750), 
        .Q(WX4728), .QN(n9679) );
  SDFFX1 DFF_711_Q_reg ( .D(WX4729), .SI(WX4728), .SE(n10278), .CLK(n10751), 
        .Q(WX4730), .QN(n9680) );
  SDFFX1 DFF_712_Q_reg ( .D(WX4731), .SI(WX4730), .SE(n10278), .CLK(n10751), 
        .Q(WX4732), .QN(n9681) );
  SDFFX1 DFF_713_Q_reg ( .D(WX4733), .SI(WX4732), .SE(n10277), .CLK(n10751), 
        .Q(WX4734), .QN(n9682) );
  SDFFX1 DFF_714_Q_reg ( .D(WX4735), .SI(WX4734), .SE(n10276), .CLK(n10752), 
        .Q(WX4736), .QN(n9683) );
  SDFFX1 DFF_715_Q_reg ( .D(WX4737), .SI(WX4736), .SE(n10275), .CLK(n10752), 
        .Q(WX4738), .QN(n9684) );
  SDFFX1 DFF_716_Q_reg ( .D(WX4739), .SI(WX4738), .SE(n10275), .CLK(n10752), 
        .Q(WX4740), .QN(n9685) );
  SDFFX1 DFF_717_Q_reg ( .D(WX4741), .SI(WX4740), .SE(n10274), .CLK(n10753), 
        .Q(WX4742), .QN(n9686) );
  SDFFX1 DFF_718_Q_reg ( .D(WX4743), .SI(WX4742), .SE(n10274), .CLK(n10753), 
        .Q(WX4744), .QN(n9687) );
  SDFFX1 DFF_719_Q_reg ( .D(WX4745), .SI(WX4744), .SE(n10273), .CLK(n10753), 
        .Q(WX4746), .QN(n9525) );
  SDFFX1 DFF_720_Q_reg ( .D(WX4747), .SI(WX4746), .SE(n10272), .CLK(n10754), 
        .Q(WX4748), .QN(n9688) );
  SDFFX1 DFF_721_Q_reg ( .D(WX4749), .SI(WX4748), .SE(n10272), .CLK(n10754), 
        .Q(WX4750), .QN(n9689) );
  SDFFX1 DFF_722_Q_reg ( .D(WX4751), .SI(WX4750), .SE(n10271), .CLK(n10754), 
        .Q(WX4752), .QN(n9690) );
  SDFFX1 DFF_723_Q_reg ( .D(WX4753), .SI(WX4752), .SE(n10270), .CLK(n10755), 
        .Q(WX4754), .QN(n9691) );
  SDFFX1 DFF_724_Q_reg ( .D(WX4755), .SI(WX4754), .SE(n10270), .CLK(n10755), 
        .Q(test_so41), .QN(n9887) );
  SDFFX1 DFF_725_Q_reg ( .D(WX4757), .SI(test_si42), .SE(n10269), .CLK(n10755), 
        .Q(WX4758), .QN(n9692) );
  SDFFX1 DFF_726_Q_reg ( .D(WX4759), .SI(WX4758), .SE(n10268), .CLK(n10755), 
        .Q(WX4760), .QN(n9693) );
  SDFFX1 DFF_727_Q_reg ( .D(WX4761), .SI(WX4760), .SE(n10268), .CLK(n10756), 
        .Q(WX4762), .QN(n9694) );
  SDFFX1 DFF_728_Q_reg ( .D(WX4763), .SI(WX4762), .SE(n10267), .CLK(n10756), 
        .Q(WX4764), .QN(n9695) );
  SDFFX1 DFF_729_Q_reg ( .D(WX4765), .SI(WX4764), .SE(n10266), .CLK(n10756), 
        .Q(WX4766), .QN(n9696) );
  SDFFX1 DFF_730_Q_reg ( .D(WX4767), .SI(WX4766), .SE(n10266), .CLK(n10757), 
        .Q(WX4768), .QN(n9697) );
  SDFFX1 DFF_731_Q_reg ( .D(WX4769), .SI(WX4768), .SE(n10265), .CLK(n10757), 
        .Q(WX4770), .QN(n9526) );
  SDFFX1 DFF_732_Q_reg ( .D(WX4771), .SI(WX4770), .SE(n10264), .CLK(n10757), 
        .Q(WX4772), .QN(n9698) );
  SDFFX1 DFF_733_Q_reg ( .D(WX4773), .SI(WX4772), .SE(n10264), .CLK(n10758), 
        .Q(WX4774), .QN(n9699) );
  SDFFX1 DFF_734_Q_reg ( .D(WX4775), .SI(WX4774), .SE(n10263), .CLK(n10758), 
        .Q(WX4776), .QN(n9700) );
  SDFFX1 DFF_735_Q_reg ( .D(WX4777), .SI(WX4776), .SE(n10262), .CLK(n10758), 
        .Q(WX4778), .QN(n9538) );
  SDFFX1 DFF_736_Q_reg ( .D(WX5143), .SI(WX4778), .SE(n10103), .CLK(n10839), 
        .Q(CRC_OUT_6_0), .QN(DFF_736_n1) );
  SDFFX1 DFF_737_Q_reg ( .D(WX5145), .SI(CRC_OUT_6_0), .SE(n10103), .CLK(
        n10839), .Q(CRC_OUT_6_1), .QN(DFF_737_n1) );
  SDFFX1 DFF_738_Q_reg ( .D(WX5147), .SI(CRC_OUT_6_1), .SE(n10103), .CLK(
        n10839), .Q(CRC_OUT_6_2), .QN(DFF_738_n1) );
  SDFFX1 DFF_739_Q_reg ( .D(WX5149), .SI(CRC_OUT_6_2), .SE(n10102), .CLK(
        n10839), .Q(CRC_OUT_6_3), .QN(DFF_739_n1) );
  SDFFX1 DFF_740_Q_reg ( .D(WX5151), .SI(CRC_OUT_6_3), .SE(n10102), .CLK(
        n10839), .Q(CRC_OUT_6_4), .QN(DFF_740_n1) );
  SDFFX1 DFF_741_Q_reg ( .D(WX5153), .SI(CRC_OUT_6_4), .SE(n10102), .CLK(
        n10839), .Q(test_so42), .QN(n9944) );
  SDFFX1 DFF_742_Q_reg ( .D(WX5155), .SI(test_si43), .SE(n10102), .CLK(n10839), 
        .Q(CRC_OUT_6_6), .QN(DFF_742_n1) );
  SDFFX1 DFF_743_Q_reg ( .D(WX5157), .SI(CRC_OUT_6_6), .SE(n10102), .CLK(
        n10839), .Q(CRC_OUT_6_7), .QN(DFF_743_n1) );
  SDFFX1 DFF_744_Q_reg ( .D(WX5159), .SI(CRC_OUT_6_7), .SE(n10102), .CLK(
        n10839), .Q(CRC_OUT_6_8), .QN(DFF_744_n1) );
  SDFFX1 DFF_745_Q_reg ( .D(WX5161), .SI(CRC_OUT_6_8), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_9), .QN(DFF_745_n1) );
  SDFFX1 DFF_746_Q_reg ( .D(WX5163), .SI(CRC_OUT_6_9), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_10), .QN(DFF_746_n1) );
  SDFFX1 DFF_747_Q_reg ( .D(WX5165), .SI(CRC_OUT_6_10), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_11), .QN(DFF_747_n1) );
  SDFFX1 DFF_748_Q_reg ( .D(WX5167), .SI(CRC_OUT_6_11), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_12), .QN(DFF_748_n1) );
  SDFFX1 DFF_749_Q_reg ( .D(WX5169), .SI(CRC_OUT_6_12), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_13), .QN(DFF_749_n1) );
  SDFFX1 DFF_750_Q_reg ( .D(WX5171), .SI(CRC_OUT_6_13), .SE(n10101), .CLK(
        n10840), .Q(CRC_OUT_6_14), .QN(DFF_750_n1) );
  SDFFX1 DFF_751_Q_reg ( .D(WX5173), .SI(CRC_OUT_6_14), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_15), .QN(DFF_751_n1) );
  SDFFX1 DFF_752_Q_reg ( .D(WX5175), .SI(CRC_OUT_6_15), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_16), .QN(DFF_752_n1) );
  SDFFX1 DFF_753_Q_reg ( .D(WX5177), .SI(CRC_OUT_6_16), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_17), .QN(DFF_753_n1) );
  SDFFX1 DFF_754_Q_reg ( .D(WX5179), .SI(CRC_OUT_6_17), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_18), .QN(DFF_754_n1) );
  SDFFX1 DFF_755_Q_reg ( .D(WX5181), .SI(CRC_OUT_6_18), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_19), .QN(DFF_755_n1) );
  SDFFX1 DFF_756_Q_reg ( .D(WX5183), .SI(CRC_OUT_6_19), .SE(n10100), .CLK(
        n10840), .Q(CRC_OUT_6_20), .QN(DFF_756_n1) );
  SDFFX1 DFF_757_Q_reg ( .D(WX5185), .SI(CRC_OUT_6_20), .SE(n10099), .CLK(
        n10841), .Q(CRC_OUT_6_21), .QN(DFF_757_n1) );
  SDFFX1 DFF_758_Q_reg ( .D(WX5187), .SI(CRC_OUT_6_21), .SE(n10099), .CLK(
        n10841), .Q(test_so43), .QN(n9943) );
  SDFFX1 DFF_759_Q_reg ( .D(WX5189), .SI(test_si44), .SE(n10099), .CLK(n10841), 
        .Q(CRC_OUT_6_23), .QN(DFF_759_n1) );
  SDFFX1 DFF_760_Q_reg ( .D(WX5191), .SI(CRC_OUT_6_23), .SE(n10099), .CLK(
        n10841), .Q(CRC_OUT_6_24), .QN(DFF_760_n1) );
  SDFFX1 DFF_761_Q_reg ( .D(WX5193), .SI(CRC_OUT_6_24), .SE(n10099), .CLK(
        n10841), .Q(CRC_OUT_6_25), .QN(DFF_761_n1) );
  SDFFX1 DFF_762_Q_reg ( .D(WX5195), .SI(CRC_OUT_6_25), .SE(n10099), .CLK(
        n10841), .Q(CRC_OUT_6_26), .QN(DFF_762_n1) );
  SDFFX1 DFF_763_Q_reg ( .D(WX5197), .SI(CRC_OUT_6_26), .SE(n10098), .CLK(
        n10841), .Q(CRC_OUT_6_27), .QN(DFF_763_n1) );
  SDFFX1 DFF_764_Q_reg ( .D(WX5199), .SI(CRC_OUT_6_27), .SE(n10098), .CLK(
        n10841), .Q(CRC_OUT_6_28), .QN(DFF_764_n1) );
  SDFFX1 DFF_765_Q_reg ( .D(WX5201), .SI(CRC_OUT_6_28), .SE(n10098), .CLK(
        n10841), .Q(CRC_OUT_6_29), .QN(DFF_765_n1) );
  SDFFX1 DFF_766_Q_reg ( .D(WX5203), .SI(CRC_OUT_6_29), .SE(n10261), .CLK(
        n10759), .Q(CRC_OUT_6_30), .QN(DFF_766_n1) );
  SDFFX1 DFF_767_Q_reg ( .D(WX5205), .SI(CRC_OUT_6_30), .SE(n10261), .CLK(
        n10759), .Q(CRC_OUT_6_31), .QN(DFF_767_n1) );
  SDFFX1 DFF_768_Q_reg ( .D(n973), .SI(CRC_OUT_6_31), .SE(n10261), .CLK(n10759), .Q(WX5657), .QN(n9847) );
  SDFFX1 DFF_769_Q_reg ( .D(n974), .SI(WX5657), .SE(n10256), .CLK(n10762), .Q(
        n8528), .QN(n3940) );
  SDFFX1 DFF_770_Q_reg ( .D(n975), .SI(n8528), .SE(n10256), .CLK(n10762), .Q(
        n8527), .QN(n3939) );
  SDFFX1 DFF_771_Q_reg ( .D(n976), .SI(n8527), .SE(n10256), .CLK(n10762), .Q(
        n8526), .QN(n3938) );
  SDFFX1 DFF_772_Q_reg ( .D(n977), .SI(n8526), .SE(n10256), .CLK(n10762), .Q(
        n8525), .QN(n3937) );
  SDFFX1 DFF_773_Q_reg ( .D(n978), .SI(n8525), .SE(n10256), .CLK(n10761), .Q(
        n8524), .QN(n3936) );
  SDFFX1 DFF_774_Q_reg ( .D(n979), .SI(n8524), .SE(n10257), .CLK(n10761), .Q(
        n8523), .QN(n3935) );
  SDFFX1 DFF_775_Q_reg ( .D(n980), .SI(n8523), .SE(n10257), .CLK(n10761), .Q(
        test_so44), .QN(n3934) );
  SDFFX1 DFF_776_Q_reg ( .D(n981), .SI(test_si45), .SE(n10257), .CLK(n10761), 
        .Q(n8520), .QN(n3933) );
  SDFFX1 DFF_777_Q_reg ( .D(n982), .SI(n8520), .SE(n10257), .CLK(n10761), .Q(
        n8519), .QN(n3932) );
  SDFFX1 DFF_778_Q_reg ( .D(n983), .SI(n8519), .SE(n10257), .CLK(n10761), .Q(
        n8518), .QN(n3931) );
  SDFFX1 DFF_779_Q_reg ( .D(n984), .SI(n8518), .SE(n10257), .CLK(n10761), .Q(
        n8517), .QN(n3930) );
  SDFFX1 DFF_780_Q_reg ( .D(n985), .SI(n8517), .SE(n10258), .CLK(n10761), .Q(
        n8516), .QN(n3929) );
  SDFFX1 DFF_781_Q_reg ( .D(n986), .SI(n8516), .SE(n10258), .CLK(n10761), .Q(
        n8515), .QN(n3928) );
  SDFFX1 DFF_782_Q_reg ( .D(n987), .SI(n8515), .SE(n10258), .CLK(n10761), .Q(
        n8514), .QN(n3927) );
  SDFFX1 DFF_783_Q_reg ( .D(n988), .SI(n8514), .SE(n10258), .CLK(n10761), .Q(
        n8513), .QN(n3926) );
  SDFFX1 DFF_784_Q_reg ( .D(n989), .SI(n8513), .SE(n10258), .CLK(n10761), .Q(
        n8512), .QN(n3925) );
  SDFFX1 DFF_785_Q_reg ( .D(n990), .SI(n8512), .SE(n10258), .CLK(n10760), .Q(
        n8511), .QN(n3924) );
  SDFFX1 DFF_786_Q_reg ( .D(n991), .SI(n8511), .SE(n10259), .CLK(n10760), .Q(
        n8510), .QN(n3923) );
  SDFFX1 DFF_787_Q_reg ( .D(n992), .SI(n8510), .SE(n10259), .CLK(n10760), .Q(
        n8509), .QN(n3922) );
  SDFFX1 DFF_788_Q_reg ( .D(n993), .SI(n8509), .SE(n10259), .CLK(n10760), .Q(
        n8508), .QN(n3921) );
  SDFFX1 DFF_789_Q_reg ( .D(n994), .SI(n8508), .SE(n10259), .CLK(n10760), .Q(
        n8507), .QN(n3920) );
  SDFFX1 DFF_790_Q_reg ( .D(n995), .SI(n8507), .SE(n10259), .CLK(n10760), .Q(
        n8506), .QN(n3919) );
  SDFFX1 DFF_791_Q_reg ( .D(n996), .SI(n8506), .SE(n10259), .CLK(n10760), .Q(
        n8505), .QN(n3918) );
  SDFFX1 DFF_792_Q_reg ( .D(n997), .SI(n8505), .SE(n10260), .CLK(n10760), .Q(
        test_so45), .QN(n3917) );
  SDFFX1 DFF_793_Q_reg ( .D(n998), .SI(test_si46), .SE(n10260), .CLK(n10760), 
        .Q(n8502), .QN(n3916) );
  SDFFX1 DFF_794_Q_reg ( .D(n999), .SI(n8502), .SE(n10260), .CLK(n10760), .Q(
        n8501), .QN(n3915) );
  SDFFX1 DFF_795_Q_reg ( .D(n1000), .SI(n8501), .SE(n10260), .CLK(n10760), .Q(
        n8500), .QN(n3914) );
  SDFFX1 DFF_796_Q_reg ( .D(n1001), .SI(n8500), .SE(n10260), .CLK(n10760), .Q(
        n8499), .QN(n3913) );
  SDFFX1 DFF_797_Q_reg ( .D(n1002), .SI(n8499), .SE(n10260), .CLK(n10759), .Q(
        n8498), .QN(n3912) );
  SDFFX1 DFF_798_Q_reg ( .D(n1003), .SI(n8498), .SE(n10261), .CLK(n10759), .Q(
        n8497), .QN(n3911) );
  SDFFX1 DFF_799_Q_reg ( .D(WX5718), .SI(n8497), .SE(n10261), .CLK(n10759), 
        .Q(n8496), .QN(n3910) );
  SDFFX1 DFF_800_Q_reg ( .D(WX5816), .SI(n8496), .SE(n10103), .CLK(n10839), 
        .Q(n8495), .QN(n17941) );
  SDFFX1 DFF_801_Q_reg ( .D(WX5818), .SI(n8495), .SE(n10256), .CLK(n10762), 
        .Q(n8494), .QN(n17940) );
  SDFFX1 DFF_802_Q_reg ( .D(WX5820), .SI(n8494), .SE(n10255), .CLK(n10762), 
        .Q(n8493), .QN(n17939) );
  SDFFX1 DFF_803_Q_reg ( .D(WX5822), .SI(n8493), .SE(n10255), .CLK(n10762), 
        .Q(n8492), .QN(n17938) );
  SDFFX1 DFF_804_Q_reg ( .D(WX5824), .SI(n8492), .SE(n10254), .CLK(n10762), 
        .Q(n8491), .QN(n17937) );
  SDFFX1 DFF_805_Q_reg ( .D(WX5826), .SI(n8491), .SE(n10254), .CLK(n10763), 
        .Q(n8490), .QN(n17936) );
  SDFFX1 DFF_806_Q_reg ( .D(WX5828), .SI(n8490), .SE(n10254), .CLK(n10763), 
        .Q(n8489), .QN(n17935) );
  SDFFX1 DFF_807_Q_reg ( .D(WX5830), .SI(n8489), .SE(n10254), .CLK(n10763), 
        .Q(n8488), .QN(n17934) );
  SDFFX1 DFF_808_Q_reg ( .D(WX5832), .SI(n8488), .SE(n10253), .CLK(n10763), 
        .Q(n8487), .QN(n17933) );
  SDFFX1 DFF_809_Q_reg ( .D(WX5834), .SI(n8487), .SE(n10253), .CLK(n10763), 
        .Q(test_so46), .QN(n9892) );
  SDFFX1 DFF_810_Q_reg ( .D(WX5836), .SI(test_si47), .SE(n10252), .CLK(n10763), 
        .Q(n8484), .QN(n17932) );
  SDFFX1 DFF_811_Q_reg ( .D(WX5838), .SI(n8484), .SE(n10252), .CLK(n10764), 
        .Q(n8483), .QN(n17931) );
  SDFFX1 DFF_812_Q_reg ( .D(WX5840), .SI(n8483), .SE(n10252), .CLK(n10764), 
        .Q(n8482), .QN(n17930) );
  SDFFX1 DFF_813_Q_reg ( .D(WX5842), .SI(n8482), .SE(n10251), .CLK(n10764), 
        .Q(n8481), .QN(n17929) );
  SDFFX1 DFF_814_Q_reg ( .D(WX5844), .SI(n8481), .SE(n10251), .CLK(n10764), 
        .Q(n8480), .QN(n17928) );
  SDFFX1 DFF_815_Q_reg ( .D(WX5846), .SI(n8480), .SE(n10250), .CLK(n10765), 
        .Q(n8479), .QN(n17927) );
  SDFFX1 DFF_816_Q_reg ( .D(WX5848), .SI(n8479), .SE(n10250), .CLK(n10765), 
        .Q(WX5849), .QN(n9419) );
  SDFFX1 DFF_817_Q_reg ( .D(WX5850), .SI(WX5849), .SE(n10249), .CLK(n10765), 
        .Q(WX5851), .QN(n9417) );
  SDFFX1 DFF_818_Q_reg ( .D(WX5852), .SI(WX5851), .SE(n10248), .CLK(n10765), 
        .Q(WX5853), .QN(n9415) );
  SDFFX1 DFF_819_Q_reg ( .D(WX5854), .SI(WX5853), .SE(n10248), .CLK(n10766), 
        .Q(WX5855), .QN(n9413) );
  SDFFX1 DFF_820_Q_reg ( .D(WX5856), .SI(WX5855), .SE(n10336), .CLK(n10722), 
        .Q(WX5857), .QN(n9411) );
  SDFFX1 DFF_821_Q_reg ( .D(WX5858), .SI(WX5857), .SE(n10246), .CLK(n10767), 
        .Q(WX5859), .QN(n9409) );
  SDFFX1 DFF_822_Q_reg ( .D(WX5860), .SI(WX5859), .SE(n10246), .CLK(n10767), 
        .Q(WX5861), .QN(n9407) );
  SDFFX1 DFF_823_Q_reg ( .D(WX5862), .SI(WX5861), .SE(n10245), .CLK(n10767), 
        .Q(WX5863), .QN(n9405) );
  SDFFX1 DFF_824_Q_reg ( .D(WX5864), .SI(WX5863), .SE(n10245), .CLK(n10767), 
        .Q(WX5865), .QN(n9403) );
  SDFFX1 DFF_825_Q_reg ( .D(WX5866), .SI(WX5865), .SE(n10244), .CLK(n10768), 
        .Q(WX5867), .QN(n9401) );
  SDFFX1 DFF_826_Q_reg ( .D(WX5868), .SI(WX5867), .SE(n10243), .CLK(n10768), 
        .Q(test_so47), .QN(n9925) );
  SDFFX1 DFF_827_Q_reg ( .D(WX5870), .SI(test_si48), .SE(n10242), .CLK(n10769), 
        .Q(WX5871), .QN(n9398) );
  SDFFX1 DFF_828_Q_reg ( .D(WX5872), .SI(WX5871), .SE(n10242), .CLK(n10769), 
        .Q(WX5873), .QN(n9396) );
  SDFFX1 DFF_829_Q_reg ( .D(WX5874), .SI(WX5873), .SE(n10241), .CLK(n10769), 
        .Q(WX5875), .QN(n9394) );
  SDFFX1 DFF_830_Q_reg ( .D(WX5876), .SI(WX5875), .SE(n10241), .CLK(n10769), 
        .Q(WX5877) );
  SDFFX1 DFF_831_Q_reg ( .D(WX5878), .SI(WX5877), .SE(n10240), .CLK(n10770), 
        .Q(WX5879), .QN(n9391) );
  SDFFX1 DFF_832_Q_reg ( .D(WX5880), .SI(WX5879), .SE(n10239), .CLK(n10770), 
        .Q(WX5881), .QN(n9036) );
  SDFFX1 DFF_833_Q_reg ( .D(WX5882), .SI(WX5881), .SE(n10255), .CLK(n10762), 
        .Q(WX5883), .QN(n9182) );
  SDFFX1 DFF_834_Q_reg ( .D(WX5884), .SI(WX5883), .SE(n10255), .CLK(n10762), 
        .Q(WX5885), .QN(n9180) );
  SDFFX1 DFF_835_Q_reg ( .D(WX5886), .SI(WX5885), .SE(n10255), .CLK(n10762), 
        .Q(WX5887), .QN(n9178) );
  SDFFX1 DFF_836_Q_reg ( .D(WX5888), .SI(WX5887), .SE(n10255), .CLK(n10762), 
        .Q(WX5889), .QN(n9176) );
  SDFFX1 DFF_837_Q_reg ( .D(WX5890), .SI(WX5889), .SE(n10254), .CLK(n10763), 
        .Q(WX5891), .QN(n9174) );
  SDFFX1 DFF_838_Q_reg ( .D(WX5892), .SI(WX5891), .SE(n10254), .CLK(n10763), 
        .Q(WX5893), .QN(n9172) );
  SDFFX1 DFF_839_Q_reg ( .D(WX5894), .SI(WX5893), .SE(n10253), .CLK(n10763), 
        .Q(WX5895), .QN(n9170) );
  SDFFX1 DFF_840_Q_reg ( .D(WX5896), .SI(WX5895), .SE(n10253), .CLK(n10763), 
        .Q(WX5897), .QN(n9168) );
  SDFFX1 DFF_841_Q_reg ( .D(WX5898), .SI(WX5897), .SE(n10253), .CLK(n10763), 
        .Q(WX5899), .QN(n9166) );
  SDFFX1 DFF_842_Q_reg ( .D(WX5900), .SI(WX5899), .SE(n10253), .CLK(n10763), 
        .Q(WX5901), .QN(n9164) );
  SDFFX1 DFF_843_Q_reg ( .D(WX5902), .SI(WX5901), .SE(n10252), .CLK(n10764), 
        .Q(test_so48), .QN(n9960) );
  SDFFX1 DFF_844_Q_reg ( .D(WX5904), .SI(test_si49), .SE(n10251), .CLK(n10764), 
        .Q(WX5905), .QN(n9161) );
  SDFFX1 DFF_845_Q_reg ( .D(WX5906), .SI(WX5905), .SE(n10251), .CLK(n10764), 
        .Q(WX5907), .QN(n9160) );
  SDFFX1 DFF_846_Q_reg ( .D(WX5908), .SI(WX5907), .SE(n10251), .CLK(n10764), 
        .Q(WX5909), .QN(n9158) );
  SDFFX1 DFF_847_Q_reg ( .D(WX5910), .SI(WX5909), .SE(n10250), .CLK(n10765), 
        .Q(WX5911), .QN(n9156) );
  SDFFX1 DFF_848_Q_reg ( .D(WX5912), .SI(WX5911), .SE(n10250), .CLK(n10765), 
        .Q(WX5913), .QN(n3689) );
  SDFFX1 DFF_849_Q_reg ( .D(WX5914), .SI(WX5913), .SE(n10249), .CLK(n10765), 
        .Q(WX5915), .QN(n3687) );
  SDFFX1 DFF_850_Q_reg ( .D(WX5916), .SI(WX5915), .SE(n10248), .CLK(n10766), 
        .Q(WX5917), .QN(n3685) );
  SDFFX1 DFF_851_Q_reg ( .D(WX5918), .SI(WX5917), .SE(n10248), .CLK(n10766), 
        .Q(WX5919), .QN(n3683) );
  SDFFX1 DFF_852_Q_reg ( .D(WX5920), .SI(WX5919), .SE(n10247), .CLK(n10766), 
        .Q(WX5921), .QN(n3681) );
  SDFFX1 DFF_853_Q_reg ( .D(WX5922), .SI(WX5921), .SE(n10247), .CLK(n10766), 
        .Q(WX5923), .QN(n3679) );
  SDFFX1 DFF_854_Q_reg ( .D(WX5924), .SI(WX5923), .SE(n10246), .CLK(n10767), 
        .Q(WX5925), .QN(n3677) );
  SDFFX1 DFF_855_Q_reg ( .D(WX5926), .SI(WX5925), .SE(n10245), .CLK(n10767), 
        .Q(WX5927), .QN(n3675) );
  SDFFX1 DFF_856_Q_reg ( .D(WX5928), .SI(WX5927), .SE(n10244), .CLK(n10767), 
        .Q(WX5929), .QN(n3673) );
  SDFFX1 DFF_857_Q_reg ( .D(WX5930), .SI(WX5929), .SE(n10244), .CLK(n10768), 
        .Q(WX5931), .QN(n3671) );
  SDFFX1 DFF_858_Q_reg ( .D(WX5932), .SI(WX5931), .SE(n10243), .CLK(n10768), 
        .Q(WX5933), .QN(n3669) );
  SDFFX1 DFF_859_Q_reg ( .D(WX5934), .SI(WX5933), .SE(n10243), .CLK(n10768), 
        .Q(WX5935), .QN(n3667) );
  SDFFX1 DFF_860_Q_reg ( .D(WX5936), .SI(WX5935), .SE(n10242), .CLK(n10769), 
        .Q(test_so49), .QN(n9924) );
  SDFFX1 DFF_861_Q_reg ( .D(WX5938), .SI(test_si50), .SE(n10241), .CLK(n10769), 
        .Q(WX5939), .QN(n3663) );
  SDFFX1 DFF_862_Q_reg ( .D(WX5940), .SI(WX5939), .SE(n10240), .CLK(n10769), 
        .Q(WX5941), .QN(n3661) );
  SDFFX1 DFF_863_Q_reg ( .D(WX5942), .SI(WX5941), .SE(n10240), .CLK(n10770), 
        .Q(WX5943), .QN(n3659) );
  SDFFX1 DFF_864_Q_reg ( .D(WX5944), .SI(WX5943), .SE(n10239), .CLK(n10770), 
        .Q(WX5945), .QN(n9037) );
  SDFFX1 DFF_865_Q_reg ( .D(WX5946), .SI(WX5945), .SE(n10239), .CLK(n10770), 
        .Q(WX5947), .QN(n9183) );
  SDFFX1 DFF_866_Q_reg ( .D(WX5948), .SI(WX5947), .SE(n10238), .CLK(n10770), 
        .Q(WX5949), .QN(n9181) );
  SDFFX1 DFF_867_Q_reg ( .D(WX5950), .SI(WX5949), .SE(n10238), .CLK(n10771), 
        .Q(WX5951), .QN(n9179) );
  SDFFX1 DFF_868_Q_reg ( .D(WX5952), .SI(WX5951), .SE(n10238), .CLK(n10771), 
        .Q(WX5953), .QN(n9177) );
  SDFFX1 DFF_869_Q_reg ( .D(WX5954), .SI(WX5953), .SE(n10237), .CLK(n10771), 
        .Q(WX5955), .QN(n9175) );
  SDFFX1 DFF_870_Q_reg ( .D(WX5956), .SI(WX5955), .SE(n10237), .CLK(n10771), 
        .Q(WX5957), .QN(n9173) );
  SDFFX1 DFF_871_Q_reg ( .D(WX5958), .SI(WX5957), .SE(n10237), .CLK(n10771), 
        .Q(WX5959), .QN(n9171) );
  SDFFX1 DFF_872_Q_reg ( .D(WX5960), .SI(WX5959), .SE(n10236), .CLK(n10771), 
        .Q(WX5961), .QN(n9169) );
  SDFFX1 DFF_873_Q_reg ( .D(WX5962), .SI(WX5961), .SE(n10236), .CLK(n10772), 
        .Q(WX5963), .QN(n9167) );
  SDFFX1 DFF_874_Q_reg ( .D(WX5964), .SI(WX5963), .SE(n10236), .CLK(n10772), 
        .Q(WX5965), .QN(n9165) );
  SDFFX1 DFF_875_Q_reg ( .D(WX5966), .SI(WX5965), .SE(n10252), .CLK(n10764), 
        .Q(WX5967), .QN(n9163) );
  SDFFX1 DFF_876_Q_reg ( .D(WX5968), .SI(WX5967), .SE(n10252), .CLK(n10764), 
        .Q(WX5969), .QN(n9162) );
  SDFFX1 DFF_877_Q_reg ( .D(WX5970), .SI(WX5969), .SE(n10251), .CLK(n10764), 
        .Q(test_so50), .QN(n9959) );
  SDFFX1 DFF_878_Q_reg ( .D(WX5972), .SI(test_si51), .SE(n10250), .CLK(n10764), 
        .Q(WX5973), .QN(n9159) );
  SDFFX1 DFF_879_Q_reg ( .D(WX5974), .SI(WX5973), .SE(n10250), .CLK(n10765), 
        .Q(WX5975) );
  SDFFX1 DFF_880_Q_reg ( .D(WX5976), .SI(WX5975), .SE(n10249), .CLK(n10765), 
        .Q(WX5977), .QN(n9420) );
  SDFFX1 DFF_881_Q_reg ( .D(WX5978), .SI(WX5977), .SE(n10249), .CLK(n10765), 
        .Q(WX5979), .QN(n9418) );
  SDFFX1 DFF_882_Q_reg ( .D(WX5980), .SI(WX5979), .SE(n10248), .CLK(n10766), 
        .Q(WX5981), .QN(n9416) );
  SDFFX1 DFF_883_Q_reg ( .D(WX5982), .SI(WX5981), .SE(n10247), .CLK(n10766), 
        .Q(WX5983), .QN(n9414) );
  SDFFX1 DFF_884_Q_reg ( .D(WX5984), .SI(WX5983), .SE(n10247), .CLK(n10766), 
        .Q(WX5985), .QN(n9412) );
  SDFFX1 DFF_885_Q_reg ( .D(WX5986), .SI(WX5985), .SE(n10246), .CLK(n10766), 
        .Q(WX5987), .QN(n9410) );
  SDFFX1 DFF_886_Q_reg ( .D(WX5988), .SI(WX5987), .SE(n10246), .CLK(n10767), 
        .Q(WX5989), .QN(n9408) );
  SDFFX1 DFF_887_Q_reg ( .D(WX5990), .SI(WX5989), .SE(n10245), .CLK(n10767), 
        .Q(WX5991), .QN(n9406) );
  SDFFX1 DFF_888_Q_reg ( .D(WX5992), .SI(WX5991), .SE(n10244), .CLK(n10768), 
        .Q(WX5993), .QN(n9404) );
  SDFFX1 DFF_889_Q_reg ( .D(WX5994), .SI(WX5993), .SE(n10244), .CLK(n10768), 
        .Q(WX5995), .QN(n9402) );
  SDFFX1 DFF_890_Q_reg ( .D(WX5996), .SI(WX5995), .SE(n10243), .CLK(n10768), 
        .Q(WX5997) );
  SDFFX1 DFF_891_Q_reg ( .D(WX5998), .SI(WX5997), .SE(n10242), .CLK(n10768), 
        .Q(WX5999), .QN(n9399) );
  SDFFX1 DFF_892_Q_reg ( .D(WX6000), .SI(WX5999), .SE(n10242), .CLK(n10769), 
        .Q(WX6001) );
  SDFFX1 DFF_893_Q_reg ( .D(WX6002), .SI(WX6001), .SE(n10241), .CLK(n10769), 
        .Q(WX6003), .QN(n9395) );
  SDFFX1 DFF_894_Q_reg ( .D(WX6004), .SI(WX6003), .SE(n10240), .CLK(n10770), 
        .Q(test_so51), .QN(n9923) );
  SDFFX1 DFF_895_Q_reg ( .D(WX6006), .SI(test_si52), .SE(n10240), .CLK(n10770), 
        .Q(WX6007), .QN(n9392) );
  SDFFX1 DFF_896_Q_reg ( .D(WX6008), .SI(WX6007), .SE(n10239), .CLK(n10770), 
        .Q(WX6009), .QN(n9646) );
  SDFFX1 DFF_897_Q_reg ( .D(WX6010), .SI(WX6009), .SE(n10239), .CLK(n10770), 
        .Q(WX6011), .QN(n9647) );
  SDFFX1 DFF_898_Q_reg ( .D(WX6012), .SI(WX6011), .SE(n10238), .CLK(n10771), 
        .Q(WX6013), .QN(n9648) );
  SDFFX1 DFF_899_Q_reg ( .D(WX6014), .SI(WX6013), .SE(n10238), .CLK(n10771), 
        .Q(WX6015), .QN(n9649) );
  SDFFX1 DFF_900_Q_reg ( .D(WX6016), .SI(WX6015), .SE(n10238), .CLK(n10771), 
        .Q(WX6017), .QN(n9650) );
  SDFFX1 DFF_901_Q_reg ( .D(WX6018), .SI(WX6017), .SE(n10237), .CLK(n10771), 
        .Q(WX6019), .QN(n9651) );
  SDFFX1 DFF_902_Q_reg ( .D(WX6020), .SI(WX6019), .SE(n10237), .CLK(n10771), 
        .Q(WX6021), .QN(n9652) );
  SDFFX1 DFF_903_Q_reg ( .D(WX6022), .SI(WX6021), .SE(n10237), .CLK(n10771), 
        .Q(WX6023), .QN(n9653) );
  SDFFX1 DFF_904_Q_reg ( .D(WX6024), .SI(WX6023), .SE(n10236), .CLK(n10772), 
        .Q(WX6025), .QN(n9654) );
  SDFFX1 DFF_905_Q_reg ( .D(WX6026), .SI(WX6025), .SE(n10236), .CLK(n10772), 
        .Q(WX6027), .QN(n9655) );
  SDFFX1 DFF_906_Q_reg ( .D(WX6028), .SI(WX6027), .SE(n10236), .CLK(n10772), 
        .Q(WX6029), .QN(n9656) );
  SDFFX1 DFF_907_Q_reg ( .D(WX6030), .SI(WX6029), .SE(n10235), .CLK(n10772), 
        .Q(WX6031), .QN(n9657) );
  SDFFX1 DFF_908_Q_reg ( .D(WX6032), .SI(WX6031), .SE(n10235), .CLK(n10772), 
        .Q(WX6033), .QN(n9658) );
  SDFFX1 DFF_909_Q_reg ( .D(WX6034), .SI(WX6033), .SE(n10235), .CLK(n10772), 
        .Q(WX6035), .QN(n9659) );
  SDFFX1 DFF_910_Q_reg ( .D(WX6036), .SI(WX6035), .SE(n10235), .CLK(n10772), 
        .Q(WX6037), .QN(n9660) );
  SDFFX1 DFF_911_Q_reg ( .D(WX6038), .SI(WX6037), .SE(n10235), .CLK(n10772), 
        .Q(test_so52), .QN(n9888) );
  SDFFX1 DFF_912_Q_reg ( .D(WX6040), .SI(test_si53), .SE(n10249), .CLK(n10765), 
        .Q(WX6041), .QN(n9661) );
  SDFFX1 DFF_913_Q_reg ( .D(WX6042), .SI(WX6041), .SE(n10249), .CLK(n10765), 
        .Q(WX6043), .QN(n9662) );
  SDFFX1 DFF_914_Q_reg ( .D(WX6044), .SI(WX6043), .SE(n10248), .CLK(n10766), 
        .Q(WX6045), .QN(n9663) );
  SDFFX1 DFF_915_Q_reg ( .D(WX6046), .SI(WX6045), .SE(n10247), .CLK(n10766), 
        .Q(WX6047), .QN(n9664) );
  SDFFX1 DFF_916_Q_reg ( .D(WX6048), .SI(WX6047), .SE(n10247), .CLK(n10766), 
        .Q(WX6049), .QN(n9523) );
  SDFFX1 DFF_917_Q_reg ( .D(WX6050), .SI(WX6049), .SE(n10246), .CLK(n10767), 
        .Q(WX6051), .QN(n9665) );
  SDFFX1 DFF_918_Q_reg ( .D(WX6052), .SI(WX6051), .SE(n10245), .CLK(n10767), 
        .Q(WX6053), .QN(n9666) );
  SDFFX1 DFF_919_Q_reg ( .D(WX6054), .SI(WX6053), .SE(n10245), .CLK(n10767), 
        .Q(WX6055), .QN(n9667) );
  SDFFX1 DFF_920_Q_reg ( .D(WX6056), .SI(WX6055), .SE(n10244), .CLK(n10768), 
        .Q(WX6057), .QN(n9668) );
  SDFFX1 DFF_921_Q_reg ( .D(WX6058), .SI(WX6057), .SE(n10243), .CLK(n10768), 
        .Q(WX6059), .QN(n9669) );
  SDFFX1 DFF_922_Q_reg ( .D(WX6060), .SI(WX6059), .SE(n10243), .CLK(n10768), 
        .Q(WX6061), .QN(n9670) );
  SDFFX1 DFF_923_Q_reg ( .D(WX6062), .SI(WX6061), .SE(n10242), .CLK(n10769), 
        .Q(WX6063), .QN(n9524) );
  SDFFX1 DFF_924_Q_reg ( .D(WX6064), .SI(WX6063), .SE(n10241), .CLK(n10769), 
        .Q(WX6065), .QN(n9671) );
  SDFFX1 DFF_925_Q_reg ( .D(WX6066), .SI(WX6065), .SE(n10241), .CLK(n10769), 
        .Q(WX6067), .QN(n9672) );
  SDFFX1 DFF_926_Q_reg ( .D(WX6068), .SI(WX6067), .SE(n10240), .CLK(n10770), 
        .Q(WX6069), .QN(n9673) );
  SDFFX1 DFF_927_Q_reg ( .D(WX6070), .SI(WX6069), .SE(n10239), .CLK(n10770), 
        .Q(WX6071), .QN(n9537) );
  SDFFX1 DFF_928_Q_reg ( .D(WX6436), .SI(WX6071), .SE(n10107), .CLK(n10837), 
        .Q(test_so53), .QN(n9942) );
  SDFFX1 DFF_929_Q_reg ( .D(WX6438), .SI(test_si54), .SE(n10106), .CLK(n10837), 
        .Q(CRC_OUT_5_1), .QN(DFF_929_n1) );
  SDFFX1 DFF_930_Q_reg ( .D(WX6440), .SI(CRC_OUT_5_1), .SE(n10106), .CLK(
        n10837), .Q(CRC_OUT_5_2), .QN(DFF_930_n1) );
  SDFFX1 DFF_931_Q_reg ( .D(WX6442), .SI(CRC_OUT_5_2), .SE(n10106), .CLK(
        n10837), .Q(CRC_OUT_5_3), .QN(DFF_931_n1) );
  SDFFX1 DFF_932_Q_reg ( .D(WX6444), .SI(CRC_OUT_5_3), .SE(n10106), .CLK(
        n10837), .Q(CRC_OUT_5_4), .QN(DFF_932_n1) );
  SDFFX1 DFF_933_Q_reg ( .D(WX6446), .SI(CRC_OUT_5_4), .SE(n10106), .CLK(
        n10837), .Q(CRC_OUT_5_5), .QN(DFF_933_n1) );
  SDFFX1 DFF_934_Q_reg ( .D(WX6448), .SI(CRC_OUT_5_5), .SE(n10106), .CLK(
        n10837), .Q(CRC_OUT_5_6), .QN(DFF_934_n1) );
  SDFFX1 DFF_935_Q_reg ( .D(WX6450), .SI(CRC_OUT_5_6), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_7), .QN(DFF_935_n1) );
  SDFFX1 DFF_936_Q_reg ( .D(WX6452), .SI(CRC_OUT_5_7), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_8), .QN(DFF_936_n1) );
  SDFFX1 DFF_937_Q_reg ( .D(WX6454), .SI(CRC_OUT_5_8), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_9), .QN(DFF_937_n1) );
  SDFFX1 DFF_938_Q_reg ( .D(WX6456), .SI(CRC_OUT_5_9), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_10), .QN(DFF_938_n1) );
  SDFFX1 DFF_939_Q_reg ( .D(WX6458), .SI(CRC_OUT_5_10), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_11), .QN(DFF_939_n1) );
  SDFFX1 DFF_940_Q_reg ( .D(WX6460), .SI(CRC_OUT_5_11), .SE(n10105), .CLK(
        n10838), .Q(CRC_OUT_5_12), .QN(DFF_940_n1) );
  SDFFX1 DFF_941_Q_reg ( .D(WX6462), .SI(CRC_OUT_5_12), .SE(n10104), .CLK(
        n10838), .Q(CRC_OUT_5_13), .QN(DFF_941_n1) );
  SDFFX1 DFF_942_Q_reg ( .D(WX6464), .SI(CRC_OUT_5_13), .SE(n10104), .CLK(
        n10838), .Q(CRC_OUT_5_14), .QN(DFF_942_n1) );
  SDFFX1 DFF_943_Q_reg ( .D(WX6466), .SI(CRC_OUT_5_14), .SE(n10104), .CLK(
        n10838), .Q(CRC_OUT_5_15), .QN(DFF_943_n1) );
  SDFFX1 DFF_944_Q_reg ( .D(WX6468), .SI(CRC_OUT_5_15), .SE(n10104), .CLK(
        n10838), .Q(CRC_OUT_5_16), .QN(DFF_944_n1) );
  SDFFX1 DFF_945_Q_reg ( .D(WX6470), .SI(CRC_OUT_5_16), .SE(n10104), .CLK(
        n10838), .Q(test_so54), .QN(n9941) );
  SDFFX1 DFF_946_Q_reg ( .D(WX6472), .SI(test_si55), .SE(n10104), .CLK(n10838), 
        .Q(CRC_OUT_5_18), .QN(DFF_946_n1) );
  SDFFX1 DFF_947_Q_reg ( .D(WX6474), .SI(CRC_OUT_5_18), .SE(n10103), .CLK(
        n10839), .Q(CRC_OUT_5_19), .QN(DFF_947_n1) );
  SDFFX1 DFF_948_Q_reg ( .D(WX6476), .SI(CRC_OUT_5_19), .SE(n10103), .CLK(
        n10839), .Q(CRC_OUT_5_20), .QN(DFF_948_n1) );
  SDFFX1 DFF_949_Q_reg ( .D(WX6478), .SI(CRC_OUT_5_20), .SE(n10235), .CLK(
        n10772), .Q(CRC_OUT_5_21), .QN(DFF_949_n1) );
  SDFFX1 DFF_950_Q_reg ( .D(WX6480), .SI(CRC_OUT_5_21), .SE(n10234), .CLK(
        n10772), .Q(CRC_OUT_5_22), .QN(DFF_950_n1) );
  SDFFX1 DFF_951_Q_reg ( .D(WX6482), .SI(CRC_OUT_5_22), .SE(n10234), .CLK(
        n10773), .Q(CRC_OUT_5_23), .QN(DFF_951_n1) );
  SDFFX1 DFF_952_Q_reg ( .D(WX6484), .SI(CRC_OUT_5_23), .SE(n10234), .CLK(
        n10773), .Q(CRC_OUT_5_24), .QN(DFF_952_n1) );
  SDFFX1 DFF_953_Q_reg ( .D(WX6486), .SI(CRC_OUT_5_24), .SE(n10234), .CLK(
        n10773), .Q(CRC_OUT_5_25), .QN(DFF_953_n1) );
  SDFFX1 DFF_954_Q_reg ( .D(WX6488), .SI(CRC_OUT_5_25), .SE(n10234), .CLK(
        n10773), .Q(CRC_OUT_5_26), .QN(DFF_954_n1) );
  SDFFX1 DFF_955_Q_reg ( .D(WX6490), .SI(CRC_OUT_5_26), .SE(n10234), .CLK(
        n10773), .Q(CRC_OUT_5_27), .QN(DFF_955_n1) );
  SDFFX1 DFF_956_Q_reg ( .D(WX6492), .SI(CRC_OUT_5_27), .SE(n10233), .CLK(
        n10773), .Q(CRC_OUT_5_28), .QN(DFF_956_n1) );
  SDFFX1 DFF_957_Q_reg ( .D(WX6494), .SI(CRC_OUT_5_28), .SE(n10233), .CLK(
        n10773), .Q(CRC_OUT_5_29), .QN(DFF_957_n1) );
  SDFFX1 DFF_958_Q_reg ( .D(WX6496), .SI(CRC_OUT_5_29), .SE(n10233), .CLK(
        n10773), .Q(CRC_OUT_5_30), .QN(DFF_958_n1) );
  SDFFX1 DFF_959_Q_reg ( .D(WX6498), .SI(CRC_OUT_5_30), .SE(n10233), .CLK(
        n10773), .Q(CRC_OUT_5_31), .QN(DFF_959_n1) );
  SDFFX1 DFF_960_Q_reg ( .D(n1214), .SI(CRC_OUT_5_31), .SE(n10233), .CLK(
        n10773), .Q(WX6950), .QN(n9848) );
  SDFFX1 DFF_961_Q_reg ( .D(n1215), .SI(WX6950), .SE(n10228), .CLK(n10776), 
        .Q(n8470), .QN(n3909) );
  SDFFX1 DFF_962_Q_reg ( .D(n1216), .SI(n8470), .SE(n10228), .CLK(n10776), .Q(
        test_so55), .QN(n3908) );
  SDFFX1 DFF_963_Q_reg ( .D(n1217), .SI(test_si56), .SE(n10228), .CLK(n10776), 
        .Q(n8467), .QN(n3907) );
  SDFFX1 DFF_964_Q_reg ( .D(n1218), .SI(n8467), .SE(n10228), .CLK(n10776), .Q(
        n8466), .QN(n3906) );
  SDFFX1 DFF_965_Q_reg ( .D(n1219), .SI(n8466), .SE(n10228), .CLK(n10776), .Q(
        n8465), .QN(n3905) );
  SDFFX1 DFF_966_Q_reg ( .D(n1220), .SI(n8465), .SE(n10228), .CLK(n10775), .Q(
        n8464), .QN(n3904) );
  SDFFX1 DFF_967_Q_reg ( .D(n1221), .SI(n8464), .SE(n10229), .CLK(n10775), .Q(
        n8463), .QN(n3903) );
  SDFFX1 DFF_968_Q_reg ( .D(n1222), .SI(n8463), .SE(n10229), .CLK(n10775), .Q(
        n8462), .QN(n3902) );
  SDFFX1 DFF_969_Q_reg ( .D(n1223), .SI(n8462), .SE(n10229), .CLK(n10775), .Q(
        n8461), .QN(n3901) );
  SDFFX1 DFF_970_Q_reg ( .D(n1224), .SI(n8461), .SE(n10229), .CLK(n10775), .Q(
        n8460), .QN(n3900) );
  SDFFX1 DFF_971_Q_reg ( .D(n1225), .SI(n8460), .SE(n10229), .CLK(n10775), .Q(
        n8459), .QN(n3899) );
  SDFFX1 DFF_972_Q_reg ( .D(n1226), .SI(n8459), .SE(n10229), .CLK(n10775), .Q(
        n8458), .QN(n3898) );
  SDFFX1 DFF_973_Q_reg ( .D(n1227), .SI(n8458), .SE(n10230), .CLK(n10775), .Q(
        n8457), .QN(n3897) );
  SDFFX1 DFF_974_Q_reg ( .D(n1228), .SI(n8457), .SE(n10230), .CLK(n10775), .Q(
        n8456), .QN(n3896) );
  SDFFX1 DFF_975_Q_reg ( .D(n1229), .SI(n8456), .SE(n10230), .CLK(n10775), .Q(
        n8455), .QN(n3895) );
  SDFFX1 DFF_976_Q_reg ( .D(n1230), .SI(n8455), .SE(n10230), .CLK(n10775), .Q(
        n8454), .QN(n3894) );
  SDFFX1 DFF_977_Q_reg ( .D(n1231), .SI(n8454), .SE(n10230), .CLK(n10775), .Q(
        n8453), .QN(n3893) );
  SDFFX1 DFF_978_Q_reg ( .D(n1232), .SI(n8453), .SE(n10230), .CLK(n10774), .Q(
        n8452), .QN(n3892) );
  SDFFX1 DFF_979_Q_reg ( .D(n1233), .SI(n8452), .SE(n10231), .CLK(n10774), .Q(
        test_so56), .QN(n3891) );
  SDFFX1 DFF_980_Q_reg ( .D(n1234), .SI(test_si57), .SE(n10231), .CLK(n10774), 
        .Q(n8449), .QN(n3890) );
  SDFFX1 DFF_981_Q_reg ( .D(n1235), .SI(n8449), .SE(n10231), .CLK(n10774), .Q(
        n8448), .QN(n3889) );
  SDFFX1 DFF_982_Q_reg ( .D(n1236), .SI(n8448), .SE(n10231), .CLK(n10774), .Q(
        n8447), .QN(n3888) );
  SDFFX1 DFF_983_Q_reg ( .D(n1237), .SI(n8447), .SE(n10231), .CLK(n10774), .Q(
        n8446), .QN(n3887) );
  SDFFX1 DFF_984_Q_reg ( .D(n1238), .SI(n8446), .SE(n10231), .CLK(n10774), .Q(
        n8445), .QN(n3886) );
  SDFFX1 DFF_985_Q_reg ( .D(n1239), .SI(n8445), .SE(n10232), .CLK(n10774), .Q(
        n8444), .QN(n3885) );
  SDFFX1 DFF_986_Q_reg ( .D(n1240), .SI(n8444), .SE(n10232), .CLK(n10774), .Q(
        n8443), .QN(n3884) );
  SDFFX1 DFF_987_Q_reg ( .D(n1241), .SI(n8443), .SE(n10232), .CLK(n10774), .Q(
        n8442), .QN(n3883) );
  SDFFX1 DFF_988_Q_reg ( .D(n1242), .SI(n8442), .SE(n10232), .CLK(n10774), .Q(
        n8441), .QN(n3882) );
  SDFFX1 DFF_989_Q_reg ( .D(n1243), .SI(n8441), .SE(n10232), .CLK(n10774), .Q(
        n8440), .QN(n3881) );
  SDFFX1 DFF_990_Q_reg ( .D(n1244), .SI(n8440), .SE(n10232), .CLK(n10773), .Q(
        n8439), .QN(n3880) );
  SDFFX1 DFF_991_Q_reg ( .D(WX7011), .SI(n8439), .SE(n10233), .CLK(n10773), 
        .Q(n8438), .QN(n3879) );
  SDFFX1 DFF_992_Q_reg ( .D(WX7109), .SI(n8438), .SE(n10107), .CLK(n10837), 
        .Q(n8437), .QN(n17926) );
  SDFFX1 DFF_993_Q_reg ( .D(WX7111), .SI(n8437), .SE(n10227), .CLK(n10776), 
        .Q(n8436), .QN(n17925) );
  SDFFX1 DFF_994_Q_reg ( .D(WX7113), .SI(n8436), .SE(n10227), .CLK(n10776), 
        .Q(n8435), .QN(n17924) );
  SDFFX1 DFF_995_Q_reg ( .D(WX7115), .SI(n8435), .SE(n10227), .CLK(n10776), 
        .Q(n8434), .QN(n17923) );
  SDFFX1 DFF_996_Q_reg ( .D(WX7117), .SI(n8434), .SE(n10107), .CLK(n10837), 
        .Q(test_so57), .QN(n9891) );
  SDFFX1 DFF_997_Q_reg ( .D(WX7119), .SI(test_si58), .SE(n10226), .CLK(n10777), 
        .Q(n8431), .QN(n17922) );
  SDFFX1 DFF_998_Q_reg ( .D(WX7121), .SI(n8431), .SE(n10226), .CLK(n10777), 
        .Q(n8430), .QN(n17921) );
  SDFFX1 DFF_999_Q_reg ( .D(WX7123), .SI(n8430), .SE(n10225), .CLK(n10777), 
        .Q(n8429), .QN(n17920) );
  SDFFX1 DFF_1000_Q_reg ( .D(WX7125), .SI(n8429), .SE(n10225), .CLK(n10777), 
        .Q(n8428), .QN(n17919) );
  SDFFX1 DFF_1001_Q_reg ( .D(WX7127), .SI(n8428), .SE(n10224), .CLK(n10777), 
        .Q(n8427), .QN(n17918) );
  SDFFX1 DFF_1002_Q_reg ( .D(WX7129), .SI(n8427), .SE(n10224), .CLK(n10778), 
        .Q(n8426), .QN(n17917) );
  SDFFX1 DFF_1003_Q_reg ( .D(WX7131), .SI(n8426), .SE(n10223), .CLK(n10778), 
        .Q(n8425), .QN(n17916) );
  SDFFX1 DFF_1004_Q_reg ( .D(WX7133), .SI(n8425), .SE(n10222), .CLK(n10779), 
        .Q(n8424), .QN(n17915) );
  SDFFX1 DFF_1005_Q_reg ( .D(WX7135), .SI(n8424), .SE(n10222), .CLK(n10779), 
        .Q(n8423), .QN(n17914) );
  SDFFX1 DFF_1006_Q_reg ( .D(WX7137), .SI(n8423), .SE(n10221), .CLK(n10779), 
        .Q(n8422), .QN(n17913) );
  SDFFX1 DFF_1007_Q_reg ( .D(WX7139), .SI(n8422), .SE(n10221), .CLK(n10779), 
        .Q(n8421), .QN(n17912) );
  SDFFX1 DFF_1008_Q_reg ( .D(WX7141), .SI(n8421), .SE(n10220), .CLK(n10780), 
        .Q(WX7142), .QN(n9389) );
  SDFFX1 DFF_1009_Q_reg ( .D(WX7143), .SI(WX7142), .SE(n10219), .CLK(n10780), 
        .Q(WX7144), .QN(n9387) );
  SDFFX1 DFF_1010_Q_reg ( .D(WX7145), .SI(WX7144), .SE(n10219), .CLK(n10780), 
        .Q(WX7146), .QN(n9385) );
  SDFFX1 DFF_1011_Q_reg ( .D(WX7147), .SI(WX7146), .SE(n10218), .CLK(n10781), 
        .Q(WX7148), .QN(n9383) );
  SDFFX1 DFF_1012_Q_reg ( .D(WX7149), .SI(WX7148), .SE(n10336), .CLK(n10722), 
        .Q(WX7150), .QN(n9381) );
  SDFFX1 DFF_1013_Q_reg ( .D(WX7151), .SI(WX7150), .SE(n10107), .CLK(n10837), 
        .Q(test_so58), .QN(n9922) );
  SDFFX1 DFF_1014_Q_reg ( .D(WX7153), .SI(test_si59), .SE(n10216), .CLK(n10782), .Q(WX7154), .QN(n9378) );
  SDFFX1 DFF_1015_Q_reg ( .D(WX7155), .SI(WX7154), .SE(n10216), .CLK(n10782), 
        .Q(WX7156), .QN(n9376) );
  SDFFX1 DFF_1016_Q_reg ( .D(WX7157), .SI(WX7156), .SE(n10215), .CLK(n10782), 
        .Q(WX7158), .QN(n9374) );
  SDFFX1 DFF_1017_Q_reg ( .D(WX7159), .SI(WX7158), .SE(n10214), .CLK(n10782), 
        .Q(WX7160) );
  SDFFX1 DFF_1018_Q_reg ( .D(WX7161), .SI(WX7160), .SE(n10214), .CLK(n10783), 
        .Q(WX7162), .QN(n9371) );
  SDFFX1 DFF_1019_Q_reg ( .D(WX7163), .SI(WX7162), .SE(n10213), .CLK(n10783), 
        .Q(WX7164) );
  SDFFX1 DFF_1020_Q_reg ( .D(WX7165), .SI(WX7164), .SE(n10212), .CLK(n10783), 
        .Q(WX7166), .QN(n9367) );
  SDFFX1 DFF_1021_Q_reg ( .D(WX7167), .SI(WX7166), .SE(n10212), .CLK(n10784), 
        .Q(WX7168), .QN(n9365) );
  SDFFX1 DFF_1022_Q_reg ( .D(WX7169), .SI(WX7168), .SE(n10211), .CLK(n10784), 
        .Q(WX7170), .QN(n9363) );
  SDFFX1 DFF_1023_Q_reg ( .D(WX7171), .SI(WX7170), .SE(n10210), .CLK(n10784), 
        .Q(WX7172), .QN(n9361) );
  SDFFX1 DFF_1024_Q_reg ( .D(WX7173), .SI(WX7172), .SE(n10210), .CLK(n10785), 
        .Q(WX7174), .QN(n9034) );
  SDFFX1 DFF_1025_Q_reg ( .D(WX7175), .SI(WX7174), .SE(n10227), .CLK(n10776), 
        .Q(WX7176), .QN(n9154) );
  SDFFX1 DFF_1026_Q_reg ( .D(WX7177), .SI(WX7176), .SE(n10227), .CLK(n10776), 
        .Q(WX7178), .QN(n9152) );
  SDFFX1 DFF_1027_Q_reg ( .D(WX7179), .SI(WX7178), .SE(n10227), .CLK(n10776), 
        .Q(WX7180), .QN(n9150) );
  SDFFX1 DFF_1028_Q_reg ( .D(WX7181), .SI(WX7180), .SE(n10226), .CLK(n10776), 
        .Q(WX7182), .QN(n9148) );
  SDFFX1 DFF_1029_Q_reg ( .D(WX7183), .SI(WX7182), .SE(n10226), .CLK(n10777), 
        .Q(WX7184), .QN(n9146) );
  SDFFX1 DFF_1030_Q_reg ( .D(WX7185), .SI(WX7184), .SE(n10226), .CLK(n10777), 
        .Q(test_so59), .QN(n9958) );
  SDFFX1 DFF_1031_Q_reg ( .D(WX7187), .SI(test_si60), .SE(n10225), .CLK(n10777), .Q(WX7188), .QN(n9143) );
  SDFFX1 DFF_1032_Q_reg ( .D(WX7189), .SI(WX7188), .SE(n10225), .CLK(n10777), 
        .Q(WX7190), .QN(n9142) );
  SDFFX1 DFF_1033_Q_reg ( .D(WX7191), .SI(WX7190), .SE(n10224), .CLK(n10778), 
        .Q(WX7192), .QN(n9140) );
  SDFFX1 DFF_1034_Q_reg ( .D(WX7193), .SI(WX7192), .SE(n10224), .CLK(n10778), 
        .Q(WX7194), .QN(n9138) );
  SDFFX1 DFF_1035_Q_reg ( .D(WX7195), .SI(WX7194), .SE(n10223), .CLK(n10778), 
        .Q(WX7196), .QN(n9136) );
  SDFFX1 DFF_1036_Q_reg ( .D(WX7197), .SI(WX7196), .SE(n10223), .CLK(n10778), 
        .Q(WX7198), .QN(n9134) );
  SDFFX1 DFF_1037_Q_reg ( .D(WX7199), .SI(WX7198), .SE(n10222), .CLK(n10779), 
        .Q(WX7200), .QN(n9132) );
  SDFFX1 DFF_1038_Q_reg ( .D(WX7201), .SI(WX7200), .SE(n10221), .CLK(n10779), 
        .Q(WX7202), .QN(n9130) );
  SDFFX1 DFF_1039_Q_reg ( .D(WX7203), .SI(WX7202), .SE(n10221), .CLK(n10779), 
        .Q(WX7204), .QN(n9128) );
  SDFFX1 DFF_1040_Q_reg ( .D(WX7205), .SI(WX7204), .SE(n10220), .CLK(n10780), 
        .Q(WX7206), .QN(n3657) );
  SDFFX1 DFF_1041_Q_reg ( .D(WX7207), .SI(WX7206), .SE(n10219), .CLK(n10780), 
        .Q(WX7208), .QN(n3655) );
  SDFFX1 DFF_1042_Q_reg ( .D(WX7209), .SI(WX7208), .SE(n10219), .CLK(n10780), 
        .Q(WX7210), .QN(n3653) );
  SDFFX1 DFF_1043_Q_reg ( .D(WX7211), .SI(WX7210), .SE(n10218), .CLK(n10781), 
        .Q(WX7212), .QN(n3651) );
  SDFFX1 DFF_1044_Q_reg ( .D(WX7213), .SI(WX7212), .SE(n10217), .CLK(n10781), 
        .Q(WX7214), .QN(n3649) );
  SDFFX1 DFF_1045_Q_reg ( .D(WX7215), .SI(WX7214), .SE(n10217), .CLK(n10781), 
        .Q(WX7216), .QN(n3647) );
  SDFFX1 DFF_1046_Q_reg ( .D(WX7217), .SI(WX7216), .SE(n10216), .CLK(n10781), 
        .Q(WX7218), .QN(n3645) );
  SDFFX1 DFF_1047_Q_reg ( .D(WX7219), .SI(WX7218), .SE(n10216), .CLK(n10782), 
        .Q(test_so60), .QN(n9921) );
  SDFFX1 DFF_1048_Q_reg ( .D(WX7221), .SI(test_si61), .SE(n10215), .CLK(n10782), .Q(WX7222), .QN(n3641) );
  SDFFX1 DFF_1049_Q_reg ( .D(WX7223), .SI(WX7222), .SE(n10214), .CLK(n10783), 
        .Q(WX7224), .QN(n3639) );
  SDFFX1 DFF_1050_Q_reg ( .D(WX7225), .SI(WX7224), .SE(n10214), .CLK(n10783), 
        .Q(WX7226), .QN(n3637) );
  SDFFX1 DFF_1051_Q_reg ( .D(WX7227), .SI(WX7226), .SE(n10213), .CLK(n10783), 
        .Q(WX7228), .QN(n3635) );
  SDFFX1 DFF_1052_Q_reg ( .D(WX7229), .SI(WX7228), .SE(n10212), .CLK(n10784), 
        .Q(WX7230), .QN(n3633) );
  SDFFX1 DFF_1053_Q_reg ( .D(WX7231), .SI(WX7230), .SE(n10212), .CLK(n10784), 
        .Q(WX7232), .QN(n3631) );
  SDFFX1 DFF_1054_Q_reg ( .D(WX7233), .SI(WX7232), .SE(n10211), .CLK(n10784), 
        .Q(WX7234), .QN(n3629) );
  SDFFX1 DFF_1055_Q_reg ( .D(WX7235), .SI(WX7234), .SE(n10210), .CLK(n10785), 
        .Q(WX7236), .QN(n3627) );
  SDFFX1 DFF_1056_Q_reg ( .D(WX7237), .SI(WX7236), .SE(n10210), .CLK(n10785), 
        .Q(WX7238), .QN(n9035) );
  SDFFX1 DFF_1057_Q_reg ( .D(WX7239), .SI(WX7238), .SE(n10209), .CLK(n10785), 
        .Q(WX7240), .QN(n9155) );
  SDFFX1 DFF_1058_Q_reg ( .D(WX7241), .SI(WX7240), .SE(n10209), .CLK(n10785), 
        .Q(WX7242), .QN(n9153) );
  SDFFX1 DFF_1059_Q_reg ( .D(WX7243), .SI(WX7242), .SE(n10209), .CLK(n10785), 
        .Q(WX7244), .QN(n9151) );
  SDFFX1 DFF_1060_Q_reg ( .D(WX7245), .SI(WX7244), .SE(n10208), .CLK(n10786), 
        .Q(WX7246), .QN(n9149) );
  SDFFX1 DFF_1061_Q_reg ( .D(WX7247), .SI(WX7246), .SE(n10208), .CLK(n10786), 
        .Q(WX7248), .QN(n9147) );
  SDFFX1 DFF_1062_Q_reg ( .D(WX7249), .SI(WX7248), .SE(n10226), .CLK(n10777), 
        .Q(WX7250), .QN(n9145) );
  SDFFX1 DFF_1063_Q_reg ( .D(WX7251), .SI(WX7250), .SE(n10225), .CLK(n10777), 
        .Q(WX7252), .QN(n9144) );
  SDFFX1 DFF_1064_Q_reg ( .D(WX7253), .SI(WX7252), .SE(n10225), .CLK(n10777), 
        .Q(test_so61), .QN(n9957) );
  SDFFX1 DFF_1065_Q_reg ( .D(WX7255), .SI(test_si62), .SE(n10224), .CLK(n10778), .Q(WX7256), .QN(n9141) );
  SDFFX1 DFF_1066_Q_reg ( .D(WX7257), .SI(WX7256), .SE(n10224), .CLK(n10778), 
        .Q(WX7258) );
  SDFFX1 DFF_1067_Q_reg ( .D(WX7259), .SI(WX7258), .SE(n10223), .CLK(n10778), 
        .Q(WX7260), .QN(n9137) );
  SDFFX1 DFF_1068_Q_reg ( .D(WX7261), .SI(WX7260), .SE(n10223), .CLK(n10778), 
        .Q(WX7262), .QN(n9135) );
  SDFFX1 DFF_1069_Q_reg ( .D(WX7263), .SI(WX7262), .SE(n10222), .CLK(n10779), 
        .Q(WX7264), .QN(n9133) );
  SDFFX1 DFF_1070_Q_reg ( .D(WX7265), .SI(WX7264), .SE(n10221), .CLK(n10779), 
        .Q(WX7266), .QN(n9131) );
  SDFFX1 DFF_1071_Q_reg ( .D(WX7267), .SI(WX7266), .SE(n10220), .CLK(n10779), 
        .Q(WX7268), .QN(n9129) );
  SDFFX1 DFF_1072_Q_reg ( .D(WX7269), .SI(WX7268), .SE(n10220), .CLK(n10780), 
        .Q(WX7270), .QN(n9390) );
  SDFFX1 DFF_1073_Q_reg ( .D(WX7271), .SI(WX7270), .SE(n10219), .CLK(n10780), 
        .Q(WX7272), .QN(n9388) );
  SDFFX1 DFF_1074_Q_reg ( .D(WX7273), .SI(WX7272), .SE(n10218), .CLK(n10780), 
        .Q(WX7274), .QN(n9386) );
  SDFFX1 DFF_1075_Q_reg ( .D(WX7275), .SI(WX7274), .SE(n10218), .CLK(n10781), 
        .Q(WX7276), .QN(n9384) );
  SDFFX1 DFF_1076_Q_reg ( .D(WX7277), .SI(WX7276), .SE(n10217), .CLK(n10781), 
        .Q(WX7278), .QN(n9382) );
  SDFFX1 DFF_1077_Q_reg ( .D(WX7279), .SI(WX7278), .SE(n10217), .CLK(n10781), 
        .Q(WX7280) );
  SDFFX1 DFF_1078_Q_reg ( .D(WX7281), .SI(WX7280), .SE(n10216), .CLK(n10782), 
        .Q(WX7282), .QN(n9379) );
  SDFFX1 DFF_1079_Q_reg ( .D(WX7283), .SI(WX7282), .SE(n10215), .CLK(n10782), 
        .Q(WX7284) );
  SDFFX1 DFF_1080_Q_reg ( .D(WX7285), .SI(WX7284), .SE(n10215), .CLK(n10782), 
        .Q(WX7286), .QN(n9375) );
  SDFFX1 DFF_1081_Q_reg ( .D(WX7287), .SI(WX7286), .SE(n10214), .CLK(n10783), 
        .Q(test_so62), .QN(n9920) );
  SDFFX1 DFF_1082_Q_reg ( .D(WX7289), .SI(test_si63), .SE(n10213), .CLK(n10783), .Q(WX7290), .QN(n9372) );
  SDFFX1 DFF_1083_Q_reg ( .D(WX7291), .SI(WX7290), .SE(n10213), .CLK(n10783), 
        .Q(WX7292), .QN(n9370) );
  SDFFX1 DFF_1084_Q_reg ( .D(WX7293), .SI(WX7292), .SE(n10212), .CLK(n10784), 
        .Q(WX7294), .QN(n9368) );
  SDFFX1 DFF_1085_Q_reg ( .D(WX7295), .SI(WX7294), .SE(n10211), .CLK(n10784), 
        .Q(WX7296), .QN(n9366) );
  SDFFX1 DFF_1086_Q_reg ( .D(WX7297), .SI(WX7296), .SE(n10211), .CLK(n10784), 
        .Q(WX7298), .QN(n9364) );
  SDFFX1 DFF_1087_Q_reg ( .D(WX7299), .SI(WX7298), .SE(n10210), .CLK(n10785), 
        .Q(WX7300), .QN(n9362) );
  SDFFX1 DFF_1088_Q_reg ( .D(WX7301), .SI(WX7300), .SE(n10209), .CLK(n10785), 
        .Q(WX7302), .QN(n9619) );
  SDFFX1 DFF_1089_Q_reg ( .D(WX7303), .SI(WX7302), .SE(n10209), .CLK(n10785), 
        .Q(WX7304), .QN(n9620) );
  SDFFX1 DFF_1090_Q_reg ( .D(WX7305), .SI(WX7304), .SE(n10209), .CLK(n10785), 
        .Q(WX7306), .QN(n9621) );
  SDFFX1 DFF_1091_Q_reg ( .D(WX7307), .SI(WX7306), .SE(n10208), .CLK(n10785), 
        .Q(WX7308), .QN(n9622) );
  SDFFX1 DFF_1092_Q_reg ( .D(WX7309), .SI(WX7308), .SE(n10208), .CLK(n10786), 
        .Q(WX7310), .QN(n9623) );
  SDFFX1 DFF_1093_Q_reg ( .D(WX7311), .SI(WX7310), .SE(n10208), .CLK(n10786), 
        .Q(WX7312), .QN(n9624) );
  SDFFX1 DFF_1094_Q_reg ( .D(WX7313), .SI(WX7312), .SE(n10208), .CLK(n10786), 
        .Q(WX7314), .QN(n9625) );
  SDFFX1 DFF_1095_Q_reg ( .D(WX7315), .SI(WX7314), .SE(n10207), .CLK(n10786), 
        .Q(WX7316), .QN(n9626) );
  SDFFX1 DFF_1096_Q_reg ( .D(WX7317), .SI(WX7316), .SE(n10207), .CLK(n10786), 
        .Q(WX7318), .QN(n9627) );
  SDFFX1 DFF_1097_Q_reg ( .D(WX7319), .SI(WX7318), .SE(n10207), .CLK(n10786), 
        .Q(WX7320), .QN(n9628) );
  SDFFX1 DFF_1098_Q_reg ( .D(WX7321), .SI(WX7320), .SE(n10207), .CLK(n10786), 
        .Q(test_so63), .QN(n9909) );
  SDFFX1 DFF_1099_Q_reg ( .D(WX7323), .SI(test_si64), .SE(n10223), .CLK(n10778), .Q(WX7324), .QN(n9629) );
  SDFFX1 DFF_1100_Q_reg ( .D(WX7325), .SI(WX7324), .SE(n10222), .CLK(n10778), 
        .Q(WX7326), .QN(n9630) );
  SDFFX1 DFF_1101_Q_reg ( .D(WX7327), .SI(WX7326), .SE(n10222), .CLK(n10779), 
        .Q(WX7328), .QN(n9631) );
  SDFFX1 DFF_1102_Q_reg ( .D(WX7329), .SI(WX7328), .SE(n10221), .CLK(n10779), 
        .Q(WX7330), .QN(n9632) );
  SDFFX1 DFF_1103_Q_reg ( .D(WX7331), .SI(WX7330), .SE(n10220), .CLK(n10780), 
        .Q(WX7332), .QN(n9521) );
  SDFFX1 DFF_1104_Q_reg ( .D(WX7333), .SI(WX7332), .SE(n10220), .CLK(n10780), 
        .Q(WX7334), .QN(n9633) );
  SDFFX1 DFF_1105_Q_reg ( .D(WX7335), .SI(WX7334), .SE(n10219), .CLK(n10780), 
        .Q(WX7336), .QN(n9634) );
  SDFFX1 DFF_1106_Q_reg ( .D(WX7337), .SI(WX7336), .SE(n10218), .CLK(n10781), 
        .Q(WX7338), .QN(n9635) );
  SDFFX1 DFF_1107_Q_reg ( .D(WX7339), .SI(WX7338), .SE(n10218), .CLK(n10781), 
        .Q(WX7340), .QN(n9636) );
  SDFFX1 DFF_1108_Q_reg ( .D(WX7341), .SI(WX7340), .SE(n10217), .CLK(n10781), 
        .Q(WX7342), .QN(n9522) );
  SDFFX1 DFF_1109_Q_reg ( .D(WX7343), .SI(WX7342), .SE(n10217), .CLK(n10781), 
        .Q(WX7344), .QN(n9637) );
  SDFFX1 DFF_1110_Q_reg ( .D(WX7345), .SI(WX7344), .SE(n10216), .CLK(n10782), 
        .Q(WX7346), .QN(n9638) );
  SDFFX1 DFF_1111_Q_reg ( .D(WX7347), .SI(WX7346), .SE(n10215), .CLK(n10782), 
        .Q(WX7348), .QN(n9639) );
  SDFFX1 DFF_1112_Q_reg ( .D(WX7349), .SI(WX7348), .SE(n10215), .CLK(n10782), 
        .Q(WX7350), .QN(n9640) );
  SDFFX1 DFF_1113_Q_reg ( .D(WX7351), .SI(WX7350), .SE(n10214), .CLK(n10783), 
        .Q(WX7352), .QN(n9641) );
  SDFFX1 DFF_1114_Q_reg ( .D(WX7353), .SI(WX7352), .SE(n10213), .CLK(n10783), 
        .Q(WX7354), .QN(n9642) );
  SDFFX1 DFF_1115_Q_reg ( .D(WX7355), .SI(WX7354), .SE(n10213), .CLK(n10783), 
        .Q(test_so64), .QN(n9886) );
  SDFFX1 DFF_1116_Q_reg ( .D(WX7357), .SI(test_si65), .SE(n10212), .CLK(n10784), .Q(WX7358), .QN(n9643) );
  SDFFX1 DFF_1117_Q_reg ( .D(WX7359), .SI(WX7358), .SE(n10211), .CLK(n10784), 
        .Q(WX7360), .QN(n9644) );
  SDFFX1 DFF_1118_Q_reg ( .D(WX7361), .SI(WX7360), .SE(n10211), .CLK(n10784), 
        .Q(WX7362), .QN(n9645) );
  SDFFX1 DFF_1119_Q_reg ( .D(WX7363), .SI(WX7362), .SE(n10210), .CLK(n10785), 
        .Q(WX7364), .QN(n9536) );
  SDFFX1 DFF_1120_Q_reg ( .D(WX7729), .SI(WX7364), .SE(n10111), .CLK(n10835), 
        .Q(CRC_OUT_4_0), .QN(DFF_1120_n1) );
  SDFFX1 DFF_1121_Q_reg ( .D(WX7731), .SI(CRC_OUT_4_0), .SE(n10111), .CLK(
        n10835), .Q(CRC_OUT_4_1), .QN(DFF_1121_n1) );
  SDFFX1 DFF_1122_Q_reg ( .D(WX7733), .SI(CRC_OUT_4_1), .SE(n10111), .CLK(
        n10835), .Q(CRC_OUT_4_2), .QN(DFF_1122_n1) );
  SDFFX1 DFF_1123_Q_reg ( .D(WX7735), .SI(CRC_OUT_4_2), .SE(n10111), .CLK(
        n10835), .Q(CRC_OUT_4_3), .QN(DFF_1123_n1) );
  SDFFX1 DFF_1124_Q_reg ( .D(WX7737), .SI(CRC_OUT_4_3), .SE(n10111), .CLK(
        n10835), .Q(CRC_OUT_4_4), .QN(DFF_1124_n1) );
  SDFFX1 DFF_1125_Q_reg ( .D(WX7739), .SI(CRC_OUT_4_4), .SE(n10111), .CLK(
        n10835), .Q(CRC_OUT_4_5), .QN(DFF_1125_n1) );
  SDFFX1 DFF_1126_Q_reg ( .D(WX7741), .SI(CRC_OUT_4_5), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_6), .QN(DFF_1126_n1) );
  SDFFX1 DFF_1127_Q_reg ( .D(WX7743), .SI(CRC_OUT_4_6), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_7), .QN(DFF_1127_n1) );
  SDFFX1 DFF_1128_Q_reg ( .D(WX7745), .SI(CRC_OUT_4_7), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_8), .QN(DFF_1128_n1) );
  SDFFX1 DFF_1129_Q_reg ( .D(WX7747), .SI(CRC_OUT_4_8), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_9), .QN(DFF_1129_n1) );
  SDFFX1 DFF_1130_Q_reg ( .D(WX7749), .SI(CRC_OUT_4_9), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_10), .QN(DFF_1130_n1) );
  SDFFX1 DFF_1131_Q_reg ( .D(WX7751), .SI(CRC_OUT_4_10), .SE(n10110), .CLK(
        n10835), .Q(CRC_OUT_4_11), .QN(DFF_1131_n1) );
  SDFFX1 DFF_1132_Q_reg ( .D(WX7753), .SI(CRC_OUT_4_11), .SE(n10109), .CLK(
        n10836), .Q(test_so65), .QN(n9940) );
  SDFFX1 DFF_1133_Q_reg ( .D(WX7755), .SI(test_si66), .SE(n10109), .CLK(n10836), .Q(CRC_OUT_4_13), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1134_Q_reg ( .D(WX7757), .SI(CRC_OUT_4_13), .SE(n10109), .CLK(
        n10836), .Q(CRC_OUT_4_14), .QN(DFF_1134_n1) );
  SDFFX1 DFF_1135_Q_reg ( .D(WX7759), .SI(CRC_OUT_4_14), .SE(n10109), .CLK(
        n10836), .Q(CRC_OUT_4_15), .QN(DFF_1135_n1) );
  SDFFX1 DFF_1136_Q_reg ( .D(WX7761), .SI(CRC_OUT_4_15), .SE(n10109), .CLK(
        n10836), .Q(CRC_OUT_4_16), .QN(DFF_1136_n1) );
  SDFFX1 DFF_1137_Q_reg ( .D(WX7763), .SI(CRC_OUT_4_16), .SE(n10109), .CLK(
        n10836), .Q(CRC_OUT_4_17), .QN(DFF_1137_n1) );
  SDFFX1 DFF_1138_Q_reg ( .D(WX7765), .SI(CRC_OUT_4_17), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_18), .QN(DFF_1138_n1) );
  SDFFX1 DFF_1139_Q_reg ( .D(WX7767), .SI(CRC_OUT_4_18), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_19), .QN(DFF_1139_n1) );
  SDFFX1 DFF_1140_Q_reg ( .D(WX7769), .SI(CRC_OUT_4_19), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_20), .QN(DFF_1140_n1) );
  SDFFX1 DFF_1141_Q_reg ( .D(WX7771), .SI(CRC_OUT_4_20), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_21), .QN(DFF_1141_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(WX7773), .SI(CRC_OUT_4_21), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_22), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(WX7775), .SI(CRC_OUT_4_22), .SE(n10108), .CLK(
        n10836), .Q(CRC_OUT_4_23), .QN(DFF_1143_n1) );
  SDFFX1 DFF_1144_Q_reg ( .D(WX7777), .SI(CRC_OUT_4_23), .SE(n10107), .CLK(
        n10837), .Q(CRC_OUT_4_24), .QN(DFF_1144_n1) );
  SDFFX1 DFF_1145_Q_reg ( .D(WX7779), .SI(CRC_OUT_4_24), .SE(n10107), .CLK(
        n10837), .Q(CRC_OUT_4_25), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(WX7781), .SI(CRC_OUT_4_25), .SE(n10207), .CLK(
        n10786), .Q(CRC_OUT_4_26), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(WX7783), .SI(CRC_OUT_4_26), .SE(n10207), .CLK(
        n10786), .Q(CRC_OUT_4_27), .QN(DFF_1147_n1) );
  SDFFX1 DFF_1148_Q_reg ( .D(WX7785), .SI(CRC_OUT_4_27), .SE(n10206), .CLK(
        n10786), .Q(CRC_OUT_4_28), .QN(DFF_1148_n1) );
  SDFFX1 DFF_1149_Q_reg ( .D(WX7787), .SI(CRC_OUT_4_28), .SE(n10206), .CLK(
        n10787), .Q(test_so66), .QN(n9939) );
  SDFFX1 DFF_1150_Q_reg ( .D(WX7789), .SI(test_si67), .SE(n10206), .CLK(n10787), .Q(CRC_OUT_4_30), .QN(DFF_1150_n1) );
  SDFFX1 DFF_1151_Q_reg ( .D(WX7791), .SI(CRC_OUT_4_30), .SE(n10206), .CLK(
        n10787), .Q(CRC_OUT_4_31), .QN(DFF_1151_n1) );
  SDFFX1 DFF_1152_Q_reg ( .D(n1455), .SI(CRC_OUT_4_31), .SE(n10206), .CLK(
        n10787), .Q(WX8243), .QN(n9849) );
  SDFFX1 DFF_1153_Q_reg ( .D(n1456), .SI(WX8243), .SE(n10201), .CLK(n10789), 
        .Q(n8411), .QN(n3878) );
  SDFFX1 DFF_1154_Q_reg ( .D(n1457), .SI(n8411), .SE(n10201), .CLK(n10789), 
        .Q(n8410), .QN(n3877) );
  SDFFX1 DFF_1155_Q_reg ( .D(n1458), .SI(n8410), .SE(n10201), .CLK(n10789), 
        .Q(n8409), .QN(n3876) );
  SDFFX1 DFF_1156_Q_reg ( .D(n1459), .SI(n8409), .SE(n10201), .CLK(n10789), 
        .Q(n8408), .QN(n3875) );
  SDFFX1 DFF_1157_Q_reg ( .D(n1460), .SI(n8408), .SE(n10201), .CLK(n10789), 
        .Q(n8407), .QN(n3874) );
  SDFFX1 DFF_1158_Q_reg ( .D(n1461), .SI(n8407), .SE(n10201), .CLK(n10789), 
        .Q(n8406), .QN(n3873) );
  SDFFX1 DFF_1159_Q_reg ( .D(n1462), .SI(n8406), .SE(n10202), .CLK(n10789), 
        .Q(n8405), .QN(n3872) );
  SDFFX1 DFF_1160_Q_reg ( .D(n1463), .SI(n8405), .SE(n10202), .CLK(n10789), 
        .Q(n8404), .QN(n3871) );
  SDFFX1 DFF_1161_Q_reg ( .D(n1464), .SI(n8404), .SE(n10202), .CLK(n10789), 
        .Q(n8403), .QN(n3870) );
  SDFFX1 DFF_1162_Q_reg ( .D(n1465), .SI(n8403), .SE(n10202), .CLK(n10789), 
        .Q(n8402), .QN(n3869) );
  SDFFX1 DFF_1163_Q_reg ( .D(n1466), .SI(n8402), .SE(n10202), .CLK(n10789), 
        .Q(n8401), .QN(n3868) );
  SDFFX1 DFF_1164_Q_reg ( .D(n1467), .SI(n8401), .SE(n10202), .CLK(n10788), 
        .Q(n8400), .QN(n3867) );
  SDFFX1 DFF_1165_Q_reg ( .D(n1468), .SI(n8400), .SE(n10203), .CLK(n10788), 
        .Q(n8399), .QN(n3866) );
  SDFFX1 DFF_1166_Q_reg ( .D(n1469), .SI(n8399), .SE(n10203), .CLK(n10788), 
        .Q(test_so67), .QN(n3865) );
  SDFFX1 DFF_1167_Q_reg ( .D(n1470), .SI(test_si68), .SE(n10203), .CLK(n10788), 
        .Q(n8396), .QN(n3864) );
  SDFFX1 DFF_1168_Q_reg ( .D(n1471), .SI(n8396), .SE(n10203), .CLK(n10788), 
        .Q(n8395), .QN(n3863) );
  SDFFX1 DFF_1169_Q_reg ( .D(n1472), .SI(n8395), .SE(n10203), .CLK(n10788), 
        .Q(n8394), .QN(n3862) );
  SDFFX1 DFF_1170_Q_reg ( .D(n1473), .SI(n8394), .SE(n10203), .CLK(n10788), 
        .Q(n8393), .QN(n3861) );
  SDFFX1 DFF_1171_Q_reg ( .D(n1474), .SI(n8393), .SE(n10204), .CLK(n10788), 
        .Q(n8392), .QN(n3860) );
  SDFFX1 DFF_1172_Q_reg ( .D(n1475), .SI(n8392), .SE(n10204), .CLK(n10788), 
        .Q(n8391), .QN(n3859) );
  SDFFX1 DFF_1173_Q_reg ( .D(n1476), .SI(n8391), .SE(n10204), .CLK(n10788), 
        .Q(n8390), .QN(n3858) );
  SDFFX1 DFF_1174_Q_reg ( .D(n1477), .SI(n8390), .SE(n10204), .CLK(n10788), 
        .Q(n8389), .QN(n3857) );
  SDFFX1 DFF_1175_Q_reg ( .D(n1478), .SI(n8389), .SE(n10204), .CLK(n10788), 
        .Q(n8388), .QN(n3856) );
  SDFFX1 DFF_1176_Q_reg ( .D(n1479), .SI(n8388), .SE(n10204), .CLK(n10787), 
        .Q(n8387), .QN(n3855) );
  SDFFX1 DFF_1177_Q_reg ( .D(n1480), .SI(n8387), .SE(n10205), .CLK(n10787), 
        .Q(n8386), .QN(n3854) );
  SDFFX1 DFF_1178_Q_reg ( .D(n1481), .SI(n8386), .SE(n10205), .CLK(n10787), 
        .Q(n8385), .QN(n3853) );
  SDFFX1 DFF_1179_Q_reg ( .D(n1482), .SI(n8385), .SE(n10205), .CLK(n10787), 
        .Q(n8384), .QN(n3852) );
  SDFFX1 DFF_1180_Q_reg ( .D(n1483), .SI(n8384), .SE(n10205), .CLK(n10787), 
        .Q(n8383), .QN(n3851) );
  SDFFX1 DFF_1181_Q_reg ( .D(n1484), .SI(n8383), .SE(n10205), .CLK(n10787), 
        .Q(n8382), .QN(n3850) );
  SDFFX1 DFF_1182_Q_reg ( .D(n1485), .SI(n8382), .SE(n10205), .CLK(n10787), 
        .Q(n8381), .QN(n3849) );
  SDFFX1 DFF_1183_Q_reg ( .D(WX8304), .SI(n8381), .SE(n10206), .CLK(n10787), 
        .Q(test_so68), .QN(n3848) );
  SDFFX1 DFF_1184_Q_reg ( .D(WX8402), .SI(test_si69), .SE(n10112), .CLK(n10834), .Q(n8378), .QN(n17911) );
  SDFFX1 DFF_1185_Q_reg ( .D(WX8404), .SI(n8378), .SE(n10200), .CLK(n10789), 
        .Q(n8377), .QN(n17910) );
  SDFFX1 DFF_1186_Q_reg ( .D(WX8406), .SI(n8377), .SE(n10200), .CLK(n10790), 
        .Q(n8376), .QN(n17909) );
  SDFFX1 DFF_1187_Q_reg ( .D(WX8408), .SI(n8376), .SE(n10199), .CLK(n10790), 
        .Q(n8375), .QN(n17908) );
  SDFFX1 DFF_1188_Q_reg ( .D(WX8410), .SI(n8375), .SE(n10199), .CLK(n10790), 
        .Q(n8374), .QN(n17907) );
  SDFFX1 DFF_1189_Q_reg ( .D(WX8412), .SI(n8374), .SE(n10198), .CLK(n10791), 
        .Q(n8373), .QN(n17906) );
  SDFFX1 DFF_1190_Q_reg ( .D(WX8414), .SI(n8373), .SE(n10198), .CLK(n10791), 
        .Q(n8372), .QN(n17905) );
  SDFFX1 DFF_1191_Q_reg ( .D(WX8416), .SI(n8372), .SE(n10197), .CLK(n10791), 
        .Q(n8371), .QN(n17904) );
  SDFFX1 DFF_1192_Q_reg ( .D(WX8418), .SI(n8371), .SE(n10197), .CLK(n10791), 
        .Q(n8370), .QN(n17903) );
  SDFFX1 DFF_1193_Q_reg ( .D(WX8420), .SI(n8370), .SE(n10195), .CLK(n10792), 
        .Q(n8369), .QN(n17902) );
  SDFFX1 DFF_1194_Q_reg ( .D(WX8422), .SI(n8369), .SE(n10195), .CLK(n10792), 
        .Q(n8368), .QN(n17901) );
  SDFFX1 DFF_1195_Q_reg ( .D(WX8424), .SI(n8368), .SE(n10194), .CLK(n10793), 
        .Q(n8367), .QN(n17900) );
  SDFFX1 DFF_1196_Q_reg ( .D(WX8426), .SI(n8367), .SE(n10194), .CLK(n10793), 
        .Q(n8366), .QN(n17899) );
  SDFFX1 DFF_1197_Q_reg ( .D(WX8428), .SI(n8366), .SE(n10193), .CLK(n10793), 
        .Q(n8365), .QN(n17898) );
  SDFFX1 DFF_1198_Q_reg ( .D(WX8430), .SI(n8365), .SE(n10193), .CLK(n10793), 
        .Q(n8364), .QN(n17897) );
  SDFFX1 DFF_1199_Q_reg ( .D(WX8432), .SI(n8364), .SE(n10191), .CLK(n10794), 
        .Q(n8363), .QN(n17896) );
  SDFFX1 DFF_1200_Q_reg ( .D(WX8434), .SI(n8363), .SE(n10191), .CLK(n10794), 
        .Q(test_so69), .QN(n9919) );
  SDFFX1 DFF_1201_Q_reg ( .D(WX8436), .SI(test_si70), .SE(n10190), .CLK(n10795), .Q(WX8437), .QN(n9358) );
  SDFFX1 DFF_1202_Q_reg ( .D(WX8438), .SI(WX8437), .SE(n10190), .CLK(n10795), 
        .Q(WX8439), .QN(n9356) );
  SDFFX1 DFF_1203_Q_reg ( .D(WX8440), .SI(WX8439), .SE(n10189), .CLK(n10795), 
        .Q(WX8441), .QN(n9354) );
  SDFFX1 DFF_1204_Q_reg ( .D(WX8442), .SI(WX8441), .SE(n10336), .CLK(n10722), 
        .Q(WX8443) );
  SDFFX1 DFF_1205_Q_reg ( .D(WX8444), .SI(WX8443), .SE(n10188), .CLK(n10796), 
        .Q(WX8445), .QN(n9351) );
  SDFFX1 DFF_1206_Q_reg ( .D(WX8446), .SI(WX8445), .SE(n10187), .CLK(n10796), 
        .Q(WX8447) );
  SDFFX1 DFF_1207_Q_reg ( .D(WX8448), .SI(WX8447), .SE(n10187), .CLK(n10796), 
        .Q(WX8449), .QN(n9347) );
  SDFFX1 DFF_1208_Q_reg ( .D(WX8450), .SI(WX8449), .SE(n10186), .CLK(n10797), 
        .Q(WX8451), .QN(n9345) );
  SDFFX1 DFF_1209_Q_reg ( .D(WX8452), .SI(WX8451), .SE(n10185), .CLK(n10797), 
        .Q(WX8453), .QN(n9343) );
  SDFFX1 DFF_1210_Q_reg ( .D(WX8454), .SI(WX8453), .SE(n10185), .CLK(n10797), 
        .Q(WX8455), .QN(n9341) );
  SDFFX1 DFF_1211_Q_reg ( .D(WX8456), .SI(WX8455), .SE(n10184), .CLK(n10798), 
        .Q(WX8457), .QN(n9339) );
  SDFFX1 DFF_1212_Q_reg ( .D(WX8458), .SI(WX8457), .SE(n10183), .CLK(n10798), 
        .Q(WX8459), .QN(n9337) );
  SDFFX1 DFF_1213_Q_reg ( .D(WX8460), .SI(WX8459), .SE(n10183), .CLK(n10798), 
        .Q(WX8461), .QN(n9335) );
  SDFFX1 DFF_1214_Q_reg ( .D(WX8462), .SI(WX8461), .SE(n10182), .CLK(n10799), 
        .Q(WX8463), .QN(n9333) );
  SDFFX1 DFF_1215_Q_reg ( .D(WX8464), .SI(WX8463), .SE(n10181), .CLK(n10799), 
        .Q(WX8465), .QN(n9331) );
  SDFFX1 DFF_1216_Q_reg ( .D(WX8466), .SI(WX8465), .SE(n10181), .CLK(n10799), 
        .Q(WX8467), .QN(n9032) );
  SDFFX1 DFF_1217_Q_reg ( .D(WX8468), .SI(WX8467), .SE(n10200), .CLK(n10790), 
        .Q(test_so70), .QN(n9956) );
  SDFFX1 DFF_1218_Q_reg ( .D(WX8470), .SI(test_si71), .SE(n10200), .CLK(n10790), .Q(WX8471), .QN(n9125) );
  SDFFX1 DFF_1219_Q_reg ( .D(WX8472), .SI(WX8471), .SE(n10199), .CLK(n10790), 
        .Q(WX8473), .QN(n9124) );
  SDFFX1 DFF_1220_Q_reg ( .D(WX8474), .SI(WX8473), .SE(n10199), .CLK(n10790), 
        .Q(WX8475), .QN(n9122) );
  SDFFX1 DFF_1221_Q_reg ( .D(WX8476), .SI(WX8475), .SE(n10198), .CLK(n10790), 
        .Q(WX8477), .QN(n9120) );
  SDFFX1 DFF_1222_Q_reg ( .D(WX8478), .SI(WX8477), .SE(n10198), .CLK(n10791), 
        .Q(WX8479), .QN(n9118) );
  SDFFX1 DFF_1223_Q_reg ( .D(WX8480), .SI(WX8479), .SE(n10197), .CLK(n10791), 
        .Q(WX8481), .QN(n9116) );
  SDFFX1 DFF_1224_Q_reg ( .D(WX8482), .SI(WX8481), .SE(n10196), .CLK(n10791), 
        .Q(WX8483), .QN(n9114) );
  SDFFX1 DFF_1225_Q_reg ( .D(WX8484), .SI(WX8483), .SE(n10196), .CLK(n10792), 
        .Q(WX8485), .QN(n9112) );
  SDFFX1 DFF_1226_Q_reg ( .D(WX8486), .SI(WX8485), .SE(n10195), .CLK(n10792), 
        .Q(WX8487), .QN(n9110) );
  SDFFX1 DFF_1227_Q_reg ( .D(WX8488), .SI(WX8487), .SE(n10195), .CLK(n10792), 
        .Q(WX8489), .QN(n9108) );
  SDFFX1 DFF_1228_Q_reg ( .D(WX8490), .SI(WX8489), .SE(n10194), .CLK(n10793), 
        .Q(WX8491), .QN(n9106) );
  SDFFX1 DFF_1229_Q_reg ( .D(WX8492), .SI(WX8491), .SE(n10193), .CLK(n10793), 
        .Q(WX8493), .QN(n9104) );
  SDFFX1 DFF_1230_Q_reg ( .D(WX8494), .SI(WX8493), .SE(n10192), .CLK(n10793), 
        .Q(WX8495), .QN(n9102) );
  SDFFX1 DFF_1231_Q_reg ( .D(WX8496), .SI(WX8495), .SE(n10192), .CLK(n10794), 
        .Q(WX8497), .QN(n9100) );
  SDFFX1 DFF_1232_Q_reg ( .D(WX8498), .SI(WX8497), .SE(n10191), .CLK(n10794), 
        .Q(WX8499), .QN(n3625) );
  SDFFX1 DFF_1233_Q_reg ( .D(WX8500), .SI(WX8499), .SE(n10191), .CLK(n10794), 
        .Q(WX8501), .QN(n3623) );
  SDFFX1 DFF_1234_Q_reg ( .D(WX8502), .SI(WX8501), .SE(n10190), .CLK(n10795), 
        .Q(test_so71), .QN(n9918) );
  SDFFX1 DFF_1235_Q_reg ( .D(WX8504), .SI(test_si72), .SE(n10189), .CLK(n10795), .Q(WX8505), .QN(n3619) );
  SDFFX1 DFF_1236_Q_reg ( .D(WX8506), .SI(WX8505), .SE(n10189), .CLK(n10795), 
        .Q(WX8507), .QN(n3617) );
  SDFFX1 DFF_1237_Q_reg ( .D(WX8508), .SI(WX8507), .SE(n10188), .CLK(n10796), 
        .Q(WX8509), .QN(n3615) );
  SDFFX1 DFF_1238_Q_reg ( .D(WX8510), .SI(WX8509), .SE(n10187), .CLK(n10796), 
        .Q(WX8511), .QN(n3613) );
  SDFFX1 DFF_1239_Q_reg ( .D(WX8512), .SI(WX8511), .SE(n10187), .CLK(n10796), 
        .Q(WX8513), .QN(n3611) );
  SDFFX1 DFF_1240_Q_reg ( .D(WX8514), .SI(WX8513), .SE(n10186), .CLK(n10797), 
        .Q(WX8515), .QN(n3609) );
  SDFFX1 DFF_1241_Q_reg ( .D(WX8516), .SI(WX8515), .SE(n10185), .CLK(n10797), 
        .Q(WX8517), .QN(n3607) );
  SDFFX1 DFF_1242_Q_reg ( .D(WX8518), .SI(WX8517), .SE(n10185), .CLK(n10797), 
        .Q(WX8519), .QN(n3605) );
  SDFFX1 DFF_1243_Q_reg ( .D(WX8520), .SI(WX8519), .SE(n10184), .CLK(n10798), 
        .Q(WX8521), .QN(n3603) );
  SDFFX1 DFF_1244_Q_reg ( .D(WX8522), .SI(WX8521), .SE(n10183), .CLK(n10798), 
        .Q(WX8523), .QN(n3601) );
  SDFFX1 DFF_1245_Q_reg ( .D(WX8524), .SI(WX8523), .SE(n10183), .CLK(n10798), 
        .Q(WX8525), .QN(n3599) );
  SDFFX1 DFF_1246_Q_reg ( .D(WX8526), .SI(WX8525), .SE(n10182), .CLK(n10799), 
        .Q(WX8527), .QN(n3597) );
  SDFFX1 DFF_1247_Q_reg ( .D(WX8528), .SI(WX8527), .SE(n10181), .CLK(n10799), 
        .Q(WX8529), .QN(n3595) );
  SDFFX1 DFF_1248_Q_reg ( .D(WX8530), .SI(WX8529), .SE(n10181), .CLK(n10799), 
        .Q(WX8531), .QN(n9033) );
  SDFFX1 DFF_1249_Q_reg ( .D(WX8532), .SI(WX8531), .SE(n10200), .CLK(n10790), 
        .Q(WX8533), .QN(n9127) );
  SDFFX1 DFF_1250_Q_reg ( .D(WX8534), .SI(WX8533), .SE(n10200), .CLK(n10790), 
        .Q(WX8535), .QN(n9126) );
  SDFFX1 DFF_1251_Q_reg ( .D(WX8536), .SI(WX8535), .SE(n10199), .CLK(n10790), 
        .Q(test_so72), .QN(n9955) );
  SDFFX1 DFF_1252_Q_reg ( .D(WX8538), .SI(test_si73), .SE(n10199), .CLK(n10790), .Q(WX8539), .QN(n9123) );
  SDFFX1 DFF_1253_Q_reg ( .D(WX8540), .SI(WX8539), .SE(n10198), .CLK(n10791), 
        .Q(WX8541) );
  SDFFX1 DFF_1254_Q_reg ( .D(WX8542), .SI(WX8541), .SE(n10198), .CLK(n10791), 
        .Q(WX8543), .QN(n9119) );
  SDFFX1 DFF_1255_Q_reg ( .D(WX8544), .SI(WX8543), .SE(n10197), .CLK(n10791), 
        .Q(WX8545), .QN(n9117) );
  SDFFX1 DFF_1256_Q_reg ( .D(WX8546), .SI(WX8545), .SE(n10196), .CLK(n10792), 
        .Q(WX8547), .QN(n9115) );
  SDFFX1 DFF_1257_Q_reg ( .D(WX8548), .SI(WX8547), .SE(n10196), .CLK(n10792), 
        .Q(WX8549), .QN(n9113) );
  SDFFX1 DFF_1258_Q_reg ( .D(WX8550), .SI(WX8549), .SE(n10195), .CLK(n10792), 
        .Q(WX8551), .QN(n9111) );
  SDFFX1 DFF_1259_Q_reg ( .D(WX8552), .SI(WX8551), .SE(n10194), .CLK(n10792), 
        .Q(WX8553), .QN(n9109) );
  SDFFX1 DFF_1260_Q_reg ( .D(WX8554), .SI(WX8553), .SE(n10194), .CLK(n10793), 
        .Q(WX8555), .QN(n9107) );
  SDFFX1 DFF_1261_Q_reg ( .D(WX8556), .SI(WX8555), .SE(n10193), .CLK(n10793), 
        .Q(WX8557), .QN(n9105) );
  SDFFX1 DFF_1262_Q_reg ( .D(WX8558), .SI(WX8557), .SE(n10192), .CLK(n10794), 
        .Q(WX8559), .QN(n9103) );
  SDFFX1 DFF_1263_Q_reg ( .D(WX8560), .SI(WX8559), .SE(n10192), .CLK(n10794), 
        .Q(WX8561), .QN(n9101) );
  SDFFX1 DFF_1264_Q_reg ( .D(WX8562), .SI(WX8561), .SE(n10191), .CLK(n10794), 
        .Q(WX8563) );
  SDFFX1 DFF_1265_Q_reg ( .D(WX8564), .SI(WX8563), .SE(n10190), .CLK(n10794), 
        .Q(WX8565), .QN(n9359) );
  SDFFX1 DFF_1266_Q_reg ( .D(WX8566), .SI(WX8565), .SE(n10190), .CLK(n10795), 
        .Q(WX8567) );
  SDFFX1 DFF_1267_Q_reg ( .D(WX8568), .SI(WX8567), .SE(n10189), .CLK(n10795), 
        .Q(WX8569), .QN(n9355) );
  SDFFX1 DFF_1268_Q_reg ( .D(WX8570), .SI(WX8569), .SE(n10188), .CLK(n10795), 
        .Q(test_so73), .QN(n9917) );
  SDFFX1 DFF_1269_Q_reg ( .D(WX8572), .SI(test_si74), .SE(n10188), .CLK(n10796), .Q(WX8573), .QN(n9352) );
  SDFFX1 DFF_1270_Q_reg ( .D(WX8574), .SI(WX8573), .SE(n10187), .CLK(n10796), 
        .Q(WX8575), .QN(n9350) );
  SDFFX1 DFF_1271_Q_reg ( .D(WX8576), .SI(WX8575), .SE(n10186), .CLK(n10796), 
        .Q(WX8577), .QN(n9348) );
  SDFFX1 DFF_1272_Q_reg ( .D(WX8578), .SI(WX8577), .SE(n10186), .CLK(n10797), 
        .Q(WX8579), .QN(n9346) );
  SDFFX1 DFF_1273_Q_reg ( .D(WX8580), .SI(WX8579), .SE(n10185), .CLK(n10797), 
        .Q(WX8581), .QN(n9344) );
  SDFFX1 DFF_1274_Q_reg ( .D(WX8582), .SI(WX8581), .SE(n10184), .CLK(n10797), 
        .Q(WX8583), .QN(n9342) );
  SDFFX1 DFF_1275_Q_reg ( .D(WX8584), .SI(WX8583), .SE(n10184), .CLK(n10798), 
        .Q(WX8585), .QN(n9340) );
  SDFFX1 DFF_1276_Q_reg ( .D(WX8586), .SI(WX8585), .SE(n10183), .CLK(n10798), 
        .Q(WX8587), .QN(n9338) );
  SDFFX1 DFF_1277_Q_reg ( .D(WX8588), .SI(WX8587), .SE(n10182), .CLK(n10798), 
        .Q(WX8589), .QN(n9336) );
  SDFFX1 DFF_1278_Q_reg ( .D(WX8590), .SI(WX8589), .SE(n10182), .CLK(n10799), 
        .Q(WX8591), .QN(n9334) );
  SDFFX1 DFF_1279_Q_reg ( .D(WX8592), .SI(WX8591), .SE(n10181), .CLK(n10799), 
        .Q(WX8593), .QN(n9332) );
  SDFFX1 DFF_1280_Q_reg ( .D(WX8594), .SI(WX8593), .SE(n10180), .CLK(n10799), 
        .Q(WX8595), .QN(n9593) );
  SDFFX1 DFF_1281_Q_reg ( .D(WX8596), .SI(WX8595), .SE(n10180), .CLK(n10800), 
        .Q(WX8597), .QN(n9594) );
  SDFFX1 DFF_1282_Q_reg ( .D(WX8598), .SI(WX8597), .SE(n10180), .CLK(n10800), 
        .Q(WX8599), .QN(n9595) );
  SDFFX1 DFF_1283_Q_reg ( .D(WX8600), .SI(WX8599), .SE(n10180), .CLK(n10800), 
        .Q(WX8601), .QN(n9596) );
  SDFFX1 DFF_1284_Q_reg ( .D(WX8602), .SI(WX8601), .SE(n10180), .CLK(n10800), 
        .Q(WX8603), .QN(n9597) );
  SDFFX1 DFF_1285_Q_reg ( .D(WX8604), .SI(WX8603), .SE(n10180), .CLK(n10800), 
        .Q(test_so74), .QN(n9908) );
  SDFFX1 DFF_1286_Q_reg ( .D(WX8606), .SI(test_si75), .SE(n10197), .CLK(n10791), .Q(WX8607), .QN(n9598) );
  SDFFX1 DFF_1287_Q_reg ( .D(WX8608), .SI(WX8607), .SE(n10197), .CLK(n10791), 
        .Q(WX8609), .QN(n9599) );
  SDFFX1 DFF_1288_Q_reg ( .D(WX8610), .SI(WX8609), .SE(n10196), .CLK(n10792), 
        .Q(WX8611), .QN(n9600) );
  SDFFX1 DFF_1289_Q_reg ( .D(WX8612), .SI(WX8611), .SE(n10196), .CLK(n10792), 
        .Q(WX8613), .QN(n9601) );
  SDFFX1 DFF_1290_Q_reg ( .D(WX8614), .SI(WX8613), .SE(n10195), .CLK(n10792), 
        .Q(WX8615), .QN(n9602) );
  SDFFX1 DFF_1291_Q_reg ( .D(WX8616), .SI(WX8615), .SE(n10194), .CLK(n10793), 
        .Q(WX8617), .QN(n9603) );
  SDFFX1 DFF_1292_Q_reg ( .D(WX8618), .SI(WX8617), .SE(n10193), .CLK(n10793), 
        .Q(WX8619), .QN(n9604) );
  SDFFX1 DFF_1293_Q_reg ( .D(WX8620), .SI(WX8619), .SE(n10193), .CLK(n10793), 
        .Q(WX8621), .QN(n9605) );
  SDFFX1 DFF_1294_Q_reg ( .D(WX8622), .SI(WX8621), .SE(n10192), .CLK(n10794), 
        .Q(WX8623), .QN(n9606) );
  SDFFX1 DFF_1295_Q_reg ( .D(WX8624), .SI(WX8623), .SE(n10192), .CLK(n10794), 
        .Q(WX8625), .QN(n9518) );
  SDFFX1 DFF_1296_Q_reg ( .D(WX8626), .SI(WX8625), .SE(n10191), .CLK(n10794), 
        .Q(WX8627), .QN(n9607) );
  SDFFX1 DFF_1297_Q_reg ( .D(WX8628), .SI(WX8627), .SE(n10190), .CLK(n10795), 
        .Q(WX8629), .QN(n9608) );
  SDFFX1 DFF_1298_Q_reg ( .D(WX8630), .SI(WX8629), .SE(n10189), .CLK(n10795), 
        .Q(WX8631), .QN(n9609) );
  SDFFX1 DFF_1299_Q_reg ( .D(WX8632), .SI(WX8631), .SE(n10189), .CLK(n10795), 
        .Q(WX8633), .QN(n9610) );
  SDFFX1 DFF_1300_Q_reg ( .D(WX8634), .SI(WX8633), .SE(n10188), .CLK(n10796), 
        .Q(WX8635), .QN(n9519) );
  SDFFX1 DFF_1301_Q_reg ( .D(WX8636), .SI(WX8635), .SE(n10188), .CLK(n10796), 
        .Q(WX8637), .QN(n9611) );
  SDFFX1 DFF_1302_Q_reg ( .D(WX8638), .SI(WX8637), .SE(n10187), .CLK(n10796), 
        .Q(test_so75), .QN(n9903) );
  SDFFX1 DFF_1303_Q_reg ( .D(WX8640), .SI(test_si76), .SE(n10186), .CLK(n10797), .Q(WX8641), .QN(n9612) );
  SDFFX1 DFF_1304_Q_reg ( .D(WX8642), .SI(WX8641), .SE(n10186), .CLK(n10797), 
        .Q(WX8643), .QN(n9613) );
  SDFFX1 DFF_1305_Q_reg ( .D(WX8644), .SI(WX8643), .SE(n10185), .CLK(n10797), 
        .Q(WX8645), .QN(n9614) );
  SDFFX1 DFF_1306_Q_reg ( .D(WX8646), .SI(WX8645), .SE(n10184), .CLK(n10798), 
        .Q(WX8647), .QN(n9615) );
  SDFFX1 DFF_1307_Q_reg ( .D(WX8648), .SI(WX8647), .SE(n10184), .CLK(n10798), 
        .Q(WX8649), .QN(n9520) );
  SDFFX1 DFF_1308_Q_reg ( .D(WX8650), .SI(WX8649), .SE(n10183), .CLK(n10798), 
        .Q(WX8651), .QN(n9616) );
  SDFFX1 DFF_1309_Q_reg ( .D(WX8652), .SI(WX8651), .SE(n10182), .CLK(n10799), 
        .Q(WX8653), .QN(n9617) );
  SDFFX1 DFF_1310_Q_reg ( .D(WX8654), .SI(WX8653), .SE(n10182), .CLK(n10799), 
        .Q(WX8655), .QN(n9618) );
  SDFFX1 DFF_1311_Q_reg ( .D(WX8656), .SI(WX8655), .SE(n10181), .CLK(n10799), 
        .Q(WX8657), .QN(n9535) );
  SDFFX1 DFF_1312_Q_reg ( .D(WX9022), .SI(WX8657), .SE(n10117), .CLK(n10832), 
        .Q(CRC_OUT_3_0), .QN(DFF_1312_n1) );
  SDFFX1 DFF_1313_Q_reg ( .D(WX9024), .SI(CRC_OUT_3_0), .SE(n10117), .CLK(
        n10832), .Q(CRC_OUT_3_1), .QN(DFF_1313_n1) );
  SDFFX1 DFF_1314_Q_reg ( .D(WX9026), .SI(CRC_OUT_3_1), .SE(n10116), .CLK(
        n10832), .Q(CRC_OUT_3_2), .QN(DFF_1314_n1) );
  SDFFX1 DFF_1315_Q_reg ( .D(WX9028), .SI(CRC_OUT_3_2), .SE(n10116), .CLK(
        n10832), .Q(CRC_OUT_3_3), .QN(DFF_1315_n1) );
  SDFFX1 DFF_1316_Q_reg ( .D(WX9030), .SI(CRC_OUT_3_3), .SE(n10116), .CLK(
        n10832), .Q(CRC_OUT_3_4), .QN(DFF_1316_n1) );
  SDFFX1 DFF_1317_Q_reg ( .D(WX9032), .SI(CRC_OUT_3_4), .SE(n10116), .CLK(
        n10832), .Q(CRC_OUT_3_5), .QN(DFF_1317_n1) );
  SDFFX1 DFF_1318_Q_reg ( .D(WX9034), .SI(CRC_OUT_3_5), .SE(n10116), .CLK(
        n10832), .Q(CRC_OUT_3_6), .QN(DFF_1318_n1) );
  SDFFX1 DFF_1319_Q_reg ( .D(WX9036), .SI(CRC_OUT_3_6), .SE(n10116), .CLK(
        n10832), .Q(test_so76), .QN(n9938) );
  SDFFX1 DFF_1320_Q_reg ( .D(WX9038), .SI(test_si77), .SE(n10115), .CLK(n10833), .Q(CRC_OUT_3_8), .QN(DFF_1320_n1) );
  SDFFX1 DFF_1321_Q_reg ( .D(WX9040), .SI(CRC_OUT_3_8), .SE(n10115), .CLK(
        n10833), .Q(CRC_OUT_3_9), .QN(DFF_1321_n1) );
  SDFFX1 DFF_1322_Q_reg ( .D(WX9042), .SI(CRC_OUT_3_9), .SE(n10115), .CLK(
        n10833), .Q(CRC_OUT_3_10), .QN(DFF_1322_n1) );
  SDFFX1 DFF_1323_Q_reg ( .D(WX9044), .SI(CRC_OUT_3_10), .SE(n10115), .CLK(
        n10833), .Q(CRC_OUT_3_11), .QN(DFF_1323_n1) );
  SDFFX1 DFF_1324_Q_reg ( .D(WX9046), .SI(CRC_OUT_3_11), .SE(n10115), .CLK(
        n10833), .Q(CRC_OUT_3_12), .QN(DFF_1324_n1) );
  SDFFX1 DFF_1325_Q_reg ( .D(WX9048), .SI(CRC_OUT_3_12), .SE(n10115), .CLK(
        n10833), .Q(CRC_OUT_3_13), .QN(DFF_1325_n1) );
  SDFFX1 DFF_1326_Q_reg ( .D(WX9050), .SI(CRC_OUT_3_13), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_14), .QN(DFF_1326_n1) );
  SDFFX1 DFF_1327_Q_reg ( .D(WX9052), .SI(CRC_OUT_3_14), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_15), .QN(DFF_1327_n1) );
  SDFFX1 DFF_1328_Q_reg ( .D(WX9054), .SI(CRC_OUT_3_15), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_16), .QN(DFF_1328_n1) );
  SDFFX1 DFF_1329_Q_reg ( .D(WX9056), .SI(CRC_OUT_3_16), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_17), .QN(DFF_1329_n1) );
  SDFFX1 DFF_1330_Q_reg ( .D(WX9058), .SI(CRC_OUT_3_17), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_18), .QN(DFF_1330_n1) );
  SDFFX1 DFF_1331_Q_reg ( .D(WX9060), .SI(CRC_OUT_3_18), .SE(n10114), .CLK(
        n10833), .Q(CRC_OUT_3_19), .QN(DFF_1331_n1) );
  SDFFX1 DFF_1332_Q_reg ( .D(WX9062), .SI(CRC_OUT_3_19), .SE(n10113), .CLK(
        n10834), .Q(CRC_OUT_3_20), .QN(DFF_1332_n1) );
  SDFFX1 DFF_1333_Q_reg ( .D(WX9064), .SI(CRC_OUT_3_20), .SE(n10113), .CLK(
        n10834), .Q(CRC_OUT_3_21), .QN(DFF_1333_n1) );
  SDFFX1 DFF_1334_Q_reg ( .D(WX9066), .SI(CRC_OUT_3_21), .SE(n10113), .CLK(
        n10834), .Q(CRC_OUT_3_22), .QN(DFF_1334_n1) );
  SDFFX1 DFF_1335_Q_reg ( .D(WX9068), .SI(CRC_OUT_3_22), .SE(n10113), .CLK(
        n10834), .Q(CRC_OUT_3_23), .QN(DFF_1335_n1) );
  SDFFX1 DFF_1336_Q_reg ( .D(WX9070), .SI(CRC_OUT_3_23), .SE(n10113), .CLK(
        n10834), .Q(test_so77), .QN(n9937) );
  SDFFX1 DFF_1337_Q_reg ( .D(WX9072), .SI(test_si78), .SE(n10113), .CLK(n10834), .Q(CRC_OUT_3_25), .QN(DFF_1337_n1) );
  SDFFX1 DFF_1338_Q_reg ( .D(WX9074), .SI(CRC_OUT_3_25), .SE(n10112), .CLK(
        n10834), .Q(CRC_OUT_3_26), .QN(DFF_1338_n1) );
  SDFFX1 DFF_1339_Q_reg ( .D(WX9076), .SI(CRC_OUT_3_26), .SE(n10112), .CLK(
        n10834), .Q(CRC_OUT_3_27), .QN(DFF_1339_n1) );
  SDFFX1 DFF_1340_Q_reg ( .D(WX9078), .SI(CRC_OUT_3_27), .SE(n10112), .CLK(
        n10834), .Q(CRC_OUT_3_28), .QN(DFF_1340_n1) );
  SDFFX1 DFF_1341_Q_reg ( .D(WX9080), .SI(CRC_OUT_3_28), .SE(n10112), .CLK(
        n10834), .Q(CRC_OUT_3_29), .QN(DFF_1341_n1) );
  SDFFX1 DFF_1342_Q_reg ( .D(WX9082), .SI(CRC_OUT_3_29), .SE(n10112), .CLK(
        n10834), .Q(CRC_OUT_3_30), .QN(DFF_1342_n1) );
  SDFFX1 DFF_1343_Q_reg ( .D(WX9084), .SI(CRC_OUT_3_30), .SE(n10179), .CLK(
        n10800), .Q(CRC_OUT_3_31), .QN(DFF_1343_n1) );
  SDFFX1 DFF_1344_Q_reg ( .D(n1697), .SI(CRC_OUT_3_31), .SE(n10179), .CLK(
        n10800), .Q(WX9536), .QN(n9850) );
  SDFFX1 DFF_1345_Q_reg ( .D(n1698), .SI(WX9536), .SE(n10174), .CLK(n10803), 
        .Q(n8353), .QN(n3847) );
  SDFFX1 DFF_1346_Q_reg ( .D(n1699), .SI(n8353), .SE(n10174), .CLK(n10803), 
        .Q(n8352), .QN(n3846) );
  SDFFX1 DFF_1347_Q_reg ( .D(n1700), .SI(n8352), .SE(n10174), .CLK(n10802), 
        .Q(n8351), .QN(n3845) );
  SDFFX1 DFF_1348_Q_reg ( .D(n1701), .SI(n8351), .SE(n10175), .CLK(n10802), 
        .Q(n8350), .QN(n3844) );
  SDFFX1 DFF_1349_Q_reg ( .D(n1702), .SI(n8350), .SE(n10175), .CLK(n10802), 
        .Q(n8349), .QN(n3843) );
  SDFFX1 DFF_1350_Q_reg ( .D(n1703), .SI(n8349), .SE(n10175), .CLK(n10802), 
        .Q(n8348), .QN(n3842) );
  SDFFX1 DFF_1351_Q_reg ( .D(n1704), .SI(n8348), .SE(n10175), .CLK(n10802), 
        .Q(n8347), .QN(n3841) );
  SDFFX1 DFF_1352_Q_reg ( .D(n1705), .SI(n8347), .SE(n10175), .CLK(n10802), 
        .Q(n8346), .QN(n3840) );
  SDFFX1 DFF_1353_Q_reg ( .D(n1706), .SI(n8346), .SE(n10175), .CLK(n10802), 
        .Q(test_so78), .QN(n3839) );
  SDFFX1 DFF_1354_Q_reg ( .D(n1707), .SI(test_si79), .SE(n10176), .CLK(n10802), 
        .Q(n8343), .QN(n3838) );
  SDFFX1 DFF_1355_Q_reg ( .D(n1708), .SI(n8343), .SE(n10176), .CLK(n10802), 
        .Q(n8342), .QN(n3837) );
  SDFFX1 DFF_1356_Q_reg ( .D(n1709), .SI(n8342), .SE(n10176), .CLK(n10802), 
        .Q(n8341), .QN(n3836) );
  SDFFX1 DFF_1357_Q_reg ( .D(n1710), .SI(n8341), .SE(n10176), .CLK(n10802), 
        .Q(n8340), .QN(n3835) );
  SDFFX1 DFF_1358_Q_reg ( .D(n1711), .SI(n8340), .SE(n10176), .CLK(n10802), 
        .Q(n8339), .QN(n3834) );
  SDFFX1 DFF_1359_Q_reg ( .D(n1712), .SI(n8339), .SE(n10176), .CLK(n10801), 
        .Q(n8338), .QN(n3833) );
  SDFFX1 DFF_1360_Q_reg ( .D(n1713), .SI(n8338), .SE(n10177), .CLK(n10801), 
        .Q(n8337), .QN(n3832) );
  SDFFX1 DFF_1361_Q_reg ( .D(n1714), .SI(n8337), .SE(n10177), .CLK(n10801), 
        .Q(n8336), .QN(n3831) );
  SDFFX1 DFF_1362_Q_reg ( .D(n1715), .SI(n8336), .SE(n10177), .CLK(n10801), 
        .Q(n8335), .QN(n3830) );
  SDFFX1 DFF_1363_Q_reg ( .D(n1716), .SI(n8335), .SE(n10177), .CLK(n10801), 
        .Q(n8334), .QN(n3829) );
  SDFFX1 DFF_1364_Q_reg ( .D(n1717), .SI(n8334), .SE(n10177), .CLK(n10801), 
        .Q(n8333), .QN(n3828) );
  SDFFX1 DFF_1365_Q_reg ( .D(n1718), .SI(n8333), .SE(n10177), .CLK(n10801), 
        .Q(n8332), .QN(n3827) );
  SDFFX1 DFF_1366_Q_reg ( .D(n1719), .SI(n8332), .SE(n10178), .CLK(n10801), 
        .Q(n8331), .QN(n3826) );
  SDFFX1 DFF_1367_Q_reg ( .D(n1720), .SI(n8331), .SE(n10178), .CLK(n10801), 
        .Q(n8330), .QN(n3825) );
  SDFFX1 DFF_1368_Q_reg ( .D(n1721), .SI(n8330), .SE(n10178), .CLK(n10801), 
        .Q(n8329), .QN(n3824) );
  SDFFX1 DFF_1369_Q_reg ( .D(n1722), .SI(n8329), .SE(n10178), .CLK(n10801), 
        .Q(n8328), .QN(n3823) );
  SDFFX1 DFF_1370_Q_reg ( .D(n1723), .SI(n8328), .SE(n10178), .CLK(n10801), 
        .Q(test_so79), .QN(n3822) );
  SDFFX1 DFF_1371_Q_reg ( .D(n1724), .SI(test_si80), .SE(n10178), .CLK(n10800), 
        .Q(n8325), .QN(n3821) );
  SDFFX1 DFF_1372_Q_reg ( .D(n1725), .SI(n8325), .SE(n10179), .CLK(n10800), 
        .Q(n8324), .QN(n3820) );
  SDFFX1 DFF_1373_Q_reg ( .D(n1726), .SI(n8324), .SE(n10179), .CLK(n10800), 
        .Q(n8323), .QN(n3819) );
  SDFFX1 DFF_1374_Q_reg ( .D(n1727), .SI(n8323), .SE(n10179), .CLK(n10800), 
        .Q(n8322), .QN(n3818) );
  SDFFX1 DFF_1375_Q_reg ( .D(WX9597), .SI(n8322), .SE(n10179), .CLK(n10800), 
        .Q(n8321), .QN(n3817) );
  SDFFX1 DFF_1376_Q_reg ( .D(WX9695), .SI(n8321), .SE(n10117), .CLK(n10832), 
        .Q(n8320), .QN(n17895) );
  SDFFX1 DFF_1377_Q_reg ( .D(WX9697), .SI(n8320), .SE(n10174), .CLK(n10803), 
        .Q(n8319), .QN(n17894) );
  SDFFX1 DFF_1378_Q_reg ( .D(WX9699), .SI(n8319), .SE(n10173), .CLK(n10803), 
        .Q(n8318), .QN(n17893) );
  SDFFX1 DFF_1379_Q_reg ( .D(WX9701), .SI(n8318), .SE(n10173), .CLK(n10803), 
        .Q(n8317), .QN(n17892) );
  SDFFX1 DFF_1380_Q_reg ( .D(WX9703), .SI(n8317), .SE(n10173), .CLK(n10803), 
        .Q(n8316), .QN(n17891) );
  SDFFX1 DFF_1381_Q_reg ( .D(WX9705), .SI(n8316), .SE(n10173), .CLK(n10803), 
        .Q(n8315), .QN(n17890) );
  SDFFX1 DFF_1382_Q_reg ( .D(WX9707), .SI(n8315), .SE(n10172), .CLK(n10804), 
        .Q(n8314), .QN(n17889) );
  SDFFX1 DFF_1383_Q_reg ( .D(WX9709), .SI(n8314), .SE(n10172), .CLK(n10804), 
        .Q(n8313), .QN(n17888) );
  SDFFX1 DFF_1384_Q_reg ( .D(WX9711), .SI(n8313), .SE(n10171), .CLK(n10804), 
        .Q(n8312), .QN(n17887) );
  SDFFX1 DFF_1385_Q_reg ( .D(WX9713), .SI(n8312), .SE(n10171), .CLK(n10804), 
        .Q(n8311), .QN(n17886) );
  SDFFX1 DFF_1386_Q_reg ( .D(WX9715), .SI(n8311), .SE(n10171), .CLK(n10804), 
        .Q(n8310), .QN(n17885) );
  SDFFX1 DFF_1387_Q_reg ( .D(WX9717), .SI(n8310), .SE(n10171), .CLK(n10804), 
        .Q(test_so80), .QN(n9890) );
  SDFFX1 DFF_1388_Q_reg ( .D(WX9719), .SI(test_si81), .SE(n10170), .CLK(n10805), .Q(n8307), .QN(n17884) );
  SDFFX1 DFF_1389_Q_reg ( .D(WX9721), .SI(n8307), .SE(n10170), .CLK(n10805), 
        .Q(n8306), .QN(n17883) );
  SDFFX1 DFF_1390_Q_reg ( .D(WX9723), .SI(n8306), .SE(n10169), .CLK(n10805), 
        .Q(n8305), .QN(n17882) );
  SDFFX1 DFF_1391_Q_reg ( .D(WX9725), .SI(n8305), .SE(n10169), .CLK(n10805), 
        .Q(n8304), .QN(n17881) );
  SDFFX1 DFF_1392_Q_reg ( .D(WX9727), .SI(n8304), .SE(n10168), .CLK(n10805), 
        .Q(WX9728), .QN(n9329) );
  SDFFX1 DFF_1393_Q_reg ( .D(WX9729), .SI(WX9728), .SE(n10168), .CLK(n10806), 
        .Q(WX9730) );
  SDFFX1 DFF_1394_Q_reg ( .D(WX9731), .SI(WX9730), .SE(n10167), .CLK(n10806), 
        .Q(WX9732), .QN(n9325) );
  SDFFX1 DFF_1395_Q_reg ( .D(WX9733), .SI(WX9732), .SE(n10167), .CLK(n10806), 
        .Q(WX9734), .QN(n9323) );
  SDFFX1 DFF_1396_Q_reg ( .D(WX9735), .SI(WX9734), .SE(n10336), .CLK(n10722), 
        .Q(WX9736), .QN(n9321) );
  SDFFX1 DFF_1397_Q_reg ( .D(WX9737), .SI(WX9736), .SE(n10165), .CLK(n10807), 
        .Q(WX9738), .QN(n9319) );
  SDFFX1 DFF_1398_Q_reg ( .D(WX9739), .SI(WX9738), .SE(n10165), .CLK(n10807), 
        .Q(WX9740), .QN(n9317) );
  SDFFX1 DFF_1399_Q_reg ( .D(WX9741), .SI(WX9740), .SE(n10164), .CLK(n10808), 
        .Q(WX9742), .QN(n9315) );
  SDFFX1 DFF_1400_Q_reg ( .D(WX9743), .SI(WX9742), .SE(n10164), .CLK(n10808), 
        .Q(WX9744), .QN(n9313) );
  SDFFX1 DFF_1401_Q_reg ( .D(WX9745), .SI(WX9744), .SE(n10163), .CLK(n10808), 
        .Q(WX9746), .QN(n9311) );
  SDFFX1 DFF_1402_Q_reg ( .D(WX9747), .SI(WX9746), .SE(n10162), .CLK(n10809), 
        .Q(WX9748), .QN(n9309) );
  SDFFX1 DFF_1403_Q_reg ( .D(WX9749), .SI(WX9748), .SE(n10162), .CLK(n10809), 
        .Q(WX9750), .QN(n9307) );
  SDFFX1 DFF_1404_Q_reg ( .D(WX9751), .SI(WX9750), .SE(n10161), .CLK(n10809), 
        .Q(test_so81), .QN(n9916) );
  SDFFX1 DFF_1405_Q_reg ( .D(WX9753), .SI(test_si82), .SE(n10160), .CLK(n10810), .Q(WX9754), .QN(n9304) );
  SDFFX1 DFF_1406_Q_reg ( .D(WX9755), .SI(WX9754), .SE(n10160), .CLK(n10810), 
        .Q(WX9756), .QN(n9302) );
  SDFFX1 DFF_1407_Q_reg ( .D(WX9757), .SI(WX9756), .SE(n10159), .CLK(n10810), 
        .Q(WX9758), .QN(n9300) );
  SDFFX1 DFF_1408_Q_reg ( .D(WX9759), .SI(WX9758), .SE(n10158), .CLK(n10811), 
        .Q(WX9760), .QN(n9030) );
  SDFFX1 DFF_1409_Q_reg ( .D(WX9761), .SI(WX9760), .SE(n10174), .CLK(n10803), 
        .Q(WX9762), .QN(n9098) );
  SDFFX1 DFF_1410_Q_reg ( .D(WX9763), .SI(WX9762), .SE(n10174), .CLK(n10803), 
        .Q(WX9764), .QN(n9096) );
  SDFFX1 DFF_1411_Q_reg ( .D(WX9765), .SI(WX9764), .SE(n10173), .CLK(n10803), 
        .Q(WX9766), .QN(n9094) );
  SDFFX1 DFF_1412_Q_reg ( .D(WX9767), .SI(WX9766), .SE(n10173), .CLK(n10803), 
        .Q(WX9768), .QN(n9092) );
  SDFFX1 DFF_1413_Q_reg ( .D(WX9769), .SI(WX9768), .SE(n10172), .CLK(n10803), 
        .Q(WX9770), .QN(n9090) );
  SDFFX1 DFF_1414_Q_reg ( .D(WX9771), .SI(WX9770), .SE(n10172), .CLK(n10804), 
        .Q(WX9772), .QN(n9088) );
  SDFFX1 DFF_1415_Q_reg ( .D(WX9773), .SI(WX9772), .SE(n10172), .CLK(n10804), 
        .Q(WX9774), .QN(n9086) );
  SDFFX1 DFF_1416_Q_reg ( .D(WX9775), .SI(WX9774), .SE(n10172), .CLK(n10804), 
        .Q(WX9776), .QN(n9084) );
  SDFFX1 DFF_1417_Q_reg ( .D(WX9777), .SI(WX9776), .SE(n10171), .CLK(n10804), 
        .Q(WX9778), .QN(n9082) );
  SDFFX1 DFF_1418_Q_reg ( .D(WX9779), .SI(WX9778), .SE(n10171), .CLK(n10804), 
        .Q(WX9780), .QN(n9080) );
  SDFFX1 DFF_1419_Q_reg ( .D(WX9781), .SI(WX9780), .SE(n10170), .CLK(n10804), 
        .Q(WX9782), .QN(n9078) );
  SDFFX1 DFF_1420_Q_reg ( .D(WX9783), .SI(WX9782), .SE(n10170), .CLK(n10805), 
        .Q(WX9784), .QN(n9076) );
  SDFFX1 DFF_1421_Q_reg ( .D(WX9785), .SI(WX9784), .SE(n10170), .CLK(n10805), 
        .Q(test_so82), .QN(n9954) );
  SDFFX1 DFF_1422_Q_reg ( .D(WX9787), .SI(test_si83), .SE(n10169), .CLK(n10805), .Q(WX9788), .QN(n9073) );
  SDFFX1 DFF_1423_Q_reg ( .D(WX9789), .SI(WX9788), .SE(n10169), .CLK(n10805), 
        .Q(WX9790), .QN(n9072) );
  SDFFX1 DFF_1424_Q_reg ( .D(WX9791), .SI(WX9790), .SE(n10168), .CLK(n10806), 
        .Q(WX9792), .QN(n3593) );
  SDFFX1 DFF_1425_Q_reg ( .D(WX9793), .SI(WX9792), .SE(n10168), .CLK(n10806), 
        .Q(WX9794), .QN(n3591) );
  SDFFX1 DFF_1426_Q_reg ( .D(WX9795), .SI(WX9794), .SE(n10167), .CLK(n10806), 
        .Q(WX9796), .QN(n3589) );
  SDFFX1 DFF_1427_Q_reg ( .D(WX9797), .SI(WX9796), .SE(n10167), .CLK(n10806), 
        .Q(WX9798), .QN(n3587) );
  SDFFX1 DFF_1428_Q_reg ( .D(WX9799), .SI(WX9798), .SE(n10166), .CLK(n10807), 
        .Q(WX9800), .QN(n3585) );
  SDFFX1 DFF_1429_Q_reg ( .D(WX9801), .SI(WX9800), .SE(n10166), .CLK(n10807), 
        .Q(WX9802), .QN(n3583) );
  SDFFX1 DFF_1430_Q_reg ( .D(WX9803), .SI(WX9802), .SE(n10165), .CLK(n10807), 
        .Q(WX9804), .QN(n3581) );
  SDFFX1 DFF_1431_Q_reg ( .D(WX9805), .SI(WX9804), .SE(n10164), .CLK(n10808), 
        .Q(WX9806), .QN(n3579) );
  SDFFX1 DFF_1432_Q_reg ( .D(WX9807), .SI(WX9806), .SE(n10163), .CLK(n10808), 
        .Q(WX9808), .QN(n3577) );
  SDFFX1 DFF_1433_Q_reg ( .D(WX9809), .SI(WX9808), .SE(n10163), .CLK(n10808), 
        .Q(WX9810), .QN(n3575) );
  SDFFX1 DFF_1434_Q_reg ( .D(WX9811), .SI(WX9810), .SE(n10162), .CLK(n10809), 
        .Q(WX9812), .QN(n3573) );
  SDFFX1 DFF_1435_Q_reg ( .D(WX9813), .SI(WX9812), .SE(n10161), .CLK(n10809), 
        .Q(WX9814), .QN(n3571) );
  SDFFX1 DFF_1436_Q_reg ( .D(WX9815), .SI(WX9814), .SE(n10161), .CLK(n10809), 
        .Q(WX9816), .QN(n3569) );
  SDFFX1 DFF_1437_Q_reg ( .D(WX9817), .SI(WX9816), .SE(n10160), .CLK(n10810), 
        .Q(WX9818), .QN(n3567) );
  SDFFX1 DFF_1438_Q_reg ( .D(WX9819), .SI(WX9818), .SE(n10159), .CLK(n10810), 
        .Q(test_so83), .QN(n9915) );
  SDFFX1 DFF_1439_Q_reg ( .D(WX9821), .SI(test_si84), .SE(n10159), .CLK(n10810), .Q(WX9822), .QN(n3563) );
  SDFFX1 DFF_1440_Q_reg ( .D(WX9823), .SI(WX9822), .SE(n10158), .CLK(n10811), 
        .Q(WX9824) );
  SDFFX1 DFF_1441_Q_reg ( .D(WX9825), .SI(WX9824), .SE(n10158), .CLK(n10811), 
        .Q(WX9826), .QN(n9099) );
  SDFFX1 DFF_1442_Q_reg ( .D(WX9827), .SI(WX9826), .SE(n10157), .CLK(n10811), 
        .Q(WX9828), .QN(n9097) );
  SDFFX1 DFF_1443_Q_reg ( .D(WX9829), .SI(WX9828), .SE(n10157), .CLK(n10811), 
        .Q(WX9830), .QN(n9095) );
  SDFFX1 DFF_1444_Q_reg ( .D(WX9831), .SI(WX9830), .SE(n10157), .CLK(n10811), 
        .Q(WX9832), .QN(n9093) );
  SDFFX1 DFF_1445_Q_reg ( .D(WX9833), .SI(WX9832), .SE(n10156), .CLK(n10811), 
        .Q(WX9834), .QN(n9091) );
  SDFFX1 DFF_1446_Q_reg ( .D(WX9835), .SI(WX9834), .SE(n10156), .CLK(n10812), 
        .Q(WX9836), .QN(n9089) );
  SDFFX1 DFF_1447_Q_reg ( .D(WX9837), .SI(WX9836), .SE(n10156), .CLK(n10812), 
        .Q(WX9838), .QN(n9087) );
  SDFFX1 DFF_1448_Q_reg ( .D(WX9839), .SI(WX9838), .SE(n10155), .CLK(n10812), 
        .Q(WX9840), .QN(n9085) );
  SDFFX1 DFF_1449_Q_reg ( .D(WX9841), .SI(WX9840), .SE(n10155), .CLK(n10812), 
        .Q(WX9842), .QN(n9083) );
  SDFFX1 DFF_1450_Q_reg ( .D(WX9843), .SI(WX9842), .SE(n10155), .CLK(n10812), 
        .Q(WX9844), .QN(n9081) );
  SDFFX1 DFF_1451_Q_reg ( .D(WX9845), .SI(WX9844), .SE(n10154), .CLK(n10812), 
        .Q(WX9846), .QN(n9079) );
  SDFFX1 DFF_1452_Q_reg ( .D(WX9847), .SI(WX9846), .SE(n10154), .CLK(n10813), 
        .Q(WX9848), .QN(n9077) );
  SDFFX1 DFF_1453_Q_reg ( .D(WX9849), .SI(WX9848), .SE(n10170), .CLK(n10805), 
        .Q(WX9850), .QN(n9075) );
  SDFFX1 DFF_1454_Q_reg ( .D(WX9851), .SI(WX9850), .SE(n10169), .CLK(n10805), 
        .Q(WX9852), .QN(n9074) );
  SDFFX1 DFF_1455_Q_reg ( .D(WX9853), .SI(WX9852), .SE(n10169), .CLK(n10805), 
        .Q(test_so84), .QN(n9953) );
  SDFFX1 DFF_1456_Q_reg ( .D(WX9855), .SI(test_si85), .SE(n10168), .CLK(n10806), .Q(WX9856), .QN(n9330) );
  SDFFX1 DFF_1457_Q_reg ( .D(WX9857), .SI(WX9856), .SE(n10168), .CLK(n10806), 
        .Q(WX9858), .QN(n9328) );
  SDFFX1 DFF_1458_Q_reg ( .D(WX9859), .SI(WX9858), .SE(n10167), .CLK(n10806), 
        .Q(WX9860), .QN(n9326) );
  SDFFX1 DFF_1459_Q_reg ( .D(WX9861), .SI(WX9860), .SE(n10166), .CLK(n10806), 
        .Q(WX9862), .QN(n9324) );
  SDFFX1 DFF_1460_Q_reg ( .D(WX9863), .SI(WX9862), .SE(n10166), .CLK(n10807), 
        .Q(WX9864), .QN(n9322) );
  SDFFX1 DFF_1461_Q_reg ( .D(WX9865), .SI(WX9864), .SE(n10165), .CLK(n10807), 
        .Q(WX9866), .QN(n9320) );
  SDFFX1 DFF_1462_Q_reg ( .D(WX9867), .SI(WX9866), .SE(n10165), .CLK(n10807), 
        .Q(WX9868), .QN(n9318) );
  SDFFX1 DFF_1463_Q_reg ( .D(WX9869), .SI(WX9868), .SE(n10164), .CLK(n10808), 
        .Q(WX9870), .QN(n9316) );
  SDFFX1 DFF_1464_Q_reg ( .D(WX9871), .SI(WX9870), .SE(n10163), .CLK(n10808), 
        .Q(WX9872), .QN(n9314) );
  SDFFX1 DFF_1465_Q_reg ( .D(WX9873), .SI(WX9872), .SE(n10163), .CLK(n10808), 
        .Q(WX9874), .QN(n9312) );
  SDFFX1 DFF_1466_Q_reg ( .D(WX9875), .SI(WX9874), .SE(n10162), .CLK(n10809), 
        .Q(WX9876), .QN(n9310) );
  SDFFX1 DFF_1467_Q_reg ( .D(WX9877), .SI(WX9876), .SE(n10161), .CLK(n10809), 
        .Q(WX9878), .QN(n9308) );
  SDFFX1 DFF_1468_Q_reg ( .D(WX9879), .SI(WX9878), .SE(n10161), .CLK(n10809), 
        .Q(WX9880) );
  SDFFX1 DFF_1469_Q_reg ( .D(WX9881), .SI(WX9880), .SE(n10160), .CLK(n10810), 
        .Q(WX9882), .QN(n9305) );
  SDFFX1 DFF_1470_Q_reg ( .D(WX9883), .SI(WX9882), .SE(n10159), .CLK(n10810), 
        .Q(WX9884) );
  SDFFX1 DFF_1471_Q_reg ( .D(WX9885), .SI(WX9884), .SE(n10159), .CLK(n10810), 
        .Q(WX9886), .QN(n9301) );
  SDFFX1 DFF_1472_Q_reg ( .D(WX9887), .SI(WX9886), .SE(n10158), .CLK(n10811), 
        .Q(test_so85), .QN(n9914) );
  SDFFX1 DFF_1473_Q_reg ( .D(WX9889), .SI(test_si86), .SE(n10158), .CLK(n10811), .Q(WX9890), .QN(n9567) );
  SDFFX1 DFF_1474_Q_reg ( .D(WX9891), .SI(WX9890), .SE(n10157), .CLK(n10811), 
        .Q(WX9892), .QN(n9568) );
  SDFFX1 DFF_1475_Q_reg ( .D(WX9893), .SI(WX9892), .SE(n10157), .CLK(n10811), 
        .Q(WX9894), .QN(n9569) );
  SDFFX1 DFF_1476_Q_reg ( .D(WX9895), .SI(WX9894), .SE(n10157), .CLK(n10811), 
        .Q(WX9896), .QN(n9570) );
  SDFFX1 DFF_1477_Q_reg ( .D(WX9897), .SI(WX9896), .SE(n10156), .CLK(n10812), 
        .Q(WX9898), .QN(n9571) );
  SDFFX1 DFF_1478_Q_reg ( .D(WX9899), .SI(WX9898), .SE(n10156), .CLK(n10812), 
        .Q(WX9900), .QN(n9572) );
  SDFFX1 DFF_1479_Q_reg ( .D(WX9901), .SI(WX9900), .SE(n10156), .CLK(n10812), 
        .Q(WX9902), .QN(n9573) );
  SDFFX1 DFF_1480_Q_reg ( .D(WX9903), .SI(WX9902), .SE(n10155), .CLK(n10812), 
        .Q(WX9904), .QN(n9574) );
  SDFFX1 DFF_1481_Q_reg ( .D(WX9905), .SI(WX9904), .SE(n10155), .CLK(n10812), 
        .Q(WX9906), .QN(n9575) );
  SDFFX1 DFF_1482_Q_reg ( .D(WX9907), .SI(WX9906), .SE(n10155), .CLK(n10812), 
        .Q(WX9908), .QN(n9576) );
  SDFFX1 DFF_1483_Q_reg ( .D(WX9909), .SI(WX9908), .SE(n10154), .CLK(n10813), 
        .Q(WX9910), .QN(n9577) );
  SDFFX1 DFF_1484_Q_reg ( .D(WX9911), .SI(WX9910), .SE(n10154), .CLK(n10813), 
        .Q(WX9912), .QN(n9578) );
  SDFFX1 DFF_1485_Q_reg ( .D(WX9913), .SI(WX9912), .SE(n10154), .CLK(n10813), 
        .Q(WX9914), .QN(n9579) );
  SDFFX1 DFF_1486_Q_reg ( .D(WX9915), .SI(WX9914), .SE(n10154), .CLK(n10813), 
        .Q(WX9916), .QN(n9580) );
  SDFFX1 DFF_1487_Q_reg ( .D(WX9917), .SI(WX9916), .SE(n10153), .CLK(n10813), 
        .Q(WX9918), .QN(n9515) );
  SDFFX1 DFF_1488_Q_reg ( .D(WX9919), .SI(WX9918), .SE(n10153), .CLK(n10813), 
        .Q(WX9920), .QN(n9581) );
  SDFFX1 DFF_1489_Q_reg ( .D(WX9921), .SI(WX9920), .SE(n10153), .CLK(n10813), 
        .Q(test_so86), .QN(n9907) );
  SDFFX1 DFF_1490_Q_reg ( .D(WX9923), .SI(test_si87), .SE(n10167), .CLK(n10806), .Q(WX9924), .QN(n9582) );
  SDFFX1 DFF_1491_Q_reg ( .D(WX9925), .SI(WX9924), .SE(n10166), .CLK(n10807), 
        .Q(WX9926), .QN(n9583) );
  SDFFX1 DFF_1492_Q_reg ( .D(WX9927), .SI(WX9926), .SE(n10166), .CLK(n10807), 
        .Q(WX9928), .QN(n9516) );
  SDFFX1 DFF_1493_Q_reg ( .D(WX9929), .SI(WX9928), .SE(n10165), .CLK(n10807), 
        .Q(WX9930), .QN(n9584) );
  SDFFX1 DFF_1494_Q_reg ( .D(WX9931), .SI(WX9930), .SE(n10164), .CLK(n10807), 
        .Q(WX9932), .QN(n9585) );
  SDFFX1 DFF_1495_Q_reg ( .D(WX9933), .SI(WX9932), .SE(n10164), .CLK(n10808), 
        .Q(WX9934), .QN(n9586) );
  SDFFX1 DFF_1496_Q_reg ( .D(WX9935), .SI(WX9934), .SE(n10163), .CLK(n10808), 
        .Q(WX9936), .QN(n9587) );
  SDFFX1 DFF_1497_Q_reg ( .D(WX9937), .SI(WX9936), .SE(n10162), .CLK(n10808), 
        .Q(WX9938), .QN(n9588) );
  SDFFX1 DFF_1498_Q_reg ( .D(WX9939), .SI(WX9938), .SE(n10162), .CLK(n10809), 
        .Q(WX9940), .QN(n9589) );
  SDFFX1 DFF_1499_Q_reg ( .D(WX9941), .SI(WX9940), .SE(n10161), .CLK(n10809), 
        .Q(WX9942), .QN(n9517) );
  SDFFX1 DFF_1500_Q_reg ( .D(WX9943), .SI(WX9942), .SE(n10160), .CLK(n10809), 
        .Q(WX9944), .QN(n9590) );
  SDFFX1 DFF_1501_Q_reg ( .D(WX9945), .SI(WX9944), .SE(n10160), .CLK(n10810), 
        .Q(WX9946), .QN(n9591) );
  SDFFX1 DFF_1502_Q_reg ( .D(WX9947), .SI(WX9946), .SE(n10159), .CLK(n10810), 
        .Q(WX9948), .QN(n9592) );
  SDFFX1 DFF_1503_Q_reg ( .D(WX9949), .SI(WX9948), .SE(n10158), .CLK(n10810), 
        .Q(WX9950), .QN(n9534) );
  SDFFX1 DFF_1504_Q_reg ( .D(WX10315), .SI(WX9950), .SE(n10120), .CLK(n10830), 
        .Q(CRC_OUT_2_0), .QN(DFF_1504_n1) );
  SDFFX1 DFF_1505_Q_reg ( .D(WX10317), .SI(CRC_OUT_2_0), .SE(n10120), .CLK(
        n10830), .Q(CRC_OUT_2_1), .QN(DFF_1505_n1) );
  SDFFX1 DFF_1506_Q_reg ( .D(WX10319), .SI(CRC_OUT_2_1), .SE(n10120), .CLK(
        n10830), .Q(test_so87), .QN(n9952) );
  SDFFX1 DFF_1507_Q_reg ( .D(WX10321), .SI(test_si88), .SE(n10120), .CLK(
        n10830), .Q(CRC_OUT_2_3), .QN(DFF_1507_n1) );
  SDFFX1 DFF_1508_Q_reg ( .D(WX10323), .SI(CRC_OUT_2_3), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_4), .QN(DFF_1508_n1) );
  SDFFX1 DFF_1509_Q_reg ( .D(WX10325), .SI(CRC_OUT_2_4), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_5), .QN(DFF_1509_n1) );
  SDFFX1 DFF_1510_Q_reg ( .D(WX10327), .SI(CRC_OUT_2_5), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_6), .QN(DFF_1510_n1) );
  SDFFX1 DFF_1511_Q_reg ( .D(WX10329), .SI(CRC_OUT_2_6), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_7), .QN(DFF_1511_n1) );
  SDFFX1 DFF_1512_Q_reg ( .D(WX10331), .SI(CRC_OUT_2_7), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_8), .QN(DFF_1512_n1) );
  SDFFX1 DFF_1513_Q_reg ( .D(WX10333), .SI(CRC_OUT_2_8), .SE(n10119), .CLK(
        n10831), .Q(CRC_OUT_2_9), .QN(DFF_1513_n1) );
  SDFFX1 DFF_1514_Q_reg ( .D(WX10335), .SI(CRC_OUT_2_9), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_10), .QN(DFF_1514_n1) );
  SDFFX1 DFF_1515_Q_reg ( .D(WX10337), .SI(CRC_OUT_2_10), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_11), .QN(DFF_1515_n1) );
  SDFFX1 DFF_1516_Q_reg ( .D(WX10339), .SI(CRC_OUT_2_11), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_12), .QN(DFF_1516_n1) );
  SDFFX1 DFF_1517_Q_reg ( .D(WX10341), .SI(CRC_OUT_2_12), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_13), .QN(DFF_1517_n1) );
  SDFFX1 DFF_1518_Q_reg ( .D(WX10343), .SI(CRC_OUT_2_13), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_14), .QN(DFF_1518_n1) );
  SDFFX1 DFF_1519_Q_reg ( .D(WX10345), .SI(CRC_OUT_2_14), .SE(n10118), .CLK(
        n10831), .Q(CRC_OUT_2_15), .QN(DFF_1519_n1) );
  SDFFX1 DFF_1520_Q_reg ( .D(WX10347), .SI(CRC_OUT_2_15), .SE(n10117), .CLK(
        n10832), .Q(CRC_OUT_2_16), .QN(DFF_1520_n1) );
  SDFFX1 DFF_1521_Q_reg ( .D(WX10349), .SI(CRC_OUT_2_16), .SE(n10117), .CLK(
        n10832), .Q(CRC_OUT_2_17), .QN(DFF_1521_n1) );
  SDFFX1 DFF_1522_Q_reg ( .D(WX10351), .SI(CRC_OUT_2_17), .SE(n10117), .CLK(
        n10832), .Q(CRC_OUT_2_18), .QN(DFF_1522_n1) );
  SDFFX1 DFF_1523_Q_reg ( .D(WX10353), .SI(CRC_OUT_2_18), .SE(n10153), .CLK(
        n10813), .Q(test_so88), .QN(n9951) );
  SDFFX1 DFF_1524_Q_reg ( .D(WX10355), .SI(test_si89), .SE(n10153), .CLK(
        n10813), .Q(CRC_OUT_2_20), .QN(DFF_1524_n1) );
  SDFFX1 DFF_1525_Q_reg ( .D(WX10357), .SI(CRC_OUT_2_20), .SE(n10153), .CLK(
        n10813), .Q(CRC_OUT_2_21), .QN(DFF_1525_n1) );
  SDFFX1 DFF_1526_Q_reg ( .D(WX10359), .SI(CRC_OUT_2_21), .SE(n10152), .CLK(
        n10813), .Q(CRC_OUT_2_22), .QN(DFF_1526_n1) );
  SDFFX1 DFF_1527_Q_reg ( .D(WX10361), .SI(CRC_OUT_2_22), .SE(n10152), .CLK(
        n10814), .Q(CRC_OUT_2_23), .QN(DFF_1527_n1) );
  SDFFX1 DFF_1528_Q_reg ( .D(WX10363), .SI(CRC_OUT_2_23), .SE(n10152), .CLK(
        n10814), .Q(CRC_OUT_2_24), .QN(DFF_1528_n1) );
  SDFFX1 DFF_1529_Q_reg ( .D(WX10365), .SI(CRC_OUT_2_24), .SE(n10152), .CLK(
        n10814), .Q(CRC_OUT_2_25), .QN(DFF_1529_n1) );
  SDFFX1 DFF_1530_Q_reg ( .D(WX10367), .SI(CRC_OUT_2_25), .SE(n10152), .CLK(
        n10814), .Q(CRC_OUT_2_26), .QN(DFF_1530_n1) );
  SDFFX1 DFF_1531_Q_reg ( .D(WX10369), .SI(CRC_OUT_2_26), .SE(n10152), .CLK(
        n10814), .Q(CRC_OUT_2_27), .QN(DFF_1531_n1) );
  SDFFX1 DFF_1532_Q_reg ( .D(WX10371), .SI(CRC_OUT_2_27), .SE(n10151), .CLK(
        n10814), .Q(CRC_OUT_2_28), .QN(DFF_1532_n1) );
  SDFFX1 DFF_1533_Q_reg ( .D(WX10373), .SI(CRC_OUT_2_28), .SE(n10151), .CLK(
        n10814), .Q(CRC_OUT_2_29), .QN(DFF_1533_n1) );
  SDFFX1 DFF_1534_Q_reg ( .D(WX10375), .SI(CRC_OUT_2_29), .SE(n10151), .CLK(
        n10814), .Q(CRC_OUT_2_30), .QN(DFF_1534_n1) );
  SDFFX1 DFF_1535_Q_reg ( .D(WX10377), .SI(CRC_OUT_2_30), .SE(n10151), .CLK(
        n10814), .Q(CRC_OUT_2_31), .QN(DFF_1535_n1) );
  SDFFX1 DFF_1536_Q_reg ( .D(n1938), .SI(CRC_OUT_2_31), .SE(n10151), .CLK(
        n10814), .Q(WX10829), .QN(n9851) );
  SDFFX1 DFF_1537_Q_reg ( .D(n1939), .SI(WX10829), .SE(n10146), .CLK(n10817), 
        .Q(n8295), .QN(n3816) );
  SDFFX1 DFF_1538_Q_reg ( .D(n1940), .SI(n8295), .SE(n10146), .CLK(n10817), 
        .Q(n8294), .QN(n3815) );
  SDFFX1 DFF_1539_Q_reg ( .D(n1941), .SI(n8294), .SE(n10146), .CLK(n10817), 
        .Q(n8293), .QN(n3814) );
  SDFFX1 DFF_1540_Q_reg ( .D(n1942), .SI(n8293), .SE(n10146), .CLK(n10817), 
        .Q(test_so89), .QN(n3813) );
  SDFFX1 DFF_1541_Q_reg ( .D(n1943), .SI(test_si90), .SE(n10146), .CLK(n10817), 
        .Q(n8290), .QN(n3812) );
  SDFFX1 DFF_1542_Q_reg ( .D(n1944), .SI(n8290), .SE(n10146), .CLK(n10816), 
        .Q(n8289), .QN(n3811) );
  SDFFX1 DFF_1543_Q_reg ( .D(n1945), .SI(n8289), .SE(n10147), .CLK(n10816), 
        .Q(n8288), .QN(n3810) );
  SDFFX1 DFF_1544_Q_reg ( .D(n1946), .SI(n8288), .SE(n10147), .CLK(n10816), 
        .Q(n8287), .QN(n3809) );
  SDFFX1 DFF_1545_Q_reg ( .D(n1947), .SI(n8287), .SE(n10147), .CLK(n10816), 
        .Q(n8286), .QN(n3808) );
  SDFFX1 DFF_1546_Q_reg ( .D(n1948), .SI(n8286), .SE(n10147), .CLK(n10816), 
        .Q(n8285), .QN(n3807) );
  SDFFX1 DFF_1547_Q_reg ( .D(n1949), .SI(n8285), .SE(n10147), .CLK(n10816), 
        .Q(n8284), .QN(n3806) );
  SDFFX1 DFF_1548_Q_reg ( .D(n1950), .SI(n8284), .SE(n10147), .CLK(n10816), 
        .Q(n8283), .QN(n3805) );
  SDFFX1 DFF_1549_Q_reg ( .D(n1951), .SI(n8283), .SE(n10148), .CLK(n10816), 
        .Q(n8282), .QN(n3804) );
  SDFFX1 DFF_1550_Q_reg ( .D(n1952), .SI(n8282), .SE(n10148), .CLK(n10816), 
        .Q(n8281), .QN(n3803) );
  SDFFX1 DFF_1551_Q_reg ( .D(n1953), .SI(n8281), .SE(n10148), .CLK(n10816), 
        .Q(n8280), .QN(n3802) );
  SDFFX1 DFF_1552_Q_reg ( .D(n1954), .SI(n8280), .SE(n10148), .CLK(n10816), 
        .Q(n8279), .QN(n3801) );
  SDFFX1 DFF_1553_Q_reg ( .D(n1955), .SI(n8279), .SE(n10148), .CLK(n10816), 
        .Q(n8278), .QN(n3800) );
  SDFFX1 DFF_1554_Q_reg ( .D(n1956), .SI(n8278), .SE(n10148), .CLK(n10815), 
        .Q(n8277), .QN(n3799) );
  SDFFX1 DFF_1555_Q_reg ( .D(n1957), .SI(n8277), .SE(n10149), .CLK(n10815), 
        .Q(n8276), .QN(n3798) );
  SDFFX1 DFF_1556_Q_reg ( .D(n1958), .SI(n8276), .SE(n10149), .CLK(n10815), 
        .Q(n8275), .QN(n3797) );
  SDFFX1 DFF_1557_Q_reg ( .D(n1959), .SI(n8275), .SE(n10149), .CLK(n10815), 
        .Q(test_so90), .QN(n3796) );
  SDFFX1 DFF_1558_Q_reg ( .D(n1960), .SI(test_si91), .SE(n10149), .CLK(n10815), 
        .Q(n8272), .QN(n3795) );
  SDFFX1 DFF_1559_Q_reg ( .D(n1961), .SI(n8272), .SE(n10149), .CLK(n10815), 
        .Q(n8271), .QN(n3794) );
  SDFFX1 DFF_1560_Q_reg ( .D(n1962), .SI(n8271), .SE(n10149), .CLK(n10815), 
        .Q(n8270), .QN(n3793) );
  SDFFX1 DFF_1561_Q_reg ( .D(n1963), .SI(n8270), .SE(n10150), .CLK(n10815), 
        .Q(n8269), .QN(n3792) );
  SDFFX1 DFF_1562_Q_reg ( .D(n1964), .SI(n8269), .SE(n10150), .CLK(n10815), 
        .Q(n8268), .QN(n3791) );
  SDFFX1 DFF_1563_Q_reg ( .D(n1965), .SI(n8268), .SE(n10150), .CLK(n10815), 
        .Q(n8267), .QN(n3790) );
  SDFFX1 DFF_1564_Q_reg ( .D(n1966), .SI(n8267), .SE(n10150), .CLK(n10815), 
        .Q(n8266), .QN(n3789) );
  SDFFX1 DFF_1565_Q_reg ( .D(n1967), .SI(n8266), .SE(n10150), .CLK(n10815), 
        .Q(n8265), .QN(n3788) );
  SDFFX1 DFF_1566_Q_reg ( .D(n1968), .SI(n8265), .SE(n10150), .CLK(n10814), 
        .Q(n8264), .QN(n3787) );
  SDFFX1 DFF_1567_Q_reg ( .D(WX10890), .SI(n8264), .SE(n10151), .CLK(n10814), 
        .Q(n8263), .QN(n3786) );
  SDFFX1 DFF_1568_Q_reg ( .D(WX10988), .SI(n8263), .SE(n10120), .CLK(n10830), 
        .Q(n8262), .QN(n18001) );
  SDFFX1 DFF_1569_Q_reg ( .D(WX10990), .SI(n8262), .SE(n10145), .CLK(n10817), 
        .Q(n8261), .QN(n18000) );
  SDFFX1 DFF_1570_Q_reg ( .D(WX10992), .SI(n8261), .SE(n10145), .CLK(n10817), 
        .Q(n8260), .QN(n17999) );
  SDFFX1 DFF_1571_Q_reg ( .D(WX10994), .SI(n8260), .SE(n10145), .CLK(n10817), 
        .Q(n8259), .QN(n17998) );
  SDFFX1 DFF_1572_Q_reg ( .D(WX10996), .SI(n8259), .SE(n10144), .CLK(n10818), 
        .Q(n8258), .QN(n17997) );
  SDFFX1 DFF_1573_Q_reg ( .D(WX10998), .SI(n8258), .SE(n10144), .CLK(n10818), 
        .Q(n8257), .QN(n17996) );
  SDFFX1 DFF_1574_Q_reg ( .D(WX11000), .SI(n8257), .SE(n10120), .CLK(n10830), 
        .Q(test_so91), .QN(n9896) );
  SDFFX1 DFF_1575_Q_reg ( .D(WX11002), .SI(test_si92), .SE(n10143), .CLK(
        n10818), .Q(n8254), .QN(n17995) );
  SDFFX1 DFF_1576_Q_reg ( .D(WX11004), .SI(n8254), .SE(n10143), .CLK(n10818), 
        .Q(n8253), .QN(n17994) );
  SDFFX1 DFF_1577_Q_reg ( .D(WX11006), .SI(n8253), .SE(n10143), .CLK(n10818), 
        .Q(n8252), .QN(n17993) );
  SDFFX1 DFF_1578_Q_reg ( .D(WX11008), .SI(n8252), .SE(n10142), .CLK(n10819), 
        .Q(n8251), .QN(n17992) );
  SDFFX1 DFF_1579_Q_reg ( .D(WX11010), .SI(n8251), .SE(n10142), .CLK(n10819), 
        .Q(n8250), .QN(n17991) );
  SDFFX1 DFF_1580_Q_reg ( .D(WX11012), .SI(n8250), .SE(n10141), .CLK(n10819), 
        .Q(n8249), .QN(n17990) );
  SDFFX1 DFF_1581_Q_reg ( .D(WX11014), .SI(n8249), .SE(n10141), .CLK(n10819), 
        .Q(n8248), .QN(n17989) );
  SDFFX1 DFF_1582_Q_reg ( .D(WX11016), .SI(n8248), .SE(n10140), .CLK(n10820), 
        .Q(n8247), .QN(n17988) );
  SDFFX1 DFF_1583_Q_reg ( .D(WX11018), .SI(n8247), .SE(n10139), .CLK(n10820), 
        .Q(n8246), .QN(n17987) );
  SDFFX1 DFF_1584_Q_reg ( .D(WX11020), .SI(n8246), .SE(n10138), .CLK(n10821), 
        .Q(WX11021), .QN(n9298) );
  SDFFX1 DFF_1585_Q_reg ( .D(WX11022), .SI(WX11021), .SE(n10138), .CLK(n10821), 
        .Q(WX11023), .QN(n9296) );
  SDFFX1 DFF_1586_Q_reg ( .D(WX11024), .SI(WX11023), .SE(n10137), .CLK(n10821), 
        .Q(WX11025), .QN(n9294) );
  SDFFX1 DFF_1587_Q_reg ( .D(WX11026), .SI(WX11025), .SE(n10137), .CLK(n10821), 
        .Q(WX11027), .QN(n9292) );
  SDFFX1 DFF_1588_Q_reg ( .D(WX11028), .SI(WX11027), .SE(n10136), .CLK(n10822), 
        .Q(WX11029), .QN(n9290) );
  SDFFX1 DFF_1589_Q_reg ( .D(WX11030), .SI(WX11029), .SE(n10136), .CLK(n10822), 
        .Q(WX11031), .QN(n9288) );
  SDFFX1 DFF_1590_Q_reg ( .D(WX11032), .SI(WX11031), .SE(n10135), .CLK(n10822), 
        .Q(WX11033), .QN(n9286) );
  SDFFX1 DFF_1591_Q_reg ( .D(WX11034), .SI(WX11033), .SE(n10135), .CLK(n10823), 
        .Q(test_so92), .QN(n9936) );
  SDFFX1 DFF_1592_Q_reg ( .D(WX11036), .SI(test_si93), .SE(n10134), .CLK(
        n10823), .Q(WX11037), .QN(n9283) );
  SDFFX1 DFF_1593_Q_reg ( .D(WX11038), .SI(WX11037), .SE(n10134), .CLK(n10823), 
        .Q(WX11039), .QN(n9281) );
  SDFFX1 DFF_1594_Q_reg ( .D(WX11040), .SI(WX11039), .SE(n10133), .CLK(n10824), 
        .Q(WX11041), .QN(n9279) );
  SDFFX1 DFF_1595_Q_reg ( .D(WX11042), .SI(WX11041), .SE(n10133), .CLK(n10824), 
        .Q(WX11043) );
  SDFFX1 DFF_1596_Q_reg ( .D(WX11044), .SI(WX11043), .SE(n10132), .CLK(n10824), 
        .Q(WX11045), .QN(n9276) );
  SDFFX1 DFF_1597_Q_reg ( .D(WX11046), .SI(WX11045), .SE(n10131), .CLK(n10825), 
        .Q(WX11047) );
  SDFFX1 DFF_1598_Q_reg ( .D(WX11048), .SI(WX11047), .SE(n10131), .CLK(n10825), 
        .Q(WX11049), .QN(n9272) );
  SDFFX1 DFF_1599_Q_reg ( .D(WX11050), .SI(WX11049), .SE(n10130), .CLK(n10825), 
        .Q(WX11051), .QN(n9270) );
  SDFFX1 DFF_1600_Q_reg ( .D(WX11052), .SI(WX11051), .SE(n10129), .CLK(n10826), 
        .Q(WX11053), .QN(n9028) );
  SDFFX1 DFF_1601_Q_reg ( .D(WX11054), .SI(WX11053), .SE(n10145), .CLK(n10817), 
        .Q(WX11055), .QN(n9070) );
  SDFFX1 DFF_1602_Q_reg ( .D(WX11056), .SI(WX11055), .SE(n10145), .CLK(n10817), 
        .Q(WX11057), .QN(n9068) );
  SDFFX1 DFF_1603_Q_reg ( .D(WX11058), .SI(WX11057), .SE(n10145), .CLK(n10817), 
        .Q(WX11059), .QN(n9066) );
  SDFFX1 DFF_1604_Q_reg ( .D(WX11060), .SI(WX11059), .SE(n10144), .CLK(n10817), 
        .Q(WX11061), .QN(n9064) );
  SDFFX1 DFF_1605_Q_reg ( .D(WX11062), .SI(WX11061), .SE(n10144), .CLK(n10818), 
        .Q(WX11063), .QN(n9062) );
  SDFFX1 DFF_1606_Q_reg ( .D(WX11064), .SI(WX11063), .SE(n10144), .CLK(n10818), 
        .Q(WX11065), .QN(n9060) );
  SDFFX1 DFF_1607_Q_reg ( .D(WX11066), .SI(WX11065), .SE(n10144), .CLK(n10818), 
        .Q(WX11067), .QN(n9058) );
  SDFFX1 DFF_1608_Q_reg ( .D(WX11068), .SI(WX11067), .SE(n10143), .CLK(n10818), 
        .Q(test_so93), .QN(n9966) );
  SDFFX1 DFF_1609_Q_reg ( .D(WX11070), .SI(test_si94), .SE(n10142), .CLK(
        n10818), .Q(WX11071), .QN(n9055) );
  SDFFX1 DFF_1610_Q_reg ( .D(WX11072), .SI(WX11071), .SE(n10142), .CLK(n10819), 
        .Q(WX11073), .QN(n9054) );
  SDFFX1 DFF_1611_Q_reg ( .D(WX11074), .SI(WX11073), .SE(n10142), .CLK(n10819), 
        .Q(WX11075), .QN(n9052) );
  SDFFX1 DFF_1612_Q_reg ( .D(WX11076), .SI(WX11075), .SE(n10141), .CLK(n10819), 
        .Q(WX11077), .QN(n9050) );
  SDFFX1 DFF_1613_Q_reg ( .D(WX11078), .SI(WX11077), .SE(n10141), .CLK(n10819), 
        .Q(WX11079), .QN(n9048) );
  SDFFX1 DFF_1614_Q_reg ( .D(WX11080), .SI(WX11079), .SE(n10140), .CLK(n10820), 
        .Q(WX11081), .QN(n9046) );
  SDFFX1 DFF_1615_Q_reg ( .D(WX11082), .SI(WX11081), .SE(n10139), .CLK(n10820), 
        .Q(WX11083), .QN(n9044) );
  SDFFX1 DFF_1616_Q_reg ( .D(WX11084), .SI(WX11083), .SE(n10139), .CLK(n10820), 
        .Q(WX11085), .QN(n3561) );
  SDFFX1 DFF_1617_Q_reg ( .D(WX11086), .SI(WX11085), .SE(n10138), .CLK(n10821), 
        .Q(WX11087), .QN(n3559) );
  SDFFX1 DFF_1618_Q_reg ( .D(WX11088), .SI(WX11087), .SE(n10137), .CLK(n10821), 
        .Q(WX11089), .QN(n3557) );
  SDFFX1 DFF_1619_Q_reg ( .D(WX11090), .SI(WX11089), .SE(n10137), .CLK(n10821), 
        .Q(WX11091), .QN(n3555) );
  SDFFX1 DFF_1620_Q_reg ( .D(WX11092), .SI(WX11091), .SE(n10136), .CLK(n10822), 
        .Q(WX11093), .QN(n3553) );
  SDFFX1 DFF_1621_Q_reg ( .D(WX11094), .SI(WX11093), .SE(n10135), .CLK(n10822), 
        .Q(WX11095), .QN(n3551) );
  SDFFX1 DFF_1622_Q_reg ( .D(WX11096), .SI(WX11095), .SE(n10135), .CLK(n10822), 
        .Q(WX11097), .QN(n3549) );
  SDFFX1 DFF_1623_Q_reg ( .D(WX11098), .SI(WX11097), .SE(n10134), .CLK(n10823), 
        .Q(WX11099), .QN(n3547) );
  SDFFX1 DFF_1624_Q_reg ( .D(WX11100), .SI(WX11099), .SE(n10134), .CLK(n10823), 
        .Q(WX11101), .QN(n3545) );
  SDFFX1 DFF_1625_Q_reg ( .D(WX11102), .SI(WX11101), .SE(n10133), .CLK(n10823), 
        .Q(test_so94), .QN(n9935) );
  SDFFX1 DFF_1626_Q_reg ( .D(WX11104), .SI(test_si95), .SE(n10133), .CLK(
        n10824), .Q(WX11105), .QN(n3541) );
  SDFFX1 DFF_1627_Q_reg ( .D(WX11106), .SI(WX11105), .SE(n10132), .CLK(n10824), 
        .Q(WX11107), .QN(n3539) );
  SDFFX1 DFF_1628_Q_reg ( .D(WX11108), .SI(WX11107), .SE(n10132), .CLK(n10824), 
        .Q(WX11109), .QN(n3537) );
  SDFFX1 DFF_1629_Q_reg ( .D(WX11110), .SI(WX11109), .SE(n10131), .CLK(n10825), 
        .Q(WX11111), .QN(n3535) );
  SDFFX1 DFF_1630_Q_reg ( .D(WX11112), .SI(WX11111), .SE(n10131), .CLK(n10825), 
        .Q(WX11113), .QN(n3533) );
  SDFFX1 DFF_1631_Q_reg ( .D(WX11114), .SI(WX11113), .SE(n10130), .CLK(n10825), 
        .Q(WX11115), .QN(n3531) );
  SDFFX1 DFF_1632_Q_reg ( .D(WX11116), .SI(WX11115), .SE(n10129), .CLK(n10826), 
        .Q(WX11117), .QN(n9029) );
  SDFFX1 DFF_1633_Q_reg ( .D(WX11118), .SI(WX11117), .SE(n10129), .CLK(n10826), 
        .Q(WX11119), .QN(n9071) );
  SDFFX1 DFF_1634_Q_reg ( .D(WX11120), .SI(WX11119), .SE(n10129), .CLK(n10826), 
        .Q(WX11121), .QN(n9069) );
  SDFFX1 DFF_1635_Q_reg ( .D(WX11122), .SI(WX11121), .SE(n10128), .CLK(n10826), 
        .Q(WX11123), .QN(n9067) );
  SDFFX1 DFF_1636_Q_reg ( .D(WX11124), .SI(WX11123), .SE(n10128), .CLK(n10826), 
        .Q(WX11125), .QN(n9065) );
  SDFFX1 DFF_1637_Q_reg ( .D(WX11126), .SI(WX11125), .SE(n10128), .CLK(n10826), 
        .Q(WX11127), .QN(n9063) );
  SDFFX1 DFF_1638_Q_reg ( .D(WX11128), .SI(WX11127), .SE(n10127), .CLK(n10827), 
        .Q(WX11129), .QN(n9061) );
  SDFFX1 DFF_1639_Q_reg ( .D(WX11130), .SI(WX11129), .SE(n10127), .CLK(n10827), 
        .Q(WX11131), .QN(n9059) );
  SDFFX1 DFF_1640_Q_reg ( .D(WX11132), .SI(WX11131), .SE(n10143), .CLK(n10818), 
        .Q(WX11133), .QN(n9057) );
  SDFFX1 DFF_1641_Q_reg ( .D(WX11134), .SI(WX11133), .SE(n10143), .CLK(n10818), 
        .Q(WX11135), .QN(n9056) );
  SDFFX1 DFF_1642_Q_reg ( .D(WX11136), .SI(WX11135), .SE(n10142), .CLK(n10819), 
        .Q(test_so95), .QN(n9965) );
  SDFFX1 DFF_1643_Q_reg ( .D(WX11138), .SI(test_si96), .SE(n10141), .CLK(
        n10819), .Q(WX11139), .QN(n9053) );
  SDFFX1 DFF_1644_Q_reg ( .D(WX11140), .SI(WX11139), .SE(n10141), .CLK(n10819), 
        .Q(WX11141) );
  SDFFX1 DFF_1645_Q_reg ( .D(WX11142), .SI(WX11141), .SE(n10140), .CLK(n10819), 
        .Q(WX11143), .QN(n9049) );
  SDFFX1 DFF_1646_Q_reg ( .D(WX11144), .SI(WX11143), .SE(n10140), .CLK(n10820), 
        .Q(WX11145), .QN(n9047) );
  SDFFX1 DFF_1647_Q_reg ( .D(WX11146), .SI(WX11145), .SE(n10139), .CLK(n10820), 
        .Q(WX11147), .QN(n9045) );
  SDFFX1 DFF_1648_Q_reg ( .D(WX11148), .SI(WX11147), .SE(n10139), .CLK(n10820), 
        .Q(WX11149), .QN(n9299) );
  SDFFX1 DFF_1649_Q_reg ( .D(WX11150), .SI(WX11149), .SE(n10138), .CLK(n10821), 
        .Q(WX11151), .QN(n9297) );
  SDFFX1 DFF_1650_Q_reg ( .D(WX11152), .SI(WX11151), .SE(n10137), .CLK(n10821), 
        .Q(WX11153), .QN(n9295) );
  SDFFX1 DFF_1651_Q_reg ( .D(WX11154), .SI(WX11153), .SE(n10136), .CLK(n10821), 
        .Q(WX11155), .QN(n9293) );
  SDFFX1 DFF_1652_Q_reg ( .D(WX11156), .SI(WX11155_Tj_Payload), .SE(
        test_se_Trojan), .CLK(n10722), .Q(WX11157), .QN(n9291) );
  SDFFX1 DFF_1653_Q_reg ( .D(WX11158), .SI(WX11157), .SE(test_se_Trojan), 
        .CLK(n10822), .Q(WX11159), .QN(n9289) );
  SDFFX1 DFF_1654_Q_reg ( .D(WX11160), .SI(WX11159), .SE(test_se_Trojan), 
        .CLK(n10822), .Q(WX11161), .QN(n9287) );
  SDFFX1 DFF_1655_Q_reg ( .D(WX11162), .SI(WX11161), .SE(test_se_Trojan), 
        .CLK(n10823), .Q(WX11163) );
  SDFFX1 DFF_1656_Q_reg ( .D(WX11164), .SI(WX11163), .SE(test_se_Trojan), 
        .CLK(n10823), .Q(WX11165), .QN(n9284) );
  SDFFX1 DFF_1657_Q_reg ( .D(WX11166), .SI(WX11165), .SE(test_se_Trojan), 
        .CLK(n10823), .Q(WX11167) );
  SDFFX1 DFF_1658_Q_reg ( .D(WX11168), .SI(WX11167), .SE(test_se_Trojan), 
        .CLK(n10824), .Q(WX11169), .QN(n9280) );
  SDFFX1 DFF_1659_Q_reg ( .D(WX11170), .SI(WX11169), .SE(test_se_Trojan), 
        .CLK(n10824), .Q(test_so96), .QN(n9934) );
  SDFFX1 DFF_1660_Q_reg ( .D(WX11172), .SI(test_si97), .SE(n10132), .CLK(
        n10824), .Q(WX11173), .QN(n9277) );
  SDFFX1 DFF_1661_Q_reg ( .D(WX11174), .SI(WX11173), .SE(n10131), .CLK(n10825), 
        .Q(WX11175), .QN(n9275) );
  SDFFX1 DFF_1662_Q_reg ( .D(WX11176), .SI(WX11175), .SE(n10130), .CLK(n10825), 
        .Q(WX11177), .QN(n9273) );
  SDFFX1 DFF_1663_Q_reg ( .D(WX11178), .SI(WX11177), .SE(n10130), .CLK(n10825), 
        .Q(WX11179), .QN(n9271) );
  SDFFX1 DFF_1664_Q_reg ( .D(WX11180), .SI(WX11179), .SE(n10129), .CLK(n10826), 
        .Q(WX11181), .QN(n9541) );
  SDFFX1 DFF_1665_Q_reg ( .D(WX11182), .SI(WX11181), .SE(n10129), .CLK(n10826), 
        .Q(WX11183), .QN(n9542) );
  SDFFX1 DFF_1666_Q_reg ( .D(WX11184), .SI(WX11183), .SE(n10128), .CLK(n10826), 
        .Q(WX11185), .QN(n9543) );
  SDFFX1 DFF_1667_Q_reg ( .D(WX11186), .SI(WX11185), .SE(n10128), .CLK(n10826), 
        .Q(WX11187), .QN(n9544) );
  SDFFX1 DFF_1668_Q_reg ( .D(WX11188), .SI(WX11187), .SE(n10128), .CLK(n10826), 
        .Q(WX11189), .QN(n9545) );
  SDFFX1 DFF_1669_Q_reg ( .D(WX11190), .SI(WX11189), .SE(n10127), .CLK(n10827), 
        .Q(WX11191), .QN(n9546) );
  SDFFX1 DFF_1670_Q_reg ( .D(WX11192), .SI(WX11191), .SE(n10127), .CLK(n10827), 
        .Q(WX11193), .QN(n9547) );
  SDFFX1 DFF_1671_Q_reg ( .D(WX11194), .SI(WX11193), .SE(n10127), .CLK(n10827), 
        .Q(WX11195), .QN(n9548) );
  SDFFX1 DFF_1672_Q_reg ( .D(WX11196), .SI(WX11195), .SE(n10127), .CLK(n10827), 
        .Q(WX11197), .QN(n9549) );
  SDFFX1 DFF_1673_Q_reg ( .D(WX11198), .SI(WX11197), .SE(n10126), .CLK(n10827), 
        .Q(WX11199), .QN(n9550) );
  SDFFX1 DFF_1674_Q_reg ( .D(WX11200), .SI(WX11199), .SE(n10126), .CLK(n10827), 
        .Q(WX11201), .QN(n9551) );
  SDFFX1 DFF_1675_Q_reg ( .D(WX11202), .SI(WX11201), .SE(n10126), .CLK(n10827), 
        .Q(WX11203), .QN(n9552) );
  SDFFX1 DFF_1676_Q_reg ( .D(WX11204), .SI(WX11203), .SE(n10126), .CLK(n10827), 
        .Q(test_so97), .QN(n9913) );
  SDFFX1 DFF_1677_Q_reg ( .D(WX11206), .SI(test_si98), .SE(n10140), .CLK(
        n10820), .Q(WX11207), .QN(n9553) );
  SDFFX1 DFF_1678_Q_reg ( .D(WX11208), .SI(WX11207), .SE(n10140), .CLK(n10820), 
        .Q(WX11209), .QN(n9554) );
  SDFFX1 DFF_1679_Q_reg ( .D(WX11210), .SI(WX11209), .SE(n10139), .CLK(n10820), 
        .Q(WX11211), .QN(n9512) );
  SDFFX1 DFF_1680_Q_reg ( .D(WX11212), .SI(WX11211), .SE(n10138), .CLK(n10820), 
        .Q(WX11213), .QN(n9555) );
  SDFFX1 DFF_1681_Q_reg ( .D(WX11214), .SI(WX11213), .SE(n10138), .CLK(n10821), 
        .Q(WX11215), .QN(n9556) );
  SDFFX1 DFF_1682_Q_reg ( .D(WX11216), .SI(WX11215), .SE(n10137), .CLK(n10821), 
        .Q(WX11217), .QN(n9557) );
  SDFFX1 DFF_1683_Q_reg ( .D(WX11218), .SI(WX11217), .SE(n10136), .CLK(n10822), 
        .Q(WX11219), .QN(n9558) );
  SDFFX1 DFF_1684_Q_reg ( .D(WX11220), .SI(WX11219), .SE(n10136), .CLK(n10822), 
        .Q(WX11221), .QN(n9513) );
  SDFFX1 DFF_1685_Q_reg ( .D(WX11222), .SI(WX11221), .SE(n10135), .CLK(n10822), 
        .Q(WX11223), .QN(n9559) );
  SDFFX1 DFF_1686_Q_reg ( .D(WX11224), .SI(WX11223), .SE(n10135), .CLK(n10822), 
        .Q(WX11225), .QN(n9560) );
  SDFFX1 DFF_1687_Q_reg ( .D(WX11226), .SI(WX11225), .SE(n10134), .CLK(n10823), 
        .Q(WX11227), .QN(n9561) );
  SDFFX1 DFF_1688_Q_reg ( .D(WX11228), .SI(WX11227), .SE(n10134), .CLK(n10823), 
        .Q(WX11229), .QN(n9562) );
  SDFFX1 DFF_1689_Q_reg ( .D(WX11230), .SI(WX11229), .SE(n10133), .CLK(n10823), 
        .Q(WX11231), .QN(n9563) );
  SDFFX1 DFF_1690_Q_reg ( .D(WX11232), .SI(WX11231), .SE(n10133), .CLK(n10824), 
        .Q(WX11233), .QN(n9564) );
  SDFFX1 DFF_1691_Q_reg ( .D(WX11234), .SI(WX11233), .SE(n10132), .CLK(n10824), 
        .Q(WX11235), .QN(n9514) );
  SDFFX1 DFF_1692_Q_reg ( .D(WX11236), .SI(WX11235), .SE(n10132), .CLK(n10824), 
        .Q(WX11237), .QN(n9565) );
  SDFFX1 DFF_1693_Q_reg ( .D(WX11238), .SI(WX11237), .SE(n10131), .CLK(n10825), 
        .Q(test_so98), .QN(n9906) );
  SDFFX1 DFF_1694_Q_reg ( .D(WX11240), .SI(test_si99), .SE(n10130), .CLK(
        n10825), .Q(WX11241), .QN(n9566) );
  SDFFX1 DFF_1695_Q_reg ( .D(WX11242), .SI(WX11241), .SE(n10130), .CLK(n10825), 
        .Q(WX11243), .QN(n9533) );
  SDFFX1 DFF_1696_Q_reg ( .D(WX11608), .SI(WX11243), .SE(n10124), .CLK(n10828), 
        .Q(CRC_OUT_1_0), .QN(DFF_1696_n1) );
  SDFFX1 DFF_1697_Q_reg ( .D(WX11610), .SI(CRC_OUT_1_0), .SE(n10124), .CLK(
        n10828), .Q(CRC_OUT_1_1), .QN(DFF_1697_n1) );
  SDFFX1 DFF_1698_Q_reg ( .D(WX11612), .SI(CRC_OUT_1_1), .SE(n10124), .CLK(
        n10828), .Q(CRC_OUT_1_2), .QN(DFF_1698_n1) );
  SDFFX1 DFF_1699_Q_reg ( .D(WX11614), .SI(CRC_OUT_1_2), .SE(n10124), .CLK(
        n10828), .Q(CRC_OUT_1_3), .QN(DFF_1699_n1) );
  SDFFX1 DFF_1700_Q_reg ( .D(WX11616), .SI(CRC_OUT_1_3), .SE(n10124), .CLK(
        n10828), .Q(CRC_OUT_1_4), .QN(DFF_1700_n1) );
  SDFFX1 DFF_1701_Q_reg ( .D(WX11618), .SI(CRC_OUT_1_4), .SE(n10124), .CLK(
        n10828), .Q(CRC_OUT_1_5), .QN(DFF_1701_n1) );
  SDFFX1 DFF_1702_Q_reg ( .D(WX11620), .SI(CRC_OUT_1_5), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_6), .QN(DFF_1702_n1) );
  SDFFX1 DFF_1703_Q_reg ( .D(WX11622), .SI(CRC_OUT_1_6), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_7), .QN(DFF_1703_n1) );
  SDFFX1 DFF_1704_Q_reg ( .D(WX11624), .SI(CRC_OUT_1_7), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_8), .QN(DFF_1704_n1) );
  SDFFX1 DFF_1705_Q_reg ( .D(WX11626), .SI(CRC_OUT_1_8), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_9), .QN(DFF_1705_n1) );
  SDFFX1 DFF_1706_Q_reg ( .D(WX11628), .SI(CRC_OUT_1_9), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_10), .QN(DFF_1706_n1) );
  SDFFX1 DFF_1707_Q_reg ( .D(WX11630), .SI(CRC_OUT_1_10), .SE(n10123), .CLK(
        n10829), .Q(CRC_OUT_1_11), .QN(DFF_1707_n1) );
  SDFFX1 DFF_1708_Q_reg ( .D(WX11632), .SI(CRC_OUT_1_11), .SE(n10122), .CLK(
        n10829), .Q(CRC_OUT_1_12), .QN(DFF_1708_n1) );
  SDFFX1 DFF_1709_Q_reg ( .D(WX11634), .SI(CRC_OUT_1_12), .SE(n10122), .CLK(
        n10829), .Q(CRC_OUT_1_13), .QN(DFF_1709_n1) );
  SDFFX1 DFF_1710_Q_reg ( .D(WX11636), .SI(CRC_OUT_1_13), .SE(n10122), .CLK(
        n10829), .Q(test_so99), .QN(n9950) );
  SDFFX1 DFF_1711_Q_reg ( .D(WX11638), .SI(test_si100), .SE(n10122), .CLK(
        n10829), .Q(CRC_OUT_1_15), .QN(DFF_1711_n1) );
  SDFFX1 DFF_1712_Q_reg ( .D(WX11640), .SI(CRC_OUT_1_15), .SE(n10122), .CLK(
        n10829), .Q(CRC_OUT_1_16), .QN(DFF_1712_n1) );
  SDFFX1 DFF_1713_Q_reg ( .D(WX11642), .SI(CRC_OUT_1_16), .SE(n10122), .CLK(
        n10829), .Q(CRC_OUT_1_17), .QN(DFF_1713_n1) );
  SDFFX1 DFF_1714_Q_reg ( .D(WX11644), .SI(CRC_OUT_1_17), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_18), .QN(DFF_1714_n1) );
  SDFFX1 DFF_1715_Q_reg ( .D(WX11646), .SI(CRC_OUT_1_18), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_19), .QN(DFF_1715_n1) );
  SDFFX1 DFF_1716_Q_reg ( .D(WX11648), .SI(CRC_OUT_1_19), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_20), .QN(DFF_1716_n1) );
  SDFFX1 DFF_1717_Q_reg ( .D(WX11650), .SI(CRC_OUT_1_20), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_21), .QN(DFF_1717_n1) );
  SDFFX1 DFF_1718_Q_reg ( .D(WX11652), .SI(CRC_OUT_1_21), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_22), .QN(DFF_1718_n1) );
  SDFFX1 DFF_1719_Q_reg ( .D(WX11654), .SI(CRC_OUT_1_22), .SE(n10121), .CLK(
        n10830), .Q(CRC_OUT_1_23), .QN(DFF_1719_n1) );
  SDFFX1 DFF_1720_Q_reg ( .D(WX11656), .SI(CRC_OUT_1_23), .SE(n10126), .CLK(
        n10827), .Q(CRC_OUT_1_24), .QN(DFF_1720_n1) );
  SDFFX1 DFF_1721_Q_reg ( .D(WX11658), .SI(CRC_OUT_1_24), .SE(n10126), .CLK(
        n10827), .Q(CRC_OUT_1_25), .QN(DFF_1721_n1) );
  SDFFX1 DFF_1722_Q_reg ( .D(WX11660), .SI(CRC_OUT_1_25), .SE(n10125), .CLK(
        n10828), .Q(CRC_OUT_1_26), .QN(DFF_1722_n1) );
  SDFFX1 DFF_1723_Q_reg ( .D(WX11662), .SI(CRC_OUT_1_26), .SE(n10125), .CLK(
        n10828), .Q(CRC_OUT_1_27), .QN(DFF_1723_n1) );
  SDFFX1 DFF_1724_Q_reg ( .D(WX11664), .SI(CRC_OUT_1_27), .SE(n10125), .CLK(
        n10828), .Q(CRC_OUT_1_28), .QN(DFF_1724_n1) );
  SDFFX1 DFF_1725_Q_reg ( .D(WX11666), .SI(CRC_OUT_1_28), .SE(n10125), .CLK(
        n10828), .Q(CRC_OUT_1_29), .QN(DFF_1725_n1) );
  SDFFX1 DFF_1726_Q_reg ( .D(WX11668), .SI(CRC_OUT_1_29), .SE(n10125), .CLK(
        n10828), .Q(CRC_OUT_1_30), .QN(DFF_1726_n1) );
  SDFFX1 DFF_1727_Q_reg ( .D(WX11670), .SI(CRC_OUT_1_30), .SE(n10125), .CLK(
        n10828), .Q(test_so100), .QN(n9884) );
  AND2X1 Trojan1 ( .IN1(WX742), .IN2(WX7249), .Q(Tj_OUT1) );
  AND2X1 Trojan2 ( .IN1(WX5922), .IN2(WX5960), .Q(Tj_OUT2) );
  AND2X1 Trojan3 ( .IN1(WX4697), .IN2(WX9032), .Q(Tj_OUT3) );
  AND2X1 Trojan4 ( .IN1(n1483), .IN2(n1947), .Q(Tj_OUT4) );
  NOR4X0 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .QN(Tj_OUT1234) );
  AND2X1 Trojan5 ( .IN1(WX3340), .IN2(WX6476), .Q(Tj_OUT5) );
  AND2X1 Trojan6 ( .IN1(WX9819), .IN2(n268), .Q(Tj_OUT6) );
  AND2X1 Trojan7 ( .IN1(n1000), .IN2(WX3458), .Q(Tj_OUT7) );
  AND2X1 Trojan8 ( .IN1(WX9060), .IN2(WX7749), .Q(Tj_OUT8) );
  NOR4X0 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .QN(Tj_OUT5678) );
  INVX0 TrojanINV_test_se ( .INP(n10370), .ZN(test_se_NOT) );
  AND3X1 Trojan_Trigger ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .IN3(test_se_NOT), .Q(Tj_Trigger) );
  DFFX2 TrojanScanEnable ( .D(1'b1), .CLK(Tj_Trigger), .Q(Trojan_SE) );
  MUX21X1 Trojan_Payload1 ( .IN1(n10370), .IN2(1'b1), .S(Trojan_SE), .Q(
        test_se_Trojan) );
  MUX21X1 Trojan_Payload2 ( .IN1(WX11155), .IN2(WX3442), .S(Trojan_SE), .Q(
        WX11155_Tj_Payload) );
  INVX2 U9790 ( .INP(TM0), .ZN(n2182) );
  NBUFFX2 U9791 ( .INP(n10053), .Z(n10027) );
  NBUFFX2 U9792 ( .INP(n10053), .Z(n10028) );
  NBUFFX2 U9793 ( .INP(n10051), .Z(n10036) );
  NBUFFX2 U9794 ( .INP(n10051), .Z(n10038) );
  NBUFFX2 U9795 ( .INP(n10050), .Z(n10039) );
  NBUFFX2 U9796 ( .INP(n10050), .Z(n10040) );
  NBUFFX2 U9797 ( .INP(n10050), .Z(n10041) );
  NBUFFX2 U9798 ( .INP(n10050), .Z(n10042) );
  NBUFFX2 U9799 ( .INP(n10050), .Z(n10043) );
  NBUFFX2 U9800 ( .INP(n10049), .Z(n10047) );
  NBUFFX2 U9801 ( .INP(n10052), .Z(n10029) );
  NBUFFX2 U9802 ( .INP(n10052), .Z(n10030) );
  NBUFFX2 U9803 ( .INP(n10052), .Z(n10031) );
  NBUFFX2 U9804 ( .INP(n10051), .Z(n10037) );
  NBUFFX2 U9805 ( .INP(n10052), .Z(n10032) );
  NBUFFX2 U9806 ( .INP(n10052), .Z(n10033) );
  NBUFFX2 U9807 ( .INP(n10051), .Z(n10034) );
  NBUFFX2 U9808 ( .INP(n10051), .Z(n10035) );
  NBUFFX2 U9809 ( .INP(n10049), .Z(n10044) );
  NBUFFX2 U9810 ( .INP(n10049), .Z(n10045) );
  NBUFFX2 U9811 ( .INP(n10049), .Z(n10046) );
  NBUFFX2 U9812 ( .INP(n10053), .Z(n10026) );
  NBUFFX2 U9813 ( .INP(n10877), .Z(n10708) );
  NBUFFX2 U9814 ( .INP(n10877), .Z(n10706) );
  NBUFFX2 U9815 ( .INP(n10877), .Z(n10707) );
  NBUFFX2 U9816 ( .INP(n10877), .Z(n10705) );
  NBUFFX2 U9817 ( .INP(n10852), .Z(n10829) );
  NBUFFX2 U9818 ( .INP(n10853), .Z(n10828) );
  NBUFFX2 U9819 ( .INP(n10853), .Z(n10827) );
  NBUFFX2 U9820 ( .INP(n10853), .Z(n10826) );
  NBUFFX2 U9821 ( .INP(n10853), .Z(n10825) );
  NBUFFX2 U9822 ( .INP(n10853), .Z(n10824) );
  NBUFFX2 U9823 ( .INP(n10854), .Z(n10823) );
  NBUFFX2 U9824 ( .INP(n10854), .Z(n10822) );
  NBUFFX2 U9825 ( .INP(n10854), .Z(n10821) );
  NBUFFX2 U9826 ( .INP(n10854), .Z(n10820) );
  NBUFFX2 U9827 ( .INP(n10854), .Z(n10819) );
  NBUFFX2 U9828 ( .INP(n10855), .Z(n10818) );
  NBUFFX2 U9829 ( .INP(n10855), .Z(n10815) );
  NBUFFX2 U9830 ( .INP(n10855), .Z(n10816) );
  NBUFFX2 U9831 ( .INP(n10855), .Z(n10817) );
  NBUFFX2 U9832 ( .INP(n10855), .Z(n10814) );
  NBUFFX2 U9833 ( .INP(n10852), .Z(n10831) );
  NBUFFX2 U9834 ( .INP(n10852), .Z(n10830) );
  NBUFFX2 U9835 ( .INP(n10856), .Z(n10813) );
  NBUFFX2 U9836 ( .INP(n10856), .Z(n10812) );
  NBUFFX2 U9837 ( .INP(n10856), .Z(n10811) );
  NBUFFX2 U9838 ( .INP(n10856), .Z(n10810) );
  NBUFFX2 U9839 ( .INP(n10856), .Z(n10809) );
  NBUFFX2 U9840 ( .INP(n10857), .Z(n10808) );
  NBUFFX2 U9841 ( .INP(n10857), .Z(n10807) );
  NBUFFX2 U9842 ( .INP(n10857), .Z(n10806) );
  NBUFFX2 U9843 ( .INP(n10857), .Z(n10805) );
  NBUFFX2 U9844 ( .INP(n10857), .Z(n10804) );
  NBUFFX2 U9845 ( .INP(n10858), .Z(n10801) );
  NBUFFX2 U9846 ( .INP(n10858), .Z(n10802) );
  NBUFFX2 U9847 ( .INP(n10858), .Z(n10803) );
  NBUFFX2 U9848 ( .INP(n10852), .Z(n10833) );
  NBUFFX2 U9849 ( .INP(n10852), .Z(n10832) );
  NBUFFX2 U9850 ( .INP(n10858), .Z(n10800) );
  NBUFFX2 U9851 ( .INP(n10858), .Z(n10799) );
  NBUFFX2 U9852 ( .INP(n10859), .Z(n10798) );
  NBUFFX2 U9853 ( .INP(n10859), .Z(n10797) );
  NBUFFX2 U9854 ( .INP(n10859), .Z(n10796) );
  NBUFFX2 U9855 ( .INP(n10859), .Z(n10795) );
  NBUFFX2 U9856 ( .INP(n10859), .Z(n10794) );
  NBUFFX2 U9857 ( .INP(n10860), .Z(n10793) );
  NBUFFX2 U9858 ( .INP(n10860), .Z(n10792) );
  NBUFFX2 U9859 ( .INP(n10860), .Z(n10791) );
  NBUFFX2 U9860 ( .INP(n10860), .Z(n10790) );
  NBUFFX2 U9861 ( .INP(n10851), .Z(n10834) );
  NBUFFX2 U9862 ( .INP(n10861), .Z(n10788) );
  NBUFFX2 U9863 ( .INP(n10860), .Z(n10789) );
  NBUFFX2 U9864 ( .INP(n10861), .Z(n10787) );
  NBUFFX2 U9865 ( .INP(n10851), .Z(n10836) );
  NBUFFX2 U9866 ( .INP(n10851), .Z(n10835) );
  NBUFFX2 U9867 ( .INP(n10861), .Z(n10786) );
  NBUFFX2 U9868 ( .INP(n10861), .Z(n10785) );
  NBUFFX2 U9869 ( .INP(n10861), .Z(n10784) );
  NBUFFX2 U9870 ( .INP(n10862), .Z(n10783) );
  NBUFFX2 U9871 ( .INP(n10862), .Z(n10782) );
  NBUFFX2 U9872 ( .INP(n10862), .Z(n10781) );
  NBUFFX2 U9873 ( .INP(n10862), .Z(n10780) );
  NBUFFX2 U9874 ( .INP(n10862), .Z(n10779) );
  NBUFFX2 U9875 ( .INP(n10863), .Z(n10778) );
  NBUFFX2 U9876 ( .INP(n10863), .Z(n10777) );
  NBUFFX2 U9877 ( .INP(n10863), .Z(n10774) );
  NBUFFX2 U9878 ( .INP(n10863), .Z(n10775) );
  NBUFFX2 U9879 ( .INP(n10863), .Z(n10776) );
  NBUFFX2 U9880 ( .INP(n10864), .Z(n10773) );
  NBUFFX2 U9881 ( .INP(n10851), .Z(n10838) );
  NBUFFX2 U9882 ( .INP(n10851), .Z(n10837) );
  NBUFFX2 U9883 ( .INP(n10864), .Z(n10772) );
  NBUFFX2 U9884 ( .INP(n10864), .Z(n10771) );
  NBUFFX2 U9885 ( .INP(n10864), .Z(n10770) );
  NBUFFX2 U9886 ( .INP(n10864), .Z(n10769) );
  NBUFFX2 U9887 ( .INP(n10865), .Z(n10768) );
  NBUFFX2 U9888 ( .INP(n10865), .Z(n10767) );
  NBUFFX2 U9889 ( .INP(n10865), .Z(n10766) );
  NBUFFX2 U9890 ( .INP(n10865), .Z(n10765) );
  NBUFFX2 U9891 ( .INP(n10865), .Z(n10764) );
  NBUFFX2 U9892 ( .INP(n10866), .Z(n10763) );
  NBUFFX2 U9893 ( .INP(n10866), .Z(n10760) );
  NBUFFX2 U9894 ( .INP(n10866), .Z(n10761) );
  NBUFFX2 U9895 ( .INP(n10866), .Z(n10762) );
  NBUFFX2 U9896 ( .INP(n10850), .Z(n10840) );
  NBUFFX2 U9897 ( .INP(n10850), .Z(n10839) );
  NBUFFX2 U9898 ( .INP(n10866), .Z(n10759) );
  NBUFFX2 U9899 ( .INP(n10867), .Z(n10758) );
  NBUFFX2 U9900 ( .INP(n10867), .Z(n10757) );
  NBUFFX2 U9901 ( .INP(n10867), .Z(n10756) );
  NBUFFX2 U9902 ( .INP(n10867), .Z(n10755) );
  NBUFFX2 U9903 ( .INP(n10867), .Z(n10754) );
  NBUFFX2 U9904 ( .INP(n10868), .Z(n10753) );
  NBUFFX2 U9905 ( .INP(n10868), .Z(n10752) );
  NBUFFX2 U9906 ( .INP(n10868), .Z(n10751) );
  NBUFFX2 U9907 ( .INP(n10868), .Z(n10750) );
  NBUFFX2 U9908 ( .INP(n10850), .Z(n10841) );
  NBUFFX2 U9909 ( .INP(n10869), .Z(n10747) );
  NBUFFX2 U9910 ( .INP(n10869), .Z(n10748) );
  NBUFFX2 U9911 ( .INP(n10868), .Z(n10749) );
  NBUFFX2 U9912 ( .INP(n10850), .Z(n10843) );
  NBUFFX2 U9913 ( .INP(n10850), .Z(n10842) );
  NBUFFX2 U9914 ( .INP(n10869), .Z(n10746) );
  NBUFFX2 U9915 ( .INP(n10869), .Z(n10745) );
  NBUFFX2 U9916 ( .INP(n10869), .Z(n10744) );
  NBUFFX2 U9917 ( .INP(n10870), .Z(n10743) );
  NBUFFX2 U9918 ( .INP(n10870), .Z(n10742) );
  NBUFFX2 U9919 ( .INP(n10870), .Z(n10741) );
  NBUFFX2 U9920 ( .INP(n10870), .Z(n10740) );
  NBUFFX2 U9921 ( .INP(n10870), .Z(n10739) );
  NBUFFX2 U9922 ( .INP(n10871), .Z(n10738) );
  NBUFFX2 U9923 ( .INP(n10871), .Z(n10737) );
  NBUFFX2 U9924 ( .INP(n10871), .Z(n10734) );
  NBUFFX2 U9925 ( .INP(n10871), .Z(n10735) );
  NBUFFX2 U9926 ( .INP(n10871), .Z(n10736) );
  NBUFFX2 U9927 ( .INP(n10849), .Z(n10846) );
  NBUFFX2 U9928 ( .INP(n10849), .Z(n10845) );
  NBUFFX2 U9929 ( .INP(n10849), .Z(n10844) );
  NBUFFX2 U9930 ( .INP(n10872), .Z(n10733) );
  NBUFFX2 U9931 ( .INP(n10872), .Z(n10732) );
  NBUFFX2 U9932 ( .INP(n10872), .Z(n10731) );
  NBUFFX2 U9933 ( .INP(n10874), .Z(n10723) );
  NBUFFX2 U9934 ( .INP(n10874), .Z(n10722) );
  NBUFFX2 U9935 ( .INP(n10872), .Z(n10730) );
  NBUFFX2 U9936 ( .INP(n10872), .Z(n10729) );
  NBUFFX2 U9937 ( .INP(n10873), .Z(n10728) );
  NBUFFX2 U9938 ( .INP(n10873), .Z(n10727) );
  NBUFFX2 U9939 ( .INP(n10873), .Z(n10726) );
  NBUFFX2 U9940 ( .INP(n10873), .Z(n10725) );
  NBUFFX2 U9941 ( .INP(n10873), .Z(n10724) );
  NBUFFX2 U9942 ( .INP(n10874), .Z(n10720) );
  NBUFFX2 U9943 ( .INP(n10874), .Z(n10721) );
  NBUFFX2 U9944 ( .INP(n10874), .Z(n10719) );
  NBUFFX2 U9945 ( .INP(n10849), .Z(n10848) );
  NBUFFX2 U9946 ( .INP(n10849), .Z(n10847) );
  NBUFFX2 U9947 ( .INP(n10875), .Z(n10718) );
  NBUFFX2 U9948 ( .INP(n10875), .Z(n10717) );
  NBUFFX2 U9949 ( .INP(n10875), .Z(n10716) );
  NBUFFX2 U9950 ( .INP(n10875), .Z(n10715) );
  NBUFFX2 U9951 ( .INP(n10875), .Z(n10714) );
  NBUFFX2 U9952 ( .INP(n10876), .Z(n10713) );
  NBUFFX2 U9953 ( .INP(n10876), .Z(n10712) );
  NBUFFX2 U9954 ( .INP(n10876), .Z(n10711) );
  NBUFFX2 U9955 ( .INP(n10876), .Z(n10710) );
  NBUFFX2 U9956 ( .INP(n10876), .Z(n10709) );
  NBUFFX2 U9957 ( .INP(n10049), .Z(n10048) );
  NBUFFX2 U9958 ( .INP(n10082), .Z(n10063) );
  NBUFFX2 U9959 ( .INP(n9968), .Z(n9977) );
  NBUFFX2 U9960 ( .INP(n9971), .Z(n9993) );
  NBUFFX2 U9961 ( .INP(n9971), .Z(n9992) );
  NBUFFX2 U9962 ( .INP(n10080), .Z(n10070) );
  NBUFFX2 U9963 ( .INP(n10080), .Z(n10071) );
  NBUFFX2 U9964 ( .INP(n10080), .Z(n10072) );
  NBUFFX2 U9965 ( .INP(n10080), .Z(n10073) );
  NBUFFX2 U9966 ( .INP(n10079), .Z(n10077) );
  NBUFFX2 U9967 ( .INP(n10081), .Z(n10065) );
  NBUFFX2 U9968 ( .INP(n10081), .Z(n10066) );
  NBUFFX2 U9969 ( .INP(n10081), .Z(n10067) );
  NBUFFX2 U9970 ( .INP(n10081), .Z(n10064) );
  NBUFFX2 U9971 ( .INP(n10080), .Z(n10069) );
  NBUFFX2 U9972 ( .INP(n10081), .Z(n10068) );
  NBUFFX2 U9973 ( .INP(n10079), .Z(n10074) );
  NBUFFX2 U9974 ( .INP(n10079), .Z(n10075) );
  NBUFFX2 U9975 ( .INP(n10079), .Z(n10076) );
  NBUFFX2 U9976 ( .INP(n9969), .Z(n9985) );
  NBUFFX2 U9977 ( .INP(n9969), .Z(n9984) );
  NBUFFX2 U9978 ( .INP(n9969), .Z(n9983) );
  NBUFFX2 U9979 ( .INP(n9969), .Z(n9982) );
  NBUFFX2 U9980 ( .INP(n9968), .Z(n9981) );
  NBUFFX2 U9981 ( .INP(n9970), .Z(n9991) );
  NBUFFX2 U9982 ( .INP(n9970), .Z(n9990) );
  NBUFFX2 U9983 ( .INP(n9970), .Z(n9989) );
  NBUFFX2 U9984 ( .INP(n9970), .Z(n9988) );
  NBUFFX2 U9985 ( .INP(n9970), .Z(n9987) );
  NBUFFX2 U9986 ( .INP(n9969), .Z(n9986) );
  NBUFFX2 U9987 ( .INP(n9968), .Z(n9978) );
  NBUFFX2 U9988 ( .INP(n9968), .Z(n9979) );
  NBUFFX2 U9989 ( .INP(n9968), .Z(n9980) );
  NBUFFX2 U9990 ( .INP(n10083), .Z(n10056) );
  NBUFFX2 U9991 ( .INP(n10083), .Z(n10058) );
  NBUFFX2 U9992 ( .INP(n10083), .Z(n10057) );
  NBUFFX2 U9993 ( .INP(n10082), .Z(n10062) );
  NBUFFX2 U9994 ( .INP(n10082), .Z(n10061) );
  NBUFFX2 U9995 ( .INP(n10082), .Z(n10059) );
  NBUFFX2 U9996 ( .INP(n10082), .Z(n10060) );
  NBUFFX2 U9997 ( .INP(n9967), .Z(n9976) );
  NBUFFX2 U9998 ( .INP(n9967), .Z(n9975) );
  NBUFFX2 U9999 ( .INP(n9967), .Z(n9974) );
  NBUFFX2 U10000 ( .INP(n9967), .Z(n9973) );
  NBUFFX2 U10001 ( .INP(n9967), .Z(n9972) );
  NBUFFX2 U10002 ( .INP(n10079), .Z(n10078) );
  NBUFFX2 U10003 ( .INP(n9971), .Z(n9994) );
  NBUFFX2 U10004 ( .INP(n9999), .Z(n10022) );
  NBUFFX2 U10005 ( .INP(n9999), .Z(n10020) );
  NBUFFX2 U10006 ( .INP(n9999), .Z(n10021) );
  NBUFFX2 U10007 ( .INP(n9997), .Z(n10010) );
  NBUFFX2 U10008 ( .INP(n9997), .Z(n10011) );
  NBUFFX2 U10009 ( .INP(n9997), .Z(n10012) );
  NBUFFX2 U10010 ( .INP(n9997), .Z(n10013) );
  NBUFFX2 U10011 ( .INP(n9997), .Z(n10014) );
  NBUFFX2 U10012 ( .INP(n9998), .Z(n10015) );
  NBUFFX2 U10013 ( .INP(n9998), .Z(n10016) );
  NBUFFX2 U10014 ( .INP(n9998), .Z(n10017) );
  NBUFFX2 U10015 ( .INP(n9998), .Z(n10018) );
  NBUFFX2 U10016 ( .INP(n9995), .Z(n10000) );
  NBUFFX2 U10017 ( .INP(n9995), .Z(n10001) );
  NBUFFX2 U10018 ( .INP(n9995), .Z(n10002) );
  NBUFFX2 U10019 ( .INP(n9995), .Z(n10003) );
  NBUFFX2 U10020 ( .INP(n9995), .Z(n10004) );
  NBUFFX2 U10021 ( .INP(n9996), .Z(n10005) );
  NBUFFX2 U10022 ( .INP(n9996), .Z(n10006) );
  NBUFFX2 U10023 ( .INP(n9996), .Z(n10007) );
  NBUFFX2 U10024 ( .INP(n9996), .Z(n10008) );
  NBUFFX2 U10025 ( .INP(n9996), .Z(n10009) );
  NBUFFX2 U10026 ( .INP(n9998), .Z(n10019) );
  NBUFFX2 U10027 ( .INP(n9999), .Z(n10023) );
  NBUFFX2 U10028 ( .INP(n10896), .Z(n9967) );
  NBUFFX2 U10029 ( .INP(n10896), .Z(n9968) );
  NBUFFX2 U10030 ( .INP(n10896), .Z(n9969) );
  NBUFFX2 U10031 ( .INP(n10896), .Z(n9970) );
  NBUFFX2 U10032 ( .INP(n10896), .Z(n9971) );
  NBUFFX2 U10033 ( .INP(n2148), .Z(n9995) );
  NBUFFX2 U10034 ( .INP(n2148), .Z(n9996) );
  NBUFFX2 U10035 ( .INP(n2148), .Z(n9997) );
  NBUFFX2 U10036 ( .INP(n2148), .Z(n9998) );
  NBUFFX2 U10037 ( .INP(n2148), .Z(n9999) );
  NBUFFX2 U10038 ( .INP(n2152), .Z(n10024) );
  NBUFFX2 U10039 ( .INP(n2152), .Z(n10025) );
  NBUFFX2 U10040 ( .INP(n10024), .Z(n10049) );
  NBUFFX2 U10041 ( .INP(n10024), .Z(n10050) );
  NBUFFX2 U10042 ( .INP(n10024), .Z(n10051) );
  NBUFFX2 U10043 ( .INP(n10025), .Z(n10052) );
  NBUFFX2 U10044 ( .INP(n10025), .Z(n10053) );
  NBUFFX2 U10045 ( .INP(n2153), .Z(n10054) );
  NBUFFX2 U10046 ( .INP(n2153), .Z(n10055) );
  NBUFFX2 U10047 ( .INP(n10054), .Z(n10079) );
  NBUFFX2 U10048 ( .INP(n10054), .Z(n10080) );
  NBUFFX2 U10049 ( .INP(n10054), .Z(n10081) );
  NBUFFX2 U10050 ( .INP(n10055), .Z(n10082) );
  NBUFFX2 U10051 ( .INP(n10055), .Z(n10083) );
  NBUFFX2 U10052 ( .INP(n10466), .Z(n10084) );
  NBUFFX2 U10053 ( .INP(n10466), .Z(n10085) );
  NBUFFX2 U10054 ( .INP(n10465), .Z(n10086) );
  NBUFFX2 U10055 ( .INP(n10465), .Z(n10087) );
  NBUFFX2 U10056 ( .INP(n10465), .Z(n10088) );
  NBUFFX2 U10057 ( .INP(n10464), .Z(n10089) );
  NBUFFX2 U10058 ( .INP(n10464), .Z(n10090) );
  NBUFFX2 U10059 ( .INP(n10464), .Z(n10091) );
  NBUFFX2 U10060 ( .INP(n10463), .Z(n10092) );
  NBUFFX2 U10061 ( .INP(n10463), .Z(n10093) );
  NBUFFX2 U10062 ( .INP(n10463), .Z(n10094) );
  NBUFFX2 U10063 ( .INP(n10462), .Z(n10095) );
  NBUFFX2 U10064 ( .INP(n10462), .Z(n10096) );
  NBUFFX2 U10065 ( .INP(n10462), .Z(n10097) );
  NBUFFX2 U10066 ( .INP(n10461), .Z(n10098) );
  NBUFFX2 U10067 ( .INP(n10461), .Z(n10099) );
  NBUFFX2 U10068 ( .INP(n10461), .Z(n10100) );
  NBUFFX2 U10069 ( .INP(n10460), .Z(n10101) );
  NBUFFX2 U10070 ( .INP(n10460), .Z(n10102) );
  NBUFFX2 U10071 ( .INP(n10460), .Z(n10103) );
  NBUFFX2 U10072 ( .INP(n10459), .Z(n10104) );
  NBUFFX2 U10073 ( .INP(n10459), .Z(n10105) );
  NBUFFX2 U10074 ( .INP(n10459), .Z(n10106) );
  NBUFFX2 U10075 ( .INP(n10458), .Z(n10107) );
  NBUFFX2 U10076 ( .INP(n10458), .Z(n10108) );
  NBUFFX2 U10077 ( .INP(n10458), .Z(n10109) );
  NBUFFX2 U10078 ( .INP(n10457), .Z(n10110) );
  NBUFFX2 U10079 ( .INP(n10457), .Z(n10111) );
  NBUFFX2 U10080 ( .INP(n10457), .Z(n10112) );
  NBUFFX2 U10081 ( .INP(n10456), .Z(n10113) );
  NBUFFX2 U10082 ( .INP(n10456), .Z(n10114) );
  NBUFFX2 U10083 ( .INP(n10456), .Z(n10115) );
  NBUFFX2 U10084 ( .INP(n10455), .Z(n10116) );
  NBUFFX2 U10085 ( .INP(n10455), .Z(n10117) );
  NBUFFX2 U10086 ( .INP(n10455), .Z(n10118) );
  NBUFFX2 U10087 ( .INP(n10454), .Z(n10119) );
  NBUFFX2 U10088 ( .INP(n10454), .Z(n10120) );
  NBUFFX2 U10089 ( .INP(n10454), .Z(n10121) );
  NBUFFX2 U10090 ( .INP(n10453), .Z(n10122) );
  NBUFFX2 U10091 ( .INP(n10453), .Z(n10123) );
  NBUFFX2 U10092 ( .INP(n10453), .Z(n10124) );
  NBUFFX2 U10093 ( .INP(n10452), .Z(n10125) );
  NBUFFX2 U10094 ( .INP(n10452), .Z(n10126) );
  NBUFFX2 U10095 ( .INP(n10452), .Z(n10127) );
  NBUFFX2 U10096 ( .INP(n10451), .Z(n10128) );
  NBUFFX2 U10097 ( .INP(n10451), .Z(n10129) );
  NBUFFX2 U10098 ( .INP(n10451), .Z(n10130) );
  NBUFFX2 U10099 ( .INP(n10450), .Z(n10131) );
  NBUFFX2 U10100 ( .INP(n10450), .Z(n10132) );
  NBUFFX2 U10101 ( .INP(n10450), .Z(n10133) );
  NBUFFX2 U10102 ( .INP(n10449), .Z(n10134) );
  NBUFFX2 U10103 ( .INP(n10449), .Z(n10135) );
  NBUFFX2 U10104 ( .INP(n10449), .Z(n10136) );
  NBUFFX2 U10105 ( .INP(n10448), .Z(n10137) );
  NBUFFX2 U10106 ( .INP(n10448), .Z(n10138) );
  NBUFFX2 U10107 ( .INP(n10448), .Z(n10139) );
  NBUFFX2 U10108 ( .INP(n10447), .Z(n10140) );
  NBUFFX2 U10109 ( .INP(n10447), .Z(n10141) );
  NBUFFX2 U10110 ( .INP(n10447), .Z(n10142) );
  NBUFFX2 U10111 ( .INP(n10446), .Z(n10143) );
  NBUFFX2 U10112 ( .INP(n10446), .Z(n10144) );
  NBUFFX2 U10113 ( .INP(n10446), .Z(n10145) );
  NBUFFX2 U10114 ( .INP(n10445), .Z(n10146) );
  NBUFFX2 U10115 ( .INP(n10445), .Z(n10147) );
  NBUFFX2 U10116 ( .INP(n10445), .Z(n10148) );
  NBUFFX2 U10117 ( .INP(n10444), .Z(n10149) );
  NBUFFX2 U10118 ( .INP(n10444), .Z(n10150) );
  NBUFFX2 U10119 ( .INP(n10444), .Z(n10151) );
  NBUFFX2 U10120 ( .INP(n10443), .Z(n10152) );
  NBUFFX2 U10121 ( .INP(n10443), .Z(n10153) );
  NBUFFX2 U10122 ( .INP(n10443), .Z(n10154) );
  NBUFFX2 U10123 ( .INP(n10442), .Z(n10155) );
  NBUFFX2 U10124 ( .INP(n10442), .Z(n10156) );
  NBUFFX2 U10125 ( .INP(n10442), .Z(n10157) );
  NBUFFX2 U10126 ( .INP(n10441), .Z(n10158) );
  NBUFFX2 U10127 ( .INP(n10441), .Z(n10159) );
  NBUFFX2 U10128 ( .INP(n10441), .Z(n10160) );
  NBUFFX2 U10129 ( .INP(n10440), .Z(n10161) );
  NBUFFX2 U10130 ( .INP(n10440), .Z(n10162) );
  NBUFFX2 U10131 ( .INP(n10440), .Z(n10163) );
  NBUFFX2 U10132 ( .INP(n10439), .Z(n10164) );
  NBUFFX2 U10133 ( .INP(n10439), .Z(n10165) );
  NBUFFX2 U10134 ( .INP(n10439), .Z(n10166) );
  NBUFFX2 U10135 ( .INP(n10438), .Z(n10167) );
  NBUFFX2 U10136 ( .INP(n10438), .Z(n10168) );
  NBUFFX2 U10137 ( .INP(n10438), .Z(n10169) );
  NBUFFX2 U10138 ( .INP(n10437), .Z(n10170) );
  NBUFFX2 U10139 ( .INP(n10437), .Z(n10171) );
  NBUFFX2 U10140 ( .INP(n10437), .Z(n10172) );
  NBUFFX2 U10141 ( .INP(n10436), .Z(n10173) );
  NBUFFX2 U10142 ( .INP(n10436), .Z(n10174) );
  NBUFFX2 U10143 ( .INP(n10436), .Z(n10175) );
  NBUFFX2 U10144 ( .INP(n10435), .Z(n10176) );
  NBUFFX2 U10145 ( .INP(n10435), .Z(n10177) );
  NBUFFX2 U10146 ( .INP(n10435), .Z(n10178) );
  NBUFFX2 U10147 ( .INP(n10434), .Z(n10179) );
  NBUFFX2 U10148 ( .INP(n10434), .Z(n10180) );
  NBUFFX2 U10149 ( .INP(n10434), .Z(n10181) );
  NBUFFX2 U10150 ( .INP(n10433), .Z(n10182) );
  NBUFFX2 U10151 ( .INP(n10433), .Z(n10183) );
  NBUFFX2 U10152 ( .INP(n10433), .Z(n10184) );
  NBUFFX2 U10153 ( .INP(n10432), .Z(n10185) );
  NBUFFX2 U10154 ( .INP(n10432), .Z(n10186) );
  NBUFFX2 U10155 ( .INP(n10432), .Z(n10187) );
  NBUFFX2 U10156 ( .INP(n10431), .Z(n10188) );
  NBUFFX2 U10157 ( .INP(n10431), .Z(n10189) );
  NBUFFX2 U10158 ( .INP(n10431), .Z(n10190) );
  NBUFFX2 U10159 ( .INP(n10430), .Z(n10191) );
  NBUFFX2 U10160 ( .INP(n10430), .Z(n10192) );
  NBUFFX2 U10161 ( .INP(n10430), .Z(n10193) );
  NBUFFX2 U10162 ( .INP(n10429), .Z(n10194) );
  NBUFFX2 U10163 ( .INP(n10429), .Z(n10195) );
  NBUFFX2 U10164 ( .INP(n10429), .Z(n10196) );
  NBUFFX2 U10165 ( .INP(n10428), .Z(n10197) );
  NBUFFX2 U10166 ( .INP(n10428), .Z(n10198) );
  NBUFFX2 U10167 ( .INP(n10428), .Z(n10199) );
  NBUFFX2 U10168 ( .INP(n10427), .Z(n10200) );
  NBUFFX2 U10169 ( .INP(n10427), .Z(n10201) );
  NBUFFX2 U10170 ( .INP(n10427), .Z(n10202) );
  NBUFFX2 U10171 ( .INP(n10426), .Z(n10203) );
  NBUFFX2 U10172 ( .INP(n10426), .Z(n10204) );
  NBUFFX2 U10173 ( .INP(n10426), .Z(n10205) );
  NBUFFX2 U10174 ( .INP(n10425), .Z(n10206) );
  NBUFFX2 U10175 ( .INP(n10425), .Z(n10207) );
  NBUFFX2 U10176 ( .INP(n10425), .Z(n10208) );
  NBUFFX2 U10177 ( .INP(n10424), .Z(n10209) );
  NBUFFX2 U10178 ( .INP(n10424), .Z(n10210) );
  NBUFFX2 U10179 ( .INP(n10424), .Z(n10211) );
  NBUFFX2 U10180 ( .INP(n10423), .Z(n10212) );
  NBUFFX2 U10181 ( .INP(n10423), .Z(n10213) );
  NBUFFX2 U10182 ( .INP(n10423), .Z(n10214) );
  NBUFFX2 U10183 ( .INP(n10422), .Z(n10215) );
  NBUFFX2 U10184 ( .INP(n10422), .Z(n10216) );
  NBUFFX2 U10185 ( .INP(n10422), .Z(n10217) );
  NBUFFX2 U10186 ( .INP(n10421), .Z(n10218) );
  NBUFFX2 U10187 ( .INP(n10421), .Z(n10219) );
  NBUFFX2 U10188 ( .INP(n10421), .Z(n10220) );
  NBUFFX2 U10189 ( .INP(n10420), .Z(n10221) );
  NBUFFX2 U10190 ( .INP(n10420), .Z(n10222) );
  NBUFFX2 U10191 ( .INP(n10420), .Z(n10223) );
  NBUFFX2 U10192 ( .INP(n10419), .Z(n10224) );
  NBUFFX2 U10193 ( .INP(n10419), .Z(n10225) );
  NBUFFX2 U10194 ( .INP(n10419), .Z(n10226) );
  NBUFFX2 U10195 ( .INP(n10418), .Z(n10227) );
  NBUFFX2 U10196 ( .INP(n10418), .Z(n10228) );
  NBUFFX2 U10197 ( .INP(n10418), .Z(n10229) );
  NBUFFX2 U10198 ( .INP(n10417), .Z(n10230) );
  NBUFFX2 U10199 ( .INP(n10417), .Z(n10231) );
  NBUFFX2 U10200 ( .INP(n10417), .Z(n10232) );
  NBUFFX2 U10201 ( .INP(n10416), .Z(n10233) );
  NBUFFX2 U10202 ( .INP(n10416), .Z(n10234) );
  NBUFFX2 U10203 ( .INP(n10416), .Z(n10235) );
  NBUFFX2 U10204 ( .INP(n10415), .Z(n10236) );
  NBUFFX2 U10205 ( .INP(n10415), .Z(n10237) );
  NBUFFX2 U10206 ( .INP(n10415), .Z(n10238) );
  NBUFFX2 U10207 ( .INP(n10414), .Z(n10239) );
  NBUFFX2 U10208 ( .INP(n10414), .Z(n10240) );
  NBUFFX2 U10209 ( .INP(n10414), .Z(n10241) );
  NBUFFX2 U10210 ( .INP(n10413), .Z(n10242) );
  NBUFFX2 U10211 ( .INP(n10413), .Z(n10243) );
  NBUFFX2 U10212 ( .INP(n10413), .Z(n10244) );
  NBUFFX2 U10213 ( .INP(n10412), .Z(n10245) );
  NBUFFX2 U10214 ( .INP(n10412), .Z(n10246) );
  NBUFFX2 U10215 ( .INP(n10412), .Z(n10247) );
  NBUFFX2 U10216 ( .INP(n10411), .Z(n10248) );
  NBUFFX2 U10217 ( .INP(n10411), .Z(n10249) );
  NBUFFX2 U10218 ( .INP(n10411), .Z(n10250) );
  NBUFFX2 U10219 ( .INP(n10410), .Z(n10251) );
  NBUFFX2 U10220 ( .INP(n10410), .Z(n10252) );
  NBUFFX2 U10221 ( .INP(n10410), .Z(n10253) );
  NBUFFX2 U10222 ( .INP(n10409), .Z(n10254) );
  NBUFFX2 U10223 ( .INP(n10409), .Z(n10255) );
  NBUFFX2 U10224 ( .INP(n10409), .Z(n10256) );
  NBUFFX2 U10225 ( .INP(n10408), .Z(n10257) );
  NBUFFX2 U10226 ( .INP(n10408), .Z(n10258) );
  NBUFFX2 U10227 ( .INP(n10408), .Z(n10259) );
  NBUFFX2 U10228 ( .INP(n10407), .Z(n10260) );
  NBUFFX2 U10229 ( .INP(n10407), .Z(n10261) );
  NBUFFX2 U10230 ( .INP(n10407), .Z(n10262) );
  NBUFFX2 U10231 ( .INP(n10406), .Z(n10263) );
  NBUFFX2 U10232 ( .INP(n10406), .Z(n10264) );
  NBUFFX2 U10233 ( .INP(n10406), .Z(n10265) );
  NBUFFX2 U10234 ( .INP(n10405), .Z(n10266) );
  NBUFFX2 U10235 ( .INP(n10405), .Z(n10267) );
  NBUFFX2 U10236 ( .INP(n10405), .Z(n10268) );
  NBUFFX2 U10237 ( .INP(n10404), .Z(n10269) );
  NBUFFX2 U10238 ( .INP(n10404), .Z(n10270) );
  NBUFFX2 U10239 ( .INP(n10404), .Z(n10271) );
  NBUFFX2 U10240 ( .INP(n10403), .Z(n10272) );
  NBUFFX2 U10241 ( .INP(n10403), .Z(n10273) );
  NBUFFX2 U10242 ( .INP(n10403), .Z(n10274) );
  NBUFFX2 U10243 ( .INP(n10402), .Z(n10275) );
  NBUFFX2 U10244 ( .INP(n10402), .Z(n10276) );
  NBUFFX2 U10245 ( .INP(n10402), .Z(n10277) );
  NBUFFX2 U10246 ( .INP(n10401), .Z(n10278) );
  NBUFFX2 U10247 ( .INP(n10401), .Z(n10279) );
  NBUFFX2 U10248 ( .INP(n10401), .Z(n10280) );
  NBUFFX2 U10249 ( .INP(n10400), .Z(n10281) );
  NBUFFX2 U10250 ( .INP(n10400), .Z(n10282) );
  NBUFFX2 U10251 ( .INP(n10400), .Z(n10283) );
  NBUFFX2 U10252 ( .INP(n10399), .Z(n10284) );
  NBUFFX2 U10253 ( .INP(n10399), .Z(n10285) );
  NBUFFX2 U10254 ( .INP(n10399), .Z(n10286) );
  NBUFFX2 U10255 ( .INP(n10398), .Z(n10287) );
  NBUFFX2 U10256 ( .INP(n10398), .Z(n10288) );
  NBUFFX2 U10257 ( .INP(n10398), .Z(n10289) );
  NBUFFX2 U10258 ( .INP(n10397), .Z(n10290) );
  NBUFFX2 U10259 ( .INP(n10397), .Z(n10291) );
  NBUFFX2 U10260 ( .INP(n10397), .Z(n10292) );
  NBUFFX2 U10261 ( .INP(n10396), .Z(n10293) );
  NBUFFX2 U10262 ( .INP(n10396), .Z(n10294) );
  NBUFFX2 U10263 ( .INP(n10396), .Z(n10295) );
  NBUFFX2 U10264 ( .INP(n10395), .Z(n10296) );
  NBUFFX2 U10265 ( .INP(n10395), .Z(n10297) );
  NBUFFX2 U10266 ( .INP(n10395), .Z(n10298) );
  NBUFFX2 U10267 ( .INP(n10394), .Z(n10299) );
  NBUFFX2 U10268 ( .INP(n10394), .Z(n10300) );
  NBUFFX2 U10269 ( .INP(n10394), .Z(n10301) );
  NBUFFX2 U10270 ( .INP(n10393), .Z(n10302) );
  NBUFFX2 U10271 ( .INP(n10393), .Z(n10303) );
  NBUFFX2 U10272 ( .INP(n10393), .Z(n10304) );
  NBUFFX2 U10273 ( .INP(n10392), .Z(n10305) );
  NBUFFX2 U10274 ( .INP(n10392), .Z(n10306) );
  NBUFFX2 U10275 ( .INP(n10392), .Z(n10307) );
  NBUFFX2 U10276 ( .INP(n10391), .Z(n10308) );
  NBUFFX2 U10277 ( .INP(n10391), .Z(n10309) );
  NBUFFX2 U10278 ( .INP(n10391), .Z(n10310) );
  NBUFFX2 U10279 ( .INP(n10390), .Z(n10311) );
  NBUFFX2 U10280 ( .INP(n10390), .Z(n10312) );
  NBUFFX2 U10281 ( .INP(n10390), .Z(n10313) );
  NBUFFX2 U10282 ( .INP(n10389), .Z(n10314) );
  NBUFFX2 U10283 ( .INP(n10389), .Z(n10315) );
  NBUFFX2 U10284 ( .INP(n10389), .Z(n10316) );
  NBUFFX2 U10285 ( .INP(n10388), .Z(n10317) );
  NBUFFX2 U10286 ( .INP(n10388), .Z(n10318) );
  NBUFFX2 U10287 ( .INP(n10388), .Z(n10319) );
  NBUFFX2 U10288 ( .INP(n10387), .Z(n10320) );
  NBUFFX2 U10289 ( .INP(n10387), .Z(n10321) );
  NBUFFX2 U10290 ( .INP(n10387), .Z(n10322) );
  NBUFFX2 U10291 ( .INP(n10386), .Z(n10323) );
  NBUFFX2 U10292 ( .INP(n10386), .Z(n10324) );
  NBUFFX2 U10293 ( .INP(n10386), .Z(n10325) );
  NBUFFX2 U10294 ( .INP(n10385), .Z(n10326) );
  NBUFFX2 U10295 ( .INP(n10385), .Z(n10327) );
  NBUFFX2 U10296 ( .INP(n10385), .Z(n10328) );
  NBUFFX2 U10297 ( .INP(n10384), .Z(n10329) );
  NBUFFX2 U10298 ( .INP(n10384), .Z(n10330) );
  NBUFFX2 U10299 ( .INP(n10384), .Z(n10331) );
  NBUFFX2 U10300 ( .INP(n10383), .Z(n10332) );
  NBUFFX2 U10301 ( .INP(n10383), .Z(n10333) );
  NBUFFX2 U10302 ( .INP(n10383), .Z(n10334) );
  NBUFFX2 U10303 ( .INP(n10382), .Z(n10335) );
  NBUFFX2 U10304 ( .INP(n10382), .Z(n10336) );
  NBUFFX2 U10305 ( .INP(n10382), .Z(n10337) );
  NBUFFX2 U10306 ( .INP(n10381), .Z(n10338) );
  NBUFFX2 U10307 ( .INP(n10381), .Z(n10339) );
  NBUFFX2 U10308 ( .INP(n10381), .Z(n10340) );
  NBUFFX2 U10309 ( .INP(n10380), .Z(n10341) );
  NBUFFX2 U10310 ( .INP(n10380), .Z(n10342) );
  NBUFFX2 U10311 ( .INP(n10380), .Z(n10343) );
  NBUFFX2 U10312 ( .INP(n10379), .Z(n10344) );
  NBUFFX2 U10313 ( .INP(n10379), .Z(n10345) );
  NBUFFX2 U10314 ( .INP(n10379), .Z(n10346) );
  NBUFFX2 U10315 ( .INP(n10378), .Z(n10347) );
  NBUFFX2 U10316 ( .INP(n10378), .Z(n10348) );
  NBUFFX2 U10317 ( .INP(n10378), .Z(n10349) );
  NBUFFX2 U10318 ( .INP(n10377), .Z(n10350) );
  NBUFFX2 U10319 ( .INP(n10377), .Z(n10351) );
  NBUFFX2 U10320 ( .INP(n10377), .Z(n10352) );
  NBUFFX2 U10321 ( .INP(n10376), .Z(n10353) );
  NBUFFX2 U10322 ( .INP(n10376), .Z(n10354) );
  NBUFFX2 U10323 ( .INP(n10376), .Z(n10355) );
  NBUFFX2 U10324 ( .INP(n10375), .Z(n10356) );
  NBUFFX2 U10325 ( .INP(n10375), .Z(n10357) );
  NBUFFX2 U10326 ( .INP(n10375), .Z(n10358) );
  NBUFFX2 U10327 ( .INP(n10374), .Z(n10359) );
  NBUFFX2 U10328 ( .INP(n10374), .Z(n10360) );
  NBUFFX2 U10329 ( .INP(n10374), .Z(n10361) );
  NBUFFX2 U10330 ( .INP(n10373), .Z(n10362) );
  NBUFFX2 U10331 ( .INP(n10373), .Z(n10363) );
  NBUFFX2 U10332 ( .INP(n10373), .Z(n10364) );
  NBUFFX2 U10333 ( .INP(n10372), .Z(n10365) );
  NBUFFX2 U10334 ( .INP(n10372), .Z(n10366) );
  NBUFFX2 U10335 ( .INP(n10372), .Z(n10367) );
  NBUFFX2 U10336 ( .INP(n10371), .Z(n10368) );
  NBUFFX2 U10337 ( .INP(n10371), .Z(n10369) );
  NBUFFX2 U10338 ( .INP(n10371), .Z(n10370) );
  NBUFFX2 U10339 ( .INP(n10498), .Z(n10371) );
  NBUFFX2 U10340 ( .INP(n10498), .Z(n10372) );
  NBUFFX2 U10341 ( .INP(n10498), .Z(n10373) );
  NBUFFX2 U10342 ( .INP(n10497), .Z(n10374) );
  NBUFFX2 U10343 ( .INP(n10497), .Z(n10375) );
  NBUFFX2 U10344 ( .INP(n10497), .Z(n10376) );
  NBUFFX2 U10345 ( .INP(n10496), .Z(n10377) );
  NBUFFX2 U10346 ( .INP(n10496), .Z(n10378) );
  NBUFFX2 U10347 ( .INP(n10496), .Z(n10379) );
  NBUFFX2 U10348 ( .INP(n10495), .Z(n10380) );
  NBUFFX2 U10349 ( .INP(n10495), .Z(n10381) );
  NBUFFX2 U10350 ( .INP(n10495), .Z(n10382) );
  NBUFFX2 U10351 ( .INP(n10494), .Z(n10383) );
  NBUFFX2 U10352 ( .INP(n10494), .Z(n10384) );
  NBUFFX2 U10353 ( .INP(n10494), .Z(n10385) );
  NBUFFX2 U10354 ( .INP(n10493), .Z(n10386) );
  NBUFFX2 U10355 ( .INP(n10493), .Z(n10387) );
  NBUFFX2 U10356 ( .INP(n10493), .Z(n10388) );
  NBUFFX2 U10357 ( .INP(n10492), .Z(n10389) );
  NBUFFX2 U10358 ( .INP(n10492), .Z(n10390) );
  NBUFFX2 U10359 ( .INP(n10492), .Z(n10391) );
  NBUFFX2 U10360 ( .INP(n10491), .Z(n10392) );
  NBUFFX2 U10361 ( .INP(n10491), .Z(n10393) );
  NBUFFX2 U10362 ( .INP(n10491), .Z(n10394) );
  NBUFFX2 U10363 ( .INP(n10490), .Z(n10395) );
  NBUFFX2 U10364 ( .INP(n10490), .Z(n10396) );
  NBUFFX2 U10365 ( .INP(n10490), .Z(n10397) );
  NBUFFX2 U10366 ( .INP(n10489), .Z(n10398) );
  NBUFFX2 U10367 ( .INP(n10489), .Z(n10399) );
  NBUFFX2 U10368 ( .INP(n10489), .Z(n10400) );
  NBUFFX2 U10369 ( .INP(n10488), .Z(n10401) );
  NBUFFX2 U10370 ( .INP(n10488), .Z(n10402) );
  NBUFFX2 U10371 ( .INP(n10488), .Z(n10403) );
  NBUFFX2 U10372 ( .INP(n10487), .Z(n10404) );
  NBUFFX2 U10373 ( .INP(n10487), .Z(n10405) );
  NBUFFX2 U10374 ( .INP(n10487), .Z(n10406) );
  NBUFFX2 U10375 ( .INP(n10486), .Z(n10407) );
  NBUFFX2 U10376 ( .INP(n10486), .Z(n10408) );
  NBUFFX2 U10377 ( .INP(n10486), .Z(n10409) );
  NBUFFX2 U10378 ( .INP(n10485), .Z(n10410) );
  NBUFFX2 U10379 ( .INP(n10485), .Z(n10411) );
  NBUFFX2 U10380 ( .INP(n10485), .Z(n10412) );
  NBUFFX2 U10381 ( .INP(n10484), .Z(n10413) );
  NBUFFX2 U10382 ( .INP(n10484), .Z(n10414) );
  NBUFFX2 U10383 ( .INP(n10484), .Z(n10415) );
  NBUFFX2 U10384 ( .INP(n10483), .Z(n10416) );
  NBUFFX2 U10385 ( .INP(n10483), .Z(n10417) );
  NBUFFX2 U10386 ( .INP(n10483), .Z(n10418) );
  NBUFFX2 U10387 ( .INP(n10482), .Z(n10419) );
  NBUFFX2 U10388 ( .INP(n10482), .Z(n10420) );
  NBUFFX2 U10389 ( .INP(n10482), .Z(n10421) );
  NBUFFX2 U10390 ( .INP(n10481), .Z(n10422) );
  NBUFFX2 U10391 ( .INP(n10481), .Z(n10423) );
  NBUFFX2 U10392 ( .INP(n10481), .Z(n10424) );
  NBUFFX2 U10393 ( .INP(n10480), .Z(n10425) );
  NBUFFX2 U10394 ( .INP(n10480), .Z(n10426) );
  NBUFFX2 U10395 ( .INP(n10480), .Z(n10427) );
  NBUFFX2 U10396 ( .INP(n10479), .Z(n10428) );
  NBUFFX2 U10397 ( .INP(n10479), .Z(n10429) );
  NBUFFX2 U10398 ( .INP(n10479), .Z(n10430) );
  NBUFFX2 U10399 ( .INP(n10478), .Z(n10431) );
  NBUFFX2 U10400 ( .INP(n10478), .Z(n10432) );
  NBUFFX2 U10401 ( .INP(n10478), .Z(n10433) );
  NBUFFX2 U10402 ( .INP(n10477), .Z(n10434) );
  NBUFFX2 U10403 ( .INP(n10477), .Z(n10435) );
  NBUFFX2 U10404 ( .INP(n10477), .Z(n10436) );
  NBUFFX2 U10405 ( .INP(n10476), .Z(n10437) );
  NBUFFX2 U10406 ( .INP(n10476), .Z(n10438) );
  NBUFFX2 U10407 ( .INP(n10476), .Z(n10439) );
  NBUFFX2 U10408 ( .INP(n10475), .Z(n10440) );
  NBUFFX2 U10409 ( .INP(n10475), .Z(n10441) );
  NBUFFX2 U10410 ( .INP(n10475), .Z(n10442) );
  NBUFFX2 U10411 ( .INP(n10474), .Z(n10443) );
  NBUFFX2 U10412 ( .INP(n10474), .Z(n10444) );
  NBUFFX2 U10413 ( .INP(n10474), .Z(n10445) );
  NBUFFX2 U10414 ( .INP(n10473), .Z(n10446) );
  NBUFFX2 U10415 ( .INP(n10473), .Z(n10447) );
  NBUFFX2 U10416 ( .INP(n10473), .Z(n10448) );
  NBUFFX2 U10417 ( .INP(n10472), .Z(n10449) );
  NBUFFX2 U10418 ( .INP(n10472), .Z(n10450) );
  NBUFFX2 U10419 ( .INP(n10472), .Z(n10451) );
  NBUFFX2 U10420 ( .INP(n10471), .Z(n10452) );
  NBUFFX2 U10421 ( .INP(n10471), .Z(n10453) );
  NBUFFX2 U10422 ( .INP(n10471), .Z(n10454) );
  NBUFFX2 U10423 ( .INP(n10470), .Z(n10455) );
  NBUFFX2 U10424 ( .INP(n10470), .Z(n10456) );
  NBUFFX2 U10425 ( .INP(n10470), .Z(n10457) );
  NBUFFX2 U10426 ( .INP(n10469), .Z(n10458) );
  NBUFFX2 U10427 ( .INP(n10469), .Z(n10459) );
  NBUFFX2 U10428 ( .INP(n10469), .Z(n10460) );
  NBUFFX2 U10429 ( .INP(n10468), .Z(n10461) );
  NBUFFX2 U10430 ( .INP(n10468), .Z(n10462) );
  NBUFFX2 U10431 ( .INP(n10468), .Z(n10463) );
  NBUFFX2 U10432 ( .INP(n10467), .Z(n10464) );
  NBUFFX2 U10433 ( .INP(n10467), .Z(n10465) );
  NBUFFX2 U10434 ( .INP(n10467), .Z(n10466) );
  NBUFFX2 U10435 ( .INP(n10509), .Z(n10467) );
  NBUFFX2 U10436 ( .INP(n10509), .Z(n10468) );
  NBUFFX2 U10437 ( .INP(n10508), .Z(n10469) );
  NBUFFX2 U10438 ( .INP(n10508), .Z(n10470) );
  NBUFFX2 U10439 ( .INP(n10508), .Z(n10471) );
  NBUFFX2 U10440 ( .INP(n10507), .Z(n10472) );
  NBUFFX2 U10441 ( .INP(n10507), .Z(n10473) );
  NBUFFX2 U10442 ( .INP(n10507), .Z(n10474) );
  NBUFFX2 U10443 ( .INP(n10506), .Z(n10475) );
  NBUFFX2 U10444 ( .INP(n10506), .Z(n10476) );
  NBUFFX2 U10445 ( .INP(n10506), .Z(n10477) );
  NBUFFX2 U10446 ( .INP(n10505), .Z(n10478) );
  NBUFFX2 U10447 ( .INP(n10505), .Z(n10479) );
  NBUFFX2 U10448 ( .INP(n10505), .Z(n10480) );
  NBUFFX2 U10449 ( .INP(n10504), .Z(n10481) );
  NBUFFX2 U10450 ( .INP(n10504), .Z(n10482) );
  NBUFFX2 U10451 ( .INP(n10504), .Z(n10483) );
  NBUFFX2 U10452 ( .INP(n10503), .Z(n10484) );
  NBUFFX2 U10453 ( .INP(n10503), .Z(n10485) );
  NBUFFX2 U10454 ( .INP(n10503), .Z(n10486) );
  NBUFFX2 U10455 ( .INP(n10502), .Z(n10487) );
  NBUFFX2 U10456 ( .INP(n10502), .Z(n10488) );
  NBUFFX2 U10457 ( .INP(n10502), .Z(n10489) );
  NBUFFX2 U10458 ( .INP(n10501), .Z(n10490) );
  NBUFFX2 U10459 ( .INP(n10501), .Z(n10491) );
  NBUFFX2 U10460 ( .INP(n10501), .Z(n10492) );
  NBUFFX2 U10461 ( .INP(n10500), .Z(n10493) );
  NBUFFX2 U10462 ( .INP(n10500), .Z(n10494) );
  NBUFFX2 U10463 ( .INP(n10500), .Z(n10495) );
  NBUFFX2 U10464 ( .INP(n10499), .Z(n10496) );
  NBUFFX2 U10465 ( .INP(n10499), .Z(n10497) );
  NBUFFX2 U10466 ( .INP(n10499), .Z(n10498) );
  NBUFFX2 U10467 ( .INP(n10513), .Z(n10499) );
  NBUFFX2 U10468 ( .INP(n10513), .Z(n10500) );
  NBUFFX2 U10469 ( .INP(n10512), .Z(n10501) );
  NBUFFX2 U10470 ( .INP(n10512), .Z(n10502) );
  NBUFFX2 U10471 ( .INP(n10512), .Z(n10503) );
  NBUFFX2 U10472 ( .INP(n10511), .Z(n10504) );
  NBUFFX2 U10473 ( .INP(n10511), .Z(n10505) );
  NBUFFX2 U10474 ( .INP(n10511), .Z(n10506) );
  NBUFFX2 U10475 ( .INP(n10510), .Z(n10507) );
  NBUFFX2 U10476 ( .INP(n10510), .Z(n10508) );
  NBUFFX2 U10477 ( .INP(n10510), .Z(n10509) );
  NBUFFX2 U10478 ( .INP(test_se), .Z(n10510) );
  NBUFFX2 U10479 ( .INP(test_se), .Z(n10511) );
  NBUFFX2 U10480 ( .INP(test_se), .Z(n10512) );
  NBUFFX2 U10481 ( .INP(test_se), .Z(n10513) );
  NBUFFX2 U10482 ( .INP(n10536), .Z(n10514) );
  NBUFFX2 U10483 ( .INP(n10536), .Z(n10515) );
  NBUFFX2 U10484 ( .INP(n10535), .Z(n10516) );
  NBUFFX2 U10485 ( .INP(n10535), .Z(n10517) );
  NBUFFX2 U10486 ( .INP(n10535), .Z(n10518) );
  NBUFFX2 U10487 ( .INP(n10534), .Z(n10519) );
  NBUFFX2 U10488 ( .INP(n10534), .Z(n10520) );
  NBUFFX2 U10489 ( .INP(n10534), .Z(n10521) );
  NBUFFX2 U10490 ( .INP(n10533), .Z(n10522) );
  NBUFFX2 U10491 ( .INP(n10533), .Z(n10523) );
  NBUFFX2 U10492 ( .INP(n10533), .Z(n10524) );
  NBUFFX2 U10493 ( .INP(n10532), .Z(n10525) );
  NBUFFX2 U10494 ( .INP(n10532), .Z(n10526) );
  NBUFFX2 U10495 ( .INP(n10532), .Z(n10527) );
  NBUFFX2 U10496 ( .INP(n10531), .Z(n10528) );
  NBUFFX2 U10497 ( .INP(n10531), .Z(n10529) );
  NBUFFX2 U10498 ( .INP(n10531), .Z(n10530) );
  NBUFFX2 U10499 ( .INP(TM1), .Z(n10531) );
  NBUFFX2 U10500 ( .INP(TM1), .Z(n10532) );
  NBUFFX2 U10501 ( .INP(TM1), .Z(n10533) );
  NBUFFX2 U10502 ( .INP(TM1), .Z(n10534) );
  NBUFFX2 U10503 ( .INP(TM1), .Z(n10535) );
  NBUFFX2 U10504 ( .INP(TM1), .Z(n10536) );
  INVX0 U10505 ( .INP(n10517), .ZN(n10537) );
  INVX0 U10506 ( .INP(n10517), .ZN(n10538) );
  INVX0 U10507 ( .INP(n10517), .ZN(n10539) );
  INVX0 U10508 ( .INP(n10516), .ZN(n10540) );
  INVX0 U10509 ( .INP(n10517), .ZN(n10541) );
  INVX0 U10510 ( .INP(n10517), .ZN(n10542) );
  INVX0 U10511 ( .INP(n10516), .ZN(n10543) );
  INVX0 U10512 ( .INP(n10516), .ZN(n10544) );
  INVX0 U10513 ( .INP(n10517), .ZN(n10545) );
  NBUFFX2 U10514 ( .INP(n10621), .Z(n10546) );
  NBUFFX2 U10515 ( .INP(n10621), .Z(n10547) );
  NBUFFX2 U10516 ( .INP(n10621), .Z(n10548) );
  NBUFFX2 U10517 ( .INP(n10620), .Z(n10549) );
  NBUFFX2 U10518 ( .INP(n10620), .Z(n10550) );
  NBUFFX2 U10519 ( .INP(n10620), .Z(n10551) );
  NBUFFX2 U10520 ( .INP(n10619), .Z(n10552) );
  NBUFFX2 U10521 ( .INP(n10619), .Z(n10553) );
  NBUFFX2 U10522 ( .INP(n10619), .Z(n10554) );
  NBUFFX2 U10523 ( .INP(n10618), .Z(n10555) );
  NBUFFX2 U10524 ( .INP(n10618), .Z(n10556) );
  NBUFFX2 U10525 ( .INP(n10618), .Z(n10557) );
  NBUFFX2 U10526 ( .INP(n10617), .Z(n10558) );
  NBUFFX2 U10527 ( .INP(n10617), .Z(n10559) );
  NBUFFX2 U10528 ( .INP(n10617), .Z(n10560) );
  NBUFFX2 U10529 ( .INP(n10616), .Z(n10561) );
  NBUFFX2 U10530 ( .INP(n10616), .Z(n10562) );
  NBUFFX2 U10531 ( .INP(n10616), .Z(n10563) );
  NBUFFX2 U10532 ( .INP(n10615), .Z(n10564) );
  NBUFFX2 U10533 ( .INP(n10615), .Z(n10565) );
  NBUFFX2 U10534 ( .INP(n10615), .Z(n10566) );
  NBUFFX2 U10535 ( .INP(n10614), .Z(n10567) );
  NBUFFX2 U10536 ( .INP(n10614), .Z(n10568) );
  NBUFFX2 U10537 ( .INP(n10614), .Z(n10569) );
  NBUFFX2 U10538 ( .INP(n10613), .Z(n10570) );
  NBUFFX2 U10539 ( .INP(n10613), .Z(n10571) );
  NBUFFX2 U10540 ( .INP(n10613), .Z(n10572) );
  NBUFFX2 U10541 ( .INP(n10612), .Z(n10573) );
  NBUFFX2 U10542 ( .INP(n10612), .Z(n10574) );
  NBUFFX2 U10543 ( .INP(n10612), .Z(n10575) );
  NBUFFX2 U10544 ( .INP(n10611), .Z(n10576) );
  NBUFFX2 U10545 ( .INP(n10611), .Z(n10577) );
  NBUFFX2 U10546 ( .INP(n10611), .Z(n10578) );
  NBUFFX2 U10547 ( .INP(n10610), .Z(n10579) );
  NBUFFX2 U10548 ( .INP(n10610), .Z(n10580) );
  NBUFFX2 U10549 ( .INP(n10610), .Z(n10581) );
  NBUFFX2 U10550 ( .INP(n10609), .Z(n10582) );
  NBUFFX2 U10551 ( .INP(n10609), .Z(n10583) );
  NBUFFX2 U10552 ( .INP(n10609), .Z(n10584) );
  NBUFFX2 U10553 ( .INP(n10608), .Z(n10585) );
  NBUFFX2 U10554 ( .INP(n10608), .Z(n10586) );
  NBUFFX2 U10555 ( .INP(n10608), .Z(n10587) );
  NBUFFX2 U10556 ( .INP(n10607), .Z(n10588) );
  NBUFFX2 U10557 ( .INP(n10607), .Z(n10589) );
  NBUFFX2 U10558 ( .INP(n10607), .Z(n10590) );
  NBUFFX2 U10559 ( .INP(n10606), .Z(n10591) );
  NBUFFX2 U10560 ( .INP(n10606), .Z(n10592) );
  NBUFFX2 U10561 ( .INP(n10606), .Z(n10593) );
  NBUFFX2 U10562 ( .INP(n10605), .Z(n10594) );
  NBUFFX2 U10563 ( .INP(n10605), .Z(n10595) );
  NBUFFX2 U10564 ( .INP(n10605), .Z(n10596) );
  NBUFFX2 U10565 ( .INP(n10604), .Z(n10597) );
  NBUFFX2 U10566 ( .INP(n10604), .Z(n10598) );
  NBUFFX2 U10567 ( .INP(n10604), .Z(n10599) );
  NBUFFX2 U10568 ( .INP(n10603), .Z(n10600) );
  NBUFFX2 U10569 ( .INP(n10603), .Z(n10601) );
  NBUFFX2 U10570 ( .INP(n10603), .Z(n10602) );
  NBUFFX2 U10571 ( .INP(n10628), .Z(n10603) );
  NBUFFX2 U10572 ( .INP(n10627), .Z(n10604) );
  NBUFFX2 U10573 ( .INP(n10627), .Z(n10605) );
  NBUFFX2 U10574 ( .INP(n10627), .Z(n10606) );
  NBUFFX2 U10575 ( .INP(n10626), .Z(n10607) );
  NBUFFX2 U10576 ( .INP(n10626), .Z(n10608) );
  NBUFFX2 U10577 ( .INP(n10626), .Z(n10609) );
  NBUFFX2 U10578 ( .INP(n10625), .Z(n10610) );
  NBUFFX2 U10579 ( .INP(n10625), .Z(n10611) );
  NBUFFX2 U10580 ( .INP(n10625), .Z(n10612) );
  NBUFFX2 U10581 ( .INP(n10624), .Z(n10613) );
  NBUFFX2 U10582 ( .INP(n10624), .Z(n10614) );
  NBUFFX2 U10583 ( .INP(n10624), .Z(n10615) );
  NBUFFX2 U10584 ( .INP(n10623), .Z(n10616) );
  NBUFFX2 U10585 ( .INP(n10623), .Z(n10617) );
  NBUFFX2 U10586 ( .INP(n10623), .Z(n10618) );
  NBUFFX2 U10587 ( .INP(n10622), .Z(n10619) );
  NBUFFX2 U10588 ( .INP(n10622), .Z(n10620) );
  NBUFFX2 U10589 ( .INP(n10622), .Z(n10621) );
  NBUFFX2 U10590 ( .INP(RESET), .Z(n10622) );
  NBUFFX2 U10591 ( .INP(RESET), .Z(n10623) );
  NBUFFX2 U10592 ( .INP(RESET), .Z(n10624) );
  NBUFFX2 U10593 ( .INP(RESET), .Z(n10625) );
  NBUFFX2 U10594 ( .INP(RESET), .Z(n10626) );
  NBUFFX2 U10595 ( .INP(RESET), .Z(n10627) );
  NBUFFX2 U10596 ( .INP(RESET), .Z(n10628) );
  INVX0 U10597 ( .INP(n10546), .ZN(n10629) );
  INVX0 U10598 ( .INP(n10546), .ZN(n10630) );
  INVX0 U10599 ( .INP(n10546), .ZN(n10631) );
  INVX0 U10600 ( .INP(n10546), .ZN(n10632) );
  INVX0 U10601 ( .INP(n10546), .ZN(n10633) );
  INVX0 U10602 ( .INP(n10546), .ZN(n10634) );
  INVX0 U10603 ( .INP(n10546), .ZN(n10635) );
  INVX0 U10604 ( .INP(n10546), .ZN(n10636) );
  INVX0 U10605 ( .INP(n10547), .ZN(n10637) );
  INVX0 U10606 ( .INP(n10547), .ZN(n10638) );
  INVX0 U10607 ( .INP(n10547), .ZN(n10639) );
  INVX0 U10608 ( .INP(n10547), .ZN(n10640) );
  INVX0 U10609 ( .INP(n10547), .ZN(n10641) );
  INVX0 U10610 ( .INP(n10547), .ZN(n10642) );
  INVX0 U10611 ( .INP(n10547), .ZN(n10643) );
  INVX0 U10612 ( .INP(n10547), .ZN(n10644) );
  INVX0 U10613 ( .INP(n10548), .ZN(n10645) );
  INVX0 U10614 ( .INP(n10548), .ZN(n10646) );
  INVX0 U10615 ( .INP(n10548), .ZN(n10647) );
  INVX0 U10616 ( .INP(n10548), .ZN(n10648) );
  INVX0 U10617 ( .INP(n10548), .ZN(n10649) );
  INVX0 U10618 ( .INP(n10548), .ZN(n10650) );
  INVX0 U10619 ( .INP(n10548), .ZN(n10651) );
  INVX0 U10620 ( .INP(n10548), .ZN(n10652) );
  INVX0 U10621 ( .INP(n10549), .ZN(n10653) );
  INVX0 U10622 ( .INP(n10549), .ZN(n10654) );
  INVX0 U10623 ( .INP(n10549), .ZN(n10655) );
  INVX0 U10624 ( .INP(n10549), .ZN(n10656) );
  INVX0 U10625 ( .INP(n10549), .ZN(n10657) );
  INVX0 U10626 ( .INP(n10549), .ZN(n10658) );
  INVX0 U10627 ( .INP(n10549), .ZN(n10659) );
  INVX0 U10628 ( .INP(n10549), .ZN(n10660) );
  INVX0 U10629 ( .INP(n10550), .ZN(n10661) );
  INVX0 U10630 ( .INP(n10550), .ZN(n10662) );
  INVX0 U10631 ( .INP(n10550), .ZN(n10663) );
  INVX0 U10632 ( .INP(n10550), .ZN(n10664) );
  INVX0 U10633 ( .INP(n10550), .ZN(n10665) );
  INVX0 U10634 ( .INP(n10550), .ZN(n10666) );
  INVX0 U10635 ( .INP(n10550), .ZN(n10667) );
  INVX0 U10636 ( .INP(n10551), .ZN(n10668) );
  INVX0 U10637 ( .INP(n10551), .ZN(n10669) );
  INVX0 U10638 ( .INP(n10551), .ZN(n10670) );
  INVX0 U10639 ( .INP(n10551), .ZN(n10671) );
  INVX0 U10640 ( .INP(n10551), .ZN(n10672) );
  INVX0 U10641 ( .INP(n10551), .ZN(n10673) );
  INVX0 U10642 ( .INP(n10551), .ZN(n10674) );
  INVX0 U10643 ( .INP(n10551), .ZN(n10675) );
  INVX0 U10644 ( .INP(n10552), .ZN(n10676) );
  INVX0 U10645 ( .INP(n10552), .ZN(n10677) );
  INVX0 U10646 ( .INP(n10552), .ZN(n10678) );
  INVX0 U10647 ( .INP(n10552), .ZN(n10679) );
  INVX0 U10648 ( .INP(n10552), .ZN(n10680) );
  INVX0 U10649 ( .INP(n10552), .ZN(n10681) );
  INVX0 U10650 ( .INP(n10552), .ZN(n10682) );
  INVX0 U10651 ( .INP(n10552), .ZN(n10683) );
  INVX0 U10652 ( .INP(n10553), .ZN(n10684) );
  INVX0 U10653 ( .INP(n10553), .ZN(n10685) );
  INVX0 U10654 ( .INP(n10553), .ZN(n10686) );
  INVX0 U10655 ( .INP(n10553), .ZN(n10687) );
  INVX0 U10656 ( .INP(n10553), .ZN(n10688) );
  INVX0 U10657 ( .INP(n10553), .ZN(n10689) );
  INVX0 U10658 ( .INP(n10553), .ZN(n10690) );
  INVX0 U10659 ( .INP(n10553), .ZN(n10691) );
  INVX0 U10660 ( .INP(n10554), .ZN(n10692) );
  INVX0 U10661 ( .INP(n10554), .ZN(n10693) );
  INVX0 U10662 ( .INP(n10554), .ZN(n10694) );
  INVX0 U10663 ( .INP(n10554), .ZN(n10695) );
  INVX0 U10664 ( .INP(n10554), .ZN(n10696) );
  INVX0 U10665 ( .INP(n10554), .ZN(n10697) );
  INVX0 U10666 ( .INP(n10554), .ZN(n10698) );
  INVX0 U10667 ( .INP(n10554), .ZN(n10699) );
  INVX0 U10668 ( .INP(n10555), .ZN(n10700) );
  INVX0 U10669 ( .INP(n10555), .ZN(n10701) );
  INVX0 U10670 ( .INP(n10555), .ZN(n10702) );
  INVX0 U10671 ( .INP(n10555), .ZN(n10703) );
  INVX0 U10672 ( .INP(n10550), .ZN(n10704) );
  NBUFFX2 U10673 ( .INP(n10887), .Z(n10849) );
  NBUFFX2 U10674 ( .INP(n10887), .Z(n10850) );
  NBUFFX2 U10675 ( .INP(n10886), .Z(n10851) );
  NBUFFX2 U10676 ( .INP(n10886), .Z(n10852) );
  NBUFFX2 U10677 ( .INP(n10886), .Z(n10853) );
  NBUFFX2 U10678 ( .INP(n10885), .Z(n10854) );
  NBUFFX2 U10679 ( .INP(n10885), .Z(n10855) );
  NBUFFX2 U10680 ( .INP(n10885), .Z(n10856) );
  NBUFFX2 U10681 ( .INP(n10884), .Z(n10857) );
  NBUFFX2 U10682 ( .INP(n10884), .Z(n10858) );
  NBUFFX2 U10683 ( .INP(n10884), .Z(n10859) );
  NBUFFX2 U10684 ( .INP(n10883), .Z(n10860) );
  NBUFFX2 U10685 ( .INP(n10883), .Z(n10861) );
  NBUFFX2 U10686 ( .INP(n10883), .Z(n10862) );
  NBUFFX2 U10687 ( .INP(n10882), .Z(n10863) );
  NBUFFX2 U10688 ( .INP(n10882), .Z(n10864) );
  NBUFFX2 U10689 ( .INP(n10882), .Z(n10865) );
  NBUFFX2 U10690 ( .INP(n10881), .Z(n10866) );
  NBUFFX2 U10691 ( .INP(n10881), .Z(n10867) );
  NBUFFX2 U10692 ( .INP(n10881), .Z(n10868) );
  NBUFFX2 U10693 ( .INP(n10880), .Z(n10869) );
  NBUFFX2 U10694 ( .INP(n10880), .Z(n10870) );
  NBUFFX2 U10695 ( .INP(n10880), .Z(n10871) );
  NBUFFX2 U10696 ( .INP(n10879), .Z(n10872) );
  NBUFFX2 U10697 ( .INP(n10879), .Z(n10873) );
  NBUFFX2 U10698 ( .INP(n10879), .Z(n10874) );
  NBUFFX2 U10699 ( .INP(n10878), .Z(n10875) );
  NBUFFX2 U10700 ( .INP(n10878), .Z(n10876) );
  NBUFFX2 U10701 ( .INP(n10878), .Z(n10877) );
  NBUFFX2 U10702 ( .INP(CK), .Z(n10878) );
  NBUFFX2 U10703 ( .INP(CK), .Z(n10879) );
  NBUFFX2 U10704 ( .INP(n10887), .Z(n10880) );
  NBUFFX2 U10705 ( .INP(CK), .Z(n10881) );
  NBUFFX2 U10706 ( .INP(n10883), .Z(n10882) );
  NBUFFX2 U10707 ( .INP(CK), .Z(n10883) );
  NBUFFX2 U10708 ( .INP(n10878), .Z(n10884) );
  NBUFFX2 U10709 ( .INP(n10879), .Z(n10885) );
  NBUFFX2 U10710 ( .INP(n10881), .Z(n10886) );
  NBUFFX2 U10711 ( .INP(n10718), .Z(n10887) );
  AND2X1 U10712 ( .IN1(n10594), .IN2(n10545), .Q(n3278) );
  AND2X1 U10713 ( .IN1(n10594), .IN2(n8304), .Q(WX9789) );
  AND2X1 U10714 ( .IN1(n10594), .IN2(n8305), .Q(WX9787) );
  AND2X1 U10715 ( .IN1(n10594), .IN2(n8306), .Q(WX9785) );
  AND2X1 U10716 ( .IN1(n10594), .IN2(n8307), .Q(WX9783) );
  AND2X1 U10717 ( .IN1(test_so80), .IN2(n10570), .Q(WX9781) );
  AND2X1 U10718 ( .IN1(n10594), .IN2(n8310), .Q(WX9779) );
  AND2X1 U10719 ( .IN1(n10594), .IN2(n8311), .Q(WX9777) );
  AND2X1 U10720 ( .IN1(n10595), .IN2(n8312), .Q(WX9775) );
  AND2X1 U10721 ( .IN1(n10595), .IN2(n8313), .Q(WX9773) );
  AND2X1 U10722 ( .IN1(n10595), .IN2(n8314), .Q(WX9771) );
  AND2X1 U10723 ( .IN1(n10595), .IN2(n8315), .Q(WX9769) );
  AND2X1 U10724 ( .IN1(n10595), .IN2(n8316), .Q(WX9767) );
  AND2X1 U10725 ( .IN1(n10595), .IN2(n8317), .Q(WX9765) );
  AND2X1 U10726 ( .IN1(n10595), .IN2(n8318), .Q(WX9763) );
  AND2X1 U10727 ( .IN1(n10595), .IN2(n8319), .Q(WX9761) );
  AND2X1 U10728 ( .IN1(n10595), .IN2(n8320), .Q(WX9759) );
  OR2X1 U10729 ( .IN1(n10888), .IN2(n10889), .Q(WX9757) );
  OR2X1 U10730 ( .IN1(n10890), .IN2(n10891), .Q(n10889) );
  AND2X1 U10731 ( .IN1(n10028), .IN2(CRC_OUT_2_0), .Q(n10891) );
  AND2X1 U10732 ( .IN1(n10023), .IN2(n1727), .Q(n10890) );
  INVX0 U10733 ( .INP(n10892), .ZN(n1727) );
  OR2X1 U10734 ( .IN1(n10649), .IN2(n3817), .Q(n10892) );
  OR2X1 U10735 ( .IN1(n10893), .IN2(n10894), .Q(n10888) );
  AND2X1 U10736 ( .IN1(n10065), .IN2(n10895), .Q(n10894) );
  AND2X1 U10737 ( .IN1(n9984), .IN2(n10897), .Q(n10893) );
  OR2X1 U10738 ( .IN1(n10898), .IN2(n10899), .Q(WX9755) );
  OR2X1 U10739 ( .IN1(n10900), .IN2(n10901), .Q(n10899) );
  AND2X1 U10740 ( .IN1(n10042), .IN2(CRC_OUT_2_1), .Q(n10901) );
  AND2X1 U10741 ( .IN1(n1726), .IN2(n10011), .Q(n10900) );
  INVX0 U10742 ( .INP(n10902), .ZN(n1726) );
  OR2X1 U10743 ( .IN1(n10649), .IN2(n3818), .Q(n10902) );
  OR2X1 U10744 ( .IN1(n10903), .IN2(n10904), .Q(n10898) );
  AND2X1 U10745 ( .IN1(n10073), .IN2(n10905), .Q(n10904) );
  AND2X1 U10746 ( .IN1(n10906), .IN2(n9972), .Q(n10903) );
  OR2X1 U10747 ( .IN1(n10907), .IN2(n10908), .Q(WX9753) );
  OR2X1 U10748 ( .IN1(n10909), .IN2(n10910), .Q(n10908) );
  AND2X1 U10749 ( .IN1(test_so87), .IN2(n10026), .Q(n10910) );
  AND2X1 U10750 ( .IN1(n1725), .IN2(n10011), .Q(n10909) );
  INVX0 U10751 ( .INP(n10911), .ZN(n1725) );
  OR2X1 U10752 ( .IN1(n10649), .IN2(n3819), .Q(n10911) );
  OR2X1 U10753 ( .IN1(n10912), .IN2(n10913), .Q(n10907) );
  AND2X1 U10754 ( .IN1(n10914), .IN2(n10060), .Q(n10913) );
  AND2X1 U10755 ( .IN1(n9984), .IN2(n10915), .Q(n10912) );
  OR2X1 U10756 ( .IN1(n10916), .IN2(n10917), .Q(WX9751) );
  OR2X1 U10757 ( .IN1(n10918), .IN2(n10919), .Q(n10917) );
  AND2X1 U10758 ( .IN1(n10037), .IN2(CRC_OUT_2_3), .Q(n10919) );
  AND2X1 U10759 ( .IN1(n1724), .IN2(n10011), .Q(n10918) );
  INVX0 U10760 ( .INP(n10920), .ZN(n1724) );
  OR2X1 U10761 ( .IN1(n10649), .IN2(n3820), .Q(n10920) );
  OR2X1 U10762 ( .IN1(n10921), .IN2(n10922), .Q(n10916) );
  AND2X1 U10763 ( .IN1(n10069), .IN2(n10923), .Q(n10922) );
  AND2X1 U10764 ( .IN1(n10924), .IN2(n9972), .Q(n10921) );
  OR2X1 U10765 ( .IN1(n10925), .IN2(n10926), .Q(WX9749) );
  OR2X1 U10766 ( .IN1(n10927), .IN2(n10928), .Q(n10926) );
  AND2X1 U10767 ( .IN1(n10037), .IN2(CRC_OUT_2_4), .Q(n10928) );
  AND2X1 U10768 ( .IN1(n1723), .IN2(n10011), .Q(n10927) );
  INVX0 U10769 ( .INP(n10929), .ZN(n1723) );
  OR2X1 U10770 ( .IN1(n10649), .IN2(n3821), .Q(n10929) );
  OR2X1 U10771 ( .IN1(n10930), .IN2(n10931), .Q(n10925) );
  AND2X1 U10772 ( .IN1(n10932), .IN2(n10060), .Q(n10931) );
  AND2X1 U10773 ( .IN1(n9984), .IN2(n10933), .Q(n10930) );
  OR2X1 U10774 ( .IN1(n10934), .IN2(n10935), .Q(WX9747) );
  OR2X1 U10775 ( .IN1(n10936), .IN2(n10937), .Q(n10935) );
  AND2X1 U10776 ( .IN1(n10037), .IN2(CRC_OUT_2_5), .Q(n10937) );
  AND2X1 U10777 ( .IN1(n1722), .IN2(n10012), .Q(n10936) );
  INVX0 U10778 ( .INP(n10938), .ZN(n1722) );
  OR2X1 U10779 ( .IN1(n10649), .IN2(n3822), .Q(n10938) );
  OR2X1 U10780 ( .IN1(n10939), .IN2(n10940), .Q(n10934) );
  AND2X1 U10781 ( .IN1(n10069), .IN2(n10941), .Q(n10940) );
  AND2X1 U10782 ( .IN1(n9984), .IN2(n10942), .Q(n10939) );
  OR2X1 U10783 ( .IN1(n10943), .IN2(n10944), .Q(WX9745) );
  OR2X1 U10784 ( .IN1(n10945), .IN2(n10946), .Q(n10944) );
  AND2X1 U10785 ( .IN1(n10037), .IN2(CRC_OUT_2_6), .Q(n10946) );
  AND2X1 U10786 ( .IN1(n1721), .IN2(n10012), .Q(n10945) );
  INVX0 U10787 ( .INP(n10947), .ZN(n1721) );
  OR2X1 U10788 ( .IN1(n10649), .IN2(n3823), .Q(n10947) );
  OR2X1 U10789 ( .IN1(n10948), .IN2(n10949), .Q(n10943) );
  AND2X1 U10790 ( .IN1(n10950), .IN2(n10061), .Q(n10949) );
  AND2X1 U10791 ( .IN1(n9984), .IN2(n10951), .Q(n10948) );
  OR2X1 U10792 ( .IN1(n10952), .IN2(n10953), .Q(WX9743) );
  OR2X1 U10793 ( .IN1(n10954), .IN2(n10955), .Q(n10953) );
  AND2X1 U10794 ( .IN1(n10037), .IN2(CRC_OUT_2_7), .Q(n10955) );
  AND2X1 U10795 ( .IN1(n1720), .IN2(n10012), .Q(n10954) );
  INVX0 U10796 ( .INP(n10956), .ZN(n1720) );
  OR2X1 U10797 ( .IN1(n10649), .IN2(n3824), .Q(n10956) );
  OR2X1 U10798 ( .IN1(n10957), .IN2(n10958), .Q(n10952) );
  AND2X1 U10799 ( .IN1(n10069), .IN2(n10959), .Q(n10958) );
  AND2X1 U10800 ( .IN1(n9984), .IN2(n10960), .Q(n10957) );
  OR2X1 U10801 ( .IN1(n10961), .IN2(n10962), .Q(WX9741) );
  OR2X1 U10802 ( .IN1(n10963), .IN2(n10964), .Q(n10962) );
  AND2X1 U10803 ( .IN1(n10038), .IN2(CRC_OUT_2_8), .Q(n10964) );
  AND2X1 U10804 ( .IN1(n1719), .IN2(n10012), .Q(n10963) );
  INVX0 U10805 ( .INP(n10965), .ZN(n1719) );
  OR2X1 U10806 ( .IN1(n10648), .IN2(n3825), .Q(n10965) );
  OR2X1 U10807 ( .IN1(n10966), .IN2(n10967), .Q(n10961) );
  AND2X1 U10808 ( .IN1(n10968), .IN2(n10061), .Q(n10967) );
  AND2X1 U10809 ( .IN1(n9984), .IN2(n10969), .Q(n10966) );
  OR2X1 U10810 ( .IN1(n10970), .IN2(n10971), .Q(WX9739) );
  OR2X1 U10811 ( .IN1(n10972), .IN2(n10973), .Q(n10971) );
  AND2X1 U10812 ( .IN1(n10038), .IN2(CRC_OUT_2_9), .Q(n10973) );
  AND2X1 U10813 ( .IN1(n1718), .IN2(n10012), .Q(n10972) );
  INVX0 U10814 ( .INP(n10974), .ZN(n1718) );
  OR2X1 U10815 ( .IN1(n10648), .IN2(n3826), .Q(n10974) );
  OR2X1 U10816 ( .IN1(n10975), .IN2(n10976), .Q(n10970) );
  AND2X1 U10817 ( .IN1(n10069), .IN2(n10977), .Q(n10976) );
  AND2X1 U10818 ( .IN1(n9984), .IN2(n10978), .Q(n10975) );
  OR2X1 U10819 ( .IN1(n10979), .IN2(n10980), .Q(WX9737) );
  OR2X1 U10820 ( .IN1(n10981), .IN2(n10982), .Q(n10980) );
  AND2X1 U10821 ( .IN1(n10038), .IN2(CRC_OUT_2_10), .Q(n10982) );
  AND2X1 U10822 ( .IN1(n1717), .IN2(n10012), .Q(n10981) );
  INVX0 U10823 ( .INP(n10983), .ZN(n1717) );
  OR2X1 U10824 ( .IN1(n10648), .IN2(n3827), .Q(n10983) );
  OR2X1 U10825 ( .IN1(n10984), .IN2(n10985), .Q(n10979) );
  AND2X1 U10826 ( .IN1(n10069), .IN2(n10986), .Q(n10985) );
  AND2X1 U10827 ( .IN1(n9984), .IN2(n10987), .Q(n10984) );
  OR2X1 U10828 ( .IN1(n10988), .IN2(n10989), .Q(WX9735) );
  OR2X1 U10829 ( .IN1(n10990), .IN2(n10991), .Q(n10989) );
  AND2X1 U10830 ( .IN1(n10038), .IN2(CRC_OUT_2_11), .Q(n10991) );
  AND2X1 U10831 ( .IN1(n1716), .IN2(n10012), .Q(n10990) );
  INVX0 U10832 ( .INP(n10992), .ZN(n1716) );
  OR2X1 U10833 ( .IN1(n10648), .IN2(n3828), .Q(n10992) );
  OR2X1 U10834 ( .IN1(n10993), .IN2(n10994), .Q(n10988) );
  AND2X1 U10835 ( .IN1(n10069), .IN2(n10995), .Q(n10994) );
  AND2X1 U10836 ( .IN1(n9984), .IN2(n10996), .Q(n10993) );
  OR2X1 U10837 ( .IN1(n10997), .IN2(n10998), .Q(WX9733) );
  OR2X1 U10838 ( .IN1(n10999), .IN2(n11000), .Q(n10998) );
  AND2X1 U10839 ( .IN1(n10038), .IN2(CRC_OUT_2_12), .Q(n11000) );
  AND2X1 U10840 ( .IN1(n1715), .IN2(n10012), .Q(n10999) );
  INVX0 U10841 ( .INP(n11001), .ZN(n1715) );
  OR2X1 U10842 ( .IN1(n10648), .IN2(n3829), .Q(n11001) );
  OR2X1 U10843 ( .IN1(n11002), .IN2(n11003), .Q(n10997) );
  AND2X1 U10844 ( .IN1(n10069), .IN2(n11004), .Q(n11003) );
  AND2X1 U10845 ( .IN1(n9984), .IN2(n11005), .Q(n11002) );
  OR2X1 U10846 ( .IN1(n11006), .IN2(n11007), .Q(WX9731) );
  OR2X1 U10847 ( .IN1(n11008), .IN2(n11009), .Q(n11007) );
  AND2X1 U10848 ( .IN1(n10038), .IN2(CRC_OUT_2_13), .Q(n11009) );
  AND2X1 U10849 ( .IN1(n1714), .IN2(n10012), .Q(n11008) );
  INVX0 U10850 ( .INP(n11010), .ZN(n1714) );
  OR2X1 U10851 ( .IN1(n10648), .IN2(n3830), .Q(n11010) );
  OR2X1 U10852 ( .IN1(n11011), .IN2(n11012), .Q(n11006) );
  AND2X1 U10853 ( .IN1(n10069), .IN2(n11013), .Q(n11012) );
  AND2X1 U10854 ( .IN1(n9984), .IN2(n11014), .Q(n11011) );
  OR2X1 U10855 ( .IN1(n11015), .IN2(n11016), .Q(WX9729) );
  OR2X1 U10856 ( .IN1(n11017), .IN2(n11018), .Q(n11016) );
  AND2X1 U10857 ( .IN1(n10038), .IN2(CRC_OUT_2_14), .Q(n11018) );
  AND2X1 U10858 ( .IN1(n1713), .IN2(n10012), .Q(n11017) );
  INVX0 U10859 ( .INP(n11019), .ZN(n1713) );
  OR2X1 U10860 ( .IN1(n10648), .IN2(n3831), .Q(n11019) );
  OR2X1 U10861 ( .IN1(n11020), .IN2(n11021), .Q(n11015) );
  AND2X1 U10862 ( .IN1(n10069), .IN2(n11022), .Q(n11021) );
  AND2X1 U10863 ( .IN1(n11023), .IN2(n9973), .Q(n11020) );
  OR2X1 U10864 ( .IN1(n11024), .IN2(n11025), .Q(WX9727) );
  OR2X1 U10865 ( .IN1(n11026), .IN2(n11027), .Q(n11025) );
  AND2X1 U10866 ( .IN1(n10038), .IN2(CRC_OUT_2_15), .Q(n11027) );
  AND2X1 U10867 ( .IN1(n1712), .IN2(n10012), .Q(n11026) );
  INVX0 U10868 ( .INP(n11028), .ZN(n1712) );
  OR2X1 U10869 ( .IN1(n10648), .IN2(n3832), .Q(n11028) );
  OR2X1 U10870 ( .IN1(n11029), .IN2(n11030), .Q(n11024) );
  AND2X1 U10871 ( .IN1(n10069), .IN2(n11031), .Q(n11030) );
  AND2X1 U10872 ( .IN1(n9983), .IN2(n11032), .Q(n11029) );
  OR2X1 U10873 ( .IN1(n11033), .IN2(n11034), .Q(WX9725) );
  OR2X1 U10874 ( .IN1(n11035), .IN2(n11036), .Q(n11034) );
  AND2X1 U10875 ( .IN1(n10038), .IN2(CRC_OUT_2_16), .Q(n11036) );
  AND2X1 U10876 ( .IN1(n1711), .IN2(n10012), .Q(n11035) );
  INVX0 U10877 ( .INP(n11037), .ZN(n1711) );
  OR2X1 U10878 ( .IN1(n10648), .IN2(n3833), .Q(n11037) );
  OR2X1 U10879 ( .IN1(n11038), .IN2(n11039), .Q(n11033) );
  AND2X1 U10880 ( .IN1(n10069), .IN2(n11040), .Q(n11039) );
  AND2X1 U10881 ( .IN1(n11041), .IN2(n9973), .Q(n11038) );
  OR2X1 U10882 ( .IN1(n11042), .IN2(n11043), .Q(WX9723) );
  OR2X1 U10883 ( .IN1(n11044), .IN2(n11045), .Q(n11043) );
  AND2X1 U10884 ( .IN1(n10038), .IN2(CRC_OUT_2_17), .Q(n11045) );
  AND2X1 U10885 ( .IN1(n1710), .IN2(n10013), .Q(n11044) );
  INVX0 U10886 ( .INP(n11046), .ZN(n1710) );
  OR2X1 U10887 ( .IN1(n10648), .IN2(n3834), .Q(n11046) );
  OR2X1 U10888 ( .IN1(n11047), .IN2(n11048), .Q(n11042) );
  AND2X1 U10889 ( .IN1(n10070), .IN2(n11049), .Q(n11048) );
  AND2X1 U10890 ( .IN1(n9983), .IN2(n11050), .Q(n11047) );
  OR2X1 U10891 ( .IN1(n11051), .IN2(n11052), .Q(WX9721) );
  OR2X1 U10892 ( .IN1(n11053), .IN2(n11054), .Q(n11052) );
  AND2X1 U10893 ( .IN1(n10038), .IN2(CRC_OUT_2_18), .Q(n11054) );
  AND2X1 U10894 ( .IN1(n1709), .IN2(n10013), .Q(n11053) );
  INVX0 U10895 ( .INP(n11055), .ZN(n1709) );
  OR2X1 U10896 ( .IN1(n10648), .IN2(n3835), .Q(n11055) );
  OR2X1 U10897 ( .IN1(n11056), .IN2(n11057), .Q(n11051) );
  AND2X1 U10898 ( .IN1(n10070), .IN2(n11058), .Q(n11057) );
  AND2X1 U10899 ( .IN1(n11059), .IN2(n9973), .Q(n11056) );
  OR2X1 U10900 ( .IN1(n11060), .IN2(n11061), .Q(WX9719) );
  OR2X1 U10901 ( .IN1(n11062), .IN2(n11063), .Q(n11061) );
  AND2X1 U10902 ( .IN1(test_so88), .IN2(n10026), .Q(n11063) );
  AND2X1 U10903 ( .IN1(n1708), .IN2(n10013), .Q(n11062) );
  INVX0 U10904 ( .INP(n11064), .ZN(n1708) );
  OR2X1 U10905 ( .IN1(n10648), .IN2(n3836), .Q(n11064) );
  OR2X1 U10906 ( .IN1(n11065), .IN2(n11066), .Q(n11060) );
  AND2X1 U10907 ( .IN1(n11067), .IN2(n10063), .Q(n11066) );
  AND2X1 U10908 ( .IN1(n9983), .IN2(n11068), .Q(n11065) );
  OR2X1 U10909 ( .IN1(n11069), .IN2(n11070), .Q(WX9717) );
  OR2X1 U10910 ( .IN1(n11071), .IN2(n11072), .Q(n11070) );
  AND2X1 U10911 ( .IN1(n10038), .IN2(CRC_OUT_2_20), .Q(n11072) );
  AND2X1 U10912 ( .IN1(n1707), .IN2(n10013), .Q(n11071) );
  INVX0 U10913 ( .INP(n11073), .ZN(n1707) );
  OR2X1 U10914 ( .IN1(n10647), .IN2(n3837), .Q(n11073) );
  OR2X1 U10915 ( .IN1(n11074), .IN2(n11075), .Q(n11069) );
  AND2X1 U10916 ( .IN1(n10070), .IN2(n11076), .Q(n11075) );
  AND2X1 U10917 ( .IN1(n11077), .IN2(n9973), .Q(n11074) );
  OR2X1 U10918 ( .IN1(n11078), .IN2(n11079), .Q(WX9715) );
  OR2X1 U10919 ( .IN1(n11080), .IN2(n11081), .Q(n11079) );
  AND2X1 U10920 ( .IN1(n10038), .IN2(CRC_OUT_2_21), .Q(n11081) );
  AND2X1 U10921 ( .IN1(n1706), .IN2(n10013), .Q(n11080) );
  INVX0 U10922 ( .INP(n11082), .ZN(n1706) );
  OR2X1 U10923 ( .IN1(n10647), .IN2(n3838), .Q(n11082) );
  OR2X1 U10924 ( .IN1(n11083), .IN2(n11084), .Q(n11078) );
  AND2X1 U10925 ( .IN1(n11085), .IN2(n10062), .Q(n11084) );
  AND2X1 U10926 ( .IN1(n9983), .IN2(n11086), .Q(n11083) );
  OR2X1 U10927 ( .IN1(n11087), .IN2(n11088), .Q(WX9713) );
  OR2X1 U10928 ( .IN1(n11089), .IN2(n11090), .Q(n11088) );
  AND2X1 U10929 ( .IN1(n10039), .IN2(CRC_OUT_2_22), .Q(n11090) );
  AND2X1 U10930 ( .IN1(n1705), .IN2(n10013), .Q(n11089) );
  INVX0 U10931 ( .INP(n11091), .ZN(n1705) );
  OR2X1 U10932 ( .IN1(n10647), .IN2(n3839), .Q(n11091) );
  OR2X1 U10933 ( .IN1(n11092), .IN2(n11093), .Q(n11087) );
  AND2X1 U10934 ( .IN1(n10070), .IN2(n11094), .Q(n11093) );
  AND2X1 U10935 ( .IN1(n9983), .IN2(n11095), .Q(n11092) );
  OR2X1 U10936 ( .IN1(n11096), .IN2(n11097), .Q(WX9711) );
  OR2X1 U10937 ( .IN1(n11098), .IN2(n11099), .Q(n11097) );
  AND2X1 U10938 ( .IN1(n10039), .IN2(CRC_OUT_2_23), .Q(n11099) );
  AND2X1 U10939 ( .IN1(n1704), .IN2(n10013), .Q(n11098) );
  INVX0 U10940 ( .INP(n11100), .ZN(n1704) );
  OR2X1 U10941 ( .IN1(n10647), .IN2(n3840), .Q(n11100) );
  OR2X1 U10942 ( .IN1(n11101), .IN2(n11102), .Q(n11096) );
  AND2X1 U10943 ( .IN1(n11103), .IN2(n10063), .Q(n11102) );
  AND2X1 U10944 ( .IN1(n9983), .IN2(n11104), .Q(n11101) );
  OR2X1 U10945 ( .IN1(n11105), .IN2(n11106), .Q(WX9709) );
  OR2X1 U10946 ( .IN1(n11107), .IN2(n11108), .Q(n11106) );
  AND2X1 U10947 ( .IN1(n10039), .IN2(CRC_OUT_2_24), .Q(n11108) );
  AND2X1 U10948 ( .IN1(n1703), .IN2(n10013), .Q(n11107) );
  INVX0 U10949 ( .INP(n11109), .ZN(n1703) );
  OR2X1 U10950 ( .IN1(n10647), .IN2(n3841), .Q(n11109) );
  OR2X1 U10951 ( .IN1(n11110), .IN2(n11111), .Q(n11105) );
  AND2X1 U10952 ( .IN1(n10070), .IN2(n11112), .Q(n11111) );
  AND2X1 U10953 ( .IN1(n9983), .IN2(n11113), .Q(n11110) );
  OR2X1 U10954 ( .IN1(n11114), .IN2(n11115), .Q(WX9707) );
  OR2X1 U10955 ( .IN1(n11116), .IN2(n11117), .Q(n11115) );
  AND2X1 U10956 ( .IN1(n10039), .IN2(CRC_OUT_2_25), .Q(n11117) );
  AND2X1 U10957 ( .IN1(n1702), .IN2(n10013), .Q(n11116) );
  INVX0 U10958 ( .INP(n11118), .ZN(n1702) );
  OR2X1 U10959 ( .IN1(n10647), .IN2(n3842), .Q(n11118) );
  OR2X1 U10960 ( .IN1(n11119), .IN2(n11120), .Q(n11114) );
  AND2X1 U10961 ( .IN1(n11121), .IN2(n10062), .Q(n11120) );
  AND2X1 U10962 ( .IN1(n9983), .IN2(n11122), .Q(n11119) );
  OR2X1 U10963 ( .IN1(n11123), .IN2(n11124), .Q(WX9705) );
  OR2X1 U10964 ( .IN1(n11125), .IN2(n11126), .Q(n11124) );
  AND2X1 U10965 ( .IN1(n10039), .IN2(CRC_OUT_2_26), .Q(n11126) );
  AND2X1 U10966 ( .IN1(n1701), .IN2(n10013), .Q(n11125) );
  INVX0 U10967 ( .INP(n11127), .ZN(n1701) );
  OR2X1 U10968 ( .IN1(n10647), .IN2(n3843), .Q(n11127) );
  OR2X1 U10969 ( .IN1(n11128), .IN2(n11129), .Q(n11123) );
  AND2X1 U10970 ( .IN1(n10070), .IN2(n11130), .Q(n11129) );
  AND2X1 U10971 ( .IN1(n9983), .IN2(n11131), .Q(n11128) );
  OR2X1 U10972 ( .IN1(n11132), .IN2(n11133), .Q(WX9703) );
  OR2X1 U10973 ( .IN1(n11134), .IN2(n11135), .Q(n11133) );
  AND2X1 U10974 ( .IN1(n10039), .IN2(CRC_OUT_2_27), .Q(n11135) );
  AND2X1 U10975 ( .IN1(n1700), .IN2(n10013), .Q(n11134) );
  INVX0 U10976 ( .INP(n11136), .ZN(n1700) );
  OR2X1 U10977 ( .IN1(n10647), .IN2(n3844), .Q(n11136) );
  OR2X1 U10978 ( .IN1(n11137), .IN2(n11138), .Q(n11132) );
  AND2X1 U10979 ( .IN1(n10070), .IN2(n11139), .Q(n11138) );
  AND2X1 U10980 ( .IN1(n9983), .IN2(n11140), .Q(n11137) );
  OR2X1 U10981 ( .IN1(n11141), .IN2(n11142), .Q(WX9701) );
  OR2X1 U10982 ( .IN1(n11143), .IN2(n11144), .Q(n11142) );
  AND2X1 U10983 ( .IN1(n10039), .IN2(CRC_OUT_2_28), .Q(n11144) );
  AND2X1 U10984 ( .IN1(n1699), .IN2(n10013), .Q(n11143) );
  INVX0 U10985 ( .INP(n11145), .ZN(n1699) );
  OR2X1 U10986 ( .IN1(n10647), .IN2(n3845), .Q(n11145) );
  OR2X1 U10987 ( .IN1(n11146), .IN2(n11147), .Q(n11141) );
  AND2X1 U10988 ( .IN1(n10070), .IN2(n11148), .Q(n11147) );
  AND2X1 U10989 ( .IN1(n9983), .IN2(n11149), .Q(n11146) );
  OR2X1 U10990 ( .IN1(n11150), .IN2(n11151), .Q(WX9699) );
  OR2X1 U10991 ( .IN1(n11152), .IN2(n11153), .Q(n11151) );
  AND2X1 U10992 ( .IN1(n10039), .IN2(CRC_OUT_2_29), .Q(n11153) );
  AND2X1 U10993 ( .IN1(n1698), .IN2(n10014), .Q(n11152) );
  INVX0 U10994 ( .INP(n11154), .ZN(n1698) );
  OR2X1 U10995 ( .IN1(n10647), .IN2(n3846), .Q(n11154) );
  OR2X1 U10996 ( .IN1(n11155), .IN2(n11156), .Q(n11150) );
  AND2X1 U10997 ( .IN1(n10070), .IN2(n11157), .Q(n11156) );
  AND2X1 U10998 ( .IN1(n9983), .IN2(n11158), .Q(n11155) );
  OR2X1 U10999 ( .IN1(n11159), .IN2(n11160), .Q(WX9697) );
  OR2X1 U11000 ( .IN1(n11161), .IN2(n11162), .Q(n11160) );
  AND2X1 U11001 ( .IN1(n10039), .IN2(CRC_OUT_2_30), .Q(n11162) );
  AND2X1 U11002 ( .IN1(n1697), .IN2(n10014), .Q(n11161) );
  INVX0 U11003 ( .INP(n11163), .ZN(n1697) );
  OR2X1 U11004 ( .IN1(n10647), .IN2(n3847), .Q(n11163) );
  OR2X1 U11005 ( .IN1(n11164), .IN2(n11165), .Q(n11159) );
  AND2X1 U11006 ( .IN1(n10070), .IN2(n11166), .Q(n11165) );
  AND2X1 U11007 ( .IN1(n9983), .IN2(n11167), .Q(n11164) );
  OR2X1 U11008 ( .IN1(n11168), .IN2(n11169), .Q(WX9695) );
  OR2X1 U11009 ( .IN1(n11170), .IN2(n11171), .Q(n11169) );
  AND2X1 U11010 ( .IN1(n2245), .IN2(WX9536), .Q(n11171) );
  AND2X1 U11011 ( .IN1(n10039), .IN2(CRC_OUT_2_31), .Q(n11170) );
  OR2X1 U11012 ( .IN1(n11172), .IN2(n11173), .Q(n11168) );
  AND2X1 U11013 ( .IN1(n10070), .IN2(n11174), .Q(n11173) );
  AND2X1 U11014 ( .IN1(n11175), .IN2(n9975), .Q(n11172) );
  AND2X1 U11015 ( .IN1(n9850), .IN2(n10570), .Q(WX9597) );
  AND2X1 U11016 ( .IN1(n11176), .IN2(n10570), .Q(WX9084) );
  AND2X1 U11017 ( .IN1(n11177), .IN2(n11178), .Q(n11176) );
  OR2X1 U11018 ( .IN1(DFF_1342_n1), .IN2(WX8595), .Q(n11178) );
  OR2X1 U11019 ( .IN1(n9593), .IN2(CRC_OUT_3_30), .Q(n11177) );
  AND2X1 U11020 ( .IN1(n11179), .IN2(n10570), .Q(WX9082) );
  AND2X1 U11021 ( .IN1(n11180), .IN2(n11181), .Q(n11179) );
  OR2X1 U11022 ( .IN1(DFF_1341_n1), .IN2(WX8597), .Q(n11181) );
  OR2X1 U11023 ( .IN1(n9594), .IN2(CRC_OUT_3_29), .Q(n11180) );
  AND2X1 U11024 ( .IN1(n11182), .IN2(n10570), .Q(WX9080) );
  AND2X1 U11025 ( .IN1(n11183), .IN2(n11184), .Q(n11182) );
  OR2X1 U11026 ( .IN1(DFF_1340_n1), .IN2(WX8599), .Q(n11184) );
  OR2X1 U11027 ( .IN1(n9595), .IN2(CRC_OUT_3_28), .Q(n11183) );
  AND2X1 U11028 ( .IN1(n11185), .IN2(n10570), .Q(WX9078) );
  AND2X1 U11029 ( .IN1(n11186), .IN2(n11187), .Q(n11185) );
  OR2X1 U11030 ( .IN1(DFF_1339_n1), .IN2(WX8601), .Q(n11187) );
  OR2X1 U11031 ( .IN1(n9596), .IN2(CRC_OUT_3_27), .Q(n11186) );
  AND2X1 U11032 ( .IN1(n11188), .IN2(n10570), .Q(WX9076) );
  AND2X1 U11033 ( .IN1(n11189), .IN2(n11190), .Q(n11188) );
  OR2X1 U11034 ( .IN1(DFF_1338_n1), .IN2(WX8603), .Q(n11190) );
  OR2X1 U11035 ( .IN1(n9597), .IN2(CRC_OUT_3_26), .Q(n11189) );
  AND2X1 U11036 ( .IN1(n11191), .IN2(n10569), .Q(WX9074) );
  OR2X1 U11037 ( .IN1(n11192), .IN2(n11193), .Q(n11191) );
  AND2X1 U11038 ( .IN1(DFF_1337_n1), .IN2(n9908), .Q(n11193) );
  AND2X1 U11039 ( .IN1(test_so74), .IN2(CRC_OUT_3_25), .Q(n11192) );
  AND2X1 U11040 ( .IN1(n11194), .IN2(n10569), .Q(WX9072) );
  OR2X1 U11041 ( .IN1(n11195), .IN2(n11196), .Q(n11194) );
  AND2X1 U11042 ( .IN1(n9598), .IN2(n9937), .Q(n11196) );
  AND2X1 U11043 ( .IN1(test_so77), .IN2(WX8607), .Q(n11195) );
  AND2X1 U11044 ( .IN1(n11197), .IN2(n10569), .Q(WX9070) );
  AND2X1 U11045 ( .IN1(n11198), .IN2(n11199), .Q(n11197) );
  OR2X1 U11046 ( .IN1(DFF_1335_n1), .IN2(WX8609), .Q(n11199) );
  OR2X1 U11047 ( .IN1(n9599), .IN2(CRC_OUT_3_23), .Q(n11198) );
  AND2X1 U11048 ( .IN1(n11200), .IN2(n10569), .Q(WX9068) );
  AND2X1 U11049 ( .IN1(n11201), .IN2(n11202), .Q(n11200) );
  OR2X1 U11050 ( .IN1(DFF_1334_n1), .IN2(WX8611), .Q(n11202) );
  OR2X1 U11051 ( .IN1(n9600), .IN2(CRC_OUT_3_22), .Q(n11201) );
  AND2X1 U11052 ( .IN1(n11203), .IN2(n10569), .Q(WX9066) );
  AND2X1 U11053 ( .IN1(n11204), .IN2(n11205), .Q(n11203) );
  OR2X1 U11054 ( .IN1(DFF_1333_n1), .IN2(WX8613), .Q(n11205) );
  OR2X1 U11055 ( .IN1(n9601), .IN2(CRC_OUT_3_21), .Q(n11204) );
  AND2X1 U11056 ( .IN1(n11206), .IN2(n10569), .Q(WX9064) );
  AND2X1 U11057 ( .IN1(n11207), .IN2(n11208), .Q(n11206) );
  OR2X1 U11058 ( .IN1(DFF_1332_n1), .IN2(WX8615), .Q(n11208) );
  OR2X1 U11059 ( .IN1(n9602), .IN2(CRC_OUT_3_20), .Q(n11207) );
  AND2X1 U11060 ( .IN1(n11209), .IN2(n10569), .Q(WX9062) );
  AND2X1 U11061 ( .IN1(n11210), .IN2(n11211), .Q(n11209) );
  OR2X1 U11062 ( .IN1(DFF_1331_n1), .IN2(WX8617), .Q(n11211) );
  OR2X1 U11063 ( .IN1(n9603), .IN2(CRC_OUT_3_19), .Q(n11210) );
  AND2X1 U11064 ( .IN1(n11212), .IN2(n10569), .Q(WX9060) );
  AND2X1 U11065 ( .IN1(n11213), .IN2(n11214), .Q(n11212) );
  OR2X1 U11066 ( .IN1(DFF_1330_n1), .IN2(WX8619), .Q(n11214) );
  OR2X1 U11067 ( .IN1(n9604), .IN2(CRC_OUT_3_18), .Q(n11213) );
  AND2X1 U11068 ( .IN1(n11215), .IN2(n10569), .Q(WX9058) );
  AND2X1 U11069 ( .IN1(n11216), .IN2(n11217), .Q(n11215) );
  OR2X1 U11070 ( .IN1(DFF_1329_n1), .IN2(WX8621), .Q(n11217) );
  OR2X1 U11071 ( .IN1(n9605), .IN2(CRC_OUT_3_17), .Q(n11216) );
  AND2X1 U11072 ( .IN1(n11218), .IN2(n10568), .Q(WX9056) );
  AND2X1 U11073 ( .IN1(n11219), .IN2(n11220), .Q(n11218) );
  OR2X1 U11074 ( .IN1(DFF_1328_n1), .IN2(WX8623), .Q(n11220) );
  OR2X1 U11075 ( .IN1(n9606), .IN2(CRC_OUT_3_16), .Q(n11219) );
  AND2X1 U11076 ( .IN1(n11221), .IN2(n10568), .Q(WX9054) );
  OR2X1 U11077 ( .IN1(n11222), .IN2(n11223), .Q(n11221) );
  AND2X1 U11078 ( .IN1(n11224), .IN2(CRC_OUT_3_15), .Q(n11223) );
  AND2X1 U11079 ( .IN1(DFF_1327_n1), .IN2(n11225), .Q(n11222) );
  INVX0 U11080 ( .INP(n11224), .ZN(n11225) );
  OR2X1 U11081 ( .IN1(n11226), .IN2(n11227), .Q(n11224) );
  AND2X1 U11082 ( .IN1(DFF_1343_n1), .IN2(WX8625), .Q(n11227) );
  AND2X1 U11083 ( .IN1(n9518), .IN2(CRC_OUT_3_31), .Q(n11226) );
  AND2X1 U11084 ( .IN1(n11228), .IN2(n10568), .Q(WX9052) );
  AND2X1 U11085 ( .IN1(n11229), .IN2(n11230), .Q(n11228) );
  OR2X1 U11086 ( .IN1(DFF_1326_n1), .IN2(WX8627), .Q(n11230) );
  OR2X1 U11087 ( .IN1(n9607), .IN2(CRC_OUT_3_14), .Q(n11229) );
  AND2X1 U11088 ( .IN1(n11231), .IN2(n10568), .Q(WX9050) );
  AND2X1 U11089 ( .IN1(n11232), .IN2(n11233), .Q(n11231) );
  OR2X1 U11090 ( .IN1(DFF_1325_n1), .IN2(WX8629), .Q(n11233) );
  OR2X1 U11091 ( .IN1(n9608), .IN2(CRC_OUT_3_13), .Q(n11232) );
  AND2X1 U11092 ( .IN1(n11234), .IN2(n10568), .Q(WX9048) );
  AND2X1 U11093 ( .IN1(n11235), .IN2(n11236), .Q(n11234) );
  OR2X1 U11094 ( .IN1(DFF_1324_n1), .IN2(WX8631), .Q(n11236) );
  OR2X1 U11095 ( .IN1(n9609), .IN2(CRC_OUT_3_12), .Q(n11235) );
  AND2X1 U11096 ( .IN1(n11237), .IN2(n10568), .Q(WX9046) );
  AND2X1 U11097 ( .IN1(n11238), .IN2(n11239), .Q(n11237) );
  OR2X1 U11098 ( .IN1(DFF_1323_n1), .IN2(WX8633), .Q(n11239) );
  OR2X1 U11099 ( .IN1(n9610), .IN2(CRC_OUT_3_11), .Q(n11238) );
  AND2X1 U11100 ( .IN1(n11240), .IN2(n10568), .Q(WX9044) );
  OR2X1 U11101 ( .IN1(n11241), .IN2(n11242), .Q(n11240) );
  AND2X1 U11102 ( .IN1(n11243), .IN2(CRC_OUT_3_10), .Q(n11242) );
  AND2X1 U11103 ( .IN1(DFF_1322_n1), .IN2(n11244), .Q(n11241) );
  INVX0 U11104 ( .INP(n11243), .ZN(n11244) );
  OR2X1 U11105 ( .IN1(n11245), .IN2(n11246), .Q(n11243) );
  AND2X1 U11106 ( .IN1(DFF_1343_n1), .IN2(WX8635), .Q(n11246) );
  AND2X1 U11107 ( .IN1(n9519), .IN2(CRC_OUT_3_31), .Q(n11245) );
  AND2X1 U11108 ( .IN1(n11247), .IN2(n10568), .Q(WX9042) );
  AND2X1 U11109 ( .IN1(n11248), .IN2(n11249), .Q(n11247) );
  OR2X1 U11110 ( .IN1(DFF_1321_n1), .IN2(WX8637), .Q(n11249) );
  OR2X1 U11111 ( .IN1(n9611), .IN2(CRC_OUT_3_9), .Q(n11248) );
  AND2X1 U11112 ( .IN1(n11250), .IN2(n10568), .Q(WX9040) );
  OR2X1 U11113 ( .IN1(n11251), .IN2(n11252), .Q(n11250) );
  AND2X1 U11114 ( .IN1(DFF_1320_n1), .IN2(n9903), .Q(n11252) );
  AND2X1 U11115 ( .IN1(test_so75), .IN2(CRC_OUT_3_8), .Q(n11251) );
  AND2X1 U11116 ( .IN1(n11253), .IN2(n10567), .Q(WX9038) );
  OR2X1 U11117 ( .IN1(n11254), .IN2(n11255), .Q(n11253) );
  AND2X1 U11118 ( .IN1(n9612), .IN2(n9938), .Q(n11255) );
  AND2X1 U11119 ( .IN1(test_so76), .IN2(WX8641), .Q(n11254) );
  AND2X1 U11120 ( .IN1(n11256), .IN2(n10567), .Q(WX9036) );
  AND2X1 U11121 ( .IN1(n11257), .IN2(n11258), .Q(n11256) );
  OR2X1 U11122 ( .IN1(DFF_1318_n1), .IN2(WX8643), .Q(n11258) );
  OR2X1 U11123 ( .IN1(n9613), .IN2(CRC_OUT_3_6), .Q(n11257) );
  AND2X1 U11124 ( .IN1(n11259), .IN2(n10567), .Q(WX9034) );
  AND2X1 U11125 ( .IN1(n11260), .IN2(n11261), .Q(n11259) );
  OR2X1 U11126 ( .IN1(DFF_1317_n1), .IN2(WX8645), .Q(n11261) );
  OR2X1 U11127 ( .IN1(n9614), .IN2(CRC_OUT_3_5), .Q(n11260) );
  AND2X1 U11128 ( .IN1(n11262), .IN2(n10567), .Q(WX9032) );
  AND2X1 U11129 ( .IN1(n11263), .IN2(n11264), .Q(n11262) );
  OR2X1 U11130 ( .IN1(DFF_1316_n1), .IN2(WX8647), .Q(n11264) );
  OR2X1 U11131 ( .IN1(n9615), .IN2(CRC_OUT_3_4), .Q(n11263) );
  AND2X1 U11132 ( .IN1(n11265), .IN2(n10567), .Q(WX9030) );
  OR2X1 U11133 ( .IN1(n11266), .IN2(n11267), .Q(n11265) );
  AND2X1 U11134 ( .IN1(n11268), .IN2(CRC_OUT_3_3), .Q(n11267) );
  AND2X1 U11135 ( .IN1(DFF_1315_n1), .IN2(n11269), .Q(n11266) );
  INVX0 U11136 ( .INP(n11268), .ZN(n11269) );
  OR2X1 U11137 ( .IN1(n11270), .IN2(n11271), .Q(n11268) );
  AND2X1 U11138 ( .IN1(DFF_1343_n1), .IN2(WX8649), .Q(n11271) );
  AND2X1 U11139 ( .IN1(n9520), .IN2(CRC_OUT_3_31), .Q(n11270) );
  AND2X1 U11140 ( .IN1(n11272), .IN2(n10567), .Q(WX9028) );
  AND2X1 U11141 ( .IN1(n11273), .IN2(n11274), .Q(n11272) );
  OR2X1 U11142 ( .IN1(DFF_1314_n1), .IN2(WX8651), .Q(n11274) );
  OR2X1 U11143 ( .IN1(n9616), .IN2(CRC_OUT_3_2), .Q(n11273) );
  AND2X1 U11144 ( .IN1(n11275), .IN2(n10567), .Q(WX9026) );
  AND2X1 U11145 ( .IN1(n11276), .IN2(n11277), .Q(n11275) );
  OR2X1 U11146 ( .IN1(DFF_1313_n1), .IN2(WX8653), .Q(n11277) );
  OR2X1 U11147 ( .IN1(n9617), .IN2(CRC_OUT_3_1), .Q(n11276) );
  AND2X1 U11148 ( .IN1(n11278), .IN2(n10567), .Q(WX9024) );
  AND2X1 U11149 ( .IN1(n11279), .IN2(n11280), .Q(n11278) );
  OR2X1 U11150 ( .IN1(DFF_1312_n1), .IN2(WX8655), .Q(n11280) );
  OR2X1 U11151 ( .IN1(n9618), .IN2(CRC_OUT_3_0), .Q(n11279) );
  AND2X1 U11152 ( .IN1(n11281), .IN2(n10567), .Q(WX9022) );
  AND2X1 U11153 ( .IN1(n11282), .IN2(n11283), .Q(n11281) );
  OR2X1 U11154 ( .IN1(DFF_1343_n1), .IN2(WX8657), .Q(n11283) );
  OR2X1 U11155 ( .IN1(n9535), .IN2(CRC_OUT_3_31), .Q(n11282) );
  AND2X1 U11156 ( .IN1(n10597), .IN2(n8363), .Q(WX8496) );
  AND2X1 U11157 ( .IN1(n10598), .IN2(n8364), .Q(WX8494) );
  AND2X1 U11158 ( .IN1(n10598), .IN2(n8365), .Q(WX8492) );
  AND2X1 U11159 ( .IN1(n10598), .IN2(n8366), .Q(WX8490) );
  AND2X1 U11160 ( .IN1(n10598), .IN2(n8367), .Q(WX8488) );
  AND2X1 U11161 ( .IN1(n10598), .IN2(n8368), .Q(WX8486) );
  AND2X1 U11162 ( .IN1(n10598), .IN2(n8369), .Q(WX8484) );
  AND2X1 U11163 ( .IN1(n10598), .IN2(n8370), .Q(WX8482) );
  AND2X1 U11164 ( .IN1(n10598), .IN2(n8371), .Q(WX8480) );
  AND2X1 U11165 ( .IN1(n10598), .IN2(n8372), .Q(WX8478) );
  AND2X1 U11166 ( .IN1(n10599), .IN2(n8373), .Q(WX8476) );
  AND2X1 U11167 ( .IN1(n10599), .IN2(n8374), .Q(WX8474) );
  AND2X1 U11168 ( .IN1(n10599), .IN2(n8375), .Q(WX8472) );
  AND2X1 U11169 ( .IN1(n10599), .IN2(n8376), .Q(WX8470) );
  AND2X1 U11170 ( .IN1(n10599), .IN2(n8377), .Q(WX8468) );
  AND2X1 U11171 ( .IN1(n10599), .IN2(n8378), .Q(WX8466) );
  OR2X1 U11172 ( .IN1(n11284), .IN2(n11285), .Q(WX8464) );
  OR2X1 U11173 ( .IN1(n11286), .IN2(n11287), .Q(n11285) );
  AND2X1 U11174 ( .IN1(n10039), .IN2(CRC_OUT_3_0), .Q(n11287) );
  AND2X1 U11175 ( .IN1(n1485), .IN2(n10014), .Q(n11286) );
  INVX0 U11176 ( .INP(n11288), .ZN(n1485) );
  OR2X1 U11177 ( .IN1(n10647), .IN2(n3848), .Q(n11288) );
  OR2X1 U11178 ( .IN1(n11289), .IN2(n11290), .Q(n11284) );
  AND2X1 U11179 ( .IN1(n9982), .IN2(n11291), .Q(n11290) );
  AND2X1 U11180 ( .IN1(n10070), .IN2(n10897), .Q(n11289) );
  OR2X1 U11181 ( .IN1(n11292), .IN2(n11293), .Q(n10897) );
  INVX0 U11182 ( .INP(n11294), .ZN(n11293) );
  OR2X1 U11183 ( .IN1(n11295), .IN2(n11296), .Q(n11294) );
  AND2X1 U11184 ( .IN1(n11296), .IN2(n11295), .Q(n11292) );
  AND2X1 U11185 ( .IN1(n11297), .IN2(n11298), .Q(n11295) );
  OR2X1 U11186 ( .IN1(WX9822), .IN2(n9300), .Q(n11298) );
  OR2X1 U11187 ( .IN1(WX9758), .IN2(n3563), .Q(n11297) );
  OR2X1 U11188 ( .IN1(n11299), .IN2(n11300), .Q(n11296) );
  AND2X1 U11189 ( .IN1(n9301), .IN2(WX9950), .Q(n11300) );
  AND2X1 U11190 ( .IN1(n9534), .IN2(WX9886), .Q(n11299) );
  OR2X1 U11191 ( .IN1(n11301), .IN2(n11302), .Q(WX8462) );
  OR2X1 U11192 ( .IN1(n11303), .IN2(n11304), .Q(n11302) );
  AND2X1 U11193 ( .IN1(n10039), .IN2(CRC_OUT_3_1), .Q(n11304) );
  AND2X1 U11194 ( .IN1(n1484), .IN2(n10014), .Q(n11303) );
  INVX0 U11195 ( .INP(n11305), .ZN(n1484) );
  OR2X1 U11196 ( .IN1(n10646), .IN2(n3849), .Q(n11305) );
  OR2X1 U11197 ( .IN1(n11306), .IN2(n11307), .Q(n11301) );
  AND2X1 U11198 ( .IN1(n9982), .IN2(n11308), .Q(n11307) );
  AND2X1 U11199 ( .IN1(n10906), .IN2(n10061), .Q(n11306) );
  AND2X1 U11200 ( .IN1(n11309), .IN2(n11310), .Q(n10906) );
  INVX0 U11201 ( .INP(n11311), .ZN(n11310) );
  AND2X1 U11202 ( .IN1(n11312), .IN2(n11313), .Q(n11311) );
  OR2X1 U11203 ( .IN1(n11313), .IN2(n11312), .Q(n11309) );
  OR2X1 U11204 ( .IN1(n11314), .IN2(n11315), .Q(n11312) );
  AND2X1 U11205 ( .IN1(n9302), .IN2(WX9884), .Q(n11315) );
  INVX0 U11206 ( .INP(n11316), .ZN(n11314) );
  OR2X1 U11207 ( .IN1(WX9884), .IN2(n9302), .Q(n11316) );
  AND2X1 U11208 ( .IN1(n11317), .IN2(n11318), .Q(n11313) );
  OR2X1 U11209 ( .IN1(WX9948), .IN2(test_so83), .Q(n11318) );
  OR2X1 U11210 ( .IN1(n9915), .IN2(n9592), .Q(n11317) );
  OR2X1 U11211 ( .IN1(n11319), .IN2(n11320), .Q(WX8460) );
  OR2X1 U11212 ( .IN1(n11321), .IN2(n11322), .Q(n11320) );
  AND2X1 U11213 ( .IN1(n10039), .IN2(CRC_OUT_3_2), .Q(n11322) );
  AND2X1 U11214 ( .IN1(n1483), .IN2(n10017), .Q(n11321) );
  INVX0 U11215 ( .INP(n11323), .ZN(n1483) );
  OR2X1 U11216 ( .IN1(n10646), .IN2(n3850), .Q(n11323) );
  OR2X1 U11217 ( .IN1(n11324), .IN2(n11325), .Q(n11319) );
  AND2X1 U11218 ( .IN1(n9982), .IN2(n11326), .Q(n11325) );
  AND2X1 U11219 ( .IN1(n10070), .IN2(n10915), .Q(n11324) );
  OR2X1 U11220 ( .IN1(n11327), .IN2(n11328), .Q(n10915) );
  INVX0 U11221 ( .INP(n11329), .ZN(n11328) );
  OR2X1 U11222 ( .IN1(n11330), .IN2(n11331), .Q(n11329) );
  AND2X1 U11223 ( .IN1(n11331), .IN2(n11330), .Q(n11327) );
  AND2X1 U11224 ( .IN1(n11332), .IN2(n11333), .Q(n11330) );
  OR2X1 U11225 ( .IN1(WX9818), .IN2(n9304), .Q(n11333) );
  OR2X1 U11226 ( .IN1(WX9754), .IN2(n3567), .Q(n11332) );
  OR2X1 U11227 ( .IN1(n11334), .IN2(n11335), .Q(n11331) );
  AND2X1 U11228 ( .IN1(n9305), .IN2(WX9946), .Q(n11335) );
  AND2X1 U11229 ( .IN1(n9591), .IN2(WX9882), .Q(n11334) );
  OR2X1 U11230 ( .IN1(n11336), .IN2(n11337), .Q(WX8458) );
  OR2X1 U11231 ( .IN1(n11338), .IN2(n11339), .Q(n11337) );
  AND2X1 U11232 ( .IN1(n10040), .IN2(CRC_OUT_3_3), .Q(n11339) );
  AND2X1 U11233 ( .IN1(n1482), .IN2(n10014), .Q(n11338) );
  INVX0 U11234 ( .INP(n11340), .ZN(n1482) );
  OR2X1 U11235 ( .IN1(n10646), .IN2(n3851), .Q(n11340) );
  OR2X1 U11236 ( .IN1(n11341), .IN2(n11342), .Q(n11336) );
  AND2X1 U11237 ( .IN1(n9982), .IN2(n11343), .Q(n11342) );
  AND2X1 U11238 ( .IN1(n10924), .IN2(n10060), .Q(n11341) );
  AND2X1 U11239 ( .IN1(n11344), .IN2(n11345), .Q(n10924) );
  INVX0 U11240 ( .INP(n11346), .ZN(n11345) );
  AND2X1 U11241 ( .IN1(n11347), .IN2(n11348), .Q(n11346) );
  OR2X1 U11242 ( .IN1(n11348), .IN2(n11347), .Q(n11344) );
  OR2X1 U11243 ( .IN1(n11349), .IN2(n11350), .Q(n11347) );
  AND2X1 U11244 ( .IN1(n3569), .IN2(WX9880), .Q(n11350) );
  INVX0 U11245 ( .INP(n11351), .ZN(n11349) );
  OR2X1 U11246 ( .IN1(WX9880), .IN2(n3569), .Q(n11351) );
  AND2X1 U11247 ( .IN1(n11352), .IN2(n11353), .Q(n11348) );
  OR2X1 U11248 ( .IN1(WX9944), .IN2(test_so81), .Q(n11353) );
  OR2X1 U11249 ( .IN1(n9916), .IN2(n9590), .Q(n11352) );
  OR2X1 U11250 ( .IN1(n11354), .IN2(n11355), .Q(WX8456) );
  OR2X1 U11251 ( .IN1(n11356), .IN2(n11357), .Q(n11355) );
  AND2X1 U11252 ( .IN1(n10040), .IN2(CRC_OUT_3_4), .Q(n11357) );
  AND2X1 U11253 ( .IN1(n1481), .IN2(n10014), .Q(n11356) );
  INVX0 U11254 ( .INP(n11358), .ZN(n1481) );
  OR2X1 U11255 ( .IN1(n10646), .IN2(n3852), .Q(n11358) );
  OR2X1 U11256 ( .IN1(n11359), .IN2(n11360), .Q(n11354) );
  AND2X1 U11257 ( .IN1(n9982), .IN2(n11361), .Q(n11360) );
  AND2X1 U11258 ( .IN1(n10071), .IN2(n10933), .Q(n11359) );
  OR2X1 U11259 ( .IN1(n11362), .IN2(n11363), .Q(n10933) );
  INVX0 U11260 ( .INP(n11364), .ZN(n11363) );
  OR2X1 U11261 ( .IN1(n11365), .IN2(n11366), .Q(n11364) );
  AND2X1 U11262 ( .IN1(n11366), .IN2(n11365), .Q(n11362) );
  AND2X1 U11263 ( .IN1(n11367), .IN2(n11368), .Q(n11365) );
  OR2X1 U11264 ( .IN1(WX9814), .IN2(n9307), .Q(n11368) );
  OR2X1 U11265 ( .IN1(WX9750), .IN2(n3571), .Q(n11367) );
  OR2X1 U11266 ( .IN1(n11369), .IN2(n11370), .Q(n11366) );
  AND2X1 U11267 ( .IN1(n9308), .IN2(WX9942), .Q(n11370) );
  AND2X1 U11268 ( .IN1(n9517), .IN2(WX9878), .Q(n11369) );
  OR2X1 U11269 ( .IN1(n11371), .IN2(n11372), .Q(WX8454) );
  OR2X1 U11270 ( .IN1(n11373), .IN2(n11374), .Q(n11372) );
  AND2X1 U11271 ( .IN1(n10040), .IN2(CRC_OUT_3_5), .Q(n11374) );
  AND2X1 U11272 ( .IN1(n1480), .IN2(n10014), .Q(n11373) );
  INVX0 U11273 ( .INP(n11375), .ZN(n1480) );
  OR2X1 U11274 ( .IN1(n10646), .IN2(n3853), .Q(n11375) );
  OR2X1 U11275 ( .IN1(n11376), .IN2(n11377), .Q(n11371) );
  AND2X1 U11276 ( .IN1(n9982), .IN2(n11378), .Q(n11377) );
  AND2X1 U11277 ( .IN1(n10071), .IN2(n10942), .Q(n11376) );
  OR2X1 U11278 ( .IN1(n11379), .IN2(n11380), .Q(n10942) );
  INVX0 U11279 ( .INP(n11381), .ZN(n11380) );
  OR2X1 U11280 ( .IN1(n11382), .IN2(n11383), .Q(n11381) );
  AND2X1 U11281 ( .IN1(n11383), .IN2(n11382), .Q(n11379) );
  AND2X1 U11282 ( .IN1(n11384), .IN2(n11385), .Q(n11382) );
  OR2X1 U11283 ( .IN1(WX9812), .IN2(n9309), .Q(n11385) );
  OR2X1 U11284 ( .IN1(WX9748), .IN2(n3573), .Q(n11384) );
  OR2X1 U11285 ( .IN1(n11386), .IN2(n11387), .Q(n11383) );
  AND2X1 U11286 ( .IN1(n9310), .IN2(WX9940), .Q(n11387) );
  AND2X1 U11287 ( .IN1(n9589), .IN2(WX9876), .Q(n11386) );
  OR2X1 U11288 ( .IN1(n11388), .IN2(n11389), .Q(WX8452) );
  OR2X1 U11289 ( .IN1(n11390), .IN2(n11391), .Q(n11389) );
  AND2X1 U11290 ( .IN1(n10040), .IN2(CRC_OUT_3_6), .Q(n11391) );
  AND2X1 U11291 ( .IN1(n1479), .IN2(n10014), .Q(n11390) );
  INVX0 U11292 ( .INP(n11392), .ZN(n1479) );
  OR2X1 U11293 ( .IN1(n10646), .IN2(n3854), .Q(n11392) );
  OR2X1 U11294 ( .IN1(n11393), .IN2(n11394), .Q(n11388) );
  AND2X1 U11295 ( .IN1(n9982), .IN2(n11395), .Q(n11394) );
  AND2X1 U11296 ( .IN1(n10071), .IN2(n10951), .Q(n11393) );
  OR2X1 U11297 ( .IN1(n11396), .IN2(n11397), .Q(n10951) );
  INVX0 U11298 ( .INP(n11398), .ZN(n11397) );
  OR2X1 U11299 ( .IN1(n11399), .IN2(n11400), .Q(n11398) );
  AND2X1 U11300 ( .IN1(n11400), .IN2(n11399), .Q(n11396) );
  AND2X1 U11301 ( .IN1(n11401), .IN2(n11402), .Q(n11399) );
  OR2X1 U11302 ( .IN1(WX9810), .IN2(n9311), .Q(n11402) );
  OR2X1 U11303 ( .IN1(WX9746), .IN2(n3575), .Q(n11401) );
  OR2X1 U11304 ( .IN1(n11403), .IN2(n11404), .Q(n11400) );
  AND2X1 U11305 ( .IN1(n9312), .IN2(WX9938), .Q(n11404) );
  AND2X1 U11306 ( .IN1(n9588), .IN2(WX9874), .Q(n11403) );
  OR2X1 U11307 ( .IN1(n11405), .IN2(n11406), .Q(WX8450) );
  OR2X1 U11308 ( .IN1(n11407), .IN2(n11408), .Q(n11406) );
  AND2X1 U11309 ( .IN1(test_so76), .IN2(n10027), .Q(n11408) );
  AND2X1 U11310 ( .IN1(n1478), .IN2(n10014), .Q(n11407) );
  INVX0 U11311 ( .INP(n11409), .ZN(n1478) );
  OR2X1 U11312 ( .IN1(n10646), .IN2(n3855), .Q(n11409) );
  OR2X1 U11313 ( .IN1(n11410), .IN2(n11411), .Q(n11405) );
  AND2X1 U11314 ( .IN1(n9982), .IN2(n11412), .Q(n11411) );
  AND2X1 U11315 ( .IN1(n10071), .IN2(n10960), .Q(n11410) );
  OR2X1 U11316 ( .IN1(n11413), .IN2(n11414), .Q(n10960) );
  INVX0 U11317 ( .INP(n11415), .ZN(n11414) );
  OR2X1 U11318 ( .IN1(n11416), .IN2(n11417), .Q(n11415) );
  AND2X1 U11319 ( .IN1(n11417), .IN2(n11416), .Q(n11413) );
  AND2X1 U11320 ( .IN1(n11418), .IN2(n11419), .Q(n11416) );
  OR2X1 U11321 ( .IN1(WX9808), .IN2(n9313), .Q(n11419) );
  OR2X1 U11322 ( .IN1(WX9744), .IN2(n3577), .Q(n11418) );
  OR2X1 U11323 ( .IN1(n11420), .IN2(n11421), .Q(n11417) );
  AND2X1 U11324 ( .IN1(n9314), .IN2(WX9936), .Q(n11421) );
  AND2X1 U11325 ( .IN1(n9587), .IN2(WX9872), .Q(n11420) );
  OR2X1 U11326 ( .IN1(n11422), .IN2(n11423), .Q(WX8448) );
  OR2X1 U11327 ( .IN1(n11424), .IN2(n11425), .Q(n11423) );
  AND2X1 U11328 ( .IN1(n10040), .IN2(CRC_OUT_3_8), .Q(n11425) );
  AND2X1 U11329 ( .IN1(n1477), .IN2(n10014), .Q(n11424) );
  INVX0 U11330 ( .INP(n11426), .ZN(n1477) );
  OR2X1 U11331 ( .IN1(n10646), .IN2(n3856), .Q(n11426) );
  OR2X1 U11332 ( .IN1(n11427), .IN2(n11428), .Q(n11422) );
  AND2X1 U11333 ( .IN1(n9982), .IN2(n11429), .Q(n11428) );
  AND2X1 U11334 ( .IN1(n10071), .IN2(n10969), .Q(n11427) );
  OR2X1 U11335 ( .IN1(n11430), .IN2(n11431), .Q(n10969) );
  INVX0 U11336 ( .INP(n11432), .ZN(n11431) );
  OR2X1 U11337 ( .IN1(n11433), .IN2(n11434), .Q(n11432) );
  AND2X1 U11338 ( .IN1(n11434), .IN2(n11433), .Q(n11430) );
  AND2X1 U11339 ( .IN1(n11435), .IN2(n11436), .Q(n11433) );
  OR2X1 U11340 ( .IN1(WX9806), .IN2(n9315), .Q(n11436) );
  OR2X1 U11341 ( .IN1(WX9742), .IN2(n3579), .Q(n11435) );
  OR2X1 U11342 ( .IN1(n11437), .IN2(n11438), .Q(n11434) );
  AND2X1 U11343 ( .IN1(n9316), .IN2(WX9934), .Q(n11438) );
  AND2X1 U11344 ( .IN1(n9586), .IN2(WX9870), .Q(n11437) );
  OR2X1 U11345 ( .IN1(n11439), .IN2(n11440), .Q(WX8446) );
  OR2X1 U11346 ( .IN1(n11441), .IN2(n11442), .Q(n11440) );
  AND2X1 U11347 ( .IN1(n10040), .IN2(CRC_OUT_3_9), .Q(n11442) );
  AND2X1 U11348 ( .IN1(n1476), .IN2(n10014), .Q(n11441) );
  INVX0 U11349 ( .INP(n11443), .ZN(n1476) );
  OR2X1 U11350 ( .IN1(n10646), .IN2(n3857), .Q(n11443) );
  OR2X1 U11351 ( .IN1(n11444), .IN2(n11445), .Q(n11439) );
  AND2X1 U11352 ( .IN1(n11446), .IN2(n9976), .Q(n11445) );
  AND2X1 U11353 ( .IN1(n10071), .IN2(n10978), .Q(n11444) );
  OR2X1 U11354 ( .IN1(n11447), .IN2(n11448), .Q(n10978) );
  INVX0 U11355 ( .INP(n11449), .ZN(n11448) );
  OR2X1 U11356 ( .IN1(n11450), .IN2(n11451), .Q(n11449) );
  AND2X1 U11357 ( .IN1(n11451), .IN2(n11450), .Q(n11447) );
  AND2X1 U11358 ( .IN1(n11452), .IN2(n11453), .Q(n11450) );
  OR2X1 U11359 ( .IN1(WX9804), .IN2(n9317), .Q(n11453) );
  OR2X1 U11360 ( .IN1(WX9740), .IN2(n3581), .Q(n11452) );
  OR2X1 U11361 ( .IN1(n11454), .IN2(n11455), .Q(n11451) );
  AND2X1 U11362 ( .IN1(n9318), .IN2(WX9932), .Q(n11455) );
  AND2X1 U11363 ( .IN1(n9585), .IN2(WX9868), .Q(n11454) );
  OR2X1 U11364 ( .IN1(n11456), .IN2(n11457), .Q(WX8444) );
  OR2X1 U11365 ( .IN1(n11458), .IN2(n11459), .Q(n11457) );
  AND2X1 U11366 ( .IN1(n10040), .IN2(CRC_OUT_3_10), .Q(n11459) );
  AND2X1 U11367 ( .IN1(n1475), .IN2(n10014), .Q(n11458) );
  INVX0 U11368 ( .INP(n11460), .ZN(n1475) );
  OR2X1 U11369 ( .IN1(n10646), .IN2(n3858), .Q(n11460) );
  OR2X1 U11370 ( .IN1(n11461), .IN2(n11462), .Q(n11456) );
  AND2X1 U11371 ( .IN1(n9982), .IN2(n11463), .Q(n11462) );
  AND2X1 U11372 ( .IN1(n10071), .IN2(n10987), .Q(n11461) );
  OR2X1 U11373 ( .IN1(n11464), .IN2(n11465), .Q(n10987) );
  INVX0 U11374 ( .INP(n11466), .ZN(n11465) );
  OR2X1 U11375 ( .IN1(n11467), .IN2(n11468), .Q(n11466) );
  AND2X1 U11376 ( .IN1(n11468), .IN2(n11467), .Q(n11464) );
  AND2X1 U11377 ( .IN1(n11469), .IN2(n11470), .Q(n11467) );
  OR2X1 U11378 ( .IN1(WX9802), .IN2(n9319), .Q(n11470) );
  OR2X1 U11379 ( .IN1(WX9738), .IN2(n3583), .Q(n11469) );
  OR2X1 U11380 ( .IN1(n11471), .IN2(n11472), .Q(n11468) );
  AND2X1 U11381 ( .IN1(n9320), .IN2(WX9930), .Q(n11472) );
  AND2X1 U11382 ( .IN1(n9584), .IN2(WX9866), .Q(n11471) );
  OR2X1 U11383 ( .IN1(n11473), .IN2(n11474), .Q(WX8442) );
  OR2X1 U11384 ( .IN1(n11475), .IN2(n11476), .Q(n11474) );
  AND2X1 U11385 ( .IN1(n10040), .IN2(CRC_OUT_3_11), .Q(n11476) );
  AND2X1 U11386 ( .IN1(n1474), .IN2(n10015), .Q(n11475) );
  INVX0 U11387 ( .INP(n11477), .ZN(n1474) );
  OR2X1 U11388 ( .IN1(n10646), .IN2(n3859), .Q(n11477) );
  OR2X1 U11389 ( .IN1(n11478), .IN2(n11479), .Q(n11473) );
  AND2X1 U11390 ( .IN1(n11480), .IN2(n9976), .Q(n11479) );
  AND2X1 U11391 ( .IN1(n10071), .IN2(n10996), .Q(n11478) );
  OR2X1 U11392 ( .IN1(n11481), .IN2(n11482), .Q(n10996) );
  INVX0 U11393 ( .INP(n11483), .ZN(n11482) );
  OR2X1 U11394 ( .IN1(n11484), .IN2(n11485), .Q(n11483) );
  AND2X1 U11395 ( .IN1(n11485), .IN2(n11484), .Q(n11481) );
  AND2X1 U11396 ( .IN1(n11486), .IN2(n11487), .Q(n11484) );
  OR2X1 U11397 ( .IN1(WX9800), .IN2(n9321), .Q(n11487) );
  OR2X1 U11398 ( .IN1(WX9736), .IN2(n3585), .Q(n11486) );
  OR2X1 U11399 ( .IN1(n11488), .IN2(n11489), .Q(n11485) );
  AND2X1 U11400 ( .IN1(n9322), .IN2(WX9928), .Q(n11489) );
  AND2X1 U11401 ( .IN1(n9516), .IN2(WX9864), .Q(n11488) );
  OR2X1 U11402 ( .IN1(n11490), .IN2(n11491), .Q(WX8440) );
  OR2X1 U11403 ( .IN1(n11492), .IN2(n11493), .Q(n11491) );
  AND2X1 U11404 ( .IN1(n10040), .IN2(CRC_OUT_3_12), .Q(n11493) );
  AND2X1 U11405 ( .IN1(n1473), .IN2(n10015), .Q(n11492) );
  INVX0 U11406 ( .INP(n11494), .ZN(n1473) );
  OR2X1 U11407 ( .IN1(n10646), .IN2(n3860), .Q(n11494) );
  OR2X1 U11408 ( .IN1(n11495), .IN2(n11496), .Q(n11490) );
  AND2X1 U11409 ( .IN1(n9982), .IN2(n11497), .Q(n11496) );
  AND2X1 U11410 ( .IN1(n10071), .IN2(n11005), .Q(n11495) );
  OR2X1 U11411 ( .IN1(n11498), .IN2(n11499), .Q(n11005) );
  INVX0 U11412 ( .INP(n11500), .ZN(n11499) );
  OR2X1 U11413 ( .IN1(n11501), .IN2(n11502), .Q(n11500) );
  AND2X1 U11414 ( .IN1(n11502), .IN2(n11501), .Q(n11498) );
  AND2X1 U11415 ( .IN1(n11503), .IN2(n11504), .Q(n11501) );
  OR2X1 U11416 ( .IN1(WX9798), .IN2(n9323), .Q(n11504) );
  OR2X1 U11417 ( .IN1(WX9734), .IN2(n3587), .Q(n11503) );
  OR2X1 U11418 ( .IN1(n11505), .IN2(n11506), .Q(n11502) );
  AND2X1 U11419 ( .IN1(n9324), .IN2(WX9926), .Q(n11506) );
  AND2X1 U11420 ( .IN1(n9583), .IN2(WX9862), .Q(n11505) );
  OR2X1 U11421 ( .IN1(n11507), .IN2(n11508), .Q(WX8438) );
  OR2X1 U11422 ( .IN1(n11509), .IN2(n11510), .Q(n11508) );
  AND2X1 U11423 ( .IN1(n10040), .IN2(CRC_OUT_3_13), .Q(n11510) );
  AND2X1 U11424 ( .IN1(n1472), .IN2(n10015), .Q(n11509) );
  INVX0 U11425 ( .INP(n11511), .ZN(n1472) );
  OR2X1 U11426 ( .IN1(n10645), .IN2(n3861), .Q(n11511) );
  OR2X1 U11427 ( .IN1(n11512), .IN2(n11513), .Q(n11507) );
  AND2X1 U11428 ( .IN1(n11514), .IN2(n9976), .Q(n11513) );
  AND2X1 U11429 ( .IN1(n10071), .IN2(n11014), .Q(n11512) );
  OR2X1 U11430 ( .IN1(n11515), .IN2(n11516), .Q(n11014) );
  INVX0 U11431 ( .INP(n11517), .ZN(n11516) );
  OR2X1 U11432 ( .IN1(n11518), .IN2(n11519), .Q(n11517) );
  AND2X1 U11433 ( .IN1(n11519), .IN2(n11518), .Q(n11515) );
  AND2X1 U11434 ( .IN1(n11520), .IN2(n11521), .Q(n11518) );
  OR2X1 U11435 ( .IN1(WX9796), .IN2(n9325), .Q(n11521) );
  OR2X1 U11436 ( .IN1(WX9732), .IN2(n3589), .Q(n11520) );
  OR2X1 U11437 ( .IN1(n11522), .IN2(n11523), .Q(n11519) );
  AND2X1 U11438 ( .IN1(n9326), .IN2(WX9924), .Q(n11523) );
  AND2X1 U11439 ( .IN1(n9582), .IN2(WX9860), .Q(n11522) );
  OR2X1 U11440 ( .IN1(n11524), .IN2(n11525), .Q(WX8436) );
  OR2X1 U11441 ( .IN1(n11526), .IN2(n11527), .Q(n11525) );
  AND2X1 U11442 ( .IN1(n10040), .IN2(CRC_OUT_3_14), .Q(n11527) );
  AND2X1 U11443 ( .IN1(n1471), .IN2(n10015), .Q(n11526) );
  INVX0 U11444 ( .INP(n11528), .ZN(n1471) );
  OR2X1 U11445 ( .IN1(n10645), .IN2(n3862), .Q(n11528) );
  OR2X1 U11446 ( .IN1(n11529), .IN2(n11530), .Q(n11524) );
  AND2X1 U11447 ( .IN1(n9982), .IN2(n11531), .Q(n11530) );
  AND2X1 U11448 ( .IN1(n11023), .IN2(n10060), .Q(n11529) );
  AND2X1 U11449 ( .IN1(n11532), .IN2(n11533), .Q(n11023) );
  INVX0 U11450 ( .INP(n11534), .ZN(n11533) );
  AND2X1 U11451 ( .IN1(n11535), .IN2(n11536), .Q(n11534) );
  OR2X1 U11452 ( .IN1(n11536), .IN2(n11535), .Q(n11532) );
  OR2X1 U11453 ( .IN1(n11537), .IN2(n11538), .Q(n11535) );
  AND2X1 U11454 ( .IN1(n3591), .IN2(WX9730), .Q(n11538) );
  INVX0 U11455 ( .INP(n11539), .ZN(n11537) );
  OR2X1 U11456 ( .IN1(WX9730), .IN2(n3591), .Q(n11539) );
  AND2X1 U11457 ( .IN1(n11540), .IN2(n11541), .Q(n11536) );
  OR2X1 U11458 ( .IN1(WX9858), .IN2(test_so86), .Q(n11541) );
  OR2X1 U11459 ( .IN1(n9907), .IN2(n9328), .Q(n11540) );
  OR2X1 U11460 ( .IN1(n11542), .IN2(n11543), .Q(WX8434) );
  OR2X1 U11461 ( .IN1(n11544), .IN2(n11545), .Q(n11543) );
  AND2X1 U11462 ( .IN1(n10040), .IN2(CRC_OUT_3_15), .Q(n11545) );
  AND2X1 U11463 ( .IN1(n1470), .IN2(n10015), .Q(n11544) );
  INVX0 U11464 ( .INP(n11546), .ZN(n1470) );
  OR2X1 U11465 ( .IN1(n10645), .IN2(n3863), .Q(n11546) );
  OR2X1 U11466 ( .IN1(n11547), .IN2(n11548), .Q(n11542) );
  AND2X1 U11467 ( .IN1(n11549), .IN2(n9975), .Q(n11548) );
  AND2X1 U11468 ( .IN1(n10071), .IN2(n11032), .Q(n11547) );
  OR2X1 U11469 ( .IN1(n11550), .IN2(n11551), .Q(n11032) );
  INVX0 U11470 ( .INP(n11552), .ZN(n11551) );
  OR2X1 U11471 ( .IN1(n11553), .IN2(n11554), .Q(n11552) );
  AND2X1 U11472 ( .IN1(n11554), .IN2(n11553), .Q(n11550) );
  AND2X1 U11473 ( .IN1(n11555), .IN2(n11556), .Q(n11553) );
  OR2X1 U11474 ( .IN1(WX9792), .IN2(n9329), .Q(n11556) );
  OR2X1 U11475 ( .IN1(WX9728), .IN2(n3593), .Q(n11555) );
  OR2X1 U11476 ( .IN1(n11557), .IN2(n11558), .Q(n11554) );
  AND2X1 U11477 ( .IN1(n9330), .IN2(WX9920), .Q(n11558) );
  AND2X1 U11478 ( .IN1(n9581), .IN2(WX9856), .Q(n11557) );
  OR2X1 U11479 ( .IN1(n11559), .IN2(n11560), .Q(WX8432) );
  OR2X1 U11480 ( .IN1(n11561), .IN2(n11562), .Q(n11560) );
  AND2X1 U11481 ( .IN1(n10040), .IN2(CRC_OUT_3_16), .Q(n11562) );
  AND2X1 U11482 ( .IN1(n1469), .IN2(n10015), .Q(n11561) );
  INVX0 U11483 ( .INP(n11563), .ZN(n1469) );
  OR2X1 U11484 ( .IN1(n10645), .IN2(n3864), .Q(n11563) );
  OR2X1 U11485 ( .IN1(n11564), .IN2(n11565), .Q(n11559) );
  AND2X1 U11486 ( .IN1(n9982), .IN2(n11566), .Q(n11565) );
  AND2X1 U11487 ( .IN1(n11041), .IN2(n10059), .Q(n11564) );
  AND2X1 U11488 ( .IN1(n11567), .IN2(n11568), .Q(n11041) );
  INVX0 U11489 ( .INP(n11569), .ZN(n11568) );
  AND2X1 U11490 ( .IN1(n11570), .IN2(n11571), .Q(n11569) );
  OR2X1 U11491 ( .IN1(n11571), .IN2(n11570), .Q(n11567) );
  OR2X1 U11492 ( .IN1(n11572), .IN2(n11573), .Q(n11570) );
  AND2X1 U11493 ( .IN1(n10515), .IN2(WX9790), .Q(n11573) );
  AND2X1 U11494 ( .IN1(n9072), .IN2(n10545), .Q(n11572) );
  AND2X1 U11495 ( .IN1(n11574), .IN2(n11575), .Q(n11571) );
  OR2X1 U11496 ( .IN1(n11576), .IN2(n9515), .Q(n11575) );
  INVX0 U11497 ( .INP(n11577), .ZN(n11576) );
  OR2X1 U11498 ( .IN1(WX9918), .IN2(n11577), .Q(n11574) );
  OR2X1 U11499 ( .IN1(n11578), .IN2(n11579), .Q(n11577) );
  AND2X1 U11500 ( .IN1(n17881), .IN2(n9953), .Q(n11579) );
  AND2X1 U11501 ( .IN1(test_so84), .IN2(n8304), .Q(n11578) );
  OR2X1 U11502 ( .IN1(n11580), .IN2(n11581), .Q(WX8430) );
  OR2X1 U11503 ( .IN1(n11582), .IN2(n11583), .Q(n11581) );
  AND2X1 U11504 ( .IN1(n10041), .IN2(CRC_OUT_3_17), .Q(n11583) );
  AND2X1 U11505 ( .IN1(n1468), .IN2(n10015), .Q(n11582) );
  INVX0 U11506 ( .INP(n11584), .ZN(n1468) );
  OR2X1 U11507 ( .IN1(n10645), .IN2(n3865), .Q(n11584) );
  OR2X1 U11508 ( .IN1(n11585), .IN2(n11586), .Q(n11580) );
  AND2X1 U11509 ( .IN1(n9981), .IN2(n11587), .Q(n11586) );
  AND2X1 U11510 ( .IN1(n10071), .IN2(n11050), .Q(n11585) );
  OR2X1 U11511 ( .IN1(n11588), .IN2(n11589), .Q(n11050) );
  INVX0 U11512 ( .INP(n11590), .ZN(n11589) );
  OR2X1 U11513 ( .IN1(n11591), .IN2(n11592), .Q(n11590) );
  AND2X1 U11514 ( .IN1(n11592), .IN2(n11591), .Q(n11588) );
  INVX0 U11515 ( .INP(n11593), .ZN(n11591) );
  OR2X1 U11516 ( .IN1(n11594), .IN2(n11595), .Q(n11593) );
  AND2X1 U11517 ( .IN1(n10517), .IN2(n8305), .Q(n11595) );
  AND2X1 U11518 ( .IN1(n17882), .IN2(n10545), .Q(n11594) );
  OR2X1 U11519 ( .IN1(n11596), .IN2(n11597), .Q(n11592) );
  AND2X1 U11520 ( .IN1(n9580), .IN2(n11598), .Q(n11597) );
  AND2X1 U11521 ( .IN1(n11599), .IN2(n11600), .Q(n11598) );
  OR2X1 U11522 ( .IN1(n9073), .IN2(WX9852), .Q(n11600) );
  OR2X1 U11523 ( .IN1(n9074), .IN2(WX9788), .Q(n11599) );
  AND2X1 U11524 ( .IN1(n11601), .IN2(WX9916), .Q(n11596) );
  OR2X1 U11525 ( .IN1(n11602), .IN2(n11603), .Q(n11601) );
  AND2X1 U11526 ( .IN1(n9073), .IN2(WX9852), .Q(n11603) );
  AND2X1 U11527 ( .IN1(n9074), .IN2(WX9788), .Q(n11602) );
  OR2X1 U11528 ( .IN1(n11604), .IN2(n11605), .Q(WX8428) );
  OR2X1 U11529 ( .IN1(n11606), .IN2(n11607), .Q(n11605) );
  AND2X1 U11530 ( .IN1(n10041), .IN2(CRC_OUT_3_18), .Q(n11607) );
  AND2X1 U11531 ( .IN1(n1467), .IN2(n10015), .Q(n11606) );
  INVX0 U11532 ( .INP(n11608), .ZN(n1467) );
  OR2X1 U11533 ( .IN1(n10645), .IN2(n3866), .Q(n11608) );
  OR2X1 U11534 ( .IN1(n11609), .IN2(n11610), .Q(n11604) );
  AND2X1 U11535 ( .IN1(n9981), .IN2(n11611), .Q(n11610) );
  AND2X1 U11536 ( .IN1(n11059), .IN2(n10059), .Q(n11609) );
  AND2X1 U11537 ( .IN1(n11612), .IN2(n11613), .Q(n11059) );
  INVX0 U11538 ( .INP(n11614), .ZN(n11613) );
  AND2X1 U11539 ( .IN1(n11615), .IN2(n11616), .Q(n11614) );
  OR2X1 U11540 ( .IN1(n11616), .IN2(n11615), .Q(n11612) );
  OR2X1 U11541 ( .IN1(n11617), .IN2(n11618), .Q(n11615) );
  AND2X1 U11542 ( .IN1(n10518), .IN2(WX9850), .Q(n11618) );
  AND2X1 U11543 ( .IN1(n9075), .IN2(n10545), .Q(n11617) );
  AND2X1 U11544 ( .IN1(n11619), .IN2(n11620), .Q(n11616) );
  OR2X1 U11545 ( .IN1(n11621), .IN2(n9579), .Q(n11620) );
  INVX0 U11546 ( .INP(n11622), .ZN(n11621) );
  OR2X1 U11547 ( .IN1(WX9914), .IN2(n11622), .Q(n11619) );
  OR2X1 U11548 ( .IN1(n11623), .IN2(n11624), .Q(n11622) );
  AND2X1 U11549 ( .IN1(n17883), .IN2(n9954), .Q(n11624) );
  AND2X1 U11550 ( .IN1(test_so82), .IN2(n8306), .Q(n11623) );
  OR2X1 U11551 ( .IN1(n11625), .IN2(n11626), .Q(WX8426) );
  OR2X1 U11552 ( .IN1(n11627), .IN2(n11628), .Q(n11626) );
  AND2X1 U11553 ( .IN1(n10041), .IN2(CRC_OUT_3_19), .Q(n11628) );
  AND2X1 U11554 ( .IN1(n1466), .IN2(n10015), .Q(n11627) );
  INVX0 U11555 ( .INP(n11629), .ZN(n1466) );
  OR2X1 U11556 ( .IN1(n10645), .IN2(n3867), .Q(n11629) );
  OR2X1 U11557 ( .IN1(n11630), .IN2(n11631), .Q(n11625) );
  AND2X1 U11558 ( .IN1(n9981), .IN2(n11632), .Q(n11631) );
  AND2X1 U11559 ( .IN1(n10071), .IN2(n11068), .Q(n11630) );
  OR2X1 U11560 ( .IN1(n11633), .IN2(n11634), .Q(n11068) );
  INVX0 U11561 ( .INP(n11635), .ZN(n11634) );
  OR2X1 U11562 ( .IN1(n11636), .IN2(n11637), .Q(n11635) );
  AND2X1 U11563 ( .IN1(n11637), .IN2(n11636), .Q(n11633) );
  INVX0 U11564 ( .INP(n11638), .ZN(n11636) );
  OR2X1 U11565 ( .IN1(n11639), .IN2(n11640), .Q(n11638) );
  AND2X1 U11566 ( .IN1(n10517), .IN2(n8307), .Q(n11640) );
  AND2X1 U11567 ( .IN1(n17884), .IN2(n10545), .Q(n11639) );
  OR2X1 U11568 ( .IN1(n11641), .IN2(n11642), .Q(n11637) );
  AND2X1 U11569 ( .IN1(n9578), .IN2(n11643), .Q(n11642) );
  AND2X1 U11570 ( .IN1(n11644), .IN2(n11645), .Q(n11643) );
  OR2X1 U11571 ( .IN1(n9076), .IN2(WX9848), .Q(n11645) );
  OR2X1 U11572 ( .IN1(n9077), .IN2(WX9784), .Q(n11644) );
  AND2X1 U11573 ( .IN1(n11646), .IN2(WX9912), .Q(n11641) );
  OR2X1 U11574 ( .IN1(n11647), .IN2(n11648), .Q(n11646) );
  AND2X1 U11575 ( .IN1(n9076), .IN2(WX9848), .Q(n11648) );
  AND2X1 U11576 ( .IN1(n9077), .IN2(WX9784), .Q(n11647) );
  OR2X1 U11577 ( .IN1(n11649), .IN2(n11650), .Q(WX8424) );
  OR2X1 U11578 ( .IN1(n11651), .IN2(n11652), .Q(n11650) );
  AND2X1 U11579 ( .IN1(n10041), .IN2(CRC_OUT_3_20), .Q(n11652) );
  AND2X1 U11580 ( .IN1(n1465), .IN2(n10015), .Q(n11651) );
  INVX0 U11581 ( .INP(n11653), .ZN(n1465) );
  OR2X1 U11582 ( .IN1(n10645), .IN2(n3868), .Q(n11653) );
  OR2X1 U11583 ( .IN1(n11654), .IN2(n11655), .Q(n11649) );
  AND2X1 U11584 ( .IN1(n9981), .IN2(n11656), .Q(n11655) );
  AND2X1 U11585 ( .IN1(n11077), .IN2(n10059), .Q(n11654) );
  AND2X1 U11586 ( .IN1(n11657), .IN2(n11658), .Q(n11077) );
  OR2X1 U11587 ( .IN1(n11659), .IN2(n11660), .Q(n11658) );
  INVX0 U11588 ( .INP(n11661), .ZN(n11659) );
  OR2X1 U11589 ( .IN1(n11662), .IN2(n11661), .Q(n11657) );
  OR2X1 U11590 ( .IN1(n11663), .IN2(n11664), .Q(n11661) );
  AND2X1 U11591 ( .IN1(n10518), .IN2(WX9910), .Q(n11664) );
  AND2X1 U11592 ( .IN1(n9577), .IN2(n10545), .Q(n11663) );
  INVX0 U11593 ( .INP(n11660), .ZN(n11662) );
  OR2X1 U11594 ( .IN1(n11665), .IN2(n11666), .Q(n11660) );
  AND2X1 U11595 ( .IN1(n9079), .IN2(n11667), .Q(n11666) );
  AND2X1 U11596 ( .IN1(n11668), .IN2(n11669), .Q(n11667) );
  OR2X1 U11597 ( .IN1(n9078), .IN2(n9890), .Q(n11669) );
  OR2X1 U11598 ( .IN1(test_so80), .IN2(WX9782), .Q(n11668) );
  AND2X1 U11599 ( .IN1(n11670), .IN2(WX9846), .Q(n11665) );
  OR2X1 U11600 ( .IN1(n11671), .IN2(n11672), .Q(n11670) );
  AND2X1 U11601 ( .IN1(n9078), .IN2(n9890), .Q(n11672) );
  AND2X1 U11602 ( .IN1(test_so80), .IN2(WX9782), .Q(n11671) );
  OR2X1 U11603 ( .IN1(n11673), .IN2(n11674), .Q(WX8422) );
  OR2X1 U11604 ( .IN1(n11675), .IN2(n11676), .Q(n11674) );
  AND2X1 U11605 ( .IN1(n10041), .IN2(CRC_OUT_3_21), .Q(n11676) );
  AND2X1 U11606 ( .IN1(n1464), .IN2(n10015), .Q(n11675) );
  INVX0 U11607 ( .INP(n11677), .ZN(n1464) );
  OR2X1 U11608 ( .IN1(n10645), .IN2(n3869), .Q(n11677) );
  OR2X1 U11609 ( .IN1(n11678), .IN2(n11679), .Q(n11673) );
  AND2X1 U11610 ( .IN1(n9981), .IN2(n11680), .Q(n11679) );
  AND2X1 U11611 ( .IN1(n10072), .IN2(n11086), .Q(n11678) );
  OR2X1 U11612 ( .IN1(n11681), .IN2(n11682), .Q(n11086) );
  INVX0 U11613 ( .INP(n11683), .ZN(n11682) );
  OR2X1 U11614 ( .IN1(n11684), .IN2(n11685), .Q(n11683) );
  AND2X1 U11615 ( .IN1(n11685), .IN2(n11684), .Q(n11681) );
  INVX0 U11616 ( .INP(n11686), .ZN(n11684) );
  OR2X1 U11617 ( .IN1(n11687), .IN2(n11688), .Q(n11686) );
  AND2X1 U11618 ( .IN1(n10518), .IN2(n8310), .Q(n11688) );
  AND2X1 U11619 ( .IN1(n17885), .IN2(n10545), .Q(n11687) );
  OR2X1 U11620 ( .IN1(n11689), .IN2(n11690), .Q(n11685) );
  AND2X1 U11621 ( .IN1(n9576), .IN2(n11691), .Q(n11690) );
  AND2X1 U11622 ( .IN1(n11692), .IN2(n11693), .Q(n11691) );
  OR2X1 U11623 ( .IN1(n9080), .IN2(WX9844), .Q(n11693) );
  OR2X1 U11624 ( .IN1(n9081), .IN2(WX9780), .Q(n11692) );
  AND2X1 U11625 ( .IN1(n11694), .IN2(WX9908), .Q(n11689) );
  OR2X1 U11626 ( .IN1(n11695), .IN2(n11696), .Q(n11694) );
  AND2X1 U11627 ( .IN1(n9080), .IN2(WX9844), .Q(n11696) );
  AND2X1 U11628 ( .IN1(n9081), .IN2(WX9780), .Q(n11695) );
  OR2X1 U11629 ( .IN1(n11697), .IN2(n11698), .Q(WX8420) );
  OR2X1 U11630 ( .IN1(n11699), .IN2(n11700), .Q(n11698) );
  AND2X1 U11631 ( .IN1(n10041), .IN2(CRC_OUT_3_22), .Q(n11700) );
  AND2X1 U11632 ( .IN1(n1463), .IN2(n10015), .Q(n11699) );
  INVX0 U11633 ( .INP(n11701), .ZN(n1463) );
  OR2X1 U11634 ( .IN1(n10645), .IN2(n3870), .Q(n11701) );
  OR2X1 U11635 ( .IN1(n11702), .IN2(n11703), .Q(n11697) );
  AND2X1 U11636 ( .IN1(n9981), .IN2(n11704), .Q(n11703) );
  AND2X1 U11637 ( .IN1(n10072), .IN2(n11095), .Q(n11702) );
  OR2X1 U11638 ( .IN1(n11705), .IN2(n11706), .Q(n11095) );
  INVX0 U11639 ( .INP(n11707), .ZN(n11706) );
  OR2X1 U11640 ( .IN1(n11708), .IN2(n11709), .Q(n11707) );
  AND2X1 U11641 ( .IN1(n11709), .IN2(n11708), .Q(n11705) );
  INVX0 U11642 ( .INP(n11710), .ZN(n11708) );
  OR2X1 U11643 ( .IN1(n11711), .IN2(n11712), .Q(n11710) );
  AND2X1 U11644 ( .IN1(n10518), .IN2(n8311), .Q(n11712) );
  AND2X1 U11645 ( .IN1(n17886), .IN2(n10545), .Q(n11711) );
  OR2X1 U11646 ( .IN1(n11713), .IN2(n11714), .Q(n11709) );
  AND2X1 U11647 ( .IN1(n9575), .IN2(n11715), .Q(n11714) );
  AND2X1 U11648 ( .IN1(n11716), .IN2(n11717), .Q(n11715) );
  OR2X1 U11649 ( .IN1(n9082), .IN2(WX9842), .Q(n11717) );
  OR2X1 U11650 ( .IN1(n9083), .IN2(WX9778), .Q(n11716) );
  AND2X1 U11651 ( .IN1(n11718), .IN2(WX9906), .Q(n11713) );
  OR2X1 U11652 ( .IN1(n11719), .IN2(n11720), .Q(n11718) );
  AND2X1 U11653 ( .IN1(n9082), .IN2(WX9842), .Q(n11720) );
  AND2X1 U11654 ( .IN1(n9083), .IN2(WX9778), .Q(n11719) );
  OR2X1 U11655 ( .IN1(n11721), .IN2(n11722), .Q(WX8418) );
  OR2X1 U11656 ( .IN1(n11723), .IN2(n11724), .Q(n11722) );
  AND2X1 U11657 ( .IN1(n10041), .IN2(CRC_OUT_3_23), .Q(n11724) );
  AND2X1 U11658 ( .IN1(n1462), .IN2(n10016), .Q(n11723) );
  INVX0 U11659 ( .INP(n11725), .ZN(n1462) );
  OR2X1 U11660 ( .IN1(n10645), .IN2(n3871), .Q(n11725) );
  OR2X1 U11661 ( .IN1(n11726), .IN2(n11727), .Q(n11721) );
  AND2X1 U11662 ( .IN1(n9981), .IN2(n11728), .Q(n11727) );
  AND2X1 U11663 ( .IN1(n10072), .IN2(n11104), .Q(n11726) );
  OR2X1 U11664 ( .IN1(n11729), .IN2(n11730), .Q(n11104) );
  INVX0 U11665 ( .INP(n11731), .ZN(n11730) );
  OR2X1 U11666 ( .IN1(n11732), .IN2(n11733), .Q(n11731) );
  AND2X1 U11667 ( .IN1(n11733), .IN2(n11732), .Q(n11729) );
  INVX0 U11668 ( .INP(n11734), .ZN(n11732) );
  OR2X1 U11669 ( .IN1(n11735), .IN2(n11736), .Q(n11734) );
  AND2X1 U11670 ( .IN1(n10518), .IN2(n8312), .Q(n11736) );
  AND2X1 U11671 ( .IN1(n17887), .IN2(n10545), .Q(n11735) );
  OR2X1 U11672 ( .IN1(n11737), .IN2(n11738), .Q(n11733) );
  AND2X1 U11673 ( .IN1(n9574), .IN2(n11739), .Q(n11738) );
  AND2X1 U11674 ( .IN1(n11740), .IN2(n11741), .Q(n11739) );
  OR2X1 U11675 ( .IN1(n9084), .IN2(WX9840), .Q(n11741) );
  OR2X1 U11676 ( .IN1(n9085), .IN2(WX9776), .Q(n11740) );
  AND2X1 U11677 ( .IN1(n11742), .IN2(WX9904), .Q(n11737) );
  OR2X1 U11678 ( .IN1(n11743), .IN2(n11744), .Q(n11742) );
  AND2X1 U11679 ( .IN1(n9084), .IN2(WX9840), .Q(n11744) );
  AND2X1 U11680 ( .IN1(n9085), .IN2(WX9776), .Q(n11743) );
  OR2X1 U11681 ( .IN1(n11745), .IN2(n11746), .Q(WX8416) );
  OR2X1 U11682 ( .IN1(n11747), .IN2(n11748), .Q(n11746) );
  AND2X1 U11683 ( .IN1(test_so77), .IN2(n10026), .Q(n11748) );
  AND2X1 U11684 ( .IN1(n1461), .IN2(n10016), .Q(n11747) );
  INVX0 U11685 ( .INP(n11749), .ZN(n1461) );
  OR2X1 U11686 ( .IN1(n10645), .IN2(n3872), .Q(n11749) );
  OR2X1 U11687 ( .IN1(n11750), .IN2(n11751), .Q(n11745) );
  AND2X1 U11688 ( .IN1(n9981), .IN2(n11752), .Q(n11751) );
  AND2X1 U11689 ( .IN1(n10072), .IN2(n11113), .Q(n11750) );
  OR2X1 U11690 ( .IN1(n11753), .IN2(n11754), .Q(n11113) );
  INVX0 U11691 ( .INP(n11755), .ZN(n11754) );
  OR2X1 U11692 ( .IN1(n11756), .IN2(n11757), .Q(n11755) );
  AND2X1 U11693 ( .IN1(n11757), .IN2(n11756), .Q(n11753) );
  INVX0 U11694 ( .INP(n11758), .ZN(n11756) );
  OR2X1 U11695 ( .IN1(n11759), .IN2(n11760), .Q(n11758) );
  AND2X1 U11696 ( .IN1(n10518), .IN2(n8313), .Q(n11760) );
  AND2X1 U11697 ( .IN1(n17888), .IN2(n10544), .Q(n11759) );
  OR2X1 U11698 ( .IN1(n11761), .IN2(n11762), .Q(n11757) );
  AND2X1 U11699 ( .IN1(n9573), .IN2(n11763), .Q(n11762) );
  AND2X1 U11700 ( .IN1(n11764), .IN2(n11765), .Q(n11763) );
  OR2X1 U11701 ( .IN1(n9086), .IN2(WX9838), .Q(n11765) );
  OR2X1 U11702 ( .IN1(n9087), .IN2(WX9774), .Q(n11764) );
  AND2X1 U11703 ( .IN1(n11766), .IN2(WX9902), .Q(n11761) );
  OR2X1 U11704 ( .IN1(n11767), .IN2(n11768), .Q(n11766) );
  AND2X1 U11705 ( .IN1(n9086), .IN2(WX9838), .Q(n11768) );
  AND2X1 U11706 ( .IN1(n9087), .IN2(WX9774), .Q(n11767) );
  OR2X1 U11707 ( .IN1(n11769), .IN2(n11770), .Q(WX8414) );
  OR2X1 U11708 ( .IN1(n11771), .IN2(n11772), .Q(n11770) );
  AND2X1 U11709 ( .IN1(n10041), .IN2(CRC_OUT_3_25), .Q(n11772) );
  AND2X1 U11710 ( .IN1(n1460), .IN2(n10016), .Q(n11771) );
  INVX0 U11711 ( .INP(n11773), .ZN(n1460) );
  OR2X1 U11712 ( .IN1(n10644), .IN2(n3873), .Q(n11773) );
  OR2X1 U11713 ( .IN1(n11774), .IN2(n11775), .Q(n11769) );
  AND2X1 U11714 ( .IN1(n9981), .IN2(n11776), .Q(n11775) );
  AND2X1 U11715 ( .IN1(n10072), .IN2(n11122), .Q(n11774) );
  OR2X1 U11716 ( .IN1(n11777), .IN2(n11778), .Q(n11122) );
  INVX0 U11717 ( .INP(n11779), .ZN(n11778) );
  OR2X1 U11718 ( .IN1(n11780), .IN2(n11781), .Q(n11779) );
  AND2X1 U11719 ( .IN1(n11781), .IN2(n11780), .Q(n11777) );
  INVX0 U11720 ( .INP(n11782), .ZN(n11780) );
  OR2X1 U11721 ( .IN1(n11783), .IN2(n11784), .Q(n11782) );
  AND2X1 U11722 ( .IN1(n10518), .IN2(n8314), .Q(n11784) );
  AND2X1 U11723 ( .IN1(n17889), .IN2(n10544), .Q(n11783) );
  OR2X1 U11724 ( .IN1(n11785), .IN2(n11786), .Q(n11781) );
  AND2X1 U11725 ( .IN1(n9572), .IN2(n11787), .Q(n11786) );
  AND2X1 U11726 ( .IN1(n11788), .IN2(n11789), .Q(n11787) );
  OR2X1 U11727 ( .IN1(n9088), .IN2(WX9836), .Q(n11789) );
  OR2X1 U11728 ( .IN1(n9089), .IN2(WX9772), .Q(n11788) );
  AND2X1 U11729 ( .IN1(n11790), .IN2(WX9900), .Q(n11785) );
  OR2X1 U11730 ( .IN1(n11791), .IN2(n11792), .Q(n11790) );
  AND2X1 U11731 ( .IN1(n9088), .IN2(WX9836), .Q(n11792) );
  AND2X1 U11732 ( .IN1(n9089), .IN2(WX9772), .Q(n11791) );
  OR2X1 U11733 ( .IN1(n11793), .IN2(n11794), .Q(WX8412) );
  OR2X1 U11734 ( .IN1(n11795), .IN2(n11796), .Q(n11794) );
  AND2X1 U11735 ( .IN1(n10041), .IN2(CRC_OUT_3_26), .Q(n11796) );
  AND2X1 U11736 ( .IN1(n1459), .IN2(n10016), .Q(n11795) );
  INVX0 U11737 ( .INP(n11797), .ZN(n1459) );
  OR2X1 U11738 ( .IN1(n10644), .IN2(n3874), .Q(n11797) );
  OR2X1 U11739 ( .IN1(n11798), .IN2(n11799), .Q(n11793) );
  AND2X1 U11740 ( .IN1(n11800), .IN2(n9976), .Q(n11799) );
  AND2X1 U11741 ( .IN1(n10072), .IN2(n11131), .Q(n11798) );
  OR2X1 U11742 ( .IN1(n11801), .IN2(n11802), .Q(n11131) );
  INVX0 U11743 ( .INP(n11803), .ZN(n11802) );
  OR2X1 U11744 ( .IN1(n11804), .IN2(n11805), .Q(n11803) );
  AND2X1 U11745 ( .IN1(n11805), .IN2(n11804), .Q(n11801) );
  INVX0 U11746 ( .INP(n11806), .ZN(n11804) );
  OR2X1 U11747 ( .IN1(n11807), .IN2(n11808), .Q(n11806) );
  AND2X1 U11748 ( .IN1(n10518), .IN2(n8315), .Q(n11808) );
  AND2X1 U11749 ( .IN1(n17890), .IN2(n10544), .Q(n11807) );
  OR2X1 U11750 ( .IN1(n11809), .IN2(n11810), .Q(n11805) );
  AND2X1 U11751 ( .IN1(n9571), .IN2(n11811), .Q(n11810) );
  AND2X1 U11752 ( .IN1(n11812), .IN2(n11813), .Q(n11811) );
  OR2X1 U11753 ( .IN1(n9090), .IN2(WX9834), .Q(n11813) );
  OR2X1 U11754 ( .IN1(n9091), .IN2(WX9770), .Q(n11812) );
  AND2X1 U11755 ( .IN1(n11814), .IN2(WX9898), .Q(n11809) );
  OR2X1 U11756 ( .IN1(n11815), .IN2(n11816), .Q(n11814) );
  AND2X1 U11757 ( .IN1(n9090), .IN2(WX9834), .Q(n11816) );
  AND2X1 U11758 ( .IN1(n9091), .IN2(WX9770), .Q(n11815) );
  OR2X1 U11759 ( .IN1(n11817), .IN2(n11818), .Q(WX8410) );
  OR2X1 U11760 ( .IN1(n11819), .IN2(n11820), .Q(n11818) );
  AND2X1 U11761 ( .IN1(n10041), .IN2(CRC_OUT_3_27), .Q(n11820) );
  AND2X1 U11762 ( .IN1(n1458), .IN2(n10016), .Q(n11819) );
  INVX0 U11763 ( .INP(n11821), .ZN(n1458) );
  OR2X1 U11764 ( .IN1(n10644), .IN2(n3875), .Q(n11821) );
  OR2X1 U11765 ( .IN1(n11822), .IN2(n11823), .Q(n11817) );
  AND2X1 U11766 ( .IN1(n9981), .IN2(n11824), .Q(n11823) );
  AND2X1 U11767 ( .IN1(n10072), .IN2(n11140), .Q(n11822) );
  OR2X1 U11768 ( .IN1(n11825), .IN2(n11826), .Q(n11140) );
  INVX0 U11769 ( .INP(n11827), .ZN(n11826) );
  OR2X1 U11770 ( .IN1(n11828), .IN2(n11829), .Q(n11827) );
  AND2X1 U11771 ( .IN1(n11829), .IN2(n11828), .Q(n11825) );
  INVX0 U11772 ( .INP(n11830), .ZN(n11828) );
  OR2X1 U11773 ( .IN1(n11831), .IN2(n11832), .Q(n11830) );
  AND2X1 U11774 ( .IN1(n10519), .IN2(n8316), .Q(n11832) );
  AND2X1 U11775 ( .IN1(n17891), .IN2(n10544), .Q(n11831) );
  OR2X1 U11776 ( .IN1(n11833), .IN2(n11834), .Q(n11829) );
  AND2X1 U11777 ( .IN1(n9570), .IN2(n11835), .Q(n11834) );
  AND2X1 U11778 ( .IN1(n11836), .IN2(n11837), .Q(n11835) );
  OR2X1 U11779 ( .IN1(n9092), .IN2(WX9832), .Q(n11837) );
  OR2X1 U11780 ( .IN1(n9093), .IN2(WX9768), .Q(n11836) );
  AND2X1 U11781 ( .IN1(n11838), .IN2(WX9896), .Q(n11833) );
  OR2X1 U11782 ( .IN1(n11839), .IN2(n11840), .Q(n11838) );
  AND2X1 U11783 ( .IN1(n9092), .IN2(WX9832), .Q(n11840) );
  AND2X1 U11784 ( .IN1(n9093), .IN2(WX9768), .Q(n11839) );
  OR2X1 U11785 ( .IN1(n11841), .IN2(n11842), .Q(WX8408) );
  OR2X1 U11786 ( .IN1(n11843), .IN2(n11844), .Q(n11842) );
  AND2X1 U11787 ( .IN1(n10041), .IN2(CRC_OUT_3_28), .Q(n11844) );
  AND2X1 U11788 ( .IN1(n1457), .IN2(n10016), .Q(n11843) );
  INVX0 U11789 ( .INP(n11845), .ZN(n1457) );
  OR2X1 U11790 ( .IN1(n10644), .IN2(n3876), .Q(n11845) );
  OR2X1 U11791 ( .IN1(n11846), .IN2(n11847), .Q(n11841) );
  AND2X1 U11792 ( .IN1(n11848), .IN2(n9977), .Q(n11847) );
  AND2X1 U11793 ( .IN1(n10072), .IN2(n11149), .Q(n11846) );
  OR2X1 U11794 ( .IN1(n11849), .IN2(n11850), .Q(n11149) );
  INVX0 U11795 ( .INP(n11851), .ZN(n11850) );
  OR2X1 U11796 ( .IN1(n11852), .IN2(n11853), .Q(n11851) );
  AND2X1 U11797 ( .IN1(n11853), .IN2(n11852), .Q(n11849) );
  INVX0 U11798 ( .INP(n11854), .ZN(n11852) );
  OR2X1 U11799 ( .IN1(n11855), .IN2(n11856), .Q(n11854) );
  AND2X1 U11800 ( .IN1(n10518), .IN2(n8317), .Q(n11856) );
  AND2X1 U11801 ( .IN1(n17892), .IN2(n10544), .Q(n11855) );
  OR2X1 U11802 ( .IN1(n11857), .IN2(n11858), .Q(n11853) );
  AND2X1 U11803 ( .IN1(n9569), .IN2(n11859), .Q(n11858) );
  AND2X1 U11804 ( .IN1(n11860), .IN2(n11861), .Q(n11859) );
  OR2X1 U11805 ( .IN1(n9094), .IN2(WX9830), .Q(n11861) );
  OR2X1 U11806 ( .IN1(n9095), .IN2(WX9766), .Q(n11860) );
  AND2X1 U11807 ( .IN1(n11862), .IN2(WX9894), .Q(n11857) );
  OR2X1 U11808 ( .IN1(n11863), .IN2(n11864), .Q(n11862) );
  AND2X1 U11809 ( .IN1(n9094), .IN2(WX9830), .Q(n11864) );
  AND2X1 U11810 ( .IN1(n9095), .IN2(WX9766), .Q(n11863) );
  OR2X1 U11811 ( .IN1(n11865), .IN2(n11866), .Q(WX8406) );
  OR2X1 U11812 ( .IN1(n11867), .IN2(n11868), .Q(n11866) );
  AND2X1 U11813 ( .IN1(n10041), .IN2(CRC_OUT_3_29), .Q(n11868) );
  AND2X1 U11814 ( .IN1(n1456), .IN2(n10016), .Q(n11867) );
  INVX0 U11815 ( .INP(n11869), .ZN(n1456) );
  OR2X1 U11816 ( .IN1(n10644), .IN2(n3877), .Q(n11869) );
  OR2X1 U11817 ( .IN1(n11870), .IN2(n11871), .Q(n11865) );
  AND2X1 U11818 ( .IN1(n9981), .IN2(n11872), .Q(n11871) );
  AND2X1 U11819 ( .IN1(n10072), .IN2(n11158), .Q(n11870) );
  OR2X1 U11820 ( .IN1(n11873), .IN2(n11874), .Q(n11158) );
  INVX0 U11821 ( .INP(n11875), .ZN(n11874) );
  OR2X1 U11822 ( .IN1(n11876), .IN2(n11877), .Q(n11875) );
  AND2X1 U11823 ( .IN1(n11877), .IN2(n11876), .Q(n11873) );
  INVX0 U11824 ( .INP(n11878), .ZN(n11876) );
  OR2X1 U11825 ( .IN1(n11879), .IN2(n11880), .Q(n11878) );
  AND2X1 U11826 ( .IN1(n10518), .IN2(n8318), .Q(n11880) );
  AND2X1 U11827 ( .IN1(n17893), .IN2(n10544), .Q(n11879) );
  OR2X1 U11828 ( .IN1(n11881), .IN2(n11882), .Q(n11877) );
  AND2X1 U11829 ( .IN1(n9568), .IN2(n11883), .Q(n11882) );
  AND2X1 U11830 ( .IN1(n11884), .IN2(n11885), .Q(n11883) );
  OR2X1 U11831 ( .IN1(n9096), .IN2(WX9828), .Q(n11885) );
  OR2X1 U11832 ( .IN1(n9097), .IN2(WX9764), .Q(n11884) );
  AND2X1 U11833 ( .IN1(n11886), .IN2(WX9892), .Q(n11881) );
  OR2X1 U11834 ( .IN1(n11887), .IN2(n11888), .Q(n11886) );
  AND2X1 U11835 ( .IN1(n9096), .IN2(WX9828), .Q(n11888) );
  AND2X1 U11836 ( .IN1(n9097), .IN2(WX9764), .Q(n11887) );
  OR2X1 U11837 ( .IN1(n11889), .IN2(n11890), .Q(WX8404) );
  OR2X1 U11838 ( .IN1(n11891), .IN2(n11892), .Q(n11890) );
  AND2X1 U11839 ( .IN1(n10041), .IN2(CRC_OUT_3_30), .Q(n11892) );
  AND2X1 U11840 ( .IN1(n1455), .IN2(n10016), .Q(n11891) );
  INVX0 U11841 ( .INP(n11893), .ZN(n1455) );
  OR2X1 U11842 ( .IN1(n10644), .IN2(n3878), .Q(n11893) );
  OR2X1 U11843 ( .IN1(n11894), .IN2(n11895), .Q(n11889) );
  AND2X1 U11844 ( .IN1(n11896), .IN2(n9976), .Q(n11895) );
  AND2X1 U11845 ( .IN1(n10072), .IN2(n11167), .Q(n11894) );
  OR2X1 U11846 ( .IN1(n11897), .IN2(n11898), .Q(n11167) );
  INVX0 U11847 ( .INP(n11899), .ZN(n11898) );
  OR2X1 U11848 ( .IN1(n11900), .IN2(n11901), .Q(n11899) );
  AND2X1 U11849 ( .IN1(n11901), .IN2(n11900), .Q(n11897) );
  INVX0 U11850 ( .INP(n11902), .ZN(n11900) );
  OR2X1 U11851 ( .IN1(n11903), .IN2(n11904), .Q(n11902) );
  AND2X1 U11852 ( .IN1(n10519), .IN2(n8319), .Q(n11904) );
  AND2X1 U11853 ( .IN1(n17894), .IN2(n10544), .Q(n11903) );
  OR2X1 U11854 ( .IN1(n11905), .IN2(n11906), .Q(n11901) );
  AND2X1 U11855 ( .IN1(n9567), .IN2(n11907), .Q(n11906) );
  AND2X1 U11856 ( .IN1(n11908), .IN2(n11909), .Q(n11907) );
  OR2X1 U11857 ( .IN1(n9098), .IN2(WX9826), .Q(n11909) );
  OR2X1 U11858 ( .IN1(n9099), .IN2(WX9762), .Q(n11908) );
  AND2X1 U11859 ( .IN1(n11910), .IN2(WX9890), .Q(n11905) );
  OR2X1 U11860 ( .IN1(n11911), .IN2(n11912), .Q(n11910) );
  AND2X1 U11861 ( .IN1(n9098), .IN2(WX9826), .Q(n11912) );
  AND2X1 U11862 ( .IN1(n9099), .IN2(WX9762), .Q(n11911) );
  OR2X1 U11863 ( .IN1(n11913), .IN2(n11914), .Q(WX8402) );
  OR2X1 U11864 ( .IN1(n11915), .IN2(n11916), .Q(n11914) );
  AND2X1 U11865 ( .IN1(n2245), .IN2(WX8243), .Q(n11916) );
  AND2X1 U11866 ( .IN1(n10042), .IN2(CRC_OUT_3_31), .Q(n11915) );
  OR2X1 U11867 ( .IN1(n11917), .IN2(n11918), .Q(n11913) );
  AND2X1 U11868 ( .IN1(n9981), .IN2(n11919), .Q(n11918) );
  AND2X1 U11869 ( .IN1(n11175), .IN2(n10059), .Q(n11917) );
  AND2X1 U11870 ( .IN1(n11920), .IN2(n11921), .Q(n11175) );
  INVX0 U11871 ( .INP(n11922), .ZN(n11921) );
  AND2X1 U11872 ( .IN1(n11923), .IN2(n11924), .Q(n11922) );
  OR2X1 U11873 ( .IN1(n11924), .IN2(n11923), .Q(n11920) );
  OR2X1 U11874 ( .IN1(n11925), .IN2(n11926), .Q(n11923) );
  AND2X1 U11875 ( .IN1(n10519), .IN2(WX9760), .Q(n11926) );
  AND2X1 U11876 ( .IN1(n9030), .IN2(n10544), .Q(n11925) );
  AND2X1 U11877 ( .IN1(n11927), .IN2(n11928), .Q(n11924) );
  INVX0 U11878 ( .INP(n11929), .ZN(n11928) );
  AND2X1 U11879 ( .IN1(n11930), .IN2(WX9824), .Q(n11929) );
  OR2X1 U11880 ( .IN1(WX9824), .IN2(n11930), .Q(n11927) );
  OR2X1 U11881 ( .IN1(n11931), .IN2(n11932), .Q(n11930) );
  AND2X1 U11882 ( .IN1(n17895), .IN2(n9914), .Q(n11932) );
  AND2X1 U11883 ( .IN1(test_so85), .IN2(n8320), .Q(n11931) );
  AND2X1 U11884 ( .IN1(n9849), .IN2(n10566), .Q(WX8304) );
  AND2X1 U11885 ( .IN1(n11933), .IN2(n10566), .Q(WX7791) );
  AND2X1 U11886 ( .IN1(n11934), .IN2(n11935), .Q(n11933) );
  OR2X1 U11887 ( .IN1(DFF_1150_n1), .IN2(WX7302), .Q(n11935) );
  OR2X1 U11888 ( .IN1(n9619), .IN2(CRC_OUT_4_30), .Q(n11934) );
  AND2X1 U11889 ( .IN1(n11936), .IN2(n10566), .Q(WX7789) );
  OR2X1 U11890 ( .IN1(n11937), .IN2(n11938), .Q(n11936) );
  AND2X1 U11891 ( .IN1(n9620), .IN2(n9939), .Q(n11938) );
  AND2X1 U11892 ( .IN1(test_so66), .IN2(WX7304), .Q(n11937) );
  AND2X1 U11893 ( .IN1(n11939), .IN2(n10566), .Q(WX7787) );
  AND2X1 U11894 ( .IN1(n11940), .IN2(n11941), .Q(n11939) );
  OR2X1 U11895 ( .IN1(DFF_1148_n1), .IN2(WX7306), .Q(n11941) );
  OR2X1 U11896 ( .IN1(n9621), .IN2(CRC_OUT_4_28), .Q(n11940) );
  AND2X1 U11897 ( .IN1(n11942), .IN2(n10566), .Q(WX7785) );
  AND2X1 U11898 ( .IN1(n11943), .IN2(n11944), .Q(n11942) );
  OR2X1 U11899 ( .IN1(DFF_1147_n1), .IN2(WX7308), .Q(n11944) );
  OR2X1 U11900 ( .IN1(n9622), .IN2(CRC_OUT_4_27), .Q(n11943) );
  AND2X1 U11901 ( .IN1(n11945), .IN2(n10566), .Q(WX7783) );
  AND2X1 U11902 ( .IN1(n11946), .IN2(n11947), .Q(n11945) );
  OR2X1 U11903 ( .IN1(DFF_1146_n1), .IN2(WX7310), .Q(n11947) );
  OR2X1 U11904 ( .IN1(n9623), .IN2(CRC_OUT_4_26), .Q(n11946) );
  AND2X1 U11905 ( .IN1(n11948), .IN2(n10566), .Q(WX7781) );
  AND2X1 U11906 ( .IN1(n11949), .IN2(n11950), .Q(n11948) );
  OR2X1 U11907 ( .IN1(DFF_1145_n1), .IN2(WX7312), .Q(n11950) );
  OR2X1 U11908 ( .IN1(n9624), .IN2(CRC_OUT_4_25), .Q(n11949) );
  AND2X1 U11909 ( .IN1(n11951), .IN2(n10566), .Q(WX7779) );
  AND2X1 U11910 ( .IN1(n11952), .IN2(n11953), .Q(n11951) );
  OR2X1 U11911 ( .IN1(DFF_1144_n1), .IN2(WX7314), .Q(n11953) );
  OR2X1 U11912 ( .IN1(n9625), .IN2(CRC_OUT_4_24), .Q(n11952) );
  AND2X1 U11913 ( .IN1(n11954), .IN2(n10566), .Q(WX7777) );
  AND2X1 U11914 ( .IN1(n11955), .IN2(n11956), .Q(n11954) );
  OR2X1 U11915 ( .IN1(DFF_1143_n1), .IN2(WX7316), .Q(n11956) );
  OR2X1 U11916 ( .IN1(n9626), .IN2(CRC_OUT_4_23), .Q(n11955) );
  AND2X1 U11917 ( .IN1(n11957), .IN2(n10565), .Q(WX7775) );
  AND2X1 U11918 ( .IN1(n11958), .IN2(n11959), .Q(n11957) );
  OR2X1 U11919 ( .IN1(DFF_1142_n1), .IN2(WX7318), .Q(n11959) );
  OR2X1 U11920 ( .IN1(n9627), .IN2(CRC_OUT_4_22), .Q(n11958) );
  AND2X1 U11921 ( .IN1(n11960), .IN2(n10565), .Q(WX7773) );
  AND2X1 U11922 ( .IN1(n11961), .IN2(n11962), .Q(n11960) );
  OR2X1 U11923 ( .IN1(DFF_1141_n1), .IN2(WX7320), .Q(n11962) );
  OR2X1 U11924 ( .IN1(n9628), .IN2(CRC_OUT_4_21), .Q(n11961) );
  AND2X1 U11925 ( .IN1(n11963), .IN2(n10565), .Q(WX7771) );
  OR2X1 U11926 ( .IN1(n11964), .IN2(n11965), .Q(n11963) );
  AND2X1 U11927 ( .IN1(DFF_1140_n1), .IN2(n9909), .Q(n11965) );
  AND2X1 U11928 ( .IN1(test_so63), .IN2(CRC_OUT_4_20), .Q(n11964) );
  AND2X1 U11929 ( .IN1(n11966), .IN2(n10565), .Q(WX7769) );
  AND2X1 U11930 ( .IN1(n11967), .IN2(n11968), .Q(n11966) );
  OR2X1 U11931 ( .IN1(DFF_1139_n1), .IN2(WX7324), .Q(n11968) );
  OR2X1 U11932 ( .IN1(n9629), .IN2(CRC_OUT_4_19), .Q(n11967) );
  AND2X1 U11933 ( .IN1(n11969), .IN2(n10565), .Q(WX7767) );
  AND2X1 U11934 ( .IN1(n11970), .IN2(n11971), .Q(n11969) );
  OR2X1 U11935 ( .IN1(DFF_1138_n1), .IN2(WX7326), .Q(n11971) );
  OR2X1 U11936 ( .IN1(n9630), .IN2(CRC_OUT_4_18), .Q(n11970) );
  AND2X1 U11937 ( .IN1(n11972), .IN2(n10565), .Q(WX7765) );
  AND2X1 U11938 ( .IN1(n11973), .IN2(n11974), .Q(n11972) );
  OR2X1 U11939 ( .IN1(DFF_1137_n1), .IN2(WX7328), .Q(n11974) );
  OR2X1 U11940 ( .IN1(n9631), .IN2(CRC_OUT_4_17), .Q(n11973) );
  AND2X1 U11941 ( .IN1(n11975), .IN2(n10565), .Q(WX7763) );
  AND2X1 U11942 ( .IN1(n11976), .IN2(n11977), .Q(n11975) );
  OR2X1 U11943 ( .IN1(DFF_1136_n1), .IN2(WX7330), .Q(n11977) );
  OR2X1 U11944 ( .IN1(n9632), .IN2(CRC_OUT_4_16), .Q(n11976) );
  AND2X1 U11945 ( .IN1(n11978), .IN2(n10565), .Q(WX7761) );
  OR2X1 U11946 ( .IN1(n11979), .IN2(n11980), .Q(n11978) );
  AND2X1 U11947 ( .IN1(n11981), .IN2(CRC_OUT_4_15), .Q(n11980) );
  AND2X1 U11948 ( .IN1(DFF_1135_n1), .IN2(n11982), .Q(n11979) );
  INVX0 U11949 ( .INP(n11981), .ZN(n11982) );
  OR2X1 U11950 ( .IN1(n11983), .IN2(n11984), .Q(n11981) );
  AND2X1 U11951 ( .IN1(DFF_1151_n1), .IN2(WX7332), .Q(n11984) );
  AND2X1 U11952 ( .IN1(n9521), .IN2(CRC_OUT_4_31), .Q(n11983) );
  AND2X1 U11953 ( .IN1(n11985), .IN2(n10565), .Q(WX7759) );
  AND2X1 U11954 ( .IN1(n11986), .IN2(n11987), .Q(n11985) );
  OR2X1 U11955 ( .IN1(DFF_1134_n1), .IN2(WX7334), .Q(n11987) );
  OR2X1 U11956 ( .IN1(n9633), .IN2(CRC_OUT_4_14), .Q(n11986) );
  AND2X1 U11957 ( .IN1(n11988), .IN2(n10564), .Q(WX7757) );
  AND2X1 U11958 ( .IN1(n11989), .IN2(n11990), .Q(n11988) );
  OR2X1 U11959 ( .IN1(DFF_1133_n1), .IN2(WX7336), .Q(n11990) );
  OR2X1 U11960 ( .IN1(n9634), .IN2(CRC_OUT_4_13), .Q(n11989) );
  AND2X1 U11961 ( .IN1(n11991), .IN2(n10564), .Q(WX7755) );
  OR2X1 U11962 ( .IN1(n11992), .IN2(n11993), .Q(n11991) );
  AND2X1 U11963 ( .IN1(n9635), .IN2(n9940), .Q(n11993) );
  AND2X1 U11964 ( .IN1(test_so65), .IN2(WX7338), .Q(n11992) );
  AND2X1 U11965 ( .IN1(n11994), .IN2(n10564), .Q(WX7753) );
  AND2X1 U11966 ( .IN1(n11995), .IN2(n11996), .Q(n11994) );
  OR2X1 U11967 ( .IN1(DFF_1131_n1), .IN2(WX7340), .Q(n11996) );
  OR2X1 U11968 ( .IN1(n9636), .IN2(CRC_OUT_4_11), .Q(n11995) );
  AND2X1 U11969 ( .IN1(n11997), .IN2(n10564), .Q(WX7751) );
  OR2X1 U11970 ( .IN1(n11998), .IN2(n11999), .Q(n11997) );
  AND2X1 U11971 ( .IN1(n12000), .IN2(CRC_OUT_4_10), .Q(n11999) );
  AND2X1 U11972 ( .IN1(DFF_1130_n1), .IN2(n12001), .Q(n11998) );
  INVX0 U11973 ( .INP(n12000), .ZN(n12001) );
  OR2X1 U11974 ( .IN1(n12002), .IN2(n12003), .Q(n12000) );
  AND2X1 U11975 ( .IN1(DFF_1151_n1), .IN2(WX7342), .Q(n12003) );
  AND2X1 U11976 ( .IN1(n9522), .IN2(CRC_OUT_4_31), .Q(n12002) );
  AND2X1 U11977 ( .IN1(n12004), .IN2(n10564), .Q(WX7749) );
  AND2X1 U11978 ( .IN1(n12005), .IN2(n12006), .Q(n12004) );
  OR2X1 U11979 ( .IN1(DFF_1129_n1), .IN2(WX7344), .Q(n12006) );
  OR2X1 U11980 ( .IN1(n9637), .IN2(CRC_OUT_4_9), .Q(n12005) );
  AND2X1 U11981 ( .IN1(n12007), .IN2(n10564), .Q(WX7747) );
  AND2X1 U11982 ( .IN1(n12008), .IN2(n12009), .Q(n12007) );
  OR2X1 U11983 ( .IN1(DFF_1128_n1), .IN2(WX7346), .Q(n12009) );
  OR2X1 U11984 ( .IN1(n9638), .IN2(CRC_OUT_4_8), .Q(n12008) );
  AND2X1 U11985 ( .IN1(n12010), .IN2(n10564), .Q(WX7745) );
  AND2X1 U11986 ( .IN1(n12011), .IN2(n12012), .Q(n12010) );
  OR2X1 U11987 ( .IN1(DFF_1127_n1), .IN2(WX7348), .Q(n12012) );
  OR2X1 U11988 ( .IN1(n9639), .IN2(CRC_OUT_4_7), .Q(n12011) );
  AND2X1 U11989 ( .IN1(n12013), .IN2(n10564), .Q(WX7743) );
  AND2X1 U11990 ( .IN1(n12014), .IN2(n12015), .Q(n12013) );
  OR2X1 U11991 ( .IN1(DFF_1126_n1), .IN2(WX7350), .Q(n12015) );
  OR2X1 U11992 ( .IN1(n9640), .IN2(CRC_OUT_4_6), .Q(n12014) );
  AND2X1 U11993 ( .IN1(n12016), .IN2(n10564), .Q(WX7741) );
  AND2X1 U11994 ( .IN1(n12017), .IN2(n12018), .Q(n12016) );
  OR2X1 U11995 ( .IN1(DFF_1125_n1), .IN2(WX7352), .Q(n12018) );
  OR2X1 U11996 ( .IN1(n9641), .IN2(CRC_OUT_4_5), .Q(n12017) );
  AND2X1 U11997 ( .IN1(n12019), .IN2(n10563), .Q(WX7739) );
  AND2X1 U11998 ( .IN1(n12020), .IN2(n12021), .Q(n12019) );
  OR2X1 U11999 ( .IN1(DFF_1124_n1), .IN2(WX7354), .Q(n12021) );
  OR2X1 U12000 ( .IN1(n9642), .IN2(CRC_OUT_4_4), .Q(n12020) );
  AND2X1 U12001 ( .IN1(n12022), .IN2(n10563), .Q(WX7737) );
  AND2X1 U12002 ( .IN1(n12023), .IN2(n12024), .Q(n12022) );
  OR2X1 U12003 ( .IN1(DFF_1123_n1), .IN2(n12025), .Q(n12024) );
  AND2X1 U12004 ( .IN1(n12026), .IN2(n12027), .Q(n12025) );
  OR2X1 U12005 ( .IN1(DFF_1151_n1), .IN2(n9886), .Q(n12027) );
  OR2X1 U12006 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .Q(n12026) );
  OR2X1 U12007 ( .IN1(n12028), .IN2(CRC_OUT_4_3), .Q(n12023) );
  OR2X1 U12008 ( .IN1(n12029), .IN2(n12030), .Q(n12028) );
  AND2X1 U12009 ( .IN1(DFF_1151_n1), .IN2(n9886), .Q(n12030) );
  AND2X1 U12010 ( .IN1(test_so64), .IN2(CRC_OUT_4_31), .Q(n12029) );
  AND2X1 U12011 ( .IN1(n12031), .IN2(n10563), .Q(WX7735) );
  AND2X1 U12012 ( .IN1(n12032), .IN2(n12033), .Q(n12031) );
  OR2X1 U12013 ( .IN1(DFF_1122_n1), .IN2(WX7358), .Q(n12033) );
  OR2X1 U12014 ( .IN1(n9643), .IN2(CRC_OUT_4_2), .Q(n12032) );
  AND2X1 U12015 ( .IN1(n12034), .IN2(n10563), .Q(WX7733) );
  AND2X1 U12016 ( .IN1(n12035), .IN2(n12036), .Q(n12034) );
  OR2X1 U12017 ( .IN1(DFF_1121_n1), .IN2(WX7360), .Q(n12036) );
  OR2X1 U12018 ( .IN1(n9644), .IN2(CRC_OUT_4_1), .Q(n12035) );
  AND2X1 U12019 ( .IN1(n12037), .IN2(n10563), .Q(WX7731) );
  AND2X1 U12020 ( .IN1(n12038), .IN2(n12039), .Q(n12037) );
  OR2X1 U12021 ( .IN1(DFF_1120_n1), .IN2(WX7362), .Q(n12039) );
  OR2X1 U12022 ( .IN1(n9645), .IN2(CRC_OUT_4_0), .Q(n12038) );
  AND2X1 U12023 ( .IN1(n12040), .IN2(n10563), .Q(WX7729) );
  AND2X1 U12024 ( .IN1(n12041), .IN2(n12042), .Q(n12040) );
  OR2X1 U12025 ( .IN1(DFF_1151_n1), .IN2(WX7364), .Q(n12042) );
  OR2X1 U12026 ( .IN1(n9536), .IN2(CRC_OUT_4_31), .Q(n12041) );
  AND2X1 U12027 ( .IN1(n10591), .IN2(n8421), .Q(WX7203) );
  AND2X1 U12028 ( .IN1(n10602), .IN2(n8422), .Q(WX7201) );
  AND2X1 U12029 ( .IN1(n10602), .IN2(n8423), .Q(WX7199) );
  AND2X1 U12030 ( .IN1(n10602), .IN2(n8424), .Q(WX7197) );
  AND2X1 U12031 ( .IN1(n10602), .IN2(n8425), .Q(WX7195) );
  AND2X1 U12032 ( .IN1(n10602), .IN2(n8426), .Q(WX7193) );
  AND2X1 U12033 ( .IN1(n10602), .IN2(n8427), .Q(WX7191) );
  AND2X1 U12034 ( .IN1(n10602), .IN2(n8428), .Q(WX7189) );
  AND2X1 U12035 ( .IN1(n10602), .IN2(n8429), .Q(WX7187) );
  AND2X1 U12036 ( .IN1(n10601), .IN2(n8430), .Q(WX7185) );
  AND2X1 U12037 ( .IN1(n10601), .IN2(n8431), .Q(WX7183) );
  AND2X1 U12038 ( .IN1(test_so57), .IN2(n10563), .Q(WX7181) );
  AND2X1 U12039 ( .IN1(n10601), .IN2(n8434), .Q(WX7179) );
  AND2X1 U12040 ( .IN1(n10601), .IN2(n8435), .Q(WX7177) );
  AND2X1 U12041 ( .IN1(n10600), .IN2(n8436), .Q(WX7175) );
  AND2X1 U12042 ( .IN1(n10599), .IN2(n8437), .Q(WX7173) );
  OR2X1 U12043 ( .IN1(n12043), .IN2(n12044), .Q(WX7171) );
  OR2X1 U12044 ( .IN1(n12045), .IN2(n12046), .Q(n12044) );
  AND2X1 U12045 ( .IN1(n10042), .IN2(CRC_OUT_4_0), .Q(n12046) );
  AND2X1 U12046 ( .IN1(n1244), .IN2(n10016), .Q(n12045) );
  INVX0 U12047 ( .INP(n12047), .ZN(n1244) );
  OR2X1 U12048 ( .IN1(n10644), .IN2(n3879), .Q(n12047) );
  OR2X1 U12049 ( .IN1(n12048), .IN2(n12049), .Q(n12043) );
  AND2X1 U12050 ( .IN1(n9981), .IN2(n12050), .Q(n12049) );
  AND2X1 U12051 ( .IN1(n10072), .IN2(n11291), .Q(n12048) );
  OR2X1 U12052 ( .IN1(n12051), .IN2(n12052), .Q(n11291) );
  INVX0 U12053 ( .INP(n12053), .ZN(n12052) );
  OR2X1 U12054 ( .IN1(n12054), .IN2(n12055), .Q(n12053) );
  AND2X1 U12055 ( .IN1(n12055), .IN2(n12054), .Q(n12051) );
  AND2X1 U12056 ( .IN1(n12056), .IN2(n12057), .Q(n12054) );
  OR2X1 U12057 ( .IN1(WX8529), .IN2(n9331), .Q(n12057) );
  OR2X1 U12058 ( .IN1(WX8465), .IN2(n3595), .Q(n12056) );
  OR2X1 U12059 ( .IN1(n12058), .IN2(n12059), .Q(n12055) );
  AND2X1 U12060 ( .IN1(n9332), .IN2(WX8657), .Q(n12059) );
  AND2X1 U12061 ( .IN1(n9535), .IN2(WX8593), .Q(n12058) );
  OR2X1 U12062 ( .IN1(n12060), .IN2(n12061), .Q(WX7169) );
  OR2X1 U12063 ( .IN1(n12062), .IN2(n12063), .Q(n12061) );
  AND2X1 U12064 ( .IN1(n10042), .IN2(CRC_OUT_4_1), .Q(n12063) );
  AND2X1 U12065 ( .IN1(n1243), .IN2(n10016), .Q(n12062) );
  INVX0 U12066 ( .INP(n12064), .ZN(n1243) );
  OR2X1 U12067 ( .IN1(n10644), .IN2(n3880), .Q(n12064) );
  OR2X1 U12068 ( .IN1(n12065), .IN2(n12066), .Q(n12060) );
  AND2X1 U12069 ( .IN1(n9980), .IN2(n12067), .Q(n12066) );
  AND2X1 U12070 ( .IN1(n10072), .IN2(n11308), .Q(n12065) );
  OR2X1 U12071 ( .IN1(n12068), .IN2(n12069), .Q(n11308) );
  INVX0 U12072 ( .INP(n12070), .ZN(n12069) );
  OR2X1 U12073 ( .IN1(n12071), .IN2(n12072), .Q(n12070) );
  AND2X1 U12074 ( .IN1(n12072), .IN2(n12071), .Q(n12068) );
  AND2X1 U12075 ( .IN1(n12073), .IN2(n12074), .Q(n12071) );
  OR2X1 U12076 ( .IN1(WX8527), .IN2(n9333), .Q(n12074) );
  OR2X1 U12077 ( .IN1(WX8463), .IN2(n3597), .Q(n12073) );
  OR2X1 U12078 ( .IN1(n12075), .IN2(n12076), .Q(n12072) );
  AND2X1 U12079 ( .IN1(n9334), .IN2(WX8655), .Q(n12076) );
  AND2X1 U12080 ( .IN1(n9618), .IN2(WX8591), .Q(n12075) );
  OR2X1 U12081 ( .IN1(n12077), .IN2(n12078), .Q(WX7167) );
  OR2X1 U12082 ( .IN1(n12079), .IN2(n12080), .Q(n12078) );
  AND2X1 U12083 ( .IN1(n10042), .IN2(CRC_OUT_4_2), .Q(n12080) );
  AND2X1 U12084 ( .IN1(n1242), .IN2(n10016), .Q(n12079) );
  INVX0 U12085 ( .INP(n12081), .ZN(n1242) );
  OR2X1 U12086 ( .IN1(n10644), .IN2(n3881), .Q(n12081) );
  OR2X1 U12087 ( .IN1(n12082), .IN2(n12083), .Q(n12077) );
  AND2X1 U12088 ( .IN1(n9980), .IN2(n12084), .Q(n12083) );
  AND2X1 U12089 ( .IN1(n10072), .IN2(n11326), .Q(n12082) );
  OR2X1 U12090 ( .IN1(n12085), .IN2(n12086), .Q(n11326) );
  INVX0 U12091 ( .INP(n12087), .ZN(n12086) );
  OR2X1 U12092 ( .IN1(n12088), .IN2(n12089), .Q(n12087) );
  AND2X1 U12093 ( .IN1(n12089), .IN2(n12088), .Q(n12085) );
  AND2X1 U12094 ( .IN1(n12090), .IN2(n12091), .Q(n12088) );
  OR2X1 U12095 ( .IN1(WX8525), .IN2(n9335), .Q(n12091) );
  OR2X1 U12096 ( .IN1(WX8461), .IN2(n3599), .Q(n12090) );
  OR2X1 U12097 ( .IN1(n12092), .IN2(n12093), .Q(n12089) );
  AND2X1 U12098 ( .IN1(n9336), .IN2(WX8653), .Q(n12093) );
  AND2X1 U12099 ( .IN1(n9617), .IN2(WX8589), .Q(n12092) );
  OR2X1 U12100 ( .IN1(n12094), .IN2(n12095), .Q(WX7165) );
  OR2X1 U12101 ( .IN1(n12096), .IN2(n12097), .Q(n12095) );
  AND2X1 U12102 ( .IN1(n10042), .IN2(CRC_OUT_4_3), .Q(n12097) );
  AND2X1 U12103 ( .IN1(n1241), .IN2(n10016), .Q(n12096) );
  INVX0 U12104 ( .INP(n12098), .ZN(n1241) );
  OR2X1 U12105 ( .IN1(n10644), .IN2(n3882), .Q(n12098) );
  OR2X1 U12106 ( .IN1(n12099), .IN2(n12100), .Q(n12094) );
  AND2X1 U12107 ( .IN1(n9980), .IN2(n12101), .Q(n12100) );
  AND2X1 U12108 ( .IN1(n10073), .IN2(n11343), .Q(n12099) );
  OR2X1 U12109 ( .IN1(n12102), .IN2(n12103), .Q(n11343) );
  INVX0 U12110 ( .INP(n12104), .ZN(n12103) );
  OR2X1 U12111 ( .IN1(n12105), .IN2(n12106), .Q(n12104) );
  AND2X1 U12112 ( .IN1(n12106), .IN2(n12105), .Q(n12102) );
  AND2X1 U12113 ( .IN1(n12107), .IN2(n12108), .Q(n12105) );
  OR2X1 U12114 ( .IN1(WX8523), .IN2(n9337), .Q(n12108) );
  OR2X1 U12115 ( .IN1(WX8459), .IN2(n3601), .Q(n12107) );
  OR2X1 U12116 ( .IN1(n12109), .IN2(n12110), .Q(n12106) );
  AND2X1 U12117 ( .IN1(n9338), .IN2(WX8651), .Q(n12110) );
  AND2X1 U12118 ( .IN1(n9616), .IN2(WX8587), .Q(n12109) );
  OR2X1 U12119 ( .IN1(n12111), .IN2(n12112), .Q(WX7163) );
  OR2X1 U12120 ( .IN1(n12113), .IN2(n12114), .Q(n12112) );
  AND2X1 U12121 ( .IN1(n10042), .IN2(CRC_OUT_4_4), .Q(n12114) );
  AND2X1 U12122 ( .IN1(n1240), .IN2(n10017), .Q(n12113) );
  INVX0 U12123 ( .INP(n12115), .ZN(n1240) );
  OR2X1 U12124 ( .IN1(n10644), .IN2(n3883), .Q(n12115) );
  OR2X1 U12125 ( .IN1(n12116), .IN2(n12117), .Q(n12111) );
  AND2X1 U12126 ( .IN1(n12118), .IN2(n9974), .Q(n12117) );
  AND2X1 U12127 ( .IN1(n10073), .IN2(n11361), .Q(n12116) );
  OR2X1 U12128 ( .IN1(n12119), .IN2(n12120), .Q(n11361) );
  INVX0 U12129 ( .INP(n12121), .ZN(n12120) );
  OR2X1 U12130 ( .IN1(n12122), .IN2(n12123), .Q(n12121) );
  AND2X1 U12131 ( .IN1(n12123), .IN2(n12122), .Q(n12119) );
  AND2X1 U12132 ( .IN1(n12124), .IN2(n12125), .Q(n12122) );
  OR2X1 U12133 ( .IN1(WX8521), .IN2(n9339), .Q(n12125) );
  OR2X1 U12134 ( .IN1(WX8457), .IN2(n3603), .Q(n12124) );
  OR2X1 U12135 ( .IN1(n12126), .IN2(n12127), .Q(n12123) );
  AND2X1 U12136 ( .IN1(n9340), .IN2(WX8649), .Q(n12127) );
  AND2X1 U12137 ( .IN1(n9520), .IN2(WX8585), .Q(n12126) );
  OR2X1 U12138 ( .IN1(n12128), .IN2(n12129), .Q(WX7161) );
  OR2X1 U12139 ( .IN1(n12130), .IN2(n12131), .Q(n12129) );
  AND2X1 U12140 ( .IN1(n10042), .IN2(CRC_OUT_4_5), .Q(n12131) );
  AND2X1 U12141 ( .IN1(n1239), .IN2(n10017), .Q(n12130) );
  INVX0 U12142 ( .INP(n12132), .ZN(n1239) );
  OR2X1 U12143 ( .IN1(n10644), .IN2(n3884), .Q(n12132) );
  OR2X1 U12144 ( .IN1(n12133), .IN2(n12134), .Q(n12128) );
  AND2X1 U12145 ( .IN1(n9980), .IN2(n12135), .Q(n12134) );
  AND2X1 U12146 ( .IN1(n10073), .IN2(n11378), .Q(n12133) );
  OR2X1 U12147 ( .IN1(n12136), .IN2(n12137), .Q(n11378) );
  INVX0 U12148 ( .INP(n12138), .ZN(n12137) );
  OR2X1 U12149 ( .IN1(n12139), .IN2(n12140), .Q(n12138) );
  AND2X1 U12150 ( .IN1(n12140), .IN2(n12139), .Q(n12136) );
  AND2X1 U12151 ( .IN1(n12141), .IN2(n12142), .Q(n12139) );
  OR2X1 U12152 ( .IN1(WX8519), .IN2(n9341), .Q(n12142) );
  OR2X1 U12153 ( .IN1(WX8455), .IN2(n3605), .Q(n12141) );
  OR2X1 U12154 ( .IN1(n12143), .IN2(n12144), .Q(n12140) );
  AND2X1 U12155 ( .IN1(n9342), .IN2(WX8647), .Q(n12144) );
  AND2X1 U12156 ( .IN1(n9615), .IN2(WX8583), .Q(n12143) );
  OR2X1 U12157 ( .IN1(n12145), .IN2(n12146), .Q(WX7159) );
  OR2X1 U12158 ( .IN1(n12147), .IN2(n12148), .Q(n12146) );
  AND2X1 U12159 ( .IN1(n10042), .IN2(CRC_OUT_4_6), .Q(n12148) );
  AND2X1 U12160 ( .IN1(n1238), .IN2(n10017), .Q(n12147) );
  INVX0 U12161 ( .INP(n12149), .ZN(n1238) );
  OR2X1 U12162 ( .IN1(n10643), .IN2(n3885), .Q(n12149) );
  OR2X1 U12163 ( .IN1(n12150), .IN2(n12151), .Q(n12145) );
  AND2X1 U12164 ( .IN1(n12152), .IN2(n9974), .Q(n12151) );
  AND2X1 U12165 ( .IN1(n10073), .IN2(n11395), .Q(n12150) );
  OR2X1 U12166 ( .IN1(n12153), .IN2(n12154), .Q(n11395) );
  INVX0 U12167 ( .INP(n12155), .ZN(n12154) );
  OR2X1 U12168 ( .IN1(n12156), .IN2(n12157), .Q(n12155) );
  AND2X1 U12169 ( .IN1(n12157), .IN2(n12156), .Q(n12153) );
  AND2X1 U12170 ( .IN1(n12158), .IN2(n12159), .Q(n12156) );
  OR2X1 U12171 ( .IN1(WX8517), .IN2(n9343), .Q(n12159) );
  OR2X1 U12172 ( .IN1(WX8453), .IN2(n3607), .Q(n12158) );
  OR2X1 U12173 ( .IN1(n12160), .IN2(n12161), .Q(n12157) );
  AND2X1 U12174 ( .IN1(n9344), .IN2(WX8645), .Q(n12161) );
  AND2X1 U12175 ( .IN1(n9614), .IN2(WX8581), .Q(n12160) );
  OR2X1 U12176 ( .IN1(n12162), .IN2(n12163), .Q(WX7157) );
  OR2X1 U12177 ( .IN1(n12164), .IN2(n12165), .Q(n12163) );
  AND2X1 U12178 ( .IN1(n10042), .IN2(CRC_OUT_4_7), .Q(n12165) );
  AND2X1 U12179 ( .IN1(n1237), .IN2(n10017), .Q(n12164) );
  INVX0 U12180 ( .INP(n12166), .ZN(n1237) );
  OR2X1 U12181 ( .IN1(n10643), .IN2(n3886), .Q(n12166) );
  OR2X1 U12182 ( .IN1(n12167), .IN2(n12168), .Q(n12162) );
  AND2X1 U12183 ( .IN1(n9980), .IN2(n12169), .Q(n12168) );
  AND2X1 U12184 ( .IN1(n10073), .IN2(n11412), .Q(n12167) );
  OR2X1 U12185 ( .IN1(n12170), .IN2(n12171), .Q(n11412) );
  INVX0 U12186 ( .INP(n12172), .ZN(n12171) );
  OR2X1 U12187 ( .IN1(n12173), .IN2(n12174), .Q(n12172) );
  AND2X1 U12188 ( .IN1(n12174), .IN2(n12173), .Q(n12170) );
  AND2X1 U12189 ( .IN1(n12175), .IN2(n12176), .Q(n12173) );
  OR2X1 U12190 ( .IN1(WX8515), .IN2(n9345), .Q(n12176) );
  OR2X1 U12191 ( .IN1(WX8451), .IN2(n3609), .Q(n12175) );
  OR2X1 U12192 ( .IN1(n12177), .IN2(n12178), .Q(n12174) );
  AND2X1 U12193 ( .IN1(n9346), .IN2(WX8643), .Q(n12178) );
  AND2X1 U12194 ( .IN1(n9613), .IN2(WX8579), .Q(n12177) );
  OR2X1 U12195 ( .IN1(n12179), .IN2(n12180), .Q(WX7155) );
  OR2X1 U12196 ( .IN1(n12181), .IN2(n12182), .Q(n12180) );
  AND2X1 U12197 ( .IN1(n10042), .IN2(CRC_OUT_4_8), .Q(n12182) );
  AND2X1 U12198 ( .IN1(n1236), .IN2(n10017), .Q(n12181) );
  INVX0 U12199 ( .INP(n12183), .ZN(n1236) );
  OR2X1 U12200 ( .IN1(n10643), .IN2(n3887), .Q(n12183) );
  OR2X1 U12201 ( .IN1(n12184), .IN2(n12185), .Q(n12179) );
  AND2X1 U12202 ( .IN1(n12186), .IN2(n9973), .Q(n12185) );
  AND2X1 U12203 ( .IN1(n10073), .IN2(n11429), .Q(n12184) );
  OR2X1 U12204 ( .IN1(n12187), .IN2(n12188), .Q(n11429) );
  INVX0 U12205 ( .INP(n12189), .ZN(n12188) );
  OR2X1 U12206 ( .IN1(n12190), .IN2(n12191), .Q(n12189) );
  AND2X1 U12207 ( .IN1(n12191), .IN2(n12190), .Q(n12187) );
  AND2X1 U12208 ( .IN1(n12192), .IN2(n12193), .Q(n12190) );
  OR2X1 U12209 ( .IN1(WX8513), .IN2(n9347), .Q(n12193) );
  OR2X1 U12210 ( .IN1(WX8449), .IN2(n3611), .Q(n12192) );
  OR2X1 U12211 ( .IN1(n12194), .IN2(n12195), .Q(n12191) );
  AND2X1 U12212 ( .IN1(n9348), .IN2(WX8641), .Q(n12195) );
  AND2X1 U12213 ( .IN1(n9612), .IN2(WX8577), .Q(n12194) );
  OR2X1 U12214 ( .IN1(n12196), .IN2(n12197), .Q(WX7153) );
  OR2X1 U12215 ( .IN1(n12198), .IN2(n12199), .Q(n12197) );
  AND2X1 U12216 ( .IN1(n10042), .IN2(CRC_OUT_4_9), .Q(n12199) );
  AND2X1 U12217 ( .IN1(n1235), .IN2(n10017), .Q(n12198) );
  INVX0 U12218 ( .INP(n12200), .ZN(n1235) );
  OR2X1 U12219 ( .IN1(n10643), .IN2(n3888), .Q(n12200) );
  OR2X1 U12220 ( .IN1(n12201), .IN2(n12202), .Q(n12196) );
  AND2X1 U12221 ( .IN1(n9980), .IN2(n12203), .Q(n12202) );
  AND2X1 U12222 ( .IN1(n11446), .IN2(n10058), .Q(n12201) );
  AND2X1 U12223 ( .IN1(n12204), .IN2(n12205), .Q(n11446) );
  INVX0 U12224 ( .INP(n12206), .ZN(n12205) );
  AND2X1 U12225 ( .IN1(n12207), .IN2(n12208), .Q(n12206) );
  OR2X1 U12226 ( .IN1(n12208), .IN2(n12207), .Q(n12204) );
  OR2X1 U12227 ( .IN1(n12209), .IN2(n12210), .Q(n12207) );
  AND2X1 U12228 ( .IN1(n3613), .IN2(WX8447), .Q(n12210) );
  INVX0 U12229 ( .INP(n12211), .ZN(n12209) );
  OR2X1 U12230 ( .IN1(WX8447), .IN2(n3613), .Q(n12211) );
  AND2X1 U12231 ( .IN1(n12212), .IN2(n12213), .Q(n12208) );
  OR2X1 U12232 ( .IN1(WX8575), .IN2(test_so75), .Q(n12213) );
  OR2X1 U12233 ( .IN1(n9903), .IN2(n9350), .Q(n12212) );
  OR2X1 U12234 ( .IN1(n12214), .IN2(n12215), .Q(WX7151) );
  OR2X1 U12235 ( .IN1(n12216), .IN2(n12217), .Q(n12215) );
  AND2X1 U12236 ( .IN1(n10042), .IN2(CRC_OUT_4_10), .Q(n12217) );
  AND2X1 U12237 ( .IN1(n1234), .IN2(n10017), .Q(n12216) );
  INVX0 U12238 ( .INP(n12218), .ZN(n1234) );
  OR2X1 U12239 ( .IN1(n10643), .IN2(n3889), .Q(n12218) );
  OR2X1 U12240 ( .IN1(n12219), .IN2(n12220), .Q(n12214) );
  AND2X1 U12241 ( .IN1(n12221), .IN2(n9973), .Q(n12220) );
  AND2X1 U12242 ( .IN1(n10073), .IN2(n11463), .Q(n12219) );
  OR2X1 U12243 ( .IN1(n12222), .IN2(n12223), .Q(n11463) );
  INVX0 U12244 ( .INP(n12224), .ZN(n12223) );
  OR2X1 U12245 ( .IN1(n12225), .IN2(n12226), .Q(n12224) );
  AND2X1 U12246 ( .IN1(n12226), .IN2(n12225), .Q(n12222) );
  AND2X1 U12247 ( .IN1(n12227), .IN2(n12228), .Q(n12225) );
  OR2X1 U12248 ( .IN1(WX8509), .IN2(n9351), .Q(n12228) );
  OR2X1 U12249 ( .IN1(WX8445), .IN2(n3615), .Q(n12227) );
  OR2X1 U12250 ( .IN1(n12229), .IN2(n12230), .Q(n12226) );
  AND2X1 U12251 ( .IN1(n9352), .IN2(WX8637), .Q(n12230) );
  AND2X1 U12252 ( .IN1(n9611), .IN2(WX8573), .Q(n12229) );
  OR2X1 U12253 ( .IN1(n12231), .IN2(n12232), .Q(WX7149) );
  OR2X1 U12254 ( .IN1(n12233), .IN2(n12234), .Q(n12232) );
  AND2X1 U12255 ( .IN1(n10043), .IN2(CRC_OUT_4_11), .Q(n12234) );
  AND2X1 U12256 ( .IN1(n1233), .IN2(n10017), .Q(n12233) );
  INVX0 U12257 ( .INP(n12235), .ZN(n1233) );
  OR2X1 U12258 ( .IN1(n10643), .IN2(n3890), .Q(n12235) );
  OR2X1 U12259 ( .IN1(n12236), .IN2(n12237), .Q(n12231) );
  AND2X1 U12260 ( .IN1(n9980), .IN2(n12238), .Q(n12237) );
  AND2X1 U12261 ( .IN1(n11480), .IN2(n10058), .Q(n12236) );
  AND2X1 U12262 ( .IN1(n12239), .IN2(n12240), .Q(n11480) );
  INVX0 U12263 ( .INP(n12241), .ZN(n12240) );
  AND2X1 U12264 ( .IN1(n12242), .IN2(n12243), .Q(n12241) );
  OR2X1 U12265 ( .IN1(n12243), .IN2(n12242), .Q(n12239) );
  OR2X1 U12266 ( .IN1(n12244), .IN2(n12245), .Q(n12242) );
  AND2X1 U12267 ( .IN1(n3617), .IN2(WX8443), .Q(n12245) );
  INVX0 U12268 ( .INP(n12246), .ZN(n12244) );
  OR2X1 U12269 ( .IN1(WX8443), .IN2(n3617), .Q(n12246) );
  AND2X1 U12270 ( .IN1(n12247), .IN2(n12248), .Q(n12243) );
  OR2X1 U12271 ( .IN1(WX8635), .IN2(test_so73), .Q(n12248) );
  OR2X1 U12272 ( .IN1(n9917), .IN2(n9519), .Q(n12247) );
  OR2X1 U12273 ( .IN1(n12249), .IN2(n12250), .Q(WX7147) );
  OR2X1 U12274 ( .IN1(n12251), .IN2(n12252), .Q(n12250) );
  AND2X1 U12275 ( .IN1(test_so65), .IN2(n10026), .Q(n12252) );
  AND2X1 U12276 ( .IN1(n1232), .IN2(n10017), .Q(n12251) );
  INVX0 U12277 ( .INP(n12253), .ZN(n1232) );
  OR2X1 U12278 ( .IN1(n10643), .IN2(n3891), .Q(n12253) );
  OR2X1 U12279 ( .IN1(n12254), .IN2(n12255), .Q(n12249) );
  AND2X1 U12280 ( .IN1(n9980), .IN2(n12256), .Q(n12255) );
  AND2X1 U12281 ( .IN1(n10073), .IN2(n11497), .Q(n12254) );
  OR2X1 U12282 ( .IN1(n12257), .IN2(n12258), .Q(n11497) );
  INVX0 U12283 ( .INP(n12259), .ZN(n12258) );
  OR2X1 U12284 ( .IN1(n12260), .IN2(n12261), .Q(n12259) );
  AND2X1 U12285 ( .IN1(n12261), .IN2(n12260), .Q(n12257) );
  AND2X1 U12286 ( .IN1(n12262), .IN2(n12263), .Q(n12260) );
  OR2X1 U12287 ( .IN1(WX8505), .IN2(n9354), .Q(n12263) );
  OR2X1 U12288 ( .IN1(WX8441), .IN2(n3619), .Q(n12262) );
  OR2X1 U12289 ( .IN1(n12264), .IN2(n12265), .Q(n12261) );
  AND2X1 U12290 ( .IN1(n9355), .IN2(WX8633), .Q(n12265) );
  AND2X1 U12291 ( .IN1(n9610), .IN2(WX8569), .Q(n12264) );
  OR2X1 U12292 ( .IN1(n12266), .IN2(n12267), .Q(WX7145) );
  OR2X1 U12293 ( .IN1(n12268), .IN2(n12269), .Q(n12267) );
  AND2X1 U12294 ( .IN1(n10043), .IN2(CRC_OUT_4_13), .Q(n12269) );
  AND2X1 U12295 ( .IN1(n1231), .IN2(n10017), .Q(n12268) );
  INVX0 U12296 ( .INP(n12270), .ZN(n1231) );
  OR2X1 U12297 ( .IN1(n10643), .IN2(n3892), .Q(n12270) );
  OR2X1 U12298 ( .IN1(n12271), .IN2(n12272), .Q(n12266) );
  AND2X1 U12299 ( .IN1(n9980), .IN2(n12273), .Q(n12272) );
  AND2X1 U12300 ( .IN1(n11514), .IN2(n10058), .Q(n12271) );
  AND2X1 U12301 ( .IN1(n12274), .IN2(n12275), .Q(n11514) );
  INVX0 U12302 ( .INP(n12276), .ZN(n12275) );
  AND2X1 U12303 ( .IN1(n12277), .IN2(n12278), .Q(n12276) );
  OR2X1 U12304 ( .IN1(n12278), .IN2(n12277), .Q(n12274) );
  OR2X1 U12305 ( .IN1(n12279), .IN2(n12280), .Q(n12277) );
  AND2X1 U12306 ( .IN1(n9356), .IN2(WX8567), .Q(n12280) );
  INVX0 U12307 ( .INP(n12281), .ZN(n12279) );
  OR2X1 U12308 ( .IN1(WX8567), .IN2(n9356), .Q(n12281) );
  AND2X1 U12309 ( .IN1(n12282), .IN2(n12283), .Q(n12278) );
  OR2X1 U12310 ( .IN1(WX8631), .IN2(test_so71), .Q(n12283) );
  OR2X1 U12311 ( .IN1(n9918), .IN2(n9609), .Q(n12282) );
  OR2X1 U12312 ( .IN1(n12284), .IN2(n12285), .Q(WX7143) );
  OR2X1 U12313 ( .IN1(n12286), .IN2(n12287), .Q(n12285) );
  AND2X1 U12314 ( .IN1(n10043), .IN2(CRC_OUT_4_14), .Q(n12287) );
  AND2X1 U12315 ( .IN1(n1230), .IN2(n10017), .Q(n12286) );
  INVX0 U12316 ( .INP(n12288), .ZN(n1230) );
  OR2X1 U12317 ( .IN1(n10643), .IN2(n3893), .Q(n12288) );
  OR2X1 U12318 ( .IN1(n12289), .IN2(n12290), .Q(n12284) );
  AND2X1 U12319 ( .IN1(n9977), .IN2(n12291), .Q(n12290) );
  AND2X1 U12320 ( .IN1(n10073), .IN2(n11531), .Q(n12289) );
  OR2X1 U12321 ( .IN1(n12292), .IN2(n12293), .Q(n11531) );
  INVX0 U12322 ( .INP(n12294), .ZN(n12293) );
  OR2X1 U12323 ( .IN1(n12295), .IN2(n12296), .Q(n12294) );
  AND2X1 U12324 ( .IN1(n12296), .IN2(n12295), .Q(n12292) );
  AND2X1 U12325 ( .IN1(n12297), .IN2(n12298), .Q(n12295) );
  OR2X1 U12326 ( .IN1(WX8501), .IN2(n9358), .Q(n12298) );
  OR2X1 U12327 ( .IN1(WX8437), .IN2(n3623), .Q(n12297) );
  OR2X1 U12328 ( .IN1(n12299), .IN2(n12300), .Q(n12296) );
  AND2X1 U12329 ( .IN1(n9359), .IN2(WX8629), .Q(n12300) );
  AND2X1 U12330 ( .IN1(n9608), .IN2(WX8565), .Q(n12299) );
  OR2X1 U12331 ( .IN1(n12301), .IN2(n12302), .Q(WX7141) );
  OR2X1 U12332 ( .IN1(n12303), .IN2(n12304), .Q(n12302) );
  AND2X1 U12333 ( .IN1(n10043), .IN2(CRC_OUT_4_15), .Q(n12304) );
  AND2X1 U12334 ( .IN1(n1229), .IN2(n10018), .Q(n12303) );
  INVX0 U12335 ( .INP(n12305), .ZN(n1229) );
  OR2X1 U12336 ( .IN1(n10643), .IN2(n3894), .Q(n12305) );
  OR2X1 U12337 ( .IN1(n12306), .IN2(n12307), .Q(n12301) );
  AND2X1 U12338 ( .IN1(n9977), .IN2(n12308), .Q(n12307) );
  AND2X1 U12339 ( .IN1(n11549), .IN2(n10058), .Q(n12306) );
  AND2X1 U12340 ( .IN1(n12309), .IN2(n12310), .Q(n11549) );
  INVX0 U12341 ( .INP(n12311), .ZN(n12310) );
  AND2X1 U12342 ( .IN1(n12312), .IN2(n12313), .Q(n12311) );
  OR2X1 U12343 ( .IN1(n12313), .IN2(n12312), .Q(n12309) );
  OR2X1 U12344 ( .IN1(n12314), .IN2(n12315), .Q(n12312) );
  AND2X1 U12345 ( .IN1(n3625), .IN2(WX8563), .Q(n12315) );
  INVX0 U12346 ( .INP(n12316), .ZN(n12314) );
  OR2X1 U12347 ( .IN1(WX8563), .IN2(n3625), .Q(n12316) );
  AND2X1 U12348 ( .IN1(n12317), .IN2(n12318), .Q(n12313) );
  OR2X1 U12349 ( .IN1(WX8627), .IN2(test_so69), .Q(n12318) );
  OR2X1 U12350 ( .IN1(n9919), .IN2(n9607), .Q(n12317) );
  OR2X1 U12351 ( .IN1(n12319), .IN2(n12320), .Q(WX7139) );
  OR2X1 U12352 ( .IN1(n12321), .IN2(n12322), .Q(n12320) );
  AND2X1 U12353 ( .IN1(n10043), .IN2(CRC_OUT_4_16), .Q(n12322) );
  AND2X1 U12354 ( .IN1(n1228), .IN2(n10018), .Q(n12321) );
  INVX0 U12355 ( .INP(n12323), .ZN(n1228) );
  OR2X1 U12356 ( .IN1(n10643), .IN2(n3895), .Q(n12323) );
  OR2X1 U12357 ( .IN1(n12324), .IN2(n12325), .Q(n12319) );
  AND2X1 U12358 ( .IN1(n9977), .IN2(n12326), .Q(n12325) );
  AND2X1 U12359 ( .IN1(n10073), .IN2(n11566), .Q(n12324) );
  OR2X1 U12360 ( .IN1(n12327), .IN2(n12328), .Q(n11566) );
  INVX0 U12361 ( .INP(n12329), .ZN(n12328) );
  OR2X1 U12362 ( .IN1(n12330), .IN2(n12331), .Q(n12329) );
  AND2X1 U12363 ( .IN1(n12331), .IN2(n12330), .Q(n12327) );
  INVX0 U12364 ( .INP(n12332), .ZN(n12330) );
  OR2X1 U12365 ( .IN1(n12333), .IN2(n12334), .Q(n12332) );
  AND2X1 U12366 ( .IN1(n10519), .IN2(n8363), .Q(n12334) );
  AND2X1 U12367 ( .IN1(n17896), .IN2(n10544), .Q(n12333) );
  OR2X1 U12368 ( .IN1(n12335), .IN2(n12336), .Q(n12331) );
  AND2X1 U12369 ( .IN1(n9518), .IN2(n12337), .Q(n12336) );
  AND2X1 U12370 ( .IN1(n12338), .IN2(n12339), .Q(n12337) );
  OR2X1 U12371 ( .IN1(n9100), .IN2(WX8561), .Q(n12339) );
  OR2X1 U12372 ( .IN1(n9101), .IN2(WX8497), .Q(n12338) );
  AND2X1 U12373 ( .IN1(n12340), .IN2(WX8625), .Q(n12335) );
  OR2X1 U12374 ( .IN1(n12341), .IN2(n12342), .Q(n12340) );
  AND2X1 U12375 ( .IN1(n9100), .IN2(WX8561), .Q(n12342) );
  AND2X1 U12376 ( .IN1(n9101), .IN2(WX8497), .Q(n12341) );
  OR2X1 U12377 ( .IN1(n12343), .IN2(n12344), .Q(WX7137) );
  OR2X1 U12378 ( .IN1(n12345), .IN2(n12346), .Q(n12344) );
  AND2X1 U12379 ( .IN1(n10043), .IN2(CRC_OUT_4_17), .Q(n12346) );
  AND2X1 U12380 ( .IN1(n1227), .IN2(n10018), .Q(n12345) );
  INVX0 U12381 ( .INP(n12347), .ZN(n1227) );
  OR2X1 U12382 ( .IN1(n10643), .IN2(n3896), .Q(n12347) );
  OR2X1 U12383 ( .IN1(n12348), .IN2(n12349), .Q(n12343) );
  AND2X1 U12384 ( .IN1(n9977), .IN2(n12350), .Q(n12349) );
  AND2X1 U12385 ( .IN1(n10073), .IN2(n11587), .Q(n12348) );
  OR2X1 U12386 ( .IN1(n12351), .IN2(n12352), .Q(n11587) );
  INVX0 U12387 ( .INP(n12353), .ZN(n12352) );
  OR2X1 U12388 ( .IN1(n12354), .IN2(n12355), .Q(n12353) );
  AND2X1 U12389 ( .IN1(n12355), .IN2(n12354), .Q(n12351) );
  INVX0 U12390 ( .INP(n12356), .ZN(n12354) );
  OR2X1 U12391 ( .IN1(n12357), .IN2(n12358), .Q(n12356) );
  AND2X1 U12392 ( .IN1(n10519), .IN2(n8364), .Q(n12358) );
  AND2X1 U12393 ( .IN1(n17897), .IN2(n10544), .Q(n12357) );
  OR2X1 U12394 ( .IN1(n12359), .IN2(n12360), .Q(n12355) );
  AND2X1 U12395 ( .IN1(n9606), .IN2(n12361), .Q(n12360) );
  AND2X1 U12396 ( .IN1(n12362), .IN2(n12363), .Q(n12361) );
  OR2X1 U12397 ( .IN1(n9102), .IN2(WX8559), .Q(n12363) );
  OR2X1 U12398 ( .IN1(n9103), .IN2(WX8495), .Q(n12362) );
  AND2X1 U12399 ( .IN1(n12364), .IN2(WX8623), .Q(n12359) );
  OR2X1 U12400 ( .IN1(n12365), .IN2(n12366), .Q(n12364) );
  AND2X1 U12401 ( .IN1(n9102), .IN2(WX8559), .Q(n12366) );
  AND2X1 U12402 ( .IN1(n9103), .IN2(WX8495), .Q(n12365) );
  OR2X1 U12403 ( .IN1(n12367), .IN2(n12368), .Q(WX7135) );
  OR2X1 U12404 ( .IN1(n12369), .IN2(n12370), .Q(n12368) );
  AND2X1 U12405 ( .IN1(n10043), .IN2(CRC_OUT_4_18), .Q(n12370) );
  AND2X1 U12406 ( .IN1(n1226), .IN2(n10018), .Q(n12369) );
  INVX0 U12407 ( .INP(n12371), .ZN(n1226) );
  OR2X1 U12408 ( .IN1(n10642), .IN2(n3897), .Q(n12371) );
  OR2X1 U12409 ( .IN1(n12372), .IN2(n12373), .Q(n12367) );
  AND2X1 U12410 ( .IN1(n9977), .IN2(n12374), .Q(n12373) );
  AND2X1 U12411 ( .IN1(n10073), .IN2(n11611), .Q(n12372) );
  OR2X1 U12412 ( .IN1(n12375), .IN2(n12376), .Q(n11611) );
  INVX0 U12413 ( .INP(n12377), .ZN(n12376) );
  OR2X1 U12414 ( .IN1(n12378), .IN2(n12379), .Q(n12377) );
  AND2X1 U12415 ( .IN1(n12379), .IN2(n12378), .Q(n12375) );
  INVX0 U12416 ( .INP(n12380), .ZN(n12378) );
  OR2X1 U12417 ( .IN1(n12381), .IN2(n12382), .Q(n12380) );
  AND2X1 U12418 ( .IN1(n10519), .IN2(n8365), .Q(n12382) );
  AND2X1 U12419 ( .IN1(n17898), .IN2(n10544), .Q(n12381) );
  OR2X1 U12420 ( .IN1(n12383), .IN2(n12384), .Q(n12379) );
  AND2X1 U12421 ( .IN1(n9605), .IN2(n12385), .Q(n12384) );
  AND2X1 U12422 ( .IN1(n12386), .IN2(n12387), .Q(n12385) );
  OR2X1 U12423 ( .IN1(n9104), .IN2(WX8557), .Q(n12387) );
  OR2X1 U12424 ( .IN1(n9105), .IN2(WX8493), .Q(n12386) );
  AND2X1 U12425 ( .IN1(n12388), .IN2(WX8621), .Q(n12383) );
  OR2X1 U12426 ( .IN1(n12389), .IN2(n12390), .Q(n12388) );
  AND2X1 U12427 ( .IN1(n9104), .IN2(WX8557), .Q(n12390) );
  AND2X1 U12428 ( .IN1(n9105), .IN2(WX8493), .Q(n12389) );
  OR2X1 U12429 ( .IN1(n12391), .IN2(n12392), .Q(WX7133) );
  OR2X1 U12430 ( .IN1(n12393), .IN2(n12394), .Q(n12392) );
  AND2X1 U12431 ( .IN1(n10043), .IN2(CRC_OUT_4_19), .Q(n12394) );
  AND2X1 U12432 ( .IN1(n1225), .IN2(n10018), .Q(n12393) );
  INVX0 U12433 ( .INP(n12395), .ZN(n1225) );
  OR2X1 U12434 ( .IN1(n10642), .IN2(n3898), .Q(n12395) );
  OR2X1 U12435 ( .IN1(n12396), .IN2(n12397), .Q(n12391) );
  AND2X1 U12436 ( .IN1(n9978), .IN2(n12398), .Q(n12397) );
  AND2X1 U12437 ( .IN1(n10074), .IN2(n11632), .Q(n12396) );
  OR2X1 U12438 ( .IN1(n12399), .IN2(n12400), .Q(n11632) );
  INVX0 U12439 ( .INP(n12401), .ZN(n12400) );
  OR2X1 U12440 ( .IN1(n12402), .IN2(n12403), .Q(n12401) );
  AND2X1 U12441 ( .IN1(n12403), .IN2(n12402), .Q(n12399) );
  INVX0 U12442 ( .INP(n12404), .ZN(n12402) );
  OR2X1 U12443 ( .IN1(n12405), .IN2(n12406), .Q(n12404) );
  AND2X1 U12444 ( .IN1(n10519), .IN2(n8366), .Q(n12406) );
  AND2X1 U12445 ( .IN1(n17899), .IN2(n10544), .Q(n12405) );
  OR2X1 U12446 ( .IN1(n12407), .IN2(n12408), .Q(n12403) );
  AND2X1 U12447 ( .IN1(n9604), .IN2(n12409), .Q(n12408) );
  AND2X1 U12448 ( .IN1(n12410), .IN2(n12411), .Q(n12409) );
  OR2X1 U12449 ( .IN1(n9106), .IN2(WX8555), .Q(n12411) );
  OR2X1 U12450 ( .IN1(n9107), .IN2(WX8491), .Q(n12410) );
  AND2X1 U12451 ( .IN1(n12412), .IN2(WX8619), .Q(n12407) );
  OR2X1 U12452 ( .IN1(n12413), .IN2(n12414), .Q(n12412) );
  AND2X1 U12453 ( .IN1(n9106), .IN2(WX8555), .Q(n12414) );
  AND2X1 U12454 ( .IN1(n9107), .IN2(WX8491), .Q(n12413) );
  OR2X1 U12455 ( .IN1(n12415), .IN2(n12416), .Q(WX7131) );
  OR2X1 U12456 ( .IN1(n12417), .IN2(n12418), .Q(n12416) );
  AND2X1 U12457 ( .IN1(n10043), .IN2(CRC_OUT_4_20), .Q(n12418) );
  AND2X1 U12458 ( .IN1(n1224), .IN2(n10018), .Q(n12417) );
  INVX0 U12459 ( .INP(n12419), .ZN(n1224) );
  OR2X1 U12460 ( .IN1(n10642), .IN2(n3899), .Q(n12419) );
  OR2X1 U12461 ( .IN1(n12420), .IN2(n12421), .Q(n12415) );
  AND2X1 U12462 ( .IN1(n9977), .IN2(n12422), .Q(n12421) );
  AND2X1 U12463 ( .IN1(n10074), .IN2(n11656), .Q(n12420) );
  OR2X1 U12464 ( .IN1(n12423), .IN2(n12424), .Q(n11656) );
  INVX0 U12465 ( .INP(n12425), .ZN(n12424) );
  OR2X1 U12466 ( .IN1(n12426), .IN2(n12427), .Q(n12425) );
  AND2X1 U12467 ( .IN1(n12427), .IN2(n12426), .Q(n12423) );
  INVX0 U12468 ( .INP(n12428), .ZN(n12426) );
  OR2X1 U12469 ( .IN1(n12429), .IN2(n12430), .Q(n12428) );
  AND2X1 U12470 ( .IN1(n10519), .IN2(n8367), .Q(n12430) );
  AND2X1 U12471 ( .IN1(n17900), .IN2(n10544), .Q(n12429) );
  OR2X1 U12472 ( .IN1(n12431), .IN2(n12432), .Q(n12427) );
  AND2X1 U12473 ( .IN1(n9603), .IN2(n12433), .Q(n12432) );
  AND2X1 U12474 ( .IN1(n12434), .IN2(n12435), .Q(n12433) );
  OR2X1 U12475 ( .IN1(n9108), .IN2(WX8553), .Q(n12435) );
  OR2X1 U12476 ( .IN1(n9109), .IN2(WX8489), .Q(n12434) );
  AND2X1 U12477 ( .IN1(n12436), .IN2(WX8617), .Q(n12431) );
  OR2X1 U12478 ( .IN1(n12437), .IN2(n12438), .Q(n12436) );
  AND2X1 U12479 ( .IN1(n9108), .IN2(WX8553), .Q(n12438) );
  AND2X1 U12480 ( .IN1(n9109), .IN2(WX8489), .Q(n12437) );
  OR2X1 U12481 ( .IN1(n12439), .IN2(n12440), .Q(WX7129) );
  OR2X1 U12482 ( .IN1(n12441), .IN2(n12442), .Q(n12440) );
  AND2X1 U12483 ( .IN1(n10043), .IN2(CRC_OUT_4_21), .Q(n12442) );
  AND2X1 U12484 ( .IN1(n1223), .IN2(n10018), .Q(n12441) );
  INVX0 U12485 ( .INP(n12443), .ZN(n1223) );
  OR2X1 U12486 ( .IN1(n10642), .IN2(n3900), .Q(n12443) );
  OR2X1 U12487 ( .IN1(n12444), .IN2(n12445), .Q(n12439) );
  AND2X1 U12488 ( .IN1(n12446), .IN2(n9975), .Q(n12445) );
  AND2X1 U12489 ( .IN1(n10074), .IN2(n11680), .Q(n12444) );
  OR2X1 U12490 ( .IN1(n12447), .IN2(n12448), .Q(n11680) );
  INVX0 U12491 ( .INP(n12449), .ZN(n12448) );
  OR2X1 U12492 ( .IN1(n12450), .IN2(n12451), .Q(n12449) );
  AND2X1 U12493 ( .IN1(n12451), .IN2(n12450), .Q(n12447) );
  INVX0 U12494 ( .INP(n12452), .ZN(n12450) );
  OR2X1 U12495 ( .IN1(n12453), .IN2(n12454), .Q(n12452) );
  AND2X1 U12496 ( .IN1(n10519), .IN2(n8368), .Q(n12454) );
  AND2X1 U12497 ( .IN1(n17901), .IN2(n10544), .Q(n12453) );
  OR2X1 U12498 ( .IN1(n12455), .IN2(n12456), .Q(n12451) );
  AND2X1 U12499 ( .IN1(n9602), .IN2(n12457), .Q(n12456) );
  AND2X1 U12500 ( .IN1(n12458), .IN2(n12459), .Q(n12457) );
  OR2X1 U12501 ( .IN1(n9110), .IN2(WX8551), .Q(n12459) );
  OR2X1 U12502 ( .IN1(n9111), .IN2(WX8487), .Q(n12458) );
  AND2X1 U12503 ( .IN1(n12460), .IN2(WX8615), .Q(n12455) );
  OR2X1 U12504 ( .IN1(n12461), .IN2(n12462), .Q(n12460) );
  AND2X1 U12505 ( .IN1(n9110), .IN2(WX8551), .Q(n12462) );
  AND2X1 U12506 ( .IN1(n9111), .IN2(WX8487), .Q(n12461) );
  OR2X1 U12507 ( .IN1(n12463), .IN2(n12464), .Q(WX7127) );
  OR2X1 U12508 ( .IN1(n12465), .IN2(n12466), .Q(n12464) );
  AND2X1 U12509 ( .IN1(n10043), .IN2(CRC_OUT_4_22), .Q(n12466) );
  AND2X1 U12510 ( .IN1(n1222), .IN2(n10018), .Q(n12465) );
  INVX0 U12511 ( .INP(n12467), .ZN(n1222) );
  OR2X1 U12512 ( .IN1(n10642), .IN2(n3901), .Q(n12467) );
  OR2X1 U12513 ( .IN1(n12468), .IN2(n12469), .Q(n12463) );
  AND2X1 U12514 ( .IN1(n9977), .IN2(n12470), .Q(n12469) );
  AND2X1 U12515 ( .IN1(n10074), .IN2(n11704), .Q(n12468) );
  OR2X1 U12516 ( .IN1(n12471), .IN2(n12472), .Q(n11704) );
  INVX0 U12517 ( .INP(n12473), .ZN(n12472) );
  OR2X1 U12518 ( .IN1(n12474), .IN2(n12475), .Q(n12473) );
  AND2X1 U12519 ( .IN1(n12475), .IN2(n12474), .Q(n12471) );
  INVX0 U12520 ( .INP(n12476), .ZN(n12474) );
  OR2X1 U12521 ( .IN1(n12477), .IN2(n12478), .Q(n12476) );
  AND2X1 U12522 ( .IN1(n10519), .IN2(n8369), .Q(n12478) );
  AND2X1 U12523 ( .IN1(n17902), .IN2(n10544), .Q(n12477) );
  OR2X1 U12524 ( .IN1(n12479), .IN2(n12480), .Q(n12475) );
  AND2X1 U12525 ( .IN1(n9601), .IN2(n12481), .Q(n12480) );
  AND2X1 U12526 ( .IN1(n12482), .IN2(n12483), .Q(n12481) );
  OR2X1 U12527 ( .IN1(n9112), .IN2(WX8549), .Q(n12483) );
  OR2X1 U12528 ( .IN1(n9113), .IN2(WX8485), .Q(n12482) );
  AND2X1 U12529 ( .IN1(n12484), .IN2(WX8613), .Q(n12479) );
  OR2X1 U12530 ( .IN1(n12485), .IN2(n12486), .Q(n12484) );
  AND2X1 U12531 ( .IN1(n9112), .IN2(WX8549), .Q(n12486) );
  AND2X1 U12532 ( .IN1(n9113), .IN2(WX8485), .Q(n12485) );
  OR2X1 U12533 ( .IN1(n12487), .IN2(n12488), .Q(WX7125) );
  OR2X1 U12534 ( .IN1(n12489), .IN2(n12490), .Q(n12488) );
  AND2X1 U12535 ( .IN1(n10043), .IN2(CRC_OUT_4_23), .Q(n12490) );
  AND2X1 U12536 ( .IN1(n1221), .IN2(n10018), .Q(n12489) );
  INVX0 U12537 ( .INP(n12491), .ZN(n1221) );
  OR2X1 U12538 ( .IN1(n10642), .IN2(n3902), .Q(n12491) );
  OR2X1 U12539 ( .IN1(n12492), .IN2(n12493), .Q(n12487) );
  AND2X1 U12540 ( .IN1(n12494), .IN2(n9976), .Q(n12493) );
  AND2X1 U12541 ( .IN1(n10074), .IN2(n11728), .Q(n12492) );
  OR2X1 U12542 ( .IN1(n12495), .IN2(n12496), .Q(n11728) );
  INVX0 U12543 ( .INP(n12497), .ZN(n12496) );
  OR2X1 U12544 ( .IN1(n12498), .IN2(n12499), .Q(n12497) );
  AND2X1 U12545 ( .IN1(n12499), .IN2(n12498), .Q(n12495) );
  INVX0 U12546 ( .INP(n12500), .ZN(n12498) );
  OR2X1 U12547 ( .IN1(n12501), .IN2(n12502), .Q(n12500) );
  AND2X1 U12548 ( .IN1(n10520), .IN2(n8370), .Q(n12502) );
  AND2X1 U12549 ( .IN1(n17903), .IN2(n10544), .Q(n12501) );
  OR2X1 U12550 ( .IN1(n12503), .IN2(n12504), .Q(n12499) );
  AND2X1 U12551 ( .IN1(n9600), .IN2(n12505), .Q(n12504) );
  AND2X1 U12552 ( .IN1(n12506), .IN2(n12507), .Q(n12505) );
  OR2X1 U12553 ( .IN1(n9114), .IN2(WX8547), .Q(n12507) );
  OR2X1 U12554 ( .IN1(n9115), .IN2(WX8483), .Q(n12506) );
  AND2X1 U12555 ( .IN1(n12508), .IN2(WX8611), .Q(n12503) );
  OR2X1 U12556 ( .IN1(n12509), .IN2(n12510), .Q(n12508) );
  AND2X1 U12557 ( .IN1(n9114), .IN2(WX8547), .Q(n12510) );
  AND2X1 U12558 ( .IN1(n9115), .IN2(WX8483), .Q(n12509) );
  OR2X1 U12559 ( .IN1(n12511), .IN2(n12512), .Q(WX7123) );
  OR2X1 U12560 ( .IN1(n12513), .IN2(n12514), .Q(n12512) );
  AND2X1 U12561 ( .IN1(n10043), .IN2(CRC_OUT_4_24), .Q(n12514) );
  AND2X1 U12562 ( .IN1(n1220), .IN2(n10018), .Q(n12513) );
  INVX0 U12563 ( .INP(n12515), .ZN(n1220) );
  OR2X1 U12564 ( .IN1(n10642), .IN2(n3903), .Q(n12515) );
  OR2X1 U12565 ( .IN1(n12516), .IN2(n12517), .Q(n12511) );
  AND2X1 U12566 ( .IN1(n9977), .IN2(n12518), .Q(n12517) );
  AND2X1 U12567 ( .IN1(n10074), .IN2(n11752), .Q(n12516) );
  OR2X1 U12568 ( .IN1(n12519), .IN2(n12520), .Q(n11752) );
  INVX0 U12569 ( .INP(n12521), .ZN(n12520) );
  OR2X1 U12570 ( .IN1(n12522), .IN2(n12523), .Q(n12521) );
  AND2X1 U12571 ( .IN1(n12523), .IN2(n12522), .Q(n12519) );
  INVX0 U12572 ( .INP(n12524), .ZN(n12522) );
  OR2X1 U12573 ( .IN1(n12525), .IN2(n12526), .Q(n12524) );
  AND2X1 U12574 ( .IN1(n10520), .IN2(n8371), .Q(n12526) );
  AND2X1 U12575 ( .IN1(n17904), .IN2(n10544), .Q(n12525) );
  OR2X1 U12576 ( .IN1(n12527), .IN2(n12528), .Q(n12523) );
  AND2X1 U12577 ( .IN1(n9599), .IN2(n12529), .Q(n12528) );
  AND2X1 U12578 ( .IN1(n12530), .IN2(n12531), .Q(n12529) );
  OR2X1 U12579 ( .IN1(n9116), .IN2(WX8545), .Q(n12531) );
  OR2X1 U12580 ( .IN1(n9117), .IN2(WX8481), .Q(n12530) );
  AND2X1 U12581 ( .IN1(n12532), .IN2(WX8609), .Q(n12527) );
  OR2X1 U12582 ( .IN1(n12533), .IN2(n12534), .Q(n12532) );
  AND2X1 U12583 ( .IN1(n9116), .IN2(WX8545), .Q(n12534) );
  AND2X1 U12584 ( .IN1(n9117), .IN2(WX8481), .Q(n12533) );
  OR2X1 U12585 ( .IN1(n12535), .IN2(n12536), .Q(WX7121) );
  OR2X1 U12586 ( .IN1(n12537), .IN2(n12538), .Q(n12536) );
  AND2X1 U12587 ( .IN1(n10044), .IN2(CRC_OUT_4_25), .Q(n12538) );
  AND2X1 U12588 ( .IN1(n1219), .IN2(n10018), .Q(n12537) );
  INVX0 U12589 ( .INP(n12539), .ZN(n1219) );
  OR2X1 U12590 ( .IN1(n10642), .IN2(n3904), .Q(n12539) );
  OR2X1 U12591 ( .IN1(n12540), .IN2(n12541), .Q(n12535) );
  AND2X1 U12592 ( .IN1(n12542), .IN2(n9976), .Q(n12541) );
  AND2X1 U12593 ( .IN1(n10074), .IN2(n11776), .Q(n12540) );
  OR2X1 U12594 ( .IN1(n12543), .IN2(n12544), .Q(n11776) );
  INVX0 U12595 ( .INP(n12545), .ZN(n12544) );
  OR2X1 U12596 ( .IN1(n12546), .IN2(n12547), .Q(n12545) );
  AND2X1 U12597 ( .IN1(n12547), .IN2(n12546), .Q(n12543) );
  INVX0 U12598 ( .INP(n12548), .ZN(n12546) );
  OR2X1 U12599 ( .IN1(n12549), .IN2(n12550), .Q(n12548) );
  AND2X1 U12600 ( .IN1(n10520), .IN2(n8372), .Q(n12550) );
  AND2X1 U12601 ( .IN1(n17905), .IN2(n10544), .Q(n12549) );
  OR2X1 U12602 ( .IN1(n12551), .IN2(n12552), .Q(n12547) );
  AND2X1 U12603 ( .IN1(n9598), .IN2(n12553), .Q(n12552) );
  AND2X1 U12604 ( .IN1(n12554), .IN2(n12555), .Q(n12553) );
  OR2X1 U12605 ( .IN1(n9118), .IN2(WX8543), .Q(n12555) );
  OR2X1 U12606 ( .IN1(n9119), .IN2(WX8479), .Q(n12554) );
  AND2X1 U12607 ( .IN1(n12556), .IN2(WX8607), .Q(n12551) );
  OR2X1 U12608 ( .IN1(n12557), .IN2(n12558), .Q(n12556) );
  AND2X1 U12609 ( .IN1(n9118), .IN2(WX8543), .Q(n12558) );
  AND2X1 U12610 ( .IN1(n9119), .IN2(WX8479), .Q(n12557) );
  OR2X1 U12611 ( .IN1(n12559), .IN2(n12560), .Q(WX7119) );
  OR2X1 U12612 ( .IN1(n12561), .IN2(n12562), .Q(n12560) );
  AND2X1 U12613 ( .IN1(n10044), .IN2(CRC_OUT_4_26), .Q(n12562) );
  AND2X1 U12614 ( .IN1(n1218), .IN2(n10018), .Q(n12561) );
  INVX0 U12615 ( .INP(n12563), .ZN(n1218) );
  OR2X1 U12616 ( .IN1(n10642), .IN2(n3905), .Q(n12563) );
  OR2X1 U12617 ( .IN1(n12564), .IN2(n12565), .Q(n12559) );
  AND2X1 U12618 ( .IN1(n9978), .IN2(n12566), .Q(n12565) );
  AND2X1 U12619 ( .IN1(n11800), .IN2(n10058), .Q(n12564) );
  AND2X1 U12620 ( .IN1(n12567), .IN2(n12568), .Q(n11800) );
  INVX0 U12621 ( .INP(n12569), .ZN(n12568) );
  AND2X1 U12622 ( .IN1(n12570), .IN2(n12571), .Q(n12569) );
  OR2X1 U12623 ( .IN1(n12571), .IN2(n12570), .Q(n12567) );
  OR2X1 U12624 ( .IN1(n12572), .IN2(n12573), .Q(n12570) );
  AND2X1 U12625 ( .IN1(n10520), .IN2(WX8477), .Q(n12573) );
  AND2X1 U12626 ( .IN1(n9120), .IN2(n10543), .Q(n12572) );
  AND2X1 U12627 ( .IN1(n12574), .IN2(n12575), .Q(n12571) );
  INVX0 U12628 ( .INP(n12576), .ZN(n12575) );
  AND2X1 U12629 ( .IN1(n12577), .IN2(WX8541), .Q(n12576) );
  OR2X1 U12630 ( .IN1(WX8541), .IN2(n12577), .Q(n12574) );
  OR2X1 U12631 ( .IN1(n12578), .IN2(n12579), .Q(n12577) );
  AND2X1 U12632 ( .IN1(n17906), .IN2(n9908), .Q(n12579) );
  AND2X1 U12633 ( .IN1(test_so74), .IN2(n8373), .Q(n12578) );
  OR2X1 U12634 ( .IN1(n12580), .IN2(n12581), .Q(WX7117) );
  OR2X1 U12635 ( .IN1(n12582), .IN2(n12583), .Q(n12581) );
  AND2X1 U12636 ( .IN1(n10044), .IN2(CRC_OUT_4_27), .Q(n12583) );
  AND2X1 U12637 ( .IN1(n1217), .IN2(n10019), .Q(n12582) );
  INVX0 U12638 ( .INP(n12584), .ZN(n1217) );
  OR2X1 U12639 ( .IN1(n10642), .IN2(n3906), .Q(n12584) );
  OR2X1 U12640 ( .IN1(n12585), .IN2(n12586), .Q(n12580) );
  AND2X1 U12641 ( .IN1(n12587), .IN2(n9977), .Q(n12586) );
  AND2X1 U12642 ( .IN1(n10074), .IN2(n11824), .Q(n12585) );
  OR2X1 U12643 ( .IN1(n12588), .IN2(n12589), .Q(n11824) );
  INVX0 U12644 ( .INP(n12590), .ZN(n12589) );
  OR2X1 U12645 ( .IN1(n12591), .IN2(n12592), .Q(n12590) );
  AND2X1 U12646 ( .IN1(n12592), .IN2(n12591), .Q(n12588) );
  INVX0 U12647 ( .INP(n12593), .ZN(n12591) );
  OR2X1 U12648 ( .IN1(n12594), .IN2(n12595), .Q(n12593) );
  AND2X1 U12649 ( .IN1(n10520), .IN2(n8374), .Q(n12595) );
  AND2X1 U12650 ( .IN1(n17907), .IN2(n10543), .Q(n12594) );
  OR2X1 U12651 ( .IN1(n12596), .IN2(n12597), .Q(n12592) );
  AND2X1 U12652 ( .IN1(n9597), .IN2(n12598), .Q(n12597) );
  AND2X1 U12653 ( .IN1(n12599), .IN2(n12600), .Q(n12598) );
  OR2X1 U12654 ( .IN1(n9122), .IN2(WX8539), .Q(n12600) );
  OR2X1 U12655 ( .IN1(n9123), .IN2(WX8475), .Q(n12599) );
  AND2X1 U12656 ( .IN1(n12601), .IN2(WX8603), .Q(n12596) );
  OR2X1 U12657 ( .IN1(n12602), .IN2(n12603), .Q(n12601) );
  AND2X1 U12658 ( .IN1(n9122), .IN2(WX8539), .Q(n12603) );
  AND2X1 U12659 ( .IN1(n9123), .IN2(WX8475), .Q(n12602) );
  OR2X1 U12660 ( .IN1(n12604), .IN2(n12605), .Q(WX7115) );
  OR2X1 U12661 ( .IN1(n12606), .IN2(n12607), .Q(n12605) );
  AND2X1 U12662 ( .IN1(n10044), .IN2(CRC_OUT_4_28), .Q(n12607) );
  AND2X1 U12663 ( .IN1(n1216), .IN2(n10019), .Q(n12606) );
  INVX0 U12664 ( .INP(n12608), .ZN(n1216) );
  OR2X1 U12665 ( .IN1(n10642), .IN2(n3907), .Q(n12608) );
  OR2X1 U12666 ( .IN1(n12609), .IN2(n12610), .Q(n12604) );
  AND2X1 U12667 ( .IN1(n9978), .IN2(n12611), .Q(n12610) );
  AND2X1 U12668 ( .IN1(n11848), .IN2(n10058), .Q(n12609) );
  AND2X1 U12669 ( .IN1(n12612), .IN2(n12613), .Q(n11848) );
  INVX0 U12670 ( .INP(n12614), .ZN(n12613) );
  AND2X1 U12671 ( .IN1(n12615), .IN2(n12616), .Q(n12614) );
  OR2X1 U12672 ( .IN1(n12616), .IN2(n12615), .Q(n12612) );
  OR2X1 U12673 ( .IN1(n12617), .IN2(n12618), .Q(n12615) );
  AND2X1 U12674 ( .IN1(n10520), .IN2(WX8473), .Q(n12618) );
  AND2X1 U12675 ( .IN1(n9124), .IN2(n10543), .Q(n12617) );
  AND2X1 U12676 ( .IN1(n12619), .IN2(n12620), .Q(n12616) );
  OR2X1 U12677 ( .IN1(n12621), .IN2(n9596), .Q(n12620) );
  INVX0 U12678 ( .INP(n12622), .ZN(n12621) );
  OR2X1 U12679 ( .IN1(WX8601), .IN2(n12622), .Q(n12619) );
  OR2X1 U12680 ( .IN1(n12623), .IN2(n12624), .Q(n12622) );
  AND2X1 U12681 ( .IN1(n17908), .IN2(n9955), .Q(n12624) );
  AND2X1 U12682 ( .IN1(test_so72), .IN2(n8375), .Q(n12623) );
  OR2X1 U12683 ( .IN1(n12625), .IN2(n12626), .Q(WX7113) );
  OR2X1 U12684 ( .IN1(n12627), .IN2(n12628), .Q(n12626) );
  AND2X1 U12685 ( .IN1(test_so66), .IN2(n10026), .Q(n12628) );
  AND2X1 U12686 ( .IN1(n1215), .IN2(n10019), .Q(n12627) );
  INVX0 U12687 ( .INP(n12629), .ZN(n1215) );
  OR2X1 U12688 ( .IN1(n10642), .IN2(n3908), .Q(n12629) );
  OR2X1 U12689 ( .IN1(n12630), .IN2(n12631), .Q(n12625) );
  AND2X1 U12690 ( .IN1(n9978), .IN2(n12632), .Q(n12631) );
  AND2X1 U12691 ( .IN1(n10074), .IN2(n11872), .Q(n12630) );
  OR2X1 U12692 ( .IN1(n12633), .IN2(n12634), .Q(n11872) );
  INVX0 U12693 ( .INP(n12635), .ZN(n12634) );
  OR2X1 U12694 ( .IN1(n12636), .IN2(n12637), .Q(n12635) );
  AND2X1 U12695 ( .IN1(n12637), .IN2(n12636), .Q(n12633) );
  INVX0 U12696 ( .INP(n12638), .ZN(n12636) );
  OR2X1 U12697 ( .IN1(n12639), .IN2(n12640), .Q(n12638) );
  AND2X1 U12698 ( .IN1(n10523), .IN2(n8376), .Q(n12640) );
  AND2X1 U12699 ( .IN1(n17909), .IN2(n10543), .Q(n12639) );
  OR2X1 U12700 ( .IN1(n12641), .IN2(n12642), .Q(n12637) );
  AND2X1 U12701 ( .IN1(n9595), .IN2(n12643), .Q(n12642) );
  AND2X1 U12702 ( .IN1(n12644), .IN2(n12645), .Q(n12643) );
  OR2X1 U12703 ( .IN1(n9125), .IN2(WX8535), .Q(n12645) );
  OR2X1 U12704 ( .IN1(n9126), .IN2(WX8471), .Q(n12644) );
  AND2X1 U12705 ( .IN1(n12646), .IN2(WX8599), .Q(n12641) );
  OR2X1 U12706 ( .IN1(n12647), .IN2(n12648), .Q(n12646) );
  AND2X1 U12707 ( .IN1(n9125), .IN2(WX8535), .Q(n12648) );
  AND2X1 U12708 ( .IN1(n9126), .IN2(WX8471), .Q(n12647) );
  OR2X1 U12709 ( .IN1(n12649), .IN2(n12650), .Q(WX7111) );
  OR2X1 U12710 ( .IN1(n12651), .IN2(n12652), .Q(n12650) );
  AND2X1 U12711 ( .IN1(n10044), .IN2(CRC_OUT_4_30), .Q(n12652) );
  AND2X1 U12712 ( .IN1(n1214), .IN2(n10019), .Q(n12651) );
  INVX0 U12713 ( .INP(n12653), .ZN(n1214) );
  OR2X1 U12714 ( .IN1(n10641), .IN2(n3909), .Q(n12653) );
  OR2X1 U12715 ( .IN1(n12654), .IN2(n12655), .Q(n12649) );
  AND2X1 U12716 ( .IN1(n9978), .IN2(n12656), .Q(n12655) );
  AND2X1 U12717 ( .IN1(n11896), .IN2(n10058), .Q(n12654) );
  AND2X1 U12718 ( .IN1(n12657), .IN2(n12658), .Q(n11896) );
  INVX0 U12719 ( .INP(n12659), .ZN(n12658) );
  AND2X1 U12720 ( .IN1(n12660), .IN2(n12661), .Q(n12659) );
  OR2X1 U12721 ( .IN1(n12661), .IN2(n12660), .Q(n12657) );
  OR2X1 U12722 ( .IN1(n12662), .IN2(n12663), .Q(n12660) );
  AND2X1 U12723 ( .IN1(n10520), .IN2(WX8533), .Q(n12663) );
  AND2X1 U12724 ( .IN1(n9127), .IN2(n10543), .Q(n12662) );
  AND2X1 U12725 ( .IN1(n12664), .IN2(n12665), .Q(n12661) );
  OR2X1 U12726 ( .IN1(n12666), .IN2(n9594), .Q(n12665) );
  INVX0 U12727 ( .INP(n12667), .ZN(n12666) );
  OR2X1 U12728 ( .IN1(WX8597), .IN2(n12667), .Q(n12664) );
  OR2X1 U12729 ( .IN1(n12668), .IN2(n12669), .Q(n12667) );
  AND2X1 U12730 ( .IN1(n17910), .IN2(n9956), .Q(n12669) );
  AND2X1 U12731 ( .IN1(test_so70), .IN2(n8377), .Q(n12668) );
  OR2X1 U12732 ( .IN1(n12670), .IN2(n12671), .Q(WX7109) );
  OR2X1 U12733 ( .IN1(n12672), .IN2(n12673), .Q(n12671) );
  AND2X1 U12734 ( .IN1(n2245), .IN2(WX6950), .Q(n12673) );
  AND2X1 U12735 ( .IN1(n10044), .IN2(CRC_OUT_4_31), .Q(n12672) );
  OR2X1 U12736 ( .IN1(n12674), .IN2(n12675), .Q(n12670) );
  AND2X1 U12737 ( .IN1(n9978), .IN2(n12676), .Q(n12675) );
  AND2X1 U12738 ( .IN1(n10074), .IN2(n11919), .Q(n12674) );
  OR2X1 U12739 ( .IN1(n12677), .IN2(n12678), .Q(n11919) );
  INVX0 U12740 ( .INP(n12679), .ZN(n12678) );
  OR2X1 U12741 ( .IN1(n12680), .IN2(n12681), .Q(n12679) );
  AND2X1 U12742 ( .IN1(n12681), .IN2(n12680), .Q(n12677) );
  INVX0 U12743 ( .INP(n12682), .ZN(n12680) );
  OR2X1 U12744 ( .IN1(n12683), .IN2(n12684), .Q(n12682) );
  AND2X1 U12745 ( .IN1(n10520), .IN2(n8378), .Q(n12684) );
  AND2X1 U12746 ( .IN1(n17911), .IN2(n10543), .Q(n12683) );
  OR2X1 U12747 ( .IN1(n12685), .IN2(n12686), .Q(n12681) );
  AND2X1 U12748 ( .IN1(n9593), .IN2(n12687), .Q(n12686) );
  AND2X1 U12749 ( .IN1(n12688), .IN2(n12689), .Q(n12687) );
  OR2X1 U12750 ( .IN1(n9032), .IN2(WX8531), .Q(n12689) );
  OR2X1 U12751 ( .IN1(n9033), .IN2(WX8467), .Q(n12688) );
  AND2X1 U12752 ( .IN1(n12690), .IN2(WX8595), .Q(n12685) );
  OR2X1 U12753 ( .IN1(n12691), .IN2(n12692), .Q(n12690) );
  AND2X1 U12754 ( .IN1(n9032), .IN2(WX8531), .Q(n12692) );
  AND2X1 U12755 ( .IN1(n9033), .IN2(WX8467), .Q(n12691) );
  OR2X1 U12756 ( .IN1(n12693), .IN2(n12694), .Q(WX706) );
  OR2X1 U12757 ( .IN1(n12695), .IN2(n12696), .Q(n12694) );
  AND2X1 U12758 ( .IN1(n10044), .IN2(CRC_OUT_9_0), .Q(n12696) );
  AND2X1 U12759 ( .IN1(WX544), .IN2(n10019), .Q(n12695) );
  OR2X1 U12760 ( .IN1(n12697), .IN2(n12698), .Q(n12693) );
  AND2X1 U12761 ( .IN1(n9978), .IN2(n12699), .Q(n12698) );
  AND2X1 U12762 ( .IN1(n12700), .IN2(n10058), .Q(n12697) );
  OR2X1 U12763 ( .IN1(n12701), .IN2(n12702), .Q(WX704) );
  OR2X1 U12764 ( .IN1(n12703), .IN2(n12704), .Q(n12702) );
  AND2X1 U12765 ( .IN1(test_so9), .IN2(n10027), .Q(n12704) );
  AND2X1 U12766 ( .IN1(WX542), .IN2(n10019), .Q(n12703) );
  OR2X1 U12767 ( .IN1(n12705), .IN2(n12706), .Q(n12701) );
  AND2X1 U12768 ( .IN1(n9978), .IN2(n12707), .Q(n12706) );
  AND2X1 U12769 ( .IN1(n10074), .IN2(n12708), .Q(n12705) );
  OR2X1 U12770 ( .IN1(n12709), .IN2(n12710), .Q(WX702) );
  OR2X1 U12771 ( .IN1(n12711), .IN2(n12712), .Q(n12710) );
  AND2X1 U12772 ( .IN1(n10044), .IN2(CRC_OUT_9_2), .Q(n12712) );
  AND2X1 U12773 ( .IN1(WX540), .IN2(n10019), .Q(n12711) );
  OR2X1 U12774 ( .IN1(n12713), .IN2(n12714), .Q(n12709) );
  AND2X1 U12775 ( .IN1(n12715), .IN2(n9975), .Q(n12714) );
  AND2X1 U12776 ( .IN1(n10074), .IN2(n12716), .Q(n12713) );
  AND2X1 U12777 ( .IN1(n9848), .IN2(n10559), .Q(WX7011) );
  OR2X1 U12778 ( .IN1(n12717), .IN2(n12718), .Q(WX700) );
  OR2X1 U12779 ( .IN1(n12719), .IN2(n12720), .Q(n12718) );
  AND2X1 U12780 ( .IN1(n10044), .IN2(CRC_OUT_9_3), .Q(n12720) );
  AND2X1 U12781 ( .IN1(WX538), .IN2(n10019), .Q(n12719) );
  OR2X1 U12782 ( .IN1(n12721), .IN2(n12722), .Q(n12717) );
  AND2X1 U12783 ( .IN1(n9978), .IN2(n12723), .Q(n12722) );
  AND2X1 U12784 ( .IN1(n10074), .IN2(n12724), .Q(n12721) );
  OR2X1 U12785 ( .IN1(n12725), .IN2(n12726), .Q(WX698) );
  OR2X1 U12786 ( .IN1(n12727), .IN2(n12728), .Q(n12726) );
  AND2X1 U12787 ( .IN1(n10044), .IN2(CRC_OUT_9_4), .Q(n12728) );
  AND2X1 U12788 ( .IN1(WX536), .IN2(n10019), .Q(n12727) );
  OR2X1 U12789 ( .IN1(n12729), .IN2(n12730), .Q(n12725) );
  AND2X1 U12790 ( .IN1(n9978), .IN2(n12731), .Q(n12730) );
  AND2X1 U12791 ( .IN1(n12732), .IN2(n10058), .Q(n12729) );
  OR2X1 U12792 ( .IN1(n12733), .IN2(n12734), .Q(WX696) );
  OR2X1 U12793 ( .IN1(n12735), .IN2(n12736), .Q(n12734) );
  AND2X1 U12794 ( .IN1(n10044), .IN2(CRC_OUT_9_5), .Q(n12736) );
  AND2X1 U12795 ( .IN1(WX534), .IN2(n10019), .Q(n12735) );
  OR2X1 U12796 ( .IN1(n12737), .IN2(n12738), .Q(n12733) );
  AND2X1 U12797 ( .IN1(n9978), .IN2(n12739), .Q(n12738) );
  AND2X1 U12798 ( .IN1(n10075), .IN2(n12740), .Q(n12737) );
  OR2X1 U12799 ( .IN1(n12741), .IN2(n12742), .Q(WX694) );
  OR2X1 U12800 ( .IN1(n12743), .IN2(n12744), .Q(n12742) );
  AND2X1 U12801 ( .IN1(n10044), .IN2(CRC_OUT_9_6), .Q(n12744) );
  AND2X1 U12802 ( .IN1(WX532), .IN2(n10019), .Q(n12743) );
  OR2X1 U12803 ( .IN1(n12745), .IN2(n12746), .Q(n12741) );
  AND2X1 U12804 ( .IN1(n12747), .IN2(n9975), .Q(n12746) );
  AND2X1 U12805 ( .IN1(n10075), .IN2(n12748), .Q(n12745) );
  OR2X1 U12806 ( .IN1(n12749), .IN2(n12750), .Q(WX692) );
  OR2X1 U12807 ( .IN1(n12751), .IN2(n12752), .Q(n12750) );
  AND2X1 U12808 ( .IN1(n10044), .IN2(CRC_OUT_9_7), .Q(n12752) );
  AND2X1 U12809 ( .IN1(WX530), .IN2(n10019), .Q(n12751) );
  OR2X1 U12810 ( .IN1(n12753), .IN2(n12754), .Q(n12749) );
  AND2X1 U12811 ( .IN1(n9978), .IN2(n12755), .Q(n12754) );
  AND2X1 U12812 ( .IN1(n10075), .IN2(n12756), .Q(n12753) );
  OR2X1 U12813 ( .IN1(n12757), .IN2(n12758), .Q(WX690) );
  OR2X1 U12814 ( .IN1(n12759), .IN2(n12760), .Q(n12758) );
  AND2X1 U12815 ( .IN1(n10045), .IN2(CRC_OUT_9_8), .Q(n12760) );
  AND2X1 U12816 ( .IN1(WX528), .IN2(n10020), .Q(n12759) );
  OR2X1 U12817 ( .IN1(n12761), .IN2(n12762), .Q(n12757) );
  AND2X1 U12818 ( .IN1(n9979), .IN2(n12763), .Q(n12762) );
  AND2X1 U12819 ( .IN1(n10075), .IN2(n12764), .Q(n12761) );
  OR2X1 U12820 ( .IN1(n12765), .IN2(n12766), .Q(WX688) );
  OR2X1 U12821 ( .IN1(n12767), .IN2(n12768), .Q(n12766) );
  AND2X1 U12822 ( .IN1(n10045), .IN2(CRC_OUT_9_9), .Q(n12768) );
  AND2X1 U12823 ( .IN1(WX526), .IN2(n10020), .Q(n12767) );
  OR2X1 U12824 ( .IN1(n12769), .IN2(n12770), .Q(n12765) );
  AND2X1 U12825 ( .IN1(n9979), .IN2(n12771), .Q(n12770) );
  AND2X1 U12826 ( .IN1(n10075), .IN2(n12772), .Q(n12769) );
  OR2X1 U12827 ( .IN1(n12773), .IN2(n12774), .Q(WX686) );
  OR2X1 U12828 ( .IN1(n12775), .IN2(n12776), .Q(n12774) );
  AND2X1 U12829 ( .IN1(n10045), .IN2(CRC_OUT_9_10), .Q(n12776) );
  AND2X1 U12830 ( .IN1(WX524), .IN2(n10020), .Q(n12775) );
  OR2X1 U12831 ( .IN1(n12777), .IN2(n12778), .Q(n12773) );
  AND2X1 U12832 ( .IN1(n12779), .IN2(n9974), .Q(n12778) );
  AND2X1 U12833 ( .IN1(n12780), .IN2(n10057), .Q(n12777) );
  OR2X1 U12834 ( .IN1(n12781), .IN2(n12782), .Q(WX684) );
  OR2X1 U12835 ( .IN1(n12783), .IN2(n12784), .Q(n12782) );
  AND2X1 U12836 ( .IN1(n10045), .IN2(CRC_OUT_9_11), .Q(n12784) );
  AND2X1 U12837 ( .IN1(WX522), .IN2(n10020), .Q(n12783) );
  OR2X1 U12838 ( .IN1(n12785), .IN2(n12786), .Q(n12781) );
  AND2X1 U12839 ( .IN1(n9979), .IN2(n12787), .Q(n12786) );
  AND2X1 U12840 ( .IN1(n10075), .IN2(n12788), .Q(n12785) );
  OR2X1 U12841 ( .IN1(n12789), .IN2(n12790), .Q(WX682) );
  OR2X1 U12842 ( .IN1(n12791), .IN2(n12792), .Q(n12790) );
  AND2X1 U12843 ( .IN1(n10045), .IN2(CRC_OUT_9_12), .Q(n12792) );
  AND2X1 U12844 ( .IN1(WX520), .IN2(n10020), .Q(n12791) );
  OR2X1 U12845 ( .IN1(n12793), .IN2(n12794), .Q(n12789) );
  AND2X1 U12846 ( .IN1(n9979), .IN2(n12795), .Q(n12794) );
  AND2X1 U12847 ( .IN1(n10075), .IN2(n12796), .Q(n12793) );
  OR2X1 U12848 ( .IN1(n12797), .IN2(n12798), .Q(WX680) );
  OR2X1 U12849 ( .IN1(n12799), .IN2(n12800), .Q(n12798) );
  AND2X1 U12850 ( .IN1(n10045), .IN2(CRC_OUT_9_13), .Q(n12800) );
  AND2X1 U12851 ( .IN1(WX518), .IN2(n10020), .Q(n12799) );
  OR2X1 U12852 ( .IN1(n12801), .IN2(n12802), .Q(n12797) );
  AND2X1 U12853 ( .IN1(n9979), .IN2(n12803), .Q(n12802) );
  AND2X1 U12854 ( .IN1(n10075), .IN2(n12804), .Q(n12801) );
  OR2X1 U12855 ( .IN1(n12805), .IN2(n12806), .Q(WX678) );
  OR2X1 U12856 ( .IN1(n12807), .IN2(n12808), .Q(n12806) );
  AND2X1 U12857 ( .IN1(n10045), .IN2(CRC_OUT_9_14), .Q(n12808) );
  AND2X1 U12858 ( .IN1(WX516), .IN2(n10020), .Q(n12807) );
  OR2X1 U12859 ( .IN1(n12809), .IN2(n12810), .Q(n12805) );
  AND2X1 U12860 ( .IN1(n9979), .IN2(n12811), .Q(n12810) );
  AND2X1 U12861 ( .IN1(n12812), .IN2(n10057), .Q(n12809) );
  OR2X1 U12862 ( .IN1(n12813), .IN2(n12814), .Q(WX676) );
  OR2X1 U12863 ( .IN1(n12815), .IN2(n12816), .Q(n12814) );
  AND2X1 U12864 ( .IN1(n10045), .IN2(CRC_OUT_9_15), .Q(n12816) );
  AND2X1 U12865 ( .IN1(WX514), .IN2(n10020), .Q(n12815) );
  OR2X1 U12866 ( .IN1(n12817), .IN2(n12818), .Q(n12813) );
  AND2X1 U12867 ( .IN1(n9979), .IN2(n12819), .Q(n12818) );
  AND2X1 U12868 ( .IN1(n10075), .IN2(n12820), .Q(n12817) );
  OR2X1 U12869 ( .IN1(n12821), .IN2(n12822), .Q(WX674) );
  OR2X1 U12870 ( .IN1(n12823), .IN2(n12824), .Q(n12822) );
  AND2X1 U12871 ( .IN1(n10045), .IN2(CRC_OUT_9_16), .Q(n12824) );
  AND2X1 U12872 ( .IN1(WX512), .IN2(n10020), .Q(n12823) );
  OR2X1 U12873 ( .IN1(n12825), .IN2(n12826), .Q(n12821) );
  AND2X1 U12874 ( .IN1(n12827), .IN2(n9974), .Q(n12826) );
  AND2X1 U12875 ( .IN1(n10075), .IN2(n12828), .Q(n12825) );
  OR2X1 U12876 ( .IN1(n12829), .IN2(n12830), .Q(WX672) );
  OR2X1 U12877 ( .IN1(n12831), .IN2(n12832), .Q(n12830) );
  AND2X1 U12878 ( .IN1(n10045), .IN2(CRC_OUT_9_17), .Q(n12832) );
  AND2X1 U12879 ( .IN1(WX510), .IN2(n10020), .Q(n12831) );
  OR2X1 U12880 ( .IN1(n12833), .IN2(n12834), .Q(n12829) );
  AND2X1 U12881 ( .IN1(n9979), .IN2(n12835), .Q(n12834) );
  AND2X1 U12882 ( .IN1(n10075), .IN2(n12836), .Q(n12833) );
  OR2X1 U12883 ( .IN1(n12837), .IN2(n12838), .Q(WX670) );
  OR2X1 U12884 ( .IN1(n12839), .IN2(n12840), .Q(n12838) );
  AND2X1 U12885 ( .IN1(n10045), .IN2(CRC_OUT_9_18), .Q(n12840) );
  AND2X1 U12886 ( .IN1(WX508), .IN2(n10020), .Q(n12839) );
  OR2X1 U12887 ( .IN1(n12841), .IN2(n12842), .Q(n12837) );
  AND2X1 U12888 ( .IN1(n9979), .IN2(n12843), .Q(n12842) );
  AND2X1 U12889 ( .IN1(n12844), .IN2(n10057), .Q(n12841) );
  OR2X1 U12890 ( .IN1(n12845), .IN2(n12846), .Q(WX668) );
  OR2X1 U12891 ( .IN1(n12847), .IN2(n12848), .Q(n12846) );
  AND2X1 U12892 ( .IN1(test_so10), .IN2(n10026), .Q(n12848) );
  AND2X1 U12893 ( .IN1(WX506), .IN2(n10021), .Q(n12847) );
  OR2X1 U12894 ( .IN1(n12849), .IN2(n12850), .Q(n12845) );
  AND2X1 U12895 ( .IN1(n9979), .IN2(n12851), .Q(n12850) );
  AND2X1 U12896 ( .IN1(n10075), .IN2(n12852), .Q(n12849) );
  OR2X1 U12897 ( .IN1(n12853), .IN2(n12854), .Q(WX666) );
  OR2X1 U12898 ( .IN1(n12855), .IN2(n12856), .Q(n12854) );
  AND2X1 U12899 ( .IN1(n10045), .IN2(CRC_OUT_9_20), .Q(n12856) );
  AND2X1 U12900 ( .IN1(WX504), .IN2(n10020), .Q(n12855) );
  OR2X1 U12901 ( .IN1(n12857), .IN2(n12858), .Q(n12853) );
  AND2X1 U12902 ( .IN1(n12859), .IN2(n9973), .Q(n12858) );
  AND2X1 U12903 ( .IN1(n10075), .IN2(n12860), .Q(n12857) );
  OR2X1 U12904 ( .IN1(n12861), .IN2(n12862), .Q(WX664) );
  OR2X1 U12905 ( .IN1(n12863), .IN2(n12864), .Q(n12862) );
  AND2X1 U12906 ( .IN1(n10045), .IN2(CRC_OUT_9_21), .Q(n12864) );
  AND2X1 U12907 ( .IN1(WX502), .IN2(n10021), .Q(n12863) );
  OR2X1 U12908 ( .IN1(n12865), .IN2(n12866), .Q(n12861) );
  AND2X1 U12909 ( .IN1(n9979), .IN2(n12867), .Q(n12866) );
  AND2X1 U12910 ( .IN1(n10076), .IN2(n12868), .Q(n12865) );
  OR2X1 U12911 ( .IN1(n12869), .IN2(n12870), .Q(WX662) );
  OR2X1 U12912 ( .IN1(n12871), .IN2(n12872), .Q(n12870) );
  AND2X1 U12913 ( .IN1(n10046), .IN2(CRC_OUT_9_22), .Q(n12872) );
  AND2X1 U12914 ( .IN1(WX500), .IN2(n10021), .Q(n12871) );
  OR2X1 U12915 ( .IN1(n12873), .IN2(n12874), .Q(n12869) );
  AND2X1 U12916 ( .IN1(n9979), .IN2(n12875), .Q(n12874) );
  AND2X1 U12917 ( .IN1(n12876), .IN2(n10057), .Q(n12873) );
  OR2X1 U12918 ( .IN1(n12877), .IN2(n12878), .Q(WX660) );
  OR2X1 U12919 ( .IN1(n12879), .IN2(n12880), .Q(n12878) );
  AND2X1 U12920 ( .IN1(n10046), .IN2(CRC_OUT_9_23), .Q(n12880) );
  AND2X1 U12921 ( .IN1(WX498), .IN2(n10021), .Q(n12879) );
  OR2X1 U12922 ( .IN1(n12881), .IN2(n12882), .Q(n12877) );
  AND2X1 U12923 ( .IN1(n9979), .IN2(n12883), .Q(n12882) );
  AND2X1 U12924 ( .IN1(n10076), .IN2(n12884), .Q(n12881) );
  OR2X1 U12925 ( .IN1(n12885), .IN2(n12886), .Q(WX658) );
  OR2X1 U12926 ( .IN1(n12887), .IN2(n12888), .Q(n12886) );
  AND2X1 U12927 ( .IN1(n10046), .IN2(CRC_OUT_9_24), .Q(n12888) );
  AND2X1 U12928 ( .IN1(WX496), .IN2(n10021), .Q(n12887) );
  OR2X1 U12929 ( .IN1(n12889), .IN2(n12890), .Q(n12885) );
  AND2X1 U12930 ( .IN1(n12891), .IN2(n9973), .Q(n12890) );
  AND2X1 U12931 ( .IN1(n10076), .IN2(n12892), .Q(n12889) );
  OR2X1 U12932 ( .IN1(n12893), .IN2(n12894), .Q(WX656) );
  OR2X1 U12933 ( .IN1(n12895), .IN2(n12896), .Q(n12894) );
  AND2X1 U12934 ( .IN1(n10046), .IN2(CRC_OUT_9_25), .Q(n12896) );
  AND2X1 U12935 ( .IN1(WX494), .IN2(n10021), .Q(n12895) );
  OR2X1 U12936 ( .IN1(n12897), .IN2(n12898), .Q(n12893) );
  AND2X1 U12937 ( .IN1(n9980), .IN2(n12899), .Q(n12898) );
  AND2X1 U12938 ( .IN1(n10076), .IN2(n12900), .Q(n12897) );
  OR2X1 U12939 ( .IN1(n12901), .IN2(n12902), .Q(WX654) );
  OR2X1 U12940 ( .IN1(n12903), .IN2(n12904), .Q(n12902) );
  AND2X1 U12941 ( .IN1(n10046), .IN2(CRC_OUT_9_26), .Q(n12904) );
  AND2X1 U12942 ( .IN1(WX492), .IN2(n10021), .Q(n12903) );
  OR2X1 U12943 ( .IN1(n12905), .IN2(n12906), .Q(n12901) );
  AND2X1 U12944 ( .IN1(n9980), .IN2(n12907), .Q(n12906) );
  AND2X1 U12945 ( .IN1(n10076), .IN2(n12908), .Q(n12905) );
  OR2X1 U12946 ( .IN1(n12909), .IN2(n12910), .Q(WX652) );
  OR2X1 U12947 ( .IN1(n12911), .IN2(n12912), .Q(n12910) );
  AND2X1 U12948 ( .IN1(n10046), .IN2(CRC_OUT_9_27), .Q(n12912) );
  AND2X1 U12949 ( .IN1(WX490), .IN2(n10021), .Q(n12911) );
  OR2X1 U12950 ( .IN1(n12913), .IN2(n12914), .Q(n12909) );
  AND2X1 U12951 ( .IN1(n9980), .IN2(n12915), .Q(n12914) );
  AND2X1 U12952 ( .IN1(n10076), .IN2(n12916), .Q(n12913) );
  OR2X1 U12953 ( .IN1(n12917), .IN2(n12918), .Q(WX650) );
  OR2X1 U12954 ( .IN1(n12919), .IN2(n12920), .Q(n12918) );
  AND2X1 U12955 ( .IN1(n10046), .IN2(CRC_OUT_9_28), .Q(n12920) );
  AND2X1 U12956 ( .IN1(WX488), .IN2(n10021), .Q(n12919) );
  OR2X1 U12957 ( .IN1(n12921), .IN2(n12922), .Q(n12917) );
  AND2X1 U12958 ( .IN1(n12923), .IN2(n9972), .Q(n12922) );
  AND2X1 U12959 ( .IN1(n12924), .IN2(n10057), .Q(n12921) );
  AND2X1 U12960 ( .IN1(n12925), .IN2(n10555), .Q(WX6498) );
  AND2X1 U12961 ( .IN1(n12926), .IN2(n12927), .Q(n12925) );
  OR2X1 U12962 ( .IN1(DFF_958_n1), .IN2(WX6009), .Q(n12927) );
  OR2X1 U12963 ( .IN1(n9646), .IN2(CRC_OUT_5_30), .Q(n12926) );
  AND2X1 U12964 ( .IN1(n12928), .IN2(n10555), .Q(WX6496) );
  AND2X1 U12965 ( .IN1(n12929), .IN2(n12930), .Q(n12928) );
  OR2X1 U12966 ( .IN1(DFF_957_n1), .IN2(WX6011), .Q(n12930) );
  OR2X1 U12967 ( .IN1(n9647), .IN2(CRC_OUT_5_29), .Q(n12929) );
  AND2X1 U12968 ( .IN1(n12931), .IN2(n10555), .Q(WX6494) );
  AND2X1 U12969 ( .IN1(n12932), .IN2(n12933), .Q(n12931) );
  OR2X1 U12970 ( .IN1(DFF_956_n1), .IN2(WX6013), .Q(n12933) );
  OR2X1 U12971 ( .IN1(n9648), .IN2(CRC_OUT_5_28), .Q(n12932) );
  AND2X1 U12972 ( .IN1(n12934), .IN2(n10555), .Q(WX6492) );
  AND2X1 U12973 ( .IN1(n12935), .IN2(n12936), .Q(n12934) );
  OR2X1 U12974 ( .IN1(DFF_955_n1), .IN2(WX6015), .Q(n12936) );
  OR2X1 U12975 ( .IN1(n9649), .IN2(CRC_OUT_5_27), .Q(n12935) );
  AND2X1 U12976 ( .IN1(n12937), .IN2(n10556), .Q(WX6490) );
  AND2X1 U12977 ( .IN1(n12938), .IN2(n12939), .Q(n12937) );
  OR2X1 U12978 ( .IN1(DFF_954_n1), .IN2(WX6017), .Q(n12939) );
  OR2X1 U12979 ( .IN1(n9650), .IN2(CRC_OUT_5_26), .Q(n12938) );
  AND2X1 U12980 ( .IN1(n12940), .IN2(n10556), .Q(WX6488) );
  AND2X1 U12981 ( .IN1(n12941), .IN2(n12942), .Q(n12940) );
  OR2X1 U12982 ( .IN1(DFF_953_n1), .IN2(WX6019), .Q(n12942) );
  OR2X1 U12983 ( .IN1(n9651), .IN2(CRC_OUT_5_25), .Q(n12941) );
  AND2X1 U12984 ( .IN1(n12943), .IN2(n10556), .Q(WX6486) );
  AND2X1 U12985 ( .IN1(n12944), .IN2(n12945), .Q(n12943) );
  OR2X1 U12986 ( .IN1(DFF_952_n1), .IN2(WX6021), .Q(n12945) );
  OR2X1 U12987 ( .IN1(n9652), .IN2(CRC_OUT_5_24), .Q(n12944) );
  AND2X1 U12988 ( .IN1(n12946), .IN2(n10556), .Q(WX6484) );
  AND2X1 U12989 ( .IN1(n12947), .IN2(n12948), .Q(n12946) );
  OR2X1 U12990 ( .IN1(DFF_951_n1), .IN2(WX6023), .Q(n12948) );
  OR2X1 U12991 ( .IN1(n9653), .IN2(CRC_OUT_5_23), .Q(n12947) );
  AND2X1 U12992 ( .IN1(n12949), .IN2(n10556), .Q(WX6482) );
  AND2X1 U12993 ( .IN1(n12950), .IN2(n12951), .Q(n12949) );
  OR2X1 U12994 ( .IN1(DFF_950_n1), .IN2(WX6025), .Q(n12951) );
  OR2X1 U12995 ( .IN1(n9654), .IN2(CRC_OUT_5_22), .Q(n12950) );
  AND2X1 U12996 ( .IN1(n12952), .IN2(n10556), .Q(WX6480) );
  AND2X1 U12997 ( .IN1(n12953), .IN2(n12954), .Q(n12952) );
  OR2X1 U12998 ( .IN1(DFF_949_n1), .IN2(WX6027), .Q(n12954) );
  OR2X1 U12999 ( .IN1(n9655), .IN2(CRC_OUT_5_21), .Q(n12953) );
  OR2X1 U13000 ( .IN1(n12955), .IN2(n12956), .Q(WX648) );
  OR2X1 U13001 ( .IN1(n12957), .IN2(n12958), .Q(n12956) );
  AND2X1 U13002 ( .IN1(n10046), .IN2(CRC_OUT_9_29), .Q(n12958) );
  AND2X1 U13003 ( .IN1(WX486), .IN2(n10021), .Q(n12957) );
  OR2X1 U13004 ( .IN1(n12959), .IN2(n12960), .Q(n12955) );
  AND2X1 U13005 ( .IN1(n9980), .IN2(n12961), .Q(n12960) );
  AND2X1 U13006 ( .IN1(n10076), .IN2(n12962), .Q(n12959) );
  AND2X1 U13007 ( .IN1(n12963), .IN2(n10556), .Q(WX6478) );
  AND2X1 U13008 ( .IN1(n12964), .IN2(n12965), .Q(n12963) );
  OR2X1 U13009 ( .IN1(DFF_948_n1), .IN2(WX6029), .Q(n12965) );
  OR2X1 U13010 ( .IN1(n9656), .IN2(CRC_OUT_5_20), .Q(n12964) );
  AND2X1 U13011 ( .IN1(n12966), .IN2(n10556), .Q(WX6476) );
  AND2X1 U13012 ( .IN1(n12967), .IN2(n12968), .Q(n12966) );
  OR2X1 U13013 ( .IN1(DFF_947_n1), .IN2(WX6031), .Q(n12968) );
  OR2X1 U13014 ( .IN1(n9657), .IN2(CRC_OUT_5_19), .Q(n12967) );
  AND2X1 U13015 ( .IN1(n12969), .IN2(n10556), .Q(WX6474) );
  AND2X1 U13016 ( .IN1(n12970), .IN2(n12971), .Q(n12969) );
  OR2X1 U13017 ( .IN1(DFF_946_n1), .IN2(WX6033), .Q(n12971) );
  OR2X1 U13018 ( .IN1(n9658), .IN2(CRC_OUT_5_18), .Q(n12970) );
  AND2X1 U13019 ( .IN1(n12972), .IN2(n10557), .Q(WX6472) );
  OR2X1 U13020 ( .IN1(n12973), .IN2(n12974), .Q(n12972) );
  AND2X1 U13021 ( .IN1(n9659), .IN2(n9941), .Q(n12974) );
  AND2X1 U13022 ( .IN1(test_so54), .IN2(WX6035), .Q(n12973) );
  AND2X1 U13023 ( .IN1(n12975), .IN2(n10557), .Q(WX6470) );
  AND2X1 U13024 ( .IN1(n12976), .IN2(n12977), .Q(n12975) );
  OR2X1 U13025 ( .IN1(DFF_944_n1), .IN2(WX6037), .Q(n12977) );
  OR2X1 U13026 ( .IN1(n9660), .IN2(CRC_OUT_5_16), .Q(n12976) );
  AND2X1 U13027 ( .IN1(n12978), .IN2(n10557), .Q(WX6468) );
  AND2X1 U13028 ( .IN1(n12979), .IN2(n12980), .Q(n12978) );
  OR2X1 U13029 ( .IN1(DFF_943_n1), .IN2(n12981), .Q(n12980) );
  AND2X1 U13030 ( .IN1(n12982), .IN2(n12983), .Q(n12981) );
  OR2X1 U13031 ( .IN1(DFF_959_n1), .IN2(n9888), .Q(n12983) );
  OR2X1 U13032 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .Q(n12982) );
  OR2X1 U13033 ( .IN1(n12984), .IN2(CRC_OUT_5_15), .Q(n12979) );
  OR2X1 U13034 ( .IN1(n12985), .IN2(n12986), .Q(n12984) );
  AND2X1 U13035 ( .IN1(DFF_959_n1), .IN2(n9888), .Q(n12986) );
  AND2X1 U13036 ( .IN1(test_so52), .IN2(CRC_OUT_5_31), .Q(n12985) );
  AND2X1 U13037 ( .IN1(n12987), .IN2(n10557), .Q(WX6466) );
  AND2X1 U13038 ( .IN1(n12988), .IN2(n12989), .Q(n12987) );
  OR2X1 U13039 ( .IN1(DFF_942_n1), .IN2(WX6041), .Q(n12989) );
  OR2X1 U13040 ( .IN1(n9661), .IN2(CRC_OUT_5_14), .Q(n12988) );
  AND2X1 U13041 ( .IN1(n12990), .IN2(n10557), .Q(WX6464) );
  AND2X1 U13042 ( .IN1(n12991), .IN2(n12992), .Q(n12990) );
  OR2X1 U13043 ( .IN1(DFF_941_n1), .IN2(WX6043), .Q(n12992) );
  OR2X1 U13044 ( .IN1(n9662), .IN2(CRC_OUT_5_13), .Q(n12991) );
  AND2X1 U13045 ( .IN1(n12993), .IN2(n10557), .Q(WX6462) );
  AND2X1 U13046 ( .IN1(n12994), .IN2(n12995), .Q(n12993) );
  OR2X1 U13047 ( .IN1(DFF_940_n1), .IN2(WX6045), .Q(n12995) );
  OR2X1 U13048 ( .IN1(n9663), .IN2(CRC_OUT_5_12), .Q(n12994) );
  AND2X1 U13049 ( .IN1(n12996), .IN2(n10557), .Q(WX6460) );
  AND2X1 U13050 ( .IN1(n12997), .IN2(n12998), .Q(n12996) );
  OR2X1 U13051 ( .IN1(DFF_939_n1), .IN2(WX6047), .Q(n12998) );
  OR2X1 U13052 ( .IN1(n9664), .IN2(CRC_OUT_5_11), .Q(n12997) );
  OR2X1 U13053 ( .IN1(n12999), .IN2(n13000), .Q(WX646) );
  OR2X1 U13054 ( .IN1(n13001), .IN2(n13002), .Q(n13000) );
  AND2X1 U13055 ( .IN1(n10046), .IN2(CRC_OUT_9_30), .Q(n13002) );
  AND2X1 U13056 ( .IN1(WX484), .IN2(n10021), .Q(n13001) );
  OR2X1 U13057 ( .IN1(n13003), .IN2(n13004), .Q(n12999) );
  AND2X1 U13058 ( .IN1(n9994), .IN2(n13005), .Q(n13004) );
  AND2X1 U13059 ( .IN1(n10076), .IN2(n13006), .Q(n13003) );
  AND2X1 U13060 ( .IN1(n13007), .IN2(n10557), .Q(WX6458) );
  OR2X1 U13061 ( .IN1(n13008), .IN2(n13009), .Q(n13007) );
  AND2X1 U13062 ( .IN1(n13010), .IN2(CRC_OUT_5_10), .Q(n13009) );
  AND2X1 U13063 ( .IN1(DFF_938_n1), .IN2(n13011), .Q(n13008) );
  INVX0 U13064 ( .INP(n13010), .ZN(n13011) );
  OR2X1 U13065 ( .IN1(n13012), .IN2(n13013), .Q(n13010) );
  AND2X1 U13066 ( .IN1(DFF_959_n1), .IN2(WX6049), .Q(n13013) );
  AND2X1 U13067 ( .IN1(n9523), .IN2(CRC_OUT_5_31), .Q(n13012) );
  AND2X1 U13068 ( .IN1(n13014), .IN2(n10557), .Q(WX6456) );
  AND2X1 U13069 ( .IN1(n13015), .IN2(n13016), .Q(n13014) );
  OR2X1 U13070 ( .IN1(DFF_937_n1), .IN2(WX6051), .Q(n13016) );
  OR2X1 U13071 ( .IN1(n9665), .IN2(CRC_OUT_5_9), .Q(n13015) );
  AND2X1 U13072 ( .IN1(n13017), .IN2(n10558), .Q(WX6454) );
  AND2X1 U13073 ( .IN1(n13018), .IN2(n13019), .Q(n13017) );
  OR2X1 U13074 ( .IN1(DFF_936_n1), .IN2(WX6053), .Q(n13019) );
  OR2X1 U13075 ( .IN1(n9666), .IN2(CRC_OUT_5_8), .Q(n13018) );
  AND2X1 U13076 ( .IN1(n13020), .IN2(n10558), .Q(WX6452) );
  AND2X1 U13077 ( .IN1(n13021), .IN2(n13022), .Q(n13020) );
  OR2X1 U13078 ( .IN1(DFF_935_n1), .IN2(WX6055), .Q(n13022) );
  OR2X1 U13079 ( .IN1(n9667), .IN2(CRC_OUT_5_7), .Q(n13021) );
  AND2X1 U13080 ( .IN1(n13023), .IN2(n10558), .Q(WX6450) );
  AND2X1 U13081 ( .IN1(n13024), .IN2(n13025), .Q(n13023) );
  OR2X1 U13082 ( .IN1(DFF_934_n1), .IN2(WX6057), .Q(n13025) );
  OR2X1 U13083 ( .IN1(n9668), .IN2(CRC_OUT_5_6), .Q(n13024) );
  AND2X1 U13084 ( .IN1(n13026), .IN2(n10558), .Q(WX6448) );
  AND2X1 U13085 ( .IN1(n13027), .IN2(n13028), .Q(n13026) );
  OR2X1 U13086 ( .IN1(DFF_933_n1), .IN2(WX6059), .Q(n13028) );
  OR2X1 U13087 ( .IN1(n9669), .IN2(CRC_OUT_5_5), .Q(n13027) );
  AND2X1 U13088 ( .IN1(n13029), .IN2(n10558), .Q(WX6446) );
  AND2X1 U13089 ( .IN1(n13030), .IN2(n13031), .Q(n13029) );
  OR2X1 U13090 ( .IN1(DFF_932_n1), .IN2(WX6061), .Q(n13031) );
  OR2X1 U13091 ( .IN1(n9670), .IN2(CRC_OUT_5_4), .Q(n13030) );
  AND2X1 U13092 ( .IN1(n13032), .IN2(n10558), .Q(WX6444) );
  OR2X1 U13093 ( .IN1(n13033), .IN2(n13034), .Q(n13032) );
  AND2X1 U13094 ( .IN1(n13035), .IN2(CRC_OUT_5_3), .Q(n13034) );
  AND2X1 U13095 ( .IN1(DFF_931_n1), .IN2(n13036), .Q(n13033) );
  INVX0 U13096 ( .INP(n13035), .ZN(n13036) );
  OR2X1 U13097 ( .IN1(n13037), .IN2(n13038), .Q(n13035) );
  AND2X1 U13098 ( .IN1(DFF_959_n1), .IN2(WX6063), .Q(n13038) );
  AND2X1 U13099 ( .IN1(n9524), .IN2(CRC_OUT_5_31), .Q(n13037) );
  AND2X1 U13100 ( .IN1(n13039), .IN2(n10558), .Q(WX6442) );
  AND2X1 U13101 ( .IN1(n13040), .IN2(n13041), .Q(n13039) );
  OR2X1 U13102 ( .IN1(DFF_930_n1), .IN2(WX6065), .Q(n13041) );
  OR2X1 U13103 ( .IN1(n9671), .IN2(CRC_OUT_5_2), .Q(n13040) );
  AND2X1 U13104 ( .IN1(n13042), .IN2(n10558), .Q(WX6440) );
  AND2X1 U13105 ( .IN1(n13043), .IN2(n13044), .Q(n13042) );
  OR2X1 U13106 ( .IN1(DFF_929_n1), .IN2(WX6067), .Q(n13044) );
  OR2X1 U13107 ( .IN1(n9672), .IN2(CRC_OUT_5_1), .Q(n13043) );
  OR2X1 U13108 ( .IN1(n13045), .IN2(n13046), .Q(WX644) );
  OR2X1 U13109 ( .IN1(n13047), .IN2(n13048), .Q(n13046) );
  AND2X1 U13110 ( .IN1(n2245), .IN2(WX485), .Q(n13048) );
  AND2X1 U13111 ( .IN1(n10046), .IN2(CRC_OUT_9_31), .Q(n13047) );
  OR2X1 U13112 ( .IN1(n13049), .IN2(n13050), .Q(n13045) );
  AND2X1 U13113 ( .IN1(n9994), .IN2(n13051), .Q(n13050) );
  AND2X1 U13114 ( .IN1(n10076), .IN2(n13052), .Q(n13049) );
  AND2X1 U13115 ( .IN1(n13053), .IN2(n10558), .Q(WX6438) );
  OR2X1 U13116 ( .IN1(n13054), .IN2(n13055), .Q(n13053) );
  AND2X1 U13117 ( .IN1(n9673), .IN2(n9942), .Q(n13055) );
  AND2X1 U13118 ( .IN1(test_so53), .IN2(WX6069), .Q(n13054) );
  AND2X1 U13119 ( .IN1(n13056), .IN2(n10559), .Q(WX6436) );
  AND2X1 U13120 ( .IN1(n13057), .IN2(n13058), .Q(n13056) );
  OR2X1 U13121 ( .IN1(DFF_959_n1), .IN2(WX6071), .Q(n13058) );
  OR2X1 U13122 ( .IN1(n9537), .IN2(CRC_OUT_5_31), .Q(n13057) );
  AND2X1 U13123 ( .IN1(n10596), .IN2(n8479), .Q(WX5910) );
  AND2X1 U13124 ( .IN1(n10596), .IN2(n8480), .Q(WX5908) );
  AND2X1 U13125 ( .IN1(n10594), .IN2(n8481), .Q(WX5906) );
  AND2X1 U13126 ( .IN1(n10593), .IN2(n8482), .Q(WX5904) );
  AND2X1 U13127 ( .IN1(n10593), .IN2(n8483), .Q(WX5902) );
  AND2X1 U13128 ( .IN1(n10593), .IN2(n8484), .Q(WX5900) );
  AND2X1 U13129 ( .IN1(test_so46), .IN2(n10559), .Q(WX5898) );
  AND2X1 U13130 ( .IN1(n10593), .IN2(n8487), .Q(WX5896) );
  AND2X1 U13131 ( .IN1(n10593), .IN2(n8488), .Q(WX5894) );
  AND2X1 U13132 ( .IN1(n10593), .IN2(n8489), .Q(WX5892) );
  AND2X1 U13133 ( .IN1(n10593), .IN2(n8490), .Q(WX5890) );
  AND2X1 U13134 ( .IN1(n10593), .IN2(n8491), .Q(WX5888) );
  AND2X1 U13135 ( .IN1(n10593), .IN2(n8492), .Q(WX5886) );
  AND2X1 U13136 ( .IN1(n10592), .IN2(n8493), .Q(WX5884) );
  AND2X1 U13137 ( .IN1(n10592), .IN2(n8494), .Q(WX5882) );
  AND2X1 U13138 ( .IN1(n10592), .IN2(n8495), .Q(WX5880) );
  OR2X1 U13139 ( .IN1(n13059), .IN2(n13060), .Q(WX5878) );
  OR2X1 U13140 ( .IN1(n13061), .IN2(n13062), .Q(n13060) );
  AND2X1 U13141 ( .IN1(test_so53), .IN2(n10027), .Q(n13062) );
  AND2X1 U13142 ( .IN1(n1003), .IN2(n10022), .Q(n13061) );
  INVX0 U13143 ( .INP(n13063), .ZN(n1003) );
  OR2X1 U13144 ( .IN1(n10641), .IN2(n3910), .Q(n13063) );
  OR2X1 U13145 ( .IN1(n13064), .IN2(n13065), .Q(n13059) );
  AND2X1 U13146 ( .IN1(n9994), .IN2(n13066), .Q(n13065) );
  AND2X1 U13147 ( .IN1(n10076), .IN2(n12050), .Q(n13064) );
  OR2X1 U13148 ( .IN1(n13067), .IN2(n13068), .Q(n12050) );
  INVX0 U13149 ( .INP(n13069), .ZN(n13068) );
  OR2X1 U13150 ( .IN1(n13070), .IN2(n13071), .Q(n13069) );
  AND2X1 U13151 ( .IN1(n13071), .IN2(n13070), .Q(n13067) );
  AND2X1 U13152 ( .IN1(n13072), .IN2(n13073), .Q(n13070) );
  OR2X1 U13153 ( .IN1(WX7236), .IN2(n9361), .Q(n13073) );
  OR2X1 U13154 ( .IN1(WX7172), .IN2(n3627), .Q(n13072) );
  OR2X1 U13155 ( .IN1(n13074), .IN2(n13075), .Q(n13071) );
  AND2X1 U13156 ( .IN1(n9362), .IN2(WX7364), .Q(n13075) );
  AND2X1 U13157 ( .IN1(n9536), .IN2(WX7300), .Q(n13074) );
  OR2X1 U13158 ( .IN1(n13076), .IN2(n13077), .Q(WX5876) );
  OR2X1 U13159 ( .IN1(n13078), .IN2(n13079), .Q(n13077) );
  AND2X1 U13160 ( .IN1(n10046), .IN2(CRC_OUT_5_1), .Q(n13079) );
  AND2X1 U13161 ( .IN1(n1002), .IN2(n10021), .Q(n13078) );
  INVX0 U13162 ( .INP(n13080), .ZN(n1002) );
  OR2X1 U13163 ( .IN1(n10641), .IN2(n3911), .Q(n13080) );
  OR2X1 U13164 ( .IN1(n13081), .IN2(n13082), .Q(n13076) );
  AND2X1 U13165 ( .IN1(n13083), .IN2(n9972), .Q(n13082) );
  AND2X1 U13166 ( .IN1(n10076), .IN2(n12067), .Q(n13081) );
  OR2X1 U13167 ( .IN1(n13084), .IN2(n13085), .Q(n12067) );
  INVX0 U13168 ( .INP(n13086), .ZN(n13085) );
  OR2X1 U13169 ( .IN1(n13087), .IN2(n13088), .Q(n13086) );
  AND2X1 U13170 ( .IN1(n13088), .IN2(n13087), .Q(n13084) );
  AND2X1 U13171 ( .IN1(n13089), .IN2(n13090), .Q(n13087) );
  OR2X1 U13172 ( .IN1(WX7234), .IN2(n9363), .Q(n13090) );
  OR2X1 U13173 ( .IN1(WX7170), .IN2(n3629), .Q(n13089) );
  OR2X1 U13174 ( .IN1(n13091), .IN2(n13092), .Q(n13088) );
  AND2X1 U13175 ( .IN1(n9364), .IN2(WX7362), .Q(n13092) );
  AND2X1 U13176 ( .IN1(n9645), .IN2(WX7298), .Q(n13091) );
  OR2X1 U13177 ( .IN1(n13093), .IN2(n13094), .Q(WX5874) );
  OR2X1 U13178 ( .IN1(n13095), .IN2(n13096), .Q(n13094) );
  AND2X1 U13179 ( .IN1(n10046), .IN2(CRC_OUT_5_2), .Q(n13096) );
  AND2X1 U13180 ( .IN1(n1001), .IN2(n10022), .Q(n13095) );
  INVX0 U13181 ( .INP(n13097), .ZN(n1001) );
  OR2X1 U13182 ( .IN1(n10641), .IN2(n3912), .Q(n13097) );
  OR2X1 U13183 ( .IN1(n13098), .IN2(n13099), .Q(n13093) );
  AND2X1 U13184 ( .IN1(n9994), .IN2(n13100), .Q(n13099) );
  AND2X1 U13185 ( .IN1(n10076), .IN2(n12084), .Q(n13098) );
  OR2X1 U13186 ( .IN1(n13101), .IN2(n13102), .Q(n12084) );
  INVX0 U13187 ( .INP(n13103), .ZN(n13102) );
  OR2X1 U13188 ( .IN1(n13104), .IN2(n13105), .Q(n13103) );
  AND2X1 U13189 ( .IN1(n13105), .IN2(n13104), .Q(n13101) );
  AND2X1 U13190 ( .IN1(n13106), .IN2(n13107), .Q(n13104) );
  OR2X1 U13191 ( .IN1(WX7232), .IN2(n9365), .Q(n13107) );
  OR2X1 U13192 ( .IN1(WX7168), .IN2(n3631), .Q(n13106) );
  OR2X1 U13193 ( .IN1(n13108), .IN2(n13109), .Q(n13105) );
  AND2X1 U13194 ( .IN1(n9366), .IN2(WX7360), .Q(n13109) );
  AND2X1 U13195 ( .IN1(n9644), .IN2(WX7296), .Q(n13108) );
  OR2X1 U13196 ( .IN1(n13110), .IN2(n13111), .Q(WX5872) );
  OR2X1 U13197 ( .IN1(n13112), .IN2(n13113), .Q(n13111) );
  AND2X1 U13198 ( .IN1(n10046), .IN2(CRC_OUT_5_3), .Q(n13113) );
  AND2X1 U13199 ( .IN1(n1000), .IN2(n10022), .Q(n13112) );
  INVX0 U13200 ( .INP(n13114), .ZN(n1000) );
  OR2X1 U13201 ( .IN1(n10641), .IN2(n3913), .Q(n13114) );
  OR2X1 U13202 ( .IN1(n13115), .IN2(n13116), .Q(n13110) );
  AND2X1 U13203 ( .IN1(n13117), .IN2(n9972), .Q(n13116) );
  AND2X1 U13204 ( .IN1(n10076), .IN2(n12101), .Q(n13115) );
  OR2X1 U13205 ( .IN1(n13118), .IN2(n13119), .Q(n12101) );
  INVX0 U13206 ( .INP(n13120), .ZN(n13119) );
  OR2X1 U13207 ( .IN1(n13121), .IN2(n13122), .Q(n13120) );
  AND2X1 U13208 ( .IN1(n13122), .IN2(n13121), .Q(n13118) );
  AND2X1 U13209 ( .IN1(n13123), .IN2(n13124), .Q(n13121) );
  OR2X1 U13210 ( .IN1(WX7230), .IN2(n9367), .Q(n13124) );
  OR2X1 U13211 ( .IN1(WX7166), .IN2(n3633), .Q(n13123) );
  OR2X1 U13212 ( .IN1(n13125), .IN2(n13126), .Q(n13122) );
  AND2X1 U13213 ( .IN1(n9368), .IN2(WX7358), .Q(n13126) );
  AND2X1 U13214 ( .IN1(n9643), .IN2(WX7294), .Q(n13125) );
  OR2X1 U13215 ( .IN1(n13127), .IN2(n13128), .Q(WX5870) );
  OR2X1 U13216 ( .IN1(n13129), .IN2(n13130), .Q(n13128) );
  AND2X1 U13217 ( .IN1(n10047), .IN2(CRC_OUT_5_4), .Q(n13130) );
  AND2X1 U13218 ( .IN1(n999), .IN2(n10022), .Q(n13129) );
  INVX0 U13219 ( .INP(n13131), .ZN(n999) );
  OR2X1 U13220 ( .IN1(n10641), .IN2(n3914), .Q(n13131) );
  OR2X1 U13221 ( .IN1(n13132), .IN2(n13133), .Q(n13127) );
  AND2X1 U13222 ( .IN1(n9994), .IN2(n13134), .Q(n13133) );
  AND2X1 U13223 ( .IN1(n12118), .IN2(n10057), .Q(n13132) );
  AND2X1 U13224 ( .IN1(n13135), .IN2(n13136), .Q(n12118) );
  INVX0 U13225 ( .INP(n13137), .ZN(n13136) );
  AND2X1 U13226 ( .IN1(n13138), .IN2(n13139), .Q(n13137) );
  OR2X1 U13227 ( .IN1(n13139), .IN2(n13138), .Q(n13135) );
  OR2X1 U13228 ( .IN1(n13140), .IN2(n13141), .Q(n13138) );
  AND2X1 U13229 ( .IN1(n3635), .IN2(WX7164), .Q(n13141) );
  INVX0 U13230 ( .INP(n13142), .ZN(n13140) );
  OR2X1 U13231 ( .IN1(WX7164), .IN2(n3635), .Q(n13142) );
  AND2X1 U13232 ( .IN1(n13143), .IN2(n13144), .Q(n13139) );
  OR2X1 U13233 ( .IN1(WX7292), .IN2(test_so64), .Q(n13144) );
  OR2X1 U13234 ( .IN1(n9886), .IN2(n9370), .Q(n13143) );
  OR2X1 U13235 ( .IN1(n13145), .IN2(n13146), .Q(WX5868) );
  OR2X1 U13236 ( .IN1(n13147), .IN2(n13148), .Q(n13146) );
  AND2X1 U13237 ( .IN1(n10047), .IN2(CRC_OUT_5_5), .Q(n13148) );
  AND2X1 U13238 ( .IN1(n998), .IN2(n10022), .Q(n13147) );
  INVX0 U13239 ( .INP(n13149), .ZN(n998) );
  OR2X1 U13240 ( .IN1(n10641), .IN2(n3915), .Q(n13149) );
  OR2X1 U13241 ( .IN1(n13150), .IN2(n13151), .Q(n13145) );
  AND2X1 U13242 ( .IN1(n13152), .IN2(n9972), .Q(n13151) );
  AND2X1 U13243 ( .IN1(n10077), .IN2(n12135), .Q(n13150) );
  OR2X1 U13244 ( .IN1(n13153), .IN2(n13154), .Q(n12135) );
  INVX0 U13245 ( .INP(n13155), .ZN(n13154) );
  OR2X1 U13246 ( .IN1(n13156), .IN2(n13157), .Q(n13155) );
  AND2X1 U13247 ( .IN1(n13157), .IN2(n13156), .Q(n13153) );
  AND2X1 U13248 ( .IN1(n13158), .IN2(n13159), .Q(n13156) );
  OR2X1 U13249 ( .IN1(WX7226), .IN2(n9371), .Q(n13159) );
  OR2X1 U13250 ( .IN1(WX7162), .IN2(n3637), .Q(n13158) );
  OR2X1 U13251 ( .IN1(n13160), .IN2(n13161), .Q(n13157) );
  AND2X1 U13252 ( .IN1(n9372), .IN2(WX7354), .Q(n13161) );
  AND2X1 U13253 ( .IN1(n9642), .IN2(WX7290), .Q(n13160) );
  OR2X1 U13254 ( .IN1(n13162), .IN2(n13163), .Q(WX5866) );
  OR2X1 U13255 ( .IN1(n13164), .IN2(n13165), .Q(n13163) );
  AND2X1 U13256 ( .IN1(n10047), .IN2(CRC_OUT_5_6), .Q(n13165) );
  AND2X1 U13257 ( .IN1(n997), .IN2(n10022), .Q(n13164) );
  INVX0 U13258 ( .INP(n13166), .ZN(n997) );
  OR2X1 U13259 ( .IN1(n10641), .IN2(n3916), .Q(n13166) );
  OR2X1 U13260 ( .IN1(n13167), .IN2(n13168), .Q(n13162) );
  AND2X1 U13261 ( .IN1(n9994), .IN2(n13169), .Q(n13168) );
  AND2X1 U13262 ( .IN1(n12152), .IN2(n10057), .Q(n13167) );
  AND2X1 U13263 ( .IN1(n13170), .IN2(n13171), .Q(n12152) );
  INVX0 U13264 ( .INP(n13172), .ZN(n13171) );
  AND2X1 U13265 ( .IN1(n13173), .IN2(n13174), .Q(n13172) );
  OR2X1 U13266 ( .IN1(n13174), .IN2(n13173), .Q(n13170) );
  OR2X1 U13267 ( .IN1(n13175), .IN2(n13176), .Q(n13173) );
  AND2X1 U13268 ( .IN1(n3639), .IN2(WX7160), .Q(n13176) );
  INVX0 U13269 ( .INP(n13177), .ZN(n13175) );
  OR2X1 U13270 ( .IN1(WX7160), .IN2(n3639), .Q(n13177) );
  AND2X1 U13271 ( .IN1(n13178), .IN2(n13179), .Q(n13174) );
  OR2X1 U13272 ( .IN1(WX7352), .IN2(test_so62), .Q(n13179) );
  OR2X1 U13273 ( .IN1(n9920), .IN2(n9641), .Q(n13178) );
  OR2X1 U13274 ( .IN1(n13180), .IN2(n13181), .Q(WX5864) );
  OR2X1 U13275 ( .IN1(n13182), .IN2(n13183), .Q(n13181) );
  AND2X1 U13276 ( .IN1(n10047), .IN2(CRC_OUT_5_7), .Q(n13183) );
  AND2X1 U13277 ( .IN1(n996), .IN2(n10022), .Q(n13182) );
  INVX0 U13278 ( .INP(n13184), .ZN(n996) );
  OR2X1 U13279 ( .IN1(n10641), .IN2(n3917), .Q(n13184) );
  OR2X1 U13280 ( .IN1(n13185), .IN2(n13186), .Q(n13180) );
  AND2X1 U13281 ( .IN1(n9994), .IN2(n13187), .Q(n13186) );
  AND2X1 U13282 ( .IN1(n10077), .IN2(n12169), .Q(n13185) );
  OR2X1 U13283 ( .IN1(n13188), .IN2(n13189), .Q(n12169) );
  INVX0 U13284 ( .INP(n13190), .ZN(n13189) );
  OR2X1 U13285 ( .IN1(n13191), .IN2(n13192), .Q(n13190) );
  AND2X1 U13286 ( .IN1(n13192), .IN2(n13191), .Q(n13188) );
  AND2X1 U13287 ( .IN1(n13193), .IN2(n13194), .Q(n13191) );
  OR2X1 U13288 ( .IN1(WX7222), .IN2(n9374), .Q(n13194) );
  OR2X1 U13289 ( .IN1(WX7158), .IN2(n3641), .Q(n13193) );
  OR2X1 U13290 ( .IN1(n13195), .IN2(n13196), .Q(n13192) );
  AND2X1 U13291 ( .IN1(n9375), .IN2(WX7350), .Q(n13196) );
  AND2X1 U13292 ( .IN1(n9640), .IN2(WX7286), .Q(n13195) );
  OR2X1 U13293 ( .IN1(n13197), .IN2(n13198), .Q(WX5862) );
  OR2X1 U13294 ( .IN1(n13199), .IN2(n13200), .Q(n13198) );
  AND2X1 U13295 ( .IN1(n10047), .IN2(CRC_OUT_5_8), .Q(n13200) );
  AND2X1 U13296 ( .IN1(n995), .IN2(n10022), .Q(n13199) );
  INVX0 U13297 ( .INP(n13201), .ZN(n995) );
  OR2X1 U13298 ( .IN1(n10641), .IN2(n3918), .Q(n13201) );
  OR2X1 U13299 ( .IN1(n13202), .IN2(n13203), .Q(n13197) );
  AND2X1 U13300 ( .IN1(n9993), .IN2(n13204), .Q(n13203) );
  AND2X1 U13301 ( .IN1(n12186), .IN2(n10056), .Q(n13202) );
  AND2X1 U13302 ( .IN1(n13205), .IN2(n13206), .Q(n12186) );
  INVX0 U13303 ( .INP(n13207), .ZN(n13206) );
  AND2X1 U13304 ( .IN1(n13208), .IN2(n13209), .Q(n13207) );
  OR2X1 U13305 ( .IN1(n13209), .IN2(n13208), .Q(n13205) );
  OR2X1 U13306 ( .IN1(n13210), .IN2(n13211), .Q(n13208) );
  AND2X1 U13307 ( .IN1(n9376), .IN2(WX7284), .Q(n13211) );
  INVX0 U13308 ( .INP(n13212), .ZN(n13210) );
  OR2X1 U13309 ( .IN1(WX7284), .IN2(n9376), .Q(n13212) );
  AND2X1 U13310 ( .IN1(n13213), .IN2(n13214), .Q(n13209) );
  OR2X1 U13311 ( .IN1(WX7348), .IN2(test_so60), .Q(n13214) );
  OR2X1 U13312 ( .IN1(n9921), .IN2(n9639), .Q(n13213) );
  OR2X1 U13313 ( .IN1(n13215), .IN2(n13216), .Q(WX5860) );
  OR2X1 U13314 ( .IN1(n13217), .IN2(n13218), .Q(n13216) );
  AND2X1 U13315 ( .IN1(n10047), .IN2(CRC_OUT_5_9), .Q(n13218) );
  AND2X1 U13316 ( .IN1(n994), .IN2(n10022), .Q(n13217) );
  INVX0 U13317 ( .INP(n13219), .ZN(n994) );
  OR2X1 U13318 ( .IN1(n10641), .IN2(n3919), .Q(n13219) );
  OR2X1 U13319 ( .IN1(n13220), .IN2(n13221), .Q(n13215) );
  AND2X1 U13320 ( .IN1(n9993), .IN2(n13222), .Q(n13221) );
  AND2X1 U13321 ( .IN1(n10077), .IN2(n12203), .Q(n13220) );
  OR2X1 U13322 ( .IN1(n13223), .IN2(n13224), .Q(n12203) );
  INVX0 U13323 ( .INP(n13225), .ZN(n13224) );
  OR2X1 U13324 ( .IN1(n13226), .IN2(n13227), .Q(n13225) );
  AND2X1 U13325 ( .IN1(n13227), .IN2(n13226), .Q(n13223) );
  AND2X1 U13326 ( .IN1(n13228), .IN2(n13229), .Q(n13226) );
  OR2X1 U13327 ( .IN1(WX7218), .IN2(n9378), .Q(n13229) );
  OR2X1 U13328 ( .IN1(WX7154), .IN2(n3645), .Q(n13228) );
  OR2X1 U13329 ( .IN1(n13230), .IN2(n13231), .Q(n13227) );
  AND2X1 U13330 ( .IN1(n9379), .IN2(WX7346), .Q(n13231) );
  AND2X1 U13331 ( .IN1(n9638), .IN2(WX7282), .Q(n13230) );
  OR2X1 U13332 ( .IN1(n13232), .IN2(n13233), .Q(WX5858) );
  OR2X1 U13333 ( .IN1(n13234), .IN2(n13235), .Q(n13233) );
  AND2X1 U13334 ( .IN1(n10047), .IN2(CRC_OUT_5_10), .Q(n13235) );
  AND2X1 U13335 ( .IN1(n993), .IN2(n10022), .Q(n13234) );
  INVX0 U13336 ( .INP(n13236), .ZN(n993) );
  OR2X1 U13337 ( .IN1(n10641), .IN2(n3920), .Q(n13236) );
  OR2X1 U13338 ( .IN1(n13237), .IN2(n13238), .Q(n13232) );
  AND2X1 U13339 ( .IN1(n9993), .IN2(n13239), .Q(n13238) );
  AND2X1 U13340 ( .IN1(n12221), .IN2(n10056), .Q(n13237) );
  AND2X1 U13341 ( .IN1(n13240), .IN2(n13241), .Q(n12221) );
  INVX0 U13342 ( .INP(n13242), .ZN(n13241) );
  AND2X1 U13343 ( .IN1(n13243), .IN2(n13244), .Q(n13242) );
  OR2X1 U13344 ( .IN1(n13244), .IN2(n13243), .Q(n13240) );
  OR2X1 U13345 ( .IN1(n13245), .IN2(n13246), .Q(n13243) );
  AND2X1 U13346 ( .IN1(n3647), .IN2(WX7280), .Q(n13246) );
  INVX0 U13347 ( .INP(n13247), .ZN(n13245) );
  OR2X1 U13348 ( .IN1(WX7280), .IN2(n3647), .Q(n13247) );
  AND2X1 U13349 ( .IN1(n13248), .IN2(n13249), .Q(n13244) );
  OR2X1 U13350 ( .IN1(WX7344), .IN2(test_so58), .Q(n13249) );
  OR2X1 U13351 ( .IN1(n9922), .IN2(n9637), .Q(n13248) );
  OR2X1 U13352 ( .IN1(n13250), .IN2(n13251), .Q(WX5856) );
  OR2X1 U13353 ( .IN1(n13252), .IN2(n13253), .Q(n13251) );
  AND2X1 U13354 ( .IN1(n10047), .IN2(CRC_OUT_5_11), .Q(n13253) );
  AND2X1 U13355 ( .IN1(n992), .IN2(n10022), .Q(n13252) );
  INVX0 U13356 ( .INP(n13254), .ZN(n992) );
  OR2X1 U13357 ( .IN1(n10640), .IN2(n3921), .Q(n13254) );
  OR2X1 U13358 ( .IN1(n13255), .IN2(n13256), .Q(n13250) );
  AND2X1 U13359 ( .IN1(n9993), .IN2(n13257), .Q(n13256) );
  AND2X1 U13360 ( .IN1(n10077), .IN2(n12238), .Q(n13255) );
  OR2X1 U13361 ( .IN1(n13258), .IN2(n13259), .Q(n12238) );
  INVX0 U13362 ( .INP(n13260), .ZN(n13259) );
  OR2X1 U13363 ( .IN1(n13261), .IN2(n13262), .Q(n13260) );
  AND2X1 U13364 ( .IN1(n13262), .IN2(n13261), .Q(n13258) );
  AND2X1 U13365 ( .IN1(n13263), .IN2(n13264), .Q(n13261) );
  OR2X1 U13366 ( .IN1(WX7214), .IN2(n9381), .Q(n13264) );
  OR2X1 U13367 ( .IN1(WX7150), .IN2(n3649), .Q(n13263) );
  OR2X1 U13368 ( .IN1(n13265), .IN2(n13266), .Q(n13262) );
  AND2X1 U13369 ( .IN1(n9382), .IN2(WX7342), .Q(n13266) );
  AND2X1 U13370 ( .IN1(n9522), .IN2(WX7278), .Q(n13265) );
  OR2X1 U13371 ( .IN1(n13267), .IN2(n13268), .Q(WX5854) );
  OR2X1 U13372 ( .IN1(n13269), .IN2(n13270), .Q(n13268) );
  AND2X1 U13373 ( .IN1(n10047), .IN2(CRC_OUT_5_12), .Q(n13270) );
  AND2X1 U13374 ( .IN1(n991), .IN2(n10023), .Q(n13269) );
  INVX0 U13375 ( .INP(n13271), .ZN(n991) );
  OR2X1 U13376 ( .IN1(n10640), .IN2(n3922), .Q(n13271) );
  OR2X1 U13377 ( .IN1(n13272), .IN2(n13273), .Q(n13267) );
  AND2X1 U13378 ( .IN1(n9993), .IN2(n13274), .Q(n13273) );
  AND2X1 U13379 ( .IN1(n10077), .IN2(n12256), .Q(n13272) );
  OR2X1 U13380 ( .IN1(n13275), .IN2(n13276), .Q(n12256) );
  INVX0 U13381 ( .INP(n13277), .ZN(n13276) );
  OR2X1 U13382 ( .IN1(n13278), .IN2(n13279), .Q(n13277) );
  AND2X1 U13383 ( .IN1(n13279), .IN2(n13278), .Q(n13275) );
  AND2X1 U13384 ( .IN1(n13280), .IN2(n13281), .Q(n13278) );
  OR2X1 U13385 ( .IN1(WX7212), .IN2(n9383), .Q(n13281) );
  OR2X1 U13386 ( .IN1(WX7148), .IN2(n3651), .Q(n13280) );
  OR2X1 U13387 ( .IN1(n13282), .IN2(n13283), .Q(n13279) );
  AND2X1 U13388 ( .IN1(n9384), .IN2(WX7340), .Q(n13283) );
  AND2X1 U13389 ( .IN1(n9636), .IN2(WX7276), .Q(n13282) );
  OR2X1 U13390 ( .IN1(n13284), .IN2(n13285), .Q(WX5852) );
  OR2X1 U13391 ( .IN1(n13286), .IN2(n13287), .Q(n13285) );
  AND2X1 U13392 ( .IN1(n10047), .IN2(CRC_OUT_5_13), .Q(n13287) );
  AND2X1 U13393 ( .IN1(n990), .IN2(n10022), .Q(n13286) );
  INVX0 U13394 ( .INP(n13288), .ZN(n990) );
  OR2X1 U13395 ( .IN1(n10640), .IN2(n3923), .Q(n13288) );
  OR2X1 U13396 ( .IN1(n13289), .IN2(n13290), .Q(n13284) );
  AND2X1 U13397 ( .IN1(n9993), .IN2(n13291), .Q(n13290) );
  AND2X1 U13398 ( .IN1(n10077), .IN2(n12273), .Q(n13289) );
  OR2X1 U13399 ( .IN1(n13292), .IN2(n13293), .Q(n12273) );
  INVX0 U13400 ( .INP(n13294), .ZN(n13293) );
  OR2X1 U13401 ( .IN1(n13295), .IN2(n13296), .Q(n13294) );
  AND2X1 U13402 ( .IN1(n13296), .IN2(n13295), .Q(n13292) );
  AND2X1 U13403 ( .IN1(n13297), .IN2(n13298), .Q(n13295) );
  OR2X1 U13404 ( .IN1(WX7210), .IN2(n9385), .Q(n13298) );
  OR2X1 U13405 ( .IN1(WX7146), .IN2(n3653), .Q(n13297) );
  OR2X1 U13406 ( .IN1(n13299), .IN2(n13300), .Q(n13296) );
  AND2X1 U13407 ( .IN1(n9386), .IN2(WX7338), .Q(n13300) );
  AND2X1 U13408 ( .IN1(n9635), .IN2(WX7274), .Q(n13299) );
  OR2X1 U13409 ( .IN1(n13301), .IN2(n13302), .Q(WX5850) );
  OR2X1 U13410 ( .IN1(n13303), .IN2(n13304), .Q(n13302) );
  AND2X1 U13411 ( .IN1(n10047), .IN2(CRC_OUT_5_14), .Q(n13304) );
  AND2X1 U13412 ( .IN1(n989), .IN2(n10023), .Q(n13303) );
  INVX0 U13413 ( .INP(n13305), .ZN(n989) );
  OR2X1 U13414 ( .IN1(n10640), .IN2(n3924), .Q(n13305) );
  OR2X1 U13415 ( .IN1(n13306), .IN2(n13307), .Q(n13301) );
  AND2X1 U13416 ( .IN1(n9993), .IN2(n13308), .Q(n13307) );
  AND2X1 U13417 ( .IN1(n10077), .IN2(n12291), .Q(n13306) );
  OR2X1 U13418 ( .IN1(n13309), .IN2(n13310), .Q(n12291) );
  INVX0 U13419 ( .INP(n13311), .ZN(n13310) );
  OR2X1 U13420 ( .IN1(n13312), .IN2(n13313), .Q(n13311) );
  AND2X1 U13421 ( .IN1(n13313), .IN2(n13312), .Q(n13309) );
  AND2X1 U13422 ( .IN1(n13314), .IN2(n13315), .Q(n13312) );
  OR2X1 U13423 ( .IN1(WX7208), .IN2(n9387), .Q(n13315) );
  OR2X1 U13424 ( .IN1(WX7144), .IN2(n3655), .Q(n13314) );
  OR2X1 U13425 ( .IN1(n13316), .IN2(n13317), .Q(n13313) );
  AND2X1 U13426 ( .IN1(n9388), .IN2(WX7336), .Q(n13317) );
  AND2X1 U13427 ( .IN1(n9634), .IN2(WX7272), .Q(n13316) );
  OR2X1 U13428 ( .IN1(n13318), .IN2(n13319), .Q(WX5848) );
  OR2X1 U13429 ( .IN1(n13320), .IN2(n13321), .Q(n13319) );
  AND2X1 U13430 ( .IN1(n10047), .IN2(CRC_OUT_5_15), .Q(n13321) );
  AND2X1 U13431 ( .IN1(n988), .IN2(n10005), .Q(n13320) );
  INVX0 U13432 ( .INP(n13322), .ZN(n988) );
  OR2X1 U13433 ( .IN1(n10640), .IN2(n3925), .Q(n13322) );
  OR2X1 U13434 ( .IN1(n13323), .IN2(n13324), .Q(n13318) );
  AND2X1 U13435 ( .IN1(n9993), .IN2(n13325), .Q(n13324) );
  AND2X1 U13436 ( .IN1(n10077), .IN2(n12308), .Q(n13323) );
  OR2X1 U13437 ( .IN1(n13326), .IN2(n13327), .Q(n12308) );
  INVX0 U13438 ( .INP(n13328), .ZN(n13327) );
  OR2X1 U13439 ( .IN1(n13329), .IN2(n13330), .Q(n13328) );
  AND2X1 U13440 ( .IN1(n13330), .IN2(n13329), .Q(n13326) );
  AND2X1 U13441 ( .IN1(n13331), .IN2(n13332), .Q(n13329) );
  OR2X1 U13442 ( .IN1(WX7206), .IN2(n9389), .Q(n13332) );
  OR2X1 U13443 ( .IN1(WX7142), .IN2(n3657), .Q(n13331) );
  OR2X1 U13444 ( .IN1(n13333), .IN2(n13334), .Q(n13330) );
  AND2X1 U13445 ( .IN1(n9390), .IN2(WX7334), .Q(n13334) );
  AND2X1 U13446 ( .IN1(n9633), .IN2(WX7270), .Q(n13333) );
  OR2X1 U13447 ( .IN1(n13335), .IN2(n13336), .Q(WX5846) );
  OR2X1 U13448 ( .IN1(n13337), .IN2(n13338), .Q(n13336) );
  AND2X1 U13449 ( .IN1(n10047), .IN2(CRC_OUT_5_16), .Q(n13338) );
  AND2X1 U13450 ( .IN1(n987), .IN2(n10000), .Q(n13337) );
  INVX0 U13451 ( .INP(n13339), .ZN(n987) );
  OR2X1 U13452 ( .IN1(n10640), .IN2(n3926), .Q(n13339) );
  OR2X1 U13453 ( .IN1(n13340), .IN2(n13341), .Q(n13335) );
  AND2X1 U13454 ( .IN1(n13342), .IN2(n9974), .Q(n13341) );
  AND2X1 U13455 ( .IN1(n10077), .IN2(n12326), .Q(n13340) );
  OR2X1 U13456 ( .IN1(n13343), .IN2(n13344), .Q(n12326) );
  INVX0 U13457 ( .INP(n13345), .ZN(n13344) );
  OR2X1 U13458 ( .IN1(n13346), .IN2(n13347), .Q(n13345) );
  AND2X1 U13459 ( .IN1(n13347), .IN2(n13346), .Q(n13343) );
  INVX0 U13460 ( .INP(n13348), .ZN(n13346) );
  OR2X1 U13461 ( .IN1(n13349), .IN2(n13350), .Q(n13348) );
  AND2X1 U13462 ( .IN1(n10520), .IN2(n8421), .Q(n13350) );
  AND2X1 U13463 ( .IN1(n17912), .IN2(n10543), .Q(n13349) );
  OR2X1 U13464 ( .IN1(n13351), .IN2(n13352), .Q(n13347) );
  AND2X1 U13465 ( .IN1(n9521), .IN2(n13353), .Q(n13352) );
  AND2X1 U13466 ( .IN1(n13354), .IN2(n13355), .Q(n13353) );
  OR2X1 U13467 ( .IN1(n9128), .IN2(WX7268), .Q(n13355) );
  OR2X1 U13468 ( .IN1(n9129), .IN2(WX7204), .Q(n13354) );
  AND2X1 U13469 ( .IN1(n13356), .IN2(WX7332), .Q(n13351) );
  OR2X1 U13470 ( .IN1(n13357), .IN2(n13358), .Q(n13356) );
  AND2X1 U13471 ( .IN1(n9128), .IN2(WX7268), .Q(n13358) );
  AND2X1 U13472 ( .IN1(n9129), .IN2(WX7204), .Q(n13357) );
  OR2X1 U13473 ( .IN1(n13359), .IN2(n13360), .Q(WX5844) );
  OR2X1 U13474 ( .IN1(n13361), .IN2(n13362), .Q(n13360) );
  AND2X1 U13475 ( .IN1(test_so54), .IN2(n10026), .Q(n13362) );
  AND2X1 U13476 ( .IN1(n986), .IN2(n10000), .Q(n13361) );
  INVX0 U13477 ( .INP(n13363), .ZN(n986) );
  OR2X1 U13478 ( .IN1(n10640), .IN2(n3927), .Q(n13363) );
  OR2X1 U13479 ( .IN1(n13364), .IN2(n13365), .Q(n13359) );
  AND2X1 U13480 ( .IN1(n9993), .IN2(n13366), .Q(n13365) );
  AND2X1 U13481 ( .IN1(n10077), .IN2(n12350), .Q(n13364) );
  OR2X1 U13482 ( .IN1(n13367), .IN2(n13368), .Q(n12350) );
  INVX0 U13483 ( .INP(n13369), .ZN(n13368) );
  OR2X1 U13484 ( .IN1(n13370), .IN2(n13371), .Q(n13369) );
  AND2X1 U13485 ( .IN1(n13371), .IN2(n13370), .Q(n13367) );
  INVX0 U13486 ( .INP(n13372), .ZN(n13370) );
  OR2X1 U13487 ( .IN1(n13373), .IN2(n13374), .Q(n13372) );
  AND2X1 U13488 ( .IN1(n10520), .IN2(n8422), .Q(n13374) );
  AND2X1 U13489 ( .IN1(n17913), .IN2(n10543), .Q(n13373) );
  OR2X1 U13490 ( .IN1(n13375), .IN2(n13376), .Q(n13371) );
  AND2X1 U13491 ( .IN1(n9632), .IN2(n13377), .Q(n13376) );
  AND2X1 U13492 ( .IN1(n13378), .IN2(n13379), .Q(n13377) );
  OR2X1 U13493 ( .IN1(n9130), .IN2(WX7266), .Q(n13379) );
  OR2X1 U13494 ( .IN1(n9131), .IN2(WX7202), .Q(n13378) );
  AND2X1 U13495 ( .IN1(n13380), .IN2(WX7330), .Q(n13375) );
  OR2X1 U13496 ( .IN1(n13381), .IN2(n13382), .Q(n13380) );
  AND2X1 U13497 ( .IN1(n9130), .IN2(WX7266), .Q(n13382) );
  AND2X1 U13498 ( .IN1(n9131), .IN2(WX7202), .Q(n13381) );
  OR2X1 U13499 ( .IN1(n13383), .IN2(n13384), .Q(WX5842) );
  OR2X1 U13500 ( .IN1(n13385), .IN2(n13386), .Q(n13384) );
  AND2X1 U13501 ( .IN1(n10048), .IN2(CRC_OUT_5_18), .Q(n13386) );
  AND2X1 U13502 ( .IN1(n985), .IN2(n10000), .Q(n13385) );
  INVX0 U13503 ( .INP(n13387), .ZN(n985) );
  OR2X1 U13504 ( .IN1(n10640), .IN2(n3928), .Q(n13387) );
  OR2X1 U13505 ( .IN1(n13388), .IN2(n13389), .Q(n13383) );
  AND2X1 U13506 ( .IN1(n13390), .IN2(n9974), .Q(n13389) );
  AND2X1 U13507 ( .IN1(n10077), .IN2(n12374), .Q(n13388) );
  OR2X1 U13508 ( .IN1(n13391), .IN2(n13392), .Q(n12374) );
  INVX0 U13509 ( .INP(n13393), .ZN(n13392) );
  OR2X1 U13510 ( .IN1(n13394), .IN2(n13395), .Q(n13393) );
  AND2X1 U13511 ( .IN1(n13395), .IN2(n13394), .Q(n13391) );
  INVX0 U13512 ( .INP(n13396), .ZN(n13394) );
  OR2X1 U13513 ( .IN1(n13397), .IN2(n13398), .Q(n13396) );
  AND2X1 U13514 ( .IN1(n10521), .IN2(n8423), .Q(n13398) );
  AND2X1 U13515 ( .IN1(n17914), .IN2(n10543), .Q(n13397) );
  OR2X1 U13516 ( .IN1(n13399), .IN2(n13400), .Q(n13395) );
  AND2X1 U13517 ( .IN1(n9631), .IN2(n13401), .Q(n13400) );
  AND2X1 U13518 ( .IN1(n13402), .IN2(n13403), .Q(n13401) );
  OR2X1 U13519 ( .IN1(n9132), .IN2(WX7264), .Q(n13403) );
  OR2X1 U13520 ( .IN1(n9133), .IN2(WX7200), .Q(n13402) );
  AND2X1 U13521 ( .IN1(n13404), .IN2(WX7328), .Q(n13399) );
  OR2X1 U13522 ( .IN1(n13405), .IN2(n13406), .Q(n13404) );
  AND2X1 U13523 ( .IN1(n9132), .IN2(WX7264), .Q(n13406) );
  AND2X1 U13524 ( .IN1(n9133), .IN2(WX7200), .Q(n13405) );
  OR2X1 U13525 ( .IN1(n13407), .IN2(n13408), .Q(WX5840) );
  OR2X1 U13526 ( .IN1(n13409), .IN2(n13410), .Q(n13408) );
  AND2X1 U13527 ( .IN1(n10048), .IN2(CRC_OUT_5_19), .Q(n13410) );
  AND2X1 U13528 ( .IN1(n984), .IN2(n10000), .Q(n13409) );
  INVX0 U13529 ( .INP(n13411), .ZN(n984) );
  OR2X1 U13530 ( .IN1(n10640), .IN2(n3929), .Q(n13411) );
  OR2X1 U13531 ( .IN1(n13412), .IN2(n13413), .Q(n13407) );
  AND2X1 U13532 ( .IN1(n9993), .IN2(n13414), .Q(n13413) );
  AND2X1 U13533 ( .IN1(n10077), .IN2(n12398), .Q(n13412) );
  OR2X1 U13534 ( .IN1(n13415), .IN2(n13416), .Q(n12398) );
  INVX0 U13535 ( .INP(n13417), .ZN(n13416) );
  OR2X1 U13536 ( .IN1(n13418), .IN2(n13419), .Q(n13417) );
  AND2X1 U13537 ( .IN1(n13419), .IN2(n13418), .Q(n13415) );
  INVX0 U13538 ( .INP(n13420), .ZN(n13418) );
  OR2X1 U13539 ( .IN1(n13421), .IN2(n13422), .Q(n13420) );
  AND2X1 U13540 ( .IN1(n10521), .IN2(n8424), .Q(n13422) );
  AND2X1 U13541 ( .IN1(n17915), .IN2(n10543), .Q(n13421) );
  OR2X1 U13542 ( .IN1(n13423), .IN2(n13424), .Q(n13419) );
  AND2X1 U13543 ( .IN1(n9630), .IN2(n13425), .Q(n13424) );
  AND2X1 U13544 ( .IN1(n13426), .IN2(n13427), .Q(n13425) );
  OR2X1 U13545 ( .IN1(n9134), .IN2(WX7262), .Q(n13427) );
  OR2X1 U13546 ( .IN1(n9135), .IN2(WX7198), .Q(n13426) );
  AND2X1 U13547 ( .IN1(n13428), .IN2(WX7326), .Q(n13423) );
  OR2X1 U13548 ( .IN1(n13429), .IN2(n13430), .Q(n13428) );
  AND2X1 U13549 ( .IN1(n9134), .IN2(WX7262), .Q(n13430) );
  AND2X1 U13550 ( .IN1(n9135), .IN2(WX7198), .Q(n13429) );
  OR2X1 U13551 ( .IN1(n13431), .IN2(n13432), .Q(WX5838) );
  OR2X1 U13552 ( .IN1(n13433), .IN2(n13434), .Q(n13432) );
  AND2X1 U13553 ( .IN1(n10048), .IN2(CRC_OUT_5_20), .Q(n13434) );
  AND2X1 U13554 ( .IN1(n983), .IN2(n10000), .Q(n13433) );
  INVX0 U13555 ( .INP(n13435), .ZN(n983) );
  OR2X1 U13556 ( .IN1(n10640), .IN2(n3930), .Q(n13435) );
  OR2X1 U13557 ( .IN1(n13436), .IN2(n13437), .Q(n13431) );
  AND2X1 U13558 ( .IN1(n13438), .IN2(n9974), .Q(n13437) );
  AND2X1 U13559 ( .IN1(n10077), .IN2(n12422), .Q(n13436) );
  OR2X1 U13560 ( .IN1(n13439), .IN2(n13440), .Q(n12422) );
  INVX0 U13561 ( .INP(n13441), .ZN(n13440) );
  OR2X1 U13562 ( .IN1(n13442), .IN2(n13443), .Q(n13441) );
  AND2X1 U13563 ( .IN1(n13443), .IN2(n13442), .Q(n13439) );
  INVX0 U13564 ( .INP(n13444), .ZN(n13442) );
  OR2X1 U13565 ( .IN1(n13445), .IN2(n13446), .Q(n13444) );
  AND2X1 U13566 ( .IN1(n10521), .IN2(n8425), .Q(n13446) );
  AND2X1 U13567 ( .IN1(n17916), .IN2(n10543), .Q(n13445) );
  OR2X1 U13568 ( .IN1(n13447), .IN2(n13448), .Q(n13443) );
  AND2X1 U13569 ( .IN1(n9629), .IN2(n13449), .Q(n13448) );
  AND2X1 U13570 ( .IN1(n13450), .IN2(n13451), .Q(n13449) );
  OR2X1 U13571 ( .IN1(n9136), .IN2(WX7260), .Q(n13451) );
  OR2X1 U13572 ( .IN1(n9137), .IN2(WX7196), .Q(n13450) );
  AND2X1 U13573 ( .IN1(n13452), .IN2(WX7324), .Q(n13447) );
  OR2X1 U13574 ( .IN1(n13453), .IN2(n13454), .Q(n13452) );
  AND2X1 U13575 ( .IN1(n9136), .IN2(WX7260), .Q(n13454) );
  AND2X1 U13576 ( .IN1(n9137), .IN2(WX7196), .Q(n13453) );
  OR2X1 U13577 ( .IN1(n13455), .IN2(n13456), .Q(WX5836) );
  OR2X1 U13578 ( .IN1(n13457), .IN2(n13458), .Q(n13456) );
  AND2X1 U13579 ( .IN1(n10032), .IN2(CRC_OUT_5_21), .Q(n13458) );
  AND2X1 U13580 ( .IN1(n982), .IN2(n10000), .Q(n13457) );
  INVX0 U13581 ( .INP(n13459), .ZN(n982) );
  OR2X1 U13582 ( .IN1(n10640), .IN2(n3931), .Q(n13459) );
  OR2X1 U13583 ( .IN1(n13460), .IN2(n13461), .Q(n13455) );
  AND2X1 U13584 ( .IN1(n9993), .IN2(n13462), .Q(n13461) );
  AND2X1 U13585 ( .IN1(n12446), .IN2(n10056), .Q(n13460) );
  AND2X1 U13586 ( .IN1(n13463), .IN2(n13464), .Q(n12446) );
  INVX0 U13587 ( .INP(n13465), .ZN(n13464) );
  AND2X1 U13588 ( .IN1(n13466), .IN2(n13467), .Q(n13465) );
  OR2X1 U13589 ( .IN1(n13467), .IN2(n13466), .Q(n13463) );
  OR2X1 U13590 ( .IN1(n13468), .IN2(n13469), .Q(n13466) );
  AND2X1 U13591 ( .IN1(n10521), .IN2(WX7194), .Q(n13469) );
  AND2X1 U13592 ( .IN1(n9138), .IN2(n10543), .Q(n13468) );
  AND2X1 U13593 ( .IN1(n13470), .IN2(n13471), .Q(n13467) );
  INVX0 U13594 ( .INP(n13472), .ZN(n13471) );
  AND2X1 U13595 ( .IN1(n13473), .IN2(WX7258), .Q(n13472) );
  OR2X1 U13596 ( .IN1(WX7258), .IN2(n13473), .Q(n13470) );
  OR2X1 U13597 ( .IN1(n13474), .IN2(n13475), .Q(n13473) );
  AND2X1 U13598 ( .IN1(n17917), .IN2(n9909), .Q(n13475) );
  AND2X1 U13599 ( .IN1(test_so63), .IN2(n8426), .Q(n13474) );
  OR2X1 U13600 ( .IN1(n13476), .IN2(n13477), .Q(WX5834) );
  OR2X1 U13601 ( .IN1(n13478), .IN2(n13479), .Q(n13477) );
  AND2X1 U13602 ( .IN1(n10027), .IN2(CRC_OUT_5_22), .Q(n13479) );
  AND2X1 U13603 ( .IN1(n981), .IN2(n10000), .Q(n13478) );
  INVX0 U13604 ( .INP(n13480), .ZN(n981) );
  OR2X1 U13605 ( .IN1(n10640), .IN2(n3932), .Q(n13480) );
  OR2X1 U13606 ( .IN1(n13481), .IN2(n13482), .Q(n13476) );
  AND2X1 U13607 ( .IN1(n13483), .IN2(n9974), .Q(n13482) );
  AND2X1 U13608 ( .IN1(n10078), .IN2(n12470), .Q(n13481) );
  OR2X1 U13609 ( .IN1(n13484), .IN2(n13485), .Q(n12470) );
  INVX0 U13610 ( .INP(n13486), .ZN(n13485) );
  OR2X1 U13611 ( .IN1(n13487), .IN2(n13488), .Q(n13486) );
  AND2X1 U13612 ( .IN1(n13488), .IN2(n13487), .Q(n13484) );
  INVX0 U13613 ( .INP(n13489), .ZN(n13487) );
  OR2X1 U13614 ( .IN1(n13490), .IN2(n13491), .Q(n13489) );
  AND2X1 U13615 ( .IN1(n10521), .IN2(n8427), .Q(n13491) );
  AND2X1 U13616 ( .IN1(n17918), .IN2(n10543), .Q(n13490) );
  OR2X1 U13617 ( .IN1(n13492), .IN2(n13493), .Q(n13488) );
  AND2X1 U13618 ( .IN1(n9628), .IN2(n13494), .Q(n13493) );
  AND2X1 U13619 ( .IN1(n13495), .IN2(n13496), .Q(n13494) );
  OR2X1 U13620 ( .IN1(n9140), .IN2(WX7256), .Q(n13496) );
  OR2X1 U13621 ( .IN1(n9141), .IN2(WX7192), .Q(n13495) );
  AND2X1 U13622 ( .IN1(n13497), .IN2(WX7320), .Q(n13492) );
  OR2X1 U13623 ( .IN1(n13498), .IN2(n13499), .Q(n13497) );
  AND2X1 U13624 ( .IN1(n9140), .IN2(WX7256), .Q(n13499) );
  AND2X1 U13625 ( .IN1(n9141), .IN2(WX7192), .Q(n13498) );
  OR2X1 U13626 ( .IN1(n13500), .IN2(n13501), .Q(WX5832) );
  OR2X1 U13627 ( .IN1(n13502), .IN2(n13503), .Q(n13501) );
  AND2X1 U13628 ( .IN1(n10029), .IN2(CRC_OUT_5_23), .Q(n13503) );
  AND2X1 U13629 ( .IN1(n980), .IN2(n10000), .Q(n13502) );
  INVX0 U13630 ( .INP(n13504), .ZN(n980) );
  OR2X1 U13631 ( .IN1(n10639), .IN2(n3933), .Q(n13504) );
  OR2X1 U13632 ( .IN1(n13505), .IN2(n13506), .Q(n13500) );
  AND2X1 U13633 ( .IN1(n9993), .IN2(n13507), .Q(n13506) );
  AND2X1 U13634 ( .IN1(n12494), .IN2(n10056), .Q(n13505) );
  AND2X1 U13635 ( .IN1(n13508), .IN2(n13509), .Q(n12494) );
  INVX0 U13636 ( .INP(n13510), .ZN(n13509) );
  AND2X1 U13637 ( .IN1(n13511), .IN2(n13512), .Q(n13510) );
  OR2X1 U13638 ( .IN1(n13512), .IN2(n13511), .Q(n13508) );
  OR2X1 U13639 ( .IN1(n13513), .IN2(n13514), .Q(n13511) );
  AND2X1 U13640 ( .IN1(n10521), .IN2(WX7190), .Q(n13514) );
  AND2X1 U13641 ( .IN1(n9142), .IN2(n10543), .Q(n13513) );
  AND2X1 U13642 ( .IN1(n13515), .IN2(n13516), .Q(n13512) );
  OR2X1 U13643 ( .IN1(n13517), .IN2(n9627), .Q(n13516) );
  INVX0 U13644 ( .INP(n13518), .ZN(n13517) );
  OR2X1 U13645 ( .IN1(WX7318), .IN2(n13518), .Q(n13515) );
  OR2X1 U13646 ( .IN1(n13519), .IN2(n13520), .Q(n13518) );
  AND2X1 U13647 ( .IN1(n17919), .IN2(n9957), .Q(n13520) );
  AND2X1 U13648 ( .IN1(test_so61), .IN2(n8428), .Q(n13519) );
  OR2X1 U13649 ( .IN1(n13521), .IN2(n13522), .Q(WX5830) );
  OR2X1 U13650 ( .IN1(n13523), .IN2(n13524), .Q(n13522) );
  AND2X1 U13651 ( .IN1(n10027), .IN2(CRC_OUT_5_24), .Q(n13524) );
  AND2X1 U13652 ( .IN1(n979), .IN2(n10000), .Q(n13523) );
  INVX0 U13653 ( .INP(n13525), .ZN(n979) );
  OR2X1 U13654 ( .IN1(n10639), .IN2(n3934), .Q(n13525) );
  OR2X1 U13655 ( .IN1(n13526), .IN2(n13527), .Q(n13521) );
  AND2X1 U13656 ( .IN1(n9993), .IN2(n13528), .Q(n13527) );
  AND2X1 U13657 ( .IN1(n10078), .IN2(n12518), .Q(n13526) );
  OR2X1 U13658 ( .IN1(n13529), .IN2(n13530), .Q(n12518) );
  INVX0 U13659 ( .INP(n13531), .ZN(n13530) );
  OR2X1 U13660 ( .IN1(n13532), .IN2(n13533), .Q(n13531) );
  AND2X1 U13661 ( .IN1(n13533), .IN2(n13532), .Q(n13529) );
  INVX0 U13662 ( .INP(n13534), .ZN(n13532) );
  OR2X1 U13663 ( .IN1(n13535), .IN2(n13536), .Q(n13534) );
  AND2X1 U13664 ( .IN1(n10521), .IN2(n8429), .Q(n13536) );
  AND2X1 U13665 ( .IN1(n17920), .IN2(n10543), .Q(n13535) );
  OR2X1 U13666 ( .IN1(n13537), .IN2(n13538), .Q(n13533) );
  AND2X1 U13667 ( .IN1(n9626), .IN2(n13539), .Q(n13538) );
  AND2X1 U13668 ( .IN1(n13540), .IN2(n13541), .Q(n13539) );
  OR2X1 U13669 ( .IN1(n9143), .IN2(WX7252), .Q(n13541) );
  OR2X1 U13670 ( .IN1(n9144), .IN2(WX7188), .Q(n13540) );
  AND2X1 U13671 ( .IN1(n13542), .IN2(WX7316), .Q(n13537) );
  OR2X1 U13672 ( .IN1(n13543), .IN2(n13544), .Q(n13542) );
  AND2X1 U13673 ( .IN1(n9143), .IN2(WX7252), .Q(n13544) );
  AND2X1 U13674 ( .IN1(n9144), .IN2(WX7188), .Q(n13543) );
  OR2X1 U13675 ( .IN1(n13545), .IN2(n13546), .Q(WX5828) );
  OR2X1 U13676 ( .IN1(n13547), .IN2(n13548), .Q(n13546) );
  AND2X1 U13677 ( .IN1(n10028), .IN2(CRC_OUT_5_25), .Q(n13548) );
  AND2X1 U13678 ( .IN1(n978), .IN2(n10000), .Q(n13547) );
  INVX0 U13679 ( .INP(n13549), .ZN(n978) );
  OR2X1 U13680 ( .IN1(n10639), .IN2(n3935), .Q(n13549) );
  OR2X1 U13681 ( .IN1(n13550), .IN2(n13551), .Q(n13545) );
  AND2X1 U13682 ( .IN1(n9992), .IN2(n13552), .Q(n13551) );
  AND2X1 U13683 ( .IN1(n12542), .IN2(n10056), .Q(n13550) );
  AND2X1 U13684 ( .IN1(n13553), .IN2(n13554), .Q(n12542) );
  INVX0 U13685 ( .INP(n13555), .ZN(n13554) );
  AND2X1 U13686 ( .IN1(n13556), .IN2(n13557), .Q(n13555) );
  OR2X1 U13687 ( .IN1(n13557), .IN2(n13556), .Q(n13553) );
  OR2X1 U13688 ( .IN1(n13558), .IN2(n13559), .Q(n13556) );
  AND2X1 U13689 ( .IN1(n10521), .IN2(WX7250), .Q(n13559) );
  AND2X1 U13690 ( .IN1(n9145), .IN2(n10543), .Q(n13558) );
  AND2X1 U13691 ( .IN1(n13560), .IN2(n13561), .Q(n13557) );
  OR2X1 U13692 ( .IN1(n13562), .IN2(n9625), .Q(n13561) );
  INVX0 U13693 ( .INP(n13563), .ZN(n13562) );
  OR2X1 U13694 ( .IN1(WX7314), .IN2(n13563), .Q(n13560) );
  OR2X1 U13695 ( .IN1(n13564), .IN2(n13565), .Q(n13563) );
  AND2X1 U13696 ( .IN1(n17921), .IN2(n9958), .Q(n13565) );
  AND2X1 U13697 ( .IN1(test_so59), .IN2(n8430), .Q(n13564) );
  OR2X1 U13698 ( .IN1(n13566), .IN2(n13567), .Q(WX5826) );
  OR2X1 U13699 ( .IN1(n13568), .IN2(n13569), .Q(n13567) );
  AND2X1 U13700 ( .IN1(n10027), .IN2(CRC_OUT_5_26), .Q(n13569) );
  AND2X1 U13701 ( .IN1(n977), .IN2(n10000), .Q(n13568) );
  INVX0 U13702 ( .INP(n13570), .ZN(n977) );
  OR2X1 U13703 ( .IN1(n10639), .IN2(n3936), .Q(n13570) );
  OR2X1 U13704 ( .IN1(n13571), .IN2(n13572), .Q(n13566) );
  AND2X1 U13705 ( .IN1(n9992), .IN2(n13573), .Q(n13572) );
  AND2X1 U13706 ( .IN1(n10078), .IN2(n12566), .Q(n13571) );
  OR2X1 U13707 ( .IN1(n13574), .IN2(n13575), .Q(n12566) );
  INVX0 U13708 ( .INP(n13576), .ZN(n13575) );
  OR2X1 U13709 ( .IN1(n13577), .IN2(n13578), .Q(n13576) );
  AND2X1 U13710 ( .IN1(n13578), .IN2(n13577), .Q(n13574) );
  INVX0 U13711 ( .INP(n13579), .ZN(n13577) );
  OR2X1 U13712 ( .IN1(n13580), .IN2(n13581), .Q(n13579) );
  AND2X1 U13713 ( .IN1(n10521), .IN2(n8431), .Q(n13581) );
  AND2X1 U13714 ( .IN1(n17922), .IN2(n10543), .Q(n13580) );
  OR2X1 U13715 ( .IN1(n13582), .IN2(n13583), .Q(n13578) );
  AND2X1 U13716 ( .IN1(n9624), .IN2(n13584), .Q(n13583) );
  AND2X1 U13717 ( .IN1(n13585), .IN2(n13586), .Q(n13584) );
  OR2X1 U13718 ( .IN1(n9146), .IN2(WX7248), .Q(n13586) );
  OR2X1 U13719 ( .IN1(n9147), .IN2(WX7184), .Q(n13585) );
  AND2X1 U13720 ( .IN1(n13587), .IN2(WX7312), .Q(n13582) );
  OR2X1 U13721 ( .IN1(n13588), .IN2(n13589), .Q(n13587) );
  AND2X1 U13722 ( .IN1(n9146), .IN2(WX7248), .Q(n13589) );
  AND2X1 U13723 ( .IN1(n9147), .IN2(WX7184), .Q(n13588) );
  OR2X1 U13724 ( .IN1(n13590), .IN2(n13591), .Q(WX5824) );
  OR2X1 U13725 ( .IN1(n13592), .IN2(n13593), .Q(n13591) );
  AND2X1 U13726 ( .IN1(n10028), .IN2(CRC_OUT_5_27), .Q(n13593) );
  AND2X1 U13727 ( .IN1(n976), .IN2(n10001), .Q(n13592) );
  INVX0 U13728 ( .INP(n13594), .ZN(n976) );
  OR2X1 U13729 ( .IN1(n10639), .IN2(n3937), .Q(n13594) );
  OR2X1 U13730 ( .IN1(n13595), .IN2(n13596), .Q(n13590) );
  AND2X1 U13731 ( .IN1(n9992), .IN2(n13597), .Q(n13596) );
  AND2X1 U13732 ( .IN1(n12587), .IN2(n10056), .Q(n13595) );
  AND2X1 U13733 ( .IN1(n13598), .IN2(n13599), .Q(n12587) );
  OR2X1 U13734 ( .IN1(n13600), .IN2(n13601), .Q(n13599) );
  INVX0 U13735 ( .INP(n13602), .ZN(n13600) );
  OR2X1 U13736 ( .IN1(n13603), .IN2(n13602), .Q(n13598) );
  OR2X1 U13737 ( .IN1(n13604), .IN2(n13605), .Q(n13602) );
  AND2X1 U13738 ( .IN1(n10521), .IN2(WX7310), .Q(n13605) );
  AND2X1 U13739 ( .IN1(n9623), .IN2(n10543), .Q(n13604) );
  INVX0 U13740 ( .INP(n13601), .ZN(n13603) );
  OR2X1 U13741 ( .IN1(n13606), .IN2(n13607), .Q(n13601) );
  AND2X1 U13742 ( .IN1(n9149), .IN2(n13608), .Q(n13607) );
  AND2X1 U13743 ( .IN1(n13609), .IN2(n13610), .Q(n13608) );
  OR2X1 U13744 ( .IN1(n9148), .IN2(n9891), .Q(n13610) );
  OR2X1 U13745 ( .IN1(test_so57), .IN2(WX7182), .Q(n13609) );
  AND2X1 U13746 ( .IN1(n13611), .IN2(WX7246), .Q(n13606) );
  OR2X1 U13747 ( .IN1(n13612), .IN2(n13613), .Q(n13611) );
  AND2X1 U13748 ( .IN1(n9148), .IN2(n9891), .Q(n13613) );
  AND2X1 U13749 ( .IN1(test_so57), .IN2(WX7182), .Q(n13612) );
  OR2X1 U13750 ( .IN1(n13614), .IN2(n13615), .Q(WX5822) );
  OR2X1 U13751 ( .IN1(n13616), .IN2(n13617), .Q(n13615) );
  AND2X1 U13752 ( .IN1(n10027), .IN2(CRC_OUT_5_28), .Q(n13617) );
  AND2X1 U13753 ( .IN1(n975), .IN2(n10001), .Q(n13616) );
  INVX0 U13754 ( .INP(n13618), .ZN(n975) );
  OR2X1 U13755 ( .IN1(n10639), .IN2(n3938), .Q(n13618) );
  OR2X1 U13756 ( .IN1(n13619), .IN2(n13620), .Q(n13614) );
  AND2X1 U13757 ( .IN1(n9992), .IN2(n13621), .Q(n13620) );
  AND2X1 U13758 ( .IN1(n10078), .IN2(n12611), .Q(n13619) );
  OR2X1 U13759 ( .IN1(n13622), .IN2(n13623), .Q(n12611) );
  INVX0 U13760 ( .INP(n13624), .ZN(n13623) );
  OR2X1 U13761 ( .IN1(n13625), .IN2(n13626), .Q(n13624) );
  AND2X1 U13762 ( .IN1(n13626), .IN2(n13625), .Q(n13622) );
  INVX0 U13763 ( .INP(n13627), .ZN(n13625) );
  OR2X1 U13764 ( .IN1(n13628), .IN2(n13629), .Q(n13627) );
  AND2X1 U13765 ( .IN1(n10522), .IN2(n8434), .Q(n13629) );
  AND2X1 U13766 ( .IN1(n17923), .IN2(n10542), .Q(n13628) );
  OR2X1 U13767 ( .IN1(n13630), .IN2(n13631), .Q(n13626) );
  AND2X1 U13768 ( .IN1(n9622), .IN2(n13632), .Q(n13631) );
  AND2X1 U13769 ( .IN1(n13633), .IN2(n13634), .Q(n13632) );
  OR2X1 U13770 ( .IN1(n9150), .IN2(WX7244), .Q(n13634) );
  OR2X1 U13771 ( .IN1(n9151), .IN2(WX7180), .Q(n13633) );
  AND2X1 U13772 ( .IN1(n13635), .IN2(WX7308), .Q(n13630) );
  OR2X1 U13773 ( .IN1(n13636), .IN2(n13637), .Q(n13635) );
  AND2X1 U13774 ( .IN1(n9150), .IN2(WX7244), .Q(n13637) );
  AND2X1 U13775 ( .IN1(n9151), .IN2(WX7180), .Q(n13636) );
  OR2X1 U13776 ( .IN1(n13638), .IN2(n13639), .Q(WX5820) );
  OR2X1 U13777 ( .IN1(n13640), .IN2(n13641), .Q(n13639) );
  AND2X1 U13778 ( .IN1(n10028), .IN2(CRC_OUT_5_29), .Q(n13641) );
  AND2X1 U13779 ( .IN1(n974), .IN2(n10001), .Q(n13640) );
  INVX0 U13780 ( .INP(n13642), .ZN(n974) );
  OR2X1 U13781 ( .IN1(n10639), .IN2(n3939), .Q(n13642) );
  OR2X1 U13782 ( .IN1(n13643), .IN2(n13644), .Q(n13638) );
  AND2X1 U13783 ( .IN1(n9992), .IN2(n13645), .Q(n13644) );
  AND2X1 U13784 ( .IN1(n10078), .IN2(n12632), .Q(n13643) );
  OR2X1 U13785 ( .IN1(n13646), .IN2(n13647), .Q(n12632) );
  INVX0 U13786 ( .INP(n13648), .ZN(n13647) );
  OR2X1 U13787 ( .IN1(n13649), .IN2(n13650), .Q(n13648) );
  AND2X1 U13788 ( .IN1(n13650), .IN2(n13649), .Q(n13646) );
  INVX0 U13789 ( .INP(n13651), .ZN(n13649) );
  OR2X1 U13790 ( .IN1(n13652), .IN2(n13653), .Q(n13651) );
  AND2X1 U13791 ( .IN1(n10522), .IN2(n8435), .Q(n13653) );
  AND2X1 U13792 ( .IN1(n17924), .IN2(n10542), .Q(n13652) );
  OR2X1 U13793 ( .IN1(n13654), .IN2(n13655), .Q(n13650) );
  AND2X1 U13794 ( .IN1(n9621), .IN2(n13656), .Q(n13655) );
  AND2X1 U13795 ( .IN1(n13657), .IN2(n13658), .Q(n13656) );
  OR2X1 U13796 ( .IN1(n9152), .IN2(WX7242), .Q(n13658) );
  OR2X1 U13797 ( .IN1(n9153), .IN2(WX7178), .Q(n13657) );
  AND2X1 U13798 ( .IN1(n13659), .IN2(WX7306), .Q(n13654) );
  OR2X1 U13799 ( .IN1(n13660), .IN2(n13661), .Q(n13659) );
  AND2X1 U13800 ( .IN1(n9152), .IN2(WX7242), .Q(n13661) );
  AND2X1 U13801 ( .IN1(n9153), .IN2(WX7178), .Q(n13660) );
  OR2X1 U13802 ( .IN1(n13662), .IN2(n13663), .Q(WX5818) );
  OR2X1 U13803 ( .IN1(n13664), .IN2(n13665), .Q(n13663) );
  AND2X1 U13804 ( .IN1(n10027), .IN2(CRC_OUT_5_30), .Q(n13665) );
  AND2X1 U13805 ( .IN1(n973), .IN2(n10001), .Q(n13664) );
  INVX0 U13806 ( .INP(n13666), .ZN(n973) );
  OR2X1 U13807 ( .IN1(n10639), .IN2(n3940), .Q(n13666) );
  OR2X1 U13808 ( .IN1(n13667), .IN2(n13668), .Q(n13662) );
  AND2X1 U13809 ( .IN1(n9992), .IN2(n13669), .Q(n13668) );
  AND2X1 U13810 ( .IN1(n10078), .IN2(n12656), .Q(n13667) );
  OR2X1 U13811 ( .IN1(n13670), .IN2(n13671), .Q(n12656) );
  INVX0 U13812 ( .INP(n13672), .ZN(n13671) );
  OR2X1 U13813 ( .IN1(n13673), .IN2(n13674), .Q(n13672) );
  AND2X1 U13814 ( .IN1(n13674), .IN2(n13673), .Q(n13670) );
  INVX0 U13815 ( .INP(n13675), .ZN(n13673) );
  OR2X1 U13816 ( .IN1(n13676), .IN2(n13677), .Q(n13675) );
  AND2X1 U13817 ( .IN1(n10522), .IN2(n8436), .Q(n13677) );
  AND2X1 U13818 ( .IN1(n17925), .IN2(n10542), .Q(n13676) );
  OR2X1 U13819 ( .IN1(n13678), .IN2(n13679), .Q(n13674) );
  AND2X1 U13820 ( .IN1(n9620), .IN2(n13680), .Q(n13679) );
  AND2X1 U13821 ( .IN1(n13681), .IN2(n13682), .Q(n13680) );
  OR2X1 U13822 ( .IN1(n9154), .IN2(WX7240), .Q(n13682) );
  OR2X1 U13823 ( .IN1(n9155), .IN2(WX7176), .Q(n13681) );
  AND2X1 U13824 ( .IN1(n13683), .IN2(WX7304), .Q(n13678) );
  OR2X1 U13825 ( .IN1(n13684), .IN2(n13685), .Q(n13683) );
  AND2X1 U13826 ( .IN1(n9154), .IN2(WX7240), .Q(n13685) );
  AND2X1 U13827 ( .IN1(n9155), .IN2(WX7176), .Q(n13684) );
  OR2X1 U13828 ( .IN1(n13686), .IN2(n13687), .Q(WX5816) );
  OR2X1 U13829 ( .IN1(n13688), .IN2(n13689), .Q(n13687) );
  AND2X1 U13830 ( .IN1(n2245), .IN2(WX5657), .Q(n13689) );
  AND2X1 U13831 ( .IN1(n10029), .IN2(CRC_OUT_5_31), .Q(n13688) );
  OR2X1 U13832 ( .IN1(n13690), .IN2(n13691), .Q(n13686) );
  AND2X1 U13833 ( .IN1(n9992), .IN2(n13692), .Q(n13691) );
  AND2X1 U13834 ( .IN1(n10078), .IN2(n12676), .Q(n13690) );
  OR2X1 U13835 ( .IN1(n13693), .IN2(n13694), .Q(n12676) );
  INVX0 U13836 ( .INP(n13695), .ZN(n13694) );
  OR2X1 U13837 ( .IN1(n13696), .IN2(n13697), .Q(n13695) );
  AND2X1 U13838 ( .IN1(n13697), .IN2(n13696), .Q(n13693) );
  INVX0 U13839 ( .INP(n13698), .ZN(n13696) );
  OR2X1 U13840 ( .IN1(n13699), .IN2(n13700), .Q(n13698) );
  AND2X1 U13841 ( .IN1(n10522), .IN2(n8437), .Q(n13700) );
  AND2X1 U13842 ( .IN1(n17926), .IN2(n10542), .Q(n13699) );
  OR2X1 U13843 ( .IN1(n13701), .IN2(n13702), .Q(n13697) );
  AND2X1 U13844 ( .IN1(n9619), .IN2(n13703), .Q(n13702) );
  AND2X1 U13845 ( .IN1(n13704), .IN2(n13705), .Q(n13703) );
  OR2X1 U13846 ( .IN1(n9034), .IN2(WX7238), .Q(n13705) );
  OR2X1 U13847 ( .IN1(n9035), .IN2(WX7174), .Q(n13704) );
  AND2X1 U13848 ( .IN1(n13706), .IN2(WX7302), .Q(n13701) );
  OR2X1 U13849 ( .IN1(n13707), .IN2(n13708), .Q(n13706) );
  AND2X1 U13850 ( .IN1(n9034), .IN2(WX7238), .Q(n13708) );
  AND2X1 U13851 ( .IN1(n9035), .IN2(WX7174), .Q(n13707) );
  AND2X1 U13852 ( .IN1(n9847), .IN2(n10559), .Q(WX5718) );
  AND2X1 U13853 ( .IN1(n9877), .IN2(n10559), .Q(WX546) );
  AND2X1 U13854 ( .IN1(n13709), .IN2(n10559), .Q(WX5205) );
  AND2X1 U13855 ( .IN1(n13710), .IN2(n13711), .Q(n13709) );
  OR2X1 U13856 ( .IN1(DFF_766_n1), .IN2(WX4716), .Q(n13711) );
  OR2X1 U13857 ( .IN1(n9674), .IN2(CRC_OUT_6_30), .Q(n13710) );
  AND2X1 U13858 ( .IN1(n13712), .IN2(n10559), .Q(WX5203) );
  AND2X1 U13859 ( .IN1(n13713), .IN2(n13714), .Q(n13712) );
  OR2X1 U13860 ( .IN1(DFF_765_n1), .IN2(WX4718), .Q(n13714) );
  OR2X1 U13861 ( .IN1(n9675), .IN2(CRC_OUT_6_29), .Q(n13713) );
  AND2X1 U13862 ( .IN1(n13715), .IN2(n10559), .Q(WX5201) );
  AND2X1 U13863 ( .IN1(n13716), .IN2(n13717), .Q(n13715) );
  OR2X1 U13864 ( .IN1(DFF_764_n1), .IN2(WX4720), .Q(n13717) );
  OR2X1 U13865 ( .IN1(n9676), .IN2(CRC_OUT_6_28), .Q(n13716) );
  AND2X1 U13866 ( .IN1(n13718), .IN2(n10559), .Q(WX5199) );
  OR2X1 U13867 ( .IN1(n13719), .IN2(n13720), .Q(n13718) );
  AND2X1 U13868 ( .IN1(DFF_763_n1), .IN2(n9910), .Q(n13720) );
  AND2X1 U13869 ( .IN1(test_so40), .IN2(CRC_OUT_6_27), .Q(n13719) );
  AND2X1 U13870 ( .IN1(n13721), .IN2(n10560), .Q(WX5197) );
  AND2X1 U13871 ( .IN1(n13722), .IN2(n13723), .Q(n13721) );
  OR2X1 U13872 ( .IN1(DFF_762_n1), .IN2(WX4724), .Q(n13723) );
  OR2X1 U13873 ( .IN1(n9677), .IN2(CRC_OUT_6_26), .Q(n13722) );
  AND2X1 U13874 ( .IN1(n13724), .IN2(n10560), .Q(WX5195) );
  AND2X1 U13875 ( .IN1(n13725), .IN2(n13726), .Q(n13724) );
  OR2X1 U13876 ( .IN1(DFF_761_n1), .IN2(WX4726), .Q(n13726) );
  OR2X1 U13877 ( .IN1(n9678), .IN2(CRC_OUT_6_25), .Q(n13725) );
  AND2X1 U13878 ( .IN1(n13727), .IN2(n10560), .Q(WX5193) );
  AND2X1 U13879 ( .IN1(n13728), .IN2(n13729), .Q(n13727) );
  OR2X1 U13880 ( .IN1(DFF_760_n1), .IN2(WX4728), .Q(n13729) );
  OR2X1 U13881 ( .IN1(n9679), .IN2(CRC_OUT_6_24), .Q(n13728) );
  AND2X1 U13882 ( .IN1(n13730), .IN2(n10560), .Q(WX5191) );
  AND2X1 U13883 ( .IN1(n13731), .IN2(n13732), .Q(n13730) );
  OR2X1 U13884 ( .IN1(DFF_759_n1), .IN2(WX4730), .Q(n13732) );
  OR2X1 U13885 ( .IN1(n9680), .IN2(CRC_OUT_6_23), .Q(n13731) );
  AND2X1 U13886 ( .IN1(n13733), .IN2(n10560), .Q(WX5189) );
  OR2X1 U13887 ( .IN1(n13734), .IN2(n13735), .Q(n13733) );
  AND2X1 U13888 ( .IN1(n9681), .IN2(n9943), .Q(n13735) );
  AND2X1 U13889 ( .IN1(test_so43), .IN2(WX4732), .Q(n13734) );
  AND2X1 U13890 ( .IN1(n13736), .IN2(n10560), .Q(WX5187) );
  AND2X1 U13891 ( .IN1(n13737), .IN2(n13738), .Q(n13736) );
  OR2X1 U13892 ( .IN1(DFF_757_n1), .IN2(WX4734), .Q(n13738) );
  OR2X1 U13893 ( .IN1(n9682), .IN2(CRC_OUT_6_21), .Q(n13737) );
  AND2X1 U13894 ( .IN1(n13739), .IN2(n10560), .Q(WX5185) );
  AND2X1 U13895 ( .IN1(n13740), .IN2(n13741), .Q(n13739) );
  OR2X1 U13896 ( .IN1(DFF_756_n1), .IN2(WX4736), .Q(n13741) );
  OR2X1 U13897 ( .IN1(n9683), .IN2(CRC_OUT_6_20), .Q(n13740) );
  AND2X1 U13898 ( .IN1(n13742), .IN2(n10560), .Q(WX5183) );
  AND2X1 U13899 ( .IN1(n13743), .IN2(n13744), .Q(n13742) );
  OR2X1 U13900 ( .IN1(DFF_755_n1), .IN2(WX4738), .Q(n13744) );
  OR2X1 U13901 ( .IN1(n9684), .IN2(CRC_OUT_6_19), .Q(n13743) );
  AND2X1 U13902 ( .IN1(n13745), .IN2(n10560), .Q(WX5181) );
  AND2X1 U13903 ( .IN1(n13746), .IN2(n13747), .Q(n13745) );
  OR2X1 U13904 ( .IN1(DFF_754_n1), .IN2(WX4740), .Q(n13747) );
  OR2X1 U13905 ( .IN1(n9685), .IN2(CRC_OUT_6_18), .Q(n13746) );
  AND2X1 U13906 ( .IN1(n13748), .IN2(n10561), .Q(WX5179) );
  AND2X1 U13907 ( .IN1(n13749), .IN2(n13750), .Q(n13748) );
  OR2X1 U13908 ( .IN1(DFF_753_n1), .IN2(WX4742), .Q(n13750) );
  OR2X1 U13909 ( .IN1(n9686), .IN2(CRC_OUT_6_17), .Q(n13749) );
  AND2X1 U13910 ( .IN1(n13751), .IN2(n10561), .Q(WX5177) );
  AND2X1 U13911 ( .IN1(n13752), .IN2(n13753), .Q(n13751) );
  OR2X1 U13912 ( .IN1(DFF_752_n1), .IN2(WX4744), .Q(n13753) );
  OR2X1 U13913 ( .IN1(n9687), .IN2(CRC_OUT_6_16), .Q(n13752) );
  AND2X1 U13914 ( .IN1(n13754), .IN2(n10561), .Q(WX5175) );
  OR2X1 U13915 ( .IN1(n13755), .IN2(n13756), .Q(n13754) );
  AND2X1 U13916 ( .IN1(n13757), .IN2(CRC_OUT_6_15), .Q(n13756) );
  AND2X1 U13917 ( .IN1(DFF_751_n1), .IN2(n13758), .Q(n13755) );
  INVX0 U13918 ( .INP(n13757), .ZN(n13758) );
  OR2X1 U13919 ( .IN1(n13759), .IN2(n13760), .Q(n13757) );
  AND2X1 U13920 ( .IN1(DFF_767_n1), .IN2(WX4746), .Q(n13760) );
  AND2X1 U13921 ( .IN1(n9525), .IN2(CRC_OUT_6_31), .Q(n13759) );
  AND2X1 U13922 ( .IN1(n13761), .IN2(n10561), .Q(WX5173) );
  AND2X1 U13923 ( .IN1(n13762), .IN2(n13763), .Q(n13761) );
  OR2X1 U13924 ( .IN1(DFF_750_n1), .IN2(WX4748), .Q(n13763) );
  OR2X1 U13925 ( .IN1(n9688), .IN2(CRC_OUT_6_14), .Q(n13762) );
  AND2X1 U13926 ( .IN1(n13764), .IN2(n10561), .Q(WX5171) );
  AND2X1 U13927 ( .IN1(n13765), .IN2(n13766), .Q(n13764) );
  OR2X1 U13928 ( .IN1(DFF_749_n1), .IN2(WX4750), .Q(n13766) );
  OR2X1 U13929 ( .IN1(n9689), .IN2(CRC_OUT_6_13), .Q(n13765) );
  AND2X1 U13930 ( .IN1(n13767), .IN2(n10561), .Q(WX5169) );
  AND2X1 U13931 ( .IN1(n13768), .IN2(n13769), .Q(n13767) );
  OR2X1 U13932 ( .IN1(DFF_748_n1), .IN2(WX4752), .Q(n13769) );
  OR2X1 U13933 ( .IN1(n9690), .IN2(CRC_OUT_6_12), .Q(n13768) );
  AND2X1 U13934 ( .IN1(n13770), .IN2(n10561), .Q(WX5167) );
  AND2X1 U13935 ( .IN1(n13771), .IN2(n13772), .Q(n13770) );
  OR2X1 U13936 ( .IN1(DFF_747_n1), .IN2(WX4754), .Q(n13772) );
  OR2X1 U13937 ( .IN1(n9691), .IN2(CRC_OUT_6_11), .Q(n13771) );
  AND2X1 U13938 ( .IN1(n13773), .IN2(n10561), .Q(WX5165) );
  AND2X1 U13939 ( .IN1(n13774), .IN2(n13775), .Q(n13773) );
  OR2X1 U13940 ( .IN1(DFF_746_n1), .IN2(n13776), .Q(n13775) );
  AND2X1 U13941 ( .IN1(n13777), .IN2(n13778), .Q(n13776) );
  OR2X1 U13942 ( .IN1(DFF_767_n1), .IN2(n9887), .Q(n13778) );
  OR2X1 U13943 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .Q(n13777) );
  OR2X1 U13944 ( .IN1(n13779), .IN2(CRC_OUT_6_10), .Q(n13774) );
  OR2X1 U13945 ( .IN1(n13780), .IN2(n13781), .Q(n13779) );
  AND2X1 U13946 ( .IN1(DFF_767_n1), .IN2(n9887), .Q(n13781) );
  AND2X1 U13947 ( .IN1(test_so41), .IN2(CRC_OUT_6_31), .Q(n13780) );
  AND2X1 U13948 ( .IN1(n13782), .IN2(n10561), .Q(WX5163) );
  AND2X1 U13949 ( .IN1(n13783), .IN2(n13784), .Q(n13782) );
  OR2X1 U13950 ( .IN1(DFF_745_n1), .IN2(WX4758), .Q(n13784) );
  OR2X1 U13951 ( .IN1(n9692), .IN2(CRC_OUT_6_9), .Q(n13783) );
  AND2X1 U13952 ( .IN1(n13785), .IN2(n10562), .Q(WX5161) );
  AND2X1 U13953 ( .IN1(n13786), .IN2(n13787), .Q(n13785) );
  OR2X1 U13954 ( .IN1(DFF_744_n1), .IN2(WX4760), .Q(n13787) );
  OR2X1 U13955 ( .IN1(n9693), .IN2(CRC_OUT_6_8), .Q(n13786) );
  AND2X1 U13956 ( .IN1(n13788), .IN2(n10562), .Q(WX5159) );
  AND2X1 U13957 ( .IN1(n13789), .IN2(n13790), .Q(n13788) );
  OR2X1 U13958 ( .IN1(DFF_743_n1), .IN2(WX4762), .Q(n13790) );
  OR2X1 U13959 ( .IN1(n9694), .IN2(CRC_OUT_6_7), .Q(n13789) );
  AND2X1 U13960 ( .IN1(n13791), .IN2(n10562), .Q(WX5157) );
  AND2X1 U13961 ( .IN1(n13792), .IN2(n13793), .Q(n13791) );
  OR2X1 U13962 ( .IN1(DFF_742_n1), .IN2(WX4764), .Q(n13793) );
  OR2X1 U13963 ( .IN1(n9695), .IN2(CRC_OUT_6_6), .Q(n13792) );
  AND2X1 U13964 ( .IN1(n13794), .IN2(n10562), .Q(WX5155) );
  OR2X1 U13965 ( .IN1(n13795), .IN2(n13796), .Q(n13794) );
  AND2X1 U13966 ( .IN1(n9696), .IN2(n9944), .Q(n13796) );
  AND2X1 U13967 ( .IN1(test_so42), .IN2(WX4766), .Q(n13795) );
  AND2X1 U13968 ( .IN1(n13797), .IN2(n10562), .Q(WX5153) );
  AND2X1 U13969 ( .IN1(n13798), .IN2(n13799), .Q(n13797) );
  OR2X1 U13970 ( .IN1(DFF_740_n1), .IN2(WX4768), .Q(n13799) );
  OR2X1 U13971 ( .IN1(n9697), .IN2(CRC_OUT_6_4), .Q(n13798) );
  AND2X1 U13972 ( .IN1(n13800), .IN2(n10562), .Q(WX5151) );
  OR2X1 U13973 ( .IN1(n13801), .IN2(n13802), .Q(n13800) );
  AND2X1 U13974 ( .IN1(n13803), .IN2(CRC_OUT_6_3), .Q(n13802) );
  AND2X1 U13975 ( .IN1(DFF_739_n1), .IN2(n13804), .Q(n13801) );
  INVX0 U13976 ( .INP(n13803), .ZN(n13804) );
  OR2X1 U13977 ( .IN1(n13805), .IN2(n13806), .Q(n13803) );
  AND2X1 U13978 ( .IN1(DFF_767_n1), .IN2(WX4770), .Q(n13806) );
  AND2X1 U13979 ( .IN1(n9526), .IN2(CRC_OUT_6_31), .Q(n13805) );
  AND2X1 U13980 ( .IN1(n13807), .IN2(n10562), .Q(WX5149) );
  AND2X1 U13981 ( .IN1(n13808), .IN2(n13809), .Q(n13807) );
  OR2X1 U13982 ( .IN1(DFF_738_n1), .IN2(WX4772), .Q(n13809) );
  OR2X1 U13983 ( .IN1(n9698), .IN2(CRC_OUT_6_2), .Q(n13808) );
  AND2X1 U13984 ( .IN1(n13810), .IN2(n10562), .Q(WX5147) );
  AND2X1 U13985 ( .IN1(n13811), .IN2(n13812), .Q(n13810) );
  OR2X1 U13986 ( .IN1(DFF_737_n1), .IN2(WX4774), .Q(n13812) );
  OR2X1 U13987 ( .IN1(n9699), .IN2(CRC_OUT_6_1), .Q(n13811) );
  AND2X1 U13988 ( .IN1(n13813), .IN2(n10562), .Q(WX5145) );
  AND2X1 U13989 ( .IN1(n13814), .IN2(n13815), .Q(n13813) );
  OR2X1 U13990 ( .IN1(DFF_736_n1), .IN2(WX4776), .Q(n13815) );
  OR2X1 U13991 ( .IN1(n9700), .IN2(CRC_OUT_6_0), .Q(n13814) );
  AND2X1 U13992 ( .IN1(n13816), .IN2(n10563), .Q(WX5143) );
  AND2X1 U13993 ( .IN1(n13817), .IN2(n13818), .Q(n13816) );
  OR2X1 U13994 ( .IN1(DFF_767_n1), .IN2(WX4778), .Q(n13818) );
  OR2X1 U13995 ( .IN1(n9538), .IN2(CRC_OUT_6_31), .Q(n13817) );
  AND2X1 U13996 ( .IN1(n10590), .IN2(n8537), .Q(WX4617) );
  AND2X1 U13997 ( .IN1(test_so35), .IN2(n10563), .Q(WX4615) );
  AND2X1 U13998 ( .IN1(n10591), .IN2(n8540), .Q(WX4613) );
  AND2X1 U13999 ( .IN1(n10590), .IN2(n8541), .Q(WX4611) );
  AND2X1 U14000 ( .IN1(n10589), .IN2(n8542), .Q(WX4609) );
  AND2X1 U14001 ( .IN1(n10592), .IN2(n8543), .Q(WX4607) );
  AND2X1 U14002 ( .IN1(n10589), .IN2(n8544), .Q(WX4605) );
  AND2X1 U14003 ( .IN1(n10592), .IN2(n8545), .Q(WX4603) );
  AND2X1 U14004 ( .IN1(n10589), .IN2(n8546), .Q(WX4601) );
  AND2X1 U14005 ( .IN1(n10591), .IN2(n8547), .Q(WX4599) );
  AND2X1 U14006 ( .IN1(n10589), .IN2(n8548), .Q(WX4597) );
  AND2X1 U14007 ( .IN1(n10589), .IN2(n8549), .Q(WX4595) );
  AND2X1 U14008 ( .IN1(n10589), .IN2(n8550), .Q(WX4593) );
  AND2X1 U14009 ( .IN1(n10594), .IN2(n8551), .Q(WX4591) );
  AND2X1 U14010 ( .IN1(n10590), .IN2(n8552), .Q(WX4589) );
  AND2X1 U14011 ( .IN1(n10592), .IN2(n8553), .Q(WX4587) );
  OR2X1 U14012 ( .IN1(n13819), .IN2(n13820), .Q(WX4585) );
  OR2X1 U14013 ( .IN1(n13821), .IN2(n13822), .Q(n13820) );
  AND2X1 U14014 ( .IN1(n10027), .IN2(CRC_OUT_6_0), .Q(n13822) );
  AND2X1 U14015 ( .IN1(n762), .IN2(n10001), .Q(n13821) );
  INVX0 U14016 ( .INP(n13823), .ZN(n762) );
  OR2X1 U14017 ( .IN1(n10639), .IN2(n3941), .Q(n13823) );
  OR2X1 U14018 ( .IN1(n13824), .IN2(n13825), .Q(n13819) );
  AND2X1 U14019 ( .IN1(n13826), .IN2(n9975), .Q(n13825) );
  AND2X1 U14020 ( .IN1(n10078), .IN2(n13066), .Q(n13824) );
  OR2X1 U14021 ( .IN1(n13827), .IN2(n13828), .Q(n13066) );
  INVX0 U14022 ( .INP(n13829), .ZN(n13828) );
  OR2X1 U14023 ( .IN1(n13830), .IN2(n13831), .Q(n13829) );
  AND2X1 U14024 ( .IN1(n13831), .IN2(n13830), .Q(n13827) );
  AND2X1 U14025 ( .IN1(n13832), .IN2(n13833), .Q(n13830) );
  OR2X1 U14026 ( .IN1(WX5943), .IN2(n9391), .Q(n13833) );
  OR2X1 U14027 ( .IN1(WX5879), .IN2(n3659), .Q(n13832) );
  OR2X1 U14028 ( .IN1(n13834), .IN2(n13835), .Q(n13831) );
  AND2X1 U14029 ( .IN1(n9392), .IN2(WX6071), .Q(n13835) );
  AND2X1 U14030 ( .IN1(n9537), .IN2(WX6007), .Q(n13834) );
  OR2X1 U14031 ( .IN1(n13836), .IN2(n13837), .Q(WX4583) );
  OR2X1 U14032 ( .IN1(n13838), .IN2(n13839), .Q(n13837) );
  AND2X1 U14033 ( .IN1(n10028), .IN2(CRC_OUT_6_1), .Q(n13839) );
  AND2X1 U14034 ( .IN1(n761), .IN2(n10001), .Q(n13838) );
  INVX0 U14035 ( .INP(n13840), .ZN(n761) );
  OR2X1 U14036 ( .IN1(n10639), .IN2(n3942), .Q(n13840) );
  OR2X1 U14037 ( .IN1(n13841), .IN2(n13842), .Q(n13836) );
  AND2X1 U14038 ( .IN1(n9992), .IN2(n13843), .Q(n13842) );
  AND2X1 U14039 ( .IN1(n13083), .IN2(n10056), .Q(n13841) );
  AND2X1 U14040 ( .IN1(n13844), .IN2(n13845), .Q(n13083) );
  INVX0 U14041 ( .INP(n13846), .ZN(n13845) );
  AND2X1 U14042 ( .IN1(n13847), .IN2(n13848), .Q(n13846) );
  OR2X1 U14043 ( .IN1(n13848), .IN2(n13847), .Q(n13844) );
  OR2X1 U14044 ( .IN1(n13849), .IN2(n13850), .Q(n13847) );
  AND2X1 U14045 ( .IN1(n3661), .IN2(WX5877), .Q(n13850) );
  INVX0 U14046 ( .INP(n13851), .ZN(n13849) );
  OR2X1 U14047 ( .IN1(WX5877), .IN2(n3661), .Q(n13851) );
  AND2X1 U14048 ( .IN1(n13852), .IN2(n13853), .Q(n13848) );
  OR2X1 U14049 ( .IN1(WX6069), .IN2(test_so51), .Q(n13853) );
  OR2X1 U14050 ( .IN1(n9923), .IN2(n9673), .Q(n13852) );
  OR2X1 U14051 ( .IN1(n13854), .IN2(n13855), .Q(WX4581) );
  OR2X1 U14052 ( .IN1(n13856), .IN2(n13857), .Q(n13855) );
  AND2X1 U14053 ( .IN1(n10027), .IN2(CRC_OUT_6_2), .Q(n13857) );
  AND2X1 U14054 ( .IN1(n760), .IN2(n10001), .Q(n13856) );
  INVX0 U14055 ( .INP(n13858), .ZN(n760) );
  OR2X1 U14056 ( .IN1(n10639), .IN2(n3943), .Q(n13858) );
  OR2X1 U14057 ( .IN1(n13859), .IN2(n13860), .Q(n13854) );
  AND2X1 U14058 ( .IN1(n9992), .IN2(n13861), .Q(n13860) );
  AND2X1 U14059 ( .IN1(n10078), .IN2(n13100), .Q(n13859) );
  OR2X1 U14060 ( .IN1(n13862), .IN2(n13863), .Q(n13100) );
  INVX0 U14061 ( .INP(n13864), .ZN(n13863) );
  OR2X1 U14062 ( .IN1(n13865), .IN2(n13866), .Q(n13864) );
  AND2X1 U14063 ( .IN1(n13866), .IN2(n13865), .Q(n13862) );
  AND2X1 U14064 ( .IN1(n13867), .IN2(n13868), .Q(n13865) );
  OR2X1 U14065 ( .IN1(WX5939), .IN2(n9394), .Q(n13868) );
  OR2X1 U14066 ( .IN1(WX5875), .IN2(n3663), .Q(n13867) );
  OR2X1 U14067 ( .IN1(n13869), .IN2(n13870), .Q(n13866) );
  AND2X1 U14068 ( .IN1(n9395), .IN2(WX6067), .Q(n13870) );
  AND2X1 U14069 ( .IN1(n9672), .IN2(WX6003), .Q(n13869) );
  OR2X1 U14070 ( .IN1(n13871), .IN2(n13872), .Q(WX4579) );
  OR2X1 U14071 ( .IN1(n13873), .IN2(n13874), .Q(n13872) );
  AND2X1 U14072 ( .IN1(n10028), .IN2(CRC_OUT_6_3), .Q(n13874) );
  AND2X1 U14073 ( .IN1(n759), .IN2(n10001), .Q(n13873) );
  INVX0 U14074 ( .INP(n13875), .ZN(n759) );
  OR2X1 U14075 ( .IN1(n10639), .IN2(n3944), .Q(n13875) );
  OR2X1 U14076 ( .IN1(n13876), .IN2(n13877), .Q(n13871) );
  AND2X1 U14077 ( .IN1(n9992), .IN2(n13878), .Q(n13877) );
  AND2X1 U14078 ( .IN1(n13117), .IN2(n10056), .Q(n13876) );
  AND2X1 U14079 ( .IN1(n13879), .IN2(n13880), .Q(n13117) );
  INVX0 U14080 ( .INP(n13881), .ZN(n13880) );
  AND2X1 U14081 ( .IN1(n13882), .IN2(n13883), .Q(n13881) );
  OR2X1 U14082 ( .IN1(n13883), .IN2(n13882), .Q(n13879) );
  OR2X1 U14083 ( .IN1(n13884), .IN2(n13885), .Q(n13882) );
  AND2X1 U14084 ( .IN1(n9396), .IN2(WX6001), .Q(n13885) );
  INVX0 U14085 ( .INP(n13886), .ZN(n13884) );
  OR2X1 U14086 ( .IN1(WX6001), .IN2(n9396), .Q(n13886) );
  AND2X1 U14087 ( .IN1(n13887), .IN2(n13888), .Q(n13883) );
  OR2X1 U14088 ( .IN1(WX6065), .IN2(test_so49), .Q(n13888) );
  OR2X1 U14089 ( .IN1(n9924), .IN2(n9671), .Q(n13887) );
  OR2X1 U14090 ( .IN1(n13889), .IN2(n13890), .Q(WX4577) );
  OR2X1 U14091 ( .IN1(n13891), .IN2(n13892), .Q(n13890) );
  AND2X1 U14092 ( .IN1(n10028), .IN2(CRC_OUT_6_4), .Q(n13892) );
  AND2X1 U14093 ( .IN1(n758), .IN2(n10001), .Q(n13891) );
  INVX0 U14094 ( .INP(n13893), .ZN(n758) );
  OR2X1 U14095 ( .IN1(n10638), .IN2(n3945), .Q(n13893) );
  OR2X1 U14096 ( .IN1(n13894), .IN2(n13895), .Q(n13889) );
  AND2X1 U14097 ( .IN1(n9992), .IN2(n13896), .Q(n13895) );
  AND2X1 U14098 ( .IN1(n10063), .IN2(n13134), .Q(n13894) );
  OR2X1 U14099 ( .IN1(n13897), .IN2(n13898), .Q(n13134) );
  INVX0 U14100 ( .INP(n13899), .ZN(n13898) );
  OR2X1 U14101 ( .IN1(n13900), .IN2(n13901), .Q(n13899) );
  AND2X1 U14102 ( .IN1(n13901), .IN2(n13900), .Q(n13897) );
  AND2X1 U14103 ( .IN1(n13902), .IN2(n13903), .Q(n13900) );
  OR2X1 U14104 ( .IN1(WX5935), .IN2(n9398), .Q(n13903) );
  OR2X1 U14105 ( .IN1(WX5871), .IN2(n3667), .Q(n13902) );
  OR2X1 U14106 ( .IN1(n13904), .IN2(n13905), .Q(n13901) );
  AND2X1 U14107 ( .IN1(n9399), .IN2(WX6063), .Q(n13905) );
  AND2X1 U14108 ( .IN1(n9524), .IN2(WX5999), .Q(n13904) );
  OR2X1 U14109 ( .IN1(n13906), .IN2(n13907), .Q(WX4575) );
  OR2X1 U14110 ( .IN1(n13908), .IN2(n13909), .Q(n13907) );
  AND2X1 U14111 ( .IN1(test_so42), .IN2(n10026), .Q(n13909) );
  AND2X1 U14112 ( .IN1(n757), .IN2(n10001), .Q(n13908) );
  INVX0 U14113 ( .INP(n13910), .ZN(n757) );
  OR2X1 U14114 ( .IN1(n10638), .IN2(n3946), .Q(n13910) );
  OR2X1 U14115 ( .IN1(n13911), .IN2(n13912), .Q(n13906) );
  AND2X1 U14116 ( .IN1(n9992), .IN2(n13913), .Q(n13912) );
  AND2X1 U14117 ( .IN1(n13152), .IN2(n10056), .Q(n13911) );
  AND2X1 U14118 ( .IN1(n13914), .IN2(n13915), .Q(n13152) );
  INVX0 U14119 ( .INP(n13916), .ZN(n13915) );
  AND2X1 U14120 ( .IN1(n13917), .IN2(n13918), .Q(n13916) );
  OR2X1 U14121 ( .IN1(n13918), .IN2(n13917), .Q(n13914) );
  OR2X1 U14122 ( .IN1(n13919), .IN2(n13920), .Q(n13917) );
  AND2X1 U14123 ( .IN1(n3669), .IN2(WX5997), .Q(n13920) );
  INVX0 U14124 ( .INP(n13921), .ZN(n13919) );
  OR2X1 U14125 ( .IN1(WX5997), .IN2(n3669), .Q(n13921) );
  AND2X1 U14126 ( .IN1(n13922), .IN2(n13923), .Q(n13918) );
  OR2X1 U14127 ( .IN1(WX6061), .IN2(test_so47), .Q(n13923) );
  OR2X1 U14128 ( .IN1(n9925), .IN2(n9670), .Q(n13922) );
  OR2X1 U14129 ( .IN1(n13924), .IN2(n13925), .Q(WX4573) );
  OR2X1 U14130 ( .IN1(n13926), .IN2(n13927), .Q(n13925) );
  AND2X1 U14131 ( .IN1(n10028), .IN2(CRC_OUT_6_6), .Q(n13927) );
  AND2X1 U14132 ( .IN1(n756), .IN2(n10001), .Q(n13926) );
  INVX0 U14133 ( .INP(n13928), .ZN(n756) );
  OR2X1 U14134 ( .IN1(n10638), .IN2(n3947), .Q(n13928) );
  OR2X1 U14135 ( .IN1(n13929), .IN2(n13930), .Q(n13924) );
  AND2X1 U14136 ( .IN1(n9992), .IN2(n13931), .Q(n13930) );
  AND2X1 U14137 ( .IN1(n10065), .IN2(n13169), .Q(n13929) );
  OR2X1 U14138 ( .IN1(n13932), .IN2(n13933), .Q(n13169) );
  INVX0 U14139 ( .INP(n13934), .ZN(n13933) );
  OR2X1 U14140 ( .IN1(n13935), .IN2(n13936), .Q(n13934) );
  AND2X1 U14141 ( .IN1(n13936), .IN2(n13935), .Q(n13932) );
  AND2X1 U14142 ( .IN1(n13937), .IN2(n13938), .Q(n13935) );
  OR2X1 U14143 ( .IN1(WX5931), .IN2(n9401), .Q(n13938) );
  OR2X1 U14144 ( .IN1(WX5867), .IN2(n3671), .Q(n13937) );
  OR2X1 U14145 ( .IN1(n13939), .IN2(n13940), .Q(n13936) );
  AND2X1 U14146 ( .IN1(n9402), .IN2(WX6059), .Q(n13940) );
  AND2X1 U14147 ( .IN1(n9669), .IN2(WX5995), .Q(n13939) );
  OR2X1 U14148 ( .IN1(n13941), .IN2(n13942), .Q(WX4571) );
  OR2X1 U14149 ( .IN1(n13943), .IN2(n13944), .Q(n13942) );
  AND2X1 U14150 ( .IN1(n10028), .IN2(CRC_OUT_6_7), .Q(n13944) );
  AND2X1 U14151 ( .IN1(n755), .IN2(n10001), .Q(n13943) );
  INVX0 U14152 ( .INP(n13945), .ZN(n755) );
  OR2X1 U14153 ( .IN1(n10638), .IN2(n3948), .Q(n13945) );
  OR2X1 U14154 ( .IN1(n13946), .IN2(n13947), .Q(n13941) );
  AND2X1 U14155 ( .IN1(n9991), .IN2(n13948), .Q(n13947) );
  AND2X1 U14156 ( .IN1(n10063), .IN2(n13187), .Q(n13946) );
  OR2X1 U14157 ( .IN1(n13949), .IN2(n13950), .Q(n13187) );
  INVX0 U14158 ( .INP(n13951), .ZN(n13950) );
  OR2X1 U14159 ( .IN1(n13952), .IN2(n13953), .Q(n13951) );
  AND2X1 U14160 ( .IN1(n13953), .IN2(n13952), .Q(n13949) );
  AND2X1 U14161 ( .IN1(n13954), .IN2(n13955), .Q(n13952) );
  OR2X1 U14162 ( .IN1(WX5929), .IN2(n9403), .Q(n13955) );
  OR2X1 U14163 ( .IN1(WX5865), .IN2(n3673), .Q(n13954) );
  OR2X1 U14164 ( .IN1(n13956), .IN2(n13957), .Q(n13953) );
  AND2X1 U14165 ( .IN1(n9404), .IN2(WX6057), .Q(n13957) );
  AND2X1 U14166 ( .IN1(n9668), .IN2(WX5993), .Q(n13956) );
  OR2X1 U14167 ( .IN1(n13958), .IN2(n13959), .Q(WX4569) );
  OR2X1 U14168 ( .IN1(n13960), .IN2(n13961), .Q(n13959) );
  AND2X1 U14169 ( .IN1(n10030), .IN2(CRC_OUT_6_8), .Q(n13961) );
  AND2X1 U14170 ( .IN1(n754), .IN2(n10002), .Q(n13960) );
  INVX0 U14171 ( .INP(n13962), .ZN(n754) );
  OR2X1 U14172 ( .IN1(n10638), .IN2(n3949), .Q(n13962) );
  OR2X1 U14173 ( .IN1(n13963), .IN2(n13964), .Q(n13958) );
  AND2X1 U14174 ( .IN1(n9991), .IN2(n13965), .Q(n13964) );
  AND2X1 U14175 ( .IN1(n10063), .IN2(n13204), .Q(n13963) );
  OR2X1 U14176 ( .IN1(n13966), .IN2(n13967), .Q(n13204) );
  INVX0 U14177 ( .INP(n13968), .ZN(n13967) );
  OR2X1 U14178 ( .IN1(n13969), .IN2(n13970), .Q(n13968) );
  AND2X1 U14179 ( .IN1(n13970), .IN2(n13969), .Q(n13966) );
  AND2X1 U14180 ( .IN1(n13971), .IN2(n13972), .Q(n13969) );
  OR2X1 U14181 ( .IN1(WX5927), .IN2(n9405), .Q(n13972) );
  OR2X1 U14182 ( .IN1(WX5863), .IN2(n3675), .Q(n13971) );
  OR2X1 U14183 ( .IN1(n13973), .IN2(n13974), .Q(n13970) );
  AND2X1 U14184 ( .IN1(n9406), .IN2(WX6055), .Q(n13974) );
  AND2X1 U14185 ( .IN1(n9667), .IN2(WX5991), .Q(n13973) );
  OR2X1 U14186 ( .IN1(n13975), .IN2(n13976), .Q(WX4567) );
  OR2X1 U14187 ( .IN1(n13977), .IN2(n13978), .Q(n13976) );
  AND2X1 U14188 ( .IN1(n10028), .IN2(CRC_OUT_6_9), .Q(n13978) );
  AND2X1 U14189 ( .IN1(n753), .IN2(n10002), .Q(n13977) );
  INVX0 U14190 ( .INP(n13979), .ZN(n753) );
  OR2X1 U14191 ( .IN1(n10638), .IN2(n3950), .Q(n13979) );
  OR2X1 U14192 ( .IN1(n13980), .IN2(n13981), .Q(n13975) );
  AND2X1 U14193 ( .IN1(n9991), .IN2(n13982), .Q(n13981) );
  AND2X1 U14194 ( .IN1(n10064), .IN2(n13222), .Q(n13980) );
  OR2X1 U14195 ( .IN1(n13983), .IN2(n13984), .Q(n13222) );
  INVX0 U14196 ( .INP(n13985), .ZN(n13984) );
  OR2X1 U14197 ( .IN1(n13986), .IN2(n13987), .Q(n13985) );
  AND2X1 U14198 ( .IN1(n13987), .IN2(n13986), .Q(n13983) );
  AND2X1 U14199 ( .IN1(n13988), .IN2(n13989), .Q(n13986) );
  OR2X1 U14200 ( .IN1(WX5925), .IN2(n9407), .Q(n13989) );
  OR2X1 U14201 ( .IN1(WX5861), .IN2(n3677), .Q(n13988) );
  OR2X1 U14202 ( .IN1(n13990), .IN2(n13991), .Q(n13987) );
  AND2X1 U14203 ( .IN1(n9408), .IN2(WX6053), .Q(n13991) );
  AND2X1 U14204 ( .IN1(n9666), .IN2(WX5989), .Q(n13990) );
  OR2X1 U14205 ( .IN1(n13992), .IN2(n13993), .Q(WX4565) );
  OR2X1 U14206 ( .IN1(n13994), .IN2(n13995), .Q(n13993) );
  AND2X1 U14207 ( .IN1(n10029), .IN2(CRC_OUT_6_10), .Q(n13995) );
  AND2X1 U14208 ( .IN1(n752), .IN2(n10002), .Q(n13994) );
  INVX0 U14209 ( .INP(n13996), .ZN(n752) );
  OR2X1 U14210 ( .IN1(n10638), .IN2(n3951), .Q(n13996) );
  OR2X1 U14211 ( .IN1(n13997), .IN2(n13998), .Q(n13992) );
  AND2X1 U14212 ( .IN1(n9991), .IN2(n13999), .Q(n13998) );
  AND2X1 U14213 ( .IN1(n10064), .IN2(n13239), .Q(n13997) );
  OR2X1 U14214 ( .IN1(n14000), .IN2(n14001), .Q(n13239) );
  INVX0 U14215 ( .INP(n14002), .ZN(n14001) );
  OR2X1 U14216 ( .IN1(n14003), .IN2(n14004), .Q(n14002) );
  AND2X1 U14217 ( .IN1(n14004), .IN2(n14003), .Q(n14000) );
  AND2X1 U14218 ( .IN1(n14005), .IN2(n14006), .Q(n14003) );
  OR2X1 U14219 ( .IN1(WX5923), .IN2(n9409), .Q(n14006) );
  OR2X1 U14220 ( .IN1(WX5859), .IN2(n3679), .Q(n14005) );
  OR2X1 U14221 ( .IN1(n14007), .IN2(n14008), .Q(n14004) );
  AND2X1 U14222 ( .IN1(n9410), .IN2(WX6051), .Q(n14008) );
  AND2X1 U14223 ( .IN1(n9665), .IN2(WX5987), .Q(n14007) );
  OR2X1 U14224 ( .IN1(n14009), .IN2(n14010), .Q(WX4563) );
  OR2X1 U14225 ( .IN1(n14011), .IN2(n14012), .Q(n14010) );
  AND2X1 U14226 ( .IN1(n10028), .IN2(CRC_OUT_6_11), .Q(n14012) );
  AND2X1 U14227 ( .IN1(n751), .IN2(n10002), .Q(n14011) );
  INVX0 U14228 ( .INP(n14013), .ZN(n751) );
  OR2X1 U14229 ( .IN1(n10638), .IN2(n3952), .Q(n14013) );
  OR2X1 U14230 ( .IN1(n14014), .IN2(n14015), .Q(n14009) );
  AND2X1 U14231 ( .IN1(n14016), .IN2(n9977), .Q(n14015) );
  AND2X1 U14232 ( .IN1(n10063), .IN2(n13257), .Q(n14014) );
  OR2X1 U14233 ( .IN1(n14017), .IN2(n14018), .Q(n13257) );
  INVX0 U14234 ( .INP(n14019), .ZN(n14018) );
  OR2X1 U14235 ( .IN1(n14020), .IN2(n14021), .Q(n14019) );
  AND2X1 U14236 ( .IN1(n14021), .IN2(n14020), .Q(n14017) );
  AND2X1 U14237 ( .IN1(n14022), .IN2(n14023), .Q(n14020) );
  OR2X1 U14238 ( .IN1(WX5921), .IN2(n9411), .Q(n14023) );
  OR2X1 U14239 ( .IN1(WX5857), .IN2(n3681), .Q(n14022) );
  OR2X1 U14240 ( .IN1(n14024), .IN2(n14025), .Q(n14021) );
  AND2X1 U14241 ( .IN1(n9412), .IN2(WX6049), .Q(n14025) );
  AND2X1 U14242 ( .IN1(n9523), .IN2(WX5985), .Q(n14024) );
  OR2X1 U14243 ( .IN1(n14026), .IN2(n14027), .Q(WX4561) );
  OR2X1 U14244 ( .IN1(n14028), .IN2(n14029), .Q(n14027) );
  AND2X1 U14245 ( .IN1(n10029), .IN2(CRC_OUT_6_12), .Q(n14029) );
  AND2X1 U14246 ( .IN1(n750), .IN2(n10002), .Q(n14028) );
  INVX0 U14247 ( .INP(n14030), .ZN(n750) );
  OR2X1 U14248 ( .IN1(n10638), .IN2(n3953), .Q(n14030) );
  OR2X1 U14249 ( .IN1(n14031), .IN2(n14032), .Q(n14026) );
  AND2X1 U14250 ( .IN1(n9991), .IN2(n14033), .Q(n14032) );
  AND2X1 U14251 ( .IN1(n10064), .IN2(n13274), .Q(n14031) );
  OR2X1 U14252 ( .IN1(n14034), .IN2(n14035), .Q(n13274) );
  INVX0 U14253 ( .INP(n14036), .ZN(n14035) );
  OR2X1 U14254 ( .IN1(n14037), .IN2(n14038), .Q(n14036) );
  AND2X1 U14255 ( .IN1(n14038), .IN2(n14037), .Q(n14034) );
  AND2X1 U14256 ( .IN1(n14039), .IN2(n14040), .Q(n14037) );
  OR2X1 U14257 ( .IN1(WX5919), .IN2(n9413), .Q(n14040) );
  OR2X1 U14258 ( .IN1(WX5855), .IN2(n3683), .Q(n14039) );
  OR2X1 U14259 ( .IN1(n14041), .IN2(n14042), .Q(n14038) );
  AND2X1 U14260 ( .IN1(n9414), .IN2(WX6047), .Q(n14042) );
  AND2X1 U14261 ( .IN1(n9664), .IN2(WX5983), .Q(n14041) );
  OR2X1 U14262 ( .IN1(n14043), .IN2(n14044), .Q(WX4559) );
  OR2X1 U14263 ( .IN1(n14045), .IN2(n14046), .Q(n14044) );
  AND2X1 U14264 ( .IN1(n10028), .IN2(CRC_OUT_6_13), .Q(n14046) );
  AND2X1 U14265 ( .IN1(n749), .IN2(n10002), .Q(n14045) );
  INVX0 U14266 ( .INP(n14047), .ZN(n749) );
  OR2X1 U14267 ( .IN1(n10638), .IN2(n3954), .Q(n14047) );
  OR2X1 U14268 ( .IN1(n14048), .IN2(n14049), .Q(n14043) );
  AND2X1 U14269 ( .IN1(n14050), .IN2(n9977), .Q(n14049) );
  AND2X1 U14270 ( .IN1(n10064), .IN2(n13291), .Q(n14048) );
  OR2X1 U14271 ( .IN1(n14051), .IN2(n14052), .Q(n13291) );
  INVX0 U14272 ( .INP(n14053), .ZN(n14052) );
  OR2X1 U14273 ( .IN1(n14054), .IN2(n14055), .Q(n14053) );
  AND2X1 U14274 ( .IN1(n14055), .IN2(n14054), .Q(n14051) );
  AND2X1 U14275 ( .IN1(n14056), .IN2(n14057), .Q(n14054) );
  OR2X1 U14276 ( .IN1(WX5917), .IN2(n9415), .Q(n14057) );
  OR2X1 U14277 ( .IN1(WX5853), .IN2(n3685), .Q(n14056) );
  OR2X1 U14278 ( .IN1(n14058), .IN2(n14059), .Q(n14055) );
  AND2X1 U14279 ( .IN1(n9416), .IN2(WX6045), .Q(n14059) );
  AND2X1 U14280 ( .IN1(n9663), .IN2(WX5981), .Q(n14058) );
  OR2X1 U14281 ( .IN1(n14060), .IN2(n14061), .Q(WX4557) );
  OR2X1 U14282 ( .IN1(n14062), .IN2(n14063), .Q(n14061) );
  AND2X1 U14283 ( .IN1(n10030), .IN2(CRC_OUT_6_14), .Q(n14063) );
  AND2X1 U14284 ( .IN1(n748), .IN2(n10002), .Q(n14062) );
  INVX0 U14285 ( .INP(n14064), .ZN(n748) );
  OR2X1 U14286 ( .IN1(n10638), .IN2(n3955), .Q(n14064) );
  OR2X1 U14287 ( .IN1(n14065), .IN2(n14066), .Q(n14060) );
  AND2X1 U14288 ( .IN1(n9991), .IN2(n14067), .Q(n14066) );
  AND2X1 U14289 ( .IN1(n10063), .IN2(n13308), .Q(n14065) );
  OR2X1 U14290 ( .IN1(n14068), .IN2(n14069), .Q(n13308) );
  INVX0 U14291 ( .INP(n14070), .ZN(n14069) );
  OR2X1 U14292 ( .IN1(n14071), .IN2(n14072), .Q(n14070) );
  AND2X1 U14293 ( .IN1(n14072), .IN2(n14071), .Q(n14068) );
  AND2X1 U14294 ( .IN1(n14073), .IN2(n14074), .Q(n14071) );
  OR2X1 U14295 ( .IN1(WX5915), .IN2(n9417), .Q(n14074) );
  OR2X1 U14296 ( .IN1(WX5851), .IN2(n3687), .Q(n14073) );
  OR2X1 U14297 ( .IN1(n14075), .IN2(n14076), .Q(n14072) );
  AND2X1 U14298 ( .IN1(n9418), .IN2(WX6043), .Q(n14076) );
  AND2X1 U14299 ( .IN1(n9662), .IN2(WX5979), .Q(n14075) );
  OR2X1 U14300 ( .IN1(n14077), .IN2(n14078), .Q(WX4555) );
  OR2X1 U14301 ( .IN1(n14079), .IN2(n14080), .Q(n14078) );
  AND2X1 U14302 ( .IN1(n10028), .IN2(CRC_OUT_6_15), .Q(n14080) );
  AND2X1 U14303 ( .IN1(n747), .IN2(n10002), .Q(n14079) );
  INVX0 U14304 ( .INP(n14081), .ZN(n747) );
  OR2X1 U14305 ( .IN1(n10638), .IN2(n3956), .Q(n14081) );
  OR2X1 U14306 ( .IN1(n14082), .IN2(n14083), .Q(n14077) );
  AND2X1 U14307 ( .IN1(n14084), .IN2(n9975), .Q(n14083) );
  AND2X1 U14308 ( .IN1(n10064), .IN2(n13325), .Q(n14082) );
  OR2X1 U14309 ( .IN1(n14085), .IN2(n14086), .Q(n13325) );
  INVX0 U14310 ( .INP(n14087), .ZN(n14086) );
  OR2X1 U14311 ( .IN1(n14088), .IN2(n14089), .Q(n14087) );
  AND2X1 U14312 ( .IN1(n14089), .IN2(n14088), .Q(n14085) );
  AND2X1 U14313 ( .IN1(n14090), .IN2(n14091), .Q(n14088) );
  OR2X1 U14314 ( .IN1(WX5913), .IN2(n9419), .Q(n14091) );
  OR2X1 U14315 ( .IN1(WX5849), .IN2(n3689), .Q(n14090) );
  OR2X1 U14316 ( .IN1(n14092), .IN2(n14093), .Q(n14089) );
  AND2X1 U14317 ( .IN1(n9420), .IN2(WX6041), .Q(n14093) );
  AND2X1 U14318 ( .IN1(n9661), .IN2(WX5977), .Q(n14092) );
  OR2X1 U14319 ( .IN1(n14094), .IN2(n14095), .Q(WX4553) );
  OR2X1 U14320 ( .IN1(n14096), .IN2(n14097), .Q(n14095) );
  AND2X1 U14321 ( .IN1(n10029), .IN2(CRC_OUT_6_16), .Q(n14097) );
  AND2X1 U14322 ( .IN1(n746), .IN2(n10002), .Q(n14096) );
  INVX0 U14323 ( .INP(n14098), .ZN(n746) );
  OR2X1 U14324 ( .IN1(n10637), .IN2(n3957), .Q(n14098) );
  OR2X1 U14325 ( .IN1(n14099), .IN2(n14100), .Q(n14094) );
  AND2X1 U14326 ( .IN1(n9991), .IN2(n14101), .Q(n14100) );
  AND2X1 U14327 ( .IN1(n13342), .IN2(n10056), .Q(n14099) );
  AND2X1 U14328 ( .IN1(n14102), .IN2(n14103), .Q(n13342) );
  INVX0 U14329 ( .INP(n14104), .ZN(n14103) );
  AND2X1 U14330 ( .IN1(n14105), .IN2(n14106), .Q(n14104) );
  OR2X1 U14331 ( .IN1(n14106), .IN2(n14105), .Q(n14102) );
  OR2X1 U14332 ( .IN1(n14107), .IN2(n14108), .Q(n14105) );
  AND2X1 U14333 ( .IN1(n10522), .IN2(WX5911), .Q(n14108) );
  AND2X1 U14334 ( .IN1(n9156), .IN2(n10542), .Q(n14107) );
  AND2X1 U14335 ( .IN1(n14109), .IN2(n14110), .Q(n14106) );
  INVX0 U14336 ( .INP(n14111), .ZN(n14110) );
  AND2X1 U14337 ( .IN1(n14112), .IN2(WX5975), .Q(n14111) );
  OR2X1 U14338 ( .IN1(WX5975), .IN2(n14112), .Q(n14109) );
  OR2X1 U14339 ( .IN1(n14113), .IN2(n14114), .Q(n14112) );
  AND2X1 U14340 ( .IN1(n17927), .IN2(n9888), .Q(n14114) );
  AND2X1 U14341 ( .IN1(test_so52), .IN2(n8479), .Q(n14113) );
  OR2X1 U14342 ( .IN1(n14115), .IN2(n14116), .Q(WX4551) );
  OR2X1 U14343 ( .IN1(n14117), .IN2(n14118), .Q(n14116) );
  AND2X1 U14344 ( .IN1(n10029), .IN2(CRC_OUT_6_17), .Q(n14118) );
  AND2X1 U14345 ( .IN1(n745), .IN2(n10002), .Q(n14117) );
  INVX0 U14346 ( .INP(n14119), .ZN(n745) );
  OR2X1 U14347 ( .IN1(n10637), .IN2(n3958), .Q(n14119) );
  OR2X1 U14348 ( .IN1(n14120), .IN2(n14121), .Q(n14115) );
  AND2X1 U14349 ( .IN1(n14122), .IN2(n9975), .Q(n14121) );
  AND2X1 U14350 ( .IN1(n10063), .IN2(n13366), .Q(n14120) );
  OR2X1 U14351 ( .IN1(n14123), .IN2(n14124), .Q(n13366) );
  INVX0 U14352 ( .INP(n14125), .ZN(n14124) );
  OR2X1 U14353 ( .IN1(n14126), .IN2(n14127), .Q(n14125) );
  AND2X1 U14354 ( .IN1(n14127), .IN2(n14126), .Q(n14123) );
  INVX0 U14355 ( .INP(n14128), .ZN(n14126) );
  OR2X1 U14356 ( .IN1(n14129), .IN2(n14130), .Q(n14128) );
  AND2X1 U14357 ( .IN1(n10522), .IN2(n8480), .Q(n14130) );
  AND2X1 U14358 ( .IN1(n17928), .IN2(n10542), .Q(n14129) );
  OR2X1 U14359 ( .IN1(n14131), .IN2(n14132), .Q(n14127) );
  AND2X1 U14360 ( .IN1(n9660), .IN2(n14133), .Q(n14132) );
  AND2X1 U14361 ( .IN1(n14134), .IN2(n14135), .Q(n14133) );
  OR2X1 U14362 ( .IN1(n9158), .IN2(WX5973), .Q(n14135) );
  OR2X1 U14363 ( .IN1(n9159), .IN2(WX5909), .Q(n14134) );
  AND2X1 U14364 ( .IN1(n14136), .IN2(WX6037), .Q(n14131) );
  OR2X1 U14365 ( .IN1(n14137), .IN2(n14138), .Q(n14136) );
  AND2X1 U14366 ( .IN1(n9158), .IN2(WX5973), .Q(n14138) );
  AND2X1 U14367 ( .IN1(n9159), .IN2(WX5909), .Q(n14137) );
  OR2X1 U14368 ( .IN1(n14139), .IN2(n14140), .Q(WX4549) );
  OR2X1 U14369 ( .IN1(n14141), .IN2(n14142), .Q(n14140) );
  AND2X1 U14370 ( .IN1(n10029), .IN2(CRC_OUT_6_18), .Q(n14142) );
  AND2X1 U14371 ( .IN1(n744), .IN2(n10002), .Q(n14141) );
  INVX0 U14372 ( .INP(n14143), .ZN(n744) );
  OR2X1 U14373 ( .IN1(n10637), .IN2(n3959), .Q(n14143) );
  OR2X1 U14374 ( .IN1(n14144), .IN2(n14145), .Q(n14139) );
  AND2X1 U14375 ( .IN1(n9991), .IN2(n14146), .Q(n14145) );
  AND2X1 U14376 ( .IN1(n13390), .IN2(n10059), .Q(n14144) );
  AND2X1 U14377 ( .IN1(n14147), .IN2(n14148), .Q(n13390) );
  INVX0 U14378 ( .INP(n14149), .ZN(n14148) );
  AND2X1 U14379 ( .IN1(n14150), .IN2(n14151), .Q(n14149) );
  OR2X1 U14380 ( .IN1(n14151), .IN2(n14150), .Q(n14147) );
  OR2X1 U14381 ( .IN1(n14152), .IN2(n14153), .Q(n14150) );
  AND2X1 U14382 ( .IN1(n10522), .IN2(WX5907), .Q(n14153) );
  AND2X1 U14383 ( .IN1(n9160), .IN2(n10542), .Q(n14152) );
  AND2X1 U14384 ( .IN1(n14154), .IN2(n14155), .Q(n14151) );
  OR2X1 U14385 ( .IN1(n14156), .IN2(n9659), .Q(n14155) );
  INVX0 U14386 ( .INP(n14157), .ZN(n14156) );
  OR2X1 U14387 ( .IN1(WX6035), .IN2(n14157), .Q(n14154) );
  OR2X1 U14388 ( .IN1(n14158), .IN2(n14159), .Q(n14157) );
  AND2X1 U14389 ( .IN1(n17929), .IN2(n9959), .Q(n14159) );
  AND2X1 U14390 ( .IN1(test_so50), .IN2(n8481), .Q(n14158) );
  OR2X1 U14391 ( .IN1(n14160), .IN2(n14161), .Q(WX4547) );
  OR2X1 U14392 ( .IN1(n14162), .IN2(n14163), .Q(n14161) );
  AND2X1 U14393 ( .IN1(n10029), .IN2(CRC_OUT_6_19), .Q(n14163) );
  AND2X1 U14394 ( .IN1(n743), .IN2(n10002), .Q(n14162) );
  INVX0 U14395 ( .INP(n14164), .ZN(n743) );
  OR2X1 U14396 ( .IN1(n10637), .IN2(n3960), .Q(n14164) );
  OR2X1 U14397 ( .IN1(n14165), .IN2(n14166), .Q(n14160) );
  AND2X1 U14398 ( .IN1(n9991), .IN2(n14167), .Q(n14166) );
  AND2X1 U14399 ( .IN1(n10063), .IN2(n13414), .Q(n14165) );
  OR2X1 U14400 ( .IN1(n14168), .IN2(n14169), .Q(n13414) );
  INVX0 U14401 ( .INP(n14170), .ZN(n14169) );
  OR2X1 U14402 ( .IN1(n14171), .IN2(n14172), .Q(n14170) );
  AND2X1 U14403 ( .IN1(n14172), .IN2(n14171), .Q(n14168) );
  INVX0 U14404 ( .INP(n14173), .ZN(n14171) );
  OR2X1 U14405 ( .IN1(n14174), .IN2(n14175), .Q(n14173) );
  AND2X1 U14406 ( .IN1(n10522), .IN2(n8482), .Q(n14175) );
  AND2X1 U14407 ( .IN1(n17930), .IN2(n10542), .Q(n14174) );
  OR2X1 U14408 ( .IN1(n14176), .IN2(n14177), .Q(n14172) );
  AND2X1 U14409 ( .IN1(n9658), .IN2(n14178), .Q(n14177) );
  AND2X1 U14410 ( .IN1(n14179), .IN2(n14180), .Q(n14178) );
  OR2X1 U14411 ( .IN1(n9161), .IN2(WX5969), .Q(n14180) );
  OR2X1 U14412 ( .IN1(n9162), .IN2(WX5905), .Q(n14179) );
  AND2X1 U14413 ( .IN1(n14181), .IN2(WX6033), .Q(n14176) );
  OR2X1 U14414 ( .IN1(n14182), .IN2(n14183), .Q(n14181) );
  AND2X1 U14415 ( .IN1(n9161), .IN2(WX5969), .Q(n14183) );
  AND2X1 U14416 ( .IN1(n9162), .IN2(WX5905), .Q(n14182) );
  OR2X1 U14417 ( .IN1(n14184), .IN2(n14185), .Q(WX4545) );
  OR2X1 U14418 ( .IN1(n14186), .IN2(n14187), .Q(n14185) );
  AND2X1 U14419 ( .IN1(n10029), .IN2(CRC_OUT_6_20), .Q(n14187) );
  AND2X1 U14420 ( .IN1(n742), .IN2(n10003), .Q(n14186) );
  INVX0 U14421 ( .INP(n14188), .ZN(n742) );
  OR2X1 U14422 ( .IN1(n10637), .IN2(n3961), .Q(n14188) );
  OR2X1 U14423 ( .IN1(n14189), .IN2(n14190), .Q(n14184) );
  AND2X1 U14424 ( .IN1(n9991), .IN2(n14191), .Q(n14190) );
  AND2X1 U14425 ( .IN1(n13438), .IN2(n10056), .Q(n14189) );
  AND2X1 U14426 ( .IN1(n14192), .IN2(n14193), .Q(n13438) );
  INVX0 U14427 ( .INP(n14194), .ZN(n14193) );
  AND2X1 U14428 ( .IN1(n14195), .IN2(n14196), .Q(n14194) );
  OR2X1 U14429 ( .IN1(n14196), .IN2(n14195), .Q(n14192) );
  OR2X1 U14430 ( .IN1(n14197), .IN2(n14198), .Q(n14195) );
  AND2X1 U14431 ( .IN1(n10522), .IN2(WX5967), .Q(n14198) );
  AND2X1 U14432 ( .IN1(n9163), .IN2(n10542), .Q(n14197) );
  AND2X1 U14433 ( .IN1(n14199), .IN2(n14200), .Q(n14196) );
  OR2X1 U14434 ( .IN1(n14201), .IN2(n9657), .Q(n14200) );
  INVX0 U14435 ( .INP(n14202), .ZN(n14201) );
  OR2X1 U14436 ( .IN1(WX6031), .IN2(n14202), .Q(n14199) );
  OR2X1 U14437 ( .IN1(n14203), .IN2(n14204), .Q(n14202) );
  AND2X1 U14438 ( .IN1(n17931), .IN2(n9960), .Q(n14204) );
  AND2X1 U14439 ( .IN1(test_so48), .IN2(n8483), .Q(n14203) );
  OR2X1 U14440 ( .IN1(n14205), .IN2(n14206), .Q(WX4543) );
  OR2X1 U14441 ( .IN1(n14207), .IN2(n14208), .Q(n14206) );
  AND2X1 U14442 ( .IN1(n10029), .IN2(CRC_OUT_6_21), .Q(n14208) );
  AND2X1 U14443 ( .IN1(n741), .IN2(n10003), .Q(n14207) );
  INVX0 U14444 ( .INP(n14209), .ZN(n741) );
  OR2X1 U14445 ( .IN1(n10637), .IN2(n3962), .Q(n14209) );
  OR2X1 U14446 ( .IN1(n14210), .IN2(n14211), .Q(n14205) );
  AND2X1 U14447 ( .IN1(n9991), .IN2(n14212), .Q(n14211) );
  AND2X1 U14448 ( .IN1(n10064), .IN2(n13462), .Q(n14210) );
  OR2X1 U14449 ( .IN1(n14213), .IN2(n14214), .Q(n13462) );
  INVX0 U14450 ( .INP(n14215), .ZN(n14214) );
  OR2X1 U14451 ( .IN1(n14216), .IN2(n14217), .Q(n14215) );
  AND2X1 U14452 ( .IN1(n14217), .IN2(n14216), .Q(n14213) );
  INVX0 U14453 ( .INP(n14218), .ZN(n14216) );
  OR2X1 U14454 ( .IN1(n14219), .IN2(n14220), .Q(n14218) );
  AND2X1 U14455 ( .IN1(n10522), .IN2(n8484), .Q(n14220) );
  AND2X1 U14456 ( .IN1(n17932), .IN2(n10542), .Q(n14219) );
  OR2X1 U14457 ( .IN1(n14221), .IN2(n14222), .Q(n14217) );
  AND2X1 U14458 ( .IN1(n9656), .IN2(n14223), .Q(n14222) );
  AND2X1 U14459 ( .IN1(n14224), .IN2(n14225), .Q(n14223) );
  OR2X1 U14460 ( .IN1(n9164), .IN2(WX5965), .Q(n14225) );
  OR2X1 U14461 ( .IN1(n9165), .IN2(WX5901), .Q(n14224) );
  AND2X1 U14462 ( .IN1(n14226), .IN2(WX6029), .Q(n14221) );
  OR2X1 U14463 ( .IN1(n14227), .IN2(n14228), .Q(n14226) );
  AND2X1 U14464 ( .IN1(n9164), .IN2(WX5965), .Q(n14228) );
  AND2X1 U14465 ( .IN1(n9165), .IN2(WX5901), .Q(n14227) );
  OR2X1 U14466 ( .IN1(n14229), .IN2(n14230), .Q(WX4541) );
  OR2X1 U14467 ( .IN1(n14231), .IN2(n14232), .Q(n14230) );
  AND2X1 U14468 ( .IN1(test_so43), .IN2(n10026), .Q(n14232) );
  AND2X1 U14469 ( .IN1(n740), .IN2(n10003), .Q(n14231) );
  INVX0 U14470 ( .INP(n14233), .ZN(n740) );
  OR2X1 U14471 ( .IN1(n10637), .IN2(n3963), .Q(n14233) );
  OR2X1 U14472 ( .IN1(n14234), .IN2(n14235), .Q(n14229) );
  AND2X1 U14473 ( .IN1(n9991), .IN2(n14236), .Q(n14235) );
  AND2X1 U14474 ( .IN1(n13483), .IN2(n10056), .Q(n14234) );
  AND2X1 U14475 ( .IN1(n14237), .IN2(n14238), .Q(n13483) );
  OR2X1 U14476 ( .IN1(n14239), .IN2(n14240), .Q(n14238) );
  INVX0 U14477 ( .INP(n14241), .ZN(n14239) );
  OR2X1 U14478 ( .IN1(n14242), .IN2(n14241), .Q(n14237) );
  OR2X1 U14479 ( .IN1(n14243), .IN2(n14244), .Q(n14241) );
  AND2X1 U14480 ( .IN1(n10523), .IN2(WX6027), .Q(n14244) );
  AND2X1 U14481 ( .IN1(n9655), .IN2(n10542), .Q(n14243) );
  INVX0 U14482 ( .INP(n14240), .ZN(n14242) );
  OR2X1 U14483 ( .IN1(n14245), .IN2(n14246), .Q(n14240) );
  AND2X1 U14484 ( .IN1(n9167), .IN2(n14247), .Q(n14246) );
  AND2X1 U14485 ( .IN1(n14248), .IN2(n14249), .Q(n14247) );
  OR2X1 U14486 ( .IN1(n9166), .IN2(n9892), .Q(n14249) );
  OR2X1 U14487 ( .IN1(test_so46), .IN2(WX5899), .Q(n14248) );
  AND2X1 U14488 ( .IN1(n14250), .IN2(WX5963), .Q(n14245) );
  OR2X1 U14489 ( .IN1(n14251), .IN2(n14252), .Q(n14250) );
  AND2X1 U14490 ( .IN1(n9166), .IN2(n9892), .Q(n14252) );
  AND2X1 U14491 ( .IN1(test_so46), .IN2(WX5899), .Q(n14251) );
  OR2X1 U14492 ( .IN1(n14253), .IN2(n14254), .Q(WX4539) );
  OR2X1 U14493 ( .IN1(n14255), .IN2(n14256), .Q(n14254) );
  AND2X1 U14494 ( .IN1(n10030), .IN2(CRC_OUT_6_23), .Q(n14256) );
  AND2X1 U14495 ( .IN1(n739), .IN2(n10003), .Q(n14255) );
  INVX0 U14496 ( .INP(n14257), .ZN(n739) );
  OR2X1 U14497 ( .IN1(n10637), .IN2(n3964), .Q(n14257) );
  OR2X1 U14498 ( .IN1(n14258), .IN2(n14259), .Q(n14253) );
  AND2X1 U14499 ( .IN1(n9991), .IN2(n14260), .Q(n14259) );
  AND2X1 U14500 ( .IN1(n10064), .IN2(n13507), .Q(n14258) );
  OR2X1 U14501 ( .IN1(n14261), .IN2(n14262), .Q(n13507) );
  INVX0 U14502 ( .INP(n14263), .ZN(n14262) );
  OR2X1 U14503 ( .IN1(n14264), .IN2(n14265), .Q(n14263) );
  AND2X1 U14504 ( .IN1(n14265), .IN2(n14264), .Q(n14261) );
  INVX0 U14505 ( .INP(n14266), .ZN(n14264) );
  OR2X1 U14506 ( .IN1(n14267), .IN2(n14268), .Q(n14266) );
  AND2X1 U14507 ( .IN1(n10523), .IN2(n8487), .Q(n14268) );
  AND2X1 U14508 ( .IN1(n17933), .IN2(n10542), .Q(n14267) );
  OR2X1 U14509 ( .IN1(n14269), .IN2(n14270), .Q(n14265) );
  AND2X1 U14510 ( .IN1(n9654), .IN2(n14271), .Q(n14270) );
  AND2X1 U14511 ( .IN1(n14272), .IN2(n14273), .Q(n14271) );
  OR2X1 U14512 ( .IN1(n9168), .IN2(WX5961), .Q(n14273) );
  OR2X1 U14513 ( .IN1(n9169), .IN2(WX5897), .Q(n14272) );
  AND2X1 U14514 ( .IN1(n14274), .IN2(WX6025), .Q(n14269) );
  OR2X1 U14515 ( .IN1(n14275), .IN2(n14276), .Q(n14274) );
  AND2X1 U14516 ( .IN1(n9168), .IN2(WX5961), .Q(n14276) );
  AND2X1 U14517 ( .IN1(n9169), .IN2(WX5897), .Q(n14275) );
  OR2X1 U14518 ( .IN1(n14277), .IN2(n14278), .Q(WX4537) );
  OR2X1 U14519 ( .IN1(n14279), .IN2(n14280), .Q(n14278) );
  AND2X1 U14520 ( .IN1(n10029), .IN2(CRC_OUT_6_24), .Q(n14280) );
  AND2X1 U14521 ( .IN1(n738), .IN2(n10003), .Q(n14279) );
  INVX0 U14522 ( .INP(n14281), .ZN(n738) );
  OR2X1 U14523 ( .IN1(n10637), .IN2(n3965), .Q(n14281) );
  OR2X1 U14524 ( .IN1(n14282), .IN2(n14283), .Q(n14277) );
  AND2X1 U14525 ( .IN1(n9990), .IN2(n14284), .Q(n14283) );
  AND2X1 U14526 ( .IN1(n10064), .IN2(n13528), .Q(n14282) );
  OR2X1 U14527 ( .IN1(n14285), .IN2(n14286), .Q(n13528) );
  INVX0 U14528 ( .INP(n14287), .ZN(n14286) );
  OR2X1 U14529 ( .IN1(n14288), .IN2(n14289), .Q(n14287) );
  AND2X1 U14530 ( .IN1(n14289), .IN2(n14288), .Q(n14285) );
  INVX0 U14531 ( .INP(n14290), .ZN(n14288) );
  OR2X1 U14532 ( .IN1(n14291), .IN2(n14292), .Q(n14290) );
  AND2X1 U14533 ( .IN1(n10523), .IN2(n8488), .Q(n14292) );
  AND2X1 U14534 ( .IN1(n17934), .IN2(n10542), .Q(n14291) );
  OR2X1 U14535 ( .IN1(n14293), .IN2(n14294), .Q(n14289) );
  AND2X1 U14536 ( .IN1(n9653), .IN2(n14295), .Q(n14294) );
  AND2X1 U14537 ( .IN1(n14296), .IN2(n14297), .Q(n14295) );
  OR2X1 U14538 ( .IN1(n9170), .IN2(WX5959), .Q(n14297) );
  OR2X1 U14539 ( .IN1(n9171), .IN2(WX5895), .Q(n14296) );
  AND2X1 U14540 ( .IN1(n14298), .IN2(WX6023), .Q(n14293) );
  OR2X1 U14541 ( .IN1(n14299), .IN2(n14300), .Q(n14298) );
  AND2X1 U14542 ( .IN1(n9170), .IN2(WX5959), .Q(n14300) );
  AND2X1 U14543 ( .IN1(n9171), .IN2(WX5895), .Q(n14299) );
  OR2X1 U14544 ( .IN1(n14301), .IN2(n14302), .Q(WX4535) );
  OR2X1 U14545 ( .IN1(n14303), .IN2(n14304), .Q(n14302) );
  AND2X1 U14546 ( .IN1(n10030), .IN2(CRC_OUT_6_25), .Q(n14304) );
  AND2X1 U14547 ( .IN1(n737), .IN2(n10003), .Q(n14303) );
  INVX0 U14548 ( .INP(n14305), .ZN(n737) );
  OR2X1 U14549 ( .IN1(n10637), .IN2(n3966), .Q(n14305) );
  OR2X1 U14550 ( .IN1(n14306), .IN2(n14307), .Q(n14301) );
  AND2X1 U14551 ( .IN1(n9990), .IN2(n14308), .Q(n14307) );
  AND2X1 U14552 ( .IN1(n10064), .IN2(n13552), .Q(n14306) );
  OR2X1 U14553 ( .IN1(n14309), .IN2(n14310), .Q(n13552) );
  INVX0 U14554 ( .INP(n14311), .ZN(n14310) );
  OR2X1 U14555 ( .IN1(n14312), .IN2(n14313), .Q(n14311) );
  AND2X1 U14556 ( .IN1(n14313), .IN2(n14312), .Q(n14309) );
  INVX0 U14557 ( .INP(n14314), .ZN(n14312) );
  OR2X1 U14558 ( .IN1(n14315), .IN2(n14316), .Q(n14314) );
  AND2X1 U14559 ( .IN1(n10523), .IN2(n8489), .Q(n14316) );
  AND2X1 U14560 ( .IN1(n17935), .IN2(n10542), .Q(n14315) );
  OR2X1 U14561 ( .IN1(n14317), .IN2(n14318), .Q(n14313) );
  AND2X1 U14562 ( .IN1(n9652), .IN2(n14319), .Q(n14318) );
  AND2X1 U14563 ( .IN1(n14320), .IN2(n14321), .Q(n14319) );
  OR2X1 U14564 ( .IN1(n9172), .IN2(WX5957), .Q(n14321) );
  OR2X1 U14565 ( .IN1(n9173), .IN2(WX5893), .Q(n14320) );
  AND2X1 U14566 ( .IN1(n14322), .IN2(WX6021), .Q(n14317) );
  OR2X1 U14567 ( .IN1(n14323), .IN2(n14324), .Q(n14322) );
  AND2X1 U14568 ( .IN1(n9172), .IN2(WX5957), .Q(n14324) );
  AND2X1 U14569 ( .IN1(n9173), .IN2(WX5893), .Q(n14323) );
  OR2X1 U14570 ( .IN1(n14325), .IN2(n14326), .Q(WX4533) );
  OR2X1 U14571 ( .IN1(n14327), .IN2(n14328), .Q(n14326) );
  AND2X1 U14572 ( .IN1(n10029), .IN2(CRC_OUT_6_26), .Q(n14328) );
  AND2X1 U14573 ( .IN1(n736), .IN2(n10003), .Q(n14327) );
  INVX0 U14574 ( .INP(n14329), .ZN(n736) );
  OR2X1 U14575 ( .IN1(n10637), .IN2(n3967), .Q(n14329) );
  OR2X1 U14576 ( .IN1(n14330), .IN2(n14331), .Q(n14325) );
  AND2X1 U14577 ( .IN1(n9990), .IN2(n14332), .Q(n14331) );
  AND2X1 U14578 ( .IN1(n10064), .IN2(n13573), .Q(n14330) );
  OR2X1 U14579 ( .IN1(n14333), .IN2(n14334), .Q(n13573) );
  INVX0 U14580 ( .INP(n14335), .ZN(n14334) );
  OR2X1 U14581 ( .IN1(n14336), .IN2(n14337), .Q(n14335) );
  AND2X1 U14582 ( .IN1(n14337), .IN2(n14336), .Q(n14333) );
  INVX0 U14583 ( .INP(n14338), .ZN(n14336) );
  OR2X1 U14584 ( .IN1(n14339), .IN2(n14340), .Q(n14338) );
  AND2X1 U14585 ( .IN1(n10523), .IN2(n8490), .Q(n14340) );
  AND2X1 U14586 ( .IN1(n17936), .IN2(n10542), .Q(n14339) );
  OR2X1 U14587 ( .IN1(n14341), .IN2(n14342), .Q(n14337) );
  AND2X1 U14588 ( .IN1(n9651), .IN2(n14343), .Q(n14342) );
  AND2X1 U14589 ( .IN1(n14344), .IN2(n14345), .Q(n14343) );
  OR2X1 U14590 ( .IN1(n9174), .IN2(WX5955), .Q(n14345) );
  OR2X1 U14591 ( .IN1(n9175), .IN2(WX5891), .Q(n14344) );
  AND2X1 U14592 ( .IN1(n14346), .IN2(WX6019), .Q(n14341) );
  OR2X1 U14593 ( .IN1(n14347), .IN2(n14348), .Q(n14346) );
  AND2X1 U14594 ( .IN1(n9174), .IN2(WX5955), .Q(n14348) );
  AND2X1 U14595 ( .IN1(n9175), .IN2(WX5891), .Q(n14347) );
  OR2X1 U14596 ( .IN1(n14349), .IN2(n14350), .Q(WX4531) );
  OR2X1 U14597 ( .IN1(n14351), .IN2(n14352), .Q(n14350) );
  AND2X1 U14598 ( .IN1(n10030), .IN2(CRC_OUT_6_27), .Q(n14352) );
  AND2X1 U14599 ( .IN1(n735), .IN2(n10003), .Q(n14351) );
  INVX0 U14600 ( .INP(n14353), .ZN(n735) );
  OR2X1 U14601 ( .IN1(n10637), .IN2(n3968), .Q(n14353) );
  OR2X1 U14602 ( .IN1(n14354), .IN2(n14355), .Q(n14349) );
  AND2X1 U14603 ( .IN1(n9990), .IN2(n14356), .Q(n14355) );
  AND2X1 U14604 ( .IN1(n10064), .IN2(n13597), .Q(n14354) );
  OR2X1 U14605 ( .IN1(n14357), .IN2(n14358), .Q(n13597) );
  INVX0 U14606 ( .INP(n14359), .ZN(n14358) );
  OR2X1 U14607 ( .IN1(n14360), .IN2(n14361), .Q(n14359) );
  AND2X1 U14608 ( .IN1(n14361), .IN2(n14360), .Q(n14357) );
  INVX0 U14609 ( .INP(n14362), .ZN(n14360) );
  OR2X1 U14610 ( .IN1(n14363), .IN2(n14364), .Q(n14362) );
  AND2X1 U14611 ( .IN1(n10523), .IN2(n8491), .Q(n14364) );
  AND2X1 U14612 ( .IN1(n17937), .IN2(n10542), .Q(n14363) );
  OR2X1 U14613 ( .IN1(n14365), .IN2(n14366), .Q(n14361) );
  AND2X1 U14614 ( .IN1(n9650), .IN2(n14367), .Q(n14366) );
  AND2X1 U14615 ( .IN1(n14368), .IN2(n14369), .Q(n14367) );
  OR2X1 U14616 ( .IN1(n9176), .IN2(WX5953), .Q(n14369) );
  OR2X1 U14617 ( .IN1(n9177), .IN2(WX5889), .Q(n14368) );
  AND2X1 U14618 ( .IN1(n14370), .IN2(WX6017), .Q(n14365) );
  OR2X1 U14619 ( .IN1(n14371), .IN2(n14372), .Q(n14370) );
  AND2X1 U14620 ( .IN1(n9176), .IN2(WX5953), .Q(n14372) );
  AND2X1 U14621 ( .IN1(n9177), .IN2(WX5889), .Q(n14371) );
  OR2X1 U14622 ( .IN1(n14373), .IN2(n14374), .Q(WX4529) );
  OR2X1 U14623 ( .IN1(n14375), .IN2(n14376), .Q(n14374) );
  AND2X1 U14624 ( .IN1(n10029), .IN2(CRC_OUT_6_28), .Q(n14376) );
  AND2X1 U14625 ( .IN1(n734), .IN2(n10003), .Q(n14375) );
  INVX0 U14626 ( .INP(n14377), .ZN(n734) );
  OR2X1 U14627 ( .IN1(n10636), .IN2(n3969), .Q(n14377) );
  OR2X1 U14628 ( .IN1(n14378), .IN2(n14379), .Q(n14373) );
  AND2X1 U14629 ( .IN1(n14380), .IN2(n9972), .Q(n14379) );
  AND2X1 U14630 ( .IN1(n10065), .IN2(n13621), .Q(n14378) );
  OR2X1 U14631 ( .IN1(n14381), .IN2(n14382), .Q(n13621) );
  INVX0 U14632 ( .INP(n14383), .ZN(n14382) );
  OR2X1 U14633 ( .IN1(n14384), .IN2(n14385), .Q(n14383) );
  AND2X1 U14634 ( .IN1(n14385), .IN2(n14384), .Q(n14381) );
  INVX0 U14635 ( .INP(n14386), .ZN(n14384) );
  OR2X1 U14636 ( .IN1(n14387), .IN2(n14388), .Q(n14386) );
  AND2X1 U14637 ( .IN1(n10523), .IN2(n8492), .Q(n14388) );
  AND2X1 U14638 ( .IN1(n17938), .IN2(n10542), .Q(n14387) );
  OR2X1 U14639 ( .IN1(n14389), .IN2(n14390), .Q(n14385) );
  AND2X1 U14640 ( .IN1(n9649), .IN2(n14391), .Q(n14390) );
  AND2X1 U14641 ( .IN1(n14392), .IN2(n14393), .Q(n14391) );
  OR2X1 U14642 ( .IN1(n9178), .IN2(WX5951), .Q(n14393) );
  OR2X1 U14643 ( .IN1(n9179), .IN2(WX5887), .Q(n14392) );
  AND2X1 U14644 ( .IN1(n14394), .IN2(WX6015), .Q(n14389) );
  OR2X1 U14645 ( .IN1(n14395), .IN2(n14396), .Q(n14394) );
  AND2X1 U14646 ( .IN1(n9178), .IN2(WX5951), .Q(n14396) );
  AND2X1 U14647 ( .IN1(n9179), .IN2(WX5887), .Q(n14395) );
  OR2X1 U14648 ( .IN1(n14397), .IN2(n14398), .Q(WX4527) );
  OR2X1 U14649 ( .IN1(n14399), .IN2(n14400), .Q(n14398) );
  AND2X1 U14650 ( .IN1(n10031), .IN2(CRC_OUT_6_29), .Q(n14400) );
  AND2X1 U14651 ( .IN1(n733), .IN2(n10003), .Q(n14399) );
  INVX0 U14652 ( .INP(n14401), .ZN(n733) );
  OR2X1 U14653 ( .IN1(n10636), .IN2(n3970), .Q(n14401) );
  OR2X1 U14654 ( .IN1(n14402), .IN2(n14403), .Q(n14397) );
  AND2X1 U14655 ( .IN1(n9990), .IN2(n14404), .Q(n14403) );
  AND2X1 U14656 ( .IN1(n10064), .IN2(n13645), .Q(n14402) );
  OR2X1 U14657 ( .IN1(n14405), .IN2(n14406), .Q(n13645) );
  INVX0 U14658 ( .INP(n14407), .ZN(n14406) );
  OR2X1 U14659 ( .IN1(n14408), .IN2(n14409), .Q(n14407) );
  AND2X1 U14660 ( .IN1(n14409), .IN2(n14408), .Q(n14405) );
  INVX0 U14661 ( .INP(n14410), .ZN(n14408) );
  OR2X1 U14662 ( .IN1(n14411), .IN2(n14412), .Q(n14410) );
  AND2X1 U14663 ( .IN1(n10523), .IN2(n8493), .Q(n14412) );
  AND2X1 U14664 ( .IN1(n17939), .IN2(n10542), .Q(n14411) );
  OR2X1 U14665 ( .IN1(n14413), .IN2(n14414), .Q(n14409) );
  AND2X1 U14666 ( .IN1(n9648), .IN2(n14415), .Q(n14414) );
  AND2X1 U14667 ( .IN1(n14416), .IN2(n14417), .Q(n14415) );
  OR2X1 U14668 ( .IN1(n9180), .IN2(WX5949), .Q(n14417) );
  OR2X1 U14669 ( .IN1(n9181), .IN2(WX5885), .Q(n14416) );
  AND2X1 U14670 ( .IN1(n14418), .IN2(WX6013), .Q(n14413) );
  OR2X1 U14671 ( .IN1(n14419), .IN2(n14420), .Q(n14418) );
  AND2X1 U14672 ( .IN1(n9180), .IN2(WX5949), .Q(n14420) );
  AND2X1 U14673 ( .IN1(n9181), .IN2(WX5885), .Q(n14419) );
  OR2X1 U14674 ( .IN1(n14421), .IN2(n14422), .Q(WX4525) );
  OR2X1 U14675 ( .IN1(n14423), .IN2(n14424), .Q(n14422) );
  AND2X1 U14676 ( .IN1(n10030), .IN2(CRC_OUT_6_30), .Q(n14424) );
  AND2X1 U14677 ( .IN1(n732), .IN2(n10003), .Q(n14423) );
  INVX0 U14678 ( .INP(n14425), .ZN(n732) );
  OR2X1 U14679 ( .IN1(n10636), .IN2(n3971), .Q(n14425) );
  OR2X1 U14680 ( .IN1(n14426), .IN2(n14427), .Q(n14421) );
  AND2X1 U14681 ( .IN1(n14428), .IN2(n9972), .Q(n14427) );
  AND2X1 U14682 ( .IN1(n10065), .IN2(n13669), .Q(n14426) );
  OR2X1 U14683 ( .IN1(n14429), .IN2(n14430), .Q(n13669) );
  INVX0 U14684 ( .INP(n14431), .ZN(n14430) );
  OR2X1 U14685 ( .IN1(n14432), .IN2(n14433), .Q(n14431) );
  AND2X1 U14686 ( .IN1(n14433), .IN2(n14432), .Q(n14429) );
  INVX0 U14687 ( .INP(n14434), .ZN(n14432) );
  OR2X1 U14688 ( .IN1(n14435), .IN2(n14436), .Q(n14434) );
  AND2X1 U14689 ( .IN1(n10523), .IN2(n8494), .Q(n14436) );
  AND2X1 U14690 ( .IN1(n17940), .IN2(n10541), .Q(n14435) );
  OR2X1 U14691 ( .IN1(n14437), .IN2(n14438), .Q(n14433) );
  AND2X1 U14692 ( .IN1(n9647), .IN2(n14439), .Q(n14438) );
  AND2X1 U14693 ( .IN1(n14440), .IN2(n14441), .Q(n14439) );
  OR2X1 U14694 ( .IN1(n9182), .IN2(WX5947), .Q(n14441) );
  OR2X1 U14695 ( .IN1(n9183), .IN2(WX5883), .Q(n14440) );
  AND2X1 U14696 ( .IN1(n14442), .IN2(WX6011), .Q(n14437) );
  OR2X1 U14697 ( .IN1(n14443), .IN2(n14444), .Q(n14442) );
  AND2X1 U14698 ( .IN1(n9182), .IN2(WX5947), .Q(n14444) );
  AND2X1 U14699 ( .IN1(n9183), .IN2(WX5883), .Q(n14443) );
  OR2X1 U14700 ( .IN1(n14445), .IN2(n14446), .Q(WX4523) );
  OR2X1 U14701 ( .IN1(n14447), .IN2(n14448), .Q(n14446) );
  AND2X1 U14702 ( .IN1(n2245), .IN2(WX4364), .Q(n14448) );
  AND2X1 U14703 ( .IN1(n10030), .IN2(CRC_OUT_6_31), .Q(n14447) );
  OR2X1 U14704 ( .IN1(n14449), .IN2(n14450), .Q(n14445) );
  AND2X1 U14705 ( .IN1(n9990), .IN2(n14451), .Q(n14450) );
  AND2X1 U14706 ( .IN1(n10065), .IN2(n13692), .Q(n14449) );
  OR2X1 U14707 ( .IN1(n14452), .IN2(n14453), .Q(n13692) );
  INVX0 U14708 ( .INP(n14454), .ZN(n14453) );
  OR2X1 U14709 ( .IN1(n14455), .IN2(n14456), .Q(n14454) );
  AND2X1 U14710 ( .IN1(n14456), .IN2(n14455), .Q(n14452) );
  INVX0 U14711 ( .INP(n14457), .ZN(n14455) );
  OR2X1 U14712 ( .IN1(n14458), .IN2(n14459), .Q(n14457) );
  AND2X1 U14713 ( .IN1(n10524), .IN2(n8495), .Q(n14459) );
  AND2X1 U14714 ( .IN1(n17941), .IN2(n10541), .Q(n14458) );
  OR2X1 U14715 ( .IN1(n14460), .IN2(n14461), .Q(n14456) );
  AND2X1 U14716 ( .IN1(n9646), .IN2(n14462), .Q(n14461) );
  AND2X1 U14717 ( .IN1(n14463), .IN2(n14464), .Q(n14462) );
  OR2X1 U14718 ( .IN1(n9036), .IN2(WX5945), .Q(n14464) );
  OR2X1 U14719 ( .IN1(n9037), .IN2(WX5881), .Q(n14463) );
  AND2X1 U14720 ( .IN1(n14465), .IN2(WX6009), .Q(n14460) );
  OR2X1 U14721 ( .IN1(n14466), .IN2(n14467), .Q(n14465) );
  AND2X1 U14722 ( .IN1(n9036), .IN2(WX5945), .Q(n14467) );
  AND2X1 U14723 ( .IN1(n9037), .IN2(WX5881), .Q(n14466) );
  AND2X1 U14724 ( .IN1(n9846), .IN2(n10583), .Q(WX4425) );
  AND2X1 U14725 ( .IN1(n14468), .IN2(n10584), .Q(WX3912) );
  AND2X1 U14726 ( .IN1(n14469), .IN2(n14470), .Q(n14468) );
  OR2X1 U14727 ( .IN1(DFF_574_n1), .IN2(WX3423), .Q(n14470) );
  OR2X1 U14728 ( .IN1(n9701), .IN2(CRC_OUT_7_30), .Q(n14469) );
  AND2X1 U14729 ( .IN1(n14471), .IN2(n10584), .Q(WX3910) );
  AND2X1 U14730 ( .IN1(n14472), .IN2(n14473), .Q(n14471) );
  OR2X1 U14731 ( .IN1(DFF_573_n1), .IN2(WX3425), .Q(n14473) );
  OR2X1 U14732 ( .IN1(n9702), .IN2(CRC_OUT_7_29), .Q(n14472) );
  AND2X1 U14733 ( .IN1(n14474), .IN2(n10584), .Q(WX3908) );
  AND2X1 U14734 ( .IN1(n14475), .IN2(n14476), .Q(n14474) );
  OR2X1 U14735 ( .IN1(DFF_572_n1), .IN2(WX3427), .Q(n14476) );
  OR2X1 U14736 ( .IN1(n9703), .IN2(CRC_OUT_7_28), .Q(n14475) );
  AND2X1 U14737 ( .IN1(n14477), .IN2(n10583), .Q(WX3906) );
  OR2X1 U14738 ( .IN1(n14478), .IN2(n14479), .Q(n14477) );
  AND2X1 U14739 ( .IN1(n9704), .IN2(n9945), .Q(n14479) );
  AND2X1 U14740 ( .IN1(test_so32), .IN2(WX3429), .Q(n14478) );
  AND2X1 U14741 ( .IN1(n14480), .IN2(n10584), .Q(WX3904) );
  AND2X1 U14742 ( .IN1(n14481), .IN2(n14482), .Q(n14480) );
  OR2X1 U14743 ( .IN1(DFF_570_n1), .IN2(WX3431), .Q(n14482) );
  OR2X1 U14744 ( .IN1(n9705), .IN2(CRC_OUT_7_26), .Q(n14481) );
  AND2X1 U14745 ( .IN1(n14483), .IN2(n10584), .Q(WX3902) );
  AND2X1 U14746 ( .IN1(n14484), .IN2(n14485), .Q(n14483) );
  OR2X1 U14747 ( .IN1(DFF_569_n1), .IN2(WX3433), .Q(n14485) );
  OR2X1 U14748 ( .IN1(n9706), .IN2(CRC_OUT_7_25), .Q(n14484) );
  AND2X1 U14749 ( .IN1(n14486), .IN2(n10585), .Q(WX3900) );
  AND2X1 U14750 ( .IN1(n14487), .IN2(n14488), .Q(n14486) );
  OR2X1 U14751 ( .IN1(DFF_568_n1), .IN2(WX3435), .Q(n14488) );
  OR2X1 U14752 ( .IN1(n9707), .IN2(CRC_OUT_7_24), .Q(n14487) );
  AND2X1 U14753 ( .IN1(n14489), .IN2(n10583), .Q(WX3898) );
  AND2X1 U14754 ( .IN1(n14490), .IN2(n14491), .Q(n14489) );
  OR2X1 U14755 ( .IN1(DFF_567_n1), .IN2(WX3437), .Q(n14491) );
  OR2X1 U14756 ( .IN1(n9708), .IN2(CRC_OUT_7_23), .Q(n14490) );
  AND2X1 U14757 ( .IN1(n14492), .IN2(n10585), .Q(WX3896) );
  OR2X1 U14758 ( .IN1(n14493), .IN2(n14494), .Q(n14492) );
  AND2X1 U14759 ( .IN1(DFF_566_n1), .IN2(n9911), .Q(n14494) );
  AND2X1 U14760 ( .IN1(test_so29), .IN2(CRC_OUT_7_22), .Q(n14493) );
  AND2X1 U14761 ( .IN1(n14495), .IN2(n10585), .Q(WX3894) );
  AND2X1 U14762 ( .IN1(n14496), .IN2(n14497), .Q(n14495) );
  OR2X1 U14763 ( .IN1(DFF_565_n1), .IN2(WX3441), .Q(n14497) );
  OR2X1 U14764 ( .IN1(n9709), .IN2(CRC_OUT_7_21), .Q(n14496) );
  AND2X1 U14765 ( .IN1(n14498), .IN2(n10585), .Q(WX3892) );
  AND2X1 U14766 ( .IN1(n14499), .IN2(n14500), .Q(n14498) );
  OR2X1 U14767 ( .IN1(DFF_564_n1), .IN2(WX3443), .Q(n14500) );
  OR2X1 U14768 ( .IN1(n9710), .IN2(CRC_OUT_7_20), .Q(n14499) );
  AND2X1 U14769 ( .IN1(n14501), .IN2(n10584), .Q(WX3890) );
  AND2X1 U14770 ( .IN1(n14502), .IN2(n14503), .Q(n14501) );
  OR2X1 U14771 ( .IN1(DFF_563_n1), .IN2(WX3445), .Q(n14503) );
  OR2X1 U14772 ( .IN1(n9711), .IN2(CRC_OUT_7_19), .Q(n14502) );
  AND2X1 U14773 ( .IN1(n14504), .IN2(n10585), .Q(WX3888) );
  AND2X1 U14774 ( .IN1(n14505), .IN2(n14506), .Q(n14504) );
  OR2X1 U14775 ( .IN1(DFF_562_n1), .IN2(WX3447), .Q(n14506) );
  OR2X1 U14776 ( .IN1(n9712), .IN2(CRC_OUT_7_18), .Q(n14505) );
  AND2X1 U14777 ( .IN1(n14507), .IN2(n10585), .Q(WX3886) );
  AND2X1 U14778 ( .IN1(n14508), .IN2(n14509), .Q(n14507) );
  OR2X1 U14779 ( .IN1(DFF_561_n1), .IN2(WX3449), .Q(n14509) );
  OR2X1 U14780 ( .IN1(n9713), .IN2(CRC_OUT_7_17), .Q(n14508) );
  AND2X1 U14781 ( .IN1(n14510), .IN2(n10584), .Q(WX3884) );
  AND2X1 U14782 ( .IN1(n14511), .IN2(n14512), .Q(n14510) );
  OR2X1 U14783 ( .IN1(DFF_560_n1), .IN2(WX3451), .Q(n14512) );
  OR2X1 U14784 ( .IN1(n9714), .IN2(CRC_OUT_7_16), .Q(n14511) );
  AND2X1 U14785 ( .IN1(n14513), .IN2(n10586), .Q(WX3882) );
  OR2X1 U14786 ( .IN1(n14514), .IN2(n14515), .Q(n14513) );
  AND2X1 U14787 ( .IN1(n14516), .IN2(CRC_OUT_7_15), .Q(n14515) );
  AND2X1 U14788 ( .IN1(DFF_559_n1), .IN2(n14517), .Q(n14514) );
  INVX0 U14789 ( .INP(n14516), .ZN(n14517) );
  OR2X1 U14790 ( .IN1(n14518), .IN2(n14519), .Q(n14516) );
  AND2X1 U14791 ( .IN1(DFF_575_n1), .IN2(WX3453), .Q(n14519) );
  AND2X1 U14792 ( .IN1(n9527), .IN2(CRC_OUT_7_31), .Q(n14518) );
  AND2X1 U14793 ( .IN1(n14520), .IN2(n10586), .Q(WX3880) );
  AND2X1 U14794 ( .IN1(n14521), .IN2(n14522), .Q(n14520) );
  OR2X1 U14795 ( .IN1(DFF_558_n1), .IN2(WX3455), .Q(n14522) );
  OR2X1 U14796 ( .IN1(n9715), .IN2(CRC_OUT_7_14), .Q(n14521) );
  AND2X1 U14797 ( .IN1(n14523), .IN2(n10588), .Q(WX3878) );
  AND2X1 U14798 ( .IN1(n14524), .IN2(n14525), .Q(n14523) );
  OR2X1 U14799 ( .IN1(DFF_557_n1), .IN2(WX3457), .Q(n14525) );
  OR2X1 U14800 ( .IN1(n9716), .IN2(CRC_OUT_7_13), .Q(n14524) );
  AND2X1 U14801 ( .IN1(n14526), .IN2(n10586), .Q(WX3876) );
  AND2X1 U14802 ( .IN1(n14527), .IN2(n14528), .Q(n14526) );
  OR2X1 U14803 ( .IN1(DFF_556_n1), .IN2(WX3459), .Q(n14528) );
  OR2X1 U14804 ( .IN1(n9717), .IN2(CRC_OUT_7_12), .Q(n14527) );
  AND2X1 U14805 ( .IN1(n14529), .IN2(n10586), .Q(WX3874) );
  AND2X1 U14806 ( .IN1(n14530), .IN2(n14531), .Q(n14529) );
  OR2X1 U14807 ( .IN1(DFF_555_n1), .IN2(WX3461), .Q(n14531) );
  OR2X1 U14808 ( .IN1(n9718), .IN2(CRC_OUT_7_11), .Q(n14530) );
  AND2X1 U14809 ( .IN1(n14532), .IN2(n10588), .Q(WX3872) );
  AND2X1 U14810 ( .IN1(n14533), .IN2(n14534), .Q(n14532) );
  OR2X1 U14811 ( .IN1(DFF_575_n1), .IN2(n14535), .Q(n14534) );
  AND2X1 U14812 ( .IN1(n14536), .IN2(n14537), .Q(n14535) );
  OR2X1 U14813 ( .IN1(n9528), .IN2(n9889), .Q(n14537) );
  OR2X1 U14814 ( .IN1(test_so31), .IN2(WX3463), .Q(n14536) );
  OR2X1 U14815 ( .IN1(n14538), .IN2(CRC_OUT_7_31), .Q(n14533) );
  OR2X1 U14816 ( .IN1(n14539), .IN2(n14540), .Q(n14538) );
  AND2X1 U14817 ( .IN1(n9528), .IN2(n9889), .Q(n14540) );
  AND2X1 U14818 ( .IN1(test_so31), .IN2(WX3463), .Q(n14539) );
  AND2X1 U14819 ( .IN1(n14541), .IN2(n10588), .Q(WX3870) );
  AND2X1 U14820 ( .IN1(n14542), .IN2(n14543), .Q(n14541) );
  OR2X1 U14821 ( .IN1(DFF_553_n1), .IN2(WX3465), .Q(n14543) );
  OR2X1 U14822 ( .IN1(n9719), .IN2(CRC_OUT_7_9), .Q(n14542) );
  AND2X1 U14823 ( .IN1(n14544), .IN2(n10586), .Q(WX3868) );
  AND2X1 U14824 ( .IN1(n14545), .IN2(n14546), .Q(n14544) );
  OR2X1 U14825 ( .IN1(DFF_552_n1), .IN2(WX3467), .Q(n14546) );
  OR2X1 U14826 ( .IN1(n9720), .IN2(CRC_OUT_7_8), .Q(n14545) );
  AND2X1 U14827 ( .IN1(n14547), .IN2(n10588), .Q(WX3866) );
  AND2X1 U14828 ( .IN1(n14548), .IN2(n14549), .Q(n14547) );
  OR2X1 U14829 ( .IN1(DFF_551_n1), .IN2(WX3469), .Q(n14549) );
  OR2X1 U14830 ( .IN1(n9721), .IN2(CRC_OUT_7_7), .Q(n14548) );
  AND2X1 U14831 ( .IN1(n14550), .IN2(n10588), .Q(WX3864) );
  AND2X1 U14832 ( .IN1(n14551), .IN2(n14552), .Q(n14550) );
  OR2X1 U14833 ( .IN1(DFF_550_n1), .IN2(WX3471), .Q(n14552) );
  OR2X1 U14834 ( .IN1(n9722), .IN2(CRC_OUT_7_6), .Q(n14551) );
  AND2X1 U14835 ( .IN1(n14553), .IN2(n10588), .Q(WX3862) );
  OR2X1 U14836 ( .IN1(n14554), .IN2(n14555), .Q(n14553) );
  AND2X1 U14837 ( .IN1(DFF_549_n1), .IN2(n9904), .Q(n14555) );
  AND2X1 U14838 ( .IN1(test_so30), .IN2(CRC_OUT_7_5), .Q(n14554) );
  AND2X1 U14839 ( .IN1(n14556), .IN2(n10585), .Q(WX3860) );
  AND2X1 U14840 ( .IN1(n14557), .IN2(n14558), .Q(n14556) );
  OR2X1 U14841 ( .IN1(DFF_548_n1), .IN2(WX3475), .Q(n14558) );
  OR2X1 U14842 ( .IN1(n9723), .IN2(CRC_OUT_7_4), .Q(n14557) );
  AND2X1 U14843 ( .IN1(n14559), .IN2(n10588), .Q(WX3858) );
  OR2X1 U14844 ( .IN1(n14560), .IN2(n14561), .Q(n14559) );
  AND2X1 U14845 ( .IN1(n14562), .IN2(CRC_OUT_7_3), .Q(n14561) );
  AND2X1 U14846 ( .IN1(DFF_547_n1), .IN2(n14563), .Q(n14560) );
  INVX0 U14847 ( .INP(n14562), .ZN(n14563) );
  OR2X1 U14848 ( .IN1(n14564), .IN2(n14565), .Q(n14562) );
  AND2X1 U14849 ( .IN1(DFF_575_n1), .IN2(WX3477), .Q(n14565) );
  AND2X1 U14850 ( .IN1(n9529), .IN2(CRC_OUT_7_31), .Q(n14564) );
  AND2X1 U14851 ( .IN1(n14566), .IN2(n10587), .Q(WX3856) );
  AND2X1 U14852 ( .IN1(n14567), .IN2(n14568), .Q(n14566) );
  OR2X1 U14853 ( .IN1(DFF_546_n1), .IN2(WX3479), .Q(n14568) );
  OR2X1 U14854 ( .IN1(n9724), .IN2(CRC_OUT_7_2), .Q(n14567) );
  AND2X1 U14855 ( .IN1(n14569), .IN2(n10589), .Q(WX3854) );
  AND2X1 U14856 ( .IN1(n14570), .IN2(n14571), .Q(n14569) );
  OR2X1 U14857 ( .IN1(DFF_545_n1), .IN2(WX3481), .Q(n14571) );
  OR2X1 U14858 ( .IN1(n9725), .IN2(CRC_OUT_7_1), .Q(n14570) );
  AND2X1 U14859 ( .IN1(n14572), .IN2(n10586), .Q(WX3852) );
  AND2X1 U14860 ( .IN1(n14573), .IN2(n14574), .Q(n14572) );
  OR2X1 U14861 ( .IN1(DFF_544_n1), .IN2(WX3483), .Q(n14574) );
  OR2X1 U14862 ( .IN1(n9726), .IN2(CRC_OUT_7_0), .Q(n14573) );
  AND2X1 U14863 ( .IN1(n14575), .IN2(n10589), .Q(WX3850) );
  AND2X1 U14864 ( .IN1(n14576), .IN2(n14577), .Q(n14575) );
  OR2X1 U14865 ( .IN1(DFF_575_n1), .IN2(WX3485), .Q(n14577) );
  OR2X1 U14866 ( .IN1(n9539), .IN2(CRC_OUT_7_31), .Q(n14576) );
  AND2X1 U14867 ( .IN1(test_so24), .IN2(n10589), .Q(WX3324) );
  AND2X1 U14868 ( .IN1(n10596), .IN2(n8597), .Q(WX3322) );
  AND2X1 U14869 ( .IN1(n10596), .IN2(n8598), .Q(WX3320) );
  AND2X1 U14870 ( .IN1(n10596), .IN2(n8599), .Q(WX3318) );
  AND2X1 U14871 ( .IN1(n10596), .IN2(n8600), .Q(WX3316) );
  AND2X1 U14872 ( .IN1(n10596), .IN2(n8601), .Q(WX3314) );
  AND2X1 U14873 ( .IN1(n10596), .IN2(n8602), .Q(WX3312) );
  AND2X1 U14874 ( .IN1(n10596), .IN2(n8603), .Q(WX3310) );
  AND2X1 U14875 ( .IN1(n10597), .IN2(n8604), .Q(WX3308) );
  AND2X1 U14876 ( .IN1(n10597), .IN2(n8605), .Q(WX3306) );
  AND2X1 U14877 ( .IN1(n10597), .IN2(n8606), .Q(WX3304) );
  AND2X1 U14878 ( .IN1(n10597), .IN2(n8607), .Q(WX3302) );
  AND2X1 U14879 ( .IN1(n10597), .IN2(n8608), .Q(WX3300) );
  AND2X1 U14880 ( .IN1(n10597), .IN2(n8609), .Q(WX3298) );
  AND2X1 U14881 ( .IN1(n10597), .IN2(n8610), .Q(WX3296) );
  AND2X1 U14882 ( .IN1(n10597), .IN2(n8611), .Q(WX3294) );
  OR2X1 U14883 ( .IN1(n14578), .IN2(n14579), .Q(WX3292) );
  OR2X1 U14884 ( .IN1(n14580), .IN2(n14581), .Q(n14579) );
  AND2X1 U14885 ( .IN1(n10030), .IN2(CRC_OUT_7_0), .Q(n14581) );
  AND2X1 U14886 ( .IN1(n521), .IN2(n10003), .Q(n14580) );
  INVX0 U14887 ( .INP(n14582), .ZN(n521) );
  OR2X1 U14888 ( .IN1(n10636), .IN2(n3972), .Q(n14582) );
  OR2X1 U14889 ( .IN1(n14583), .IN2(n14584), .Q(n14578) );
  AND2X1 U14890 ( .IN1(n9990), .IN2(n14585), .Q(n14584) );
  AND2X1 U14891 ( .IN1(n13826), .IN2(n10057), .Q(n14583) );
  AND2X1 U14892 ( .IN1(n14586), .IN2(n14587), .Q(n13826) );
  INVX0 U14893 ( .INP(n14588), .ZN(n14587) );
  AND2X1 U14894 ( .IN1(n14589), .IN2(n14590), .Q(n14588) );
  OR2X1 U14895 ( .IN1(n14590), .IN2(n14589), .Q(n14586) );
  OR2X1 U14896 ( .IN1(n14591), .IN2(n14592), .Q(n14589) );
  AND2X1 U14897 ( .IN1(n3691), .IN2(WX4714), .Q(n14592) );
  INVX0 U14898 ( .INP(n14593), .ZN(n14591) );
  OR2X1 U14899 ( .IN1(WX4714), .IN2(n3691), .Q(n14593) );
  AND2X1 U14900 ( .IN1(n14594), .IN2(n14595), .Q(n14590) );
  OR2X1 U14901 ( .IN1(WX4778), .IN2(test_so36), .Q(n14595) );
  OR2X1 U14902 ( .IN1(n9926), .IN2(n9538), .Q(n14594) );
  OR2X1 U14903 ( .IN1(n14596), .IN2(n14597), .Q(WX3290) );
  OR2X1 U14904 ( .IN1(n14598), .IN2(n14599), .Q(n14597) );
  AND2X1 U14905 ( .IN1(n10030), .IN2(CRC_OUT_7_1), .Q(n14599) );
  AND2X1 U14906 ( .IN1(n520), .IN2(n10004), .Q(n14598) );
  INVX0 U14907 ( .INP(n14600), .ZN(n520) );
  OR2X1 U14908 ( .IN1(n10636), .IN2(n3973), .Q(n14600) );
  OR2X1 U14909 ( .IN1(n14601), .IN2(n14602), .Q(n14596) );
  AND2X1 U14910 ( .IN1(n9990), .IN2(n14603), .Q(n14602) );
  AND2X1 U14911 ( .IN1(n10065), .IN2(n13843), .Q(n14601) );
  OR2X1 U14912 ( .IN1(n14604), .IN2(n14605), .Q(n13843) );
  INVX0 U14913 ( .INP(n14606), .ZN(n14605) );
  OR2X1 U14914 ( .IN1(n14607), .IN2(n14608), .Q(n14606) );
  AND2X1 U14915 ( .IN1(n14608), .IN2(n14607), .Q(n14604) );
  AND2X1 U14916 ( .IN1(n14609), .IN2(n14610), .Q(n14607) );
  OR2X1 U14917 ( .IN1(WX4648), .IN2(n9422), .Q(n14610) );
  OR2X1 U14918 ( .IN1(WX4584), .IN2(n3693), .Q(n14609) );
  OR2X1 U14919 ( .IN1(n14611), .IN2(n14612), .Q(n14608) );
  AND2X1 U14920 ( .IN1(n9423), .IN2(WX4776), .Q(n14612) );
  AND2X1 U14921 ( .IN1(n9700), .IN2(WX4712), .Q(n14611) );
  OR2X1 U14922 ( .IN1(n14613), .IN2(n14614), .Q(WX3288) );
  OR2X1 U14923 ( .IN1(n14615), .IN2(n14616), .Q(n14614) );
  AND2X1 U14924 ( .IN1(n10030), .IN2(CRC_OUT_7_2), .Q(n14616) );
  AND2X1 U14925 ( .IN1(n519), .IN2(n10004), .Q(n14615) );
  INVX0 U14926 ( .INP(n14617), .ZN(n519) );
  OR2X1 U14927 ( .IN1(n10636), .IN2(n3974), .Q(n14617) );
  OR2X1 U14928 ( .IN1(n14618), .IN2(n14619), .Q(n14613) );
  AND2X1 U14929 ( .IN1(n9990), .IN2(n14620), .Q(n14619) );
  AND2X1 U14930 ( .IN1(n10065), .IN2(n13861), .Q(n14618) );
  OR2X1 U14931 ( .IN1(n14621), .IN2(n14622), .Q(n13861) );
  INVX0 U14932 ( .INP(n14623), .ZN(n14622) );
  OR2X1 U14933 ( .IN1(n14624), .IN2(n14625), .Q(n14623) );
  AND2X1 U14934 ( .IN1(n14625), .IN2(n14624), .Q(n14621) );
  AND2X1 U14935 ( .IN1(n14626), .IN2(n14627), .Q(n14624) );
  OR2X1 U14936 ( .IN1(WX4646), .IN2(n9424), .Q(n14627) );
  OR2X1 U14937 ( .IN1(WX4582), .IN2(n3695), .Q(n14626) );
  OR2X1 U14938 ( .IN1(n14628), .IN2(n14629), .Q(n14625) );
  AND2X1 U14939 ( .IN1(n9425), .IN2(WX4774), .Q(n14629) );
  AND2X1 U14940 ( .IN1(n9699), .IN2(WX4710), .Q(n14628) );
  OR2X1 U14941 ( .IN1(n14630), .IN2(n14631), .Q(WX3286) );
  OR2X1 U14942 ( .IN1(n14632), .IN2(n14633), .Q(n14631) );
  AND2X1 U14943 ( .IN1(n10031), .IN2(CRC_OUT_7_3), .Q(n14633) );
  AND2X1 U14944 ( .IN1(n518), .IN2(n10004), .Q(n14632) );
  INVX0 U14945 ( .INP(n14634), .ZN(n518) );
  OR2X1 U14946 ( .IN1(n10636), .IN2(n3975), .Q(n14634) );
  OR2X1 U14947 ( .IN1(n14635), .IN2(n14636), .Q(n14630) );
  AND2X1 U14948 ( .IN1(n9990), .IN2(n14637), .Q(n14636) );
  AND2X1 U14949 ( .IN1(n10065), .IN2(n13878), .Q(n14635) );
  OR2X1 U14950 ( .IN1(n14638), .IN2(n14639), .Q(n13878) );
  INVX0 U14951 ( .INP(n14640), .ZN(n14639) );
  OR2X1 U14952 ( .IN1(n14641), .IN2(n14642), .Q(n14640) );
  AND2X1 U14953 ( .IN1(n14642), .IN2(n14641), .Q(n14638) );
  AND2X1 U14954 ( .IN1(n14643), .IN2(n14644), .Q(n14641) );
  OR2X1 U14955 ( .IN1(WX4644), .IN2(n9426), .Q(n14644) );
  OR2X1 U14956 ( .IN1(WX4580), .IN2(n3697), .Q(n14643) );
  OR2X1 U14957 ( .IN1(n14645), .IN2(n14646), .Q(n14642) );
  AND2X1 U14958 ( .IN1(n9427), .IN2(WX4772), .Q(n14646) );
  AND2X1 U14959 ( .IN1(n9698), .IN2(WX4708), .Q(n14645) );
  OR2X1 U14960 ( .IN1(n14647), .IN2(n14648), .Q(WX3284) );
  OR2X1 U14961 ( .IN1(n14649), .IN2(n14650), .Q(n14648) );
  AND2X1 U14962 ( .IN1(n10030), .IN2(CRC_OUT_7_4), .Q(n14650) );
  AND2X1 U14963 ( .IN1(n517), .IN2(n10004), .Q(n14649) );
  INVX0 U14964 ( .INP(n14651), .ZN(n517) );
  OR2X1 U14965 ( .IN1(n10636), .IN2(n3976), .Q(n14651) );
  OR2X1 U14966 ( .IN1(n14652), .IN2(n14653), .Q(n14647) );
  AND2X1 U14967 ( .IN1(n9990), .IN2(n14654), .Q(n14653) );
  AND2X1 U14968 ( .IN1(n10065), .IN2(n13896), .Q(n14652) );
  OR2X1 U14969 ( .IN1(n14655), .IN2(n14656), .Q(n13896) );
  INVX0 U14970 ( .INP(n14657), .ZN(n14656) );
  OR2X1 U14971 ( .IN1(n14658), .IN2(n14659), .Q(n14657) );
  AND2X1 U14972 ( .IN1(n14659), .IN2(n14658), .Q(n14655) );
  AND2X1 U14973 ( .IN1(n14660), .IN2(n14661), .Q(n14658) );
  OR2X1 U14974 ( .IN1(WX4642), .IN2(n9428), .Q(n14661) );
  OR2X1 U14975 ( .IN1(WX4578), .IN2(n3699), .Q(n14660) );
  OR2X1 U14976 ( .IN1(n14662), .IN2(n14663), .Q(n14659) );
  AND2X1 U14977 ( .IN1(n9429), .IN2(WX4770), .Q(n14663) );
  AND2X1 U14978 ( .IN1(n9526), .IN2(WX4706), .Q(n14662) );
  OR2X1 U14979 ( .IN1(n14664), .IN2(n14665), .Q(WX3282) );
  OR2X1 U14980 ( .IN1(n14666), .IN2(n14667), .Q(n14665) );
  AND2X1 U14981 ( .IN1(n10031), .IN2(CRC_OUT_7_5), .Q(n14667) );
  AND2X1 U14982 ( .IN1(n516), .IN2(n10004), .Q(n14666) );
  INVX0 U14983 ( .INP(n14668), .ZN(n516) );
  OR2X1 U14984 ( .IN1(n10636), .IN2(n3977), .Q(n14668) );
  OR2X1 U14985 ( .IN1(n14669), .IN2(n14670), .Q(n14664) );
  AND2X1 U14986 ( .IN1(n9990), .IN2(n14671), .Q(n14670) );
  AND2X1 U14987 ( .IN1(n10065), .IN2(n13913), .Q(n14669) );
  OR2X1 U14988 ( .IN1(n14672), .IN2(n14673), .Q(n13913) );
  INVX0 U14989 ( .INP(n14674), .ZN(n14673) );
  OR2X1 U14990 ( .IN1(n14675), .IN2(n14676), .Q(n14674) );
  AND2X1 U14991 ( .IN1(n14676), .IN2(n14675), .Q(n14672) );
  AND2X1 U14992 ( .IN1(n14677), .IN2(n14678), .Q(n14675) );
  OR2X1 U14993 ( .IN1(WX4640), .IN2(n9430), .Q(n14678) );
  OR2X1 U14994 ( .IN1(WX4576), .IN2(n3701), .Q(n14677) );
  OR2X1 U14995 ( .IN1(n14679), .IN2(n14680), .Q(n14676) );
  AND2X1 U14996 ( .IN1(n9431), .IN2(WX4768), .Q(n14680) );
  AND2X1 U14997 ( .IN1(n9697), .IN2(WX4704), .Q(n14679) );
  OR2X1 U14998 ( .IN1(n14681), .IN2(n14682), .Q(WX3280) );
  OR2X1 U14999 ( .IN1(n14683), .IN2(n14684), .Q(n14682) );
  AND2X1 U15000 ( .IN1(n10030), .IN2(CRC_OUT_7_6), .Q(n14684) );
  AND2X1 U15001 ( .IN1(n515), .IN2(n10004), .Q(n14683) );
  INVX0 U15002 ( .INP(n14685), .ZN(n515) );
  OR2X1 U15003 ( .IN1(n10636), .IN2(n3978), .Q(n14685) );
  OR2X1 U15004 ( .IN1(n14686), .IN2(n14687), .Q(n14681) );
  AND2X1 U15005 ( .IN1(n14688), .IN2(n9974), .Q(n14687) );
  AND2X1 U15006 ( .IN1(n10065), .IN2(n13931), .Q(n14686) );
  OR2X1 U15007 ( .IN1(n14689), .IN2(n14690), .Q(n13931) );
  INVX0 U15008 ( .INP(n14691), .ZN(n14690) );
  OR2X1 U15009 ( .IN1(n14692), .IN2(n14693), .Q(n14691) );
  AND2X1 U15010 ( .IN1(n14693), .IN2(n14692), .Q(n14689) );
  AND2X1 U15011 ( .IN1(n14694), .IN2(n14695), .Q(n14692) );
  OR2X1 U15012 ( .IN1(WX4638), .IN2(n9432), .Q(n14695) );
  OR2X1 U15013 ( .IN1(WX4574), .IN2(n3703), .Q(n14694) );
  OR2X1 U15014 ( .IN1(n14696), .IN2(n14697), .Q(n14693) );
  AND2X1 U15015 ( .IN1(n9433), .IN2(WX4766), .Q(n14697) );
  AND2X1 U15016 ( .IN1(n9696), .IN2(WX4702), .Q(n14696) );
  OR2X1 U15017 ( .IN1(n14698), .IN2(n14699), .Q(WX3278) );
  OR2X1 U15018 ( .IN1(n14700), .IN2(n14701), .Q(n14699) );
  AND2X1 U15019 ( .IN1(n10030), .IN2(CRC_OUT_7_7), .Q(n14701) );
  AND2X1 U15020 ( .IN1(n514), .IN2(n10004), .Q(n14700) );
  INVX0 U15021 ( .INP(n14702), .ZN(n514) );
  OR2X1 U15022 ( .IN1(n10636), .IN2(n3979), .Q(n14702) );
  OR2X1 U15023 ( .IN1(n14703), .IN2(n14704), .Q(n14698) );
  AND2X1 U15024 ( .IN1(n9990), .IN2(n14705), .Q(n14704) );
  AND2X1 U15025 ( .IN1(n10065), .IN2(n13948), .Q(n14703) );
  OR2X1 U15026 ( .IN1(n14706), .IN2(n14707), .Q(n13948) );
  INVX0 U15027 ( .INP(n14708), .ZN(n14707) );
  OR2X1 U15028 ( .IN1(n14709), .IN2(n14710), .Q(n14708) );
  AND2X1 U15029 ( .IN1(n14710), .IN2(n14709), .Q(n14706) );
  AND2X1 U15030 ( .IN1(n14711), .IN2(n14712), .Q(n14709) );
  OR2X1 U15031 ( .IN1(WX4636), .IN2(n9434), .Q(n14712) );
  OR2X1 U15032 ( .IN1(WX4572), .IN2(n3705), .Q(n14711) );
  OR2X1 U15033 ( .IN1(n14713), .IN2(n14714), .Q(n14710) );
  AND2X1 U15034 ( .IN1(n9435), .IN2(WX4764), .Q(n14714) );
  AND2X1 U15035 ( .IN1(n9695), .IN2(WX4700), .Q(n14713) );
  OR2X1 U15036 ( .IN1(n14715), .IN2(n14716), .Q(WX3276) );
  OR2X1 U15037 ( .IN1(n14717), .IN2(n14718), .Q(n14716) );
  AND2X1 U15038 ( .IN1(n10031), .IN2(CRC_OUT_7_8), .Q(n14718) );
  AND2X1 U15039 ( .IN1(n513), .IN2(n10004), .Q(n14717) );
  INVX0 U15040 ( .INP(n14719), .ZN(n513) );
  OR2X1 U15041 ( .IN1(n10636), .IN2(n3980), .Q(n14719) );
  OR2X1 U15042 ( .IN1(n14720), .IN2(n14721), .Q(n14715) );
  AND2X1 U15043 ( .IN1(n14722), .IN2(n9975), .Q(n14721) );
  AND2X1 U15044 ( .IN1(n10065), .IN2(n13965), .Q(n14720) );
  OR2X1 U15045 ( .IN1(n14723), .IN2(n14724), .Q(n13965) );
  INVX0 U15046 ( .INP(n14725), .ZN(n14724) );
  OR2X1 U15047 ( .IN1(n14726), .IN2(n14727), .Q(n14725) );
  AND2X1 U15048 ( .IN1(n14727), .IN2(n14726), .Q(n14723) );
  AND2X1 U15049 ( .IN1(n14728), .IN2(n14729), .Q(n14726) );
  OR2X1 U15050 ( .IN1(WX4634), .IN2(n9436), .Q(n14729) );
  OR2X1 U15051 ( .IN1(WX4570), .IN2(n3707), .Q(n14728) );
  OR2X1 U15052 ( .IN1(n14730), .IN2(n14731), .Q(n14727) );
  AND2X1 U15053 ( .IN1(n9437), .IN2(WX4762), .Q(n14731) );
  AND2X1 U15054 ( .IN1(n9694), .IN2(WX4698), .Q(n14730) );
  OR2X1 U15055 ( .IN1(n14732), .IN2(n14733), .Q(WX3274) );
  OR2X1 U15056 ( .IN1(n14734), .IN2(n14735), .Q(n14733) );
  AND2X1 U15057 ( .IN1(n10031), .IN2(CRC_OUT_7_9), .Q(n14735) );
  AND2X1 U15058 ( .IN1(n512), .IN2(n10004), .Q(n14734) );
  INVX0 U15059 ( .INP(n14736), .ZN(n512) );
  OR2X1 U15060 ( .IN1(n10635), .IN2(n3981), .Q(n14736) );
  OR2X1 U15061 ( .IN1(n14737), .IN2(n14738), .Q(n14732) );
  AND2X1 U15062 ( .IN1(n9989), .IN2(n14739), .Q(n14738) );
  AND2X1 U15063 ( .IN1(n10066), .IN2(n13982), .Q(n14737) );
  OR2X1 U15064 ( .IN1(n14740), .IN2(n14741), .Q(n13982) );
  INVX0 U15065 ( .INP(n14742), .ZN(n14741) );
  OR2X1 U15066 ( .IN1(n14743), .IN2(n14744), .Q(n14742) );
  AND2X1 U15067 ( .IN1(n14744), .IN2(n14743), .Q(n14740) );
  AND2X1 U15068 ( .IN1(n14745), .IN2(n14746), .Q(n14743) );
  OR2X1 U15069 ( .IN1(WX4632), .IN2(n9438), .Q(n14746) );
  OR2X1 U15070 ( .IN1(WX4568), .IN2(n3709), .Q(n14745) );
  OR2X1 U15071 ( .IN1(n14747), .IN2(n14748), .Q(n14744) );
  AND2X1 U15072 ( .IN1(n9439), .IN2(WX4760), .Q(n14748) );
  AND2X1 U15073 ( .IN1(n9693), .IN2(WX4696), .Q(n14747) );
  OR2X1 U15074 ( .IN1(n14749), .IN2(n14750), .Q(WX3272) );
  OR2X1 U15075 ( .IN1(n14751), .IN2(n14752), .Q(n14750) );
  AND2X1 U15076 ( .IN1(test_so31), .IN2(n10027), .Q(n14752) );
  AND2X1 U15077 ( .IN1(n511), .IN2(n10004), .Q(n14751) );
  INVX0 U15078 ( .INP(n14753), .ZN(n511) );
  OR2X1 U15079 ( .IN1(n10635), .IN2(n3982), .Q(n14753) );
  OR2X1 U15080 ( .IN1(n14754), .IN2(n14755), .Q(n14749) );
  AND2X1 U15081 ( .IN1(n9989), .IN2(n14756), .Q(n14755) );
  AND2X1 U15082 ( .IN1(n10066), .IN2(n13999), .Q(n14754) );
  OR2X1 U15083 ( .IN1(n14757), .IN2(n14758), .Q(n13999) );
  INVX0 U15084 ( .INP(n14759), .ZN(n14758) );
  OR2X1 U15085 ( .IN1(n14760), .IN2(n14761), .Q(n14759) );
  AND2X1 U15086 ( .IN1(n14761), .IN2(n14760), .Q(n14757) );
  AND2X1 U15087 ( .IN1(n14762), .IN2(n14763), .Q(n14760) );
  OR2X1 U15088 ( .IN1(WX4630), .IN2(n9440), .Q(n14763) );
  OR2X1 U15089 ( .IN1(WX4566), .IN2(n3711), .Q(n14762) );
  OR2X1 U15090 ( .IN1(n14764), .IN2(n14765), .Q(n14761) );
  AND2X1 U15091 ( .IN1(n9441), .IN2(WX4758), .Q(n14765) );
  AND2X1 U15092 ( .IN1(n9692), .IN2(WX4694), .Q(n14764) );
  OR2X1 U15093 ( .IN1(n14766), .IN2(n14767), .Q(WX3270) );
  OR2X1 U15094 ( .IN1(n14768), .IN2(n14769), .Q(n14767) );
  AND2X1 U15095 ( .IN1(n10031), .IN2(CRC_OUT_7_11), .Q(n14769) );
  AND2X1 U15096 ( .IN1(n510), .IN2(n10004), .Q(n14768) );
  INVX0 U15097 ( .INP(n14770), .ZN(n510) );
  OR2X1 U15098 ( .IN1(n10635), .IN2(n3983), .Q(n14770) );
  OR2X1 U15099 ( .IN1(n14771), .IN2(n14772), .Q(n14766) );
  AND2X1 U15100 ( .IN1(n9989), .IN2(n14773), .Q(n14772) );
  AND2X1 U15101 ( .IN1(n14016), .IN2(n10057), .Q(n14771) );
  AND2X1 U15102 ( .IN1(n14774), .IN2(n14775), .Q(n14016) );
  INVX0 U15103 ( .INP(n14776), .ZN(n14775) );
  AND2X1 U15104 ( .IN1(n14777), .IN2(n14778), .Q(n14776) );
  OR2X1 U15105 ( .IN1(n14778), .IN2(n14777), .Q(n14774) );
  OR2X1 U15106 ( .IN1(n14779), .IN2(n14780), .Q(n14777) );
  AND2X1 U15107 ( .IN1(n3713), .IN2(WX4564), .Q(n14780) );
  INVX0 U15108 ( .INP(n14781), .ZN(n14779) );
  OR2X1 U15109 ( .IN1(WX4564), .IN2(n3713), .Q(n14781) );
  AND2X1 U15110 ( .IN1(n14782), .IN2(n14783), .Q(n14778) );
  OR2X1 U15111 ( .IN1(WX4692), .IN2(test_so41), .Q(n14783) );
  OR2X1 U15112 ( .IN1(n9887), .IN2(n9443), .Q(n14782) );
  OR2X1 U15113 ( .IN1(n14784), .IN2(n14785), .Q(WX3268) );
  OR2X1 U15114 ( .IN1(n14786), .IN2(n14787), .Q(n14785) );
  AND2X1 U15115 ( .IN1(n10031), .IN2(CRC_OUT_7_12), .Q(n14787) );
  AND2X1 U15116 ( .IN1(n509), .IN2(n10004), .Q(n14786) );
  INVX0 U15117 ( .INP(n14788), .ZN(n509) );
  OR2X1 U15118 ( .IN1(n10635), .IN2(n3984), .Q(n14788) );
  OR2X1 U15119 ( .IN1(n14789), .IN2(n14790), .Q(n14784) );
  AND2X1 U15120 ( .IN1(n14791), .IN2(n9975), .Q(n14790) );
  AND2X1 U15121 ( .IN1(n10066), .IN2(n14033), .Q(n14789) );
  OR2X1 U15122 ( .IN1(n14792), .IN2(n14793), .Q(n14033) );
  INVX0 U15123 ( .INP(n14794), .ZN(n14793) );
  OR2X1 U15124 ( .IN1(n14795), .IN2(n14796), .Q(n14794) );
  AND2X1 U15125 ( .IN1(n14796), .IN2(n14795), .Q(n14792) );
  AND2X1 U15126 ( .IN1(n14797), .IN2(n14798), .Q(n14795) );
  OR2X1 U15127 ( .IN1(WX4626), .IN2(n9444), .Q(n14798) );
  OR2X1 U15128 ( .IN1(WX4562), .IN2(n3715), .Q(n14797) );
  OR2X1 U15129 ( .IN1(n14799), .IN2(n14800), .Q(n14796) );
  AND2X1 U15130 ( .IN1(n9445), .IN2(WX4754), .Q(n14800) );
  AND2X1 U15131 ( .IN1(n9691), .IN2(WX4690), .Q(n14799) );
  OR2X1 U15132 ( .IN1(n14801), .IN2(n14802), .Q(WX3266) );
  OR2X1 U15133 ( .IN1(n14803), .IN2(n14804), .Q(n14802) );
  AND2X1 U15134 ( .IN1(n10031), .IN2(CRC_OUT_7_13), .Q(n14804) );
  AND2X1 U15135 ( .IN1(n508), .IN2(n10005), .Q(n14803) );
  INVX0 U15136 ( .INP(n14805), .ZN(n508) );
  OR2X1 U15137 ( .IN1(n10635), .IN2(n3985), .Q(n14805) );
  OR2X1 U15138 ( .IN1(n14806), .IN2(n14807), .Q(n14801) );
  AND2X1 U15139 ( .IN1(n9989), .IN2(n14808), .Q(n14807) );
  AND2X1 U15140 ( .IN1(n14050), .IN2(n10057), .Q(n14806) );
  AND2X1 U15141 ( .IN1(n14809), .IN2(n14810), .Q(n14050) );
  INVX0 U15142 ( .INP(n14811), .ZN(n14810) );
  AND2X1 U15143 ( .IN1(n14812), .IN2(n14813), .Q(n14811) );
  OR2X1 U15144 ( .IN1(n14813), .IN2(n14812), .Q(n14809) );
  OR2X1 U15145 ( .IN1(n14814), .IN2(n14815), .Q(n14812) );
  AND2X1 U15146 ( .IN1(n3717), .IN2(WX4560), .Q(n14815) );
  INVX0 U15147 ( .INP(n14816), .ZN(n14814) );
  OR2X1 U15148 ( .IN1(WX4560), .IN2(n3717), .Q(n14816) );
  AND2X1 U15149 ( .IN1(n14817), .IN2(n14818), .Q(n14813) );
  OR2X1 U15150 ( .IN1(WX4752), .IN2(test_so39), .Q(n14818) );
  OR2X1 U15151 ( .IN1(n9927), .IN2(n9690), .Q(n14817) );
  OR2X1 U15152 ( .IN1(n14819), .IN2(n14820), .Q(WX3264) );
  OR2X1 U15153 ( .IN1(n14821), .IN2(n14822), .Q(n14820) );
  AND2X1 U15154 ( .IN1(n10031), .IN2(CRC_OUT_7_14), .Q(n14822) );
  AND2X1 U15155 ( .IN1(n507), .IN2(n10005), .Q(n14821) );
  INVX0 U15156 ( .INP(n14823), .ZN(n507) );
  OR2X1 U15157 ( .IN1(n10635), .IN2(n3986), .Q(n14823) );
  OR2X1 U15158 ( .IN1(n14824), .IN2(n14825), .Q(n14819) );
  AND2X1 U15159 ( .IN1(n9989), .IN2(n14826), .Q(n14825) );
  AND2X1 U15160 ( .IN1(n10066), .IN2(n14067), .Q(n14824) );
  OR2X1 U15161 ( .IN1(n14827), .IN2(n14828), .Q(n14067) );
  INVX0 U15162 ( .INP(n14829), .ZN(n14828) );
  OR2X1 U15163 ( .IN1(n14830), .IN2(n14831), .Q(n14829) );
  AND2X1 U15164 ( .IN1(n14831), .IN2(n14830), .Q(n14827) );
  AND2X1 U15165 ( .IN1(n14832), .IN2(n14833), .Q(n14830) );
  OR2X1 U15166 ( .IN1(WX4622), .IN2(n9447), .Q(n14833) );
  OR2X1 U15167 ( .IN1(WX4558), .IN2(n3719), .Q(n14832) );
  OR2X1 U15168 ( .IN1(n14834), .IN2(n14835), .Q(n14831) );
  AND2X1 U15169 ( .IN1(n9448), .IN2(WX4750), .Q(n14835) );
  AND2X1 U15170 ( .IN1(n9689), .IN2(WX4686), .Q(n14834) );
  OR2X1 U15171 ( .IN1(n14836), .IN2(n14837), .Q(WX3262) );
  OR2X1 U15172 ( .IN1(n14838), .IN2(n14839), .Q(n14837) );
  AND2X1 U15173 ( .IN1(n10031), .IN2(CRC_OUT_7_15), .Q(n14839) );
  AND2X1 U15174 ( .IN1(n506), .IN2(n10005), .Q(n14838) );
  INVX0 U15175 ( .INP(n14840), .ZN(n506) );
  OR2X1 U15176 ( .IN1(n10635), .IN2(n3987), .Q(n14840) );
  OR2X1 U15177 ( .IN1(n14841), .IN2(n14842), .Q(n14836) );
  AND2X1 U15178 ( .IN1(n9989), .IN2(n14843), .Q(n14842) );
  AND2X1 U15179 ( .IN1(n14084), .IN2(n10057), .Q(n14841) );
  AND2X1 U15180 ( .IN1(n14844), .IN2(n14845), .Q(n14084) );
  INVX0 U15181 ( .INP(n14846), .ZN(n14845) );
  AND2X1 U15182 ( .IN1(n14847), .IN2(n14848), .Q(n14846) );
  OR2X1 U15183 ( .IN1(n14848), .IN2(n14847), .Q(n14844) );
  OR2X1 U15184 ( .IN1(n14849), .IN2(n14850), .Q(n14847) );
  AND2X1 U15185 ( .IN1(n9449), .IN2(WX4684), .Q(n14850) );
  INVX0 U15186 ( .INP(n14851), .ZN(n14849) );
  OR2X1 U15187 ( .IN1(WX4684), .IN2(n9449), .Q(n14851) );
  AND2X1 U15188 ( .IN1(n14852), .IN2(n14853), .Q(n14848) );
  OR2X1 U15189 ( .IN1(WX4748), .IN2(test_so37), .Q(n14853) );
  OR2X1 U15190 ( .IN1(n9928), .IN2(n9688), .Q(n14852) );
  OR2X1 U15191 ( .IN1(n14854), .IN2(n14855), .Q(WX3260) );
  OR2X1 U15192 ( .IN1(n14856), .IN2(n14857), .Q(n14855) );
  AND2X1 U15193 ( .IN1(n10031), .IN2(CRC_OUT_7_16), .Q(n14857) );
  AND2X1 U15194 ( .IN1(n505), .IN2(n10005), .Q(n14856) );
  INVX0 U15195 ( .INP(n14858), .ZN(n505) );
  OR2X1 U15196 ( .IN1(n10635), .IN2(n3988), .Q(n14858) );
  OR2X1 U15197 ( .IN1(n14859), .IN2(n14860), .Q(n14854) );
  AND2X1 U15198 ( .IN1(n14861), .IN2(n9976), .Q(n14860) );
  AND2X1 U15199 ( .IN1(n10066), .IN2(n14101), .Q(n14859) );
  OR2X1 U15200 ( .IN1(n14862), .IN2(n14863), .Q(n14101) );
  INVX0 U15201 ( .INP(n14864), .ZN(n14863) );
  OR2X1 U15202 ( .IN1(n14865), .IN2(n14866), .Q(n14864) );
  AND2X1 U15203 ( .IN1(n14866), .IN2(n14865), .Q(n14862) );
  INVX0 U15204 ( .INP(n14867), .ZN(n14865) );
  OR2X1 U15205 ( .IN1(n14868), .IN2(n14869), .Q(n14867) );
  AND2X1 U15206 ( .IN1(n10524), .IN2(n8537), .Q(n14869) );
  AND2X1 U15207 ( .IN1(n17942), .IN2(n10541), .Q(n14868) );
  OR2X1 U15208 ( .IN1(n14870), .IN2(n14871), .Q(n14866) );
  AND2X1 U15209 ( .IN1(n9525), .IN2(n14872), .Q(n14871) );
  AND2X1 U15210 ( .IN1(n14873), .IN2(n14874), .Q(n14872) );
  OR2X1 U15211 ( .IN1(n9184), .IN2(WX4682), .Q(n14874) );
  OR2X1 U15212 ( .IN1(n9185), .IN2(WX4618), .Q(n14873) );
  AND2X1 U15213 ( .IN1(n14875), .IN2(WX4746), .Q(n14870) );
  OR2X1 U15214 ( .IN1(n14876), .IN2(n14877), .Q(n14875) );
  AND2X1 U15215 ( .IN1(n9184), .IN2(WX4682), .Q(n14877) );
  AND2X1 U15216 ( .IN1(n9185), .IN2(WX4618), .Q(n14876) );
  OR2X1 U15217 ( .IN1(n14878), .IN2(n14879), .Q(WX3258) );
  OR2X1 U15218 ( .IN1(n14880), .IN2(n14881), .Q(n14879) );
  AND2X1 U15219 ( .IN1(n10031), .IN2(CRC_OUT_7_17), .Q(n14881) );
  AND2X1 U15220 ( .IN1(n504), .IN2(n10005), .Q(n14880) );
  INVX0 U15221 ( .INP(n14882), .ZN(n504) );
  OR2X1 U15222 ( .IN1(n10635), .IN2(n3989), .Q(n14882) );
  OR2X1 U15223 ( .IN1(n14883), .IN2(n14884), .Q(n14878) );
  AND2X1 U15224 ( .IN1(n9989), .IN2(n14885), .Q(n14884) );
  AND2X1 U15225 ( .IN1(n14122), .IN2(n10057), .Q(n14883) );
  AND2X1 U15226 ( .IN1(n14886), .IN2(n14887), .Q(n14122) );
  OR2X1 U15227 ( .IN1(n14888), .IN2(n14889), .Q(n14887) );
  INVX0 U15228 ( .INP(n14890), .ZN(n14888) );
  OR2X1 U15229 ( .IN1(n14891), .IN2(n14890), .Q(n14886) );
  OR2X1 U15230 ( .IN1(n14892), .IN2(n14893), .Q(n14890) );
  AND2X1 U15231 ( .IN1(n10524), .IN2(WX4744), .Q(n14893) );
  AND2X1 U15232 ( .IN1(n9687), .IN2(n10541), .Q(n14892) );
  INVX0 U15233 ( .INP(n14889), .ZN(n14891) );
  OR2X1 U15234 ( .IN1(n14894), .IN2(n14895), .Q(n14889) );
  AND2X1 U15235 ( .IN1(n9187), .IN2(n14896), .Q(n14895) );
  AND2X1 U15236 ( .IN1(n14897), .IN2(n14898), .Q(n14896) );
  OR2X1 U15237 ( .IN1(n9186), .IN2(n9893), .Q(n14898) );
  OR2X1 U15238 ( .IN1(test_so35), .IN2(WX4616), .Q(n14897) );
  AND2X1 U15239 ( .IN1(n14899), .IN2(WX4680), .Q(n14894) );
  OR2X1 U15240 ( .IN1(n14900), .IN2(n14901), .Q(n14899) );
  AND2X1 U15241 ( .IN1(n9186), .IN2(n9893), .Q(n14901) );
  AND2X1 U15242 ( .IN1(test_so35), .IN2(WX4616), .Q(n14900) );
  OR2X1 U15243 ( .IN1(n14902), .IN2(n14903), .Q(WX3256) );
  OR2X1 U15244 ( .IN1(n14904), .IN2(n14905), .Q(n14903) );
  AND2X1 U15245 ( .IN1(n10032), .IN2(CRC_OUT_7_18), .Q(n14905) );
  AND2X1 U15246 ( .IN1(n503), .IN2(n10005), .Q(n14904) );
  INVX0 U15247 ( .INP(n14906), .ZN(n503) );
  OR2X1 U15248 ( .IN1(n10635), .IN2(n3990), .Q(n14906) );
  OR2X1 U15249 ( .IN1(n14907), .IN2(n14908), .Q(n14902) );
  AND2X1 U15250 ( .IN1(n9989), .IN2(n14909), .Q(n14908) );
  AND2X1 U15251 ( .IN1(n10066), .IN2(n14146), .Q(n14907) );
  OR2X1 U15252 ( .IN1(n14910), .IN2(n14911), .Q(n14146) );
  INVX0 U15253 ( .INP(n14912), .ZN(n14911) );
  OR2X1 U15254 ( .IN1(n14913), .IN2(n14914), .Q(n14912) );
  AND2X1 U15255 ( .IN1(n14914), .IN2(n14913), .Q(n14910) );
  INVX0 U15256 ( .INP(n14915), .ZN(n14913) );
  OR2X1 U15257 ( .IN1(n14916), .IN2(n14917), .Q(n14915) );
  AND2X1 U15258 ( .IN1(n10524), .IN2(n8540), .Q(n14917) );
  AND2X1 U15259 ( .IN1(n17943), .IN2(n10541), .Q(n14916) );
  OR2X1 U15260 ( .IN1(n14918), .IN2(n14919), .Q(n14914) );
  AND2X1 U15261 ( .IN1(n9686), .IN2(n14920), .Q(n14919) );
  AND2X1 U15262 ( .IN1(n14921), .IN2(n14922), .Q(n14920) );
  OR2X1 U15263 ( .IN1(n9188), .IN2(WX4678), .Q(n14922) );
  OR2X1 U15264 ( .IN1(n9189), .IN2(WX4614), .Q(n14921) );
  AND2X1 U15265 ( .IN1(n14923), .IN2(WX4742), .Q(n14918) );
  OR2X1 U15266 ( .IN1(n14924), .IN2(n14925), .Q(n14923) );
  AND2X1 U15267 ( .IN1(n9188), .IN2(WX4678), .Q(n14925) );
  AND2X1 U15268 ( .IN1(n9189), .IN2(WX4614), .Q(n14924) );
  OR2X1 U15269 ( .IN1(n14926), .IN2(n14927), .Q(WX3254) );
  OR2X1 U15270 ( .IN1(n14928), .IN2(n14929), .Q(n14927) );
  AND2X1 U15271 ( .IN1(n10031), .IN2(CRC_OUT_7_19), .Q(n14929) );
  AND2X1 U15272 ( .IN1(n502), .IN2(n10005), .Q(n14928) );
  INVX0 U15273 ( .INP(n14930), .ZN(n502) );
  OR2X1 U15274 ( .IN1(n10635), .IN2(n3991), .Q(n14930) );
  OR2X1 U15275 ( .IN1(n14931), .IN2(n14932), .Q(n14926) );
  AND2X1 U15276 ( .IN1(n9989), .IN2(n14933), .Q(n14932) );
  AND2X1 U15277 ( .IN1(n10066), .IN2(n14167), .Q(n14931) );
  OR2X1 U15278 ( .IN1(n14934), .IN2(n14935), .Q(n14167) );
  INVX0 U15279 ( .INP(n14936), .ZN(n14935) );
  OR2X1 U15280 ( .IN1(n14937), .IN2(n14938), .Q(n14936) );
  AND2X1 U15281 ( .IN1(n14938), .IN2(n14937), .Q(n14934) );
  INVX0 U15282 ( .INP(n14939), .ZN(n14937) );
  OR2X1 U15283 ( .IN1(n14940), .IN2(n14941), .Q(n14939) );
  AND2X1 U15284 ( .IN1(n10524), .IN2(n8541), .Q(n14941) );
  AND2X1 U15285 ( .IN1(n17944), .IN2(n10541), .Q(n14940) );
  OR2X1 U15286 ( .IN1(n14942), .IN2(n14943), .Q(n14938) );
  AND2X1 U15287 ( .IN1(n9685), .IN2(n14944), .Q(n14943) );
  AND2X1 U15288 ( .IN1(n14945), .IN2(n14946), .Q(n14944) );
  OR2X1 U15289 ( .IN1(n9190), .IN2(WX4676), .Q(n14946) );
  OR2X1 U15290 ( .IN1(n9191), .IN2(WX4612), .Q(n14945) );
  AND2X1 U15291 ( .IN1(n14947), .IN2(WX4740), .Q(n14942) );
  OR2X1 U15292 ( .IN1(n14948), .IN2(n14949), .Q(n14947) );
  AND2X1 U15293 ( .IN1(n9190), .IN2(WX4676), .Q(n14949) );
  AND2X1 U15294 ( .IN1(n9191), .IN2(WX4612), .Q(n14948) );
  OR2X1 U15295 ( .IN1(n14950), .IN2(n14951), .Q(WX3252) );
  OR2X1 U15296 ( .IN1(n14952), .IN2(n14953), .Q(n14951) );
  AND2X1 U15297 ( .IN1(n10032), .IN2(CRC_OUT_7_20), .Q(n14953) );
  AND2X1 U15298 ( .IN1(n501), .IN2(n10005), .Q(n14952) );
  INVX0 U15299 ( .INP(n14954), .ZN(n501) );
  OR2X1 U15300 ( .IN1(n10635), .IN2(n3992), .Q(n14954) );
  OR2X1 U15301 ( .IN1(n14955), .IN2(n14956), .Q(n14950) );
  AND2X1 U15302 ( .IN1(n9989), .IN2(n14957), .Q(n14956) );
  AND2X1 U15303 ( .IN1(n10066), .IN2(n14191), .Q(n14955) );
  OR2X1 U15304 ( .IN1(n14958), .IN2(n14959), .Q(n14191) );
  INVX0 U15305 ( .INP(n14960), .ZN(n14959) );
  OR2X1 U15306 ( .IN1(n14961), .IN2(n14962), .Q(n14960) );
  AND2X1 U15307 ( .IN1(n14962), .IN2(n14961), .Q(n14958) );
  INVX0 U15308 ( .INP(n14963), .ZN(n14961) );
  OR2X1 U15309 ( .IN1(n14964), .IN2(n14965), .Q(n14963) );
  AND2X1 U15310 ( .IN1(n10524), .IN2(n8542), .Q(n14965) );
  AND2X1 U15311 ( .IN1(n17945), .IN2(n10541), .Q(n14964) );
  OR2X1 U15312 ( .IN1(n14966), .IN2(n14967), .Q(n14962) );
  AND2X1 U15313 ( .IN1(n9684), .IN2(n14968), .Q(n14967) );
  AND2X1 U15314 ( .IN1(n14969), .IN2(n14970), .Q(n14968) );
  OR2X1 U15315 ( .IN1(n9192), .IN2(WX4674), .Q(n14970) );
  OR2X1 U15316 ( .IN1(n9193), .IN2(WX4610), .Q(n14969) );
  AND2X1 U15317 ( .IN1(n14971), .IN2(WX4738), .Q(n14966) );
  OR2X1 U15318 ( .IN1(n14972), .IN2(n14973), .Q(n14971) );
  AND2X1 U15319 ( .IN1(n9192), .IN2(WX4674), .Q(n14973) );
  AND2X1 U15320 ( .IN1(n9193), .IN2(WX4610), .Q(n14972) );
  OR2X1 U15321 ( .IN1(n14974), .IN2(n14975), .Q(WX3250) );
  OR2X1 U15322 ( .IN1(n14976), .IN2(n14977), .Q(n14975) );
  AND2X1 U15323 ( .IN1(n10032), .IN2(CRC_OUT_7_21), .Q(n14977) );
  AND2X1 U15324 ( .IN1(n500), .IN2(n10005), .Q(n14976) );
  INVX0 U15325 ( .INP(n14978), .ZN(n500) );
  OR2X1 U15326 ( .IN1(n10634), .IN2(n3993), .Q(n14978) );
  OR2X1 U15327 ( .IN1(n14979), .IN2(n14980), .Q(n14974) );
  AND2X1 U15328 ( .IN1(n9989), .IN2(n14981), .Q(n14980) );
  AND2X1 U15329 ( .IN1(n10066), .IN2(n14212), .Q(n14979) );
  OR2X1 U15330 ( .IN1(n14982), .IN2(n14983), .Q(n14212) );
  INVX0 U15331 ( .INP(n14984), .ZN(n14983) );
  OR2X1 U15332 ( .IN1(n14985), .IN2(n14986), .Q(n14984) );
  AND2X1 U15333 ( .IN1(n14986), .IN2(n14985), .Q(n14982) );
  INVX0 U15334 ( .INP(n14987), .ZN(n14985) );
  OR2X1 U15335 ( .IN1(n14988), .IN2(n14989), .Q(n14987) );
  AND2X1 U15336 ( .IN1(n10524), .IN2(n8543), .Q(n14989) );
  AND2X1 U15337 ( .IN1(n17946), .IN2(n10541), .Q(n14988) );
  OR2X1 U15338 ( .IN1(n14990), .IN2(n14991), .Q(n14986) );
  AND2X1 U15339 ( .IN1(n9683), .IN2(n14992), .Q(n14991) );
  AND2X1 U15340 ( .IN1(n14993), .IN2(n14994), .Q(n14992) );
  OR2X1 U15341 ( .IN1(n9194), .IN2(WX4672), .Q(n14994) );
  OR2X1 U15342 ( .IN1(n9195), .IN2(WX4608), .Q(n14993) );
  AND2X1 U15343 ( .IN1(n14995), .IN2(WX4736), .Q(n14990) );
  OR2X1 U15344 ( .IN1(n14996), .IN2(n14997), .Q(n14995) );
  AND2X1 U15345 ( .IN1(n9194), .IN2(WX4672), .Q(n14997) );
  AND2X1 U15346 ( .IN1(n9195), .IN2(WX4608), .Q(n14996) );
  OR2X1 U15347 ( .IN1(n14998), .IN2(n14999), .Q(WX3248) );
  OR2X1 U15348 ( .IN1(n15000), .IN2(n15001), .Q(n14999) );
  AND2X1 U15349 ( .IN1(n10032), .IN2(CRC_OUT_7_22), .Q(n15001) );
  AND2X1 U15350 ( .IN1(n499), .IN2(n10005), .Q(n15000) );
  INVX0 U15351 ( .INP(n15002), .ZN(n499) );
  OR2X1 U15352 ( .IN1(n10634), .IN2(n3994), .Q(n15002) );
  OR2X1 U15353 ( .IN1(n15003), .IN2(n15004), .Q(n14998) );
  AND2X1 U15354 ( .IN1(n9989), .IN2(n15005), .Q(n15004) );
  AND2X1 U15355 ( .IN1(n10066), .IN2(n14236), .Q(n15003) );
  OR2X1 U15356 ( .IN1(n15006), .IN2(n15007), .Q(n14236) );
  INVX0 U15357 ( .INP(n15008), .ZN(n15007) );
  OR2X1 U15358 ( .IN1(n15009), .IN2(n15010), .Q(n15008) );
  AND2X1 U15359 ( .IN1(n15010), .IN2(n15009), .Q(n15006) );
  INVX0 U15360 ( .INP(n15011), .ZN(n15009) );
  OR2X1 U15361 ( .IN1(n15012), .IN2(n15013), .Q(n15011) );
  AND2X1 U15362 ( .IN1(n10524), .IN2(n8544), .Q(n15013) );
  AND2X1 U15363 ( .IN1(n17947), .IN2(n10541), .Q(n15012) );
  OR2X1 U15364 ( .IN1(n15014), .IN2(n15015), .Q(n15010) );
  AND2X1 U15365 ( .IN1(n9682), .IN2(n15016), .Q(n15015) );
  AND2X1 U15366 ( .IN1(n15017), .IN2(n15018), .Q(n15016) );
  OR2X1 U15367 ( .IN1(n9196), .IN2(WX4670), .Q(n15018) );
  OR2X1 U15368 ( .IN1(n9197), .IN2(WX4606), .Q(n15017) );
  AND2X1 U15369 ( .IN1(n15019), .IN2(WX4734), .Q(n15014) );
  OR2X1 U15370 ( .IN1(n15020), .IN2(n15021), .Q(n15019) );
  AND2X1 U15371 ( .IN1(n9196), .IN2(WX4670), .Q(n15021) );
  AND2X1 U15372 ( .IN1(n9197), .IN2(WX4606), .Q(n15020) );
  OR2X1 U15373 ( .IN1(n15022), .IN2(n15023), .Q(WX3246) );
  OR2X1 U15374 ( .IN1(n15024), .IN2(n15025), .Q(n15023) );
  AND2X1 U15375 ( .IN1(n10037), .IN2(CRC_OUT_7_23), .Q(n15025) );
  AND2X1 U15376 ( .IN1(n498), .IN2(n10005), .Q(n15024) );
  INVX0 U15377 ( .INP(n15026), .ZN(n498) );
  OR2X1 U15378 ( .IN1(n10634), .IN2(n3995), .Q(n15026) );
  OR2X1 U15379 ( .IN1(n15027), .IN2(n15028), .Q(n15022) );
  AND2X1 U15380 ( .IN1(n15029), .IN2(n9977), .Q(n15028) );
  AND2X1 U15381 ( .IN1(n10069), .IN2(n14260), .Q(n15027) );
  OR2X1 U15382 ( .IN1(n15030), .IN2(n15031), .Q(n14260) );
  INVX0 U15383 ( .INP(n15032), .ZN(n15031) );
  OR2X1 U15384 ( .IN1(n15033), .IN2(n15034), .Q(n15032) );
  AND2X1 U15385 ( .IN1(n15034), .IN2(n15033), .Q(n15030) );
  INVX0 U15386 ( .INP(n15035), .ZN(n15033) );
  OR2X1 U15387 ( .IN1(n15036), .IN2(n15037), .Q(n15035) );
  AND2X1 U15388 ( .IN1(n10524), .IN2(n8545), .Q(n15037) );
  AND2X1 U15389 ( .IN1(n17948), .IN2(n10541), .Q(n15036) );
  OR2X1 U15390 ( .IN1(n15038), .IN2(n15039), .Q(n15034) );
  AND2X1 U15391 ( .IN1(n9681), .IN2(n15040), .Q(n15039) );
  AND2X1 U15392 ( .IN1(n15041), .IN2(n15042), .Q(n15040) );
  OR2X1 U15393 ( .IN1(n9198), .IN2(WX4668), .Q(n15042) );
  OR2X1 U15394 ( .IN1(n9199), .IN2(WX4604), .Q(n15041) );
  AND2X1 U15395 ( .IN1(n15043), .IN2(WX4732), .Q(n15038) );
  OR2X1 U15396 ( .IN1(n15044), .IN2(n15045), .Q(n15043) );
  AND2X1 U15397 ( .IN1(n9198), .IN2(WX4668), .Q(n15045) );
  AND2X1 U15398 ( .IN1(n9199), .IN2(WX4604), .Q(n15044) );
  OR2X1 U15399 ( .IN1(n15046), .IN2(n15047), .Q(WX3244) );
  OR2X1 U15400 ( .IN1(n15048), .IN2(n15049), .Q(n15047) );
  AND2X1 U15401 ( .IN1(n10032), .IN2(CRC_OUT_7_24), .Q(n15049) );
  AND2X1 U15402 ( .IN1(n497), .IN2(n10006), .Q(n15048) );
  INVX0 U15403 ( .INP(n15050), .ZN(n497) );
  OR2X1 U15404 ( .IN1(n10634), .IN2(n3996), .Q(n15050) );
  OR2X1 U15405 ( .IN1(n15051), .IN2(n15052), .Q(n15046) );
  AND2X1 U15406 ( .IN1(n9988), .IN2(n15053), .Q(n15052) );
  AND2X1 U15407 ( .IN1(n10066), .IN2(n14284), .Q(n15051) );
  OR2X1 U15408 ( .IN1(n15054), .IN2(n15055), .Q(n14284) );
  INVX0 U15409 ( .INP(n15056), .ZN(n15055) );
  OR2X1 U15410 ( .IN1(n15057), .IN2(n15058), .Q(n15056) );
  AND2X1 U15411 ( .IN1(n15058), .IN2(n15057), .Q(n15054) );
  INVX0 U15412 ( .INP(n15059), .ZN(n15057) );
  OR2X1 U15413 ( .IN1(n15060), .IN2(n15061), .Q(n15059) );
  AND2X1 U15414 ( .IN1(n10524), .IN2(n8546), .Q(n15061) );
  AND2X1 U15415 ( .IN1(n17949), .IN2(n10541), .Q(n15060) );
  OR2X1 U15416 ( .IN1(n15062), .IN2(n15063), .Q(n15058) );
  AND2X1 U15417 ( .IN1(n9680), .IN2(n15064), .Q(n15063) );
  AND2X1 U15418 ( .IN1(n15065), .IN2(n15066), .Q(n15064) );
  OR2X1 U15419 ( .IN1(n9200), .IN2(WX4666), .Q(n15066) );
  OR2X1 U15420 ( .IN1(n9201), .IN2(WX4602), .Q(n15065) );
  AND2X1 U15421 ( .IN1(n15067), .IN2(WX4730), .Q(n15062) );
  OR2X1 U15422 ( .IN1(n15068), .IN2(n15069), .Q(n15067) );
  AND2X1 U15423 ( .IN1(n9200), .IN2(WX4666), .Q(n15069) );
  AND2X1 U15424 ( .IN1(n9201), .IN2(WX4602), .Q(n15068) );
  OR2X1 U15425 ( .IN1(n15070), .IN2(n15071), .Q(WX3242) );
  OR2X1 U15426 ( .IN1(n15072), .IN2(n15073), .Q(n15071) );
  AND2X1 U15427 ( .IN1(n10032), .IN2(CRC_OUT_7_25), .Q(n15073) );
  AND2X1 U15428 ( .IN1(n496), .IN2(n10006), .Q(n15072) );
  INVX0 U15429 ( .INP(n15074), .ZN(n496) );
  OR2X1 U15430 ( .IN1(n10634), .IN2(n3997), .Q(n15074) );
  OR2X1 U15431 ( .IN1(n15075), .IN2(n15076), .Q(n15070) );
  AND2X1 U15432 ( .IN1(n9988), .IN2(n15077), .Q(n15076) );
  AND2X1 U15433 ( .IN1(n10066), .IN2(n14308), .Q(n15075) );
  OR2X1 U15434 ( .IN1(n15078), .IN2(n15079), .Q(n14308) );
  INVX0 U15435 ( .INP(n15080), .ZN(n15079) );
  OR2X1 U15436 ( .IN1(n15081), .IN2(n15082), .Q(n15080) );
  AND2X1 U15437 ( .IN1(n15082), .IN2(n15081), .Q(n15078) );
  INVX0 U15438 ( .INP(n15083), .ZN(n15081) );
  OR2X1 U15439 ( .IN1(n15084), .IN2(n15085), .Q(n15083) );
  AND2X1 U15440 ( .IN1(n10525), .IN2(n8547), .Q(n15085) );
  AND2X1 U15441 ( .IN1(n17950), .IN2(n10541), .Q(n15084) );
  OR2X1 U15442 ( .IN1(n15086), .IN2(n15087), .Q(n15082) );
  AND2X1 U15443 ( .IN1(n9679), .IN2(n15088), .Q(n15087) );
  AND2X1 U15444 ( .IN1(n15089), .IN2(n15090), .Q(n15088) );
  OR2X1 U15445 ( .IN1(n9202), .IN2(WX4664), .Q(n15090) );
  OR2X1 U15446 ( .IN1(n9203), .IN2(WX4600), .Q(n15089) );
  AND2X1 U15447 ( .IN1(n15091), .IN2(WX4728), .Q(n15086) );
  OR2X1 U15448 ( .IN1(n15092), .IN2(n15093), .Q(n15091) );
  AND2X1 U15449 ( .IN1(n9202), .IN2(WX4664), .Q(n15093) );
  AND2X1 U15450 ( .IN1(n9203), .IN2(WX4600), .Q(n15092) );
  OR2X1 U15451 ( .IN1(n15094), .IN2(n15095), .Q(WX3240) );
  OR2X1 U15452 ( .IN1(n15096), .IN2(n15097), .Q(n15095) );
  AND2X1 U15453 ( .IN1(n10032), .IN2(CRC_OUT_7_26), .Q(n15097) );
  AND2X1 U15454 ( .IN1(n495), .IN2(n10006), .Q(n15096) );
  INVX0 U15455 ( .INP(n15098), .ZN(n495) );
  OR2X1 U15456 ( .IN1(n10634), .IN2(n3998), .Q(n15098) );
  OR2X1 U15457 ( .IN1(n15099), .IN2(n15100), .Q(n15094) );
  AND2X1 U15458 ( .IN1(n15101), .IN2(n9976), .Q(n15100) );
  AND2X1 U15459 ( .IN1(n10066), .IN2(n14332), .Q(n15099) );
  OR2X1 U15460 ( .IN1(n15102), .IN2(n15103), .Q(n14332) );
  INVX0 U15461 ( .INP(n15104), .ZN(n15103) );
  OR2X1 U15462 ( .IN1(n15105), .IN2(n15106), .Q(n15104) );
  AND2X1 U15463 ( .IN1(n15106), .IN2(n15105), .Q(n15102) );
  INVX0 U15464 ( .INP(n15107), .ZN(n15105) );
  OR2X1 U15465 ( .IN1(n15108), .IN2(n15109), .Q(n15107) );
  AND2X1 U15466 ( .IN1(n10525), .IN2(n8548), .Q(n15109) );
  AND2X1 U15467 ( .IN1(n17951), .IN2(n10541), .Q(n15108) );
  OR2X1 U15468 ( .IN1(n15110), .IN2(n15111), .Q(n15106) );
  AND2X1 U15469 ( .IN1(n9678), .IN2(n15112), .Q(n15111) );
  AND2X1 U15470 ( .IN1(n15113), .IN2(n15114), .Q(n15112) );
  OR2X1 U15471 ( .IN1(n9204), .IN2(WX4662), .Q(n15114) );
  OR2X1 U15472 ( .IN1(n9205), .IN2(WX4598), .Q(n15113) );
  AND2X1 U15473 ( .IN1(n15115), .IN2(WX4726), .Q(n15110) );
  OR2X1 U15474 ( .IN1(n15116), .IN2(n15117), .Q(n15115) );
  AND2X1 U15475 ( .IN1(n9204), .IN2(WX4662), .Q(n15117) );
  AND2X1 U15476 ( .IN1(n9205), .IN2(WX4598), .Q(n15116) );
  OR2X1 U15477 ( .IN1(n15118), .IN2(n15119), .Q(WX3238) );
  OR2X1 U15478 ( .IN1(n15120), .IN2(n15121), .Q(n15119) );
  AND2X1 U15479 ( .IN1(test_so32), .IN2(n10026), .Q(n15121) );
  AND2X1 U15480 ( .IN1(n494), .IN2(n10006), .Q(n15120) );
  INVX0 U15481 ( .INP(n15122), .ZN(n494) );
  OR2X1 U15482 ( .IN1(n10634), .IN2(n3999), .Q(n15122) );
  OR2X1 U15483 ( .IN1(n15123), .IN2(n15124), .Q(n15118) );
  AND2X1 U15484 ( .IN1(n9988), .IN2(n15125), .Q(n15124) );
  AND2X1 U15485 ( .IN1(n10067), .IN2(n14356), .Q(n15123) );
  OR2X1 U15486 ( .IN1(n15126), .IN2(n15127), .Q(n14356) );
  INVX0 U15487 ( .INP(n15128), .ZN(n15127) );
  OR2X1 U15488 ( .IN1(n15129), .IN2(n15130), .Q(n15128) );
  AND2X1 U15489 ( .IN1(n15130), .IN2(n15129), .Q(n15126) );
  INVX0 U15490 ( .INP(n15131), .ZN(n15129) );
  OR2X1 U15491 ( .IN1(n15132), .IN2(n15133), .Q(n15131) );
  AND2X1 U15492 ( .IN1(n10525), .IN2(n8549), .Q(n15133) );
  AND2X1 U15493 ( .IN1(n17952), .IN2(n10541), .Q(n15132) );
  OR2X1 U15494 ( .IN1(n15134), .IN2(n15135), .Q(n15130) );
  AND2X1 U15495 ( .IN1(n9677), .IN2(n15136), .Q(n15135) );
  AND2X1 U15496 ( .IN1(n15137), .IN2(n15138), .Q(n15136) );
  OR2X1 U15497 ( .IN1(n9206), .IN2(WX4660), .Q(n15138) );
  OR2X1 U15498 ( .IN1(n9207), .IN2(WX4596), .Q(n15137) );
  AND2X1 U15499 ( .IN1(n15139), .IN2(WX4724), .Q(n15134) );
  OR2X1 U15500 ( .IN1(n15140), .IN2(n15141), .Q(n15139) );
  AND2X1 U15501 ( .IN1(n9206), .IN2(WX4660), .Q(n15141) );
  AND2X1 U15502 ( .IN1(n9207), .IN2(WX4596), .Q(n15140) );
  OR2X1 U15503 ( .IN1(n15142), .IN2(n15143), .Q(WX3236) );
  OR2X1 U15504 ( .IN1(n15144), .IN2(n15145), .Q(n15143) );
  AND2X1 U15505 ( .IN1(n10032), .IN2(CRC_OUT_7_28), .Q(n15145) );
  AND2X1 U15506 ( .IN1(n493), .IN2(n10006), .Q(n15144) );
  INVX0 U15507 ( .INP(n15146), .ZN(n493) );
  OR2X1 U15508 ( .IN1(n10634), .IN2(n4000), .Q(n15146) );
  OR2X1 U15509 ( .IN1(n15147), .IN2(n15148), .Q(n15142) );
  AND2X1 U15510 ( .IN1(n9988), .IN2(n15149), .Q(n15148) );
  AND2X1 U15511 ( .IN1(n14380), .IN2(n10058), .Q(n15147) );
  AND2X1 U15512 ( .IN1(n15150), .IN2(n15151), .Q(n14380) );
  INVX0 U15513 ( .INP(n15152), .ZN(n15151) );
  AND2X1 U15514 ( .IN1(n15153), .IN2(n15154), .Q(n15152) );
  OR2X1 U15515 ( .IN1(n15154), .IN2(n15153), .Q(n15150) );
  OR2X1 U15516 ( .IN1(n15155), .IN2(n15156), .Q(n15153) );
  AND2X1 U15517 ( .IN1(n10525), .IN2(WX4594), .Q(n15156) );
  AND2X1 U15518 ( .IN1(n9208), .IN2(n10541), .Q(n15155) );
  AND2X1 U15519 ( .IN1(n15157), .IN2(n15158), .Q(n15154) );
  INVX0 U15520 ( .INP(n15159), .ZN(n15158) );
  AND2X1 U15521 ( .IN1(n15160), .IN2(WX4658), .Q(n15159) );
  OR2X1 U15522 ( .IN1(WX4658), .IN2(n15160), .Q(n15157) );
  OR2X1 U15523 ( .IN1(n15161), .IN2(n15162), .Q(n15160) );
  AND2X1 U15524 ( .IN1(n17953), .IN2(n9910), .Q(n15162) );
  AND2X1 U15525 ( .IN1(test_so40), .IN2(n8550), .Q(n15161) );
  OR2X1 U15526 ( .IN1(n15163), .IN2(n15164), .Q(WX3234) );
  OR2X1 U15527 ( .IN1(n15165), .IN2(n15166), .Q(n15164) );
  AND2X1 U15528 ( .IN1(n10032), .IN2(CRC_OUT_7_29), .Q(n15166) );
  AND2X1 U15529 ( .IN1(n492), .IN2(n10006), .Q(n15165) );
  INVX0 U15530 ( .INP(n15167), .ZN(n492) );
  OR2X1 U15531 ( .IN1(n10634), .IN2(n4001), .Q(n15167) );
  OR2X1 U15532 ( .IN1(n15168), .IN2(n15169), .Q(n15163) );
  AND2X1 U15533 ( .IN1(n9988), .IN2(n15170), .Q(n15169) );
  AND2X1 U15534 ( .IN1(n10067), .IN2(n14404), .Q(n15168) );
  OR2X1 U15535 ( .IN1(n15171), .IN2(n15172), .Q(n14404) );
  INVX0 U15536 ( .INP(n15173), .ZN(n15172) );
  OR2X1 U15537 ( .IN1(n15174), .IN2(n15175), .Q(n15173) );
  AND2X1 U15538 ( .IN1(n15175), .IN2(n15174), .Q(n15171) );
  INVX0 U15539 ( .INP(n15176), .ZN(n15174) );
  OR2X1 U15540 ( .IN1(n15177), .IN2(n15178), .Q(n15176) );
  AND2X1 U15541 ( .IN1(n10525), .IN2(n8551), .Q(n15178) );
  AND2X1 U15542 ( .IN1(n17954), .IN2(n10541), .Q(n15177) );
  OR2X1 U15543 ( .IN1(n15179), .IN2(n15180), .Q(n15175) );
  AND2X1 U15544 ( .IN1(n9676), .IN2(n15181), .Q(n15180) );
  AND2X1 U15545 ( .IN1(n15182), .IN2(n15183), .Q(n15181) );
  OR2X1 U15546 ( .IN1(n9210), .IN2(WX4656), .Q(n15183) );
  OR2X1 U15547 ( .IN1(n9211), .IN2(WX4592), .Q(n15182) );
  AND2X1 U15548 ( .IN1(n15184), .IN2(WX4720), .Q(n15179) );
  OR2X1 U15549 ( .IN1(n15185), .IN2(n15186), .Q(n15184) );
  AND2X1 U15550 ( .IN1(n9210), .IN2(WX4656), .Q(n15186) );
  AND2X1 U15551 ( .IN1(n9211), .IN2(WX4592), .Q(n15185) );
  OR2X1 U15552 ( .IN1(n15187), .IN2(n15188), .Q(WX3232) );
  OR2X1 U15553 ( .IN1(n15189), .IN2(n15190), .Q(n15188) );
  AND2X1 U15554 ( .IN1(n10032), .IN2(CRC_OUT_7_30), .Q(n15190) );
  AND2X1 U15555 ( .IN1(n491), .IN2(n10006), .Q(n15189) );
  INVX0 U15556 ( .INP(n15191), .ZN(n491) );
  OR2X1 U15557 ( .IN1(n10634), .IN2(n4002), .Q(n15191) );
  OR2X1 U15558 ( .IN1(n15192), .IN2(n15193), .Q(n15187) );
  AND2X1 U15559 ( .IN1(n15194), .IN2(n9976), .Q(n15193) );
  AND2X1 U15560 ( .IN1(n14428), .IN2(n10058), .Q(n15192) );
  AND2X1 U15561 ( .IN1(n15195), .IN2(n15196), .Q(n14428) );
  INVX0 U15562 ( .INP(n15197), .ZN(n15196) );
  AND2X1 U15563 ( .IN1(n15198), .IN2(n15199), .Q(n15197) );
  OR2X1 U15564 ( .IN1(n15199), .IN2(n15198), .Q(n15195) );
  OR2X1 U15565 ( .IN1(n15200), .IN2(n15201), .Q(n15198) );
  AND2X1 U15566 ( .IN1(n10525), .IN2(WX4590), .Q(n15201) );
  AND2X1 U15567 ( .IN1(n9212), .IN2(n10541), .Q(n15200) );
  AND2X1 U15568 ( .IN1(n15202), .IN2(n15203), .Q(n15199) );
  OR2X1 U15569 ( .IN1(n15204), .IN2(n9675), .Q(n15203) );
  INVX0 U15570 ( .INP(n15205), .ZN(n15204) );
  OR2X1 U15571 ( .IN1(WX4718), .IN2(n15205), .Q(n15202) );
  OR2X1 U15572 ( .IN1(n15206), .IN2(n15207), .Q(n15205) );
  AND2X1 U15573 ( .IN1(n17955), .IN2(n9961), .Q(n15207) );
  AND2X1 U15574 ( .IN1(test_so38), .IN2(n8552), .Q(n15206) );
  OR2X1 U15575 ( .IN1(n15208), .IN2(n15209), .Q(WX3230) );
  OR2X1 U15576 ( .IN1(n15210), .IN2(n15211), .Q(n15209) );
  AND2X1 U15577 ( .IN1(n2245), .IN2(WX3071), .Q(n15211) );
  AND2X1 U15578 ( .IN1(n10032), .IN2(CRC_OUT_7_31), .Q(n15210) );
  OR2X1 U15579 ( .IN1(n15212), .IN2(n15213), .Q(n15208) );
  AND2X1 U15580 ( .IN1(n9988), .IN2(n15214), .Q(n15213) );
  AND2X1 U15581 ( .IN1(n10067), .IN2(n14451), .Q(n15212) );
  OR2X1 U15582 ( .IN1(n15215), .IN2(n15216), .Q(n14451) );
  INVX0 U15583 ( .INP(n15217), .ZN(n15216) );
  OR2X1 U15584 ( .IN1(n15218), .IN2(n15219), .Q(n15217) );
  AND2X1 U15585 ( .IN1(n15219), .IN2(n15218), .Q(n15215) );
  INVX0 U15586 ( .INP(n15220), .ZN(n15218) );
  OR2X1 U15587 ( .IN1(n15221), .IN2(n15222), .Q(n15220) );
  AND2X1 U15588 ( .IN1(n10525), .IN2(n8553), .Q(n15222) );
  AND2X1 U15589 ( .IN1(n17956), .IN2(n10541), .Q(n15221) );
  OR2X1 U15590 ( .IN1(n15223), .IN2(n15224), .Q(n15219) );
  AND2X1 U15591 ( .IN1(n9674), .IN2(n15225), .Q(n15224) );
  AND2X1 U15592 ( .IN1(n15226), .IN2(n15227), .Q(n15225) );
  OR2X1 U15593 ( .IN1(n9038), .IN2(WX4652), .Q(n15227) );
  OR2X1 U15594 ( .IN1(n9039), .IN2(WX4588), .Q(n15226) );
  AND2X1 U15595 ( .IN1(n15228), .IN2(WX4716), .Q(n15223) );
  OR2X1 U15596 ( .IN1(n15229), .IN2(n15230), .Q(n15228) );
  AND2X1 U15597 ( .IN1(n9038), .IN2(WX4652), .Q(n15230) );
  AND2X1 U15598 ( .IN1(n9039), .IN2(WX4588), .Q(n15229) );
  AND2X1 U15599 ( .IN1(n9845), .IN2(n10586), .Q(WX3132) );
  AND2X1 U15600 ( .IN1(n15231), .IN2(n10588), .Q(WX2619) );
  AND2X1 U15601 ( .IN1(n15232), .IN2(n15233), .Q(n15231) );
  OR2X1 U15602 ( .IN1(DFF_382_n1), .IN2(WX2130), .Q(n15233) );
  OR2X1 U15603 ( .IN1(n9727), .IN2(CRC_OUT_8_30), .Q(n15232) );
  AND2X1 U15604 ( .IN1(n15234), .IN2(n10588), .Q(WX2617) );
  AND2X1 U15605 ( .IN1(n15235), .IN2(n15236), .Q(n15234) );
  OR2X1 U15606 ( .IN1(DFF_381_n1), .IN2(WX2132), .Q(n15236) );
  OR2X1 U15607 ( .IN1(n9728), .IN2(CRC_OUT_8_29), .Q(n15235) );
  AND2X1 U15608 ( .IN1(n15237), .IN2(n10587), .Q(WX2615) );
  AND2X1 U15609 ( .IN1(n15238), .IN2(n15239), .Q(n15237) );
  OR2X1 U15610 ( .IN1(DFF_380_n1), .IN2(WX2134), .Q(n15239) );
  OR2X1 U15611 ( .IN1(n9729), .IN2(CRC_OUT_8_28), .Q(n15238) );
  AND2X1 U15612 ( .IN1(n15240), .IN2(n10586), .Q(WX2613) );
  OR2X1 U15613 ( .IN1(n15241), .IN2(n15242), .Q(n15240) );
  AND2X1 U15614 ( .IN1(DFF_379_n1), .IN2(n9912), .Q(n15242) );
  AND2X1 U15615 ( .IN1(test_so18), .IN2(CRC_OUT_8_27), .Q(n15241) );
  AND2X1 U15616 ( .IN1(n15243), .IN2(n10587), .Q(WX2611) );
  AND2X1 U15617 ( .IN1(n15244), .IN2(n15245), .Q(n15243) );
  OR2X1 U15618 ( .IN1(DFF_378_n1), .IN2(WX2138), .Q(n15245) );
  OR2X1 U15619 ( .IN1(n9730), .IN2(CRC_OUT_8_26), .Q(n15244) );
  AND2X1 U15620 ( .IN1(n15246), .IN2(n10587), .Q(WX2609) );
  OR2X1 U15621 ( .IN1(n15247), .IN2(n15248), .Q(n15246) );
  AND2X1 U15622 ( .IN1(n9731), .IN2(n9946), .Q(n15248) );
  AND2X1 U15623 ( .IN1(test_so21), .IN2(WX2140), .Q(n15247) );
  AND2X1 U15624 ( .IN1(n15249), .IN2(n10587), .Q(WX2607) );
  AND2X1 U15625 ( .IN1(n15250), .IN2(n15251), .Q(n15249) );
  OR2X1 U15626 ( .IN1(DFF_376_n1), .IN2(WX2142), .Q(n15251) );
  OR2X1 U15627 ( .IN1(n9732), .IN2(CRC_OUT_8_24), .Q(n15250) );
  AND2X1 U15628 ( .IN1(n15252), .IN2(n10585), .Q(WX2605) );
  AND2X1 U15629 ( .IN1(n15253), .IN2(n15254), .Q(n15252) );
  OR2X1 U15630 ( .IN1(DFF_375_n1), .IN2(WX2144), .Q(n15254) );
  OR2X1 U15631 ( .IN1(n9733), .IN2(CRC_OUT_8_23), .Q(n15253) );
  AND2X1 U15632 ( .IN1(n15255), .IN2(n10587), .Q(WX2603) );
  AND2X1 U15633 ( .IN1(n15256), .IN2(n15257), .Q(n15255) );
  OR2X1 U15634 ( .IN1(DFF_374_n1), .IN2(WX2146), .Q(n15257) );
  OR2X1 U15635 ( .IN1(n9734), .IN2(CRC_OUT_8_22), .Q(n15256) );
  AND2X1 U15636 ( .IN1(n15258), .IN2(n10587), .Q(WX2601) );
  AND2X1 U15637 ( .IN1(n15259), .IN2(n15260), .Q(n15258) );
  OR2X1 U15638 ( .IN1(DFF_373_n1), .IN2(WX2148), .Q(n15260) );
  OR2X1 U15639 ( .IN1(n9735), .IN2(CRC_OUT_8_21), .Q(n15259) );
  AND2X1 U15640 ( .IN1(n15261), .IN2(n10587), .Q(WX2599) );
  AND2X1 U15641 ( .IN1(n15262), .IN2(n15263), .Q(n15261) );
  OR2X1 U15642 ( .IN1(DFF_372_n1), .IN2(WX2150), .Q(n15263) );
  OR2X1 U15643 ( .IN1(n9736), .IN2(CRC_OUT_8_20), .Q(n15262) );
  AND2X1 U15644 ( .IN1(n15264), .IN2(n10583), .Q(WX2597) );
  AND2X1 U15645 ( .IN1(n15265), .IN2(n15266), .Q(n15264) );
  OR2X1 U15646 ( .IN1(DFF_371_n1), .IN2(WX2152), .Q(n15266) );
  OR2X1 U15647 ( .IN1(n9737), .IN2(CRC_OUT_8_19), .Q(n15265) );
  AND2X1 U15648 ( .IN1(n15267), .IN2(n10584), .Q(WX2595) );
  AND2X1 U15649 ( .IN1(n15268), .IN2(n15269), .Q(n15267) );
  OR2X1 U15650 ( .IN1(DFF_370_n1), .IN2(WX2154), .Q(n15269) );
  OR2X1 U15651 ( .IN1(n9738), .IN2(CRC_OUT_8_18), .Q(n15268) );
  AND2X1 U15652 ( .IN1(n15270), .IN2(n10587), .Q(WX2593) );
  AND2X1 U15653 ( .IN1(n15271), .IN2(n15272), .Q(n15270) );
  OR2X1 U15654 ( .IN1(DFF_369_n1), .IN2(WX2156), .Q(n15272) );
  OR2X1 U15655 ( .IN1(n9739), .IN2(CRC_OUT_8_17), .Q(n15271) );
  AND2X1 U15656 ( .IN1(n15273), .IN2(n10586), .Q(WX2591) );
  AND2X1 U15657 ( .IN1(n15274), .IN2(n15275), .Q(n15273) );
  OR2X1 U15658 ( .IN1(DFF_368_n1), .IN2(WX2158), .Q(n15275) );
  OR2X1 U15659 ( .IN1(n9740), .IN2(CRC_OUT_8_16), .Q(n15274) );
  AND2X1 U15660 ( .IN1(n15276), .IN2(n10584), .Q(WX2589) );
  OR2X1 U15661 ( .IN1(n15277), .IN2(n15278), .Q(n15276) );
  AND2X1 U15662 ( .IN1(n15279), .IN2(CRC_OUT_8_15), .Q(n15278) );
  AND2X1 U15663 ( .IN1(DFF_367_n1), .IN2(n15280), .Q(n15277) );
  INVX0 U15664 ( .INP(n15279), .ZN(n15280) );
  OR2X1 U15665 ( .IN1(n15281), .IN2(n15282), .Q(n15279) );
  AND2X1 U15666 ( .IN1(DFF_383_n1), .IN2(WX2160), .Q(n15282) );
  AND2X1 U15667 ( .IN1(n9530), .IN2(CRC_OUT_8_31), .Q(n15281) );
  AND2X1 U15668 ( .IN1(n15283), .IN2(n10585), .Q(WX2587) );
  AND2X1 U15669 ( .IN1(n15284), .IN2(n15285), .Q(n15283) );
  OR2X1 U15670 ( .IN1(DFF_366_n1), .IN2(WX2162), .Q(n15285) );
  OR2X1 U15671 ( .IN1(n9741), .IN2(CRC_OUT_8_14), .Q(n15284) );
  AND2X1 U15672 ( .IN1(n15286), .IN2(n10583), .Q(WX2585) );
  AND2X1 U15673 ( .IN1(n15287), .IN2(n15288), .Q(n15286) );
  OR2X1 U15674 ( .IN1(DFF_365_n1), .IN2(WX2164), .Q(n15288) );
  OR2X1 U15675 ( .IN1(n9742), .IN2(CRC_OUT_8_13), .Q(n15287) );
  AND2X1 U15676 ( .IN1(n15289), .IN2(n10577), .Q(WX2583) );
  AND2X1 U15677 ( .IN1(n15290), .IN2(n15291), .Q(n15289) );
  OR2X1 U15678 ( .IN1(DFF_364_n1), .IN2(WX2166), .Q(n15291) );
  OR2X1 U15679 ( .IN1(n9743), .IN2(CRC_OUT_8_12), .Q(n15290) );
  AND2X1 U15680 ( .IN1(n15292), .IN2(n10570), .Q(WX2581) );
  AND2X1 U15681 ( .IN1(n15293), .IN2(n15294), .Q(n15292) );
  OR2X1 U15682 ( .IN1(DFF_363_n1), .IN2(WX2168), .Q(n15294) );
  OR2X1 U15683 ( .IN1(n9744), .IN2(CRC_OUT_8_11), .Q(n15293) );
  AND2X1 U15684 ( .IN1(n15295), .IN2(n10571), .Q(WX2579) );
  OR2X1 U15685 ( .IN1(n15296), .IN2(n15297), .Q(n15295) );
  AND2X1 U15686 ( .IN1(n15298), .IN2(CRC_OUT_8_10), .Q(n15297) );
  AND2X1 U15687 ( .IN1(DFF_362_n1), .IN2(n15299), .Q(n15296) );
  INVX0 U15688 ( .INP(n15298), .ZN(n15299) );
  OR2X1 U15689 ( .IN1(n15300), .IN2(n15301), .Q(n15298) );
  AND2X1 U15690 ( .IN1(DFF_383_n1), .IN2(WX2170), .Q(n15301) );
  AND2X1 U15691 ( .IN1(n9531), .IN2(CRC_OUT_8_31), .Q(n15300) );
  AND2X1 U15692 ( .IN1(n15302), .IN2(n10571), .Q(WX2577) );
  OR2X1 U15693 ( .IN1(n15303), .IN2(n15304), .Q(n15302) );
  AND2X1 U15694 ( .IN1(DFF_361_n1), .IN2(n9905), .Q(n15304) );
  AND2X1 U15695 ( .IN1(test_so19), .IN2(CRC_OUT_8_9), .Q(n15303) );
  AND2X1 U15696 ( .IN1(n15305), .IN2(n10571), .Q(WX2575) );
  AND2X1 U15697 ( .IN1(n15306), .IN2(n15307), .Q(n15305) );
  OR2X1 U15698 ( .IN1(DFF_360_n1), .IN2(WX2174), .Q(n15307) );
  OR2X1 U15699 ( .IN1(n9745), .IN2(CRC_OUT_8_8), .Q(n15306) );
  AND2X1 U15700 ( .IN1(n15308), .IN2(n10571), .Q(WX2573) );
  OR2X1 U15701 ( .IN1(n15309), .IN2(n15310), .Q(n15308) );
  AND2X1 U15702 ( .IN1(n9746), .IN2(n9947), .Q(n15310) );
  AND2X1 U15703 ( .IN1(test_so20), .IN2(WX2176), .Q(n15309) );
  AND2X1 U15704 ( .IN1(n15311), .IN2(n10571), .Q(WX2571) );
  AND2X1 U15705 ( .IN1(n15312), .IN2(n15313), .Q(n15311) );
  OR2X1 U15706 ( .IN1(DFF_358_n1), .IN2(WX2178), .Q(n15313) );
  OR2X1 U15707 ( .IN1(n9747), .IN2(CRC_OUT_8_6), .Q(n15312) );
  AND2X1 U15708 ( .IN1(n15314), .IN2(n10571), .Q(WX2569) );
  AND2X1 U15709 ( .IN1(n15315), .IN2(n15316), .Q(n15314) );
  OR2X1 U15710 ( .IN1(DFF_357_n1), .IN2(WX2180), .Q(n15316) );
  OR2X1 U15711 ( .IN1(n9748), .IN2(CRC_OUT_8_5), .Q(n15315) );
  AND2X1 U15712 ( .IN1(n15317), .IN2(n10571), .Q(WX2567) );
  AND2X1 U15713 ( .IN1(n15318), .IN2(n15319), .Q(n15317) );
  OR2X1 U15714 ( .IN1(DFF_356_n1), .IN2(WX2182), .Q(n15319) );
  OR2X1 U15715 ( .IN1(n9749), .IN2(CRC_OUT_8_4), .Q(n15318) );
  AND2X1 U15716 ( .IN1(n15320), .IN2(n10571), .Q(WX2565) );
  OR2X1 U15717 ( .IN1(n15321), .IN2(n15322), .Q(n15320) );
  AND2X1 U15718 ( .IN1(n15323), .IN2(CRC_OUT_8_3), .Q(n15322) );
  AND2X1 U15719 ( .IN1(DFF_355_n1), .IN2(n15324), .Q(n15321) );
  INVX0 U15720 ( .INP(n15323), .ZN(n15324) );
  OR2X1 U15721 ( .IN1(n15325), .IN2(n15326), .Q(n15323) );
  AND2X1 U15722 ( .IN1(DFF_383_n1), .IN2(WX2184), .Q(n15326) );
  AND2X1 U15723 ( .IN1(n9532), .IN2(CRC_OUT_8_31), .Q(n15325) );
  AND2X1 U15724 ( .IN1(n15327), .IN2(n10571), .Q(WX2563) );
  AND2X1 U15725 ( .IN1(n15328), .IN2(n15329), .Q(n15327) );
  OR2X1 U15726 ( .IN1(DFF_354_n1), .IN2(WX2186), .Q(n15329) );
  OR2X1 U15727 ( .IN1(n9750), .IN2(CRC_OUT_8_2), .Q(n15328) );
  AND2X1 U15728 ( .IN1(n15330), .IN2(n10572), .Q(WX2561) );
  AND2X1 U15729 ( .IN1(n15331), .IN2(n15332), .Q(n15330) );
  OR2X1 U15730 ( .IN1(DFF_353_n1), .IN2(WX2188), .Q(n15332) );
  OR2X1 U15731 ( .IN1(n9751), .IN2(CRC_OUT_8_1), .Q(n15331) );
  AND2X1 U15732 ( .IN1(n15333), .IN2(n10572), .Q(WX2559) );
  AND2X1 U15733 ( .IN1(n15334), .IN2(n15335), .Q(n15333) );
  OR2X1 U15734 ( .IN1(DFF_352_n1), .IN2(WX2190), .Q(n15335) );
  OR2X1 U15735 ( .IN1(n9752), .IN2(CRC_OUT_8_0), .Q(n15334) );
  AND2X1 U15736 ( .IN1(n15336), .IN2(n10572), .Q(WX2557) );
  AND2X1 U15737 ( .IN1(n15337), .IN2(n15338), .Q(n15336) );
  OR2X1 U15738 ( .IN1(DFF_383_n1), .IN2(WX2192), .Q(n15338) );
  OR2X1 U15739 ( .IN1(n9540), .IN2(CRC_OUT_8_31), .Q(n15337) );
  AND2X1 U15740 ( .IN1(n10601), .IN2(n8653), .Q(WX2031) );
  AND2X1 U15741 ( .IN1(n10601), .IN2(n8654), .Q(WX2029) );
  AND2X1 U15742 ( .IN1(n10601), .IN2(n8655), .Q(WX2027) );
  AND2X1 U15743 ( .IN1(n10601), .IN2(n8656), .Q(WX2025) );
  AND2X1 U15744 ( .IN1(n10601), .IN2(n8657), .Q(WX2023) );
  AND2X1 U15745 ( .IN1(n10600), .IN2(n8658), .Q(WX2021) );
  AND2X1 U15746 ( .IN1(test_so13), .IN2(n10572), .Q(WX2019) );
  AND2X1 U15747 ( .IN1(n10600), .IN2(n8661), .Q(WX2017) );
  AND2X1 U15748 ( .IN1(n10600), .IN2(n8662), .Q(WX2015) );
  AND2X1 U15749 ( .IN1(n10600), .IN2(n8663), .Q(WX2013) );
  AND2X1 U15750 ( .IN1(n10600), .IN2(n8664), .Q(WX2011) );
  AND2X1 U15751 ( .IN1(n10600), .IN2(n8665), .Q(WX2009) );
  AND2X1 U15752 ( .IN1(n10600), .IN2(n8666), .Q(WX2007) );
  AND2X1 U15753 ( .IN1(n10600), .IN2(n8667), .Q(WX2005) );
  AND2X1 U15754 ( .IN1(n10599), .IN2(n8668), .Q(WX2003) );
  AND2X1 U15755 ( .IN1(n10599), .IN2(n8669), .Q(WX2001) );
  OR2X1 U15756 ( .IN1(n15339), .IN2(n15340), .Q(WX1999) );
  OR2X1 U15757 ( .IN1(n15341), .IN2(n15342), .Q(n15340) );
  AND2X1 U15758 ( .IN1(n10032), .IN2(CRC_OUT_8_0), .Q(n15342) );
  AND2X1 U15759 ( .IN1(n280), .IN2(n10006), .Q(n15341) );
  INVX0 U15760 ( .INP(n15343), .ZN(n280) );
  OR2X1 U15761 ( .IN1(n10634), .IN2(n4003), .Q(n15343) );
  OR2X1 U15762 ( .IN1(n15344), .IN2(n15345), .Q(n15339) );
  AND2X1 U15763 ( .IN1(n10067), .IN2(n14585), .Q(n15345) );
  OR2X1 U15764 ( .IN1(n15346), .IN2(n15347), .Q(n14585) );
  INVX0 U15765 ( .INP(n15348), .ZN(n15347) );
  OR2X1 U15766 ( .IN1(n15349), .IN2(n15350), .Q(n15348) );
  AND2X1 U15767 ( .IN1(n15350), .IN2(n15349), .Q(n15346) );
  AND2X1 U15768 ( .IN1(n15351), .IN2(n15352), .Q(n15349) );
  OR2X1 U15769 ( .IN1(WX3357), .IN2(n9451), .Q(n15352) );
  OR2X1 U15770 ( .IN1(WX3293), .IN2(n3723), .Q(n15351) );
  OR2X1 U15771 ( .IN1(n15353), .IN2(n15354), .Q(n15350) );
  AND2X1 U15772 ( .IN1(n9452), .IN2(WX3485), .Q(n15354) );
  AND2X1 U15773 ( .IN1(n9539), .IN2(WX3421), .Q(n15353) );
  AND2X1 U15774 ( .IN1(n12700), .IN2(n9976), .Q(n15344) );
  AND2X1 U15775 ( .IN1(n15355), .IN2(n15356), .Q(n12700) );
  INVX0 U15776 ( .INP(n15357), .ZN(n15356) );
  AND2X1 U15777 ( .IN1(n15358), .IN2(n15359), .Q(n15357) );
  OR2X1 U15778 ( .IN1(n15359), .IN2(n15358), .Q(n15355) );
  OR2X1 U15779 ( .IN1(n15360), .IN2(n15361), .Q(n15358) );
  AND2X1 U15780 ( .IN1(n9482), .IN2(WX2128), .Q(n15361) );
  INVX0 U15781 ( .INP(n15362), .ZN(n15360) );
  OR2X1 U15782 ( .IN1(WX2128), .IN2(n9482), .Q(n15362) );
  AND2X1 U15783 ( .IN1(n15363), .IN2(n15364), .Q(n15359) );
  OR2X1 U15784 ( .IN1(WX2192), .IN2(test_so16), .Q(n15364) );
  OR2X1 U15785 ( .IN1(n9929), .IN2(n9540), .Q(n15363) );
  OR2X1 U15786 ( .IN1(n15365), .IN2(n15366), .Q(WX1997) );
  OR2X1 U15787 ( .IN1(n15367), .IN2(n15368), .Q(n15366) );
  AND2X1 U15788 ( .IN1(n10033), .IN2(CRC_OUT_8_1), .Q(n15368) );
  AND2X1 U15789 ( .IN1(n279), .IN2(n10006), .Q(n15367) );
  INVX0 U15790 ( .INP(n15369), .ZN(n279) );
  OR2X1 U15791 ( .IN1(n10634), .IN2(n4004), .Q(n15369) );
  OR2X1 U15792 ( .IN1(n15370), .IN2(n15371), .Q(n15365) );
  AND2X1 U15793 ( .IN1(n10067), .IN2(n14603), .Q(n15371) );
  OR2X1 U15794 ( .IN1(n15372), .IN2(n15373), .Q(n14603) );
  INVX0 U15795 ( .INP(n15374), .ZN(n15373) );
  OR2X1 U15796 ( .IN1(n15375), .IN2(n15376), .Q(n15374) );
  AND2X1 U15797 ( .IN1(n15376), .IN2(n15375), .Q(n15372) );
  AND2X1 U15798 ( .IN1(n15377), .IN2(n15378), .Q(n15375) );
  OR2X1 U15799 ( .IN1(WX3355), .IN2(n9453), .Q(n15378) );
  OR2X1 U15800 ( .IN1(WX3291), .IN2(n3725), .Q(n15377) );
  OR2X1 U15801 ( .IN1(n15379), .IN2(n15380), .Q(n15376) );
  AND2X1 U15802 ( .IN1(n9454), .IN2(WX3483), .Q(n15380) );
  AND2X1 U15803 ( .IN1(n9726), .IN2(WX3419), .Q(n15379) );
  AND2X1 U15804 ( .IN1(n9988), .IN2(n12708), .Q(n15370) );
  OR2X1 U15805 ( .IN1(n15381), .IN2(n15382), .Q(n12708) );
  INVX0 U15806 ( .INP(n15383), .ZN(n15382) );
  OR2X1 U15807 ( .IN1(n15384), .IN2(n15385), .Q(n15383) );
  AND2X1 U15808 ( .IN1(n15385), .IN2(n15384), .Q(n15381) );
  AND2X1 U15809 ( .IN1(n15386), .IN2(n15387), .Q(n15384) );
  OR2X1 U15810 ( .IN1(WX2062), .IN2(n9484), .Q(n15387) );
  OR2X1 U15811 ( .IN1(WX1998), .IN2(n3757), .Q(n15386) );
  OR2X1 U15812 ( .IN1(n15388), .IN2(n15389), .Q(n15385) );
  AND2X1 U15813 ( .IN1(n9485), .IN2(WX2190), .Q(n15389) );
  AND2X1 U15814 ( .IN1(n9752), .IN2(WX2126), .Q(n15388) );
  OR2X1 U15815 ( .IN1(n15390), .IN2(n15391), .Q(WX1995) );
  OR2X1 U15816 ( .IN1(n15392), .IN2(n15393), .Q(n15391) );
  AND2X1 U15817 ( .IN1(n10033), .IN2(CRC_OUT_8_2), .Q(n15393) );
  AND2X1 U15818 ( .IN1(n278), .IN2(n10006), .Q(n15392) );
  INVX0 U15819 ( .INP(n15394), .ZN(n278) );
  OR2X1 U15820 ( .IN1(n10633), .IN2(n4005), .Q(n15394) );
  OR2X1 U15821 ( .IN1(n15395), .IN2(n15396), .Q(n15390) );
  AND2X1 U15822 ( .IN1(n10067), .IN2(n14620), .Q(n15396) );
  OR2X1 U15823 ( .IN1(n15397), .IN2(n15398), .Q(n14620) );
  INVX0 U15824 ( .INP(n15399), .ZN(n15398) );
  OR2X1 U15825 ( .IN1(n15400), .IN2(n15401), .Q(n15399) );
  AND2X1 U15826 ( .IN1(n15401), .IN2(n15400), .Q(n15397) );
  AND2X1 U15827 ( .IN1(n15402), .IN2(n15403), .Q(n15400) );
  OR2X1 U15828 ( .IN1(WX3353), .IN2(n9455), .Q(n15403) );
  OR2X1 U15829 ( .IN1(WX3289), .IN2(n3727), .Q(n15402) );
  OR2X1 U15830 ( .IN1(n15404), .IN2(n15405), .Q(n15401) );
  AND2X1 U15831 ( .IN1(n9456), .IN2(WX3481), .Q(n15405) );
  AND2X1 U15832 ( .IN1(n9725), .IN2(WX3417), .Q(n15404) );
  AND2X1 U15833 ( .IN1(n9988), .IN2(n12716), .Q(n15395) );
  OR2X1 U15834 ( .IN1(n15406), .IN2(n15407), .Q(n12716) );
  INVX0 U15835 ( .INP(n15408), .ZN(n15407) );
  OR2X1 U15836 ( .IN1(n15409), .IN2(n15410), .Q(n15408) );
  AND2X1 U15837 ( .IN1(n15410), .IN2(n15409), .Q(n15406) );
  AND2X1 U15838 ( .IN1(n15411), .IN2(n15412), .Q(n15409) );
  OR2X1 U15839 ( .IN1(WX2060), .IN2(n9486), .Q(n15412) );
  OR2X1 U15840 ( .IN1(WX1996), .IN2(n3759), .Q(n15411) );
  OR2X1 U15841 ( .IN1(n15413), .IN2(n15414), .Q(n15410) );
  AND2X1 U15842 ( .IN1(n9487), .IN2(WX2188), .Q(n15414) );
  AND2X1 U15843 ( .IN1(n9751), .IN2(WX2124), .Q(n15413) );
  OR2X1 U15844 ( .IN1(n15415), .IN2(n15416), .Q(WX1993) );
  OR2X1 U15845 ( .IN1(n15417), .IN2(n15418), .Q(n15416) );
  AND2X1 U15846 ( .IN1(n10033), .IN2(CRC_OUT_8_3), .Q(n15418) );
  AND2X1 U15847 ( .IN1(n277), .IN2(n10006), .Q(n15417) );
  INVX0 U15848 ( .INP(n15419), .ZN(n277) );
  OR2X1 U15849 ( .IN1(n10633), .IN2(n4006), .Q(n15419) );
  OR2X1 U15850 ( .IN1(n15420), .IN2(n15421), .Q(n15415) );
  AND2X1 U15851 ( .IN1(n10067), .IN2(n14637), .Q(n15421) );
  OR2X1 U15852 ( .IN1(n15422), .IN2(n15423), .Q(n14637) );
  INVX0 U15853 ( .INP(n15424), .ZN(n15423) );
  OR2X1 U15854 ( .IN1(n15425), .IN2(n15426), .Q(n15424) );
  AND2X1 U15855 ( .IN1(n15426), .IN2(n15425), .Q(n15422) );
  AND2X1 U15856 ( .IN1(n15427), .IN2(n15428), .Q(n15425) );
  OR2X1 U15857 ( .IN1(WX3351), .IN2(n9457), .Q(n15428) );
  OR2X1 U15858 ( .IN1(WX3287), .IN2(n3729), .Q(n15427) );
  OR2X1 U15859 ( .IN1(n15429), .IN2(n15430), .Q(n15426) );
  AND2X1 U15860 ( .IN1(n9458), .IN2(WX3479), .Q(n15430) );
  AND2X1 U15861 ( .IN1(n9724), .IN2(WX3415), .Q(n15429) );
  AND2X1 U15862 ( .IN1(n9988), .IN2(n12724), .Q(n15420) );
  OR2X1 U15863 ( .IN1(n15431), .IN2(n15432), .Q(n12724) );
  INVX0 U15864 ( .INP(n15433), .ZN(n15432) );
  OR2X1 U15865 ( .IN1(n15434), .IN2(n15435), .Q(n15433) );
  AND2X1 U15866 ( .IN1(n15435), .IN2(n15434), .Q(n15431) );
  AND2X1 U15867 ( .IN1(n15436), .IN2(n15437), .Q(n15434) );
  OR2X1 U15868 ( .IN1(WX2058), .IN2(n9488), .Q(n15437) );
  OR2X1 U15869 ( .IN1(WX1994), .IN2(n3761), .Q(n15436) );
  OR2X1 U15870 ( .IN1(n15438), .IN2(n15439), .Q(n15435) );
  AND2X1 U15871 ( .IN1(n9489), .IN2(WX2186), .Q(n15439) );
  AND2X1 U15872 ( .IN1(n9750), .IN2(WX2122), .Q(n15438) );
  OR2X1 U15873 ( .IN1(n15440), .IN2(n15441), .Q(WX1991) );
  OR2X1 U15874 ( .IN1(n15442), .IN2(n15443), .Q(n15441) );
  AND2X1 U15875 ( .IN1(n10033), .IN2(CRC_OUT_8_4), .Q(n15443) );
  AND2X1 U15876 ( .IN1(n276), .IN2(n10006), .Q(n15442) );
  INVX0 U15877 ( .INP(n15444), .ZN(n276) );
  OR2X1 U15878 ( .IN1(n10633), .IN2(n4007), .Q(n15444) );
  OR2X1 U15879 ( .IN1(n15445), .IN2(n15446), .Q(n15440) );
  AND2X1 U15880 ( .IN1(n10067), .IN2(n14654), .Q(n15446) );
  OR2X1 U15881 ( .IN1(n15447), .IN2(n15448), .Q(n14654) );
  INVX0 U15882 ( .INP(n15449), .ZN(n15448) );
  OR2X1 U15883 ( .IN1(n15450), .IN2(n15451), .Q(n15449) );
  AND2X1 U15884 ( .IN1(n15451), .IN2(n15450), .Q(n15447) );
  AND2X1 U15885 ( .IN1(n15452), .IN2(n15453), .Q(n15450) );
  OR2X1 U15886 ( .IN1(WX3349), .IN2(n9459), .Q(n15453) );
  OR2X1 U15887 ( .IN1(WX3285), .IN2(n3731), .Q(n15452) );
  OR2X1 U15888 ( .IN1(n15454), .IN2(n15455), .Q(n15451) );
  AND2X1 U15889 ( .IN1(n9460), .IN2(WX3477), .Q(n15455) );
  AND2X1 U15890 ( .IN1(n9529), .IN2(WX3413), .Q(n15454) );
  AND2X1 U15891 ( .IN1(n12732), .IN2(n9976), .Q(n15445) );
  AND2X1 U15892 ( .IN1(n15456), .IN2(n15457), .Q(n12732) );
  INVX0 U15893 ( .INP(n15458), .ZN(n15457) );
  AND2X1 U15894 ( .IN1(n15459), .IN2(n15460), .Q(n15458) );
  OR2X1 U15895 ( .IN1(n15460), .IN2(n15459), .Q(n15456) );
  OR2X1 U15896 ( .IN1(n15461), .IN2(n15462), .Q(n15459) );
  AND2X1 U15897 ( .IN1(n3763), .IN2(WX2120), .Q(n15462) );
  INVX0 U15898 ( .INP(n15463), .ZN(n15461) );
  OR2X1 U15899 ( .IN1(WX2120), .IN2(n3763), .Q(n15463) );
  AND2X1 U15900 ( .IN1(n15464), .IN2(n15465), .Q(n15460) );
  OR2X1 U15901 ( .IN1(WX2184), .IN2(test_so14), .Q(n15465) );
  OR2X1 U15902 ( .IN1(n9930), .IN2(n9532), .Q(n15464) );
  OR2X1 U15903 ( .IN1(n15466), .IN2(n15467), .Q(WX1989) );
  OR2X1 U15904 ( .IN1(n15468), .IN2(n15469), .Q(n15467) );
  AND2X1 U15905 ( .IN1(n10033), .IN2(CRC_OUT_8_5), .Q(n15469) );
  AND2X1 U15906 ( .IN1(n275), .IN2(n10007), .Q(n15468) );
  INVX0 U15907 ( .INP(n15470), .ZN(n275) );
  OR2X1 U15908 ( .IN1(n10633), .IN2(n4008), .Q(n15470) );
  OR2X1 U15909 ( .IN1(n15471), .IN2(n15472), .Q(n15466) );
  AND2X1 U15910 ( .IN1(n10067), .IN2(n14671), .Q(n15472) );
  OR2X1 U15911 ( .IN1(n15473), .IN2(n15474), .Q(n14671) );
  INVX0 U15912 ( .INP(n15475), .ZN(n15474) );
  OR2X1 U15913 ( .IN1(n15476), .IN2(n15477), .Q(n15475) );
  AND2X1 U15914 ( .IN1(n15477), .IN2(n15476), .Q(n15473) );
  AND2X1 U15915 ( .IN1(n15478), .IN2(n15479), .Q(n15476) );
  OR2X1 U15916 ( .IN1(WX3347), .IN2(n9461), .Q(n15479) );
  OR2X1 U15917 ( .IN1(WX3283), .IN2(n3733), .Q(n15478) );
  OR2X1 U15918 ( .IN1(n15480), .IN2(n15481), .Q(n15477) );
  AND2X1 U15919 ( .IN1(n9462), .IN2(WX3475), .Q(n15481) );
  AND2X1 U15920 ( .IN1(n9723), .IN2(WX3411), .Q(n15480) );
  AND2X1 U15921 ( .IN1(n9988), .IN2(n12740), .Q(n15471) );
  OR2X1 U15922 ( .IN1(n15482), .IN2(n15483), .Q(n12740) );
  INVX0 U15923 ( .INP(n15484), .ZN(n15483) );
  OR2X1 U15924 ( .IN1(n15485), .IN2(n15486), .Q(n15484) );
  AND2X1 U15925 ( .IN1(n15486), .IN2(n15485), .Q(n15482) );
  AND2X1 U15926 ( .IN1(n15487), .IN2(n15488), .Q(n15485) );
  OR2X1 U15927 ( .IN1(WX2054), .IN2(n9491), .Q(n15488) );
  OR2X1 U15928 ( .IN1(WX1990), .IN2(n3765), .Q(n15487) );
  OR2X1 U15929 ( .IN1(n15489), .IN2(n15490), .Q(n15486) );
  AND2X1 U15930 ( .IN1(n9492), .IN2(WX2182), .Q(n15490) );
  AND2X1 U15931 ( .IN1(n9749), .IN2(WX2118), .Q(n15489) );
  OR2X1 U15932 ( .IN1(n15491), .IN2(n15492), .Q(WX1987) );
  OR2X1 U15933 ( .IN1(n15493), .IN2(n15494), .Q(n15492) );
  AND2X1 U15934 ( .IN1(n10033), .IN2(CRC_OUT_8_6), .Q(n15494) );
  AND2X1 U15935 ( .IN1(n274), .IN2(n10007), .Q(n15493) );
  INVX0 U15936 ( .INP(n15495), .ZN(n274) );
  OR2X1 U15937 ( .IN1(n10633), .IN2(n4009), .Q(n15495) );
  OR2X1 U15938 ( .IN1(n15496), .IN2(n15497), .Q(n15491) );
  AND2X1 U15939 ( .IN1(n14688), .IN2(n10059), .Q(n15497) );
  AND2X1 U15940 ( .IN1(n15498), .IN2(n15499), .Q(n14688) );
  INVX0 U15941 ( .INP(n15500), .ZN(n15499) );
  AND2X1 U15942 ( .IN1(n15501), .IN2(n15502), .Q(n15500) );
  OR2X1 U15943 ( .IN1(n15502), .IN2(n15501), .Q(n15498) );
  OR2X1 U15944 ( .IN1(n15503), .IN2(n15504), .Q(n15501) );
  AND2X1 U15945 ( .IN1(n3735), .IN2(WX3281), .Q(n15504) );
  INVX0 U15946 ( .INP(n15505), .ZN(n15503) );
  OR2X1 U15947 ( .IN1(WX3281), .IN2(n3735), .Q(n15505) );
  AND2X1 U15948 ( .IN1(n15506), .IN2(n15507), .Q(n15502) );
  OR2X1 U15949 ( .IN1(WX3409), .IN2(test_so30), .Q(n15507) );
  OR2X1 U15950 ( .IN1(n9904), .IN2(n9464), .Q(n15506) );
  AND2X1 U15951 ( .IN1(n9988), .IN2(n12748), .Q(n15496) );
  OR2X1 U15952 ( .IN1(n15508), .IN2(n15509), .Q(n12748) );
  INVX0 U15953 ( .INP(n15510), .ZN(n15509) );
  OR2X1 U15954 ( .IN1(n15511), .IN2(n15512), .Q(n15510) );
  AND2X1 U15955 ( .IN1(n15512), .IN2(n15511), .Q(n15508) );
  AND2X1 U15956 ( .IN1(n15513), .IN2(n15514), .Q(n15511) );
  OR2X1 U15957 ( .IN1(WX2052), .IN2(n9493), .Q(n15514) );
  OR2X1 U15958 ( .IN1(WX1988), .IN2(n3767), .Q(n15513) );
  OR2X1 U15959 ( .IN1(n15515), .IN2(n15516), .Q(n15512) );
  AND2X1 U15960 ( .IN1(n9494), .IN2(WX2180), .Q(n15516) );
  AND2X1 U15961 ( .IN1(n9748), .IN2(WX2116), .Q(n15515) );
  OR2X1 U15962 ( .IN1(n15517), .IN2(n15518), .Q(WX1985) );
  OR2X1 U15963 ( .IN1(n15519), .IN2(n15520), .Q(n15518) );
  AND2X1 U15964 ( .IN1(test_so20), .IN2(n10026), .Q(n15520) );
  AND2X1 U15965 ( .IN1(n273), .IN2(n10007), .Q(n15519) );
  INVX0 U15966 ( .INP(n15521), .ZN(n273) );
  OR2X1 U15967 ( .IN1(n10633), .IN2(n4010), .Q(n15521) );
  OR2X1 U15968 ( .IN1(n15522), .IN2(n15523), .Q(n15517) );
  AND2X1 U15969 ( .IN1(n10067), .IN2(n14705), .Q(n15523) );
  OR2X1 U15970 ( .IN1(n15524), .IN2(n15525), .Q(n14705) );
  INVX0 U15971 ( .INP(n15526), .ZN(n15525) );
  OR2X1 U15972 ( .IN1(n15527), .IN2(n15528), .Q(n15526) );
  AND2X1 U15973 ( .IN1(n15528), .IN2(n15527), .Q(n15524) );
  AND2X1 U15974 ( .IN1(n15529), .IN2(n15530), .Q(n15527) );
  OR2X1 U15975 ( .IN1(WX3343), .IN2(n9465), .Q(n15530) );
  OR2X1 U15976 ( .IN1(WX3279), .IN2(n3737), .Q(n15529) );
  OR2X1 U15977 ( .IN1(n15531), .IN2(n15532), .Q(n15528) );
  AND2X1 U15978 ( .IN1(n9466), .IN2(WX3471), .Q(n15532) );
  AND2X1 U15979 ( .IN1(n9722), .IN2(WX3407), .Q(n15531) );
  AND2X1 U15980 ( .IN1(n9988), .IN2(n12756), .Q(n15522) );
  OR2X1 U15981 ( .IN1(n15533), .IN2(n15534), .Q(n12756) );
  INVX0 U15982 ( .INP(n15535), .ZN(n15534) );
  OR2X1 U15983 ( .IN1(n15536), .IN2(n15537), .Q(n15535) );
  AND2X1 U15984 ( .IN1(n15537), .IN2(n15536), .Q(n15533) );
  AND2X1 U15985 ( .IN1(n15538), .IN2(n15539), .Q(n15536) );
  OR2X1 U15986 ( .IN1(WX2050), .IN2(n9495), .Q(n15539) );
  OR2X1 U15987 ( .IN1(WX1986), .IN2(n3769), .Q(n15538) );
  OR2X1 U15988 ( .IN1(n15540), .IN2(n15541), .Q(n15537) );
  AND2X1 U15989 ( .IN1(n9496), .IN2(WX2178), .Q(n15541) );
  AND2X1 U15990 ( .IN1(n9747), .IN2(WX2114), .Q(n15540) );
  OR2X1 U15991 ( .IN1(n15542), .IN2(n15543), .Q(WX1983) );
  OR2X1 U15992 ( .IN1(n15544), .IN2(n15545), .Q(n15543) );
  AND2X1 U15993 ( .IN1(n10033), .IN2(CRC_OUT_8_8), .Q(n15545) );
  AND2X1 U15994 ( .IN1(n272), .IN2(n10007), .Q(n15544) );
  INVX0 U15995 ( .INP(n15546), .ZN(n272) );
  OR2X1 U15996 ( .IN1(n10633), .IN2(n4011), .Q(n15546) );
  OR2X1 U15997 ( .IN1(n15547), .IN2(n15548), .Q(n15542) );
  AND2X1 U15998 ( .IN1(n14722), .IN2(n10059), .Q(n15548) );
  AND2X1 U15999 ( .IN1(n15549), .IN2(n15550), .Q(n14722) );
  INVX0 U16000 ( .INP(n15551), .ZN(n15550) );
  AND2X1 U16001 ( .IN1(n15552), .IN2(n15553), .Q(n15551) );
  OR2X1 U16002 ( .IN1(n15553), .IN2(n15552), .Q(n15549) );
  OR2X1 U16003 ( .IN1(n15554), .IN2(n15555), .Q(n15552) );
  AND2X1 U16004 ( .IN1(n3739), .IN2(WX3277), .Q(n15555) );
  INVX0 U16005 ( .INP(n15556), .ZN(n15554) );
  OR2X1 U16006 ( .IN1(WX3277), .IN2(n3739), .Q(n15556) );
  AND2X1 U16007 ( .IN1(n15557), .IN2(n15558), .Q(n15553) );
  OR2X1 U16008 ( .IN1(WX3469), .IN2(test_so28), .Q(n15558) );
  OR2X1 U16009 ( .IN1(n9931), .IN2(n9721), .Q(n15557) );
  AND2X1 U16010 ( .IN1(n9988), .IN2(n12764), .Q(n15547) );
  OR2X1 U16011 ( .IN1(n15559), .IN2(n15560), .Q(n12764) );
  INVX0 U16012 ( .INP(n15561), .ZN(n15560) );
  OR2X1 U16013 ( .IN1(n15562), .IN2(n15563), .Q(n15561) );
  AND2X1 U16014 ( .IN1(n15563), .IN2(n15562), .Q(n15559) );
  AND2X1 U16015 ( .IN1(n15564), .IN2(n15565), .Q(n15562) );
  OR2X1 U16016 ( .IN1(WX2048), .IN2(n9497), .Q(n15565) );
  OR2X1 U16017 ( .IN1(WX1984), .IN2(n3771), .Q(n15564) );
  OR2X1 U16018 ( .IN1(n15566), .IN2(n15567), .Q(n15563) );
  AND2X1 U16019 ( .IN1(n9498), .IN2(WX2176), .Q(n15567) );
  AND2X1 U16020 ( .IN1(n9746), .IN2(WX2112), .Q(n15566) );
  OR2X1 U16021 ( .IN1(n15568), .IN2(n15569), .Q(WX1981) );
  OR2X1 U16022 ( .IN1(n15570), .IN2(n15571), .Q(n15569) );
  AND2X1 U16023 ( .IN1(n10033), .IN2(CRC_OUT_8_9), .Q(n15571) );
  AND2X1 U16024 ( .IN1(n271), .IN2(n10007), .Q(n15570) );
  INVX0 U16025 ( .INP(n15572), .ZN(n271) );
  OR2X1 U16026 ( .IN1(n10633), .IN2(n4012), .Q(n15572) );
  OR2X1 U16027 ( .IN1(n15573), .IN2(n15574), .Q(n15568) );
  AND2X1 U16028 ( .IN1(n10067), .IN2(n14739), .Q(n15574) );
  OR2X1 U16029 ( .IN1(n15575), .IN2(n15576), .Q(n14739) );
  INVX0 U16030 ( .INP(n15577), .ZN(n15576) );
  OR2X1 U16031 ( .IN1(n15578), .IN2(n15579), .Q(n15577) );
  AND2X1 U16032 ( .IN1(n15579), .IN2(n15578), .Q(n15575) );
  AND2X1 U16033 ( .IN1(n15580), .IN2(n15581), .Q(n15578) );
  OR2X1 U16034 ( .IN1(WX3339), .IN2(n9468), .Q(n15581) );
  OR2X1 U16035 ( .IN1(WX3275), .IN2(n3741), .Q(n15580) );
  OR2X1 U16036 ( .IN1(n15582), .IN2(n15583), .Q(n15579) );
  AND2X1 U16037 ( .IN1(n9469), .IN2(WX3467), .Q(n15583) );
  AND2X1 U16038 ( .IN1(n9720), .IN2(WX3403), .Q(n15582) );
  AND2X1 U16039 ( .IN1(n9987), .IN2(n12772), .Q(n15573) );
  OR2X1 U16040 ( .IN1(n15584), .IN2(n15585), .Q(n12772) );
  INVX0 U16041 ( .INP(n15586), .ZN(n15585) );
  OR2X1 U16042 ( .IN1(n15587), .IN2(n15588), .Q(n15586) );
  AND2X1 U16043 ( .IN1(n15588), .IN2(n15587), .Q(n15584) );
  AND2X1 U16044 ( .IN1(n15589), .IN2(n15590), .Q(n15587) );
  OR2X1 U16045 ( .IN1(WX2046), .IN2(n9499), .Q(n15590) );
  OR2X1 U16046 ( .IN1(WX1982), .IN2(n3773), .Q(n15589) );
  OR2X1 U16047 ( .IN1(n15591), .IN2(n15592), .Q(n15588) );
  AND2X1 U16048 ( .IN1(n9500), .IN2(WX2174), .Q(n15592) );
  AND2X1 U16049 ( .IN1(n9745), .IN2(WX2110), .Q(n15591) );
  OR2X1 U16050 ( .IN1(n15593), .IN2(n15594), .Q(WX1979) );
  OR2X1 U16051 ( .IN1(n15595), .IN2(n15596), .Q(n15594) );
  AND2X1 U16052 ( .IN1(n10033), .IN2(CRC_OUT_8_10), .Q(n15596) );
  AND2X1 U16053 ( .IN1(n270), .IN2(n10007), .Q(n15595) );
  INVX0 U16054 ( .INP(n15597), .ZN(n270) );
  OR2X1 U16055 ( .IN1(n10633), .IN2(n4013), .Q(n15597) );
  OR2X1 U16056 ( .IN1(n15598), .IN2(n15599), .Q(n15593) );
  AND2X1 U16057 ( .IN1(n10067), .IN2(n14756), .Q(n15599) );
  OR2X1 U16058 ( .IN1(n15600), .IN2(n15601), .Q(n14756) );
  INVX0 U16059 ( .INP(n15602), .ZN(n15601) );
  OR2X1 U16060 ( .IN1(n15603), .IN2(n15604), .Q(n15602) );
  AND2X1 U16061 ( .IN1(n15604), .IN2(n15603), .Q(n15600) );
  AND2X1 U16062 ( .IN1(n15605), .IN2(n15606), .Q(n15603) );
  OR2X1 U16063 ( .IN1(WX3337), .IN2(n9470), .Q(n15606) );
  OR2X1 U16064 ( .IN1(WX3273), .IN2(n3743), .Q(n15605) );
  OR2X1 U16065 ( .IN1(n15607), .IN2(n15608), .Q(n15604) );
  AND2X1 U16066 ( .IN1(n9471), .IN2(WX3465), .Q(n15608) );
  AND2X1 U16067 ( .IN1(n9719), .IN2(WX3401), .Q(n15607) );
  AND2X1 U16068 ( .IN1(n12780), .IN2(n9975), .Q(n15598) );
  AND2X1 U16069 ( .IN1(n15609), .IN2(n15610), .Q(n12780) );
  INVX0 U16070 ( .INP(n15611), .ZN(n15610) );
  AND2X1 U16071 ( .IN1(n15612), .IN2(n15613), .Q(n15611) );
  OR2X1 U16072 ( .IN1(n15613), .IN2(n15612), .Q(n15609) );
  OR2X1 U16073 ( .IN1(n15614), .IN2(n15615), .Q(n15612) );
  AND2X1 U16074 ( .IN1(n3775), .IN2(WX1980), .Q(n15615) );
  INVX0 U16075 ( .INP(n15616), .ZN(n15614) );
  OR2X1 U16076 ( .IN1(WX1980), .IN2(n3775), .Q(n15616) );
  AND2X1 U16077 ( .IN1(n15617), .IN2(n15618), .Q(n15613) );
  OR2X1 U16078 ( .IN1(WX2108), .IN2(test_so19), .Q(n15618) );
  OR2X1 U16079 ( .IN1(n9905), .IN2(n9502), .Q(n15617) );
  OR2X1 U16080 ( .IN1(n15619), .IN2(n15620), .Q(WX1977) );
  OR2X1 U16081 ( .IN1(n15621), .IN2(n15622), .Q(n15620) );
  AND2X1 U16082 ( .IN1(n10033), .IN2(CRC_OUT_8_11), .Q(n15622) );
  AND2X1 U16083 ( .IN1(n269), .IN2(n10007), .Q(n15621) );
  INVX0 U16084 ( .INP(n15623), .ZN(n269) );
  OR2X1 U16085 ( .IN1(n10633), .IN2(n4014), .Q(n15623) );
  OR2X1 U16086 ( .IN1(n15624), .IN2(n15625), .Q(n15619) );
  AND2X1 U16087 ( .IN1(n10067), .IN2(n14773), .Q(n15625) );
  OR2X1 U16088 ( .IN1(n15626), .IN2(n15627), .Q(n14773) );
  INVX0 U16089 ( .INP(n15628), .ZN(n15627) );
  OR2X1 U16090 ( .IN1(n15629), .IN2(n15630), .Q(n15628) );
  AND2X1 U16091 ( .IN1(n15630), .IN2(n15629), .Q(n15626) );
  AND2X1 U16092 ( .IN1(n15631), .IN2(n15632), .Q(n15629) );
  OR2X1 U16093 ( .IN1(WX3335), .IN2(n9472), .Q(n15632) );
  OR2X1 U16094 ( .IN1(WX3271), .IN2(n3745), .Q(n15631) );
  OR2X1 U16095 ( .IN1(n15633), .IN2(n15634), .Q(n15630) );
  AND2X1 U16096 ( .IN1(n9473), .IN2(WX3463), .Q(n15634) );
  AND2X1 U16097 ( .IN1(n9528), .IN2(WX3399), .Q(n15633) );
  AND2X1 U16098 ( .IN1(n9987), .IN2(n12788), .Q(n15624) );
  OR2X1 U16099 ( .IN1(n15635), .IN2(n15636), .Q(n12788) );
  INVX0 U16100 ( .INP(n15637), .ZN(n15636) );
  OR2X1 U16101 ( .IN1(n15638), .IN2(n15639), .Q(n15637) );
  AND2X1 U16102 ( .IN1(n15639), .IN2(n15638), .Q(n15635) );
  AND2X1 U16103 ( .IN1(n15640), .IN2(n15641), .Q(n15638) );
  OR2X1 U16104 ( .IN1(WX2042), .IN2(n9503), .Q(n15641) );
  OR2X1 U16105 ( .IN1(WX1978), .IN2(n3777), .Q(n15640) );
  OR2X1 U16106 ( .IN1(n15642), .IN2(n15643), .Q(n15639) );
  AND2X1 U16107 ( .IN1(n9504), .IN2(WX2170), .Q(n15643) );
  AND2X1 U16108 ( .IN1(n9531), .IN2(WX2106), .Q(n15642) );
  OR2X1 U16109 ( .IN1(n15644), .IN2(n15645), .Q(WX1975) );
  OR2X1 U16110 ( .IN1(n15646), .IN2(n15647), .Q(n15645) );
  AND2X1 U16111 ( .IN1(n10033), .IN2(CRC_OUT_8_12), .Q(n15647) );
  AND2X1 U16112 ( .IN1(n268), .IN2(n10007), .Q(n15646) );
  INVX0 U16113 ( .INP(n15648), .ZN(n268) );
  OR2X1 U16114 ( .IN1(n10633), .IN2(n4015), .Q(n15648) );
  OR2X1 U16115 ( .IN1(n15649), .IN2(n15650), .Q(n15644) );
  AND2X1 U16116 ( .IN1(n14791), .IN2(n10059), .Q(n15650) );
  AND2X1 U16117 ( .IN1(n15651), .IN2(n15652), .Q(n14791) );
  INVX0 U16118 ( .INP(n15653), .ZN(n15652) );
  AND2X1 U16119 ( .IN1(n15654), .IN2(n15655), .Q(n15653) );
  OR2X1 U16120 ( .IN1(n15655), .IN2(n15654), .Q(n15651) );
  OR2X1 U16121 ( .IN1(n15656), .IN2(n15657), .Q(n15654) );
  AND2X1 U16122 ( .IN1(n9474), .IN2(WX3397), .Q(n15657) );
  INVX0 U16123 ( .INP(n15658), .ZN(n15656) );
  OR2X1 U16124 ( .IN1(WX3397), .IN2(n9474), .Q(n15658) );
  AND2X1 U16125 ( .IN1(n15659), .IN2(n15660), .Q(n15655) );
  OR2X1 U16126 ( .IN1(WX3461), .IN2(test_so26), .Q(n15660) );
  OR2X1 U16127 ( .IN1(n9932), .IN2(n9718), .Q(n15659) );
  AND2X1 U16128 ( .IN1(n9987), .IN2(n12796), .Q(n15649) );
  OR2X1 U16129 ( .IN1(n15661), .IN2(n15662), .Q(n12796) );
  INVX0 U16130 ( .INP(n15663), .ZN(n15662) );
  OR2X1 U16131 ( .IN1(n15664), .IN2(n15665), .Q(n15663) );
  AND2X1 U16132 ( .IN1(n15665), .IN2(n15664), .Q(n15661) );
  AND2X1 U16133 ( .IN1(n15666), .IN2(n15667), .Q(n15664) );
  OR2X1 U16134 ( .IN1(WX2040), .IN2(n9505), .Q(n15667) );
  OR2X1 U16135 ( .IN1(WX1976), .IN2(n3779), .Q(n15666) );
  OR2X1 U16136 ( .IN1(n15668), .IN2(n15669), .Q(n15665) );
  AND2X1 U16137 ( .IN1(n9506), .IN2(WX2168), .Q(n15669) );
  AND2X1 U16138 ( .IN1(n9744), .IN2(WX2104), .Q(n15668) );
  OR2X1 U16139 ( .IN1(n15670), .IN2(n15671), .Q(WX1973) );
  OR2X1 U16140 ( .IN1(n15672), .IN2(n15673), .Q(n15671) );
  AND2X1 U16141 ( .IN1(n10033), .IN2(CRC_OUT_8_13), .Q(n15673) );
  AND2X1 U16142 ( .IN1(n267), .IN2(n10007), .Q(n15672) );
  INVX0 U16143 ( .INP(n15674), .ZN(n267) );
  OR2X1 U16144 ( .IN1(n10633), .IN2(n4016), .Q(n15674) );
  OR2X1 U16145 ( .IN1(n15675), .IN2(n15676), .Q(n15670) );
  AND2X1 U16146 ( .IN1(n10068), .IN2(n14808), .Q(n15676) );
  OR2X1 U16147 ( .IN1(n15677), .IN2(n15678), .Q(n14808) );
  INVX0 U16148 ( .INP(n15679), .ZN(n15678) );
  OR2X1 U16149 ( .IN1(n15680), .IN2(n15681), .Q(n15679) );
  AND2X1 U16150 ( .IN1(n15681), .IN2(n15680), .Q(n15677) );
  AND2X1 U16151 ( .IN1(n15682), .IN2(n15683), .Q(n15680) );
  OR2X1 U16152 ( .IN1(WX3331), .IN2(n9476), .Q(n15683) );
  OR2X1 U16153 ( .IN1(WX3267), .IN2(n3749), .Q(n15682) );
  OR2X1 U16154 ( .IN1(n15684), .IN2(n15685), .Q(n15681) );
  AND2X1 U16155 ( .IN1(n9477), .IN2(WX3459), .Q(n15685) );
  AND2X1 U16156 ( .IN1(n9717), .IN2(WX3395), .Q(n15684) );
  AND2X1 U16157 ( .IN1(n9987), .IN2(n12804), .Q(n15675) );
  OR2X1 U16158 ( .IN1(n15686), .IN2(n15687), .Q(n12804) );
  INVX0 U16159 ( .INP(n15688), .ZN(n15687) );
  OR2X1 U16160 ( .IN1(n15689), .IN2(n15690), .Q(n15688) );
  AND2X1 U16161 ( .IN1(n15690), .IN2(n15689), .Q(n15686) );
  AND2X1 U16162 ( .IN1(n15691), .IN2(n15692), .Q(n15689) );
  OR2X1 U16163 ( .IN1(WX2038), .IN2(n9507), .Q(n15692) );
  OR2X1 U16164 ( .IN1(WX1974), .IN2(n3781), .Q(n15691) );
  OR2X1 U16165 ( .IN1(n15693), .IN2(n15694), .Q(n15690) );
  AND2X1 U16166 ( .IN1(n9508), .IN2(WX2166), .Q(n15694) );
  AND2X1 U16167 ( .IN1(n9743), .IN2(WX2102), .Q(n15693) );
  OR2X1 U16168 ( .IN1(n15695), .IN2(n15696), .Q(WX1971) );
  OR2X1 U16169 ( .IN1(n15697), .IN2(n15698), .Q(n15696) );
  AND2X1 U16170 ( .IN1(n10033), .IN2(CRC_OUT_8_14), .Q(n15698) );
  AND2X1 U16171 ( .IN1(n266), .IN2(n10007), .Q(n15697) );
  INVX0 U16172 ( .INP(n15699), .ZN(n266) );
  OR2X1 U16173 ( .IN1(n10632), .IN2(n4017), .Q(n15699) );
  OR2X1 U16174 ( .IN1(n15700), .IN2(n15701), .Q(n15695) );
  AND2X1 U16175 ( .IN1(n10068), .IN2(n14826), .Q(n15701) );
  OR2X1 U16176 ( .IN1(n15702), .IN2(n15703), .Q(n14826) );
  INVX0 U16177 ( .INP(n15704), .ZN(n15703) );
  OR2X1 U16178 ( .IN1(n15705), .IN2(n15706), .Q(n15704) );
  AND2X1 U16179 ( .IN1(n15706), .IN2(n15705), .Q(n15702) );
  AND2X1 U16180 ( .IN1(n15707), .IN2(n15708), .Q(n15705) );
  OR2X1 U16181 ( .IN1(WX3329), .IN2(n9478), .Q(n15708) );
  OR2X1 U16182 ( .IN1(WX3265), .IN2(n3751), .Q(n15707) );
  OR2X1 U16183 ( .IN1(n15709), .IN2(n15710), .Q(n15706) );
  AND2X1 U16184 ( .IN1(n9479), .IN2(WX3457), .Q(n15710) );
  AND2X1 U16185 ( .IN1(n9716), .IN2(WX3393), .Q(n15709) );
  AND2X1 U16186 ( .IN1(n12812), .IN2(n9974), .Q(n15700) );
  AND2X1 U16187 ( .IN1(n15711), .IN2(n15712), .Q(n12812) );
  INVX0 U16188 ( .INP(n15713), .ZN(n15712) );
  AND2X1 U16189 ( .IN1(n15714), .IN2(n15715), .Q(n15713) );
  OR2X1 U16190 ( .IN1(n15715), .IN2(n15714), .Q(n15711) );
  OR2X1 U16191 ( .IN1(n15716), .IN2(n15717), .Q(n15714) );
  AND2X1 U16192 ( .IN1(n3783), .IN2(WX1972), .Q(n15717) );
  INVX0 U16193 ( .INP(n15718), .ZN(n15716) );
  OR2X1 U16194 ( .IN1(WX1972), .IN2(n3783), .Q(n15718) );
  AND2X1 U16195 ( .IN1(n15719), .IN2(n15720), .Q(n15715) );
  OR2X1 U16196 ( .IN1(WX2164), .IN2(test_so17), .Q(n15720) );
  OR2X1 U16197 ( .IN1(n9933), .IN2(n9742), .Q(n15719) );
  OR2X1 U16198 ( .IN1(n15721), .IN2(n15722), .Q(WX1969) );
  OR2X1 U16199 ( .IN1(n15723), .IN2(n15724), .Q(n15722) );
  AND2X1 U16200 ( .IN1(n10034), .IN2(CRC_OUT_8_15), .Q(n15724) );
  AND2X1 U16201 ( .IN1(n265), .IN2(n10007), .Q(n15723) );
  INVX0 U16202 ( .INP(n15725), .ZN(n265) );
  OR2X1 U16203 ( .IN1(n10632), .IN2(n4018), .Q(n15725) );
  OR2X1 U16204 ( .IN1(n15726), .IN2(n15727), .Q(n15721) );
  AND2X1 U16205 ( .IN1(n10068), .IN2(n14843), .Q(n15727) );
  OR2X1 U16206 ( .IN1(n15728), .IN2(n15729), .Q(n14843) );
  INVX0 U16207 ( .INP(n15730), .ZN(n15729) );
  OR2X1 U16208 ( .IN1(n15731), .IN2(n15732), .Q(n15730) );
  AND2X1 U16209 ( .IN1(n15732), .IN2(n15731), .Q(n15728) );
  AND2X1 U16210 ( .IN1(n15733), .IN2(n15734), .Q(n15731) );
  OR2X1 U16211 ( .IN1(WX3327), .IN2(n9480), .Q(n15734) );
  OR2X1 U16212 ( .IN1(WX3263), .IN2(n3753), .Q(n15733) );
  OR2X1 U16213 ( .IN1(n15735), .IN2(n15736), .Q(n15732) );
  AND2X1 U16214 ( .IN1(n9481), .IN2(WX3455), .Q(n15736) );
  AND2X1 U16215 ( .IN1(n9715), .IN2(WX3391), .Q(n15735) );
  AND2X1 U16216 ( .IN1(n9987), .IN2(n12820), .Q(n15726) );
  OR2X1 U16217 ( .IN1(n15737), .IN2(n15738), .Q(n12820) );
  INVX0 U16218 ( .INP(n15739), .ZN(n15738) );
  OR2X1 U16219 ( .IN1(n15740), .IN2(n15741), .Q(n15739) );
  AND2X1 U16220 ( .IN1(n15741), .IN2(n15740), .Q(n15737) );
  AND2X1 U16221 ( .IN1(n15742), .IN2(n15743), .Q(n15740) );
  OR2X1 U16222 ( .IN1(WX2034), .IN2(n9510), .Q(n15743) );
  OR2X1 U16223 ( .IN1(WX1970), .IN2(n3785), .Q(n15742) );
  OR2X1 U16224 ( .IN1(n15744), .IN2(n15745), .Q(n15741) );
  AND2X1 U16225 ( .IN1(n9511), .IN2(WX2162), .Q(n15745) );
  AND2X1 U16226 ( .IN1(n9741), .IN2(WX2098), .Q(n15744) );
  OR2X1 U16227 ( .IN1(n15746), .IN2(n15747), .Q(WX1967) );
  OR2X1 U16228 ( .IN1(n15748), .IN2(n15749), .Q(n15747) );
  AND2X1 U16229 ( .IN1(n10034), .IN2(CRC_OUT_8_16), .Q(n15749) );
  AND2X1 U16230 ( .IN1(n264), .IN2(n10007), .Q(n15748) );
  INVX0 U16231 ( .INP(n15750), .ZN(n264) );
  OR2X1 U16232 ( .IN1(n10632), .IN2(n4019), .Q(n15750) );
  OR2X1 U16233 ( .IN1(n15751), .IN2(n15752), .Q(n15746) );
  AND2X1 U16234 ( .IN1(n14861), .IN2(n10059), .Q(n15752) );
  AND2X1 U16235 ( .IN1(n15753), .IN2(n15754), .Q(n14861) );
  OR2X1 U16236 ( .IN1(n15755), .IN2(n15756), .Q(n15754) );
  INVX0 U16237 ( .INP(n15757), .ZN(n15755) );
  OR2X1 U16238 ( .IN1(n15758), .IN2(n15757), .Q(n15753) );
  OR2X1 U16239 ( .IN1(n15759), .IN2(n15760), .Q(n15757) );
  AND2X1 U16240 ( .IN1(n10525), .IN2(WX3453), .Q(n15760) );
  AND2X1 U16241 ( .IN1(n9527), .IN2(n10540), .Q(n15759) );
  INVX0 U16242 ( .INP(n15756), .ZN(n15758) );
  OR2X1 U16243 ( .IN1(n15761), .IN2(n15762), .Q(n15756) );
  AND2X1 U16244 ( .IN1(n9214), .IN2(n15763), .Q(n15762) );
  AND2X1 U16245 ( .IN1(n15764), .IN2(n15765), .Q(n15763) );
  OR2X1 U16246 ( .IN1(n9213), .IN2(n9894), .Q(n15765) );
  OR2X1 U16247 ( .IN1(test_so24), .IN2(WX3325), .Q(n15764) );
  AND2X1 U16248 ( .IN1(n15766), .IN2(WX3389), .Q(n15761) );
  OR2X1 U16249 ( .IN1(n15767), .IN2(n15768), .Q(n15766) );
  AND2X1 U16250 ( .IN1(n9213), .IN2(n9894), .Q(n15768) );
  AND2X1 U16251 ( .IN1(test_so24), .IN2(WX3325), .Q(n15767) );
  AND2X1 U16252 ( .IN1(n9987), .IN2(n12828), .Q(n15751) );
  OR2X1 U16253 ( .IN1(n15769), .IN2(n15770), .Q(n12828) );
  INVX0 U16254 ( .INP(n15771), .ZN(n15770) );
  OR2X1 U16255 ( .IN1(n15772), .IN2(n15773), .Q(n15771) );
  AND2X1 U16256 ( .IN1(n15773), .IN2(n15772), .Q(n15769) );
  INVX0 U16257 ( .INP(n15774), .ZN(n15772) );
  OR2X1 U16258 ( .IN1(n15775), .IN2(n15776), .Q(n15774) );
  AND2X1 U16259 ( .IN1(n10525), .IN2(n8653), .Q(n15776) );
  AND2X1 U16260 ( .IN1(n17957), .IN2(n10540), .Q(n15775) );
  OR2X1 U16261 ( .IN1(n15777), .IN2(n15778), .Q(n15773) );
  AND2X1 U16262 ( .IN1(n9530), .IN2(n15779), .Q(n15778) );
  AND2X1 U16263 ( .IN1(n15780), .IN2(n15781), .Q(n15779) );
  OR2X1 U16264 ( .IN1(n9241), .IN2(WX2096), .Q(n15781) );
  OR2X1 U16265 ( .IN1(n9242), .IN2(WX2032), .Q(n15780) );
  AND2X1 U16266 ( .IN1(n15782), .IN2(WX2160), .Q(n15777) );
  OR2X1 U16267 ( .IN1(n15783), .IN2(n15784), .Q(n15782) );
  AND2X1 U16268 ( .IN1(n9241), .IN2(WX2096), .Q(n15784) );
  AND2X1 U16269 ( .IN1(n9242), .IN2(WX2032), .Q(n15783) );
  OR2X1 U16270 ( .IN1(n15785), .IN2(n15786), .Q(WX1965) );
  OR2X1 U16271 ( .IN1(n15787), .IN2(n15788), .Q(n15786) );
  AND2X1 U16272 ( .IN1(n10034), .IN2(CRC_OUT_8_17), .Q(n15788) );
  AND2X1 U16273 ( .IN1(n263), .IN2(n10008), .Q(n15787) );
  INVX0 U16274 ( .INP(n15789), .ZN(n263) );
  OR2X1 U16275 ( .IN1(n10632), .IN2(n4020), .Q(n15789) );
  OR2X1 U16276 ( .IN1(n15790), .IN2(n15791), .Q(n15785) );
  AND2X1 U16277 ( .IN1(n10068), .IN2(n14885), .Q(n15791) );
  OR2X1 U16278 ( .IN1(n15792), .IN2(n15793), .Q(n14885) );
  INVX0 U16279 ( .INP(n15794), .ZN(n15793) );
  OR2X1 U16280 ( .IN1(n15795), .IN2(n15796), .Q(n15794) );
  AND2X1 U16281 ( .IN1(n15796), .IN2(n15795), .Q(n15792) );
  INVX0 U16282 ( .INP(n15797), .ZN(n15795) );
  OR2X1 U16283 ( .IN1(n15798), .IN2(n15799), .Q(n15797) );
  AND2X1 U16284 ( .IN1(n10525), .IN2(n8597), .Q(n15799) );
  AND2X1 U16285 ( .IN1(n17959), .IN2(n10540), .Q(n15798) );
  OR2X1 U16286 ( .IN1(n15800), .IN2(n15801), .Q(n15796) );
  AND2X1 U16287 ( .IN1(n9714), .IN2(n15802), .Q(n15801) );
  AND2X1 U16288 ( .IN1(n15803), .IN2(n15804), .Q(n15802) );
  OR2X1 U16289 ( .IN1(n9215), .IN2(WX3387), .Q(n15804) );
  OR2X1 U16290 ( .IN1(n9216), .IN2(WX3323), .Q(n15803) );
  AND2X1 U16291 ( .IN1(n15805), .IN2(WX3451), .Q(n15800) );
  OR2X1 U16292 ( .IN1(n15806), .IN2(n15807), .Q(n15805) );
  AND2X1 U16293 ( .IN1(n9215), .IN2(WX3387), .Q(n15807) );
  AND2X1 U16294 ( .IN1(n9216), .IN2(WX3323), .Q(n15806) );
  AND2X1 U16295 ( .IN1(n9987), .IN2(n12836), .Q(n15790) );
  OR2X1 U16296 ( .IN1(n15808), .IN2(n15809), .Q(n12836) );
  INVX0 U16297 ( .INP(n15810), .ZN(n15809) );
  OR2X1 U16298 ( .IN1(n15811), .IN2(n15812), .Q(n15810) );
  AND2X1 U16299 ( .IN1(n15812), .IN2(n15811), .Q(n15808) );
  INVX0 U16300 ( .INP(n15813), .ZN(n15811) );
  OR2X1 U16301 ( .IN1(n15814), .IN2(n15815), .Q(n15813) );
  AND2X1 U16302 ( .IN1(n10526), .IN2(n8654), .Q(n15815) );
  AND2X1 U16303 ( .IN1(n17958), .IN2(n10540), .Q(n15814) );
  OR2X1 U16304 ( .IN1(n15816), .IN2(n15817), .Q(n15812) );
  AND2X1 U16305 ( .IN1(n9740), .IN2(n15818), .Q(n15817) );
  AND2X1 U16306 ( .IN1(n15819), .IN2(n15820), .Q(n15818) );
  OR2X1 U16307 ( .IN1(n9243), .IN2(WX2094), .Q(n15820) );
  OR2X1 U16308 ( .IN1(n9244), .IN2(WX2030), .Q(n15819) );
  AND2X1 U16309 ( .IN1(n15821), .IN2(WX2158), .Q(n15816) );
  OR2X1 U16310 ( .IN1(n15822), .IN2(n15823), .Q(n15821) );
  AND2X1 U16311 ( .IN1(n9243), .IN2(WX2094), .Q(n15823) );
  AND2X1 U16312 ( .IN1(n9244), .IN2(WX2030), .Q(n15822) );
  OR2X1 U16313 ( .IN1(n15824), .IN2(n15825), .Q(WX1963) );
  OR2X1 U16314 ( .IN1(n15826), .IN2(n15827), .Q(n15825) );
  AND2X1 U16315 ( .IN1(n10034), .IN2(CRC_OUT_8_18), .Q(n15827) );
  AND2X1 U16316 ( .IN1(n262), .IN2(n10008), .Q(n15826) );
  INVX0 U16317 ( .INP(n15828), .ZN(n262) );
  OR2X1 U16318 ( .IN1(n10632), .IN2(n4021), .Q(n15828) );
  OR2X1 U16319 ( .IN1(n15829), .IN2(n15830), .Q(n15824) );
  AND2X1 U16320 ( .IN1(n10068), .IN2(n14909), .Q(n15830) );
  OR2X1 U16321 ( .IN1(n15831), .IN2(n15832), .Q(n14909) );
  INVX0 U16322 ( .INP(n15833), .ZN(n15832) );
  OR2X1 U16323 ( .IN1(n15834), .IN2(n15835), .Q(n15833) );
  AND2X1 U16324 ( .IN1(n15835), .IN2(n15834), .Q(n15831) );
  INVX0 U16325 ( .INP(n15836), .ZN(n15834) );
  OR2X1 U16326 ( .IN1(n15837), .IN2(n15838), .Q(n15836) );
  AND2X1 U16327 ( .IN1(n10526), .IN2(n8598), .Q(n15838) );
  AND2X1 U16328 ( .IN1(n17961), .IN2(n10540), .Q(n15837) );
  OR2X1 U16329 ( .IN1(n15839), .IN2(n15840), .Q(n15835) );
  AND2X1 U16330 ( .IN1(n9713), .IN2(n15841), .Q(n15840) );
  AND2X1 U16331 ( .IN1(n15842), .IN2(n15843), .Q(n15841) );
  OR2X1 U16332 ( .IN1(n9217), .IN2(WX3385), .Q(n15843) );
  OR2X1 U16333 ( .IN1(n9218), .IN2(WX3321), .Q(n15842) );
  AND2X1 U16334 ( .IN1(n15844), .IN2(WX3449), .Q(n15839) );
  OR2X1 U16335 ( .IN1(n15845), .IN2(n15846), .Q(n15844) );
  AND2X1 U16336 ( .IN1(n9217), .IN2(WX3385), .Q(n15846) );
  AND2X1 U16337 ( .IN1(n9218), .IN2(WX3321), .Q(n15845) );
  AND2X1 U16338 ( .IN1(n12844), .IN2(n9975), .Q(n15829) );
  AND2X1 U16339 ( .IN1(n15847), .IN2(n15848), .Q(n12844) );
  INVX0 U16340 ( .INP(n15849), .ZN(n15848) );
  AND2X1 U16341 ( .IN1(n15850), .IN2(n15851), .Q(n15849) );
  OR2X1 U16342 ( .IN1(n15851), .IN2(n15850), .Q(n15847) );
  OR2X1 U16343 ( .IN1(n15852), .IN2(n15853), .Q(n15850) );
  AND2X1 U16344 ( .IN1(n10526), .IN2(WX2092), .Q(n15853) );
  AND2X1 U16345 ( .IN1(n9245), .IN2(n10540), .Q(n15852) );
  AND2X1 U16346 ( .IN1(n15854), .IN2(n15855), .Q(n15851) );
  OR2X1 U16347 ( .IN1(n15856), .IN2(n9739), .Q(n15855) );
  INVX0 U16348 ( .INP(n15857), .ZN(n15856) );
  OR2X1 U16349 ( .IN1(WX2156), .IN2(n15857), .Q(n15854) );
  OR2X1 U16350 ( .IN1(n15858), .IN2(n15859), .Q(n15857) );
  AND2X1 U16351 ( .IN1(n17960), .IN2(n9962), .Q(n15859) );
  AND2X1 U16352 ( .IN1(test_so15), .IN2(n8655), .Q(n15858) );
  OR2X1 U16353 ( .IN1(n15860), .IN2(n15861), .Q(WX1961) );
  OR2X1 U16354 ( .IN1(n15862), .IN2(n15863), .Q(n15861) );
  AND2X1 U16355 ( .IN1(n10034), .IN2(CRC_OUT_8_19), .Q(n15863) );
  AND2X1 U16356 ( .IN1(n261), .IN2(n10008), .Q(n15862) );
  INVX0 U16357 ( .INP(n15864), .ZN(n261) );
  OR2X1 U16358 ( .IN1(n10632), .IN2(n4022), .Q(n15864) );
  OR2X1 U16359 ( .IN1(n15865), .IN2(n15866), .Q(n15860) );
  AND2X1 U16360 ( .IN1(n10068), .IN2(n14933), .Q(n15866) );
  OR2X1 U16361 ( .IN1(n15867), .IN2(n15868), .Q(n14933) );
  INVX0 U16362 ( .INP(n15869), .ZN(n15868) );
  OR2X1 U16363 ( .IN1(n15870), .IN2(n15871), .Q(n15869) );
  AND2X1 U16364 ( .IN1(n15871), .IN2(n15870), .Q(n15867) );
  INVX0 U16365 ( .INP(n15872), .ZN(n15870) );
  OR2X1 U16366 ( .IN1(n15873), .IN2(n15874), .Q(n15872) );
  AND2X1 U16367 ( .IN1(n10526), .IN2(n8599), .Q(n15874) );
  AND2X1 U16368 ( .IN1(n17963), .IN2(n10540), .Q(n15873) );
  OR2X1 U16369 ( .IN1(n15875), .IN2(n15876), .Q(n15871) );
  AND2X1 U16370 ( .IN1(n9712), .IN2(n15877), .Q(n15876) );
  AND2X1 U16371 ( .IN1(n15878), .IN2(n15879), .Q(n15877) );
  OR2X1 U16372 ( .IN1(n9219), .IN2(WX3383), .Q(n15879) );
  OR2X1 U16373 ( .IN1(n9220), .IN2(WX3319), .Q(n15878) );
  AND2X1 U16374 ( .IN1(n15880), .IN2(WX3447), .Q(n15875) );
  OR2X1 U16375 ( .IN1(n15881), .IN2(n15882), .Q(n15880) );
  AND2X1 U16376 ( .IN1(n9219), .IN2(WX3383), .Q(n15882) );
  AND2X1 U16377 ( .IN1(n9220), .IN2(WX3319), .Q(n15881) );
  AND2X1 U16378 ( .IN1(n9987), .IN2(n12852), .Q(n15865) );
  OR2X1 U16379 ( .IN1(n15883), .IN2(n15884), .Q(n12852) );
  INVX0 U16380 ( .INP(n15885), .ZN(n15884) );
  OR2X1 U16381 ( .IN1(n15886), .IN2(n15887), .Q(n15885) );
  AND2X1 U16382 ( .IN1(n15887), .IN2(n15886), .Q(n15883) );
  INVX0 U16383 ( .INP(n15888), .ZN(n15886) );
  OR2X1 U16384 ( .IN1(n15889), .IN2(n15890), .Q(n15888) );
  AND2X1 U16385 ( .IN1(n10526), .IN2(n8656), .Q(n15890) );
  AND2X1 U16386 ( .IN1(n17962), .IN2(n10540), .Q(n15889) );
  OR2X1 U16387 ( .IN1(n15891), .IN2(n15892), .Q(n15887) );
  AND2X1 U16388 ( .IN1(n9738), .IN2(n15893), .Q(n15892) );
  AND2X1 U16389 ( .IN1(n15894), .IN2(n15895), .Q(n15893) );
  OR2X1 U16390 ( .IN1(n9246), .IN2(WX2090), .Q(n15895) );
  OR2X1 U16391 ( .IN1(n9247), .IN2(WX2026), .Q(n15894) );
  AND2X1 U16392 ( .IN1(n15896), .IN2(WX2154), .Q(n15891) );
  OR2X1 U16393 ( .IN1(n15897), .IN2(n15898), .Q(n15896) );
  AND2X1 U16394 ( .IN1(n9246), .IN2(WX2090), .Q(n15898) );
  AND2X1 U16395 ( .IN1(n9247), .IN2(WX2026), .Q(n15897) );
  OR2X1 U16396 ( .IN1(n15899), .IN2(n15900), .Q(WX1959) );
  OR2X1 U16397 ( .IN1(n15901), .IN2(n15902), .Q(n15900) );
  AND2X1 U16398 ( .IN1(n10034), .IN2(CRC_OUT_8_20), .Q(n15902) );
  AND2X1 U16399 ( .IN1(n260), .IN2(n10008), .Q(n15901) );
  INVX0 U16400 ( .INP(n15903), .ZN(n260) );
  OR2X1 U16401 ( .IN1(n10632), .IN2(n4023), .Q(n15903) );
  OR2X1 U16402 ( .IN1(n15904), .IN2(n15905), .Q(n15899) );
  AND2X1 U16403 ( .IN1(n10068), .IN2(n14957), .Q(n15905) );
  OR2X1 U16404 ( .IN1(n15906), .IN2(n15907), .Q(n14957) );
  INVX0 U16405 ( .INP(n15908), .ZN(n15907) );
  OR2X1 U16406 ( .IN1(n15909), .IN2(n15910), .Q(n15908) );
  AND2X1 U16407 ( .IN1(n15910), .IN2(n15909), .Q(n15906) );
  INVX0 U16408 ( .INP(n15911), .ZN(n15909) );
  OR2X1 U16409 ( .IN1(n15912), .IN2(n15913), .Q(n15911) );
  AND2X1 U16410 ( .IN1(n10526), .IN2(n8600), .Q(n15913) );
  AND2X1 U16411 ( .IN1(n17965), .IN2(n10540), .Q(n15912) );
  OR2X1 U16412 ( .IN1(n15914), .IN2(n15915), .Q(n15910) );
  AND2X1 U16413 ( .IN1(n9711), .IN2(n15916), .Q(n15915) );
  AND2X1 U16414 ( .IN1(n15917), .IN2(n15918), .Q(n15916) );
  OR2X1 U16415 ( .IN1(n9221), .IN2(WX3381), .Q(n15918) );
  OR2X1 U16416 ( .IN1(n9222), .IN2(WX3317), .Q(n15917) );
  AND2X1 U16417 ( .IN1(n15919), .IN2(WX3445), .Q(n15914) );
  OR2X1 U16418 ( .IN1(n15920), .IN2(n15921), .Q(n15919) );
  AND2X1 U16419 ( .IN1(n9221), .IN2(WX3381), .Q(n15921) );
  AND2X1 U16420 ( .IN1(n9222), .IN2(WX3317), .Q(n15920) );
  AND2X1 U16421 ( .IN1(n9987), .IN2(n12860), .Q(n15904) );
  OR2X1 U16422 ( .IN1(n15922), .IN2(n15923), .Q(n12860) );
  INVX0 U16423 ( .INP(n15924), .ZN(n15923) );
  OR2X1 U16424 ( .IN1(n15925), .IN2(n15926), .Q(n15924) );
  AND2X1 U16425 ( .IN1(n15926), .IN2(n15925), .Q(n15922) );
  INVX0 U16426 ( .INP(n15927), .ZN(n15925) );
  OR2X1 U16427 ( .IN1(n15928), .IN2(n15929), .Q(n15927) );
  AND2X1 U16428 ( .IN1(n10526), .IN2(n8657), .Q(n15929) );
  AND2X1 U16429 ( .IN1(n17964), .IN2(n10540), .Q(n15928) );
  OR2X1 U16430 ( .IN1(n15930), .IN2(n15931), .Q(n15926) );
  AND2X1 U16431 ( .IN1(n9737), .IN2(n15932), .Q(n15931) );
  AND2X1 U16432 ( .IN1(n15933), .IN2(n15934), .Q(n15932) );
  OR2X1 U16433 ( .IN1(n9248), .IN2(WX2088), .Q(n15934) );
  OR2X1 U16434 ( .IN1(n9249), .IN2(WX2024), .Q(n15933) );
  AND2X1 U16435 ( .IN1(n15935), .IN2(WX2152), .Q(n15930) );
  OR2X1 U16436 ( .IN1(n15936), .IN2(n15937), .Q(n15935) );
  AND2X1 U16437 ( .IN1(n9248), .IN2(WX2088), .Q(n15937) );
  AND2X1 U16438 ( .IN1(n9249), .IN2(WX2024), .Q(n15936) );
  OR2X1 U16439 ( .IN1(n15938), .IN2(n15939), .Q(WX1957) );
  OR2X1 U16440 ( .IN1(n15940), .IN2(n15941), .Q(n15939) );
  AND2X1 U16441 ( .IN1(n10034), .IN2(CRC_OUT_8_21), .Q(n15941) );
  AND2X1 U16442 ( .IN1(n259), .IN2(n10008), .Q(n15940) );
  INVX0 U16443 ( .INP(n15942), .ZN(n259) );
  OR2X1 U16444 ( .IN1(n10632), .IN2(n4024), .Q(n15942) );
  OR2X1 U16445 ( .IN1(n15943), .IN2(n15944), .Q(n15938) );
  AND2X1 U16446 ( .IN1(n10068), .IN2(n14981), .Q(n15944) );
  OR2X1 U16447 ( .IN1(n15945), .IN2(n15946), .Q(n14981) );
  INVX0 U16448 ( .INP(n15947), .ZN(n15946) );
  OR2X1 U16449 ( .IN1(n15948), .IN2(n15949), .Q(n15947) );
  AND2X1 U16450 ( .IN1(n15949), .IN2(n15948), .Q(n15945) );
  INVX0 U16451 ( .INP(n15950), .ZN(n15948) );
  OR2X1 U16452 ( .IN1(n15951), .IN2(n15952), .Q(n15950) );
  AND2X1 U16453 ( .IN1(n10526), .IN2(n8601), .Q(n15952) );
  AND2X1 U16454 ( .IN1(n17967), .IN2(n10540), .Q(n15951) );
  OR2X1 U16455 ( .IN1(n15953), .IN2(n15954), .Q(n15949) );
  AND2X1 U16456 ( .IN1(n9710), .IN2(n15955), .Q(n15954) );
  AND2X1 U16457 ( .IN1(n15956), .IN2(n15957), .Q(n15955) );
  OR2X1 U16458 ( .IN1(n9223), .IN2(WX3379), .Q(n15957) );
  OR2X1 U16459 ( .IN1(n9224), .IN2(WX3315), .Q(n15956) );
  AND2X1 U16460 ( .IN1(n15958), .IN2(WX3443), .Q(n15953) );
  OR2X1 U16461 ( .IN1(n15959), .IN2(n15960), .Q(n15958) );
  AND2X1 U16462 ( .IN1(n9223), .IN2(WX3379), .Q(n15960) );
  AND2X1 U16463 ( .IN1(n9224), .IN2(WX3315), .Q(n15959) );
  AND2X1 U16464 ( .IN1(n9987), .IN2(n12868), .Q(n15943) );
  OR2X1 U16465 ( .IN1(n15961), .IN2(n15962), .Q(n12868) );
  INVX0 U16466 ( .INP(n15963), .ZN(n15962) );
  OR2X1 U16467 ( .IN1(n15964), .IN2(n15965), .Q(n15963) );
  AND2X1 U16468 ( .IN1(n15965), .IN2(n15964), .Q(n15961) );
  INVX0 U16469 ( .INP(n15966), .ZN(n15964) );
  OR2X1 U16470 ( .IN1(n15967), .IN2(n15968), .Q(n15966) );
  AND2X1 U16471 ( .IN1(n10526), .IN2(n8658), .Q(n15968) );
  AND2X1 U16472 ( .IN1(n17966), .IN2(n10540), .Q(n15967) );
  OR2X1 U16473 ( .IN1(n15969), .IN2(n15970), .Q(n15965) );
  AND2X1 U16474 ( .IN1(n9736), .IN2(n15971), .Q(n15970) );
  AND2X1 U16475 ( .IN1(n15972), .IN2(n15973), .Q(n15971) );
  OR2X1 U16476 ( .IN1(n9250), .IN2(WX2086), .Q(n15973) );
  OR2X1 U16477 ( .IN1(n9251), .IN2(WX2022), .Q(n15972) );
  AND2X1 U16478 ( .IN1(n15974), .IN2(WX2150), .Q(n15969) );
  OR2X1 U16479 ( .IN1(n15975), .IN2(n15976), .Q(n15974) );
  AND2X1 U16480 ( .IN1(n9250), .IN2(WX2086), .Q(n15976) );
  AND2X1 U16481 ( .IN1(n9251), .IN2(WX2022), .Q(n15975) );
  OR2X1 U16482 ( .IN1(n15977), .IN2(n15978), .Q(WX1955) );
  OR2X1 U16483 ( .IN1(n15979), .IN2(n15980), .Q(n15978) );
  AND2X1 U16484 ( .IN1(n10034), .IN2(CRC_OUT_8_22), .Q(n15980) );
  AND2X1 U16485 ( .IN1(n258), .IN2(n10008), .Q(n15979) );
  INVX0 U16486 ( .INP(n15981), .ZN(n258) );
  OR2X1 U16487 ( .IN1(n10632), .IN2(n4025), .Q(n15981) );
  OR2X1 U16488 ( .IN1(n15982), .IN2(n15983), .Q(n15977) );
  AND2X1 U16489 ( .IN1(n10068), .IN2(n15005), .Q(n15983) );
  OR2X1 U16490 ( .IN1(n15984), .IN2(n15985), .Q(n15005) );
  INVX0 U16491 ( .INP(n15986), .ZN(n15985) );
  OR2X1 U16492 ( .IN1(n15987), .IN2(n15988), .Q(n15986) );
  AND2X1 U16493 ( .IN1(n15988), .IN2(n15987), .Q(n15984) );
  INVX0 U16494 ( .INP(n15989), .ZN(n15987) );
  OR2X1 U16495 ( .IN1(n15990), .IN2(n15991), .Q(n15989) );
  AND2X1 U16496 ( .IN1(n10526), .IN2(n8602), .Q(n15991) );
  AND2X1 U16497 ( .IN1(n17968), .IN2(n10540), .Q(n15990) );
  OR2X1 U16498 ( .IN1(n15992), .IN2(n15993), .Q(n15988) );
  AND2X1 U16499 ( .IN1(n9709), .IN2(n15994), .Q(n15993) );
  AND2X1 U16500 ( .IN1(n15995), .IN2(n15996), .Q(n15994) );
  OR2X1 U16501 ( .IN1(n9225), .IN2(WX3377), .Q(n15996) );
  OR2X1 U16502 ( .IN1(n9226), .IN2(WX3313), .Q(n15995) );
  AND2X1 U16503 ( .IN1(n15997), .IN2(WX3441), .Q(n15992) );
  OR2X1 U16504 ( .IN1(n15998), .IN2(n15999), .Q(n15997) );
  AND2X1 U16505 ( .IN1(n9225), .IN2(WX3377), .Q(n15999) );
  AND2X1 U16506 ( .IN1(n9226), .IN2(WX3313), .Q(n15998) );
  AND2X1 U16507 ( .IN1(n12876), .IN2(n9974), .Q(n15982) );
  AND2X1 U16508 ( .IN1(n16000), .IN2(n16001), .Q(n12876) );
  OR2X1 U16509 ( .IN1(n16002), .IN2(n16003), .Q(n16001) );
  INVX0 U16510 ( .INP(n16004), .ZN(n16002) );
  OR2X1 U16511 ( .IN1(n16005), .IN2(n16004), .Q(n16000) );
  OR2X1 U16512 ( .IN1(n16006), .IN2(n16007), .Q(n16004) );
  AND2X1 U16513 ( .IN1(n10527), .IN2(WX2148), .Q(n16007) );
  AND2X1 U16514 ( .IN1(n9735), .IN2(n10540), .Q(n16006) );
  INVX0 U16515 ( .INP(n16003), .ZN(n16005) );
  OR2X1 U16516 ( .IN1(n16008), .IN2(n16009), .Q(n16003) );
  AND2X1 U16517 ( .IN1(n9253), .IN2(n16010), .Q(n16009) );
  AND2X1 U16518 ( .IN1(n16011), .IN2(n16012), .Q(n16010) );
  OR2X1 U16519 ( .IN1(n9252), .IN2(n9895), .Q(n16012) );
  OR2X1 U16520 ( .IN1(test_so13), .IN2(WX2020), .Q(n16011) );
  AND2X1 U16521 ( .IN1(n16013), .IN2(WX2084), .Q(n16008) );
  OR2X1 U16522 ( .IN1(n16014), .IN2(n16015), .Q(n16013) );
  AND2X1 U16523 ( .IN1(n9252), .IN2(n9895), .Q(n16015) );
  AND2X1 U16524 ( .IN1(test_so13), .IN2(WX2020), .Q(n16014) );
  OR2X1 U16525 ( .IN1(n16016), .IN2(n16017), .Q(WX1953) );
  OR2X1 U16526 ( .IN1(n16018), .IN2(n16019), .Q(n16017) );
  AND2X1 U16527 ( .IN1(n10034), .IN2(CRC_OUT_8_23), .Q(n16019) );
  AND2X1 U16528 ( .IN1(n257), .IN2(n10008), .Q(n16018) );
  INVX0 U16529 ( .INP(n16020), .ZN(n257) );
  OR2X1 U16530 ( .IN1(n10632), .IN2(n4026), .Q(n16020) );
  OR2X1 U16531 ( .IN1(n16021), .IN2(n16022), .Q(n16016) );
  AND2X1 U16532 ( .IN1(n15029), .IN2(n10059), .Q(n16022) );
  AND2X1 U16533 ( .IN1(n16023), .IN2(n16024), .Q(n15029) );
  INVX0 U16534 ( .INP(n16025), .ZN(n16024) );
  AND2X1 U16535 ( .IN1(n16026), .IN2(n16027), .Q(n16025) );
  OR2X1 U16536 ( .IN1(n16027), .IN2(n16026), .Q(n16023) );
  OR2X1 U16537 ( .IN1(n16028), .IN2(n16029), .Q(n16026) );
  AND2X1 U16538 ( .IN1(n10527), .IN2(WX3311), .Q(n16029) );
  AND2X1 U16539 ( .IN1(n9227), .IN2(n10540), .Q(n16028) );
  AND2X1 U16540 ( .IN1(n16030), .IN2(n16031), .Q(n16027) );
  INVX0 U16541 ( .INP(n16032), .ZN(n16031) );
  AND2X1 U16542 ( .IN1(n16033), .IN2(WX3375), .Q(n16032) );
  OR2X1 U16543 ( .IN1(WX3375), .IN2(n16033), .Q(n16030) );
  OR2X1 U16544 ( .IN1(n16034), .IN2(n16035), .Q(n16033) );
  AND2X1 U16545 ( .IN1(n17970), .IN2(n9911), .Q(n16035) );
  AND2X1 U16546 ( .IN1(test_so29), .IN2(n8603), .Q(n16034) );
  AND2X1 U16547 ( .IN1(n9987), .IN2(n12884), .Q(n16021) );
  OR2X1 U16548 ( .IN1(n16036), .IN2(n16037), .Q(n12884) );
  INVX0 U16549 ( .INP(n16038), .ZN(n16037) );
  OR2X1 U16550 ( .IN1(n16039), .IN2(n16040), .Q(n16038) );
  AND2X1 U16551 ( .IN1(n16040), .IN2(n16039), .Q(n16036) );
  INVX0 U16552 ( .INP(n16041), .ZN(n16039) );
  OR2X1 U16553 ( .IN1(n16042), .IN2(n16043), .Q(n16041) );
  AND2X1 U16554 ( .IN1(n10527), .IN2(n8661), .Q(n16043) );
  AND2X1 U16555 ( .IN1(n17969), .IN2(n10540), .Q(n16042) );
  OR2X1 U16556 ( .IN1(n16044), .IN2(n16045), .Q(n16040) );
  AND2X1 U16557 ( .IN1(n9734), .IN2(n16046), .Q(n16045) );
  AND2X1 U16558 ( .IN1(n16047), .IN2(n16048), .Q(n16046) );
  OR2X1 U16559 ( .IN1(n9254), .IN2(WX2082), .Q(n16048) );
  OR2X1 U16560 ( .IN1(n9255), .IN2(WX2018), .Q(n16047) );
  AND2X1 U16561 ( .IN1(n16049), .IN2(WX2146), .Q(n16044) );
  OR2X1 U16562 ( .IN1(n16050), .IN2(n16051), .Q(n16049) );
  AND2X1 U16563 ( .IN1(n9254), .IN2(WX2082), .Q(n16051) );
  AND2X1 U16564 ( .IN1(n9255), .IN2(WX2018), .Q(n16050) );
  OR2X1 U16565 ( .IN1(n16052), .IN2(n16053), .Q(WX1951) );
  OR2X1 U16566 ( .IN1(n16054), .IN2(n16055), .Q(n16053) );
  AND2X1 U16567 ( .IN1(n10034), .IN2(CRC_OUT_8_24), .Q(n16055) );
  AND2X1 U16568 ( .IN1(n256), .IN2(n10008), .Q(n16054) );
  INVX0 U16569 ( .INP(n16056), .ZN(n256) );
  OR2X1 U16570 ( .IN1(n10632), .IN2(n4027), .Q(n16056) );
  OR2X1 U16571 ( .IN1(n16057), .IN2(n16058), .Q(n16052) );
  AND2X1 U16572 ( .IN1(n10068), .IN2(n15053), .Q(n16058) );
  OR2X1 U16573 ( .IN1(n16059), .IN2(n16060), .Q(n15053) );
  INVX0 U16574 ( .INP(n16061), .ZN(n16060) );
  OR2X1 U16575 ( .IN1(n16062), .IN2(n16063), .Q(n16061) );
  AND2X1 U16576 ( .IN1(n16063), .IN2(n16062), .Q(n16059) );
  INVX0 U16577 ( .INP(n16064), .ZN(n16062) );
  OR2X1 U16578 ( .IN1(n16065), .IN2(n16066), .Q(n16064) );
  AND2X1 U16579 ( .IN1(n10527), .IN2(n8604), .Q(n16066) );
  AND2X1 U16580 ( .IN1(n17972), .IN2(n10540), .Q(n16065) );
  OR2X1 U16581 ( .IN1(n16067), .IN2(n16068), .Q(n16063) );
  AND2X1 U16582 ( .IN1(n9708), .IN2(n16069), .Q(n16068) );
  AND2X1 U16583 ( .IN1(n16070), .IN2(n16071), .Q(n16069) );
  OR2X1 U16584 ( .IN1(n9229), .IN2(WX3373), .Q(n16071) );
  OR2X1 U16585 ( .IN1(n9230), .IN2(WX3309), .Q(n16070) );
  AND2X1 U16586 ( .IN1(n16072), .IN2(WX3437), .Q(n16067) );
  OR2X1 U16587 ( .IN1(n16073), .IN2(n16074), .Q(n16072) );
  AND2X1 U16588 ( .IN1(n9229), .IN2(WX3373), .Q(n16074) );
  AND2X1 U16589 ( .IN1(n9230), .IN2(WX3309), .Q(n16073) );
  AND2X1 U16590 ( .IN1(n9987), .IN2(n12892), .Q(n16057) );
  OR2X1 U16591 ( .IN1(n16075), .IN2(n16076), .Q(n12892) );
  INVX0 U16592 ( .INP(n16077), .ZN(n16076) );
  OR2X1 U16593 ( .IN1(n16078), .IN2(n16079), .Q(n16077) );
  AND2X1 U16594 ( .IN1(n16079), .IN2(n16078), .Q(n16075) );
  INVX0 U16595 ( .INP(n16080), .ZN(n16078) );
  OR2X1 U16596 ( .IN1(n16081), .IN2(n16082), .Q(n16080) );
  AND2X1 U16597 ( .IN1(n10527), .IN2(n8662), .Q(n16082) );
  AND2X1 U16598 ( .IN1(n17971), .IN2(n10540), .Q(n16081) );
  OR2X1 U16599 ( .IN1(n16083), .IN2(n16084), .Q(n16079) );
  AND2X1 U16600 ( .IN1(n9733), .IN2(n16085), .Q(n16084) );
  AND2X1 U16601 ( .IN1(n16086), .IN2(n16087), .Q(n16085) );
  OR2X1 U16602 ( .IN1(n9256), .IN2(WX2080), .Q(n16087) );
  OR2X1 U16603 ( .IN1(n9257), .IN2(WX2016), .Q(n16086) );
  AND2X1 U16604 ( .IN1(n16088), .IN2(WX2144), .Q(n16083) );
  OR2X1 U16605 ( .IN1(n16089), .IN2(n16090), .Q(n16088) );
  AND2X1 U16606 ( .IN1(n9256), .IN2(WX2080), .Q(n16090) );
  AND2X1 U16607 ( .IN1(n9257), .IN2(WX2016), .Q(n16089) );
  OR2X1 U16608 ( .IN1(n16091), .IN2(n16092), .Q(WX1949) );
  OR2X1 U16609 ( .IN1(n16093), .IN2(n16094), .Q(n16092) );
  AND2X1 U16610 ( .IN1(test_so21), .IN2(n10027), .Q(n16094) );
  AND2X1 U16611 ( .IN1(n255), .IN2(n10008), .Q(n16093) );
  INVX0 U16612 ( .INP(n16095), .ZN(n255) );
  OR2X1 U16613 ( .IN1(n10632), .IN2(n4028), .Q(n16095) );
  OR2X1 U16614 ( .IN1(n16096), .IN2(n16097), .Q(n16091) );
  AND2X1 U16615 ( .IN1(n10068), .IN2(n15077), .Q(n16097) );
  OR2X1 U16616 ( .IN1(n16098), .IN2(n16099), .Q(n15077) );
  INVX0 U16617 ( .INP(n16100), .ZN(n16099) );
  OR2X1 U16618 ( .IN1(n16101), .IN2(n16102), .Q(n16100) );
  AND2X1 U16619 ( .IN1(n16102), .IN2(n16101), .Q(n16098) );
  INVX0 U16620 ( .INP(n16103), .ZN(n16101) );
  OR2X1 U16621 ( .IN1(n16104), .IN2(n16105), .Q(n16103) );
  AND2X1 U16622 ( .IN1(n10527), .IN2(n8605), .Q(n16105) );
  AND2X1 U16623 ( .IN1(n17974), .IN2(n10539), .Q(n16104) );
  OR2X1 U16624 ( .IN1(n16106), .IN2(n16107), .Q(n16102) );
  AND2X1 U16625 ( .IN1(n9707), .IN2(n16108), .Q(n16107) );
  AND2X1 U16626 ( .IN1(n16109), .IN2(n16110), .Q(n16108) );
  OR2X1 U16627 ( .IN1(n9231), .IN2(WX3371), .Q(n16110) );
  OR2X1 U16628 ( .IN1(n9232), .IN2(WX3307), .Q(n16109) );
  AND2X1 U16629 ( .IN1(n16111), .IN2(WX3435), .Q(n16106) );
  OR2X1 U16630 ( .IN1(n16112), .IN2(n16113), .Q(n16111) );
  AND2X1 U16631 ( .IN1(n9231), .IN2(WX3371), .Q(n16113) );
  AND2X1 U16632 ( .IN1(n9232), .IN2(WX3307), .Q(n16112) );
  AND2X1 U16633 ( .IN1(n9987), .IN2(n12900), .Q(n16096) );
  OR2X1 U16634 ( .IN1(n16114), .IN2(n16115), .Q(n12900) );
  INVX0 U16635 ( .INP(n16116), .ZN(n16115) );
  OR2X1 U16636 ( .IN1(n16117), .IN2(n16118), .Q(n16116) );
  AND2X1 U16637 ( .IN1(n16118), .IN2(n16117), .Q(n16114) );
  INVX0 U16638 ( .INP(n16119), .ZN(n16117) );
  OR2X1 U16639 ( .IN1(n16120), .IN2(n16121), .Q(n16119) );
  AND2X1 U16640 ( .IN1(n10527), .IN2(n8663), .Q(n16121) );
  AND2X1 U16641 ( .IN1(n17973), .IN2(n10539), .Q(n16120) );
  OR2X1 U16642 ( .IN1(n16122), .IN2(n16123), .Q(n16118) );
  AND2X1 U16643 ( .IN1(n9732), .IN2(n16124), .Q(n16123) );
  AND2X1 U16644 ( .IN1(n16125), .IN2(n16126), .Q(n16124) );
  OR2X1 U16645 ( .IN1(n9258), .IN2(WX2078), .Q(n16126) );
  OR2X1 U16646 ( .IN1(n9259), .IN2(WX2014), .Q(n16125) );
  AND2X1 U16647 ( .IN1(n16127), .IN2(WX2142), .Q(n16122) );
  OR2X1 U16648 ( .IN1(n16128), .IN2(n16129), .Q(n16127) );
  AND2X1 U16649 ( .IN1(n9258), .IN2(WX2078), .Q(n16129) );
  AND2X1 U16650 ( .IN1(n9259), .IN2(WX2014), .Q(n16128) );
  OR2X1 U16651 ( .IN1(n16130), .IN2(n16131), .Q(WX1947) );
  OR2X1 U16652 ( .IN1(n16132), .IN2(n16133), .Q(n16131) );
  AND2X1 U16653 ( .IN1(n10034), .IN2(CRC_OUT_8_26), .Q(n16133) );
  AND2X1 U16654 ( .IN1(n254), .IN2(n10008), .Q(n16132) );
  INVX0 U16655 ( .INP(n16134), .ZN(n254) );
  OR2X1 U16656 ( .IN1(n10631), .IN2(n4029), .Q(n16134) );
  OR2X1 U16657 ( .IN1(n16135), .IN2(n16136), .Q(n16130) );
  AND2X1 U16658 ( .IN1(n15101), .IN2(n10059), .Q(n16136) );
  AND2X1 U16659 ( .IN1(n16137), .IN2(n16138), .Q(n15101) );
  INVX0 U16660 ( .INP(n16139), .ZN(n16138) );
  AND2X1 U16661 ( .IN1(n16140), .IN2(n16141), .Q(n16139) );
  OR2X1 U16662 ( .IN1(n16141), .IN2(n16140), .Q(n16137) );
  OR2X1 U16663 ( .IN1(n16142), .IN2(n16143), .Q(n16140) );
  AND2X1 U16664 ( .IN1(n10527), .IN2(WX3305), .Q(n16143) );
  AND2X1 U16665 ( .IN1(n9233), .IN2(n10539), .Q(n16142) );
  AND2X1 U16666 ( .IN1(n16144), .IN2(n16145), .Q(n16141) );
  OR2X1 U16667 ( .IN1(n16146), .IN2(n9706), .Q(n16145) );
  INVX0 U16668 ( .INP(n16147), .ZN(n16146) );
  OR2X1 U16669 ( .IN1(WX3433), .IN2(n16147), .Q(n16144) );
  OR2X1 U16670 ( .IN1(n16148), .IN2(n16149), .Q(n16147) );
  AND2X1 U16671 ( .IN1(n17976), .IN2(n9963), .Q(n16149) );
  AND2X1 U16672 ( .IN1(test_so27), .IN2(n8606), .Q(n16148) );
  AND2X1 U16673 ( .IN1(n9986), .IN2(n12908), .Q(n16135) );
  OR2X1 U16674 ( .IN1(n16150), .IN2(n16151), .Q(n12908) );
  INVX0 U16675 ( .INP(n16152), .ZN(n16151) );
  OR2X1 U16676 ( .IN1(n16153), .IN2(n16154), .Q(n16152) );
  AND2X1 U16677 ( .IN1(n16154), .IN2(n16153), .Q(n16150) );
  INVX0 U16678 ( .INP(n16155), .ZN(n16153) );
  OR2X1 U16679 ( .IN1(n16156), .IN2(n16157), .Q(n16155) );
  AND2X1 U16680 ( .IN1(n10527), .IN2(n8664), .Q(n16157) );
  AND2X1 U16681 ( .IN1(n17975), .IN2(n10539), .Q(n16156) );
  OR2X1 U16682 ( .IN1(n16158), .IN2(n16159), .Q(n16154) );
  AND2X1 U16683 ( .IN1(n9731), .IN2(n16160), .Q(n16159) );
  AND2X1 U16684 ( .IN1(n16161), .IN2(n16162), .Q(n16160) );
  OR2X1 U16685 ( .IN1(n9260), .IN2(WX2076), .Q(n16162) );
  OR2X1 U16686 ( .IN1(n9261), .IN2(WX2012), .Q(n16161) );
  AND2X1 U16687 ( .IN1(n16163), .IN2(WX2140), .Q(n16158) );
  OR2X1 U16688 ( .IN1(n16164), .IN2(n16165), .Q(n16163) );
  AND2X1 U16689 ( .IN1(n9260), .IN2(WX2076), .Q(n16165) );
  AND2X1 U16690 ( .IN1(n9261), .IN2(WX2012), .Q(n16164) );
  OR2X1 U16691 ( .IN1(n16166), .IN2(n16167), .Q(WX1945) );
  OR2X1 U16692 ( .IN1(n16168), .IN2(n16169), .Q(n16167) );
  AND2X1 U16693 ( .IN1(n10034), .IN2(CRC_OUT_8_27), .Q(n16169) );
  AND2X1 U16694 ( .IN1(n253), .IN2(n10008), .Q(n16168) );
  INVX0 U16695 ( .INP(n16170), .ZN(n253) );
  OR2X1 U16696 ( .IN1(n10631), .IN2(n4030), .Q(n16170) );
  OR2X1 U16697 ( .IN1(n16171), .IN2(n16172), .Q(n16166) );
  AND2X1 U16698 ( .IN1(n10064), .IN2(n15125), .Q(n16172) );
  OR2X1 U16699 ( .IN1(n16173), .IN2(n16174), .Q(n15125) );
  INVX0 U16700 ( .INP(n16175), .ZN(n16174) );
  OR2X1 U16701 ( .IN1(n16176), .IN2(n16177), .Q(n16175) );
  AND2X1 U16702 ( .IN1(n16177), .IN2(n16176), .Q(n16173) );
  INVX0 U16703 ( .INP(n16178), .ZN(n16176) );
  OR2X1 U16704 ( .IN1(n16179), .IN2(n16180), .Q(n16178) );
  AND2X1 U16705 ( .IN1(n10527), .IN2(n8607), .Q(n16180) );
  AND2X1 U16706 ( .IN1(n17978), .IN2(n10539), .Q(n16179) );
  OR2X1 U16707 ( .IN1(n16181), .IN2(n16182), .Q(n16177) );
  AND2X1 U16708 ( .IN1(n9705), .IN2(n16183), .Q(n16182) );
  AND2X1 U16709 ( .IN1(n16184), .IN2(n16185), .Q(n16183) );
  OR2X1 U16710 ( .IN1(n9234), .IN2(WX3367), .Q(n16185) );
  OR2X1 U16711 ( .IN1(n9235), .IN2(WX3303), .Q(n16184) );
  AND2X1 U16712 ( .IN1(n16186), .IN2(WX3431), .Q(n16181) );
  OR2X1 U16713 ( .IN1(n16187), .IN2(n16188), .Q(n16186) );
  AND2X1 U16714 ( .IN1(n9234), .IN2(WX3367), .Q(n16188) );
  AND2X1 U16715 ( .IN1(n9235), .IN2(WX3303), .Q(n16187) );
  AND2X1 U16716 ( .IN1(n9986), .IN2(n12916), .Q(n16171) );
  OR2X1 U16717 ( .IN1(n16189), .IN2(n16190), .Q(n12916) );
  INVX0 U16718 ( .INP(n16191), .ZN(n16190) );
  OR2X1 U16719 ( .IN1(n16192), .IN2(n16193), .Q(n16191) );
  AND2X1 U16720 ( .IN1(n16193), .IN2(n16192), .Q(n16189) );
  INVX0 U16721 ( .INP(n16194), .ZN(n16192) );
  OR2X1 U16722 ( .IN1(n16195), .IN2(n16196), .Q(n16194) );
  AND2X1 U16723 ( .IN1(n10528), .IN2(n8665), .Q(n16196) );
  AND2X1 U16724 ( .IN1(n17977), .IN2(n10539), .Q(n16195) );
  OR2X1 U16725 ( .IN1(n16197), .IN2(n16198), .Q(n16193) );
  AND2X1 U16726 ( .IN1(n9730), .IN2(n16199), .Q(n16198) );
  AND2X1 U16727 ( .IN1(n16200), .IN2(n16201), .Q(n16199) );
  OR2X1 U16728 ( .IN1(n9262), .IN2(WX2074), .Q(n16201) );
  OR2X1 U16729 ( .IN1(n9263), .IN2(WX2010), .Q(n16200) );
  AND2X1 U16730 ( .IN1(n16202), .IN2(WX2138), .Q(n16197) );
  OR2X1 U16731 ( .IN1(n16203), .IN2(n16204), .Q(n16202) );
  AND2X1 U16732 ( .IN1(n9262), .IN2(WX2074), .Q(n16204) );
  AND2X1 U16733 ( .IN1(n9263), .IN2(WX2010), .Q(n16203) );
  OR2X1 U16734 ( .IN1(n16205), .IN2(n16206), .Q(WX1943) );
  OR2X1 U16735 ( .IN1(n16207), .IN2(n16208), .Q(n16206) );
  AND2X1 U16736 ( .IN1(n10034), .IN2(CRC_OUT_8_28), .Q(n16208) );
  AND2X1 U16737 ( .IN1(n252), .IN2(n10008), .Q(n16207) );
  INVX0 U16738 ( .INP(n16209), .ZN(n252) );
  OR2X1 U16739 ( .IN1(n10631), .IN2(n4031), .Q(n16209) );
  OR2X1 U16740 ( .IN1(n16210), .IN2(n16211), .Q(n16205) );
  AND2X1 U16741 ( .IN1(n10069), .IN2(n15149), .Q(n16211) );
  OR2X1 U16742 ( .IN1(n16212), .IN2(n16213), .Q(n15149) );
  INVX0 U16743 ( .INP(n16214), .ZN(n16213) );
  OR2X1 U16744 ( .IN1(n16215), .IN2(n16216), .Q(n16214) );
  AND2X1 U16745 ( .IN1(n16216), .IN2(n16215), .Q(n16212) );
  INVX0 U16746 ( .INP(n16217), .ZN(n16215) );
  OR2X1 U16747 ( .IN1(n16218), .IN2(n16219), .Q(n16217) );
  AND2X1 U16748 ( .IN1(n10528), .IN2(n8608), .Q(n16219) );
  AND2X1 U16749 ( .IN1(n17980), .IN2(n10539), .Q(n16218) );
  OR2X1 U16750 ( .IN1(n16220), .IN2(n16221), .Q(n16216) );
  AND2X1 U16751 ( .IN1(n9704), .IN2(n16222), .Q(n16221) );
  AND2X1 U16752 ( .IN1(n16223), .IN2(n16224), .Q(n16222) );
  OR2X1 U16753 ( .IN1(n9236), .IN2(WX3365), .Q(n16224) );
  OR2X1 U16754 ( .IN1(n9237), .IN2(WX3301), .Q(n16223) );
  AND2X1 U16755 ( .IN1(n16225), .IN2(WX3429), .Q(n16220) );
  OR2X1 U16756 ( .IN1(n16226), .IN2(n16227), .Q(n16225) );
  AND2X1 U16757 ( .IN1(n9236), .IN2(WX3365), .Q(n16227) );
  AND2X1 U16758 ( .IN1(n9237), .IN2(WX3301), .Q(n16226) );
  AND2X1 U16759 ( .IN1(n12924), .IN2(n9974), .Q(n16210) );
  AND2X1 U16760 ( .IN1(n16228), .IN2(n16229), .Q(n12924) );
  INVX0 U16761 ( .INP(n16230), .ZN(n16229) );
  AND2X1 U16762 ( .IN1(n16231), .IN2(n16232), .Q(n16230) );
  OR2X1 U16763 ( .IN1(n16232), .IN2(n16231), .Q(n16228) );
  OR2X1 U16764 ( .IN1(n16233), .IN2(n16234), .Q(n16231) );
  AND2X1 U16765 ( .IN1(n10528), .IN2(WX2008), .Q(n16234) );
  AND2X1 U16766 ( .IN1(n9264), .IN2(n10539), .Q(n16233) );
  AND2X1 U16767 ( .IN1(n16235), .IN2(n16236), .Q(n16232) );
  INVX0 U16768 ( .INP(n16237), .ZN(n16236) );
  AND2X1 U16769 ( .IN1(n16238), .IN2(WX2072), .Q(n16237) );
  OR2X1 U16770 ( .IN1(WX2072), .IN2(n16238), .Q(n16235) );
  OR2X1 U16771 ( .IN1(n16239), .IN2(n16240), .Q(n16238) );
  AND2X1 U16772 ( .IN1(n17979), .IN2(n9912), .Q(n16240) );
  AND2X1 U16773 ( .IN1(test_so18), .IN2(n8666), .Q(n16239) );
  OR2X1 U16774 ( .IN1(n16241), .IN2(n16242), .Q(WX1941) );
  OR2X1 U16775 ( .IN1(n16243), .IN2(n16244), .Q(n16242) );
  AND2X1 U16776 ( .IN1(n10035), .IN2(CRC_OUT_8_29), .Q(n16244) );
  AND2X1 U16777 ( .IN1(n251), .IN2(n10009), .Q(n16243) );
  INVX0 U16778 ( .INP(n16245), .ZN(n251) );
  OR2X1 U16779 ( .IN1(n10631), .IN2(n4032), .Q(n16245) );
  OR2X1 U16780 ( .IN1(n16246), .IN2(n16247), .Q(n16241) );
  AND2X1 U16781 ( .IN1(n10068), .IN2(n15170), .Q(n16247) );
  OR2X1 U16782 ( .IN1(n16248), .IN2(n16249), .Q(n15170) );
  INVX0 U16783 ( .INP(n16250), .ZN(n16249) );
  OR2X1 U16784 ( .IN1(n16251), .IN2(n16252), .Q(n16250) );
  AND2X1 U16785 ( .IN1(n16252), .IN2(n16251), .Q(n16248) );
  INVX0 U16786 ( .INP(n16253), .ZN(n16251) );
  OR2X1 U16787 ( .IN1(n16254), .IN2(n16255), .Q(n16253) );
  AND2X1 U16788 ( .IN1(n10528), .IN2(n8609), .Q(n16255) );
  AND2X1 U16789 ( .IN1(n17982), .IN2(n10539), .Q(n16254) );
  OR2X1 U16790 ( .IN1(n16256), .IN2(n16257), .Q(n16252) );
  AND2X1 U16791 ( .IN1(n9703), .IN2(n16258), .Q(n16257) );
  AND2X1 U16792 ( .IN1(n16259), .IN2(n16260), .Q(n16258) );
  OR2X1 U16793 ( .IN1(n9238), .IN2(WX3363), .Q(n16260) );
  OR2X1 U16794 ( .IN1(n9239), .IN2(WX3299), .Q(n16259) );
  AND2X1 U16795 ( .IN1(n16261), .IN2(WX3427), .Q(n16256) );
  OR2X1 U16796 ( .IN1(n16262), .IN2(n16263), .Q(n16261) );
  AND2X1 U16797 ( .IN1(n9238), .IN2(WX3363), .Q(n16263) );
  AND2X1 U16798 ( .IN1(n9239), .IN2(WX3299), .Q(n16262) );
  AND2X1 U16799 ( .IN1(n9986), .IN2(n12962), .Q(n16246) );
  OR2X1 U16800 ( .IN1(n16264), .IN2(n16265), .Q(n12962) );
  INVX0 U16801 ( .INP(n16266), .ZN(n16265) );
  OR2X1 U16802 ( .IN1(n16267), .IN2(n16268), .Q(n16266) );
  AND2X1 U16803 ( .IN1(n16268), .IN2(n16267), .Q(n16264) );
  INVX0 U16804 ( .INP(n16269), .ZN(n16267) );
  OR2X1 U16805 ( .IN1(n16270), .IN2(n16271), .Q(n16269) );
  AND2X1 U16806 ( .IN1(n10528), .IN2(n8667), .Q(n16271) );
  AND2X1 U16807 ( .IN1(n17981), .IN2(n10539), .Q(n16270) );
  OR2X1 U16808 ( .IN1(n16272), .IN2(n16273), .Q(n16268) );
  AND2X1 U16809 ( .IN1(n9729), .IN2(n16274), .Q(n16273) );
  AND2X1 U16810 ( .IN1(n16275), .IN2(n16276), .Q(n16274) );
  OR2X1 U16811 ( .IN1(n9266), .IN2(WX2070), .Q(n16276) );
  OR2X1 U16812 ( .IN1(n9267), .IN2(WX2006), .Q(n16275) );
  AND2X1 U16813 ( .IN1(n16277), .IN2(WX2134), .Q(n16272) );
  OR2X1 U16814 ( .IN1(n16278), .IN2(n16279), .Q(n16277) );
  AND2X1 U16815 ( .IN1(n9266), .IN2(WX2070), .Q(n16279) );
  AND2X1 U16816 ( .IN1(n9267), .IN2(WX2006), .Q(n16278) );
  OR2X1 U16817 ( .IN1(n16280), .IN2(n16281), .Q(WX1939) );
  OR2X1 U16818 ( .IN1(n16282), .IN2(n16283), .Q(n16281) );
  AND2X1 U16819 ( .IN1(n10035), .IN2(CRC_OUT_8_30), .Q(n16283) );
  AND2X1 U16820 ( .IN1(n250), .IN2(n10009), .Q(n16282) );
  INVX0 U16821 ( .INP(n16284), .ZN(n250) );
  OR2X1 U16822 ( .IN1(n10631), .IN2(n4033), .Q(n16284) );
  OR2X1 U16823 ( .IN1(n16285), .IN2(n16286), .Q(n16280) );
  AND2X1 U16824 ( .IN1(n15194), .IN2(n10060), .Q(n16286) );
  AND2X1 U16825 ( .IN1(n16287), .IN2(n16288), .Q(n15194) );
  INVX0 U16826 ( .INP(n16289), .ZN(n16288) );
  AND2X1 U16827 ( .IN1(n16290), .IN2(n16291), .Q(n16289) );
  OR2X1 U16828 ( .IN1(n16291), .IN2(n16290), .Q(n16287) );
  OR2X1 U16829 ( .IN1(n16292), .IN2(n16293), .Q(n16290) );
  AND2X1 U16830 ( .IN1(n10528), .IN2(WX3361), .Q(n16293) );
  AND2X1 U16831 ( .IN1(n9240), .IN2(n10539), .Q(n16292) );
  AND2X1 U16832 ( .IN1(n16294), .IN2(n16295), .Q(n16291) );
  OR2X1 U16833 ( .IN1(n16296), .IN2(n9702), .Q(n16295) );
  INVX0 U16834 ( .INP(n16297), .ZN(n16296) );
  OR2X1 U16835 ( .IN1(WX3425), .IN2(n16297), .Q(n16294) );
  OR2X1 U16836 ( .IN1(n16298), .IN2(n16299), .Q(n16297) );
  AND2X1 U16837 ( .IN1(n17984), .IN2(n9964), .Q(n16299) );
  AND2X1 U16838 ( .IN1(test_so25), .IN2(n8610), .Q(n16298) );
  AND2X1 U16839 ( .IN1(n9986), .IN2(n13006), .Q(n16285) );
  OR2X1 U16840 ( .IN1(n16300), .IN2(n16301), .Q(n13006) );
  INVX0 U16841 ( .INP(n16302), .ZN(n16301) );
  OR2X1 U16842 ( .IN1(n16303), .IN2(n16304), .Q(n16302) );
  AND2X1 U16843 ( .IN1(n16304), .IN2(n16303), .Q(n16300) );
  INVX0 U16844 ( .INP(n16305), .ZN(n16303) );
  OR2X1 U16845 ( .IN1(n16306), .IN2(n16307), .Q(n16305) );
  AND2X1 U16846 ( .IN1(n10528), .IN2(n8668), .Q(n16307) );
  AND2X1 U16847 ( .IN1(n17983), .IN2(n10539), .Q(n16306) );
  OR2X1 U16848 ( .IN1(n16308), .IN2(n16309), .Q(n16304) );
  AND2X1 U16849 ( .IN1(n9728), .IN2(n16310), .Q(n16309) );
  AND2X1 U16850 ( .IN1(n16311), .IN2(n16312), .Q(n16310) );
  OR2X1 U16851 ( .IN1(n9268), .IN2(WX2068), .Q(n16312) );
  OR2X1 U16852 ( .IN1(n9269), .IN2(WX2004), .Q(n16311) );
  AND2X1 U16853 ( .IN1(n16313), .IN2(WX2132), .Q(n16308) );
  OR2X1 U16854 ( .IN1(n16314), .IN2(n16315), .Q(n16313) );
  AND2X1 U16855 ( .IN1(n9268), .IN2(WX2068), .Q(n16315) );
  AND2X1 U16856 ( .IN1(n9269), .IN2(WX2004), .Q(n16314) );
  OR2X1 U16857 ( .IN1(n16316), .IN2(n16317), .Q(WX1937) );
  OR2X1 U16858 ( .IN1(n16318), .IN2(n16319), .Q(n16317) );
  AND2X1 U16859 ( .IN1(n2245), .IN2(WX1778), .Q(n16319) );
  AND2X1 U16860 ( .IN1(n10035), .IN2(CRC_OUT_8_31), .Q(n16318) );
  OR2X1 U16861 ( .IN1(n16320), .IN2(n16321), .Q(n16316) );
  AND2X1 U16862 ( .IN1(n9986), .IN2(n13052), .Q(n16321) );
  OR2X1 U16863 ( .IN1(n16322), .IN2(n16323), .Q(n13052) );
  INVX0 U16864 ( .INP(n16324), .ZN(n16323) );
  OR2X1 U16865 ( .IN1(n16325), .IN2(n16326), .Q(n16324) );
  AND2X1 U16866 ( .IN1(n16326), .IN2(n16325), .Q(n16322) );
  INVX0 U16867 ( .INP(n16327), .ZN(n16325) );
  OR2X1 U16868 ( .IN1(n16328), .IN2(n16329), .Q(n16327) );
  AND2X1 U16869 ( .IN1(n10528), .IN2(n8669), .Q(n16329) );
  AND2X1 U16870 ( .IN1(n17986), .IN2(n10539), .Q(n16328) );
  OR2X1 U16871 ( .IN1(n16330), .IN2(n16331), .Q(n16326) );
  AND2X1 U16872 ( .IN1(n9727), .IN2(n16332), .Q(n16331) );
  AND2X1 U16873 ( .IN1(n16333), .IN2(n16334), .Q(n16332) );
  OR2X1 U16874 ( .IN1(n9042), .IN2(WX2066), .Q(n16334) );
  OR2X1 U16875 ( .IN1(n9043), .IN2(WX2002), .Q(n16333) );
  AND2X1 U16876 ( .IN1(n16335), .IN2(WX2130), .Q(n16330) );
  OR2X1 U16877 ( .IN1(n16336), .IN2(n16337), .Q(n16335) );
  AND2X1 U16878 ( .IN1(n9042), .IN2(WX2066), .Q(n16337) );
  AND2X1 U16879 ( .IN1(n9043), .IN2(WX2002), .Q(n16336) );
  AND2X1 U16880 ( .IN1(n10068), .IN2(n15214), .Q(n16320) );
  OR2X1 U16881 ( .IN1(n16338), .IN2(n16339), .Q(n15214) );
  INVX0 U16882 ( .INP(n16340), .ZN(n16339) );
  OR2X1 U16883 ( .IN1(n16341), .IN2(n16342), .Q(n16340) );
  AND2X1 U16884 ( .IN1(n16342), .IN2(n16341), .Q(n16338) );
  INVX0 U16885 ( .INP(n16343), .ZN(n16341) );
  OR2X1 U16886 ( .IN1(n16344), .IN2(n16345), .Q(n16343) );
  AND2X1 U16887 ( .IN1(n10528), .IN2(n8611), .Q(n16345) );
  AND2X1 U16888 ( .IN1(n17985), .IN2(n10539), .Q(n16344) );
  OR2X1 U16889 ( .IN1(n16346), .IN2(n16347), .Q(n16342) );
  AND2X1 U16890 ( .IN1(n9701), .IN2(n16348), .Q(n16347) );
  AND2X1 U16891 ( .IN1(n16349), .IN2(n16350), .Q(n16348) );
  OR2X1 U16892 ( .IN1(n9040), .IN2(WX3359), .Q(n16350) );
  OR2X1 U16893 ( .IN1(n9041), .IN2(WX3295), .Q(n16349) );
  AND2X1 U16894 ( .IN1(n16351), .IN2(WX3423), .Q(n16346) );
  OR2X1 U16895 ( .IN1(n16352), .IN2(n16353), .Q(n16351) );
  AND2X1 U16896 ( .IN1(n9040), .IN2(WX3359), .Q(n16353) );
  AND2X1 U16897 ( .IN1(n9041), .IN2(WX3295), .Q(n16352) );
  AND2X1 U16898 ( .IN1(n9844), .IN2(n10572), .Q(WX1839) );
  AND2X1 U16899 ( .IN1(n16354), .IN2(n10572), .Q(WX1326) );
  AND2X1 U16900 ( .IN1(n16355), .IN2(n16356), .Q(n16354) );
  OR2X1 U16901 ( .IN1(DFF_190_n1), .IN2(WX837), .Q(n16356) );
  OR2X1 U16902 ( .IN1(n9829), .IN2(CRC_OUT_9_30), .Q(n16355) );
  AND2X1 U16903 ( .IN1(n16357), .IN2(n10572), .Q(WX1324) );
  AND2X1 U16904 ( .IN1(n16358), .IN2(n16359), .Q(n16357) );
  OR2X1 U16905 ( .IN1(DFF_189_n1), .IN2(WX839), .Q(n16359) );
  OR2X1 U16906 ( .IN1(n9755), .IN2(CRC_OUT_9_29), .Q(n16358) );
  AND2X1 U16907 ( .IN1(n16360), .IN2(n10572), .Q(WX1322) );
  AND2X1 U16908 ( .IN1(n16361), .IN2(n16362), .Q(n16360) );
  OR2X1 U16909 ( .IN1(DFF_188_n1), .IN2(WX841), .Q(n16362) );
  OR2X1 U16910 ( .IN1(n9763), .IN2(CRC_OUT_9_28), .Q(n16361) );
  AND2X1 U16911 ( .IN1(n16363), .IN2(n10572), .Q(WX1320) );
  AND2X1 U16912 ( .IN1(n16364), .IN2(n16365), .Q(n16363) );
  OR2X1 U16913 ( .IN1(DFF_187_n1), .IN2(WX843), .Q(n16365) );
  OR2X1 U16914 ( .IN1(n9772), .IN2(CRC_OUT_9_27), .Q(n16364) );
  AND2X1 U16915 ( .IN1(n16366), .IN2(n10573), .Q(WX1318) );
  AND2X1 U16916 ( .IN1(n16367), .IN2(n16368), .Q(n16366) );
  OR2X1 U16917 ( .IN1(DFF_186_n1), .IN2(WX845), .Q(n16368) );
  OR2X1 U16918 ( .IN1(n9778), .IN2(CRC_OUT_9_26), .Q(n16367) );
  AND2X1 U16919 ( .IN1(n16369), .IN2(n10573), .Q(WX1316) );
  AND2X1 U16920 ( .IN1(n16370), .IN2(n16371), .Q(n16369) );
  OR2X1 U16921 ( .IN1(DFF_185_n1), .IN2(WX847), .Q(n16371) );
  OR2X1 U16922 ( .IN1(n9781), .IN2(CRC_OUT_9_25), .Q(n16370) );
  AND2X1 U16923 ( .IN1(n16372), .IN2(n10573), .Q(WX1314) );
  AND2X1 U16924 ( .IN1(n16373), .IN2(n16374), .Q(n16372) );
  OR2X1 U16925 ( .IN1(DFF_184_n1), .IN2(WX849), .Q(n16374) );
  OR2X1 U16926 ( .IN1(n9790), .IN2(CRC_OUT_9_24), .Q(n16373) );
  AND2X1 U16927 ( .IN1(n16375), .IN2(n10573), .Q(WX1312) );
  AND2X1 U16928 ( .IN1(n16376), .IN2(n16377), .Q(n16375) );
  OR2X1 U16929 ( .IN1(DFF_183_n1), .IN2(WX851), .Q(n16377) );
  OR2X1 U16930 ( .IN1(n9799), .IN2(CRC_OUT_9_23), .Q(n16376) );
  AND2X1 U16931 ( .IN1(n16378), .IN2(n10573), .Q(WX1310) );
  AND2X1 U16932 ( .IN1(n16379), .IN2(n16380), .Q(n16378) );
  OR2X1 U16933 ( .IN1(DFF_182_n1), .IN2(WX853), .Q(n16380) );
  OR2X1 U16934 ( .IN1(n9801), .IN2(CRC_OUT_9_22), .Q(n16379) );
  AND2X1 U16935 ( .IN1(n16381), .IN2(n10573), .Q(WX1308) );
  AND2X1 U16936 ( .IN1(n16382), .IN2(n16383), .Q(n16381) );
  OR2X1 U16937 ( .IN1(DFF_181_n1), .IN2(WX855), .Q(n16383) );
  OR2X1 U16938 ( .IN1(n9816), .IN2(CRC_OUT_9_21), .Q(n16382) );
  AND2X1 U16939 ( .IN1(n16384), .IN2(n10573), .Q(WX1306) );
  AND2X1 U16940 ( .IN1(n16385), .IN2(n16386), .Q(n16384) );
  OR2X1 U16941 ( .IN1(DFF_180_n1), .IN2(WX857), .Q(n16386) );
  OR2X1 U16942 ( .IN1(n9822), .IN2(CRC_OUT_9_20), .Q(n16385) );
  AND2X1 U16943 ( .IN1(n16387), .IN2(n10573), .Q(WX1304) );
  OR2X1 U16944 ( .IN1(n16388), .IN2(n16389), .Q(n16387) );
  AND2X1 U16945 ( .IN1(n9825), .IN2(n9948), .Q(n16389) );
  AND2X1 U16946 ( .IN1(test_so10), .IN2(WX859), .Q(n16388) );
  AND2X1 U16947 ( .IN1(n16390), .IN2(n10573), .Q(WX1302) );
  AND2X1 U16948 ( .IN1(n16391), .IN2(n16392), .Q(n16390) );
  OR2X1 U16949 ( .IN1(DFF_178_n1), .IN2(WX861), .Q(n16392) );
  OR2X1 U16950 ( .IN1(n9760), .IN2(CRC_OUT_9_18), .Q(n16391) );
  AND2X1 U16951 ( .IN1(n16393), .IN2(n10574), .Q(WX1300) );
  AND2X1 U16952 ( .IN1(n16394), .IN2(n16395), .Q(n16393) );
  OR2X1 U16953 ( .IN1(DFF_177_n1), .IN2(WX863), .Q(n16395) );
  OR2X1 U16954 ( .IN1(n9775), .IN2(CRC_OUT_9_17), .Q(n16394) );
  AND2X1 U16955 ( .IN1(n16396), .IN2(n10574), .Q(WX1298) );
  AND2X1 U16956 ( .IN1(n16397), .IN2(n16398), .Q(n16396) );
  OR2X1 U16957 ( .IN1(DFF_176_n1), .IN2(WX865), .Q(n16398) );
  OR2X1 U16958 ( .IN1(n9787), .IN2(CRC_OUT_9_16), .Q(n16397) );
  AND2X1 U16959 ( .IN1(n16399), .IN2(n10574), .Q(WX1296) );
  AND2X1 U16960 ( .IN1(n16400), .IN2(n16401), .Q(n16399) );
  OR2X1 U16961 ( .IN1(DFF_175_n1), .IN2(n16402), .Q(n16401) );
  AND2X1 U16962 ( .IN1(n16403), .IN2(n16404), .Q(n16402) );
  OR2X1 U16963 ( .IN1(DFF_191_n1), .IN2(n9885), .Q(n16404) );
  OR2X1 U16964 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .Q(n16403) );
  OR2X1 U16965 ( .IN1(n16405), .IN2(CRC_OUT_9_15), .Q(n16400) );
  OR2X1 U16966 ( .IN1(n16406), .IN2(n16407), .Q(n16405) );
  AND2X1 U16967 ( .IN1(DFF_191_n1), .IN2(n9885), .Q(n16407) );
  AND2X1 U16968 ( .IN1(test_so8), .IN2(CRC_OUT_9_31), .Q(n16406) );
  AND2X1 U16969 ( .IN1(n16408), .IN2(n10574), .Q(WX1294) );
  AND2X1 U16970 ( .IN1(n16409), .IN2(n16410), .Q(n16408) );
  OR2X1 U16971 ( .IN1(DFF_174_n1), .IN2(WX869), .Q(n16410) );
  OR2X1 U16972 ( .IN1(n9819), .IN2(CRC_OUT_9_14), .Q(n16409) );
  AND2X1 U16973 ( .IN1(n16411), .IN2(n10574), .Q(WX1292) );
  AND2X1 U16974 ( .IN1(n16412), .IN2(n16413), .Q(n16411) );
  OR2X1 U16975 ( .IN1(DFF_173_n1), .IN2(WX871), .Q(n16413) );
  OR2X1 U16976 ( .IN1(n9831), .IN2(CRC_OUT_9_13), .Q(n16412) );
  AND2X1 U16977 ( .IN1(n16414), .IN2(n10574), .Q(WX1290) );
  AND2X1 U16978 ( .IN1(n16415), .IN2(n16416), .Q(n16414) );
  OR2X1 U16979 ( .IN1(DFF_172_n1), .IN2(WX873), .Q(n16416) );
  OR2X1 U16980 ( .IN1(n9766), .IN2(CRC_OUT_9_12), .Q(n16415) );
  AND2X1 U16981 ( .IN1(n16417), .IN2(n10574), .Q(WX1288) );
  AND2X1 U16982 ( .IN1(n16418), .IN2(n16419), .Q(n16417) );
  OR2X1 U16983 ( .IN1(DFF_171_n1), .IN2(WX875), .Q(n16419) );
  OR2X1 U16984 ( .IN1(n9793), .IN2(CRC_OUT_9_11), .Q(n16418) );
  AND2X1 U16985 ( .IN1(n16420), .IN2(n10574), .Q(WX1286) );
  OR2X1 U16986 ( .IN1(n16421), .IN2(n16422), .Q(n16420) );
  AND2X1 U16987 ( .IN1(n16423), .IN2(CRC_OUT_9_10), .Q(n16422) );
  AND2X1 U16988 ( .IN1(DFF_170_n1), .IN2(n16424), .Q(n16421) );
  INVX0 U16989 ( .INP(n16423), .ZN(n16424) );
  OR2X1 U16990 ( .IN1(n16425), .IN2(n16426), .Q(n16423) );
  AND2X1 U16991 ( .IN1(DFF_191_n1), .IN2(WX877), .Q(n16426) );
  AND2X1 U16992 ( .IN1(n9839), .IN2(CRC_OUT_9_31), .Q(n16425) );
  AND2X1 U16993 ( .IN1(n16427), .IN2(n10574), .Q(WX1284) );
  AND2X1 U16994 ( .IN1(n16428), .IN2(n16429), .Q(n16427) );
  OR2X1 U16995 ( .IN1(DFF_169_n1), .IN2(WX879), .Q(n16429) );
  OR2X1 U16996 ( .IN1(n9784), .IN2(CRC_OUT_9_9), .Q(n16428) );
  AND2X1 U16997 ( .IN1(n16430), .IN2(n10575), .Q(WX1282) );
  AND2X1 U16998 ( .IN1(n16431), .IN2(n16432), .Q(n16430) );
  OR2X1 U16999 ( .IN1(DFF_168_n1), .IN2(WX881), .Q(n16432) );
  OR2X1 U17000 ( .IN1(n9797), .IN2(CRC_OUT_9_8), .Q(n16431) );
  AND2X1 U17001 ( .IN1(n16433), .IN2(n10575), .Q(WX1280) );
  AND2X1 U17002 ( .IN1(n16434), .IN2(n16435), .Q(n16433) );
  OR2X1 U17003 ( .IN1(DFF_167_n1), .IN2(WX883), .Q(n16435) );
  OR2X1 U17004 ( .IN1(n9806), .IN2(CRC_OUT_9_7), .Q(n16434) );
  AND2X1 U17005 ( .IN1(n16436), .IN2(n10575), .Q(WX1278) );
  AND2X1 U17006 ( .IN1(n16437), .IN2(n16438), .Q(n16436) );
  OR2X1 U17007 ( .IN1(DFF_166_n1), .IN2(WX885), .Q(n16438) );
  OR2X1 U17008 ( .IN1(n9837), .IN2(CRC_OUT_9_6), .Q(n16437) );
  AND2X1 U17009 ( .IN1(n16439), .IN2(n10575), .Q(WX1276) );
  AND2X1 U17010 ( .IN1(n16440), .IN2(n16441), .Q(n16439) );
  OR2X1 U17011 ( .IN1(DFF_165_n1), .IN2(WX887), .Q(n16441) );
  OR2X1 U17012 ( .IN1(n9824), .IN2(CRC_OUT_9_5), .Q(n16440) );
  AND2X1 U17013 ( .IN1(n16442), .IN2(n10575), .Q(WX1274) );
  AND2X1 U17014 ( .IN1(n16443), .IN2(n16444), .Q(n16442) );
  OR2X1 U17015 ( .IN1(DFF_164_n1), .IN2(WX889), .Q(n16444) );
  OR2X1 U17016 ( .IN1(n9809), .IN2(CRC_OUT_9_4), .Q(n16443) );
  AND2X1 U17017 ( .IN1(n16445), .IN2(n10575), .Q(WX1272) );
  OR2X1 U17018 ( .IN1(n16446), .IN2(n16447), .Q(n16445) );
  AND2X1 U17019 ( .IN1(n16448), .IN2(CRC_OUT_9_3), .Q(n16447) );
  AND2X1 U17020 ( .IN1(DFF_163_n1), .IN2(n16449), .Q(n16446) );
  INVX0 U17021 ( .INP(n16448), .ZN(n16449) );
  OR2X1 U17022 ( .IN1(n16450), .IN2(n16451), .Q(n16448) );
  AND2X1 U17023 ( .IN1(DFF_191_n1), .IN2(WX891), .Q(n16451) );
  AND2X1 U17024 ( .IN1(n9812), .IN2(CRC_OUT_9_31), .Q(n16450) );
  AND2X1 U17025 ( .IN1(n16452), .IN2(n10575), .Q(WX1270) );
  AND2X1 U17026 ( .IN1(n16453), .IN2(n16454), .Q(n16452) );
  OR2X1 U17027 ( .IN1(DFF_162_n1), .IN2(WX893), .Q(n16454) );
  OR2X1 U17028 ( .IN1(n9757), .IN2(CRC_OUT_9_2), .Q(n16453) );
  AND2X1 U17029 ( .IN1(n16455), .IN2(n10575), .Q(WX1268) );
  OR2X1 U17030 ( .IN1(n16456), .IN2(n16457), .Q(n16455) );
  AND2X1 U17031 ( .IN1(n9834), .IN2(n9949), .Q(n16457) );
  AND2X1 U17032 ( .IN1(test_so9), .IN2(WX895), .Q(n16456) );
  AND2X1 U17033 ( .IN1(n16458), .IN2(n10575), .Q(WX1266) );
  AND2X1 U17034 ( .IN1(n16459), .IN2(n16460), .Q(n16458) );
  INVX0 U17035 ( .INP(n16461), .ZN(n16460) );
  AND2X1 U17036 ( .IN1(CRC_OUT_9_0), .IN2(n9768), .Q(n16461) );
  OR2X1 U17037 ( .IN1(n9768), .IN2(CRC_OUT_9_0), .Q(n16459) );
  AND2X1 U17038 ( .IN1(n16462), .IN2(n10576), .Q(WX1264) );
  AND2X1 U17039 ( .IN1(n16463), .IN2(n16464), .Q(n16462) );
  OR2X1 U17040 ( .IN1(DFF_191_n1), .IN2(WX899), .Q(n16464) );
  OR2X1 U17041 ( .IN1(n9843), .IN2(CRC_OUT_9_31), .Q(n16463) );
  AND2X1 U17042 ( .IN1(n16465), .IN2(n10576), .Q(WX11670) );
  AND2X1 U17043 ( .IN1(n16466), .IN2(n16467), .Q(n16465) );
  OR2X1 U17044 ( .IN1(DFF_1726_n1), .IN2(WX11181), .Q(n16467) );
  OR2X1 U17045 ( .IN1(n9541), .IN2(CRC_OUT_1_30), .Q(n16466) );
  AND2X1 U17046 ( .IN1(n16468), .IN2(n10576), .Q(WX11668) );
  AND2X1 U17047 ( .IN1(n16469), .IN2(n16470), .Q(n16468) );
  OR2X1 U17048 ( .IN1(DFF_1725_n1), .IN2(WX11183), .Q(n16470) );
  OR2X1 U17049 ( .IN1(n9542), .IN2(CRC_OUT_1_29), .Q(n16469) );
  AND2X1 U17050 ( .IN1(n16471), .IN2(n10576), .Q(WX11666) );
  AND2X1 U17051 ( .IN1(n16472), .IN2(n16473), .Q(n16471) );
  OR2X1 U17052 ( .IN1(DFF_1724_n1), .IN2(WX11185), .Q(n16473) );
  OR2X1 U17053 ( .IN1(n9543), .IN2(CRC_OUT_1_28), .Q(n16472) );
  AND2X1 U17054 ( .IN1(n16474), .IN2(n10576), .Q(WX11664) );
  AND2X1 U17055 ( .IN1(n16475), .IN2(n16476), .Q(n16474) );
  OR2X1 U17056 ( .IN1(DFF_1723_n1), .IN2(WX11187), .Q(n16476) );
  OR2X1 U17057 ( .IN1(n9544), .IN2(CRC_OUT_1_27), .Q(n16475) );
  AND2X1 U17058 ( .IN1(n16477), .IN2(n10576), .Q(WX11662) );
  AND2X1 U17059 ( .IN1(n16478), .IN2(n16479), .Q(n16477) );
  OR2X1 U17060 ( .IN1(DFF_1722_n1), .IN2(WX11189), .Q(n16479) );
  OR2X1 U17061 ( .IN1(n9545), .IN2(CRC_OUT_1_26), .Q(n16478) );
  AND2X1 U17062 ( .IN1(n16480), .IN2(n10576), .Q(WX11660) );
  AND2X1 U17063 ( .IN1(n16481), .IN2(n16482), .Q(n16480) );
  OR2X1 U17064 ( .IN1(DFF_1721_n1), .IN2(WX11191), .Q(n16482) );
  OR2X1 U17065 ( .IN1(n9546), .IN2(CRC_OUT_1_25), .Q(n16481) );
  AND2X1 U17066 ( .IN1(n16483), .IN2(n10576), .Q(WX11658) );
  AND2X1 U17067 ( .IN1(n16484), .IN2(n16485), .Q(n16483) );
  OR2X1 U17068 ( .IN1(DFF_1720_n1), .IN2(WX11193), .Q(n16485) );
  OR2X1 U17069 ( .IN1(n9547), .IN2(CRC_OUT_1_24), .Q(n16484) );
  AND2X1 U17070 ( .IN1(n16486), .IN2(n10576), .Q(WX11656) );
  AND2X1 U17071 ( .IN1(n16487), .IN2(n16488), .Q(n16486) );
  OR2X1 U17072 ( .IN1(DFF_1719_n1), .IN2(WX11195), .Q(n16488) );
  OR2X1 U17073 ( .IN1(n9548), .IN2(CRC_OUT_1_23), .Q(n16487) );
  AND2X1 U17074 ( .IN1(n16489), .IN2(n10577), .Q(WX11654) );
  AND2X1 U17075 ( .IN1(n16490), .IN2(n16491), .Q(n16489) );
  OR2X1 U17076 ( .IN1(DFF_1718_n1), .IN2(WX11197), .Q(n16491) );
  OR2X1 U17077 ( .IN1(n9549), .IN2(CRC_OUT_1_22), .Q(n16490) );
  AND2X1 U17078 ( .IN1(n16492), .IN2(n10577), .Q(WX11652) );
  AND2X1 U17079 ( .IN1(n16493), .IN2(n16494), .Q(n16492) );
  OR2X1 U17080 ( .IN1(DFF_1717_n1), .IN2(WX11199), .Q(n16494) );
  OR2X1 U17081 ( .IN1(n9550), .IN2(CRC_OUT_1_21), .Q(n16493) );
  AND2X1 U17082 ( .IN1(n16495), .IN2(n10577), .Q(WX11650) );
  AND2X1 U17083 ( .IN1(n16496), .IN2(n16497), .Q(n16495) );
  OR2X1 U17084 ( .IN1(DFF_1716_n1), .IN2(WX11201), .Q(n16497) );
  OR2X1 U17085 ( .IN1(n9551), .IN2(CRC_OUT_1_20), .Q(n16496) );
  AND2X1 U17086 ( .IN1(n16498), .IN2(n10577), .Q(WX11648) );
  AND2X1 U17087 ( .IN1(n16499), .IN2(n16500), .Q(n16498) );
  OR2X1 U17088 ( .IN1(DFF_1715_n1), .IN2(WX11203), .Q(n16500) );
  OR2X1 U17089 ( .IN1(n9552), .IN2(CRC_OUT_1_19), .Q(n16499) );
  AND2X1 U17090 ( .IN1(n16501), .IN2(n10577), .Q(WX11646) );
  OR2X1 U17091 ( .IN1(n16502), .IN2(n16503), .Q(n16501) );
  AND2X1 U17092 ( .IN1(DFF_1714_n1), .IN2(n9913), .Q(n16503) );
  AND2X1 U17093 ( .IN1(test_so97), .IN2(CRC_OUT_1_18), .Q(n16502) );
  AND2X1 U17094 ( .IN1(n16504), .IN2(n10577), .Q(WX11644) );
  AND2X1 U17095 ( .IN1(n16505), .IN2(n16506), .Q(n16504) );
  OR2X1 U17096 ( .IN1(DFF_1713_n1), .IN2(WX11207), .Q(n16506) );
  OR2X1 U17097 ( .IN1(n9553), .IN2(CRC_OUT_1_17), .Q(n16505) );
  AND2X1 U17098 ( .IN1(n16507), .IN2(n10577), .Q(WX11642) );
  AND2X1 U17099 ( .IN1(n16508), .IN2(n16509), .Q(n16507) );
  OR2X1 U17100 ( .IN1(DFF_1712_n1), .IN2(WX11209), .Q(n16509) );
  OR2X1 U17101 ( .IN1(n9554), .IN2(CRC_OUT_1_16), .Q(n16508) );
  AND2X1 U17102 ( .IN1(n16510), .IN2(n10577), .Q(WX11640) );
  AND2X1 U17103 ( .IN1(n16511), .IN2(n16512), .Q(n16510) );
  OR2X1 U17104 ( .IN1(DFF_1711_n1), .IN2(n16513), .Q(n16512) );
  AND2X1 U17105 ( .IN1(n16514), .IN2(n16515), .Q(n16513) );
  OR2X1 U17106 ( .IN1(n9512), .IN2(n9884), .Q(n16515) );
  OR2X1 U17107 ( .IN1(test_so100), .IN2(WX11211), .Q(n16514) );
  OR2X1 U17108 ( .IN1(n16516), .IN2(CRC_OUT_1_15), .Q(n16511) );
  OR2X1 U17109 ( .IN1(n16517), .IN2(n16518), .Q(n16516) );
  AND2X1 U17110 ( .IN1(n9512), .IN2(n9884), .Q(n16518) );
  AND2X1 U17111 ( .IN1(test_so100), .IN2(WX11211), .Q(n16517) );
  AND2X1 U17112 ( .IN1(n16519), .IN2(n10578), .Q(WX11638) );
  OR2X1 U17113 ( .IN1(n16520), .IN2(n16521), .Q(n16519) );
  AND2X1 U17114 ( .IN1(n9555), .IN2(n9950), .Q(n16521) );
  AND2X1 U17115 ( .IN1(test_so99), .IN2(WX11213), .Q(n16520) );
  AND2X1 U17116 ( .IN1(n16522), .IN2(n10578), .Q(WX11636) );
  AND2X1 U17117 ( .IN1(n16523), .IN2(n16524), .Q(n16522) );
  OR2X1 U17118 ( .IN1(DFF_1709_n1), .IN2(WX11215), .Q(n16524) );
  OR2X1 U17119 ( .IN1(n9556), .IN2(CRC_OUT_1_13), .Q(n16523) );
  AND2X1 U17120 ( .IN1(n16525), .IN2(n10578), .Q(WX11634) );
  AND2X1 U17121 ( .IN1(n16526), .IN2(n16527), .Q(n16525) );
  OR2X1 U17122 ( .IN1(DFF_1708_n1), .IN2(WX11217), .Q(n16527) );
  OR2X1 U17123 ( .IN1(n9557), .IN2(CRC_OUT_1_12), .Q(n16526) );
  AND2X1 U17124 ( .IN1(n16528), .IN2(n10578), .Q(WX11632) );
  AND2X1 U17125 ( .IN1(n16529), .IN2(n16530), .Q(n16528) );
  OR2X1 U17126 ( .IN1(DFF_1707_n1), .IN2(WX11219), .Q(n16530) );
  OR2X1 U17127 ( .IN1(n9558), .IN2(CRC_OUT_1_11), .Q(n16529) );
  AND2X1 U17128 ( .IN1(n16531), .IN2(n10578), .Q(WX11630) );
  AND2X1 U17129 ( .IN1(n16532), .IN2(n16533), .Q(n16531) );
  OR2X1 U17130 ( .IN1(DFF_1706_n1), .IN2(n16534), .Q(n16533) );
  AND2X1 U17131 ( .IN1(n16535), .IN2(n16536), .Q(n16534) );
  OR2X1 U17132 ( .IN1(n9513), .IN2(n9884), .Q(n16536) );
  OR2X1 U17133 ( .IN1(test_so100), .IN2(WX11221), .Q(n16535) );
  OR2X1 U17134 ( .IN1(n16537), .IN2(CRC_OUT_1_10), .Q(n16532) );
  OR2X1 U17135 ( .IN1(n16538), .IN2(n16539), .Q(n16537) );
  AND2X1 U17136 ( .IN1(n9513), .IN2(n9884), .Q(n16539) );
  AND2X1 U17137 ( .IN1(test_so100), .IN2(WX11221), .Q(n16538) );
  AND2X1 U17138 ( .IN1(n16540), .IN2(n10578), .Q(WX11628) );
  AND2X1 U17139 ( .IN1(n16541), .IN2(n16542), .Q(n16540) );
  OR2X1 U17140 ( .IN1(DFF_1705_n1), .IN2(WX11223), .Q(n16542) );
  OR2X1 U17141 ( .IN1(n9559), .IN2(CRC_OUT_1_9), .Q(n16541) );
  AND2X1 U17142 ( .IN1(n16543), .IN2(n10578), .Q(WX11626) );
  AND2X1 U17143 ( .IN1(n16544), .IN2(n16545), .Q(n16543) );
  OR2X1 U17144 ( .IN1(DFF_1704_n1), .IN2(WX11225), .Q(n16545) );
  OR2X1 U17145 ( .IN1(n9560), .IN2(CRC_OUT_1_8), .Q(n16544) );
  AND2X1 U17146 ( .IN1(n16546), .IN2(n10578), .Q(WX11624) );
  AND2X1 U17147 ( .IN1(n16547), .IN2(n16548), .Q(n16546) );
  OR2X1 U17148 ( .IN1(DFF_1703_n1), .IN2(WX11227), .Q(n16548) );
  OR2X1 U17149 ( .IN1(n9561), .IN2(CRC_OUT_1_7), .Q(n16547) );
  AND2X1 U17150 ( .IN1(n16549), .IN2(n10578), .Q(WX11622) );
  AND2X1 U17151 ( .IN1(n16550), .IN2(n16551), .Q(n16549) );
  OR2X1 U17152 ( .IN1(DFF_1702_n1), .IN2(WX11229), .Q(n16551) );
  OR2X1 U17153 ( .IN1(n9562), .IN2(CRC_OUT_1_6), .Q(n16550) );
  AND2X1 U17154 ( .IN1(n16552), .IN2(n10579), .Q(WX11620) );
  AND2X1 U17155 ( .IN1(n16553), .IN2(n16554), .Q(n16552) );
  OR2X1 U17156 ( .IN1(DFF_1701_n1), .IN2(WX11231), .Q(n16554) );
  OR2X1 U17157 ( .IN1(n9563), .IN2(CRC_OUT_1_5), .Q(n16553) );
  AND2X1 U17158 ( .IN1(n16555), .IN2(n10579), .Q(WX11618) );
  AND2X1 U17159 ( .IN1(n16556), .IN2(n16557), .Q(n16555) );
  OR2X1 U17160 ( .IN1(DFF_1700_n1), .IN2(WX11233), .Q(n16557) );
  OR2X1 U17161 ( .IN1(n9564), .IN2(CRC_OUT_1_4), .Q(n16556) );
  AND2X1 U17162 ( .IN1(n16558), .IN2(n10579), .Q(WX11616) );
  AND2X1 U17163 ( .IN1(n16559), .IN2(n16560), .Q(n16558) );
  OR2X1 U17164 ( .IN1(DFF_1699_n1), .IN2(n16561), .Q(n16560) );
  AND2X1 U17165 ( .IN1(n16562), .IN2(n16563), .Q(n16561) );
  OR2X1 U17166 ( .IN1(n9514), .IN2(n9884), .Q(n16563) );
  OR2X1 U17167 ( .IN1(test_so100), .IN2(WX11235), .Q(n16562) );
  OR2X1 U17168 ( .IN1(n16564), .IN2(CRC_OUT_1_3), .Q(n16559) );
  OR2X1 U17169 ( .IN1(n16565), .IN2(n16566), .Q(n16564) );
  AND2X1 U17170 ( .IN1(n9514), .IN2(n9884), .Q(n16566) );
  AND2X1 U17171 ( .IN1(test_so100), .IN2(WX11235), .Q(n16565) );
  AND2X1 U17172 ( .IN1(n16567), .IN2(n10579), .Q(WX11614) );
  AND2X1 U17173 ( .IN1(n16568), .IN2(n16569), .Q(n16567) );
  OR2X1 U17174 ( .IN1(DFF_1698_n1), .IN2(WX11237), .Q(n16569) );
  OR2X1 U17175 ( .IN1(n9565), .IN2(CRC_OUT_1_2), .Q(n16568) );
  AND2X1 U17176 ( .IN1(n16570), .IN2(n10579), .Q(WX11612) );
  OR2X1 U17177 ( .IN1(n16571), .IN2(n16572), .Q(n16570) );
  AND2X1 U17178 ( .IN1(DFF_1697_n1), .IN2(n9906), .Q(n16572) );
  AND2X1 U17179 ( .IN1(test_so98), .IN2(CRC_OUT_1_1), .Q(n16571) );
  AND2X1 U17180 ( .IN1(n16573), .IN2(n10579), .Q(WX11610) );
  AND2X1 U17181 ( .IN1(n16574), .IN2(n16575), .Q(n16573) );
  OR2X1 U17182 ( .IN1(DFF_1696_n1), .IN2(WX11241), .Q(n16575) );
  OR2X1 U17183 ( .IN1(n9566), .IN2(CRC_OUT_1_0), .Q(n16574) );
  AND2X1 U17184 ( .IN1(n16576), .IN2(n10579), .Q(WX11608) );
  OR2X1 U17185 ( .IN1(n16577), .IN2(n16578), .Q(n16576) );
  AND2X1 U17186 ( .IN1(n9533), .IN2(n9884), .Q(n16578) );
  AND2X1 U17187 ( .IN1(test_so100), .IN2(WX11243), .Q(n16577) );
  AND2X1 U17188 ( .IN1(n10591), .IN2(n8246), .Q(WX11082) );
  AND2X1 U17189 ( .IN1(n10591), .IN2(n8247), .Q(WX11080) );
  AND2X1 U17190 ( .IN1(n10592), .IN2(n8248), .Q(WX11078) );
  AND2X1 U17191 ( .IN1(n10591), .IN2(n8249), .Q(WX11076) );
  AND2X1 U17192 ( .IN1(n10591), .IN2(n8250), .Q(WX11074) );
  AND2X1 U17193 ( .IN1(n10590), .IN2(n8251), .Q(WX11072) );
  AND2X1 U17194 ( .IN1(n10591), .IN2(n8252), .Q(WX11070) );
  AND2X1 U17195 ( .IN1(n10590), .IN2(n8253), .Q(WX11068) );
  AND2X1 U17196 ( .IN1(n10592), .IN2(n8254), .Q(WX11066) );
  AND2X1 U17197 ( .IN1(test_so91), .IN2(n10579), .Q(WX11064) );
  AND2X1 U17198 ( .IN1(n10591), .IN2(n8257), .Q(WX11062) );
  AND2X1 U17199 ( .IN1(n10590), .IN2(n8258), .Q(WX11060) );
  AND2X1 U17200 ( .IN1(n10590), .IN2(n8259), .Q(WX11058) );
  AND2X1 U17201 ( .IN1(n10590), .IN2(n8260), .Q(WX11056) );
  AND2X1 U17202 ( .IN1(n10592), .IN2(n8261), .Q(WX11054) );
  AND2X1 U17203 ( .IN1(n10590), .IN2(n8262), .Q(WX11052) );
  OR2X1 U17204 ( .IN1(n16579), .IN2(n16580), .Q(WX11050) );
  OR2X1 U17205 ( .IN1(n16581), .IN2(n16582), .Q(n16580) );
  AND2X1 U17206 ( .IN1(n10035), .IN2(CRC_OUT_1_0), .Q(n16582) );
  AND2X1 U17207 ( .IN1(DATA_0_0), .IN2(n10059), .Q(n16581) );
  OR2X1 U17208 ( .IN1(n16583), .IN2(n16584), .Q(n16579) );
  AND2X1 U17209 ( .IN1(n1968), .IN2(n10009), .Q(n16584) );
  INVX0 U17210 ( .INP(n16585), .ZN(n1968) );
  OR2X1 U17211 ( .IN1(n10631), .IN2(n3786), .Q(n16585) );
  AND2X1 U17212 ( .IN1(n9986), .IN2(n10895), .Q(n16583) );
  OR2X1 U17213 ( .IN1(n16586), .IN2(n16587), .Q(n10895) );
  INVX0 U17214 ( .INP(n16588), .ZN(n16587) );
  OR2X1 U17215 ( .IN1(n16589), .IN2(n16590), .Q(n16588) );
  AND2X1 U17216 ( .IN1(n16590), .IN2(n16589), .Q(n16586) );
  AND2X1 U17217 ( .IN1(n16591), .IN2(n16592), .Q(n16589) );
  OR2X1 U17218 ( .IN1(WX11115), .IN2(n9270), .Q(n16592) );
  OR2X1 U17219 ( .IN1(WX11051), .IN2(n3531), .Q(n16591) );
  OR2X1 U17220 ( .IN1(n16593), .IN2(n16594), .Q(n16590) );
  AND2X1 U17221 ( .IN1(n9271), .IN2(WX11243), .Q(n16594) );
  AND2X1 U17222 ( .IN1(n9533), .IN2(WX11179), .Q(n16593) );
  OR2X1 U17223 ( .IN1(n16595), .IN2(n16596), .Q(WX11048) );
  OR2X1 U17224 ( .IN1(n16597), .IN2(n16598), .Q(n16596) );
  AND2X1 U17225 ( .IN1(n10035), .IN2(CRC_OUT_1_1), .Q(n16598) );
  AND2X1 U17226 ( .IN1(DATA_0_1), .IN2(n10060), .Q(n16597) );
  OR2X1 U17227 ( .IN1(n16599), .IN2(n16600), .Q(n16595) );
  AND2X1 U17228 ( .IN1(n1967), .IN2(n10009), .Q(n16600) );
  INVX0 U17229 ( .INP(n16601), .ZN(n1967) );
  OR2X1 U17230 ( .IN1(n10631), .IN2(n3787), .Q(n16601) );
  AND2X1 U17231 ( .IN1(n9986), .IN2(n10905), .Q(n16599) );
  OR2X1 U17232 ( .IN1(n16602), .IN2(n16603), .Q(n10905) );
  INVX0 U17233 ( .INP(n16604), .ZN(n16603) );
  OR2X1 U17234 ( .IN1(n16605), .IN2(n16606), .Q(n16604) );
  AND2X1 U17235 ( .IN1(n16606), .IN2(n16605), .Q(n16602) );
  AND2X1 U17236 ( .IN1(n16607), .IN2(n16608), .Q(n16605) );
  OR2X1 U17237 ( .IN1(WX11113), .IN2(n9272), .Q(n16608) );
  OR2X1 U17238 ( .IN1(WX11049), .IN2(n3533), .Q(n16607) );
  OR2X1 U17239 ( .IN1(n16609), .IN2(n16610), .Q(n16606) );
  AND2X1 U17240 ( .IN1(n9273), .IN2(WX11241), .Q(n16610) );
  AND2X1 U17241 ( .IN1(n9566), .IN2(WX11177), .Q(n16609) );
  OR2X1 U17242 ( .IN1(n16611), .IN2(n16612), .Q(WX11046) );
  OR2X1 U17243 ( .IN1(n16613), .IN2(n16614), .Q(n16612) );
  AND2X1 U17244 ( .IN1(n10035), .IN2(CRC_OUT_1_2), .Q(n16614) );
  AND2X1 U17245 ( .IN1(DATA_0_2), .IN2(n10061), .Q(n16613) );
  OR2X1 U17246 ( .IN1(n16615), .IN2(n16616), .Q(n16611) );
  AND2X1 U17247 ( .IN1(n1966), .IN2(n10009), .Q(n16616) );
  INVX0 U17248 ( .INP(n16617), .ZN(n1966) );
  OR2X1 U17249 ( .IN1(n10631), .IN2(n3788), .Q(n16617) );
  AND2X1 U17250 ( .IN1(n10914), .IN2(n9973), .Q(n16615) );
  AND2X1 U17251 ( .IN1(n16618), .IN2(n16619), .Q(n10914) );
  INVX0 U17252 ( .INP(n16620), .ZN(n16619) );
  AND2X1 U17253 ( .IN1(n16621), .IN2(n16622), .Q(n16620) );
  OR2X1 U17254 ( .IN1(n16622), .IN2(n16621), .Q(n16618) );
  OR2X1 U17255 ( .IN1(n16623), .IN2(n16624), .Q(n16621) );
  AND2X1 U17256 ( .IN1(n3535), .IN2(WX11047), .Q(n16624) );
  INVX0 U17257 ( .INP(n16625), .ZN(n16623) );
  OR2X1 U17258 ( .IN1(WX11047), .IN2(n3535), .Q(n16625) );
  AND2X1 U17259 ( .IN1(n16626), .IN2(n16627), .Q(n16622) );
  OR2X1 U17260 ( .IN1(WX11175), .IN2(test_so98), .Q(n16627) );
  OR2X1 U17261 ( .IN1(n9906), .IN2(n9275), .Q(n16626) );
  OR2X1 U17262 ( .IN1(n16628), .IN2(n16629), .Q(WX11044) );
  OR2X1 U17263 ( .IN1(n16630), .IN2(n16631), .Q(n16629) );
  AND2X1 U17264 ( .IN1(n10035), .IN2(CRC_OUT_1_3), .Q(n16631) );
  AND2X1 U17265 ( .IN1(DATA_0_3), .IN2(n10061), .Q(n16630) );
  OR2X1 U17266 ( .IN1(n16632), .IN2(n16633), .Q(n16628) );
  AND2X1 U17267 ( .IN1(n1965), .IN2(n10009), .Q(n16633) );
  INVX0 U17268 ( .INP(n16634), .ZN(n1965) );
  OR2X1 U17269 ( .IN1(n10631), .IN2(n3789), .Q(n16634) );
  AND2X1 U17270 ( .IN1(n9986), .IN2(n10923), .Q(n16632) );
  OR2X1 U17271 ( .IN1(n16635), .IN2(n16636), .Q(n10923) );
  INVX0 U17272 ( .INP(n16637), .ZN(n16636) );
  OR2X1 U17273 ( .IN1(n16638), .IN2(n16639), .Q(n16637) );
  AND2X1 U17274 ( .IN1(n16639), .IN2(n16638), .Q(n16635) );
  AND2X1 U17275 ( .IN1(n16640), .IN2(n16641), .Q(n16638) );
  OR2X1 U17276 ( .IN1(WX11109), .IN2(n9276), .Q(n16641) );
  OR2X1 U17277 ( .IN1(WX11045), .IN2(n3537), .Q(n16640) );
  OR2X1 U17278 ( .IN1(n16642), .IN2(n16643), .Q(n16639) );
  AND2X1 U17279 ( .IN1(n9277), .IN2(WX11237), .Q(n16643) );
  AND2X1 U17280 ( .IN1(n9565), .IN2(WX11173), .Q(n16642) );
  OR2X1 U17281 ( .IN1(n16644), .IN2(n16645), .Q(WX11042) );
  OR2X1 U17282 ( .IN1(n16646), .IN2(n16647), .Q(n16645) );
  AND2X1 U17283 ( .IN1(n10035), .IN2(CRC_OUT_1_4), .Q(n16647) );
  AND2X1 U17284 ( .IN1(DATA_0_4), .IN2(n10061), .Q(n16646) );
  OR2X1 U17285 ( .IN1(n16648), .IN2(n16649), .Q(n16644) );
  AND2X1 U17286 ( .IN1(n1964), .IN2(n10009), .Q(n16649) );
  INVX0 U17287 ( .INP(n16650), .ZN(n1964) );
  OR2X1 U17288 ( .IN1(n10631), .IN2(n3790), .Q(n16650) );
  AND2X1 U17289 ( .IN1(n10932), .IN2(n9973), .Q(n16648) );
  AND2X1 U17290 ( .IN1(n16651), .IN2(n16652), .Q(n10932) );
  INVX0 U17291 ( .INP(n16653), .ZN(n16652) );
  AND2X1 U17292 ( .IN1(n16654), .IN2(n16655), .Q(n16653) );
  OR2X1 U17293 ( .IN1(n16655), .IN2(n16654), .Q(n16651) );
  OR2X1 U17294 ( .IN1(n16656), .IN2(n16657), .Q(n16654) );
  AND2X1 U17295 ( .IN1(n3539), .IN2(WX11043), .Q(n16657) );
  INVX0 U17296 ( .INP(n16658), .ZN(n16656) );
  OR2X1 U17297 ( .IN1(WX11043), .IN2(n3539), .Q(n16658) );
  AND2X1 U17298 ( .IN1(n16659), .IN2(n16660), .Q(n16655) );
  OR2X1 U17299 ( .IN1(WX11235), .IN2(test_so96), .Q(n16660) );
  OR2X1 U17300 ( .IN1(n9934), .IN2(n9514), .Q(n16659) );
  OR2X1 U17301 ( .IN1(n16661), .IN2(n16662), .Q(WX11040) );
  OR2X1 U17302 ( .IN1(n16663), .IN2(n16664), .Q(n16662) );
  AND2X1 U17303 ( .IN1(n10035), .IN2(CRC_OUT_1_5), .Q(n16664) );
  AND2X1 U17304 ( .IN1(DATA_0_5), .IN2(n10061), .Q(n16663) );
  OR2X1 U17305 ( .IN1(n16665), .IN2(n16666), .Q(n16661) );
  AND2X1 U17306 ( .IN1(n1963), .IN2(n10009), .Q(n16666) );
  INVX0 U17307 ( .INP(n16667), .ZN(n1963) );
  OR2X1 U17308 ( .IN1(n10631), .IN2(n3791), .Q(n16667) );
  AND2X1 U17309 ( .IN1(n9986), .IN2(n10941), .Q(n16665) );
  OR2X1 U17310 ( .IN1(n16668), .IN2(n16669), .Q(n10941) );
  INVX0 U17311 ( .INP(n16670), .ZN(n16669) );
  OR2X1 U17312 ( .IN1(n16671), .IN2(n16672), .Q(n16670) );
  AND2X1 U17313 ( .IN1(n16672), .IN2(n16671), .Q(n16668) );
  AND2X1 U17314 ( .IN1(n16673), .IN2(n16674), .Q(n16671) );
  OR2X1 U17315 ( .IN1(WX11105), .IN2(n9279), .Q(n16674) );
  OR2X1 U17316 ( .IN1(WX11041), .IN2(n3541), .Q(n16673) );
  OR2X1 U17317 ( .IN1(n16675), .IN2(n16676), .Q(n16672) );
  AND2X1 U17318 ( .IN1(n9280), .IN2(WX11233), .Q(n16676) );
  AND2X1 U17319 ( .IN1(n9564), .IN2(WX11169), .Q(n16675) );
  OR2X1 U17320 ( .IN1(n16677), .IN2(n16678), .Q(WX11038) );
  OR2X1 U17321 ( .IN1(n16679), .IN2(n16680), .Q(n16678) );
  AND2X1 U17322 ( .IN1(n10035), .IN2(CRC_OUT_1_6), .Q(n16680) );
  AND2X1 U17323 ( .IN1(DATA_0_6), .IN2(n10061), .Q(n16679) );
  OR2X1 U17324 ( .IN1(n16681), .IN2(n16682), .Q(n16677) );
  AND2X1 U17325 ( .IN1(n1962), .IN2(n10009), .Q(n16682) );
  INVX0 U17326 ( .INP(n16683), .ZN(n1962) );
  OR2X1 U17327 ( .IN1(n10631), .IN2(n3792), .Q(n16683) );
  AND2X1 U17328 ( .IN1(n10950), .IN2(n9973), .Q(n16681) );
  AND2X1 U17329 ( .IN1(n16684), .IN2(n16685), .Q(n10950) );
  INVX0 U17330 ( .INP(n16686), .ZN(n16685) );
  AND2X1 U17331 ( .IN1(n16687), .IN2(n16688), .Q(n16686) );
  OR2X1 U17332 ( .IN1(n16688), .IN2(n16687), .Q(n16684) );
  OR2X1 U17333 ( .IN1(n16689), .IN2(n16690), .Q(n16687) );
  AND2X1 U17334 ( .IN1(n9281), .IN2(WX11167), .Q(n16690) );
  INVX0 U17335 ( .INP(n16691), .ZN(n16689) );
  OR2X1 U17336 ( .IN1(WX11167), .IN2(n9281), .Q(n16691) );
  AND2X1 U17337 ( .IN1(n16692), .IN2(n16693), .Q(n16688) );
  OR2X1 U17338 ( .IN1(WX11231), .IN2(test_so94), .Q(n16693) );
  OR2X1 U17339 ( .IN1(n9935), .IN2(n9563), .Q(n16692) );
  OR2X1 U17340 ( .IN1(n16694), .IN2(n16695), .Q(WX11036) );
  OR2X1 U17341 ( .IN1(n16696), .IN2(n16697), .Q(n16695) );
  AND2X1 U17342 ( .IN1(n10035), .IN2(CRC_OUT_1_7), .Q(n16697) );
  AND2X1 U17343 ( .IN1(DATA_0_7), .IN2(n10062), .Q(n16696) );
  OR2X1 U17344 ( .IN1(n16698), .IN2(n16699), .Q(n16694) );
  AND2X1 U17345 ( .IN1(n1961), .IN2(n10009), .Q(n16699) );
  INVX0 U17346 ( .INP(n16700), .ZN(n1961) );
  OR2X1 U17347 ( .IN1(n10630), .IN2(n3793), .Q(n16700) );
  AND2X1 U17348 ( .IN1(n9986), .IN2(n10959), .Q(n16698) );
  OR2X1 U17349 ( .IN1(n16701), .IN2(n16702), .Q(n10959) );
  INVX0 U17350 ( .INP(n16703), .ZN(n16702) );
  OR2X1 U17351 ( .IN1(n16704), .IN2(n16705), .Q(n16703) );
  AND2X1 U17352 ( .IN1(n16705), .IN2(n16704), .Q(n16701) );
  AND2X1 U17353 ( .IN1(n16706), .IN2(n16707), .Q(n16704) );
  OR2X1 U17354 ( .IN1(WX11101), .IN2(n9283), .Q(n16707) );
  OR2X1 U17355 ( .IN1(WX11037), .IN2(n3545), .Q(n16706) );
  OR2X1 U17356 ( .IN1(n16708), .IN2(n16709), .Q(n16705) );
  AND2X1 U17357 ( .IN1(n9284), .IN2(WX11229), .Q(n16709) );
  AND2X1 U17358 ( .IN1(n9562), .IN2(WX11165), .Q(n16708) );
  OR2X1 U17359 ( .IN1(n16710), .IN2(n16711), .Q(WX11034) );
  OR2X1 U17360 ( .IN1(n16712), .IN2(n16713), .Q(n16711) );
  AND2X1 U17361 ( .IN1(n10035), .IN2(CRC_OUT_1_8), .Q(n16713) );
  AND2X1 U17362 ( .IN1(DATA_0_8), .IN2(n10062), .Q(n16712) );
  OR2X1 U17363 ( .IN1(n16714), .IN2(n16715), .Q(n16710) );
  AND2X1 U17364 ( .IN1(n1960), .IN2(n10009), .Q(n16715) );
  INVX0 U17365 ( .INP(n16716), .ZN(n1960) );
  OR2X1 U17366 ( .IN1(n10630), .IN2(n3794), .Q(n16716) );
  AND2X1 U17367 ( .IN1(n10968), .IN2(n9973), .Q(n16714) );
  AND2X1 U17368 ( .IN1(n16717), .IN2(n16718), .Q(n10968) );
  INVX0 U17369 ( .INP(n16719), .ZN(n16718) );
  AND2X1 U17370 ( .IN1(n16720), .IN2(n16721), .Q(n16719) );
  OR2X1 U17371 ( .IN1(n16721), .IN2(n16720), .Q(n16717) );
  OR2X1 U17372 ( .IN1(n16722), .IN2(n16723), .Q(n16720) );
  AND2X1 U17373 ( .IN1(n3547), .IN2(WX11163), .Q(n16723) );
  INVX0 U17374 ( .INP(n16724), .ZN(n16722) );
  OR2X1 U17375 ( .IN1(WX11163), .IN2(n3547), .Q(n16724) );
  AND2X1 U17376 ( .IN1(n16725), .IN2(n16726), .Q(n16721) );
  OR2X1 U17377 ( .IN1(WX11227), .IN2(test_so92), .Q(n16726) );
  OR2X1 U17378 ( .IN1(n9936), .IN2(n9561), .Q(n16725) );
  OR2X1 U17379 ( .IN1(n16727), .IN2(n16728), .Q(WX11032) );
  OR2X1 U17380 ( .IN1(n16729), .IN2(n16730), .Q(n16728) );
  AND2X1 U17381 ( .IN1(n10035), .IN2(CRC_OUT_1_9), .Q(n16730) );
  AND2X1 U17382 ( .IN1(DATA_0_9), .IN2(n10062), .Q(n16729) );
  OR2X1 U17383 ( .IN1(n16731), .IN2(n16732), .Q(n16727) );
  AND2X1 U17384 ( .IN1(n1959), .IN2(n10009), .Q(n16732) );
  INVX0 U17385 ( .INP(n16733), .ZN(n1959) );
  OR2X1 U17386 ( .IN1(n10630), .IN2(n3795), .Q(n16733) );
  AND2X1 U17387 ( .IN1(n9986), .IN2(n10977), .Q(n16731) );
  OR2X1 U17388 ( .IN1(n16734), .IN2(n16735), .Q(n10977) );
  INVX0 U17389 ( .INP(n16736), .ZN(n16735) );
  OR2X1 U17390 ( .IN1(n16737), .IN2(n16738), .Q(n16736) );
  AND2X1 U17391 ( .IN1(n16738), .IN2(n16737), .Q(n16734) );
  AND2X1 U17392 ( .IN1(n16739), .IN2(n16740), .Q(n16737) );
  OR2X1 U17393 ( .IN1(WX11097), .IN2(n9286), .Q(n16740) );
  OR2X1 U17394 ( .IN1(WX11033), .IN2(n3549), .Q(n16739) );
  OR2X1 U17395 ( .IN1(n16741), .IN2(n16742), .Q(n16738) );
  AND2X1 U17396 ( .IN1(n9287), .IN2(WX11225), .Q(n16742) );
  AND2X1 U17397 ( .IN1(n9560), .IN2(WX11161), .Q(n16741) );
  OR2X1 U17398 ( .IN1(n16743), .IN2(n16744), .Q(WX11030) );
  OR2X1 U17399 ( .IN1(n16745), .IN2(n16746), .Q(n16744) );
  AND2X1 U17400 ( .IN1(n10036), .IN2(CRC_OUT_1_10), .Q(n16746) );
  AND2X1 U17401 ( .IN1(DATA_0_10), .IN2(n10062), .Q(n16745) );
  OR2X1 U17402 ( .IN1(n16747), .IN2(n16748), .Q(n16743) );
  AND2X1 U17403 ( .IN1(n1958), .IN2(n10010), .Q(n16748) );
  INVX0 U17404 ( .INP(n16749), .ZN(n1958) );
  OR2X1 U17405 ( .IN1(n10630), .IN2(n3796), .Q(n16749) );
  AND2X1 U17406 ( .IN1(n9986), .IN2(n10986), .Q(n16747) );
  OR2X1 U17407 ( .IN1(n16750), .IN2(n16751), .Q(n10986) );
  INVX0 U17408 ( .INP(n16752), .ZN(n16751) );
  OR2X1 U17409 ( .IN1(n16753), .IN2(n16754), .Q(n16752) );
  AND2X1 U17410 ( .IN1(n16754), .IN2(n16753), .Q(n16750) );
  AND2X1 U17411 ( .IN1(n16755), .IN2(n16756), .Q(n16753) );
  OR2X1 U17412 ( .IN1(WX11095), .IN2(n9288), .Q(n16756) );
  OR2X1 U17413 ( .IN1(WX11031), .IN2(n3551), .Q(n16755) );
  OR2X1 U17414 ( .IN1(n16757), .IN2(n16758), .Q(n16754) );
  AND2X1 U17415 ( .IN1(n9289), .IN2(WX11223), .Q(n16758) );
  AND2X1 U17416 ( .IN1(n9559), .IN2(WX11159), .Q(n16757) );
  OR2X1 U17417 ( .IN1(n16759), .IN2(n16760), .Q(WX11028) );
  OR2X1 U17418 ( .IN1(n16761), .IN2(n16762), .Q(n16760) );
  AND2X1 U17419 ( .IN1(n10036), .IN2(CRC_OUT_1_11), .Q(n16762) );
  AND2X1 U17420 ( .IN1(DATA_0_11), .IN2(n10060), .Q(n16761) );
  OR2X1 U17421 ( .IN1(n16763), .IN2(n16764), .Q(n16759) );
  AND2X1 U17422 ( .IN1(n1957), .IN2(n10010), .Q(n16764) );
  INVX0 U17423 ( .INP(n16765), .ZN(n1957) );
  OR2X1 U17424 ( .IN1(n10630), .IN2(n3797), .Q(n16765) );
  AND2X1 U17425 ( .IN1(n9986), .IN2(n10995), .Q(n16763) );
  OR2X1 U17426 ( .IN1(n16766), .IN2(n16767), .Q(n10995) );
  INVX0 U17427 ( .INP(n16768), .ZN(n16767) );
  OR2X1 U17428 ( .IN1(n16769), .IN2(n16770), .Q(n16768) );
  AND2X1 U17429 ( .IN1(n16770), .IN2(n16769), .Q(n16766) );
  AND2X1 U17430 ( .IN1(n16771), .IN2(n16772), .Q(n16769) );
  OR2X1 U17431 ( .IN1(WX11093), .IN2(n9290), .Q(n16772) );
  OR2X1 U17432 ( .IN1(WX11029), .IN2(n3553), .Q(n16771) );
  OR2X1 U17433 ( .IN1(n16773), .IN2(n16774), .Q(n16770) );
  AND2X1 U17434 ( .IN1(n9291), .IN2(WX11221), .Q(n16774) );
  AND2X1 U17435 ( .IN1(n9513), .IN2(WX11157), .Q(n16773) );
  OR2X1 U17436 ( .IN1(n16775), .IN2(n16776), .Q(WX11026) );
  OR2X1 U17437 ( .IN1(n16777), .IN2(n16778), .Q(n16776) );
  AND2X1 U17438 ( .IN1(n10036), .IN2(CRC_OUT_1_12), .Q(n16778) );
  AND2X1 U17439 ( .IN1(DATA_0_12), .IN2(n10062), .Q(n16777) );
  OR2X1 U17440 ( .IN1(n16779), .IN2(n16780), .Q(n16775) );
  AND2X1 U17441 ( .IN1(n1956), .IN2(n10010), .Q(n16780) );
  INVX0 U17442 ( .INP(n16781), .ZN(n1956) );
  OR2X1 U17443 ( .IN1(n10630), .IN2(n3798), .Q(n16781) );
  AND2X1 U17444 ( .IN1(n9985), .IN2(n11004), .Q(n16779) );
  OR2X1 U17445 ( .IN1(n16782), .IN2(n16783), .Q(n11004) );
  INVX0 U17446 ( .INP(n16784), .ZN(n16783) );
  OR2X1 U17447 ( .IN1(n16785), .IN2(n16786), .Q(n16784) );
  AND2X1 U17448 ( .IN1(n16786), .IN2(n16785), .Q(n16782) );
  AND2X1 U17449 ( .IN1(n16787), .IN2(n16788), .Q(n16785) );
  OR2X1 U17450 ( .IN1(WX11091), .IN2(n9292), .Q(n16788) );
  OR2X1 U17451 ( .IN1(WX11027), .IN2(n3555), .Q(n16787) );
  OR2X1 U17452 ( .IN1(n16789), .IN2(n16790), .Q(n16786) );
  AND2X1 U17453 ( .IN1(n9293), .IN2(WX11219), .Q(n16790) );
  AND2X1 U17454 ( .IN1(n9558), .IN2(WX11155), .Q(n16789) );
  OR2X1 U17455 ( .IN1(n16791), .IN2(n16792), .Q(WX11024) );
  OR2X1 U17456 ( .IN1(n16793), .IN2(n16794), .Q(n16792) );
  AND2X1 U17457 ( .IN1(n10036), .IN2(CRC_OUT_1_13), .Q(n16794) );
  AND2X1 U17458 ( .IN1(DATA_0_13), .IN2(n10062), .Q(n16793) );
  OR2X1 U17459 ( .IN1(n16795), .IN2(n16796), .Q(n16791) );
  AND2X1 U17460 ( .IN1(n1955), .IN2(n10010), .Q(n16796) );
  INVX0 U17461 ( .INP(n16797), .ZN(n1955) );
  OR2X1 U17462 ( .IN1(n10630), .IN2(n3799), .Q(n16797) );
  AND2X1 U17463 ( .IN1(n9985), .IN2(n11013), .Q(n16795) );
  OR2X1 U17464 ( .IN1(n16798), .IN2(n16799), .Q(n11013) );
  INVX0 U17465 ( .INP(n16800), .ZN(n16799) );
  OR2X1 U17466 ( .IN1(n16801), .IN2(n16802), .Q(n16800) );
  AND2X1 U17467 ( .IN1(n16802), .IN2(n16801), .Q(n16798) );
  AND2X1 U17468 ( .IN1(n16803), .IN2(n16804), .Q(n16801) );
  OR2X1 U17469 ( .IN1(WX11089), .IN2(n9294), .Q(n16804) );
  OR2X1 U17470 ( .IN1(WX11025), .IN2(n3557), .Q(n16803) );
  OR2X1 U17471 ( .IN1(n16805), .IN2(n16806), .Q(n16802) );
  AND2X1 U17472 ( .IN1(n9295), .IN2(WX11217), .Q(n16806) );
  AND2X1 U17473 ( .IN1(n9557), .IN2(WX11153), .Q(n16805) );
  OR2X1 U17474 ( .IN1(n16807), .IN2(n16808), .Q(WX11022) );
  OR2X1 U17475 ( .IN1(n16809), .IN2(n16810), .Q(n16808) );
  AND2X1 U17476 ( .IN1(test_so99), .IN2(n10026), .Q(n16810) );
  AND2X1 U17477 ( .IN1(DATA_0_14), .IN2(n10063), .Q(n16809) );
  OR2X1 U17478 ( .IN1(n16811), .IN2(n16812), .Q(n16807) );
  AND2X1 U17479 ( .IN1(n1954), .IN2(n10010), .Q(n16812) );
  INVX0 U17480 ( .INP(n16813), .ZN(n1954) );
  OR2X1 U17481 ( .IN1(n10630), .IN2(n3800), .Q(n16813) );
  AND2X1 U17482 ( .IN1(n9985), .IN2(n11022), .Q(n16811) );
  OR2X1 U17483 ( .IN1(n16814), .IN2(n16815), .Q(n11022) );
  INVX0 U17484 ( .INP(n16816), .ZN(n16815) );
  OR2X1 U17485 ( .IN1(n16817), .IN2(n16818), .Q(n16816) );
  AND2X1 U17486 ( .IN1(n16818), .IN2(n16817), .Q(n16814) );
  AND2X1 U17487 ( .IN1(n16819), .IN2(n16820), .Q(n16817) );
  OR2X1 U17488 ( .IN1(WX11087), .IN2(n9296), .Q(n16820) );
  OR2X1 U17489 ( .IN1(WX11023), .IN2(n3559), .Q(n16819) );
  OR2X1 U17490 ( .IN1(n16821), .IN2(n16822), .Q(n16818) );
  AND2X1 U17491 ( .IN1(n9297), .IN2(WX11215), .Q(n16822) );
  AND2X1 U17492 ( .IN1(n9556), .IN2(WX11151), .Q(n16821) );
  OR2X1 U17493 ( .IN1(n16823), .IN2(n16824), .Q(WX11020) );
  OR2X1 U17494 ( .IN1(n16825), .IN2(n16826), .Q(n16824) );
  AND2X1 U17495 ( .IN1(n10036), .IN2(CRC_OUT_1_15), .Q(n16826) );
  AND2X1 U17496 ( .IN1(DATA_0_15), .IN2(n10063), .Q(n16825) );
  OR2X1 U17497 ( .IN1(n16827), .IN2(n16828), .Q(n16823) );
  AND2X1 U17498 ( .IN1(n1953), .IN2(n10010), .Q(n16828) );
  INVX0 U17499 ( .INP(n16829), .ZN(n1953) );
  OR2X1 U17500 ( .IN1(n10630), .IN2(n3801), .Q(n16829) );
  AND2X1 U17501 ( .IN1(n9985), .IN2(n11031), .Q(n16827) );
  OR2X1 U17502 ( .IN1(n16830), .IN2(n16831), .Q(n11031) );
  INVX0 U17503 ( .INP(n16832), .ZN(n16831) );
  OR2X1 U17504 ( .IN1(n16833), .IN2(n16834), .Q(n16832) );
  AND2X1 U17505 ( .IN1(n16834), .IN2(n16833), .Q(n16830) );
  AND2X1 U17506 ( .IN1(n16835), .IN2(n16836), .Q(n16833) );
  OR2X1 U17507 ( .IN1(WX11085), .IN2(n9298), .Q(n16836) );
  OR2X1 U17508 ( .IN1(WX11021), .IN2(n3561), .Q(n16835) );
  OR2X1 U17509 ( .IN1(n16837), .IN2(n16838), .Q(n16834) );
  AND2X1 U17510 ( .IN1(n9299), .IN2(WX11213), .Q(n16838) );
  AND2X1 U17511 ( .IN1(n9555), .IN2(WX11149), .Q(n16837) );
  OR2X1 U17512 ( .IN1(n16839), .IN2(n16840), .Q(WX11018) );
  OR2X1 U17513 ( .IN1(n16841), .IN2(n16842), .Q(n16840) );
  AND2X1 U17514 ( .IN1(n10036), .IN2(CRC_OUT_1_16), .Q(n16842) );
  AND2X1 U17515 ( .IN1(DATA_0_16), .IN2(n10062), .Q(n16841) );
  OR2X1 U17516 ( .IN1(n16843), .IN2(n16844), .Q(n16839) );
  AND2X1 U17517 ( .IN1(n1952), .IN2(n10010), .Q(n16844) );
  INVX0 U17518 ( .INP(n16845), .ZN(n1952) );
  OR2X1 U17519 ( .IN1(n10630), .IN2(n3802), .Q(n16845) );
  AND2X1 U17520 ( .IN1(n9985), .IN2(n11040), .Q(n16843) );
  OR2X1 U17521 ( .IN1(n16846), .IN2(n16847), .Q(n11040) );
  INVX0 U17522 ( .INP(n16848), .ZN(n16847) );
  OR2X1 U17523 ( .IN1(n16849), .IN2(n16850), .Q(n16848) );
  AND2X1 U17524 ( .IN1(n16850), .IN2(n16849), .Q(n16846) );
  INVX0 U17525 ( .INP(n16851), .ZN(n16849) );
  OR2X1 U17526 ( .IN1(n16852), .IN2(n16853), .Q(n16851) );
  AND2X1 U17527 ( .IN1(n10528), .IN2(n8246), .Q(n16853) );
  AND2X1 U17528 ( .IN1(n17987), .IN2(n10539), .Q(n16852) );
  OR2X1 U17529 ( .IN1(n16854), .IN2(n16855), .Q(n16850) );
  AND2X1 U17530 ( .IN1(n9512), .IN2(n16856), .Q(n16855) );
  AND2X1 U17531 ( .IN1(n16857), .IN2(n16858), .Q(n16856) );
  OR2X1 U17532 ( .IN1(n9044), .IN2(WX11147), .Q(n16858) );
  OR2X1 U17533 ( .IN1(n9045), .IN2(WX11083), .Q(n16857) );
  AND2X1 U17534 ( .IN1(n16859), .IN2(WX11211), .Q(n16854) );
  OR2X1 U17535 ( .IN1(n16860), .IN2(n16861), .Q(n16859) );
  AND2X1 U17536 ( .IN1(n9044), .IN2(WX11147), .Q(n16861) );
  AND2X1 U17537 ( .IN1(n9045), .IN2(WX11083), .Q(n16860) );
  OR2X1 U17538 ( .IN1(n16862), .IN2(n16863), .Q(WX11016) );
  OR2X1 U17539 ( .IN1(n16864), .IN2(n16865), .Q(n16863) );
  AND2X1 U17540 ( .IN1(n10036), .IN2(CRC_OUT_1_17), .Q(n16865) );
  AND2X1 U17541 ( .IN1(DATA_0_17), .IN2(n10063), .Q(n16864) );
  OR2X1 U17542 ( .IN1(n16866), .IN2(n16867), .Q(n16862) );
  AND2X1 U17543 ( .IN1(n1951), .IN2(n10010), .Q(n16867) );
  INVX0 U17544 ( .INP(n16868), .ZN(n1951) );
  OR2X1 U17545 ( .IN1(n10630), .IN2(n3803), .Q(n16868) );
  AND2X1 U17546 ( .IN1(n9985), .IN2(n11049), .Q(n16866) );
  OR2X1 U17547 ( .IN1(n16869), .IN2(n16870), .Q(n11049) );
  INVX0 U17548 ( .INP(n16871), .ZN(n16870) );
  OR2X1 U17549 ( .IN1(n16872), .IN2(n16873), .Q(n16871) );
  AND2X1 U17550 ( .IN1(n16873), .IN2(n16872), .Q(n16869) );
  INVX0 U17551 ( .INP(n16874), .ZN(n16872) );
  OR2X1 U17552 ( .IN1(n16875), .IN2(n16876), .Q(n16874) );
  AND2X1 U17553 ( .IN1(n10529), .IN2(n8247), .Q(n16876) );
  AND2X1 U17554 ( .IN1(n17988), .IN2(n10539), .Q(n16875) );
  OR2X1 U17555 ( .IN1(n16877), .IN2(n16878), .Q(n16873) );
  AND2X1 U17556 ( .IN1(n9554), .IN2(n16879), .Q(n16878) );
  AND2X1 U17557 ( .IN1(n16880), .IN2(n16881), .Q(n16879) );
  OR2X1 U17558 ( .IN1(n9046), .IN2(WX11145), .Q(n16881) );
  OR2X1 U17559 ( .IN1(n9047), .IN2(WX11081), .Q(n16880) );
  AND2X1 U17560 ( .IN1(n16882), .IN2(WX11209), .Q(n16877) );
  OR2X1 U17561 ( .IN1(n16883), .IN2(n16884), .Q(n16882) );
  AND2X1 U17562 ( .IN1(n9046), .IN2(WX11145), .Q(n16884) );
  AND2X1 U17563 ( .IN1(n9047), .IN2(WX11081), .Q(n16883) );
  OR2X1 U17564 ( .IN1(n16885), .IN2(n16886), .Q(WX11014) );
  OR2X1 U17565 ( .IN1(n16887), .IN2(n16888), .Q(n16886) );
  AND2X1 U17566 ( .IN1(n10036), .IN2(CRC_OUT_1_18), .Q(n16888) );
  AND2X1 U17567 ( .IN1(DATA_0_18), .IN2(n10061), .Q(n16887) );
  OR2X1 U17568 ( .IN1(n16889), .IN2(n16890), .Q(n16885) );
  AND2X1 U17569 ( .IN1(n1950), .IN2(n10010), .Q(n16890) );
  INVX0 U17570 ( .INP(n16891), .ZN(n1950) );
  OR2X1 U17571 ( .IN1(n10630), .IN2(n3804), .Q(n16891) );
  AND2X1 U17572 ( .IN1(n9985), .IN2(n11058), .Q(n16889) );
  OR2X1 U17573 ( .IN1(n16892), .IN2(n16893), .Q(n11058) );
  INVX0 U17574 ( .INP(n16894), .ZN(n16893) );
  OR2X1 U17575 ( .IN1(n16895), .IN2(n16896), .Q(n16894) );
  AND2X1 U17576 ( .IN1(n16896), .IN2(n16895), .Q(n16892) );
  INVX0 U17577 ( .INP(n16897), .ZN(n16895) );
  OR2X1 U17578 ( .IN1(n16898), .IN2(n16899), .Q(n16897) );
  AND2X1 U17579 ( .IN1(n10529), .IN2(n8248), .Q(n16899) );
  AND2X1 U17580 ( .IN1(n17989), .IN2(n10539), .Q(n16898) );
  OR2X1 U17581 ( .IN1(n16900), .IN2(n16901), .Q(n16896) );
  AND2X1 U17582 ( .IN1(n9553), .IN2(n16902), .Q(n16901) );
  AND2X1 U17583 ( .IN1(n16903), .IN2(n16904), .Q(n16902) );
  OR2X1 U17584 ( .IN1(n9048), .IN2(WX11143), .Q(n16904) );
  OR2X1 U17585 ( .IN1(n9049), .IN2(WX11079), .Q(n16903) );
  AND2X1 U17586 ( .IN1(n16905), .IN2(WX11207), .Q(n16900) );
  OR2X1 U17587 ( .IN1(n16906), .IN2(n16907), .Q(n16905) );
  AND2X1 U17588 ( .IN1(n9048), .IN2(WX11143), .Q(n16907) );
  AND2X1 U17589 ( .IN1(n9049), .IN2(WX11079), .Q(n16906) );
  OR2X1 U17590 ( .IN1(n16908), .IN2(n16909), .Q(WX11012) );
  OR2X1 U17591 ( .IN1(n16910), .IN2(n16911), .Q(n16909) );
  AND2X1 U17592 ( .IN1(n10036), .IN2(CRC_OUT_1_19), .Q(n16911) );
  AND2X1 U17593 ( .IN1(DATA_0_19), .IN2(n10060), .Q(n16910) );
  OR2X1 U17594 ( .IN1(n16912), .IN2(n16913), .Q(n16908) );
  AND2X1 U17595 ( .IN1(n1949), .IN2(n10010), .Q(n16913) );
  INVX0 U17596 ( .INP(n16914), .ZN(n1949) );
  OR2X1 U17597 ( .IN1(n10629), .IN2(n3805), .Q(n16914) );
  AND2X1 U17598 ( .IN1(n11067), .IN2(n9972), .Q(n16912) );
  AND2X1 U17599 ( .IN1(n16915), .IN2(n16916), .Q(n11067) );
  INVX0 U17600 ( .INP(n16917), .ZN(n16916) );
  AND2X1 U17601 ( .IN1(n16918), .IN2(n16919), .Q(n16917) );
  OR2X1 U17602 ( .IN1(n16919), .IN2(n16918), .Q(n16915) );
  OR2X1 U17603 ( .IN1(n16920), .IN2(n16921), .Q(n16918) );
  AND2X1 U17604 ( .IN1(n10529), .IN2(WX11077), .Q(n16921) );
  AND2X1 U17605 ( .IN1(n9050), .IN2(n10539), .Q(n16920) );
  AND2X1 U17606 ( .IN1(n16922), .IN2(n16923), .Q(n16919) );
  INVX0 U17607 ( .INP(n16924), .ZN(n16923) );
  AND2X1 U17608 ( .IN1(n16925), .IN2(WX11141), .Q(n16924) );
  OR2X1 U17609 ( .IN1(WX11141), .IN2(n16925), .Q(n16922) );
  OR2X1 U17610 ( .IN1(n16926), .IN2(n16927), .Q(n16925) );
  AND2X1 U17611 ( .IN1(n17990), .IN2(n9913), .Q(n16927) );
  AND2X1 U17612 ( .IN1(test_so97), .IN2(n8249), .Q(n16926) );
  OR2X1 U17613 ( .IN1(n16928), .IN2(n16929), .Q(WX11010) );
  OR2X1 U17614 ( .IN1(n16930), .IN2(n16931), .Q(n16929) );
  AND2X1 U17615 ( .IN1(n10036), .IN2(CRC_OUT_1_20), .Q(n16931) );
  AND2X1 U17616 ( .IN1(DATA_0_20), .IN2(n10063), .Q(n16930) );
  OR2X1 U17617 ( .IN1(n16932), .IN2(n16933), .Q(n16928) );
  AND2X1 U17618 ( .IN1(n1948), .IN2(n10010), .Q(n16933) );
  INVX0 U17619 ( .INP(n16934), .ZN(n1948) );
  OR2X1 U17620 ( .IN1(n10629), .IN2(n3806), .Q(n16934) );
  AND2X1 U17621 ( .IN1(n9985), .IN2(n11076), .Q(n16932) );
  OR2X1 U17622 ( .IN1(n16935), .IN2(n16936), .Q(n11076) );
  INVX0 U17623 ( .INP(n16937), .ZN(n16936) );
  OR2X1 U17624 ( .IN1(n16938), .IN2(n16939), .Q(n16937) );
  AND2X1 U17625 ( .IN1(n16939), .IN2(n16938), .Q(n16935) );
  INVX0 U17626 ( .INP(n16940), .ZN(n16938) );
  OR2X1 U17627 ( .IN1(n16941), .IN2(n16942), .Q(n16940) );
  AND2X1 U17628 ( .IN1(n10529), .IN2(n8250), .Q(n16942) );
  AND2X1 U17629 ( .IN1(n17991), .IN2(n10538), .Q(n16941) );
  OR2X1 U17630 ( .IN1(n16943), .IN2(n16944), .Q(n16939) );
  AND2X1 U17631 ( .IN1(n9552), .IN2(n16945), .Q(n16944) );
  AND2X1 U17632 ( .IN1(n16946), .IN2(n16947), .Q(n16945) );
  OR2X1 U17633 ( .IN1(n9052), .IN2(WX11139), .Q(n16947) );
  OR2X1 U17634 ( .IN1(n9053), .IN2(WX11075), .Q(n16946) );
  AND2X1 U17635 ( .IN1(n16948), .IN2(WX11203), .Q(n16943) );
  OR2X1 U17636 ( .IN1(n16949), .IN2(n16950), .Q(n16948) );
  AND2X1 U17637 ( .IN1(n9052), .IN2(WX11139), .Q(n16950) );
  AND2X1 U17638 ( .IN1(n9053), .IN2(WX11075), .Q(n16949) );
  OR2X1 U17639 ( .IN1(n16951), .IN2(n16952), .Q(WX11008) );
  OR2X1 U17640 ( .IN1(n16953), .IN2(n16954), .Q(n16952) );
  AND2X1 U17641 ( .IN1(n10036), .IN2(CRC_OUT_1_21), .Q(n16954) );
  AND2X1 U17642 ( .IN1(DATA_0_21), .IN2(n10061), .Q(n16953) );
  OR2X1 U17643 ( .IN1(n16955), .IN2(n16956), .Q(n16951) );
  AND2X1 U17644 ( .IN1(n1947), .IN2(n10010), .Q(n16956) );
  INVX0 U17645 ( .INP(n16957), .ZN(n1947) );
  OR2X1 U17646 ( .IN1(n10629), .IN2(n3807), .Q(n16957) );
  AND2X1 U17647 ( .IN1(n11085), .IN2(n9972), .Q(n16955) );
  AND2X1 U17648 ( .IN1(n16958), .IN2(n16959), .Q(n11085) );
  INVX0 U17649 ( .INP(n16960), .ZN(n16959) );
  AND2X1 U17650 ( .IN1(n16961), .IN2(n16962), .Q(n16960) );
  OR2X1 U17651 ( .IN1(n16962), .IN2(n16961), .Q(n16958) );
  OR2X1 U17652 ( .IN1(n16963), .IN2(n16964), .Q(n16961) );
  AND2X1 U17653 ( .IN1(n10529), .IN2(WX11073), .Q(n16964) );
  AND2X1 U17654 ( .IN1(n9054), .IN2(n10538), .Q(n16963) );
  AND2X1 U17655 ( .IN1(n16965), .IN2(n16966), .Q(n16962) );
  OR2X1 U17656 ( .IN1(n16967), .IN2(n9551), .Q(n16966) );
  INVX0 U17657 ( .INP(n16968), .ZN(n16967) );
  OR2X1 U17658 ( .IN1(WX11201), .IN2(n16968), .Q(n16965) );
  OR2X1 U17659 ( .IN1(n16969), .IN2(n16970), .Q(n16968) );
  AND2X1 U17660 ( .IN1(n17992), .IN2(n9965), .Q(n16970) );
  AND2X1 U17661 ( .IN1(test_so95), .IN2(n8251), .Q(n16969) );
  OR2X1 U17662 ( .IN1(n16971), .IN2(n16972), .Q(WX11006) );
  OR2X1 U17663 ( .IN1(n16973), .IN2(n16974), .Q(n16972) );
  AND2X1 U17664 ( .IN1(n10036), .IN2(CRC_OUT_1_22), .Q(n16974) );
  AND2X1 U17665 ( .IN1(DATA_0_22), .IN2(n10062), .Q(n16973) );
  OR2X1 U17666 ( .IN1(n16975), .IN2(n16976), .Q(n16971) );
  AND2X1 U17667 ( .IN1(n1946), .IN2(n10011), .Q(n16976) );
  INVX0 U17668 ( .INP(n16977), .ZN(n1946) );
  OR2X1 U17669 ( .IN1(n10629), .IN2(n3808), .Q(n16977) );
  AND2X1 U17670 ( .IN1(n9985), .IN2(n11094), .Q(n16975) );
  OR2X1 U17671 ( .IN1(n16978), .IN2(n16979), .Q(n11094) );
  INVX0 U17672 ( .INP(n16980), .ZN(n16979) );
  OR2X1 U17673 ( .IN1(n16981), .IN2(n16982), .Q(n16980) );
  AND2X1 U17674 ( .IN1(n16982), .IN2(n16981), .Q(n16978) );
  INVX0 U17675 ( .INP(n16983), .ZN(n16981) );
  OR2X1 U17676 ( .IN1(n16984), .IN2(n16985), .Q(n16983) );
  AND2X1 U17677 ( .IN1(n10529), .IN2(n8252), .Q(n16985) );
  AND2X1 U17678 ( .IN1(n17993), .IN2(n10538), .Q(n16984) );
  OR2X1 U17679 ( .IN1(n16986), .IN2(n16987), .Q(n16982) );
  AND2X1 U17680 ( .IN1(n9550), .IN2(n16988), .Q(n16987) );
  AND2X1 U17681 ( .IN1(n16989), .IN2(n16990), .Q(n16988) );
  OR2X1 U17682 ( .IN1(n9055), .IN2(WX11135), .Q(n16990) );
  OR2X1 U17683 ( .IN1(n9056), .IN2(WX11071), .Q(n16989) );
  AND2X1 U17684 ( .IN1(n16991), .IN2(WX11199), .Q(n16986) );
  OR2X1 U17685 ( .IN1(n16992), .IN2(n16993), .Q(n16991) );
  AND2X1 U17686 ( .IN1(n9055), .IN2(WX11135), .Q(n16993) );
  AND2X1 U17687 ( .IN1(n9056), .IN2(WX11071), .Q(n16992) );
  OR2X1 U17688 ( .IN1(n16994), .IN2(n16995), .Q(WX11004) );
  OR2X1 U17689 ( .IN1(n16996), .IN2(n16997), .Q(n16995) );
  AND2X1 U17690 ( .IN1(n10036), .IN2(CRC_OUT_1_23), .Q(n16997) );
  AND2X1 U17691 ( .IN1(DATA_0_23), .IN2(n10060), .Q(n16996) );
  OR2X1 U17692 ( .IN1(n16998), .IN2(n16999), .Q(n16994) );
  AND2X1 U17693 ( .IN1(n1945), .IN2(n10011), .Q(n16999) );
  INVX0 U17694 ( .INP(n17000), .ZN(n1945) );
  OR2X1 U17695 ( .IN1(n10629), .IN2(n3809), .Q(n17000) );
  AND2X1 U17696 ( .IN1(n11103), .IN2(n9972), .Q(n16998) );
  AND2X1 U17697 ( .IN1(n17001), .IN2(n17002), .Q(n11103) );
  INVX0 U17698 ( .INP(n17003), .ZN(n17002) );
  AND2X1 U17699 ( .IN1(n17004), .IN2(n17005), .Q(n17003) );
  OR2X1 U17700 ( .IN1(n17005), .IN2(n17004), .Q(n17001) );
  OR2X1 U17701 ( .IN1(n17006), .IN2(n17007), .Q(n17004) );
  AND2X1 U17702 ( .IN1(n10529), .IN2(WX11133), .Q(n17007) );
  AND2X1 U17703 ( .IN1(n9057), .IN2(n10538), .Q(n17006) );
  AND2X1 U17704 ( .IN1(n17008), .IN2(n17009), .Q(n17005) );
  OR2X1 U17705 ( .IN1(n17010), .IN2(n9549), .Q(n17009) );
  INVX0 U17706 ( .INP(n17011), .ZN(n17010) );
  OR2X1 U17707 ( .IN1(WX11197), .IN2(n17011), .Q(n17008) );
  OR2X1 U17708 ( .IN1(n17012), .IN2(n17013), .Q(n17011) );
  AND2X1 U17709 ( .IN1(n17994), .IN2(n9966), .Q(n17013) );
  AND2X1 U17710 ( .IN1(test_so93), .IN2(n8253), .Q(n17012) );
  OR2X1 U17711 ( .IN1(n17014), .IN2(n17015), .Q(WX11002) );
  OR2X1 U17712 ( .IN1(n17016), .IN2(n17017), .Q(n17015) );
  AND2X1 U17713 ( .IN1(n10037), .IN2(CRC_OUT_1_24), .Q(n17017) );
  AND2X1 U17714 ( .IN1(DATA_0_24), .IN2(n10061), .Q(n17016) );
  OR2X1 U17715 ( .IN1(n17018), .IN2(n17019), .Q(n17014) );
  AND2X1 U17716 ( .IN1(n1944), .IN2(n10011), .Q(n17019) );
  INVX0 U17717 ( .INP(n17020), .ZN(n1944) );
  OR2X1 U17718 ( .IN1(n10629), .IN2(n3810), .Q(n17020) );
  AND2X1 U17719 ( .IN1(n9985), .IN2(n11112), .Q(n17018) );
  OR2X1 U17720 ( .IN1(n17021), .IN2(n17022), .Q(n11112) );
  INVX0 U17721 ( .INP(n17023), .ZN(n17022) );
  OR2X1 U17722 ( .IN1(n17024), .IN2(n17025), .Q(n17023) );
  AND2X1 U17723 ( .IN1(n17025), .IN2(n17024), .Q(n17021) );
  INVX0 U17724 ( .INP(n17026), .ZN(n17024) );
  OR2X1 U17725 ( .IN1(n17027), .IN2(n17028), .Q(n17026) );
  AND2X1 U17726 ( .IN1(n10529), .IN2(n8254), .Q(n17028) );
  AND2X1 U17727 ( .IN1(n17995), .IN2(n10538), .Q(n17027) );
  OR2X1 U17728 ( .IN1(n17029), .IN2(n17030), .Q(n17025) );
  AND2X1 U17729 ( .IN1(n9548), .IN2(n17031), .Q(n17030) );
  AND2X1 U17730 ( .IN1(n17032), .IN2(n17033), .Q(n17031) );
  OR2X1 U17731 ( .IN1(n9058), .IN2(WX11131), .Q(n17033) );
  OR2X1 U17732 ( .IN1(n9059), .IN2(WX11067), .Q(n17032) );
  AND2X1 U17733 ( .IN1(n17034), .IN2(WX11195), .Q(n17029) );
  OR2X1 U17734 ( .IN1(n17035), .IN2(n17036), .Q(n17034) );
  AND2X1 U17735 ( .IN1(n9058), .IN2(WX11131), .Q(n17036) );
  AND2X1 U17736 ( .IN1(n9059), .IN2(WX11067), .Q(n17035) );
  OR2X1 U17737 ( .IN1(n17037), .IN2(n17038), .Q(WX11000) );
  OR2X1 U17738 ( .IN1(n17039), .IN2(n17040), .Q(n17038) );
  AND2X1 U17739 ( .IN1(n10037), .IN2(CRC_OUT_1_25), .Q(n17040) );
  AND2X1 U17740 ( .IN1(DATA_0_25), .IN2(n10062), .Q(n17039) );
  OR2X1 U17741 ( .IN1(n17041), .IN2(n17042), .Q(n17037) );
  AND2X1 U17742 ( .IN1(n1943), .IN2(n10011), .Q(n17042) );
  INVX0 U17743 ( .INP(n17043), .ZN(n1943) );
  OR2X1 U17744 ( .IN1(n10629), .IN2(n3811), .Q(n17043) );
  AND2X1 U17745 ( .IN1(n11121), .IN2(n9972), .Q(n17041) );
  AND2X1 U17746 ( .IN1(n17044), .IN2(n17045), .Q(n11121) );
  OR2X1 U17747 ( .IN1(n17046), .IN2(n17047), .Q(n17045) );
  INVX0 U17748 ( .INP(n17048), .ZN(n17046) );
  OR2X1 U17749 ( .IN1(n17049), .IN2(n17048), .Q(n17044) );
  OR2X1 U17750 ( .IN1(n17050), .IN2(n17051), .Q(n17048) );
  AND2X1 U17751 ( .IN1(n10529), .IN2(WX11193), .Q(n17051) );
  AND2X1 U17752 ( .IN1(n9547), .IN2(n10538), .Q(n17050) );
  INVX0 U17753 ( .INP(n17047), .ZN(n17049) );
  OR2X1 U17754 ( .IN1(n17052), .IN2(n17053), .Q(n17047) );
  AND2X1 U17755 ( .IN1(n9061), .IN2(n17054), .Q(n17053) );
  AND2X1 U17756 ( .IN1(n17055), .IN2(n17056), .Q(n17054) );
  OR2X1 U17757 ( .IN1(n9060), .IN2(n9896), .Q(n17056) );
  OR2X1 U17758 ( .IN1(test_so91), .IN2(WX11065), .Q(n17055) );
  AND2X1 U17759 ( .IN1(n17057), .IN2(WX11129), .Q(n17052) );
  OR2X1 U17760 ( .IN1(n17058), .IN2(n17059), .Q(n17057) );
  AND2X1 U17761 ( .IN1(n9060), .IN2(n9896), .Q(n17059) );
  AND2X1 U17762 ( .IN1(test_so91), .IN2(WX11065), .Q(n17058) );
  OR2X1 U17763 ( .IN1(n17060), .IN2(n17061), .Q(WX10998) );
  OR2X1 U17764 ( .IN1(n17062), .IN2(n17063), .Q(n17061) );
  AND2X1 U17765 ( .IN1(n10037), .IN2(CRC_OUT_1_26), .Q(n17063) );
  AND2X1 U17766 ( .IN1(DATA_0_26), .IN2(n10062), .Q(n17062) );
  OR2X1 U17767 ( .IN1(n17064), .IN2(n17065), .Q(n17060) );
  AND2X1 U17768 ( .IN1(n1942), .IN2(n10011), .Q(n17065) );
  INVX0 U17769 ( .INP(n17066), .ZN(n1942) );
  OR2X1 U17770 ( .IN1(n10629), .IN2(n3812), .Q(n17066) );
  AND2X1 U17771 ( .IN1(n9985), .IN2(n11130), .Q(n17064) );
  OR2X1 U17772 ( .IN1(n17067), .IN2(n17068), .Q(n11130) );
  INVX0 U17773 ( .INP(n17069), .ZN(n17068) );
  OR2X1 U17774 ( .IN1(n17070), .IN2(n17071), .Q(n17069) );
  AND2X1 U17775 ( .IN1(n17071), .IN2(n17070), .Q(n17067) );
  INVX0 U17776 ( .INP(n17072), .ZN(n17070) );
  OR2X1 U17777 ( .IN1(n17073), .IN2(n17074), .Q(n17072) );
  AND2X1 U17778 ( .IN1(n10529), .IN2(n8257), .Q(n17074) );
  AND2X1 U17779 ( .IN1(n17996), .IN2(n10538), .Q(n17073) );
  OR2X1 U17780 ( .IN1(n17075), .IN2(n17076), .Q(n17071) );
  AND2X1 U17781 ( .IN1(n9546), .IN2(n17077), .Q(n17076) );
  AND2X1 U17782 ( .IN1(n17078), .IN2(n17079), .Q(n17077) );
  OR2X1 U17783 ( .IN1(n9062), .IN2(WX11127), .Q(n17079) );
  OR2X1 U17784 ( .IN1(n9063), .IN2(WX11063), .Q(n17078) );
  AND2X1 U17785 ( .IN1(n17080), .IN2(WX11191), .Q(n17075) );
  OR2X1 U17786 ( .IN1(n17081), .IN2(n17082), .Q(n17080) );
  AND2X1 U17787 ( .IN1(n9062), .IN2(WX11127), .Q(n17082) );
  AND2X1 U17788 ( .IN1(n9063), .IN2(WX11063), .Q(n17081) );
  OR2X1 U17789 ( .IN1(n17083), .IN2(n17084), .Q(WX10996) );
  OR2X1 U17790 ( .IN1(n17085), .IN2(n17086), .Q(n17084) );
  AND2X1 U17791 ( .IN1(n10037), .IN2(CRC_OUT_1_27), .Q(n17086) );
  AND2X1 U17792 ( .IN1(DATA_0_27), .IN2(n10061), .Q(n17085) );
  OR2X1 U17793 ( .IN1(n17087), .IN2(n17088), .Q(n17083) );
  AND2X1 U17794 ( .IN1(n1941), .IN2(n10011), .Q(n17088) );
  INVX0 U17795 ( .INP(n17089), .ZN(n1941) );
  OR2X1 U17796 ( .IN1(n10629), .IN2(n3813), .Q(n17089) );
  AND2X1 U17797 ( .IN1(n9985), .IN2(n11139), .Q(n17087) );
  OR2X1 U17798 ( .IN1(n17090), .IN2(n17091), .Q(n11139) );
  INVX0 U17799 ( .INP(n17092), .ZN(n17091) );
  OR2X1 U17800 ( .IN1(n17093), .IN2(n17094), .Q(n17092) );
  AND2X1 U17801 ( .IN1(n17094), .IN2(n17093), .Q(n17090) );
  INVX0 U17802 ( .INP(n17095), .ZN(n17093) );
  OR2X1 U17803 ( .IN1(n17096), .IN2(n17097), .Q(n17095) );
  AND2X1 U17804 ( .IN1(n10530), .IN2(n8258), .Q(n17097) );
  AND2X1 U17805 ( .IN1(n17997), .IN2(n10538), .Q(n17096) );
  OR2X1 U17806 ( .IN1(n17098), .IN2(n17099), .Q(n17094) );
  AND2X1 U17807 ( .IN1(n9545), .IN2(n17100), .Q(n17099) );
  AND2X1 U17808 ( .IN1(n17101), .IN2(n17102), .Q(n17100) );
  OR2X1 U17809 ( .IN1(n9064), .IN2(WX11125), .Q(n17102) );
  OR2X1 U17810 ( .IN1(n9065), .IN2(WX11061), .Q(n17101) );
  AND2X1 U17811 ( .IN1(n17103), .IN2(WX11189), .Q(n17098) );
  OR2X1 U17812 ( .IN1(n17104), .IN2(n17105), .Q(n17103) );
  AND2X1 U17813 ( .IN1(n9064), .IN2(WX11125), .Q(n17105) );
  AND2X1 U17814 ( .IN1(n9065), .IN2(WX11061), .Q(n17104) );
  OR2X1 U17815 ( .IN1(n17106), .IN2(n17107), .Q(WX10994) );
  OR2X1 U17816 ( .IN1(n17108), .IN2(n17109), .Q(n17107) );
  AND2X1 U17817 ( .IN1(n10037), .IN2(CRC_OUT_1_28), .Q(n17109) );
  AND2X1 U17818 ( .IN1(DATA_0_28), .IN2(n10060), .Q(n17108) );
  OR2X1 U17819 ( .IN1(n17110), .IN2(n17111), .Q(n17106) );
  AND2X1 U17820 ( .IN1(n1940), .IN2(n10011), .Q(n17111) );
  INVX0 U17821 ( .INP(n17112), .ZN(n1940) );
  OR2X1 U17822 ( .IN1(n10629), .IN2(n3814), .Q(n17112) );
  AND2X1 U17823 ( .IN1(n9985), .IN2(n11148), .Q(n17110) );
  OR2X1 U17824 ( .IN1(n17113), .IN2(n17114), .Q(n11148) );
  INVX0 U17825 ( .INP(n17115), .ZN(n17114) );
  OR2X1 U17826 ( .IN1(n17116), .IN2(n17117), .Q(n17115) );
  AND2X1 U17827 ( .IN1(n17117), .IN2(n17116), .Q(n17113) );
  INVX0 U17828 ( .INP(n17118), .ZN(n17116) );
  OR2X1 U17829 ( .IN1(n17119), .IN2(n17120), .Q(n17118) );
  AND2X1 U17830 ( .IN1(n10530), .IN2(n8259), .Q(n17120) );
  AND2X1 U17831 ( .IN1(n17998), .IN2(n10538), .Q(n17119) );
  OR2X1 U17832 ( .IN1(n17121), .IN2(n17122), .Q(n17117) );
  AND2X1 U17833 ( .IN1(n9544), .IN2(n17123), .Q(n17122) );
  AND2X1 U17834 ( .IN1(n17124), .IN2(n17125), .Q(n17123) );
  OR2X1 U17835 ( .IN1(n9066), .IN2(WX11123), .Q(n17125) );
  OR2X1 U17836 ( .IN1(n9067), .IN2(WX11059), .Q(n17124) );
  AND2X1 U17837 ( .IN1(n17126), .IN2(WX11187), .Q(n17121) );
  OR2X1 U17838 ( .IN1(n17127), .IN2(n17128), .Q(n17126) );
  AND2X1 U17839 ( .IN1(n9066), .IN2(WX11123), .Q(n17128) );
  AND2X1 U17840 ( .IN1(n9067), .IN2(WX11059), .Q(n17127) );
  OR2X1 U17841 ( .IN1(n17129), .IN2(n17130), .Q(WX10992) );
  OR2X1 U17842 ( .IN1(n17131), .IN2(n17132), .Q(n17130) );
  AND2X1 U17843 ( .IN1(n10037), .IN2(CRC_OUT_1_29), .Q(n17132) );
  AND2X1 U17844 ( .IN1(DATA_0_29), .IN2(n10060), .Q(n17131) );
  OR2X1 U17845 ( .IN1(n17133), .IN2(n17134), .Q(n17129) );
  AND2X1 U17846 ( .IN1(n1939), .IN2(n10000), .Q(n17134) );
  INVX0 U17847 ( .INP(n17135), .ZN(n1939) );
  OR2X1 U17848 ( .IN1(n10629), .IN2(n3815), .Q(n17135) );
  AND2X1 U17849 ( .IN1(n9984), .IN2(n11157), .Q(n17133) );
  OR2X1 U17850 ( .IN1(n17136), .IN2(n17137), .Q(n11157) );
  INVX0 U17851 ( .INP(n17138), .ZN(n17137) );
  OR2X1 U17852 ( .IN1(n17139), .IN2(n17140), .Q(n17138) );
  AND2X1 U17853 ( .IN1(n17140), .IN2(n17139), .Q(n17136) );
  INVX0 U17854 ( .INP(n17141), .ZN(n17139) );
  OR2X1 U17855 ( .IN1(n17142), .IN2(n17143), .Q(n17141) );
  AND2X1 U17856 ( .IN1(n10530), .IN2(n8260), .Q(n17143) );
  AND2X1 U17857 ( .IN1(n17999), .IN2(n10538), .Q(n17142) );
  OR2X1 U17858 ( .IN1(n17144), .IN2(n17145), .Q(n17140) );
  AND2X1 U17859 ( .IN1(n9543), .IN2(n17146), .Q(n17145) );
  AND2X1 U17860 ( .IN1(n17147), .IN2(n17148), .Q(n17146) );
  OR2X1 U17861 ( .IN1(n9068), .IN2(WX11121), .Q(n17148) );
  OR2X1 U17862 ( .IN1(n9069), .IN2(WX11057), .Q(n17147) );
  AND2X1 U17863 ( .IN1(n17149), .IN2(WX11185), .Q(n17144) );
  OR2X1 U17864 ( .IN1(n17150), .IN2(n17151), .Q(n17149) );
  AND2X1 U17865 ( .IN1(n9068), .IN2(WX11121), .Q(n17151) );
  AND2X1 U17866 ( .IN1(n9069), .IN2(WX11057), .Q(n17150) );
  OR2X1 U17867 ( .IN1(n17152), .IN2(n17153), .Q(WX10990) );
  OR2X1 U17868 ( .IN1(n17154), .IN2(n17155), .Q(n17153) );
  AND2X1 U17869 ( .IN1(n10037), .IN2(CRC_OUT_1_30), .Q(n17155) );
  AND2X1 U17870 ( .IN1(DATA_0_30), .IN2(n10060), .Q(n17154) );
  OR2X1 U17871 ( .IN1(n17156), .IN2(n17157), .Q(n17152) );
  AND2X1 U17872 ( .IN1(n1938), .IN2(n10011), .Q(n17157) );
  AND2X1 U17873 ( .IN1(TM0), .IN2(n10514), .Q(n2148) );
  INVX0 U17874 ( .INP(n17158), .ZN(n1938) );
  OR2X1 U17875 ( .IN1(n10629), .IN2(n3816), .Q(n17158) );
  AND2X1 U17876 ( .IN1(n9989), .IN2(n11166), .Q(n17156) );
  OR2X1 U17877 ( .IN1(n17159), .IN2(n17160), .Q(n11166) );
  INVX0 U17878 ( .INP(n17161), .ZN(n17160) );
  OR2X1 U17879 ( .IN1(n17162), .IN2(n17163), .Q(n17161) );
  AND2X1 U17880 ( .IN1(n17163), .IN2(n17162), .Q(n17159) );
  INVX0 U17881 ( .INP(n17164), .ZN(n17162) );
  OR2X1 U17882 ( .IN1(n17165), .IN2(n17166), .Q(n17164) );
  AND2X1 U17883 ( .IN1(n10530), .IN2(n8261), .Q(n17166) );
  AND2X1 U17884 ( .IN1(n18000), .IN2(n10538), .Q(n17165) );
  OR2X1 U17885 ( .IN1(n17167), .IN2(n17168), .Q(n17163) );
  AND2X1 U17886 ( .IN1(n9542), .IN2(n17169), .Q(n17168) );
  AND2X1 U17887 ( .IN1(n17170), .IN2(n17171), .Q(n17169) );
  OR2X1 U17888 ( .IN1(n9070), .IN2(WX11119), .Q(n17171) );
  OR2X1 U17889 ( .IN1(n9071), .IN2(WX11055), .Q(n17170) );
  AND2X1 U17890 ( .IN1(n17172), .IN2(WX11183), .Q(n17167) );
  OR2X1 U17891 ( .IN1(n17173), .IN2(n17174), .Q(n17172) );
  AND2X1 U17892 ( .IN1(n9070), .IN2(WX11119), .Q(n17174) );
  AND2X1 U17893 ( .IN1(n9071), .IN2(WX11055), .Q(n17173) );
  OR2X1 U17894 ( .IN1(n17175), .IN2(n17176), .Q(WX10988) );
  OR2X1 U17895 ( .IN1(n17177), .IN2(n17178), .Q(n17176) );
  AND2X1 U17896 ( .IN1(n2245), .IN2(WX10829), .Q(n17178) );
  AND2X1 U17897 ( .IN1(test_so100), .IN2(n10027), .Q(n17177) );
  OR2X1 U17898 ( .IN1(n17179), .IN2(n17180), .Q(n17175) );
  AND2X1 U17899 ( .IN1(DATA_0_31), .IN2(n10058), .Q(n17180) );
  AND2X1 U17900 ( .IN1(n9978), .IN2(n11174), .Q(n17179) );
  OR2X1 U17901 ( .IN1(n17181), .IN2(n17182), .Q(n11174) );
  INVX0 U17902 ( .INP(n17183), .ZN(n17182) );
  OR2X1 U17903 ( .IN1(n17184), .IN2(n17185), .Q(n17183) );
  AND2X1 U17904 ( .IN1(n17185), .IN2(n17184), .Q(n17181) );
  INVX0 U17905 ( .INP(n17186), .ZN(n17184) );
  OR2X1 U17906 ( .IN1(n17187), .IN2(n17188), .Q(n17186) );
  AND2X1 U17907 ( .IN1(n10530), .IN2(n8262), .Q(n17188) );
  AND2X1 U17908 ( .IN1(n18001), .IN2(n10538), .Q(n17187) );
  OR2X1 U17909 ( .IN1(n17189), .IN2(n17190), .Q(n17185) );
  AND2X1 U17910 ( .IN1(n9541), .IN2(n17191), .Q(n17190) );
  AND2X1 U17911 ( .IN1(n17192), .IN2(n17193), .Q(n17191) );
  OR2X1 U17912 ( .IN1(n9028), .IN2(WX11117), .Q(n17193) );
  OR2X1 U17913 ( .IN1(n9029), .IN2(WX11053), .Q(n17192) );
  AND2X1 U17914 ( .IN1(n17194), .IN2(WX11181), .Q(n17189) );
  OR2X1 U17915 ( .IN1(n17195), .IN2(n17196), .Q(n17194) );
  AND2X1 U17916 ( .IN1(n9028), .IN2(WX11117), .Q(n17196) );
  AND2X1 U17917 ( .IN1(n9029), .IN2(WX11053), .Q(n17195) );
  AND2X1 U17918 ( .IN1(n10517), .IN2(n17197), .Q(n10896) );
  AND2X1 U17919 ( .IN1(n2182), .IN2(n10579), .Q(n17197) );
  AND2X1 U17920 ( .IN1(n9851), .IN2(n10580), .Q(WX10890) );
  AND2X1 U17921 ( .IN1(n17198), .IN2(n10580), .Q(WX10377) );
  OR2X1 U17922 ( .IN1(n17199), .IN2(n17200), .Q(n17198) );
  AND2X1 U17923 ( .IN1(DFF_1534_n1), .IN2(n9914), .Q(n17200) );
  AND2X1 U17924 ( .IN1(test_so85), .IN2(CRC_OUT_2_30), .Q(n17199) );
  AND2X1 U17925 ( .IN1(n17201), .IN2(n10580), .Q(WX10375) );
  AND2X1 U17926 ( .IN1(n17202), .IN2(n17203), .Q(n17201) );
  OR2X1 U17927 ( .IN1(DFF_1533_n1), .IN2(WX9890), .Q(n17203) );
  OR2X1 U17928 ( .IN1(n9567), .IN2(CRC_OUT_2_29), .Q(n17202) );
  AND2X1 U17929 ( .IN1(n17204), .IN2(n10580), .Q(WX10373) );
  AND2X1 U17930 ( .IN1(n17205), .IN2(n17206), .Q(n17204) );
  OR2X1 U17931 ( .IN1(DFF_1532_n1), .IN2(WX9892), .Q(n17206) );
  OR2X1 U17932 ( .IN1(n9568), .IN2(CRC_OUT_2_28), .Q(n17205) );
  AND2X1 U17933 ( .IN1(n17207), .IN2(n10580), .Q(WX10371) );
  AND2X1 U17934 ( .IN1(n17208), .IN2(n17209), .Q(n17207) );
  OR2X1 U17935 ( .IN1(DFF_1531_n1), .IN2(WX9894), .Q(n17209) );
  OR2X1 U17936 ( .IN1(n9569), .IN2(CRC_OUT_2_27), .Q(n17208) );
  AND2X1 U17937 ( .IN1(n17210), .IN2(n10580), .Q(WX10369) );
  AND2X1 U17938 ( .IN1(n17211), .IN2(n17212), .Q(n17210) );
  OR2X1 U17939 ( .IN1(DFF_1530_n1), .IN2(WX9896), .Q(n17212) );
  OR2X1 U17940 ( .IN1(n9570), .IN2(CRC_OUT_2_26), .Q(n17211) );
  AND2X1 U17941 ( .IN1(n17213), .IN2(n10580), .Q(WX10367) );
  AND2X1 U17942 ( .IN1(n17214), .IN2(n17215), .Q(n17213) );
  OR2X1 U17943 ( .IN1(DFF_1529_n1), .IN2(WX9898), .Q(n17215) );
  OR2X1 U17944 ( .IN1(n9571), .IN2(CRC_OUT_2_25), .Q(n17214) );
  AND2X1 U17945 ( .IN1(n17216), .IN2(n10580), .Q(WX10365) );
  AND2X1 U17946 ( .IN1(n17217), .IN2(n17218), .Q(n17216) );
  OR2X1 U17947 ( .IN1(DFF_1528_n1), .IN2(WX9900), .Q(n17218) );
  OR2X1 U17948 ( .IN1(n9572), .IN2(CRC_OUT_2_24), .Q(n17217) );
  AND2X1 U17949 ( .IN1(n17219), .IN2(n10580), .Q(WX10363) );
  AND2X1 U17950 ( .IN1(n17220), .IN2(n17221), .Q(n17219) );
  OR2X1 U17951 ( .IN1(DFF_1527_n1), .IN2(WX9902), .Q(n17221) );
  OR2X1 U17952 ( .IN1(n9573), .IN2(CRC_OUT_2_23), .Q(n17220) );
  AND2X1 U17953 ( .IN1(n17222), .IN2(n10581), .Q(WX10361) );
  AND2X1 U17954 ( .IN1(n17223), .IN2(n17224), .Q(n17222) );
  OR2X1 U17955 ( .IN1(DFF_1526_n1), .IN2(WX9904), .Q(n17224) );
  OR2X1 U17956 ( .IN1(n9574), .IN2(CRC_OUT_2_22), .Q(n17223) );
  AND2X1 U17957 ( .IN1(n17225), .IN2(n10581), .Q(WX10359) );
  AND2X1 U17958 ( .IN1(n17226), .IN2(n17227), .Q(n17225) );
  OR2X1 U17959 ( .IN1(DFF_1525_n1), .IN2(WX9906), .Q(n17227) );
  OR2X1 U17960 ( .IN1(n9575), .IN2(CRC_OUT_2_21), .Q(n17226) );
  AND2X1 U17961 ( .IN1(n17228), .IN2(n10581), .Q(WX10357) );
  AND2X1 U17962 ( .IN1(n17229), .IN2(n17230), .Q(n17228) );
  OR2X1 U17963 ( .IN1(DFF_1524_n1), .IN2(WX9908), .Q(n17230) );
  OR2X1 U17964 ( .IN1(n9576), .IN2(CRC_OUT_2_20), .Q(n17229) );
  AND2X1 U17965 ( .IN1(n17231), .IN2(n10581), .Q(WX10355) );
  OR2X1 U17966 ( .IN1(n17232), .IN2(n17233), .Q(n17231) );
  AND2X1 U17967 ( .IN1(n9577), .IN2(n9951), .Q(n17233) );
  AND2X1 U17968 ( .IN1(test_so88), .IN2(WX9910), .Q(n17232) );
  AND2X1 U17969 ( .IN1(n17234), .IN2(n10581), .Q(WX10353) );
  AND2X1 U17970 ( .IN1(n17235), .IN2(n17236), .Q(n17234) );
  OR2X1 U17971 ( .IN1(DFF_1522_n1), .IN2(WX9912), .Q(n17236) );
  OR2X1 U17972 ( .IN1(n9578), .IN2(CRC_OUT_2_18), .Q(n17235) );
  AND2X1 U17973 ( .IN1(n17237), .IN2(n10581), .Q(WX10351) );
  AND2X1 U17974 ( .IN1(n17238), .IN2(n17239), .Q(n17237) );
  OR2X1 U17975 ( .IN1(DFF_1521_n1), .IN2(WX9914), .Q(n17239) );
  OR2X1 U17976 ( .IN1(n9579), .IN2(CRC_OUT_2_17), .Q(n17238) );
  AND2X1 U17977 ( .IN1(n17240), .IN2(n10581), .Q(WX10349) );
  AND2X1 U17978 ( .IN1(n17241), .IN2(n17242), .Q(n17240) );
  OR2X1 U17979 ( .IN1(DFF_1520_n1), .IN2(WX9916), .Q(n17242) );
  OR2X1 U17980 ( .IN1(n9580), .IN2(CRC_OUT_2_16), .Q(n17241) );
  AND2X1 U17981 ( .IN1(n17243), .IN2(n10581), .Q(WX10347) );
  OR2X1 U17982 ( .IN1(n17244), .IN2(n17245), .Q(n17243) );
  AND2X1 U17983 ( .IN1(n17246), .IN2(CRC_OUT_2_15), .Q(n17245) );
  INVX0 U17984 ( .INP(n17247), .ZN(n17246) );
  AND2X1 U17985 ( .IN1(DFF_1519_n1), .IN2(n17247), .Q(n17244) );
  AND2X1 U17986 ( .IN1(n17248), .IN2(n17249), .Q(n17247) );
  OR2X1 U17987 ( .IN1(CRC_OUT_2_31), .IN2(n9515), .Q(n17249) );
  OR2X1 U17988 ( .IN1(WX9918), .IN2(DFF_1535_n1), .Q(n17248) );
  AND2X1 U17989 ( .IN1(n17250), .IN2(n10581), .Q(WX10345) );
  AND2X1 U17990 ( .IN1(n17251), .IN2(n17252), .Q(n17250) );
  OR2X1 U17991 ( .IN1(DFF_1518_n1), .IN2(WX9920), .Q(n17252) );
  OR2X1 U17992 ( .IN1(n9581), .IN2(CRC_OUT_2_14), .Q(n17251) );
  AND2X1 U17993 ( .IN1(n17253), .IN2(n10582), .Q(WX10343) );
  OR2X1 U17994 ( .IN1(n17254), .IN2(n17255), .Q(n17253) );
  AND2X1 U17995 ( .IN1(DFF_1517_n1), .IN2(n9907), .Q(n17255) );
  AND2X1 U17996 ( .IN1(test_so86), .IN2(CRC_OUT_2_13), .Q(n17254) );
  AND2X1 U17997 ( .IN1(n17256), .IN2(n10582), .Q(WX10341) );
  AND2X1 U17998 ( .IN1(n17257), .IN2(n17258), .Q(n17256) );
  OR2X1 U17999 ( .IN1(DFF_1516_n1), .IN2(WX9924), .Q(n17258) );
  OR2X1 U18000 ( .IN1(n9582), .IN2(CRC_OUT_2_12), .Q(n17257) );
  AND2X1 U18001 ( .IN1(n17259), .IN2(n10582), .Q(WX10339) );
  AND2X1 U18002 ( .IN1(n17260), .IN2(n17261), .Q(n17259) );
  OR2X1 U18003 ( .IN1(DFF_1515_n1), .IN2(WX9926), .Q(n17261) );
  OR2X1 U18004 ( .IN1(n9583), .IN2(CRC_OUT_2_11), .Q(n17260) );
  AND2X1 U18005 ( .IN1(n17262), .IN2(n10582), .Q(WX10337) );
  OR2X1 U18006 ( .IN1(n17263), .IN2(n17264), .Q(n17262) );
  AND2X1 U18007 ( .IN1(n17265), .IN2(CRC_OUT_2_10), .Q(n17264) );
  AND2X1 U18008 ( .IN1(DFF_1514_n1), .IN2(n17266), .Q(n17263) );
  INVX0 U18009 ( .INP(n17265), .ZN(n17266) );
  OR2X1 U18010 ( .IN1(n17267), .IN2(n17268), .Q(n17265) );
  AND2X1 U18011 ( .IN1(DFF_1535_n1), .IN2(WX9928), .Q(n17268) );
  AND2X1 U18012 ( .IN1(n9516), .IN2(CRC_OUT_2_31), .Q(n17267) );
  AND2X1 U18013 ( .IN1(n17269), .IN2(n10582), .Q(WX10335) );
  AND2X1 U18014 ( .IN1(n17270), .IN2(n17271), .Q(n17269) );
  OR2X1 U18015 ( .IN1(DFF_1513_n1), .IN2(WX9930), .Q(n17271) );
  OR2X1 U18016 ( .IN1(n9584), .IN2(CRC_OUT_2_9), .Q(n17270) );
  AND2X1 U18017 ( .IN1(n17272), .IN2(n10582), .Q(WX10333) );
  AND2X1 U18018 ( .IN1(n17273), .IN2(n17274), .Q(n17272) );
  OR2X1 U18019 ( .IN1(DFF_1512_n1), .IN2(WX9932), .Q(n17274) );
  OR2X1 U18020 ( .IN1(n9585), .IN2(CRC_OUT_2_8), .Q(n17273) );
  AND2X1 U18021 ( .IN1(n17275), .IN2(n10582), .Q(WX10331) );
  AND2X1 U18022 ( .IN1(n17276), .IN2(n17277), .Q(n17275) );
  OR2X1 U18023 ( .IN1(DFF_1511_n1), .IN2(WX9934), .Q(n17277) );
  OR2X1 U18024 ( .IN1(n9586), .IN2(CRC_OUT_2_7), .Q(n17276) );
  AND2X1 U18025 ( .IN1(n17278), .IN2(n10582), .Q(WX10329) );
  AND2X1 U18026 ( .IN1(n17279), .IN2(n17280), .Q(n17278) );
  OR2X1 U18027 ( .IN1(DFF_1510_n1), .IN2(WX9936), .Q(n17280) );
  OR2X1 U18028 ( .IN1(n9587), .IN2(CRC_OUT_2_6), .Q(n17279) );
  AND2X1 U18029 ( .IN1(n17281), .IN2(n10582), .Q(WX10327) );
  AND2X1 U18030 ( .IN1(n17282), .IN2(n17283), .Q(n17281) );
  OR2X1 U18031 ( .IN1(DFF_1509_n1), .IN2(WX9938), .Q(n17283) );
  OR2X1 U18032 ( .IN1(n9588), .IN2(CRC_OUT_2_5), .Q(n17282) );
  AND2X1 U18033 ( .IN1(n17284), .IN2(n10583), .Q(WX10325) );
  AND2X1 U18034 ( .IN1(n17285), .IN2(n17286), .Q(n17284) );
  OR2X1 U18035 ( .IN1(DFF_1508_n1), .IN2(WX9940), .Q(n17286) );
  OR2X1 U18036 ( .IN1(n9589), .IN2(CRC_OUT_2_4), .Q(n17285) );
  AND2X1 U18037 ( .IN1(n17287), .IN2(n10583), .Q(WX10323) );
  OR2X1 U18038 ( .IN1(n17288), .IN2(n17289), .Q(n17287) );
  AND2X1 U18039 ( .IN1(n17290), .IN2(CRC_OUT_2_3), .Q(n17289) );
  AND2X1 U18040 ( .IN1(DFF_1507_n1), .IN2(n17291), .Q(n17288) );
  INVX0 U18041 ( .INP(n17290), .ZN(n17291) );
  OR2X1 U18042 ( .IN1(n17292), .IN2(n17293), .Q(n17290) );
  AND2X1 U18043 ( .IN1(DFF_1535_n1), .IN2(WX9942), .Q(n17293) );
  AND2X1 U18044 ( .IN1(n9517), .IN2(CRC_OUT_2_31), .Q(n17292) );
  AND2X1 U18045 ( .IN1(n17294), .IN2(n10583), .Q(WX10321) );
  OR2X1 U18046 ( .IN1(n17295), .IN2(n17296), .Q(n17294) );
  AND2X1 U18047 ( .IN1(n9590), .IN2(n9952), .Q(n17296) );
  AND2X1 U18048 ( .IN1(test_so87), .IN2(WX9944), .Q(n17295) );
  AND2X1 U18049 ( .IN1(n17297), .IN2(n10583), .Q(WX10319) );
  AND2X1 U18050 ( .IN1(n17298), .IN2(n17299), .Q(n17297) );
  OR2X1 U18051 ( .IN1(DFF_1505_n1), .IN2(WX9946), .Q(n17299) );
  OR2X1 U18052 ( .IN1(n9591), .IN2(CRC_OUT_2_1), .Q(n17298) );
  AND2X1 U18053 ( .IN1(n17300), .IN2(n10555), .Q(WX10317) );
  AND2X1 U18054 ( .IN1(n17301), .IN2(n17302), .Q(n17300) );
  OR2X1 U18055 ( .IN1(DFF_1504_n1), .IN2(WX9948), .Q(n17302) );
  OR2X1 U18056 ( .IN1(n9592), .IN2(CRC_OUT_2_0), .Q(n17301) );
  AND2X1 U18057 ( .IN1(n17303), .IN2(n10570), .Q(WX10315) );
  AND2X1 U18058 ( .IN1(n17304), .IN2(n17305), .Q(n17303) );
  OR2X1 U18059 ( .IN1(DFF_1535_n1), .IN2(WX9950), .Q(n17305) );
  OR2X1 U18060 ( .IN1(n9534), .IN2(CRC_OUT_2_31), .Q(n17304) );
  OR2X1 U18061 ( .IN1(n17306), .IN2(n17307), .Q(DATA_9_9) );
  AND2X1 U18062 ( .IN1(n12771), .IN2(n17308), .Q(n17307) );
  INVX0 U18063 ( .INP(n17309), .ZN(n17306) );
  OR2X1 U18064 ( .IN1(n17308), .IN2(n12771), .Q(n17309) );
  OR2X1 U18065 ( .IN1(n17310), .IN2(n17311), .Q(n12771) );
  INVX0 U18066 ( .INP(n17312), .ZN(n17311) );
  OR2X1 U18067 ( .IN1(n17313), .IN2(n17314), .Q(n17312) );
  AND2X1 U18068 ( .IN1(n17314), .IN2(n17313), .Q(n17310) );
  AND2X1 U18069 ( .IN1(n17315), .IN2(n17316), .Q(n17313) );
  OR2X1 U18070 ( .IN1(n2182), .IN2(n3485), .Q(n17316) );
  OR2X1 U18071 ( .IN1(WX689), .IN2(TM0), .Q(n17315) );
  OR2X1 U18072 ( .IN1(n17317), .IN2(n17318), .Q(n17314) );
  AND2X1 U18073 ( .IN1(n9797), .IN2(n17319), .Q(n17318) );
  AND2X1 U18074 ( .IN1(n17320), .IN2(n17321), .Q(n17319) );
  OR2X1 U18075 ( .IN1(n9795), .IN2(WX817), .Q(n17321) );
  OR2X1 U18076 ( .IN1(n9796), .IN2(WX753), .Q(n17320) );
  AND2X1 U18077 ( .IN1(n17322), .IN2(WX881), .Q(n17317) );
  OR2X1 U18078 ( .IN1(n17323), .IN2(n17324), .Q(n17322) );
  AND2X1 U18079 ( .IN1(n9795), .IN2(WX817), .Q(n17324) );
  AND2X1 U18080 ( .IN1(n9796), .IN2(WX753), .Q(n17323) );
  OR2X1 U18081 ( .IN1(n9883), .IN2(n2182), .Q(n17308) );
  OR2X1 U18082 ( .IN1(n17325), .IN2(n17326), .Q(DATA_9_8) );
  AND2X1 U18083 ( .IN1(n12763), .IN2(n17327), .Q(n17326) );
  INVX0 U18084 ( .INP(n17328), .ZN(n17325) );
  OR2X1 U18085 ( .IN1(n17327), .IN2(n12763), .Q(n17328) );
  OR2X1 U18086 ( .IN1(n17329), .IN2(n17330), .Q(n12763) );
  INVX0 U18087 ( .INP(n17331), .ZN(n17330) );
  OR2X1 U18088 ( .IN1(n17332), .IN2(n17333), .Q(n17331) );
  AND2X1 U18089 ( .IN1(n17333), .IN2(n17332), .Q(n17329) );
  AND2X1 U18090 ( .IN1(n17334), .IN2(n17335), .Q(n17332) );
  OR2X1 U18091 ( .IN1(n2182), .IN2(n3483), .Q(n17335) );
  OR2X1 U18092 ( .IN1(WX691), .IN2(TM0), .Q(n17334) );
  OR2X1 U18093 ( .IN1(n17336), .IN2(n17337), .Q(n17333) );
  INVX0 U18094 ( .INP(n17338), .ZN(n17337) );
  OR2X1 U18095 ( .IN1(n17339), .IN2(n9805), .Q(n17338) );
  AND2X1 U18096 ( .IN1(n9805), .IN2(n17339), .Q(n17336) );
  AND2X1 U18097 ( .IN1(n17340), .IN2(n17341), .Q(n17339) );
  OR2X1 U18098 ( .IN1(WX883), .IN2(n9807), .Q(n17341) );
  OR2X1 U18099 ( .IN1(WX755), .IN2(n9806), .Q(n17340) );
  OR2X1 U18100 ( .IN1(n9882), .IN2(n2182), .Q(n17327) );
  OR2X1 U18101 ( .IN1(n17342), .IN2(n17343), .Q(DATA_9_7) );
  AND2X1 U18102 ( .IN1(n12755), .IN2(n17344), .Q(n17343) );
  INVX0 U18103 ( .INP(n17345), .ZN(n17342) );
  OR2X1 U18104 ( .IN1(n17344), .IN2(n12755), .Q(n17345) );
  OR2X1 U18105 ( .IN1(n17346), .IN2(n17347), .Q(n12755) );
  INVX0 U18106 ( .INP(n17348), .ZN(n17347) );
  OR2X1 U18107 ( .IN1(n17349), .IN2(n17350), .Q(n17348) );
  AND2X1 U18108 ( .IN1(n17350), .IN2(n17349), .Q(n17346) );
  AND2X1 U18109 ( .IN1(n17351), .IN2(n17352), .Q(n17349) );
  OR2X1 U18110 ( .IN1(n2182), .IN2(n3481), .Q(n17352) );
  OR2X1 U18111 ( .IN1(WX693), .IN2(TM0), .Q(n17351) );
  OR2X1 U18112 ( .IN1(n17353), .IN2(n17354), .Q(n17350) );
  AND2X1 U18113 ( .IN1(n9837), .IN2(n17355), .Q(n17354) );
  AND2X1 U18114 ( .IN1(n17356), .IN2(n17357), .Q(n17355) );
  OR2X1 U18115 ( .IN1(n9835), .IN2(WX821), .Q(n17357) );
  OR2X1 U18116 ( .IN1(n9836), .IN2(WX757), .Q(n17356) );
  AND2X1 U18117 ( .IN1(n17358), .IN2(WX885), .Q(n17353) );
  OR2X1 U18118 ( .IN1(n17359), .IN2(n17360), .Q(n17358) );
  AND2X1 U18119 ( .IN1(n9835), .IN2(WX821), .Q(n17360) );
  AND2X1 U18120 ( .IN1(n9836), .IN2(WX757), .Q(n17359) );
  OR2X1 U18121 ( .IN1(n9881), .IN2(n2182), .Q(n17344) );
  OR2X1 U18122 ( .IN1(n17361), .IN2(n17362), .Q(DATA_9_6) );
  AND2X1 U18123 ( .IN1(n12747), .IN2(n17363), .Q(n17362) );
  INVX0 U18124 ( .INP(n17364), .ZN(n17361) );
  OR2X1 U18125 ( .IN1(n17363), .IN2(n12747), .Q(n17364) );
  AND2X1 U18126 ( .IN1(n17365), .IN2(n17366), .Q(n12747) );
  OR2X1 U18127 ( .IN1(n17367), .IN2(n17368), .Q(n17366) );
  INVX0 U18128 ( .INP(n17369), .ZN(n17365) );
  AND2X1 U18129 ( .IN1(n17368), .IN2(n17367), .Q(n17369) );
  AND2X1 U18130 ( .IN1(n17370), .IN2(n17371), .Q(n17367) );
  OR2X1 U18131 ( .IN1(n2182), .IN2(n3479), .Q(n17371) );
  OR2X1 U18132 ( .IN1(WX695), .IN2(TM0), .Q(n17370) );
  OR2X1 U18133 ( .IN1(n17372), .IN2(n17373), .Q(n17368) );
  AND2X1 U18134 ( .IN1(n9824), .IN2(n17374), .Q(n17373) );
  AND2X1 U18135 ( .IN1(n17375), .IN2(n17376), .Q(n17374) );
  OR2X1 U18136 ( .IN1(n9823), .IN2(n9897), .Q(n17376) );
  OR2X1 U18137 ( .IN1(test_so5), .IN2(WX823), .Q(n17375) );
  AND2X1 U18138 ( .IN1(n17377), .IN2(WX887), .Q(n17372) );
  OR2X1 U18139 ( .IN1(n17378), .IN2(n17379), .Q(n17377) );
  AND2X1 U18140 ( .IN1(n9823), .IN2(n9897), .Q(n17379) );
  AND2X1 U18141 ( .IN1(test_so5), .IN2(WX823), .Q(n17378) );
  OR2X1 U18142 ( .IN1(n9880), .IN2(n2182), .Q(n17363) );
  OR2X1 U18143 ( .IN1(n17380), .IN2(n17381), .Q(DATA_9_5) );
  AND2X1 U18144 ( .IN1(n12739), .IN2(n17382), .Q(n17381) );
  INVX0 U18145 ( .INP(n17383), .ZN(n17380) );
  OR2X1 U18146 ( .IN1(n17382), .IN2(n12739), .Q(n17383) );
  OR2X1 U18147 ( .IN1(n17384), .IN2(n17385), .Q(n12739) );
  INVX0 U18148 ( .INP(n17386), .ZN(n17385) );
  OR2X1 U18149 ( .IN1(n17387), .IN2(n17388), .Q(n17386) );
  AND2X1 U18150 ( .IN1(n17388), .IN2(n17387), .Q(n17384) );
  AND2X1 U18151 ( .IN1(n17389), .IN2(n17390), .Q(n17387) );
  OR2X1 U18152 ( .IN1(n2182), .IN2(n3477), .Q(n17390) );
  OR2X1 U18153 ( .IN1(WX697), .IN2(TM0), .Q(n17389) );
  OR2X1 U18154 ( .IN1(n17391), .IN2(n17392), .Q(n17388) );
  INVX0 U18155 ( .INP(n17393), .ZN(n17392) );
  OR2X1 U18156 ( .IN1(n17394), .IN2(n9808), .Q(n17393) );
  AND2X1 U18157 ( .IN1(n9808), .IN2(n17394), .Q(n17391) );
  AND2X1 U18158 ( .IN1(n17395), .IN2(n17396), .Q(n17394) );
  OR2X1 U18159 ( .IN1(WX889), .IN2(n9810), .Q(n17396) );
  OR2X1 U18160 ( .IN1(WX761), .IN2(n9809), .Q(n17395) );
  OR2X1 U18161 ( .IN1(n9879), .IN2(n2182), .Q(n17382) );
  OR2X1 U18162 ( .IN1(n17397), .IN2(n17398), .Q(DATA_9_4) );
  AND2X1 U18163 ( .IN1(n12731), .IN2(n17399), .Q(n17398) );
  INVX0 U18164 ( .INP(n17400), .ZN(n17397) );
  OR2X1 U18165 ( .IN1(n17399), .IN2(n12731), .Q(n17400) );
  OR2X1 U18166 ( .IN1(n17401), .IN2(n17402), .Q(n12731) );
  INVX0 U18167 ( .INP(n17403), .ZN(n17402) );
  OR2X1 U18168 ( .IN1(n17404), .IN2(n17405), .Q(n17403) );
  AND2X1 U18169 ( .IN1(n17405), .IN2(n17404), .Q(n17401) );
  AND2X1 U18170 ( .IN1(n17406), .IN2(n17407), .Q(n17404) );
  OR2X1 U18171 ( .IN1(n2182), .IN2(n3475), .Q(n17407) );
  OR2X1 U18172 ( .IN1(WX699), .IN2(TM0), .Q(n17406) );
  OR2X1 U18173 ( .IN1(n17408), .IN2(n17409), .Q(n17405) );
  INVX0 U18174 ( .INP(n17410), .ZN(n17409) );
  OR2X1 U18175 ( .IN1(n17411), .IN2(n9811), .Q(n17410) );
  AND2X1 U18176 ( .IN1(n9811), .IN2(n17411), .Q(n17408) );
  AND2X1 U18177 ( .IN1(n17412), .IN2(n17413), .Q(n17411) );
  OR2X1 U18178 ( .IN1(WX891), .IN2(n9813), .Q(n17413) );
  OR2X1 U18179 ( .IN1(WX763), .IN2(n9812), .Q(n17412) );
  OR2X1 U18180 ( .IN1(n9878), .IN2(n2182), .Q(n17399) );
  OR2X1 U18181 ( .IN1(n17414), .IN2(n17415), .Q(DATA_9_31) );
  AND2X1 U18182 ( .IN1(n13051), .IN2(n17416), .Q(n17415) );
  INVX0 U18183 ( .INP(n17417), .ZN(n17414) );
  OR2X1 U18184 ( .IN1(n17416), .IN2(n13051), .Q(n17417) );
  OR2X1 U18185 ( .IN1(n17418), .IN2(n17419), .Q(n13051) );
  INVX0 U18186 ( .INP(n17420), .ZN(n17419) );
  OR2X1 U18187 ( .IN1(n17421), .IN2(n17422), .Q(n17420) );
  AND2X1 U18188 ( .IN1(n17422), .IN2(n17421), .Q(n17418) );
  AND2X1 U18189 ( .IN1(n17423), .IN2(n17424), .Q(n17421) );
  OR2X1 U18190 ( .IN1(n10538), .IN2(n3529), .Q(n17424) );
  OR2X1 U18191 ( .IN1(WX645), .IN2(n10516), .Q(n17423) );
  OR2X1 U18192 ( .IN1(n17425), .IN2(n17426), .Q(n17422) );
  AND2X1 U18193 ( .IN1(n9829), .IN2(n17427), .Q(n17426) );
  AND2X1 U18194 ( .IN1(n17428), .IN2(n17429), .Q(n17427) );
  OR2X1 U18195 ( .IN1(n9827), .IN2(WX773), .Q(n17429) );
  OR2X1 U18196 ( .IN1(n9828), .IN2(WX709), .Q(n17428) );
  AND2X1 U18197 ( .IN1(n17430), .IN2(WX837), .Q(n17425) );
  OR2X1 U18198 ( .IN1(n17431), .IN2(n17432), .Q(n17430) );
  AND2X1 U18199 ( .IN1(n9827), .IN2(WX773), .Q(n17432) );
  AND2X1 U18200 ( .IN1(n9828), .IN2(WX709), .Q(n17431) );
  OR2X1 U18201 ( .IN1(n9877), .IN2(n2182), .Q(n17416) );
  OR2X1 U18202 ( .IN1(n17433), .IN2(n17434), .Q(DATA_9_30) );
  AND2X1 U18203 ( .IN1(n13005), .IN2(n17435), .Q(n17434) );
  INVX0 U18204 ( .INP(n17436), .ZN(n17433) );
  OR2X1 U18205 ( .IN1(n17435), .IN2(n13005), .Q(n17436) );
  OR2X1 U18206 ( .IN1(n17437), .IN2(n17438), .Q(n13005) );
  INVX0 U18207 ( .INP(n17439), .ZN(n17438) );
  OR2X1 U18208 ( .IN1(n17440), .IN2(n17441), .Q(n17439) );
  AND2X1 U18209 ( .IN1(n17441), .IN2(n17440), .Q(n17437) );
  AND2X1 U18210 ( .IN1(n17442), .IN2(n17443), .Q(n17440) );
  OR2X1 U18211 ( .IN1(n10538), .IN2(n3527), .Q(n17443) );
  OR2X1 U18212 ( .IN1(WX647), .IN2(n10516), .Q(n17442) );
  OR2X1 U18213 ( .IN1(n17444), .IN2(n17445), .Q(n17441) );
  AND2X1 U18214 ( .IN1(n9755), .IN2(n17446), .Q(n17445) );
  AND2X1 U18215 ( .IN1(n17447), .IN2(n17448), .Q(n17446) );
  OR2X1 U18216 ( .IN1(n9753), .IN2(WX775), .Q(n17448) );
  OR2X1 U18217 ( .IN1(n9754), .IN2(WX711), .Q(n17447) );
  AND2X1 U18218 ( .IN1(n17449), .IN2(WX839), .Q(n17444) );
  OR2X1 U18219 ( .IN1(n17450), .IN2(n17451), .Q(n17449) );
  AND2X1 U18220 ( .IN1(n9753), .IN2(WX775), .Q(n17451) );
  AND2X1 U18221 ( .IN1(n9754), .IN2(WX711), .Q(n17450) );
  OR2X1 U18222 ( .IN1(n9876), .IN2(n2182), .Q(n17435) );
  OR2X1 U18223 ( .IN1(n17452), .IN2(n17453), .Q(DATA_9_3) );
  AND2X1 U18224 ( .IN1(n12723), .IN2(n17454), .Q(n17453) );
  INVX0 U18225 ( .INP(n17455), .ZN(n17452) );
  OR2X1 U18226 ( .IN1(n17454), .IN2(n12723), .Q(n17455) );
  OR2X1 U18227 ( .IN1(n17456), .IN2(n17457), .Q(n12723) );
  INVX0 U18228 ( .INP(n17458), .ZN(n17457) );
  OR2X1 U18229 ( .IN1(n17459), .IN2(n17460), .Q(n17458) );
  AND2X1 U18230 ( .IN1(n17460), .IN2(n17459), .Q(n17456) );
  AND2X1 U18231 ( .IN1(n17461), .IN2(n17462), .Q(n17459) );
  OR2X1 U18232 ( .IN1(n2182), .IN2(n3473), .Q(n17462) );
  OR2X1 U18233 ( .IN1(WX701), .IN2(TM0), .Q(n17461) );
  OR2X1 U18234 ( .IN1(n17463), .IN2(n17464), .Q(n17460) );
  INVX0 U18235 ( .INP(n17465), .ZN(n17464) );
  OR2X1 U18236 ( .IN1(n17466), .IN2(n9756), .Q(n17465) );
  AND2X1 U18237 ( .IN1(n9756), .IN2(n17466), .Q(n17463) );
  AND2X1 U18238 ( .IN1(n17467), .IN2(n17468), .Q(n17466) );
  OR2X1 U18239 ( .IN1(WX893), .IN2(n9758), .Q(n17468) );
  OR2X1 U18240 ( .IN1(WX765), .IN2(n9757), .Q(n17467) );
  OR2X1 U18241 ( .IN1(n9875), .IN2(n2182), .Q(n17454) );
  OR2X1 U18242 ( .IN1(n17469), .IN2(n17470), .Q(DATA_9_29) );
  AND2X1 U18243 ( .IN1(n12961), .IN2(n17471), .Q(n17470) );
  INVX0 U18244 ( .INP(n17472), .ZN(n17469) );
  OR2X1 U18245 ( .IN1(n17471), .IN2(n12961), .Q(n17472) );
  OR2X1 U18246 ( .IN1(n17473), .IN2(n17474), .Q(n12961) );
  INVX0 U18247 ( .INP(n17475), .ZN(n17474) );
  OR2X1 U18248 ( .IN1(n17476), .IN2(n17477), .Q(n17475) );
  AND2X1 U18249 ( .IN1(n17477), .IN2(n17476), .Q(n17473) );
  AND2X1 U18250 ( .IN1(n17478), .IN2(n17479), .Q(n17476) );
  OR2X1 U18251 ( .IN1(n10538), .IN2(n3525), .Q(n17479) );
  OR2X1 U18252 ( .IN1(WX649), .IN2(n10516), .Q(n17478) );
  OR2X1 U18253 ( .IN1(n17480), .IN2(n17481), .Q(n17477) );
  INVX0 U18254 ( .INP(n17482), .ZN(n17481) );
  OR2X1 U18255 ( .IN1(n17483), .IN2(n9762), .Q(n17482) );
  AND2X1 U18256 ( .IN1(n9762), .IN2(n17483), .Q(n17480) );
  AND2X1 U18257 ( .IN1(n17484), .IN2(n17485), .Q(n17483) );
  OR2X1 U18258 ( .IN1(WX841), .IN2(n9764), .Q(n17485) );
  OR2X1 U18259 ( .IN1(WX713), .IN2(n9763), .Q(n17484) );
  OR2X1 U18260 ( .IN1(n9874), .IN2(n2182), .Q(n17471) );
  OR2X1 U18261 ( .IN1(n17486), .IN2(n17487), .Q(DATA_9_28) );
  AND2X1 U18262 ( .IN1(n12923), .IN2(n17488), .Q(n17487) );
  INVX0 U18263 ( .INP(n17489), .ZN(n17486) );
  OR2X1 U18264 ( .IN1(n17488), .IN2(n12923), .Q(n17489) );
  AND2X1 U18265 ( .IN1(n17490), .IN2(n17491), .Q(n12923) );
  OR2X1 U18266 ( .IN1(n17492), .IN2(n17493), .Q(n17491) );
  INVX0 U18267 ( .INP(n17494), .ZN(n17490) );
  AND2X1 U18268 ( .IN1(n17493), .IN2(n17492), .Q(n17494) );
  AND2X1 U18269 ( .IN1(n17495), .IN2(n17496), .Q(n17492) );
  OR2X1 U18270 ( .IN1(n10538), .IN2(n9773), .Q(n17496) );
  OR2X1 U18271 ( .IN1(WX715), .IN2(n10516), .Q(n17495) );
  OR2X1 U18272 ( .IN1(n17497), .IN2(n17498), .Q(n17493) );
  AND2X1 U18273 ( .IN1(n9772), .IN2(n17499), .Q(n17498) );
  AND2X1 U18274 ( .IN1(n17500), .IN2(n17501), .Q(n17499) );
  OR2X1 U18275 ( .IN1(n9771), .IN2(n9898), .Q(n17501) );
  OR2X1 U18276 ( .IN1(test_so2), .IN2(WX779), .Q(n17500) );
  AND2X1 U18277 ( .IN1(n17502), .IN2(WX843), .Q(n17497) );
  OR2X1 U18278 ( .IN1(n17503), .IN2(n17504), .Q(n17502) );
  AND2X1 U18279 ( .IN1(n9771), .IN2(n9898), .Q(n17504) );
  AND2X1 U18280 ( .IN1(test_so2), .IN2(WX779), .Q(n17503) );
  OR2X1 U18281 ( .IN1(n9873), .IN2(n2182), .Q(n17488) );
  OR2X1 U18282 ( .IN1(n17505), .IN2(n17506), .Q(DATA_9_27) );
  AND2X1 U18283 ( .IN1(n12915), .IN2(n17507), .Q(n17506) );
  INVX0 U18284 ( .INP(n17508), .ZN(n17505) );
  OR2X1 U18285 ( .IN1(n17507), .IN2(n12915), .Q(n17508) );
  OR2X1 U18286 ( .IN1(n17509), .IN2(n17510), .Q(n12915) );
  INVX0 U18287 ( .INP(n17511), .ZN(n17510) );
  OR2X1 U18288 ( .IN1(n17512), .IN2(n17513), .Q(n17511) );
  AND2X1 U18289 ( .IN1(n17513), .IN2(n17512), .Q(n17509) );
  AND2X1 U18290 ( .IN1(n17514), .IN2(n17515), .Q(n17512) );
  OR2X1 U18291 ( .IN1(n10537), .IN2(n3521), .Q(n17515) );
  OR2X1 U18292 ( .IN1(WX653), .IN2(n10515), .Q(n17514) );
  OR2X1 U18293 ( .IN1(n17516), .IN2(n17517), .Q(n17513) );
  INVX0 U18294 ( .INP(n17518), .ZN(n17517) );
  OR2X1 U18295 ( .IN1(n17519), .IN2(n9777), .Q(n17518) );
  AND2X1 U18296 ( .IN1(n9777), .IN2(n17519), .Q(n17516) );
  AND2X1 U18297 ( .IN1(n17520), .IN2(n17521), .Q(n17519) );
  OR2X1 U18298 ( .IN1(WX845), .IN2(n9779), .Q(n17521) );
  OR2X1 U18299 ( .IN1(WX717), .IN2(n9778), .Q(n17520) );
  OR2X1 U18300 ( .IN1(n9872), .IN2(n2182), .Q(n17507) );
  OR2X1 U18301 ( .IN1(n17522), .IN2(n17523), .Q(DATA_9_26) );
  AND2X1 U18302 ( .IN1(n12907), .IN2(n17524), .Q(n17523) );
  INVX0 U18303 ( .INP(n17525), .ZN(n17522) );
  OR2X1 U18304 ( .IN1(n17524), .IN2(n12907), .Q(n17525) );
  OR2X1 U18305 ( .IN1(n17526), .IN2(n17527), .Q(n12907) );
  INVX0 U18306 ( .INP(n17528), .ZN(n17527) );
  OR2X1 U18307 ( .IN1(n17529), .IN2(n17530), .Q(n17528) );
  AND2X1 U18308 ( .IN1(n17530), .IN2(n17529), .Q(n17526) );
  AND2X1 U18309 ( .IN1(n17531), .IN2(n17532), .Q(n17529) );
  OR2X1 U18310 ( .IN1(n10537), .IN2(n3519), .Q(n17532) );
  OR2X1 U18311 ( .IN1(WX655), .IN2(n10515), .Q(n17531) );
  OR2X1 U18312 ( .IN1(n17533), .IN2(n17534), .Q(n17530) );
  INVX0 U18313 ( .INP(n17535), .ZN(n17534) );
  OR2X1 U18314 ( .IN1(n17536), .IN2(n9780), .Q(n17535) );
  AND2X1 U18315 ( .IN1(n9780), .IN2(n17536), .Q(n17533) );
  AND2X1 U18316 ( .IN1(n17537), .IN2(n17538), .Q(n17536) );
  OR2X1 U18317 ( .IN1(WX847), .IN2(n9782), .Q(n17538) );
  OR2X1 U18318 ( .IN1(WX719), .IN2(n9781), .Q(n17537) );
  OR2X1 U18319 ( .IN1(n9871), .IN2(n2182), .Q(n17524) );
  OR2X1 U18320 ( .IN1(n17539), .IN2(n17540), .Q(DATA_9_25) );
  AND2X1 U18321 ( .IN1(n12899), .IN2(n17541), .Q(n17540) );
  INVX0 U18322 ( .INP(n17542), .ZN(n17539) );
  OR2X1 U18323 ( .IN1(n17541), .IN2(n12899), .Q(n17542) );
  OR2X1 U18324 ( .IN1(n17543), .IN2(n17544), .Q(n12899) );
  INVX0 U18325 ( .INP(n17545), .ZN(n17544) );
  OR2X1 U18326 ( .IN1(n17546), .IN2(n17547), .Q(n17545) );
  AND2X1 U18327 ( .IN1(n17547), .IN2(n17546), .Q(n17543) );
  AND2X1 U18328 ( .IN1(n17548), .IN2(n17549), .Q(n17546) );
  OR2X1 U18329 ( .IN1(n10537), .IN2(n3517), .Q(n17549) );
  OR2X1 U18330 ( .IN1(WX657), .IN2(n10515), .Q(n17548) );
  OR2X1 U18331 ( .IN1(n17550), .IN2(n17551), .Q(n17547) );
  INVX0 U18332 ( .INP(n17552), .ZN(n17551) );
  OR2X1 U18333 ( .IN1(n17553), .IN2(n9789), .Q(n17552) );
  AND2X1 U18334 ( .IN1(n9789), .IN2(n17553), .Q(n17550) );
  AND2X1 U18335 ( .IN1(n17554), .IN2(n17555), .Q(n17553) );
  OR2X1 U18336 ( .IN1(WX849), .IN2(n9791), .Q(n17555) );
  OR2X1 U18337 ( .IN1(WX721), .IN2(n9790), .Q(n17554) );
  OR2X1 U18338 ( .IN1(n9870), .IN2(n2182), .Q(n17541) );
  OR2X1 U18339 ( .IN1(n17556), .IN2(n17557), .Q(DATA_9_24) );
  AND2X1 U18340 ( .IN1(n12891), .IN2(n17558), .Q(n17557) );
  INVX0 U18341 ( .INP(n17559), .ZN(n17556) );
  OR2X1 U18342 ( .IN1(n17558), .IN2(n12891), .Q(n17559) );
  AND2X1 U18343 ( .IN1(n17560), .IN2(n17561), .Q(n12891) );
  OR2X1 U18344 ( .IN1(n17562), .IN2(n17563), .Q(n17561) );
  INVX0 U18345 ( .INP(n17564), .ZN(n17560) );
  AND2X1 U18346 ( .IN1(n17563), .IN2(n17562), .Q(n17564) );
  AND2X1 U18347 ( .IN1(n17565), .IN2(n17566), .Q(n17562) );
  OR2X1 U18348 ( .IN1(n10537), .IN2(n3515), .Q(n17566) );
  OR2X1 U18349 ( .IN1(WX659), .IN2(n10515), .Q(n17565) );
  OR2X1 U18350 ( .IN1(n17567), .IN2(n17568), .Q(n17563) );
  AND2X1 U18351 ( .IN1(n9799), .IN2(n17569), .Q(n17568) );
  AND2X1 U18352 ( .IN1(n17570), .IN2(n17571), .Q(n17569) );
  OR2X1 U18353 ( .IN1(n9798), .IN2(n9899), .Q(n17571) );
  OR2X1 U18354 ( .IN1(test_so4), .IN2(WX787), .Q(n17570) );
  AND2X1 U18355 ( .IN1(n17572), .IN2(WX851), .Q(n17567) );
  OR2X1 U18356 ( .IN1(n17573), .IN2(n17574), .Q(n17572) );
  AND2X1 U18357 ( .IN1(n9798), .IN2(n9899), .Q(n17574) );
  AND2X1 U18358 ( .IN1(test_so4), .IN2(WX787), .Q(n17573) );
  OR2X1 U18359 ( .IN1(n9869), .IN2(n2182), .Q(n17558) );
  OR2X1 U18360 ( .IN1(n17575), .IN2(n17576), .Q(DATA_9_23) );
  AND2X1 U18361 ( .IN1(n12883), .IN2(n17577), .Q(n17576) );
  INVX0 U18362 ( .INP(n17578), .ZN(n17575) );
  OR2X1 U18363 ( .IN1(n17577), .IN2(n12883), .Q(n17578) );
  OR2X1 U18364 ( .IN1(n17579), .IN2(n17580), .Q(n12883) );
  INVX0 U18365 ( .INP(n17581), .ZN(n17580) );
  OR2X1 U18366 ( .IN1(n17582), .IN2(n17583), .Q(n17581) );
  AND2X1 U18367 ( .IN1(n17583), .IN2(n17582), .Q(n17579) );
  AND2X1 U18368 ( .IN1(n17584), .IN2(n17585), .Q(n17582) );
  OR2X1 U18369 ( .IN1(n10537), .IN2(n3513), .Q(n17585) );
  OR2X1 U18370 ( .IN1(WX661), .IN2(n10515), .Q(n17584) );
  OR2X1 U18371 ( .IN1(n17586), .IN2(n17587), .Q(n17583) );
  INVX0 U18372 ( .INP(n17588), .ZN(n17587) );
  OR2X1 U18373 ( .IN1(n17589), .IN2(n9800), .Q(n17588) );
  AND2X1 U18374 ( .IN1(n9800), .IN2(n17589), .Q(n17586) );
  AND2X1 U18375 ( .IN1(n17590), .IN2(n17591), .Q(n17589) );
  OR2X1 U18376 ( .IN1(WX853), .IN2(n9802), .Q(n17591) );
  OR2X1 U18377 ( .IN1(WX725), .IN2(n9801), .Q(n17590) );
  OR2X1 U18378 ( .IN1(n9868), .IN2(n2182), .Q(n17577) );
  OR2X1 U18379 ( .IN1(n17592), .IN2(n17593), .Q(DATA_9_22) );
  AND2X1 U18380 ( .IN1(n12875), .IN2(n17594), .Q(n17593) );
  INVX0 U18381 ( .INP(n17595), .ZN(n17592) );
  OR2X1 U18382 ( .IN1(n17594), .IN2(n12875), .Q(n17595) );
  OR2X1 U18383 ( .IN1(n17596), .IN2(n17597), .Q(n12875) );
  INVX0 U18384 ( .INP(n17598), .ZN(n17597) );
  OR2X1 U18385 ( .IN1(n17599), .IN2(n17600), .Q(n17598) );
  AND2X1 U18386 ( .IN1(n17600), .IN2(n17599), .Q(n17596) );
  AND2X1 U18387 ( .IN1(n17601), .IN2(n17602), .Q(n17599) );
  OR2X1 U18388 ( .IN1(n10537), .IN2(n3511), .Q(n17602) );
  OR2X1 U18389 ( .IN1(WX663), .IN2(n10515), .Q(n17601) );
  OR2X1 U18390 ( .IN1(n17603), .IN2(n17604), .Q(n17600) );
  AND2X1 U18391 ( .IN1(n9816), .IN2(n17605), .Q(n17604) );
  AND2X1 U18392 ( .IN1(n17606), .IN2(n17607), .Q(n17605) );
  OR2X1 U18393 ( .IN1(n9814), .IN2(WX791), .Q(n17607) );
  OR2X1 U18394 ( .IN1(n9815), .IN2(WX727), .Q(n17606) );
  AND2X1 U18395 ( .IN1(n17608), .IN2(WX855), .Q(n17603) );
  OR2X1 U18396 ( .IN1(n17609), .IN2(n17610), .Q(n17608) );
  AND2X1 U18397 ( .IN1(n9814), .IN2(WX791), .Q(n17610) );
  AND2X1 U18398 ( .IN1(n9815), .IN2(WX727), .Q(n17609) );
  OR2X1 U18399 ( .IN1(n9867), .IN2(n2182), .Q(n17594) );
  OR2X1 U18400 ( .IN1(n17611), .IN2(n17612), .Q(DATA_9_21) );
  AND2X1 U18401 ( .IN1(n12867), .IN2(n17613), .Q(n17612) );
  INVX0 U18402 ( .INP(n17614), .ZN(n17611) );
  OR2X1 U18403 ( .IN1(n17613), .IN2(n12867), .Q(n17614) );
  OR2X1 U18404 ( .IN1(n17615), .IN2(n17616), .Q(n12867) );
  INVX0 U18405 ( .INP(n17617), .ZN(n17616) );
  OR2X1 U18406 ( .IN1(n17618), .IN2(n17619), .Q(n17617) );
  AND2X1 U18407 ( .IN1(n17619), .IN2(n17618), .Q(n17615) );
  AND2X1 U18408 ( .IN1(n17620), .IN2(n17621), .Q(n17618) );
  OR2X1 U18409 ( .IN1(n10537), .IN2(n3509), .Q(n17621) );
  OR2X1 U18410 ( .IN1(WX665), .IN2(n10514), .Q(n17620) );
  OR2X1 U18411 ( .IN1(n17622), .IN2(n17623), .Q(n17619) );
  AND2X1 U18412 ( .IN1(n9822), .IN2(n17624), .Q(n17623) );
  AND2X1 U18413 ( .IN1(n17625), .IN2(n17626), .Q(n17624) );
  OR2X1 U18414 ( .IN1(n9820), .IN2(WX793), .Q(n17626) );
  OR2X1 U18415 ( .IN1(n9821), .IN2(WX729), .Q(n17625) );
  AND2X1 U18416 ( .IN1(n17627), .IN2(WX857), .Q(n17622) );
  OR2X1 U18417 ( .IN1(n17628), .IN2(n17629), .Q(n17627) );
  AND2X1 U18418 ( .IN1(n9820), .IN2(WX793), .Q(n17629) );
  AND2X1 U18419 ( .IN1(n9821), .IN2(WX729), .Q(n17628) );
  OR2X1 U18420 ( .IN1(n9866), .IN2(n2182), .Q(n17613) );
  OR2X1 U18421 ( .IN1(n17630), .IN2(n17631), .Q(DATA_9_20) );
  AND2X1 U18422 ( .IN1(n12859), .IN2(n17632), .Q(n17631) );
  INVX0 U18423 ( .INP(n17633), .ZN(n17630) );
  OR2X1 U18424 ( .IN1(n17632), .IN2(n12859), .Q(n17633) );
  AND2X1 U18425 ( .IN1(n17634), .IN2(n17635), .Q(n12859) );
  OR2X1 U18426 ( .IN1(n17636), .IN2(n17637), .Q(n17635) );
  INVX0 U18427 ( .INP(n17638), .ZN(n17634) );
  AND2X1 U18428 ( .IN1(n17637), .IN2(n17636), .Q(n17638) );
  AND2X1 U18429 ( .IN1(n17639), .IN2(n17640), .Q(n17636) );
  OR2X1 U18430 ( .IN1(n10537), .IN2(n3507), .Q(n17640) );
  OR2X1 U18431 ( .IN1(WX667), .IN2(n10514), .Q(n17639) );
  OR2X1 U18432 ( .IN1(n17641), .IN2(n17642), .Q(n17637) );
  AND2X1 U18433 ( .IN1(n9826), .IN2(n17643), .Q(n17642) );
  AND2X1 U18434 ( .IN1(n17644), .IN2(n17645), .Q(n17643) );
  OR2X1 U18435 ( .IN1(n9825), .IN2(n9900), .Q(n17645) );
  OR2X1 U18436 ( .IN1(test_so6), .IN2(WX859), .Q(n17644) );
  AND2X1 U18437 ( .IN1(n17646), .IN2(WX731), .Q(n17641) );
  OR2X1 U18438 ( .IN1(n17647), .IN2(n17648), .Q(n17646) );
  AND2X1 U18439 ( .IN1(n9825), .IN2(n9900), .Q(n17648) );
  AND2X1 U18440 ( .IN1(test_so6), .IN2(WX859), .Q(n17647) );
  OR2X1 U18441 ( .IN1(n9865), .IN2(n2182), .Q(n17632) );
  OR2X1 U18442 ( .IN1(n17649), .IN2(n17650), .Q(DATA_9_2) );
  AND2X1 U18443 ( .IN1(n12715), .IN2(n17651), .Q(n17650) );
  INVX0 U18444 ( .INP(n17652), .ZN(n17649) );
  OR2X1 U18445 ( .IN1(n17651), .IN2(n12715), .Q(n17652) );
  AND2X1 U18446 ( .IN1(n17653), .IN2(n17654), .Q(n12715) );
  OR2X1 U18447 ( .IN1(n17655), .IN2(n17656), .Q(n17654) );
  INVX0 U18448 ( .INP(n17657), .ZN(n17653) );
  AND2X1 U18449 ( .IN1(n17656), .IN2(n17655), .Q(n17657) );
  AND2X1 U18450 ( .IN1(n17658), .IN2(n17659), .Q(n17655) );
  OR2X1 U18451 ( .IN1(n2182), .IN2(n3471), .Q(n17659) );
  OR2X1 U18452 ( .IN1(WX703), .IN2(TM0), .Q(n17658) );
  OR2X1 U18453 ( .IN1(n17660), .IN2(n17661), .Q(n17656) );
  AND2X1 U18454 ( .IN1(n9834), .IN2(n17662), .Q(n17661) );
  AND2X1 U18455 ( .IN1(n17663), .IN2(n17664), .Q(n17662) );
  OR2X1 U18456 ( .IN1(n9833), .IN2(n9901), .Q(n17664) );
  OR2X1 U18457 ( .IN1(test_so7), .IN2(WX767), .Q(n17663) );
  AND2X1 U18458 ( .IN1(n17665), .IN2(WX895), .Q(n17660) );
  OR2X1 U18459 ( .IN1(n17666), .IN2(n17667), .Q(n17665) );
  AND2X1 U18460 ( .IN1(n9833), .IN2(n9901), .Q(n17667) );
  AND2X1 U18461 ( .IN1(test_so7), .IN2(WX767), .Q(n17666) );
  OR2X1 U18462 ( .IN1(n9864), .IN2(n2182), .Q(n17651) );
  OR2X1 U18463 ( .IN1(n17668), .IN2(n17669), .Q(DATA_9_19) );
  AND2X1 U18464 ( .IN1(n12851), .IN2(n17670), .Q(n17669) );
  INVX0 U18465 ( .INP(n17671), .ZN(n17668) );
  OR2X1 U18466 ( .IN1(n17670), .IN2(n12851), .Q(n17671) );
  OR2X1 U18467 ( .IN1(n17672), .IN2(n17673), .Q(n12851) );
  INVX0 U18468 ( .INP(n17674), .ZN(n17673) );
  OR2X1 U18469 ( .IN1(n17675), .IN2(n17676), .Q(n17674) );
  AND2X1 U18470 ( .IN1(n17676), .IN2(n17675), .Q(n17672) );
  AND2X1 U18471 ( .IN1(n17677), .IN2(n17678), .Q(n17675) );
  OR2X1 U18472 ( .IN1(n10537), .IN2(n3505), .Q(n17678) );
  OR2X1 U18473 ( .IN1(WX669), .IN2(n10514), .Q(n17677) );
  OR2X1 U18474 ( .IN1(n17679), .IN2(n17680), .Q(n17676) );
  INVX0 U18475 ( .INP(n17681), .ZN(n17680) );
  OR2X1 U18476 ( .IN1(n17682), .IN2(n9759), .Q(n17681) );
  AND2X1 U18477 ( .IN1(n9759), .IN2(n17682), .Q(n17679) );
  AND2X1 U18478 ( .IN1(n17683), .IN2(n17684), .Q(n17682) );
  OR2X1 U18479 ( .IN1(WX861), .IN2(n9761), .Q(n17684) );
  OR2X1 U18480 ( .IN1(WX733), .IN2(n9760), .Q(n17683) );
  OR2X1 U18481 ( .IN1(n9863), .IN2(n2182), .Q(n17670) );
  OR2X1 U18482 ( .IN1(n17685), .IN2(n17686), .Q(DATA_9_18) );
  AND2X1 U18483 ( .IN1(n12843), .IN2(n17687), .Q(n17686) );
  INVX0 U18484 ( .INP(n17688), .ZN(n17685) );
  OR2X1 U18485 ( .IN1(n17687), .IN2(n12843), .Q(n17688) );
  OR2X1 U18486 ( .IN1(n17689), .IN2(n17690), .Q(n12843) );
  INVX0 U18487 ( .INP(n17691), .ZN(n17690) );
  OR2X1 U18488 ( .IN1(n17692), .IN2(n17693), .Q(n17691) );
  AND2X1 U18489 ( .IN1(n17693), .IN2(n17692), .Q(n17689) );
  AND2X1 U18490 ( .IN1(n17694), .IN2(n17695), .Q(n17692) );
  OR2X1 U18491 ( .IN1(n10537), .IN2(n3503), .Q(n17695) );
  OR2X1 U18492 ( .IN1(WX671), .IN2(n10514), .Q(n17694) );
  OR2X1 U18493 ( .IN1(n17696), .IN2(n17697), .Q(n17693) );
  INVX0 U18494 ( .INP(n17698), .ZN(n17697) );
  OR2X1 U18495 ( .IN1(n17699), .IN2(n9774), .Q(n17698) );
  AND2X1 U18496 ( .IN1(n9774), .IN2(n17699), .Q(n17696) );
  AND2X1 U18497 ( .IN1(n17700), .IN2(n17701), .Q(n17699) );
  OR2X1 U18498 ( .IN1(WX863), .IN2(n9776), .Q(n17701) );
  OR2X1 U18499 ( .IN1(WX735), .IN2(n9775), .Q(n17700) );
  OR2X1 U18500 ( .IN1(n9862), .IN2(n2182), .Q(n17687) );
  OR2X1 U18501 ( .IN1(n17702), .IN2(n17703), .Q(DATA_9_17) );
  AND2X1 U18502 ( .IN1(n12835), .IN2(n17704), .Q(n17703) );
  INVX0 U18503 ( .INP(n17705), .ZN(n17702) );
  OR2X1 U18504 ( .IN1(n17704), .IN2(n12835), .Q(n17705) );
  OR2X1 U18505 ( .IN1(n17706), .IN2(n17707), .Q(n12835) );
  INVX0 U18506 ( .INP(n17708), .ZN(n17707) );
  OR2X1 U18507 ( .IN1(n17709), .IN2(n17710), .Q(n17708) );
  AND2X1 U18508 ( .IN1(n17710), .IN2(n17709), .Q(n17706) );
  AND2X1 U18509 ( .IN1(n17711), .IN2(n17712), .Q(n17709) );
  OR2X1 U18510 ( .IN1(n10537), .IN2(n3501), .Q(n17712) );
  OR2X1 U18511 ( .IN1(WX673), .IN2(n10514), .Q(n17711) );
  OR2X1 U18512 ( .IN1(n17713), .IN2(n17714), .Q(n17710) );
  INVX0 U18513 ( .INP(n17715), .ZN(n17714) );
  OR2X1 U18514 ( .IN1(n17716), .IN2(n9786), .Q(n17715) );
  AND2X1 U18515 ( .IN1(n9786), .IN2(n17716), .Q(n17713) );
  AND2X1 U18516 ( .IN1(n17717), .IN2(n17718), .Q(n17716) );
  OR2X1 U18517 ( .IN1(WX865), .IN2(n9788), .Q(n17718) );
  OR2X1 U18518 ( .IN1(WX737), .IN2(n9787), .Q(n17717) );
  OR2X1 U18519 ( .IN1(n9861), .IN2(n2182), .Q(n17704) );
  OR2X1 U18520 ( .IN1(n17719), .IN2(n17720), .Q(DATA_9_16) );
  AND2X1 U18521 ( .IN1(n12827), .IN2(n17721), .Q(n17720) );
  INVX0 U18522 ( .INP(n17722), .ZN(n17719) );
  OR2X1 U18523 ( .IN1(n17721), .IN2(n12827), .Q(n17722) );
  AND2X1 U18524 ( .IN1(n17723), .IN2(n17724), .Q(n12827) );
  OR2X1 U18525 ( .IN1(n17725), .IN2(n17726), .Q(n17724) );
  INVX0 U18526 ( .INP(n17727), .ZN(n17723) );
  AND2X1 U18527 ( .IN1(n17726), .IN2(n17725), .Q(n17727) );
  AND2X1 U18528 ( .IN1(n17728), .IN2(n17729), .Q(n17725) );
  OR2X1 U18529 ( .IN1(n10537), .IN2(n3499), .Q(n17729) );
  OR2X1 U18530 ( .IN1(WX675), .IN2(n10514), .Q(n17728) );
  OR2X1 U18531 ( .IN1(n17730), .IN2(n17731), .Q(n17726) );
  AND2X1 U18532 ( .IN1(n9804), .IN2(n17732), .Q(n17731) );
  AND2X1 U18533 ( .IN1(n17733), .IN2(n17734), .Q(n17732) );
  OR2X1 U18534 ( .IN1(n9803), .IN2(n9885), .Q(n17734) );
  OR2X1 U18535 ( .IN1(test_so8), .IN2(WX739), .Q(n17733) );
  AND2X1 U18536 ( .IN1(n17735), .IN2(WX803), .Q(n17730) );
  OR2X1 U18537 ( .IN1(n17736), .IN2(n17737), .Q(n17735) );
  AND2X1 U18538 ( .IN1(n9803), .IN2(n9885), .Q(n17737) );
  AND2X1 U18539 ( .IN1(test_so8), .IN2(WX739), .Q(n17736) );
  OR2X1 U18540 ( .IN1(n9860), .IN2(n2182), .Q(n17721) );
  OR2X1 U18541 ( .IN1(n17738), .IN2(n17739), .Q(DATA_9_15) );
  AND2X1 U18542 ( .IN1(n12819), .IN2(n17740), .Q(n17739) );
  INVX0 U18543 ( .INP(n17741), .ZN(n17738) );
  OR2X1 U18544 ( .IN1(n17740), .IN2(n12819), .Q(n17741) );
  OR2X1 U18545 ( .IN1(n17742), .IN2(n17743), .Q(n12819) );
  INVX0 U18546 ( .INP(n17744), .ZN(n17743) );
  OR2X1 U18547 ( .IN1(n17745), .IN2(n17746), .Q(n17744) );
  AND2X1 U18548 ( .IN1(n17746), .IN2(n17745), .Q(n17742) );
  AND2X1 U18549 ( .IN1(n17747), .IN2(n17748), .Q(n17745) );
  OR2X1 U18550 ( .IN1(n2182), .IN2(n3497), .Q(n17748) );
  OR2X1 U18551 ( .IN1(WX677), .IN2(TM0), .Q(n17747) );
  OR2X1 U18552 ( .IN1(n17749), .IN2(n17750), .Q(n17746) );
  AND2X1 U18553 ( .IN1(n9819), .IN2(n17751), .Q(n17750) );
  AND2X1 U18554 ( .IN1(n17752), .IN2(n17753), .Q(n17751) );
  OR2X1 U18555 ( .IN1(n9817), .IN2(WX805), .Q(n17753) );
  OR2X1 U18556 ( .IN1(n9818), .IN2(WX741), .Q(n17752) );
  AND2X1 U18557 ( .IN1(n17754), .IN2(WX869), .Q(n17749) );
  OR2X1 U18558 ( .IN1(n17755), .IN2(n17756), .Q(n17754) );
  AND2X1 U18559 ( .IN1(n9817), .IN2(WX805), .Q(n17756) );
  AND2X1 U18560 ( .IN1(n9818), .IN2(WX741), .Q(n17755) );
  OR2X1 U18561 ( .IN1(n9859), .IN2(n2182), .Q(n17740) );
  OR2X1 U18562 ( .IN1(n17757), .IN2(n17758), .Q(DATA_9_14) );
  AND2X1 U18563 ( .IN1(n12811), .IN2(n17759), .Q(n17758) );
  INVX0 U18564 ( .INP(n17760), .ZN(n17757) );
  OR2X1 U18565 ( .IN1(n17759), .IN2(n12811), .Q(n17760) );
  OR2X1 U18566 ( .IN1(n17761), .IN2(n17762), .Q(n12811) );
  INVX0 U18567 ( .INP(n17763), .ZN(n17762) );
  OR2X1 U18568 ( .IN1(n17764), .IN2(n17765), .Q(n17763) );
  AND2X1 U18569 ( .IN1(n17765), .IN2(n17764), .Q(n17761) );
  AND2X1 U18570 ( .IN1(n17766), .IN2(n17767), .Q(n17764) );
  OR2X1 U18571 ( .IN1(n2182), .IN2(n3495), .Q(n17767) );
  OR2X1 U18572 ( .IN1(WX679), .IN2(TM0), .Q(n17766) );
  OR2X1 U18573 ( .IN1(n17768), .IN2(n17769), .Q(n17765) );
  INVX0 U18574 ( .INP(n17770), .ZN(n17769) );
  OR2X1 U18575 ( .IN1(n17771), .IN2(n9830), .Q(n17770) );
  AND2X1 U18576 ( .IN1(n9830), .IN2(n17771), .Q(n17768) );
  AND2X1 U18577 ( .IN1(n17772), .IN2(n17773), .Q(n17771) );
  OR2X1 U18578 ( .IN1(WX871), .IN2(n9832), .Q(n17773) );
  OR2X1 U18579 ( .IN1(WX743), .IN2(n9831), .Q(n17772) );
  OR2X1 U18580 ( .IN1(n2182), .IN2(n9858), .Q(n17759) );
  OR2X1 U18581 ( .IN1(n17774), .IN2(n17775), .Q(DATA_9_13) );
  AND2X1 U18582 ( .IN1(n12803), .IN2(n17776), .Q(n17775) );
  INVX0 U18583 ( .INP(n17777), .ZN(n17774) );
  OR2X1 U18584 ( .IN1(n17776), .IN2(n12803), .Q(n17777) );
  OR2X1 U18585 ( .IN1(n17778), .IN2(n17779), .Q(n12803) );
  INVX0 U18586 ( .INP(n17780), .ZN(n17779) );
  OR2X1 U18587 ( .IN1(n17781), .IN2(n17782), .Q(n17780) );
  AND2X1 U18588 ( .IN1(n17782), .IN2(n17781), .Q(n17778) );
  AND2X1 U18589 ( .IN1(n17783), .IN2(n17784), .Q(n17781) );
  OR2X1 U18590 ( .IN1(n2182), .IN2(n3493), .Q(n17784) );
  OR2X1 U18591 ( .IN1(WX681), .IN2(TM0), .Q(n17783) );
  OR2X1 U18592 ( .IN1(n17785), .IN2(n17786), .Q(n17782) );
  INVX0 U18593 ( .INP(n17787), .ZN(n17786) );
  OR2X1 U18594 ( .IN1(n17788), .IN2(n9765), .Q(n17787) );
  AND2X1 U18595 ( .IN1(n9765), .IN2(n17788), .Q(n17785) );
  AND2X1 U18596 ( .IN1(n17789), .IN2(n17790), .Q(n17788) );
  OR2X1 U18597 ( .IN1(WX873), .IN2(n9767), .Q(n17790) );
  OR2X1 U18598 ( .IN1(WX745), .IN2(n9766), .Q(n17789) );
  OR2X1 U18599 ( .IN1(n9857), .IN2(n2182), .Q(n17776) );
  OR2X1 U18600 ( .IN1(n17791), .IN2(n17792), .Q(DATA_9_12) );
  AND2X1 U18601 ( .IN1(n12795), .IN2(n17793), .Q(n17792) );
  INVX0 U18602 ( .INP(n17794), .ZN(n17791) );
  OR2X1 U18603 ( .IN1(n17793), .IN2(n12795), .Q(n17794) );
  OR2X1 U18604 ( .IN1(n17795), .IN2(n17796), .Q(n12795) );
  INVX0 U18605 ( .INP(n17797), .ZN(n17796) );
  OR2X1 U18606 ( .IN1(n17798), .IN2(n17799), .Q(n17797) );
  AND2X1 U18607 ( .IN1(n17799), .IN2(n17798), .Q(n17795) );
  AND2X1 U18608 ( .IN1(n17800), .IN2(n17801), .Q(n17798) );
  OR2X1 U18609 ( .IN1(n2182), .IN2(n3491), .Q(n17801) );
  OR2X1 U18610 ( .IN1(WX683), .IN2(TM0), .Q(n17800) );
  OR2X1 U18611 ( .IN1(n17802), .IN2(n17803), .Q(n17799) );
  INVX0 U18612 ( .INP(n17804), .ZN(n17803) );
  OR2X1 U18613 ( .IN1(n17805), .IN2(n9792), .Q(n17804) );
  AND2X1 U18614 ( .IN1(n9792), .IN2(n17805), .Q(n17802) );
  AND2X1 U18615 ( .IN1(n17806), .IN2(n17807), .Q(n17805) );
  OR2X1 U18616 ( .IN1(WX875), .IN2(n9794), .Q(n17807) );
  OR2X1 U18617 ( .IN1(WX747), .IN2(n9793), .Q(n17806) );
  OR2X1 U18618 ( .IN1(n9856), .IN2(n2182), .Q(n17793) );
  OR2X1 U18619 ( .IN1(n17808), .IN2(n17809), .Q(DATA_9_11) );
  AND2X1 U18620 ( .IN1(n12787), .IN2(n17810), .Q(n17809) );
  INVX0 U18621 ( .INP(n17811), .ZN(n17808) );
  OR2X1 U18622 ( .IN1(n17810), .IN2(n12787), .Q(n17811) );
  OR2X1 U18623 ( .IN1(n17812), .IN2(n17813), .Q(n12787) );
  INVX0 U18624 ( .INP(n17814), .ZN(n17813) );
  OR2X1 U18625 ( .IN1(n17815), .IN2(n17816), .Q(n17814) );
  AND2X1 U18626 ( .IN1(n17816), .IN2(n17815), .Q(n17812) );
  AND2X1 U18627 ( .IN1(n17817), .IN2(n17818), .Q(n17815) );
  OR2X1 U18628 ( .IN1(n2182), .IN2(n3489), .Q(n17818) );
  OR2X1 U18629 ( .IN1(WX685), .IN2(TM0), .Q(n17817) );
  OR2X1 U18630 ( .IN1(n17819), .IN2(n17820), .Q(n17816) );
  INVX0 U18631 ( .INP(n17821), .ZN(n17820) );
  OR2X1 U18632 ( .IN1(n17822), .IN2(n9838), .Q(n17821) );
  AND2X1 U18633 ( .IN1(n9838), .IN2(n17822), .Q(n17819) );
  AND2X1 U18634 ( .IN1(n17823), .IN2(n17824), .Q(n17822) );
  OR2X1 U18635 ( .IN1(WX877), .IN2(n9840), .Q(n17824) );
  OR2X1 U18636 ( .IN1(WX749), .IN2(n9839), .Q(n17823) );
  OR2X1 U18637 ( .IN1(n9855), .IN2(n2182), .Q(n17810) );
  OR2X1 U18638 ( .IN1(n17825), .IN2(n17826), .Q(DATA_9_10) );
  AND2X1 U18639 ( .IN1(n12779), .IN2(n17827), .Q(n17826) );
  INVX0 U18640 ( .INP(n17828), .ZN(n17825) );
  OR2X1 U18641 ( .IN1(n17827), .IN2(n12779), .Q(n17828) );
  AND2X1 U18642 ( .IN1(n17829), .IN2(n17830), .Q(n12779) );
  OR2X1 U18643 ( .IN1(n17831), .IN2(n17832), .Q(n17830) );
  INVX0 U18644 ( .INP(n17833), .ZN(n17829) );
  AND2X1 U18645 ( .IN1(n17832), .IN2(n17831), .Q(n17833) );
  AND2X1 U18646 ( .IN1(n17834), .IN2(n17835), .Q(n17831) );
  OR2X1 U18647 ( .IN1(n2182), .IN2(n9785), .Q(n17835) );
  OR2X1 U18648 ( .IN1(WX751), .IN2(TM0), .Q(n17834) );
  OR2X1 U18649 ( .IN1(n17836), .IN2(n17837), .Q(n17832) );
  AND2X1 U18650 ( .IN1(n9784), .IN2(n17838), .Q(n17837) );
  AND2X1 U18651 ( .IN1(n17839), .IN2(n17840), .Q(n17838) );
  OR2X1 U18652 ( .IN1(n9783), .IN2(n9902), .Q(n17840) );
  OR2X1 U18653 ( .IN1(test_so3), .IN2(WX815), .Q(n17839) );
  AND2X1 U18654 ( .IN1(n17841), .IN2(WX879), .Q(n17836) );
  OR2X1 U18655 ( .IN1(n17842), .IN2(n17843), .Q(n17841) );
  AND2X1 U18656 ( .IN1(n9783), .IN2(n9902), .Q(n17843) );
  AND2X1 U18657 ( .IN1(test_so3), .IN2(WX815), .Q(n17842) );
  OR2X1 U18658 ( .IN1(n9854), .IN2(n2182), .Q(n17827) );
  OR2X1 U18659 ( .IN1(n17844), .IN2(n17845), .Q(DATA_9_1) );
  AND2X1 U18660 ( .IN1(n12707), .IN2(n17846), .Q(n17845) );
  INVX0 U18661 ( .INP(n17847), .ZN(n17844) );
  OR2X1 U18662 ( .IN1(n17846), .IN2(n12707), .Q(n17847) );
  OR2X1 U18663 ( .IN1(n17848), .IN2(n17849), .Q(n12707) );
  AND2X1 U18664 ( .IN1(n17850), .IN2(n17851), .Q(n17849) );
  INVX0 U18665 ( .INP(n17852), .ZN(n17848) );
  OR2X1 U18666 ( .IN1(n17851), .IN2(n17850), .Q(n17852) );
  OR2X1 U18667 ( .IN1(n17853), .IN2(n17854), .Q(n17850) );
  AND2X1 U18668 ( .IN1(TM0), .IN2(WX705), .Q(n17854) );
  AND2X1 U18669 ( .IN1(n3469), .IN2(n2182), .Q(n17853) );
  AND2X1 U18670 ( .IN1(n17855), .IN2(n17856), .Q(n17851) );
  OR2X1 U18671 ( .IN1(n17857), .IN2(n9768), .Q(n17856) );
  INVX0 U18672 ( .INP(n17858), .ZN(n17855) );
  AND2X1 U18673 ( .IN1(n9768), .IN2(n17857), .Q(n17858) );
  AND2X1 U18674 ( .IN1(n17859), .IN2(n17860), .Q(n17857) );
  OR2X1 U18675 ( .IN1(WX769), .IN2(n9770), .Q(n17860) );
  INVX0 U18676 ( .INP(n17861), .ZN(n17859) );
  AND2X1 U18677 ( .IN1(n9770), .IN2(WX769), .Q(n17861) );
  OR2X1 U18678 ( .IN1(n9853), .IN2(n2182), .Q(n17846) );
  OR2X1 U18679 ( .IN1(n17862), .IN2(n17863), .Q(DATA_9_0) );
  AND2X1 U18680 ( .IN1(n12699), .IN2(n17864), .Q(n17863) );
  INVX0 U18681 ( .INP(n17865), .ZN(n17862) );
  OR2X1 U18682 ( .IN1(n17864), .IN2(n12699), .Q(n17865) );
  OR2X1 U18683 ( .IN1(n17866), .IN2(n17867), .Q(n12699) );
  INVX0 U18684 ( .INP(n17868), .ZN(n17867) );
  OR2X1 U18685 ( .IN1(n17869), .IN2(n17870), .Q(n17868) );
  AND2X1 U18686 ( .IN1(n17870), .IN2(n17869), .Q(n17866) );
  AND2X1 U18687 ( .IN1(n17871), .IN2(n17872), .Q(n17869) );
  OR2X1 U18688 ( .IN1(n2182), .IN2(n3467), .Q(n17872) );
  OR2X1 U18689 ( .IN1(WX707), .IN2(TM0), .Q(n17871) );
  OR2X1 U18690 ( .IN1(n17873), .IN2(n17874), .Q(n17870) );
  AND2X1 U18691 ( .IN1(n9843), .IN2(n17875), .Q(n17874) );
  AND2X1 U18692 ( .IN1(n17876), .IN2(n17877), .Q(n17875) );
  OR2X1 U18693 ( .IN1(n9841), .IN2(WX835), .Q(n17877) );
  OR2X1 U18694 ( .IN1(n9842), .IN2(WX771), .Q(n17876) );
  AND2X1 U18695 ( .IN1(n17878), .IN2(WX899), .Q(n17873) );
  OR2X1 U18696 ( .IN1(n17879), .IN2(n17880), .Q(n17878) );
  AND2X1 U18697 ( .IN1(n9841), .IN2(WX835), .Q(n17880) );
  AND2X1 U18698 ( .IN1(n9842), .IN2(WX771), .Q(n17879) );
  OR2X1 U18699 ( .IN1(n9852), .IN2(n2182), .Q(n17864) );
  AND2X1 U3558_U2 ( .IN1(n10023), .IN2(U3558_n1), .Q(n2245) );
  INVX0 U3558_U1 ( .INP(n10649), .ZN(U3558_n1) );
  INVX0 U3871_U2 ( .INP(TM0), .ZN(U3871_n1) );
  AND2X1 U3871_U1 ( .IN1(n3278), .IN2(U3871_n1), .Q(n2153) );
  INVX0 U3991_U2 ( .INP(n2182), .ZN(U3991_n1) );
  AND2X1 U3991_U1 ( .IN1(n3278), .IN2(U3991_n1), .Q(n2152) );
  AND2X1 U5716_U2 ( .IN1(WX547), .IN2(U5716_n1), .Q(WX544) );
  INVX0 U5716_U1 ( .INP(n10704), .ZN(U5716_n1) );
  AND2X1 U5717_U2 ( .IN1(WX545), .IN2(U5717_n1), .Q(WX542) );
  INVX0 U5717_U1 ( .INP(n10704), .ZN(U5717_n1) );
  AND2X1 U5718_U2 ( .IN1(WX543), .IN2(U5718_n1), .Q(WX540) );
  INVX0 U5718_U1 ( .INP(n10704), .ZN(U5718_n1) );
  AND2X1 U5719_U2 ( .IN1(WX541), .IN2(U5719_n1), .Q(WX538) );
  INVX0 U5719_U1 ( .INP(n10704), .ZN(U5719_n1) );
  AND2X1 U5720_U2 ( .IN1(WX539), .IN2(U5720_n1), .Q(WX536) );
  INVX0 U5720_U1 ( .INP(n10704), .ZN(U5720_n1) );
  AND2X1 U5721_U2 ( .IN1(WX537), .IN2(U5721_n1), .Q(WX534) );
  INVX0 U5721_U1 ( .INP(n10704), .ZN(U5721_n1) );
  AND2X1 U5722_U2 ( .IN1(WX535), .IN2(U5722_n1), .Q(WX532) );
  INVX0 U5722_U1 ( .INP(n10704), .ZN(U5722_n1) );
  AND2X1 U5723_U2 ( .IN1(WX533), .IN2(U5723_n1), .Q(WX530) );
  INVX0 U5723_U1 ( .INP(n10704), .ZN(U5723_n1) );
  AND2X1 U5724_U2 ( .IN1(WX531), .IN2(U5724_n1), .Q(WX528) );
  INVX0 U5724_U1 ( .INP(n10703), .ZN(U5724_n1) );
  AND2X1 U5725_U2 ( .IN1(WX529), .IN2(U5725_n1), .Q(WX526) );
  INVX0 U5725_U1 ( .INP(n10703), .ZN(U5725_n1) );
  AND2X1 U5726_U2 ( .IN1(WX527), .IN2(U5726_n1), .Q(WX524) );
  INVX0 U5726_U1 ( .INP(n10703), .ZN(U5726_n1) );
  AND2X1 U5727_U2 ( .IN1(WX525), .IN2(U5727_n1), .Q(WX522) );
  INVX0 U5727_U1 ( .INP(n10703), .ZN(U5727_n1) );
  AND2X1 U5728_U2 ( .IN1(WX523), .IN2(U5728_n1), .Q(WX520) );
  INVX0 U5728_U1 ( .INP(n10703), .ZN(U5728_n1) );
  AND2X1 U5729_U2 ( .IN1(WX521), .IN2(U5729_n1), .Q(WX518) );
  INVX0 U5729_U1 ( .INP(n10703), .ZN(U5729_n1) );
  AND2X1 U5730_U2 ( .IN1(test_so1), .IN2(U5730_n1), .Q(WX516) );
  INVX0 U5730_U1 ( .INP(n10703), .ZN(U5730_n1) );
  AND2X1 U5731_U2 ( .IN1(WX517), .IN2(U5731_n1), .Q(WX514) );
  INVX0 U5731_U1 ( .INP(n10703), .ZN(U5731_n1) );
  AND2X1 U5732_U2 ( .IN1(WX515), .IN2(U5732_n1), .Q(WX512) );
  INVX0 U5732_U1 ( .INP(n10703), .ZN(U5732_n1) );
  AND2X1 U5733_U2 ( .IN1(WX513), .IN2(U5733_n1), .Q(WX510) );
  INVX0 U5733_U1 ( .INP(n10703), .ZN(U5733_n1) );
  AND2X1 U5734_U2 ( .IN1(WX511), .IN2(U5734_n1), .Q(WX508) );
  INVX0 U5734_U1 ( .INP(n10703), .ZN(U5734_n1) );
  AND2X1 U5735_U2 ( .IN1(WX509), .IN2(U5735_n1), .Q(WX506) );
  INVX0 U5735_U1 ( .INP(n10703), .ZN(U5735_n1) );
  AND2X1 U5736_U2 ( .IN1(WX507), .IN2(U5736_n1), .Q(WX504) );
  INVX0 U5736_U1 ( .INP(n10703), .ZN(U5736_n1) );
  AND2X1 U5737_U2 ( .IN1(WX505), .IN2(U5737_n1), .Q(WX502) );
  INVX0 U5737_U1 ( .INP(n10703), .ZN(U5737_n1) );
  AND2X1 U5738_U2 ( .IN1(WX503), .IN2(U5738_n1), .Q(WX500) );
  INVX0 U5738_U1 ( .INP(n10702), .ZN(U5738_n1) );
  AND2X1 U5739_U2 ( .IN1(WX501), .IN2(U5739_n1), .Q(WX498) );
  INVX0 U5739_U1 ( .INP(n10702), .ZN(U5739_n1) );
  AND2X1 U5740_U2 ( .IN1(WX499), .IN2(U5740_n1), .Q(WX496) );
  INVX0 U5740_U1 ( .INP(n10702), .ZN(U5740_n1) );
  AND2X1 U5741_U2 ( .IN1(WX497), .IN2(U5741_n1), .Q(WX494) );
  INVX0 U5741_U1 ( .INP(n10702), .ZN(U5741_n1) );
  AND2X1 U5742_U2 ( .IN1(WX495), .IN2(U5742_n1), .Q(WX492) );
  INVX0 U5742_U1 ( .INP(n10702), .ZN(U5742_n1) );
  AND2X1 U5743_U2 ( .IN1(WX493), .IN2(U5743_n1), .Q(WX490) );
  INVX0 U5743_U1 ( .INP(n10702), .ZN(U5743_n1) );
  AND2X1 U5744_U2 ( .IN1(WX491), .IN2(U5744_n1), .Q(WX488) );
  INVX0 U5744_U1 ( .INP(n10702), .ZN(U5744_n1) );
  AND2X1 U5745_U2 ( .IN1(WX489), .IN2(U5745_n1), .Q(WX486) );
  INVX0 U5745_U1 ( .INP(n10702), .ZN(U5745_n1) );
  AND2X1 U5746_U2 ( .IN1(WX487), .IN2(U5746_n1), .Q(WX484) );
  INVX0 U5746_U1 ( .INP(n10702), .ZN(U5746_n1) );
  AND2X1 U5747_U2 ( .IN1(WX5939), .IN2(U5747_n1), .Q(WX6002) );
  INVX0 U5747_U1 ( .INP(n10702), .ZN(U5747_n1) );
  AND2X1 U5748_U2 ( .IN1(test_so49), .IN2(U5748_n1), .Q(WX6000) );
  INVX0 U5748_U1 ( .INP(n10702), .ZN(U5748_n1) );
  AND2X1 U5749_U2 ( .IN1(WX5935), .IN2(U5749_n1), .Q(WX5998) );
  INVX0 U5749_U1 ( .INP(n10702), .ZN(U5749_n1) );
  AND2X1 U5750_U2 ( .IN1(WX5933), .IN2(U5750_n1), .Q(WX5996) );
  INVX0 U5750_U1 ( .INP(n10702), .ZN(U5750_n1) );
  AND2X1 U5751_U2 ( .IN1(WX5931), .IN2(U5751_n1), .Q(WX5994) );
  INVX0 U5751_U1 ( .INP(n10702), .ZN(U5751_n1) );
  AND2X1 U5752_U2 ( .IN1(WX3269), .IN2(U5752_n1), .Q(WX3332) );
  INVX0 U5752_U1 ( .INP(n10701), .ZN(U5752_n1) );
  AND2X1 U5753_U2 ( .IN1(WX3265), .IN2(U5753_n1), .Q(WX3328) );
  INVX0 U5753_U1 ( .INP(n10701), .ZN(U5753_n1) );
  AND2X1 U5754_U2 ( .IN1(WX3263), .IN2(U5754_n1), .Q(WX3326) );
  INVX0 U5754_U1 ( .INP(n10701), .ZN(U5754_n1) );
  AND2X1 U5755_U2 ( .IN1(WX11179), .IN2(U5755_n1), .Q(WX11242) );
  INVX0 U5755_U1 ( .INP(n10701), .ZN(U5755_n1) );
  AND2X1 U5756_U2 ( .IN1(WX11177), .IN2(U5756_n1), .Q(WX11240) );
  INVX0 U5756_U1 ( .INP(n10701), .ZN(U5756_n1) );
  AND2X1 U5757_U2 ( .IN1(WX11175), .IN2(U5757_n1), .Q(WX11238) );
  INVX0 U5757_U1 ( .INP(n10701), .ZN(U5757_n1) );
  AND2X1 U5758_U2 ( .IN1(WX11173), .IN2(U5758_n1), .Q(WX11236) );
  INVX0 U5758_U1 ( .INP(n10701), .ZN(U5758_n1) );
  AND2X1 U5759_U2 ( .IN1(test_so96), .IN2(U5759_n1), .Q(WX11234) );
  INVX0 U5759_U1 ( .INP(n10701), .ZN(U5759_n1) );
  AND2X1 U5760_U2 ( .IN1(WX11169), .IN2(U5760_n1), .Q(WX11232) );
  INVX0 U5760_U1 ( .INP(n10701), .ZN(U5760_n1) );
  AND2X1 U5761_U2 ( .IN1(WX11167), .IN2(U5761_n1), .Q(WX11230) );
  INVX0 U5761_U1 ( .INP(n10701), .ZN(U5761_n1) );
  AND2X1 U5762_U2 ( .IN1(WX11165), .IN2(U5762_n1), .Q(WX11228) );
  INVX0 U5762_U1 ( .INP(n10701), .ZN(U5762_n1) );
  AND2X1 U5763_U2 ( .IN1(WX11163), .IN2(U5763_n1), .Q(WX11226) );
  INVX0 U5763_U1 ( .INP(n10701), .ZN(U5763_n1) );
  AND2X1 U5764_U2 ( .IN1(WX11161), .IN2(U5764_n1), .Q(WX11224) );
  INVX0 U5764_U1 ( .INP(n10701), .ZN(U5764_n1) );
  AND2X1 U5765_U2 ( .IN1(WX11159), .IN2(U5765_n1), .Q(WX11222) );
  INVX0 U5765_U1 ( .INP(n10701), .ZN(U5765_n1) );
  AND2X1 U5766_U2 ( .IN1(WX11157), .IN2(U5766_n1), .Q(WX11220) );
  INVX0 U5766_U1 ( .INP(n10700), .ZN(U5766_n1) );
  AND2X1 U5767_U2 ( .IN1(WX11155), .IN2(U5767_n1), .Q(WX11218) );
  INVX0 U5767_U1 ( .INP(n10700), .ZN(U5767_n1) );
  AND2X1 U5768_U2 ( .IN1(WX11153), .IN2(U5768_n1), .Q(WX11216) );
  INVX0 U5768_U1 ( .INP(n10700), .ZN(U5768_n1) );
  AND2X1 U5769_U2 ( .IN1(WX11151), .IN2(U5769_n1), .Q(WX11214) );
  INVX0 U5769_U1 ( .INP(n10700), .ZN(U5769_n1) );
  AND2X1 U5770_U2 ( .IN1(WX11149), .IN2(U5770_n1), .Q(WX11212) );
  INVX0 U5770_U1 ( .INP(n10700), .ZN(U5770_n1) );
  AND2X1 U5771_U2 ( .IN1(WX11147), .IN2(U5771_n1), .Q(WX11210) );
  INVX0 U5771_U1 ( .INP(n10700), .ZN(U5771_n1) );
  AND2X1 U5772_U2 ( .IN1(WX11145), .IN2(U5772_n1), .Q(WX11208) );
  INVX0 U5772_U1 ( .INP(n10700), .ZN(U5772_n1) );
  AND2X1 U5773_U2 ( .IN1(WX11143), .IN2(U5773_n1), .Q(WX11206) );
  INVX0 U5773_U1 ( .INP(n10700), .ZN(U5773_n1) );
  AND2X1 U5774_U2 ( .IN1(WX11141), .IN2(U5774_n1), .Q(WX11204) );
  INVX0 U5774_U1 ( .INP(n10700), .ZN(U5774_n1) );
  AND2X1 U5775_U2 ( .IN1(WX11139), .IN2(U5775_n1), .Q(WX11202) );
  INVX0 U5775_U1 ( .INP(n10700), .ZN(U5775_n1) );
  AND2X1 U5776_U2 ( .IN1(test_so95), .IN2(U5776_n1), .Q(WX11200) );
  INVX0 U5776_U1 ( .INP(n10700), .ZN(U5776_n1) );
  AND2X1 U5777_U2 ( .IN1(WX11135), .IN2(U5777_n1), .Q(WX11198) );
  INVX0 U5777_U1 ( .INP(n10700), .ZN(U5777_n1) );
  AND2X1 U5778_U2 ( .IN1(WX11133), .IN2(U5778_n1), .Q(WX11196) );
  INVX0 U5778_U1 ( .INP(n10700), .ZN(U5778_n1) );
  AND2X1 U5779_U2 ( .IN1(WX11131), .IN2(U5779_n1), .Q(WX11194) );
  INVX0 U5779_U1 ( .INP(n10700), .ZN(U5779_n1) );
  AND2X1 U5780_U2 ( .IN1(WX11129), .IN2(U5780_n1), .Q(WX11192) );
  INVX0 U5780_U1 ( .INP(n10699), .ZN(U5780_n1) );
  AND2X1 U5781_U2 ( .IN1(WX11127), .IN2(U5781_n1), .Q(WX11190) );
  INVX0 U5781_U1 ( .INP(n10699), .ZN(U5781_n1) );
  AND2X1 U5782_U2 ( .IN1(WX11125), .IN2(U5782_n1), .Q(WX11188) );
  INVX0 U5782_U1 ( .INP(n10699), .ZN(U5782_n1) );
  AND2X1 U5783_U2 ( .IN1(WX11123), .IN2(U5783_n1), .Q(WX11186) );
  INVX0 U5783_U1 ( .INP(n10699), .ZN(U5783_n1) );
  AND2X1 U5784_U2 ( .IN1(WX11121), .IN2(U5784_n1), .Q(WX11184) );
  INVX0 U5784_U1 ( .INP(n10699), .ZN(U5784_n1) );
  AND2X1 U5785_U2 ( .IN1(WX11119), .IN2(U5785_n1), .Q(WX11182) );
  INVX0 U5785_U1 ( .INP(n10699), .ZN(U5785_n1) );
  AND2X1 U5786_U2 ( .IN1(WX11117), .IN2(U5786_n1), .Q(WX11180) );
  INVX0 U5786_U1 ( .INP(n10699), .ZN(U5786_n1) );
  AND2X1 U5787_U2 ( .IN1(WX11115), .IN2(U5787_n1), .Q(WX11178) );
  INVX0 U5787_U1 ( .INP(n10699), .ZN(U5787_n1) );
  AND2X1 U5788_U2 ( .IN1(WX11113), .IN2(U5788_n1), .Q(WX11176) );
  INVX0 U5788_U1 ( .INP(n10699), .ZN(U5788_n1) );
  AND2X1 U5789_U2 ( .IN1(WX11111), .IN2(U5789_n1), .Q(WX11174) );
  INVX0 U5789_U1 ( .INP(n10699), .ZN(U5789_n1) );
  AND2X1 U5790_U2 ( .IN1(WX11109), .IN2(U5790_n1), .Q(WX11172) );
  INVX0 U5790_U1 ( .INP(n10699), .ZN(U5790_n1) );
  AND2X1 U5791_U2 ( .IN1(WX11107), .IN2(U5791_n1), .Q(WX11170) );
  INVX0 U5791_U1 ( .INP(n10699), .ZN(U5791_n1) );
  AND2X1 U5792_U2 ( .IN1(WX11105), .IN2(U5792_n1), .Q(WX11168) );
  INVX0 U5792_U1 ( .INP(n10699), .ZN(U5792_n1) );
  AND2X1 U5793_U2 ( .IN1(test_so94), .IN2(U5793_n1), .Q(WX11166) );
  INVX0 U5793_U1 ( .INP(n10699), .ZN(U5793_n1) );
  AND2X1 U5794_U2 ( .IN1(WX11101), .IN2(U5794_n1), .Q(WX11164) );
  INVX0 U5794_U1 ( .INP(n10698), .ZN(U5794_n1) );
  AND2X1 U5795_U2 ( .IN1(WX11099), .IN2(U5795_n1), .Q(WX11162) );
  INVX0 U5795_U1 ( .INP(n10698), .ZN(U5795_n1) );
  AND2X1 U5796_U2 ( .IN1(WX11097), .IN2(U5796_n1), .Q(WX11160) );
  INVX0 U5796_U1 ( .INP(n10698), .ZN(U5796_n1) );
  AND2X1 U5797_U2 ( .IN1(WX11095), .IN2(U5797_n1), .Q(WX11158) );
  INVX0 U5797_U1 ( .INP(n10698), .ZN(U5797_n1) );
  AND2X1 U5798_U2 ( .IN1(WX11093), .IN2(U5798_n1), .Q(WX11156) );
  INVX0 U5798_U1 ( .INP(n10698), .ZN(U5798_n1) );
  AND2X1 U5799_U2 ( .IN1(WX11091), .IN2(U5799_n1), .Q(WX11154) );
  INVX0 U5799_U1 ( .INP(n10698), .ZN(U5799_n1) );
  AND2X1 U5800_U2 ( .IN1(WX11089), .IN2(U5800_n1), .Q(WX11152) );
  INVX0 U5800_U1 ( .INP(n10698), .ZN(U5800_n1) );
  AND2X1 U5801_U2 ( .IN1(WX11087), .IN2(U5801_n1), .Q(WX11150) );
  INVX0 U5801_U1 ( .INP(n10698), .ZN(U5801_n1) );
  AND2X1 U5802_U2 ( .IN1(WX11085), .IN2(U5802_n1), .Q(WX11148) );
  INVX0 U5802_U1 ( .INP(n10698), .ZN(U5802_n1) );
  AND2X1 U5803_U2 ( .IN1(WX11083), .IN2(U5803_n1), .Q(WX11146) );
  INVX0 U5803_U1 ( .INP(n10698), .ZN(U5803_n1) );
  AND2X1 U5804_U2 ( .IN1(WX11081), .IN2(U5804_n1), .Q(WX11144) );
  INVX0 U5804_U1 ( .INP(n10698), .ZN(U5804_n1) );
  AND2X1 U5805_U2 ( .IN1(WX11079), .IN2(U5805_n1), .Q(WX11142) );
  INVX0 U5805_U1 ( .INP(n10698), .ZN(U5805_n1) );
  AND2X1 U5806_U2 ( .IN1(WX11077), .IN2(U5806_n1), .Q(WX11140) );
  INVX0 U5806_U1 ( .INP(n10698), .ZN(U5806_n1) );
  AND2X1 U5807_U2 ( .IN1(WX11075), .IN2(U5807_n1), .Q(WX11138) );
  INVX0 U5807_U1 ( .INP(n10698), .ZN(U5807_n1) );
  AND2X1 U5808_U2 ( .IN1(WX11073), .IN2(U5808_n1), .Q(WX11136) );
  INVX0 U5808_U1 ( .INP(n10697), .ZN(U5808_n1) );
  AND2X1 U5809_U2 ( .IN1(WX11071), .IN2(U5809_n1), .Q(WX11134) );
  INVX0 U5809_U1 ( .INP(n10697), .ZN(U5809_n1) );
  AND2X1 U5810_U2 ( .IN1(test_so93), .IN2(U5810_n1), .Q(WX11132) );
  INVX0 U5810_U1 ( .INP(n10697), .ZN(U5810_n1) );
  AND2X1 U5811_U2 ( .IN1(WX11067), .IN2(U5811_n1), .Q(WX11130) );
  INVX0 U5811_U1 ( .INP(n10697), .ZN(U5811_n1) );
  AND2X1 U5812_U2 ( .IN1(WX11065), .IN2(U5812_n1), .Q(WX11128) );
  INVX0 U5812_U1 ( .INP(n10697), .ZN(U5812_n1) );
  AND2X1 U5813_U2 ( .IN1(WX11063), .IN2(U5813_n1), .Q(WX11126) );
  INVX0 U5813_U1 ( .INP(n10697), .ZN(U5813_n1) );
  AND2X1 U5814_U2 ( .IN1(WX11061), .IN2(U5814_n1), .Q(WX11124) );
  INVX0 U5814_U1 ( .INP(n10697), .ZN(U5814_n1) );
  AND2X1 U5815_U2 ( .IN1(WX11059), .IN2(U5815_n1), .Q(WX11122) );
  INVX0 U5815_U1 ( .INP(n10697), .ZN(U5815_n1) );
  AND2X1 U5816_U2 ( .IN1(WX11057), .IN2(U5816_n1), .Q(WX11120) );
  INVX0 U5816_U1 ( .INP(n10697), .ZN(U5816_n1) );
  AND2X1 U5817_U2 ( .IN1(WX11055), .IN2(U5817_n1), .Q(WX11118) );
  INVX0 U5817_U1 ( .INP(n10697), .ZN(U5817_n1) );
  AND2X1 U5818_U2 ( .IN1(WX11053), .IN2(U5818_n1), .Q(WX11116) );
  INVX0 U5818_U1 ( .INP(n10697), .ZN(U5818_n1) );
  AND2X1 U5819_U2 ( .IN1(WX11051), .IN2(U5819_n1), .Q(WX11114) );
  INVX0 U5819_U1 ( .INP(n10697), .ZN(U5819_n1) );
  AND2X1 U5820_U2 ( .IN1(WX11049), .IN2(U5820_n1), .Q(WX11112) );
  INVX0 U5820_U1 ( .INP(n10697), .ZN(U5820_n1) );
  AND2X1 U5821_U2 ( .IN1(WX11047), .IN2(U5821_n1), .Q(WX11110) );
  INVX0 U5821_U1 ( .INP(n10697), .ZN(U5821_n1) );
  AND2X1 U5822_U2 ( .IN1(WX11045), .IN2(U5822_n1), .Q(WX11108) );
  INVX0 U5822_U1 ( .INP(n10696), .ZN(U5822_n1) );
  AND2X1 U5823_U2 ( .IN1(WX11043), .IN2(U5823_n1), .Q(WX11106) );
  INVX0 U5823_U1 ( .INP(n10696), .ZN(U5823_n1) );
  AND2X1 U5824_U2 ( .IN1(WX11041), .IN2(U5824_n1), .Q(WX11104) );
  INVX0 U5824_U1 ( .INP(n10696), .ZN(U5824_n1) );
  AND2X1 U5825_U2 ( .IN1(WX11039), .IN2(U5825_n1), .Q(WX11102) );
  INVX0 U5825_U1 ( .INP(n10696), .ZN(U5825_n1) );
  AND2X1 U5826_U2 ( .IN1(WX11037), .IN2(U5826_n1), .Q(WX11100) );
  INVX0 U5826_U1 ( .INP(n10696), .ZN(U5826_n1) );
  AND2X1 U5827_U2 ( .IN1(test_so92), .IN2(U5827_n1), .Q(WX11098) );
  INVX0 U5827_U1 ( .INP(n10696), .ZN(U5827_n1) );
  AND2X1 U5828_U2 ( .IN1(WX11033), .IN2(U5828_n1), .Q(WX11096) );
  INVX0 U5828_U1 ( .INP(n10696), .ZN(U5828_n1) );
  AND2X1 U5829_U2 ( .IN1(WX11031), .IN2(U5829_n1), .Q(WX11094) );
  INVX0 U5829_U1 ( .INP(n10696), .ZN(U5829_n1) );
  AND2X1 U5830_U2 ( .IN1(WX11029), .IN2(U5830_n1), .Q(WX11092) );
  INVX0 U5830_U1 ( .INP(n10696), .ZN(U5830_n1) );
  AND2X1 U5831_U2 ( .IN1(WX11027), .IN2(U5831_n1), .Q(WX11090) );
  INVX0 U5831_U1 ( .INP(n10696), .ZN(U5831_n1) );
  AND2X1 U5832_U2 ( .IN1(WX11025), .IN2(U5832_n1), .Q(WX11088) );
  INVX0 U5832_U1 ( .INP(n10696), .ZN(U5832_n1) );
  AND2X1 U5833_U2 ( .IN1(WX11023), .IN2(U5833_n1), .Q(WX11086) );
  INVX0 U5833_U1 ( .INP(n10696), .ZN(U5833_n1) );
  AND2X1 U5834_U2 ( .IN1(WX11021), .IN2(U5834_n1), .Q(WX11084) );
  INVX0 U5834_U1 ( .INP(n10696), .ZN(U5834_n1) );
  AND2X1 U5835_U2 ( .IN1(WX9886), .IN2(U5835_n1), .Q(WX9949) );
  INVX0 U5835_U1 ( .INP(n10696), .ZN(U5835_n1) );
  AND2X1 U5836_U2 ( .IN1(WX9884), .IN2(U5836_n1), .Q(WX9947) );
  INVX0 U5836_U1 ( .INP(n10695), .ZN(U5836_n1) );
  AND2X1 U5837_U2 ( .IN1(WX9882), .IN2(U5837_n1), .Q(WX9945) );
  INVX0 U5837_U1 ( .INP(n10695), .ZN(U5837_n1) );
  AND2X1 U5838_U2 ( .IN1(WX9880), .IN2(U5838_n1), .Q(WX9943) );
  INVX0 U5838_U1 ( .INP(n10695), .ZN(U5838_n1) );
  AND2X1 U5839_U2 ( .IN1(WX9878), .IN2(U5839_n1), .Q(WX9941) );
  INVX0 U5839_U1 ( .INP(n10695), .ZN(U5839_n1) );
  AND2X1 U5840_U2 ( .IN1(WX9876), .IN2(U5840_n1), .Q(WX9939) );
  INVX0 U5840_U1 ( .INP(n10695), .ZN(U5840_n1) );
  AND2X1 U5841_U2 ( .IN1(WX9874), .IN2(U5841_n1), .Q(WX9937) );
  INVX0 U5841_U1 ( .INP(n10695), .ZN(U5841_n1) );
  AND2X1 U5842_U2 ( .IN1(WX9872), .IN2(U5842_n1), .Q(WX9935) );
  INVX0 U5842_U1 ( .INP(n10695), .ZN(U5842_n1) );
  AND2X1 U5843_U2 ( .IN1(WX9870), .IN2(U5843_n1), .Q(WX9933) );
  INVX0 U5843_U1 ( .INP(n10695), .ZN(U5843_n1) );
  AND2X1 U5844_U2 ( .IN1(WX9868), .IN2(U5844_n1), .Q(WX9931) );
  INVX0 U5844_U1 ( .INP(n10695), .ZN(U5844_n1) );
  AND2X1 U5845_U2 ( .IN1(WX9866), .IN2(U5845_n1), .Q(WX9929) );
  INVX0 U5845_U1 ( .INP(n10695), .ZN(U5845_n1) );
  AND2X1 U5846_U2 ( .IN1(WX9864), .IN2(U5846_n1), .Q(WX9927) );
  INVX0 U5846_U1 ( .INP(n10695), .ZN(U5846_n1) );
  AND2X1 U5847_U2 ( .IN1(WX9862), .IN2(U5847_n1), .Q(WX9925) );
  INVX0 U5847_U1 ( .INP(n10695), .ZN(U5847_n1) );
  AND2X1 U5848_U2 ( .IN1(WX9860), .IN2(U5848_n1), .Q(WX9923) );
  INVX0 U5848_U1 ( .INP(n10695), .ZN(U5848_n1) );
  AND2X1 U5849_U2 ( .IN1(WX9858), .IN2(U5849_n1), .Q(WX9921) );
  INVX0 U5849_U1 ( .INP(n10695), .ZN(U5849_n1) );
  AND2X1 U5850_U2 ( .IN1(WX9856), .IN2(U5850_n1), .Q(WX9919) );
  INVX0 U5850_U1 ( .INP(n10694), .ZN(U5850_n1) );
  AND2X1 U5851_U2 ( .IN1(test_so84), .IN2(U5851_n1), .Q(WX9917) );
  INVX0 U5851_U1 ( .INP(n10694), .ZN(U5851_n1) );
  AND2X1 U5852_U2 ( .IN1(WX9852), .IN2(U5852_n1), .Q(WX9915) );
  INVX0 U5852_U1 ( .INP(n10694), .ZN(U5852_n1) );
  AND2X1 U5853_U2 ( .IN1(WX9850), .IN2(U5853_n1), .Q(WX9913) );
  INVX0 U5853_U1 ( .INP(n10694), .ZN(U5853_n1) );
  AND2X1 U5854_U2 ( .IN1(WX9848), .IN2(U5854_n1), .Q(WX9911) );
  INVX0 U5854_U1 ( .INP(n10694), .ZN(U5854_n1) );
  AND2X1 U5855_U2 ( .IN1(WX9846), .IN2(U5855_n1), .Q(WX9909) );
  INVX0 U5855_U1 ( .INP(n10694), .ZN(U5855_n1) );
  AND2X1 U5856_U2 ( .IN1(WX9844), .IN2(U5856_n1), .Q(WX9907) );
  INVX0 U5856_U1 ( .INP(n10694), .ZN(U5856_n1) );
  AND2X1 U5857_U2 ( .IN1(WX9842), .IN2(U5857_n1), .Q(WX9905) );
  INVX0 U5857_U1 ( .INP(n10694), .ZN(U5857_n1) );
  AND2X1 U5858_U2 ( .IN1(WX9840), .IN2(U5858_n1), .Q(WX9903) );
  INVX0 U5858_U1 ( .INP(n10694), .ZN(U5858_n1) );
  AND2X1 U5859_U2 ( .IN1(WX9838), .IN2(U5859_n1), .Q(WX9901) );
  INVX0 U5859_U1 ( .INP(n10694), .ZN(U5859_n1) );
  AND2X1 U5860_U2 ( .IN1(WX9836), .IN2(U5860_n1), .Q(WX9899) );
  INVX0 U5860_U1 ( .INP(n10694), .ZN(U5860_n1) );
  AND2X1 U5861_U2 ( .IN1(WX9834), .IN2(U5861_n1), .Q(WX9897) );
  INVX0 U5861_U1 ( .INP(n10694), .ZN(U5861_n1) );
  AND2X1 U5862_U2 ( .IN1(WX9832), .IN2(U5862_n1), .Q(WX9895) );
  INVX0 U5862_U1 ( .INP(n10694), .ZN(U5862_n1) );
  AND2X1 U5863_U2 ( .IN1(WX9830), .IN2(U5863_n1), .Q(WX9893) );
  INVX0 U5863_U1 ( .INP(n10694), .ZN(U5863_n1) );
  AND2X1 U5864_U2 ( .IN1(WX9828), .IN2(U5864_n1), .Q(WX9891) );
  INVX0 U5864_U1 ( .INP(n10693), .ZN(U5864_n1) );
  AND2X1 U5865_U2 ( .IN1(WX9826), .IN2(U5865_n1), .Q(WX9889) );
  INVX0 U5865_U1 ( .INP(n10693), .ZN(U5865_n1) );
  AND2X1 U5866_U2 ( .IN1(WX9824), .IN2(U5866_n1), .Q(WX9887) );
  INVX0 U5866_U1 ( .INP(n10693), .ZN(U5866_n1) );
  AND2X1 U5867_U2 ( .IN1(WX9822), .IN2(U5867_n1), .Q(WX9885) );
  INVX0 U5867_U1 ( .INP(n10693), .ZN(U5867_n1) );
  AND2X1 U5868_U2 ( .IN1(test_so83), .IN2(U5868_n1), .Q(WX9883) );
  INVX0 U5868_U1 ( .INP(n10693), .ZN(U5868_n1) );
  AND2X1 U5869_U2 ( .IN1(WX9818), .IN2(U5869_n1), .Q(WX9881) );
  INVX0 U5869_U1 ( .INP(n10693), .ZN(U5869_n1) );
  AND2X1 U5870_U2 ( .IN1(WX9816), .IN2(U5870_n1), .Q(WX9879) );
  INVX0 U5870_U1 ( .INP(n10693), .ZN(U5870_n1) );
  AND2X1 U5871_U2 ( .IN1(WX9814), .IN2(U5871_n1), .Q(WX9877) );
  INVX0 U5871_U1 ( .INP(n10693), .ZN(U5871_n1) );
  AND2X1 U5872_U2 ( .IN1(WX9812), .IN2(U5872_n1), .Q(WX9875) );
  INVX0 U5872_U1 ( .INP(n10693), .ZN(U5872_n1) );
  AND2X1 U5873_U2 ( .IN1(WX9810), .IN2(U5873_n1), .Q(WX9873) );
  INVX0 U5873_U1 ( .INP(n10693), .ZN(U5873_n1) );
  AND2X1 U5874_U2 ( .IN1(WX9808), .IN2(U5874_n1), .Q(WX9871) );
  INVX0 U5874_U1 ( .INP(n10693), .ZN(U5874_n1) );
  AND2X1 U5875_U2 ( .IN1(WX9806), .IN2(U5875_n1), .Q(WX9869) );
  INVX0 U5875_U1 ( .INP(n10693), .ZN(U5875_n1) );
  AND2X1 U5876_U2 ( .IN1(WX9804), .IN2(U5876_n1), .Q(WX9867) );
  INVX0 U5876_U1 ( .INP(n10693), .ZN(U5876_n1) );
  AND2X1 U5877_U2 ( .IN1(WX9802), .IN2(U5877_n1), .Q(WX9865) );
  INVX0 U5877_U1 ( .INP(n10693), .ZN(U5877_n1) );
  AND2X1 U5878_U2 ( .IN1(WX9800), .IN2(U5878_n1), .Q(WX9863) );
  INVX0 U5878_U1 ( .INP(n10692), .ZN(U5878_n1) );
  AND2X1 U5879_U2 ( .IN1(WX9798), .IN2(U5879_n1), .Q(WX9861) );
  INVX0 U5879_U1 ( .INP(n10692), .ZN(U5879_n1) );
  AND2X1 U5880_U2 ( .IN1(WX9796), .IN2(U5880_n1), .Q(WX9859) );
  INVX0 U5880_U1 ( .INP(n10692), .ZN(U5880_n1) );
  AND2X1 U5881_U2 ( .IN1(WX9794), .IN2(U5881_n1), .Q(WX9857) );
  INVX0 U5881_U1 ( .INP(n10692), .ZN(U5881_n1) );
  AND2X1 U5882_U2 ( .IN1(WX9792), .IN2(U5882_n1), .Q(WX9855) );
  INVX0 U5882_U1 ( .INP(n10692), .ZN(U5882_n1) );
  AND2X1 U5883_U2 ( .IN1(WX9790), .IN2(U5883_n1), .Q(WX9853) );
  INVX0 U5883_U1 ( .INP(n10692), .ZN(U5883_n1) );
  AND2X1 U5884_U2 ( .IN1(WX9788), .IN2(U5884_n1), .Q(WX9851) );
  INVX0 U5884_U1 ( .INP(n10692), .ZN(U5884_n1) );
  AND2X1 U5885_U2 ( .IN1(test_so82), .IN2(U5885_n1), .Q(WX9849) );
  INVX0 U5885_U1 ( .INP(n10692), .ZN(U5885_n1) );
  AND2X1 U5886_U2 ( .IN1(WX9784), .IN2(U5886_n1), .Q(WX9847) );
  INVX0 U5886_U1 ( .INP(n10692), .ZN(U5886_n1) );
  AND2X1 U5887_U2 ( .IN1(WX9782), .IN2(U5887_n1), .Q(WX9845) );
  INVX0 U5887_U1 ( .INP(n10692), .ZN(U5887_n1) );
  AND2X1 U5888_U2 ( .IN1(WX9780), .IN2(U5888_n1), .Q(WX9843) );
  INVX0 U5888_U1 ( .INP(n10692), .ZN(U5888_n1) );
  AND2X1 U5889_U2 ( .IN1(WX9778), .IN2(U5889_n1), .Q(WX9841) );
  INVX0 U5889_U1 ( .INP(n10692), .ZN(U5889_n1) );
  AND2X1 U5890_U2 ( .IN1(WX9776), .IN2(U5890_n1), .Q(WX9839) );
  INVX0 U5890_U1 ( .INP(n10692), .ZN(U5890_n1) );
  AND2X1 U5891_U2 ( .IN1(WX9774), .IN2(U5891_n1), .Q(WX9837) );
  INVX0 U5891_U1 ( .INP(n10692), .ZN(U5891_n1) );
  AND2X1 U5892_U2 ( .IN1(WX9772), .IN2(U5892_n1), .Q(WX9835) );
  INVX0 U5892_U1 ( .INP(n10691), .ZN(U5892_n1) );
  AND2X1 U5893_U2 ( .IN1(WX9770), .IN2(U5893_n1), .Q(WX9833) );
  INVX0 U5893_U1 ( .INP(n10691), .ZN(U5893_n1) );
  AND2X1 U5894_U2 ( .IN1(WX9768), .IN2(U5894_n1), .Q(WX9831) );
  INVX0 U5894_U1 ( .INP(n10691), .ZN(U5894_n1) );
  AND2X1 U5895_U2 ( .IN1(WX9766), .IN2(U5895_n1), .Q(WX9829) );
  INVX0 U5895_U1 ( .INP(n10691), .ZN(U5895_n1) );
  AND2X1 U5896_U2 ( .IN1(WX9764), .IN2(U5896_n1), .Q(WX9827) );
  INVX0 U5896_U1 ( .INP(n10691), .ZN(U5896_n1) );
  AND2X1 U5897_U2 ( .IN1(WX9762), .IN2(U5897_n1), .Q(WX9825) );
  INVX0 U5897_U1 ( .INP(n10691), .ZN(U5897_n1) );
  AND2X1 U5898_U2 ( .IN1(WX9760), .IN2(U5898_n1), .Q(WX9823) );
  INVX0 U5898_U1 ( .INP(n10691), .ZN(U5898_n1) );
  AND2X1 U5899_U2 ( .IN1(WX9758), .IN2(U5899_n1), .Q(WX9821) );
  INVX0 U5899_U1 ( .INP(n10691), .ZN(U5899_n1) );
  AND2X1 U5900_U2 ( .IN1(WX9756), .IN2(U5900_n1), .Q(WX9819) );
  INVX0 U5900_U1 ( .INP(n10691), .ZN(U5900_n1) );
  AND2X1 U5901_U2 ( .IN1(WX9754), .IN2(U5901_n1), .Q(WX9817) );
  INVX0 U5901_U1 ( .INP(n10691), .ZN(U5901_n1) );
  AND2X1 U5902_U2 ( .IN1(test_so81), .IN2(U5902_n1), .Q(WX9815) );
  INVX0 U5902_U1 ( .INP(n10691), .ZN(U5902_n1) );
  AND2X1 U5903_U2 ( .IN1(WX9750), .IN2(U5903_n1), .Q(WX9813) );
  INVX0 U5903_U1 ( .INP(n10691), .ZN(U5903_n1) );
  AND2X1 U5904_U2 ( .IN1(WX9748), .IN2(U5904_n1), .Q(WX9811) );
  INVX0 U5904_U1 ( .INP(n10691), .ZN(U5904_n1) );
  AND2X1 U5905_U2 ( .IN1(WX9746), .IN2(U5905_n1), .Q(WX9809) );
  INVX0 U5905_U1 ( .INP(n10691), .ZN(U5905_n1) );
  AND2X1 U5906_U2 ( .IN1(WX9744), .IN2(U5906_n1), .Q(WX9807) );
  INVX0 U5906_U1 ( .INP(n10690), .ZN(U5906_n1) );
  AND2X1 U5907_U2 ( .IN1(WX9742), .IN2(U5907_n1), .Q(WX9805) );
  INVX0 U5907_U1 ( .INP(n10690), .ZN(U5907_n1) );
  AND2X1 U5908_U2 ( .IN1(WX9740), .IN2(U5908_n1), .Q(WX9803) );
  INVX0 U5908_U1 ( .INP(n10690), .ZN(U5908_n1) );
  AND2X1 U5909_U2 ( .IN1(WX9738), .IN2(U5909_n1), .Q(WX9801) );
  INVX0 U5909_U1 ( .INP(n10690), .ZN(U5909_n1) );
  AND2X1 U5910_U2 ( .IN1(WX9736), .IN2(U5910_n1), .Q(WX9799) );
  INVX0 U5910_U1 ( .INP(n10690), .ZN(U5910_n1) );
  AND2X1 U5911_U2 ( .IN1(WX9734), .IN2(U5911_n1), .Q(WX9797) );
  INVX0 U5911_U1 ( .INP(n10690), .ZN(U5911_n1) );
  AND2X1 U5912_U2 ( .IN1(WX9732), .IN2(U5912_n1), .Q(WX9795) );
  INVX0 U5912_U1 ( .INP(n10690), .ZN(U5912_n1) );
  AND2X1 U5913_U2 ( .IN1(WX9730), .IN2(U5913_n1), .Q(WX9793) );
  INVX0 U5913_U1 ( .INP(n10690), .ZN(U5913_n1) );
  AND2X1 U5914_U2 ( .IN1(WX9728), .IN2(U5914_n1), .Q(WX9791) );
  INVX0 U5914_U1 ( .INP(n10690), .ZN(U5914_n1) );
  AND2X1 U5915_U2 ( .IN1(WX8593), .IN2(U5915_n1), .Q(WX8656) );
  INVX0 U5915_U1 ( .INP(n10690), .ZN(U5915_n1) );
  AND2X1 U5916_U2 ( .IN1(WX8591), .IN2(U5916_n1), .Q(WX8654) );
  INVX0 U5916_U1 ( .INP(n10690), .ZN(U5916_n1) );
  AND2X1 U5917_U2 ( .IN1(WX8589), .IN2(U5917_n1), .Q(WX8652) );
  INVX0 U5917_U1 ( .INP(n10690), .ZN(U5917_n1) );
  AND2X1 U5918_U2 ( .IN1(WX8587), .IN2(U5918_n1), .Q(WX8650) );
  INVX0 U5918_U1 ( .INP(n10690), .ZN(U5918_n1) );
  AND2X1 U5919_U2 ( .IN1(WX8585), .IN2(U5919_n1), .Q(WX8648) );
  INVX0 U5919_U1 ( .INP(n10690), .ZN(U5919_n1) );
  AND2X1 U5920_U2 ( .IN1(WX8583), .IN2(U5920_n1), .Q(WX8646) );
  INVX0 U5920_U1 ( .INP(n10689), .ZN(U5920_n1) );
  AND2X1 U5921_U2 ( .IN1(WX8581), .IN2(U5921_n1), .Q(WX8644) );
  INVX0 U5921_U1 ( .INP(n10689), .ZN(U5921_n1) );
  AND2X1 U5922_U2 ( .IN1(WX8579), .IN2(U5922_n1), .Q(WX8642) );
  INVX0 U5922_U1 ( .INP(n10689), .ZN(U5922_n1) );
  AND2X1 U5923_U2 ( .IN1(WX8577), .IN2(U5923_n1), .Q(WX8640) );
  INVX0 U5923_U1 ( .INP(n10689), .ZN(U5923_n1) );
  AND2X1 U5924_U2 ( .IN1(WX8575), .IN2(U5924_n1), .Q(WX8638) );
  INVX0 U5924_U1 ( .INP(n10689), .ZN(U5924_n1) );
  AND2X1 U5925_U2 ( .IN1(WX8573), .IN2(U5925_n1), .Q(WX8636) );
  INVX0 U5925_U1 ( .INP(n10689), .ZN(U5925_n1) );
  AND2X1 U5926_U2 ( .IN1(test_so73), .IN2(U5926_n1), .Q(WX8634) );
  INVX0 U5926_U1 ( .INP(n10689), .ZN(U5926_n1) );
  AND2X1 U5927_U2 ( .IN1(WX8569), .IN2(U5927_n1), .Q(WX8632) );
  INVX0 U5927_U1 ( .INP(n10689), .ZN(U5927_n1) );
  AND2X1 U5928_U2 ( .IN1(WX8567), .IN2(U5928_n1), .Q(WX8630) );
  INVX0 U5928_U1 ( .INP(n10689), .ZN(U5928_n1) );
  AND2X1 U5929_U2 ( .IN1(WX8565), .IN2(U5929_n1), .Q(WX8628) );
  INVX0 U5929_U1 ( .INP(n10689), .ZN(U5929_n1) );
  AND2X1 U5930_U2 ( .IN1(WX8563), .IN2(U5930_n1), .Q(WX8626) );
  INVX0 U5930_U1 ( .INP(n10689), .ZN(U5930_n1) );
  AND2X1 U5931_U2 ( .IN1(WX8561), .IN2(U5931_n1), .Q(WX8624) );
  INVX0 U5931_U1 ( .INP(n10689), .ZN(U5931_n1) );
  AND2X1 U5932_U2 ( .IN1(WX8559), .IN2(U5932_n1), .Q(WX8622) );
  INVX0 U5932_U1 ( .INP(n10689), .ZN(U5932_n1) );
  AND2X1 U5933_U2 ( .IN1(WX8557), .IN2(U5933_n1), .Q(WX8620) );
  INVX0 U5933_U1 ( .INP(n10689), .ZN(U5933_n1) );
  AND2X1 U5934_U2 ( .IN1(WX8555), .IN2(U5934_n1), .Q(WX8618) );
  INVX0 U5934_U1 ( .INP(n10688), .ZN(U5934_n1) );
  AND2X1 U5935_U2 ( .IN1(WX8553), .IN2(U5935_n1), .Q(WX8616) );
  INVX0 U5935_U1 ( .INP(n10688), .ZN(U5935_n1) );
  AND2X1 U5936_U2 ( .IN1(WX8551), .IN2(U5936_n1), .Q(WX8614) );
  INVX0 U5936_U1 ( .INP(n10688), .ZN(U5936_n1) );
  AND2X1 U5937_U2 ( .IN1(WX8549), .IN2(U5937_n1), .Q(WX8612) );
  INVX0 U5937_U1 ( .INP(n10688), .ZN(U5937_n1) );
  AND2X1 U5938_U2 ( .IN1(WX8547), .IN2(U5938_n1), .Q(WX8610) );
  INVX0 U5938_U1 ( .INP(n10688), .ZN(U5938_n1) );
  AND2X1 U5939_U2 ( .IN1(WX8545), .IN2(U5939_n1), .Q(WX8608) );
  INVX0 U5939_U1 ( .INP(n10688), .ZN(U5939_n1) );
  AND2X1 U5940_U2 ( .IN1(WX8543), .IN2(U5940_n1), .Q(WX8606) );
  INVX0 U5940_U1 ( .INP(n10688), .ZN(U5940_n1) );
  AND2X1 U5941_U2 ( .IN1(WX8541), .IN2(U5941_n1), .Q(WX8604) );
  INVX0 U5941_U1 ( .INP(n10688), .ZN(U5941_n1) );
  AND2X1 U5942_U2 ( .IN1(WX8539), .IN2(U5942_n1), .Q(WX8602) );
  INVX0 U5942_U1 ( .INP(n10688), .ZN(U5942_n1) );
  AND2X1 U5943_U2 ( .IN1(test_so72), .IN2(U5943_n1), .Q(WX8600) );
  INVX0 U5943_U1 ( .INP(n10688), .ZN(U5943_n1) );
  AND2X1 U5944_U2 ( .IN1(WX8535), .IN2(U5944_n1), .Q(WX8598) );
  INVX0 U5944_U1 ( .INP(n10688), .ZN(U5944_n1) );
  AND2X1 U5945_U2 ( .IN1(WX8533), .IN2(U5945_n1), .Q(WX8596) );
  INVX0 U5945_U1 ( .INP(n10688), .ZN(U5945_n1) );
  AND2X1 U5946_U2 ( .IN1(WX8531), .IN2(U5946_n1), .Q(WX8594) );
  INVX0 U5946_U1 ( .INP(n10688), .ZN(U5946_n1) );
  AND2X1 U5947_U2 ( .IN1(WX8529), .IN2(U5947_n1), .Q(WX8592) );
  INVX0 U5947_U1 ( .INP(n10688), .ZN(U5947_n1) );
  AND2X1 U5948_U2 ( .IN1(WX8527), .IN2(U5948_n1), .Q(WX8590) );
  INVX0 U5948_U1 ( .INP(n10687), .ZN(U5948_n1) );
  AND2X1 U5949_U2 ( .IN1(WX8525), .IN2(U5949_n1), .Q(WX8588) );
  INVX0 U5949_U1 ( .INP(n10687), .ZN(U5949_n1) );
  AND2X1 U5950_U2 ( .IN1(WX8523), .IN2(U5950_n1), .Q(WX8586) );
  INVX0 U5950_U1 ( .INP(n10687), .ZN(U5950_n1) );
  AND2X1 U5951_U2 ( .IN1(WX8521), .IN2(U5951_n1), .Q(WX8584) );
  INVX0 U5951_U1 ( .INP(n10687), .ZN(U5951_n1) );
  AND2X1 U5952_U2 ( .IN1(WX8519), .IN2(U5952_n1), .Q(WX8582) );
  INVX0 U5952_U1 ( .INP(n10687), .ZN(U5952_n1) );
  AND2X1 U5953_U2 ( .IN1(WX8517), .IN2(U5953_n1), .Q(WX8580) );
  INVX0 U5953_U1 ( .INP(n10687), .ZN(U5953_n1) );
  AND2X1 U5954_U2 ( .IN1(WX8515), .IN2(U5954_n1), .Q(WX8578) );
  INVX0 U5954_U1 ( .INP(n10687), .ZN(U5954_n1) );
  AND2X1 U5955_U2 ( .IN1(WX8513), .IN2(U5955_n1), .Q(WX8576) );
  INVX0 U5955_U1 ( .INP(n10687), .ZN(U5955_n1) );
  AND2X1 U5956_U2 ( .IN1(WX8511), .IN2(U5956_n1), .Q(WX8574) );
  INVX0 U5956_U1 ( .INP(n10687), .ZN(U5956_n1) );
  AND2X1 U5957_U2 ( .IN1(WX8509), .IN2(U5957_n1), .Q(WX8572) );
  INVX0 U5957_U1 ( .INP(n10687), .ZN(U5957_n1) );
  AND2X1 U5958_U2 ( .IN1(WX8507), .IN2(U5958_n1), .Q(WX8570) );
  INVX0 U5958_U1 ( .INP(n10687), .ZN(U5958_n1) );
  AND2X1 U5959_U2 ( .IN1(WX8505), .IN2(U5959_n1), .Q(WX8568) );
  INVX0 U5959_U1 ( .INP(n10687), .ZN(U5959_n1) );
  AND2X1 U5960_U2 ( .IN1(test_so71), .IN2(U5960_n1), .Q(WX8566) );
  INVX0 U5960_U1 ( .INP(n10687), .ZN(U5960_n1) );
  AND2X1 U5961_U2 ( .IN1(WX8501), .IN2(U5961_n1), .Q(WX8564) );
  INVX0 U5961_U1 ( .INP(n10687), .ZN(U5961_n1) );
  AND2X1 U5962_U2 ( .IN1(WX8499), .IN2(U5962_n1), .Q(WX8562) );
  INVX0 U5962_U1 ( .INP(n10686), .ZN(U5962_n1) );
  AND2X1 U5963_U2 ( .IN1(WX8497), .IN2(U5963_n1), .Q(WX8560) );
  INVX0 U5963_U1 ( .INP(n10686), .ZN(U5963_n1) );
  AND2X1 U5964_U2 ( .IN1(WX8495), .IN2(U5964_n1), .Q(WX8558) );
  INVX0 U5964_U1 ( .INP(n10686), .ZN(U5964_n1) );
  AND2X1 U5965_U2 ( .IN1(WX8493), .IN2(U5965_n1), .Q(WX8556) );
  INVX0 U5965_U1 ( .INP(n10686), .ZN(U5965_n1) );
  AND2X1 U5966_U2 ( .IN1(WX8491), .IN2(U5966_n1), .Q(WX8554) );
  INVX0 U5966_U1 ( .INP(n10686), .ZN(U5966_n1) );
  AND2X1 U5967_U2 ( .IN1(WX8489), .IN2(U5967_n1), .Q(WX8552) );
  INVX0 U5967_U1 ( .INP(n10686), .ZN(U5967_n1) );
  AND2X1 U5968_U2 ( .IN1(WX8487), .IN2(U5968_n1), .Q(WX8550) );
  INVX0 U5968_U1 ( .INP(n10686), .ZN(U5968_n1) );
  AND2X1 U5969_U2 ( .IN1(WX8485), .IN2(U5969_n1), .Q(WX8548) );
  INVX0 U5969_U1 ( .INP(n10686), .ZN(U5969_n1) );
  AND2X1 U5970_U2 ( .IN1(WX8483), .IN2(U5970_n1), .Q(WX8546) );
  INVX0 U5970_U1 ( .INP(n10686), .ZN(U5970_n1) );
  AND2X1 U5971_U2 ( .IN1(WX8481), .IN2(U5971_n1), .Q(WX8544) );
  INVX0 U5971_U1 ( .INP(n10686), .ZN(U5971_n1) );
  AND2X1 U5972_U2 ( .IN1(WX8479), .IN2(U5972_n1), .Q(WX8542) );
  INVX0 U5972_U1 ( .INP(n10686), .ZN(U5972_n1) );
  AND2X1 U5973_U2 ( .IN1(WX8477), .IN2(U5973_n1), .Q(WX8540) );
  INVX0 U5973_U1 ( .INP(n10686), .ZN(U5973_n1) );
  AND2X1 U5974_U2 ( .IN1(WX8475), .IN2(U5974_n1), .Q(WX8538) );
  INVX0 U5974_U1 ( .INP(n10686), .ZN(U5974_n1) );
  AND2X1 U5975_U2 ( .IN1(WX8473), .IN2(U5975_n1), .Q(WX8536) );
  INVX0 U5975_U1 ( .INP(n10686), .ZN(U5975_n1) );
  AND2X1 U5976_U2 ( .IN1(WX8471), .IN2(U5976_n1), .Q(WX8534) );
  INVX0 U5976_U1 ( .INP(n10685), .ZN(U5976_n1) );
  AND2X1 U5977_U2 ( .IN1(test_so70), .IN2(U5977_n1), .Q(WX8532) );
  INVX0 U5977_U1 ( .INP(n10685), .ZN(U5977_n1) );
  AND2X1 U5978_U2 ( .IN1(WX8467), .IN2(U5978_n1), .Q(WX8530) );
  INVX0 U5978_U1 ( .INP(n10685), .ZN(U5978_n1) );
  AND2X1 U5979_U2 ( .IN1(WX8465), .IN2(U5979_n1), .Q(WX8528) );
  INVX0 U5979_U1 ( .INP(n10685), .ZN(U5979_n1) );
  AND2X1 U5980_U2 ( .IN1(WX8463), .IN2(U5980_n1), .Q(WX8526) );
  INVX0 U5980_U1 ( .INP(n10685), .ZN(U5980_n1) );
  AND2X1 U5981_U2 ( .IN1(WX8461), .IN2(U5981_n1), .Q(WX8524) );
  INVX0 U5981_U1 ( .INP(n10685), .ZN(U5981_n1) );
  AND2X1 U5982_U2 ( .IN1(WX8459), .IN2(U5982_n1), .Q(WX8522) );
  INVX0 U5982_U1 ( .INP(n10685), .ZN(U5982_n1) );
  AND2X1 U5983_U2 ( .IN1(WX8457), .IN2(U5983_n1), .Q(WX8520) );
  INVX0 U5983_U1 ( .INP(n10685), .ZN(U5983_n1) );
  AND2X1 U5984_U2 ( .IN1(WX8455), .IN2(U5984_n1), .Q(WX8518) );
  INVX0 U5984_U1 ( .INP(n10685), .ZN(U5984_n1) );
  AND2X1 U5985_U2 ( .IN1(WX8453), .IN2(U5985_n1), .Q(WX8516) );
  INVX0 U5985_U1 ( .INP(n10685), .ZN(U5985_n1) );
  AND2X1 U5986_U2 ( .IN1(WX8451), .IN2(U5986_n1), .Q(WX8514) );
  INVX0 U5986_U1 ( .INP(n10685), .ZN(U5986_n1) );
  AND2X1 U5987_U2 ( .IN1(WX8449), .IN2(U5987_n1), .Q(WX8512) );
  INVX0 U5987_U1 ( .INP(n10685), .ZN(U5987_n1) );
  AND2X1 U5988_U2 ( .IN1(WX8447), .IN2(U5988_n1), .Q(WX8510) );
  INVX0 U5988_U1 ( .INP(n10685), .ZN(U5988_n1) );
  AND2X1 U5989_U2 ( .IN1(WX8445), .IN2(U5989_n1), .Q(WX8508) );
  INVX0 U5989_U1 ( .INP(n10685), .ZN(U5989_n1) );
  AND2X1 U5990_U2 ( .IN1(WX8443), .IN2(U5990_n1), .Q(WX8506) );
  INVX0 U5990_U1 ( .INP(n10684), .ZN(U5990_n1) );
  AND2X1 U5991_U2 ( .IN1(WX8441), .IN2(U5991_n1), .Q(WX8504) );
  INVX0 U5991_U1 ( .INP(n10684), .ZN(U5991_n1) );
  AND2X1 U5992_U2 ( .IN1(WX8439), .IN2(U5992_n1), .Q(WX8502) );
  INVX0 U5992_U1 ( .INP(n10684), .ZN(U5992_n1) );
  AND2X1 U5993_U2 ( .IN1(WX8437), .IN2(U5993_n1), .Q(WX8500) );
  INVX0 U5993_U1 ( .INP(n10684), .ZN(U5993_n1) );
  AND2X1 U5994_U2 ( .IN1(test_so69), .IN2(U5994_n1), .Q(WX8498) );
  INVX0 U5994_U1 ( .INP(n10684), .ZN(U5994_n1) );
  AND2X1 U5995_U2 ( .IN1(WX7300), .IN2(U5995_n1), .Q(WX7363) );
  INVX0 U5995_U1 ( .INP(n10684), .ZN(U5995_n1) );
  AND2X1 U5996_U2 ( .IN1(WX7298), .IN2(U5996_n1), .Q(WX7361) );
  INVX0 U5996_U1 ( .INP(n10684), .ZN(U5996_n1) );
  AND2X1 U5997_U2 ( .IN1(WX7296), .IN2(U5997_n1), .Q(WX7359) );
  INVX0 U5997_U1 ( .INP(n10684), .ZN(U5997_n1) );
  AND2X1 U5998_U2 ( .IN1(WX7294), .IN2(U5998_n1), .Q(WX7357) );
  INVX0 U5998_U1 ( .INP(n10684), .ZN(U5998_n1) );
  AND2X1 U5999_U2 ( .IN1(WX7292), .IN2(U5999_n1), .Q(WX7355) );
  INVX0 U5999_U1 ( .INP(n10684), .ZN(U5999_n1) );
  AND2X1 U6000_U2 ( .IN1(WX7290), .IN2(U6000_n1), .Q(WX7353) );
  INVX0 U6000_U1 ( .INP(n10684), .ZN(U6000_n1) );
  AND2X1 U6001_U2 ( .IN1(test_so62), .IN2(U6001_n1), .Q(WX7351) );
  INVX0 U6001_U1 ( .INP(n10684), .ZN(U6001_n1) );
  AND2X1 U6002_U2 ( .IN1(WX7286), .IN2(U6002_n1), .Q(WX7349) );
  INVX0 U6002_U1 ( .INP(n10684), .ZN(U6002_n1) );
  AND2X1 U6003_U2 ( .IN1(WX7284), .IN2(U6003_n1), .Q(WX7347) );
  INVX0 U6003_U1 ( .INP(n10684), .ZN(U6003_n1) );
  AND2X1 U6004_U2 ( .IN1(WX7282), .IN2(U6004_n1), .Q(WX7345) );
  INVX0 U6004_U1 ( .INP(n10683), .ZN(U6004_n1) );
  AND2X1 U6005_U2 ( .IN1(WX7280), .IN2(U6005_n1), .Q(WX7343) );
  INVX0 U6005_U1 ( .INP(n10683), .ZN(U6005_n1) );
  AND2X1 U6006_U2 ( .IN1(WX7278), .IN2(U6006_n1), .Q(WX7341) );
  INVX0 U6006_U1 ( .INP(n10683), .ZN(U6006_n1) );
  AND2X1 U6007_U2 ( .IN1(WX7276), .IN2(U6007_n1), .Q(WX7339) );
  INVX0 U6007_U1 ( .INP(n10683), .ZN(U6007_n1) );
  AND2X1 U6008_U2 ( .IN1(WX7274), .IN2(U6008_n1), .Q(WX7337) );
  INVX0 U6008_U1 ( .INP(n10683), .ZN(U6008_n1) );
  AND2X1 U6009_U2 ( .IN1(WX7272), .IN2(U6009_n1), .Q(WX7335) );
  INVX0 U6009_U1 ( .INP(n10683), .ZN(U6009_n1) );
  AND2X1 U6010_U2 ( .IN1(WX7270), .IN2(U6010_n1), .Q(WX7333) );
  INVX0 U6010_U1 ( .INP(n10683), .ZN(U6010_n1) );
  AND2X1 U6011_U2 ( .IN1(WX7268), .IN2(U6011_n1), .Q(WX7331) );
  INVX0 U6011_U1 ( .INP(n10683), .ZN(U6011_n1) );
  AND2X1 U6012_U2 ( .IN1(WX7266), .IN2(U6012_n1), .Q(WX7329) );
  INVX0 U6012_U1 ( .INP(n10683), .ZN(U6012_n1) );
  AND2X1 U6013_U2 ( .IN1(WX7264), .IN2(U6013_n1), .Q(WX7327) );
  INVX0 U6013_U1 ( .INP(n10683), .ZN(U6013_n1) );
  AND2X1 U6014_U2 ( .IN1(WX7262), .IN2(U6014_n1), .Q(WX7325) );
  INVX0 U6014_U1 ( .INP(n10683), .ZN(U6014_n1) );
  AND2X1 U6015_U2 ( .IN1(WX7260), .IN2(U6015_n1), .Q(WX7323) );
  INVX0 U6015_U1 ( .INP(n10683), .ZN(U6015_n1) );
  AND2X1 U6016_U2 ( .IN1(WX7258), .IN2(U6016_n1), .Q(WX7321) );
  INVX0 U6016_U1 ( .INP(n10683), .ZN(U6016_n1) );
  AND2X1 U6017_U2 ( .IN1(WX7256), .IN2(U6017_n1), .Q(WX7319) );
  INVX0 U6017_U1 ( .INP(n10683), .ZN(U6017_n1) );
  AND2X1 U6018_U2 ( .IN1(test_so61), .IN2(U6018_n1), .Q(WX7317) );
  INVX0 U6018_U1 ( .INP(n10682), .ZN(U6018_n1) );
  AND2X1 U6019_U2 ( .IN1(WX7252), .IN2(U6019_n1), .Q(WX7315) );
  INVX0 U6019_U1 ( .INP(n10682), .ZN(U6019_n1) );
  AND2X1 U6020_U2 ( .IN1(WX7250), .IN2(U6020_n1), .Q(WX7313) );
  INVX0 U6020_U1 ( .INP(n10682), .ZN(U6020_n1) );
  AND2X1 U6021_U2 ( .IN1(WX7248), .IN2(U6021_n1), .Q(WX7311) );
  INVX0 U6021_U1 ( .INP(n10682), .ZN(U6021_n1) );
  AND2X1 U6022_U2 ( .IN1(WX7246), .IN2(U6022_n1), .Q(WX7309) );
  INVX0 U6022_U1 ( .INP(n10682), .ZN(U6022_n1) );
  AND2X1 U6023_U2 ( .IN1(WX7244), .IN2(U6023_n1), .Q(WX7307) );
  INVX0 U6023_U1 ( .INP(n10682), .ZN(U6023_n1) );
  AND2X1 U6024_U2 ( .IN1(WX7242), .IN2(U6024_n1), .Q(WX7305) );
  INVX0 U6024_U1 ( .INP(n10682), .ZN(U6024_n1) );
  AND2X1 U6025_U2 ( .IN1(WX7240), .IN2(U6025_n1), .Q(WX7303) );
  INVX0 U6025_U1 ( .INP(n10682), .ZN(U6025_n1) );
  AND2X1 U6026_U2 ( .IN1(WX7238), .IN2(U6026_n1), .Q(WX7301) );
  INVX0 U6026_U1 ( .INP(n10682), .ZN(U6026_n1) );
  AND2X1 U6027_U2 ( .IN1(WX7236), .IN2(U6027_n1), .Q(WX7299) );
  INVX0 U6027_U1 ( .INP(n10682), .ZN(U6027_n1) );
  AND2X1 U6028_U2 ( .IN1(WX7234), .IN2(U6028_n1), .Q(WX7297) );
  INVX0 U6028_U1 ( .INP(n10682), .ZN(U6028_n1) );
  AND2X1 U6029_U2 ( .IN1(WX7232), .IN2(U6029_n1), .Q(WX7295) );
  INVX0 U6029_U1 ( .INP(n10682), .ZN(U6029_n1) );
  AND2X1 U6030_U2 ( .IN1(WX7230), .IN2(U6030_n1), .Q(WX7293) );
  INVX0 U6030_U1 ( .INP(n10682), .ZN(U6030_n1) );
  AND2X1 U6031_U2 ( .IN1(WX7228), .IN2(U6031_n1), .Q(WX7291) );
  INVX0 U6031_U1 ( .INP(n10682), .ZN(U6031_n1) );
  AND2X1 U6032_U2 ( .IN1(WX7226), .IN2(U6032_n1), .Q(WX7289) );
  INVX0 U6032_U1 ( .INP(n10681), .ZN(U6032_n1) );
  AND2X1 U6033_U2 ( .IN1(WX7224), .IN2(U6033_n1), .Q(WX7287) );
  INVX0 U6033_U1 ( .INP(n10681), .ZN(U6033_n1) );
  AND2X1 U6034_U2 ( .IN1(WX7222), .IN2(U6034_n1), .Q(WX7285) );
  INVX0 U6034_U1 ( .INP(n10681), .ZN(U6034_n1) );
  AND2X1 U6035_U2 ( .IN1(test_so60), .IN2(U6035_n1), .Q(WX7283) );
  INVX0 U6035_U1 ( .INP(n10681), .ZN(U6035_n1) );
  AND2X1 U6036_U2 ( .IN1(WX7218), .IN2(U6036_n1), .Q(WX7281) );
  INVX0 U6036_U1 ( .INP(n10681), .ZN(U6036_n1) );
  AND2X1 U6037_U2 ( .IN1(WX7216), .IN2(U6037_n1), .Q(WX7279) );
  INVX0 U6037_U1 ( .INP(n10681), .ZN(U6037_n1) );
  AND2X1 U6038_U2 ( .IN1(WX7214), .IN2(U6038_n1), .Q(WX7277) );
  INVX0 U6038_U1 ( .INP(n10681), .ZN(U6038_n1) );
  AND2X1 U6039_U2 ( .IN1(WX7212), .IN2(U6039_n1), .Q(WX7275) );
  INVX0 U6039_U1 ( .INP(n10681), .ZN(U6039_n1) );
  AND2X1 U6040_U2 ( .IN1(WX7210), .IN2(U6040_n1), .Q(WX7273) );
  INVX0 U6040_U1 ( .INP(n10681), .ZN(U6040_n1) );
  AND2X1 U6041_U2 ( .IN1(WX7208), .IN2(U6041_n1), .Q(WX7271) );
  INVX0 U6041_U1 ( .INP(n10681), .ZN(U6041_n1) );
  AND2X1 U6042_U2 ( .IN1(WX7206), .IN2(U6042_n1), .Q(WX7269) );
  INVX0 U6042_U1 ( .INP(n10681), .ZN(U6042_n1) );
  AND2X1 U6043_U2 ( .IN1(WX7204), .IN2(U6043_n1), .Q(WX7267) );
  INVX0 U6043_U1 ( .INP(n10681), .ZN(U6043_n1) );
  AND2X1 U6044_U2 ( .IN1(WX7202), .IN2(U6044_n1), .Q(WX7265) );
  INVX0 U6044_U1 ( .INP(n10681), .ZN(U6044_n1) );
  AND2X1 U6045_U2 ( .IN1(WX7200), .IN2(U6045_n1), .Q(WX7263) );
  INVX0 U6045_U1 ( .INP(n10681), .ZN(U6045_n1) );
  AND2X1 U6046_U2 ( .IN1(WX7198), .IN2(U6046_n1), .Q(WX7261) );
  INVX0 U6046_U1 ( .INP(n10680), .ZN(U6046_n1) );
  AND2X1 U6047_U2 ( .IN1(WX7196), .IN2(U6047_n1), .Q(WX7259) );
  INVX0 U6047_U1 ( .INP(n10680), .ZN(U6047_n1) );
  AND2X1 U6048_U2 ( .IN1(WX7194), .IN2(U6048_n1), .Q(WX7257) );
  INVX0 U6048_U1 ( .INP(n10680), .ZN(U6048_n1) );
  AND2X1 U6049_U2 ( .IN1(WX7192), .IN2(U6049_n1), .Q(WX7255) );
  INVX0 U6049_U1 ( .INP(n10680), .ZN(U6049_n1) );
  AND2X1 U6050_U2 ( .IN1(WX7190), .IN2(U6050_n1), .Q(WX7253) );
  INVX0 U6050_U1 ( .INP(n10680), .ZN(U6050_n1) );
  AND2X1 U6051_U2 ( .IN1(WX7188), .IN2(U6051_n1), .Q(WX7251) );
  INVX0 U6051_U1 ( .INP(n10680), .ZN(U6051_n1) );
  AND2X1 U6052_U2 ( .IN1(test_so59), .IN2(U6052_n1), .Q(WX7249) );
  INVX0 U6052_U1 ( .INP(n10680), .ZN(U6052_n1) );
  AND2X1 U6053_U2 ( .IN1(WX7184), .IN2(U6053_n1), .Q(WX7247) );
  INVX0 U6053_U1 ( .INP(n10680), .ZN(U6053_n1) );
  AND2X1 U6054_U2 ( .IN1(WX7182), .IN2(U6054_n1), .Q(WX7245) );
  INVX0 U6054_U1 ( .INP(n10680), .ZN(U6054_n1) );
  AND2X1 U6055_U2 ( .IN1(WX7180), .IN2(U6055_n1), .Q(WX7243) );
  INVX0 U6055_U1 ( .INP(n10680), .ZN(U6055_n1) );
  AND2X1 U6056_U2 ( .IN1(WX7178), .IN2(U6056_n1), .Q(WX7241) );
  INVX0 U6056_U1 ( .INP(n10680), .ZN(U6056_n1) );
  AND2X1 U6057_U2 ( .IN1(WX7176), .IN2(U6057_n1), .Q(WX7239) );
  INVX0 U6057_U1 ( .INP(n10680), .ZN(U6057_n1) );
  AND2X1 U6058_U2 ( .IN1(WX7174), .IN2(U6058_n1), .Q(WX7237) );
  INVX0 U6058_U1 ( .INP(n10680), .ZN(U6058_n1) );
  AND2X1 U6059_U2 ( .IN1(WX7172), .IN2(U6059_n1), .Q(WX7235) );
  INVX0 U6059_U1 ( .INP(n10680), .ZN(U6059_n1) );
  AND2X1 U6060_U2 ( .IN1(WX7170), .IN2(U6060_n1), .Q(WX7233) );
  INVX0 U6060_U1 ( .INP(n10679), .ZN(U6060_n1) );
  AND2X1 U6061_U2 ( .IN1(WX7168), .IN2(U6061_n1), .Q(WX7231) );
  INVX0 U6061_U1 ( .INP(n10679), .ZN(U6061_n1) );
  AND2X1 U6062_U2 ( .IN1(WX7166), .IN2(U6062_n1), .Q(WX7229) );
  INVX0 U6062_U1 ( .INP(n10679), .ZN(U6062_n1) );
  AND2X1 U6063_U2 ( .IN1(WX7164), .IN2(U6063_n1), .Q(WX7227) );
  INVX0 U6063_U1 ( .INP(n10679), .ZN(U6063_n1) );
  AND2X1 U6064_U2 ( .IN1(WX7162), .IN2(U6064_n1), .Q(WX7225) );
  INVX0 U6064_U1 ( .INP(n10679), .ZN(U6064_n1) );
  AND2X1 U6065_U2 ( .IN1(WX7160), .IN2(U6065_n1), .Q(WX7223) );
  INVX0 U6065_U1 ( .INP(n10679), .ZN(U6065_n1) );
  AND2X1 U6066_U2 ( .IN1(WX7158), .IN2(U6066_n1), .Q(WX7221) );
  INVX0 U6066_U1 ( .INP(n10679), .ZN(U6066_n1) );
  AND2X1 U6067_U2 ( .IN1(WX7156), .IN2(U6067_n1), .Q(WX7219) );
  INVX0 U6067_U1 ( .INP(n10679), .ZN(U6067_n1) );
  AND2X1 U6068_U2 ( .IN1(WX7154), .IN2(U6068_n1), .Q(WX7217) );
  INVX0 U6068_U1 ( .INP(n10679), .ZN(U6068_n1) );
  AND2X1 U6069_U2 ( .IN1(test_so58), .IN2(U6069_n1), .Q(WX7215) );
  INVX0 U6069_U1 ( .INP(n10679), .ZN(U6069_n1) );
  AND2X1 U6070_U2 ( .IN1(WX7150), .IN2(U6070_n1), .Q(WX7213) );
  INVX0 U6070_U1 ( .INP(n10679), .ZN(U6070_n1) );
  AND2X1 U6071_U2 ( .IN1(WX7148), .IN2(U6071_n1), .Q(WX7211) );
  INVX0 U6071_U1 ( .INP(n10679), .ZN(U6071_n1) );
  AND2X1 U6072_U2 ( .IN1(WX7146), .IN2(U6072_n1), .Q(WX7209) );
  INVX0 U6072_U1 ( .INP(n10679), .ZN(U6072_n1) );
  AND2X1 U6073_U2 ( .IN1(WX7144), .IN2(U6073_n1), .Q(WX7207) );
  INVX0 U6073_U1 ( .INP(n10679), .ZN(U6073_n1) );
  AND2X1 U6074_U2 ( .IN1(WX7142), .IN2(U6074_n1), .Q(WX7205) );
  INVX0 U6074_U1 ( .INP(n10678), .ZN(U6074_n1) );
  AND2X1 U6075_U2 ( .IN1(WX6007), .IN2(U6075_n1), .Q(WX6070) );
  INVX0 U6075_U1 ( .INP(n10678), .ZN(U6075_n1) );
  AND2X1 U6076_U2 ( .IN1(test_so51), .IN2(U6076_n1), .Q(WX6068) );
  INVX0 U6076_U1 ( .INP(n10678), .ZN(U6076_n1) );
  AND2X1 U6077_U2 ( .IN1(WX6003), .IN2(U6077_n1), .Q(WX6066) );
  INVX0 U6077_U1 ( .INP(n10678), .ZN(U6077_n1) );
  AND2X1 U6078_U2 ( .IN1(WX6001), .IN2(U6078_n1), .Q(WX6064) );
  INVX0 U6078_U1 ( .INP(n10678), .ZN(U6078_n1) );
  AND2X1 U6079_U2 ( .IN1(WX5999), .IN2(U6079_n1), .Q(WX6062) );
  INVX0 U6079_U1 ( .INP(n10678), .ZN(U6079_n1) );
  AND2X1 U6080_U2 ( .IN1(WX5997), .IN2(U6080_n1), .Q(WX6060) );
  INVX0 U6080_U1 ( .INP(n10678), .ZN(U6080_n1) );
  AND2X1 U6081_U2 ( .IN1(WX5995), .IN2(U6081_n1), .Q(WX6058) );
  INVX0 U6081_U1 ( .INP(n10678), .ZN(U6081_n1) );
  AND2X1 U6082_U2 ( .IN1(WX5993), .IN2(U6082_n1), .Q(WX6056) );
  INVX0 U6082_U1 ( .INP(n10678), .ZN(U6082_n1) );
  AND2X1 U6083_U2 ( .IN1(WX5991), .IN2(U6083_n1), .Q(WX6054) );
  INVX0 U6083_U1 ( .INP(n10678), .ZN(U6083_n1) );
  AND2X1 U6084_U2 ( .IN1(WX5989), .IN2(U6084_n1), .Q(WX6052) );
  INVX0 U6084_U1 ( .INP(n10678), .ZN(U6084_n1) );
  AND2X1 U6085_U2 ( .IN1(WX5987), .IN2(U6085_n1), .Q(WX6050) );
  INVX0 U6085_U1 ( .INP(n10678), .ZN(U6085_n1) );
  AND2X1 U6086_U2 ( .IN1(WX5985), .IN2(U6086_n1), .Q(WX6048) );
  INVX0 U6086_U1 ( .INP(n10678), .ZN(U6086_n1) );
  AND2X1 U6087_U2 ( .IN1(WX5983), .IN2(U6087_n1), .Q(WX6046) );
  INVX0 U6087_U1 ( .INP(n10678), .ZN(U6087_n1) );
  AND2X1 U6088_U2 ( .IN1(WX5981), .IN2(U6088_n1), .Q(WX6044) );
  INVX0 U6088_U1 ( .INP(n10677), .ZN(U6088_n1) );
  AND2X1 U6089_U2 ( .IN1(WX5979), .IN2(U6089_n1), .Q(WX6042) );
  INVX0 U6089_U1 ( .INP(n10677), .ZN(U6089_n1) );
  AND2X1 U6090_U2 ( .IN1(WX5977), .IN2(U6090_n1), .Q(WX6040) );
  INVX0 U6090_U1 ( .INP(n10677), .ZN(U6090_n1) );
  AND2X1 U6091_U2 ( .IN1(WX5975), .IN2(U6091_n1), .Q(WX6038) );
  INVX0 U6091_U1 ( .INP(n10677), .ZN(U6091_n1) );
  AND2X1 U6092_U2 ( .IN1(WX5973), .IN2(U6092_n1), .Q(WX6036) );
  INVX0 U6092_U1 ( .INP(n10677), .ZN(U6092_n1) );
  AND2X1 U6093_U2 ( .IN1(test_so50), .IN2(U6093_n1), .Q(WX6034) );
  INVX0 U6093_U1 ( .INP(n10677), .ZN(U6093_n1) );
  AND2X1 U6094_U2 ( .IN1(WX5969), .IN2(U6094_n1), .Q(WX6032) );
  INVX0 U6094_U1 ( .INP(n10677), .ZN(U6094_n1) );
  AND2X1 U6095_U2 ( .IN1(WX5967), .IN2(U6095_n1), .Q(WX6030) );
  INVX0 U6095_U1 ( .INP(n10677), .ZN(U6095_n1) );
  AND2X1 U6096_U2 ( .IN1(WX5965), .IN2(U6096_n1), .Q(WX6028) );
  INVX0 U6096_U1 ( .INP(n10677), .ZN(U6096_n1) );
  AND2X1 U6097_U2 ( .IN1(WX5963), .IN2(U6097_n1), .Q(WX6026) );
  INVX0 U6097_U1 ( .INP(n10677), .ZN(U6097_n1) );
  AND2X1 U6098_U2 ( .IN1(WX5961), .IN2(U6098_n1), .Q(WX6024) );
  INVX0 U6098_U1 ( .INP(n10677), .ZN(U6098_n1) );
  AND2X1 U6099_U2 ( .IN1(WX5959), .IN2(U6099_n1), .Q(WX6022) );
  INVX0 U6099_U1 ( .INP(n10677), .ZN(U6099_n1) );
  AND2X1 U6100_U2 ( .IN1(WX5957), .IN2(U6100_n1), .Q(WX6020) );
  INVX0 U6100_U1 ( .INP(n10677), .ZN(U6100_n1) );
  AND2X1 U6101_U2 ( .IN1(WX5955), .IN2(U6101_n1), .Q(WX6018) );
  INVX0 U6101_U1 ( .INP(n10677), .ZN(U6101_n1) );
  AND2X1 U6102_U2 ( .IN1(WX5953), .IN2(U6102_n1), .Q(WX6016) );
  INVX0 U6102_U1 ( .INP(n10676), .ZN(U6102_n1) );
  AND2X1 U6103_U2 ( .IN1(WX5951), .IN2(U6103_n1), .Q(WX6014) );
  INVX0 U6103_U1 ( .INP(n10676), .ZN(U6103_n1) );
  AND2X1 U6104_U2 ( .IN1(WX5949), .IN2(U6104_n1), .Q(WX6012) );
  INVX0 U6104_U1 ( .INP(n10676), .ZN(U6104_n1) );
  AND2X1 U6105_U2 ( .IN1(WX5947), .IN2(U6105_n1), .Q(WX6010) );
  INVX0 U6105_U1 ( .INP(n10676), .ZN(U6105_n1) );
  AND2X1 U6106_U2 ( .IN1(WX5945), .IN2(U6106_n1), .Q(WX6008) );
  INVX0 U6106_U1 ( .INP(n10676), .ZN(U6106_n1) );
  AND2X1 U6107_U2 ( .IN1(WX5943), .IN2(U6107_n1), .Q(WX6006) );
  INVX0 U6107_U1 ( .INP(n10676), .ZN(U6107_n1) );
  AND2X1 U6108_U2 ( .IN1(WX5941), .IN2(U6108_n1), .Q(WX6004) );
  INVX0 U6108_U1 ( .INP(n10676), .ZN(U6108_n1) );
  AND2X1 U6109_U2 ( .IN1(WX5929), .IN2(U6109_n1), .Q(WX5992) );
  INVX0 U6109_U1 ( .INP(n10676), .ZN(U6109_n1) );
  AND2X1 U6110_U2 ( .IN1(WX5927), .IN2(U6110_n1), .Q(WX5990) );
  INVX0 U6110_U1 ( .INP(n10676), .ZN(U6110_n1) );
  AND2X1 U6111_U2 ( .IN1(WX5925), .IN2(U6111_n1), .Q(WX5988) );
  INVX0 U6111_U1 ( .INP(n10676), .ZN(U6111_n1) );
  AND2X1 U6112_U2 ( .IN1(WX5923), .IN2(U6112_n1), .Q(WX5986) );
  INVX0 U6112_U1 ( .INP(n10676), .ZN(U6112_n1) );
  AND2X1 U6113_U2 ( .IN1(WX5921), .IN2(U6113_n1), .Q(WX5984) );
  INVX0 U6113_U1 ( .INP(n10676), .ZN(U6113_n1) );
  AND2X1 U6114_U2 ( .IN1(WX5919), .IN2(U6114_n1), .Q(WX5982) );
  INVX0 U6114_U1 ( .INP(n10676), .ZN(U6114_n1) );
  AND2X1 U6115_U2 ( .IN1(WX5917), .IN2(U6115_n1), .Q(WX5980) );
  INVX0 U6115_U1 ( .INP(n10676), .ZN(U6115_n1) );
  AND2X1 U6116_U2 ( .IN1(WX5915), .IN2(U6116_n1), .Q(WX5978) );
  INVX0 U6116_U1 ( .INP(n10675), .ZN(U6116_n1) );
  AND2X1 U6117_U2 ( .IN1(WX5913), .IN2(U6117_n1), .Q(WX5976) );
  INVX0 U6117_U1 ( .INP(n10675), .ZN(U6117_n1) );
  AND2X1 U6118_U2 ( .IN1(WX5911), .IN2(U6118_n1), .Q(WX5974) );
  INVX0 U6118_U1 ( .INP(n10675), .ZN(U6118_n1) );
  AND2X1 U6119_U2 ( .IN1(WX5909), .IN2(U6119_n1), .Q(WX5972) );
  INVX0 U6119_U1 ( .INP(n10675), .ZN(U6119_n1) );
  AND2X1 U6120_U2 ( .IN1(WX5907), .IN2(U6120_n1), .Q(WX5970) );
  INVX0 U6120_U1 ( .INP(n10675), .ZN(U6120_n1) );
  AND2X1 U6121_U2 ( .IN1(WX5905), .IN2(U6121_n1), .Q(WX5968) );
  INVX0 U6121_U1 ( .INP(n10675), .ZN(U6121_n1) );
  AND2X1 U6122_U2 ( .IN1(test_so48), .IN2(U6122_n1), .Q(WX5966) );
  INVX0 U6122_U1 ( .INP(n10675), .ZN(U6122_n1) );
  AND2X1 U6123_U2 ( .IN1(WX5901), .IN2(U6123_n1), .Q(WX5964) );
  INVX0 U6123_U1 ( .INP(n10675), .ZN(U6123_n1) );
  AND2X1 U6124_U2 ( .IN1(WX5899), .IN2(U6124_n1), .Q(WX5962) );
  INVX0 U6124_U1 ( .INP(n10675), .ZN(U6124_n1) );
  AND2X1 U6125_U2 ( .IN1(WX5897), .IN2(U6125_n1), .Q(WX5960) );
  INVX0 U6125_U1 ( .INP(n10675), .ZN(U6125_n1) );
  AND2X1 U6126_U2 ( .IN1(WX5895), .IN2(U6126_n1), .Q(WX5958) );
  INVX0 U6126_U1 ( .INP(n10675), .ZN(U6126_n1) );
  AND2X1 U6127_U2 ( .IN1(WX5893), .IN2(U6127_n1), .Q(WX5956) );
  INVX0 U6127_U1 ( .INP(n10675), .ZN(U6127_n1) );
  AND2X1 U6128_U2 ( .IN1(WX5891), .IN2(U6128_n1), .Q(WX5954) );
  INVX0 U6128_U1 ( .INP(n10675), .ZN(U6128_n1) );
  AND2X1 U6129_U2 ( .IN1(WX5889), .IN2(U6129_n1), .Q(WX5952) );
  INVX0 U6129_U1 ( .INP(n10675), .ZN(U6129_n1) );
  AND2X1 U6130_U2 ( .IN1(WX5887), .IN2(U6130_n1), .Q(WX5950) );
  INVX0 U6130_U1 ( .INP(n10674), .ZN(U6130_n1) );
  AND2X1 U6131_U2 ( .IN1(WX5885), .IN2(U6131_n1), .Q(WX5948) );
  INVX0 U6131_U1 ( .INP(n10674), .ZN(U6131_n1) );
  AND2X1 U6132_U2 ( .IN1(WX5883), .IN2(U6132_n1), .Q(WX5946) );
  INVX0 U6132_U1 ( .INP(n10674), .ZN(U6132_n1) );
  AND2X1 U6133_U2 ( .IN1(WX5881), .IN2(U6133_n1), .Q(WX5944) );
  INVX0 U6133_U1 ( .INP(n10674), .ZN(U6133_n1) );
  AND2X1 U6134_U2 ( .IN1(WX5879), .IN2(U6134_n1), .Q(WX5942) );
  INVX0 U6134_U1 ( .INP(n10674), .ZN(U6134_n1) );
  AND2X1 U6135_U2 ( .IN1(WX5877), .IN2(U6135_n1), .Q(WX5940) );
  INVX0 U6135_U1 ( .INP(n10674), .ZN(U6135_n1) );
  AND2X1 U6136_U2 ( .IN1(WX5875), .IN2(U6136_n1), .Q(WX5938) );
  INVX0 U6136_U1 ( .INP(n10674), .ZN(U6136_n1) );
  AND2X1 U6137_U2 ( .IN1(WX5873), .IN2(U6137_n1), .Q(WX5936) );
  INVX0 U6137_U1 ( .INP(n10674), .ZN(U6137_n1) );
  AND2X1 U6138_U2 ( .IN1(WX5871), .IN2(U6138_n1), .Q(WX5934) );
  INVX0 U6138_U1 ( .INP(n10674), .ZN(U6138_n1) );
  AND2X1 U6139_U2 ( .IN1(test_so47), .IN2(U6139_n1), .Q(WX5932) );
  INVX0 U6139_U1 ( .INP(n10674), .ZN(U6139_n1) );
  AND2X1 U6140_U2 ( .IN1(WX5867), .IN2(U6140_n1), .Q(WX5930) );
  INVX0 U6140_U1 ( .INP(n10674), .ZN(U6140_n1) );
  AND2X1 U6141_U2 ( .IN1(WX5865), .IN2(U6141_n1), .Q(WX5928) );
  INVX0 U6141_U1 ( .INP(n10674), .ZN(U6141_n1) );
  AND2X1 U6142_U2 ( .IN1(WX5863), .IN2(U6142_n1), .Q(WX5926) );
  INVX0 U6142_U1 ( .INP(n10674), .ZN(U6142_n1) );
  AND2X1 U6143_U2 ( .IN1(WX5861), .IN2(U6143_n1), .Q(WX5924) );
  INVX0 U6143_U1 ( .INP(n10674), .ZN(U6143_n1) );
  AND2X1 U6144_U2 ( .IN1(WX5859), .IN2(U6144_n1), .Q(WX5922) );
  INVX0 U6144_U1 ( .INP(n10673), .ZN(U6144_n1) );
  AND2X1 U6145_U2 ( .IN1(WX5857), .IN2(U6145_n1), .Q(WX5920) );
  INVX0 U6145_U1 ( .INP(n10673), .ZN(U6145_n1) );
  AND2X1 U6146_U2 ( .IN1(WX5855), .IN2(U6146_n1), .Q(WX5918) );
  INVX0 U6146_U1 ( .INP(n10673), .ZN(U6146_n1) );
  AND2X1 U6147_U2 ( .IN1(WX5853), .IN2(U6147_n1), .Q(WX5916) );
  INVX0 U6147_U1 ( .INP(n10673), .ZN(U6147_n1) );
  AND2X1 U6148_U2 ( .IN1(WX5851), .IN2(U6148_n1), .Q(WX5914) );
  INVX0 U6148_U1 ( .INP(n10673), .ZN(U6148_n1) );
  AND2X1 U6149_U2 ( .IN1(WX5849), .IN2(U6149_n1), .Q(WX5912) );
  INVX0 U6149_U1 ( .INP(n10673), .ZN(U6149_n1) );
  AND2X1 U6150_U2 ( .IN1(WX4714), .IN2(U6150_n1), .Q(WX4777) );
  INVX0 U6150_U1 ( .INP(n10673), .ZN(U6150_n1) );
  AND2X1 U6151_U2 ( .IN1(WX4712), .IN2(U6151_n1), .Q(WX4775) );
  INVX0 U6151_U1 ( .INP(n10673), .ZN(U6151_n1) );
  AND2X1 U6152_U2 ( .IN1(WX4710), .IN2(U6152_n1), .Q(WX4773) );
  INVX0 U6152_U1 ( .INP(n10673), .ZN(U6152_n1) );
  AND2X1 U6153_U2 ( .IN1(WX4708), .IN2(U6153_n1), .Q(WX4771) );
  INVX0 U6153_U1 ( .INP(n10673), .ZN(U6153_n1) );
  AND2X1 U6154_U2 ( .IN1(WX4706), .IN2(U6154_n1), .Q(WX4769) );
  INVX0 U6154_U1 ( .INP(n10673), .ZN(U6154_n1) );
  AND2X1 U6155_U2 ( .IN1(WX4704), .IN2(U6155_n1), .Q(WX4767) );
  INVX0 U6155_U1 ( .INP(n10673), .ZN(U6155_n1) );
  AND2X1 U6156_U2 ( .IN1(WX4702), .IN2(U6156_n1), .Q(WX4765) );
  INVX0 U6156_U1 ( .INP(n10673), .ZN(U6156_n1) );
  AND2X1 U6157_U2 ( .IN1(WX4700), .IN2(U6157_n1), .Q(WX4763) );
  INVX0 U6157_U1 ( .INP(n10673), .ZN(U6157_n1) );
  AND2X1 U6158_U2 ( .IN1(WX4698), .IN2(U6158_n1), .Q(WX4761) );
  INVX0 U6158_U1 ( .INP(n10672), .ZN(U6158_n1) );
  AND2X1 U6159_U2 ( .IN1(WX4696), .IN2(U6159_n1), .Q(WX4759) );
  INVX0 U6159_U1 ( .INP(n10672), .ZN(U6159_n1) );
  AND2X1 U6160_U2 ( .IN1(WX4694), .IN2(U6160_n1), .Q(WX4757) );
  INVX0 U6160_U1 ( .INP(n10672), .ZN(U6160_n1) );
  AND2X1 U6161_U2 ( .IN1(WX4692), .IN2(U6161_n1), .Q(WX4755) );
  INVX0 U6161_U1 ( .INP(n10672), .ZN(U6161_n1) );
  AND2X1 U6162_U2 ( .IN1(WX4690), .IN2(U6162_n1), .Q(WX4753) );
  INVX0 U6162_U1 ( .INP(n10672), .ZN(U6162_n1) );
  AND2X1 U6163_U2 ( .IN1(test_so39), .IN2(U6163_n1), .Q(WX4751) );
  INVX0 U6163_U1 ( .INP(n10672), .ZN(U6163_n1) );
  AND2X1 U6164_U2 ( .IN1(WX4686), .IN2(U6164_n1), .Q(WX4749) );
  INVX0 U6164_U1 ( .INP(n10672), .ZN(U6164_n1) );
  AND2X1 U6165_U2 ( .IN1(WX4684), .IN2(U6165_n1), .Q(WX4747) );
  INVX0 U6165_U1 ( .INP(n10672), .ZN(U6165_n1) );
  AND2X1 U6166_U2 ( .IN1(WX4682), .IN2(U6166_n1), .Q(WX4745) );
  INVX0 U6166_U1 ( .INP(n10672), .ZN(U6166_n1) );
  AND2X1 U6167_U2 ( .IN1(WX4680), .IN2(U6167_n1), .Q(WX4743) );
  INVX0 U6167_U1 ( .INP(n10672), .ZN(U6167_n1) );
  AND2X1 U6168_U2 ( .IN1(WX4678), .IN2(U6168_n1), .Q(WX4741) );
  INVX0 U6168_U1 ( .INP(n10672), .ZN(U6168_n1) );
  AND2X1 U6169_U2 ( .IN1(WX4676), .IN2(U6169_n1), .Q(WX4739) );
  INVX0 U6169_U1 ( .INP(n10672), .ZN(U6169_n1) );
  AND2X1 U6170_U2 ( .IN1(WX4674), .IN2(U6170_n1), .Q(WX4737) );
  INVX0 U6170_U1 ( .INP(n10672), .ZN(U6170_n1) );
  AND2X1 U6171_U2 ( .IN1(WX4672), .IN2(U6171_n1), .Q(WX4735) );
  INVX0 U6171_U1 ( .INP(n10672), .ZN(U6171_n1) );
  AND2X1 U6172_U2 ( .IN1(WX4670), .IN2(U6172_n1), .Q(WX4733) );
  INVX0 U6172_U1 ( .INP(n10671), .ZN(U6172_n1) );
  AND2X1 U6173_U2 ( .IN1(WX4668), .IN2(U6173_n1), .Q(WX4731) );
  INVX0 U6173_U1 ( .INP(n10671), .ZN(U6173_n1) );
  AND2X1 U6174_U2 ( .IN1(WX4666), .IN2(U6174_n1), .Q(WX4729) );
  INVX0 U6174_U1 ( .INP(n10671), .ZN(U6174_n1) );
  AND2X1 U6175_U2 ( .IN1(WX4664), .IN2(U6175_n1), .Q(WX4727) );
  INVX0 U6175_U1 ( .INP(n10671), .ZN(U6175_n1) );
  AND2X1 U6176_U2 ( .IN1(WX4662), .IN2(U6176_n1), .Q(WX4725) );
  INVX0 U6176_U1 ( .INP(n10671), .ZN(U6176_n1) );
  AND2X1 U6177_U2 ( .IN1(WX4660), .IN2(U6177_n1), .Q(WX4723) );
  INVX0 U6177_U1 ( .INP(n10671), .ZN(U6177_n1) );
  AND2X1 U6178_U2 ( .IN1(WX4658), .IN2(U6178_n1), .Q(WX4721) );
  INVX0 U6178_U1 ( .INP(n10671), .ZN(U6178_n1) );
  AND2X1 U6179_U2 ( .IN1(WX4656), .IN2(U6179_n1), .Q(WX4719) );
  INVX0 U6179_U1 ( .INP(n10671), .ZN(U6179_n1) );
  AND2X1 U6180_U2 ( .IN1(test_so38), .IN2(U6180_n1), .Q(WX4717) );
  INVX0 U6180_U1 ( .INP(n10671), .ZN(U6180_n1) );
  AND2X1 U6181_U2 ( .IN1(WX4652), .IN2(U6181_n1), .Q(WX4715) );
  INVX0 U6181_U1 ( .INP(n10671), .ZN(U6181_n1) );
  AND2X1 U6182_U2 ( .IN1(WX4650), .IN2(U6182_n1), .Q(WX4713) );
  INVX0 U6182_U1 ( .INP(n10671), .ZN(U6182_n1) );
  AND2X1 U6183_U2 ( .IN1(WX4648), .IN2(U6183_n1), .Q(WX4711) );
  INVX0 U6183_U1 ( .INP(n10671), .ZN(U6183_n1) );
  AND2X1 U6184_U2 ( .IN1(WX4646), .IN2(U6184_n1), .Q(WX4709) );
  INVX0 U6184_U1 ( .INP(n10671), .ZN(U6184_n1) );
  AND2X1 U6185_U2 ( .IN1(WX4644), .IN2(U6185_n1), .Q(WX4707) );
  INVX0 U6185_U1 ( .INP(n10671), .ZN(U6185_n1) );
  AND2X1 U6186_U2 ( .IN1(WX4642), .IN2(U6186_n1), .Q(WX4705) );
  INVX0 U6186_U1 ( .INP(n10670), .ZN(U6186_n1) );
  AND2X1 U6187_U2 ( .IN1(WX4640), .IN2(U6187_n1), .Q(WX4703) );
  INVX0 U6187_U1 ( .INP(n10670), .ZN(U6187_n1) );
  AND2X1 U6188_U2 ( .IN1(WX4638), .IN2(U6188_n1), .Q(WX4701) );
  INVX0 U6188_U1 ( .INP(n10670), .ZN(U6188_n1) );
  AND2X1 U6189_U2 ( .IN1(WX4636), .IN2(U6189_n1), .Q(WX4699) );
  INVX0 U6189_U1 ( .INP(n10670), .ZN(U6189_n1) );
  AND2X1 U6190_U2 ( .IN1(WX4634), .IN2(U6190_n1), .Q(WX4697) );
  INVX0 U6190_U1 ( .INP(n10670), .ZN(U6190_n1) );
  AND2X1 U6191_U2 ( .IN1(WX4632), .IN2(U6191_n1), .Q(WX4695) );
  INVX0 U6191_U1 ( .INP(n10670), .ZN(U6191_n1) );
  AND2X1 U6192_U2 ( .IN1(WX4630), .IN2(U6192_n1), .Q(WX4693) );
  INVX0 U6192_U1 ( .INP(n10670), .ZN(U6192_n1) );
  AND2X1 U6193_U2 ( .IN1(WX4628), .IN2(U6193_n1), .Q(WX4691) );
  INVX0 U6193_U1 ( .INP(n10670), .ZN(U6193_n1) );
  AND2X1 U6194_U2 ( .IN1(WX4626), .IN2(U6194_n1), .Q(WX4689) );
  INVX0 U6194_U1 ( .INP(n10670), .ZN(U6194_n1) );
  AND2X1 U6195_U2 ( .IN1(WX4624), .IN2(U6195_n1), .Q(WX4687) );
  INVX0 U6195_U1 ( .INP(n10670), .ZN(U6195_n1) );
  AND2X1 U6196_U2 ( .IN1(WX4622), .IN2(U6196_n1), .Q(WX4685) );
  INVX0 U6196_U1 ( .INP(n10670), .ZN(U6196_n1) );
  AND2X1 U6197_U2 ( .IN1(test_so37), .IN2(U6197_n1), .Q(WX4683) );
  INVX0 U6197_U1 ( .INP(n10670), .ZN(U6197_n1) );
  AND2X1 U6198_U2 ( .IN1(WX4618), .IN2(U6198_n1), .Q(WX4681) );
  INVX0 U6198_U1 ( .INP(n10670), .ZN(U6198_n1) );
  AND2X1 U6199_U2 ( .IN1(WX4616), .IN2(U6199_n1), .Q(WX4679) );
  INVX0 U6199_U1 ( .INP(n10670), .ZN(U6199_n1) );
  AND2X1 U6200_U2 ( .IN1(WX4614), .IN2(U6200_n1), .Q(WX4677) );
  INVX0 U6200_U1 ( .INP(n10669), .ZN(U6200_n1) );
  AND2X1 U6201_U2 ( .IN1(WX4612), .IN2(U6201_n1), .Q(WX4675) );
  INVX0 U6201_U1 ( .INP(n10669), .ZN(U6201_n1) );
  AND2X1 U6202_U2 ( .IN1(WX4610), .IN2(U6202_n1), .Q(WX4673) );
  INVX0 U6202_U1 ( .INP(n10669), .ZN(U6202_n1) );
  AND2X1 U6203_U2 ( .IN1(WX4608), .IN2(U6203_n1), .Q(WX4671) );
  INVX0 U6203_U1 ( .INP(n10669), .ZN(U6203_n1) );
  AND2X1 U6204_U2 ( .IN1(WX4606), .IN2(U6204_n1), .Q(WX4669) );
  INVX0 U6204_U1 ( .INP(n10669), .ZN(U6204_n1) );
  AND2X1 U6205_U2 ( .IN1(WX4604), .IN2(U6205_n1), .Q(WX4667) );
  INVX0 U6205_U1 ( .INP(n10669), .ZN(U6205_n1) );
  AND2X1 U6206_U2 ( .IN1(WX4602), .IN2(U6206_n1), .Q(WX4665) );
  INVX0 U6206_U1 ( .INP(n10669), .ZN(U6206_n1) );
  AND2X1 U6207_U2 ( .IN1(WX4600), .IN2(U6207_n1), .Q(WX4663) );
  INVX0 U6207_U1 ( .INP(n10669), .ZN(U6207_n1) );
  AND2X1 U6208_U2 ( .IN1(WX4598), .IN2(U6208_n1), .Q(WX4661) );
  INVX0 U6208_U1 ( .INP(n10669), .ZN(U6208_n1) );
  AND2X1 U6209_U2 ( .IN1(WX4596), .IN2(U6209_n1), .Q(WX4659) );
  INVX0 U6209_U1 ( .INP(n10669), .ZN(U6209_n1) );
  AND2X1 U6210_U2 ( .IN1(WX4594), .IN2(U6210_n1), .Q(WX4657) );
  INVX0 U6210_U1 ( .INP(n10669), .ZN(U6210_n1) );
  AND2X1 U6211_U2 ( .IN1(WX4592), .IN2(U6211_n1), .Q(WX4655) );
  INVX0 U6211_U1 ( .INP(n10669), .ZN(U6211_n1) );
  AND2X1 U6212_U2 ( .IN1(WX4590), .IN2(U6212_n1), .Q(WX4653) );
  INVX0 U6212_U1 ( .INP(n10669), .ZN(U6212_n1) );
  AND2X1 U6213_U2 ( .IN1(WX4588), .IN2(U6213_n1), .Q(WX4651) );
  INVX0 U6213_U1 ( .INP(n10669), .ZN(U6213_n1) );
  AND2X1 U6214_U2 ( .IN1(test_so36), .IN2(U6214_n1), .Q(WX4649) );
  INVX0 U6214_U1 ( .INP(n10668), .ZN(U6214_n1) );
  AND2X1 U6215_U2 ( .IN1(WX4584), .IN2(U6215_n1), .Q(WX4647) );
  INVX0 U6215_U1 ( .INP(n10668), .ZN(U6215_n1) );
  AND2X1 U6216_U2 ( .IN1(WX4582), .IN2(U6216_n1), .Q(WX4645) );
  INVX0 U6216_U1 ( .INP(n10668), .ZN(U6216_n1) );
  AND2X1 U6217_U2 ( .IN1(WX4580), .IN2(U6217_n1), .Q(WX4643) );
  INVX0 U6217_U1 ( .INP(n10668), .ZN(U6217_n1) );
  AND2X1 U6218_U2 ( .IN1(WX4578), .IN2(U6218_n1), .Q(WX4641) );
  INVX0 U6218_U1 ( .INP(n10668), .ZN(U6218_n1) );
  AND2X1 U6219_U2 ( .IN1(WX4576), .IN2(U6219_n1), .Q(WX4639) );
  INVX0 U6219_U1 ( .INP(n10668), .ZN(U6219_n1) );
  AND2X1 U6220_U2 ( .IN1(WX4574), .IN2(U6220_n1), .Q(WX4637) );
  INVX0 U6220_U1 ( .INP(n10668), .ZN(U6220_n1) );
  AND2X1 U6221_U2 ( .IN1(WX4572), .IN2(U6221_n1), .Q(WX4635) );
  INVX0 U6221_U1 ( .INP(n10668), .ZN(U6221_n1) );
  AND2X1 U6222_U2 ( .IN1(WX4570), .IN2(U6222_n1), .Q(WX4633) );
  INVX0 U6222_U1 ( .INP(n10668), .ZN(U6222_n1) );
  AND2X1 U6223_U2 ( .IN1(WX4568), .IN2(U6223_n1), .Q(WX4631) );
  INVX0 U6223_U1 ( .INP(n10668), .ZN(U6223_n1) );
  AND2X1 U6224_U2 ( .IN1(WX4566), .IN2(U6224_n1), .Q(WX4629) );
  INVX0 U6224_U1 ( .INP(n10668), .ZN(U6224_n1) );
  AND2X1 U6225_U2 ( .IN1(WX4564), .IN2(U6225_n1), .Q(WX4627) );
  INVX0 U6225_U1 ( .INP(n10668), .ZN(U6225_n1) );
  AND2X1 U6226_U2 ( .IN1(WX4562), .IN2(U6226_n1), .Q(WX4625) );
  INVX0 U6226_U1 ( .INP(n10668), .ZN(U6226_n1) );
  AND2X1 U6227_U2 ( .IN1(WX4560), .IN2(U6227_n1), .Q(WX4623) );
  INVX0 U6227_U1 ( .INP(n10668), .ZN(U6227_n1) );
  AND2X1 U6228_U2 ( .IN1(WX4558), .IN2(U6228_n1), .Q(WX4621) );
  INVX0 U6228_U1 ( .INP(n10667), .ZN(U6228_n1) );
  AND2X1 U6229_U2 ( .IN1(WX4556), .IN2(U6229_n1), .Q(WX4619) );
  INVX0 U6229_U1 ( .INP(n10667), .ZN(U6229_n1) );
  AND2X1 U6230_U2 ( .IN1(WX3421), .IN2(U6230_n1), .Q(WX3484) );
  INVX0 U6230_U1 ( .INP(n10667), .ZN(U6230_n1) );
  AND2X1 U6231_U2 ( .IN1(WX3419), .IN2(U6231_n1), .Q(WX3482) );
  INVX0 U6231_U1 ( .INP(n10667), .ZN(U6231_n1) );
  AND2X1 U6232_U2 ( .IN1(WX3417), .IN2(U6232_n1), .Q(WX3480) );
  INVX0 U6232_U1 ( .INP(n10667), .ZN(U6232_n1) );
  AND2X1 U6233_U2 ( .IN1(WX3415), .IN2(U6233_n1), .Q(WX3478) );
  INVX0 U6233_U1 ( .INP(n10667), .ZN(U6233_n1) );
  AND2X1 U6234_U2 ( .IN1(WX3413), .IN2(U6234_n1), .Q(WX3476) );
  INVX0 U6234_U1 ( .INP(n10667), .ZN(U6234_n1) );
  AND2X1 U6235_U2 ( .IN1(WX3411), .IN2(U6235_n1), .Q(WX3474) );
  INVX0 U6235_U1 ( .INP(n10667), .ZN(U6235_n1) );
  AND2X1 U6236_U2 ( .IN1(WX3409), .IN2(U6236_n1), .Q(WX3472) );
  INVX0 U6236_U1 ( .INP(n10667), .ZN(U6236_n1) );
  AND2X1 U6237_U2 ( .IN1(WX3407), .IN2(U6237_n1), .Q(WX3470) );
  INVX0 U6237_U1 ( .INP(n10667), .ZN(U6237_n1) );
  AND2X1 U6238_U2 ( .IN1(test_so28), .IN2(U6238_n1), .Q(WX3468) );
  INVX0 U6238_U1 ( .INP(n10667), .ZN(U6238_n1) );
  AND2X1 U6239_U2 ( .IN1(WX3403), .IN2(U6239_n1), .Q(WX3466) );
  INVX0 U6239_U1 ( .INP(n10667), .ZN(U6239_n1) );
  AND2X1 U6240_U2 ( .IN1(WX3401), .IN2(U6240_n1), .Q(WX3464) );
  INVX0 U6240_U1 ( .INP(n10667), .ZN(U6240_n1) );
  AND2X1 U6241_U2 ( .IN1(WX3399), .IN2(U6241_n1), .Q(WX3462) );
  INVX0 U6241_U1 ( .INP(n10667), .ZN(U6241_n1) );
  AND2X1 U6242_U2 ( .IN1(WX3397), .IN2(U6242_n1), .Q(WX3460) );
  INVX0 U6242_U1 ( .INP(n10666), .ZN(U6242_n1) );
  AND2X1 U6243_U2 ( .IN1(WX3395), .IN2(U6243_n1), .Q(WX3458) );
  INVX0 U6243_U1 ( .INP(n10666), .ZN(U6243_n1) );
  AND2X1 U6244_U2 ( .IN1(WX3393), .IN2(U6244_n1), .Q(WX3456) );
  INVX0 U6244_U1 ( .INP(n10666), .ZN(U6244_n1) );
  AND2X1 U6245_U2 ( .IN1(WX3391), .IN2(U6245_n1), .Q(WX3454) );
  INVX0 U6245_U1 ( .INP(n10666), .ZN(U6245_n1) );
  AND2X1 U6246_U2 ( .IN1(WX3389), .IN2(U6246_n1), .Q(WX3452) );
  INVX0 U6246_U1 ( .INP(n10666), .ZN(U6246_n1) );
  AND2X1 U6247_U2 ( .IN1(WX3387), .IN2(U6247_n1), .Q(WX3450) );
  INVX0 U6247_U1 ( .INP(n10666), .ZN(U6247_n1) );
  AND2X1 U6248_U2 ( .IN1(WX3385), .IN2(U6248_n1), .Q(WX3448) );
  INVX0 U6248_U1 ( .INP(n10666), .ZN(U6248_n1) );
  AND2X1 U6249_U2 ( .IN1(WX3383), .IN2(U6249_n1), .Q(WX3446) );
  INVX0 U6249_U1 ( .INP(n10666), .ZN(U6249_n1) );
  AND2X1 U6250_U2 ( .IN1(WX3381), .IN2(U6250_n1), .Q(WX3444) );
  INVX0 U6250_U1 ( .INP(n10666), .ZN(U6250_n1) );
  AND2X1 U6251_U2 ( .IN1(WX3379), .IN2(U6251_n1), .Q(WX3442) );
  INVX0 U6251_U1 ( .INP(n10666), .ZN(U6251_n1) );
  AND2X1 U6252_U2 ( .IN1(WX3377), .IN2(U6252_n1), .Q(WX3440) );
  INVX0 U6252_U1 ( .INP(n10666), .ZN(U6252_n1) );
  AND2X1 U6253_U2 ( .IN1(WX3375), .IN2(U6253_n1), .Q(WX3438) );
  INVX0 U6253_U1 ( .INP(n10666), .ZN(U6253_n1) );
  AND2X1 U6254_U2 ( .IN1(WX3373), .IN2(U6254_n1), .Q(WX3436) );
  INVX0 U6254_U1 ( .INP(n10666), .ZN(U6254_n1) );
  AND2X1 U6255_U2 ( .IN1(WX3371), .IN2(U6255_n1), .Q(WX3434) );
  INVX0 U6255_U1 ( .INP(n10666), .ZN(U6255_n1) );
  AND2X1 U6256_U2 ( .IN1(test_so27), .IN2(U6256_n1), .Q(WX3432) );
  INVX0 U6256_U1 ( .INP(n10665), .ZN(U6256_n1) );
  AND2X1 U6257_U2 ( .IN1(WX3367), .IN2(U6257_n1), .Q(WX3430) );
  INVX0 U6257_U1 ( .INP(n10665), .ZN(U6257_n1) );
  AND2X1 U6258_U2 ( .IN1(WX3365), .IN2(U6258_n1), .Q(WX3428) );
  INVX0 U6258_U1 ( .INP(n10665), .ZN(U6258_n1) );
  AND2X1 U6259_U2 ( .IN1(WX3363), .IN2(U6259_n1), .Q(WX3426) );
  INVX0 U6259_U1 ( .INP(n10665), .ZN(U6259_n1) );
  AND2X1 U6260_U2 ( .IN1(WX3361), .IN2(U6260_n1), .Q(WX3424) );
  INVX0 U6260_U1 ( .INP(n10665), .ZN(U6260_n1) );
  AND2X1 U6261_U2 ( .IN1(WX3359), .IN2(U6261_n1), .Q(WX3422) );
  INVX0 U6261_U1 ( .INP(n10665), .ZN(U6261_n1) );
  AND2X1 U6262_U2 ( .IN1(WX3357), .IN2(U6262_n1), .Q(WX3420) );
  INVX0 U6262_U1 ( .INP(n10665), .ZN(U6262_n1) );
  AND2X1 U6263_U2 ( .IN1(WX3355), .IN2(U6263_n1), .Q(WX3418) );
  INVX0 U6263_U1 ( .INP(n10665), .ZN(U6263_n1) );
  AND2X1 U6264_U2 ( .IN1(WX3353), .IN2(U6264_n1), .Q(WX3416) );
  INVX0 U6264_U1 ( .INP(n10665), .ZN(U6264_n1) );
  AND2X1 U6265_U2 ( .IN1(WX3351), .IN2(U6265_n1), .Q(WX3414) );
  INVX0 U6265_U1 ( .INP(n10665), .ZN(U6265_n1) );
  AND2X1 U6266_U2 ( .IN1(WX3349), .IN2(U6266_n1), .Q(WX3412) );
  INVX0 U6266_U1 ( .INP(n10665), .ZN(U6266_n1) );
  AND2X1 U6267_U2 ( .IN1(WX3347), .IN2(U6267_n1), .Q(WX3410) );
  INVX0 U6267_U1 ( .INP(n10665), .ZN(U6267_n1) );
  AND2X1 U6268_U2 ( .IN1(WX3345), .IN2(U6268_n1), .Q(WX3408) );
  INVX0 U6268_U1 ( .INP(n10665), .ZN(U6268_n1) );
  AND2X1 U6269_U2 ( .IN1(WX3343), .IN2(U6269_n1), .Q(WX3406) );
  INVX0 U6269_U1 ( .INP(n10665), .ZN(U6269_n1) );
  AND2X1 U6270_U2 ( .IN1(WX3341), .IN2(U6270_n1), .Q(WX3404) );
  INVX0 U6270_U1 ( .INP(n10664), .ZN(U6270_n1) );
  AND2X1 U6271_U2 ( .IN1(WX3339), .IN2(U6271_n1), .Q(WX3402) );
  INVX0 U6271_U1 ( .INP(n10664), .ZN(U6271_n1) );
  AND2X1 U6272_U2 ( .IN1(WX3337), .IN2(U6272_n1), .Q(WX3400) );
  INVX0 U6272_U1 ( .INP(n10664), .ZN(U6272_n1) );
  AND2X1 U6273_U2 ( .IN1(WX3335), .IN2(U6273_n1), .Q(WX3398) );
  INVX0 U6273_U1 ( .INP(n10664), .ZN(U6273_n1) );
  AND2X1 U6274_U2 ( .IN1(test_so26), .IN2(U6274_n1), .Q(WX3396) );
  INVX0 U6274_U1 ( .INP(n10664), .ZN(U6274_n1) );
  AND2X1 U6275_U2 ( .IN1(WX3331), .IN2(U6275_n1), .Q(WX3394) );
  INVX0 U6275_U1 ( .INP(n10664), .ZN(U6275_n1) );
  AND2X1 U6276_U2 ( .IN1(WX3329), .IN2(U6276_n1), .Q(WX3392) );
  INVX0 U6276_U1 ( .INP(n10664), .ZN(U6276_n1) );
  AND2X1 U6277_U2 ( .IN1(WX3327), .IN2(U6277_n1), .Q(WX3390) );
  INVX0 U6277_U1 ( .INP(n10664), .ZN(U6277_n1) );
  AND2X1 U6278_U2 ( .IN1(WX3325), .IN2(U6278_n1), .Q(WX3388) );
  INVX0 U6278_U1 ( .INP(n10664), .ZN(U6278_n1) );
  AND2X1 U6279_U2 ( .IN1(WX3323), .IN2(U6279_n1), .Q(WX3386) );
  INVX0 U6279_U1 ( .INP(n10664), .ZN(U6279_n1) );
  AND2X1 U6280_U2 ( .IN1(WX3321), .IN2(U6280_n1), .Q(WX3384) );
  INVX0 U6280_U1 ( .INP(n10664), .ZN(U6280_n1) );
  AND2X1 U6281_U2 ( .IN1(WX3319), .IN2(U6281_n1), .Q(WX3382) );
  INVX0 U6281_U1 ( .INP(n10664), .ZN(U6281_n1) );
  AND2X1 U6282_U2 ( .IN1(WX3317), .IN2(U6282_n1), .Q(WX3380) );
  INVX0 U6282_U1 ( .INP(n10664), .ZN(U6282_n1) );
  AND2X1 U6283_U2 ( .IN1(WX3315), .IN2(U6283_n1), .Q(WX3378) );
  INVX0 U6283_U1 ( .INP(n10664), .ZN(U6283_n1) );
  AND2X1 U6284_U2 ( .IN1(WX3313), .IN2(U6284_n1), .Q(WX3376) );
  INVX0 U6284_U1 ( .INP(n10663), .ZN(U6284_n1) );
  AND2X1 U6285_U2 ( .IN1(WX3311), .IN2(U6285_n1), .Q(WX3374) );
  INVX0 U6285_U1 ( .INP(n10663), .ZN(U6285_n1) );
  AND2X1 U6286_U2 ( .IN1(WX3309), .IN2(U6286_n1), .Q(WX3372) );
  INVX0 U6286_U1 ( .INP(n10663), .ZN(U6286_n1) );
  AND2X1 U6287_U2 ( .IN1(WX3307), .IN2(U6287_n1), .Q(WX3370) );
  INVX0 U6287_U1 ( .INP(n10663), .ZN(U6287_n1) );
  AND2X1 U6288_U2 ( .IN1(WX3305), .IN2(U6288_n1), .Q(WX3368) );
  INVX0 U6288_U1 ( .INP(n10663), .ZN(U6288_n1) );
  AND2X1 U6289_U2 ( .IN1(WX3303), .IN2(U6289_n1), .Q(WX3366) );
  INVX0 U6289_U1 ( .INP(n10663), .ZN(U6289_n1) );
  AND2X1 U6290_U2 ( .IN1(WX3301), .IN2(U6290_n1), .Q(WX3364) );
  INVX0 U6290_U1 ( .INP(n10663), .ZN(U6290_n1) );
  AND2X1 U6291_U2 ( .IN1(WX3299), .IN2(U6291_n1), .Q(WX3362) );
  INVX0 U6291_U1 ( .INP(n10663), .ZN(U6291_n1) );
  AND2X1 U6292_U2 ( .IN1(test_so25), .IN2(U6292_n1), .Q(WX3360) );
  INVX0 U6292_U1 ( .INP(n10663), .ZN(U6292_n1) );
  AND2X1 U6293_U2 ( .IN1(WX3295), .IN2(U6293_n1), .Q(WX3358) );
  INVX0 U6293_U1 ( .INP(n10663), .ZN(U6293_n1) );
  AND2X1 U6294_U2 ( .IN1(WX3293), .IN2(U6294_n1), .Q(WX3356) );
  INVX0 U6294_U1 ( .INP(n10663), .ZN(U6294_n1) );
  AND2X1 U6295_U2 ( .IN1(WX3291), .IN2(U6295_n1), .Q(WX3354) );
  INVX0 U6295_U1 ( .INP(n10663), .ZN(U6295_n1) );
  AND2X1 U6296_U2 ( .IN1(WX3289), .IN2(U6296_n1), .Q(WX3352) );
  INVX0 U6296_U1 ( .INP(n10663), .ZN(U6296_n1) );
  AND2X1 U6297_U2 ( .IN1(WX3287), .IN2(U6297_n1), .Q(WX3350) );
  INVX0 U6297_U1 ( .INP(n10663), .ZN(U6297_n1) );
  AND2X1 U6298_U2 ( .IN1(WX3285), .IN2(U6298_n1), .Q(WX3348) );
  INVX0 U6298_U1 ( .INP(n10662), .ZN(U6298_n1) );
  AND2X1 U6299_U2 ( .IN1(WX3283), .IN2(U6299_n1), .Q(WX3346) );
  INVX0 U6299_U1 ( .INP(n10662), .ZN(U6299_n1) );
  AND2X1 U6300_U2 ( .IN1(WX3281), .IN2(U6300_n1), .Q(WX3344) );
  INVX0 U6300_U1 ( .INP(n10662), .ZN(U6300_n1) );
  AND2X1 U6301_U2 ( .IN1(WX3279), .IN2(U6301_n1), .Q(WX3342) );
  INVX0 U6301_U1 ( .INP(n10662), .ZN(U6301_n1) );
  AND2X1 U6302_U2 ( .IN1(WX3277), .IN2(U6302_n1), .Q(WX3340) );
  INVX0 U6302_U1 ( .INP(n10662), .ZN(U6302_n1) );
  AND2X1 U6303_U2 ( .IN1(WX3275), .IN2(U6303_n1), .Q(WX3338) );
  INVX0 U6303_U1 ( .INP(n10662), .ZN(U6303_n1) );
  AND2X1 U6304_U2 ( .IN1(WX3273), .IN2(U6304_n1), .Q(WX3336) );
  INVX0 U6304_U1 ( .INP(n10662), .ZN(U6304_n1) );
  AND2X1 U6305_U2 ( .IN1(WX3271), .IN2(U6305_n1), .Q(WX3334) );
  INVX0 U6305_U1 ( .INP(n10662), .ZN(U6305_n1) );
  AND2X1 U6306_U2 ( .IN1(WX3267), .IN2(U6306_n1), .Q(WX3330) );
  INVX0 U6306_U1 ( .INP(n10662), .ZN(U6306_n1) );
  AND2X1 U6307_U2 ( .IN1(WX2128), .IN2(U6307_n1), .Q(WX2191) );
  INVX0 U6307_U1 ( .INP(n10662), .ZN(U6307_n1) );
  AND2X1 U6308_U2 ( .IN1(WX2126), .IN2(U6308_n1), .Q(WX2189) );
  INVX0 U6308_U1 ( .INP(n10662), .ZN(U6308_n1) );
  AND2X1 U6309_U2 ( .IN1(WX2124), .IN2(U6309_n1), .Q(WX2187) );
  INVX0 U6309_U1 ( .INP(n10662), .ZN(U6309_n1) );
  AND2X1 U6310_U2 ( .IN1(WX2122), .IN2(U6310_n1), .Q(WX2185) );
  INVX0 U6310_U1 ( .INP(n10662), .ZN(U6310_n1) );
  AND2X1 U6311_U2 ( .IN1(WX2120), .IN2(U6311_n1), .Q(WX2183) );
  INVX0 U6311_U1 ( .INP(n10662), .ZN(U6311_n1) );
  AND2X1 U6312_U2 ( .IN1(WX2118), .IN2(U6312_n1), .Q(WX2181) );
  INVX0 U6312_U1 ( .INP(n10661), .ZN(U6312_n1) );
  AND2X1 U6313_U2 ( .IN1(WX2116), .IN2(U6313_n1), .Q(WX2179) );
  INVX0 U6313_U1 ( .INP(n10661), .ZN(U6313_n1) );
  AND2X1 U6314_U2 ( .IN1(WX2114), .IN2(U6314_n1), .Q(WX2177) );
  INVX0 U6314_U1 ( .INP(n10661), .ZN(U6314_n1) );
  AND2X1 U6315_U2 ( .IN1(WX2112), .IN2(U6315_n1), .Q(WX2175) );
  INVX0 U6315_U1 ( .INP(n10661), .ZN(U6315_n1) );
  AND2X1 U6316_U2 ( .IN1(WX2110), .IN2(U6316_n1), .Q(WX2173) );
  INVX0 U6316_U1 ( .INP(n10661), .ZN(U6316_n1) );
  AND2X1 U6317_U2 ( .IN1(WX2108), .IN2(U6317_n1), .Q(WX2171) );
  INVX0 U6317_U1 ( .INP(n10661), .ZN(U6317_n1) );
  AND2X1 U6318_U2 ( .IN1(WX2106), .IN2(U6318_n1), .Q(WX2169) );
  INVX0 U6318_U1 ( .INP(n10661), .ZN(U6318_n1) );
  AND2X1 U6319_U2 ( .IN1(WX2104), .IN2(U6319_n1), .Q(WX2167) );
  INVX0 U6319_U1 ( .INP(n10661), .ZN(U6319_n1) );
  AND2X1 U6320_U2 ( .IN1(WX2102), .IN2(U6320_n1), .Q(WX2165) );
  INVX0 U6320_U1 ( .INP(n10661), .ZN(U6320_n1) );
  AND2X1 U6321_U2 ( .IN1(test_so17), .IN2(U6321_n1), .Q(WX2163) );
  INVX0 U6321_U1 ( .INP(n10661), .ZN(U6321_n1) );
  AND2X1 U6322_U2 ( .IN1(WX2098), .IN2(U6322_n1), .Q(WX2161) );
  INVX0 U6322_U1 ( .INP(n10661), .ZN(U6322_n1) );
  AND2X1 U6323_U2 ( .IN1(WX2096), .IN2(U6323_n1), .Q(WX2159) );
  INVX0 U6323_U1 ( .INP(n10661), .ZN(U6323_n1) );
  AND2X1 U6324_U2 ( .IN1(WX2094), .IN2(U6324_n1), .Q(WX2157) );
  INVX0 U6324_U1 ( .INP(n10661), .ZN(U6324_n1) );
  AND2X1 U6325_U2 ( .IN1(WX2092), .IN2(U6325_n1), .Q(WX2155) );
  INVX0 U6325_U1 ( .INP(n10661), .ZN(U6325_n1) );
  AND2X1 U6326_U2 ( .IN1(WX2090), .IN2(U6326_n1), .Q(WX2153) );
  INVX0 U6326_U1 ( .INP(n10660), .ZN(U6326_n1) );
  AND2X1 U6327_U2 ( .IN1(WX2088), .IN2(U6327_n1), .Q(WX2151) );
  INVX0 U6327_U1 ( .INP(n10660), .ZN(U6327_n1) );
  AND2X1 U6328_U2 ( .IN1(WX2086), .IN2(U6328_n1), .Q(WX2149) );
  INVX0 U6328_U1 ( .INP(n10660), .ZN(U6328_n1) );
  AND2X1 U6329_U2 ( .IN1(WX2084), .IN2(U6329_n1), .Q(WX2147) );
  INVX0 U6329_U1 ( .INP(n10660), .ZN(U6329_n1) );
  AND2X1 U6330_U2 ( .IN1(WX2082), .IN2(U6330_n1), .Q(WX2145) );
  INVX0 U6330_U1 ( .INP(n10660), .ZN(U6330_n1) );
  AND2X1 U6331_U2 ( .IN1(WX2080), .IN2(U6331_n1), .Q(WX2143) );
  INVX0 U6331_U1 ( .INP(n10660), .ZN(U6331_n1) );
  AND2X1 U6332_U2 ( .IN1(WX2078), .IN2(U6332_n1), .Q(WX2141) );
  INVX0 U6332_U1 ( .INP(n10660), .ZN(U6332_n1) );
  AND2X1 U6333_U2 ( .IN1(WX2076), .IN2(U6333_n1), .Q(WX2139) );
  INVX0 U6333_U1 ( .INP(n10660), .ZN(U6333_n1) );
  AND2X1 U6334_U2 ( .IN1(WX2074), .IN2(U6334_n1), .Q(WX2137) );
  INVX0 U6334_U1 ( .INP(n10660), .ZN(U6334_n1) );
  AND2X1 U6335_U2 ( .IN1(WX2072), .IN2(U6335_n1), .Q(WX2135) );
  INVX0 U6335_U1 ( .INP(n10660), .ZN(U6335_n1) );
  AND2X1 U6336_U2 ( .IN1(WX2070), .IN2(U6336_n1), .Q(WX2133) );
  INVX0 U6336_U1 ( .INP(n10660), .ZN(U6336_n1) );
  AND2X1 U6337_U2 ( .IN1(WX2068), .IN2(U6337_n1), .Q(WX2131) );
  INVX0 U6337_U1 ( .INP(n10660), .ZN(U6337_n1) );
  AND2X1 U6338_U2 ( .IN1(WX2066), .IN2(U6338_n1), .Q(WX2129) );
  INVX0 U6338_U1 ( .INP(n10660), .ZN(U6338_n1) );
  AND2X1 U6339_U2 ( .IN1(test_so16), .IN2(U6339_n1), .Q(WX2127) );
  INVX0 U6339_U1 ( .INP(n10660), .ZN(U6339_n1) );
  AND2X1 U6340_U2 ( .IN1(WX2062), .IN2(U6340_n1), .Q(WX2125) );
  INVX0 U6340_U1 ( .INP(n10659), .ZN(U6340_n1) );
  AND2X1 U6341_U2 ( .IN1(WX2060), .IN2(U6341_n1), .Q(WX2123) );
  INVX0 U6341_U1 ( .INP(n10659), .ZN(U6341_n1) );
  AND2X1 U6342_U2 ( .IN1(WX2058), .IN2(U6342_n1), .Q(WX2121) );
  INVX0 U6342_U1 ( .INP(n10659), .ZN(U6342_n1) );
  AND2X1 U6343_U2 ( .IN1(WX2056), .IN2(U6343_n1), .Q(WX2119) );
  INVX0 U6343_U1 ( .INP(n10659), .ZN(U6343_n1) );
  AND2X1 U6344_U2 ( .IN1(WX2054), .IN2(U6344_n1), .Q(WX2117) );
  INVX0 U6344_U1 ( .INP(n10659), .ZN(U6344_n1) );
  AND2X1 U6345_U2 ( .IN1(WX2052), .IN2(U6345_n1), .Q(WX2115) );
  INVX0 U6345_U1 ( .INP(n10659), .ZN(U6345_n1) );
  AND2X1 U6346_U2 ( .IN1(WX2050), .IN2(U6346_n1), .Q(WX2113) );
  INVX0 U6346_U1 ( .INP(n10659), .ZN(U6346_n1) );
  AND2X1 U6347_U2 ( .IN1(WX2048), .IN2(U6347_n1), .Q(WX2111) );
  INVX0 U6347_U1 ( .INP(n10659), .ZN(U6347_n1) );
  AND2X1 U6348_U2 ( .IN1(WX2046), .IN2(U6348_n1), .Q(WX2109) );
  INVX0 U6348_U1 ( .INP(n10659), .ZN(U6348_n1) );
  AND2X1 U6349_U2 ( .IN1(WX2044), .IN2(U6349_n1), .Q(WX2107) );
  INVX0 U6349_U1 ( .INP(n10659), .ZN(U6349_n1) );
  AND2X1 U6350_U2 ( .IN1(WX2042), .IN2(U6350_n1), .Q(WX2105) );
  INVX0 U6350_U1 ( .INP(n10659), .ZN(U6350_n1) );
  AND2X1 U6351_U2 ( .IN1(WX2040), .IN2(U6351_n1), .Q(WX2103) );
  INVX0 U6351_U1 ( .INP(n10659), .ZN(U6351_n1) );
  AND2X1 U6352_U2 ( .IN1(WX2038), .IN2(U6352_n1), .Q(WX2101) );
  INVX0 U6352_U1 ( .INP(n10659), .ZN(U6352_n1) );
  AND2X1 U6353_U2 ( .IN1(WX2036), .IN2(U6353_n1), .Q(WX2099) );
  INVX0 U6353_U1 ( .INP(n10659), .ZN(U6353_n1) );
  AND2X1 U6354_U2 ( .IN1(WX2034), .IN2(U6354_n1), .Q(WX2097) );
  INVX0 U6354_U1 ( .INP(n10658), .ZN(U6354_n1) );
  AND2X1 U6355_U2 ( .IN1(WX2032), .IN2(U6355_n1), .Q(WX2095) );
  INVX0 U6355_U1 ( .INP(n10658), .ZN(U6355_n1) );
  AND2X1 U6356_U2 ( .IN1(WX2030), .IN2(U6356_n1), .Q(WX2093) );
  INVX0 U6356_U1 ( .INP(n10658), .ZN(U6356_n1) );
  AND2X1 U6357_U2 ( .IN1(test_so15), .IN2(U6357_n1), .Q(WX2091) );
  INVX0 U6357_U1 ( .INP(n10658), .ZN(U6357_n1) );
  AND2X1 U6358_U2 ( .IN1(WX2026), .IN2(U6358_n1), .Q(WX2089) );
  INVX0 U6358_U1 ( .INP(n10658), .ZN(U6358_n1) );
  AND2X1 U6359_U2 ( .IN1(WX2024), .IN2(U6359_n1), .Q(WX2087) );
  INVX0 U6359_U1 ( .INP(n10658), .ZN(U6359_n1) );
  AND2X1 U6360_U2 ( .IN1(WX2022), .IN2(U6360_n1), .Q(WX2085) );
  INVX0 U6360_U1 ( .INP(n10658), .ZN(U6360_n1) );
  AND2X1 U6361_U2 ( .IN1(WX2020), .IN2(U6361_n1), .Q(WX2083) );
  INVX0 U6361_U1 ( .INP(n10658), .ZN(U6361_n1) );
  AND2X1 U6362_U2 ( .IN1(WX2018), .IN2(U6362_n1), .Q(WX2081) );
  INVX0 U6362_U1 ( .INP(n10658), .ZN(U6362_n1) );
  AND2X1 U6363_U2 ( .IN1(WX2016), .IN2(U6363_n1), .Q(WX2079) );
  INVX0 U6363_U1 ( .INP(n10658), .ZN(U6363_n1) );
  AND2X1 U6364_U2 ( .IN1(WX2014), .IN2(U6364_n1), .Q(WX2077) );
  INVX0 U6364_U1 ( .INP(n10658), .ZN(U6364_n1) );
  AND2X1 U6365_U2 ( .IN1(WX2012), .IN2(U6365_n1), .Q(WX2075) );
  INVX0 U6365_U1 ( .INP(n10658), .ZN(U6365_n1) );
  AND2X1 U6366_U2 ( .IN1(WX2010), .IN2(U6366_n1), .Q(WX2073) );
  INVX0 U6366_U1 ( .INP(n10658), .ZN(U6366_n1) );
  AND2X1 U6367_U2 ( .IN1(WX2008), .IN2(U6367_n1), .Q(WX2071) );
  INVX0 U6367_U1 ( .INP(n10658), .ZN(U6367_n1) );
  AND2X1 U6368_U2 ( .IN1(WX2006), .IN2(U6368_n1), .Q(WX2069) );
  INVX0 U6368_U1 ( .INP(n10657), .ZN(U6368_n1) );
  AND2X1 U6369_U2 ( .IN1(WX2004), .IN2(U6369_n1), .Q(WX2067) );
  INVX0 U6369_U1 ( .INP(n10657), .ZN(U6369_n1) );
  AND2X1 U6370_U2 ( .IN1(WX2002), .IN2(U6370_n1), .Q(WX2065) );
  INVX0 U6370_U1 ( .INP(n10657), .ZN(U6370_n1) );
  AND2X1 U6371_U2 ( .IN1(WX2000), .IN2(U6371_n1), .Q(WX2063) );
  INVX0 U6371_U1 ( .INP(n10657), .ZN(U6371_n1) );
  AND2X1 U6372_U2 ( .IN1(WX1998), .IN2(U6372_n1), .Q(WX2061) );
  INVX0 U6372_U1 ( .INP(n10657), .ZN(U6372_n1) );
  AND2X1 U6373_U2 ( .IN1(WX1996), .IN2(U6373_n1), .Q(WX2059) );
  INVX0 U6373_U1 ( .INP(n10657), .ZN(U6373_n1) );
  AND2X1 U6374_U2 ( .IN1(WX1994), .IN2(U6374_n1), .Q(WX2057) );
  INVX0 U6374_U1 ( .INP(n10657), .ZN(U6374_n1) );
  AND2X1 U6375_U2 ( .IN1(test_so14), .IN2(U6375_n1), .Q(WX2055) );
  INVX0 U6375_U1 ( .INP(n10657), .ZN(U6375_n1) );
  AND2X1 U6376_U2 ( .IN1(WX1990), .IN2(U6376_n1), .Q(WX2053) );
  INVX0 U6376_U1 ( .INP(n10657), .ZN(U6376_n1) );
  AND2X1 U6377_U2 ( .IN1(WX1988), .IN2(U6377_n1), .Q(WX2051) );
  INVX0 U6377_U1 ( .INP(n10657), .ZN(U6377_n1) );
  AND2X1 U6378_U2 ( .IN1(WX1986), .IN2(U6378_n1), .Q(WX2049) );
  INVX0 U6378_U1 ( .INP(n10657), .ZN(U6378_n1) );
  AND2X1 U6379_U2 ( .IN1(WX1984), .IN2(U6379_n1), .Q(WX2047) );
  INVX0 U6379_U1 ( .INP(n10657), .ZN(U6379_n1) );
  AND2X1 U6380_U2 ( .IN1(WX1982), .IN2(U6380_n1), .Q(WX2045) );
  INVX0 U6380_U1 ( .INP(n10657), .ZN(U6380_n1) );
  AND2X1 U6381_U2 ( .IN1(WX1980), .IN2(U6381_n1), .Q(WX2043) );
  INVX0 U6381_U1 ( .INP(n10657), .ZN(U6381_n1) );
  AND2X1 U6382_U2 ( .IN1(WX1978), .IN2(U6382_n1), .Q(WX2041) );
  INVX0 U6382_U1 ( .INP(n10656), .ZN(U6382_n1) );
  AND2X1 U6383_U2 ( .IN1(WX1976), .IN2(U6383_n1), .Q(WX2039) );
  INVX0 U6383_U1 ( .INP(n10656), .ZN(U6383_n1) );
  AND2X1 U6384_U2 ( .IN1(WX1974), .IN2(U6384_n1), .Q(WX2037) );
  INVX0 U6384_U1 ( .INP(n10656), .ZN(U6384_n1) );
  AND2X1 U6385_U2 ( .IN1(WX1972), .IN2(U6385_n1), .Q(WX2035) );
  INVX0 U6385_U1 ( .INP(n10656), .ZN(U6385_n1) );
  AND2X1 U6386_U2 ( .IN1(WX1970), .IN2(U6386_n1), .Q(WX2033) );
  INVX0 U6386_U1 ( .INP(n10656), .ZN(U6386_n1) );
  AND2X1 U6387_U2 ( .IN1(WX835), .IN2(U6387_n1), .Q(WX898) );
  INVX0 U6387_U1 ( .INP(n10656), .ZN(U6387_n1) );
  AND2X1 U6388_U2 ( .IN1(WX833), .IN2(U6388_n1), .Q(WX896) );
  INVX0 U6388_U1 ( .INP(n10656), .ZN(U6388_n1) );
  AND2X1 U6389_U2 ( .IN1(test_so7), .IN2(U6389_n1), .Q(WX894) );
  INVX0 U6389_U1 ( .INP(n10656), .ZN(U6389_n1) );
  AND2X1 U6390_U2 ( .IN1(WX829), .IN2(U6390_n1), .Q(WX892) );
  INVX0 U6390_U1 ( .INP(n10656), .ZN(U6390_n1) );
  AND2X1 U6391_U2 ( .IN1(WX827), .IN2(U6391_n1), .Q(WX890) );
  INVX0 U6391_U1 ( .INP(n10656), .ZN(U6391_n1) );
  AND2X1 U6392_U2 ( .IN1(WX825), .IN2(U6392_n1), .Q(WX888) );
  INVX0 U6392_U1 ( .INP(n10656), .ZN(U6392_n1) );
  AND2X1 U6393_U2 ( .IN1(WX823), .IN2(U6393_n1), .Q(WX886) );
  INVX0 U6393_U1 ( .INP(n10656), .ZN(U6393_n1) );
  AND2X1 U6394_U2 ( .IN1(WX821), .IN2(U6394_n1), .Q(WX884) );
  INVX0 U6394_U1 ( .INP(n10656), .ZN(U6394_n1) );
  AND2X1 U6395_U2 ( .IN1(WX819), .IN2(U6395_n1), .Q(WX882) );
  INVX0 U6395_U1 ( .INP(n10656), .ZN(U6395_n1) );
  AND2X1 U6396_U2 ( .IN1(WX817), .IN2(U6396_n1), .Q(WX880) );
  INVX0 U6396_U1 ( .INP(n10655), .ZN(U6396_n1) );
  AND2X1 U6397_U2 ( .IN1(WX815), .IN2(U6397_n1), .Q(WX878) );
  INVX0 U6397_U1 ( .INP(n10655), .ZN(U6397_n1) );
  AND2X1 U6398_U2 ( .IN1(WX813), .IN2(U6398_n1), .Q(WX876) );
  INVX0 U6398_U1 ( .INP(n10655), .ZN(U6398_n1) );
  AND2X1 U6399_U2 ( .IN1(WX811), .IN2(U6399_n1), .Q(WX874) );
  INVX0 U6399_U1 ( .INP(n10655), .ZN(U6399_n1) );
  AND2X1 U6400_U2 ( .IN1(WX809), .IN2(U6400_n1), .Q(WX872) );
  INVX0 U6400_U1 ( .INP(n10655), .ZN(U6400_n1) );
  AND2X1 U6401_U2 ( .IN1(WX807), .IN2(U6401_n1), .Q(WX870) );
  INVX0 U6401_U1 ( .INP(n10655), .ZN(U6401_n1) );
  AND2X1 U6402_U2 ( .IN1(WX805), .IN2(U6402_n1), .Q(WX868) );
  INVX0 U6402_U1 ( .INP(n10655), .ZN(U6402_n1) );
  AND2X1 U6403_U2 ( .IN1(WX803), .IN2(U6403_n1), .Q(WX866) );
  INVX0 U6403_U1 ( .INP(n10655), .ZN(U6403_n1) );
  AND2X1 U6404_U2 ( .IN1(WX801), .IN2(U6404_n1), .Q(WX864) );
  INVX0 U6404_U1 ( .INP(n10655), .ZN(U6404_n1) );
  AND2X1 U6405_U2 ( .IN1(WX799), .IN2(U6405_n1), .Q(WX862) );
  INVX0 U6405_U1 ( .INP(n10655), .ZN(U6405_n1) );
  AND2X1 U6406_U2 ( .IN1(WX797), .IN2(U6406_n1), .Q(WX860) );
  INVX0 U6406_U1 ( .INP(n10655), .ZN(U6406_n1) );
  AND2X1 U6407_U2 ( .IN1(test_so6), .IN2(U6407_n1), .Q(WX858) );
  INVX0 U6407_U1 ( .INP(n10655), .ZN(U6407_n1) );
  AND2X1 U6408_U2 ( .IN1(WX793), .IN2(U6408_n1), .Q(WX856) );
  INVX0 U6408_U1 ( .INP(n10655), .ZN(U6408_n1) );
  AND2X1 U6409_U2 ( .IN1(WX791), .IN2(U6409_n1), .Q(WX854) );
  INVX0 U6409_U1 ( .INP(n10655), .ZN(U6409_n1) );
  AND2X1 U6410_U2 ( .IN1(WX789), .IN2(U6410_n1), .Q(WX852) );
  INVX0 U6410_U1 ( .INP(n10654), .ZN(U6410_n1) );
  AND2X1 U6411_U2 ( .IN1(WX787), .IN2(U6411_n1), .Q(WX850) );
  INVX0 U6411_U1 ( .INP(n10654), .ZN(U6411_n1) );
  AND2X1 U6412_U2 ( .IN1(WX785), .IN2(U6412_n1), .Q(WX848) );
  INVX0 U6412_U1 ( .INP(n10654), .ZN(U6412_n1) );
  AND2X1 U6413_U2 ( .IN1(WX783), .IN2(U6413_n1), .Q(WX846) );
  INVX0 U6413_U1 ( .INP(n10654), .ZN(U6413_n1) );
  AND2X1 U6414_U2 ( .IN1(WX781), .IN2(U6414_n1), .Q(WX844) );
  INVX0 U6414_U1 ( .INP(n10654), .ZN(U6414_n1) );
  AND2X1 U6415_U2 ( .IN1(WX779), .IN2(U6415_n1), .Q(WX842) );
  INVX0 U6415_U1 ( .INP(n10654), .ZN(U6415_n1) );
  AND2X1 U6416_U2 ( .IN1(WX777), .IN2(U6416_n1), .Q(WX840) );
  INVX0 U6416_U1 ( .INP(n10654), .ZN(U6416_n1) );
  AND2X1 U6417_U2 ( .IN1(WX775), .IN2(U6417_n1), .Q(WX838) );
  INVX0 U6417_U1 ( .INP(n10654), .ZN(U6417_n1) );
  AND2X1 U6418_U2 ( .IN1(WX773), .IN2(U6418_n1), .Q(WX836) );
  INVX0 U6418_U1 ( .INP(n10654), .ZN(U6418_n1) );
  AND2X1 U6419_U2 ( .IN1(WX771), .IN2(U6419_n1), .Q(WX834) );
  INVX0 U6419_U1 ( .INP(n10654), .ZN(U6419_n1) );
  AND2X1 U6420_U2 ( .IN1(WX769), .IN2(U6420_n1), .Q(WX832) );
  INVX0 U6420_U1 ( .INP(n10654), .ZN(U6420_n1) );
  AND2X1 U6421_U2 ( .IN1(WX767), .IN2(U6421_n1), .Q(WX830) );
  INVX0 U6421_U1 ( .INP(n10654), .ZN(U6421_n1) );
  AND2X1 U6422_U2 ( .IN1(WX765), .IN2(U6422_n1), .Q(WX828) );
  INVX0 U6422_U1 ( .INP(n10654), .ZN(U6422_n1) );
  AND2X1 U6423_U2 ( .IN1(WX763), .IN2(U6423_n1), .Q(WX826) );
  INVX0 U6423_U1 ( .INP(n10654), .ZN(U6423_n1) );
  AND2X1 U6424_U2 ( .IN1(WX761), .IN2(U6424_n1), .Q(WX824) );
  INVX0 U6424_U1 ( .INP(n10653), .ZN(U6424_n1) );
  AND2X1 U6425_U2 ( .IN1(test_so5), .IN2(U6425_n1), .Q(WX822) );
  INVX0 U6425_U1 ( .INP(n10653), .ZN(U6425_n1) );
  AND2X1 U6426_U2 ( .IN1(WX757), .IN2(U6426_n1), .Q(WX820) );
  INVX0 U6426_U1 ( .INP(n10653), .ZN(U6426_n1) );
  AND2X1 U6427_U2 ( .IN1(WX755), .IN2(U6427_n1), .Q(WX818) );
  INVX0 U6427_U1 ( .INP(n10653), .ZN(U6427_n1) );
  AND2X1 U6428_U2 ( .IN1(WX753), .IN2(U6428_n1), .Q(WX816) );
  INVX0 U6428_U1 ( .INP(n10653), .ZN(U6428_n1) );
  AND2X1 U6429_U2 ( .IN1(WX751), .IN2(U6429_n1), .Q(WX814) );
  INVX0 U6429_U1 ( .INP(n10653), .ZN(U6429_n1) );
  AND2X1 U6430_U2 ( .IN1(WX749), .IN2(U6430_n1), .Q(WX812) );
  INVX0 U6430_U1 ( .INP(n10653), .ZN(U6430_n1) );
  AND2X1 U6431_U2 ( .IN1(WX747), .IN2(U6431_n1), .Q(WX810) );
  INVX0 U6431_U1 ( .INP(n10653), .ZN(U6431_n1) );
  AND2X1 U6432_U2 ( .IN1(WX745), .IN2(U6432_n1), .Q(WX808) );
  INVX0 U6432_U1 ( .INP(n10653), .ZN(U6432_n1) );
  AND2X1 U6433_U2 ( .IN1(WX743), .IN2(U6433_n1), .Q(WX806) );
  INVX0 U6433_U1 ( .INP(n10653), .ZN(U6433_n1) );
  AND2X1 U6434_U2 ( .IN1(WX741), .IN2(U6434_n1), .Q(WX804) );
  INVX0 U6434_U1 ( .INP(n10653), .ZN(U6434_n1) );
  AND2X1 U6435_U2 ( .IN1(WX739), .IN2(U6435_n1), .Q(WX802) );
  INVX0 U6435_U1 ( .INP(n10653), .ZN(U6435_n1) );
  AND2X1 U6436_U2 ( .IN1(WX737), .IN2(U6436_n1), .Q(WX800) );
  INVX0 U6436_U1 ( .INP(n10653), .ZN(U6436_n1) );
  AND2X1 U6437_U2 ( .IN1(WX735), .IN2(U6437_n1), .Q(WX798) );
  INVX0 U6437_U1 ( .INP(n10653), .ZN(U6437_n1) );
  AND2X1 U6438_U2 ( .IN1(WX733), .IN2(U6438_n1), .Q(WX796) );
  INVX0 U6438_U1 ( .INP(n10652), .ZN(U6438_n1) );
  AND2X1 U6439_U2 ( .IN1(WX731), .IN2(U6439_n1), .Q(WX794) );
  INVX0 U6439_U1 ( .INP(n10652), .ZN(U6439_n1) );
  AND2X1 U6440_U2 ( .IN1(WX729), .IN2(U6440_n1), .Q(WX792) );
  INVX0 U6440_U1 ( .INP(n10652), .ZN(U6440_n1) );
  AND2X1 U6441_U2 ( .IN1(WX727), .IN2(U6441_n1), .Q(WX790) );
  INVX0 U6441_U1 ( .INP(n10652), .ZN(U6441_n1) );
  AND2X1 U6442_U2 ( .IN1(WX725), .IN2(U6442_n1), .Q(WX788) );
  INVX0 U6442_U1 ( .INP(n10652), .ZN(U6442_n1) );
  AND2X1 U6443_U2 ( .IN1(test_so4), .IN2(U6443_n1), .Q(WX786) );
  INVX0 U6443_U1 ( .INP(n10652), .ZN(U6443_n1) );
  AND2X1 U6444_U2 ( .IN1(WX721), .IN2(U6444_n1), .Q(WX784) );
  INVX0 U6444_U1 ( .INP(n10652), .ZN(U6444_n1) );
  AND2X1 U6445_U2 ( .IN1(WX719), .IN2(U6445_n1), .Q(WX782) );
  INVX0 U6445_U1 ( .INP(n10652), .ZN(U6445_n1) );
  AND2X1 U6446_U2 ( .IN1(WX717), .IN2(U6446_n1), .Q(WX780) );
  INVX0 U6446_U1 ( .INP(n10652), .ZN(U6446_n1) );
  AND2X1 U6447_U2 ( .IN1(WX715), .IN2(U6447_n1), .Q(WX778) );
  INVX0 U6447_U1 ( .INP(n10652), .ZN(U6447_n1) );
  AND2X1 U6448_U2 ( .IN1(WX713), .IN2(U6448_n1), .Q(WX776) );
  INVX0 U6448_U1 ( .INP(n10652), .ZN(U6448_n1) );
  AND2X1 U6449_U2 ( .IN1(WX711), .IN2(U6449_n1), .Q(WX774) );
  INVX0 U6449_U1 ( .INP(n10652), .ZN(U6449_n1) );
  AND2X1 U6450_U2 ( .IN1(WX709), .IN2(U6450_n1), .Q(WX772) );
  INVX0 U6450_U1 ( .INP(n10652), .ZN(U6450_n1) );
  AND2X1 U6451_U2 ( .IN1(WX707), .IN2(U6451_n1), .Q(WX770) );
  INVX0 U6451_U1 ( .INP(n10652), .ZN(U6451_n1) );
  AND2X1 U6452_U2 ( .IN1(WX705), .IN2(U6452_n1), .Q(WX768) );
  INVX0 U6452_U1 ( .INP(n10651), .ZN(U6452_n1) );
  AND2X1 U6453_U2 ( .IN1(WX703), .IN2(U6453_n1), .Q(WX766) );
  INVX0 U6453_U1 ( .INP(n10651), .ZN(U6453_n1) );
  AND2X1 U6454_U2 ( .IN1(WX701), .IN2(U6454_n1), .Q(WX764) );
  INVX0 U6454_U1 ( .INP(n10651), .ZN(U6454_n1) );
  AND2X1 U6455_U2 ( .IN1(WX699), .IN2(U6455_n1), .Q(WX762) );
  INVX0 U6455_U1 ( .INP(n10651), .ZN(U6455_n1) );
  AND2X1 U6456_U2 ( .IN1(WX697), .IN2(U6456_n1), .Q(WX760) );
  INVX0 U6456_U1 ( .INP(n10651), .ZN(U6456_n1) );
  AND2X1 U6457_U2 ( .IN1(WX695), .IN2(U6457_n1), .Q(WX758) );
  INVX0 U6457_U1 ( .INP(n10651), .ZN(U6457_n1) );
  AND2X1 U6458_U2 ( .IN1(WX693), .IN2(U6458_n1), .Q(WX756) );
  INVX0 U6458_U1 ( .INP(n10651), .ZN(U6458_n1) );
  AND2X1 U6459_U2 ( .IN1(WX691), .IN2(U6459_n1), .Q(WX754) );
  INVX0 U6459_U1 ( .INP(n10651), .ZN(U6459_n1) );
  AND2X1 U6460_U2 ( .IN1(WX689), .IN2(U6460_n1), .Q(WX752) );
  INVX0 U6460_U1 ( .INP(n10651), .ZN(U6460_n1) );
  AND2X1 U6461_U2 ( .IN1(test_so3), .IN2(U6461_n1), .Q(WX750) );
  INVX0 U6461_U1 ( .INP(n10651), .ZN(U6461_n1) );
  AND2X1 U6462_U2 ( .IN1(WX685), .IN2(U6462_n1), .Q(WX748) );
  INVX0 U6462_U1 ( .INP(n10651), .ZN(U6462_n1) );
  AND2X1 U6463_U2 ( .IN1(WX683), .IN2(U6463_n1), .Q(WX746) );
  INVX0 U6463_U1 ( .INP(n10651), .ZN(U6463_n1) );
  AND2X1 U6464_U2 ( .IN1(WX681), .IN2(U6464_n1), .Q(WX744) );
  INVX0 U6464_U1 ( .INP(n10651), .ZN(U6464_n1) );
  AND2X1 U6465_U2 ( .IN1(WX679), .IN2(U6465_n1), .Q(WX742) );
  INVX0 U6465_U1 ( .INP(n10651), .ZN(U6465_n1) );
  AND2X1 U6466_U2 ( .IN1(WX677), .IN2(U6466_n1), .Q(WX740) );
  INVX0 U6466_U1 ( .INP(n10650), .ZN(U6466_n1) );
  AND2X1 U6467_U2 ( .IN1(WX675), .IN2(U6467_n1), .Q(WX738) );
  INVX0 U6467_U1 ( .INP(n10650), .ZN(U6467_n1) );
  AND2X1 U6468_U2 ( .IN1(WX673), .IN2(U6468_n1), .Q(WX736) );
  INVX0 U6468_U1 ( .INP(n10650), .ZN(U6468_n1) );
  AND2X1 U6469_U2 ( .IN1(WX671), .IN2(U6469_n1), .Q(WX734) );
  INVX0 U6469_U1 ( .INP(n10650), .ZN(U6469_n1) );
  AND2X1 U6470_U2 ( .IN1(WX669), .IN2(U6470_n1), .Q(WX732) );
  INVX0 U6470_U1 ( .INP(n10650), .ZN(U6470_n1) );
  AND2X1 U6471_U2 ( .IN1(WX667), .IN2(U6471_n1), .Q(WX730) );
  INVX0 U6471_U1 ( .INP(n10650), .ZN(U6471_n1) );
  AND2X1 U6472_U2 ( .IN1(WX665), .IN2(U6472_n1), .Q(WX728) );
  INVX0 U6472_U1 ( .INP(n10650), .ZN(U6472_n1) );
  AND2X1 U6473_U2 ( .IN1(WX663), .IN2(U6473_n1), .Q(WX726) );
  INVX0 U6473_U1 ( .INP(n10650), .ZN(U6473_n1) );
  AND2X1 U6474_U2 ( .IN1(WX661), .IN2(U6474_n1), .Q(WX724) );
  INVX0 U6474_U1 ( .INP(n10650), .ZN(U6474_n1) );
  AND2X1 U6475_U2 ( .IN1(WX659), .IN2(U6475_n1), .Q(WX722) );
  INVX0 U6475_U1 ( .INP(n10650), .ZN(U6475_n1) );
  AND2X1 U6476_U2 ( .IN1(WX657), .IN2(U6476_n1), .Q(WX720) );
  INVX0 U6476_U1 ( .INP(n10650), .ZN(U6476_n1) );
  AND2X1 U6477_U2 ( .IN1(WX655), .IN2(U6477_n1), .Q(WX718) );
  INVX0 U6477_U1 ( .INP(n10650), .ZN(U6477_n1) );
  AND2X1 U6478_U2 ( .IN1(WX653), .IN2(U6478_n1), .Q(WX716) );
  INVX0 U6478_U1 ( .INP(n10650), .ZN(U6478_n1) );
  AND2X1 U6479_U2 ( .IN1(test_so2), .IN2(U6479_n1), .Q(WX714) );
  INVX0 U6479_U1 ( .INP(n10650), .ZN(U6479_n1) );
  AND2X1 U6480_U2 ( .IN1(WX649), .IN2(U6480_n1), .Q(WX712) );
  INVX0 U6480_U1 ( .INP(n10649), .ZN(U6480_n1) );
  AND2X1 U6481_U2 ( .IN1(WX647), .IN2(U6481_n1), .Q(WX710) );
  INVX0 U6481_U1 ( .INP(n10649), .ZN(U6481_n1) );
  AND2X1 U6482_U2 ( .IN1(WX645), .IN2(U6482_n1), .Q(WX708) );
  INVX0 U6482_U1 ( .INP(n10649), .ZN(U6482_n1) );
endmodule

