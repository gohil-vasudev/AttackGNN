module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n170_, new_n246_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n792_, new_n1058_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n806_, new_n1016_, new_n605_, new_n1074_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n927_, new_n196_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n865_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n138_, keyIn_0_41 );
not g001 ( new_n139_, N81 );
not g002 ( new_n140_, N85 );
and g003 ( new_n141_, new_n139_, new_n140_ );
and g004 ( new_n142_, N81, N85 );
or g005 ( new_n143_, new_n141_, new_n142_ );
not g006 ( new_n144_, N89 );
not g007 ( new_n145_, N93 );
and g008 ( new_n146_, new_n144_, new_n145_ );
and g009 ( new_n147_, N89, N93 );
or g010 ( new_n148_, new_n146_, new_n147_ );
and g011 ( new_n149_, new_n143_, new_n148_ );
not g012 ( new_n150_, new_n149_ );
or g013 ( new_n151_, new_n143_, new_n148_ );
and g014 ( new_n152_, new_n150_, new_n151_ );
not g015 ( new_n153_, N73 );
not g016 ( new_n154_, N77 );
and g017 ( new_n155_, new_n153_, new_n154_ );
and g018 ( new_n156_, N73, N77 );
or g019 ( new_n157_, new_n155_, new_n156_ );
not g020 ( new_n158_, new_n157_ );
not g021 ( new_n159_, keyIn_0_5 );
not g022 ( new_n160_, N65 );
not g023 ( new_n161_, N69 );
and g024 ( new_n162_, new_n160_, new_n161_ );
not g025 ( new_n163_, new_n162_ );
and g026 ( new_n164_, N65, N69 );
not g027 ( new_n165_, new_n164_ );
and g028 ( new_n166_, new_n163_, new_n165_ );
or g029 ( new_n167_, new_n166_, new_n159_ );
and g030 ( new_n168_, new_n163_, new_n159_ );
and g031 ( new_n169_, new_n168_, new_n165_ );
not g032 ( new_n170_, new_n169_ );
and g033 ( new_n171_, new_n170_, new_n167_ );
not g034 ( new_n172_, new_n171_ );
and g035 ( new_n173_, new_n172_, keyIn_0_6 );
not g036 ( new_n174_, new_n173_ );
or g037 ( new_n175_, new_n172_, keyIn_0_6 );
and g038 ( new_n176_, new_n174_, new_n175_ );
and g039 ( new_n177_, new_n176_, new_n158_ );
not g040 ( new_n178_, new_n177_ );
or g041 ( new_n179_, new_n176_, new_n158_ );
and g042 ( new_n180_, new_n178_, new_n179_ );
not g043 ( new_n181_, new_n180_ );
and g044 ( new_n182_, new_n181_, new_n152_ );
not g045 ( new_n183_, new_n152_ );
and g046 ( new_n184_, new_n180_, new_n183_ );
or g047 ( new_n185_, new_n182_, new_n184_ );
and g048 ( new_n186_, N129, N137 );
not g049 ( new_n187_, new_n186_ );
and g050 ( new_n188_, new_n185_, new_n187_ );
not g051 ( new_n189_, new_n188_ );
or g052 ( new_n190_, new_n185_, new_n187_ );
and g053 ( new_n191_, new_n189_, new_n190_ );
not g054 ( new_n192_, N17 );
and g055 ( new_n193_, new_n192_, N1 );
not g056 ( new_n194_, N1 );
and g057 ( new_n195_, new_n194_, N17 );
or g058 ( new_n196_, new_n193_, new_n195_ );
not g059 ( new_n197_, N33 );
not g060 ( new_n198_, N49 );
and g061 ( new_n199_, new_n197_, new_n198_ );
and g062 ( new_n200_, N33, N49 );
or g063 ( new_n201_, new_n199_, new_n200_ );
and g064 ( new_n202_, new_n196_, new_n201_ );
not g065 ( new_n203_, new_n202_ );
or g066 ( new_n204_, new_n196_, new_n201_ );
and g067 ( new_n205_, new_n203_, new_n204_ );
not g068 ( new_n206_, new_n205_ );
and g069 ( new_n207_, new_n191_, new_n206_ );
not g070 ( new_n208_, new_n207_ );
or g071 ( new_n209_, new_n191_, new_n206_ );
and g072 ( new_n210_, new_n208_, new_n209_ );
not g073 ( new_n211_, new_n210_ );
not g074 ( new_n212_, keyIn_0_8 );
not g075 ( new_n213_, N101 );
and g076 ( new_n214_, new_n213_, N97 );
not g077 ( new_n215_, N97 );
and g078 ( new_n216_, new_n215_, N101 );
or g079 ( new_n217_, new_n214_, new_n216_ );
not g080 ( new_n218_, N105 );
not g081 ( new_n219_, N109 );
and g082 ( new_n220_, new_n218_, new_n219_ );
and g083 ( new_n221_, N105, N109 );
or g084 ( new_n222_, new_n220_, new_n221_ );
and g085 ( new_n223_, new_n217_, new_n222_ );
not g086 ( new_n224_, new_n223_ );
or g087 ( new_n225_, new_n217_, new_n222_ );
and g088 ( new_n226_, new_n224_, new_n225_ );
not g089 ( new_n227_, new_n226_ );
and g090 ( new_n228_, new_n227_, keyIn_0_18 );
not g091 ( new_n229_, new_n228_ );
or g092 ( new_n230_, new_n227_, keyIn_0_18 );
and g093 ( new_n231_, new_n229_, new_n230_ );
not g094 ( new_n232_, new_n231_ );
not g095 ( new_n233_, keyIn_0_19 );
not g096 ( new_n234_, keyIn_0_7 );
not g097 ( new_n235_, N121 );
not g098 ( new_n236_, N125 );
and g099 ( new_n237_, new_n235_, new_n236_ );
not g100 ( new_n238_, new_n237_ );
and g101 ( new_n239_, N121, N125 );
not g102 ( new_n240_, new_n239_ );
and g103 ( new_n241_, new_n238_, new_n240_ );
or g104 ( new_n242_, new_n241_, new_n234_ );
and g105 ( new_n243_, new_n238_, new_n234_ );
and g106 ( new_n244_, new_n243_, new_n240_ );
not g107 ( new_n245_, new_n244_ );
and g108 ( new_n246_, new_n245_, new_n242_ );
not g109 ( new_n247_, new_n246_ );
not g110 ( new_n248_, N117 );
and g111 ( new_n249_, new_n248_, N113 );
not g112 ( new_n250_, N113 );
and g113 ( new_n251_, new_n250_, N117 );
or g114 ( new_n252_, new_n249_, new_n251_ );
and g115 ( new_n253_, new_n247_, new_n252_ );
not g116 ( new_n254_, new_n253_ );
or g117 ( new_n255_, new_n247_, new_n252_ );
and g118 ( new_n256_, new_n254_, new_n255_ );
or g119 ( new_n257_, new_n256_, new_n233_ );
and g120 ( new_n258_, new_n256_, new_n233_ );
not g121 ( new_n259_, new_n258_ );
and g122 ( new_n260_, new_n259_, new_n257_ );
not g123 ( new_n261_, new_n260_ );
and g124 ( new_n262_, new_n261_, new_n232_ );
and g125 ( new_n263_, new_n260_, new_n231_ );
or g126 ( new_n264_, new_n262_, new_n263_ );
and g127 ( new_n265_, new_n264_, keyIn_0_22 );
not g128 ( new_n266_, new_n265_ );
or g129 ( new_n267_, new_n264_, keyIn_0_22 );
and g130 ( new_n268_, new_n266_, new_n267_ );
or g131 ( new_n269_, new_n268_, new_n212_ );
and g132 ( new_n270_, new_n268_, new_n212_ );
not g133 ( new_n271_, new_n270_ );
and g134 ( new_n272_, new_n271_, new_n269_ );
and g135 ( new_n273_, N130, N137 );
or g136 ( new_n274_, new_n272_, new_n273_ );
and g137 ( new_n275_, new_n272_, new_n273_ );
not g138 ( new_n276_, new_n275_ );
and g139 ( new_n277_, new_n276_, new_n274_ );
not g140 ( new_n278_, N21 );
and g141 ( new_n279_, new_n278_, N5 );
not g142 ( new_n280_, N5 );
and g143 ( new_n281_, new_n280_, N21 );
or g144 ( new_n282_, new_n279_, new_n281_ );
and g145 ( new_n283_, new_n282_, keyIn_0_12 );
not g146 ( new_n284_, new_n283_ );
or g147 ( new_n285_, new_n282_, keyIn_0_12 );
and g148 ( new_n286_, new_n284_, new_n285_ );
not g149 ( new_n287_, new_n286_ );
not g150 ( new_n288_, N53 );
and g151 ( new_n289_, new_n288_, N37 );
not g152 ( new_n290_, N37 );
and g153 ( new_n291_, new_n290_, N53 );
or g154 ( new_n292_, new_n289_, new_n291_ );
and g155 ( new_n293_, new_n292_, keyIn_0_13 );
not g156 ( new_n294_, new_n293_ );
or g157 ( new_n295_, new_n292_, keyIn_0_13 );
and g158 ( new_n296_, new_n294_, new_n295_ );
not g159 ( new_n297_, new_n296_ );
and g160 ( new_n298_, new_n287_, new_n297_ );
and g161 ( new_n299_, new_n286_, new_n296_ );
or g162 ( new_n300_, new_n298_, new_n299_ );
not g163 ( new_n301_, new_n300_ );
or g164 ( new_n302_, new_n277_, new_n301_ );
not g165 ( new_n303_, new_n272_ );
not g166 ( new_n304_, new_n273_ );
and g167 ( new_n305_, new_n303_, new_n304_ );
or g168 ( new_n306_, new_n305_, new_n275_ );
or g169 ( new_n307_, new_n306_, new_n300_ );
and g170 ( new_n308_, new_n307_, new_n302_ );
not g171 ( new_n309_, keyIn_0_24 );
and g172 ( new_n310_, new_n181_, new_n231_ );
and g173 ( new_n311_, new_n180_, new_n232_ );
or g174 ( new_n312_, new_n310_, new_n311_ );
and g175 ( new_n313_, N131, N137 );
not g176 ( new_n314_, new_n313_ );
and g177 ( new_n315_, new_n312_, new_n314_ );
not g178 ( new_n316_, new_n315_ );
or g179 ( new_n317_, new_n312_, new_n314_ );
and g180 ( new_n318_, new_n316_, new_n317_ );
not g181 ( new_n319_, N9 );
not g182 ( new_n320_, N25 );
and g183 ( new_n321_, new_n319_, new_n320_ );
and g184 ( new_n322_, N9, N25 );
or g185 ( new_n323_, new_n321_, new_n322_ );
not g186 ( new_n324_, N41 );
not g187 ( new_n325_, N57 );
and g188 ( new_n326_, new_n324_, new_n325_ );
and g189 ( new_n327_, N41, N57 );
or g190 ( new_n328_, new_n326_, new_n327_ );
and g191 ( new_n329_, new_n323_, new_n328_ );
not g192 ( new_n330_, new_n329_ );
or g193 ( new_n331_, new_n323_, new_n328_ );
and g194 ( new_n332_, new_n330_, new_n331_ );
or g195 ( new_n333_, new_n318_, new_n332_ );
and g196 ( new_n334_, new_n318_, new_n332_ );
not g197 ( new_n335_, new_n334_ );
and g198 ( new_n336_, new_n335_, new_n333_ );
or g199 ( new_n337_, new_n336_, new_n309_ );
not g200 ( new_n338_, new_n337_ );
and g201 ( new_n339_, new_n336_, new_n309_ );
or g202 ( new_n340_, new_n338_, new_n339_ );
and g203 ( new_n341_, new_n340_, new_n210_ );
and g204 ( new_n342_, new_n261_, new_n183_ );
and g205 ( new_n343_, new_n260_, new_n152_ );
or g206 ( new_n344_, new_n342_, new_n343_ );
and g207 ( new_n345_, N132, N137 );
or g208 ( new_n346_, new_n345_, keyIn_0_9 );
and g209 ( new_n347_, keyIn_0_9, N132 );
and g210 ( new_n348_, new_n347_, N137 );
not g211 ( new_n349_, new_n348_ );
and g212 ( new_n350_, new_n349_, new_n346_ );
not g213 ( new_n351_, new_n350_ );
and g214 ( new_n352_, new_n344_, new_n351_ );
not g215 ( new_n353_, new_n352_ );
or g216 ( new_n354_, new_n344_, new_n351_ );
and g217 ( new_n355_, new_n353_, new_n354_ );
or g218 ( new_n356_, new_n355_, keyIn_0_23 );
and g219 ( new_n357_, new_n355_, keyIn_0_23 );
not g220 ( new_n358_, new_n357_ );
and g221 ( new_n359_, new_n358_, new_n356_ );
not g222 ( new_n360_, new_n359_ );
not g223 ( new_n361_, N29 );
and g224 ( new_n362_, new_n361_, N13 );
not g225 ( new_n363_, N13 );
and g226 ( new_n364_, new_n363_, N29 );
or g227 ( new_n365_, new_n362_, new_n364_ );
and g228 ( new_n366_, new_n365_, keyIn_0_14 );
not g229 ( new_n367_, new_n366_ );
or g230 ( new_n368_, new_n365_, keyIn_0_14 );
and g231 ( new_n369_, new_n367_, new_n368_ );
not g232 ( new_n370_, new_n369_ );
not g233 ( new_n371_, N61 );
and g234 ( new_n372_, new_n371_, N45 );
not g235 ( new_n373_, N45 );
and g236 ( new_n374_, new_n373_, N61 );
or g237 ( new_n375_, new_n372_, new_n374_ );
and g238 ( new_n376_, new_n370_, new_n375_ );
not g239 ( new_n377_, new_n376_ );
or g240 ( new_n378_, new_n370_, new_n375_ );
and g241 ( new_n379_, new_n377_, new_n378_ );
not g242 ( new_n380_, new_n379_ );
and g243 ( new_n381_, new_n360_, new_n380_ );
and g244 ( new_n382_, new_n359_, new_n379_ );
or g245 ( new_n383_, new_n381_, new_n382_ );
and g246 ( new_n384_, new_n341_, new_n383_ );
and g247 ( new_n385_, new_n308_, new_n384_ );
and g248 ( new_n386_, new_n306_, new_n300_ );
and g249 ( new_n387_, new_n277_, new_n301_ );
or g250 ( new_n388_, new_n386_, new_n387_ );
or g251 ( new_n389_, new_n388_, new_n210_ );
and g252 ( new_n390_, new_n340_, keyIn_0_26 );
not g253 ( new_n391_, keyIn_0_26 );
not g254 ( new_n392_, new_n339_ );
and g255 ( new_n393_, new_n392_, new_n337_ );
and g256 ( new_n394_, new_n393_, new_n391_ );
or g257 ( new_n395_, new_n394_, new_n383_ );
or g258 ( new_n396_, new_n395_, new_n390_ );
or g259 ( new_n397_, new_n389_, new_n396_ );
and g260 ( new_n398_, new_n397_, keyIn_0_36 );
or g261 ( new_n399_, new_n398_, new_n385_ );
not g262 ( new_n400_, new_n383_ );
and g263 ( new_n401_, new_n210_, keyIn_0_25 );
not g264 ( new_n402_, new_n401_ );
or g265 ( new_n403_, new_n210_, keyIn_0_25 );
and g266 ( new_n404_, new_n402_, new_n403_ );
and g267 ( new_n405_, new_n404_, new_n393_ );
and g268 ( new_n406_, new_n308_, new_n405_ );
and g269 ( new_n407_, new_n388_, new_n341_ );
or g270 ( new_n408_, new_n407_, new_n406_ );
and g271 ( new_n409_, new_n408_, new_n400_ );
not g272 ( new_n410_, keyIn_0_36 );
and g273 ( new_n411_, new_n308_, new_n211_ );
not g274 ( new_n412_, new_n390_ );
or g275 ( new_n413_, new_n340_, keyIn_0_26 );
and g276 ( new_n414_, new_n413_, new_n400_ );
and g277 ( new_n415_, new_n414_, new_n412_ );
and g278 ( new_n416_, new_n415_, new_n411_ );
and g279 ( new_n417_, new_n416_, new_n410_ );
or g280 ( new_n418_, new_n409_, new_n417_ );
or g281 ( new_n419_, new_n399_, new_n418_ );
and g282 ( new_n420_, new_n419_, new_n211_ );
not g283 ( new_n421_, keyIn_0_21 );
not g284 ( new_n422_, keyIn_0_3 );
and g285 ( new_n423_, new_n324_, new_n373_ );
and g286 ( new_n424_, N41, N45 );
or g287 ( new_n425_, new_n423_, new_n424_ );
and g288 ( new_n426_, new_n425_, new_n422_ );
not g289 ( new_n427_, new_n424_ );
or g290 ( new_n428_, N41, N45 );
and g291 ( new_n429_, new_n428_, keyIn_0_3 );
and g292 ( new_n430_, new_n429_, new_n427_ );
or g293 ( new_n431_, new_n426_, new_n430_ );
and g294 ( new_n432_, new_n197_, keyIn_0_2 );
not g295 ( new_n433_, keyIn_0_2 );
and g296 ( new_n434_, new_n433_, N33 );
or g297 ( new_n435_, new_n432_, new_n434_ );
and g298 ( new_n436_, new_n435_, new_n290_ );
or g299 ( new_n437_, new_n433_, N33 );
or g300 ( new_n438_, new_n197_, keyIn_0_2 );
and g301 ( new_n439_, new_n437_, new_n438_ );
and g302 ( new_n440_, new_n439_, N37 );
or g303 ( new_n441_, new_n436_, new_n440_ );
and g304 ( new_n442_, new_n441_, new_n431_ );
and g305 ( new_n443_, new_n427_, new_n428_ );
or g306 ( new_n444_, new_n443_, keyIn_0_3 );
not g307 ( new_n445_, new_n430_ );
and g308 ( new_n446_, new_n445_, new_n444_ );
or g309 ( new_n447_, new_n439_, N37 );
or g310 ( new_n448_, new_n435_, new_n290_ );
and g311 ( new_n449_, new_n448_, new_n447_ );
and g312 ( new_n450_, new_n449_, new_n446_ );
or g313 ( new_n451_, new_n442_, new_n450_ );
and g314 ( new_n452_, new_n451_, keyIn_0_17 );
not g315 ( new_n453_, keyIn_0_17 );
or g316 ( new_n454_, new_n449_, new_n446_ );
or g317 ( new_n455_, new_n441_, new_n431_ );
and g318 ( new_n456_, new_n455_, new_n454_ );
and g319 ( new_n457_, new_n456_, new_n453_ );
or g320 ( new_n458_, new_n452_, new_n457_ );
and g321 ( new_n459_, new_n280_, N1 );
and g322 ( new_n460_, new_n194_, N5 );
or g323 ( new_n461_, new_n459_, new_n460_ );
and g324 ( new_n462_, new_n319_, new_n363_ );
and g325 ( new_n463_, N9, N13 );
or g326 ( new_n464_, new_n462_, new_n463_ );
and g327 ( new_n465_, new_n461_, new_n464_ );
not g328 ( new_n466_, new_n465_ );
or g329 ( new_n467_, new_n461_, new_n464_ );
and g330 ( new_n468_, new_n466_, new_n467_ );
not g331 ( new_n469_, new_n468_ );
and g332 ( new_n470_, new_n469_, keyIn_0_16 );
not g333 ( new_n471_, new_n470_ );
or g334 ( new_n472_, new_n469_, keyIn_0_16 );
and g335 ( new_n473_, new_n471_, new_n472_ );
and g336 ( new_n474_, new_n458_, new_n473_ );
or g337 ( new_n475_, new_n456_, new_n453_ );
or g338 ( new_n476_, new_n451_, keyIn_0_17 );
and g339 ( new_n477_, new_n476_, new_n475_ );
not g340 ( new_n478_, new_n473_ );
and g341 ( new_n479_, new_n477_, new_n478_ );
or g342 ( new_n480_, new_n474_, new_n479_ );
and g343 ( new_n481_, new_n480_, new_n421_ );
or g344 ( new_n482_, new_n477_, new_n478_ );
or g345 ( new_n483_, new_n458_, new_n473_ );
and g346 ( new_n484_, new_n483_, new_n482_ );
and g347 ( new_n485_, new_n484_, keyIn_0_21 );
or g348 ( new_n486_, new_n481_, new_n485_ );
and g349 ( new_n487_, new_n486_, keyIn_0_10 );
not g350 ( new_n488_, keyIn_0_10 );
or g351 ( new_n489_, new_n484_, keyIn_0_21 );
or g352 ( new_n490_, new_n480_, new_n421_ );
and g353 ( new_n491_, new_n490_, new_n489_ );
and g354 ( new_n492_, new_n491_, new_n488_ );
or g355 ( new_n493_, new_n487_, new_n492_ );
and g356 ( new_n494_, N135, N137 );
not g357 ( new_n495_, new_n494_ );
and g358 ( new_n496_, new_n493_, new_n495_ );
or g359 ( new_n497_, new_n491_, new_n488_ );
or g360 ( new_n498_, new_n486_, keyIn_0_10 );
and g361 ( new_n499_, new_n498_, new_n497_ );
and g362 ( new_n500_, new_n499_, new_n494_ );
or g363 ( new_n501_, new_n496_, new_n500_ );
not g364 ( new_n502_, keyIn_0_20 );
and g365 ( new_n503_, new_n144_, N73 );
and g366 ( new_n504_, new_n153_, N89 );
or g367 ( new_n505_, new_n503_, new_n504_ );
and g368 ( new_n506_, new_n218_, new_n235_ );
and g369 ( new_n507_, N105, N121 );
or g370 ( new_n508_, new_n506_, new_n507_ );
and g371 ( new_n509_, new_n505_, new_n508_ );
not g372 ( new_n510_, new_n509_ );
or g373 ( new_n511_, new_n505_, new_n508_ );
and g374 ( new_n512_, new_n510_, new_n511_ );
not g375 ( new_n513_, new_n512_ );
and g376 ( new_n514_, new_n513_, new_n502_ );
and g377 ( new_n515_, new_n512_, keyIn_0_20 );
or g378 ( new_n516_, new_n514_, new_n515_ );
and g379 ( new_n517_, new_n501_, new_n516_ );
or g380 ( new_n518_, new_n499_, new_n494_ );
or g381 ( new_n519_, new_n493_, new_n495_ );
and g382 ( new_n520_, new_n519_, new_n518_ );
not g383 ( new_n521_, new_n516_ );
and g384 ( new_n522_, new_n520_, new_n521_ );
or g385 ( new_n523_, new_n517_, new_n522_ );
not g386 ( new_n524_, keyIn_0_4 );
or g387 ( new_n525_, N49, N53 );
and g388 ( new_n526_, N49, N53 );
not g389 ( new_n527_, new_n526_ );
and g390 ( new_n528_, new_n527_, new_n525_ );
or g391 ( new_n529_, new_n528_, new_n524_ );
and g392 ( new_n530_, new_n525_, new_n524_ );
and g393 ( new_n531_, new_n530_, new_n527_ );
not g394 ( new_n532_, new_n531_ );
and g395 ( new_n533_, new_n532_, new_n529_ );
and g396 ( new_n534_, new_n325_, new_n371_ );
and g397 ( new_n535_, N57, N61 );
or g398 ( new_n536_, new_n534_, new_n535_ );
not g399 ( new_n537_, new_n536_ );
or g400 ( new_n538_, new_n533_, new_n537_ );
and g401 ( new_n539_, new_n533_, new_n537_ );
not g402 ( new_n540_, new_n539_ );
and g403 ( new_n541_, new_n540_, new_n538_ );
not g404 ( new_n542_, new_n541_ );
and g405 ( new_n543_, new_n458_, new_n542_ );
and g406 ( new_n544_, new_n477_, new_n541_ );
or g407 ( new_n545_, new_n543_, new_n544_ );
and g408 ( new_n546_, N134, N137 );
not g409 ( new_n547_, new_n546_ );
and g410 ( new_n548_, new_n545_, new_n547_ );
not g411 ( new_n549_, new_n548_ );
or g412 ( new_n550_, new_n545_, new_n547_ );
and g413 ( new_n551_, new_n549_, new_n550_ );
not g414 ( new_n552_, new_n551_ );
and g415 ( new_n553_, new_n161_, new_n140_ );
and g416 ( new_n554_, N69, N85 );
or g417 ( new_n555_, new_n553_, new_n554_ );
and g418 ( new_n556_, new_n213_, new_n248_ );
and g419 ( new_n557_, N101, N117 );
or g420 ( new_n558_, new_n556_, new_n557_ );
and g421 ( new_n559_, new_n555_, new_n558_ );
not g422 ( new_n560_, new_n559_ );
or g423 ( new_n561_, new_n555_, new_n558_ );
and g424 ( new_n562_, new_n560_, new_n561_ );
not g425 ( new_n563_, new_n562_ );
and g426 ( new_n564_, new_n552_, new_n563_ );
and g427 ( new_n565_, new_n551_, new_n562_ );
or g428 ( new_n566_, new_n564_, new_n565_ );
not g429 ( new_n567_, new_n566_ );
not g430 ( new_n568_, keyIn_0_0 );
or g431 ( new_n569_, N17, N21 );
and g432 ( new_n570_, N17, N21 );
not g433 ( new_n571_, new_n570_ );
and g434 ( new_n572_, new_n571_, new_n569_ );
or g435 ( new_n573_, new_n572_, new_n568_ );
and g436 ( new_n574_, new_n569_, new_n568_ );
and g437 ( new_n575_, new_n574_, new_n571_ );
not g438 ( new_n576_, new_n575_ );
and g439 ( new_n577_, new_n576_, new_n573_ );
not g440 ( new_n578_, keyIn_0_1 );
or g441 ( new_n579_, N25, N29 );
and g442 ( new_n580_, N25, N29 );
not g443 ( new_n581_, new_n580_ );
and g444 ( new_n582_, new_n581_, new_n579_ );
or g445 ( new_n583_, new_n582_, new_n578_ );
and g446 ( new_n584_, new_n579_, new_n578_ );
and g447 ( new_n585_, new_n584_, new_n581_ );
not g448 ( new_n586_, new_n585_ );
and g449 ( new_n587_, new_n586_, new_n583_ );
or g450 ( new_n588_, new_n577_, new_n587_ );
and g451 ( new_n589_, new_n577_, new_n587_ );
not g452 ( new_n590_, new_n589_ );
and g453 ( new_n591_, new_n590_, new_n588_ );
not g454 ( new_n592_, new_n591_ );
and g455 ( new_n593_, new_n473_, new_n592_ );
and g456 ( new_n594_, new_n478_, new_n591_ );
or g457 ( new_n595_, new_n594_, new_n593_ );
and g458 ( new_n596_, N133, N137 );
not g459 ( new_n597_, new_n596_ );
and g460 ( new_n598_, new_n595_, new_n597_ );
not g461 ( new_n599_, new_n598_ );
or g462 ( new_n600_, new_n595_, new_n597_ );
and g463 ( new_n601_, new_n599_, new_n600_ );
not g464 ( new_n602_, keyIn_0_15 );
and g465 ( new_n603_, new_n215_, new_n250_ );
and g466 ( new_n604_, N97, N113 );
or g467 ( new_n605_, new_n603_, new_n604_ );
not g468 ( new_n606_, new_n605_ );
and g469 ( new_n607_, new_n606_, new_n602_ );
and g470 ( new_n608_, new_n605_, keyIn_0_15 );
or g471 ( new_n609_, new_n607_, new_n608_ );
and g472 ( new_n610_, N65, N81 );
and g473 ( new_n611_, new_n160_, new_n139_ );
or g474 ( new_n612_, new_n611_, new_n610_ );
and g475 ( new_n613_, new_n609_, new_n612_ );
not g476 ( new_n614_, new_n613_ );
or g477 ( new_n615_, new_n609_, new_n612_ );
and g478 ( new_n616_, new_n614_, new_n615_ );
or g479 ( new_n617_, new_n601_, new_n616_ );
and g480 ( new_n618_, new_n601_, new_n616_ );
not g481 ( new_n619_, new_n618_ );
and g482 ( new_n620_, new_n619_, new_n617_ );
not g483 ( new_n621_, new_n620_ );
and g484 ( new_n622_, new_n567_, new_n621_ );
and g485 ( new_n623_, new_n592_, new_n542_ );
and g486 ( new_n624_, new_n591_, new_n541_ );
or g487 ( new_n625_, new_n623_, new_n624_ );
and g488 ( new_n626_, new_n625_, keyIn_0_11 );
not g489 ( new_n627_, new_n626_ );
or g490 ( new_n628_, new_n625_, keyIn_0_11 );
and g491 ( new_n629_, new_n627_, new_n628_ );
not g492 ( new_n630_, new_n629_ );
and g493 ( new_n631_, N136, N137 );
not g494 ( new_n632_, new_n631_ );
and g495 ( new_n633_, new_n630_, new_n632_ );
and g496 ( new_n634_, new_n629_, new_n631_ );
or g497 ( new_n635_, new_n633_, new_n634_ );
and g498 ( new_n636_, new_n154_, new_n145_ );
and g499 ( new_n637_, N77, N93 );
or g500 ( new_n638_, new_n636_, new_n637_ );
and g501 ( new_n639_, new_n219_, new_n236_ );
and g502 ( new_n640_, N109, N125 );
or g503 ( new_n641_, new_n639_, new_n640_ );
and g504 ( new_n642_, new_n638_, new_n641_ );
not g505 ( new_n643_, new_n642_ );
or g506 ( new_n644_, new_n638_, new_n641_ );
and g507 ( new_n645_, new_n643_, new_n644_ );
and g508 ( new_n646_, new_n635_, new_n645_ );
not g509 ( new_n647_, new_n646_ );
or g510 ( new_n648_, new_n635_, new_n645_ );
and g511 ( new_n649_, new_n647_, new_n648_ );
and g512 ( new_n650_, new_n622_, new_n649_ );
and g513 ( new_n651_, new_n523_, new_n650_ );
and g514 ( new_n652_, new_n420_, new_n651_ );
not g515 ( new_n653_, new_n652_ );
and g516 ( new_n654_, new_n653_, new_n138_ );
and g517 ( new_n655_, new_n652_, keyIn_0_41 );
or g518 ( new_n656_, new_n654_, new_n655_ );
and g519 ( new_n657_, new_n656_, N1 );
not g520 ( new_n658_, new_n656_ );
and g521 ( new_n659_, new_n658_, new_n194_ );
or g522 ( N724, new_n659_, new_n657_ );
not g523 ( new_n661_, keyIn_0_42 );
and g524 ( new_n662_, new_n419_, new_n388_ );
and g525 ( new_n663_, new_n662_, new_n651_ );
not g526 ( new_n664_, new_n663_ );
and g527 ( new_n665_, new_n664_, new_n661_ );
and g528 ( new_n666_, new_n663_, keyIn_0_42 );
or g529 ( new_n667_, new_n665_, new_n666_ );
and g530 ( new_n668_, new_n667_, new_n280_ );
not g531 ( new_n669_, new_n667_ );
and g532 ( new_n670_, new_n669_, N5 );
or g533 ( N725, new_n670_, new_n668_ );
and g534 ( new_n672_, new_n419_, new_n651_ );
and g535 ( new_n673_, new_n672_, new_n393_ );
not g536 ( new_n674_, new_n673_ );
and g537 ( new_n675_, new_n674_, N9 );
and g538 ( new_n676_, new_n673_, new_n319_ );
or g539 ( N726, new_n675_, new_n676_ );
and g540 ( new_n678_, new_n672_, new_n383_ );
not g541 ( new_n679_, new_n678_ );
and g542 ( new_n680_, new_n679_, N13 );
and g543 ( new_n681_, new_n678_, new_n363_ );
or g544 ( N727, new_n680_, new_n681_ );
or g545 ( new_n683_, new_n520_, new_n521_ );
or g546 ( new_n684_, new_n501_, new_n516_ );
and g547 ( new_n685_, new_n684_, new_n683_ );
not g548 ( new_n686_, new_n635_ );
not g549 ( new_n687_, new_n645_ );
and g550 ( new_n688_, new_n686_, new_n687_ );
or g551 ( new_n689_, new_n688_, new_n646_ );
and g552 ( new_n690_, new_n622_, new_n689_ );
and g553 ( new_n691_, new_n685_, new_n690_ );
and g554 ( new_n692_, new_n420_, new_n691_ );
not g555 ( new_n693_, new_n692_ );
and g556 ( new_n694_, new_n693_, N17 );
and g557 ( new_n695_, new_n692_, new_n192_ );
or g558 ( new_n696_, new_n694_, new_n695_ );
and g559 ( new_n697_, new_n696_, keyIn_0_54 );
not g560 ( new_n698_, keyIn_0_54 );
not g561 ( new_n699_, new_n696_ );
and g562 ( new_n700_, new_n699_, new_n698_ );
or g563 ( N728, new_n700_, new_n697_ );
and g564 ( new_n702_, new_n662_, new_n691_ );
not g565 ( new_n703_, new_n702_ );
and g566 ( new_n704_, new_n703_, N21 );
and g567 ( new_n705_, new_n702_, new_n278_ );
or g568 ( new_n706_, new_n704_, new_n705_ );
and g569 ( new_n707_, new_n706_, keyIn_0_55 );
not g570 ( new_n708_, keyIn_0_55 );
not g571 ( new_n709_, new_n706_ );
and g572 ( new_n710_, new_n709_, new_n708_ );
or g573 ( N729, new_n710_, new_n707_ );
and g574 ( new_n712_, new_n419_, new_n393_ );
and g575 ( new_n713_, new_n712_, new_n691_ );
not g576 ( new_n714_, new_n713_ );
and g577 ( new_n715_, new_n714_, N25 );
and g578 ( new_n716_, new_n713_, new_n320_ );
or g579 ( N730, new_n715_, new_n716_ );
not g580 ( new_n718_, keyIn_0_43 );
and g581 ( new_n719_, new_n419_, new_n383_ );
and g582 ( new_n720_, new_n719_, new_n691_ );
not g583 ( new_n721_, new_n720_ );
and g584 ( new_n722_, new_n721_, new_n718_ );
and g585 ( new_n723_, new_n720_, keyIn_0_43 );
or g586 ( new_n724_, new_n722_, new_n723_ );
and g587 ( new_n725_, new_n724_, N29 );
not g588 ( new_n726_, new_n724_ );
and g589 ( new_n727_, new_n726_, new_n361_ );
or g590 ( N731, new_n727_, new_n725_ );
and g591 ( new_n729_, new_n566_, new_n620_ );
and g592 ( new_n730_, new_n729_, new_n649_ );
and g593 ( new_n731_, new_n523_, new_n730_ );
and g594 ( new_n732_, new_n420_, new_n731_ );
not g595 ( new_n733_, new_n732_ );
and g596 ( new_n734_, new_n733_, N33 );
and g597 ( new_n735_, new_n732_, new_n197_ );
or g598 ( new_n736_, new_n734_, new_n735_ );
and g599 ( new_n737_, new_n736_, keyIn_0_56 );
not g600 ( new_n738_, keyIn_0_56 );
not g601 ( new_n739_, new_n736_ );
and g602 ( new_n740_, new_n739_, new_n738_ );
or g603 ( N732, new_n740_, new_n737_ );
and g604 ( new_n742_, new_n662_, new_n731_ );
not g605 ( new_n743_, new_n742_ );
and g606 ( new_n744_, new_n743_, new_n290_ );
and g607 ( new_n745_, new_n742_, N37 );
or g608 ( new_n746_, new_n744_, new_n745_ );
and g609 ( new_n747_, new_n746_, keyIn_0_57 );
not g610 ( new_n748_, keyIn_0_57 );
not g611 ( new_n749_, new_n746_ );
and g612 ( new_n750_, new_n749_, new_n748_ );
or g613 ( N733, new_n750_, new_n747_ );
not g614 ( new_n752_, keyIn_0_44 );
and g615 ( new_n753_, new_n712_, new_n731_ );
not g616 ( new_n754_, new_n753_ );
and g617 ( new_n755_, new_n754_, new_n752_ );
and g618 ( new_n756_, new_n753_, keyIn_0_44 );
or g619 ( new_n757_, new_n755_, new_n756_ );
and g620 ( new_n758_, new_n757_, N41 );
not g621 ( new_n759_, new_n757_ );
and g622 ( new_n760_, new_n759_, new_n324_ );
or g623 ( N734, new_n760_, new_n758_ );
not g624 ( new_n762_, keyIn_0_45 );
not g625 ( new_n763_, new_n385_ );
or g626 ( new_n764_, new_n416_, new_n410_ );
and g627 ( new_n765_, new_n764_, new_n763_ );
not g628 ( new_n766_, new_n405_ );
or g629 ( new_n767_, new_n388_, new_n766_ );
not g630 ( new_n768_, new_n341_ );
or g631 ( new_n769_, new_n308_, new_n768_ );
and g632 ( new_n770_, new_n767_, new_n769_ );
or g633 ( new_n771_, new_n770_, new_n383_ );
or g634 ( new_n772_, new_n397_, keyIn_0_36 );
and g635 ( new_n773_, new_n772_, new_n771_ );
and g636 ( new_n774_, new_n773_, new_n765_ );
or g637 ( new_n775_, new_n774_, new_n400_ );
not g638 ( new_n776_, new_n731_ );
or g639 ( new_n777_, new_n775_, new_n776_ );
and g640 ( new_n778_, new_n777_, new_n762_ );
and g641 ( new_n779_, new_n719_, new_n731_ );
and g642 ( new_n780_, new_n779_, keyIn_0_45 );
or g643 ( new_n781_, new_n780_, new_n778_ );
and g644 ( new_n782_, new_n781_, N45 );
or g645 ( new_n783_, new_n779_, keyIn_0_45 );
or g646 ( new_n784_, new_n777_, new_n762_ );
and g647 ( new_n785_, new_n783_, new_n784_ );
and g648 ( new_n786_, new_n785_, new_n373_ );
or g649 ( new_n787_, new_n782_, new_n786_ );
and g650 ( new_n788_, new_n787_, keyIn_0_58 );
not g651 ( new_n789_, keyIn_0_58 );
or g652 ( new_n790_, new_n785_, new_n373_ );
or g653 ( new_n791_, new_n781_, N45 );
and g654 ( new_n792_, new_n791_, new_n790_ );
and g655 ( new_n793_, new_n792_, new_n789_ );
or g656 ( N735, new_n788_, new_n793_ );
not g657 ( new_n795_, keyIn_0_27 );
and g658 ( new_n796_, new_n685_, new_n795_ );
and g659 ( new_n797_, new_n523_, keyIn_0_27 );
or g660 ( new_n798_, new_n797_, new_n796_ );
and g661 ( new_n799_, new_n689_, new_n620_ );
and g662 ( new_n800_, new_n799_, new_n566_ );
and g663 ( new_n801_, new_n798_, new_n800_ );
and g664 ( new_n802_, new_n419_, new_n801_ );
or g665 ( new_n803_, new_n802_, keyIn_0_39 );
not g666 ( new_n804_, keyIn_0_39 );
not g667 ( new_n805_, new_n801_ );
or g668 ( new_n806_, new_n774_, new_n805_ );
or g669 ( new_n807_, new_n806_, new_n804_ );
and g670 ( new_n808_, new_n803_, new_n807_ );
or g671 ( new_n809_, new_n808_, new_n210_ );
and g672 ( new_n810_, new_n809_, N49 );
and g673 ( new_n811_, new_n806_, new_n804_ );
and g674 ( new_n812_, new_n802_, keyIn_0_39 );
or g675 ( new_n813_, new_n812_, new_n811_ );
and g676 ( new_n814_, new_n813_, new_n211_ );
and g677 ( new_n815_, new_n814_, new_n198_ );
or g678 ( new_n816_, new_n810_, new_n815_ );
and g679 ( new_n817_, new_n816_, keyIn_0_59 );
not g680 ( new_n818_, keyIn_0_59 );
or g681 ( new_n819_, new_n814_, new_n198_ );
or g682 ( new_n820_, new_n809_, N49 );
and g683 ( new_n821_, new_n820_, new_n819_ );
and g684 ( new_n822_, new_n821_, new_n818_ );
or g685 ( N736, new_n817_, new_n822_ );
or g686 ( new_n824_, new_n808_, new_n308_ );
and g687 ( new_n825_, new_n824_, keyIn_0_46 );
not g688 ( new_n826_, keyIn_0_46 );
and g689 ( new_n827_, new_n813_, new_n388_ );
and g690 ( new_n828_, new_n827_, new_n826_ );
or g691 ( new_n829_, new_n825_, new_n828_ );
and g692 ( new_n830_, new_n829_, N53 );
or g693 ( new_n831_, new_n827_, new_n826_ );
or g694 ( new_n832_, new_n824_, keyIn_0_46 );
and g695 ( new_n833_, new_n832_, new_n831_ );
and g696 ( new_n834_, new_n833_, new_n288_ );
or g697 ( N737, new_n830_, new_n834_ );
and g698 ( new_n836_, new_n813_, new_n393_ );
not g699 ( new_n837_, new_n836_ );
and g700 ( new_n838_, new_n837_, N57 );
and g701 ( new_n839_, new_n836_, new_n325_ );
or g702 ( N738, new_n838_, new_n839_ );
and g703 ( new_n841_, new_n813_, new_n383_ );
not g704 ( new_n842_, new_n841_ );
and g705 ( new_n843_, new_n842_, N61 );
and g706 ( new_n844_, new_n841_, new_n371_ );
or g707 ( N739, new_n843_, new_n844_ );
not g708 ( new_n846_, keyIn_0_40 );
not g709 ( new_n847_, keyIn_0_38 );
not g710 ( new_n848_, keyIn_0_37 );
not g711 ( new_n849_, keyIn_0_31 );
and g712 ( new_n850_, new_n685_, new_n849_ );
not g713 ( new_n851_, new_n850_ );
or g714 ( new_n852_, new_n685_, new_n849_ );
and g715 ( new_n853_, new_n852_, new_n730_ );
and g716 ( new_n854_, new_n853_, new_n851_ );
and g717 ( new_n855_, new_n854_, new_n848_ );
not g718 ( new_n856_, new_n855_ );
or g719 ( new_n857_, new_n854_, new_n848_ );
not g720 ( new_n858_, keyIn_0_32 );
and g721 ( new_n859_, new_n685_, new_n858_ );
and g722 ( new_n860_, new_n523_, keyIn_0_32 );
not g723 ( new_n861_, keyIn_0_33 );
and g724 ( new_n862_, new_n689_, new_n861_ );
not g725 ( new_n863_, new_n622_ );
and g726 ( new_n864_, new_n649_, keyIn_0_33 );
or g727 ( new_n865_, new_n863_, new_n864_ );
or g728 ( new_n866_, new_n865_, new_n862_ );
or g729 ( new_n867_, new_n860_, new_n866_ );
or g730 ( new_n868_, new_n867_, new_n859_ );
and g731 ( new_n869_, new_n649_, keyIn_0_30 );
not g732 ( new_n870_, keyIn_0_30 );
and g733 ( new_n871_, new_n689_, new_n870_ );
or g734 ( new_n872_, new_n871_, new_n869_ );
not g735 ( new_n873_, keyIn_0_29 );
or g736 ( new_n874_, new_n620_, new_n873_ );
and g737 ( new_n875_, new_n620_, new_n873_ );
not g738 ( new_n876_, new_n875_ );
and g739 ( new_n877_, new_n876_, new_n874_ );
and g740 ( new_n878_, new_n877_, new_n567_ );
and g741 ( new_n879_, new_n872_, new_n878_ );
and g742 ( new_n880_, new_n879_, new_n523_ );
not g743 ( new_n881_, keyIn_0_28 );
and g744 ( new_n882_, new_n567_, new_n881_ );
and g745 ( new_n883_, new_n566_, keyIn_0_28 );
or g746 ( new_n884_, new_n882_, new_n883_ );
and g747 ( new_n885_, new_n884_, new_n799_ );
and g748 ( new_n886_, new_n885_, new_n685_ );
or g749 ( new_n887_, new_n880_, new_n886_ );
not g750 ( new_n888_, new_n887_ );
and g751 ( new_n889_, new_n868_, new_n888_ );
and g752 ( new_n890_, new_n889_, new_n857_ );
and g753 ( new_n891_, new_n890_, new_n856_ );
or g754 ( new_n892_, new_n891_, new_n847_ );
and g755 ( new_n893_, new_n891_, new_n847_ );
not g756 ( new_n894_, new_n893_ );
and g757 ( new_n895_, new_n894_, new_n892_ );
and g758 ( new_n896_, new_n400_, new_n393_ );
and g759 ( new_n897_, new_n411_, new_n896_ );
and g760 ( new_n898_, new_n895_, new_n897_ );
or g761 ( new_n899_, new_n898_, new_n846_ );
not g762 ( new_n900_, new_n730_ );
and g763 ( new_n901_, new_n523_, keyIn_0_31 );
or g764 ( new_n902_, new_n901_, new_n900_ );
or g765 ( new_n903_, new_n902_, new_n850_ );
and g766 ( new_n904_, new_n903_, keyIn_0_37 );
not g767 ( new_n905_, new_n859_ );
or g768 ( new_n906_, new_n685_, new_n858_ );
not g769 ( new_n907_, new_n862_ );
not g770 ( new_n908_, new_n864_ );
and g771 ( new_n909_, new_n908_, new_n622_ );
and g772 ( new_n910_, new_n909_, new_n907_ );
and g773 ( new_n911_, new_n906_, new_n910_ );
and g774 ( new_n912_, new_n911_, new_n905_ );
or g775 ( new_n913_, new_n912_, new_n887_ );
or g776 ( new_n914_, new_n904_, new_n913_ );
or g777 ( new_n915_, new_n914_, new_n855_ );
and g778 ( new_n916_, new_n915_, keyIn_0_38 );
or g779 ( new_n917_, new_n916_, new_n893_ );
not g780 ( new_n918_, new_n897_ );
or g781 ( new_n919_, new_n917_, new_n918_ );
or g782 ( new_n920_, new_n919_, keyIn_0_40 );
and g783 ( new_n921_, new_n920_, new_n899_ );
or g784 ( new_n922_, new_n921_, new_n620_ );
and g785 ( new_n923_, new_n922_, keyIn_0_47 );
not g786 ( new_n924_, keyIn_0_47 );
and g787 ( new_n925_, new_n919_, keyIn_0_40 );
and g788 ( new_n926_, new_n898_, new_n846_ );
or g789 ( new_n927_, new_n925_, new_n926_ );
and g790 ( new_n928_, new_n927_, new_n621_ );
and g791 ( new_n929_, new_n928_, new_n924_ );
or g792 ( new_n930_, new_n923_, new_n929_ );
and g793 ( new_n931_, new_n930_, new_n160_ );
or g794 ( new_n932_, new_n928_, new_n924_ );
or g795 ( new_n933_, new_n922_, keyIn_0_47 );
and g796 ( new_n934_, new_n933_, new_n932_ );
and g797 ( new_n935_, new_n934_, N65 );
or g798 ( N740, new_n931_, new_n935_ );
or g799 ( new_n937_, new_n921_, new_n567_ );
and g800 ( new_n938_, new_n937_, keyIn_0_48 );
not g801 ( new_n939_, keyIn_0_48 );
and g802 ( new_n940_, new_n927_, new_n566_ );
and g803 ( new_n941_, new_n940_, new_n939_ );
or g804 ( new_n942_, new_n938_, new_n941_ );
and g805 ( new_n943_, new_n942_, new_n161_ );
or g806 ( new_n944_, new_n940_, new_n939_ );
or g807 ( new_n945_, new_n937_, keyIn_0_48 );
and g808 ( new_n946_, new_n945_, new_n944_ );
and g809 ( new_n947_, new_n946_, N69 );
or g810 ( N741, new_n943_, new_n947_ );
and g811 ( new_n949_, new_n927_, new_n523_ );
not g812 ( new_n950_, new_n949_ );
and g813 ( new_n951_, new_n950_, N73 );
and g814 ( new_n952_, new_n949_, new_n153_ );
or g815 ( N742, new_n951_, new_n952_ );
or g816 ( new_n954_, new_n921_, new_n649_ );
and g817 ( new_n955_, new_n954_, N77 );
and g818 ( new_n956_, new_n927_, new_n689_ );
and g819 ( new_n957_, new_n956_, new_n154_ );
or g820 ( new_n958_, new_n955_, new_n957_ );
and g821 ( new_n959_, new_n958_, keyIn_0_60 );
not g822 ( new_n960_, keyIn_0_60 );
or g823 ( new_n961_, new_n956_, new_n154_ );
or g824 ( new_n962_, new_n954_, N77 );
and g825 ( new_n963_, new_n962_, new_n961_ );
and g826 ( new_n964_, new_n963_, new_n960_ );
or g827 ( N743, new_n959_, new_n964_ );
and g828 ( new_n966_, new_n388_, keyIn_0_34 );
not g829 ( new_n967_, new_n966_ );
or g830 ( new_n968_, new_n388_, keyIn_0_34 );
and g831 ( new_n969_, new_n340_, new_n211_ );
and g832 ( new_n970_, new_n969_, new_n383_ );
and g833 ( new_n971_, new_n968_, new_n970_ );
and g834 ( new_n972_, new_n971_, new_n967_ );
and g835 ( new_n973_, new_n895_, new_n972_ );
and g836 ( new_n974_, new_n973_, new_n621_ );
not g837 ( new_n975_, new_n974_ );
and g838 ( new_n976_, new_n975_, N81 );
and g839 ( new_n977_, new_n974_, new_n139_ );
or g840 ( N744, new_n976_, new_n977_ );
and g841 ( new_n979_, new_n895_, new_n566_ );
and g842 ( new_n980_, new_n979_, new_n972_ );
not g843 ( new_n981_, new_n980_ );
and g844 ( new_n982_, new_n981_, keyIn_0_49 );
not g845 ( new_n983_, keyIn_0_49 );
and g846 ( new_n984_, new_n980_, new_n983_ );
or g847 ( new_n985_, new_n982_, new_n984_ );
and g848 ( new_n986_, new_n985_, N85 );
not g849 ( new_n987_, new_n985_ );
and g850 ( new_n988_, new_n987_, new_n140_ );
or g851 ( N745, new_n988_, new_n986_ );
and g852 ( new_n990_, new_n895_, new_n523_ );
and g853 ( new_n991_, new_n990_, new_n972_ );
not g854 ( new_n992_, new_n991_ );
and g855 ( new_n993_, new_n992_, N89 );
and g856 ( new_n994_, new_n991_, new_n144_ );
or g857 ( new_n995_, new_n993_, new_n994_ );
and g858 ( new_n996_, new_n995_, keyIn_0_61 );
not g859 ( new_n997_, keyIn_0_61 );
not g860 ( new_n998_, new_n995_ );
and g861 ( new_n999_, new_n998_, new_n997_ );
or g862 ( N746, new_n999_, new_n996_ );
and g863 ( new_n1001_, new_n973_, new_n689_ );
not g864 ( new_n1002_, new_n1001_ );
and g865 ( new_n1003_, new_n1002_, N93 );
and g866 ( new_n1004_, new_n1001_, new_n145_ );
or g867 ( N747, new_n1003_, new_n1004_ );
and g868 ( new_n1006_, new_n210_, keyIn_0_35 );
not g869 ( new_n1007_, new_n1006_ );
or g870 ( new_n1008_, new_n210_, keyIn_0_35 );
and g871 ( new_n1009_, new_n1007_, new_n1008_ );
and g872 ( new_n1010_, new_n896_, new_n1009_ );
and g873 ( new_n1011_, new_n1010_, new_n388_ );
and g874 ( new_n1012_, new_n895_, new_n1011_ );
and g875 ( new_n1013_, new_n1012_, new_n621_ );
not g876 ( new_n1014_, new_n1013_ );
and g877 ( new_n1015_, new_n1014_, N97 );
and g878 ( new_n1016_, new_n1013_, new_n215_ );
or g879 ( N748, new_n1015_, new_n1016_ );
and g880 ( new_n1018_, new_n979_, new_n1011_ );
not g881 ( new_n1019_, new_n1018_ );
and g882 ( new_n1020_, new_n1019_, keyIn_0_50 );
not g883 ( new_n1021_, keyIn_0_50 );
and g884 ( new_n1022_, new_n1018_, new_n1021_ );
or g885 ( new_n1023_, new_n1020_, new_n1022_ );
and g886 ( new_n1024_, new_n1023_, N101 );
not g887 ( new_n1025_, new_n1023_ );
and g888 ( new_n1026_, new_n1025_, new_n213_ );
or g889 ( N749, new_n1026_, new_n1024_ );
and g890 ( new_n1028_, new_n1012_, new_n523_ );
not g891 ( new_n1029_, new_n1028_ );
and g892 ( new_n1030_, new_n1029_, N105 );
and g893 ( new_n1031_, new_n1028_, new_n218_ );
or g894 ( N750, new_n1030_, new_n1031_ );
and g895 ( new_n1033_, new_n1012_, new_n689_ );
not g896 ( new_n1034_, new_n1033_ );
and g897 ( new_n1035_, new_n1034_, N109 );
and g898 ( new_n1036_, new_n1033_, new_n219_ );
or g899 ( N751, new_n1035_, new_n1036_ );
and g900 ( new_n1038_, new_n407_, new_n383_ );
and g901 ( new_n1039_, new_n895_, new_n1038_ );
and g902 ( new_n1040_, new_n1039_, new_n621_ );
not g903 ( new_n1041_, new_n1040_ );
and g904 ( new_n1042_, new_n1041_, N113 );
and g905 ( new_n1043_, new_n1040_, new_n250_ );
or g906 ( N752, new_n1042_, new_n1043_ );
and g907 ( new_n1045_, new_n979_, new_n1038_ );
not g908 ( new_n1046_, new_n1045_ );
and g909 ( new_n1047_, new_n1046_, keyIn_0_51 );
not g910 ( new_n1048_, keyIn_0_51 );
and g911 ( new_n1049_, new_n1045_, new_n1048_ );
or g912 ( new_n1050_, new_n1047_, new_n1049_ );
and g913 ( new_n1051_, new_n1050_, new_n248_ );
not g914 ( new_n1052_, new_n1050_ );
and g915 ( new_n1053_, new_n1052_, N117 );
or g916 ( N753, new_n1053_, new_n1051_ );
not g917 ( new_n1055_, keyIn_0_62 );
or g918 ( new_n1056_, new_n917_, new_n685_ );
not g919 ( new_n1057_, new_n1038_ );
or g920 ( new_n1058_, new_n1056_, new_n1057_ );
and g921 ( new_n1059_, new_n1058_, keyIn_0_52 );
not g922 ( new_n1060_, keyIn_0_52 );
and g923 ( new_n1061_, new_n990_, new_n1038_ );
and g924 ( new_n1062_, new_n1061_, new_n1060_ );
or g925 ( new_n1063_, new_n1059_, new_n1062_ );
and g926 ( new_n1064_, new_n1063_, new_n235_ );
or g927 ( new_n1065_, new_n1061_, new_n1060_ );
or g928 ( new_n1066_, new_n1058_, keyIn_0_52 );
and g929 ( new_n1067_, new_n1066_, new_n1065_ );
and g930 ( new_n1068_, new_n1067_, N121 );
or g931 ( new_n1069_, new_n1064_, new_n1068_ );
and g932 ( new_n1070_, new_n1069_, new_n1055_ );
or g933 ( new_n1071_, new_n1067_, N121 );
or g934 ( new_n1072_, new_n1063_, new_n235_ );
and g935 ( new_n1073_, new_n1071_, new_n1072_ );
and g936 ( new_n1074_, new_n1073_, keyIn_0_62 );
or g937 ( N754, new_n1070_, new_n1074_ );
not g938 ( new_n1076_, keyIn_0_63 );
or g939 ( new_n1077_, new_n917_, new_n1057_ );
or g940 ( new_n1078_, new_n1077_, new_n649_ );
and g941 ( new_n1079_, new_n1078_, keyIn_0_53 );
not g942 ( new_n1080_, keyIn_0_53 );
and g943 ( new_n1081_, new_n1039_, new_n689_ );
and g944 ( new_n1082_, new_n1081_, new_n1080_ );
or g945 ( new_n1083_, new_n1079_, new_n1082_ );
and g946 ( new_n1084_, new_n1083_, N125 );
or g947 ( new_n1085_, new_n1081_, new_n1080_ );
or g948 ( new_n1086_, new_n1078_, keyIn_0_53 );
and g949 ( new_n1087_, new_n1086_, new_n1085_ );
and g950 ( new_n1088_, new_n1087_, new_n236_ );
or g951 ( new_n1089_, new_n1084_, new_n1088_ );
and g952 ( new_n1090_, new_n1089_, new_n1076_ );
or g953 ( new_n1091_, new_n1087_, new_n236_ );
or g954 ( new_n1092_, new_n1083_, N125 );
and g955 ( new_n1093_, new_n1091_, new_n1092_ );
and g956 ( new_n1094_, new_n1093_, keyIn_0_63 );
or g957 ( N755, new_n1090_, new_n1094_ );
endmodule