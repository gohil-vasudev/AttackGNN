module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736;

  INV_X2 U7417 ( .A(b_30_), .ZN(n7344) );
  INV_X2 U7418 ( .A(b_3_), .ZN(n7659) );
  INV_X2 U7419 ( .A(b_5_), .ZN(n7715) );
  INV_X2 U7420 ( .A(b_7_), .ZN(n7798) );
  INV_X2 U7421 ( .A(b_9_), .ZN(n7912) );
  INV_X2 U7422 ( .A(b_11_), .ZN(n8050) );
  XOR2_X1 U7423 ( .A(n7321), .B(n7322), .Z(Result_mul_9_) );
  AND2_X1 U7424 ( .A1(n7323), .A2(n7324), .ZN(n7322) );
  OR2_X1 U7425 ( .A1(n7325), .A2(n7326), .ZN(n7324) );
  INV_X1 U7426 ( .A(n7327), .ZN(n7323) );
  XOR2_X1 U7427 ( .A(n7328), .B(n7329), .Z(Result_mul_8_) );
  XOR2_X1 U7428 ( .A(n7330), .B(n7331), .Z(Result_mul_7_) );
  AND2_X1 U7429 ( .A1(n7332), .A2(n7333), .ZN(n7331) );
  OR2_X1 U7430 ( .A1(n7334), .A2(n7335), .ZN(n7333) );
  INV_X1 U7431 ( .A(n7336), .ZN(n7332) );
  XOR2_X1 U7432 ( .A(n7337), .B(n7338), .Z(Result_mul_6_) );
  OR2_X1 U7433 ( .A1(n7339), .A2(n7340), .ZN(Result_mul_62_) );
  AND2_X1 U7434 ( .A1(b_31_), .A2(n7341), .ZN(n7340) );
  OR2_X1 U7435 ( .A1(n7342), .A2(n7343), .ZN(n7341) );
  AND2_X1 U7436 ( .A1(a_30_), .A2(n7344), .ZN(n7342) );
  AND2_X1 U7437 ( .A1(b_30_), .A2(n7345), .ZN(n7339) );
  OR2_X1 U7438 ( .A1(n7346), .A2(n7347), .ZN(n7345) );
  AND2_X1 U7439 ( .A1(a_31_), .A2(n7348), .ZN(n7346) );
  XNOR2_X1 U7440 ( .A(n7349), .B(n7350), .ZN(Result_mul_61_) );
  XNOR2_X1 U7441 ( .A(n7351), .B(n7352), .ZN(n7349) );
  XOR2_X1 U7442 ( .A(n7353), .B(n7354), .Z(Result_mul_60_) );
  XNOR2_X1 U7443 ( .A(n7355), .B(n7356), .ZN(n7353) );
  XOR2_X1 U7444 ( .A(n7357), .B(n7358), .Z(Result_mul_5_) );
  AND2_X1 U7445 ( .A1(n7359), .A2(n7360), .ZN(n7358) );
  OR2_X1 U7446 ( .A1(n7361), .A2(n7362), .ZN(n7360) );
  INV_X1 U7447 ( .A(n7363), .ZN(n7359) );
  XNOR2_X1 U7448 ( .A(n7364), .B(n7365), .ZN(Result_mul_59_) );
  XOR2_X1 U7449 ( .A(n7366), .B(n7367), .Z(n7365) );
  XNOR2_X1 U7450 ( .A(n7368), .B(n7369), .ZN(Result_mul_58_) );
  XOR2_X1 U7451 ( .A(n7370), .B(n7371), .Z(n7369) );
  XNOR2_X1 U7452 ( .A(n7372), .B(n7373), .ZN(Result_mul_57_) );
  XOR2_X1 U7453 ( .A(n7374), .B(n7375), .Z(n7373) );
  XNOR2_X1 U7454 ( .A(n7376), .B(n7377), .ZN(Result_mul_56_) );
  XOR2_X1 U7455 ( .A(n7378), .B(n7379), .Z(n7377) );
  XNOR2_X1 U7456 ( .A(n7380), .B(n7381), .ZN(Result_mul_55_) );
  XOR2_X1 U7457 ( .A(n7382), .B(n7383), .Z(n7381) );
  XNOR2_X1 U7458 ( .A(n7384), .B(n7385), .ZN(Result_mul_54_) );
  XOR2_X1 U7459 ( .A(n7386), .B(n7387), .Z(n7385) );
  XNOR2_X1 U7460 ( .A(n7388), .B(n7389), .ZN(Result_mul_53_) );
  XOR2_X1 U7461 ( .A(n7390), .B(n7391), .Z(n7389) );
  XNOR2_X1 U7462 ( .A(n7392), .B(n7393), .ZN(Result_mul_52_) );
  XOR2_X1 U7463 ( .A(n7394), .B(n7395), .Z(n7393) );
  XNOR2_X1 U7464 ( .A(n7396), .B(n7397), .ZN(Result_mul_51_) );
  XOR2_X1 U7465 ( .A(n7398), .B(n7399), .Z(n7397) );
  XNOR2_X1 U7466 ( .A(n7400), .B(n7401), .ZN(Result_mul_50_) );
  XOR2_X1 U7467 ( .A(n7402), .B(n7403), .Z(n7401) );
  XOR2_X1 U7468 ( .A(n7404), .B(n7405), .Z(Result_mul_4_) );
  XNOR2_X1 U7469 ( .A(n7406), .B(n7407), .ZN(Result_mul_49_) );
  XOR2_X1 U7470 ( .A(n7408), .B(n7409), .Z(n7407) );
  XNOR2_X1 U7471 ( .A(n7410), .B(n7411), .ZN(Result_mul_48_) );
  XOR2_X1 U7472 ( .A(n7412), .B(n7413), .Z(n7411) );
  XNOR2_X1 U7473 ( .A(n7414), .B(n7415), .ZN(Result_mul_47_) );
  XOR2_X1 U7474 ( .A(n7416), .B(n7417), .Z(n7415) );
  XNOR2_X1 U7475 ( .A(n7418), .B(n7419), .ZN(Result_mul_46_) );
  XOR2_X1 U7476 ( .A(n7420), .B(n7421), .Z(n7419) );
  XNOR2_X1 U7477 ( .A(n7422), .B(n7423), .ZN(Result_mul_45_) );
  XOR2_X1 U7478 ( .A(n7424), .B(n7425), .Z(n7423) );
  XNOR2_X1 U7479 ( .A(n7426), .B(n7427), .ZN(Result_mul_44_) );
  XOR2_X1 U7480 ( .A(n7428), .B(n7429), .Z(n7427) );
  XNOR2_X1 U7481 ( .A(n7430), .B(n7431), .ZN(Result_mul_43_) );
  XOR2_X1 U7482 ( .A(n7432), .B(n7433), .Z(n7431) );
  XNOR2_X1 U7483 ( .A(n7434), .B(n7435), .ZN(Result_mul_42_) );
  XOR2_X1 U7484 ( .A(n7436), .B(n7437), .Z(n7435) );
  XNOR2_X1 U7485 ( .A(n7438), .B(n7439), .ZN(Result_mul_41_) );
  XOR2_X1 U7486 ( .A(n7440), .B(n7441), .Z(n7439) );
  XNOR2_X1 U7487 ( .A(n7442), .B(n7443), .ZN(Result_mul_40_) );
  XOR2_X1 U7488 ( .A(n7444), .B(n7445), .Z(n7443) );
  XOR2_X1 U7489 ( .A(n7446), .B(n7447), .Z(Result_mul_3_) );
  AND2_X1 U7490 ( .A1(n7448), .A2(n7449), .ZN(n7447) );
  OR2_X1 U7491 ( .A1(n7450), .A2(n7451), .ZN(n7449) );
  INV_X1 U7492 ( .A(n7452), .ZN(n7448) );
  XNOR2_X1 U7493 ( .A(n7453), .B(n7454), .ZN(Result_mul_39_) );
  XOR2_X1 U7494 ( .A(n7455), .B(n7456), .Z(n7454) );
  XNOR2_X1 U7495 ( .A(n7457), .B(n7458), .ZN(Result_mul_38_) );
  XOR2_X1 U7496 ( .A(n7459), .B(n7460), .Z(n7458) );
  XNOR2_X1 U7497 ( .A(n7461), .B(n7462), .ZN(Result_mul_37_) );
  XOR2_X1 U7498 ( .A(n7463), .B(n7464), .Z(n7462) );
  XNOR2_X1 U7499 ( .A(n7465), .B(n7466), .ZN(Result_mul_36_) );
  XOR2_X1 U7500 ( .A(n7467), .B(n7468), .Z(n7466) );
  XNOR2_X1 U7501 ( .A(n7469), .B(n7470), .ZN(Result_mul_35_) );
  XOR2_X1 U7502 ( .A(n7471), .B(n7472), .Z(n7470) );
  XNOR2_X1 U7503 ( .A(n7473), .B(n7474), .ZN(Result_mul_34_) );
  XOR2_X1 U7504 ( .A(n7475), .B(n7476), .Z(n7474) );
  XNOR2_X1 U7505 ( .A(n7477), .B(n7478), .ZN(Result_mul_33_) );
  XOR2_X1 U7506 ( .A(n7479), .B(n7480), .Z(n7478) );
  XNOR2_X1 U7507 ( .A(n7481), .B(n7482), .ZN(Result_mul_32_) );
  XOR2_X1 U7508 ( .A(n7483), .B(n7484), .Z(n7482) );
  XNOR2_X1 U7509 ( .A(n7485), .B(n7486), .ZN(Result_mul_31_) );
  AND2_X1 U7510 ( .A1(n7487), .A2(n7488), .ZN(Result_mul_30_) );
  OR2_X1 U7511 ( .A1(n7489), .A2(n7490), .ZN(n7487) );
  AND2_X1 U7512 ( .A1(n7491), .A2(n7486), .ZN(n7489) );
  XOR2_X1 U7513 ( .A(n7492), .B(n7493), .Z(Result_mul_2_) );
  XNOR2_X1 U7514 ( .A(n7488), .B(n7494), .ZN(Result_mul_29_) );
  AND2_X1 U7515 ( .A1(n7495), .A2(n7496), .ZN(n7494) );
  INV_X1 U7516 ( .A(n7497), .ZN(n7488) );
  XOR2_X1 U7517 ( .A(n7498), .B(n7499), .Z(Result_mul_28_) );
  AND2_X1 U7518 ( .A1(n7500), .A2(n7501), .ZN(n7499) );
  XOR2_X1 U7519 ( .A(n7502), .B(n7503), .Z(Result_mul_27_) );
  AND2_X1 U7520 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
  INV_X1 U7521 ( .A(n7506), .ZN(n7505) );
  XOR2_X1 U7522 ( .A(n7507), .B(n7508), .Z(Result_mul_26_) );
  AND2_X1 U7523 ( .A1(n7509), .A2(n7510), .ZN(n7508) );
  INV_X1 U7524 ( .A(n7511), .ZN(n7510) );
  XOR2_X1 U7525 ( .A(n7512), .B(n7513), .Z(Result_mul_25_) );
  AND2_X1 U7526 ( .A1(n7514), .A2(n7515), .ZN(n7513) );
  XOR2_X1 U7527 ( .A(n7516), .B(n7517), .Z(Result_mul_24_) );
  AND2_X1 U7528 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
  INV_X1 U7529 ( .A(n7520), .ZN(n7518) );
  XOR2_X1 U7530 ( .A(n7521), .B(n7522), .Z(Result_mul_23_) );
  AND2_X1 U7531 ( .A1(n7523), .A2(n7524), .ZN(n7522) );
  INV_X1 U7532 ( .A(n7525), .ZN(n7524) );
  XOR2_X1 U7533 ( .A(n7526), .B(n7527), .Z(Result_mul_22_) );
  AND2_X1 U7534 ( .A1(n7528), .A2(n7529), .ZN(n7527) );
  OR2_X1 U7535 ( .A1(n7530), .A2(n7531), .ZN(n7528) );
  INV_X1 U7536 ( .A(n7532), .ZN(n7530) );
  XOR2_X1 U7537 ( .A(n7533), .B(n7534), .Z(Result_mul_21_) );
  AND2_X1 U7538 ( .A1(n7535), .A2(n7536), .ZN(n7534) );
  INV_X1 U7539 ( .A(n7537), .ZN(n7536) );
  XOR2_X1 U7540 ( .A(n7538), .B(n7539), .Z(Result_mul_20_) );
  AND2_X1 U7541 ( .A1(n7540), .A2(n7541), .ZN(n7539) );
  XOR2_X1 U7542 ( .A(n7542), .B(n7543), .Z(Result_mul_1_) );
  AND2_X1 U7543 ( .A1(n7544), .A2(n7545), .ZN(n7543) );
  OR2_X1 U7544 ( .A1(n7546), .A2(n7547), .ZN(n7545) );
  AND2_X1 U7545 ( .A1(n7548), .A2(n7549), .ZN(n7546) );
  INV_X1 U7546 ( .A(n7550), .ZN(n7544) );
  XOR2_X1 U7547 ( .A(n7551), .B(n7552), .Z(Result_mul_19_) );
  AND2_X1 U7548 ( .A1(n7553), .A2(n7554), .ZN(n7552) );
  INV_X1 U7549 ( .A(n7555), .ZN(n7554) );
  XOR2_X1 U7550 ( .A(n7556), .B(n7557), .Z(Result_mul_18_) );
  AND2_X1 U7551 ( .A1(n7558), .A2(n7559), .ZN(n7557) );
  OR2_X1 U7552 ( .A1(n7560), .A2(n7561), .ZN(n7558) );
  INV_X1 U7553 ( .A(n7562), .ZN(n7560) );
  XOR2_X1 U7554 ( .A(n7563), .B(n7564), .Z(Result_mul_17_) );
  AND2_X1 U7555 ( .A1(n7565), .A2(n7566), .ZN(n7564) );
  XOR2_X1 U7556 ( .A(n7567), .B(n7568), .Z(Result_mul_16_) );
  AND2_X1 U7557 ( .A1(n7569), .A2(n7570), .ZN(n7568) );
  INV_X1 U7558 ( .A(n7571), .ZN(n7569) );
  XOR2_X1 U7559 ( .A(n7572), .B(n7573), .Z(Result_mul_15_) );
  AND2_X1 U7560 ( .A1(n7574), .A2(n7575), .ZN(n7573) );
  INV_X1 U7561 ( .A(n7576), .ZN(n7575) );
  OR2_X1 U7562 ( .A1(n7577), .A2(n7578), .ZN(Result_mul_14_) );
  AND2_X1 U7563 ( .A1(n7579), .A2(n7580), .ZN(n7578) );
  AND2_X1 U7564 ( .A1(n7581), .A2(n7582), .ZN(n7579) );
  OR2_X1 U7565 ( .A1(n7583), .A2(n7584), .ZN(n7581) );
  INV_X1 U7566 ( .A(n7585), .ZN(n7577) );
  OR2_X1 U7567 ( .A1(n7582), .A2(n7580), .ZN(n7585) );
  INV_X1 U7568 ( .A(n7586), .ZN(n7580) );
  OR2_X1 U7569 ( .A1(n7587), .A2(n7588), .ZN(n7582) );
  XOR2_X1 U7570 ( .A(n7589), .B(n7590), .Z(Result_mul_13_) );
  AND2_X1 U7571 ( .A1(n7591), .A2(n7592), .ZN(n7590) );
  OR2_X1 U7572 ( .A1(n7593), .A2(n7594), .ZN(n7592) );
  INV_X1 U7573 ( .A(n7595), .ZN(n7591) );
  OR2_X1 U7574 ( .A1(n7596), .A2(n7597), .ZN(Result_mul_12_) );
  AND2_X1 U7575 ( .A1(n7598), .A2(n7599), .ZN(n7597) );
  AND2_X1 U7576 ( .A1(n7600), .A2(n7601), .ZN(n7598) );
  OR2_X1 U7577 ( .A1(n7602), .A2(n7603), .ZN(n7600) );
  INV_X1 U7578 ( .A(n7604), .ZN(n7596) );
  OR2_X1 U7579 ( .A1(n7601), .A2(n7599), .ZN(n7604) );
  INV_X1 U7580 ( .A(n7605), .ZN(n7599) );
  OR2_X1 U7581 ( .A1(n7606), .A2(n7607), .ZN(n7601) );
  XOR2_X1 U7582 ( .A(n7608), .B(n7609), .Z(Result_mul_11_) );
  AND2_X1 U7583 ( .A1(n7610), .A2(n7611), .ZN(n7609) );
  OR2_X1 U7584 ( .A1(n7612), .A2(n7613), .ZN(n7611) );
  INV_X1 U7585 ( .A(n7614), .ZN(n7610) );
  OR2_X1 U7586 ( .A1(n7615), .A2(n7616), .ZN(Result_mul_10_) );
  AND2_X1 U7587 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  AND2_X1 U7588 ( .A1(n7619), .A2(n7620), .ZN(n7617) );
  OR2_X1 U7589 ( .A1(n7621), .A2(n7622), .ZN(n7619) );
  INV_X1 U7590 ( .A(n7623), .ZN(n7615) );
  OR2_X1 U7591 ( .A1(n7620), .A2(n7618), .ZN(n7623) );
  INV_X1 U7592 ( .A(n7624), .ZN(n7618) );
  OR2_X1 U7593 ( .A1(n7625), .A2(n7626), .ZN(n7620) );
  OR2_X1 U7594 ( .A1(n7627), .A2(n7628), .ZN(Result_mul_0_) );
  OR2_X1 U7595 ( .A1(n7550), .A2(n7629), .ZN(n7628) );
  AND2_X1 U7596 ( .A1(n7542), .A2(n7547), .ZN(n7629) );
  AND2_X1 U7597 ( .A1(n7492), .A2(n7493), .ZN(n7542) );
  XNOR2_X1 U7598 ( .A(n7549), .B(n7630), .ZN(n7493) );
  OR2_X1 U7599 ( .A1(n7631), .A2(n7632), .ZN(n7492) );
  OR2_X1 U7600 ( .A1(n7633), .A2(n7452), .ZN(n7631) );
  AND2_X1 U7601 ( .A1(n7450), .A2(n7451), .ZN(n7452) );
  AND2_X1 U7602 ( .A1(n7634), .A2(n7635), .ZN(n7451) );
  INV_X1 U7603 ( .A(n7636), .ZN(n7634) );
  AND2_X1 U7604 ( .A1(n7446), .A2(n7450), .ZN(n7633) );
  INV_X1 U7605 ( .A(n7637), .ZN(n7450) );
  OR2_X1 U7606 ( .A1(n7638), .A2(n7632), .ZN(n7637) );
  INV_X1 U7607 ( .A(n7639), .ZN(n7632) );
  OR2_X1 U7608 ( .A1(n7640), .A2(n7641), .ZN(n7639) );
  AND2_X1 U7609 ( .A1(n7640), .A2(n7641), .ZN(n7638) );
  OR2_X1 U7610 ( .A1(n7642), .A2(n7643), .ZN(n7641) );
  AND2_X1 U7611 ( .A1(n7644), .A2(n7645), .ZN(n7643) );
  AND2_X1 U7612 ( .A1(n7646), .A2(n7647), .ZN(n7642) );
  OR2_X1 U7613 ( .A1(n7645), .A2(n7644), .ZN(n7647) );
  XOR2_X1 U7614 ( .A(n7648), .B(n7649), .Z(n7640) );
  XOR2_X1 U7615 ( .A(n7650), .B(n7651), .Z(n7649) );
  AND2_X1 U7616 ( .A1(n7404), .A2(n7405), .ZN(n7446) );
  XNOR2_X1 U7617 ( .A(n7635), .B(n7636), .ZN(n7405) );
  OR2_X1 U7618 ( .A1(n7652), .A2(n7653), .ZN(n7636) );
  AND2_X1 U7619 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  AND2_X1 U7620 ( .A1(n7656), .A2(n7657), .ZN(n7652) );
  OR2_X1 U7621 ( .A1(n7655), .A2(n7654), .ZN(n7657) );
  XNOR2_X1 U7622 ( .A(n7646), .B(n7658), .ZN(n7635) );
  XOR2_X1 U7623 ( .A(n7645), .B(n7644), .Z(n7658) );
  OR2_X1 U7624 ( .A1(n7659), .A2(n7660), .ZN(n7644) );
  OR2_X1 U7625 ( .A1(n7661), .A2(n7662), .ZN(n7645) );
  AND2_X1 U7626 ( .A1(n7663), .A2(n7664), .ZN(n7662) );
  AND2_X1 U7627 ( .A1(n7665), .A2(n7666), .ZN(n7661) );
  OR2_X1 U7628 ( .A1(n7664), .A2(n7663), .ZN(n7666) );
  XOR2_X1 U7629 ( .A(n7667), .B(n7668), .Z(n7646) );
  XOR2_X1 U7630 ( .A(n7669), .B(n7670), .Z(n7668) );
  OR2_X1 U7631 ( .A1(n7671), .A2(n7672), .ZN(n7404) );
  OR2_X1 U7632 ( .A1(n7673), .A2(n7363), .ZN(n7671) );
  AND2_X1 U7633 ( .A1(n7361), .A2(n7362), .ZN(n7363) );
  AND2_X1 U7634 ( .A1(n7674), .A2(n7675), .ZN(n7362) );
  INV_X1 U7635 ( .A(n7676), .ZN(n7674) );
  AND2_X1 U7636 ( .A1(n7357), .A2(n7361), .ZN(n7673) );
  INV_X1 U7637 ( .A(n7677), .ZN(n7361) );
  OR2_X1 U7638 ( .A1(n7678), .A2(n7672), .ZN(n7677) );
  INV_X1 U7639 ( .A(n7679), .ZN(n7672) );
  OR2_X1 U7640 ( .A1(n7680), .A2(n7681), .ZN(n7679) );
  AND2_X1 U7641 ( .A1(n7680), .A2(n7681), .ZN(n7678) );
  OR2_X1 U7642 ( .A1(n7682), .A2(n7683), .ZN(n7681) );
  AND2_X1 U7643 ( .A1(n7684), .A2(n7685), .ZN(n7683) );
  AND2_X1 U7644 ( .A1(n7686), .A2(n7687), .ZN(n7682) );
  OR2_X1 U7645 ( .A1(n7685), .A2(n7684), .ZN(n7687) );
  XOR2_X1 U7646 ( .A(n7656), .B(n7688), .Z(n7680) );
  XOR2_X1 U7647 ( .A(n7655), .B(n7654), .Z(n7688) );
  OR2_X1 U7648 ( .A1(n7689), .A2(n7660), .ZN(n7654) );
  OR2_X1 U7649 ( .A1(n7690), .A2(n7691), .ZN(n7655) );
  AND2_X1 U7650 ( .A1(n7692), .A2(n7693), .ZN(n7691) );
  AND2_X1 U7651 ( .A1(n7694), .A2(n7695), .ZN(n7690) );
  OR2_X1 U7652 ( .A1(n7693), .A2(n7692), .ZN(n7695) );
  XOR2_X1 U7653 ( .A(n7665), .B(n7696), .Z(n7656) );
  XOR2_X1 U7654 ( .A(n7664), .B(n7663), .Z(n7696) );
  OR2_X1 U7655 ( .A1(n7659), .A2(n7697), .ZN(n7663) );
  OR2_X1 U7656 ( .A1(n7698), .A2(n7699), .ZN(n7664) );
  AND2_X1 U7657 ( .A1(n7700), .A2(n7701), .ZN(n7699) );
  AND2_X1 U7658 ( .A1(n7702), .A2(n7703), .ZN(n7698) );
  OR2_X1 U7659 ( .A1(n7701), .A2(n7700), .ZN(n7703) );
  XNOR2_X1 U7660 ( .A(n7704), .B(n7705), .ZN(n7665) );
  XNOR2_X1 U7661 ( .A(n7706), .B(n7707), .ZN(n7704) );
  AND2_X1 U7662 ( .A1(n7337), .A2(n7338), .ZN(n7357) );
  XNOR2_X1 U7663 ( .A(n7675), .B(n7676), .ZN(n7338) );
  OR2_X1 U7664 ( .A1(n7708), .A2(n7709), .ZN(n7676) );
  AND2_X1 U7665 ( .A1(n7710), .A2(n7711), .ZN(n7709) );
  AND2_X1 U7666 ( .A1(n7712), .A2(n7713), .ZN(n7708) );
  OR2_X1 U7667 ( .A1(n7711), .A2(n7710), .ZN(n7713) );
  XNOR2_X1 U7668 ( .A(n7686), .B(n7714), .ZN(n7675) );
  XOR2_X1 U7669 ( .A(n7685), .B(n7684), .Z(n7714) );
  OR2_X1 U7670 ( .A1(n7715), .A2(n7660), .ZN(n7684) );
  OR2_X1 U7671 ( .A1(n7716), .A2(n7717), .ZN(n7685) );
  AND2_X1 U7672 ( .A1(n7718), .A2(n7719), .ZN(n7717) );
  AND2_X1 U7673 ( .A1(n7720), .A2(n7721), .ZN(n7716) );
  OR2_X1 U7674 ( .A1(n7719), .A2(n7718), .ZN(n7721) );
  XOR2_X1 U7675 ( .A(n7694), .B(n7722), .Z(n7686) );
  XOR2_X1 U7676 ( .A(n7693), .B(n7692), .Z(n7722) );
  OR2_X1 U7677 ( .A1(n7689), .A2(n7697), .ZN(n7692) );
  OR2_X1 U7678 ( .A1(n7723), .A2(n7724), .ZN(n7693) );
  AND2_X1 U7679 ( .A1(n7725), .A2(n7726), .ZN(n7724) );
  AND2_X1 U7680 ( .A1(n7727), .A2(n7728), .ZN(n7723) );
  OR2_X1 U7681 ( .A1(n7726), .A2(n7725), .ZN(n7728) );
  XOR2_X1 U7682 ( .A(n7702), .B(n7729), .Z(n7694) );
  XOR2_X1 U7683 ( .A(n7701), .B(n7700), .Z(n7729) );
  OR2_X1 U7684 ( .A1(n7659), .A2(n7730), .ZN(n7700) );
  OR2_X1 U7685 ( .A1(n7731), .A2(n7732), .ZN(n7701) );
  AND2_X1 U7686 ( .A1(n7733), .A2(n7734), .ZN(n7732) );
  AND2_X1 U7687 ( .A1(n7735), .A2(n7736), .ZN(n7731) );
  OR2_X1 U7688 ( .A1(n7733), .A2(n7734), .ZN(n7735) );
  XOR2_X1 U7689 ( .A(n7737), .B(n7738), .Z(n7702) );
  XOR2_X1 U7690 ( .A(n7739), .B(n7740), .Z(n7738) );
  OR2_X1 U7691 ( .A1(n7741), .A2(n7742), .ZN(n7337) );
  OR2_X1 U7692 ( .A1(n7743), .A2(n7336), .ZN(n7741) );
  AND2_X1 U7693 ( .A1(n7334), .A2(n7335), .ZN(n7336) );
  AND2_X1 U7694 ( .A1(n7744), .A2(n7745), .ZN(n7335) );
  INV_X1 U7695 ( .A(n7746), .ZN(n7744) );
  AND2_X1 U7696 ( .A1(n7330), .A2(n7334), .ZN(n7743) );
  INV_X1 U7697 ( .A(n7747), .ZN(n7334) );
  OR2_X1 U7698 ( .A1(n7748), .A2(n7742), .ZN(n7747) );
  INV_X1 U7699 ( .A(n7749), .ZN(n7742) );
  OR2_X1 U7700 ( .A1(n7750), .A2(n7751), .ZN(n7749) );
  AND2_X1 U7701 ( .A1(n7750), .A2(n7751), .ZN(n7748) );
  OR2_X1 U7702 ( .A1(n7752), .A2(n7753), .ZN(n7751) );
  AND2_X1 U7703 ( .A1(n7754), .A2(n7755), .ZN(n7753) );
  AND2_X1 U7704 ( .A1(n7756), .A2(n7757), .ZN(n7752) );
  OR2_X1 U7705 ( .A1(n7755), .A2(n7754), .ZN(n7757) );
  XOR2_X1 U7706 ( .A(n7712), .B(n7758), .Z(n7750) );
  XOR2_X1 U7707 ( .A(n7711), .B(n7710), .Z(n7758) );
  OR2_X1 U7708 ( .A1(n7759), .A2(n7660), .ZN(n7710) );
  OR2_X1 U7709 ( .A1(n7760), .A2(n7761), .ZN(n7711) );
  AND2_X1 U7710 ( .A1(n7762), .A2(n7763), .ZN(n7761) );
  AND2_X1 U7711 ( .A1(n7764), .A2(n7765), .ZN(n7760) );
  OR2_X1 U7712 ( .A1(n7763), .A2(n7762), .ZN(n7765) );
  XOR2_X1 U7713 ( .A(n7720), .B(n7766), .Z(n7712) );
  XOR2_X1 U7714 ( .A(n7719), .B(n7718), .Z(n7766) );
  OR2_X1 U7715 ( .A1(n7715), .A2(n7697), .ZN(n7718) );
  OR2_X1 U7716 ( .A1(n7767), .A2(n7768), .ZN(n7719) );
  AND2_X1 U7717 ( .A1(n7769), .A2(n7770), .ZN(n7768) );
  AND2_X1 U7718 ( .A1(n7771), .A2(n7772), .ZN(n7767) );
  OR2_X1 U7719 ( .A1(n7770), .A2(n7769), .ZN(n7772) );
  XOR2_X1 U7720 ( .A(n7727), .B(n7773), .Z(n7720) );
  XOR2_X1 U7721 ( .A(n7726), .B(n7725), .Z(n7773) );
  OR2_X1 U7722 ( .A1(n7689), .A2(n7730), .ZN(n7725) );
  OR2_X1 U7723 ( .A1(n7774), .A2(n7775), .ZN(n7726) );
  AND2_X1 U7724 ( .A1(n7776), .A2(n7777), .ZN(n7775) );
  AND2_X1 U7725 ( .A1(n7778), .A2(n7779), .ZN(n7774) );
  OR2_X1 U7726 ( .A1(n7777), .A2(n7776), .ZN(n7779) );
  XNOR2_X1 U7727 ( .A(n7780), .B(n7733), .ZN(n7727) );
  XOR2_X1 U7728 ( .A(n7781), .B(n7782), .Z(n7733) );
  XOR2_X1 U7729 ( .A(n7783), .B(n7784), .Z(n7782) );
  XNOR2_X1 U7730 ( .A(n7736), .B(n7734), .ZN(n7780) );
  OR2_X1 U7731 ( .A1(n7785), .A2(n7786), .ZN(n7734) );
  AND2_X1 U7732 ( .A1(n7787), .A2(n7788), .ZN(n7786) );
  AND2_X1 U7733 ( .A1(n7789), .A2(n7790), .ZN(n7785) );
  OR2_X1 U7734 ( .A1(n7788), .A2(n7787), .ZN(n7790) );
  AND2_X1 U7735 ( .A1(n7328), .A2(n7329), .ZN(n7330) );
  XNOR2_X1 U7736 ( .A(n7745), .B(n7746), .ZN(n7329) );
  OR2_X1 U7737 ( .A1(n7791), .A2(n7792), .ZN(n7746) );
  AND2_X1 U7738 ( .A1(n7793), .A2(n7794), .ZN(n7792) );
  AND2_X1 U7739 ( .A1(n7795), .A2(n7796), .ZN(n7791) );
  OR2_X1 U7740 ( .A1(n7794), .A2(n7793), .ZN(n7796) );
  XNOR2_X1 U7741 ( .A(n7756), .B(n7797), .ZN(n7745) );
  XOR2_X1 U7742 ( .A(n7755), .B(n7754), .Z(n7797) );
  OR2_X1 U7743 ( .A1(n7798), .A2(n7660), .ZN(n7754) );
  OR2_X1 U7744 ( .A1(n7799), .A2(n7800), .ZN(n7755) );
  AND2_X1 U7745 ( .A1(n7801), .A2(n7802), .ZN(n7800) );
  AND2_X1 U7746 ( .A1(n7803), .A2(n7804), .ZN(n7799) );
  OR2_X1 U7747 ( .A1(n7802), .A2(n7801), .ZN(n7804) );
  XOR2_X1 U7748 ( .A(n7764), .B(n7805), .Z(n7756) );
  XOR2_X1 U7749 ( .A(n7763), .B(n7762), .Z(n7805) );
  OR2_X1 U7750 ( .A1(n7759), .A2(n7697), .ZN(n7762) );
  OR2_X1 U7751 ( .A1(n7806), .A2(n7807), .ZN(n7763) );
  AND2_X1 U7752 ( .A1(n7808), .A2(n7809), .ZN(n7807) );
  AND2_X1 U7753 ( .A1(n7810), .A2(n7811), .ZN(n7806) );
  OR2_X1 U7754 ( .A1(n7809), .A2(n7808), .ZN(n7811) );
  XOR2_X1 U7755 ( .A(n7771), .B(n7812), .Z(n7764) );
  XOR2_X1 U7756 ( .A(n7770), .B(n7769), .Z(n7812) );
  OR2_X1 U7757 ( .A1(n7715), .A2(n7730), .ZN(n7769) );
  OR2_X1 U7758 ( .A1(n7813), .A2(n7814), .ZN(n7770) );
  AND2_X1 U7759 ( .A1(n7815), .A2(n7816), .ZN(n7814) );
  AND2_X1 U7760 ( .A1(n7817), .A2(n7818), .ZN(n7813) );
  OR2_X1 U7761 ( .A1(n7816), .A2(n7815), .ZN(n7818) );
  XOR2_X1 U7762 ( .A(n7778), .B(n7819), .Z(n7771) );
  XOR2_X1 U7763 ( .A(n7777), .B(n7776), .Z(n7819) );
  OR2_X1 U7764 ( .A1(n7689), .A2(n7820), .ZN(n7776) );
  OR2_X1 U7765 ( .A1(n7821), .A2(n7822), .ZN(n7777) );
  AND2_X1 U7766 ( .A1(n7823), .A2(n7824), .ZN(n7822) );
  AND2_X1 U7767 ( .A1(n7825), .A2(n7826), .ZN(n7821) );
  OR2_X1 U7768 ( .A1(n7823), .A2(n7824), .ZN(n7825) );
  XOR2_X1 U7769 ( .A(n7789), .B(n7827), .Z(n7778) );
  XOR2_X1 U7770 ( .A(n7788), .B(n7787), .Z(n7827) );
  OR2_X1 U7771 ( .A1(n7659), .A2(n7828), .ZN(n7787) );
  OR2_X1 U7772 ( .A1(n7829), .A2(n7830), .ZN(n7788) );
  AND2_X1 U7773 ( .A1(n7831), .A2(n7832), .ZN(n7830) );
  AND2_X1 U7774 ( .A1(n7833), .A2(n7834), .ZN(n7829) );
  OR2_X1 U7775 ( .A1(n7832), .A2(n7831), .ZN(n7834) );
  XOR2_X1 U7776 ( .A(n7835), .B(n7836), .Z(n7789) );
  XOR2_X1 U7777 ( .A(n7837), .B(n7838), .Z(n7836) );
  OR2_X1 U7778 ( .A1(n7839), .A2(n7840), .ZN(n7328) );
  OR2_X1 U7779 ( .A1(n7841), .A2(n7327), .ZN(n7839) );
  AND2_X1 U7780 ( .A1(n7325), .A2(n7326), .ZN(n7327) );
  AND2_X1 U7781 ( .A1(n7842), .A2(n7843), .ZN(n7326) );
  INV_X1 U7782 ( .A(n7844), .ZN(n7842) );
  AND2_X1 U7783 ( .A1(n7321), .A2(n7325), .ZN(n7841) );
  INV_X1 U7784 ( .A(n7845), .ZN(n7325) );
  OR2_X1 U7785 ( .A1(n7846), .A2(n7840), .ZN(n7845) );
  INV_X1 U7786 ( .A(n7847), .ZN(n7840) );
  OR2_X1 U7787 ( .A1(n7848), .A2(n7849), .ZN(n7847) );
  AND2_X1 U7788 ( .A1(n7848), .A2(n7849), .ZN(n7846) );
  OR2_X1 U7789 ( .A1(n7850), .A2(n7851), .ZN(n7849) );
  AND2_X1 U7790 ( .A1(n7852), .A2(n7853), .ZN(n7851) );
  AND2_X1 U7791 ( .A1(n7854), .A2(n7855), .ZN(n7850) );
  OR2_X1 U7792 ( .A1(n7853), .A2(n7852), .ZN(n7855) );
  XOR2_X1 U7793 ( .A(n7795), .B(n7856), .Z(n7848) );
  XOR2_X1 U7794 ( .A(n7794), .B(n7793), .Z(n7856) );
  OR2_X1 U7795 ( .A1(n7857), .A2(n7660), .ZN(n7793) );
  OR2_X1 U7796 ( .A1(n7858), .A2(n7859), .ZN(n7794) );
  AND2_X1 U7797 ( .A1(n7860), .A2(n7861), .ZN(n7859) );
  AND2_X1 U7798 ( .A1(n7862), .A2(n7863), .ZN(n7858) );
  OR2_X1 U7799 ( .A1(n7861), .A2(n7860), .ZN(n7863) );
  XOR2_X1 U7800 ( .A(n7803), .B(n7864), .Z(n7795) );
  XOR2_X1 U7801 ( .A(n7802), .B(n7801), .Z(n7864) );
  OR2_X1 U7802 ( .A1(n7798), .A2(n7697), .ZN(n7801) );
  OR2_X1 U7803 ( .A1(n7865), .A2(n7866), .ZN(n7802) );
  AND2_X1 U7804 ( .A1(n7867), .A2(n7868), .ZN(n7866) );
  AND2_X1 U7805 ( .A1(n7869), .A2(n7870), .ZN(n7865) );
  OR2_X1 U7806 ( .A1(n7868), .A2(n7867), .ZN(n7870) );
  XOR2_X1 U7807 ( .A(n7810), .B(n7871), .Z(n7803) );
  XOR2_X1 U7808 ( .A(n7809), .B(n7808), .Z(n7871) );
  OR2_X1 U7809 ( .A1(n7759), .A2(n7730), .ZN(n7808) );
  OR2_X1 U7810 ( .A1(n7872), .A2(n7873), .ZN(n7809) );
  AND2_X1 U7811 ( .A1(n7874), .A2(n7875), .ZN(n7873) );
  AND2_X1 U7812 ( .A1(n7876), .A2(n7877), .ZN(n7872) );
  OR2_X1 U7813 ( .A1(n7875), .A2(n7874), .ZN(n7877) );
  XOR2_X1 U7814 ( .A(n7817), .B(n7878), .Z(n7810) );
  XOR2_X1 U7815 ( .A(n7816), .B(n7815), .Z(n7878) );
  OR2_X1 U7816 ( .A1(n7715), .A2(n7820), .ZN(n7815) );
  OR2_X1 U7817 ( .A1(n7879), .A2(n7880), .ZN(n7816) );
  AND2_X1 U7818 ( .A1(n7881), .A2(n7882), .ZN(n7880) );
  AND2_X1 U7819 ( .A1(n7883), .A2(n7884), .ZN(n7879) );
  OR2_X1 U7820 ( .A1(n7882), .A2(n7881), .ZN(n7884) );
  XNOR2_X1 U7821 ( .A(n7885), .B(n7823), .ZN(n7817) );
  XOR2_X1 U7822 ( .A(n7833), .B(n7886), .Z(n7823) );
  XOR2_X1 U7823 ( .A(n7832), .B(n7831), .Z(n7886) );
  OR2_X1 U7824 ( .A1(n7659), .A2(n7887), .ZN(n7831) );
  OR2_X1 U7825 ( .A1(n7888), .A2(n7889), .ZN(n7832) );
  AND2_X1 U7826 ( .A1(n7890), .A2(n7891), .ZN(n7889) );
  AND2_X1 U7827 ( .A1(n7892), .A2(n7893), .ZN(n7888) );
  OR2_X1 U7828 ( .A1(n7891), .A2(n7890), .ZN(n7893) );
  XOR2_X1 U7829 ( .A(n7894), .B(n7895), .Z(n7833) );
  XOR2_X1 U7830 ( .A(n7896), .B(n7897), .Z(n7895) );
  XNOR2_X1 U7831 ( .A(n7826), .B(n7824), .ZN(n7885) );
  OR2_X1 U7832 ( .A1(n7898), .A2(n7899), .ZN(n7824) );
  AND2_X1 U7833 ( .A1(n7900), .A2(n7901), .ZN(n7899) );
  AND2_X1 U7834 ( .A1(n7902), .A2(n7903), .ZN(n7898) );
  OR2_X1 U7835 ( .A1(n7901), .A2(n7900), .ZN(n7903) );
  AND2_X1 U7836 ( .A1(n7904), .A2(n7626), .ZN(n7321) );
  INV_X1 U7837 ( .A(n7621), .ZN(n7626) );
  XOR2_X1 U7838 ( .A(n7843), .B(n7844), .Z(n7621) );
  OR2_X1 U7839 ( .A1(n7905), .A2(n7906), .ZN(n7844) );
  AND2_X1 U7840 ( .A1(n7907), .A2(n7908), .ZN(n7906) );
  AND2_X1 U7841 ( .A1(n7909), .A2(n7910), .ZN(n7905) );
  OR2_X1 U7842 ( .A1(n7908), .A2(n7907), .ZN(n7910) );
  XNOR2_X1 U7843 ( .A(n7854), .B(n7911), .ZN(n7843) );
  XOR2_X1 U7844 ( .A(n7853), .B(n7852), .Z(n7911) );
  OR2_X1 U7845 ( .A1(n7912), .A2(n7660), .ZN(n7852) );
  OR2_X1 U7846 ( .A1(n7913), .A2(n7914), .ZN(n7853) );
  AND2_X1 U7847 ( .A1(n7915), .A2(n7916), .ZN(n7914) );
  AND2_X1 U7848 ( .A1(n7917), .A2(n7918), .ZN(n7913) );
  OR2_X1 U7849 ( .A1(n7916), .A2(n7915), .ZN(n7918) );
  XOR2_X1 U7850 ( .A(n7862), .B(n7919), .Z(n7854) );
  XOR2_X1 U7851 ( .A(n7861), .B(n7860), .Z(n7919) );
  OR2_X1 U7852 ( .A1(n7857), .A2(n7697), .ZN(n7860) );
  OR2_X1 U7853 ( .A1(n7920), .A2(n7921), .ZN(n7861) );
  AND2_X1 U7854 ( .A1(n7922), .A2(n7923), .ZN(n7921) );
  AND2_X1 U7855 ( .A1(n7924), .A2(n7925), .ZN(n7920) );
  OR2_X1 U7856 ( .A1(n7923), .A2(n7922), .ZN(n7925) );
  XOR2_X1 U7857 ( .A(n7869), .B(n7926), .Z(n7862) );
  XOR2_X1 U7858 ( .A(n7868), .B(n7867), .Z(n7926) );
  OR2_X1 U7859 ( .A1(n7798), .A2(n7730), .ZN(n7867) );
  OR2_X1 U7860 ( .A1(n7927), .A2(n7928), .ZN(n7868) );
  AND2_X1 U7861 ( .A1(n7929), .A2(n7930), .ZN(n7928) );
  AND2_X1 U7862 ( .A1(n7931), .A2(n7932), .ZN(n7927) );
  OR2_X1 U7863 ( .A1(n7930), .A2(n7929), .ZN(n7932) );
  XOR2_X1 U7864 ( .A(n7876), .B(n7933), .Z(n7869) );
  XOR2_X1 U7865 ( .A(n7875), .B(n7874), .Z(n7933) );
  OR2_X1 U7866 ( .A1(n7759), .A2(n7820), .ZN(n7874) );
  OR2_X1 U7867 ( .A1(n7934), .A2(n7935), .ZN(n7875) );
  AND2_X1 U7868 ( .A1(n7936), .A2(n7937), .ZN(n7935) );
  AND2_X1 U7869 ( .A1(n7938), .A2(n7939), .ZN(n7934) );
  OR2_X1 U7870 ( .A1(n7937), .A2(n7936), .ZN(n7939) );
  XOR2_X1 U7871 ( .A(n7883), .B(n7940), .Z(n7876) );
  XOR2_X1 U7872 ( .A(n7882), .B(n7881), .Z(n7940) );
  OR2_X1 U7873 ( .A1(n7715), .A2(n7828), .ZN(n7881) );
  OR2_X1 U7874 ( .A1(n7941), .A2(n7942), .ZN(n7882) );
  AND2_X1 U7875 ( .A1(n7943), .A2(n7944), .ZN(n7942) );
  AND2_X1 U7876 ( .A1(n7945), .A2(n7946), .ZN(n7941) );
  OR2_X1 U7877 ( .A1(n7943), .A2(n7944), .ZN(n7945) );
  XOR2_X1 U7878 ( .A(n7902), .B(n7947), .Z(n7883) );
  XOR2_X1 U7879 ( .A(n7901), .B(n7900), .Z(n7947) );
  OR2_X1 U7880 ( .A1(n7689), .A2(n7887), .ZN(n7900) );
  OR2_X1 U7881 ( .A1(n7948), .A2(n7949), .ZN(n7901) );
  AND2_X1 U7882 ( .A1(n7950), .A2(n7951), .ZN(n7949) );
  AND2_X1 U7883 ( .A1(n7952), .A2(n7953), .ZN(n7948) );
  OR2_X1 U7884 ( .A1(n7951), .A2(n7950), .ZN(n7953) );
  XOR2_X1 U7885 ( .A(n7892), .B(n7954), .Z(n7902) );
  XOR2_X1 U7886 ( .A(n7891), .B(n7890), .Z(n7954) );
  OR2_X1 U7887 ( .A1(n7659), .A2(n7955), .ZN(n7890) );
  OR2_X1 U7888 ( .A1(n7956), .A2(n7957), .ZN(n7891) );
  AND2_X1 U7889 ( .A1(n7958), .A2(n7959), .ZN(n7957) );
  AND2_X1 U7890 ( .A1(n7960), .A2(n7961), .ZN(n7956) );
  OR2_X1 U7891 ( .A1(n7959), .A2(n7958), .ZN(n7961) );
  XOR2_X1 U7892 ( .A(n7962), .B(n7963), .Z(n7892) );
  XOR2_X1 U7893 ( .A(n7964), .B(n7965), .Z(n7963) );
  OR2_X1 U7894 ( .A1(n7624), .A2(n7625), .ZN(n7904) );
  OR2_X1 U7895 ( .A1(n7966), .A2(n7614), .ZN(n7624) );
  AND2_X1 U7896 ( .A1(n7612), .A2(n7613), .ZN(n7614) );
  AND2_X1 U7897 ( .A1(n7967), .A2(n7968), .ZN(n7613) );
  INV_X1 U7898 ( .A(n7969), .ZN(n7967) );
  AND2_X1 U7899 ( .A1(n7608), .A2(n7612), .ZN(n7966) );
  INV_X1 U7900 ( .A(n7970), .ZN(n7612) );
  OR2_X1 U7901 ( .A1(n7971), .A2(n7625), .ZN(n7970) );
  INV_X1 U7902 ( .A(n7622), .ZN(n7625) );
  OR2_X1 U7903 ( .A1(n7972), .A2(n7973), .ZN(n7622) );
  AND2_X1 U7904 ( .A1(n7972), .A2(n7973), .ZN(n7971) );
  OR2_X1 U7905 ( .A1(n7974), .A2(n7975), .ZN(n7973) );
  AND2_X1 U7906 ( .A1(n7976), .A2(n7977), .ZN(n7975) );
  AND2_X1 U7907 ( .A1(n7978), .A2(n7979), .ZN(n7974) );
  OR2_X1 U7908 ( .A1(n7976), .A2(n7977), .ZN(n7979) );
  XOR2_X1 U7909 ( .A(n7909), .B(n7980), .Z(n7972) );
  XOR2_X1 U7910 ( .A(n7908), .B(n7907), .Z(n7980) );
  OR2_X1 U7911 ( .A1(n7981), .A2(n7660), .ZN(n7907) );
  OR2_X1 U7912 ( .A1(n7982), .A2(n7983), .ZN(n7908) );
  AND2_X1 U7913 ( .A1(n7984), .A2(n7985), .ZN(n7983) );
  AND2_X1 U7914 ( .A1(n7986), .A2(n7987), .ZN(n7982) );
  OR2_X1 U7915 ( .A1(n7985), .A2(n7984), .ZN(n7987) );
  XOR2_X1 U7916 ( .A(n7917), .B(n7988), .Z(n7909) );
  XOR2_X1 U7917 ( .A(n7916), .B(n7915), .Z(n7988) );
  OR2_X1 U7918 ( .A1(n7912), .A2(n7697), .ZN(n7915) );
  OR2_X1 U7919 ( .A1(n7989), .A2(n7990), .ZN(n7916) );
  AND2_X1 U7920 ( .A1(n7991), .A2(n7992), .ZN(n7990) );
  AND2_X1 U7921 ( .A1(n7993), .A2(n7994), .ZN(n7989) );
  OR2_X1 U7922 ( .A1(n7992), .A2(n7991), .ZN(n7994) );
  XOR2_X1 U7923 ( .A(n7924), .B(n7995), .Z(n7917) );
  XOR2_X1 U7924 ( .A(n7923), .B(n7922), .Z(n7995) );
  OR2_X1 U7925 ( .A1(n7857), .A2(n7730), .ZN(n7922) );
  OR2_X1 U7926 ( .A1(n7996), .A2(n7997), .ZN(n7923) );
  AND2_X1 U7927 ( .A1(n7998), .A2(n7999), .ZN(n7997) );
  AND2_X1 U7928 ( .A1(n8000), .A2(n8001), .ZN(n7996) );
  OR2_X1 U7929 ( .A1(n7999), .A2(n7998), .ZN(n8001) );
  XOR2_X1 U7930 ( .A(n7931), .B(n8002), .Z(n7924) );
  XOR2_X1 U7931 ( .A(n7930), .B(n7929), .Z(n8002) );
  OR2_X1 U7932 ( .A1(n7798), .A2(n7820), .ZN(n7929) );
  OR2_X1 U7933 ( .A1(n8003), .A2(n8004), .ZN(n7930) );
  AND2_X1 U7934 ( .A1(n8005), .A2(n8006), .ZN(n8004) );
  AND2_X1 U7935 ( .A1(n8007), .A2(n8008), .ZN(n8003) );
  OR2_X1 U7936 ( .A1(n8006), .A2(n8005), .ZN(n8008) );
  XOR2_X1 U7937 ( .A(n7938), .B(n8009), .Z(n7931) );
  XOR2_X1 U7938 ( .A(n7937), .B(n7936), .Z(n8009) );
  OR2_X1 U7939 ( .A1(n7759), .A2(n7828), .ZN(n7936) );
  OR2_X1 U7940 ( .A1(n8010), .A2(n8011), .ZN(n7937) );
  AND2_X1 U7941 ( .A1(n8012), .A2(n8013), .ZN(n8011) );
  AND2_X1 U7942 ( .A1(n8014), .A2(n8015), .ZN(n8010) );
  OR2_X1 U7943 ( .A1(n8013), .A2(n8012), .ZN(n8015) );
  XNOR2_X1 U7944 ( .A(n8016), .B(n7943), .ZN(n7938) );
  XOR2_X1 U7945 ( .A(n7952), .B(n8017), .Z(n7943) );
  XOR2_X1 U7946 ( .A(n7951), .B(n7950), .Z(n8017) );
  OR2_X1 U7947 ( .A1(n7689), .A2(n7955), .ZN(n7950) );
  OR2_X1 U7948 ( .A1(n8018), .A2(n8019), .ZN(n7951) );
  AND2_X1 U7949 ( .A1(n8020), .A2(n8021), .ZN(n8019) );
  AND2_X1 U7950 ( .A1(n8022), .A2(n8023), .ZN(n8018) );
  OR2_X1 U7951 ( .A1(n8021), .A2(n8020), .ZN(n8023) );
  XOR2_X1 U7952 ( .A(n7960), .B(n8024), .Z(n7952) );
  XOR2_X1 U7953 ( .A(n7959), .B(n7958), .Z(n8024) );
  OR2_X1 U7954 ( .A1(n7659), .A2(n8025), .ZN(n7958) );
  OR2_X1 U7955 ( .A1(n8026), .A2(n8027), .ZN(n7959) );
  AND2_X1 U7956 ( .A1(n8028), .A2(n8029), .ZN(n8027) );
  AND2_X1 U7957 ( .A1(n8030), .A2(n8031), .ZN(n8026) );
  OR2_X1 U7958 ( .A1(n8029), .A2(n8028), .ZN(n8031) );
  XOR2_X1 U7959 ( .A(n8032), .B(n8033), .Z(n7960) );
  XOR2_X1 U7960 ( .A(n8034), .B(n8035), .Z(n8033) );
  XNOR2_X1 U7961 ( .A(n7946), .B(n7944), .ZN(n8016) );
  OR2_X1 U7962 ( .A1(n8036), .A2(n8037), .ZN(n7944) );
  AND2_X1 U7963 ( .A1(n8038), .A2(n8039), .ZN(n8037) );
  AND2_X1 U7964 ( .A1(n8040), .A2(n8041), .ZN(n8036) );
  OR2_X1 U7965 ( .A1(n8039), .A2(n8038), .ZN(n8041) );
  AND2_X1 U7966 ( .A1(n8042), .A2(n7607), .ZN(n7608) );
  INV_X1 U7967 ( .A(n7602), .ZN(n7607) );
  XOR2_X1 U7968 ( .A(n7968), .B(n7969), .Z(n7602) );
  OR2_X1 U7969 ( .A1(n8043), .A2(n8044), .ZN(n7969) );
  AND2_X1 U7970 ( .A1(n8045), .A2(n8046), .ZN(n8044) );
  AND2_X1 U7971 ( .A1(n8047), .A2(n8048), .ZN(n8043) );
  OR2_X1 U7972 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  XNOR2_X1 U7973 ( .A(n7978), .B(n8049), .ZN(n7968) );
  XOR2_X1 U7974 ( .A(n7977), .B(n7976), .Z(n8049) );
  OR2_X1 U7975 ( .A1(n8050), .A2(n7660), .ZN(n7976) );
  OR2_X1 U7976 ( .A1(n8051), .A2(n8052), .ZN(n7977) );
  AND2_X1 U7977 ( .A1(n8053), .A2(n8054), .ZN(n8052) );
  AND2_X1 U7978 ( .A1(n8055), .A2(n8056), .ZN(n8051) );
  OR2_X1 U7979 ( .A1(n8053), .A2(n8054), .ZN(n8056) );
  XOR2_X1 U7980 ( .A(n7986), .B(n8057), .Z(n7978) );
  XOR2_X1 U7981 ( .A(n7985), .B(n7984), .Z(n8057) );
  OR2_X1 U7982 ( .A1(n7981), .A2(n7697), .ZN(n7984) );
  OR2_X1 U7983 ( .A1(n8058), .A2(n8059), .ZN(n7985) );
  AND2_X1 U7984 ( .A1(n8060), .A2(n8061), .ZN(n8059) );
  AND2_X1 U7985 ( .A1(n8062), .A2(n8063), .ZN(n8058) );
  OR2_X1 U7986 ( .A1(n8061), .A2(n8060), .ZN(n8063) );
  XOR2_X1 U7987 ( .A(n7993), .B(n8064), .Z(n7986) );
  XOR2_X1 U7988 ( .A(n7992), .B(n7991), .Z(n8064) );
  OR2_X1 U7989 ( .A1(n7912), .A2(n7730), .ZN(n7991) );
  OR2_X1 U7990 ( .A1(n8065), .A2(n8066), .ZN(n7992) );
  AND2_X1 U7991 ( .A1(n8067), .A2(n8068), .ZN(n8066) );
  AND2_X1 U7992 ( .A1(n8069), .A2(n8070), .ZN(n8065) );
  OR2_X1 U7993 ( .A1(n8068), .A2(n8067), .ZN(n8070) );
  XOR2_X1 U7994 ( .A(n8000), .B(n8071), .Z(n7993) );
  XOR2_X1 U7995 ( .A(n7999), .B(n7998), .Z(n8071) );
  OR2_X1 U7996 ( .A1(n7857), .A2(n7820), .ZN(n7998) );
  OR2_X1 U7997 ( .A1(n8072), .A2(n8073), .ZN(n7999) );
  AND2_X1 U7998 ( .A1(n8074), .A2(n8075), .ZN(n8073) );
  AND2_X1 U7999 ( .A1(n8076), .A2(n8077), .ZN(n8072) );
  OR2_X1 U8000 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  XOR2_X1 U8001 ( .A(n8007), .B(n8078), .Z(n8000) );
  XOR2_X1 U8002 ( .A(n8006), .B(n8005), .Z(n8078) );
  OR2_X1 U8003 ( .A1(n7798), .A2(n7828), .ZN(n8005) );
  OR2_X1 U8004 ( .A1(n8079), .A2(n8080), .ZN(n8006) );
  AND2_X1 U8005 ( .A1(n8081), .A2(n8082), .ZN(n8080) );
  AND2_X1 U8006 ( .A1(n8083), .A2(n8084), .ZN(n8079) );
  OR2_X1 U8007 ( .A1(n8082), .A2(n8081), .ZN(n8084) );
  XOR2_X1 U8008 ( .A(n8014), .B(n8085), .Z(n8007) );
  XOR2_X1 U8009 ( .A(n8013), .B(n8012), .Z(n8085) );
  OR2_X1 U8010 ( .A1(n7759), .A2(n7887), .ZN(n8012) );
  OR2_X1 U8011 ( .A1(n8086), .A2(n8087), .ZN(n8013) );
  AND2_X1 U8012 ( .A1(n8088), .A2(n8089), .ZN(n8087) );
  AND2_X1 U8013 ( .A1(n8090), .A2(n8091), .ZN(n8086) );
  OR2_X1 U8014 ( .A1(n8088), .A2(n8089), .ZN(n8090) );
  XOR2_X1 U8015 ( .A(n8040), .B(n8092), .Z(n8014) );
  XOR2_X1 U8016 ( .A(n8039), .B(n8038), .Z(n8092) );
  OR2_X1 U8017 ( .A1(n7715), .A2(n7955), .ZN(n8038) );
  OR2_X1 U8018 ( .A1(n8093), .A2(n8094), .ZN(n8039) );
  AND2_X1 U8019 ( .A1(n8095), .A2(n8096), .ZN(n8094) );
  AND2_X1 U8020 ( .A1(n8097), .A2(n8098), .ZN(n8093) );
  OR2_X1 U8021 ( .A1(n8096), .A2(n8095), .ZN(n8098) );
  XOR2_X1 U8022 ( .A(n8022), .B(n8099), .Z(n8040) );
  XOR2_X1 U8023 ( .A(n8021), .B(n8020), .Z(n8099) );
  OR2_X1 U8024 ( .A1(n7689), .A2(n8025), .ZN(n8020) );
  OR2_X1 U8025 ( .A1(n8100), .A2(n8101), .ZN(n8021) );
  AND2_X1 U8026 ( .A1(n8102), .A2(n8103), .ZN(n8101) );
  AND2_X1 U8027 ( .A1(n8104), .A2(n8105), .ZN(n8100) );
  OR2_X1 U8028 ( .A1(n8103), .A2(n8102), .ZN(n8105) );
  XOR2_X1 U8029 ( .A(n8030), .B(n8106), .Z(n8022) );
  XOR2_X1 U8030 ( .A(n8029), .B(n8028), .Z(n8106) );
  OR2_X1 U8031 ( .A1(n7659), .A2(n8107), .ZN(n8028) );
  OR2_X1 U8032 ( .A1(n8108), .A2(n8109), .ZN(n8029) );
  AND2_X1 U8033 ( .A1(n8110), .A2(n8111), .ZN(n8109) );
  AND2_X1 U8034 ( .A1(n8112), .A2(n8113), .ZN(n8108) );
  OR2_X1 U8035 ( .A1(n8111), .A2(n8110), .ZN(n8113) );
  XOR2_X1 U8036 ( .A(n8114), .B(n8115), .Z(n8030) );
  XOR2_X1 U8037 ( .A(n8116), .B(n8117), .Z(n8115) );
  OR2_X1 U8038 ( .A1(n7605), .A2(n7606), .ZN(n8042) );
  OR2_X1 U8039 ( .A1(n8118), .A2(n7595), .ZN(n7605) );
  AND2_X1 U8040 ( .A1(n7593), .A2(n7594), .ZN(n7595) );
  AND2_X1 U8041 ( .A1(n8119), .A2(n8120), .ZN(n7594) );
  INV_X1 U8042 ( .A(n8121), .ZN(n8119) );
  AND2_X1 U8043 ( .A1(n7589), .A2(n7593), .ZN(n8118) );
  INV_X1 U8044 ( .A(n8122), .ZN(n7593) );
  OR2_X1 U8045 ( .A1(n8123), .A2(n7606), .ZN(n8122) );
  INV_X1 U8046 ( .A(n7603), .ZN(n7606) );
  OR2_X1 U8047 ( .A1(n8124), .A2(n8125), .ZN(n7603) );
  AND2_X1 U8048 ( .A1(n8124), .A2(n8125), .ZN(n8123) );
  OR2_X1 U8049 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  AND2_X1 U8050 ( .A1(n8128), .A2(n8129), .ZN(n8127) );
  AND2_X1 U8051 ( .A1(n8130), .A2(n8131), .ZN(n8126) );
  OR2_X1 U8052 ( .A1(n8128), .A2(n8129), .ZN(n8131) );
  XOR2_X1 U8053 ( .A(n8047), .B(n8132), .Z(n8124) );
  XOR2_X1 U8054 ( .A(n8046), .B(n8045), .Z(n8132) );
  OR2_X1 U8055 ( .A1(n7660), .A2(n8133), .ZN(n8045) );
  OR2_X1 U8056 ( .A1(n8134), .A2(n8135), .ZN(n8046) );
  AND2_X1 U8057 ( .A1(n8136), .A2(n8137), .ZN(n8135) );
  AND2_X1 U8058 ( .A1(n8138), .A2(n8139), .ZN(n8134) );
  OR2_X1 U8059 ( .A1(n8137), .A2(n8136), .ZN(n8139) );
  XOR2_X1 U8060 ( .A(n8055), .B(n8140), .Z(n8047) );
  XOR2_X1 U8061 ( .A(n8054), .B(n8053), .Z(n8140) );
  OR2_X1 U8062 ( .A1(n8050), .A2(n7697), .ZN(n8053) );
  OR2_X1 U8063 ( .A1(n8141), .A2(n8142), .ZN(n8054) );
  AND2_X1 U8064 ( .A1(n8143), .A2(n8144), .ZN(n8142) );
  AND2_X1 U8065 ( .A1(n8145), .A2(n8146), .ZN(n8141) );
  OR2_X1 U8066 ( .A1(n8143), .A2(n8144), .ZN(n8146) );
  XOR2_X1 U8067 ( .A(n8062), .B(n8147), .Z(n8055) );
  XOR2_X1 U8068 ( .A(n8061), .B(n8060), .Z(n8147) );
  OR2_X1 U8069 ( .A1(n7981), .A2(n7730), .ZN(n8060) );
  OR2_X1 U8070 ( .A1(n8148), .A2(n8149), .ZN(n8061) );
  AND2_X1 U8071 ( .A1(n8150), .A2(n8151), .ZN(n8149) );
  AND2_X1 U8072 ( .A1(n8152), .A2(n8153), .ZN(n8148) );
  OR2_X1 U8073 ( .A1(n8151), .A2(n8150), .ZN(n8153) );
  XOR2_X1 U8074 ( .A(n8069), .B(n8154), .Z(n8062) );
  XOR2_X1 U8075 ( .A(n8068), .B(n8067), .Z(n8154) );
  OR2_X1 U8076 ( .A1(n7912), .A2(n7820), .ZN(n8067) );
  OR2_X1 U8077 ( .A1(n8155), .A2(n8156), .ZN(n8068) );
  AND2_X1 U8078 ( .A1(n8157), .A2(n8158), .ZN(n8156) );
  AND2_X1 U8079 ( .A1(n8159), .A2(n8160), .ZN(n8155) );
  OR2_X1 U8080 ( .A1(n8158), .A2(n8157), .ZN(n8160) );
  XOR2_X1 U8081 ( .A(n8076), .B(n8161), .Z(n8069) );
  XOR2_X1 U8082 ( .A(n8075), .B(n8074), .Z(n8161) );
  OR2_X1 U8083 ( .A1(n7857), .A2(n7828), .ZN(n8074) );
  OR2_X1 U8084 ( .A1(n8162), .A2(n8163), .ZN(n8075) );
  AND2_X1 U8085 ( .A1(n8164), .A2(n8165), .ZN(n8163) );
  AND2_X1 U8086 ( .A1(n8166), .A2(n8167), .ZN(n8162) );
  OR2_X1 U8087 ( .A1(n8165), .A2(n8164), .ZN(n8167) );
  XOR2_X1 U8088 ( .A(n8083), .B(n8168), .Z(n8076) );
  XOR2_X1 U8089 ( .A(n8082), .B(n8081), .Z(n8168) );
  OR2_X1 U8090 ( .A1(n7798), .A2(n7887), .ZN(n8081) );
  OR2_X1 U8091 ( .A1(n8169), .A2(n8170), .ZN(n8082) );
  AND2_X1 U8092 ( .A1(n8171), .A2(n8172), .ZN(n8170) );
  AND2_X1 U8093 ( .A1(n8173), .A2(n8174), .ZN(n8169) );
  OR2_X1 U8094 ( .A1(n8172), .A2(n8171), .ZN(n8174) );
  XNOR2_X1 U8095 ( .A(n8175), .B(n8088), .ZN(n8083) );
  XOR2_X1 U8096 ( .A(n8097), .B(n8176), .Z(n8088) );
  XOR2_X1 U8097 ( .A(n8096), .B(n8095), .Z(n8176) );
  OR2_X1 U8098 ( .A1(n7715), .A2(n8025), .ZN(n8095) );
  OR2_X1 U8099 ( .A1(n8177), .A2(n8178), .ZN(n8096) );
  AND2_X1 U8100 ( .A1(n8179), .A2(n8180), .ZN(n8178) );
  AND2_X1 U8101 ( .A1(n8181), .A2(n8182), .ZN(n8177) );
  OR2_X1 U8102 ( .A1(n8180), .A2(n8179), .ZN(n8182) );
  XOR2_X1 U8103 ( .A(n8104), .B(n8183), .Z(n8097) );
  XOR2_X1 U8104 ( .A(n8103), .B(n8102), .Z(n8183) );
  OR2_X1 U8105 ( .A1(n7689), .A2(n8107), .ZN(n8102) );
  OR2_X1 U8106 ( .A1(n8184), .A2(n8185), .ZN(n8103) );
  AND2_X1 U8107 ( .A1(n8186), .A2(n8187), .ZN(n8185) );
  AND2_X1 U8108 ( .A1(n8188), .A2(n8189), .ZN(n8184) );
  OR2_X1 U8109 ( .A1(n8187), .A2(n8186), .ZN(n8189) );
  XOR2_X1 U8110 ( .A(n8112), .B(n8190), .Z(n8104) );
  XOR2_X1 U8111 ( .A(n8111), .B(n8110), .Z(n8190) );
  OR2_X1 U8112 ( .A1(n7659), .A2(n8191), .ZN(n8110) );
  OR2_X1 U8113 ( .A1(n8192), .A2(n8193), .ZN(n8111) );
  AND2_X1 U8114 ( .A1(n8194), .A2(n8195), .ZN(n8193) );
  AND2_X1 U8115 ( .A1(n8196), .A2(n8197), .ZN(n8192) );
  OR2_X1 U8116 ( .A1(n8195), .A2(n8194), .ZN(n8197) );
  XOR2_X1 U8117 ( .A(n8198), .B(n8199), .Z(n8112) );
  XOR2_X1 U8118 ( .A(n8200), .B(n8201), .Z(n8199) );
  XNOR2_X1 U8119 ( .A(n8091), .B(n8089), .ZN(n8175) );
  OR2_X1 U8120 ( .A1(n8202), .A2(n8203), .ZN(n8089) );
  AND2_X1 U8121 ( .A1(n8204), .A2(n8205), .ZN(n8203) );
  AND2_X1 U8122 ( .A1(n8206), .A2(n8207), .ZN(n8202) );
  OR2_X1 U8123 ( .A1(n8205), .A2(n8204), .ZN(n8207) );
  AND2_X1 U8124 ( .A1(n8208), .A2(n7588), .ZN(n7589) );
  INV_X1 U8125 ( .A(n7583), .ZN(n7588) );
  XOR2_X1 U8126 ( .A(n8120), .B(n8121), .Z(n7583) );
  OR2_X1 U8127 ( .A1(n8209), .A2(n8210), .ZN(n8121) );
  AND2_X1 U8128 ( .A1(n8211), .A2(n8212), .ZN(n8210) );
  AND2_X1 U8129 ( .A1(n8213), .A2(n8214), .ZN(n8209) );
  OR2_X1 U8130 ( .A1(n8212), .A2(n8211), .ZN(n8214) );
  XNOR2_X1 U8131 ( .A(n8130), .B(n8215), .ZN(n8120) );
  XOR2_X1 U8132 ( .A(n8129), .B(n8128), .Z(n8215) );
  OR2_X1 U8133 ( .A1(n7660), .A2(n8216), .ZN(n8128) );
  OR2_X1 U8134 ( .A1(n8217), .A2(n8218), .ZN(n8129) );
  AND2_X1 U8135 ( .A1(n8219), .A2(n8220), .ZN(n8218) );
  AND2_X1 U8136 ( .A1(n8221), .A2(n8222), .ZN(n8217) );
  OR2_X1 U8137 ( .A1(n8219), .A2(n8220), .ZN(n8222) );
  XOR2_X1 U8138 ( .A(n8138), .B(n8223), .Z(n8130) );
  XOR2_X1 U8139 ( .A(n8137), .B(n8136), .Z(n8223) );
  OR2_X1 U8140 ( .A1(n7697), .A2(n8133), .ZN(n8136) );
  OR2_X1 U8141 ( .A1(n8224), .A2(n8225), .ZN(n8137) );
  AND2_X1 U8142 ( .A1(n8226), .A2(n8227), .ZN(n8225) );
  AND2_X1 U8143 ( .A1(n8228), .A2(n8229), .ZN(n8224) );
  OR2_X1 U8144 ( .A1(n8227), .A2(n8226), .ZN(n8229) );
  XOR2_X1 U8145 ( .A(n8145), .B(n8230), .Z(n8138) );
  XOR2_X1 U8146 ( .A(n8144), .B(n8143), .Z(n8230) );
  OR2_X1 U8147 ( .A1(n8050), .A2(n7730), .ZN(n8143) );
  OR2_X1 U8148 ( .A1(n8231), .A2(n8232), .ZN(n8144) );
  AND2_X1 U8149 ( .A1(n8233), .A2(n8234), .ZN(n8232) );
  AND2_X1 U8150 ( .A1(n8235), .A2(n8236), .ZN(n8231) );
  OR2_X1 U8151 ( .A1(n8233), .A2(n8234), .ZN(n8236) );
  XOR2_X1 U8152 ( .A(n8152), .B(n8237), .Z(n8145) );
  XOR2_X1 U8153 ( .A(n8151), .B(n8150), .Z(n8237) );
  OR2_X1 U8154 ( .A1(n7981), .A2(n7820), .ZN(n8150) );
  OR2_X1 U8155 ( .A1(n8238), .A2(n8239), .ZN(n8151) );
  AND2_X1 U8156 ( .A1(n8240), .A2(n8241), .ZN(n8239) );
  AND2_X1 U8157 ( .A1(n8242), .A2(n8243), .ZN(n8238) );
  OR2_X1 U8158 ( .A1(n8241), .A2(n8240), .ZN(n8243) );
  XOR2_X1 U8159 ( .A(n8159), .B(n8244), .Z(n8152) );
  XOR2_X1 U8160 ( .A(n8158), .B(n8157), .Z(n8244) );
  OR2_X1 U8161 ( .A1(n7912), .A2(n7828), .ZN(n8157) );
  OR2_X1 U8162 ( .A1(n8245), .A2(n8246), .ZN(n8158) );
  AND2_X1 U8163 ( .A1(n8247), .A2(n8248), .ZN(n8246) );
  AND2_X1 U8164 ( .A1(n8249), .A2(n8250), .ZN(n8245) );
  OR2_X1 U8165 ( .A1(n8248), .A2(n8247), .ZN(n8250) );
  XOR2_X1 U8166 ( .A(n8166), .B(n8251), .Z(n8159) );
  XOR2_X1 U8167 ( .A(n8165), .B(n8164), .Z(n8251) );
  OR2_X1 U8168 ( .A1(n7857), .A2(n7887), .ZN(n8164) );
  OR2_X1 U8169 ( .A1(n8252), .A2(n8253), .ZN(n8165) );
  AND2_X1 U8170 ( .A1(n8254), .A2(n8255), .ZN(n8253) );
  AND2_X1 U8171 ( .A1(n8256), .A2(n8257), .ZN(n8252) );
  OR2_X1 U8172 ( .A1(n8255), .A2(n8254), .ZN(n8257) );
  XOR2_X1 U8173 ( .A(n8173), .B(n8258), .Z(n8166) );
  XOR2_X1 U8174 ( .A(n8172), .B(n8171), .Z(n8258) );
  OR2_X1 U8175 ( .A1(n7798), .A2(n7955), .ZN(n8171) );
  OR2_X1 U8176 ( .A1(n8259), .A2(n8260), .ZN(n8172) );
  AND2_X1 U8177 ( .A1(n8261), .A2(n8262), .ZN(n8260) );
  AND2_X1 U8178 ( .A1(n8263), .A2(n8264), .ZN(n8259) );
  OR2_X1 U8179 ( .A1(n8261), .A2(n8262), .ZN(n8263) );
  XOR2_X1 U8180 ( .A(n8206), .B(n8265), .Z(n8173) );
  XOR2_X1 U8181 ( .A(n8205), .B(n8204), .Z(n8265) );
  OR2_X1 U8182 ( .A1(n7759), .A2(n8025), .ZN(n8204) );
  OR2_X1 U8183 ( .A1(n8266), .A2(n8267), .ZN(n8205) );
  AND2_X1 U8184 ( .A1(n8268), .A2(n8269), .ZN(n8267) );
  AND2_X1 U8185 ( .A1(n8270), .A2(n8271), .ZN(n8266) );
  OR2_X1 U8186 ( .A1(n8269), .A2(n8268), .ZN(n8271) );
  XOR2_X1 U8187 ( .A(n8181), .B(n8272), .Z(n8206) );
  XOR2_X1 U8188 ( .A(n8180), .B(n8179), .Z(n8272) );
  OR2_X1 U8189 ( .A1(n7715), .A2(n8107), .ZN(n8179) );
  OR2_X1 U8190 ( .A1(n8273), .A2(n8274), .ZN(n8180) );
  AND2_X1 U8191 ( .A1(n8275), .A2(n8276), .ZN(n8274) );
  AND2_X1 U8192 ( .A1(n8277), .A2(n8278), .ZN(n8273) );
  OR2_X1 U8193 ( .A1(n8276), .A2(n8275), .ZN(n8278) );
  XOR2_X1 U8194 ( .A(n8188), .B(n8279), .Z(n8181) );
  XOR2_X1 U8195 ( .A(n8187), .B(n8186), .Z(n8279) );
  OR2_X1 U8196 ( .A1(n7689), .A2(n8191), .ZN(n8186) );
  OR2_X1 U8197 ( .A1(n8280), .A2(n8281), .ZN(n8187) );
  AND2_X1 U8198 ( .A1(n8282), .A2(n8283), .ZN(n8281) );
  AND2_X1 U8199 ( .A1(n8284), .A2(n8285), .ZN(n8280) );
  OR2_X1 U8200 ( .A1(n8283), .A2(n8282), .ZN(n8285) );
  XOR2_X1 U8201 ( .A(n8196), .B(n8286), .Z(n8188) );
  XOR2_X1 U8202 ( .A(n8195), .B(n8194), .Z(n8286) );
  OR2_X1 U8203 ( .A1(n7659), .A2(n8287), .ZN(n8194) );
  OR2_X1 U8204 ( .A1(n8288), .A2(n8289), .ZN(n8195) );
  AND2_X1 U8205 ( .A1(n8290), .A2(n8291), .ZN(n8289) );
  AND2_X1 U8206 ( .A1(n8292), .A2(n8293), .ZN(n8288) );
  OR2_X1 U8207 ( .A1(n8291), .A2(n8290), .ZN(n8293) );
  XOR2_X1 U8208 ( .A(n8294), .B(n8295), .Z(n8196) );
  XOR2_X1 U8209 ( .A(n8296), .B(n8297), .Z(n8295) );
  OR2_X1 U8210 ( .A1(n7586), .A2(n7587), .ZN(n8208) );
  OR2_X1 U8211 ( .A1(n8298), .A2(n7576), .ZN(n7586) );
  AND2_X1 U8212 ( .A1(n8299), .A2(n8300), .ZN(n7576) );
  AND2_X1 U8213 ( .A1(n7574), .A2(n7572), .ZN(n8298) );
  OR2_X1 U8214 ( .A1(n8301), .A2(n7571), .ZN(n7572) );
  AND2_X1 U8215 ( .A1(n8302), .A2(n8303), .ZN(n7571) );
  AND2_X1 U8216 ( .A1(n7567), .A2(n7570), .ZN(n8301) );
  OR2_X1 U8217 ( .A1(n8303), .A2(n8302), .ZN(n7570) );
  XNOR2_X1 U8218 ( .A(n8304), .B(n8305), .ZN(n8302) );
  OR2_X1 U8219 ( .A1(n8306), .A2(n8307), .ZN(n7567) );
  INV_X1 U8220 ( .A(n7566), .ZN(n8307) );
  OR2_X1 U8221 ( .A1(n8308), .A2(n8309), .ZN(n7566) );
  OR2_X1 U8222 ( .A1(n8310), .A2(n8311), .ZN(n8309) );
  OR2_X1 U8223 ( .A1(n8303), .A2(n8312), .ZN(n8308) );
  AND2_X1 U8224 ( .A1(n8313), .A2(n8314), .ZN(n8312) );
  INV_X1 U8225 ( .A(n8315), .ZN(n8303) );
  OR2_X1 U8226 ( .A1(n8313), .A2(n8314), .ZN(n8315) );
  AND2_X1 U8227 ( .A1(n7565), .A2(n7563), .ZN(n8306) );
  OR2_X1 U8228 ( .A1(n8316), .A2(n8317), .ZN(n7563) );
  AND2_X1 U8229 ( .A1(n7556), .A2(n7559), .ZN(n8317) );
  OR2_X1 U8230 ( .A1(n8318), .A2(n7562), .ZN(n7559) );
  OR2_X1 U8231 ( .A1(n8319), .A2(n7555), .ZN(n7556) );
  AND2_X1 U8232 ( .A1(n8320), .A2(n8321), .ZN(n7555) );
  AND2_X1 U8233 ( .A1(n7551), .A2(n7553), .ZN(n8319) );
  OR2_X1 U8234 ( .A1(n8321), .A2(n8320), .ZN(n7553) );
  XOR2_X1 U8235 ( .A(n8322), .B(n8323), .Z(n8320) );
  OR2_X1 U8236 ( .A1(n8324), .A2(n8325), .ZN(n7551) );
  INV_X1 U8237 ( .A(n7541), .ZN(n8325) );
  OR2_X1 U8238 ( .A1(n8326), .A2(n8327), .ZN(n7541) );
  AND2_X1 U8239 ( .A1(n7538), .A2(n7540), .ZN(n8324) );
  INV_X1 U8240 ( .A(n8328), .ZN(n7540) );
  AND2_X1 U8241 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  OR2_X1 U8242 ( .A1(n8329), .A2(n8321), .ZN(n8327) );
  INV_X1 U8243 ( .A(n8330), .ZN(n8321) );
  OR2_X1 U8244 ( .A1(n8331), .A2(n8332), .ZN(n8330) );
  AND2_X1 U8245 ( .A1(n8331), .A2(n8332), .ZN(n8329) );
  OR2_X1 U8246 ( .A1(n8333), .A2(n8334), .ZN(n8332) );
  AND2_X1 U8247 ( .A1(n8335), .A2(n8336), .ZN(n8334) );
  AND2_X1 U8248 ( .A1(n8337), .A2(n8338), .ZN(n8333) );
  OR2_X1 U8249 ( .A1(n8335), .A2(n8336), .ZN(n8337) );
  XOR2_X1 U8250 ( .A(n8339), .B(n8340), .Z(n8331) );
  XOR2_X1 U8251 ( .A(n8341), .B(n8342), .Z(n8340) );
  OR2_X1 U8252 ( .A1(n8343), .A2(n7537), .ZN(n7538) );
  AND2_X1 U8253 ( .A1(n8344), .A2(n8345), .ZN(n7537) );
  AND2_X1 U8254 ( .A1(n7535), .A2(n7533), .ZN(n8343) );
  OR2_X1 U8255 ( .A1(n8346), .A2(n8347), .ZN(n7533) );
  AND2_X1 U8256 ( .A1(n7529), .A2(n7526), .ZN(n8347) );
  OR2_X1 U8257 ( .A1(n8348), .A2(n7525), .ZN(n7526) );
  AND2_X1 U8258 ( .A1(n8349), .A2(n8350), .ZN(n7525) );
  AND2_X1 U8259 ( .A1(n7523), .A2(n7521), .ZN(n8348) );
  OR2_X1 U8260 ( .A1(n8351), .A2(n7520), .ZN(n7521) );
  AND2_X1 U8261 ( .A1(n8352), .A2(n8353), .ZN(n7520) );
  AND2_X1 U8262 ( .A1(n7516), .A2(n7519), .ZN(n8351) );
  OR2_X1 U8263 ( .A1(n8353), .A2(n8352), .ZN(n7519) );
  XNOR2_X1 U8264 ( .A(n8354), .B(n8355), .ZN(n8352) );
  OR2_X1 U8265 ( .A1(n8356), .A2(n8357), .ZN(n7516) );
  INV_X1 U8266 ( .A(n7514), .ZN(n8357) );
  OR2_X1 U8267 ( .A1(n8358), .A2(n8359), .ZN(n7514) );
  AND2_X1 U8268 ( .A1(n7512), .A2(n7515), .ZN(n8356) );
  INV_X1 U8269 ( .A(n8360), .ZN(n7515) );
  AND2_X1 U8270 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  OR2_X1 U8271 ( .A1(n8361), .A2(n8353), .ZN(n8358) );
  INV_X1 U8272 ( .A(n8362), .ZN(n8353) );
  OR2_X1 U8273 ( .A1(n8363), .A2(n8364), .ZN(n8362) );
  AND2_X1 U8274 ( .A1(n8363), .A2(n8364), .ZN(n8361) );
  OR2_X1 U8275 ( .A1(n8365), .A2(n8366), .ZN(n8364) );
  AND2_X1 U8276 ( .A1(n8367), .A2(n8368), .ZN(n8366) );
  AND2_X1 U8277 ( .A1(n8369), .A2(n8370), .ZN(n8365) );
  OR2_X1 U8278 ( .A1(n8367), .A2(n8368), .ZN(n8370) );
  XOR2_X1 U8279 ( .A(n8371), .B(n8372), .Z(n8363) );
  XOR2_X1 U8280 ( .A(n8373), .B(n8374), .Z(n8372) );
  OR2_X1 U8281 ( .A1(n8375), .A2(n8376), .ZN(n8359) );
  OR2_X1 U8282 ( .A1(n8377), .A2(n7511), .ZN(n7512) );
  AND2_X1 U8283 ( .A1(n8378), .A2(n8379), .ZN(n7511) );
  AND2_X1 U8284 ( .A1(n7509), .A2(n7507), .ZN(n8377) );
  OR2_X1 U8285 ( .A1(n8380), .A2(n7506), .ZN(n7507) );
  AND2_X1 U8286 ( .A1(n8381), .A2(n8382), .ZN(n7506) );
  AND2_X1 U8287 ( .A1(n7504), .A2(n7502), .ZN(n8380) );
  OR2_X1 U8288 ( .A1(n8383), .A2(n8384), .ZN(n7502) );
  INV_X1 U8289 ( .A(n7501), .ZN(n8384) );
  OR2_X1 U8290 ( .A1(n8385), .A2(n8386), .ZN(n7501) );
  OR2_X1 U8291 ( .A1(n8387), .A2(n8388), .ZN(n8386) );
  XNOR2_X1 U8292 ( .A(n8389), .B(n8390), .ZN(n8388) );
  INV_X1 U8293 ( .A(n8391), .ZN(n8387) );
  AND2_X1 U8294 ( .A1(n7500), .A2(n7498), .ZN(n8383) );
  OR2_X1 U8295 ( .A1(n8392), .A2(n8393), .ZN(n7498) );
  INV_X1 U8296 ( .A(n7496), .ZN(n8393) );
  OR2_X1 U8297 ( .A1(n8394), .A2(n8395), .ZN(n7496) );
  OR2_X1 U8298 ( .A1(n8396), .A2(n8397), .ZN(n8395) );
  XNOR2_X1 U8299 ( .A(n8391), .B(n8398), .ZN(n8396) );
  AND2_X1 U8300 ( .A1(n7497), .A2(n7495), .ZN(n8392) );
  OR2_X1 U8301 ( .A1(n8399), .A2(n8400), .ZN(n7495) );
  XNOR2_X1 U8302 ( .A(n8385), .B(n8391), .ZN(n8400) );
  INV_X1 U8303 ( .A(n8401), .ZN(n8399) );
  OR2_X1 U8304 ( .A1(n8394), .A2(n8397), .ZN(n8401) );
  AND2_X1 U8305 ( .A1(n7491), .A2(n8402), .ZN(n7497) );
  AND2_X1 U8306 ( .A1(n7486), .A2(n7490), .ZN(n8402) );
  XOR2_X1 U8307 ( .A(n8397), .B(n8394), .Z(n7490) );
  OR2_X1 U8308 ( .A1(n8403), .A2(n8404), .ZN(n8394) );
  AND2_X1 U8309 ( .A1(n8405), .A2(n8406), .ZN(n8404) );
  AND2_X1 U8310 ( .A1(n8407), .A2(n8408), .ZN(n8403) );
  OR2_X1 U8311 ( .A1(n8405), .A2(n8406), .ZN(n8408) );
  XOR2_X1 U8312 ( .A(n8409), .B(n8410), .Z(n8397) );
  XOR2_X1 U8313 ( .A(n8411), .B(n8412), .Z(n8410) );
  XNOR2_X1 U8314 ( .A(n8407), .B(n8413), .ZN(n7486) );
  XOR2_X1 U8315 ( .A(n8406), .B(n8405), .Z(n8413) );
  OR2_X1 U8316 ( .A1(n7660), .A2(n7344), .ZN(n8405) );
  OR2_X1 U8317 ( .A1(n8414), .A2(n8415), .ZN(n8406) );
  AND2_X1 U8318 ( .A1(n8416), .A2(n8417), .ZN(n8415) );
  AND2_X1 U8319 ( .A1(n8418), .A2(n8419), .ZN(n8414) );
  OR2_X1 U8320 ( .A1(n8417), .A2(n8416), .ZN(n8418) );
  XOR2_X1 U8321 ( .A(n8420), .B(n8421), .Z(n8407) );
  XOR2_X1 U8322 ( .A(n8422), .B(n8423), .Z(n8421) );
  INV_X1 U8323 ( .A(n7485), .ZN(n7491) );
  OR2_X1 U8324 ( .A1(n8424), .A2(n8425), .ZN(n7485) );
  AND2_X1 U8325 ( .A1(n7484), .A2(n7483), .ZN(n8425) );
  AND2_X1 U8326 ( .A1(n7481), .A2(n8426), .ZN(n8424) );
  OR2_X1 U8327 ( .A1(n7484), .A2(n7483), .ZN(n8426) );
  OR2_X1 U8328 ( .A1(n8427), .A2(n8428), .ZN(n7483) );
  AND2_X1 U8329 ( .A1(n7480), .A2(n7479), .ZN(n8428) );
  AND2_X1 U8330 ( .A1(n7477), .A2(n8429), .ZN(n8427) );
  OR2_X1 U8331 ( .A1(n7480), .A2(n7479), .ZN(n8429) );
  OR2_X1 U8332 ( .A1(n8430), .A2(n8431), .ZN(n7479) );
  AND2_X1 U8333 ( .A1(n7476), .A2(n7475), .ZN(n8431) );
  AND2_X1 U8334 ( .A1(n7473), .A2(n8432), .ZN(n8430) );
  OR2_X1 U8335 ( .A1(n7476), .A2(n7475), .ZN(n8432) );
  OR2_X1 U8336 ( .A1(n8433), .A2(n8434), .ZN(n7475) );
  AND2_X1 U8337 ( .A1(n7472), .A2(n7471), .ZN(n8434) );
  AND2_X1 U8338 ( .A1(n7469), .A2(n8435), .ZN(n8433) );
  OR2_X1 U8339 ( .A1(n7472), .A2(n7471), .ZN(n8435) );
  OR2_X1 U8340 ( .A1(n8436), .A2(n8437), .ZN(n7471) );
  AND2_X1 U8341 ( .A1(n7468), .A2(n7467), .ZN(n8437) );
  AND2_X1 U8342 ( .A1(n7465), .A2(n8438), .ZN(n8436) );
  OR2_X1 U8343 ( .A1(n7468), .A2(n7467), .ZN(n8438) );
  OR2_X1 U8344 ( .A1(n8439), .A2(n8440), .ZN(n7467) );
  AND2_X1 U8345 ( .A1(n7464), .A2(n7463), .ZN(n8440) );
  AND2_X1 U8346 ( .A1(n7461), .A2(n8441), .ZN(n8439) );
  OR2_X1 U8347 ( .A1(n7464), .A2(n7463), .ZN(n8441) );
  OR2_X1 U8348 ( .A1(n8442), .A2(n8443), .ZN(n7463) );
  AND2_X1 U8349 ( .A1(n7460), .A2(n7459), .ZN(n8443) );
  AND2_X1 U8350 ( .A1(n7457), .A2(n8444), .ZN(n8442) );
  OR2_X1 U8351 ( .A1(n7460), .A2(n7459), .ZN(n8444) );
  OR2_X1 U8352 ( .A1(n8445), .A2(n8446), .ZN(n7459) );
  AND2_X1 U8353 ( .A1(n7456), .A2(n7455), .ZN(n8446) );
  AND2_X1 U8354 ( .A1(n7453), .A2(n8447), .ZN(n8445) );
  OR2_X1 U8355 ( .A1(n7456), .A2(n7455), .ZN(n8447) );
  OR2_X1 U8356 ( .A1(n8448), .A2(n8449), .ZN(n7455) );
  AND2_X1 U8357 ( .A1(n7445), .A2(n7444), .ZN(n8449) );
  AND2_X1 U8358 ( .A1(n7442), .A2(n8450), .ZN(n8448) );
  OR2_X1 U8359 ( .A1(n7445), .A2(n7444), .ZN(n8450) );
  OR2_X1 U8360 ( .A1(n8451), .A2(n8452), .ZN(n7444) );
  AND2_X1 U8361 ( .A1(n7441), .A2(n7440), .ZN(n8452) );
  AND2_X1 U8362 ( .A1(n7438), .A2(n8453), .ZN(n8451) );
  OR2_X1 U8363 ( .A1(n7441), .A2(n7440), .ZN(n8453) );
  OR2_X1 U8364 ( .A1(n8454), .A2(n8455), .ZN(n7440) );
  AND2_X1 U8365 ( .A1(n7437), .A2(n7436), .ZN(n8455) );
  AND2_X1 U8366 ( .A1(n7434), .A2(n8456), .ZN(n8454) );
  OR2_X1 U8367 ( .A1(n7437), .A2(n7436), .ZN(n8456) );
  OR2_X1 U8368 ( .A1(n8457), .A2(n8458), .ZN(n7436) );
  AND2_X1 U8369 ( .A1(n7433), .A2(n7432), .ZN(n8458) );
  AND2_X1 U8370 ( .A1(n7430), .A2(n8459), .ZN(n8457) );
  OR2_X1 U8371 ( .A1(n7433), .A2(n7432), .ZN(n8459) );
  OR2_X1 U8372 ( .A1(n8460), .A2(n8461), .ZN(n7432) );
  AND2_X1 U8373 ( .A1(n7429), .A2(n7428), .ZN(n8461) );
  AND2_X1 U8374 ( .A1(n7426), .A2(n8462), .ZN(n8460) );
  OR2_X1 U8375 ( .A1(n7429), .A2(n7428), .ZN(n8462) );
  OR2_X1 U8376 ( .A1(n8463), .A2(n8464), .ZN(n7428) );
  AND2_X1 U8377 ( .A1(n7425), .A2(n7424), .ZN(n8464) );
  AND2_X1 U8378 ( .A1(n7422), .A2(n8465), .ZN(n8463) );
  OR2_X1 U8379 ( .A1(n7425), .A2(n7424), .ZN(n8465) );
  OR2_X1 U8380 ( .A1(n8466), .A2(n8467), .ZN(n7424) );
  AND2_X1 U8381 ( .A1(n7421), .A2(n7420), .ZN(n8467) );
  AND2_X1 U8382 ( .A1(n7418), .A2(n8468), .ZN(n8466) );
  OR2_X1 U8383 ( .A1(n7421), .A2(n7420), .ZN(n8468) );
  OR2_X1 U8384 ( .A1(n8469), .A2(n8470), .ZN(n7420) );
  AND2_X1 U8385 ( .A1(n7417), .A2(n7416), .ZN(n8470) );
  AND2_X1 U8386 ( .A1(n7414), .A2(n8471), .ZN(n8469) );
  OR2_X1 U8387 ( .A1(n7417), .A2(n7416), .ZN(n8471) );
  OR2_X1 U8388 ( .A1(n8472), .A2(n8473), .ZN(n7416) );
  AND2_X1 U8389 ( .A1(n7413), .A2(n7412), .ZN(n8473) );
  AND2_X1 U8390 ( .A1(n7410), .A2(n8474), .ZN(n8472) );
  OR2_X1 U8391 ( .A1(n7413), .A2(n7412), .ZN(n8474) );
  OR2_X1 U8392 ( .A1(n8475), .A2(n8476), .ZN(n7412) );
  AND2_X1 U8393 ( .A1(n7409), .A2(n7408), .ZN(n8476) );
  AND2_X1 U8394 ( .A1(n7406), .A2(n8477), .ZN(n8475) );
  OR2_X1 U8395 ( .A1(n7409), .A2(n7408), .ZN(n8477) );
  OR2_X1 U8396 ( .A1(n8478), .A2(n8479), .ZN(n7408) );
  AND2_X1 U8397 ( .A1(n7403), .A2(n7402), .ZN(n8479) );
  AND2_X1 U8398 ( .A1(n7400), .A2(n8480), .ZN(n8478) );
  OR2_X1 U8399 ( .A1(n7403), .A2(n7402), .ZN(n8480) );
  OR2_X1 U8400 ( .A1(n8481), .A2(n8482), .ZN(n7402) );
  AND2_X1 U8401 ( .A1(n7399), .A2(n7398), .ZN(n8482) );
  AND2_X1 U8402 ( .A1(n7396), .A2(n8483), .ZN(n8481) );
  OR2_X1 U8403 ( .A1(n7399), .A2(n7398), .ZN(n8483) );
  OR2_X1 U8404 ( .A1(n8484), .A2(n8485), .ZN(n7398) );
  AND2_X1 U8405 ( .A1(n7395), .A2(n7394), .ZN(n8485) );
  AND2_X1 U8406 ( .A1(n7392), .A2(n8486), .ZN(n8484) );
  OR2_X1 U8407 ( .A1(n7395), .A2(n7394), .ZN(n8486) );
  OR2_X1 U8408 ( .A1(n8487), .A2(n8488), .ZN(n7394) );
  AND2_X1 U8409 ( .A1(n7391), .A2(n7390), .ZN(n8488) );
  AND2_X1 U8410 ( .A1(n7388), .A2(n8489), .ZN(n8487) );
  OR2_X1 U8411 ( .A1(n7391), .A2(n7390), .ZN(n8489) );
  OR2_X1 U8412 ( .A1(n8490), .A2(n8491), .ZN(n7390) );
  AND2_X1 U8413 ( .A1(n7387), .A2(n7386), .ZN(n8491) );
  AND2_X1 U8414 ( .A1(n7384), .A2(n8492), .ZN(n8490) );
  OR2_X1 U8415 ( .A1(n7387), .A2(n7386), .ZN(n8492) );
  OR2_X1 U8416 ( .A1(n8493), .A2(n8494), .ZN(n7386) );
  AND2_X1 U8417 ( .A1(n7383), .A2(n7382), .ZN(n8494) );
  AND2_X1 U8418 ( .A1(n7380), .A2(n8495), .ZN(n8493) );
  OR2_X1 U8419 ( .A1(n7383), .A2(n7382), .ZN(n8495) );
  OR2_X1 U8420 ( .A1(n8496), .A2(n8497), .ZN(n7382) );
  AND2_X1 U8421 ( .A1(n7379), .A2(n7378), .ZN(n8497) );
  AND2_X1 U8422 ( .A1(n7376), .A2(n8498), .ZN(n8496) );
  OR2_X1 U8423 ( .A1(n7379), .A2(n7378), .ZN(n8498) );
  OR2_X1 U8424 ( .A1(n8499), .A2(n8500), .ZN(n7378) );
  AND2_X1 U8425 ( .A1(n7375), .A2(n7374), .ZN(n8500) );
  AND2_X1 U8426 ( .A1(n7372), .A2(n8501), .ZN(n8499) );
  OR2_X1 U8427 ( .A1(n7375), .A2(n7374), .ZN(n8501) );
  OR2_X1 U8428 ( .A1(n8502), .A2(n8503), .ZN(n7374) );
  AND2_X1 U8429 ( .A1(n7371), .A2(n7370), .ZN(n8503) );
  AND2_X1 U8430 ( .A1(n7368), .A2(n8504), .ZN(n8502) );
  OR2_X1 U8431 ( .A1(n7371), .A2(n7370), .ZN(n8504) );
  OR2_X1 U8432 ( .A1(n8505), .A2(n8506), .ZN(n7370) );
  AND2_X1 U8433 ( .A1(n7367), .A2(n7366), .ZN(n8506) );
  AND2_X1 U8434 ( .A1(n7364), .A2(n8507), .ZN(n8505) );
  OR2_X1 U8435 ( .A1(n7367), .A2(n7366), .ZN(n8507) );
  OR2_X1 U8436 ( .A1(n8508), .A2(n8509), .ZN(n7366) );
  AND2_X1 U8437 ( .A1(n7356), .A2(n7355), .ZN(n8509) );
  AND2_X1 U8438 ( .A1(n7354), .A2(n8510), .ZN(n8508) );
  OR2_X1 U8439 ( .A1(n7356), .A2(n7355), .ZN(n8510) );
  OR2_X1 U8440 ( .A1(n8511), .A2(n8512), .ZN(n7355) );
  AND2_X1 U8441 ( .A1(n7350), .A2(n7351), .ZN(n8512) );
  AND2_X1 U8442 ( .A1(n8513), .A2(n8514), .ZN(n8511) );
  OR2_X1 U8443 ( .A1(n7350), .A2(n7351), .ZN(n8514) );
  OR2_X1 U8444 ( .A1(n8515), .A2(n7348), .ZN(n7351) );
  INV_X1 U8445 ( .A(n7352), .ZN(n8513) );
  OR2_X1 U8446 ( .A1(n8516), .A2(n8517), .ZN(n7352) );
  AND2_X1 U8447 ( .A1(b_30_), .A2(n8518), .ZN(n8517) );
  OR2_X1 U8448 ( .A1(n8519), .A2(n7343), .ZN(n8518) );
  AND2_X1 U8449 ( .A1(a_30_), .A2(n8520), .ZN(n8519) );
  AND2_X1 U8450 ( .A1(b_29_), .A2(n8521), .ZN(n8516) );
  OR2_X1 U8451 ( .A1(n8522), .A2(n7347), .ZN(n8521) );
  AND2_X1 U8452 ( .A1(a_31_), .A2(n7344), .ZN(n8522) );
  OR2_X1 U8453 ( .A1(n8523), .A2(n7348), .ZN(n7356) );
  XOR2_X1 U8454 ( .A(n8524), .B(n8525), .Z(n7354) );
  XNOR2_X1 U8455 ( .A(n8526), .B(n8527), .ZN(n8524) );
  OR2_X1 U8456 ( .A1(n8528), .A2(n7348), .ZN(n7367) );
  XOR2_X1 U8457 ( .A(n8529), .B(n8530), .Z(n7364) );
  XOR2_X1 U8458 ( .A(n8531), .B(n8532), .Z(n8530) );
  OR2_X1 U8459 ( .A1(n8533), .A2(n7348), .ZN(n7371) );
  XOR2_X1 U8460 ( .A(n8534), .B(n8535), .Z(n7368) );
  XOR2_X1 U8461 ( .A(n8536), .B(n8537), .Z(n8535) );
  OR2_X1 U8462 ( .A1(n8538), .A2(n7348), .ZN(n7375) );
  XOR2_X1 U8463 ( .A(n8539), .B(n8540), .Z(n7372) );
  XOR2_X1 U8464 ( .A(n8541), .B(n8542), .Z(n8540) );
  OR2_X1 U8465 ( .A1(n8543), .A2(n7348), .ZN(n7379) );
  XOR2_X1 U8466 ( .A(n8544), .B(n8545), .Z(n7376) );
  XOR2_X1 U8467 ( .A(n8546), .B(n8547), .Z(n8545) );
  OR2_X1 U8468 ( .A1(n8548), .A2(n7348), .ZN(n7383) );
  XOR2_X1 U8469 ( .A(n8549), .B(n8550), .Z(n7380) );
  XOR2_X1 U8470 ( .A(n8551), .B(n8552), .Z(n8550) );
  OR2_X1 U8471 ( .A1(n8553), .A2(n7348), .ZN(n7387) );
  XOR2_X1 U8472 ( .A(n8554), .B(n8555), .Z(n7384) );
  XOR2_X1 U8473 ( .A(n8556), .B(n8557), .Z(n8555) );
  OR2_X1 U8474 ( .A1(n8558), .A2(n7348), .ZN(n7391) );
  XOR2_X1 U8475 ( .A(n8559), .B(n8560), .Z(n7388) );
  XOR2_X1 U8476 ( .A(n8561), .B(n8562), .Z(n8560) );
  OR2_X1 U8477 ( .A1(n8563), .A2(n7348), .ZN(n7395) );
  XOR2_X1 U8478 ( .A(n8564), .B(n8565), .Z(n7392) );
  XOR2_X1 U8479 ( .A(n8566), .B(n8567), .Z(n8565) );
  OR2_X1 U8480 ( .A1(n8568), .A2(n7348), .ZN(n7399) );
  XOR2_X1 U8481 ( .A(n8569), .B(n8570), .Z(n7396) );
  XOR2_X1 U8482 ( .A(n8571), .B(n8572), .Z(n8570) );
  OR2_X1 U8483 ( .A1(n8573), .A2(n7348), .ZN(n7403) );
  XOR2_X1 U8484 ( .A(n8574), .B(n8575), .Z(n7400) );
  XOR2_X1 U8485 ( .A(n8576), .B(n8577), .Z(n8575) );
  OR2_X1 U8486 ( .A1(n8578), .A2(n7348), .ZN(n7409) );
  XOR2_X1 U8487 ( .A(n8579), .B(n8580), .Z(n7406) );
  XOR2_X1 U8488 ( .A(n8581), .B(n8582), .Z(n8580) );
  OR2_X1 U8489 ( .A1(n8583), .A2(n7348), .ZN(n7413) );
  XOR2_X1 U8490 ( .A(n8584), .B(n8585), .Z(n7410) );
  XOR2_X1 U8491 ( .A(n8586), .B(n8587), .Z(n8585) );
  OR2_X1 U8492 ( .A1(n8588), .A2(n7348), .ZN(n7417) );
  XOR2_X1 U8493 ( .A(n8589), .B(n8590), .Z(n7414) );
  XOR2_X1 U8494 ( .A(n8591), .B(n8592), .Z(n8590) );
  OR2_X1 U8495 ( .A1(n8593), .A2(n7348), .ZN(n7421) );
  XOR2_X1 U8496 ( .A(n8594), .B(n8595), .Z(n7418) );
  XOR2_X1 U8497 ( .A(n8596), .B(n8597), .Z(n8595) );
  OR2_X1 U8498 ( .A1(n8598), .A2(n7348), .ZN(n7425) );
  XOR2_X1 U8499 ( .A(n8599), .B(n8600), .Z(n7422) );
  XOR2_X1 U8500 ( .A(n8601), .B(n8602), .Z(n8600) );
  OR2_X1 U8501 ( .A1(n8603), .A2(n7348), .ZN(n7429) );
  XOR2_X1 U8502 ( .A(n8604), .B(n8605), .Z(n7426) );
  XOR2_X1 U8503 ( .A(n8606), .B(n8607), .Z(n8605) );
  OR2_X1 U8504 ( .A1(n8608), .A2(n7348), .ZN(n7433) );
  XOR2_X1 U8505 ( .A(n8609), .B(n8610), .Z(n7430) );
  XOR2_X1 U8506 ( .A(n8611), .B(n8612), .Z(n8610) );
  OR2_X1 U8507 ( .A1(n8287), .A2(n7348), .ZN(n7437) );
  XOR2_X1 U8508 ( .A(n8613), .B(n8614), .Z(n7434) );
  XOR2_X1 U8509 ( .A(n8615), .B(n8616), .Z(n8614) );
  OR2_X1 U8510 ( .A1(n8191), .A2(n7348), .ZN(n7441) );
  XOR2_X1 U8511 ( .A(n8617), .B(n8618), .Z(n7438) );
  XOR2_X1 U8512 ( .A(n8619), .B(n8620), .Z(n8618) );
  OR2_X1 U8513 ( .A1(n8107), .A2(n7348), .ZN(n7445) );
  XOR2_X1 U8514 ( .A(n8621), .B(n8622), .Z(n7442) );
  XOR2_X1 U8515 ( .A(n8623), .B(n8624), .Z(n8622) );
  OR2_X1 U8516 ( .A1(n8025), .A2(n7348), .ZN(n7456) );
  XOR2_X1 U8517 ( .A(n8625), .B(n8626), .Z(n7453) );
  XOR2_X1 U8518 ( .A(n8627), .B(n8628), .Z(n8626) );
  OR2_X1 U8519 ( .A1(n7955), .A2(n7348), .ZN(n7460) );
  XOR2_X1 U8520 ( .A(n8629), .B(n8630), .Z(n7457) );
  XOR2_X1 U8521 ( .A(n8631), .B(n8632), .Z(n8630) );
  OR2_X1 U8522 ( .A1(n7887), .A2(n7348), .ZN(n7464) );
  XOR2_X1 U8523 ( .A(n8633), .B(n8634), .Z(n7461) );
  XOR2_X1 U8524 ( .A(n8635), .B(n8636), .Z(n8634) );
  OR2_X1 U8525 ( .A1(n7828), .A2(n7348), .ZN(n7468) );
  XOR2_X1 U8526 ( .A(n8637), .B(n8638), .Z(n7465) );
  XOR2_X1 U8527 ( .A(n8639), .B(n8640), .Z(n8638) );
  OR2_X1 U8528 ( .A1(n7820), .A2(n7348), .ZN(n7472) );
  XOR2_X1 U8529 ( .A(n8641), .B(n8642), .Z(n7469) );
  XOR2_X1 U8530 ( .A(n8643), .B(n8644), .Z(n8642) );
  OR2_X1 U8531 ( .A1(n7730), .A2(n7348), .ZN(n7476) );
  XOR2_X1 U8532 ( .A(n8645), .B(n8646), .Z(n7473) );
  XOR2_X1 U8533 ( .A(n8647), .B(n8648), .Z(n8646) );
  OR2_X1 U8534 ( .A1(n7697), .A2(n7348), .ZN(n7480) );
  XOR2_X1 U8535 ( .A(n8649), .B(n8650), .Z(n7477) );
  XOR2_X1 U8536 ( .A(n8651), .B(n8652), .Z(n8650) );
  OR2_X1 U8537 ( .A1(n7660), .A2(n7348), .ZN(n7484) );
  XOR2_X1 U8538 ( .A(n8416), .B(n8653), .Z(n7481) );
  XOR2_X1 U8539 ( .A(n8419), .B(n8417), .Z(n8653) );
  OR2_X1 U8540 ( .A1(n7697), .A2(n7344), .ZN(n8417) );
  OR2_X1 U8541 ( .A1(n8654), .A2(n8655), .ZN(n8419) );
  AND2_X1 U8542 ( .A1(n8649), .A2(n8652), .ZN(n8655) );
  AND2_X1 U8543 ( .A1(n8656), .A2(n8651), .ZN(n8654) );
  OR2_X1 U8544 ( .A1(n8657), .A2(n8658), .ZN(n8651) );
  AND2_X1 U8545 ( .A1(n8645), .A2(n8648), .ZN(n8658) );
  AND2_X1 U8546 ( .A1(n8659), .A2(n8647), .ZN(n8657) );
  OR2_X1 U8547 ( .A1(n8660), .A2(n8661), .ZN(n8647) );
  AND2_X1 U8548 ( .A1(n8641), .A2(n8644), .ZN(n8661) );
  AND2_X1 U8549 ( .A1(n8662), .A2(n8643), .ZN(n8660) );
  OR2_X1 U8550 ( .A1(n8663), .A2(n8664), .ZN(n8643) );
  AND2_X1 U8551 ( .A1(n8637), .A2(n8640), .ZN(n8664) );
  AND2_X1 U8552 ( .A1(n8665), .A2(n8639), .ZN(n8663) );
  OR2_X1 U8553 ( .A1(n8666), .A2(n8667), .ZN(n8639) );
  AND2_X1 U8554 ( .A1(n8633), .A2(n8636), .ZN(n8667) );
  AND2_X1 U8555 ( .A1(n8668), .A2(n8635), .ZN(n8666) );
  OR2_X1 U8556 ( .A1(n8669), .A2(n8670), .ZN(n8635) );
  AND2_X1 U8557 ( .A1(n8629), .A2(n8632), .ZN(n8670) );
  AND2_X1 U8558 ( .A1(n8671), .A2(n8631), .ZN(n8669) );
  OR2_X1 U8559 ( .A1(n8672), .A2(n8673), .ZN(n8631) );
  AND2_X1 U8560 ( .A1(n8625), .A2(n8628), .ZN(n8673) );
  AND2_X1 U8561 ( .A1(n8674), .A2(n8627), .ZN(n8672) );
  OR2_X1 U8562 ( .A1(n8675), .A2(n8676), .ZN(n8627) );
  AND2_X1 U8563 ( .A1(n8621), .A2(n8624), .ZN(n8676) );
  AND2_X1 U8564 ( .A1(n8677), .A2(n8623), .ZN(n8675) );
  OR2_X1 U8565 ( .A1(n8678), .A2(n8679), .ZN(n8623) );
  AND2_X1 U8566 ( .A1(n8617), .A2(n8620), .ZN(n8679) );
  AND2_X1 U8567 ( .A1(n8680), .A2(n8619), .ZN(n8678) );
  OR2_X1 U8568 ( .A1(n8681), .A2(n8682), .ZN(n8619) );
  AND2_X1 U8569 ( .A1(n8613), .A2(n8616), .ZN(n8682) );
  AND2_X1 U8570 ( .A1(n8683), .A2(n8615), .ZN(n8681) );
  OR2_X1 U8571 ( .A1(n8684), .A2(n8685), .ZN(n8615) );
  AND2_X1 U8572 ( .A1(n8609), .A2(n8612), .ZN(n8685) );
  AND2_X1 U8573 ( .A1(n8686), .A2(n8611), .ZN(n8684) );
  OR2_X1 U8574 ( .A1(n8687), .A2(n8688), .ZN(n8611) );
  AND2_X1 U8575 ( .A1(n8604), .A2(n8607), .ZN(n8688) );
  AND2_X1 U8576 ( .A1(n8689), .A2(n8606), .ZN(n8687) );
  OR2_X1 U8577 ( .A1(n8690), .A2(n8691), .ZN(n8606) );
  AND2_X1 U8578 ( .A1(n8599), .A2(n8602), .ZN(n8691) );
  AND2_X1 U8579 ( .A1(n8692), .A2(n8601), .ZN(n8690) );
  OR2_X1 U8580 ( .A1(n8693), .A2(n8694), .ZN(n8601) );
  AND2_X1 U8581 ( .A1(n8594), .A2(n8597), .ZN(n8694) );
  AND2_X1 U8582 ( .A1(n8695), .A2(n8596), .ZN(n8693) );
  OR2_X1 U8583 ( .A1(n8696), .A2(n8697), .ZN(n8596) );
  AND2_X1 U8584 ( .A1(n8589), .A2(n8592), .ZN(n8697) );
  AND2_X1 U8585 ( .A1(n8698), .A2(n8591), .ZN(n8696) );
  OR2_X1 U8586 ( .A1(n8699), .A2(n8700), .ZN(n8591) );
  AND2_X1 U8587 ( .A1(n8584), .A2(n8587), .ZN(n8700) );
  AND2_X1 U8588 ( .A1(n8701), .A2(n8586), .ZN(n8699) );
  OR2_X1 U8589 ( .A1(n8702), .A2(n8703), .ZN(n8586) );
  AND2_X1 U8590 ( .A1(n8579), .A2(n8582), .ZN(n8703) );
  AND2_X1 U8591 ( .A1(n8704), .A2(n8581), .ZN(n8702) );
  OR2_X1 U8592 ( .A1(n8705), .A2(n8706), .ZN(n8581) );
  AND2_X1 U8593 ( .A1(n8574), .A2(n8577), .ZN(n8706) );
  AND2_X1 U8594 ( .A1(n8707), .A2(n8576), .ZN(n8705) );
  OR2_X1 U8595 ( .A1(n8708), .A2(n8709), .ZN(n8576) );
  AND2_X1 U8596 ( .A1(n8569), .A2(n8572), .ZN(n8709) );
  AND2_X1 U8597 ( .A1(n8710), .A2(n8571), .ZN(n8708) );
  OR2_X1 U8598 ( .A1(n8711), .A2(n8712), .ZN(n8571) );
  AND2_X1 U8599 ( .A1(n8564), .A2(n8567), .ZN(n8712) );
  AND2_X1 U8600 ( .A1(n8713), .A2(n8566), .ZN(n8711) );
  OR2_X1 U8601 ( .A1(n8714), .A2(n8715), .ZN(n8566) );
  AND2_X1 U8602 ( .A1(n8559), .A2(n8562), .ZN(n8715) );
  AND2_X1 U8603 ( .A1(n8716), .A2(n8561), .ZN(n8714) );
  OR2_X1 U8604 ( .A1(n8717), .A2(n8718), .ZN(n8561) );
  AND2_X1 U8605 ( .A1(n8554), .A2(n8557), .ZN(n8718) );
  AND2_X1 U8606 ( .A1(n8719), .A2(n8556), .ZN(n8717) );
  OR2_X1 U8607 ( .A1(n8720), .A2(n8721), .ZN(n8556) );
  AND2_X1 U8608 ( .A1(n8549), .A2(n8552), .ZN(n8721) );
  AND2_X1 U8609 ( .A1(n8722), .A2(n8551), .ZN(n8720) );
  OR2_X1 U8610 ( .A1(n8723), .A2(n8724), .ZN(n8551) );
  AND2_X1 U8611 ( .A1(n8544), .A2(n8547), .ZN(n8724) );
  AND2_X1 U8612 ( .A1(n8725), .A2(n8546), .ZN(n8723) );
  OR2_X1 U8613 ( .A1(n8726), .A2(n8727), .ZN(n8546) );
  AND2_X1 U8614 ( .A1(n8539), .A2(n8542), .ZN(n8727) );
  AND2_X1 U8615 ( .A1(n8728), .A2(n8541), .ZN(n8726) );
  OR2_X1 U8616 ( .A1(n8729), .A2(n8730), .ZN(n8541) );
  AND2_X1 U8617 ( .A1(n8534), .A2(n8537), .ZN(n8730) );
  AND2_X1 U8618 ( .A1(n8731), .A2(n8536), .ZN(n8729) );
  OR2_X1 U8619 ( .A1(n8732), .A2(n8733), .ZN(n8536) );
  AND2_X1 U8620 ( .A1(n8529), .A2(n8532), .ZN(n8733) );
  AND2_X1 U8621 ( .A1(n8734), .A2(n8531), .ZN(n8732) );
  OR2_X1 U8622 ( .A1(n8735), .A2(n8736), .ZN(n8531) );
  AND2_X1 U8623 ( .A1(n8525), .A2(n8526), .ZN(n8736) );
  AND2_X1 U8624 ( .A1(n8737), .A2(n8738), .ZN(n8735) );
  OR2_X1 U8625 ( .A1(n8526), .A2(n8525), .ZN(n8738) );
  OR2_X1 U8626 ( .A1(n8515), .A2(n7344), .ZN(n8525) );
  OR2_X1 U8627 ( .A1(n7344), .A2(n8739), .ZN(n8526) );
  INV_X1 U8628 ( .A(n8527), .ZN(n8737) );
  OR2_X1 U8629 ( .A1(n8740), .A2(n8741), .ZN(n8527) );
  AND2_X1 U8630 ( .A1(b_29_), .A2(n8742), .ZN(n8741) );
  OR2_X1 U8631 ( .A1(n8743), .A2(n7343), .ZN(n8742) );
  AND2_X1 U8632 ( .A1(a_30_), .A2(n8744), .ZN(n8743) );
  AND2_X1 U8633 ( .A1(b_28_), .A2(n8745), .ZN(n8740) );
  OR2_X1 U8634 ( .A1(n8746), .A2(n7347), .ZN(n8745) );
  AND2_X1 U8635 ( .A1(a_31_), .A2(n8520), .ZN(n8746) );
  OR2_X1 U8636 ( .A1(n8532), .A2(n8529), .ZN(n8734) );
  XNOR2_X1 U8637 ( .A(n8747), .B(n8748), .ZN(n8529) );
  XNOR2_X1 U8638 ( .A(n8749), .B(n8750), .ZN(n8748) );
  OR2_X1 U8639 ( .A1(n8523), .A2(n7344), .ZN(n8532) );
  OR2_X1 U8640 ( .A1(n8537), .A2(n8534), .ZN(n8731) );
  XOR2_X1 U8641 ( .A(n8751), .B(n8752), .Z(n8534) );
  XOR2_X1 U8642 ( .A(n8753), .B(n8754), .Z(n8752) );
  OR2_X1 U8643 ( .A1(n8528), .A2(n7344), .ZN(n8537) );
  OR2_X1 U8644 ( .A1(n8542), .A2(n8539), .ZN(n8728) );
  XOR2_X1 U8645 ( .A(n8755), .B(n8756), .Z(n8539) );
  XOR2_X1 U8646 ( .A(n8757), .B(n8758), .Z(n8756) );
  OR2_X1 U8647 ( .A1(n8533), .A2(n7344), .ZN(n8542) );
  OR2_X1 U8648 ( .A1(n8547), .A2(n8544), .ZN(n8725) );
  XOR2_X1 U8649 ( .A(n8759), .B(n8760), .Z(n8544) );
  XOR2_X1 U8650 ( .A(n8761), .B(n8762), .Z(n8760) );
  OR2_X1 U8651 ( .A1(n8538), .A2(n7344), .ZN(n8547) );
  OR2_X1 U8652 ( .A1(n8552), .A2(n8549), .ZN(n8722) );
  XOR2_X1 U8653 ( .A(n8763), .B(n8764), .Z(n8549) );
  XOR2_X1 U8654 ( .A(n8765), .B(n8766), .Z(n8764) );
  OR2_X1 U8655 ( .A1(n8543), .A2(n7344), .ZN(n8552) );
  OR2_X1 U8656 ( .A1(n8557), .A2(n8554), .ZN(n8719) );
  XOR2_X1 U8657 ( .A(n8767), .B(n8768), .Z(n8554) );
  XOR2_X1 U8658 ( .A(n8769), .B(n8770), .Z(n8768) );
  OR2_X1 U8659 ( .A1(n8548), .A2(n7344), .ZN(n8557) );
  OR2_X1 U8660 ( .A1(n8562), .A2(n8559), .ZN(n8716) );
  XOR2_X1 U8661 ( .A(n8771), .B(n8772), .Z(n8559) );
  XOR2_X1 U8662 ( .A(n8773), .B(n8774), .Z(n8772) );
  OR2_X1 U8663 ( .A1(n8553), .A2(n7344), .ZN(n8562) );
  OR2_X1 U8664 ( .A1(n8567), .A2(n8564), .ZN(n8713) );
  XOR2_X1 U8665 ( .A(n8775), .B(n8776), .Z(n8564) );
  XOR2_X1 U8666 ( .A(n8777), .B(n8778), .Z(n8776) );
  OR2_X1 U8667 ( .A1(n8558), .A2(n7344), .ZN(n8567) );
  OR2_X1 U8668 ( .A1(n8572), .A2(n8569), .ZN(n8710) );
  XOR2_X1 U8669 ( .A(n8779), .B(n8780), .Z(n8569) );
  XOR2_X1 U8670 ( .A(n8781), .B(n8782), .Z(n8780) );
  OR2_X1 U8671 ( .A1(n8563), .A2(n7344), .ZN(n8572) );
  OR2_X1 U8672 ( .A1(n8577), .A2(n8574), .ZN(n8707) );
  XOR2_X1 U8673 ( .A(n8783), .B(n8784), .Z(n8574) );
  XOR2_X1 U8674 ( .A(n8785), .B(n8786), .Z(n8784) );
  OR2_X1 U8675 ( .A1(n8568), .A2(n7344), .ZN(n8577) );
  OR2_X1 U8676 ( .A1(n8582), .A2(n8579), .ZN(n8704) );
  XOR2_X1 U8677 ( .A(n8787), .B(n8788), .Z(n8579) );
  XOR2_X1 U8678 ( .A(n8789), .B(n8790), .Z(n8788) );
  OR2_X1 U8679 ( .A1(n8573), .A2(n7344), .ZN(n8582) );
  OR2_X1 U8680 ( .A1(n8587), .A2(n8584), .ZN(n8701) );
  XOR2_X1 U8681 ( .A(n8791), .B(n8792), .Z(n8584) );
  XOR2_X1 U8682 ( .A(n8793), .B(n8794), .Z(n8792) );
  OR2_X1 U8683 ( .A1(n8578), .A2(n7344), .ZN(n8587) );
  OR2_X1 U8684 ( .A1(n8592), .A2(n8589), .ZN(n8698) );
  XOR2_X1 U8685 ( .A(n8795), .B(n8796), .Z(n8589) );
  XOR2_X1 U8686 ( .A(n8797), .B(n8798), .Z(n8796) );
  OR2_X1 U8687 ( .A1(n8583), .A2(n7344), .ZN(n8592) );
  OR2_X1 U8688 ( .A1(n8597), .A2(n8594), .ZN(n8695) );
  XOR2_X1 U8689 ( .A(n8799), .B(n8800), .Z(n8594) );
  XOR2_X1 U8690 ( .A(n8801), .B(n8802), .Z(n8800) );
  OR2_X1 U8691 ( .A1(n8588), .A2(n7344), .ZN(n8597) );
  OR2_X1 U8692 ( .A1(n8602), .A2(n8599), .ZN(n8692) );
  XOR2_X1 U8693 ( .A(n8803), .B(n8804), .Z(n8599) );
  XOR2_X1 U8694 ( .A(n8805), .B(n8806), .Z(n8804) );
  OR2_X1 U8695 ( .A1(n8593), .A2(n7344), .ZN(n8602) );
  OR2_X1 U8696 ( .A1(n8607), .A2(n8604), .ZN(n8689) );
  XOR2_X1 U8697 ( .A(n8807), .B(n8808), .Z(n8604) );
  XOR2_X1 U8698 ( .A(n8809), .B(n8810), .Z(n8808) );
  OR2_X1 U8699 ( .A1(n8598), .A2(n7344), .ZN(n8607) );
  OR2_X1 U8700 ( .A1(n8612), .A2(n8609), .ZN(n8686) );
  XOR2_X1 U8701 ( .A(n8811), .B(n8812), .Z(n8609) );
  XOR2_X1 U8702 ( .A(n8813), .B(n8814), .Z(n8812) );
  OR2_X1 U8703 ( .A1(n8603), .A2(n7344), .ZN(n8612) );
  OR2_X1 U8704 ( .A1(n8616), .A2(n8613), .ZN(n8683) );
  XOR2_X1 U8705 ( .A(n8815), .B(n8816), .Z(n8613) );
  XOR2_X1 U8706 ( .A(n8817), .B(n8818), .Z(n8816) );
  OR2_X1 U8707 ( .A1(n8608), .A2(n7344), .ZN(n8616) );
  OR2_X1 U8708 ( .A1(n8620), .A2(n8617), .ZN(n8680) );
  XOR2_X1 U8709 ( .A(n8819), .B(n8820), .Z(n8617) );
  XOR2_X1 U8710 ( .A(n8821), .B(n8822), .Z(n8820) );
  OR2_X1 U8711 ( .A1(n8287), .A2(n7344), .ZN(n8620) );
  OR2_X1 U8712 ( .A1(n8624), .A2(n8621), .ZN(n8677) );
  XOR2_X1 U8713 ( .A(n8823), .B(n8824), .Z(n8621) );
  XOR2_X1 U8714 ( .A(n8825), .B(n8826), .Z(n8824) );
  OR2_X1 U8715 ( .A1(n8191), .A2(n7344), .ZN(n8624) );
  OR2_X1 U8716 ( .A1(n8628), .A2(n8625), .ZN(n8674) );
  XOR2_X1 U8717 ( .A(n8827), .B(n8828), .Z(n8625) );
  XOR2_X1 U8718 ( .A(n8829), .B(n8830), .Z(n8828) );
  OR2_X1 U8719 ( .A1(n8107), .A2(n7344), .ZN(n8628) );
  OR2_X1 U8720 ( .A1(n8632), .A2(n8629), .ZN(n8671) );
  XOR2_X1 U8721 ( .A(n8831), .B(n8832), .Z(n8629) );
  XOR2_X1 U8722 ( .A(n8833), .B(n8834), .Z(n8832) );
  OR2_X1 U8723 ( .A1(n8025), .A2(n7344), .ZN(n8632) );
  OR2_X1 U8724 ( .A1(n8636), .A2(n8633), .ZN(n8668) );
  XOR2_X1 U8725 ( .A(n8835), .B(n8836), .Z(n8633) );
  XOR2_X1 U8726 ( .A(n8837), .B(n8838), .Z(n8836) );
  OR2_X1 U8727 ( .A1(n7955), .A2(n7344), .ZN(n8636) );
  OR2_X1 U8728 ( .A1(n8640), .A2(n8637), .ZN(n8665) );
  XOR2_X1 U8729 ( .A(n8839), .B(n8840), .Z(n8637) );
  XOR2_X1 U8730 ( .A(n8841), .B(n8842), .Z(n8840) );
  OR2_X1 U8731 ( .A1(n7887), .A2(n7344), .ZN(n8640) );
  OR2_X1 U8732 ( .A1(n8644), .A2(n8641), .ZN(n8662) );
  XOR2_X1 U8733 ( .A(n8843), .B(n8844), .Z(n8641) );
  XOR2_X1 U8734 ( .A(n8845), .B(n8846), .Z(n8844) );
  OR2_X1 U8735 ( .A1(n7828), .A2(n7344), .ZN(n8644) );
  OR2_X1 U8736 ( .A1(n8648), .A2(n8645), .ZN(n8659) );
  XOR2_X1 U8737 ( .A(n8847), .B(n8848), .Z(n8645) );
  XOR2_X1 U8738 ( .A(n8849), .B(n8850), .Z(n8848) );
  OR2_X1 U8739 ( .A1(n7820), .A2(n7344), .ZN(n8648) );
  OR2_X1 U8740 ( .A1(n8652), .A2(n8649), .ZN(n8656) );
  XOR2_X1 U8741 ( .A(n8851), .B(n8852), .Z(n8649) );
  XOR2_X1 U8742 ( .A(n8853), .B(n8854), .Z(n8852) );
  OR2_X1 U8743 ( .A1(n7730), .A2(n7344), .ZN(n8652) );
  XNOR2_X1 U8744 ( .A(n8855), .B(n8856), .ZN(n8416) );
  XNOR2_X1 U8745 ( .A(n8857), .B(n8858), .ZN(n8855) );
  OR2_X1 U8746 ( .A1(n8859), .A2(n8860), .ZN(n7500) );
  XNOR2_X1 U8747 ( .A(n8861), .B(n8389), .ZN(n8860) );
  AND2_X1 U8748 ( .A1(n8398), .A2(n8391), .ZN(n8859) );
  XNOR2_X1 U8749 ( .A(n8862), .B(n8863), .ZN(n8391) );
  XOR2_X1 U8750 ( .A(n8864), .B(n8865), .Z(n8863) );
  INV_X1 U8751 ( .A(n8385), .ZN(n8398) );
  OR2_X1 U8752 ( .A1(n8866), .A2(n8867), .ZN(n8385) );
  AND2_X1 U8753 ( .A1(n8412), .A2(n8411), .ZN(n8867) );
  AND2_X1 U8754 ( .A1(n8409), .A2(n8868), .ZN(n8866) );
  OR2_X1 U8755 ( .A1(n8411), .A2(n8412), .ZN(n8868) );
  OR2_X1 U8756 ( .A1(n7660), .A2(n8520), .ZN(n8412) );
  OR2_X1 U8757 ( .A1(n8869), .A2(n8870), .ZN(n8411) );
  AND2_X1 U8758 ( .A1(n8423), .A2(n8422), .ZN(n8870) );
  AND2_X1 U8759 ( .A1(n8420), .A2(n8871), .ZN(n8869) );
  OR2_X1 U8760 ( .A1(n8422), .A2(n8423), .ZN(n8871) );
  OR2_X1 U8761 ( .A1(n7697), .A2(n8520), .ZN(n8423) );
  OR2_X1 U8762 ( .A1(n8872), .A2(n8873), .ZN(n8422) );
  AND2_X1 U8763 ( .A1(n8858), .A2(n8857), .ZN(n8873) );
  AND2_X1 U8764 ( .A1(n8856), .A2(n8874), .ZN(n8872) );
  OR2_X1 U8765 ( .A1(n8857), .A2(n8858), .ZN(n8874) );
  OR2_X1 U8766 ( .A1(n8875), .A2(n8876), .ZN(n8858) );
  AND2_X1 U8767 ( .A1(n8854), .A2(n8853), .ZN(n8876) );
  AND2_X1 U8768 ( .A1(n8851), .A2(n8877), .ZN(n8875) );
  OR2_X1 U8769 ( .A1(n8853), .A2(n8854), .ZN(n8877) );
  OR2_X1 U8770 ( .A1(n7820), .A2(n8520), .ZN(n8854) );
  OR2_X1 U8771 ( .A1(n8878), .A2(n8879), .ZN(n8853) );
  AND2_X1 U8772 ( .A1(n8850), .A2(n8849), .ZN(n8879) );
  AND2_X1 U8773 ( .A1(n8847), .A2(n8880), .ZN(n8878) );
  OR2_X1 U8774 ( .A1(n8849), .A2(n8850), .ZN(n8880) );
  OR2_X1 U8775 ( .A1(n7828), .A2(n8520), .ZN(n8850) );
  OR2_X1 U8776 ( .A1(n8881), .A2(n8882), .ZN(n8849) );
  AND2_X1 U8777 ( .A1(n8846), .A2(n8845), .ZN(n8882) );
  AND2_X1 U8778 ( .A1(n8843), .A2(n8883), .ZN(n8881) );
  OR2_X1 U8779 ( .A1(n8845), .A2(n8846), .ZN(n8883) );
  OR2_X1 U8780 ( .A1(n7887), .A2(n8520), .ZN(n8846) );
  OR2_X1 U8781 ( .A1(n8884), .A2(n8885), .ZN(n8845) );
  AND2_X1 U8782 ( .A1(n8842), .A2(n8841), .ZN(n8885) );
  AND2_X1 U8783 ( .A1(n8839), .A2(n8886), .ZN(n8884) );
  OR2_X1 U8784 ( .A1(n8841), .A2(n8842), .ZN(n8886) );
  OR2_X1 U8785 ( .A1(n7955), .A2(n8520), .ZN(n8842) );
  OR2_X1 U8786 ( .A1(n8887), .A2(n8888), .ZN(n8841) );
  AND2_X1 U8787 ( .A1(n8838), .A2(n8837), .ZN(n8888) );
  AND2_X1 U8788 ( .A1(n8835), .A2(n8889), .ZN(n8887) );
  OR2_X1 U8789 ( .A1(n8837), .A2(n8838), .ZN(n8889) );
  OR2_X1 U8790 ( .A1(n8025), .A2(n8520), .ZN(n8838) );
  OR2_X1 U8791 ( .A1(n8890), .A2(n8891), .ZN(n8837) );
  AND2_X1 U8792 ( .A1(n8834), .A2(n8833), .ZN(n8891) );
  AND2_X1 U8793 ( .A1(n8831), .A2(n8892), .ZN(n8890) );
  OR2_X1 U8794 ( .A1(n8833), .A2(n8834), .ZN(n8892) );
  OR2_X1 U8795 ( .A1(n8107), .A2(n8520), .ZN(n8834) );
  OR2_X1 U8796 ( .A1(n8893), .A2(n8894), .ZN(n8833) );
  AND2_X1 U8797 ( .A1(n8830), .A2(n8829), .ZN(n8894) );
  AND2_X1 U8798 ( .A1(n8827), .A2(n8895), .ZN(n8893) );
  OR2_X1 U8799 ( .A1(n8829), .A2(n8830), .ZN(n8895) );
  OR2_X1 U8800 ( .A1(n8191), .A2(n8520), .ZN(n8830) );
  OR2_X1 U8801 ( .A1(n8896), .A2(n8897), .ZN(n8829) );
  AND2_X1 U8802 ( .A1(n8826), .A2(n8825), .ZN(n8897) );
  AND2_X1 U8803 ( .A1(n8823), .A2(n8898), .ZN(n8896) );
  OR2_X1 U8804 ( .A1(n8825), .A2(n8826), .ZN(n8898) );
  OR2_X1 U8805 ( .A1(n8287), .A2(n8520), .ZN(n8826) );
  OR2_X1 U8806 ( .A1(n8899), .A2(n8900), .ZN(n8825) );
  AND2_X1 U8807 ( .A1(n8822), .A2(n8821), .ZN(n8900) );
  AND2_X1 U8808 ( .A1(n8819), .A2(n8901), .ZN(n8899) );
  OR2_X1 U8809 ( .A1(n8821), .A2(n8822), .ZN(n8901) );
  OR2_X1 U8810 ( .A1(n8608), .A2(n8520), .ZN(n8822) );
  OR2_X1 U8811 ( .A1(n8902), .A2(n8903), .ZN(n8821) );
  AND2_X1 U8812 ( .A1(n8818), .A2(n8817), .ZN(n8903) );
  AND2_X1 U8813 ( .A1(n8815), .A2(n8904), .ZN(n8902) );
  OR2_X1 U8814 ( .A1(n8817), .A2(n8818), .ZN(n8904) );
  OR2_X1 U8815 ( .A1(n8603), .A2(n8520), .ZN(n8818) );
  OR2_X1 U8816 ( .A1(n8905), .A2(n8906), .ZN(n8817) );
  AND2_X1 U8817 ( .A1(n8814), .A2(n8813), .ZN(n8906) );
  AND2_X1 U8818 ( .A1(n8811), .A2(n8907), .ZN(n8905) );
  OR2_X1 U8819 ( .A1(n8813), .A2(n8814), .ZN(n8907) );
  OR2_X1 U8820 ( .A1(n8598), .A2(n8520), .ZN(n8814) );
  OR2_X1 U8821 ( .A1(n8908), .A2(n8909), .ZN(n8813) );
  AND2_X1 U8822 ( .A1(n8810), .A2(n8809), .ZN(n8909) );
  AND2_X1 U8823 ( .A1(n8807), .A2(n8910), .ZN(n8908) );
  OR2_X1 U8824 ( .A1(n8809), .A2(n8810), .ZN(n8910) );
  OR2_X1 U8825 ( .A1(n8593), .A2(n8520), .ZN(n8810) );
  OR2_X1 U8826 ( .A1(n8911), .A2(n8912), .ZN(n8809) );
  AND2_X1 U8827 ( .A1(n8806), .A2(n8805), .ZN(n8912) );
  AND2_X1 U8828 ( .A1(n8803), .A2(n8913), .ZN(n8911) );
  OR2_X1 U8829 ( .A1(n8805), .A2(n8806), .ZN(n8913) );
  OR2_X1 U8830 ( .A1(n8588), .A2(n8520), .ZN(n8806) );
  OR2_X1 U8831 ( .A1(n8914), .A2(n8915), .ZN(n8805) );
  AND2_X1 U8832 ( .A1(n8802), .A2(n8801), .ZN(n8915) );
  AND2_X1 U8833 ( .A1(n8799), .A2(n8916), .ZN(n8914) );
  OR2_X1 U8834 ( .A1(n8801), .A2(n8802), .ZN(n8916) );
  OR2_X1 U8835 ( .A1(n8583), .A2(n8520), .ZN(n8802) );
  OR2_X1 U8836 ( .A1(n8917), .A2(n8918), .ZN(n8801) );
  AND2_X1 U8837 ( .A1(n8798), .A2(n8797), .ZN(n8918) );
  AND2_X1 U8838 ( .A1(n8795), .A2(n8919), .ZN(n8917) );
  OR2_X1 U8839 ( .A1(n8797), .A2(n8798), .ZN(n8919) );
  OR2_X1 U8840 ( .A1(n8578), .A2(n8520), .ZN(n8798) );
  OR2_X1 U8841 ( .A1(n8920), .A2(n8921), .ZN(n8797) );
  AND2_X1 U8842 ( .A1(n8794), .A2(n8793), .ZN(n8921) );
  AND2_X1 U8843 ( .A1(n8791), .A2(n8922), .ZN(n8920) );
  OR2_X1 U8844 ( .A1(n8793), .A2(n8794), .ZN(n8922) );
  OR2_X1 U8845 ( .A1(n8573), .A2(n8520), .ZN(n8794) );
  OR2_X1 U8846 ( .A1(n8923), .A2(n8924), .ZN(n8793) );
  AND2_X1 U8847 ( .A1(n8790), .A2(n8789), .ZN(n8924) );
  AND2_X1 U8848 ( .A1(n8787), .A2(n8925), .ZN(n8923) );
  OR2_X1 U8849 ( .A1(n8789), .A2(n8790), .ZN(n8925) );
  OR2_X1 U8850 ( .A1(n8568), .A2(n8520), .ZN(n8790) );
  OR2_X1 U8851 ( .A1(n8926), .A2(n8927), .ZN(n8789) );
  AND2_X1 U8852 ( .A1(n8786), .A2(n8785), .ZN(n8927) );
  AND2_X1 U8853 ( .A1(n8783), .A2(n8928), .ZN(n8926) );
  OR2_X1 U8854 ( .A1(n8785), .A2(n8786), .ZN(n8928) );
  OR2_X1 U8855 ( .A1(n8563), .A2(n8520), .ZN(n8786) );
  OR2_X1 U8856 ( .A1(n8929), .A2(n8930), .ZN(n8785) );
  AND2_X1 U8857 ( .A1(n8782), .A2(n8781), .ZN(n8930) );
  AND2_X1 U8858 ( .A1(n8779), .A2(n8931), .ZN(n8929) );
  OR2_X1 U8859 ( .A1(n8781), .A2(n8782), .ZN(n8931) );
  OR2_X1 U8860 ( .A1(n8558), .A2(n8520), .ZN(n8782) );
  OR2_X1 U8861 ( .A1(n8932), .A2(n8933), .ZN(n8781) );
  AND2_X1 U8862 ( .A1(n8778), .A2(n8777), .ZN(n8933) );
  AND2_X1 U8863 ( .A1(n8775), .A2(n8934), .ZN(n8932) );
  OR2_X1 U8864 ( .A1(n8777), .A2(n8778), .ZN(n8934) );
  OR2_X1 U8865 ( .A1(n8553), .A2(n8520), .ZN(n8778) );
  OR2_X1 U8866 ( .A1(n8935), .A2(n8936), .ZN(n8777) );
  AND2_X1 U8867 ( .A1(n8774), .A2(n8773), .ZN(n8936) );
  AND2_X1 U8868 ( .A1(n8771), .A2(n8937), .ZN(n8935) );
  OR2_X1 U8869 ( .A1(n8773), .A2(n8774), .ZN(n8937) );
  OR2_X1 U8870 ( .A1(n8548), .A2(n8520), .ZN(n8774) );
  OR2_X1 U8871 ( .A1(n8938), .A2(n8939), .ZN(n8773) );
  AND2_X1 U8872 ( .A1(n8770), .A2(n8769), .ZN(n8939) );
  AND2_X1 U8873 ( .A1(n8767), .A2(n8940), .ZN(n8938) );
  OR2_X1 U8874 ( .A1(n8769), .A2(n8770), .ZN(n8940) );
  OR2_X1 U8875 ( .A1(n8543), .A2(n8520), .ZN(n8770) );
  OR2_X1 U8876 ( .A1(n8941), .A2(n8942), .ZN(n8769) );
  AND2_X1 U8877 ( .A1(n8766), .A2(n8765), .ZN(n8942) );
  AND2_X1 U8878 ( .A1(n8763), .A2(n8943), .ZN(n8941) );
  OR2_X1 U8879 ( .A1(n8765), .A2(n8766), .ZN(n8943) );
  OR2_X1 U8880 ( .A1(n8538), .A2(n8520), .ZN(n8766) );
  OR2_X1 U8881 ( .A1(n8944), .A2(n8945), .ZN(n8765) );
  AND2_X1 U8882 ( .A1(n8762), .A2(n8761), .ZN(n8945) );
  AND2_X1 U8883 ( .A1(n8759), .A2(n8946), .ZN(n8944) );
  OR2_X1 U8884 ( .A1(n8761), .A2(n8762), .ZN(n8946) );
  OR2_X1 U8885 ( .A1(n8533), .A2(n8520), .ZN(n8762) );
  OR2_X1 U8886 ( .A1(n8947), .A2(n8948), .ZN(n8761) );
  AND2_X1 U8887 ( .A1(n8758), .A2(n8757), .ZN(n8948) );
  AND2_X1 U8888 ( .A1(n8755), .A2(n8949), .ZN(n8947) );
  OR2_X1 U8889 ( .A1(n8757), .A2(n8758), .ZN(n8949) );
  OR2_X1 U8890 ( .A1(n8528), .A2(n8520), .ZN(n8758) );
  OR2_X1 U8891 ( .A1(n8950), .A2(n8951), .ZN(n8757) );
  AND2_X1 U8892 ( .A1(n8754), .A2(n8753), .ZN(n8951) );
  AND2_X1 U8893 ( .A1(n8751), .A2(n8952), .ZN(n8950) );
  OR2_X1 U8894 ( .A1(n8753), .A2(n8754), .ZN(n8952) );
  OR2_X1 U8895 ( .A1(n8523), .A2(n8520), .ZN(n8754) );
  OR2_X1 U8896 ( .A1(n8953), .A2(n8954), .ZN(n8753) );
  AND2_X1 U8897 ( .A1(n8750), .A2(n8747), .ZN(n8954) );
  AND2_X1 U8898 ( .A1(n8955), .A2(n8749), .ZN(n8953) );
  OR2_X1 U8899 ( .A1(n8750), .A2(n8747), .ZN(n8955) );
  OR2_X1 U8900 ( .A1(n8744), .A2(n8739), .ZN(n8747) );
  OR2_X1 U8901 ( .A1(n8956), .A2(n8520), .ZN(n8739) );
  INV_X1 U8902 ( .A(n8957), .ZN(n8750) );
  OR2_X1 U8903 ( .A1(n8958), .A2(n8959), .ZN(n8957) );
  AND2_X1 U8904 ( .A1(b_28_), .A2(n8960), .ZN(n8959) );
  OR2_X1 U8905 ( .A1(n8961), .A2(n7343), .ZN(n8960) );
  AND2_X1 U8906 ( .A1(a_30_), .A2(n8962), .ZN(n8961) );
  AND2_X1 U8907 ( .A1(b_27_), .A2(n8963), .ZN(n8958) );
  OR2_X1 U8908 ( .A1(n8964), .A2(n7347), .ZN(n8963) );
  AND2_X1 U8909 ( .A1(a_31_), .A2(n8744), .ZN(n8964) );
  XOR2_X1 U8910 ( .A(n8965), .B(n8966), .Z(n8751) );
  XNOR2_X1 U8911 ( .A(n8967), .B(n8968), .ZN(n8965) );
  XNOR2_X1 U8912 ( .A(n8969), .B(n8970), .ZN(n8755) );
  XNOR2_X1 U8913 ( .A(n8971), .B(n8972), .ZN(n8969) );
  XOR2_X1 U8914 ( .A(n8973), .B(n8974), .Z(n8759) );
  XOR2_X1 U8915 ( .A(n8975), .B(n8976), .Z(n8974) );
  XOR2_X1 U8916 ( .A(n8977), .B(n8978), .Z(n8763) );
  XOR2_X1 U8917 ( .A(n8979), .B(n8980), .Z(n8978) );
  XOR2_X1 U8918 ( .A(n8981), .B(n8982), .Z(n8767) );
  XOR2_X1 U8919 ( .A(n8983), .B(n8984), .Z(n8982) );
  XOR2_X1 U8920 ( .A(n8985), .B(n8986), .Z(n8771) );
  XOR2_X1 U8921 ( .A(n8987), .B(n8988), .Z(n8986) );
  XOR2_X1 U8922 ( .A(n8989), .B(n8990), .Z(n8775) );
  XOR2_X1 U8923 ( .A(n8991), .B(n8992), .Z(n8990) );
  XOR2_X1 U8924 ( .A(n8993), .B(n8994), .Z(n8779) );
  XOR2_X1 U8925 ( .A(n8995), .B(n8996), .Z(n8994) );
  XOR2_X1 U8926 ( .A(n8997), .B(n8998), .Z(n8783) );
  XOR2_X1 U8927 ( .A(n8999), .B(n9000), .Z(n8998) );
  XOR2_X1 U8928 ( .A(n9001), .B(n9002), .Z(n8787) );
  XOR2_X1 U8929 ( .A(n9003), .B(n9004), .Z(n9002) );
  XOR2_X1 U8930 ( .A(n9005), .B(n9006), .Z(n8791) );
  XOR2_X1 U8931 ( .A(n9007), .B(n9008), .Z(n9006) );
  XOR2_X1 U8932 ( .A(n9009), .B(n9010), .Z(n8795) );
  XOR2_X1 U8933 ( .A(n9011), .B(n9012), .Z(n9010) );
  XOR2_X1 U8934 ( .A(n9013), .B(n9014), .Z(n8799) );
  XOR2_X1 U8935 ( .A(n9015), .B(n9016), .Z(n9014) );
  XOR2_X1 U8936 ( .A(n9017), .B(n9018), .Z(n8803) );
  XOR2_X1 U8937 ( .A(n9019), .B(n9020), .Z(n9018) );
  XOR2_X1 U8938 ( .A(n9021), .B(n9022), .Z(n8807) );
  XOR2_X1 U8939 ( .A(n9023), .B(n9024), .Z(n9022) );
  XOR2_X1 U8940 ( .A(n9025), .B(n9026), .Z(n8811) );
  XOR2_X1 U8941 ( .A(n9027), .B(n9028), .Z(n9026) );
  XOR2_X1 U8942 ( .A(n9029), .B(n9030), .Z(n8815) );
  XOR2_X1 U8943 ( .A(n9031), .B(n9032), .Z(n9030) );
  XOR2_X1 U8944 ( .A(n9033), .B(n9034), .Z(n8819) );
  XOR2_X1 U8945 ( .A(n9035), .B(n9036), .Z(n9034) );
  XOR2_X1 U8946 ( .A(n9037), .B(n9038), .Z(n8823) );
  XOR2_X1 U8947 ( .A(n9039), .B(n9040), .Z(n9038) );
  XOR2_X1 U8948 ( .A(n9041), .B(n9042), .Z(n8827) );
  XOR2_X1 U8949 ( .A(n9043), .B(n9044), .Z(n9042) );
  XOR2_X1 U8950 ( .A(n9045), .B(n9046), .Z(n8831) );
  XOR2_X1 U8951 ( .A(n9047), .B(n9048), .Z(n9046) );
  XOR2_X1 U8952 ( .A(n9049), .B(n9050), .Z(n8835) );
  XOR2_X1 U8953 ( .A(n9051), .B(n9052), .Z(n9050) );
  XOR2_X1 U8954 ( .A(n9053), .B(n9054), .Z(n8839) );
  XOR2_X1 U8955 ( .A(n9055), .B(n9056), .Z(n9054) );
  XOR2_X1 U8956 ( .A(n9057), .B(n9058), .Z(n8843) );
  XOR2_X1 U8957 ( .A(n9059), .B(n9060), .Z(n9058) );
  XOR2_X1 U8958 ( .A(n9061), .B(n9062), .Z(n8847) );
  XOR2_X1 U8959 ( .A(n9063), .B(n9064), .Z(n9062) );
  XOR2_X1 U8960 ( .A(n9065), .B(n9066), .Z(n8851) );
  XOR2_X1 U8961 ( .A(n9067), .B(n9068), .Z(n9066) );
  OR2_X1 U8962 ( .A1(n7730), .A2(n8520), .ZN(n8857) );
  XOR2_X1 U8963 ( .A(n9069), .B(n9070), .Z(n8856) );
  XOR2_X1 U8964 ( .A(n9071), .B(n9072), .Z(n9070) );
  XNOR2_X1 U8965 ( .A(n9073), .B(n9074), .ZN(n8420) );
  XNOR2_X1 U8966 ( .A(n9075), .B(n9076), .ZN(n9073) );
  XOR2_X1 U8967 ( .A(n9077), .B(n9078), .Z(n8409) );
  XOR2_X1 U8968 ( .A(n9079), .B(n9080), .Z(n9078) );
  OR2_X1 U8969 ( .A1(n8382), .A2(n8381), .ZN(n7504) );
  INV_X1 U8970 ( .A(n9081), .ZN(n8381) );
  OR2_X1 U8971 ( .A1(n9082), .A2(n8379), .ZN(n9081) );
  AND2_X1 U8972 ( .A1(n9083), .A2(n9084), .ZN(n9082) );
  AND2_X1 U8973 ( .A1(n8389), .A2(n8390), .ZN(n8382) );
  INV_X1 U8974 ( .A(n8861), .ZN(n8390) );
  OR2_X1 U8975 ( .A1(n9085), .A2(n9086), .ZN(n8861) );
  AND2_X1 U8976 ( .A1(n8865), .A2(n8864), .ZN(n9086) );
  AND2_X1 U8977 ( .A1(n8862), .A2(n9087), .ZN(n9085) );
  OR2_X1 U8978 ( .A1(n8864), .A2(n8865), .ZN(n9087) );
  OR2_X1 U8979 ( .A1(n7660), .A2(n8744), .ZN(n8865) );
  OR2_X1 U8980 ( .A1(n9088), .A2(n9089), .ZN(n8864) );
  AND2_X1 U8981 ( .A1(n9080), .A2(n9079), .ZN(n9089) );
  AND2_X1 U8982 ( .A1(n9077), .A2(n9090), .ZN(n9088) );
  OR2_X1 U8983 ( .A1(n9079), .A2(n9080), .ZN(n9090) );
  OR2_X1 U8984 ( .A1(n7697), .A2(n8744), .ZN(n9080) );
  OR2_X1 U8985 ( .A1(n9091), .A2(n9092), .ZN(n9079) );
  AND2_X1 U8986 ( .A1(n9076), .A2(n9075), .ZN(n9092) );
  AND2_X1 U8987 ( .A1(n9074), .A2(n9093), .ZN(n9091) );
  OR2_X1 U8988 ( .A1(n9075), .A2(n9076), .ZN(n9093) );
  OR2_X1 U8989 ( .A1(n9094), .A2(n9095), .ZN(n9076) );
  AND2_X1 U8990 ( .A1(n9072), .A2(n9071), .ZN(n9095) );
  AND2_X1 U8991 ( .A1(n9069), .A2(n9096), .ZN(n9094) );
  OR2_X1 U8992 ( .A1(n9071), .A2(n9072), .ZN(n9096) );
  OR2_X1 U8993 ( .A1(n7820), .A2(n8744), .ZN(n9072) );
  OR2_X1 U8994 ( .A1(n9097), .A2(n9098), .ZN(n9071) );
  AND2_X1 U8995 ( .A1(n9068), .A2(n9067), .ZN(n9098) );
  AND2_X1 U8996 ( .A1(n9065), .A2(n9099), .ZN(n9097) );
  OR2_X1 U8997 ( .A1(n9067), .A2(n9068), .ZN(n9099) );
  OR2_X1 U8998 ( .A1(n7828), .A2(n8744), .ZN(n9068) );
  OR2_X1 U8999 ( .A1(n9100), .A2(n9101), .ZN(n9067) );
  AND2_X1 U9000 ( .A1(n9064), .A2(n9063), .ZN(n9101) );
  AND2_X1 U9001 ( .A1(n9061), .A2(n9102), .ZN(n9100) );
  OR2_X1 U9002 ( .A1(n9063), .A2(n9064), .ZN(n9102) );
  OR2_X1 U9003 ( .A1(n7887), .A2(n8744), .ZN(n9064) );
  OR2_X1 U9004 ( .A1(n9103), .A2(n9104), .ZN(n9063) );
  AND2_X1 U9005 ( .A1(n9060), .A2(n9059), .ZN(n9104) );
  AND2_X1 U9006 ( .A1(n9057), .A2(n9105), .ZN(n9103) );
  OR2_X1 U9007 ( .A1(n9059), .A2(n9060), .ZN(n9105) );
  OR2_X1 U9008 ( .A1(n7955), .A2(n8744), .ZN(n9060) );
  OR2_X1 U9009 ( .A1(n9106), .A2(n9107), .ZN(n9059) );
  AND2_X1 U9010 ( .A1(n9056), .A2(n9055), .ZN(n9107) );
  AND2_X1 U9011 ( .A1(n9053), .A2(n9108), .ZN(n9106) );
  OR2_X1 U9012 ( .A1(n9055), .A2(n9056), .ZN(n9108) );
  OR2_X1 U9013 ( .A1(n8025), .A2(n8744), .ZN(n9056) );
  OR2_X1 U9014 ( .A1(n9109), .A2(n9110), .ZN(n9055) );
  AND2_X1 U9015 ( .A1(n9052), .A2(n9051), .ZN(n9110) );
  AND2_X1 U9016 ( .A1(n9049), .A2(n9111), .ZN(n9109) );
  OR2_X1 U9017 ( .A1(n9051), .A2(n9052), .ZN(n9111) );
  OR2_X1 U9018 ( .A1(n8107), .A2(n8744), .ZN(n9052) );
  OR2_X1 U9019 ( .A1(n9112), .A2(n9113), .ZN(n9051) );
  AND2_X1 U9020 ( .A1(n9048), .A2(n9047), .ZN(n9113) );
  AND2_X1 U9021 ( .A1(n9045), .A2(n9114), .ZN(n9112) );
  OR2_X1 U9022 ( .A1(n9047), .A2(n9048), .ZN(n9114) );
  OR2_X1 U9023 ( .A1(n8191), .A2(n8744), .ZN(n9048) );
  OR2_X1 U9024 ( .A1(n9115), .A2(n9116), .ZN(n9047) );
  AND2_X1 U9025 ( .A1(n9044), .A2(n9043), .ZN(n9116) );
  AND2_X1 U9026 ( .A1(n9041), .A2(n9117), .ZN(n9115) );
  OR2_X1 U9027 ( .A1(n9043), .A2(n9044), .ZN(n9117) );
  OR2_X1 U9028 ( .A1(n8287), .A2(n8744), .ZN(n9044) );
  OR2_X1 U9029 ( .A1(n9118), .A2(n9119), .ZN(n9043) );
  AND2_X1 U9030 ( .A1(n9040), .A2(n9039), .ZN(n9119) );
  AND2_X1 U9031 ( .A1(n9037), .A2(n9120), .ZN(n9118) );
  OR2_X1 U9032 ( .A1(n9039), .A2(n9040), .ZN(n9120) );
  OR2_X1 U9033 ( .A1(n8608), .A2(n8744), .ZN(n9040) );
  OR2_X1 U9034 ( .A1(n9121), .A2(n9122), .ZN(n9039) );
  AND2_X1 U9035 ( .A1(n9036), .A2(n9035), .ZN(n9122) );
  AND2_X1 U9036 ( .A1(n9033), .A2(n9123), .ZN(n9121) );
  OR2_X1 U9037 ( .A1(n9035), .A2(n9036), .ZN(n9123) );
  OR2_X1 U9038 ( .A1(n8603), .A2(n8744), .ZN(n9036) );
  OR2_X1 U9039 ( .A1(n9124), .A2(n9125), .ZN(n9035) );
  AND2_X1 U9040 ( .A1(n9032), .A2(n9031), .ZN(n9125) );
  AND2_X1 U9041 ( .A1(n9029), .A2(n9126), .ZN(n9124) );
  OR2_X1 U9042 ( .A1(n9031), .A2(n9032), .ZN(n9126) );
  OR2_X1 U9043 ( .A1(n8598), .A2(n8744), .ZN(n9032) );
  OR2_X1 U9044 ( .A1(n9127), .A2(n9128), .ZN(n9031) );
  AND2_X1 U9045 ( .A1(n9028), .A2(n9027), .ZN(n9128) );
  AND2_X1 U9046 ( .A1(n9025), .A2(n9129), .ZN(n9127) );
  OR2_X1 U9047 ( .A1(n9027), .A2(n9028), .ZN(n9129) );
  OR2_X1 U9048 ( .A1(n8593), .A2(n8744), .ZN(n9028) );
  OR2_X1 U9049 ( .A1(n9130), .A2(n9131), .ZN(n9027) );
  AND2_X1 U9050 ( .A1(n9024), .A2(n9023), .ZN(n9131) );
  AND2_X1 U9051 ( .A1(n9021), .A2(n9132), .ZN(n9130) );
  OR2_X1 U9052 ( .A1(n9023), .A2(n9024), .ZN(n9132) );
  OR2_X1 U9053 ( .A1(n8588), .A2(n8744), .ZN(n9024) );
  OR2_X1 U9054 ( .A1(n9133), .A2(n9134), .ZN(n9023) );
  AND2_X1 U9055 ( .A1(n9020), .A2(n9019), .ZN(n9134) );
  AND2_X1 U9056 ( .A1(n9017), .A2(n9135), .ZN(n9133) );
  OR2_X1 U9057 ( .A1(n9019), .A2(n9020), .ZN(n9135) );
  OR2_X1 U9058 ( .A1(n8583), .A2(n8744), .ZN(n9020) );
  OR2_X1 U9059 ( .A1(n9136), .A2(n9137), .ZN(n9019) );
  AND2_X1 U9060 ( .A1(n9016), .A2(n9015), .ZN(n9137) );
  AND2_X1 U9061 ( .A1(n9013), .A2(n9138), .ZN(n9136) );
  OR2_X1 U9062 ( .A1(n9015), .A2(n9016), .ZN(n9138) );
  OR2_X1 U9063 ( .A1(n8578), .A2(n8744), .ZN(n9016) );
  OR2_X1 U9064 ( .A1(n9139), .A2(n9140), .ZN(n9015) );
  AND2_X1 U9065 ( .A1(n9012), .A2(n9011), .ZN(n9140) );
  AND2_X1 U9066 ( .A1(n9009), .A2(n9141), .ZN(n9139) );
  OR2_X1 U9067 ( .A1(n9011), .A2(n9012), .ZN(n9141) );
  OR2_X1 U9068 ( .A1(n8573), .A2(n8744), .ZN(n9012) );
  OR2_X1 U9069 ( .A1(n9142), .A2(n9143), .ZN(n9011) );
  AND2_X1 U9070 ( .A1(n9008), .A2(n9007), .ZN(n9143) );
  AND2_X1 U9071 ( .A1(n9005), .A2(n9144), .ZN(n9142) );
  OR2_X1 U9072 ( .A1(n9007), .A2(n9008), .ZN(n9144) );
  OR2_X1 U9073 ( .A1(n8568), .A2(n8744), .ZN(n9008) );
  OR2_X1 U9074 ( .A1(n9145), .A2(n9146), .ZN(n9007) );
  AND2_X1 U9075 ( .A1(n9004), .A2(n9003), .ZN(n9146) );
  AND2_X1 U9076 ( .A1(n9001), .A2(n9147), .ZN(n9145) );
  OR2_X1 U9077 ( .A1(n9003), .A2(n9004), .ZN(n9147) );
  OR2_X1 U9078 ( .A1(n8563), .A2(n8744), .ZN(n9004) );
  OR2_X1 U9079 ( .A1(n9148), .A2(n9149), .ZN(n9003) );
  AND2_X1 U9080 ( .A1(n9000), .A2(n8999), .ZN(n9149) );
  AND2_X1 U9081 ( .A1(n8997), .A2(n9150), .ZN(n9148) );
  OR2_X1 U9082 ( .A1(n8999), .A2(n9000), .ZN(n9150) );
  OR2_X1 U9083 ( .A1(n8558), .A2(n8744), .ZN(n9000) );
  OR2_X1 U9084 ( .A1(n9151), .A2(n9152), .ZN(n8999) );
  AND2_X1 U9085 ( .A1(n8996), .A2(n8995), .ZN(n9152) );
  AND2_X1 U9086 ( .A1(n8993), .A2(n9153), .ZN(n9151) );
  OR2_X1 U9087 ( .A1(n8995), .A2(n8996), .ZN(n9153) );
  OR2_X1 U9088 ( .A1(n8553), .A2(n8744), .ZN(n8996) );
  OR2_X1 U9089 ( .A1(n9154), .A2(n9155), .ZN(n8995) );
  AND2_X1 U9090 ( .A1(n8992), .A2(n8991), .ZN(n9155) );
  AND2_X1 U9091 ( .A1(n8989), .A2(n9156), .ZN(n9154) );
  OR2_X1 U9092 ( .A1(n8991), .A2(n8992), .ZN(n9156) );
  OR2_X1 U9093 ( .A1(n8548), .A2(n8744), .ZN(n8992) );
  OR2_X1 U9094 ( .A1(n9157), .A2(n9158), .ZN(n8991) );
  AND2_X1 U9095 ( .A1(n8988), .A2(n8987), .ZN(n9158) );
  AND2_X1 U9096 ( .A1(n8985), .A2(n9159), .ZN(n9157) );
  OR2_X1 U9097 ( .A1(n8987), .A2(n8988), .ZN(n9159) );
  OR2_X1 U9098 ( .A1(n8543), .A2(n8744), .ZN(n8988) );
  OR2_X1 U9099 ( .A1(n9160), .A2(n9161), .ZN(n8987) );
  AND2_X1 U9100 ( .A1(n8984), .A2(n8983), .ZN(n9161) );
  AND2_X1 U9101 ( .A1(n8981), .A2(n9162), .ZN(n9160) );
  OR2_X1 U9102 ( .A1(n8983), .A2(n8984), .ZN(n9162) );
  OR2_X1 U9103 ( .A1(n8538), .A2(n8744), .ZN(n8984) );
  OR2_X1 U9104 ( .A1(n9163), .A2(n9164), .ZN(n8983) );
  AND2_X1 U9105 ( .A1(n8980), .A2(n8979), .ZN(n9164) );
  AND2_X1 U9106 ( .A1(n8977), .A2(n9165), .ZN(n9163) );
  OR2_X1 U9107 ( .A1(n8979), .A2(n8980), .ZN(n9165) );
  OR2_X1 U9108 ( .A1(n8533), .A2(n8744), .ZN(n8980) );
  OR2_X1 U9109 ( .A1(n9166), .A2(n9167), .ZN(n8979) );
  AND2_X1 U9110 ( .A1(n8976), .A2(n8975), .ZN(n9167) );
  AND2_X1 U9111 ( .A1(n8973), .A2(n9168), .ZN(n9166) );
  OR2_X1 U9112 ( .A1(n8975), .A2(n8976), .ZN(n9168) );
  OR2_X1 U9113 ( .A1(n8528), .A2(n8744), .ZN(n8976) );
  OR2_X1 U9114 ( .A1(n9169), .A2(n9170), .ZN(n8975) );
  AND2_X1 U9115 ( .A1(n8970), .A2(n8972), .ZN(n9170) );
  AND2_X1 U9116 ( .A1(n9171), .A2(n8971), .ZN(n9169) );
  OR2_X1 U9117 ( .A1(n8972), .A2(n8970), .ZN(n9171) );
  XOR2_X1 U9118 ( .A(n9172), .B(n9173), .Z(n8970) );
  XNOR2_X1 U9119 ( .A(n9174), .B(n9175), .ZN(n9172) );
  OR2_X1 U9120 ( .A1(n9176), .A2(n9177), .ZN(n8972) );
  AND2_X1 U9121 ( .A1(n8966), .A2(n8967), .ZN(n9177) );
  AND2_X1 U9122 ( .A1(n9178), .A2(n9179), .ZN(n9176) );
  OR2_X1 U9123 ( .A1(n8967), .A2(n8966), .ZN(n9179) );
  OR2_X1 U9124 ( .A1(n8515), .A2(n8744), .ZN(n8966) );
  OR2_X1 U9125 ( .A1(n8962), .A2(n9180), .ZN(n8967) );
  OR2_X1 U9126 ( .A1(n8956), .A2(n8744), .ZN(n9180) );
  INV_X1 U9127 ( .A(n8968), .ZN(n9178) );
  OR2_X1 U9128 ( .A1(n9181), .A2(n9182), .ZN(n8968) );
  AND2_X1 U9129 ( .A1(b_27_), .A2(n9183), .ZN(n9182) );
  OR2_X1 U9130 ( .A1(n9184), .A2(n7343), .ZN(n9183) );
  AND2_X1 U9131 ( .A1(a_30_), .A2(n9185), .ZN(n9184) );
  AND2_X1 U9132 ( .A1(b_26_), .A2(n9186), .ZN(n9181) );
  OR2_X1 U9133 ( .A1(n9187), .A2(n7347), .ZN(n9186) );
  AND2_X1 U9134 ( .A1(a_31_), .A2(n8962), .ZN(n9187) );
  XOR2_X1 U9135 ( .A(n9188), .B(n9189), .Z(n8973) );
  XOR2_X1 U9136 ( .A(n9190), .B(n9191), .Z(n9189) );
  XNOR2_X1 U9137 ( .A(n9192), .B(n9193), .ZN(n8977) );
  XNOR2_X1 U9138 ( .A(n9194), .B(n9195), .ZN(n9192) );
  XOR2_X1 U9139 ( .A(n9196), .B(n9197), .Z(n8981) );
  XOR2_X1 U9140 ( .A(n9198), .B(n9199), .Z(n9197) );
  XOR2_X1 U9141 ( .A(n9200), .B(n9201), .Z(n8985) );
  XOR2_X1 U9142 ( .A(n9202), .B(n9203), .Z(n9201) );
  XOR2_X1 U9143 ( .A(n9204), .B(n9205), .Z(n8989) );
  XOR2_X1 U9144 ( .A(n9206), .B(n9207), .Z(n9205) );
  XOR2_X1 U9145 ( .A(n9208), .B(n9209), .Z(n8993) );
  XOR2_X1 U9146 ( .A(n9210), .B(n9211), .Z(n9209) );
  XOR2_X1 U9147 ( .A(n9212), .B(n9213), .Z(n8997) );
  XOR2_X1 U9148 ( .A(n9214), .B(n9215), .Z(n9213) );
  XOR2_X1 U9149 ( .A(n9216), .B(n9217), .Z(n9001) );
  XOR2_X1 U9150 ( .A(n9218), .B(n9219), .Z(n9217) );
  XOR2_X1 U9151 ( .A(n9220), .B(n9221), .Z(n9005) );
  XOR2_X1 U9152 ( .A(n9222), .B(n9223), .Z(n9221) );
  XOR2_X1 U9153 ( .A(n9224), .B(n9225), .Z(n9009) );
  XOR2_X1 U9154 ( .A(n9226), .B(n9227), .Z(n9225) );
  XOR2_X1 U9155 ( .A(n9228), .B(n9229), .Z(n9013) );
  XOR2_X1 U9156 ( .A(n9230), .B(n9231), .Z(n9229) );
  XOR2_X1 U9157 ( .A(n9232), .B(n9233), .Z(n9017) );
  XOR2_X1 U9158 ( .A(n9234), .B(n9235), .Z(n9233) );
  XOR2_X1 U9159 ( .A(n9236), .B(n9237), .Z(n9021) );
  XOR2_X1 U9160 ( .A(n9238), .B(n9239), .Z(n9237) );
  XOR2_X1 U9161 ( .A(n9240), .B(n9241), .Z(n9025) );
  XOR2_X1 U9162 ( .A(n9242), .B(n9243), .Z(n9241) );
  XOR2_X1 U9163 ( .A(n9244), .B(n9245), .Z(n9029) );
  XOR2_X1 U9164 ( .A(n9246), .B(n9247), .Z(n9245) );
  XOR2_X1 U9165 ( .A(n9248), .B(n9249), .Z(n9033) );
  XOR2_X1 U9166 ( .A(n9250), .B(n9251), .Z(n9249) );
  XOR2_X1 U9167 ( .A(n9252), .B(n9253), .Z(n9037) );
  XOR2_X1 U9168 ( .A(n9254), .B(n9255), .Z(n9253) );
  XOR2_X1 U9169 ( .A(n9256), .B(n9257), .Z(n9041) );
  XOR2_X1 U9170 ( .A(n9258), .B(n9259), .Z(n9257) );
  XOR2_X1 U9171 ( .A(n9260), .B(n9261), .Z(n9045) );
  XOR2_X1 U9172 ( .A(n9262), .B(n9263), .Z(n9261) );
  XOR2_X1 U9173 ( .A(n9264), .B(n9265), .Z(n9049) );
  XOR2_X1 U9174 ( .A(n9266), .B(n9267), .Z(n9265) );
  XOR2_X1 U9175 ( .A(n9268), .B(n9269), .Z(n9053) );
  XOR2_X1 U9176 ( .A(n9270), .B(n9271), .Z(n9269) );
  XOR2_X1 U9177 ( .A(n9272), .B(n9273), .Z(n9057) );
  XOR2_X1 U9178 ( .A(n9274), .B(n9275), .Z(n9273) );
  XNOR2_X1 U9179 ( .A(n9276), .B(n9277), .ZN(n9061) );
  XNOR2_X1 U9180 ( .A(n9278), .B(n9279), .ZN(n9276) );
  XOR2_X1 U9181 ( .A(n9280), .B(n9281), .Z(n9065) );
  XOR2_X1 U9182 ( .A(n9282), .B(n9283), .Z(n9281) );
  XOR2_X1 U9183 ( .A(n9284), .B(n9285), .Z(n9069) );
  XOR2_X1 U9184 ( .A(n9286), .B(n9287), .Z(n9285) );
  OR2_X1 U9185 ( .A1(n7730), .A2(n8744), .ZN(n9075) );
  XOR2_X1 U9186 ( .A(n9288), .B(n9289), .Z(n9074) );
  XOR2_X1 U9187 ( .A(n9290), .B(n9291), .Z(n9289) );
  XNOR2_X1 U9188 ( .A(n9292), .B(n9293), .ZN(n9077) );
  XNOR2_X1 U9189 ( .A(n9294), .B(n9295), .ZN(n9292) );
  XOR2_X1 U9190 ( .A(n9296), .B(n9297), .Z(n8862) );
  XOR2_X1 U9191 ( .A(n9298), .B(n9299), .Z(n9297) );
  XNOR2_X1 U9192 ( .A(n9300), .B(n9301), .ZN(n8389) );
  XOR2_X1 U9193 ( .A(n9302), .B(n9303), .Z(n9301) );
  OR2_X1 U9194 ( .A1(n8379), .A2(n8378), .ZN(n7509) );
  XOR2_X1 U9195 ( .A(n8375), .B(n8376), .Z(n8378) );
  OR2_X1 U9196 ( .A1(n9304), .A2(n9305), .ZN(n8376) );
  AND2_X1 U9197 ( .A1(n9306), .A2(n9307), .ZN(n9305) );
  AND2_X1 U9198 ( .A1(n9308), .A2(n9309), .ZN(n9304) );
  OR2_X1 U9199 ( .A1(n9306), .A2(n9307), .ZN(n9309) );
  XOR2_X1 U9200 ( .A(n8369), .B(n9310), .Z(n8375) );
  XOR2_X1 U9201 ( .A(n8368), .B(n8367), .Z(n9310) );
  OR2_X1 U9202 ( .A1(n7660), .A2(n9311), .ZN(n8367) );
  OR2_X1 U9203 ( .A1(n9312), .A2(n9313), .ZN(n8368) );
  AND2_X1 U9204 ( .A1(n9314), .A2(n9315), .ZN(n9313) );
  AND2_X1 U9205 ( .A1(n9316), .A2(n9317), .ZN(n9312) );
  OR2_X1 U9206 ( .A1(n9314), .A2(n9315), .ZN(n9317) );
  XNOR2_X1 U9207 ( .A(n9318), .B(n9319), .ZN(n8369) );
  XNOR2_X1 U9208 ( .A(n9320), .B(n9321), .ZN(n9318) );
  INV_X1 U9209 ( .A(n9322), .ZN(n8379) );
  OR2_X1 U9210 ( .A1(n9083), .A2(n9084), .ZN(n9322) );
  OR2_X1 U9211 ( .A1(n9323), .A2(n9324), .ZN(n9084) );
  AND2_X1 U9212 ( .A1(n9300), .A2(n9303), .ZN(n9324) );
  AND2_X1 U9213 ( .A1(n9325), .A2(n9302), .ZN(n9323) );
  OR2_X1 U9214 ( .A1(n9326), .A2(n9327), .ZN(n9302) );
  AND2_X1 U9215 ( .A1(n9299), .A2(n9298), .ZN(n9327) );
  AND2_X1 U9216 ( .A1(n9296), .A2(n9328), .ZN(n9326) );
  OR2_X1 U9217 ( .A1(n9298), .A2(n9299), .ZN(n9328) );
  OR2_X1 U9218 ( .A1(n7697), .A2(n8962), .ZN(n9299) );
  OR2_X1 U9219 ( .A1(n9329), .A2(n9330), .ZN(n9298) );
  AND2_X1 U9220 ( .A1(n9295), .A2(n9294), .ZN(n9330) );
  AND2_X1 U9221 ( .A1(n9293), .A2(n9331), .ZN(n9329) );
  OR2_X1 U9222 ( .A1(n9294), .A2(n9295), .ZN(n9331) );
  OR2_X1 U9223 ( .A1(n9332), .A2(n9333), .ZN(n9295) );
  AND2_X1 U9224 ( .A1(n9291), .A2(n9290), .ZN(n9333) );
  AND2_X1 U9225 ( .A1(n9288), .A2(n9334), .ZN(n9332) );
  OR2_X1 U9226 ( .A1(n9290), .A2(n9291), .ZN(n9334) );
  OR2_X1 U9227 ( .A1(n7820), .A2(n8962), .ZN(n9291) );
  OR2_X1 U9228 ( .A1(n9335), .A2(n9336), .ZN(n9290) );
  AND2_X1 U9229 ( .A1(n9287), .A2(n9286), .ZN(n9336) );
  AND2_X1 U9230 ( .A1(n9284), .A2(n9337), .ZN(n9335) );
  OR2_X1 U9231 ( .A1(n9286), .A2(n9287), .ZN(n9337) );
  OR2_X1 U9232 ( .A1(n7828), .A2(n8962), .ZN(n9287) );
  OR2_X1 U9233 ( .A1(n9338), .A2(n9339), .ZN(n9286) );
  AND2_X1 U9234 ( .A1(n9283), .A2(n9282), .ZN(n9339) );
  AND2_X1 U9235 ( .A1(n9280), .A2(n9340), .ZN(n9338) );
  OR2_X1 U9236 ( .A1(n9282), .A2(n9283), .ZN(n9340) );
  OR2_X1 U9237 ( .A1(n7887), .A2(n8962), .ZN(n9283) );
  OR2_X1 U9238 ( .A1(n9341), .A2(n9342), .ZN(n9282) );
  AND2_X1 U9239 ( .A1(n9279), .A2(n9278), .ZN(n9342) );
  AND2_X1 U9240 ( .A1(n9277), .A2(n9343), .ZN(n9341) );
  OR2_X1 U9241 ( .A1(n9278), .A2(n9279), .ZN(n9343) );
  OR2_X1 U9242 ( .A1(n9344), .A2(n9345), .ZN(n9279) );
  AND2_X1 U9243 ( .A1(n9275), .A2(n9274), .ZN(n9345) );
  AND2_X1 U9244 ( .A1(n9272), .A2(n9346), .ZN(n9344) );
  OR2_X1 U9245 ( .A1(n9274), .A2(n9275), .ZN(n9346) );
  OR2_X1 U9246 ( .A1(n8025), .A2(n8962), .ZN(n9275) );
  OR2_X1 U9247 ( .A1(n9347), .A2(n9348), .ZN(n9274) );
  AND2_X1 U9248 ( .A1(n9271), .A2(n9270), .ZN(n9348) );
  AND2_X1 U9249 ( .A1(n9268), .A2(n9349), .ZN(n9347) );
  OR2_X1 U9250 ( .A1(n9270), .A2(n9271), .ZN(n9349) );
  OR2_X1 U9251 ( .A1(n8107), .A2(n8962), .ZN(n9271) );
  OR2_X1 U9252 ( .A1(n9350), .A2(n9351), .ZN(n9270) );
  AND2_X1 U9253 ( .A1(n9267), .A2(n9266), .ZN(n9351) );
  AND2_X1 U9254 ( .A1(n9264), .A2(n9352), .ZN(n9350) );
  OR2_X1 U9255 ( .A1(n9266), .A2(n9267), .ZN(n9352) );
  OR2_X1 U9256 ( .A1(n8191), .A2(n8962), .ZN(n9267) );
  OR2_X1 U9257 ( .A1(n9353), .A2(n9354), .ZN(n9266) );
  AND2_X1 U9258 ( .A1(n9263), .A2(n9262), .ZN(n9354) );
  AND2_X1 U9259 ( .A1(n9260), .A2(n9355), .ZN(n9353) );
  OR2_X1 U9260 ( .A1(n9262), .A2(n9263), .ZN(n9355) );
  OR2_X1 U9261 ( .A1(n8287), .A2(n8962), .ZN(n9263) );
  OR2_X1 U9262 ( .A1(n9356), .A2(n9357), .ZN(n9262) );
  AND2_X1 U9263 ( .A1(n9259), .A2(n9258), .ZN(n9357) );
  AND2_X1 U9264 ( .A1(n9256), .A2(n9358), .ZN(n9356) );
  OR2_X1 U9265 ( .A1(n9258), .A2(n9259), .ZN(n9358) );
  OR2_X1 U9266 ( .A1(n8608), .A2(n8962), .ZN(n9259) );
  OR2_X1 U9267 ( .A1(n9359), .A2(n9360), .ZN(n9258) );
  AND2_X1 U9268 ( .A1(n9255), .A2(n9254), .ZN(n9360) );
  AND2_X1 U9269 ( .A1(n9252), .A2(n9361), .ZN(n9359) );
  OR2_X1 U9270 ( .A1(n9254), .A2(n9255), .ZN(n9361) );
  OR2_X1 U9271 ( .A1(n8603), .A2(n8962), .ZN(n9255) );
  OR2_X1 U9272 ( .A1(n9362), .A2(n9363), .ZN(n9254) );
  AND2_X1 U9273 ( .A1(n9251), .A2(n9250), .ZN(n9363) );
  AND2_X1 U9274 ( .A1(n9248), .A2(n9364), .ZN(n9362) );
  OR2_X1 U9275 ( .A1(n9250), .A2(n9251), .ZN(n9364) );
  OR2_X1 U9276 ( .A1(n8598), .A2(n8962), .ZN(n9251) );
  OR2_X1 U9277 ( .A1(n9365), .A2(n9366), .ZN(n9250) );
  AND2_X1 U9278 ( .A1(n9247), .A2(n9246), .ZN(n9366) );
  AND2_X1 U9279 ( .A1(n9244), .A2(n9367), .ZN(n9365) );
  OR2_X1 U9280 ( .A1(n9246), .A2(n9247), .ZN(n9367) );
  OR2_X1 U9281 ( .A1(n8593), .A2(n8962), .ZN(n9247) );
  OR2_X1 U9282 ( .A1(n9368), .A2(n9369), .ZN(n9246) );
  AND2_X1 U9283 ( .A1(n9243), .A2(n9242), .ZN(n9369) );
  AND2_X1 U9284 ( .A1(n9240), .A2(n9370), .ZN(n9368) );
  OR2_X1 U9285 ( .A1(n9242), .A2(n9243), .ZN(n9370) );
  OR2_X1 U9286 ( .A1(n8588), .A2(n8962), .ZN(n9243) );
  OR2_X1 U9287 ( .A1(n9371), .A2(n9372), .ZN(n9242) );
  AND2_X1 U9288 ( .A1(n9239), .A2(n9238), .ZN(n9372) );
  AND2_X1 U9289 ( .A1(n9236), .A2(n9373), .ZN(n9371) );
  OR2_X1 U9290 ( .A1(n9238), .A2(n9239), .ZN(n9373) );
  OR2_X1 U9291 ( .A1(n8583), .A2(n8962), .ZN(n9239) );
  OR2_X1 U9292 ( .A1(n9374), .A2(n9375), .ZN(n9238) );
  AND2_X1 U9293 ( .A1(n9235), .A2(n9234), .ZN(n9375) );
  AND2_X1 U9294 ( .A1(n9232), .A2(n9376), .ZN(n9374) );
  OR2_X1 U9295 ( .A1(n9234), .A2(n9235), .ZN(n9376) );
  OR2_X1 U9296 ( .A1(n8578), .A2(n8962), .ZN(n9235) );
  OR2_X1 U9297 ( .A1(n9377), .A2(n9378), .ZN(n9234) );
  AND2_X1 U9298 ( .A1(n9231), .A2(n9230), .ZN(n9378) );
  AND2_X1 U9299 ( .A1(n9228), .A2(n9379), .ZN(n9377) );
  OR2_X1 U9300 ( .A1(n9230), .A2(n9231), .ZN(n9379) );
  OR2_X1 U9301 ( .A1(n8573), .A2(n8962), .ZN(n9231) );
  OR2_X1 U9302 ( .A1(n9380), .A2(n9381), .ZN(n9230) );
  AND2_X1 U9303 ( .A1(n9227), .A2(n9226), .ZN(n9381) );
  AND2_X1 U9304 ( .A1(n9224), .A2(n9382), .ZN(n9380) );
  OR2_X1 U9305 ( .A1(n9226), .A2(n9227), .ZN(n9382) );
  OR2_X1 U9306 ( .A1(n8568), .A2(n8962), .ZN(n9227) );
  OR2_X1 U9307 ( .A1(n9383), .A2(n9384), .ZN(n9226) );
  AND2_X1 U9308 ( .A1(n9223), .A2(n9222), .ZN(n9384) );
  AND2_X1 U9309 ( .A1(n9220), .A2(n9385), .ZN(n9383) );
  OR2_X1 U9310 ( .A1(n9222), .A2(n9223), .ZN(n9385) );
  OR2_X1 U9311 ( .A1(n8563), .A2(n8962), .ZN(n9223) );
  OR2_X1 U9312 ( .A1(n9386), .A2(n9387), .ZN(n9222) );
  AND2_X1 U9313 ( .A1(n9219), .A2(n9218), .ZN(n9387) );
  AND2_X1 U9314 ( .A1(n9216), .A2(n9388), .ZN(n9386) );
  OR2_X1 U9315 ( .A1(n9218), .A2(n9219), .ZN(n9388) );
  OR2_X1 U9316 ( .A1(n8558), .A2(n8962), .ZN(n9219) );
  OR2_X1 U9317 ( .A1(n9389), .A2(n9390), .ZN(n9218) );
  AND2_X1 U9318 ( .A1(n9215), .A2(n9214), .ZN(n9390) );
  AND2_X1 U9319 ( .A1(n9212), .A2(n9391), .ZN(n9389) );
  OR2_X1 U9320 ( .A1(n9214), .A2(n9215), .ZN(n9391) );
  OR2_X1 U9321 ( .A1(n8553), .A2(n8962), .ZN(n9215) );
  OR2_X1 U9322 ( .A1(n9392), .A2(n9393), .ZN(n9214) );
  AND2_X1 U9323 ( .A1(n9211), .A2(n9210), .ZN(n9393) );
  AND2_X1 U9324 ( .A1(n9208), .A2(n9394), .ZN(n9392) );
  OR2_X1 U9325 ( .A1(n9210), .A2(n9211), .ZN(n9394) );
  OR2_X1 U9326 ( .A1(n8548), .A2(n8962), .ZN(n9211) );
  OR2_X1 U9327 ( .A1(n9395), .A2(n9396), .ZN(n9210) );
  AND2_X1 U9328 ( .A1(n9207), .A2(n9206), .ZN(n9396) );
  AND2_X1 U9329 ( .A1(n9204), .A2(n9397), .ZN(n9395) );
  OR2_X1 U9330 ( .A1(n9206), .A2(n9207), .ZN(n9397) );
  OR2_X1 U9331 ( .A1(n8543), .A2(n8962), .ZN(n9207) );
  OR2_X1 U9332 ( .A1(n9398), .A2(n9399), .ZN(n9206) );
  AND2_X1 U9333 ( .A1(n9203), .A2(n9202), .ZN(n9399) );
  AND2_X1 U9334 ( .A1(n9200), .A2(n9400), .ZN(n9398) );
  OR2_X1 U9335 ( .A1(n9202), .A2(n9203), .ZN(n9400) );
  OR2_X1 U9336 ( .A1(n8538), .A2(n8962), .ZN(n9203) );
  OR2_X1 U9337 ( .A1(n9401), .A2(n9402), .ZN(n9202) );
  AND2_X1 U9338 ( .A1(n9199), .A2(n9198), .ZN(n9402) );
  AND2_X1 U9339 ( .A1(n9196), .A2(n9403), .ZN(n9401) );
  OR2_X1 U9340 ( .A1(n9198), .A2(n9199), .ZN(n9403) );
  OR2_X1 U9341 ( .A1(n8533), .A2(n8962), .ZN(n9199) );
  OR2_X1 U9342 ( .A1(n9404), .A2(n9405), .ZN(n9198) );
  AND2_X1 U9343 ( .A1(n9193), .A2(n9195), .ZN(n9405) );
  AND2_X1 U9344 ( .A1(n9406), .A2(n9194), .ZN(n9404) );
  OR2_X1 U9345 ( .A1(n9195), .A2(n9193), .ZN(n9406) );
  XOR2_X1 U9346 ( .A(n9407), .B(n9408), .Z(n9193) );
  XOR2_X1 U9347 ( .A(n9409), .B(n9410), .Z(n9408) );
  OR2_X1 U9348 ( .A1(n9411), .A2(n9412), .ZN(n9195) );
  AND2_X1 U9349 ( .A1(n9191), .A2(n9190), .ZN(n9412) );
  AND2_X1 U9350 ( .A1(n9188), .A2(n9413), .ZN(n9411) );
  OR2_X1 U9351 ( .A1(n9190), .A2(n9191), .ZN(n9413) );
  OR2_X1 U9352 ( .A1(n8523), .A2(n8962), .ZN(n9191) );
  OR2_X1 U9353 ( .A1(n9414), .A2(n9415), .ZN(n9190) );
  AND2_X1 U9354 ( .A1(n9173), .A2(n9174), .ZN(n9415) );
  AND2_X1 U9355 ( .A1(n9416), .A2(n9417), .ZN(n9414) );
  OR2_X1 U9356 ( .A1(n9174), .A2(n9173), .ZN(n9417) );
  OR2_X1 U9357 ( .A1(n8515), .A2(n8962), .ZN(n9173) );
  OR2_X1 U9358 ( .A1(n8962), .A2(n9418), .ZN(n9174) );
  OR2_X1 U9359 ( .A1(n8956), .A2(n9185), .ZN(n9418) );
  INV_X1 U9360 ( .A(n9175), .ZN(n9416) );
  OR2_X1 U9361 ( .A1(n9419), .A2(n9420), .ZN(n9175) );
  AND2_X1 U9362 ( .A1(b_26_), .A2(n9421), .ZN(n9420) );
  OR2_X1 U9363 ( .A1(n9422), .A2(n7343), .ZN(n9421) );
  AND2_X1 U9364 ( .A1(a_30_), .A2(n9311), .ZN(n9422) );
  AND2_X1 U9365 ( .A1(b_25_), .A2(n9423), .ZN(n9419) );
  OR2_X1 U9366 ( .A1(n9424), .A2(n7347), .ZN(n9423) );
  AND2_X1 U9367 ( .A1(a_31_), .A2(n9185), .ZN(n9424) );
  XOR2_X1 U9368 ( .A(n9425), .B(n9426), .Z(n9188) );
  XNOR2_X1 U9369 ( .A(n9427), .B(n9428), .ZN(n9425) );
  XOR2_X1 U9370 ( .A(n9429), .B(n9430), .Z(n9196) );
  XOR2_X1 U9371 ( .A(n9431), .B(n9432), .Z(n9430) );
  XNOR2_X1 U9372 ( .A(n9433), .B(n9434), .ZN(n9200) );
  XNOR2_X1 U9373 ( .A(n9435), .B(n9436), .ZN(n9433) );
  XOR2_X1 U9374 ( .A(n9437), .B(n9438), .Z(n9204) );
  XOR2_X1 U9375 ( .A(n9439), .B(n9440), .Z(n9438) );
  XOR2_X1 U9376 ( .A(n9441), .B(n9442), .Z(n9208) );
  XOR2_X1 U9377 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR2_X1 U9378 ( .A(n9445), .B(n9446), .Z(n9212) );
  XOR2_X1 U9379 ( .A(n9447), .B(n9448), .Z(n9446) );
  XOR2_X1 U9380 ( .A(n9449), .B(n9450), .Z(n9216) );
  XOR2_X1 U9381 ( .A(n9451), .B(n9452), .Z(n9450) );
  XOR2_X1 U9382 ( .A(n9453), .B(n9454), .Z(n9220) );
  XOR2_X1 U9383 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR2_X1 U9384 ( .A(n9457), .B(n9458), .Z(n9224) );
  XOR2_X1 U9385 ( .A(n9459), .B(n9460), .Z(n9458) );
  XOR2_X1 U9386 ( .A(n9461), .B(n9462), .Z(n9228) );
  XOR2_X1 U9387 ( .A(n9463), .B(n9464), .Z(n9462) );
  XOR2_X1 U9388 ( .A(n9465), .B(n9466), .Z(n9232) );
  XOR2_X1 U9389 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR2_X1 U9390 ( .A(n9469), .B(n9470), .Z(n9236) );
  XOR2_X1 U9391 ( .A(n9471), .B(n9472), .Z(n9470) );
  XOR2_X1 U9392 ( .A(n9473), .B(n9474), .Z(n9240) );
  XOR2_X1 U9393 ( .A(n9475), .B(n9476), .Z(n9474) );
  XOR2_X1 U9394 ( .A(n9477), .B(n9478), .Z(n9244) );
  XOR2_X1 U9395 ( .A(n9479), .B(n9480), .Z(n9478) );
  XOR2_X1 U9396 ( .A(n9481), .B(n9482), .Z(n9248) );
  XOR2_X1 U9397 ( .A(n9483), .B(n9484), .Z(n9482) );
  XOR2_X1 U9398 ( .A(n9485), .B(n9486), .Z(n9252) );
  XOR2_X1 U9399 ( .A(n9487), .B(n9488), .Z(n9486) );
  XOR2_X1 U9400 ( .A(n9489), .B(n9490), .Z(n9256) );
  XOR2_X1 U9401 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR2_X1 U9402 ( .A(n9493), .B(n9494), .Z(n9260) );
  XOR2_X1 U9403 ( .A(n9495), .B(n9496), .Z(n9494) );
  XOR2_X1 U9404 ( .A(n9497), .B(n9498), .Z(n9264) );
  XOR2_X1 U9405 ( .A(n9499), .B(n9500), .Z(n9498) );
  XOR2_X1 U9406 ( .A(n9501), .B(n9502), .Z(n9268) );
  XOR2_X1 U9407 ( .A(n9503), .B(n9504), .Z(n9502) );
  XOR2_X1 U9408 ( .A(n9505), .B(n9506), .Z(n9272) );
  XOR2_X1 U9409 ( .A(n9507), .B(n9508), .Z(n9506) );
  OR2_X1 U9410 ( .A1(n7955), .A2(n8962), .ZN(n9278) );
  XOR2_X1 U9411 ( .A(n9509), .B(n9510), .Z(n9277) );
  XOR2_X1 U9412 ( .A(n9511), .B(n9512), .Z(n9510) );
  XNOR2_X1 U9413 ( .A(n9513), .B(n9514), .ZN(n9280) );
  XNOR2_X1 U9414 ( .A(n9515), .B(n9516), .ZN(n9513) );
  XOR2_X1 U9415 ( .A(n9517), .B(n9518), .Z(n9284) );
  XOR2_X1 U9416 ( .A(n9519), .B(n9520), .Z(n9518) );
  XOR2_X1 U9417 ( .A(n9521), .B(n9522), .Z(n9288) );
  XOR2_X1 U9418 ( .A(n9523), .B(n9524), .Z(n9522) );
  OR2_X1 U9419 ( .A1(n7730), .A2(n8962), .ZN(n9294) );
  XOR2_X1 U9420 ( .A(n9525), .B(n9526), .Z(n9293) );
  XOR2_X1 U9421 ( .A(n9527), .B(n9528), .Z(n9526) );
  XOR2_X1 U9422 ( .A(n9529), .B(n9530), .Z(n9296) );
  XOR2_X1 U9423 ( .A(n9531), .B(n9532), .Z(n9530) );
  OR2_X1 U9424 ( .A1(n9300), .A2(n9303), .ZN(n9325) );
  OR2_X1 U9425 ( .A1(n7660), .A2(n8962), .ZN(n9303) );
  XOR2_X1 U9426 ( .A(n9533), .B(n9534), .Z(n9300) );
  XOR2_X1 U9427 ( .A(n9535), .B(n9536), .Z(n9534) );
  XOR2_X1 U9428 ( .A(n9308), .B(n9537), .Z(n9083) );
  XOR2_X1 U9429 ( .A(n9307), .B(n9306), .Z(n9537) );
  OR2_X1 U9430 ( .A1(n7660), .A2(n9185), .ZN(n9306) );
  OR2_X1 U9431 ( .A1(n9538), .A2(n9539), .ZN(n9307) );
  AND2_X1 U9432 ( .A1(n9536), .A2(n9535), .ZN(n9539) );
  AND2_X1 U9433 ( .A1(n9533), .A2(n9540), .ZN(n9538) );
  OR2_X1 U9434 ( .A1(n9536), .A2(n9535), .ZN(n9540) );
  OR2_X1 U9435 ( .A1(n9541), .A2(n9542), .ZN(n9535) );
  AND2_X1 U9436 ( .A1(n9532), .A2(n9531), .ZN(n9542) );
  AND2_X1 U9437 ( .A1(n9529), .A2(n9543), .ZN(n9541) );
  OR2_X1 U9438 ( .A1(n9532), .A2(n9531), .ZN(n9543) );
  OR2_X1 U9439 ( .A1(n9544), .A2(n9545), .ZN(n9531) );
  AND2_X1 U9440 ( .A1(n9528), .A2(n9527), .ZN(n9545) );
  AND2_X1 U9441 ( .A1(n9525), .A2(n9546), .ZN(n9544) );
  OR2_X1 U9442 ( .A1(n9528), .A2(n9527), .ZN(n9546) );
  OR2_X1 U9443 ( .A1(n9547), .A2(n9548), .ZN(n9527) );
  AND2_X1 U9444 ( .A1(n9524), .A2(n9523), .ZN(n9548) );
  AND2_X1 U9445 ( .A1(n9521), .A2(n9549), .ZN(n9547) );
  OR2_X1 U9446 ( .A1(n9524), .A2(n9523), .ZN(n9549) );
  OR2_X1 U9447 ( .A1(n9550), .A2(n9551), .ZN(n9523) );
  AND2_X1 U9448 ( .A1(n9520), .A2(n9519), .ZN(n9551) );
  AND2_X1 U9449 ( .A1(n9517), .A2(n9552), .ZN(n9550) );
  OR2_X1 U9450 ( .A1(n9520), .A2(n9519), .ZN(n9552) );
  OR2_X1 U9451 ( .A1(n9553), .A2(n9554), .ZN(n9519) );
  AND2_X1 U9452 ( .A1(n9516), .A2(n9515), .ZN(n9554) );
  AND2_X1 U9453 ( .A1(n9514), .A2(n9555), .ZN(n9553) );
  OR2_X1 U9454 ( .A1(n9516), .A2(n9515), .ZN(n9555) );
  OR2_X1 U9455 ( .A1(n7955), .A2(n9185), .ZN(n9515) );
  OR2_X1 U9456 ( .A1(n9556), .A2(n9557), .ZN(n9516) );
  AND2_X1 U9457 ( .A1(n9512), .A2(n9511), .ZN(n9557) );
  AND2_X1 U9458 ( .A1(n9509), .A2(n9558), .ZN(n9556) );
  OR2_X1 U9459 ( .A1(n9512), .A2(n9511), .ZN(n9558) );
  OR2_X1 U9460 ( .A1(n9559), .A2(n9560), .ZN(n9511) );
  AND2_X1 U9461 ( .A1(n9508), .A2(n9507), .ZN(n9560) );
  AND2_X1 U9462 ( .A1(n9505), .A2(n9561), .ZN(n9559) );
  OR2_X1 U9463 ( .A1(n9508), .A2(n9507), .ZN(n9561) );
  OR2_X1 U9464 ( .A1(n9562), .A2(n9563), .ZN(n9507) );
  AND2_X1 U9465 ( .A1(n9504), .A2(n9503), .ZN(n9563) );
  AND2_X1 U9466 ( .A1(n9501), .A2(n9564), .ZN(n9562) );
  OR2_X1 U9467 ( .A1(n9504), .A2(n9503), .ZN(n9564) );
  OR2_X1 U9468 ( .A1(n9565), .A2(n9566), .ZN(n9503) );
  AND2_X1 U9469 ( .A1(n9500), .A2(n9499), .ZN(n9566) );
  AND2_X1 U9470 ( .A1(n9497), .A2(n9567), .ZN(n9565) );
  OR2_X1 U9471 ( .A1(n9500), .A2(n9499), .ZN(n9567) );
  OR2_X1 U9472 ( .A1(n9568), .A2(n9569), .ZN(n9499) );
  AND2_X1 U9473 ( .A1(n9496), .A2(n9495), .ZN(n9569) );
  AND2_X1 U9474 ( .A1(n9493), .A2(n9570), .ZN(n9568) );
  OR2_X1 U9475 ( .A1(n9496), .A2(n9495), .ZN(n9570) );
  OR2_X1 U9476 ( .A1(n9571), .A2(n9572), .ZN(n9495) );
  AND2_X1 U9477 ( .A1(n9492), .A2(n9491), .ZN(n9572) );
  AND2_X1 U9478 ( .A1(n9489), .A2(n9573), .ZN(n9571) );
  OR2_X1 U9479 ( .A1(n9492), .A2(n9491), .ZN(n9573) );
  OR2_X1 U9480 ( .A1(n9574), .A2(n9575), .ZN(n9491) );
  AND2_X1 U9481 ( .A1(n9488), .A2(n9487), .ZN(n9575) );
  AND2_X1 U9482 ( .A1(n9485), .A2(n9576), .ZN(n9574) );
  OR2_X1 U9483 ( .A1(n9488), .A2(n9487), .ZN(n9576) );
  OR2_X1 U9484 ( .A1(n9577), .A2(n9578), .ZN(n9487) );
  AND2_X1 U9485 ( .A1(n9484), .A2(n9483), .ZN(n9578) );
  AND2_X1 U9486 ( .A1(n9481), .A2(n9579), .ZN(n9577) );
  OR2_X1 U9487 ( .A1(n9484), .A2(n9483), .ZN(n9579) );
  OR2_X1 U9488 ( .A1(n9580), .A2(n9581), .ZN(n9483) );
  AND2_X1 U9489 ( .A1(n9480), .A2(n9479), .ZN(n9581) );
  AND2_X1 U9490 ( .A1(n9477), .A2(n9582), .ZN(n9580) );
  OR2_X1 U9491 ( .A1(n9480), .A2(n9479), .ZN(n9582) );
  OR2_X1 U9492 ( .A1(n9583), .A2(n9584), .ZN(n9479) );
  AND2_X1 U9493 ( .A1(n9476), .A2(n9475), .ZN(n9584) );
  AND2_X1 U9494 ( .A1(n9473), .A2(n9585), .ZN(n9583) );
  OR2_X1 U9495 ( .A1(n9476), .A2(n9475), .ZN(n9585) );
  OR2_X1 U9496 ( .A1(n9586), .A2(n9587), .ZN(n9475) );
  AND2_X1 U9497 ( .A1(n9472), .A2(n9471), .ZN(n9587) );
  AND2_X1 U9498 ( .A1(n9469), .A2(n9588), .ZN(n9586) );
  OR2_X1 U9499 ( .A1(n9472), .A2(n9471), .ZN(n9588) );
  OR2_X1 U9500 ( .A1(n9589), .A2(n9590), .ZN(n9471) );
  AND2_X1 U9501 ( .A1(n9468), .A2(n9467), .ZN(n9590) );
  AND2_X1 U9502 ( .A1(n9465), .A2(n9591), .ZN(n9589) );
  OR2_X1 U9503 ( .A1(n9468), .A2(n9467), .ZN(n9591) );
  OR2_X1 U9504 ( .A1(n9592), .A2(n9593), .ZN(n9467) );
  AND2_X1 U9505 ( .A1(n9464), .A2(n9463), .ZN(n9593) );
  AND2_X1 U9506 ( .A1(n9461), .A2(n9594), .ZN(n9592) );
  OR2_X1 U9507 ( .A1(n9464), .A2(n9463), .ZN(n9594) );
  OR2_X1 U9508 ( .A1(n9595), .A2(n9596), .ZN(n9463) );
  AND2_X1 U9509 ( .A1(n9460), .A2(n9459), .ZN(n9596) );
  AND2_X1 U9510 ( .A1(n9457), .A2(n9597), .ZN(n9595) );
  OR2_X1 U9511 ( .A1(n9460), .A2(n9459), .ZN(n9597) );
  OR2_X1 U9512 ( .A1(n9598), .A2(n9599), .ZN(n9459) );
  AND2_X1 U9513 ( .A1(n9456), .A2(n9455), .ZN(n9599) );
  AND2_X1 U9514 ( .A1(n9453), .A2(n9600), .ZN(n9598) );
  OR2_X1 U9515 ( .A1(n9456), .A2(n9455), .ZN(n9600) );
  OR2_X1 U9516 ( .A1(n9601), .A2(n9602), .ZN(n9455) );
  AND2_X1 U9517 ( .A1(n9452), .A2(n9451), .ZN(n9602) );
  AND2_X1 U9518 ( .A1(n9449), .A2(n9603), .ZN(n9601) );
  OR2_X1 U9519 ( .A1(n9452), .A2(n9451), .ZN(n9603) );
  OR2_X1 U9520 ( .A1(n9604), .A2(n9605), .ZN(n9451) );
  AND2_X1 U9521 ( .A1(n9448), .A2(n9447), .ZN(n9605) );
  AND2_X1 U9522 ( .A1(n9445), .A2(n9606), .ZN(n9604) );
  OR2_X1 U9523 ( .A1(n9448), .A2(n9447), .ZN(n9606) );
  OR2_X1 U9524 ( .A1(n9607), .A2(n9608), .ZN(n9447) );
  AND2_X1 U9525 ( .A1(n9444), .A2(n9443), .ZN(n9608) );
  AND2_X1 U9526 ( .A1(n9441), .A2(n9609), .ZN(n9607) );
  OR2_X1 U9527 ( .A1(n9444), .A2(n9443), .ZN(n9609) );
  OR2_X1 U9528 ( .A1(n9610), .A2(n9611), .ZN(n9443) );
  AND2_X1 U9529 ( .A1(n9440), .A2(n9439), .ZN(n9611) );
  AND2_X1 U9530 ( .A1(n9437), .A2(n9612), .ZN(n9610) );
  OR2_X1 U9531 ( .A1(n9440), .A2(n9439), .ZN(n9612) );
  OR2_X1 U9532 ( .A1(n9613), .A2(n9614), .ZN(n9439) );
  AND2_X1 U9533 ( .A1(n9434), .A2(n9436), .ZN(n9614) );
  AND2_X1 U9534 ( .A1(n9615), .A2(n9435), .ZN(n9613) );
  OR2_X1 U9535 ( .A1(n9434), .A2(n9436), .ZN(n9615) );
  OR2_X1 U9536 ( .A1(n9616), .A2(n9617), .ZN(n9436) );
  AND2_X1 U9537 ( .A1(n9432), .A2(n9431), .ZN(n9617) );
  AND2_X1 U9538 ( .A1(n9429), .A2(n9618), .ZN(n9616) );
  OR2_X1 U9539 ( .A1(n9432), .A2(n9431), .ZN(n9618) );
  OR2_X1 U9540 ( .A1(n9619), .A2(n9620), .ZN(n9431) );
  AND2_X1 U9541 ( .A1(n9410), .A2(n9409), .ZN(n9620) );
  AND2_X1 U9542 ( .A1(n9407), .A2(n9621), .ZN(n9619) );
  OR2_X1 U9543 ( .A1(n9410), .A2(n9409), .ZN(n9621) );
  OR2_X1 U9544 ( .A1(n9622), .A2(n9623), .ZN(n9409) );
  AND2_X1 U9545 ( .A1(n9426), .A2(n9427), .ZN(n9623) );
  AND2_X1 U9546 ( .A1(n9624), .A2(n9625), .ZN(n9622) );
  OR2_X1 U9547 ( .A1(n9426), .A2(n9427), .ZN(n9625) );
  OR2_X1 U9548 ( .A1(n9185), .A2(n9626), .ZN(n9427) );
  OR2_X1 U9549 ( .A1(n8515), .A2(n9185), .ZN(n9426) );
  INV_X1 U9550 ( .A(n9428), .ZN(n9624) );
  OR2_X1 U9551 ( .A1(n9627), .A2(n9628), .ZN(n9428) );
  AND2_X1 U9552 ( .A1(b_25_), .A2(n9629), .ZN(n9628) );
  OR2_X1 U9553 ( .A1(n9630), .A2(n7343), .ZN(n9629) );
  AND2_X1 U9554 ( .A1(a_30_), .A2(n9631), .ZN(n9630) );
  AND2_X1 U9555 ( .A1(b_24_), .A2(n9632), .ZN(n9627) );
  OR2_X1 U9556 ( .A1(n9633), .A2(n7347), .ZN(n9632) );
  AND2_X1 U9557 ( .A1(a_31_), .A2(n9311), .ZN(n9633) );
  OR2_X1 U9558 ( .A1(n8523), .A2(n9185), .ZN(n9410) );
  XOR2_X1 U9559 ( .A(n9634), .B(n9635), .Z(n9407) );
  XNOR2_X1 U9560 ( .A(n9636), .B(n9637), .ZN(n9634) );
  OR2_X1 U9561 ( .A1(n8528), .A2(n9185), .ZN(n9432) );
  XOR2_X1 U9562 ( .A(n9638), .B(n9639), .Z(n9429) );
  XOR2_X1 U9563 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR2_X1 U9564 ( .A(n9642), .B(n9643), .Z(n9434) );
  XOR2_X1 U9565 ( .A(n9644), .B(n9645), .Z(n9643) );
  OR2_X1 U9566 ( .A1(n8538), .A2(n9185), .ZN(n9440) );
  XOR2_X1 U9567 ( .A(n9646), .B(n9647), .Z(n9437) );
  XOR2_X1 U9568 ( .A(n9648), .B(n9649), .Z(n9647) );
  OR2_X1 U9569 ( .A1(n8543), .A2(n9185), .ZN(n9444) );
  XNOR2_X1 U9570 ( .A(n9650), .B(n9651), .ZN(n9441) );
  XNOR2_X1 U9571 ( .A(n9652), .B(n9653), .ZN(n9650) );
  OR2_X1 U9572 ( .A1(n8548), .A2(n9185), .ZN(n9448) );
  XOR2_X1 U9573 ( .A(n9654), .B(n9655), .Z(n9445) );
  XOR2_X1 U9574 ( .A(n9656), .B(n9657), .Z(n9655) );
  OR2_X1 U9575 ( .A1(n8553), .A2(n9185), .ZN(n9452) );
  XOR2_X1 U9576 ( .A(n9658), .B(n9659), .Z(n9449) );
  XOR2_X1 U9577 ( .A(n9660), .B(n9661), .Z(n9659) );
  OR2_X1 U9578 ( .A1(n8558), .A2(n9185), .ZN(n9456) );
  XOR2_X1 U9579 ( .A(n9662), .B(n9663), .Z(n9453) );
  XOR2_X1 U9580 ( .A(n9664), .B(n9665), .Z(n9663) );
  OR2_X1 U9581 ( .A1(n8563), .A2(n9185), .ZN(n9460) );
  XOR2_X1 U9582 ( .A(n9666), .B(n9667), .Z(n9457) );
  XOR2_X1 U9583 ( .A(n9668), .B(n9669), .Z(n9667) );
  OR2_X1 U9584 ( .A1(n8568), .A2(n9185), .ZN(n9464) );
  XOR2_X1 U9585 ( .A(n9670), .B(n9671), .Z(n9461) );
  XOR2_X1 U9586 ( .A(n9672), .B(n9673), .Z(n9671) );
  OR2_X1 U9587 ( .A1(n8573), .A2(n9185), .ZN(n9468) );
  XOR2_X1 U9588 ( .A(n9674), .B(n9675), .Z(n9465) );
  XOR2_X1 U9589 ( .A(n9676), .B(n9677), .Z(n9675) );
  OR2_X1 U9590 ( .A1(n8578), .A2(n9185), .ZN(n9472) );
  XOR2_X1 U9591 ( .A(n9678), .B(n9679), .Z(n9469) );
  XOR2_X1 U9592 ( .A(n9680), .B(n9681), .Z(n9679) );
  OR2_X1 U9593 ( .A1(n8583), .A2(n9185), .ZN(n9476) );
  XOR2_X1 U9594 ( .A(n9682), .B(n9683), .Z(n9473) );
  XOR2_X1 U9595 ( .A(n9684), .B(n9685), .Z(n9683) );
  OR2_X1 U9596 ( .A1(n8588), .A2(n9185), .ZN(n9480) );
  XOR2_X1 U9597 ( .A(n9686), .B(n9687), .Z(n9477) );
  XOR2_X1 U9598 ( .A(n9688), .B(n9689), .Z(n9687) );
  OR2_X1 U9599 ( .A1(n8593), .A2(n9185), .ZN(n9484) );
  XOR2_X1 U9600 ( .A(n9690), .B(n9691), .Z(n9481) );
  XOR2_X1 U9601 ( .A(n9692), .B(n9693), .Z(n9691) );
  OR2_X1 U9602 ( .A1(n8598), .A2(n9185), .ZN(n9488) );
  XOR2_X1 U9603 ( .A(n9694), .B(n9695), .Z(n9485) );
  XOR2_X1 U9604 ( .A(n9696), .B(n9697), .Z(n9695) );
  OR2_X1 U9605 ( .A1(n8603), .A2(n9185), .ZN(n9492) );
  XOR2_X1 U9606 ( .A(n9698), .B(n9699), .Z(n9489) );
  XOR2_X1 U9607 ( .A(n9700), .B(n9701), .Z(n9699) );
  OR2_X1 U9608 ( .A1(n8608), .A2(n9185), .ZN(n9496) );
  XOR2_X1 U9609 ( .A(n9702), .B(n9703), .Z(n9493) );
  XOR2_X1 U9610 ( .A(n9704), .B(n9705), .Z(n9703) );
  OR2_X1 U9611 ( .A1(n8287), .A2(n9185), .ZN(n9500) );
  XOR2_X1 U9612 ( .A(n9706), .B(n9707), .Z(n9497) );
  XOR2_X1 U9613 ( .A(n9708), .B(n9709), .Z(n9707) );
  OR2_X1 U9614 ( .A1(n8191), .A2(n9185), .ZN(n9504) );
  XNOR2_X1 U9615 ( .A(n9710), .B(n9711), .ZN(n9501) );
  XNOR2_X1 U9616 ( .A(n9712), .B(n9713), .ZN(n9710) );
  OR2_X1 U9617 ( .A1(n8107), .A2(n9185), .ZN(n9508) );
  XOR2_X1 U9618 ( .A(n9714), .B(n9715), .Z(n9505) );
  XOR2_X1 U9619 ( .A(n9716), .B(n9717), .Z(n9715) );
  OR2_X1 U9620 ( .A1(n8025), .A2(n9185), .ZN(n9512) );
  XOR2_X1 U9621 ( .A(n9718), .B(n9719), .Z(n9509) );
  XOR2_X1 U9622 ( .A(n9720), .B(n9721), .Z(n9719) );
  XOR2_X1 U9623 ( .A(n9722), .B(n9723), .Z(n9514) );
  XOR2_X1 U9624 ( .A(n9724), .B(n9725), .Z(n9723) );
  OR2_X1 U9625 ( .A1(n7887), .A2(n9185), .ZN(n9520) );
  XNOR2_X1 U9626 ( .A(n9726), .B(n9727), .ZN(n9517) );
  XNOR2_X1 U9627 ( .A(n9728), .B(n9729), .ZN(n9726) );
  OR2_X1 U9628 ( .A1(n7828), .A2(n9185), .ZN(n9524) );
  XOR2_X1 U9629 ( .A(n9730), .B(n9731), .Z(n9521) );
  XOR2_X1 U9630 ( .A(n9732), .B(n9733), .Z(n9731) );
  OR2_X1 U9631 ( .A1(n7820), .A2(n9185), .ZN(n9528) );
  XOR2_X1 U9632 ( .A(n9734), .B(n9735), .Z(n9525) );
  XOR2_X1 U9633 ( .A(n9736), .B(n9737), .Z(n9735) );
  OR2_X1 U9634 ( .A1(n7730), .A2(n9185), .ZN(n9532) );
  XOR2_X1 U9635 ( .A(n9738), .B(n9739), .Z(n9529) );
  XOR2_X1 U9636 ( .A(n9740), .B(n9741), .Z(n9739) );
  OR2_X1 U9637 ( .A1(n7697), .A2(n9185), .ZN(n9536) );
  XOR2_X1 U9638 ( .A(n9742), .B(n9743), .Z(n9533) );
  XOR2_X1 U9639 ( .A(n9744), .B(n9745), .Z(n9743) );
  XOR2_X1 U9640 ( .A(n9316), .B(n9746), .Z(n9308) );
  XOR2_X1 U9641 ( .A(n9315), .B(n9314), .Z(n9746) );
  OR2_X1 U9642 ( .A1(n7697), .A2(n9311), .ZN(n9314) );
  OR2_X1 U9643 ( .A1(n9747), .A2(n9748), .ZN(n9315) );
  AND2_X1 U9644 ( .A1(n9745), .A2(n9744), .ZN(n9748) );
  AND2_X1 U9645 ( .A1(n9742), .A2(n9749), .ZN(n9747) );
  OR2_X1 U9646 ( .A1(n9745), .A2(n9744), .ZN(n9749) );
  OR2_X1 U9647 ( .A1(n9750), .A2(n9751), .ZN(n9744) );
  AND2_X1 U9648 ( .A1(n9741), .A2(n9740), .ZN(n9751) );
  AND2_X1 U9649 ( .A1(n9738), .A2(n9752), .ZN(n9750) );
  OR2_X1 U9650 ( .A1(n9741), .A2(n9740), .ZN(n9752) );
  OR2_X1 U9651 ( .A1(n9753), .A2(n9754), .ZN(n9740) );
  AND2_X1 U9652 ( .A1(n9737), .A2(n9736), .ZN(n9754) );
  AND2_X1 U9653 ( .A1(n9734), .A2(n9755), .ZN(n9753) );
  OR2_X1 U9654 ( .A1(n9737), .A2(n9736), .ZN(n9755) );
  OR2_X1 U9655 ( .A1(n9756), .A2(n9757), .ZN(n9736) );
  AND2_X1 U9656 ( .A1(n9733), .A2(n9732), .ZN(n9757) );
  AND2_X1 U9657 ( .A1(n9730), .A2(n9758), .ZN(n9756) );
  OR2_X1 U9658 ( .A1(n9733), .A2(n9732), .ZN(n9758) );
  OR2_X1 U9659 ( .A1(n9759), .A2(n9760), .ZN(n9732) );
  AND2_X1 U9660 ( .A1(n9729), .A2(n9728), .ZN(n9760) );
  AND2_X1 U9661 ( .A1(n9727), .A2(n9761), .ZN(n9759) );
  OR2_X1 U9662 ( .A1(n9729), .A2(n9728), .ZN(n9761) );
  OR2_X1 U9663 ( .A1(n7955), .A2(n9311), .ZN(n9728) );
  OR2_X1 U9664 ( .A1(n9762), .A2(n9763), .ZN(n9729) );
  AND2_X1 U9665 ( .A1(n9725), .A2(n9724), .ZN(n9763) );
  AND2_X1 U9666 ( .A1(n9722), .A2(n9764), .ZN(n9762) );
  OR2_X1 U9667 ( .A1(n9725), .A2(n9724), .ZN(n9764) );
  OR2_X1 U9668 ( .A1(n9765), .A2(n9766), .ZN(n9724) );
  AND2_X1 U9669 ( .A1(n9721), .A2(n9720), .ZN(n9766) );
  AND2_X1 U9670 ( .A1(n9718), .A2(n9767), .ZN(n9765) );
  OR2_X1 U9671 ( .A1(n9721), .A2(n9720), .ZN(n9767) );
  OR2_X1 U9672 ( .A1(n9768), .A2(n9769), .ZN(n9720) );
  AND2_X1 U9673 ( .A1(n9717), .A2(n9716), .ZN(n9769) );
  AND2_X1 U9674 ( .A1(n9714), .A2(n9770), .ZN(n9768) );
  OR2_X1 U9675 ( .A1(n9717), .A2(n9716), .ZN(n9770) );
  OR2_X1 U9676 ( .A1(n9771), .A2(n9772), .ZN(n9716) );
  AND2_X1 U9677 ( .A1(n9713), .A2(n9712), .ZN(n9772) );
  AND2_X1 U9678 ( .A1(n9711), .A2(n9773), .ZN(n9771) );
  OR2_X1 U9679 ( .A1(n9713), .A2(n9712), .ZN(n9773) );
  OR2_X1 U9680 ( .A1(n8287), .A2(n9311), .ZN(n9712) );
  OR2_X1 U9681 ( .A1(n9774), .A2(n9775), .ZN(n9713) );
  AND2_X1 U9682 ( .A1(n9709), .A2(n9708), .ZN(n9775) );
  AND2_X1 U9683 ( .A1(n9706), .A2(n9776), .ZN(n9774) );
  OR2_X1 U9684 ( .A1(n9709), .A2(n9708), .ZN(n9776) );
  OR2_X1 U9685 ( .A1(n9777), .A2(n9778), .ZN(n9708) );
  AND2_X1 U9686 ( .A1(n9705), .A2(n9704), .ZN(n9778) );
  AND2_X1 U9687 ( .A1(n9702), .A2(n9779), .ZN(n9777) );
  OR2_X1 U9688 ( .A1(n9705), .A2(n9704), .ZN(n9779) );
  OR2_X1 U9689 ( .A1(n9780), .A2(n9781), .ZN(n9704) );
  AND2_X1 U9690 ( .A1(n9701), .A2(n9700), .ZN(n9781) );
  AND2_X1 U9691 ( .A1(n9698), .A2(n9782), .ZN(n9780) );
  OR2_X1 U9692 ( .A1(n9701), .A2(n9700), .ZN(n9782) );
  OR2_X1 U9693 ( .A1(n9783), .A2(n9784), .ZN(n9700) );
  AND2_X1 U9694 ( .A1(n9697), .A2(n9696), .ZN(n9784) );
  AND2_X1 U9695 ( .A1(n9694), .A2(n9785), .ZN(n9783) );
  OR2_X1 U9696 ( .A1(n9697), .A2(n9696), .ZN(n9785) );
  OR2_X1 U9697 ( .A1(n9786), .A2(n9787), .ZN(n9696) );
  AND2_X1 U9698 ( .A1(n9693), .A2(n9692), .ZN(n9787) );
  AND2_X1 U9699 ( .A1(n9690), .A2(n9788), .ZN(n9786) );
  OR2_X1 U9700 ( .A1(n9693), .A2(n9692), .ZN(n9788) );
  OR2_X1 U9701 ( .A1(n9789), .A2(n9790), .ZN(n9692) );
  AND2_X1 U9702 ( .A1(n9689), .A2(n9688), .ZN(n9790) );
  AND2_X1 U9703 ( .A1(n9686), .A2(n9791), .ZN(n9789) );
  OR2_X1 U9704 ( .A1(n9689), .A2(n9688), .ZN(n9791) );
  OR2_X1 U9705 ( .A1(n9792), .A2(n9793), .ZN(n9688) );
  AND2_X1 U9706 ( .A1(n9685), .A2(n9684), .ZN(n9793) );
  AND2_X1 U9707 ( .A1(n9682), .A2(n9794), .ZN(n9792) );
  OR2_X1 U9708 ( .A1(n9685), .A2(n9684), .ZN(n9794) );
  OR2_X1 U9709 ( .A1(n9795), .A2(n9796), .ZN(n9684) );
  AND2_X1 U9710 ( .A1(n9681), .A2(n9680), .ZN(n9796) );
  AND2_X1 U9711 ( .A1(n9678), .A2(n9797), .ZN(n9795) );
  OR2_X1 U9712 ( .A1(n9681), .A2(n9680), .ZN(n9797) );
  OR2_X1 U9713 ( .A1(n9798), .A2(n9799), .ZN(n9680) );
  AND2_X1 U9714 ( .A1(n9677), .A2(n9676), .ZN(n9799) );
  AND2_X1 U9715 ( .A1(n9674), .A2(n9800), .ZN(n9798) );
  OR2_X1 U9716 ( .A1(n9677), .A2(n9676), .ZN(n9800) );
  OR2_X1 U9717 ( .A1(n9801), .A2(n9802), .ZN(n9676) );
  AND2_X1 U9718 ( .A1(n9673), .A2(n9672), .ZN(n9802) );
  AND2_X1 U9719 ( .A1(n9670), .A2(n9803), .ZN(n9801) );
  OR2_X1 U9720 ( .A1(n9673), .A2(n9672), .ZN(n9803) );
  OR2_X1 U9721 ( .A1(n9804), .A2(n9805), .ZN(n9672) );
  AND2_X1 U9722 ( .A1(n9669), .A2(n9668), .ZN(n9805) );
  AND2_X1 U9723 ( .A1(n9666), .A2(n9806), .ZN(n9804) );
  OR2_X1 U9724 ( .A1(n9669), .A2(n9668), .ZN(n9806) );
  OR2_X1 U9725 ( .A1(n9807), .A2(n9808), .ZN(n9668) );
  AND2_X1 U9726 ( .A1(n9665), .A2(n9664), .ZN(n9808) );
  AND2_X1 U9727 ( .A1(n9662), .A2(n9809), .ZN(n9807) );
  OR2_X1 U9728 ( .A1(n9665), .A2(n9664), .ZN(n9809) );
  OR2_X1 U9729 ( .A1(n9810), .A2(n9811), .ZN(n9664) );
  AND2_X1 U9730 ( .A1(n9661), .A2(n9660), .ZN(n9811) );
  AND2_X1 U9731 ( .A1(n9658), .A2(n9812), .ZN(n9810) );
  OR2_X1 U9732 ( .A1(n9661), .A2(n9660), .ZN(n9812) );
  OR2_X1 U9733 ( .A1(n9813), .A2(n9814), .ZN(n9660) );
  AND2_X1 U9734 ( .A1(n9657), .A2(n9656), .ZN(n9814) );
  AND2_X1 U9735 ( .A1(n9654), .A2(n9815), .ZN(n9813) );
  OR2_X1 U9736 ( .A1(n9657), .A2(n9656), .ZN(n9815) );
  OR2_X1 U9737 ( .A1(n9816), .A2(n9817), .ZN(n9656) );
  AND2_X1 U9738 ( .A1(n9651), .A2(n9653), .ZN(n9817) );
  AND2_X1 U9739 ( .A1(n9818), .A2(n9652), .ZN(n9816) );
  OR2_X1 U9740 ( .A1(n9651), .A2(n9653), .ZN(n9818) );
  OR2_X1 U9741 ( .A1(n9819), .A2(n9820), .ZN(n9653) );
  AND2_X1 U9742 ( .A1(n9649), .A2(n9648), .ZN(n9820) );
  AND2_X1 U9743 ( .A1(n9646), .A2(n9821), .ZN(n9819) );
  OR2_X1 U9744 ( .A1(n9649), .A2(n9648), .ZN(n9821) );
  OR2_X1 U9745 ( .A1(n9822), .A2(n9823), .ZN(n9648) );
  AND2_X1 U9746 ( .A1(n9645), .A2(n9644), .ZN(n9823) );
  AND2_X1 U9747 ( .A1(n9642), .A2(n9824), .ZN(n9822) );
  OR2_X1 U9748 ( .A1(n9645), .A2(n9644), .ZN(n9824) );
  OR2_X1 U9749 ( .A1(n9825), .A2(n9826), .ZN(n9644) );
  AND2_X1 U9750 ( .A1(n9641), .A2(n9640), .ZN(n9826) );
  AND2_X1 U9751 ( .A1(n9638), .A2(n9827), .ZN(n9825) );
  OR2_X1 U9752 ( .A1(n9641), .A2(n9640), .ZN(n9827) );
  OR2_X1 U9753 ( .A1(n9828), .A2(n9829), .ZN(n9640) );
  AND2_X1 U9754 ( .A1(n9635), .A2(n9636), .ZN(n9829) );
  AND2_X1 U9755 ( .A1(n9830), .A2(n9831), .ZN(n9828) );
  OR2_X1 U9756 ( .A1(n9635), .A2(n9636), .ZN(n9831) );
  OR2_X1 U9757 ( .A1(n9631), .A2(n9626), .ZN(n9636) );
  OR2_X1 U9758 ( .A1(n8956), .A2(n9311), .ZN(n9626) );
  OR2_X1 U9759 ( .A1(n8515), .A2(n9311), .ZN(n9635) );
  INV_X1 U9760 ( .A(n9637), .ZN(n9830) );
  OR2_X1 U9761 ( .A1(n9832), .A2(n9833), .ZN(n9637) );
  AND2_X1 U9762 ( .A1(b_24_), .A2(n9834), .ZN(n9833) );
  OR2_X1 U9763 ( .A1(n9835), .A2(n7343), .ZN(n9834) );
  AND2_X1 U9764 ( .A1(a_30_), .A2(n9836), .ZN(n9835) );
  AND2_X1 U9765 ( .A1(b_23_), .A2(n9837), .ZN(n9832) );
  OR2_X1 U9766 ( .A1(n9838), .A2(n7347), .ZN(n9837) );
  AND2_X1 U9767 ( .A1(a_31_), .A2(n9631), .ZN(n9838) );
  OR2_X1 U9768 ( .A1(n8523), .A2(n9311), .ZN(n9641) );
  XOR2_X1 U9769 ( .A(n9839), .B(n9840), .Z(n9638) );
  XNOR2_X1 U9770 ( .A(n9841), .B(n9842), .ZN(n9839) );
  OR2_X1 U9771 ( .A1(n8528), .A2(n9311), .ZN(n9645) );
  XOR2_X1 U9772 ( .A(n9843), .B(n9844), .Z(n9642) );
  XOR2_X1 U9773 ( .A(n9845), .B(n9846), .Z(n9844) );
  OR2_X1 U9774 ( .A1(n8533), .A2(n9311), .ZN(n9649) );
  XOR2_X1 U9775 ( .A(n9847), .B(n9848), .Z(n9646) );
  XOR2_X1 U9776 ( .A(n9849), .B(n9850), .Z(n9848) );
  XOR2_X1 U9777 ( .A(n9851), .B(n9852), .Z(n9651) );
  XOR2_X1 U9778 ( .A(n9853), .B(n9854), .Z(n9852) );
  OR2_X1 U9779 ( .A1(n8543), .A2(n9311), .ZN(n9657) );
  XOR2_X1 U9780 ( .A(n9855), .B(n9856), .Z(n9654) );
  XOR2_X1 U9781 ( .A(n9857), .B(n9858), .Z(n9856) );
  OR2_X1 U9782 ( .A1(n8548), .A2(n9311), .ZN(n9661) );
  XNOR2_X1 U9783 ( .A(n9859), .B(n9860), .ZN(n9658) );
  XNOR2_X1 U9784 ( .A(n9861), .B(n9862), .ZN(n9859) );
  OR2_X1 U9785 ( .A1(n8553), .A2(n9311), .ZN(n9665) );
  XOR2_X1 U9786 ( .A(n9863), .B(n9864), .Z(n9662) );
  XOR2_X1 U9787 ( .A(n9865), .B(n9866), .Z(n9864) );
  OR2_X1 U9788 ( .A1(n8558), .A2(n9311), .ZN(n9669) );
  XOR2_X1 U9789 ( .A(n9867), .B(n9868), .Z(n9666) );
  XOR2_X1 U9790 ( .A(n9869), .B(n9870), .Z(n9868) );
  OR2_X1 U9791 ( .A1(n8563), .A2(n9311), .ZN(n9673) );
  XOR2_X1 U9792 ( .A(n9871), .B(n9872), .Z(n9670) );
  XOR2_X1 U9793 ( .A(n9873), .B(n9874), .Z(n9872) );
  OR2_X1 U9794 ( .A1(n8568), .A2(n9311), .ZN(n9677) );
  XOR2_X1 U9795 ( .A(n9875), .B(n9876), .Z(n9674) );
  XOR2_X1 U9796 ( .A(n9877), .B(n9878), .Z(n9876) );
  OR2_X1 U9797 ( .A1(n8573), .A2(n9311), .ZN(n9681) );
  XOR2_X1 U9798 ( .A(n9879), .B(n9880), .Z(n9678) );
  XOR2_X1 U9799 ( .A(n9881), .B(n9882), .Z(n9880) );
  OR2_X1 U9800 ( .A1(n8578), .A2(n9311), .ZN(n9685) );
  XOR2_X1 U9801 ( .A(n9883), .B(n9884), .Z(n9682) );
  XOR2_X1 U9802 ( .A(n9885), .B(n9886), .Z(n9884) );
  OR2_X1 U9803 ( .A1(n8583), .A2(n9311), .ZN(n9689) );
  XOR2_X1 U9804 ( .A(n9887), .B(n9888), .Z(n9686) );
  XOR2_X1 U9805 ( .A(n9889), .B(n9890), .Z(n9888) );
  OR2_X1 U9806 ( .A1(n8588), .A2(n9311), .ZN(n9693) );
  XOR2_X1 U9807 ( .A(n9891), .B(n9892), .Z(n9690) );
  XOR2_X1 U9808 ( .A(n9893), .B(n9894), .Z(n9892) );
  OR2_X1 U9809 ( .A1(n8593), .A2(n9311), .ZN(n9697) );
  XOR2_X1 U9810 ( .A(n9895), .B(n9896), .Z(n9694) );
  XOR2_X1 U9811 ( .A(n9897), .B(n9898), .Z(n9896) );
  OR2_X1 U9812 ( .A1(n8598), .A2(n9311), .ZN(n9701) );
  XOR2_X1 U9813 ( .A(n9899), .B(n9900), .Z(n9698) );
  XOR2_X1 U9814 ( .A(n9901), .B(n9902), .Z(n9900) );
  OR2_X1 U9815 ( .A1(n8603), .A2(n9311), .ZN(n9705) );
  XOR2_X1 U9816 ( .A(n9903), .B(n9904), .Z(n9702) );
  XOR2_X1 U9817 ( .A(n9905), .B(n9906), .Z(n9904) );
  OR2_X1 U9818 ( .A1(n8608), .A2(n9311), .ZN(n9709) );
  XOR2_X1 U9819 ( .A(n9907), .B(n9908), .Z(n9706) );
  XOR2_X1 U9820 ( .A(n9909), .B(n9910), .Z(n9908) );
  XOR2_X1 U9821 ( .A(n9911), .B(n9912), .Z(n9711) );
  XOR2_X1 U9822 ( .A(n9913), .B(n9914), .Z(n9912) );
  OR2_X1 U9823 ( .A1(n8191), .A2(n9311), .ZN(n9717) );
  XNOR2_X1 U9824 ( .A(n9915), .B(n9916), .ZN(n9714) );
  XNOR2_X1 U9825 ( .A(n9917), .B(n9918), .ZN(n9915) );
  OR2_X1 U9826 ( .A1(n8107), .A2(n9311), .ZN(n9721) );
  XOR2_X1 U9827 ( .A(n9919), .B(n9920), .Z(n9718) );
  XOR2_X1 U9828 ( .A(n9921), .B(n9922), .Z(n9920) );
  OR2_X1 U9829 ( .A1(n8025), .A2(n9311), .ZN(n9725) );
  XOR2_X1 U9830 ( .A(n9923), .B(n9924), .Z(n9722) );
  XOR2_X1 U9831 ( .A(n9925), .B(n9926), .Z(n9924) );
  XOR2_X1 U9832 ( .A(n9927), .B(n9928), .Z(n9727) );
  XOR2_X1 U9833 ( .A(n9929), .B(n9930), .Z(n9928) );
  OR2_X1 U9834 ( .A1(n7887), .A2(n9311), .ZN(n9733) );
  XNOR2_X1 U9835 ( .A(n9931), .B(n9932), .ZN(n9730) );
  XNOR2_X1 U9836 ( .A(n9933), .B(n9934), .ZN(n9931) );
  OR2_X1 U9837 ( .A1(n7828), .A2(n9311), .ZN(n9737) );
  XOR2_X1 U9838 ( .A(n9935), .B(n9936), .Z(n9734) );
  XOR2_X1 U9839 ( .A(n9937), .B(n9938), .Z(n9936) );
  OR2_X1 U9840 ( .A1(n7820), .A2(n9311), .ZN(n9741) );
  XOR2_X1 U9841 ( .A(n9939), .B(n9940), .Z(n9738) );
  XOR2_X1 U9842 ( .A(n9941), .B(n9942), .Z(n9940) );
  OR2_X1 U9843 ( .A1(n7730), .A2(n9311), .ZN(n9745) );
  XNOR2_X1 U9844 ( .A(n9943), .B(n9944), .ZN(n9742) );
  XNOR2_X1 U9845 ( .A(n9945), .B(n9946), .ZN(n9943) );
  XOR2_X1 U9846 ( .A(n9947), .B(n9948), .Z(n9316) );
  XOR2_X1 U9847 ( .A(n9949), .B(n9950), .Z(n9948) );
  OR2_X1 U9848 ( .A1(n8350), .A2(n8349), .ZN(n7523) );
  INV_X1 U9849 ( .A(n9951), .ZN(n8349) );
  OR2_X1 U9850 ( .A1(n9952), .A2(n9953), .ZN(n9951) );
  AND2_X1 U9851 ( .A1(n9954), .A2(n9955), .ZN(n9952) );
  AND2_X1 U9852 ( .A1(n8354), .A2(n9956), .ZN(n8350) );
  INV_X1 U9853 ( .A(n8355), .ZN(n9956) );
  OR2_X1 U9854 ( .A1(n9957), .A2(n9958), .ZN(n8355) );
  AND2_X1 U9855 ( .A1(n8374), .A2(n8373), .ZN(n9958) );
  AND2_X1 U9856 ( .A1(n8371), .A2(n9959), .ZN(n9957) );
  OR2_X1 U9857 ( .A1(n8373), .A2(n8374), .ZN(n9959) );
  OR2_X1 U9858 ( .A1(n7660), .A2(n9631), .ZN(n8374) );
  OR2_X1 U9859 ( .A1(n9960), .A2(n9961), .ZN(n8373) );
  AND2_X1 U9860 ( .A1(n9321), .A2(n9320), .ZN(n9961) );
  AND2_X1 U9861 ( .A1(n9319), .A2(n9962), .ZN(n9960) );
  OR2_X1 U9862 ( .A1(n9320), .A2(n9321), .ZN(n9962) );
  OR2_X1 U9863 ( .A1(n9963), .A2(n9964), .ZN(n9321) );
  AND2_X1 U9864 ( .A1(n9950), .A2(n9949), .ZN(n9964) );
  AND2_X1 U9865 ( .A1(n9947), .A2(n9965), .ZN(n9963) );
  OR2_X1 U9866 ( .A1(n9949), .A2(n9950), .ZN(n9965) );
  OR2_X1 U9867 ( .A1(n7730), .A2(n9631), .ZN(n9950) );
  OR2_X1 U9868 ( .A1(n9966), .A2(n9967), .ZN(n9949) );
  AND2_X1 U9869 ( .A1(n9946), .A2(n9945), .ZN(n9967) );
  AND2_X1 U9870 ( .A1(n9944), .A2(n9968), .ZN(n9966) );
  OR2_X1 U9871 ( .A1(n9945), .A2(n9946), .ZN(n9968) );
  OR2_X1 U9872 ( .A1(n9969), .A2(n9970), .ZN(n9946) );
  AND2_X1 U9873 ( .A1(n9942), .A2(n9941), .ZN(n9970) );
  AND2_X1 U9874 ( .A1(n9939), .A2(n9971), .ZN(n9969) );
  OR2_X1 U9875 ( .A1(n9941), .A2(n9942), .ZN(n9971) );
  OR2_X1 U9876 ( .A1(n7828), .A2(n9631), .ZN(n9942) );
  OR2_X1 U9877 ( .A1(n9972), .A2(n9973), .ZN(n9941) );
  AND2_X1 U9878 ( .A1(n9938), .A2(n9937), .ZN(n9973) );
  AND2_X1 U9879 ( .A1(n9935), .A2(n9974), .ZN(n9972) );
  OR2_X1 U9880 ( .A1(n9937), .A2(n9938), .ZN(n9974) );
  OR2_X1 U9881 ( .A1(n7887), .A2(n9631), .ZN(n9938) );
  OR2_X1 U9882 ( .A1(n9975), .A2(n9976), .ZN(n9937) );
  AND2_X1 U9883 ( .A1(n9934), .A2(n9933), .ZN(n9976) );
  AND2_X1 U9884 ( .A1(n9932), .A2(n9977), .ZN(n9975) );
  OR2_X1 U9885 ( .A1(n9933), .A2(n9934), .ZN(n9977) );
  OR2_X1 U9886 ( .A1(n9978), .A2(n9979), .ZN(n9934) );
  AND2_X1 U9887 ( .A1(n9930), .A2(n9929), .ZN(n9979) );
  AND2_X1 U9888 ( .A1(n9927), .A2(n9980), .ZN(n9978) );
  OR2_X1 U9889 ( .A1(n9929), .A2(n9930), .ZN(n9980) );
  OR2_X1 U9890 ( .A1(n8025), .A2(n9631), .ZN(n9930) );
  OR2_X1 U9891 ( .A1(n9981), .A2(n9982), .ZN(n9929) );
  AND2_X1 U9892 ( .A1(n9926), .A2(n9925), .ZN(n9982) );
  AND2_X1 U9893 ( .A1(n9923), .A2(n9983), .ZN(n9981) );
  OR2_X1 U9894 ( .A1(n9925), .A2(n9926), .ZN(n9983) );
  OR2_X1 U9895 ( .A1(n8107), .A2(n9631), .ZN(n9926) );
  OR2_X1 U9896 ( .A1(n9984), .A2(n9985), .ZN(n9925) );
  AND2_X1 U9897 ( .A1(n9922), .A2(n9921), .ZN(n9985) );
  AND2_X1 U9898 ( .A1(n9919), .A2(n9986), .ZN(n9984) );
  OR2_X1 U9899 ( .A1(n9921), .A2(n9922), .ZN(n9986) );
  OR2_X1 U9900 ( .A1(n8191), .A2(n9631), .ZN(n9922) );
  OR2_X1 U9901 ( .A1(n9987), .A2(n9988), .ZN(n9921) );
  AND2_X1 U9902 ( .A1(n9918), .A2(n9917), .ZN(n9988) );
  AND2_X1 U9903 ( .A1(n9916), .A2(n9989), .ZN(n9987) );
  OR2_X1 U9904 ( .A1(n9917), .A2(n9918), .ZN(n9989) );
  OR2_X1 U9905 ( .A1(n9990), .A2(n9991), .ZN(n9918) );
  AND2_X1 U9906 ( .A1(n9914), .A2(n9913), .ZN(n9991) );
  AND2_X1 U9907 ( .A1(n9911), .A2(n9992), .ZN(n9990) );
  OR2_X1 U9908 ( .A1(n9913), .A2(n9914), .ZN(n9992) );
  OR2_X1 U9909 ( .A1(n8608), .A2(n9631), .ZN(n9914) );
  OR2_X1 U9910 ( .A1(n9993), .A2(n9994), .ZN(n9913) );
  AND2_X1 U9911 ( .A1(n9910), .A2(n9909), .ZN(n9994) );
  AND2_X1 U9912 ( .A1(n9907), .A2(n9995), .ZN(n9993) );
  OR2_X1 U9913 ( .A1(n9909), .A2(n9910), .ZN(n9995) );
  OR2_X1 U9914 ( .A1(n8603), .A2(n9631), .ZN(n9910) );
  OR2_X1 U9915 ( .A1(n9996), .A2(n9997), .ZN(n9909) );
  AND2_X1 U9916 ( .A1(n9906), .A2(n9905), .ZN(n9997) );
  AND2_X1 U9917 ( .A1(n9903), .A2(n9998), .ZN(n9996) );
  OR2_X1 U9918 ( .A1(n9905), .A2(n9906), .ZN(n9998) );
  OR2_X1 U9919 ( .A1(n8598), .A2(n9631), .ZN(n9906) );
  OR2_X1 U9920 ( .A1(n9999), .A2(n10000), .ZN(n9905) );
  AND2_X1 U9921 ( .A1(n9902), .A2(n9901), .ZN(n10000) );
  AND2_X1 U9922 ( .A1(n9899), .A2(n10001), .ZN(n9999) );
  OR2_X1 U9923 ( .A1(n9901), .A2(n9902), .ZN(n10001) );
  OR2_X1 U9924 ( .A1(n8593), .A2(n9631), .ZN(n9902) );
  OR2_X1 U9925 ( .A1(n10002), .A2(n10003), .ZN(n9901) );
  AND2_X1 U9926 ( .A1(n9898), .A2(n9897), .ZN(n10003) );
  AND2_X1 U9927 ( .A1(n9895), .A2(n10004), .ZN(n10002) );
  OR2_X1 U9928 ( .A1(n9897), .A2(n9898), .ZN(n10004) );
  OR2_X1 U9929 ( .A1(n8588), .A2(n9631), .ZN(n9898) );
  OR2_X1 U9930 ( .A1(n10005), .A2(n10006), .ZN(n9897) );
  AND2_X1 U9931 ( .A1(n9894), .A2(n9893), .ZN(n10006) );
  AND2_X1 U9932 ( .A1(n9891), .A2(n10007), .ZN(n10005) );
  OR2_X1 U9933 ( .A1(n9893), .A2(n9894), .ZN(n10007) );
  OR2_X1 U9934 ( .A1(n8583), .A2(n9631), .ZN(n9894) );
  OR2_X1 U9935 ( .A1(n10008), .A2(n10009), .ZN(n9893) );
  AND2_X1 U9936 ( .A1(n9890), .A2(n9889), .ZN(n10009) );
  AND2_X1 U9937 ( .A1(n9887), .A2(n10010), .ZN(n10008) );
  OR2_X1 U9938 ( .A1(n9889), .A2(n9890), .ZN(n10010) );
  OR2_X1 U9939 ( .A1(n8578), .A2(n9631), .ZN(n9890) );
  OR2_X1 U9940 ( .A1(n10011), .A2(n10012), .ZN(n9889) );
  AND2_X1 U9941 ( .A1(n9886), .A2(n9885), .ZN(n10012) );
  AND2_X1 U9942 ( .A1(n9883), .A2(n10013), .ZN(n10011) );
  OR2_X1 U9943 ( .A1(n9885), .A2(n9886), .ZN(n10013) );
  OR2_X1 U9944 ( .A1(n8573), .A2(n9631), .ZN(n9886) );
  OR2_X1 U9945 ( .A1(n10014), .A2(n10015), .ZN(n9885) );
  AND2_X1 U9946 ( .A1(n9882), .A2(n9881), .ZN(n10015) );
  AND2_X1 U9947 ( .A1(n9879), .A2(n10016), .ZN(n10014) );
  OR2_X1 U9948 ( .A1(n9881), .A2(n9882), .ZN(n10016) );
  OR2_X1 U9949 ( .A1(n8568), .A2(n9631), .ZN(n9882) );
  OR2_X1 U9950 ( .A1(n10017), .A2(n10018), .ZN(n9881) );
  AND2_X1 U9951 ( .A1(n9878), .A2(n9877), .ZN(n10018) );
  AND2_X1 U9952 ( .A1(n9875), .A2(n10019), .ZN(n10017) );
  OR2_X1 U9953 ( .A1(n9877), .A2(n9878), .ZN(n10019) );
  OR2_X1 U9954 ( .A1(n8563), .A2(n9631), .ZN(n9878) );
  OR2_X1 U9955 ( .A1(n10020), .A2(n10021), .ZN(n9877) );
  AND2_X1 U9956 ( .A1(n9874), .A2(n9873), .ZN(n10021) );
  AND2_X1 U9957 ( .A1(n9871), .A2(n10022), .ZN(n10020) );
  OR2_X1 U9958 ( .A1(n9873), .A2(n9874), .ZN(n10022) );
  OR2_X1 U9959 ( .A1(n8558), .A2(n9631), .ZN(n9874) );
  OR2_X1 U9960 ( .A1(n10023), .A2(n10024), .ZN(n9873) );
  AND2_X1 U9961 ( .A1(n9870), .A2(n9869), .ZN(n10024) );
  AND2_X1 U9962 ( .A1(n9867), .A2(n10025), .ZN(n10023) );
  OR2_X1 U9963 ( .A1(n9869), .A2(n9870), .ZN(n10025) );
  OR2_X1 U9964 ( .A1(n8553), .A2(n9631), .ZN(n9870) );
  OR2_X1 U9965 ( .A1(n10026), .A2(n10027), .ZN(n9869) );
  AND2_X1 U9966 ( .A1(n9866), .A2(n9865), .ZN(n10027) );
  AND2_X1 U9967 ( .A1(n9863), .A2(n10028), .ZN(n10026) );
  OR2_X1 U9968 ( .A1(n9865), .A2(n9866), .ZN(n10028) );
  OR2_X1 U9969 ( .A1(n8548), .A2(n9631), .ZN(n9866) );
  OR2_X1 U9970 ( .A1(n10029), .A2(n10030), .ZN(n9865) );
  AND2_X1 U9971 ( .A1(n9860), .A2(n9862), .ZN(n10030) );
  AND2_X1 U9972 ( .A1(n10031), .A2(n9861), .ZN(n10029) );
  OR2_X1 U9973 ( .A1(n9862), .A2(n9860), .ZN(n10031) );
  XOR2_X1 U9974 ( .A(n10032), .B(n10033), .Z(n9860) );
  XOR2_X1 U9975 ( .A(n10034), .B(n10035), .Z(n10033) );
  OR2_X1 U9976 ( .A1(n10036), .A2(n10037), .ZN(n9862) );
  AND2_X1 U9977 ( .A1(n9858), .A2(n9857), .ZN(n10037) );
  AND2_X1 U9978 ( .A1(n9855), .A2(n10038), .ZN(n10036) );
  OR2_X1 U9979 ( .A1(n9857), .A2(n9858), .ZN(n10038) );
  OR2_X1 U9980 ( .A1(n8538), .A2(n9631), .ZN(n9858) );
  OR2_X1 U9981 ( .A1(n10039), .A2(n10040), .ZN(n9857) );
  AND2_X1 U9982 ( .A1(n9854), .A2(n9853), .ZN(n10040) );
  AND2_X1 U9983 ( .A1(n9851), .A2(n10041), .ZN(n10039) );
  OR2_X1 U9984 ( .A1(n9853), .A2(n9854), .ZN(n10041) );
  OR2_X1 U9985 ( .A1(n8533), .A2(n9631), .ZN(n9854) );
  OR2_X1 U9986 ( .A1(n10042), .A2(n10043), .ZN(n9853) );
  AND2_X1 U9987 ( .A1(n9850), .A2(n9849), .ZN(n10043) );
  AND2_X1 U9988 ( .A1(n9847), .A2(n10044), .ZN(n10042) );
  OR2_X1 U9989 ( .A1(n9849), .A2(n9850), .ZN(n10044) );
  OR2_X1 U9990 ( .A1(n8528), .A2(n9631), .ZN(n9850) );
  OR2_X1 U9991 ( .A1(n10045), .A2(n10046), .ZN(n9849) );
  AND2_X1 U9992 ( .A1(n9846), .A2(n9845), .ZN(n10046) );
  AND2_X1 U9993 ( .A1(n9843), .A2(n10047), .ZN(n10045) );
  OR2_X1 U9994 ( .A1(n9845), .A2(n9846), .ZN(n10047) );
  OR2_X1 U9995 ( .A1(n8523), .A2(n9631), .ZN(n9846) );
  OR2_X1 U9996 ( .A1(n10048), .A2(n10049), .ZN(n9845) );
  AND2_X1 U9997 ( .A1(n9840), .A2(n9841), .ZN(n10049) );
  AND2_X1 U9998 ( .A1(n10050), .A2(n10051), .ZN(n10048) );
  OR2_X1 U9999 ( .A1(n9841), .A2(n9840), .ZN(n10051) );
  OR2_X1 U10000 ( .A1(n8515), .A2(n9631), .ZN(n9840) );
  OR2_X1 U10001 ( .A1(n9631), .A2(n10052), .ZN(n9841) );
  INV_X1 U10002 ( .A(n9842), .ZN(n10050) );
  OR2_X1 U10003 ( .A1(n10053), .A2(n10054), .ZN(n9842) );
  AND2_X1 U10004 ( .A1(b_23_), .A2(n10055), .ZN(n10054) );
  OR2_X1 U10005 ( .A1(n10056), .A2(n7343), .ZN(n10055) );
  AND2_X1 U10006 ( .A1(a_30_), .A2(n10057), .ZN(n10056) );
  AND2_X1 U10007 ( .A1(b_22_), .A2(n10058), .ZN(n10053) );
  OR2_X1 U10008 ( .A1(n10059), .A2(n7347), .ZN(n10058) );
  AND2_X1 U10009 ( .A1(a_31_), .A2(n9836), .ZN(n10059) );
  XOR2_X1 U10010 ( .A(n10060), .B(n10061), .Z(n9843) );
  XNOR2_X1 U10011 ( .A(n10062), .B(n10063), .ZN(n10060) );
  XOR2_X1 U10012 ( .A(n10064), .B(n10065), .Z(n9847) );
  XOR2_X1 U10013 ( .A(n10066), .B(n10067), .Z(n10065) );
  XOR2_X1 U10014 ( .A(n10068), .B(n10069), .Z(n9851) );
  XOR2_X1 U10015 ( .A(n10070), .B(n10071), .Z(n10069) );
  XOR2_X1 U10016 ( .A(n10072), .B(n10073), .Z(n9855) );
  XOR2_X1 U10017 ( .A(n10074), .B(n10075), .Z(n10073) );
  XOR2_X1 U10018 ( .A(n10076), .B(n10077), .Z(n9863) );
  XOR2_X1 U10019 ( .A(n10078), .B(n10079), .Z(n10077) );
  XNOR2_X1 U10020 ( .A(n10080), .B(n10081), .ZN(n9867) );
  XNOR2_X1 U10021 ( .A(n10082), .B(n10083), .ZN(n10080) );
  XOR2_X1 U10022 ( .A(n10084), .B(n10085), .Z(n9871) );
  XOR2_X1 U10023 ( .A(n10086), .B(n10087), .Z(n10085) );
  XOR2_X1 U10024 ( .A(n10088), .B(n10089), .Z(n9875) );
  XOR2_X1 U10025 ( .A(n10090), .B(n10091), .Z(n10089) );
  XOR2_X1 U10026 ( .A(n10092), .B(n10093), .Z(n9879) );
  XOR2_X1 U10027 ( .A(n10094), .B(n10095), .Z(n10093) );
  XOR2_X1 U10028 ( .A(n10096), .B(n10097), .Z(n9883) );
  XOR2_X1 U10029 ( .A(n10098), .B(n10099), .Z(n10097) );
  XOR2_X1 U10030 ( .A(n10100), .B(n10101), .Z(n9887) );
  XOR2_X1 U10031 ( .A(n10102), .B(n10103), .Z(n10101) );
  XOR2_X1 U10032 ( .A(n10104), .B(n10105), .Z(n9891) );
  XOR2_X1 U10033 ( .A(n10106), .B(n10107), .Z(n10105) );
  XOR2_X1 U10034 ( .A(n10108), .B(n10109), .Z(n9895) );
  XOR2_X1 U10035 ( .A(n10110), .B(n10111), .Z(n10109) );
  XOR2_X1 U10036 ( .A(n10112), .B(n10113), .Z(n9899) );
  XOR2_X1 U10037 ( .A(n10114), .B(n10115), .Z(n10113) );
  XNOR2_X1 U10038 ( .A(n10116), .B(n10117), .ZN(n9903) );
  XNOR2_X1 U10039 ( .A(n10118), .B(n10119), .ZN(n10116) );
  XOR2_X1 U10040 ( .A(n10120), .B(n10121), .Z(n9907) );
  XOR2_X1 U10041 ( .A(n10122), .B(n10123), .Z(n10121) );
  XOR2_X1 U10042 ( .A(n10124), .B(n10125), .Z(n9911) );
  XOR2_X1 U10043 ( .A(n10126), .B(n10127), .Z(n10125) );
  OR2_X1 U10044 ( .A1(n8287), .A2(n9631), .ZN(n9917) );
  XOR2_X1 U10045 ( .A(n10128), .B(n10129), .Z(n9916) );
  XOR2_X1 U10046 ( .A(n10130), .B(n10131), .Z(n10129) );
  XNOR2_X1 U10047 ( .A(n10132), .B(n10133), .ZN(n9919) );
  XNOR2_X1 U10048 ( .A(n10134), .B(n10135), .ZN(n10132) );
  XOR2_X1 U10049 ( .A(n10136), .B(n10137), .Z(n9923) );
  XOR2_X1 U10050 ( .A(n10138), .B(n10139), .Z(n10137) );
  XOR2_X1 U10051 ( .A(n10140), .B(n10141), .Z(n9927) );
  XOR2_X1 U10052 ( .A(n10142), .B(n10143), .Z(n10141) );
  OR2_X1 U10053 ( .A1(n7955), .A2(n9631), .ZN(n9933) );
  XOR2_X1 U10054 ( .A(n10144), .B(n10145), .Z(n9932) );
  XOR2_X1 U10055 ( .A(n10146), .B(n10147), .Z(n10145) );
  XNOR2_X1 U10056 ( .A(n10148), .B(n10149), .ZN(n9935) );
  XNOR2_X1 U10057 ( .A(n10150), .B(n10151), .ZN(n10148) );
  XOR2_X1 U10058 ( .A(n10152), .B(n10153), .Z(n9939) );
  XOR2_X1 U10059 ( .A(n10154), .B(n10155), .Z(n10153) );
  OR2_X1 U10060 ( .A1(n7820), .A2(n9631), .ZN(n9945) );
  XOR2_X1 U10061 ( .A(n10156), .B(n10157), .Z(n9944) );
  XOR2_X1 U10062 ( .A(n10158), .B(n10159), .Z(n10157) );
  XOR2_X1 U10063 ( .A(n10160), .B(n10161), .Z(n9947) );
  XOR2_X1 U10064 ( .A(n10162), .B(n10163), .Z(n10161) );
  OR2_X1 U10065 ( .A1(n7697), .A2(n9631), .ZN(n9320) );
  XOR2_X1 U10066 ( .A(n10164), .B(n10165), .Z(n9319) );
  XOR2_X1 U10067 ( .A(n10166), .B(n10167), .Z(n10165) );
  XOR2_X1 U10068 ( .A(n10168), .B(n10169), .Z(n8371) );
  XOR2_X1 U10069 ( .A(n10170), .B(n10171), .Z(n10169) );
  XNOR2_X1 U10070 ( .A(n10172), .B(n10173), .ZN(n8354) );
  XOR2_X1 U10071 ( .A(n10174), .B(n10175), .Z(n10173) );
  OR2_X1 U10072 ( .A1(n9953), .A2(n7532), .ZN(n7529) );
  AND2_X1 U10073 ( .A1(n9953), .A2(n7532), .ZN(n8346) );
  XNOR2_X1 U10074 ( .A(n10176), .B(n10177), .ZN(n7532) );
  INV_X1 U10075 ( .A(n7531), .ZN(n9953) );
  OR2_X1 U10076 ( .A1(n9954), .A2(n9955), .ZN(n7531) );
  OR2_X1 U10077 ( .A1(n10178), .A2(n10179), .ZN(n9955) );
  AND2_X1 U10078 ( .A1(n10172), .A2(n10175), .ZN(n10179) );
  AND2_X1 U10079 ( .A1(n10180), .A2(n10174), .ZN(n10178) );
  OR2_X1 U10080 ( .A1(n10181), .A2(n10182), .ZN(n10174) );
  AND2_X1 U10081 ( .A1(n10171), .A2(n10170), .ZN(n10182) );
  AND2_X1 U10082 ( .A1(n10168), .A2(n10183), .ZN(n10181) );
  OR2_X1 U10083 ( .A1(n10171), .A2(n10170), .ZN(n10183) );
  OR2_X1 U10084 ( .A1(n10184), .A2(n10185), .ZN(n10170) );
  AND2_X1 U10085 ( .A1(n10167), .A2(n10166), .ZN(n10185) );
  AND2_X1 U10086 ( .A1(n10164), .A2(n10186), .ZN(n10184) );
  OR2_X1 U10087 ( .A1(n10167), .A2(n10166), .ZN(n10186) );
  OR2_X1 U10088 ( .A1(n10187), .A2(n10188), .ZN(n10166) );
  AND2_X1 U10089 ( .A1(n10163), .A2(n10162), .ZN(n10188) );
  AND2_X1 U10090 ( .A1(n10160), .A2(n10189), .ZN(n10187) );
  OR2_X1 U10091 ( .A1(n10163), .A2(n10162), .ZN(n10189) );
  OR2_X1 U10092 ( .A1(n10190), .A2(n10191), .ZN(n10162) );
  AND2_X1 U10093 ( .A1(n10159), .A2(n10158), .ZN(n10191) );
  AND2_X1 U10094 ( .A1(n10156), .A2(n10192), .ZN(n10190) );
  OR2_X1 U10095 ( .A1(n10159), .A2(n10158), .ZN(n10192) );
  OR2_X1 U10096 ( .A1(n10193), .A2(n10194), .ZN(n10158) );
  AND2_X1 U10097 ( .A1(n10155), .A2(n10154), .ZN(n10194) );
  AND2_X1 U10098 ( .A1(n10152), .A2(n10195), .ZN(n10193) );
  OR2_X1 U10099 ( .A1(n10155), .A2(n10154), .ZN(n10195) );
  OR2_X1 U10100 ( .A1(n10196), .A2(n10197), .ZN(n10154) );
  AND2_X1 U10101 ( .A1(n10151), .A2(n10150), .ZN(n10197) );
  AND2_X1 U10102 ( .A1(n10149), .A2(n10198), .ZN(n10196) );
  OR2_X1 U10103 ( .A1(n10151), .A2(n10150), .ZN(n10198) );
  OR2_X1 U10104 ( .A1(n7955), .A2(n9836), .ZN(n10150) );
  OR2_X1 U10105 ( .A1(n10199), .A2(n10200), .ZN(n10151) );
  AND2_X1 U10106 ( .A1(n10147), .A2(n10146), .ZN(n10200) );
  AND2_X1 U10107 ( .A1(n10144), .A2(n10201), .ZN(n10199) );
  OR2_X1 U10108 ( .A1(n10147), .A2(n10146), .ZN(n10201) );
  OR2_X1 U10109 ( .A1(n10202), .A2(n10203), .ZN(n10146) );
  AND2_X1 U10110 ( .A1(n10143), .A2(n10142), .ZN(n10203) );
  AND2_X1 U10111 ( .A1(n10140), .A2(n10204), .ZN(n10202) );
  OR2_X1 U10112 ( .A1(n10143), .A2(n10142), .ZN(n10204) );
  OR2_X1 U10113 ( .A1(n10205), .A2(n10206), .ZN(n10142) );
  AND2_X1 U10114 ( .A1(n10139), .A2(n10138), .ZN(n10206) );
  AND2_X1 U10115 ( .A1(n10136), .A2(n10207), .ZN(n10205) );
  OR2_X1 U10116 ( .A1(n10139), .A2(n10138), .ZN(n10207) );
  OR2_X1 U10117 ( .A1(n10208), .A2(n10209), .ZN(n10138) );
  AND2_X1 U10118 ( .A1(n10135), .A2(n10134), .ZN(n10209) );
  AND2_X1 U10119 ( .A1(n10133), .A2(n10210), .ZN(n10208) );
  OR2_X1 U10120 ( .A1(n10135), .A2(n10134), .ZN(n10210) );
  OR2_X1 U10121 ( .A1(n8287), .A2(n9836), .ZN(n10134) );
  OR2_X1 U10122 ( .A1(n10211), .A2(n10212), .ZN(n10135) );
  AND2_X1 U10123 ( .A1(n10131), .A2(n10130), .ZN(n10212) );
  AND2_X1 U10124 ( .A1(n10128), .A2(n10213), .ZN(n10211) );
  OR2_X1 U10125 ( .A1(n10131), .A2(n10130), .ZN(n10213) );
  OR2_X1 U10126 ( .A1(n10214), .A2(n10215), .ZN(n10130) );
  AND2_X1 U10127 ( .A1(n10127), .A2(n10126), .ZN(n10215) );
  AND2_X1 U10128 ( .A1(n10124), .A2(n10216), .ZN(n10214) );
  OR2_X1 U10129 ( .A1(n10127), .A2(n10126), .ZN(n10216) );
  OR2_X1 U10130 ( .A1(n10217), .A2(n10218), .ZN(n10126) );
  AND2_X1 U10131 ( .A1(n10123), .A2(n10122), .ZN(n10218) );
  AND2_X1 U10132 ( .A1(n10120), .A2(n10219), .ZN(n10217) );
  OR2_X1 U10133 ( .A1(n10123), .A2(n10122), .ZN(n10219) );
  OR2_X1 U10134 ( .A1(n10220), .A2(n10221), .ZN(n10122) );
  AND2_X1 U10135 ( .A1(n10119), .A2(n10118), .ZN(n10221) );
  AND2_X1 U10136 ( .A1(n10117), .A2(n10222), .ZN(n10220) );
  OR2_X1 U10137 ( .A1(n10119), .A2(n10118), .ZN(n10222) );
  OR2_X1 U10138 ( .A1(n8593), .A2(n9836), .ZN(n10118) );
  OR2_X1 U10139 ( .A1(n10223), .A2(n10224), .ZN(n10119) );
  AND2_X1 U10140 ( .A1(n10115), .A2(n10114), .ZN(n10224) );
  AND2_X1 U10141 ( .A1(n10112), .A2(n10225), .ZN(n10223) );
  OR2_X1 U10142 ( .A1(n10115), .A2(n10114), .ZN(n10225) );
  OR2_X1 U10143 ( .A1(n10226), .A2(n10227), .ZN(n10114) );
  AND2_X1 U10144 ( .A1(n10111), .A2(n10110), .ZN(n10227) );
  AND2_X1 U10145 ( .A1(n10108), .A2(n10228), .ZN(n10226) );
  OR2_X1 U10146 ( .A1(n10111), .A2(n10110), .ZN(n10228) );
  OR2_X1 U10147 ( .A1(n10229), .A2(n10230), .ZN(n10110) );
  AND2_X1 U10148 ( .A1(n10107), .A2(n10106), .ZN(n10230) );
  AND2_X1 U10149 ( .A1(n10104), .A2(n10231), .ZN(n10229) );
  OR2_X1 U10150 ( .A1(n10107), .A2(n10106), .ZN(n10231) );
  OR2_X1 U10151 ( .A1(n10232), .A2(n10233), .ZN(n10106) );
  AND2_X1 U10152 ( .A1(n10103), .A2(n10102), .ZN(n10233) );
  AND2_X1 U10153 ( .A1(n10100), .A2(n10234), .ZN(n10232) );
  OR2_X1 U10154 ( .A1(n10103), .A2(n10102), .ZN(n10234) );
  OR2_X1 U10155 ( .A1(n10235), .A2(n10236), .ZN(n10102) );
  AND2_X1 U10156 ( .A1(n10099), .A2(n10098), .ZN(n10236) );
  AND2_X1 U10157 ( .A1(n10096), .A2(n10237), .ZN(n10235) );
  OR2_X1 U10158 ( .A1(n10099), .A2(n10098), .ZN(n10237) );
  OR2_X1 U10159 ( .A1(n10238), .A2(n10239), .ZN(n10098) );
  AND2_X1 U10160 ( .A1(n10095), .A2(n10094), .ZN(n10239) );
  AND2_X1 U10161 ( .A1(n10092), .A2(n10240), .ZN(n10238) );
  OR2_X1 U10162 ( .A1(n10095), .A2(n10094), .ZN(n10240) );
  OR2_X1 U10163 ( .A1(n10241), .A2(n10242), .ZN(n10094) );
  AND2_X1 U10164 ( .A1(n10091), .A2(n10090), .ZN(n10242) );
  AND2_X1 U10165 ( .A1(n10088), .A2(n10243), .ZN(n10241) );
  OR2_X1 U10166 ( .A1(n10091), .A2(n10090), .ZN(n10243) );
  OR2_X1 U10167 ( .A1(n10244), .A2(n10245), .ZN(n10090) );
  AND2_X1 U10168 ( .A1(n10087), .A2(n10086), .ZN(n10245) );
  AND2_X1 U10169 ( .A1(n10084), .A2(n10246), .ZN(n10244) );
  OR2_X1 U10170 ( .A1(n10087), .A2(n10086), .ZN(n10246) );
  OR2_X1 U10171 ( .A1(n10247), .A2(n10248), .ZN(n10086) );
  AND2_X1 U10172 ( .A1(n10081), .A2(n10083), .ZN(n10248) );
  AND2_X1 U10173 ( .A1(n10249), .A2(n10082), .ZN(n10247) );
  OR2_X1 U10174 ( .A1(n10081), .A2(n10083), .ZN(n10249) );
  OR2_X1 U10175 ( .A1(n10250), .A2(n10251), .ZN(n10083) );
  AND2_X1 U10176 ( .A1(n10079), .A2(n10078), .ZN(n10251) );
  AND2_X1 U10177 ( .A1(n10076), .A2(n10252), .ZN(n10250) );
  OR2_X1 U10178 ( .A1(n10079), .A2(n10078), .ZN(n10252) );
  OR2_X1 U10179 ( .A1(n10253), .A2(n10254), .ZN(n10078) );
  AND2_X1 U10180 ( .A1(n10035), .A2(n10034), .ZN(n10254) );
  AND2_X1 U10181 ( .A1(n10032), .A2(n10255), .ZN(n10253) );
  OR2_X1 U10182 ( .A1(n10035), .A2(n10034), .ZN(n10255) );
  OR2_X1 U10183 ( .A1(n10256), .A2(n10257), .ZN(n10034) );
  AND2_X1 U10184 ( .A1(n10075), .A2(n10074), .ZN(n10257) );
  AND2_X1 U10185 ( .A1(n10072), .A2(n10258), .ZN(n10256) );
  OR2_X1 U10186 ( .A1(n10075), .A2(n10074), .ZN(n10258) );
  OR2_X1 U10187 ( .A1(n10259), .A2(n10260), .ZN(n10074) );
  AND2_X1 U10188 ( .A1(n10071), .A2(n10070), .ZN(n10260) );
  AND2_X1 U10189 ( .A1(n10068), .A2(n10261), .ZN(n10259) );
  OR2_X1 U10190 ( .A1(n10071), .A2(n10070), .ZN(n10261) );
  OR2_X1 U10191 ( .A1(n10262), .A2(n10263), .ZN(n10070) );
  AND2_X1 U10192 ( .A1(n10067), .A2(n10066), .ZN(n10263) );
  AND2_X1 U10193 ( .A1(n10064), .A2(n10264), .ZN(n10262) );
  OR2_X1 U10194 ( .A1(n10067), .A2(n10066), .ZN(n10264) );
  OR2_X1 U10195 ( .A1(n10265), .A2(n10266), .ZN(n10066) );
  AND2_X1 U10196 ( .A1(n10061), .A2(n10062), .ZN(n10266) );
  AND2_X1 U10197 ( .A1(n10267), .A2(n10268), .ZN(n10265) );
  OR2_X1 U10198 ( .A1(n10061), .A2(n10062), .ZN(n10268) );
  OR2_X1 U10199 ( .A1(n10057), .A2(n10052), .ZN(n10062) );
  OR2_X1 U10200 ( .A1(n8956), .A2(n9836), .ZN(n10052) );
  OR2_X1 U10201 ( .A1(n8515), .A2(n9836), .ZN(n10061) );
  INV_X1 U10202 ( .A(n10063), .ZN(n10267) );
  OR2_X1 U10203 ( .A1(n10269), .A2(n10270), .ZN(n10063) );
  AND2_X1 U10204 ( .A1(b_22_), .A2(n10271), .ZN(n10270) );
  OR2_X1 U10205 ( .A1(n10272), .A2(n7343), .ZN(n10271) );
  AND2_X1 U10206 ( .A1(a_30_), .A2(n10273), .ZN(n10272) );
  AND2_X1 U10207 ( .A1(b_21_), .A2(n10274), .ZN(n10269) );
  OR2_X1 U10208 ( .A1(n10275), .A2(n7347), .ZN(n10274) );
  AND2_X1 U10209 ( .A1(a_31_), .A2(n10057), .ZN(n10275) );
  OR2_X1 U10210 ( .A1(n8523), .A2(n9836), .ZN(n10067) );
  XOR2_X1 U10211 ( .A(n10276), .B(n10277), .Z(n10064) );
  XNOR2_X1 U10212 ( .A(n10278), .B(n10279), .ZN(n10276) );
  OR2_X1 U10213 ( .A1(n8528), .A2(n9836), .ZN(n10071) );
  XOR2_X1 U10214 ( .A(n10280), .B(n10281), .Z(n10068) );
  XOR2_X1 U10215 ( .A(n10282), .B(n10283), .Z(n10281) );
  OR2_X1 U10216 ( .A1(n8533), .A2(n9836), .ZN(n10075) );
  XOR2_X1 U10217 ( .A(n10284), .B(n10285), .Z(n10072) );
  XOR2_X1 U10218 ( .A(n10286), .B(n10287), .Z(n10285) );
  OR2_X1 U10219 ( .A1(n8538), .A2(n9836), .ZN(n10035) );
  XOR2_X1 U10220 ( .A(n10288), .B(n10289), .Z(n10032) );
  XOR2_X1 U10221 ( .A(n10290), .B(n10291), .Z(n10289) );
  OR2_X1 U10222 ( .A1(n8543), .A2(n9836), .ZN(n10079) );
  XOR2_X1 U10223 ( .A(n10292), .B(n10293), .Z(n10076) );
  XOR2_X1 U10224 ( .A(n10294), .B(n10295), .Z(n10293) );
  XOR2_X1 U10225 ( .A(n10296), .B(n10297), .Z(n10081) );
  XOR2_X1 U10226 ( .A(n10298), .B(n10299), .Z(n10297) );
  OR2_X1 U10227 ( .A1(n8553), .A2(n9836), .ZN(n10087) );
  XOR2_X1 U10228 ( .A(n10300), .B(n10301), .Z(n10084) );
  XOR2_X1 U10229 ( .A(n10302), .B(n10303), .Z(n10301) );
  OR2_X1 U10230 ( .A1(n8558), .A2(n9836), .ZN(n10091) );
  XNOR2_X1 U10231 ( .A(n10304), .B(n10305), .ZN(n10088) );
  XNOR2_X1 U10232 ( .A(n10306), .B(n10307), .ZN(n10304) );
  OR2_X1 U10233 ( .A1(n8563), .A2(n9836), .ZN(n10095) );
  XOR2_X1 U10234 ( .A(n10308), .B(n10309), .Z(n10092) );
  XOR2_X1 U10235 ( .A(n10310), .B(n10311), .Z(n10309) );
  OR2_X1 U10236 ( .A1(n8568), .A2(n9836), .ZN(n10099) );
  XOR2_X1 U10237 ( .A(n10312), .B(n10313), .Z(n10096) );
  XOR2_X1 U10238 ( .A(n10314), .B(n10315), .Z(n10313) );
  OR2_X1 U10239 ( .A1(n8573), .A2(n9836), .ZN(n10103) );
  XOR2_X1 U10240 ( .A(n10316), .B(n10317), .Z(n10100) );
  XOR2_X1 U10241 ( .A(n10318), .B(n10319), .Z(n10317) );
  OR2_X1 U10242 ( .A1(n8578), .A2(n9836), .ZN(n10107) );
  XOR2_X1 U10243 ( .A(n10320), .B(n10321), .Z(n10104) );
  XOR2_X1 U10244 ( .A(n10322), .B(n10323), .Z(n10321) );
  OR2_X1 U10245 ( .A1(n8583), .A2(n9836), .ZN(n10111) );
  XOR2_X1 U10246 ( .A(n10324), .B(n10325), .Z(n10108) );
  XOR2_X1 U10247 ( .A(n10326), .B(n10327), .Z(n10325) );
  OR2_X1 U10248 ( .A1(n8588), .A2(n9836), .ZN(n10115) );
  XOR2_X1 U10249 ( .A(n10328), .B(n10329), .Z(n10112) );
  XOR2_X1 U10250 ( .A(n10330), .B(n10331), .Z(n10329) );
  XOR2_X1 U10251 ( .A(n10332), .B(n10333), .Z(n10117) );
  XOR2_X1 U10252 ( .A(n10334), .B(n10335), .Z(n10333) );
  OR2_X1 U10253 ( .A1(n8598), .A2(n9836), .ZN(n10123) );
  XOR2_X1 U10254 ( .A(n10336), .B(n10337), .Z(n10120) );
  XOR2_X1 U10255 ( .A(n10338), .B(n10339), .Z(n10337) );
  OR2_X1 U10256 ( .A1(n8603), .A2(n9836), .ZN(n10127) );
  XOR2_X1 U10257 ( .A(n10340), .B(n10341), .Z(n10124) );
  XOR2_X1 U10258 ( .A(n10342), .B(n10343), .Z(n10341) );
  OR2_X1 U10259 ( .A1(n8608), .A2(n9836), .ZN(n10131) );
  XOR2_X1 U10260 ( .A(n10344), .B(n10345), .Z(n10128) );
  XOR2_X1 U10261 ( .A(n10346), .B(n10347), .Z(n10345) );
  XOR2_X1 U10262 ( .A(n10348), .B(n10349), .Z(n10133) );
  XOR2_X1 U10263 ( .A(n10350), .B(n10351), .Z(n10349) );
  OR2_X1 U10264 ( .A1(n8191), .A2(n9836), .ZN(n10139) );
  XOR2_X1 U10265 ( .A(n10352), .B(n10353), .Z(n10136) );
  XOR2_X1 U10266 ( .A(n10354), .B(n10355), .Z(n10353) );
  OR2_X1 U10267 ( .A1(n8107), .A2(n9836), .ZN(n10143) );
  XOR2_X1 U10268 ( .A(n10356), .B(n10357), .Z(n10140) );
  XOR2_X1 U10269 ( .A(n10358), .B(n10359), .Z(n10357) );
  OR2_X1 U10270 ( .A1(n8025), .A2(n9836), .ZN(n10147) );
  XOR2_X1 U10271 ( .A(n10360), .B(n10361), .Z(n10144) );
  XOR2_X1 U10272 ( .A(n10362), .B(n10363), .Z(n10361) );
  XOR2_X1 U10273 ( .A(n10364), .B(n10365), .Z(n10149) );
  XOR2_X1 U10274 ( .A(n10366), .B(n10367), .Z(n10365) );
  OR2_X1 U10275 ( .A1(n7887), .A2(n9836), .ZN(n10155) );
  XOR2_X1 U10276 ( .A(n10368), .B(n10369), .Z(n10152) );
  XOR2_X1 U10277 ( .A(n10370), .B(n10371), .Z(n10369) );
  OR2_X1 U10278 ( .A1(n7828), .A2(n9836), .ZN(n10159) );
  XOR2_X1 U10279 ( .A(n10372), .B(n10373), .Z(n10156) );
  XOR2_X1 U10280 ( .A(n10374), .B(n10375), .Z(n10373) );
  OR2_X1 U10281 ( .A1(n7820), .A2(n9836), .ZN(n10163) );
  XOR2_X1 U10282 ( .A(n10376), .B(n10377), .Z(n10160) );
  XOR2_X1 U10283 ( .A(n10378), .B(n10379), .Z(n10377) );
  OR2_X1 U10284 ( .A1(n7730), .A2(n9836), .ZN(n10167) );
  XOR2_X1 U10285 ( .A(n10380), .B(n10381), .Z(n10164) );
  XOR2_X1 U10286 ( .A(n10382), .B(n10383), .Z(n10381) );
  OR2_X1 U10287 ( .A1(n7697), .A2(n9836), .ZN(n10171) );
  XOR2_X1 U10288 ( .A(n10384), .B(n10385), .Z(n10168) );
  XOR2_X1 U10289 ( .A(n10386), .B(n10387), .Z(n10385) );
  OR2_X1 U10290 ( .A1(n10172), .A2(n10175), .ZN(n10180) );
  OR2_X1 U10291 ( .A1(n7660), .A2(n9836), .ZN(n10175) );
  XOR2_X1 U10292 ( .A(n10388), .B(n10389), .Z(n10172) );
  XOR2_X1 U10293 ( .A(n10390), .B(n10391), .Z(n10389) );
  XOR2_X1 U10294 ( .A(n10392), .B(n10393), .Z(n9954) );
  XOR2_X1 U10295 ( .A(n10394), .B(n10395), .Z(n10393) );
  OR2_X1 U10296 ( .A1(n8345), .A2(n8344), .ZN(n7535) );
  AND2_X1 U10297 ( .A1(n10396), .A2(n8326), .ZN(n8344) );
  OR2_X1 U10298 ( .A1(n10397), .A2(n10398), .ZN(n8326) );
  INV_X1 U10299 ( .A(n10399), .ZN(n10396) );
  AND2_X1 U10300 ( .A1(n10397), .A2(n10398), .ZN(n10399) );
  OR2_X1 U10301 ( .A1(n10400), .A2(n10401), .ZN(n10398) );
  AND2_X1 U10302 ( .A1(n10402), .A2(n10403), .ZN(n10401) );
  AND2_X1 U10303 ( .A1(n10404), .A2(n10405), .ZN(n10400) );
  OR2_X1 U10304 ( .A1(n10402), .A2(n10403), .ZN(n10404) );
  XOR2_X1 U10305 ( .A(n8335), .B(n10406), .Z(n10397) );
  XOR2_X1 U10306 ( .A(n8338), .B(n8336), .Z(n10406) );
  OR2_X1 U10307 ( .A1(n7660), .A2(n10407), .ZN(n8336) );
  OR2_X1 U10308 ( .A1(n10408), .A2(n10409), .ZN(n8338) );
  AND2_X1 U10309 ( .A1(n10410), .A2(n10411), .ZN(n10409) );
  AND2_X1 U10310 ( .A1(n10412), .A2(n10413), .ZN(n10408) );
  OR2_X1 U10311 ( .A1(n10410), .A2(n10411), .ZN(n10412) );
  XOR2_X1 U10312 ( .A(n10414), .B(n10415), .Z(n8335) );
  XOR2_X1 U10313 ( .A(n10416), .B(n10417), .Z(n10415) );
  AND2_X1 U10314 ( .A1(n10176), .A2(n10418), .ZN(n8345) );
  INV_X1 U10315 ( .A(n10177), .ZN(n10418) );
  OR2_X1 U10316 ( .A1(n10419), .A2(n10420), .ZN(n10177) );
  AND2_X1 U10317 ( .A1(n10392), .A2(n10395), .ZN(n10420) );
  AND2_X1 U10318 ( .A1(n10421), .A2(n10394), .ZN(n10419) );
  OR2_X1 U10319 ( .A1(n10422), .A2(n10423), .ZN(n10394) );
  AND2_X1 U10320 ( .A1(n10388), .A2(n10391), .ZN(n10423) );
  AND2_X1 U10321 ( .A1(n10424), .A2(n10390), .ZN(n10422) );
  OR2_X1 U10322 ( .A1(n10425), .A2(n10426), .ZN(n10390) );
  AND2_X1 U10323 ( .A1(n10384), .A2(n10387), .ZN(n10426) );
  AND2_X1 U10324 ( .A1(n10427), .A2(n10386), .ZN(n10425) );
  OR2_X1 U10325 ( .A1(n10428), .A2(n10429), .ZN(n10386) );
  AND2_X1 U10326 ( .A1(n10383), .A2(n10382), .ZN(n10429) );
  AND2_X1 U10327 ( .A1(n10380), .A2(n10430), .ZN(n10428) );
  OR2_X1 U10328 ( .A1(n10382), .A2(n10383), .ZN(n10430) );
  OR2_X1 U10329 ( .A1(n7820), .A2(n10057), .ZN(n10383) );
  OR2_X1 U10330 ( .A1(n10431), .A2(n10432), .ZN(n10382) );
  AND2_X1 U10331 ( .A1(n10379), .A2(n10378), .ZN(n10432) );
  AND2_X1 U10332 ( .A1(n10376), .A2(n10433), .ZN(n10431) );
  OR2_X1 U10333 ( .A1(n10378), .A2(n10379), .ZN(n10433) );
  OR2_X1 U10334 ( .A1(n7828), .A2(n10057), .ZN(n10379) );
  OR2_X1 U10335 ( .A1(n10434), .A2(n10435), .ZN(n10378) );
  AND2_X1 U10336 ( .A1(n10375), .A2(n10374), .ZN(n10435) );
  AND2_X1 U10337 ( .A1(n10372), .A2(n10436), .ZN(n10434) );
  OR2_X1 U10338 ( .A1(n10374), .A2(n10375), .ZN(n10436) );
  OR2_X1 U10339 ( .A1(n7887), .A2(n10057), .ZN(n10375) );
  OR2_X1 U10340 ( .A1(n10437), .A2(n10438), .ZN(n10374) );
  AND2_X1 U10341 ( .A1(n10371), .A2(n10370), .ZN(n10438) );
  AND2_X1 U10342 ( .A1(n10368), .A2(n10439), .ZN(n10437) );
  OR2_X1 U10343 ( .A1(n10370), .A2(n10371), .ZN(n10439) );
  OR2_X1 U10344 ( .A1(n7955), .A2(n10057), .ZN(n10371) );
  OR2_X1 U10345 ( .A1(n10440), .A2(n10441), .ZN(n10370) );
  AND2_X1 U10346 ( .A1(n10367), .A2(n10366), .ZN(n10441) );
  AND2_X1 U10347 ( .A1(n10364), .A2(n10442), .ZN(n10440) );
  OR2_X1 U10348 ( .A1(n10366), .A2(n10367), .ZN(n10442) );
  OR2_X1 U10349 ( .A1(n8025), .A2(n10057), .ZN(n10367) );
  OR2_X1 U10350 ( .A1(n10443), .A2(n10444), .ZN(n10366) );
  AND2_X1 U10351 ( .A1(n10363), .A2(n10362), .ZN(n10444) );
  AND2_X1 U10352 ( .A1(n10360), .A2(n10445), .ZN(n10443) );
  OR2_X1 U10353 ( .A1(n10362), .A2(n10363), .ZN(n10445) );
  OR2_X1 U10354 ( .A1(n8107), .A2(n10057), .ZN(n10363) );
  OR2_X1 U10355 ( .A1(n10446), .A2(n10447), .ZN(n10362) );
  AND2_X1 U10356 ( .A1(n10359), .A2(n10358), .ZN(n10447) );
  AND2_X1 U10357 ( .A1(n10356), .A2(n10448), .ZN(n10446) );
  OR2_X1 U10358 ( .A1(n10358), .A2(n10359), .ZN(n10448) );
  OR2_X1 U10359 ( .A1(n8191), .A2(n10057), .ZN(n10359) );
  OR2_X1 U10360 ( .A1(n10449), .A2(n10450), .ZN(n10358) );
  AND2_X1 U10361 ( .A1(n10355), .A2(n10354), .ZN(n10450) );
  AND2_X1 U10362 ( .A1(n10352), .A2(n10451), .ZN(n10449) );
  OR2_X1 U10363 ( .A1(n10354), .A2(n10355), .ZN(n10451) );
  OR2_X1 U10364 ( .A1(n8287), .A2(n10057), .ZN(n10355) );
  OR2_X1 U10365 ( .A1(n10452), .A2(n10453), .ZN(n10354) );
  AND2_X1 U10366 ( .A1(n10351), .A2(n10350), .ZN(n10453) );
  AND2_X1 U10367 ( .A1(n10348), .A2(n10454), .ZN(n10452) );
  OR2_X1 U10368 ( .A1(n10350), .A2(n10351), .ZN(n10454) );
  OR2_X1 U10369 ( .A1(n8608), .A2(n10057), .ZN(n10351) );
  OR2_X1 U10370 ( .A1(n10455), .A2(n10456), .ZN(n10350) );
  AND2_X1 U10371 ( .A1(n10347), .A2(n10346), .ZN(n10456) );
  AND2_X1 U10372 ( .A1(n10344), .A2(n10457), .ZN(n10455) );
  OR2_X1 U10373 ( .A1(n10346), .A2(n10347), .ZN(n10457) );
  OR2_X1 U10374 ( .A1(n8603), .A2(n10057), .ZN(n10347) );
  OR2_X1 U10375 ( .A1(n10458), .A2(n10459), .ZN(n10346) );
  AND2_X1 U10376 ( .A1(n10343), .A2(n10342), .ZN(n10459) );
  AND2_X1 U10377 ( .A1(n10340), .A2(n10460), .ZN(n10458) );
  OR2_X1 U10378 ( .A1(n10342), .A2(n10343), .ZN(n10460) );
  OR2_X1 U10379 ( .A1(n8598), .A2(n10057), .ZN(n10343) );
  OR2_X1 U10380 ( .A1(n10461), .A2(n10462), .ZN(n10342) );
  AND2_X1 U10381 ( .A1(n10339), .A2(n10338), .ZN(n10462) );
  AND2_X1 U10382 ( .A1(n10336), .A2(n10463), .ZN(n10461) );
  OR2_X1 U10383 ( .A1(n10338), .A2(n10339), .ZN(n10463) );
  OR2_X1 U10384 ( .A1(n8593), .A2(n10057), .ZN(n10339) );
  OR2_X1 U10385 ( .A1(n10464), .A2(n10465), .ZN(n10338) );
  AND2_X1 U10386 ( .A1(n10335), .A2(n10334), .ZN(n10465) );
  AND2_X1 U10387 ( .A1(n10332), .A2(n10466), .ZN(n10464) );
  OR2_X1 U10388 ( .A1(n10334), .A2(n10335), .ZN(n10466) );
  OR2_X1 U10389 ( .A1(n8588), .A2(n10057), .ZN(n10335) );
  OR2_X1 U10390 ( .A1(n10467), .A2(n10468), .ZN(n10334) );
  AND2_X1 U10391 ( .A1(n10331), .A2(n10330), .ZN(n10468) );
  AND2_X1 U10392 ( .A1(n10328), .A2(n10469), .ZN(n10467) );
  OR2_X1 U10393 ( .A1(n10330), .A2(n10331), .ZN(n10469) );
  OR2_X1 U10394 ( .A1(n8583), .A2(n10057), .ZN(n10331) );
  OR2_X1 U10395 ( .A1(n10470), .A2(n10471), .ZN(n10330) );
  AND2_X1 U10396 ( .A1(n10327), .A2(n10326), .ZN(n10471) );
  AND2_X1 U10397 ( .A1(n10324), .A2(n10472), .ZN(n10470) );
  OR2_X1 U10398 ( .A1(n10326), .A2(n10327), .ZN(n10472) );
  OR2_X1 U10399 ( .A1(n8578), .A2(n10057), .ZN(n10327) );
  OR2_X1 U10400 ( .A1(n10473), .A2(n10474), .ZN(n10326) );
  AND2_X1 U10401 ( .A1(n10323), .A2(n10322), .ZN(n10474) );
  AND2_X1 U10402 ( .A1(n10320), .A2(n10475), .ZN(n10473) );
  OR2_X1 U10403 ( .A1(n10322), .A2(n10323), .ZN(n10475) );
  OR2_X1 U10404 ( .A1(n8573), .A2(n10057), .ZN(n10323) );
  OR2_X1 U10405 ( .A1(n10476), .A2(n10477), .ZN(n10322) );
  AND2_X1 U10406 ( .A1(n10319), .A2(n10318), .ZN(n10477) );
  AND2_X1 U10407 ( .A1(n10316), .A2(n10478), .ZN(n10476) );
  OR2_X1 U10408 ( .A1(n10318), .A2(n10319), .ZN(n10478) );
  OR2_X1 U10409 ( .A1(n8568), .A2(n10057), .ZN(n10319) );
  OR2_X1 U10410 ( .A1(n10479), .A2(n10480), .ZN(n10318) );
  AND2_X1 U10411 ( .A1(n10315), .A2(n10314), .ZN(n10480) );
  AND2_X1 U10412 ( .A1(n10312), .A2(n10481), .ZN(n10479) );
  OR2_X1 U10413 ( .A1(n10314), .A2(n10315), .ZN(n10481) );
  OR2_X1 U10414 ( .A1(n8563), .A2(n10057), .ZN(n10315) );
  OR2_X1 U10415 ( .A1(n10482), .A2(n10483), .ZN(n10314) );
  AND2_X1 U10416 ( .A1(n10311), .A2(n10310), .ZN(n10483) );
  AND2_X1 U10417 ( .A1(n10308), .A2(n10484), .ZN(n10482) );
  OR2_X1 U10418 ( .A1(n10310), .A2(n10311), .ZN(n10484) );
  OR2_X1 U10419 ( .A1(n8558), .A2(n10057), .ZN(n10311) );
  OR2_X1 U10420 ( .A1(n10485), .A2(n10486), .ZN(n10310) );
  AND2_X1 U10421 ( .A1(n10305), .A2(n10307), .ZN(n10486) );
  AND2_X1 U10422 ( .A1(n10487), .A2(n10306), .ZN(n10485) );
  OR2_X1 U10423 ( .A1(n10307), .A2(n10305), .ZN(n10487) );
  XOR2_X1 U10424 ( .A(n10488), .B(n10489), .Z(n10305) );
  XOR2_X1 U10425 ( .A(n10490), .B(n10491), .Z(n10489) );
  OR2_X1 U10426 ( .A1(n10492), .A2(n10493), .ZN(n10307) );
  AND2_X1 U10427 ( .A1(n10303), .A2(n10302), .ZN(n10493) );
  AND2_X1 U10428 ( .A1(n10300), .A2(n10494), .ZN(n10492) );
  OR2_X1 U10429 ( .A1(n10302), .A2(n10303), .ZN(n10494) );
  OR2_X1 U10430 ( .A1(n8548), .A2(n10057), .ZN(n10303) );
  OR2_X1 U10431 ( .A1(n10495), .A2(n10496), .ZN(n10302) );
  AND2_X1 U10432 ( .A1(n10299), .A2(n10298), .ZN(n10496) );
  AND2_X1 U10433 ( .A1(n10296), .A2(n10497), .ZN(n10495) );
  OR2_X1 U10434 ( .A1(n10298), .A2(n10299), .ZN(n10497) );
  OR2_X1 U10435 ( .A1(n8543), .A2(n10057), .ZN(n10299) );
  OR2_X1 U10436 ( .A1(n10498), .A2(n10499), .ZN(n10298) );
  AND2_X1 U10437 ( .A1(n10295), .A2(n10294), .ZN(n10499) );
  AND2_X1 U10438 ( .A1(n10292), .A2(n10500), .ZN(n10498) );
  OR2_X1 U10439 ( .A1(n10294), .A2(n10295), .ZN(n10500) );
  OR2_X1 U10440 ( .A1(n8538), .A2(n10057), .ZN(n10295) );
  OR2_X1 U10441 ( .A1(n10501), .A2(n10502), .ZN(n10294) );
  AND2_X1 U10442 ( .A1(n10291), .A2(n10290), .ZN(n10502) );
  AND2_X1 U10443 ( .A1(n10288), .A2(n10503), .ZN(n10501) );
  OR2_X1 U10444 ( .A1(n10290), .A2(n10291), .ZN(n10503) );
  OR2_X1 U10445 ( .A1(n8533), .A2(n10057), .ZN(n10291) );
  OR2_X1 U10446 ( .A1(n10504), .A2(n10505), .ZN(n10290) );
  AND2_X1 U10447 ( .A1(n10287), .A2(n10286), .ZN(n10505) );
  AND2_X1 U10448 ( .A1(n10284), .A2(n10506), .ZN(n10504) );
  OR2_X1 U10449 ( .A1(n10286), .A2(n10287), .ZN(n10506) );
  OR2_X1 U10450 ( .A1(n8528), .A2(n10057), .ZN(n10287) );
  OR2_X1 U10451 ( .A1(n10507), .A2(n10508), .ZN(n10286) );
  AND2_X1 U10452 ( .A1(n10283), .A2(n10282), .ZN(n10508) );
  AND2_X1 U10453 ( .A1(n10280), .A2(n10509), .ZN(n10507) );
  OR2_X1 U10454 ( .A1(n10282), .A2(n10283), .ZN(n10509) );
  OR2_X1 U10455 ( .A1(n8523), .A2(n10057), .ZN(n10283) );
  OR2_X1 U10456 ( .A1(n10510), .A2(n10511), .ZN(n10282) );
  AND2_X1 U10457 ( .A1(n10277), .A2(n10278), .ZN(n10511) );
  AND2_X1 U10458 ( .A1(n10512), .A2(n10513), .ZN(n10510) );
  OR2_X1 U10459 ( .A1(n10278), .A2(n10277), .ZN(n10513) );
  OR2_X1 U10460 ( .A1(n8515), .A2(n10057), .ZN(n10277) );
  OR2_X1 U10461 ( .A1(n10057), .A2(n10514), .ZN(n10278) );
  OR2_X1 U10462 ( .A1(n8956), .A2(n10273), .ZN(n10514) );
  INV_X1 U10463 ( .A(n10279), .ZN(n10512) );
  OR2_X1 U10464 ( .A1(n10515), .A2(n10516), .ZN(n10279) );
  AND2_X1 U10465 ( .A1(b_21_), .A2(n10517), .ZN(n10516) );
  OR2_X1 U10466 ( .A1(n10518), .A2(n7343), .ZN(n10517) );
  AND2_X1 U10467 ( .A1(a_30_), .A2(n10407), .ZN(n10518) );
  AND2_X1 U10468 ( .A1(b_20_), .A2(n10519), .ZN(n10515) );
  OR2_X1 U10469 ( .A1(n10520), .A2(n7347), .ZN(n10519) );
  AND2_X1 U10470 ( .A1(a_31_), .A2(n10273), .ZN(n10520) );
  XOR2_X1 U10471 ( .A(n10521), .B(n10522), .Z(n10280) );
  XNOR2_X1 U10472 ( .A(n10523), .B(n10524), .ZN(n10521) );
  XOR2_X1 U10473 ( .A(n10525), .B(n10526), .Z(n10284) );
  XOR2_X1 U10474 ( .A(n10527), .B(n10528), .Z(n10526) );
  XOR2_X1 U10475 ( .A(n10529), .B(n10530), .Z(n10288) );
  XOR2_X1 U10476 ( .A(n10531), .B(n10532), .Z(n10530) );
  XOR2_X1 U10477 ( .A(n10533), .B(n10534), .Z(n10292) );
  XOR2_X1 U10478 ( .A(n10535), .B(n10536), .Z(n10534) );
  XOR2_X1 U10479 ( .A(n10537), .B(n10538), .Z(n10296) );
  XOR2_X1 U10480 ( .A(n10539), .B(n10540), .Z(n10538) );
  XOR2_X1 U10481 ( .A(n10541), .B(n10542), .Z(n10300) );
  XOR2_X1 U10482 ( .A(n10543), .B(n10544), .Z(n10542) );
  XOR2_X1 U10483 ( .A(n10545), .B(n10546), .Z(n10308) );
  XOR2_X1 U10484 ( .A(n10547), .B(n10548), .Z(n10546) );
  XNOR2_X1 U10485 ( .A(n10549), .B(n10550), .ZN(n10312) );
  XNOR2_X1 U10486 ( .A(n10551), .B(n10552), .ZN(n10549) );
  XOR2_X1 U10487 ( .A(n10553), .B(n10554), .Z(n10316) );
  XOR2_X1 U10488 ( .A(n10555), .B(n10556), .Z(n10554) );
  XOR2_X1 U10489 ( .A(n10557), .B(n10558), .Z(n10320) );
  XOR2_X1 U10490 ( .A(n10559), .B(n10560), .Z(n10558) );
  XOR2_X1 U10491 ( .A(n10561), .B(n10562), .Z(n10324) );
  XOR2_X1 U10492 ( .A(n10563), .B(n10564), .Z(n10562) );
  XOR2_X1 U10493 ( .A(n10565), .B(n10566), .Z(n10328) );
  XOR2_X1 U10494 ( .A(n10567), .B(n10568), .Z(n10566) );
  XOR2_X1 U10495 ( .A(n10569), .B(n10570), .Z(n10332) );
  XOR2_X1 U10496 ( .A(n10571), .B(n10572), .Z(n10570) );
  XOR2_X1 U10497 ( .A(n10573), .B(n10574), .Z(n10336) );
  XOR2_X1 U10498 ( .A(n10575), .B(n10576), .Z(n10574) );
  XOR2_X1 U10499 ( .A(n10577), .B(n10578), .Z(n10340) );
  XOR2_X1 U10500 ( .A(n10579), .B(n10580), .Z(n10578) );
  XOR2_X1 U10501 ( .A(n10581), .B(n10582), .Z(n10344) );
  XOR2_X1 U10502 ( .A(n10583), .B(n10584), .Z(n10582) );
  XOR2_X1 U10503 ( .A(n10585), .B(n10586), .Z(n10348) );
  XOR2_X1 U10504 ( .A(n10587), .B(n10588), .Z(n10586) );
  XOR2_X1 U10505 ( .A(n10589), .B(n10590), .Z(n10352) );
  XOR2_X1 U10506 ( .A(n10591), .B(n10592), .Z(n10590) );
  XOR2_X1 U10507 ( .A(n10593), .B(n10594), .Z(n10356) );
  XOR2_X1 U10508 ( .A(n10595), .B(n10596), .Z(n10594) );
  XOR2_X1 U10509 ( .A(n10597), .B(n10598), .Z(n10360) );
  XOR2_X1 U10510 ( .A(n10599), .B(n10600), .Z(n10598) );
  XOR2_X1 U10511 ( .A(n10601), .B(n10602), .Z(n10364) );
  XOR2_X1 U10512 ( .A(n10603), .B(n10604), .Z(n10602) );
  XOR2_X1 U10513 ( .A(n10605), .B(n10606), .Z(n10368) );
  XOR2_X1 U10514 ( .A(n10607), .B(n10608), .Z(n10606) );
  XOR2_X1 U10515 ( .A(n10609), .B(n10610), .Z(n10372) );
  XOR2_X1 U10516 ( .A(n10611), .B(n10612), .Z(n10610) );
  XOR2_X1 U10517 ( .A(n10613), .B(n10614), .Z(n10376) );
  XOR2_X1 U10518 ( .A(n10615), .B(n10616), .Z(n10614) );
  XOR2_X1 U10519 ( .A(n10617), .B(n10618), .Z(n10380) );
  XOR2_X1 U10520 ( .A(n10619), .B(n10620), .Z(n10618) );
  OR2_X1 U10521 ( .A1(n10384), .A2(n10387), .ZN(n10427) );
  OR2_X1 U10522 ( .A1(n7730), .A2(n10057), .ZN(n10387) );
  XOR2_X1 U10523 ( .A(n10621), .B(n10622), .Z(n10384) );
  XOR2_X1 U10524 ( .A(n10623), .B(n10624), .Z(n10622) );
  OR2_X1 U10525 ( .A1(n10388), .A2(n10391), .ZN(n10424) );
  OR2_X1 U10526 ( .A1(n7697), .A2(n10057), .ZN(n10391) );
  XOR2_X1 U10527 ( .A(n10625), .B(n10626), .Z(n10388) );
  XOR2_X1 U10528 ( .A(n10627), .B(n10628), .Z(n10626) );
  OR2_X1 U10529 ( .A1(n10392), .A2(n10395), .ZN(n10421) );
  OR2_X1 U10530 ( .A1(n7660), .A2(n10057), .ZN(n10395) );
  XOR2_X1 U10531 ( .A(n10629), .B(n10630), .Z(n10392) );
  XOR2_X1 U10532 ( .A(n10631), .B(n10632), .Z(n10630) );
  XNOR2_X1 U10533 ( .A(n10402), .B(n10633), .ZN(n10176) );
  XOR2_X1 U10534 ( .A(n10405), .B(n10403), .Z(n10633) );
  OR2_X1 U10535 ( .A1(n7660), .A2(n10273), .ZN(n10403) );
  OR2_X1 U10536 ( .A1(n10634), .A2(n10635), .ZN(n10405) );
  AND2_X1 U10537 ( .A1(n10629), .A2(n10632), .ZN(n10635) );
  AND2_X1 U10538 ( .A1(n10636), .A2(n10631), .ZN(n10634) );
  OR2_X1 U10539 ( .A1(n10637), .A2(n10638), .ZN(n10631) );
  AND2_X1 U10540 ( .A1(n10625), .A2(n10628), .ZN(n10638) );
  AND2_X1 U10541 ( .A1(n10639), .A2(n10627), .ZN(n10637) );
  OR2_X1 U10542 ( .A1(n10640), .A2(n10641), .ZN(n10627) );
  AND2_X1 U10543 ( .A1(n10621), .A2(n10624), .ZN(n10641) );
  AND2_X1 U10544 ( .A1(n10642), .A2(n10623), .ZN(n10640) );
  OR2_X1 U10545 ( .A1(n10643), .A2(n10644), .ZN(n10623) );
  AND2_X1 U10546 ( .A1(n10617), .A2(n10620), .ZN(n10644) );
  AND2_X1 U10547 ( .A1(n10645), .A2(n10619), .ZN(n10643) );
  OR2_X1 U10548 ( .A1(n10646), .A2(n10647), .ZN(n10619) );
  AND2_X1 U10549 ( .A1(n10616), .A2(n10615), .ZN(n10647) );
  AND2_X1 U10550 ( .A1(n10613), .A2(n10648), .ZN(n10646) );
  OR2_X1 U10551 ( .A1(n10616), .A2(n10615), .ZN(n10648) );
  OR2_X1 U10552 ( .A1(n10649), .A2(n10650), .ZN(n10615) );
  AND2_X1 U10553 ( .A1(n10612), .A2(n10611), .ZN(n10650) );
  AND2_X1 U10554 ( .A1(n10609), .A2(n10651), .ZN(n10649) );
  OR2_X1 U10555 ( .A1(n10612), .A2(n10611), .ZN(n10651) );
  OR2_X1 U10556 ( .A1(n10652), .A2(n10653), .ZN(n10611) );
  AND2_X1 U10557 ( .A1(n10608), .A2(n10607), .ZN(n10653) );
  AND2_X1 U10558 ( .A1(n10605), .A2(n10654), .ZN(n10652) );
  OR2_X1 U10559 ( .A1(n10608), .A2(n10607), .ZN(n10654) );
  OR2_X1 U10560 ( .A1(n10655), .A2(n10656), .ZN(n10607) );
  AND2_X1 U10561 ( .A1(n10604), .A2(n10603), .ZN(n10656) );
  AND2_X1 U10562 ( .A1(n10601), .A2(n10657), .ZN(n10655) );
  OR2_X1 U10563 ( .A1(n10604), .A2(n10603), .ZN(n10657) );
  OR2_X1 U10564 ( .A1(n10658), .A2(n10659), .ZN(n10603) );
  AND2_X1 U10565 ( .A1(n10600), .A2(n10599), .ZN(n10659) );
  AND2_X1 U10566 ( .A1(n10597), .A2(n10660), .ZN(n10658) );
  OR2_X1 U10567 ( .A1(n10600), .A2(n10599), .ZN(n10660) );
  OR2_X1 U10568 ( .A1(n10661), .A2(n10662), .ZN(n10599) );
  AND2_X1 U10569 ( .A1(n10596), .A2(n10595), .ZN(n10662) );
  AND2_X1 U10570 ( .A1(n10593), .A2(n10663), .ZN(n10661) );
  OR2_X1 U10571 ( .A1(n10596), .A2(n10595), .ZN(n10663) );
  OR2_X1 U10572 ( .A1(n10664), .A2(n10665), .ZN(n10595) );
  AND2_X1 U10573 ( .A1(n10592), .A2(n10591), .ZN(n10665) );
  AND2_X1 U10574 ( .A1(n10589), .A2(n10666), .ZN(n10664) );
  OR2_X1 U10575 ( .A1(n10592), .A2(n10591), .ZN(n10666) );
  OR2_X1 U10576 ( .A1(n10667), .A2(n10668), .ZN(n10591) );
  AND2_X1 U10577 ( .A1(n10588), .A2(n10587), .ZN(n10668) );
  AND2_X1 U10578 ( .A1(n10585), .A2(n10669), .ZN(n10667) );
  OR2_X1 U10579 ( .A1(n10588), .A2(n10587), .ZN(n10669) );
  OR2_X1 U10580 ( .A1(n10670), .A2(n10671), .ZN(n10587) );
  AND2_X1 U10581 ( .A1(n10584), .A2(n10583), .ZN(n10671) );
  AND2_X1 U10582 ( .A1(n10581), .A2(n10672), .ZN(n10670) );
  OR2_X1 U10583 ( .A1(n10584), .A2(n10583), .ZN(n10672) );
  OR2_X1 U10584 ( .A1(n10673), .A2(n10674), .ZN(n10583) );
  AND2_X1 U10585 ( .A1(n10580), .A2(n10579), .ZN(n10674) );
  AND2_X1 U10586 ( .A1(n10577), .A2(n10675), .ZN(n10673) );
  OR2_X1 U10587 ( .A1(n10580), .A2(n10579), .ZN(n10675) );
  OR2_X1 U10588 ( .A1(n10676), .A2(n10677), .ZN(n10579) );
  AND2_X1 U10589 ( .A1(n10576), .A2(n10575), .ZN(n10677) );
  AND2_X1 U10590 ( .A1(n10573), .A2(n10678), .ZN(n10676) );
  OR2_X1 U10591 ( .A1(n10576), .A2(n10575), .ZN(n10678) );
  OR2_X1 U10592 ( .A1(n10679), .A2(n10680), .ZN(n10575) );
  AND2_X1 U10593 ( .A1(n10572), .A2(n10571), .ZN(n10680) );
  AND2_X1 U10594 ( .A1(n10569), .A2(n10681), .ZN(n10679) );
  OR2_X1 U10595 ( .A1(n10572), .A2(n10571), .ZN(n10681) );
  OR2_X1 U10596 ( .A1(n10682), .A2(n10683), .ZN(n10571) );
  AND2_X1 U10597 ( .A1(n10568), .A2(n10567), .ZN(n10683) );
  AND2_X1 U10598 ( .A1(n10565), .A2(n10684), .ZN(n10682) );
  OR2_X1 U10599 ( .A1(n10568), .A2(n10567), .ZN(n10684) );
  OR2_X1 U10600 ( .A1(n10685), .A2(n10686), .ZN(n10567) );
  AND2_X1 U10601 ( .A1(n10564), .A2(n10563), .ZN(n10686) );
  AND2_X1 U10602 ( .A1(n10561), .A2(n10687), .ZN(n10685) );
  OR2_X1 U10603 ( .A1(n10564), .A2(n10563), .ZN(n10687) );
  OR2_X1 U10604 ( .A1(n10688), .A2(n10689), .ZN(n10563) );
  AND2_X1 U10605 ( .A1(n10560), .A2(n10559), .ZN(n10689) );
  AND2_X1 U10606 ( .A1(n10557), .A2(n10690), .ZN(n10688) );
  OR2_X1 U10607 ( .A1(n10560), .A2(n10559), .ZN(n10690) );
  OR2_X1 U10608 ( .A1(n10691), .A2(n10692), .ZN(n10559) );
  AND2_X1 U10609 ( .A1(n10556), .A2(n10555), .ZN(n10692) );
  AND2_X1 U10610 ( .A1(n10553), .A2(n10693), .ZN(n10691) );
  OR2_X1 U10611 ( .A1(n10556), .A2(n10555), .ZN(n10693) );
  OR2_X1 U10612 ( .A1(n10694), .A2(n10695), .ZN(n10555) );
  AND2_X1 U10613 ( .A1(n10550), .A2(n10552), .ZN(n10695) );
  AND2_X1 U10614 ( .A1(n10696), .A2(n10551), .ZN(n10694) );
  OR2_X1 U10615 ( .A1(n10550), .A2(n10552), .ZN(n10696) );
  OR2_X1 U10616 ( .A1(n10697), .A2(n10698), .ZN(n10552) );
  AND2_X1 U10617 ( .A1(n10548), .A2(n10547), .ZN(n10698) );
  AND2_X1 U10618 ( .A1(n10545), .A2(n10699), .ZN(n10697) );
  OR2_X1 U10619 ( .A1(n10548), .A2(n10547), .ZN(n10699) );
  OR2_X1 U10620 ( .A1(n10700), .A2(n10701), .ZN(n10547) );
  AND2_X1 U10621 ( .A1(n10491), .A2(n10490), .ZN(n10701) );
  AND2_X1 U10622 ( .A1(n10488), .A2(n10702), .ZN(n10700) );
  OR2_X1 U10623 ( .A1(n10491), .A2(n10490), .ZN(n10702) );
  OR2_X1 U10624 ( .A1(n10703), .A2(n10704), .ZN(n10490) );
  AND2_X1 U10625 ( .A1(n10544), .A2(n10543), .ZN(n10704) );
  AND2_X1 U10626 ( .A1(n10541), .A2(n10705), .ZN(n10703) );
  OR2_X1 U10627 ( .A1(n10544), .A2(n10543), .ZN(n10705) );
  OR2_X1 U10628 ( .A1(n10706), .A2(n10707), .ZN(n10543) );
  AND2_X1 U10629 ( .A1(n10540), .A2(n10539), .ZN(n10707) );
  AND2_X1 U10630 ( .A1(n10537), .A2(n10708), .ZN(n10706) );
  OR2_X1 U10631 ( .A1(n10540), .A2(n10539), .ZN(n10708) );
  OR2_X1 U10632 ( .A1(n10709), .A2(n10710), .ZN(n10539) );
  AND2_X1 U10633 ( .A1(n10536), .A2(n10535), .ZN(n10710) );
  AND2_X1 U10634 ( .A1(n10533), .A2(n10711), .ZN(n10709) );
  OR2_X1 U10635 ( .A1(n10536), .A2(n10535), .ZN(n10711) );
  OR2_X1 U10636 ( .A1(n10712), .A2(n10713), .ZN(n10535) );
  AND2_X1 U10637 ( .A1(n10532), .A2(n10531), .ZN(n10713) );
  AND2_X1 U10638 ( .A1(n10529), .A2(n10714), .ZN(n10712) );
  OR2_X1 U10639 ( .A1(n10532), .A2(n10531), .ZN(n10714) );
  OR2_X1 U10640 ( .A1(n10715), .A2(n10716), .ZN(n10531) );
  AND2_X1 U10641 ( .A1(n10528), .A2(n10527), .ZN(n10716) );
  AND2_X1 U10642 ( .A1(n10525), .A2(n10717), .ZN(n10715) );
  OR2_X1 U10643 ( .A1(n10528), .A2(n10527), .ZN(n10717) );
  OR2_X1 U10644 ( .A1(n10718), .A2(n10719), .ZN(n10527) );
  AND2_X1 U10645 ( .A1(n10522), .A2(n10523), .ZN(n10719) );
  AND2_X1 U10646 ( .A1(n10720), .A2(n10721), .ZN(n10718) );
  OR2_X1 U10647 ( .A1(n10522), .A2(n10523), .ZN(n10721) );
  OR2_X1 U10648 ( .A1(n10273), .A2(n10722), .ZN(n10523) );
  OR2_X1 U10649 ( .A1(n8956), .A2(n10407), .ZN(n10722) );
  OR2_X1 U10650 ( .A1(n8515), .A2(n10273), .ZN(n10522) );
  INV_X1 U10651 ( .A(n10524), .ZN(n10720) );
  OR2_X1 U10652 ( .A1(n10723), .A2(n10724), .ZN(n10524) );
  AND2_X1 U10653 ( .A1(b_20_), .A2(n10725), .ZN(n10724) );
  OR2_X1 U10654 ( .A1(n10726), .A2(n7343), .ZN(n10725) );
  AND2_X1 U10655 ( .A1(a_30_), .A2(n10727), .ZN(n10726) );
  AND2_X1 U10656 ( .A1(b_19_), .A2(n10728), .ZN(n10723) );
  OR2_X1 U10657 ( .A1(n10729), .A2(n7347), .ZN(n10728) );
  AND2_X1 U10658 ( .A1(a_31_), .A2(n10407), .ZN(n10729) );
  OR2_X1 U10659 ( .A1(n8523), .A2(n10273), .ZN(n10528) );
  XOR2_X1 U10660 ( .A(n10730), .B(n10731), .Z(n10525) );
  XNOR2_X1 U10661 ( .A(n10732), .B(n10733), .ZN(n10730) );
  OR2_X1 U10662 ( .A1(n8528), .A2(n10273), .ZN(n10532) );
  XOR2_X1 U10663 ( .A(n10734), .B(n10735), .Z(n10529) );
  XOR2_X1 U10664 ( .A(n10736), .B(n10737), .Z(n10735) );
  OR2_X1 U10665 ( .A1(n8533), .A2(n10273), .ZN(n10536) );
  XOR2_X1 U10666 ( .A(n10738), .B(n10739), .Z(n10533) );
  XOR2_X1 U10667 ( .A(n10740), .B(n10741), .Z(n10739) );
  OR2_X1 U10668 ( .A1(n8538), .A2(n10273), .ZN(n10540) );
  XOR2_X1 U10669 ( .A(n10742), .B(n10743), .Z(n10537) );
  XOR2_X1 U10670 ( .A(n10744), .B(n10745), .Z(n10743) );
  OR2_X1 U10671 ( .A1(n8543), .A2(n10273), .ZN(n10544) );
  XOR2_X1 U10672 ( .A(n10746), .B(n10747), .Z(n10541) );
  XOR2_X1 U10673 ( .A(n10748), .B(n10749), .Z(n10747) );
  OR2_X1 U10674 ( .A1(n8548), .A2(n10273), .ZN(n10491) );
  XOR2_X1 U10675 ( .A(n10750), .B(n10751), .Z(n10488) );
  XOR2_X1 U10676 ( .A(n10752), .B(n10753), .Z(n10751) );
  OR2_X1 U10677 ( .A1(n8553), .A2(n10273), .ZN(n10548) );
  XOR2_X1 U10678 ( .A(n10754), .B(n10755), .Z(n10545) );
  XOR2_X1 U10679 ( .A(n10756), .B(n10757), .Z(n10755) );
  XOR2_X1 U10680 ( .A(n10758), .B(n10759), .Z(n10550) );
  XOR2_X1 U10681 ( .A(n10760), .B(n10761), .Z(n10759) );
  OR2_X1 U10682 ( .A1(n8563), .A2(n10273), .ZN(n10556) );
  XOR2_X1 U10683 ( .A(n10762), .B(n10763), .Z(n10553) );
  XOR2_X1 U10684 ( .A(n10764), .B(n10765), .Z(n10763) );
  OR2_X1 U10685 ( .A1(n8568), .A2(n10273), .ZN(n10560) );
  XNOR2_X1 U10686 ( .A(n10766), .B(n10767), .ZN(n10557) );
  XNOR2_X1 U10687 ( .A(n10768), .B(n10769), .ZN(n10766) );
  OR2_X1 U10688 ( .A1(n8573), .A2(n10273), .ZN(n10564) );
  XOR2_X1 U10689 ( .A(n10770), .B(n10771), .Z(n10561) );
  XOR2_X1 U10690 ( .A(n10772), .B(n10773), .Z(n10771) );
  OR2_X1 U10691 ( .A1(n8578), .A2(n10273), .ZN(n10568) );
  XOR2_X1 U10692 ( .A(n10774), .B(n10775), .Z(n10565) );
  XOR2_X1 U10693 ( .A(n10776), .B(n10777), .Z(n10775) );
  OR2_X1 U10694 ( .A1(n8583), .A2(n10273), .ZN(n10572) );
  XOR2_X1 U10695 ( .A(n10778), .B(n10779), .Z(n10569) );
  XOR2_X1 U10696 ( .A(n10780), .B(n10781), .Z(n10779) );
  OR2_X1 U10697 ( .A1(n8588), .A2(n10273), .ZN(n10576) );
  XOR2_X1 U10698 ( .A(n10782), .B(n10783), .Z(n10573) );
  XOR2_X1 U10699 ( .A(n10784), .B(n10785), .Z(n10783) );
  OR2_X1 U10700 ( .A1(n8593), .A2(n10273), .ZN(n10580) );
  XOR2_X1 U10701 ( .A(n10786), .B(n10787), .Z(n10577) );
  XOR2_X1 U10702 ( .A(n10788), .B(n10789), .Z(n10787) );
  OR2_X1 U10703 ( .A1(n8598), .A2(n10273), .ZN(n10584) );
  XOR2_X1 U10704 ( .A(n10790), .B(n10791), .Z(n10581) );
  XOR2_X1 U10705 ( .A(n10792), .B(n10793), .Z(n10791) );
  OR2_X1 U10706 ( .A1(n8603), .A2(n10273), .ZN(n10588) );
  XOR2_X1 U10707 ( .A(n10794), .B(n10795), .Z(n10585) );
  XOR2_X1 U10708 ( .A(n10796), .B(n10797), .Z(n10795) );
  OR2_X1 U10709 ( .A1(n8608), .A2(n10273), .ZN(n10592) );
  XOR2_X1 U10710 ( .A(n10798), .B(n10799), .Z(n10589) );
  XOR2_X1 U10711 ( .A(n10800), .B(n10801), .Z(n10799) );
  OR2_X1 U10712 ( .A1(n8287), .A2(n10273), .ZN(n10596) );
  XOR2_X1 U10713 ( .A(n10802), .B(n10803), .Z(n10593) );
  XOR2_X1 U10714 ( .A(n10804), .B(n10805), .Z(n10803) );
  OR2_X1 U10715 ( .A1(n8191), .A2(n10273), .ZN(n10600) );
  XOR2_X1 U10716 ( .A(n10806), .B(n10807), .Z(n10597) );
  XOR2_X1 U10717 ( .A(n10808), .B(n10809), .Z(n10807) );
  OR2_X1 U10718 ( .A1(n8107), .A2(n10273), .ZN(n10604) );
  XOR2_X1 U10719 ( .A(n10810), .B(n10811), .Z(n10601) );
  XOR2_X1 U10720 ( .A(n10812), .B(n10813), .Z(n10811) );
  OR2_X1 U10721 ( .A1(n8025), .A2(n10273), .ZN(n10608) );
  XOR2_X1 U10722 ( .A(n10814), .B(n10815), .Z(n10605) );
  XOR2_X1 U10723 ( .A(n10816), .B(n10817), .Z(n10815) );
  OR2_X1 U10724 ( .A1(n7955), .A2(n10273), .ZN(n10612) );
  XOR2_X1 U10725 ( .A(n10818), .B(n10819), .Z(n10609) );
  XOR2_X1 U10726 ( .A(n10820), .B(n10821), .Z(n10819) );
  OR2_X1 U10727 ( .A1(n7887), .A2(n10273), .ZN(n10616) );
  XOR2_X1 U10728 ( .A(n10822), .B(n10823), .Z(n10613) );
  XOR2_X1 U10729 ( .A(n10824), .B(n10825), .Z(n10823) );
  OR2_X1 U10730 ( .A1(n10617), .A2(n10620), .ZN(n10645) );
  OR2_X1 U10731 ( .A1(n7828), .A2(n10273), .ZN(n10620) );
  XOR2_X1 U10732 ( .A(n10826), .B(n10827), .Z(n10617) );
  XOR2_X1 U10733 ( .A(n10828), .B(n10829), .Z(n10827) );
  OR2_X1 U10734 ( .A1(n10621), .A2(n10624), .ZN(n10642) );
  OR2_X1 U10735 ( .A1(n7820), .A2(n10273), .ZN(n10624) );
  XOR2_X1 U10736 ( .A(n10830), .B(n10831), .Z(n10621) );
  XOR2_X1 U10737 ( .A(n10832), .B(n10833), .Z(n10831) );
  OR2_X1 U10738 ( .A1(n10625), .A2(n10628), .ZN(n10639) );
  OR2_X1 U10739 ( .A1(n7730), .A2(n10273), .ZN(n10628) );
  XOR2_X1 U10740 ( .A(n10834), .B(n10835), .Z(n10625) );
  XOR2_X1 U10741 ( .A(n10836), .B(n10837), .Z(n10835) );
  OR2_X1 U10742 ( .A1(n10629), .A2(n10632), .ZN(n10636) );
  OR2_X1 U10743 ( .A1(n7697), .A2(n10273), .ZN(n10632) );
  XOR2_X1 U10744 ( .A(n10838), .B(n10839), .Z(n10629) );
  XOR2_X1 U10745 ( .A(n10840), .B(n10841), .Z(n10839) );
  XOR2_X1 U10746 ( .A(n10410), .B(n10842), .Z(n10402) );
  XOR2_X1 U10747 ( .A(n10413), .B(n10411), .Z(n10842) );
  OR2_X1 U10748 ( .A1(n7697), .A2(n10407), .ZN(n10411) );
  OR2_X1 U10749 ( .A1(n10843), .A2(n10844), .ZN(n10413) );
  AND2_X1 U10750 ( .A1(n10838), .A2(n10841), .ZN(n10844) );
  AND2_X1 U10751 ( .A1(n10845), .A2(n10840), .ZN(n10843) );
  OR2_X1 U10752 ( .A1(n10846), .A2(n10847), .ZN(n10840) );
  AND2_X1 U10753 ( .A1(n10834), .A2(n10837), .ZN(n10847) );
  AND2_X1 U10754 ( .A1(n10848), .A2(n10836), .ZN(n10846) );
  OR2_X1 U10755 ( .A1(n10849), .A2(n10850), .ZN(n10836) );
  AND2_X1 U10756 ( .A1(n10830), .A2(n10833), .ZN(n10850) );
  AND2_X1 U10757 ( .A1(n10851), .A2(n10832), .ZN(n10849) );
  OR2_X1 U10758 ( .A1(n10852), .A2(n10853), .ZN(n10832) );
  AND2_X1 U10759 ( .A1(n10826), .A2(n10829), .ZN(n10853) );
  AND2_X1 U10760 ( .A1(n10854), .A2(n10828), .ZN(n10852) );
  OR2_X1 U10761 ( .A1(n10855), .A2(n10856), .ZN(n10828) );
  AND2_X1 U10762 ( .A1(n10822), .A2(n10825), .ZN(n10856) );
  AND2_X1 U10763 ( .A1(n10857), .A2(n10824), .ZN(n10855) );
  OR2_X1 U10764 ( .A1(n10858), .A2(n10859), .ZN(n10824) );
  AND2_X1 U10765 ( .A1(n10821), .A2(n10820), .ZN(n10859) );
  AND2_X1 U10766 ( .A1(n10818), .A2(n10860), .ZN(n10858) );
  OR2_X1 U10767 ( .A1(n10821), .A2(n10820), .ZN(n10860) );
  OR2_X1 U10768 ( .A1(n10861), .A2(n10862), .ZN(n10820) );
  AND2_X1 U10769 ( .A1(n10817), .A2(n10816), .ZN(n10862) );
  AND2_X1 U10770 ( .A1(n10814), .A2(n10863), .ZN(n10861) );
  OR2_X1 U10771 ( .A1(n10817), .A2(n10816), .ZN(n10863) );
  OR2_X1 U10772 ( .A1(n10864), .A2(n10865), .ZN(n10816) );
  AND2_X1 U10773 ( .A1(n10813), .A2(n10812), .ZN(n10865) );
  AND2_X1 U10774 ( .A1(n10810), .A2(n10866), .ZN(n10864) );
  OR2_X1 U10775 ( .A1(n10813), .A2(n10812), .ZN(n10866) );
  OR2_X1 U10776 ( .A1(n10867), .A2(n10868), .ZN(n10812) );
  AND2_X1 U10777 ( .A1(n10809), .A2(n10808), .ZN(n10868) );
  AND2_X1 U10778 ( .A1(n10806), .A2(n10869), .ZN(n10867) );
  OR2_X1 U10779 ( .A1(n10809), .A2(n10808), .ZN(n10869) );
  OR2_X1 U10780 ( .A1(n10870), .A2(n10871), .ZN(n10808) );
  AND2_X1 U10781 ( .A1(n10805), .A2(n10804), .ZN(n10871) );
  AND2_X1 U10782 ( .A1(n10802), .A2(n10872), .ZN(n10870) );
  OR2_X1 U10783 ( .A1(n10805), .A2(n10804), .ZN(n10872) );
  OR2_X1 U10784 ( .A1(n10873), .A2(n10874), .ZN(n10804) );
  AND2_X1 U10785 ( .A1(n10801), .A2(n10800), .ZN(n10874) );
  AND2_X1 U10786 ( .A1(n10798), .A2(n10875), .ZN(n10873) );
  OR2_X1 U10787 ( .A1(n10801), .A2(n10800), .ZN(n10875) );
  OR2_X1 U10788 ( .A1(n10876), .A2(n10877), .ZN(n10800) );
  AND2_X1 U10789 ( .A1(n10797), .A2(n10796), .ZN(n10877) );
  AND2_X1 U10790 ( .A1(n10794), .A2(n10878), .ZN(n10876) );
  OR2_X1 U10791 ( .A1(n10797), .A2(n10796), .ZN(n10878) );
  OR2_X1 U10792 ( .A1(n10879), .A2(n10880), .ZN(n10796) );
  AND2_X1 U10793 ( .A1(n10793), .A2(n10792), .ZN(n10880) );
  AND2_X1 U10794 ( .A1(n10790), .A2(n10881), .ZN(n10879) );
  OR2_X1 U10795 ( .A1(n10793), .A2(n10792), .ZN(n10881) );
  OR2_X1 U10796 ( .A1(n10882), .A2(n10883), .ZN(n10792) );
  AND2_X1 U10797 ( .A1(n10789), .A2(n10788), .ZN(n10883) );
  AND2_X1 U10798 ( .A1(n10786), .A2(n10884), .ZN(n10882) );
  OR2_X1 U10799 ( .A1(n10789), .A2(n10788), .ZN(n10884) );
  OR2_X1 U10800 ( .A1(n10885), .A2(n10886), .ZN(n10788) );
  AND2_X1 U10801 ( .A1(n10785), .A2(n10784), .ZN(n10886) );
  AND2_X1 U10802 ( .A1(n10782), .A2(n10887), .ZN(n10885) );
  OR2_X1 U10803 ( .A1(n10785), .A2(n10784), .ZN(n10887) );
  OR2_X1 U10804 ( .A1(n10888), .A2(n10889), .ZN(n10784) );
  AND2_X1 U10805 ( .A1(n10781), .A2(n10780), .ZN(n10889) );
  AND2_X1 U10806 ( .A1(n10778), .A2(n10890), .ZN(n10888) );
  OR2_X1 U10807 ( .A1(n10781), .A2(n10780), .ZN(n10890) );
  OR2_X1 U10808 ( .A1(n10891), .A2(n10892), .ZN(n10780) );
  AND2_X1 U10809 ( .A1(n10777), .A2(n10776), .ZN(n10892) );
  AND2_X1 U10810 ( .A1(n10774), .A2(n10893), .ZN(n10891) );
  OR2_X1 U10811 ( .A1(n10777), .A2(n10776), .ZN(n10893) );
  OR2_X1 U10812 ( .A1(n10894), .A2(n10895), .ZN(n10776) );
  AND2_X1 U10813 ( .A1(n10773), .A2(n10772), .ZN(n10895) );
  AND2_X1 U10814 ( .A1(n10770), .A2(n10896), .ZN(n10894) );
  OR2_X1 U10815 ( .A1(n10773), .A2(n10772), .ZN(n10896) );
  OR2_X1 U10816 ( .A1(n10897), .A2(n10898), .ZN(n10772) );
  AND2_X1 U10817 ( .A1(n10767), .A2(n10769), .ZN(n10898) );
  AND2_X1 U10818 ( .A1(n10899), .A2(n10768), .ZN(n10897) );
  OR2_X1 U10819 ( .A1(n10767), .A2(n10769), .ZN(n10899) );
  OR2_X1 U10820 ( .A1(n10900), .A2(n10901), .ZN(n10769) );
  AND2_X1 U10821 ( .A1(n10765), .A2(n10764), .ZN(n10901) );
  AND2_X1 U10822 ( .A1(n10762), .A2(n10902), .ZN(n10900) );
  OR2_X1 U10823 ( .A1(n10765), .A2(n10764), .ZN(n10902) );
  OR2_X1 U10824 ( .A1(n10903), .A2(n10904), .ZN(n10764) );
  AND2_X1 U10825 ( .A1(n10761), .A2(n10760), .ZN(n10904) );
  AND2_X1 U10826 ( .A1(n10758), .A2(n10905), .ZN(n10903) );
  OR2_X1 U10827 ( .A1(n10761), .A2(n10760), .ZN(n10905) );
  OR2_X1 U10828 ( .A1(n10906), .A2(n10907), .ZN(n10760) );
  AND2_X1 U10829 ( .A1(n10757), .A2(n10756), .ZN(n10907) );
  AND2_X1 U10830 ( .A1(n10754), .A2(n10908), .ZN(n10906) );
  OR2_X1 U10831 ( .A1(n10757), .A2(n10756), .ZN(n10908) );
  OR2_X1 U10832 ( .A1(n10909), .A2(n10910), .ZN(n10756) );
  AND2_X1 U10833 ( .A1(n10753), .A2(n10752), .ZN(n10910) );
  AND2_X1 U10834 ( .A1(n10750), .A2(n10911), .ZN(n10909) );
  OR2_X1 U10835 ( .A1(n10753), .A2(n10752), .ZN(n10911) );
  OR2_X1 U10836 ( .A1(n10912), .A2(n10913), .ZN(n10752) );
  AND2_X1 U10837 ( .A1(n10749), .A2(n10748), .ZN(n10913) );
  AND2_X1 U10838 ( .A1(n10746), .A2(n10914), .ZN(n10912) );
  OR2_X1 U10839 ( .A1(n10749), .A2(n10748), .ZN(n10914) );
  OR2_X1 U10840 ( .A1(n10915), .A2(n10916), .ZN(n10748) );
  AND2_X1 U10841 ( .A1(n10745), .A2(n10744), .ZN(n10916) );
  AND2_X1 U10842 ( .A1(n10742), .A2(n10917), .ZN(n10915) );
  OR2_X1 U10843 ( .A1(n10745), .A2(n10744), .ZN(n10917) );
  OR2_X1 U10844 ( .A1(n10918), .A2(n10919), .ZN(n10744) );
  AND2_X1 U10845 ( .A1(n10741), .A2(n10740), .ZN(n10919) );
  AND2_X1 U10846 ( .A1(n10738), .A2(n10920), .ZN(n10918) );
  OR2_X1 U10847 ( .A1(n10741), .A2(n10740), .ZN(n10920) );
  OR2_X1 U10848 ( .A1(n10921), .A2(n10922), .ZN(n10740) );
  AND2_X1 U10849 ( .A1(n10737), .A2(n10736), .ZN(n10922) );
  AND2_X1 U10850 ( .A1(n10734), .A2(n10923), .ZN(n10921) );
  OR2_X1 U10851 ( .A1(n10737), .A2(n10736), .ZN(n10923) );
  OR2_X1 U10852 ( .A1(n10924), .A2(n10925), .ZN(n10736) );
  AND2_X1 U10853 ( .A1(n10731), .A2(n10732), .ZN(n10925) );
  AND2_X1 U10854 ( .A1(n10926), .A2(n10927), .ZN(n10924) );
  OR2_X1 U10855 ( .A1(n10731), .A2(n10732), .ZN(n10927) );
  OR2_X1 U10856 ( .A1(n10407), .A2(n10928), .ZN(n10732) );
  OR2_X1 U10857 ( .A1(n8515), .A2(n10407), .ZN(n10731) );
  INV_X1 U10858 ( .A(n10733), .ZN(n10926) );
  OR2_X1 U10859 ( .A1(n10929), .A2(n10930), .ZN(n10733) );
  AND2_X1 U10860 ( .A1(b_19_), .A2(n10931), .ZN(n10930) );
  OR2_X1 U10861 ( .A1(n10932), .A2(n7343), .ZN(n10931) );
  AND2_X1 U10862 ( .A1(a_30_), .A2(n10933), .ZN(n10932) );
  AND2_X1 U10863 ( .A1(b_18_), .A2(n10934), .ZN(n10929) );
  OR2_X1 U10864 ( .A1(n10935), .A2(n7347), .ZN(n10934) );
  AND2_X1 U10865 ( .A1(a_31_), .A2(n10727), .ZN(n10935) );
  OR2_X1 U10866 ( .A1(n8523), .A2(n10407), .ZN(n10737) );
  XOR2_X1 U10867 ( .A(n10936), .B(n10937), .Z(n10734) );
  XNOR2_X1 U10868 ( .A(n10938), .B(n10939), .ZN(n10936) );
  OR2_X1 U10869 ( .A1(n8528), .A2(n10407), .ZN(n10741) );
  XOR2_X1 U10870 ( .A(n10940), .B(n10941), .Z(n10738) );
  XOR2_X1 U10871 ( .A(n10942), .B(n10943), .Z(n10941) );
  OR2_X1 U10872 ( .A1(n8533), .A2(n10407), .ZN(n10745) );
  XOR2_X1 U10873 ( .A(n10944), .B(n10945), .Z(n10742) );
  XOR2_X1 U10874 ( .A(n10946), .B(n10947), .Z(n10945) );
  OR2_X1 U10875 ( .A1(n8538), .A2(n10407), .ZN(n10749) );
  XOR2_X1 U10876 ( .A(n10948), .B(n10949), .Z(n10746) );
  XOR2_X1 U10877 ( .A(n10950), .B(n10951), .Z(n10949) );
  OR2_X1 U10878 ( .A1(n8543), .A2(n10407), .ZN(n10753) );
  XOR2_X1 U10879 ( .A(n10952), .B(n10953), .Z(n10750) );
  XOR2_X1 U10880 ( .A(n10954), .B(n10955), .Z(n10953) );
  OR2_X1 U10881 ( .A1(n8548), .A2(n10407), .ZN(n10757) );
  XOR2_X1 U10882 ( .A(n10956), .B(n10957), .Z(n10754) );
  XOR2_X1 U10883 ( .A(n10958), .B(n10959), .Z(n10957) );
  OR2_X1 U10884 ( .A1(n8553), .A2(n10407), .ZN(n10761) );
  XOR2_X1 U10885 ( .A(n10960), .B(n10961), .Z(n10758) );
  XOR2_X1 U10886 ( .A(n10962), .B(n10963), .Z(n10961) );
  OR2_X1 U10887 ( .A1(n8558), .A2(n10407), .ZN(n10765) );
  XOR2_X1 U10888 ( .A(n10964), .B(n10965), .Z(n10762) );
  XOR2_X1 U10889 ( .A(n10966), .B(n10967), .Z(n10965) );
  XOR2_X1 U10890 ( .A(n10968), .B(n10969), .Z(n10767) );
  XOR2_X1 U10891 ( .A(n10970), .B(n10971), .Z(n10969) );
  OR2_X1 U10892 ( .A1(n8568), .A2(n10407), .ZN(n10773) );
  XOR2_X1 U10893 ( .A(n10972), .B(n10973), .Z(n10770) );
  XOR2_X1 U10894 ( .A(n10974), .B(n10975), .Z(n10973) );
  OR2_X1 U10895 ( .A1(n8573), .A2(n10407), .ZN(n10777) );
  XNOR2_X1 U10896 ( .A(n10976), .B(n10977), .ZN(n10774) );
  XNOR2_X1 U10897 ( .A(n10978), .B(n10979), .ZN(n10976) );
  OR2_X1 U10898 ( .A1(n8578), .A2(n10407), .ZN(n10781) );
  XOR2_X1 U10899 ( .A(n10980), .B(n10981), .Z(n10778) );
  XOR2_X1 U10900 ( .A(n10982), .B(n10983), .Z(n10981) );
  OR2_X1 U10901 ( .A1(n8583), .A2(n10407), .ZN(n10785) );
  XOR2_X1 U10902 ( .A(n10984), .B(n10985), .Z(n10782) );
  XOR2_X1 U10903 ( .A(n10986), .B(n10987), .Z(n10985) );
  OR2_X1 U10904 ( .A1(n8588), .A2(n10407), .ZN(n10789) );
  XOR2_X1 U10905 ( .A(n10988), .B(n10989), .Z(n10786) );
  XOR2_X1 U10906 ( .A(n10990), .B(n10991), .Z(n10989) );
  OR2_X1 U10907 ( .A1(n8593), .A2(n10407), .ZN(n10793) );
  XOR2_X1 U10908 ( .A(n10992), .B(n10993), .Z(n10790) );
  XOR2_X1 U10909 ( .A(n10994), .B(n10995), .Z(n10993) );
  OR2_X1 U10910 ( .A1(n8598), .A2(n10407), .ZN(n10797) );
  XOR2_X1 U10911 ( .A(n10996), .B(n10997), .Z(n10794) );
  XOR2_X1 U10912 ( .A(n10998), .B(n10999), .Z(n10997) );
  OR2_X1 U10913 ( .A1(n8603), .A2(n10407), .ZN(n10801) );
  XOR2_X1 U10914 ( .A(n11000), .B(n11001), .Z(n10798) );
  XOR2_X1 U10915 ( .A(n11002), .B(n11003), .Z(n11001) );
  OR2_X1 U10916 ( .A1(n8608), .A2(n10407), .ZN(n10805) );
  XOR2_X1 U10917 ( .A(n11004), .B(n11005), .Z(n10802) );
  XOR2_X1 U10918 ( .A(n11006), .B(n11007), .Z(n11005) );
  OR2_X1 U10919 ( .A1(n8287), .A2(n10407), .ZN(n10809) );
  XOR2_X1 U10920 ( .A(n11008), .B(n11009), .Z(n10806) );
  XOR2_X1 U10921 ( .A(n11010), .B(n11011), .Z(n11009) );
  OR2_X1 U10922 ( .A1(n8191), .A2(n10407), .ZN(n10813) );
  XOR2_X1 U10923 ( .A(n11012), .B(n11013), .Z(n10810) );
  XOR2_X1 U10924 ( .A(n11014), .B(n11015), .Z(n11013) );
  OR2_X1 U10925 ( .A1(n8107), .A2(n10407), .ZN(n10817) );
  XOR2_X1 U10926 ( .A(n11016), .B(n11017), .Z(n10814) );
  XOR2_X1 U10927 ( .A(n11018), .B(n11019), .Z(n11017) );
  OR2_X1 U10928 ( .A1(n8025), .A2(n10407), .ZN(n10821) );
  XOR2_X1 U10929 ( .A(n11020), .B(n11021), .Z(n10818) );
  XOR2_X1 U10930 ( .A(n11022), .B(n11023), .Z(n11021) );
  OR2_X1 U10931 ( .A1(n10822), .A2(n10825), .ZN(n10857) );
  OR2_X1 U10932 ( .A1(n7955), .A2(n10407), .ZN(n10825) );
  XOR2_X1 U10933 ( .A(n11024), .B(n11025), .Z(n10822) );
  XOR2_X1 U10934 ( .A(n11026), .B(n11027), .Z(n11025) );
  OR2_X1 U10935 ( .A1(n10826), .A2(n10829), .ZN(n10854) );
  OR2_X1 U10936 ( .A1(n7887), .A2(n10407), .ZN(n10829) );
  XOR2_X1 U10937 ( .A(n11028), .B(n11029), .Z(n10826) );
  XOR2_X1 U10938 ( .A(n11030), .B(n11031), .Z(n11029) );
  OR2_X1 U10939 ( .A1(n10830), .A2(n10833), .ZN(n10851) );
  OR2_X1 U10940 ( .A1(n7828), .A2(n10407), .ZN(n10833) );
  XOR2_X1 U10941 ( .A(n11032), .B(n11033), .Z(n10830) );
  XOR2_X1 U10942 ( .A(n11034), .B(n11035), .Z(n11033) );
  OR2_X1 U10943 ( .A1(n10834), .A2(n10837), .ZN(n10848) );
  OR2_X1 U10944 ( .A1(n7820), .A2(n10407), .ZN(n10837) );
  XOR2_X1 U10945 ( .A(n11036), .B(n11037), .Z(n10834) );
  XOR2_X1 U10946 ( .A(n11038), .B(n11039), .Z(n11037) );
  OR2_X1 U10947 ( .A1(n10838), .A2(n10841), .ZN(n10845) );
  OR2_X1 U10948 ( .A1(n7730), .A2(n10407), .ZN(n10841) );
  XOR2_X1 U10949 ( .A(n11040), .B(n11041), .Z(n10838) );
  XOR2_X1 U10950 ( .A(n11042), .B(n11043), .Z(n11041) );
  XOR2_X1 U10951 ( .A(n11044), .B(n11045), .Z(n10410) );
  XOR2_X1 U10952 ( .A(n11046), .B(n11047), .Z(n11045) );
  AND2_X1 U10953 ( .A1(n8318), .A2(n7562), .ZN(n8316) );
  XNOR2_X1 U10954 ( .A(n8310), .B(n11048), .ZN(n7562) );
  INV_X1 U10955 ( .A(n7561), .ZN(n8318) );
  OR2_X1 U10956 ( .A1(n8322), .A2(n8323), .ZN(n7561) );
  OR2_X1 U10957 ( .A1(n11049), .A2(n11050), .ZN(n8323) );
  AND2_X1 U10958 ( .A1(n8339), .A2(n8342), .ZN(n11050) );
  AND2_X1 U10959 ( .A1(n11051), .A2(n8341), .ZN(n11049) );
  OR2_X1 U10960 ( .A1(n11052), .A2(n11053), .ZN(n8341) );
  AND2_X1 U10961 ( .A1(n10414), .A2(n10417), .ZN(n11053) );
  AND2_X1 U10962 ( .A1(n11054), .A2(n10416), .ZN(n11052) );
  OR2_X1 U10963 ( .A1(n11055), .A2(n11056), .ZN(n10416) );
  AND2_X1 U10964 ( .A1(n11044), .A2(n11047), .ZN(n11056) );
  AND2_X1 U10965 ( .A1(n11057), .A2(n11046), .ZN(n11055) );
  OR2_X1 U10966 ( .A1(n11058), .A2(n11059), .ZN(n11046) );
  AND2_X1 U10967 ( .A1(n11040), .A2(n11043), .ZN(n11059) );
  AND2_X1 U10968 ( .A1(n11060), .A2(n11042), .ZN(n11058) );
  OR2_X1 U10969 ( .A1(n11061), .A2(n11062), .ZN(n11042) );
  AND2_X1 U10970 ( .A1(n11036), .A2(n11039), .ZN(n11062) );
  AND2_X1 U10971 ( .A1(n11063), .A2(n11038), .ZN(n11061) );
  OR2_X1 U10972 ( .A1(n11064), .A2(n11065), .ZN(n11038) );
  AND2_X1 U10973 ( .A1(n11032), .A2(n11035), .ZN(n11065) );
  AND2_X1 U10974 ( .A1(n11066), .A2(n11034), .ZN(n11064) );
  OR2_X1 U10975 ( .A1(n11067), .A2(n11068), .ZN(n11034) );
  AND2_X1 U10976 ( .A1(n11028), .A2(n11031), .ZN(n11068) );
  AND2_X1 U10977 ( .A1(n11069), .A2(n11030), .ZN(n11067) );
  OR2_X1 U10978 ( .A1(n11070), .A2(n11071), .ZN(n11030) );
  AND2_X1 U10979 ( .A1(n11024), .A2(n11027), .ZN(n11071) );
  AND2_X1 U10980 ( .A1(n11072), .A2(n11026), .ZN(n11070) );
  OR2_X1 U10981 ( .A1(n11073), .A2(n11074), .ZN(n11026) );
  AND2_X1 U10982 ( .A1(n11020), .A2(n11023), .ZN(n11074) );
  AND2_X1 U10983 ( .A1(n11075), .A2(n11022), .ZN(n11073) );
  OR2_X1 U10984 ( .A1(n11076), .A2(n11077), .ZN(n11022) );
  AND2_X1 U10985 ( .A1(n11019), .A2(n11018), .ZN(n11077) );
  AND2_X1 U10986 ( .A1(n11016), .A2(n11078), .ZN(n11076) );
  OR2_X1 U10987 ( .A1(n11019), .A2(n11018), .ZN(n11078) );
  OR2_X1 U10988 ( .A1(n11079), .A2(n11080), .ZN(n11018) );
  AND2_X1 U10989 ( .A1(n11015), .A2(n11014), .ZN(n11080) );
  AND2_X1 U10990 ( .A1(n11012), .A2(n11081), .ZN(n11079) );
  OR2_X1 U10991 ( .A1(n11015), .A2(n11014), .ZN(n11081) );
  OR2_X1 U10992 ( .A1(n11082), .A2(n11083), .ZN(n11014) );
  AND2_X1 U10993 ( .A1(n11011), .A2(n11010), .ZN(n11083) );
  AND2_X1 U10994 ( .A1(n11008), .A2(n11084), .ZN(n11082) );
  OR2_X1 U10995 ( .A1(n11011), .A2(n11010), .ZN(n11084) );
  OR2_X1 U10996 ( .A1(n11085), .A2(n11086), .ZN(n11010) );
  AND2_X1 U10997 ( .A1(n11007), .A2(n11006), .ZN(n11086) );
  AND2_X1 U10998 ( .A1(n11004), .A2(n11087), .ZN(n11085) );
  OR2_X1 U10999 ( .A1(n11007), .A2(n11006), .ZN(n11087) );
  OR2_X1 U11000 ( .A1(n11088), .A2(n11089), .ZN(n11006) );
  AND2_X1 U11001 ( .A1(n11003), .A2(n11002), .ZN(n11089) );
  AND2_X1 U11002 ( .A1(n11000), .A2(n11090), .ZN(n11088) );
  OR2_X1 U11003 ( .A1(n11003), .A2(n11002), .ZN(n11090) );
  OR2_X1 U11004 ( .A1(n11091), .A2(n11092), .ZN(n11002) );
  AND2_X1 U11005 ( .A1(n10999), .A2(n10998), .ZN(n11092) );
  AND2_X1 U11006 ( .A1(n10996), .A2(n11093), .ZN(n11091) );
  OR2_X1 U11007 ( .A1(n10999), .A2(n10998), .ZN(n11093) );
  OR2_X1 U11008 ( .A1(n11094), .A2(n11095), .ZN(n10998) );
  AND2_X1 U11009 ( .A1(n10995), .A2(n10994), .ZN(n11095) );
  AND2_X1 U11010 ( .A1(n10992), .A2(n11096), .ZN(n11094) );
  OR2_X1 U11011 ( .A1(n10995), .A2(n10994), .ZN(n11096) );
  OR2_X1 U11012 ( .A1(n11097), .A2(n11098), .ZN(n10994) );
  AND2_X1 U11013 ( .A1(n10991), .A2(n10990), .ZN(n11098) );
  AND2_X1 U11014 ( .A1(n10988), .A2(n11099), .ZN(n11097) );
  OR2_X1 U11015 ( .A1(n10991), .A2(n10990), .ZN(n11099) );
  OR2_X1 U11016 ( .A1(n11100), .A2(n11101), .ZN(n10990) );
  AND2_X1 U11017 ( .A1(n10987), .A2(n10986), .ZN(n11101) );
  AND2_X1 U11018 ( .A1(n10984), .A2(n11102), .ZN(n11100) );
  OR2_X1 U11019 ( .A1(n10987), .A2(n10986), .ZN(n11102) );
  OR2_X1 U11020 ( .A1(n11103), .A2(n11104), .ZN(n10986) );
  AND2_X1 U11021 ( .A1(n10983), .A2(n10982), .ZN(n11104) );
  AND2_X1 U11022 ( .A1(n10980), .A2(n11105), .ZN(n11103) );
  OR2_X1 U11023 ( .A1(n10983), .A2(n10982), .ZN(n11105) );
  OR2_X1 U11024 ( .A1(n11106), .A2(n11107), .ZN(n10982) );
  AND2_X1 U11025 ( .A1(n10977), .A2(n10979), .ZN(n11107) );
  AND2_X1 U11026 ( .A1(n11108), .A2(n10978), .ZN(n11106) );
  OR2_X1 U11027 ( .A1(n10977), .A2(n10979), .ZN(n11108) );
  OR2_X1 U11028 ( .A1(n11109), .A2(n11110), .ZN(n10979) );
  AND2_X1 U11029 ( .A1(n10975), .A2(n10974), .ZN(n11110) );
  AND2_X1 U11030 ( .A1(n10972), .A2(n11111), .ZN(n11109) );
  OR2_X1 U11031 ( .A1(n10975), .A2(n10974), .ZN(n11111) );
  OR2_X1 U11032 ( .A1(n11112), .A2(n11113), .ZN(n10974) );
  AND2_X1 U11033 ( .A1(n10971), .A2(n10970), .ZN(n11113) );
  AND2_X1 U11034 ( .A1(n10968), .A2(n11114), .ZN(n11112) );
  OR2_X1 U11035 ( .A1(n10971), .A2(n10970), .ZN(n11114) );
  OR2_X1 U11036 ( .A1(n11115), .A2(n11116), .ZN(n10970) );
  AND2_X1 U11037 ( .A1(n10967), .A2(n10966), .ZN(n11116) );
  AND2_X1 U11038 ( .A1(n10964), .A2(n11117), .ZN(n11115) );
  OR2_X1 U11039 ( .A1(n10967), .A2(n10966), .ZN(n11117) );
  OR2_X1 U11040 ( .A1(n11118), .A2(n11119), .ZN(n10966) );
  AND2_X1 U11041 ( .A1(n10963), .A2(n10962), .ZN(n11119) );
  AND2_X1 U11042 ( .A1(n10960), .A2(n11120), .ZN(n11118) );
  OR2_X1 U11043 ( .A1(n10963), .A2(n10962), .ZN(n11120) );
  OR2_X1 U11044 ( .A1(n11121), .A2(n11122), .ZN(n10962) );
  AND2_X1 U11045 ( .A1(n10959), .A2(n10958), .ZN(n11122) );
  AND2_X1 U11046 ( .A1(n10956), .A2(n11123), .ZN(n11121) );
  OR2_X1 U11047 ( .A1(n10959), .A2(n10958), .ZN(n11123) );
  OR2_X1 U11048 ( .A1(n11124), .A2(n11125), .ZN(n10958) );
  AND2_X1 U11049 ( .A1(n10955), .A2(n10954), .ZN(n11125) );
  AND2_X1 U11050 ( .A1(n10952), .A2(n11126), .ZN(n11124) );
  OR2_X1 U11051 ( .A1(n10955), .A2(n10954), .ZN(n11126) );
  OR2_X1 U11052 ( .A1(n11127), .A2(n11128), .ZN(n10954) );
  AND2_X1 U11053 ( .A1(n10951), .A2(n10950), .ZN(n11128) );
  AND2_X1 U11054 ( .A1(n10948), .A2(n11129), .ZN(n11127) );
  OR2_X1 U11055 ( .A1(n10951), .A2(n10950), .ZN(n11129) );
  OR2_X1 U11056 ( .A1(n11130), .A2(n11131), .ZN(n10950) );
  AND2_X1 U11057 ( .A1(n10947), .A2(n10946), .ZN(n11131) );
  AND2_X1 U11058 ( .A1(n10944), .A2(n11132), .ZN(n11130) );
  OR2_X1 U11059 ( .A1(n10947), .A2(n10946), .ZN(n11132) );
  OR2_X1 U11060 ( .A1(n11133), .A2(n11134), .ZN(n10946) );
  AND2_X1 U11061 ( .A1(n10943), .A2(n10942), .ZN(n11134) );
  AND2_X1 U11062 ( .A1(n10940), .A2(n11135), .ZN(n11133) );
  OR2_X1 U11063 ( .A1(n10943), .A2(n10942), .ZN(n11135) );
  OR2_X1 U11064 ( .A1(n11136), .A2(n11137), .ZN(n10942) );
  AND2_X1 U11065 ( .A1(n10937), .A2(n10938), .ZN(n11137) );
  AND2_X1 U11066 ( .A1(n11138), .A2(n11139), .ZN(n11136) );
  OR2_X1 U11067 ( .A1(n10937), .A2(n10938), .ZN(n11139) );
  OR2_X1 U11068 ( .A1(n10933), .A2(n10928), .ZN(n10938) );
  OR2_X1 U11069 ( .A1(n8956), .A2(n10727), .ZN(n10928) );
  OR2_X1 U11070 ( .A1(n8515), .A2(n10727), .ZN(n10937) );
  INV_X1 U11071 ( .A(n10939), .ZN(n11138) );
  OR2_X1 U11072 ( .A1(n11140), .A2(n11141), .ZN(n10939) );
  AND2_X1 U11073 ( .A1(b_18_), .A2(n11142), .ZN(n11141) );
  OR2_X1 U11074 ( .A1(n11143), .A2(n7343), .ZN(n11142) );
  AND2_X1 U11075 ( .A1(a_30_), .A2(n11144), .ZN(n11143) );
  AND2_X1 U11076 ( .A1(b_17_), .A2(n11145), .ZN(n11140) );
  OR2_X1 U11077 ( .A1(n11146), .A2(n7347), .ZN(n11145) );
  AND2_X1 U11078 ( .A1(a_31_), .A2(n10933), .ZN(n11146) );
  OR2_X1 U11079 ( .A1(n8523), .A2(n10727), .ZN(n10943) );
  XOR2_X1 U11080 ( .A(n11147), .B(n11148), .Z(n10940) );
  XNOR2_X1 U11081 ( .A(n11149), .B(n11150), .ZN(n11147) );
  OR2_X1 U11082 ( .A1(n8528), .A2(n10727), .ZN(n10947) );
  XOR2_X1 U11083 ( .A(n11151), .B(n11152), .Z(n10944) );
  XOR2_X1 U11084 ( .A(n11153), .B(n11154), .Z(n11152) );
  OR2_X1 U11085 ( .A1(n8533), .A2(n10727), .ZN(n10951) );
  XOR2_X1 U11086 ( .A(n11155), .B(n11156), .Z(n10948) );
  XOR2_X1 U11087 ( .A(n11157), .B(n11158), .Z(n11156) );
  OR2_X1 U11088 ( .A1(n8538), .A2(n10727), .ZN(n10955) );
  XOR2_X1 U11089 ( .A(n11159), .B(n11160), .Z(n10952) );
  XOR2_X1 U11090 ( .A(n11161), .B(n11162), .Z(n11160) );
  OR2_X1 U11091 ( .A1(n8543), .A2(n10727), .ZN(n10959) );
  XOR2_X1 U11092 ( .A(n11163), .B(n11164), .Z(n10956) );
  XOR2_X1 U11093 ( .A(n11165), .B(n11166), .Z(n11164) );
  OR2_X1 U11094 ( .A1(n8548), .A2(n10727), .ZN(n10963) );
  XOR2_X1 U11095 ( .A(n11167), .B(n11168), .Z(n10960) );
  XOR2_X1 U11096 ( .A(n11169), .B(n11170), .Z(n11168) );
  OR2_X1 U11097 ( .A1(n8553), .A2(n10727), .ZN(n10967) );
  XOR2_X1 U11098 ( .A(n11171), .B(n11172), .Z(n10964) );
  XOR2_X1 U11099 ( .A(n11173), .B(n11174), .Z(n11172) );
  OR2_X1 U11100 ( .A1(n8558), .A2(n10727), .ZN(n10971) );
  XOR2_X1 U11101 ( .A(n11175), .B(n11176), .Z(n10968) );
  XOR2_X1 U11102 ( .A(n11177), .B(n11178), .Z(n11176) );
  OR2_X1 U11103 ( .A1(n8563), .A2(n10727), .ZN(n10975) );
  XOR2_X1 U11104 ( .A(n11179), .B(n11180), .Z(n10972) );
  XOR2_X1 U11105 ( .A(n11181), .B(n11182), .Z(n11180) );
  XOR2_X1 U11106 ( .A(n11183), .B(n11184), .Z(n10977) );
  XOR2_X1 U11107 ( .A(n11185), .B(n11186), .Z(n11184) );
  OR2_X1 U11108 ( .A1(n8573), .A2(n10727), .ZN(n10983) );
  XOR2_X1 U11109 ( .A(n11187), .B(n11188), .Z(n10980) );
  XOR2_X1 U11110 ( .A(n11189), .B(n11190), .Z(n11188) );
  OR2_X1 U11111 ( .A1(n8578), .A2(n10727), .ZN(n10987) );
  XNOR2_X1 U11112 ( .A(n11191), .B(n11192), .ZN(n10984) );
  XNOR2_X1 U11113 ( .A(n11193), .B(n11194), .ZN(n11191) );
  OR2_X1 U11114 ( .A1(n8583), .A2(n10727), .ZN(n10991) );
  XOR2_X1 U11115 ( .A(n11195), .B(n11196), .Z(n10988) );
  XOR2_X1 U11116 ( .A(n11197), .B(n11198), .Z(n11196) );
  OR2_X1 U11117 ( .A1(n8588), .A2(n10727), .ZN(n10995) );
  XOR2_X1 U11118 ( .A(n11199), .B(n11200), .Z(n10992) );
  XOR2_X1 U11119 ( .A(n11201), .B(n11202), .Z(n11200) );
  OR2_X1 U11120 ( .A1(n8593), .A2(n10727), .ZN(n10999) );
  XOR2_X1 U11121 ( .A(n11203), .B(n11204), .Z(n10996) );
  XOR2_X1 U11122 ( .A(n11205), .B(n11206), .Z(n11204) );
  OR2_X1 U11123 ( .A1(n8598), .A2(n10727), .ZN(n11003) );
  XOR2_X1 U11124 ( .A(n11207), .B(n11208), .Z(n11000) );
  XOR2_X1 U11125 ( .A(n11209), .B(n11210), .Z(n11208) );
  OR2_X1 U11126 ( .A1(n8603), .A2(n10727), .ZN(n11007) );
  XOR2_X1 U11127 ( .A(n11211), .B(n11212), .Z(n11004) );
  XOR2_X1 U11128 ( .A(n11213), .B(n11214), .Z(n11212) );
  OR2_X1 U11129 ( .A1(n8608), .A2(n10727), .ZN(n11011) );
  XOR2_X1 U11130 ( .A(n11215), .B(n11216), .Z(n11008) );
  XOR2_X1 U11131 ( .A(n11217), .B(n11218), .Z(n11216) );
  OR2_X1 U11132 ( .A1(n8287), .A2(n10727), .ZN(n11015) );
  XOR2_X1 U11133 ( .A(n11219), .B(n11220), .Z(n11012) );
  XOR2_X1 U11134 ( .A(n11221), .B(n11222), .Z(n11220) );
  OR2_X1 U11135 ( .A1(n8191), .A2(n10727), .ZN(n11019) );
  XOR2_X1 U11136 ( .A(n11223), .B(n11224), .Z(n11016) );
  XOR2_X1 U11137 ( .A(n11225), .B(n11226), .Z(n11224) );
  OR2_X1 U11138 ( .A1(n11020), .A2(n11023), .ZN(n11075) );
  OR2_X1 U11139 ( .A1(n8107), .A2(n10727), .ZN(n11023) );
  XOR2_X1 U11140 ( .A(n11227), .B(n11228), .Z(n11020) );
  XOR2_X1 U11141 ( .A(n11229), .B(n11230), .Z(n11228) );
  OR2_X1 U11142 ( .A1(n11024), .A2(n11027), .ZN(n11072) );
  OR2_X1 U11143 ( .A1(n8025), .A2(n10727), .ZN(n11027) );
  XOR2_X1 U11144 ( .A(n11231), .B(n11232), .Z(n11024) );
  XOR2_X1 U11145 ( .A(n11233), .B(n11234), .Z(n11232) );
  OR2_X1 U11146 ( .A1(n11028), .A2(n11031), .ZN(n11069) );
  OR2_X1 U11147 ( .A1(n7955), .A2(n10727), .ZN(n11031) );
  XOR2_X1 U11148 ( .A(n11235), .B(n11236), .Z(n11028) );
  XOR2_X1 U11149 ( .A(n11237), .B(n11238), .Z(n11236) );
  OR2_X1 U11150 ( .A1(n11032), .A2(n11035), .ZN(n11066) );
  OR2_X1 U11151 ( .A1(n7887), .A2(n10727), .ZN(n11035) );
  XOR2_X1 U11152 ( .A(n11239), .B(n11240), .Z(n11032) );
  XOR2_X1 U11153 ( .A(n11241), .B(n11242), .Z(n11240) );
  OR2_X1 U11154 ( .A1(n11036), .A2(n11039), .ZN(n11063) );
  OR2_X1 U11155 ( .A1(n7828), .A2(n10727), .ZN(n11039) );
  XOR2_X1 U11156 ( .A(n11243), .B(n11244), .Z(n11036) );
  XOR2_X1 U11157 ( .A(n11245), .B(n11246), .Z(n11244) );
  OR2_X1 U11158 ( .A1(n11040), .A2(n11043), .ZN(n11060) );
  OR2_X1 U11159 ( .A1(n7820), .A2(n10727), .ZN(n11043) );
  XOR2_X1 U11160 ( .A(n11247), .B(n11248), .Z(n11040) );
  XOR2_X1 U11161 ( .A(n11249), .B(n11250), .Z(n11248) );
  OR2_X1 U11162 ( .A1(n11044), .A2(n11047), .ZN(n11057) );
  OR2_X1 U11163 ( .A1(n7730), .A2(n10727), .ZN(n11047) );
  XOR2_X1 U11164 ( .A(n11251), .B(n11252), .Z(n11044) );
  XOR2_X1 U11165 ( .A(n11253), .B(n11254), .Z(n11252) );
  OR2_X1 U11166 ( .A1(n10414), .A2(n10417), .ZN(n11054) );
  OR2_X1 U11167 ( .A1(n7697), .A2(n10727), .ZN(n10417) );
  XOR2_X1 U11168 ( .A(n11255), .B(n11256), .Z(n10414) );
  XOR2_X1 U11169 ( .A(n11257), .B(n11258), .Z(n11256) );
  OR2_X1 U11170 ( .A1(n8339), .A2(n8342), .ZN(n11051) );
  OR2_X1 U11171 ( .A1(n7660), .A2(n10727), .ZN(n8342) );
  XOR2_X1 U11172 ( .A(n11259), .B(n11260), .Z(n8339) );
  XOR2_X1 U11173 ( .A(n11261), .B(n11262), .Z(n11260) );
  XOR2_X1 U11174 ( .A(n11263), .B(n11264), .Z(n8322) );
  XOR2_X1 U11175 ( .A(n11265), .B(n11266), .Z(n11264) );
  OR2_X1 U11176 ( .A1(n11267), .A2(n11268), .ZN(n7565) );
  XOR2_X1 U11177 ( .A(n8314), .B(n8313), .Z(n11268) );
  XOR2_X1 U11178 ( .A(n11269), .B(n11270), .Z(n8313) );
  XOR2_X1 U11179 ( .A(n11271), .B(n11272), .Z(n11270) );
  OR2_X1 U11180 ( .A1(n11273), .A2(n11274), .ZN(n8314) );
  AND2_X1 U11181 ( .A1(n11275), .A2(n11276), .ZN(n11274) );
  AND2_X1 U11182 ( .A1(n11277), .A2(n11278), .ZN(n11273) );
  OR2_X1 U11183 ( .A1(n11275), .A2(n11276), .ZN(n11278) );
  AND2_X1 U11184 ( .A1(n11048), .A2(n11279), .ZN(n11267) );
  INV_X1 U11185 ( .A(n8310), .ZN(n11279) );
  XOR2_X1 U11186 ( .A(n11277), .B(n11280), .Z(n8310) );
  XOR2_X1 U11187 ( .A(n11276), .B(n11275), .Z(n11280) );
  OR2_X1 U11188 ( .A1(n7660), .A2(n11144), .ZN(n11275) );
  OR2_X1 U11189 ( .A1(n11281), .A2(n11282), .ZN(n11276) );
  AND2_X1 U11190 ( .A1(n11283), .A2(n11284), .ZN(n11282) );
  AND2_X1 U11191 ( .A1(n11285), .A2(n11286), .ZN(n11281) );
  OR2_X1 U11192 ( .A1(n11283), .A2(n11284), .ZN(n11286) );
  XOR2_X1 U11193 ( .A(n11287), .B(n11288), .Z(n11277) );
  XOR2_X1 U11194 ( .A(n11289), .B(n11290), .Z(n11288) );
  INV_X1 U11195 ( .A(n8311), .ZN(n11048) );
  OR2_X1 U11196 ( .A1(n11291), .A2(n11292), .ZN(n8311) );
  AND2_X1 U11197 ( .A1(n11266), .A2(n11265), .ZN(n11292) );
  AND2_X1 U11198 ( .A1(n11263), .A2(n11293), .ZN(n11291) );
  OR2_X1 U11199 ( .A1(n11265), .A2(n11266), .ZN(n11293) );
  OR2_X1 U11200 ( .A1(n7660), .A2(n10933), .ZN(n11266) );
  OR2_X1 U11201 ( .A1(n11294), .A2(n11295), .ZN(n11265) );
  AND2_X1 U11202 ( .A1(n11262), .A2(n11261), .ZN(n11295) );
  AND2_X1 U11203 ( .A1(n11259), .A2(n11296), .ZN(n11294) );
  OR2_X1 U11204 ( .A1(n11261), .A2(n11262), .ZN(n11296) );
  OR2_X1 U11205 ( .A1(n7697), .A2(n10933), .ZN(n11262) );
  OR2_X1 U11206 ( .A1(n11297), .A2(n11298), .ZN(n11261) );
  AND2_X1 U11207 ( .A1(n11258), .A2(n11257), .ZN(n11298) );
  AND2_X1 U11208 ( .A1(n11255), .A2(n11299), .ZN(n11297) );
  OR2_X1 U11209 ( .A1(n11257), .A2(n11258), .ZN(n11299) );
  OR2_X1 U11210 ( .A1(n7730), .A2(n10933), .ZN(n11258) );
  OR2_X1 U11211 ( .A1(n11300), .A2(n11301), .ZN(n11257) );
  AND2_X1 U11212 ( .A1(n11254), .A2(n11253), .ZN(n11301) );
  AND2_X1 U11213 ( .A1(n11251), .A2(n11302), .ZN(n11300) );
  OR2_X1 U11214 ( .A1(n11253), .A2(n11254), .ZN(n11302) );
  OR2_X1 U11215 ( .A1(n7820), .A2(n10933), .ZN(n11254) );
  OR2_X1 U11216 ( .A1(n11303), .A2(n11304), .ZN(n11253) );
  AND2_X1 U11217 ( .A1(n11250), .A2(n11249), .ZN(n11304) );
  AND2_X1 U11218 ( .A1(n11247), .A2(n11305), .ZN(n11303) );
  OR2_X1 U11219 ( .A1(n11249), .A2(n11250), .ZN(n11305) );
  OR2_X1 U11220 ( .A1(n7828), .A2(n10933), .ZN(n11250) );
  OR2_X1 U11221 ( .A1(n11306), .A2(n11307), .ZN(n11249) );
  AND2_X1 U11222 ( .A1(n11246), .A2(n11245), .ZN(n11307) );
  AND2_X1 U11223 ( .A1(n11243), .A2(n11308), .ZN(n11306) );
  OR2_X1 U11224 ( .A1(n11245), .A2(n11246), .ZN(n11308) );
  OR2_X1 U11225 ( .A1(n7887), .A2(n10933), .ZN(n11246) );
  OR2_X1 U11226 ( .A1(n11309), .A2(n11310), .ZN(n11245) );
  AND2_X1 U11227 ( .A1(n11242), .A2(n11241), .ZN(n11310) );
  AND2_X1 U11228 ( .A1(n11239), .A2(n11311), .ZN(n11309) );
  OR2_X1 U11229 ( .A1(n11241), .A2(n11242), .ZN(n11311) );
  OR2_X1 U11230 ( .A1(n7955), .A2(n10933), .ZN(n11242) );
  OR2_X1 U11231 ( .A1(n11312), .A2(n11313), .ZN(n11241) );
  AND2_X1 U11232 ( .A1(n11238), .A2(n11237), .ZN(n11313) );
  AND2_X1 U11233 ( .A1(n11235), .A2(n11314), .ZN(n11312) );
  OR2_X1 U11234 ( .A1(n11237), .A2(n11238), .ZN(n11314) );
  OR2_X1 U11235 ( .A1(n8025), .A2(n10933), .ZN(n11238) );
  OR2_X1 U11236 ( .A1(n11315), .A2(n11316), .ZN(n11237) );
  AND2_X1 U11237 ( .A1(n11234), .A2(n11233), .ZN(n11316) );
  AND2_X1 U11238 ( .A1(n11231), .A2(n11317), .ZN(n11315) );
  OR2_X1 U11239 ( .A1(n11233), .A2(n11234), .ZN(n11317) );
  OR2_X1 U11240 ( .A1(n8107), .A2(n10933), .ZN(n11234) );
  OR2_X1 U11241 ( .A1(n11318), .A2(n11319), .ZN(n11233) );
  AND2_X1 U11242 ( .A1(n11230), .A2(n11229), .ZN(n11319) );
  AND2_X1 U11243 ( .A1(n11227), .A2(n11320), .ZN(n11318) );
  OR2_X1 U11244 ( .A1(n11229), .A2(n11230), .ZN(n11320) );
  OR2_X1 U11245 ( .A1(n8191), .A2(n10933), .ZN(n11230) );
  OR2_X1 U11246 ( .A1(n11321), .A2(n11322), .ZN(n11229) );
  AND2_X1 U11247 ( .A1(n11226), .A2(n11225), .ZN(n11322) );
  AND2_X1 U11248 ( .A1(n11223), .A2(n11323), .ZN(n11321) );
  OR2_X1 U11249 ( .A1(n11225), .A2(n11226), .ZN(n11323) );
  OR2_X1 U11250 ( .A1(n8287), .A2(n10933), .ZN(n11226) );
  OR2_X1 U11251 ( .A1(n11324), .A2(n11325), .ZN(n11225) );
  AND2_X1 U11252 ( .A1(n11222), .A2(n11221), .ZN(n11325) );
  AND2_X1 U11253 ( .A1(n11219), .A2(n11326), .ZN(n11324) );
  OR2_X1 U11254 ( .A1(n11221), .A2(n11222), .ZN(n11326) );
  OR2_X1 U11255 ( .A1(n8608), .A2(n10933), .ZN(n11222) );
  OR2_X1 U11256 ( .A1(n11327), .A2(n11328), .ZN(n11221) );
  AND2_X1 U11257 ( .A1(n11218), .A2(n11217), .ZN(n11328) );
  AND2_X1 U11258 ( .A1(n11215), .A2(n11329), .ZN(n11327) );
  OR2_X1 U11259 ( .A1(n11217), .A2(n11218), .ZN(n11329) );
  OR2_X1 U11260 ( .A1(n8603), .A2(n10933), .ZN(n11218) );
  OR2_X1 U11261 ( .A1(n11330), .A2(n11331), .ZN(n11217) );
  AND2_X1 U11262 ( .A1(n11214), .A2(n11213), .ZN(n11331) );
  AND2_X1 U11263 ( .A1(n11211), .A2(n11332), .ZN(n11330) );
  OR2_X1 U11264 ( .A1(n11213), .A2(n11214), .ZN(n11332) );
  OR2_X1 U11265 ( .A1(n8598), .A2(n10933), .ZN(n11214) );
  OR2_X1 U11266 ( .A1(n11333), .A2(n11334), .ZN(n11213) );
  AND2_X1 U11267 ( .A1(n11210), .A2(n11209), .ZN(n11334) );
  AND2_X1 U11268 ( .A1(n11207), .A2(n11335), .ZN(n11333) );
  OR2_X1 U11269 ( .A1(n11209), .A2(n11210), .ZN(n11335) );
  OR2_X1 U11270 ( .A1(n8593), .A2(n10933), .ZN(n11210) );
  OR2_X1 U11271 ( .A1(n11336), .A2(n11337), .ZN(n11209) );
  AND2_X1 U11272 ( .A1(n11206), .A2(n11205), .ZN(n11337) );
  AND2_X1 U11273 ( .A1(n11203), .A2(n11338), .ZN(n11336) );
  OR2_X1 U11274 ( .A1(n11205), .A2(n11206), .ZN(n11338) );
  OR2_X1 U11275 ( .A1(n8588), .A2(n10933), .ZN(n11206) );
  OR2_X1 U11276 ( .A1(n11339), .A2(n11340), .ZN(n11205) );
  AND2_X1 U11277 ( .A1(n11202), .A2(n11201), .ZN(n11340) );
  AND2_X1 U11278 ( .A1(n11199), .A2(n11341), .ZN(n11339) );
  OR2_X1 U11279 ( .A1(n11201), .A2(n11202), .ZN(n11341) );
  OR2_X1 U11280 ( .A1(n8583), .A2(n10933), .ZN(n11202) );
  OR2_X1 U11281 ( .A1(n11342), .A2(n11343), .ZN(n11201) );
  AND2_X1 U11282 ( .A1(n11198), .A2(n11197), .ZN(n11343) );
  AND2_X1 U11283 ( .A1(n11195), .A2(n11344), .ZN(n11342) );
  OR2_X1 U11284 ( .A1(n11197), .A2(n11198), .ZN(n11344) );
  OR2_X1 U11285 ( .A1(n8578), .A2(n10933), .ZN(n11198) );
  OR2_X1 U11286 ( .A1(n11345), .A2(n11346), .ZN(n11197) );
  AND2_X1 U11287 ( .A1(n11192), .A2(n11194), .ZN(n11346) );
  AND2_X1 U11288 ( .A1(n11347), .A2(n11193), .ZN(n11345) );
  OR2_X1 U11289 ( .A1(n11194), .A2(n11192), .ZN(n11347) );
  XOR2_X1 U11290 ( .A(n11348), .B(n11349), .Z(n11192) );
  XOR2_X1 U11291 ( .A(n11350), .B(n11351), .Z(n11349) );
  OR2_X1 U11292 ( .A1(n11352), .A2(n11353), .ZN(n11194) );
  AND2_X1 U11293 ( .A1(n11190), .A2(n11189), .ZN(n11353) );
  AND2_X1 U11294 ( .A1(n11187), .A2(n11354), .ZN(n11352) );
  OR2_X1 U11295 ( .A1(n11189), .A2(n11190), .ZN(n11354) );
  OR2_X1 U11296 ( .A1(n8568), .A2(n10933), .ZN(n11190) );
  OR2_X1 U11297 ( .A1(n11355), .A2(n11356), .ZN(n11189) );
  AND2_X1 U11298 ( .A1(n11186), .A2(n11185), .ZN(n11356) );
  AND2_X1 U11299 ( .A1(n11183), .A2(n11357), .ZN(n11355) );
  OR2_X1 U11300 ( .A1(n11185), .A2(n11186), .ZN(n11357) );
  OR2_X1 U11301 ( .A1(n8563), .A2(n10933), .ZN(n11186) );
  OR2_X1 U11302 ( .A1(n11358), .A2(n11359), .ZN(n11185) );
  AND2_X1 U11303 ( .A1(n11182), .A2(n11181), .ZN(n11359) );
  AND2_X1 U11304 ( .A1(n11179), .A2(n11360), .ZN(n11358) );
  OR2_X1 U11305 ( .A1(n11181), .A2(n11182), .ZN(n11360) );
  OR2_X1 U11306 ( .A1(n8558), .A2(n10933), .ZN(n11182) );
  OR2_X1 U11307 ( .A1(n11361), .A2(n11362), .ZN(n11181) );
  AND2_X1 U11308 ( .A1(n11178), .A2(n11177), .ZN(n11362) );
  AND2_X1 U11309 ( .A1(n11175), .A2(n11363), .ZN(n11361) );
  OR2_X1 U11310 ( .A1(n11177), .A2(n11178), .ZN(n11363) );
  OR2_X1 U11311 ( .A1(n8553), .A2(n10933), .ZN(n11178) );
  OR2_X1 U11312 ( .A1(n11364), .A2(n11365), .ZN(n11177) );
  AND2_X1 U11313 ( .A1(n11174), .A2(n11173), .ZN(n11365) );
  AND2_X1 U11314 ( .A1(n11171), .A2(n11366), .ZN(n11364) );
  OR2_X1 U11315 ( .A1(n11173), .A2(n11174), .ZN(n11366) );
  OR2_X1 U11316 ( .A1(n8548), .A2(n10933), .ZN(n11174) );
  OR2_X1 U11317 ( .A1(n11367), .A2(n11368), .ZN(n11173) );
  AND2_X1 U11318 ( .A1(n11170), .A2(n11169), .ZN(n11368) );
  AND2_X1 U11319 ( .A1(n11167), .A2(n11369), .ZN(n11367) );
  OR2_X1 U11320 ( .A1(n11169), .A2(n11170), .ZN(n11369) );
  OR2_X1 U11321 ( .A1(n8543), .A2(n10933), .ZN(n11170) );
  OR2_X1 U11322 ( .A1(n11370), .A2(n11371), .ZN(n11169) );
  AND2_X1 U11323 ( .A1(n11166), .A2(n11165), .ZN(n11371) );
  AND2_X1 U11324 ( .A1(n11163), .A2(n11372), .ZN(n11370) );
  OR2_X1 U11325 ( .A1(n11165), .A2(n11166), .ZN(n11372) );
  OR2_X1 U11326 ( .A1(n8538), .A2(n10933), .ZN(n11166) );
  OR2_X1 U11327 ( .A1(n11373), .A2(n11374), .ZN(n11165) );
  AND2_X1 U11328 ( .A1(n11162), .A2(n11161), .ZN(n11374) );
  AND2_X1 U11329 ( .A1(n11159), .A2(n11375), .ZN(n11373) );
  OR2_X1 U11330 ( .A1(n11161), .A2(n11162), .ZN(n11375) );
  OR2_X1 U11331 ( .A1(n8533), .A2(n10933), .ZN(n11162) );
  OR2_X1 U11332 ( .A1(n11376), .A2(n11377), .ZN(n11161) );
  AND2_X1 U11333 ( .A1(n11158), .A2(n11157), .ZN(n11377) );
  AND2_X1 U11334 ( .A1(n11155), .A2(n11378), .ZN(n11376) );
  OR2_X1 U11335 ( .A1(n11157), .A2(n11158), .ZN(n11378) );
  OR2_X1 U11336 ( .A1(n8528), .A2(n10933), .ZN(n11158) );
  OR2_X1 U11337 ( .A1(n11379), .A2(n11380), .ZN(n11157) );
  AND2_X1 U11338 ( .A1(n11154), .A2(n11153), .ZN(n11380) );
  AND2_X1 U11339 ( .A1(n11151), .A2(n11381), .ZN(n11379) );
  OR2_X1 U11340 ( .A1(n11153), .A2(n11154), .ZN(n11381) );
  OR2_X1 U11341 ( .A1(n8523), .A2(n10933), .ZN(n11154) );
  OR2_X1 U11342 ( .A1(n11382), .A2(n11383), .ZN(n11153) );
  AND2_X1 U11343 ( .A1(n11148), .A2(n11149), .ZN(n11383) );
  AND2_X1 U11344 ( .A1(n11384), .A2(n11385), .ZN(n11382) );
  OR2_X1 U11345 ( .A1(n11149), .A2(n11148), .ZN(n11385) );
  OR2_X1 U11346 ( .A1(n8515), .A2(n10933), .ZN(n11148) );
  OR2_X1 U11347 ( .A1(n10933), .A2(n11386), .ZN(n11149) );
  INV_X1 U11348 ( .A(n11150), .ZN(n11384) );
  OR2_X1 U11349 ( .A1(n11387), .A2(n11388), .ZN(n11150) );
  AND2_X1 U11350 ( .A1(b_17_), .A2(n11389), .ZN(n11388) );
  OR2_X1 U11351 ( .A1(n11390), .A2(n7343), .ZN(n11389) );
  AND2_X1 U11352 ( .A1(a_30_), .A2(n11391), .ZN(n11390) );
  AND2_X1 U11353 ( .A1(b_16_), .A2(n11392), .ZN(n11387) );
  OR2_X1 U11354 ( .A1(n11393), .A2(n7347), .ZN(n11392) );
  AND2_X1 U11355 ( .A1(a_31_), .A2(n11144), .ZN(n11393) );
  XOR2_X1 U11356 ( .A(n11394), .B(n11395), .Z(n11151) );
  XNOR2_X1 U11357 ( .A(n11396), .B(n11397), .ZN(n11394) );
  XOR2_X1 U11358 ( .A(n11398), .B(n11399), .Z(n11155) );
  XOR2_X1 U11359 ( .A(n11400), .B(n11401), .Z(n11399) );
  XOR2_X1 U11360 ( .A(n11402), .B(n11403), .Z(n11159) );
  XOR2_X1 U11361 ( .A(n11404), .B(n11405), .Z(n11403) );
  XOR2_X1 U11362 ( .A(n11406), .B(n11407), .Z(n11163) );
  XOR2_X1 U11363 ( .A(n11408), .B(n11409), .Z(n11407) );
  XOR2_X1 U11364 ( .A(n11410), .B(n11411), .Z(n11167) );
  XOR2_X1 U11365 ( .A(n11412), .B(n11413), .Z(n11411) );
  XOR2_X1 U11366 ( .A(n11414), .B(n11415), .Z(n11171) );
  XOR2_X1 U11367 ( .A(n11416), .B(n11417), .Z(n11415) );
  XOR2_X1 U11368 ( .A(n11418), .B(n11419), .Z(n11175) );
  XOR2_X1 U11369 ( .A(n11420), .B(n11421), .Z(n11419) );
  XOR2_X1 U11370 ( .A(n11422), .B(n11423), .Z(n11179) );
  XOR2_X1 U11371 ( .A(n11424), .B(n11425), .Z(n11423) );
  XOR2_X1 U11372 ( .A(n11426), .B(n11427), .Z(n11183) );
  XOR2_X1 U11373 ( .A(n11428), .B(n11429), .Z(n11427) );
  XOR2_X1 U11374 ( .A(n11430), .B(n11431), .Z(n11187) );
  XOR2_X1 U11375 ( .A(n11432), .B(n11433), .Z(n11431) );
  XOR2_X1 U11376 ( .A(n11434), .B(n11435), .Z(n11195) );
  XOR2_X1 U11377 ( .A(n11436), .B(n11437), .Z(n11435) );
  XNOR2_X1 U11378 ( .A(n11438), .B(n11439), .ZN(n11199) );
  XNOR2_X1 U11379 ( .A(n11440), .B(n11441), .ZN(n11438) );
  XOR2_X1 U11380 ( .A(n11442), .B(n11443), .Z(n11203) );
  XOR2_X1 U11381 ( .A(n11444), .B(n11445), .Z(n11443) );
  XOR2_X1 U11382 ( .A(n11446), .B(n11447), .Z(n11207) );
  XOR2_X1 U11383 ( .A(n11448), .B(n11449), .Z(n11447) );
  XOR2_X1 U11384 ( .A(n11450), .B(n11451), .Z(n11211) );
  XOR2_X1 U11385 ( .A(n11452), .B(n11453), .Z(n11451) );
  XOR2_X1 U11386 ( .A(n11454), .B(n11455), .Z(n11215) );
  XOR2_X1 U11387 ( .A(n11456), .B(n11457), .Z(n11455) );
  XOR2_X1 U11388 ( .A(n11458), .B(n11459), .Z(n11219) );
  XOR2_X1 U11389 ( .A(n11460), .B(n11461), .Z(n11459) );
  XOR2_X1 U11390 ( .A(n11462), .B(n11463), .Z(n11223) );
  XOR2_X1 U11391 ( .A(n11464), .B(n11465), .Z(n11463) );
  XOR2_X1 U11392 ( .A(n11466), .B(n11467), .Z(n11227) );
  XOR2_X1 U11393 ( .A(n11468), .B(n11469), .Z(n11467) );
  XOR2_X1 U11394 ( .A(n11470), .B(n11471), .Z(n11231) );
  XOR2_X1 U11395 ( .A(n11472), .B(n11473), .Z(n11471) );
  XOR2_X1 U11396 ( .A(n11474), .B(n11475), .Z(n11235) );
  XOR2_X1 U11397 ( .A(n11476), .B(n11477), .Z(n11475) );
  XOR2_X1 U11398 ( .A(n11478), .B(n11479), .Z(n11239) );
  XOR2_X1 U11399 ( .A(n11480), .B(n11481), .Z(n11479) );
  XOR2_X1 U11400 ( .A(n11482), .B(n11483), .Z(n11243) );
  XOR2_X1 U11401 ( .A(n11484), .B(n11485), .Z(n11483) );
  XOR2_X1 U11402 ( .A(n11486), .B(n11487), .Z(n11247) );
  XOR2_X1 U11403 ( .A(n11488), .B(n11489), .Z(n11487) );
  XOR2_X1 U11404 ( .A(n11490), .B(n11491), .Z(n11251) );
  XOR2_X1 U11405 ( .A(n11492), .B(n11493), .Z(n11491) );
  XOR2_X1 U11406 ( .A(n11494), .B(n11495), .Z(n11255) );
  XOR2_X1 U11407 ( .A(n11496), .B(n11497), .Z(n11495) );
  XOR2_X1 U11408 ( .A(n11498), .B(n11499), .Z(n11259) );
  XOR2_X1 U11409 ( .A(n11500), .B(n11501), .Z(n11499) );
  XOR2_X1 U11410 ( .A(n11285), .B(n11502), .Z(n11263) );
  XOR2_X1 U11411 ( .A(n11284), .B(n11283), .Z(n11502) );
  OR2_X1 U11412 ( .A1(n7697), .A2(n11144), .ZN(n11283) );
  OR2_X1 U11413 ( .A1(n11503), .A2(n11504), .ZN(n11284) );
  AND2_X1 U11414 ( .A1(n11501), .A2(n11500), .ZN(n11504) );
  AND2_X1 U11415 ( .A1(n11498), .A2(n11505), .ZN(n11503) );
  OR2_X1 U11416 ( .A1(n11501), .A2(n11500), .ZN(n11505) );
  OR2_X1 U11417 ( .A1(n11506), .A2(n11507), .ZN(n11500) );
  AND2_X1 U11418 ( .A1(n11497), .A2(n11496), .ZN(n11507) );
  AND2_X1 U11419 ( .A1(n11494), .A2(n11508), .ZN(n11506) );
  OR2_X1 U11420 ( .A1(n11497), .A2(n11496), .ZN(n11508) );
  OR2_X1 U11421 ( .A1(n11509), .A2(n11510), .ZN(n11496) );
  AND2_X1 U11422 ( .A1(n11493), .A2(n11492), .ZN(n11510) );
  AND2_X1 U11423 ( .A1(n11490), .A2(n11511), .ZN(n11509) );
  OR2_X1 U11424 ( .A1(n11493), .A2(n11492), .ZN(n11511) );
  OR2_X1 U11425 ( .A1(n11512), .A2(n11513), .ZN(n11492) );
  AND2_X1 U11426 ( .A1(n11489), .A2(n11488), .ZN(n11513) );
  AND2_X1 U11427 ( .A1(n11486), .A2(n11514), .ZN(n11512) );
  OR2_X1 U11428 ( .A1(n11489), .A2(n11488), .ZN(n11514) );
  OR2_X1 U11429 ( .A1(n11515), .A2(n11516), .ZN(n11488) );
  AND2_X1 U11430 ( .A1(n11485), .A2(n11484), .ZN(n11516) );
  AND2_X1 U11431 ( .A1(n11482), .A2(n11517), .ZN(n11515) );
  OR2_X1 U11432 ( .A1(n11485), .A2(n11484), .ZN(n11517) );
  OR2_X1 U11433 ( .A1(n11518), .A2(n11519), .ZN(n11484) );
  AND2_X1 U11434 ( .A1(n11481), .A2(n11480), .ZN(n11519) );
  AND2_X1 U11435 ( .A1(n11478), .A2(n11520), .ZN(n11518) );
  OR2_X1 U11436 ( .A1(n11481), .A2(n11480), .ZN(n11520) );
  OR2_X1 U11437 ( .A1(n11521), .A2(n11522), .ZN(n11480) );
  AND2_X1 U11438 ( .A1(n11477), .A2(n11476), .ZN(n11522) );
  AND2_X1 U11439 ( .A1(n11474), .A2(n11523), .ZN(n11521) );
  OR2_X1 U11440 ( .A1(n11477), .A2(n11476), .ZN(n11523) );
  OR2_X1 U11441 ( .A1(n11524), .A2(n11525), .ZN(n11476) );
  AND2_X1 U11442 ( .A1(n11473), .A2(n11472), .ZN(n11525) );
  AND2_X1 U11443 ( .A1(n11470), .A2(n11526), .ZN(n11524) );
  OR2_X1 U11444 ( .A1(n11473), .A2(n11472), .ZN(n11526) );
  OR2_X1 U11445 ( .A1(n11527), .A2(n11528), .ZN(n11472) );
  AND2_X1 U11446 ( .A1(n11469), .A2(n11468), .ZN(n11528) );
  AND2_X1 U11447 ( .A1(n11466), .A2(n11529), .ZN(n11527) );
  OR2_X1 U11448 ( .A1(n11469), .A2(n11468), .ZN(n11529) );
  OR2_X1 U11449 ( .A1(n11530), .A2(n11531), .ZN(n11468) );
  AND2_X1 U11450 ( .A1(n11465), .A2(n11464), .ZN(n11531) );
  AND2_X1 U11451 ( .A1(n11462), .A2(n11532), .ZN(n11530) );
  OR2_X1 U11452 ( .A1(n11465), .A2(n11464), .ZN(n11532) );
  OR2_X1 U11453 ( .A1(n11533), .A2(n11534), .ZN(n11464) );
  AND2_X1 U11454 ( .A1(n11461), .A2(n11460), .ZN(n11534) );
  AND2_X1 U11455 ( .A1(n11458), .A2(n11535), .ZN(n11533) );
  OR2_X1 U11456 ( .A1(n11461), .A2(n11460), .ZN(n11535) );
  OR2_X1 U11457 ( .A1(n11536), .A2(n11537), .ZN(n11460) );
  AND2_X1 U11458 ( .A1(n11457), .A2(n11456), .ZN(n11537) );
  AND2_X1 U11459 ( .A1(n11454), .A2(n11538), .ZN(n11536) );
  OR2_X1 U11460 ( .A1(n11457), .A2(n11456), .ZN(n11538) );
  OR2_X1 U11461 ( .A1(n11539), .A2(n11540), .ZN(n11456) );
  AND2_X1 U11462 ( .A1(n11453), .A2(n11452), .ZN(n11540) );
  AND2_X1 U11463 ( .A1(n11450), .A2(n11541), .ZN(n11539) );
  OR2_X1 U11464 ( .A1(n11453), .A2(n11452), .ZN(n11541) );
  OR2_X1 U11465 ( .A1(n11542), .A2(n11543), .ZN(n11452) );
  AND2_X1 U11466 ( .A1(n11449), .A2(n11448), .ZN(n11543) );
  AND2_X1 U11467 ( .A1(n11446), .A2(n11544), .ZN(n11542) );
  OR2_X1 U11468 ( .A1(n11449), .A2(n11448), .ZN(n11544) );
  OR2_X1 U11469 ( .A1(n11545), .A2(n11546), .ZN(n11448) );
  AND2_X1 U11470 ( .A1(n11445), .A2(n11444), .ZN(n11546) );
  AND2_X1 U11471 ( .A1(n11442), .A2(n11547), .ZN(n11545) );
  OR2_X1 U11472 ( .A1(n11445), .A2(n11444), .ZN(n11547) );
  OR2_X1 U11473 ( .A1(n11548), .A2(n11549), .ZN(n11444) );
  AND2_X1 U11474 ( .A1(n11439), .A2(n11441), .ZN(n11549) );
  AND2_X1 U11475 ( .A1(n11550), .A2(n11440), .ZN(n11548) );
  OR2_X1 U11476 ( .A1(n11439), .A2(n11441), .ZN(n11550) );
  OR2_X1 U11477 ( .A1(n11551), .A2(n11552), .ZN(n11441) );
  AND2_X1 U11478 ( .A1(n11437), .A2(n11436), .ZN(n11552) );
  AND2_X1 U11479 ( .A1(n11434), .A2(n11553), .ZN(n11551) );
  OR2_X1 U11480 ( .A1(n11437), .A2(n11436), .ZN(n11553) );
  OR2_X1 U11481 ( .A1(n11554), .A2(n11555), .ZN(n11436) );
  AND2_X1 U11482 ( .A1(n11351), .A2(n11350), .ZN(n11555) );
  AND2_X1 U11483 ( .A1(n11348), .A2(n11556), .ZN(n11554) );
  OR2_X1 U11484 ( .A1(n11351), .A2(n11350), .ZN(n11556) );
  OR2_X1 U11485 ( .A1(n11557), .A2(n11558), .ZN(n11350) );
  AND2_X1 U11486 ( .A1(n11433), .A2(n11432), .ZN(n11558) );
  AND2_X1 U11487 ( .A1(n11430), .A2(n11559), .ZN(n11557) );
  OR2_X1 U11488 ( .A1(n11433), .A2(n11432), .ZN(n11559) );
  OR2_X1 U11489 ( .A1(n11560), .A2(n11561), .ZN(n11432) );
  AND2_X1 U11490 ( .A1(n11429), .A2(n11428), .ZN(n11561) );
  AND2_X1 U11491 ( .A1(n11426), .A2(n11562), .ZN(n11560) );
  OR2_X1 U11492 ( .A1(n11429), .A2(n11428), .ZN(n11562) );
  OR2_X1 U11493 ( .A1(n11563), .A2(n11564), .ZN(n11428) );
  AND2_X1 U11494 ( .A1(n11425), .A2(n11424), .ZN(n11564) );
  AND2_X1 U11495 ( .A1(n11422), .A2(n11565), .ZN(n11563) );
  OR2_X1 U11496 ( .A1(n11425), .A2(n11424), .ZN(n11565) );
  OR2_X1 U11497 ( .A1(n11566), .A2(n11567), .ZN(n11424) );
  AND2_X1 U11498 ( .A1(n11421), .A2(n11420), .ZN(n11567) );
  AND2_X1 U11499 ( .A1(n11418), .A2(n11568), .ZN(n11566) );
  OR2_X1 U11500 ( .A1(n11421), .A2(n11420), .ZN(n11568) );
  OR2_X1 U11501 ( .A1(n11569), .A2(n11570), .ZN(n11420) );
  AND2_X1 U11502 ( .A1(n11417), .A2(n11416), .ZN(n11570) );
  AND2_X1 U11503 ( .A1(n11414), .A2(n11571), .ZN(n11569) );
  OR2_X1 U11504 ( .A1(n11417), .A2(n11416), .ZN(n11571) );
  OR2_X1 U11505 ( .A1(n11572), .A2(n11573), .ZN(n11416) );
  AND2_X1 U11506 ( .A1(n11413), .A2(n11412), .ZN(n11573) );
  AND2_X1 U11507 ( .A1(n11410), .A2(n11574), .ZN(n11572) );
  OR2_X1 U11508 ( .A1(n11413), .A2(n11412), .ZN(n11574) );
  OR2_X1 U11509 ( .A1(n11575), .A2(n11576), .ZN(n11412) );
  AND2_X1 U11510 ( .A1(n11409), .A2(n11408), .ZN(n11576) );
  AND2_X1 U11511 ( .A1(n11406), .A2(n11577), .ZN(n11575) );
  OR2_X1 U11512 ( .A1(n11409), .A2(n11408), .ZN(n11577) );
  OR2_X1 U11513 ( .A1(n11578), .A2(n11579), .ZN(n11408) );
  AND2_X1 U11514 ( .A1(n11405), .A2(n11404), .ZN(n11579) );
  AND2_X1 U11515 ( .A1(n11402), .A2(n11580), .ZN(n11578) );
  OR2_X1 U11516 ( .A1(n11405), .A2(n11404), .ZN(n11580) );
  OR2_X1 U11517 ( .A1(n11581), .A2(n11582), .ZN(n11404) );
  AND2_X1 U11518 ( .A1(n11401), .A2(n11400), .ZN(n11582) );
  AND2_X1 U11519 ( .A1(n11398), .A2(n11583), .ZN(n11581) );
  OR2_X1 U11520 ( .A1(n11401), .A2(n11400), .ZN(n11583) );
  OR2_X1 U11521 ( .A1(n11584), .A2(n11585), .ZN(n11400) );
  AND2_X1 U11522 ( .A1(n11395), .A2(n11396), .ZN(n11585) );
  AND2_X1 U11523 ( .A1(n11586), .A2(n11587), .ZN(n11584) );
  OR2_X1 U11524 ( .A1(n11395), .A2(n11396), .ZN(n11587) );
  OR2_X1 U11525 ( .A1(n11391), .A2(n11386), .ZN(n11396) );
  OR2_X1 U11526 ( .A1(n8956), .A2(n11144), .ZN(n11386) );
  OR2_X1 U11527 ( .A1(n8515), .A2(n11144), .ZN(n11395) );
  INV_X1 U11528 ( .A(n11397), .ZN(n11586) );
  OR2_X1 U11529 ( .A1(n11588), .A2(n11589), .ZN(n11397) );
  AND2_X1 U11530 ( .A1(b_16_), .A2(n11590), .ZN(n11589) );
  OR2_X1 U11531 ( .A1(n11591), .A2(n7343), .ZN(n11590) );
  AND2_X1 U11532 ( .A1(a_30_), .A2(n11592), .ZN(n11591) );
  AND2_X1 U11533 ( .A1(b_15_), .A2(n11593), .ZN(n11588) );
  OR2_X1 U11534 ( .A1(n11594), .A2(n7347), .ZN(n11593) );
  AND2_X1 U11535 ( .A1(a_31_), .A2(n11391), .ZN(n11594) );
  OR2_X1 U11536 ( .A1(n8523), .A2(n11144), .ZN(n11401) );
  XOR2_X1 U11537 ( .A(n11595), .B(n11596), .Z(n11398) );
  XNOR2_X1 U11538 ( .A(n11597), .B(n11598), .ZN(n11595) );
  OR2_X1 U11539 ( .A1(n8528), .A2(n11144), .ZN(n11405) );
  XOR2_X1 U11540 ( .A(n11599), .B(n11600), .Z(n11402) );
  XOR2_X1 U11541 ( .A(n11601), .B(n11602), .Z(n11600) );
  OR2_X1 U11542 ( .A1(n8533), .A2(n11144), .ZN(n11409) );
  XOR2_X1 U11543 ( .A(n11603), .B(n11604), .Z(n11406) );
  XOR2_X1 U11544 ( .A(n11605), .B(n11606), .Z(n11604) );
  OR2_X1 U11545 ( .A1(n8538), .A2(n11144), .ZN(n11413) );
  XOR2_X1 U11546 ( .A(n11607), .B(n11608), .Z(n11410) );
  XOR2_X1 U11547 ( .A(n11609), .B(n11610), .Z(n11608) );
  OR2_X1 U11548 ( .A1(n8543), .A2(n11144), .ZN(n11417) );
  XOR2_X1 U11549 ( .A(n11611), .B(n11612), .Z(n11414) );
  XOR2_X1 U11550 ( .A(n11613), .B(n11614), .Z(n11612) );
  OR2_X1 U11551 ( .A1(n8548), .A2(n11144), .ZN(n11421) );
  XOR2_X1 U11552 ( .A(n11615), .B(n11616), .Z(n11418) );
  XOR2_X1 U11553 ( .A(n11617), .B(n11618), .Z(n11616) );
  OR2_X1 U11554 ( .A1(n8553), .A2(n11144), .ZN(n11425) );
  XOR2_X1 U11555 ( .A(n11619), .B(n11620), .Z(n11422) );
  XOR2_X1 U11556 ( .A(n11621), .B(n11622), .Z(n11620) );
  OR2_X1 U11557 ( .A1(n8558), .A2(n11144), .ZN(n11429) );
  XOR2_X1 U11558 ( .A(n11623), .B(n11624), .Z(n11426) );
  XOR2_X1 U11559 ( .A(n11625), .B(n11626), .Z(n11624) );
  OR2_X1 U11560 ( .A1(n8563), .A2(n11144), .ZN(n11433) );
  XOR2_X1 U11561 ( .A(n11627), .B(n11628), .Z(n11430) );
  XOR2_X1 U11562 ( .A(n11629), .B(n11630), .Z(n11628) );
  OR2_X1 U11563 ( .A1(n8568), .A2(n11144), .ZN(n11351) );
  XOR2_X1 U11564 ( .A(n11631), .B(n11632), .Z(n11348) );
  XOR2_X1 U11565 ( .A(n11633), .B(n11634), .Z(n11632) );
  OR2_X1 U11566 ( .A1(n8573), .A2(n11144), .ZN(n11437) );
  XOR2_X1 U11567 ( .A(n11635), .B(n11636), .Z(n11434) );
  XOR2_X1 U11568 ( .A(n11637), .B(n11638), .Z(n11636) );
  XOR2_X1 U11569 ( .A(n11639), .B(n11640), .Z(n11439) );
  XOR2_X1 U11570 ( .A(n11641), .B(n11642), .Z(n11640) );
  OR2_X1 U11571 ( .A1(n8583), .A2(n11144), .ZN(n11445) );
  XOR2_X1 U11572 ( .A(n11643), .B(n11644), .Z(n11442) );
  XOR2_X1 U11573 ( .A(n11645), .B(n11646), .Z(n11644) );
  OR2_X1 U11574 ( .A1(n8588), .A2(n11144), .ZN(n11449) );
  XNOR2_X1 U11575 ( .A(n11647), .B(n11648), .ZN(n11446) );
  XNOR2_X1 U11576 ( .A(n11649), .B(n11650), .ZN(n11647) );
  OR2_X1 U11577 ( .A1(n8593), .A2(n11144), .ZN(n11453) );
  XOR2_X1 U11578 ( .A(n11651), .B(n11652), .Z(n11450) );
  XOR2_X1 U11579 ( .A(n11653), .B(n11654), .Z(n11652) );
  OR2_X1 U11580 ( .A1(n8598), .A2(n11144), .ZN(n11457) );
  XOR2_X1 U11581 ( .A(n11655), .B(n11656), .Z(n11454) );
  XOR2_X1 U11582 ( .A(n11657), .B(n11658), .Z(n11656) );
  OR2_X1 U11583 ( .A1(n8603), .A2(n11144), .ZN(n11461) );
  XOR2_X1 U11584 ( .A(n11659), .B(n11660), .Z(n11458) );
  XOR2_X1 U11585 ( .A(n11661), .B(n11662), .Z(n11660) );
  OR2_X1 U11586 ( .A1(n8608), .A2(n11144), .ZN(n11465) );
  XOR2_X1 U11587 ( .A(n11663), .B(n11664), .Z(n11462) );
  XOR2_X1 U11588 ( .A(n11665), .B(n11666), .Z(n11664) );
  OR2_X1 U11589 ( .A1(n8287), .A2(n11144), .ZN(n11469) );
  XOR2_X1 U11590 ( .A(n11667), .B(n11668), .Z(n11466) );
  XOR2_X1 U11591 ( .A(n11669), .B(n11670), .Z(n11668) );
  OR2_X1 U11592 ( .A1(n8191), .A2(n11144), .ZN(n11473) );
  XOR2_X1 U11593 ( .A(n11671), .B(n11672), .Z(n11470) );
  XOR2_X1 U11594 ( .A(n11673), .B(n11674), .Z(n11672) );
  OR2_X1 U11595 ( .A1(n8107), .A2(n11144), .ZN(n11477) );
  XOR2_X1 U11596 ( .A(n11675), .B(n11676), .Z(n11474) );
  XOR2_X1 U11597 ( .A(n11677), .B(n11678), .Z(n11676) );
  OR2_X1 U11598 ( .A1(n8025), .A2(n11144), .ZN(n11481) );
  XOR2_X1 U11599 ( .A(n11679), .B(n11680), .Z(n11478) );
  XOR2_X1 U11600 ( .A(n11681), .B(n11682), .Z(n11680) );
  OR2_X1 U11601 ( .A1(n7955), .A2(n11144), .ZN(n11485) );
  XOR2_X1 U11602 ( .A(n11683), .B(n11684), .Z(n11482) );
  XOR2_X1 U11603 ( .A(n11685), .B(n11686), .Z(n11684) );
  OR2_X1 U11604 ( .A1(n7887), .A2(n11144), .ZN(n11489) );
  XOR2_X1 U11605 ( .A(n11687), .B(n11688), .Z(n11486) );
  XOR2_X1 U11606 ( .A(n11689), .B(n11690), .Z(n11688) );
  OR2_X1 U11607 ( .A1(n7828), .A2(n11144), .ZN(n11493) );
  XOR2_X1 U11608 ( .A(n11691), .B(n11692), .Z(n11490) );
  XOR2_X1 U11609 ( .A(n11693), .B(n11694), .Z(n11692) );
  OR2_X1 U11610 ( .A1(n7820), .A2(n11144), .ZN(n11497) );
  XOR2_X1 U11611 ( .A(n11695), .B(n11696), .Z(n11494) );
  XOR2_X1 U11612 ( .A(n11697), .B(n11698), .Z(n11696) );
  OR2_X1 U11613 ( .A1(n7730), .A2(n11144), .ZN(n11501) );
  XOR2_X1 U11614 ( .A(n11699), .B(n11700), .Z(n11498) );
  XOR2_X1 U11615 ( .A(n11701), .B(n11702), .Z(n11700) );
  XOR2_X1 U11616 ( .A(n11703), .B(n11704), .Z(n11285) );
  XOR2_X1 U11617 ( .A(n11705), .B(n11706), .Z(n11704) );
  OR2_X1 U11618 ( .A1(n8300), .A2(n8299), .ZN(n7574) );
  INV_X1 U11619 ( .A(n11707), .ZN(n8299) );
  OR2_X1 U11620 ( .A1(n11708), .A2(n7587), .ZN(n11707) );
  INV_X1 U11621 ( .A(n7584), .ZN(n7587) );
  OR2_X1 U11622 ( .A1(n11709), .A2(n11710), .ZN(n7584) );
  AND2_X1 U11623 ( .A1(n11709), .A2(n11710), .ZN(n11708) );
  OR2_X1 U11624 ( .A1(n11711), .A2(n11712), .ZN(n11710) );
  AND2_X1 U11625 ( .A1(n11713), .A2(n11714), .ZN(n11712) );
  AND2_X1 U11626 ( .A1(n11715), .A2(n11716), .ZN(n11711) );
  OR2_X1 U11627 ( .A1(n11713), .A2(n11714), .ZN(n11716) );
  XOR2_X1 U11628 ( .A(n8213), .B(n11717), .Z(n11709) );
  XOR2_X1 U11629 ( .A(n8212), .B(n8211), .Z(n11717) );
  OR2_X1 U11630 ( .A1(n7660), .A2(n11718), .ZN(n8211) );
  OR2_X1 U11631 ( .A1(n11719), .A2(n11720), .ZN(n8212) );
  AND2_X1 U11632 ( .A1(n11721), .A2(n11722), .ZN(n11720) );
  AND2_X1 U11633 ( .A1(n11723), .A2(n11724), .ZN(n11719) );
  OR2_X1 U11634 ( .A1(n11722), .A2(n11721), .ZN(n11724) );
  XOR2_X1 U11635 ( .A(n8221), .B(n11725), .Z(n8213) );
  XOR2_X1 U11636 ( .A(n8220), .B(n8219), .Z(n11725) );
  OR2_X1 U11637 ( .A1(n7697), .A2(n8216), .ZN(n8219) );
  OR2_X1 U11638 ( .A1(n11726), .A2(n11727), .ZN(n8220) );
  AND2_X1 U11639 ( .A1(n11728), .A2(n11729), .ZN(n11727) );
  AND2_X1 U11640 ( .A1(n11730), .A2(n11731), .ZN(n11726) );
  OR2_X1 U11641 ( .A1(n11728), .A2(n11729), .ZN(n11731) );
  XOR2_X1 U11642 ( .A(n8228), .B(n11732), .Z(n8221) );
  XOR2_X1 U11643 ( .A(n8227), .B(n8226), .Z(n11732) );
  OR2_X1 U11644 ( .A1(n7730), .A2(n8133), .ZN(n8226) );
  OR2_X1 U11645 ( .A1(n11733), .A2(n11734), .ZN(n8227) );
  AND2_X1 U11646 ( .A1(n11735), .A2(n11736), .ZN(n11734) );
  AND2_X1 U11647 ( .A1(n11737), .A2(n11738), .ZN(n11733) );
  OR2_X1 U11648 ( .A1(n11736), .A2(n11735), .ZN(n11738) );
  XOR2_X1 U11649 ( .A(n8235), .B(n11739), .Z(n8228) );
  XOR2_X1 U11650 ( .A(n8234), .B(n8233), .Z(n11739) );
  OR2_X1 U11651 ( .A1(n8050), .A2(n7820), .ZN(n8233) );
  OR2_X1 U11652 ( .A1(n11740), .A2(n11741), .ZN(n8234) );
  AND2_X1 U11653 ( .A1(n11742), .A2(n11743), .ZN(n11741) );
  AND2_X1 U11654 ( .A1(n11744), .A2(n11745), .ZN(n11740) );
  OR2_X1 U11655 ( .A1(n11742), .A2(n11743), .ZN(n11745) );
  XOR2_X1 U11656 ( .A(n8242), .B(n11746), .Z(n8235) );
  XOR2_X1 U11657 ( .A(n8241), .B(n8240), .Z(n11746) );
  OR2_X1 U11658 ( .A1(n7981), .A2(n7828), .ZN(n8240) );
  OR2_X1 U11659 ( .A1(n11747), .A2(n11748), .ZN(n8241) );
  AND2_X1 U11660 ( .A1(n11749), .A2(n11750), .ZN(n11748) );
  AND2_X1 U11661 ( .A1(n11751), .A2(n11752), .ZN(n11747) );
  OR2_X1 U11662 ( .A1(n11750), .A2(n11749), .ZN(n11752) );
  XOR2_X1 U11663 ( .A(n8249), .B(n11753), .Z(n8242) );
  XOR2_X1 U11664 ( .A(n8248), .B(n8247), .Z(n11753) );
  OR2_X1 U11665 ( .A1(n7912), .A2(n7887), .ZN(n8247) );
  OR2_X1 U11666 ( .A1(n11754), .A2(n11755), .ZN(n8248) );
  AND2_X1 U11667 ( .A1(n11756), .A2(n11757), .ZN(n11755) );
  AND2_X1 U11668 ( .A1(n11758), .A2(n11759), .ZN(n11754) );
  OR2_X1 U11669 ( .A1(n11757), .A2(n11756), .ZN(n11759) );
  XOR2_X1 U11670 ( .A(n8256), .B(n11760), .Z(n8249) );
  XOR2_X1 U11671 ( .A(n8255), .B(n8254), .Z(n11760) );
  OR2_X1 U11672 ( .A1(n7857), .A2(n7955), .ZN(n8254) );
  OR2_X1 U11673 ( .A1(n11761), .A2(n11762), .ZN(n8255) );
  AND2_X1 U11674 ( .A1(n11763), .A2(n11764), .ZN(n11762) );
  AND2_X1 U11675 ( .A1(n11765), .A2(n11766), .ZN(n11761) );
  OR2_X1 U11676 ( .A1(n11764), .A2(n11763), .ZN(n11766) );
  XNOR2_X1 U11677 ( .A(n11767), .B(n8261), .ZN(n8256) );
  XOR2_X1 U11678 ( .A(n8270), .B(n11768), .Z(n8261) );
  XOR2_X1 U11679 ( .A(n8269), .B(n8268), .Z(n11768) );
  OR2_X1 U11680 ( .A1(n7759), .A2(n8107), .ZN(n8268) );
  OR2_X1 U11681 ( .A1(n11769), .A2(n11770), .ZN(n8269) );
  AND2_X1 U11682 ( .A1(n11771), .A2(n11772), .ZN(n11770) );
  AND2_X1 U11683 ( .A1(n11773), .A2(n11774), .ZN(n11769) );
  OR2_X1 U11684 ( .A1(n11772), .A2(n11771), .ZN(n11774) );
  XOR2_X1 U11685 ( .A(n8277), .B(n11775), .Z(n8270) );
  XOR2_X1 U11686 ( .A(n8276), .B(n8275), .Z(n11775) );
  OR2_X1 U11687 ( .A1(n7715), .A2(n8191), .ZN(n8275) );
  OR2_X1 U11688 ( .A1(n11776), .A2(n11777), .ZN(n8276) );
  AND2_X1 U11689 ( .A1(n11778), .A2(n11779), .ZN(n11777) );
  AND2_X1 U11690 ( .A1(n11780), .A2(n11781), .ZN(n11776) );
  OR2_X1 U11691 ( .A1(n11779), .A2(n11778), .ZN(n11781) );
  XOR2_X1 U11692 ( .A(n8284), .B(n11782), .Z(n8277) );
  XOR2_X1 U11693 ( .A(n8283), .B(n8282), .Z(n11782) );
  OR2_X1 U11694 ( .A1(n7689), .A2(n8287), .ZN(n8282) );
  OR2_X1 U11695 ( .A1(n11783), .A2(n11784), .ZN(n8283) );
  AND2_X1 U11696 ( .A1(n11785), .A2(n11786), .ZN(n11784) );
  AND2_X1 U11697 ( .A1(n11787), .A2(n11788), .ZN(n11783) );
  OR2_X1 U11698 ( .A1(n11786), .A2(n11785), .ZN(n11788) );
  XOR2_X1 U11699 ( .A(n8292), .B(n11789), .Z(n8284) );
  XOR2_X1 U11700 ( .A(n8291), .B(n8290), .Z(n11789) );
  OR2_X1 U11701 ( .A1(n8608), .A2(n7659), .ZN(n8290) );
  OR2_X1 U11702 ( .A1(n11790), .A2(n11791), .ZN(n8291) );
  AND2_X1 U11703 ( .A1(n11792), .A2(n11793), .ZN(n11791) );
  AND2_X1 U11704 ( .A1(n11794), .A2(n11795), .ZN(n11790) );
  OR2_X1 U11705 ( .A1(n11793), .A2(n11792), .ZN(n11795) );
  XOR2_X1 U11706 ( .A(n11796), .B(n11797), .Z(n8292) );
  XOR2_X1 U11707 ( .A(n11798), .B(n11799), .Z(n11797) );
  XNOR2_X1 U11708 ( .A(n8264), .B(n8262), .ZN(n11767) );
  OR2_X1 U11709 ( .A1(n11800), .A2(n11801), .ZN(n8262) );
  AND2_X1 U11710 ( .A1(n11802), .A2(n11803), .ZN(n11801) );
  AND2_X1 U11711 ( .A1(n11804), .A2(n11805), .ZN(n11800) );
  OR2_X1 U11712 ( .A1(n11803), .A2(n11802), .ZN(n11805) );
  AND2_X1 U11713 ( .A1(n8304), .A2(n11806), .ZN(n8300) );
  INV_X1 U11714 ( .A(n8305), .ZN(n11806) );
  OR2_X1 U11715 ( .A1(n11807), .A2(n11808), .ZN(n8305) );
  AND2_X1 U11716 ( .A1(n11272), .A2(n11271), .ZN(n11808) );
  AND2_X1 U11717 ( .A1(n11269), .A2(n11809), .ZN(n11807) );
  OR2_X1 U11718 ( .A1(n11271), .A2(n11272), .ZN(n11809) );
  OR2_X1 U11719 ( .A1(n7660), .A2(n11391), .ZN(n11272) );
  OR2_X1 U11720 ( .A1(n11810), .A2(n11811), .ZN(n11271) );
  AND2_X1 U11721 ( .A1(n11290), .A2(n11289), .ZN(n11811) );
  AND2_X1 U11722 ( .A1(n11287), .A2(n11812), .ZN(n11810) );
  OR2_X1 U11723 ( .A1(n11289), .A2(n11290), .ZN(n11812) );
  OR2_X1 U11724 ( .A1(n7697), .A2(n11391), .ZN(n11290) );
  OR2_X1 U11725 ( .A1(n11813), .A2(n11814), .ZN(n11289) );
  AND2_X1 U11726 ( .A1(n11706), .A2(n11705), .ZN(n11814) );
  AND2_X1 U11727 ( .A1(n11703), .A2(n11815), .ZN(n11813) );
  OR2_X1 U11728 ( .A1(n11705), .A2(n11706), .ZN(n11815) );
  OR2_X1 U11729 ( .A1(n7730), .A2(n11391), .ZN(n11706) );
  OR2_X1 U11730 ( .A1(n11816), .A2(n11817), .ZN(n11705) );
  AND2_X1 U11731 ( .A1(n11702), .A2(n11701), .ZN(n11817) );
  AND2_X1 U11732 ( .A1(n11699), .A2(n11818), .ZN(n11816) );
  OR2_X1 U11733 ( .A1(n11701), .A2(n11702), .ZN(n11818) );
  OR2_X1 U11734 ( .A1(n7820), .A2(n11391), .ZN(n11702) );
  OR2_X1 U11735 ( .A1(n11819), .A2(n11820), .ZN(n11701) );
  AND2_X1 U11736 ( .A1(n11698), .A2(n11697), .ZN(n11820) );
  AND2_X1 U11737 ( .A1(n11695), .A2(n11821), .ZN(n11819) );
  OR2_X1 U11738 ( .A1(n11697), .A2(n11698), .ZN(n11821) );
  OR2_X1 U11739 ( .A1(n7828), .A2(n11391), .ZN(n11698) );
  OR2_X1 U11740 ( .A1(n11822), .A2(n11823), .ZN(n11697) );
  AND2_X1 U11741 ( .A1(n11694), .A2(n11693), .ZN(n11823) );
  AND2_X1 U11742 ( .A1(n11691), .A2(n11824), .ZN(n11822) );
  OR2_X1 U11743 ( .A1(n11693), .A2(n11694), .ZN(n11824) );
  OR2_X1 U11744 ( .A1(n7887), .A2(n11391), .ZN(n11694) );
  OR2_X1 U11745 ( .A1(n11825), .A2(n11826), .ZN(n11693) );
  AND2_X1 U11746 ( .A1(n11690), .A2(n11689), .ZN(n11826) );
  AND2_X1 U11747 ( .A1(n11687), .A2(n11827), .ZN(n11825) );
  OR2_X1 U11748 ( .A1(n11689), .A2(n11690), .ZN(n11827) );
  OR2_X1 U11749 ( .A1(n7955), .A2(n11391), .ZN(n11690) );
  OR2_X1 U11750 ( .A1(n11828), .A2(n11829), .ZN(n11689) );
  AND2_X1 U11751 ( .A1(n11686), .A2(n11685), .ZN(n11829) );
  AND2_X1 U11752 ( .A1(n11683), .A2(n11830), .ZN(n11828) );
  OR2_X1 U11753 ( .A1(n11685), .A2(n11686), .ZN(n11830) );
  OR2_X1 U11754 ( .A1(n8025), .A2(n11391), .ZN(n11686) );
  OR2_X1 U11755 ( .A1(n11831), .A2(n11832), .ZN(n11685) );
  AND2_X1 U11756 ( .A1(n11682), .A2(n11681), .ZN(n11832) );
  AND2_X1 U11757 ( .A1(n11679), .A2(n11833), .ZN(n11831) );
  OR2_X1 U11758 ( .A1(n11681), .A2(n11682), .ZN(n11833) );
  OR2_X1 U11759 ( .A1(n8107), .A2(n11391), .ZN(n11682) );
  OR2_X1 U11760 ( .A1(n11834), .A2(n11835), .ZN(n11681) );
  AND2_X1 U11761 ( .A1(n11678), .A2(n11677), .ZN(n11835) );
  AND2_X1 U11762 ( .A1(n11675), .A2(n11836), .ZN(n11834) );
  OR2_X1 U11763 ( .A1(n11677), .A2(n11678), .ZN(n11836) );
  OR2_X1 U11764 ( .A1(n8191), .A2(n11391), .ZN(n11678) );
  OR2_X1 U11765 ( .A1(n11837), .A2(n11838), .ZN(n11677) );
  AND2_X1 U11766 ( .A1(n11674), .A2(n11673), .ZN(n11838) );
  AND2_X1 U11767 ( .A1(n11671), .A2(n11839), .ZN(n11837) );
  OR2_X1 U11768 ( .A1(n11673), .A2(n11674), .ZN(n11839) );
  OR2_X1 U11769 ( .A1(n8287), .A2(n11391), .ZN(n11674) );
  OR2_X1 U11770 ( .A1(n11840), .A2(n11841), .ZN(n11673) );
  AND2_X1 U11771 ( .A1(n11670), .A2(n11669), .ZN(n11841) );
  AND2_X1 U11772 ( .A1(n11667), .A2(n11842), .ZN(n11840) );
  OR2_X1 U11773 ( .A1(n11669), .A2(n11670), .ZN(n11842) );
  OR2_X1 U11774 ( .A1(n8608), .A2(n11391), .ZN(n11670) );
  OR2_X1 U11775 ( .A1(n11843), .A2(n11844), .ZN(n11669) );
  AND2_X1 U11776 ( .A1(n11666), .A2(n11665), .ZN(n11844) );
  AND2_X1 U11777 ( .A1(n11663), .A2(n11845), .ZN(n11843) );
  OR2_X1 U11778 ( .A1(n11665), .A2(n11666), .ZN(n11845) );
  OR2_X1 U11779 ( .A1(n8603), .A2(n11391), .ZN(n11666) );
  OR2_X1 U11780 ( .A1(n11846), .A2(n11847), .ZN(n11665) );
  AND2_X1 U11781 ( .A1(n11662), .A2(n11661), .ZN(n11847) );
  AND2_X1 U11782 ( .A1(n11659), .A2(n11848), .ZN(n11846) );
  OR2_X1 U11783 ( .A1(n11661), .A2(n11662), .ZN(n11848) );
  OR2_X1 U11784 ( .A1(n8598), .A2(n11391), .ZN(n11662) );
  OR2_X1 U11785 ( .A1(n11849), .A2(n11850), .ZN(n11661) );
  AND2_X1 U11786 ( .A1(n11658), .A2(n11657), .ZN(n11850) );
  AND2_X1 U11787 ( .A1(n11655), .A2(n11851), .ZN(n11849) );
  OR2_X1 U11788 ( .A1(n11657), .A2(n11658), .ZN(n11851) );
  OR2_X1 U11789 ( .A1(n8593), .A2(n11391), .ZN(n11658) );
  OR2_X1 U11790 ( .A1(n11852), .A2(n11853), .ZN(n11657) );
  AND2_X1 U11791 ( .A1(n11654), .A2(n11653), .ZN(n11853) );
  AND2_X1 U11792 ( .A1(n11651), .A2(n11854), .ZN(n11852) );
  OR2_X1 U11793 ( .A1(n11653), .A2(n11654), .ZN(n11854) );
  OR2_X1 U11794 ( .A1(n8588), .A2(n11391), .ZN(n11654) );
  OR2_X1 U11795 ( .A1(n11855), .A2(n11856), .ZN(n11653) );
  AND2_X1 U11796 ( .A1(n11648), .A2(n11650), .ZN(n11856) );
  AND2_X1 U11797 ( .A1(n11857), .A2(n11649), .ZN(n11855) );
  OR2_X1 U11798 ( .A1(n11650), .A2(n11648), .ZN(n11857) );
  XOR2_X1 U11799 ( .A(n11858), .B(n11859), .Z(n11648) );
  XOR2_X1 U11800 ( .A(n11860), .B(n11861), .Z(n11859) );
  OR2_X1 U11801 ( .A1(n11862), .A2(n11863), .ZN(n11650) );
  AND2_X1 U11802 ( .A1(n11646), .A2(n11645), .ZN(n11863) );
  AND2_X1 U11803 ( .A1(n11643), .A2(n11864), .ZN(n11862) );
  OR2_X1 U11804 ( .A1(n11645), .A2(n11646), .ZN(n11864) );
  OR2_X1 U11805 ( .A1(n8578), .A2(n11391), .ZN(n11646) );
  OR2_X1 U11806 ( .A1(n11865), .A2(n11866), .ZN(n11645) );
  AND2_X1 U11807 ( .A1(n11642), .A2(n11641), .ZN(n11866) );
  AND2_X1 U11808 ( .A1(n11639), .A2(n11867), .ZN(n11865) );
  OR2_X1 U11809 ( .A1(n11641), .A2(n11642), .ZN(n11867) );
  OR2_X1 U11810 ( .A1(n8573), .A2(n11391), .ZN(n11642) );
  OR2_X1 U11811 ( .A1(n11868), .A2(n11869), .ZN(n11641) );
  AND2_X1 U11812 ( .A1(n11638), .A2(n11637), .ZN(n11869) );
  AND2_X1 U11813 ( .A1(n11635), .A2(n11870), .ZN(n11868) );
  OR2_X1 U11814 ( .A1(n11637), .A2(n11638), .ZN(n11870) );
  OR2_X1 U11815 ( .A1(n8568), .A2(n11391), .ZN(n11638) );
  OR2_X1 U11816 ( .A1(n11871), .A2(n11872), .ZN(n11637) );
  AND2_X1 U11817 ( .A1(n11634), .A2(n11633), .ZN(n11872) );
  AND2_X1 U11818 ( .A1(n11631), .A2(n11873), .ZN(n11871) );
  OR2_X1 U11819 ( .A1(n11633), .A2(n11634), .ZN(n11873) );
  OR2_X1 U11820 ( .A1(n8563), .A2(n11391), .ZN(n11634) );
  OR2_X1 U11821 ( .A1(n11874), .A2(n11875), .ZN(n11633) );
  AND2_X1 U11822 ( .A1(n11630), .A2(n11629), .ZN(n11875) );
  AND2_X1 U11823 ( .A1(n11627), .A2(n11876), .ZN(n11874) );
  OR2_X1 U11824 ( .A1(n11629), .A2(n11630), .ZN(n11876) );
  OR2_X1 U11825 ( .A1(n8558), .A2(n11391), .ZN(n11630) );
  OR2_X1 U11826 ( .A1(n11877), .A2(n11878), .ZN(n11629) );
  AND2_X1 U11827 ( .A1(n11626), .A2(n11625), .ZN(n11878) );
  AND2_X1 U11828 ( .A1(n11623), .A2(n11879), .ZN(n11877) );
  OR2_X1 U11829 ( .A1(n11625), .A2(n11626), .ZN(n11879) );
  OR2_X1 U11830 ( .A1(n8553), .A2(n11391), .ZN(n11626) );
  OR2_X1 U11831 ( .A1(n11880), .A2(n11881), .ZN(n11625) );
  AND2_X1 U11832 ( .A1(n11622), .A2(n11621), .ZN(n11881) );
  AND2_X1 U11833 ( .A1(n11619), .A2(n11882), .ZN(n11880) );
  OR2_X1 U11834 ( .A1(n11621), .A2(n11622), .ZN(n11882) );
  OR2_X1 U11835 ( .A1(n8548), .A2(n11391), .ZN(n11622) );
  OR2_X1 U11836 ( .A1(n11883), .A2(n11884), .ZN(n11621) );
  AND2_X1 U11837 ( .A1(n11618), .A2(n11617), .ZN(n11884) );
  AND2_X1 U11838 ( .A1(n11615), .A2(n11885), .ZN(n11883) );
  OR2_X1 U11839 ( .A1(n11617), .A2(n11618), .ZN(n11885) );
  OR2_X1 U11840 ( .A1(n8543), .A2(n11391), .ZN(n11618) );
  OR2_X1 U11841 ( .A1(n11886), .A2(n11887), .ZN(n11617) );
  AND2_X1 U11842 ( .A1(n11614), .A2(n11613), .ZN(n11887) );
  AND2_X1 U11843 ( .A1(n11611), .A2(n11888), .ZN(n11886) );
  OR2_X1 U11844 ( .A1(n11613), .A2(n11614), .ZN(n11888) );
  OR2_X1 U11845 ( .A1(n8538), .A2(n11391), .ZN(n11614) );
  OR2_X1 U11846 ( .A1(n11889), .A2(n11890), .ZN(n11613) );
  AND2_X1 U11847 ( .A1(n11610), .A2(n11609), .ZN(n11890) );
  AND2_X1 U11848 ( .A1(n11607), .A2(n11891), .ZN(n11889) );
  OR2_X1 U11849 ( .A1(n11609), .A2(n11610), .ZN(n11891) );
  OR2_X1 U11850 ( .A1(n8533), .A2(n11391), .ZN(n11610) );
  OR2_X1 U11851 ( .A1(n11892), .A2(n11893), .ZN(n11609) );
  AND2_X1 U11852 ( .A1(n11606), .A2(n11605), .ZN(n11893) );
  AND2_X1 U11853 ( .A1(n11603), .A2(n11894), .ZN(n11892) );
  OR2_X1 U11854 ( .A1(n11605), .A2(n11606), .ZN(n11894) );
  OR2_X1 U11855 ( .A1(n8528), .A2(n11391), .ZN(n11606) );
  OR2_X1 U11856 ( .A1(n11895), .A2(n11896), .ZN(n11605) );
  AND2_X1 U11857 ( .A1(n11602), .A2(n11601), .ZN(n11896) );
  AND2_X1 U11858 ( .A1(n11599), .A2(n11897), .ZN(n11895) );
  OR2_X1 U11859 ( .A1(n11601), .A2(n11602), .ZN(n11897) );
  OR2_X1 U11860 ( .A1(n8523), .A2(n11391), .ZN(n11602) );
  OR2_X1 U11861 ( .A1(n11898), .A2(n11899), .ZN(n11601) );
  AND2_X1 U11862 ( .A1(n11596), .A2(n11597), .ZN(n11899) );
  AND2_X1 U11863 ( .A1(n11900), .A2(n11901), .ZN(n11898) );
  OR2_X1 U11864 ( .A1(n11597), .A2(n11596), .ZN(n11901) );
  OR2_X1 U11865 ( .A1(n8515), .A2(n11391), .ZN(n11596) );
  OR2_X1 U11866 ( .A1(n11391), .A2(n11902), .ZN(n11597) );
  INV_X1 U11867 ( .A(n11598), .ZN(n11900) );
  OR2_X1 U11868 ( .A1(n11903), .A2(n11904), .ZN(n11598) );
  AND2_X1 U11869 ( .A1(b_15_), .A2(n11905), .ZN(n11904) );
  OR2_X1 U11870 ( .A1(n11906), .A2(n7343), .ZN(n11905) );
  AND2_X1 U11871 ( .A1(a_30_), .A2(n11718), .ZN(n11906) );
  AND2_X1 U11872 ( .A1(b_14_), .A2(n11907), .ZN(n11903) );
  OR2_X1 U11873 ( .A1(n11908), .A2(n7347), .ZN(n11907) );
  AND2_X1 U11874 ( .A1(a_31_), .A2(n11592), .ZN(n11908) );
  XOR2_X1 U11875 ( .A(n11909), .B(n11910), .Z(n11599) );
  XNOR2_X1 U11876 ( .A(n11911), .B(n11912), .ZN(n11909) );
  XOR2_X1 U11877 ( .A(n11913), .B(n11914), .Z(n11603) );
  XOR2_X1 U11878 ( .A(n11915), .B(n11916), .Z(n11914) );
  XOR2_X1 U11879 ( .A(n11917), .B(n11918), .Z(n11607) );
  XOR2_X1 U11880 ( .A(n11919), .B(n11920), .Z(n11918) );
  XOR2_X1 U11881 ( .A(n11921), .B(n11922), .Z(n11611) );
  XOR2_X1 U11882 ( .A(n11923), .B(n11924), .Z(n11922) );
  XOR2_X1 U11883 ( .A(n11925), .B(n11926), .Z(n11615) );
  XOR2_X1 U11884 ( .A(n11927), .B(n11928), .Z(n11926) );
  XOR2_X1 U11885 ( .A(n11929), .B(n11930), .Z(n11619) );
  XOR2_X1 U11886 ( .A(n11931), .B(n11932), .Z(n11930) );
  XOR2_X1 U11887 ( .A(n11933), .B(n11934), .Z(n11623) );
  XOR2_X1 U11888 ( .A(n11935), .B(n11936), .Z(n11934) );
  XOR2_X1 U11889 ( .A(n11937), .B(n11938), .Z(n11627) );
  XOR2_X1 U11890 ( .A(n11939), .B(n11940), .Z(n11938) );
  XOR2_X1 U11891 ( .A(n11941), .B(n11942), .Z(n11631) );
  XOR2_X1 U11892 ( .A(n11943), .B(n11944), .Z(n11942) );
  XOR2_X1 U11893 ( .A(n11945), .B(n11946), .Z(n11635) );
  XOR2_X1 U11894 ( .A(n11947), .B(n11948), .Z(n11946) );
  XOR2_X1 U11895 ( .A(n11949), .B(n11950), .Z(n11639) );
  XOR2_X1 U11896 ( .A(n11951), .B(n11952), .Z(n11950) );
  XOR2_X1 U11897 ( .A(n11953), .B(n11954), .Z(n11643) );
  XOR2_X1 U11898 ( .A(n11955), .B(n11956), .Z(n11954) );
  XOR2_X1 U11899 ( .A(n11957), .B(n11958), .Z(n11651) );
  XOR2_X1 U11900 ( .A(n11959), .B(n11960), .Z(n11958) );
  XNOR2_X1 U11901 ( .A(n11961), .B(n11962), .ZN(n11655) );
  XNOR2_X1 U11902 ( .A(n11963), .B(n11964), .ZN(n11961) );
  XOR2_X1 U11903 ( .A(n11965), .B(n11966), .Z(n11659) );
  XOR2_X1 U11904 ( .A(n11967), .B(n11968), .Z(n11966) );
  XOR2_X1 U11905 ( .A(n11969), .B(n11970), .Z(n11663) );
  XOR2_X1 U11906 ( .A(n11971), .B(n11972), .Z(n11970) );
  XOR2_X1 U11907 ( .A(n11973), .B(n11974), .Z(n11667) );
  XOR2_X1 U11908 ( .A(n11975), .B(n11976), .Z(n11974) );
  XOR2_X1 U11909 ( .A(n11977), .B(n11978), .Z(n11671) );
  XOR2_X1 U11910 ( .A(n11979), .B(n11980), .Z(n11978) );
  XOR2_X1 U11911 ( .A(n11981), .B(n11982), .Z(n11675) );
  XOR2_X1 U11912 ( .A(n11983), .B(n11984), .Z(n11982) );
  XOR2_X1 U11913 ( .A(n11985), .B(n11986), .Z(n11679) );
  XOR2_X1 U11914 ( .A(n11987), .B(n11988), .Z(n11986) );
  XOR2_X1 U11915 ( .A(n11989), .B(n11990), .Z(n11683) );
  XOR2_X1 U11916 ( .A(n11991), .B(n11992), .Z(n11990) );
  XOR2_X1 U11917 ( .A(n11993), .B(n11994), .Z(n11687) );
  XOR2_X1 U11918 ( .A(n11995), .B(n11996), .Z(n11994) );
  XOR2_X1 U11919 ( .A(n11997), .B(n11998), .Z(n11691) );
  XOR2_X1 U11920 ( .A(n11999), .B(n12000), .Z(n11998) );
  XOR2_X1 U11921 ( .A(n12001), .B(n12002), .Z(n11695) );
  XOR2_X1 U11922 ( .A(n12003), .B(n12004), .Z(n12002) );
  XOR2_X1 U11923 ( .A(n12005), .B(n12006), .Z(n11699) );
  XOR2_X1 U11924 ( .A(n12007), .B(n12008), .Z(n12006) );
  XOR2_X1 U11925 ( .A(n12009), .B(n12010), .Z(n11703) );
  XOR2_X1 U11926 ( .A(n12011), .B(n12012), .Z(n12010) );
  XOR2_X1 U11927 ( .A(n12013), .B(n12014), .Z(n11287) );
  XOR2_X1 U11928 ( .A(n12015), .B(n12016), .Z(n12014) );
  XOR2_X1 U11929 ( .A(n12017), .B(n12018), .Z(n11269) );
  XOR2_X1 U11930 ( .A(n12019), .B(n12020), .Z(n12018) );
  XNOR2_X1 U11931 ( .A(n11715), .B(n12021), .ZN(n8304) );
  XOR2_X1 U11932 ( .A(n11714), .B(n11713), .Z(n12021) );
  OR2_X1 U11933 ( .A1(n7660), .A2(n11592), .ZN(n11713) );
  OR2_X1 U11934 ( .A1(n12022), .A2(n12023), .ZN(n11714) );
  AND2_X1 U11935 ( .A1(n12020), .A2(n12019), .ZN(n12023) );
  AND2_X1 U11936 ( .A1(n12017), .A2(n12024), .ZN(n12022) );
  OR2_X1 U11937 ( .A1(n12020), .A2(n12019), .ZN(n12024) );
  OR2_X1 U11938 ( .A1(n12025), .A2(n12026), .ZN(n12019) );
  AND2_X1 U11939 ( .A1(n12016), .A2(n12015), .ZN(n12026) );
  AND2_X1 U11940 ( .A1(n12013), .A2(n12027), .ZN(n12025) );
  OR2_X1 U11941 ( .A1(n12016), .A2(n12015), .ZN(n12027) );
  OR2_X1 U11942 ( .A1(n12028), .A2(n12029), .ZN(n12015) );
  AND2_X1 U11943 ( .A1(n12012), .A2(n12011), .ZN(n12029) );
  AND2_X1 U11944 ( .A1(n12009), .A2(n12030), .ZN(n12028) );
  OR2_X1 U11945 ( .A1(n12012), .A2(n12011), .ZN(n12030) );
  OR2_X1 U11946 ( .A1(n12031), .A2(n12032), .ZN(n12011) );
  AND2_X1 U11947 ( .A1(n12008), .A2(n12007), .ZN(n12032) );
  AND2_X1 U11948 ( .A1(n12005), .A2(n12033), .ZN(n12031) );
  OR2_X1 U11949 ( .A1(n12008), .A2(n12007), .ZN(n12033) );
  OR2_X1 U11950 ( .A1(n12034), .A2(n12035), .ZN(n12007) );
  AND2_X1 U11951 ( .A1(n12004), .A2(n12003), .ZN(n12035) );
  AND2_X1 U11952 ( .A1(n12001), .A2(n12036), .ZN(n12034) );
  OR2_X1 U11953 ( .A1(n12004), .A2(n12003), .ZN(n12036) );
  OR2_X1 U11954 ( .A1(n12037), .A2(n12038), .ZN(n12003) );
  AND2_X1 U11955 ( .A1(n12000), .A2(n11999), .ZN(n12038) );
  AND2_X1 U11956 ( .A1(n11997), .A2(n12039), .ZN(n12037) );
  OR2_X1 U11957 ( .A1(n12000), .A2(n11999), .ZN(n12039) );
  OR2_X1 U11958 ( .A1(n12040), .A2(n12041), .ZN(n11999) );
  AND2_X1 U11959 ( .A1(n11996), .A2(n11995), .ZN(n12041) );
  AND2_X1 U11960 ( .A1(n11993), .A2(n12042), .ZN(n12040) );
  OR2_X1 U11961 ( .A1(n11996), .A2(n11995), .ZN(n12042) );
  OR2_X1 U11962 ( .A1(n12043), .A2(n12044), .ZN(n11995) );
  AND2_X1 U11963 ( .A1(n11992), .A2(n11991), .ZN(n12044) );
  AND2_X1 U11964 ( .A1(n11989), .A2(n12045), .ZN(n12043) );
  OR2_X1 U11965 ( .A1(n11992), .A2(n11991), .ZN(n12045) );
  OR2_X1 U11966 ( .A1(n12046), .A2(n12047), .ZN(n11991) );
  AND2_X1 U11967 ( .A1(n11988), .A2(n11987), .ZN(n12047) );
  AND2_X1 U11968 ( .A1(n11985), .A2(n12048), .ZN(n12046) );
  OR2_X1 U11969 ( .A1(n11988), .A2(n11987), .ZN(n12048) );
  OR2_X1 U11970 ( .A1(n12049), .A2(n12050), .ZN(n11987) );
  AND2_X1 U11971 ( .A1(n11984), .A2(n11983), .ZN(n12050) );
  AND2_X1 U11972 ( .A1(n11981), .A2(n12051), .ZN(n12049) );
  OR2_X1 U11973 ( .A1(n11984), .A2(n11983), .ZN(n12051) );
  OR2_X1 U11974 ( .A1(n12052), .A2(n12053), .ZN(n11983) );
  AND2_X1 U11975 ( .A1(n11980), .A2(n11979), .ZN(n12053) );
  AND2_X1 U11976 ( .A1(n11977), .A2(n12054), .ZN(n12052) );
  OR2_X1 U11977 ( .A1(n11980), .A2(n11979), .ZN(n12054) );
  OR2_X1 U11978 ( .A1(n12055), .A2(n12056), .ZN(n11979) );
  AND2_X1 U11979 ( .A1(n11976), .A2(n11975), .ZN(n12056) );
  AND2_X1 U11980 ( .A1(n11973), .A2(n12057), .ZN(n12055) );
  OR2_X1 U11981 ( .A1(n11976), .A2(n11975), .ZN(n12057) );
  OR2_X1 U11982 ( .A1(n12058), .A2(n12059), .ZN(n11975) );
  AND2_X1 U11983 ( .A1(n11972), .A2(n11971), .ZN(n12059) );
  AND2_X1 U11984 ( .A1(n11969), .A2(n12060), .ZN(n12058) );
  OR2_X1 U11985 ( .A1(n11972), .A2(n11971), .ZN(n12060) );
  OR2_X1 U11986 ( .A1(n12061), .A2(n12062), .ZN(n11971) );
  AND2_X1 U11987 ( .A1(n11968), .A2(n11967), .ZN(n12062) );
  AND2_X1 U11988 ( .A1(n11965), .A2(n12063), .ZN(n12061) );
  OR2_X1 U11989 ( .A1(n11968), .A2(n11967), .ZN(n12063) );
  OR2_X1 U11990 ( .A1(n12064), .A2(n12065), .ZN(n11967) );
  AND2_X1 U11991 ( .A1(n11962), .A2(n11964), .ZN(n12065) );
  AND2_X1 U11992 ( .A1(n12066), .A2(n11963), .ZN(n12064) );
  OR2_X1 U11993 ( .A1(n11962), .A2(n11964), .ZN(n12066) );
  OR2_X1 U11994 ( .A1(n12067), .A2(n12068), .ZN(n11964) );
  AND2_X1 U11995 ( .A1(n11960), .A2(n11959), .ZN(n12068) );
  AND2_X1 U11996 ( .A1(n11957), .A2(n12069), .ZN(n12067) );
  OR2_X1 U11997 ( .A1(n11960), .A2(n11959), .ZN(n12069) );
  OR2_X1 U11998 ( .A1(n12070), .A2(n12071), .ZN(n11959) );
  AND2_X1 U11999 ( .A1(n11861), .A2(n11860), .ZN(n12071) );
  AND2_X1 U12000 ( .A1(n11858), .A2(n12072), .ZN(n12070) );
  OR2_X1 U12001 ( .A1(n11861), .A2(n11860), .ZN(n12072) );
  OR2_X1 U12002 ( .A1(n12073), .A2(n12074), .ZN(n11860) );
  AND2_X1 U12003 ( .A1(n11956), .A2(n11955), .ZN(n12074) );
  AND2_X1 U12004 ( .A1(n11953), .A2(n12075), .ZN(n12073) );
  OR2_X1 U12005 ( .A1(n11956), .A2(n11955), .ZN(n12075) );
  OR2_X1 U12006 ( .A1(n12076), .A2(n12077), .ZN(n11955) );
  AND2_X1 U12007 ( .A1(n11952), .A2(n11951), .ZN(n12077) );
  AND2_X1 U12008 ( .A1(n11949), .A2(n12078), .ZN(n12076) );
  OR2_X1 U12009 ( .A1(n11952), .A2(n11951), .ZN(n12078) );
  OR2_X1 U12010 ( .A1(n12079), .A2(n12080), .ZN(n11951) );
  AND2_X1 U12011 ( .A1(n11948), .A2(n11947), .ZN(n12080) );
  AND2_X1 U12012 ( .A1(n11945), .A2(n12081), .ZN(n12079) );
  OR2_X1 U12013 ( .A1(n11948), .A2(n11947), .ZN(n12081) );
  OR2_X1 U12014 ( .A1(n12082), .A2(n12083), .ZN(n11947) );
  AND2_X1 U12015 ( .A1(n11944), .A2(n11943), .ZN(n12083) );
  AND2_X1 U12016 ( .A1(n11941), .A2(n12084), .ZN(n12082) );
  OR2_X1 U12017 ( .A1(n11944), .A2(n11943), .ZN(n12084) );
  OR2_X1 U12018 ( .A1(n12085), .A2(n12086), .ZN(n11943) );
  AND2_X1 U12019 ( .A1(n11940), .A2(n11939), .ZN(n12086) );
  AND2_X1 U12020 ( .A1(n11937), .A2(n12087), .ZN(n12085) );
  OR2_X1 U12021 ( .A1(n11940), .A2(n11939), .ZN(n12087) );
  OR2_X1 U12022 ( .A1(n12088), .A2(n12089), .ZN(n11939) );
  AND2_X1 U12023 ( .A1(n11936), .A2(n11935), .ZN(n12089) );
  AND2_X1 U12024 ( .A1(n11933), .A2(n12090), .ZN(n12088) );
  OR2_X1 U12025 ( .A1(n11936), .A2(n11935), .ZN(n12090) );
  OR2_X1 U12026 ( .A1(n12091), .A2(n12092), .ZN(n11935) );
  AND2_X1 U12027 ( .A1(n11932), .A2(n11931), .ZN(n12092) );
  AND2_X1 U12028 ( .A1(n11929), .A2(n12093), .ZN(n12091) );
  OR2_X1 U12029 ( .A1(n11932), .A2(n11931), .ZN(n12093) );
  OR2_X1 U12030 ( .A1(n12094), .A2(n12095), .ZN(n11931) );
  AND2_X1 U12031 ( .A1(n11928), .A2(n11927), .ZN(n12095) );
  AND2_X1 U12032 ( .A1(n11925), .A2(n12096), .ZN(n12094) );
  OR2_X1 U12033 ( .A1(n11928), .A2(n11927), .ZN(n12096) );
  OR2_X1 U12034 ( .A1(n12097), .A2(n12098), .ZN(n11927) );
  AND2_X1 U12035 ( .A1(n11924), .A2(n11923), .ZN(n12098) );
  AND2_X1 U12036 ( .A1(n11921), .A2(n12099), .ZN(n12097) );
  OR2_X1 U12037 ( .A1(n11924), .A2(n11923), .ZN(n12099) );
  OR2_X1 U12038 ( .A1(n12100), .A2(n12101), .ZN(n11923) );
  AND2_X1 U12039 ( .A1(n11920), .A2(n11919), .ZN(n12101) );
  AND2_X1 U12040 ( .A1(n11917), .A2(n12102), .ZN(n12100) );
  OR2_X1 U12041 ( .A1(n11920), .A2(n11919), .ZN(n12102) );
  OR2_X1 U12042 ( .A1(n12103), .A2(n12104), .ZN(n11919) );
  AND2_X1 U12043 ( .A1(n11916), .A2(n11915), .ZN(n12104) );
  AND2_X1 U12044 ( .A1(n11913), .A2(n12105), .ZN(n12103) );
  OR2_X1 U12045 ( .A1(n11916), .A2(n11915), .ZN(n12105) );
  OR2_X1 U12046 ( .A1(n12106), .A2(n12107), .ZN(n11915) );
  AND2_X1 U12047 ( .A1(n11910), .A2(n11911), .ZN(n12107) );
  AND2_X1 U12048 ( .A1(n12108), .A2(n12109), .ZN(n12106) );
  OR2_X1 U12049 ( .A1(n11910), .A2(n11911), .ZN(n12109) );
  OR2_X1 U12050 ( .A1(n11718), .A2(n11902), .ZN(n11911) );
  OR2_X1 U12051 ( .A1(n8956), .A2(n11592), .ZN(n11902) );
  OR2_X1 U12052 ( .A1(n8515), .A2(n11592), .ZN(n11910) );
  INV_X1 U12053 ( .A(n11912), .ZN(n12108) );
  OR2_X1 U12054 ( .A1(n12110), .A2(n12111), .ZN(n11912) );
  AND2_X1 U12055 ( .A1(b_14_), .A2(n12112), .ZN(n12111) );
  OR2_X1 U12056 ( .A1(n12113), .A2(n7343), .ZN(n12112) );
  AND2_X1 U12057 ( .A1(a_30_), .A2(n8216), .ZN(n12113) );
  AND2_X1 U12058 ( .A1(b_13_), .A2(n12114), .ZN(n12110) );
  OR2_X1 U12059 ( .A1(n12115), .A2(n7347), .ZN(n12114) );
  AND2_X1 U12060 ( .A1(a_31_), .A2(n11718), .ZN(n12115) );
  OR2_X1 U12061 ( .A1(n8523), .A2(n11592), .ZN(n11916) );
  XOR2_X1 U12062 ( .A(n12116), .B(n12117), .Z(n11913) );
  XNOR2_X1 U12063 ( .A(n12118), .B(n12119), .ZN(n12116) );
  OR2_X1 U12064 ( .A1(n8528), .A2(n11592), .ZN(n11920) );
  XOR2_X1 U12065 ( .A(n12120), .B(n12121), .Z(n11917) );
  XOR2_X1 U12066 ( .A(n12122), .B(n12123), .Z(n12121) );
  OR2_X1 U12067 ( .A1(n8533), .A2(n11592), .ZN(n11924) );
  XOR2_X1 U12068 ( .A(n12124), .B(n12125), .Z(n11921) );
  XOR2_X1 U12069 ( .A(n12126), .B(n12127), .Z(n12125) );
  OR2_X1 U12070 ( .A1(n8538), .A2(n11592), .ZN(n11928) );
  XOR2_X1 U12071 ( .A(n12128), .B(n12129), .Z(n11925) );
  XOR2_X1 U12072 ( .A(n12130), .B(n12131), .Z(n12129) );
  OR2_X1 U12073 ( .A1(n8543), .A2(n11592), .ZN(n11932) );
  XOR2_X1 U12074 ( .A(n12132), .B(n12133), .Z(n11929) );
  XOR2_X1 U12075 ( .A(n12134), .B(n12135), .Z(n12133) );
  OR2_X1 U12076 ( .A1(n8548), .A2(n11592), .ZN(n11936) );
  XOR2_X1 U12077 ( .A(n12136), .B(n12137), .Z(n11933) );
  XOR2_X1 U12078 ( .A(n12138), .B(n12139), .Z(n12137) );
  OR2_X1 U12079 ( .A1(n8553), .A2(n11592), .ZN(n11940) );
  XOR2_X1 U12080 ( .A(n12140), .B(n12141), .Z(n11937) );
  XOR2_X1 U12081 ( .A(n12142), .B(n12143), .Z(n12141) );
  OR2_X1 U12082 ( .A1(n8558), .A2(n11592), .ZN(n11944) );
  XOR2_X1 U12083 ( .A(n12144), .B(n12145), .Z(n11941) );
  XOR2_X1 U12084 ( .A(n12146), .B(n12147), .Z(n12145) );
  OR2_X1 U12085 ( .A1(n8563), .A2(n11592), .ZN(n11948) );
  XOR2_X1 U12086 ( .A(n12148), .B(n12149), .Z(n11945) );
  XOR2_X1 U12087 ( .A(n12150), .B(n12151), .Z(n12149) );
  OR2_X1 U12088 ( .A1(n8568), .A2(n11592), .ZN(n11952) );
  XOR2_X1 U12089 ( .A(n12152), .B(n12153), .Z(n11949) );
  XOR2_X1 U12090 ( .A(n12154), .B(n12155), .Z(n12153) );
  OR2_X1 U12091 ( .A1(n8573), .A2(n11592), .ZN(n11956) );
  XOR2_X1 U12092 ( .A(n12156), .B(n12157), .Z(n11953) );
  XOR2_X1 U12093 ( .A(n12158), .B(n12159), .Z(n12157) );
  OR2_X1 U12094 ( .A1(n8578), .A2(n11592), .ZN(n11861) );
  XOR2_X1 U12095 ( .A(n12160), .B(n12161), .Z(n11858) );
  XOR2_X1 U12096 ( .A(n12162), .B(n12163), .Z(n12161) );
  OR2_X1 U12097 ( .A1(n8583), .A2(n11592), .ZN(n11960) );
  XOR2_X1 U12098 ( .A(n12164), .B(n12165), .Z(n11957) );
  XOR2_X1 U12099 ( .A(n12166), .B(n12167), .Z(n12165) );
  XOR2_X1 U12100 ( .A(n12168), .B(n12169), .Z(n11962) );
  XOR2_X1 U12101 ( .A(n12170), .B(n12171), .Z(n12169) );
  OR2_X1 U12102 ( .A1(n8593), .A2(n11592), .ZN(n11968) );
  XOR2_X1 U12103 ( .A(n12172), .B(n12173), .Z(n11965) );
  XOR2_X1 U12104 ( .A(n12174), .B(n12175), .Z(n12173) );
  OR2_X1 U12105 ( .A1(n8598), .A2(n11592), .ZN(n11972) );
  XNOR2_X1 U12106 ( .A(n12176), .B(n12177), .ZN(n11969) );
  XNOR2_X1 U12107 ( .A(n12178), .B(n12179), .ZN(n12176) );
  OR2_X1 U12108 ( .A1(n8603), .A2(n11592), .ZN(n11976) );
  XOR2_X1 U12109 ( .A(n12180), .B(n12181), .Z(n11973) );
  XOR2_X1 U12110 ( .A(n12182), .B(n12183), .Z(n12181) );
  OR2_X1 U12111 ( .A1(n8608), .A2(n11592), .ZN(n11980) );
  XOR2_X1 U12112 ( .A(n12184), .B(n12185), .Z(n11977) );
  XOR2_X1 U12113 ( .A(n12186), .B(n12187), .Z(n12185) );
  OR2_X1 U12114 ( .A1(n8287), .A2(n11592), .ZN(n11984) );
  XOR2_X1 U12115 ( .A(n12188), .B(n12189), .Z(n11981) );
  XOR2_X1 U12116 ( .A(n12190), .B(n12191), .Z(n12189) );
  OR2_X1 U12117 ( .A1(n8191), .A2(n11592), .ZN(n11988) );
  XOR2_X1 U12118 ( .A(n12192), .B(n12193), .Z(n11985) );
  XOR2_X1 U12119 ( .A(n12194), .B(n12195), .Z(n12193) );
  OR2_X1 U12120 ( .A1(n8107), .A2(n11592), .ZN(n11992) );
  XOR2_X1 U12121 ( .A(n12196), .B(n12197), .Z(n11989) );
  XOR2_X1 U12122 ( .A(n12198), .B(n12199), .Z(n12197) );
  OR2_X1 U12123 ( .A1(n8025), .A2(n11592), .ZN(n11996) );
  XOR2_X1 U12124 ( .A(n12200), .B(n12201), .Z(n11993) );
  XOR2_X1 U12125 ( .A(n12202), .B(n12203), .Z(n12201) );
  OR2_X1 U12126 ( .A1(n7955), .A2(n11592), .ZN(n12000) );
  XOR2_X1 U12127 ( .A(n12204), .B(n12205), .Z(n11997) );
  XOR2_X1 U12128 ( .A(n12206), .B(n12207), .Z(n12205) );
  OR2_X1 U12129 ( .A1(n7887), .A2(n11592), .ZN(n12004) );
  XOR2_X1 U12130 ( .A(n12208), .B(n12209), .Z(n12001) );
  XOR2_X1 U12131 ( .A(n12210), .B(n12211), .Z(n12209) );
  OR2_X1 U12132 ( .A1(n7828), .A2(n11592), .ZN(n12008) );
  XOR2_X1 U12133 ( .A(n12212), .B(n12213), .Z(n12005) );
  XOR2_X1 U12134 ( .A(n12214), .B(n12215), .Z(n12213) );
  OR2_X1 U12135 ( .A1(n7820), .A2(n11592), .ZN(n12012) );
  XOR2_X1 U12136 ( .A(n12216), .B(n12217), .Z(n12009) );
  XOR2_X1 U12137 ( .A(n12218), .B(n12219), .Z(n12217) );
  OR2_X1 U12138 ( .A1(n7730), .A2(n11592), .ZN(n12016) );
  XOR2_X1 U12139 ( .A(n12220), .B(n12221), .Z(n12013) );
  XOR2_X1 U12140 ( .A(n12222), .B(n12223), .Z(n12221) );
  OR2_X1 U12141 ( .A1(n7697), .A2(n11592), .ZN(n12020) );
  XOR2_X1 U12142 ( .A(n12224), .B(n12225), .Z(n12017) );
  XOR2_X1 U12143 ( .A(n12226), .B(n12227), .Z(n12225) );
  XOR2_X1 U12144 ( .A(n11723), .B(n12228), .Z(n11715) );
  XOR2_X1 U12145 ( .A(n11722), .B(n11721), .Z(n12228) );
  OR2_X1 U12146 ( .A1(n7697), .A2(n11718), .ZN(n11721) );
  OR2_X1 U12147 ( .A1(n12229), .A2(n12230), .ZN(n11722) );
  AND2_X1 U12148 ( .A1(n12227), .A2(n12226), .ZN(n12230) );
  AND2_X1 U12149 ( .A1(n12224), .A2(n12231), .ZN(n12229) );
  OR2_X1 U12150 ( .A1(n12226), .A2(n12227), .ZN(n12231) );
  OR2_X1 U12151 ( .A1(n7730), .A2(n11718), .ZN(n12227) );
  OR2_X1 U12152 ( .A1(n12232), .A2(n12233), .ZN(n12226) );
  AND2_X1 U12153 ( .A1(n12223), .A2(n12222), .ZN(n12233) );
  AND2_X1 U12154 ( .A1(n12220), .A2(n12234), .ZN(n12232) );
  OR2_X1 U12155 ( .A1(n12222), .A2(n12223), .ZN(n12234) );
  OR2_X1 U12156 ( .A1(n7820), .A2(n11718), .ZN(n12223) );
  OR2_X1 U12157 ( .A1(n12235), .A2(n12236), .ZN(n12222) );
  AND2_X1 U12158 ( .A1(n12219), .A2(n12218), .ZN(n12236) );
  AND2_X1 U12159 ( .A1(n12216), .A2(n12237), .ZN(n12235) );
  OR2_X1 U12160 ( .A1(n12218), .A2(n12219), .ZN(n12237) );
  OR2_X1 U12161 ( .A1(n7828), .A2(n11718), .ZN(n12219) );
  OR2_X1 U12162 ( .A1(n12238), .A2(n12239), .ZN(n12218) );
  AND2_X1 U12163 ( .A1(n12215), .A2(n12214), .ZN(n12239) );
  AND2_X1 U12164 ( .A1(n12212), .A2(n12240), .ZN(n12238) );
  OR2_X1 U12165 ( .A1(n12214), .A2(n12215), .ZN(n12240) );
  OR2_X1 U12166 ( .A1(n7887), .A2(n11718), .ZN(n12215) );
  OR2_X1 U12167 ( .A1(n12241), .A2(n12242), .ZN(n12214) );
  AND2_X1 U12168 ( .A1(n12211), .A2(n12210), .ZN(n12242) );
  AND2_X1 U12169 ( .A1(n12208), .A2(n12243), .ZN(n12241) );
  OR2_X1 U12170 ( .A1(n12210), .A2(n12211), .ZN(n12243) );
  OR2_X1 U12171 ( .A1(n7955), .A2(n11718), .ZN(n12211) );
  OR2_X1 U12172 ( .A1(n12244), .A2(n12245), .ZN(n12210) );
  AND2_X1 U12173 ( .A1(n12207), .A2(n12206), .ZN(n12245) );
  AND2_X1 U12174 ( .A1(n12204), .A2(n12246), .ZN(n12244) );
  OR2_X1 U12175 ( .A1(n12206), .A2(n12207), .ZN(n12246) );
  OR2_X1 U12176 ( .A1(n8025), .A2(n11718), .ZN(n12207) );
  OR2_X1 U12177 ( .A1(n12247), .A2(n12248), .ZN(n12206) );
  AND2_X1 U12178 ( .A1(n12203), .A2(n12202), .ZN(n12248) );
  AND2_X1 U12179 ( .A1(n12200), .A2(n12249), .ZN(n12247) );
  OR2_X1 U12180 ( .A1(n12202), .A2(n12203), .ZN(n12249) );
  OR2_X1 U12181 ( .A1(n8107), .A2(n11718), .ZN(n12203) );
  OR2_X1 U12182 ( .A1(n12250), .A2(n12251), .ZN(n12202) );
  AND2_X1 U12183 ( .A1(n12199), .A2(n12198), .ZN(n12251) );
  AND2_X1 U12184 ( .A1(n12196), .A2(n12252), .ZN(n12250) );
  OR2_X1 U12185 ( .A1(n12198), .A2(n12199), .ZN(n12252) );
  OR2_X1 U12186 ( .A1(n8191), .A2(n11718), .ZN(n12199) );
  OR2_X1 U12187 ( .A1(n12253), .A2(n12254), .ZN(n12198) );
  AND2_X1 U12188 ( .A1(n12195), .A2(n12194), .ZN(n12254) );
  AND2_X1 U12189 ( .A1(n12192), .A2(n12255), .ZN(n12253) );
  OR2_X1 U12190 ( .A1(n12194), .A2(n12195), .ZN(n12255) );
  OR2_X1 U12191 ( .A1(n8287), .A2(n11718), .ZN(n12195) );
  OR2_X1 U12192 ( .A1(n12256), .A2(n12257), .ZN(n12194) );
  AND2_X1 U12193 ( .A1(n12191), .A2(n12190), .ZN(n12257) );
  AND2_X1 U12194 ( .A1(n12188), .A2(n12258), .ZN(n12256) );
  OR2_X1 U12195 ( .A1(n12190), .A2(n12191), .ZN(n12258) );
  OR2_X1 U12196 ( .A1(n8608), .A2(n11718), .ZN(n12191) );
  OR2_X1 U12197 ( .A1(n12259), .A2(n12260), .ZN(n12190) );
  AND2_X1 U12198 ( .A1(n12187), .A2(n12186), .ZN(n12260) );
  AND2_X1 U12199 ( .A1(n12184), .A2(n12261), .ZN(n12259) );
  OR2_X1 U12200 ( .A1(n12186), .A2(n12187), .ZN(n12261) );
  OR2_X1 U12201 ( .A1(n8603), .A2(n11718), .ZN(n12187) );
  OR2_X1 U12202 ( .A1(n12262), .A2(n12263), .ZN(n12186) );
  AND2_X1 U12203 ( .A1(n12183), .A2(n12182), .ZN(n12263) );
  AND2_X1 U12204 ( .A1(n12180), .A2(n12264), .ZN(n12262) );
  OR2_X1 U12205 ( .A1(n12182), .A2(n12183), .ZN(n12264) );
  OR2_X1 U12206 ( .A1(n8598), .A2(n11718), .ZN(n12183) );
  OR2_X1 U12207 ( .A1(n12265), .A2(n12266), .ZN(n12182) );
  AND2_X1 U12208 ( .A1(n12177), .A2(n12179), .ZN(n12266) );
  AND2_X1 U12209 ( .A1(n12267), .A2(n12178), .ZN(n12265) );
  OR2_X1 U12210 ( .A1(n12177), .A2(n12179), .ZN(n12267) );
  OR2_X1 U12211 ( .A1(n12268), .A2(n12269), .ZN(n12179) );
  AND2_X1 U12212 ( .A1(n12175), .A2(n12174), .ZN(n12269) );
  AND2_X1 U12213 ( .A1(n12172), .A2(n12270), .ZN(n12268) );
  OR2_X1 U12214 ( .A1(n12174), .A2(n12175), .ZN(n12270) );
  OR2_X1 U12215 ( .A1(n8588), .A2(n11718), .ZN(n12175) );
  OR2_X1 U12216 ( .A1(n12271), .A2(n12272), .ZN(n12174) );
  AND2_X1 U12217 ( .A1(n12171), .A2(n12170), .ZN(n12272) );
  AND2_X1 U12218 ( .A1(n12168), .A2(n12273), .ZN(n12271) );
  OR2_X1 U12219 ( .A1(n12170), .A2(n12171), .ZN(n12273) );
  OR2_X1 U12220 ( .A1(n8583), .A2(n11718), .ZN(n12171) );
  OR2_X1 U12221 ( .A1(n12274), .A2(n12275), .ZN(n12170) );
  AND2_X1 U12222 ( .A1(n12167), .A2(n12166), .ZN(n12275) );
  AND2_X1 U12223 ( .A1(n12164), .A2(n12276), .ZN(n12274) );
  OR2_X1 U12224 ( .A1(n12166), .A2(n12167), .ZN(n12276) );
  OR2_X1 U12225 ( .A1(n8578), .A2(n11718), .ZN(n12167) );
  OR2_X1 U12226 ( .A1(n12277), .A2(n12278), .ZN(n12166) );
  AND2_X1 U12227 ( .A1(n12163), .A2(n12162), .ZN(n12278) );
  AND2_X1 U12228 ( .A1(n12160), .A2(n12279), .ZN(n12277) );
  OR2_X1 U12229 ( .A1(n12162), .A2(n12163), .ZN(n12279) );
  OR2_X1 U12230 ( .A1(n8573), .A2(n11718), .ZN(n12163) );
  OR2_X1 U12231 ( .A1(n12280), .A2(n12281), .ZN(n12162) );
  AND2_X1 U12232 ( .A1(n12159), .A2(n12158), .ZN(n12281) );
  AND2_X1 U12233 ( .A1(n12156), .A2(n12282), .ZN(n12280) );
  OR2_X1 U12234 ( .A1(n12158), .A2(n12159), .ZN(n12282) );
  OR2_X1 U12235 ( .A1(n8568), .A2(n11718), .ZN(n12159) );
  OR2_X1 U12236 ( .A1(n12283), .A2(n12284), .ZN(n12158) );
  AND2_X1 U12237 ( .A1(n12155), .A2(n12154), .ZN(n12284) );
  AND2_X1 U12238 ( .A1(n12152), .A2(n12285), .ZN(n12283) );
  OR2_X1 U12239 ( .A1(n12154), .A2(n12155), .ZN(n12285) );
  OR2_X1 U12240 ( .A1(n8563), .A2(n11718), .ZN(n12155) );
  OR2_X1 U12241 ( .A1(n12286), .A2(n12287), .ZN(n12154) );
  AND2_X1 U12242 ( .A1(n12151), .A2(n12150), .ZN(n12287) );
  AND2_X1 U12243 ( .A1(n12148), .A2(n12288), .ZN(n12286) );
  OR2_X1 U12244 ( .A1(n12150), .A2(n12151), .ZN(n12288) );
  OR2_X1 U12245 ( .A1(n8558), .A2(n11718), .ZN(n12151) );
  OR2_X1 U12246 ( .A1(n12289), .A2(n12290), .ZN(n12150) );
  AND2_X1 U12247 ( .A1(n12147), .A2(n12146), .ZN(n12290) );
  AND2_X1 U12248 ( .A1(n12144), .A2(n12291), .ZN(n12289) );
  OR2_X1 U12249 ( .A1(n12146), .A2(n12147), .ZN(n12291) );
  OR2_X1 U12250 ( .A1(n8553), .A2(n11718), .ZN(n12147) );
  OR2_X1 U12251 ( .A1(n12292), .A2(n12293), .ZN(n12146) );
  AND2_X1 U12252 ( .A1(n12143), .A2(n12142), .ZN(n12293) );
  AND2_X1 U12253 ( .A1(n12140), .A2(n12294), .ZN(n12292) );
  OR2_X1 U12254 ( .A1(n12142), .A2(n12143), .ZN(n12294) );
  OR2_X1 U12255 ( .A1(n8548), .A2(n11718), .ZN(n12143) );
  OR2_X1 U12256 ( .A1(n12295), .A2(n12296), .ZN(n12142) );
  AND2_X1 U12257 ( .A1(n12139), .A2(n12138), .ZN(n12296) );
  AND2_X1 U12258 ( .A1(n12136), .A2(n12297), .ZN(n12295) );
  OR2_X1 U12259 ( .A1(n12138), .A2(n12139), .ZN(n12297) );
  OR2_X1 U12260 ( .A1(n8543), .A2(n11718), .ZN(n12139) );
  OR2_X1 U12261 ( .A1(n12298), .A2(n12299), .ZN(n12138) );
  AND2_X1 U12262 ( .A1(n12135), .A2(n12134), .ZN(n12299) );
  AND2_X1 U12263 ( .A1(n12132), .A2(n12300), .ZN(n12298) );
  OR2_X1 U12264 ( .A1(n12134), .A2(n12135), .ZN(n12300) );
  OR2_X1 U12265 ( .A1(n8538), .A2(n11718), .ZN(n12135) );
  OR2_X1 U12266 ( .A1(n12301), .A2(n12302), .ZN(n12134) );
  AND2_X1 U12267 ( .A1(n12131), .A2(n12130), .ZN(n12302) );
  AND2_X1 U12268 ( .A1(n12128), .A2(n12303), .ZN(n12301) );
  OR2_X1 U12269 ( .A1(n12130), .A2(n12131), .ZN(n12303) );
  OR2_X1 U12270 ( .A1(n8533), .A2(n11718), .ZN(n12131) );
  OR2_X1 U12271 ( .A1(n12304), .A2(n12305), .ZN(n12130) );
  AND2_X1 U12272 ( .A1(n12127), .A2(n12126), .ZN(n12305) );
  AND2_X1 U12273 ( .A1(n12124), .A2(n12306), .ZN(n12304) );
  OR2_X1 U12274 ( .A1(n12126), .A2(n12127), .ZN(n12306) );
  OR2_X1 U12275 ( .A1(n8528), .A2(n11718), .ZN(n12127) );
  OR2_X1 U12276 ( .A1(n12307), .A2(n12308), .ZN(n12126) );
  AND2_X1 U12277 ( .A1(n12123), .A2(n12122), .ZN(n12308) );
  AND2_X1 U12278 ( .A1(n12120), .A2(n12309), .ZN(n12307) );
  OR2_X1 U12279 ( .A1(n12122), .A2(n12123), .ZN(n12309) );
  OR2_X1 U12280 ( .A1(n8523), .A2(n11718), .ZN(n12123) );
  OR2_X1 U12281 ( .A1(n12310), .A2(n12311), .ZN(n12122) );
  AND2_X1 U12282 ( .A1(n12117), .A2(n12118), .ZN(n12311) );
  AND2_X1 U12283 ( .A1(n12312), .A2(n12313), .ZN(n12310) );
  OR2_X1 U12284 ( .A1(n12118), .A2(n12117), .ZN(n12313) );
  OR2_X1 U12285 ( .A1(n8515), .A2(n11718), .ZN(n12117) );
  OR2_X1 U12286 ( .A1(n11718), .A2(n12314), .ZN(n12118) );
  INV_X1 U12287 ( .A(n12119), .ZN(n12312) );
  OR2_X1 U12288 ( .A1(n12315), .A2(n12316), .ZN(n12119) );
  AND2_X1 U12289 ( .A1(b_13_), .A2(n12317), .ZN(n12316) );
  OR2_X1 U12290 ( .A1(n12318), .A2(n7343), .ZN(n12317) );
  AND2_X1 U12291 ( .A1(a_30_), .A2(n8133), .ZN(n12318) );
  AND2_X1 U12292 ( .A1(b_12_), .A2(n12319), .ZN(n12315) );
  OR2_X1 U12293 ( .A1(n12320), .A2(n7347), .ZN(n12319) );
  AND2_X1 U12294 ( .A1(a_31_), .A2(n8216), .ZN(n12320) );
  XOR2_X1 U12295 ( .A(n12321), .B(n12322), .Z(n12120) );
  XNOR2_X1 U12296 ( .A(n12323), .B(n12324), .ZN(n12321) );
  XOR2_X1 U12297 ( .A(n12325), .B(n12326), .Z(n12124) );
  XOR2_X1 U12298 ( .A(n12327), .B(n12328), .Z(n12326) );
  XOR2_X1 U12299 ( .A(n12329), .B(n12330), .Z(n12128) );
  XOR2_X1 U12300 ( .A(n12331), .B(n12332), .Z(n12330) );
  XOR2_X1 U12301 ( .A(n12333), .B(n12334), .Z(n12132) );
  XOR2_X1 U12302 ( .A(n12335), .B(n12336), .Z(n12334) );
  XOR2_X1 U12303 ( .A(n12337), .B(n12338), .Z(n12136) );
  XOR2_X1 U12304 ( .A(n12339), .B(n12340), .Z(n12338) );
  XOR2_X1 U12305 ( .A(n12341), .B(n12342), .Z(n12140) );
  XOR2_X1 U12306 ( .A(n12343), .B(n12344), .Z(n12342) );
  XOR2_X1 U12307 ( .A(n12345), .B(n12346), .Z(n12144) );
  XOR2_X1 U12308 ( .A(n12347), .B(n12348), .Z(n12346) );
  XOR2_X1 U12309 ( .A(n12349), .B(n12350), .Z(n12148) );
  XOR2_X1 U12310 ( .A(n12351), .B(n12352), .Z(n12350) );
  XOR2_X1 U12311 ( .A(n12353), .B(n12354), .Z(n12152) );
  XOR2_X1 U12312 ( .A(n12355), .B(n12356), .Z(n12354) );
  XOR2_X1 U12313 ( .A(n12357), .B(n12358), .Z(n12156) );
  XOR2_X1 U12314 ( .A(n12359), .B(n12360), .Z(n12358) );
  XOR2_X1 U12315 ( .A(n12361), .B(n12362), .Z(n12160) );
  XOR2_X1 U12316 ( .A(n12363), .B(n12364), .Z(n12362) );
  XOR2_X1 U12317 ( .A(n12365), .B(n12366), .Z(n12164) );
  XOR2_X1 U12318 ( .A(n12367), .B(n12368), .Z(n12366) );
  XOR2_X1 U12319 ( .A(n12369), .B(n12370), .Z(n12168) );
  XOR2_X1 U12320 ( .A(n12371), .B(n12372), .Z(n12370) );
  XOR2_X1 U12321 ( .A(n12373), .B(n12374), .Z(n12172) );
  XOR2_X1 U12322 ( .A(n12375), .B(n12376), .Z(n12374) );
  XOR2_X1 U12323 ( .A(n12377), .B(n12378), .Z(n12177) );
  XOR2_X1 U12324 ( .A(n12379), .B(n12380), .Z(n12378) );
  XOR2_X1 U12325 ( .A(n12381), .B(n12382), .Z(n12180) );
  XOR2_X1 U12326 ( .A(n12383), .B(n12384), .Z(n12382) );
  XNOR2_X1 U12327 ( .A(n12385), .B(n12386), .ZN(n12184) );
  XNOR2_X1 U12328 ( .A(n12387), .B(n12388), .ZN(n12385) );
  XOR2_X1 U12329 ( .A(n12389), .B(n12390), .Z(n12188) );
  XOR2_X1 U12330 ( .A(n12391), .B(n12392), .Z(n12390) );
  XOR2_X1 U12331 ( .A(n12393), .B(n12394), .Z(n12192) );
  XOR2_X1 U12332 ( .A(n12395), .B(n12396), .Z(n12394) );
  XOR2_X1 U12333 ( .A(n12397), .B(n12398), .Z(n12196) );
  XOR2_X1 U12334 ( .A(n12399), .B(n12400), .Z(n12398) );
  XOR2_X1 U12335 ( .A(n12401), .B(n12402), .Z(n12200) );
  XOR2_X1 U12336 ( .A(n12403), .B(n12404), .Z(n12402) );
  XOR2_X1 U12337 ( .A(n12405), .B(n12406), .Z(n12204) );
  XOR2_X1 U12338 ( .A(n12407), .B(n12408), .Z(n12406) );
  XOR2_X1 U12339 ( .A(n12409), .B(n12410), .Z(n12208) );
  XOR2_X1 U12340 ( .A(n12411), .B(n12412), .Z(n12410) );
  XOR2_X1 U12341 ( .A(n12413), .B(n12414), .Z(n12212) );
  XOR2_X1 U12342 ( .A(n12415), .B(n12416), .Z(n12414) );
  XOR2_X1 U12343 ( .A(n12417), .B(n12418), .Z(n12216) );
  XOR2_X1 U12344 ( .A(n12419), .B(n12420), .Z(n12418) );
  XOR2_X1 U12345 ( .A(n12421), .B(n12422), .Z(n12220) );
  XOR2_X1 U12346 ( .A(n12423), .B(n12424), .Z(n12422) );
  XOR2_X1 U12347 ( .A(n12425), .B(n12426), .Z(n12224) );
  XOR2_X1 U12348 ( .A(n12427), .B(n12428), .Z(n12426) );
  XOR2_X1 U12349 ( .A(n11730), .B(n12429), .Z(n11723) );
  XOR2_X1 U12350 ( .A(n11729), .B(n11728), .Z(n12429) );
  OR2_X1 U12351 ( .A1(n7730), .A2(n8216), .ZN(n11728) );
  OR2_X1 U12352 ( .A1(n12430), .A2(n12431), .ZN(n11729) );
  AND2_X1 U12353 ( .A1(n12428), .A2(n12427), .ZN(n12431) );
  AND2_X1 U12354 ( .A1(n12425), .A2(n12432), .ZN(n12430) );
  OR2_X1 U12355 ( .A1(n12428), .A2(n12427), .ZN(n12432) );
  OR2_X1 U12356 ( .A1(n12433), .A2(n12434), .ZN(n12427) );
  AND2_X1 U12357 ( .A1(n12424), .A2(n12423), .ZN(n12434) );
  AND2_X1 U12358 ( .A1(n12421), .A2(n12435), .ZN(n12433) );
  OR2_X1 U12359 ( .A1(n12424), .A2(n12423), .ZN(n12435) );
  OR2_X1 U12360 ( .A1(n12436), .A2(n12437), .ZN(n12423) );
  AND2_X1 U12361 ( .A1(n12420), .A2(n12419), .ZN(n12437) );
  AND2_X1 U12362 ( .A1(n12417), .A2(n12438), .ZN(n12436) );
  OR2_X1 U12363 ( .A1(n12420), .A2(n12419), .ZN(n12438) );
  OR2_X1 U12364 ( .A1(n12439), .A2(n12440), .ZN(n12419) );
  AND2_X1 U12365 ( .A1(n12416), .A2(n12415), .ZN(n12440) );
  AND2_X1 U12366 ( .A1(n12413), .A2(n12441), .ZN(n12439) );
  OR2_X1 U12367 ( .A1(n12416), .A2(n12415), .ZN(n12441) );
  OR2_X1 U12368 ( .A1(n12442), .A2(n12443), .ZN(n12415) );
  AND2_X1 U12369 ( .A1(n12412), .A2(n12411), .ZN(n12443) );
  AND2_X1 U12370 ( .A1(n12409), .A2(n12444), .ZN(n12442) );
  OR2_X1 U12371 ( .A1(n12412), .A2(n12411), .ZN(n12444) );
  OR2_X1 U12372 ( .A1(n12445), .A2(n12446), .ZN(n12411) );
  AND2_X1 U12373 ( .A1(n12408), .A2(n12407), .ZN(n12446) );
  AND2_X1 U12374 ( .A1(n12405), .A2(n12447), .ZN(n12445) );
  OR2_X1 U12375 ( .A1(n12408), .A2(n12407), .ZN(n12447) );
  OR2_X1 U12376 ( .A1(n12448), .A2(n12449), .ZN(n12407) );
  AND2_X1 U12377 ( .A1(n12404), .A2(n12403), .ZN(n12449) );
  AND2_X1 U12378 ( .A1(n12401), .A2(n12450), .ZN(n12448) );
  OR2_X1 U12379 ( .A1(n12404), .A2(n12403), .ZN(n12450) );
  OR2_X1 U12380 ( .A1(n12451), .A2(n12452), .ZN(n12403) );
  AND2_X1 U12381 ( .A1(n12400), .A2(n12399), .ZN(n12452) );
  AND2_X1 U12382 ( .A1(n12397), .A2(n12453), .ZN(n12451) );
  OR2_X1 U12383 ( .A1(n12400), .A2(n12399), .ZN(n12453) );
  OR2_X1 U12384 ( .A1(n12454), .A2(n12455), .ZN(n12399) );
  AND2_X1 U12385 ( .A1(n12396), .A2(n12395), .ZN(n12455) );
  AND2_X1 U12386 ( .A1(n12393), .A2(n12456), .ZN(n12454) );
  OR2_X1 U12387 ( .A1(n12396), .A2(n12395), .ZN(n12456) );
  OR2_X1 U12388 ( .A1(n12457), .A2(n12458), .ZN(n12395) );
  AND2_X1 U12389 ( .A1(n12392), .A2(n12391), .ZN(n12458) );
  AND2_X1 U12390 ( .A1(n12389), .A2(n12459), .ZN(n12457) );
  OR2_X1 U12391 ( .A1(n12392), .A2(n12391), .ZN(n12459) );
  OR2_X1 U12392 ( .A1(n12460), .A2(n12461), .ZN(n12391) );
  AND2_X1 U12393 ( .A1(n12386), .A2(n12388), .ZN(n12461) );
  AND2_X1 U12394 ( .A1(n12462), .A2(n12387), .ZN(n12460) );
  OR2_X1 U12395 ( .A1(n12386), .A2(n12388), .ZN(n12462) );
  OR2_X1 U12396 ( .A1(n12463), .A2(n12464), .ZN(n12388) );
  AND2_X1 U12397 ( .A1(n12384), .A2(n12383), .ZN(n12464) );
  AND2_X1 U12398 ( .A1(n12381), .A2(n12465), .ZN(n12463) );
  OR2_X1 U12399 ( .A1(n12384), .A2(n12383), .ZN(n12465) );
  OR2_X1 U12400 ( .A1(n12466), .A2(n12467), .ZN(n12383) );
  AND2_X1 U12401 ( .A1(n12380), .A2(n12379), .ZN(n12467) );
  AND2_X1 U12402 ( .A1(n12377), .A2(n12468), .ZN(n12466) );
  OR2_X1 U12403 ( .A1(n12380), .A2(n12379), .ZN(n12468) );
  OR2_X1 U12404 ( .A1(n12469), .A2(n12470), .ZN(n12379) );
  AND2_X1 U12405 ( .A1(n12376), .A2(n12375), .ZN(n12470) );
  AND2_X1 U12406 ( .A1(n12373), .A2(n12471), .ZN(n12469) );
  OR2_X1 U12407 ( .A1(n12376), .A2(n12375), .ZN(n12471) );
  OR2_X1 U12408 ( .A1(n12472), .A2(n12473), .ZN(n12375) );
  AND2_X1 U12409 ( .A1(n12372), .A2(n12371), .ZN(n12473) );
  AND2_X1 U12410 ( .A1(n12369), .A2(n12474), .ZN(n12472) );
  OR2_X1 U12411 ( .A1(n12372), .A2(n12371), .ZN(n12474) );
  OR2_X1 U12412 ( .A1(n12475), .A2(n12476), .ZN(n12371) );
  AND2_X1 U12413 ( .A1(n12368), .A2(n12367), .ZN(n12476) );
  AND2_X1 U12414 ( .A1(n12365), .A2(n12477), .ZN(n12475) );
  OR2_X1 U12415 ( .A1(n12368), .A2(n12367), .ZN(n12477) );
  OR2_X1 U12416 ( .A1(n12478), .A2(n12479), .ZN(n12367) );
  AND2_X1 U12417 ( .A1(n12364), .A2(n12363), .ZN(n12479) );
  AND2_X1 U12418 ( .A1(n12361), .A2(n12480), .ZN(n12478) );
  OR2_X1 U12419 ( .A1(n12364), .A2(n12363), .ZN(n12480) );
  OR2_X1 U12420 ( .A1(n12481), .A2(n12482), .ZN(n12363) );
  AND2_X1 U12421 ( .A1(n12360), .A2(n12359), .ZN(n12482) );
  AND2_X1 U12422 ( .A1(n12357), .A2(n12483), .ZN(n12481) );
  OR2_X1 U12423 ( .A1(n12360), .A2(n12359), .ZN(n12483) );
  OR2_X1 U12424 ( .A1(n12484), .A2(n12485), .ZN(n12359) );
  AND2_X1 U12425 ( .A1(n12356), .A2(n12355), .ZN(n12485) );
  AND2_X1 U12426 ( .A1(n12353), .A2(n12486), .ZN(n12484) );
  OR2_X1 U12427 ( .A1(n12356), .A2(n12355), .ZN(n12486) );
  OR2_X1 U12428 ( .A1(n12487), .A2(n12488), .ZN(n12355) );
  AND2_X1 U12429 ( .A1(n12352), .A2(n12351), .ZN(n12488) );
  AND2_X1 U12430 ( .A1(n12349), .A2(n12489), .ZN(n12487) );
  OR2_X1 U12431 ( .A1(n12352), .A2(n12351), .ZN(n12489) );
  OR2_X1 U12432 ( .A1(n12490), .A2(n12491), .ZN(n12351) );
  AND2_X1 U12433 ( .A1(n12348), .A2(n12347), .ZN(n12491) );
  AND2_X1 U12434 ( .A1(n12345), .A2(n12492), .ZN(n12490) );
  OR2_X1 U12435 ( .A1(n12348), .A2(n12347), .ZN(n12492) );
  OR2_X1 U12436 ( .A1(n12493), .A2(n12494), .ZN(n12347) );
  AND2_X1 U12437 ( .A1(n12344), .A2(n12343), .ZN(n12494) );
  AND2_X1 U12438 ( .A1(n12341), .A2(n12495), .ZN(n12493) );
  OR2_X1 U12439 ( .A1(n12344), .A2(n12343), .ZN(n12495) );
  OR2_X1 U12440 ( .A1(n12496), .A2(n12497), .ZN(n12343) );
  AND2_X1 U12441 ( .A1(n12340), .A2(n12339), .ZN(n12497) );
  AND2_X1 U12442 ( .A1(n12337), .A2(n12498), .ZN(n12496) );
  OR2_X1 U12443 ( .A1(n12340), .A2(n12339), .ZN(n12498) );
  OR2_X1 U12444 ( .A1(n12499), .A2(n12500), .ZN(n12339) );
  AND2_X1 U12445 ( .A1(n12336), .A2(n12335), .ZN(n12500) );
  AND2_X1 U12446 ( .A1(n12333), .A2(n12501), .ZN(n12499) );
  OR2_X1 U12447 ( .A1(n12336), .A2(n12335), .ZN(n12501) );
  OR2_X1 U12448 ( .A1(n12502), .A2(n12503), .ZN(n12335) );
  AND2_X1 U12449 ( .A1(n12332), .A2(n12331), .ZN(n12503) );
  AND2_X1 U12450 ( .A1(n12329), .A2(n12504), .ZN(n12502) );
  OR2_X1 U12451 ( .A1(n12332), .A2(n12331), .ZN(n12504) );
  OR2_X1 U12452 ( .A1(n12505), .A2(n12506), .ZN(n12331) );
  AND2_X1 U12453 ( .A1(n12328), .A2(n12327), .ZN(n12506) );
  AND2_X1 U12454 ( .A1(n12325), .A2(n12507), .ZN(n12505) );
  OR2_X1 U12455 ( .A1(n12328), .A2(n12327), .ZN(n12507) );
  OR2_X1 U12456 ( .A1(n12508), .A2(n12509), .ZN(n12327) );
  AND2_X1 U12457 ( .A1(n12322), .A2(n12323), .ZN(n12509) );
  AND2_X1 U12458 ( .A1(n12510), .A2(n12511), .ZN(n12508) );
  OR2_X1 U12459 ( .A1(n12322), .A2(n12323), .ZN(n12511) );
  OR2_X1 U12460 ( .A1(n8133), .A2(n12314), .ZN(n12323) );
  OR2_X1 U12461 ( .A1(n8956), .A2(n8216), .ZN(n12314) );
  OR2_X1 U12462 ( .A1(n8515), .A2(n8216), .ZN(n12322) );
  INV_X1 U12463 ( .A(n12324), .ZN(n12510) );
  OR2_X1 U12464 ( .A1(n12512), .A2(n12513), .ZN(n12324) );
  AND2_X1 U12465 ( .A1(b_12_), .A2(n12514), .ZN(n12513) );
  OR2_X1 U12466 ( .A1(n12515), .A2(n7343), .ZN(n12514) );
  AND2_X1 U12467 ( .A1(a_30_), .A2(n8050), .ZN(n12515) );
  AND2_X1 U12468 ( .A1(b_11_), .A2(n12516), .ZN(n12512) );
  OR2_X1 U12469 ( .A1(n12517), .A2(n7347), .ZN(n12516) );
  AND2_X1 U12470 ( .A1(a_31_), .A2(n8133), .ZN(n12517) );
  OR2_X1 U12471 ( .A1(n8523), .A2(n8216), .ZN(n12328) );
  XOR2_X1 U12472 ( .A(n12518), .B(n12519), .Z(n12325) );
  XNOR2_X1 U12473 ( .A(n12520), .B(n12521), .ZN(n12518) );
  OR2_X1 U12474 ( .A1(n8528), .A2(n8216), .ZN(n12332) );
  XOR2_X1 U12475 ( .A(n12522), .B(n12523), .Z(n12329) );
  XOR2_X1 U12476 ( .A(n12524), .B(n12525), .Z(n12523) );
  OR2_X1 U12477 ( .A1(n8533), .A2(n8216), .ZN(n12336) );
  XOR2_X1 U12478 ( .A(n12526), .B(n12527), .Z(n12333) );
  XOR2_X1 U12479 ( .A(n12528), .B(n12529), .Z(n12527) );
  OR2_X1 U12480 ( .A1(n8538), .A2(n8216), .ZN(n12340) );
  XOR2_X1 U12481 ( .A(n12530), .B(n12531), .Z(n12337) );
  XOR2_X1 U12482 ( .A(n12532), .B(n12533), .Z(n12531) );
  OR2_X1 U12483 ( .A1(n8543), .A2(n8216), .ZN(n12344) );
  XOR2_X1 U12484 ( .A(n12534), .B(n12535), .Z(n12341) );
  XOR2_X1 U12485 ( .A(n12536), .B(n12537), .Z(n12535) );
  OR2_X1 U12486 ( .A1(n8548), .A2(n8216), .ZN(n12348) );
  XOR2_X1 U12487 ( .A(n12538), .B(n12539), .Z(n12345) );
  XOR2_X1 U12488 ( .A(n12540), .B(n12541), .Z(n12539) );
  OR2_X1 U12489 ( .A1(n8553), .A2(n8216), .ZN(n12352) );
  XOR2_X1 U12490 ( .A(n12542), .B(n12543), .Z(n12349) );
  XOR2_X1 U12491 ( .A(n12544), .B(n12545), .Z(n12543) );
  OR2_X1 U12492 ( .A1(n8558), .A2(n8216), .ZN(n12356) );
  XOR2_X1 U12493 ( .A(n12546), .B(n12547), .Z(n12353) );
  XOR2_X1 U12494 ( .A(n12548), .B(n12549), .Z(n12547) );
  OR2_X1 U12495 ( .A1(n8563), .A2(n8216), .ZN(n12360) );
  XOR2_X1 U12496 ( .A(n12550), .B(n12551), .Z(n12357) );
  XOR2_X1 U12497 ( .A(n12552), .B(n12553), .Z(n12551) );
  OR2_X1 U12498 ( .A1(n8568), .A2(n8216), .ZN(n12364) );
  XOR2_X1 U12499 ( .A(n12554), .B(n12555), .Z(n12361) );
  XOR2_X1 U12500 ( .A(n12556), .B(n12557), .Z(n12555) );
  OR2_X1 U12501 ( .A1(n8573), .A2(n8216), .ZN(n12368) );
  XOR2_X1 U12502 ( .A(n12558), .B(n12559), .Z(n12365) );
  XOR2_X1 U12503 ( .A(n12560), .B(n12561), .Z(n12559) );
  OR2_X1 U12504 ( .A1(n8578), .A2(n8216), .ZN(n12372) );
  XOR2_X1 U12505 ( .A(n12562), .B(n12563), .Z(n12369) );
  XOR2_X1 U12506 ( .A(n12564), .B(n12565), .Z(n12563) );
  OR2_X1 U12507 ( .A1(n8583), .A2(n8216), .ZN(n12376) );
  XOR2_X1 U12508 ( .A(n12566), .B(n12567), .Z(n12373) );
  XOR2_X1 U12509 ( .A(n12568), .B(n12569), .Z(n12567) );
  OR2_X1 U12510 ( .A1(n8588), .A2(n8216), .ZN(n12380) );
  XOR2_X1 U12511 ( .A(n12570), .B(n12571), .Z(n12377) );
  XOR2_X1 U12512 ( .A(n12572), .B(n12573), .Z(n12571) );
  OR2_X1 U12513 ( .A1(n8593), .A2(n8216), .ZN(n12384) );
  XOR2_X1 U12514 ( .A(n12574), .B(n12575), .Z(n12381) );
  XOR2_X1 U12515 ( .A(n12576), .B(n12577), .Z(n12575) );
  XOR2_X1 U12516 ( .A(n12578), .B(n12579), .Z(n12386) );
  XOR2_X1 U12517 ( .A(n12580), .B(n12581), .Z(n12579) );
  OR2_X1 U12518 ( .A1(n8603), .A2(n8216), .ZN(n12392) );
  XOR2_X1 U12519 ( .A(n12582), .B(n12583), .Z(n12389) );
  XOR2_X1 U12520 ( .A(n12584), .B(n12585), .Z(n12583) );
  OR2_X1 U12521 ( .A1(n8608), .A2(n8216), .ZN(n12396) );
  XNOR2_X1 U12522 ( .A(n12586), .B(n12587), .ZN(n12393) );
  XNOR2_X1 U12523 ( .A(n12588), .B(n12589), .ZN(n12586) );
  OR2_X1 U12524 ( .A1(n8287), .A2(n8216), .ZN(n12400) );
  XOR2_X1 U12525 ( .A(n12590), .B(n12591), .Z(n12397) );
  XOR2_X1 U12526 ( .A(n12592), .B(n12593), .Z(n12591) );
  OR2_X1 U12527 ( .A1(n8191), .A2(n8216), .ZN(n12404) );
  XOR2_X1 U12528 ( .A(n12594), .B(n12595), .Z(n12401) );
  XOR2_X1 U12529 ( .A(n12596), .B(n12597), .Z(n12595) );
  OR2_X1 U12530 ( .A1(n8107), .A2(n8216), .ZN(n12408) );
  XOR2_X1 U12531 ( .A(n12598), .B(n12599), .Z(n12405) );
  XOR2_X1 U12532 ( .A(n12600), .B(n12601), .Z(n12599) );
  OR2_X1 U12533 ( .A1(n8025), .A2(n8216), .ZN(n12412) );
  XOR2_X1 U12534 ( .A(n12602), .B(n12603), .Z(n12409) );
  XOR2_X1 U12535 ( .A(n12604), .B(n12605), .Z(n12603) );
  OR2_X1 U12536 ( .A1(n7955), .A2(n8216), .ZN(n12416) );
  XOR2_X1 U12537 ( .A(n12606), .B(n12607), .Z(n12413) );
  XOR2_X1 U12538 ( .A(n12608), .B(n12609), .Z(n12607) );
  OR2_X1 U12539 ( .A1(n7887), .A2(n8216), .ZN(n12420) );
  XOR2_X1 U12540 ( .A(n12610), .B(n12611), .Z(n12417) );
  XOR2_X1 U12541 ( .A(n12612), .B(n12613), .Z(n12611) );
  OR2_X1 U12542 ( .A1(n7828), .A2(n8216), .ZN(n12424) );
  XOR2_X1 U12543 ( .A(n12614), .B(n12615), .Z(n12421) );
  XOR2_X1 U12544 ( .A(n12616), .B(n12617), .Z(n12615) );
  OR2_X1 U12545 ( .A1(n7820), .A2(n8216), .ZN(n12428) );
  XOR2_X1 U12546 ( .A(n12618), .B(n12619), .Z(n12425) );
  XOR2_X1 U12547 ( .A(n12620), .B(n12621), .Z(n12619) );
  XOR2_X1 U12548 ( .A(n11737), .B(n12622), .Z(n11730) );
  XOR2_X1 U12549 ( .A(n11736), .B(n11735), .Z(n12622) );
  OR2_X1 U12550 ( .A1(n7820), .A2(n8133), .ZN(n11735) );
  OR2_X1 U12551 ( .A1(n12623), .A2(n12624), .ZN(n11736) );
  AND2_X1 U12552 ( .A1(n12621), .A2(n12620), .ZN(n12624) );
  AND2_X1 U12553 ( .A1(n12618), .A2(n12625), .ZN(n12623) );
  OR2_X1 U12554 ( .A1(n12620), .A2(n12621), .ZN(n12625) );
  OR2_X1 U12555 ( .A1(n7828), .A2(n8133), .ZN(n12621) );
  OR2_X1 U12556 ( .A1(n12626), .A2(n12627), .ZN(n12620) );
  AND2_X1 U12557 ( .A1(n12617), .A2(n12616), .ZN(n12627) );
  AND2_X1 U12558 ( .A1(n12614), .A2(n12628), .ZN(n12626) );
  OR2_X1 U12559 ( .A1(n12616), .A2(n12617), .ZN(n12628) );
  OR2_X1 U12560 ( .A1(n7887), .A2(n8133), .ZN(n12617) );
  OR2_X1 U12561 ( .A1(n12629), .A2(n12630), .ZN(n12616) );
  AND2_X1 U12562 ( .A1(n12613), .A2(n12612), .ZN(n12630) );
  AND2_X1 U12563 ( .A1(n12610), .A2(n12631), .ZN(n12629) );
  OR2_X1 U12564 ( .A1(n12612), .A2(n12613), .ZN(n12631) );
  OR2_X1 U12565 ( .A1(n7955), .A2(n8133), .ZN(n12613) );
  OR2_X1 U12566 ( .A1(n12632), .A2(n12633), .ZN(n12612) );
  AND2_X1 U12567 ( .A1(n12609), .A2(n12608), .ZN(n12633) );
  AND2_X1 U12568 ( .A1(n12606), .A2(n12634), .ZN(n12632) );
  OR2_X1 U12569 ( .A1(n12608), .A2(n12609), .ZN(n12634) );
  OR2_X1 U12570 ( .A1(n8025), .A2(n8133), .ZN(n12609) );
  OR2_X1 U12571 ( .A1(n12635), .A2(n12636), .ZN(n12608) );
  AND2_X1 U12572 ( .A1(n12605), .A2(n12604), .ZN(n12636) );
  AND2_X1 U12573 ( .A1(n12602), .A2(n12637), .ZN(n12635) );
  OR2_X1 U12574 ( .A1(n12604), .A2(n12605), .ZN(n12637) );
  OR2_X1 U12575 ( .A1(n8107), .A2(n8133), .ZN(n12605) );
  OR2_X1 U12576 ( .A1(n12638), .A2(n12639), .ZN(n12604) );
  AND2_X1 U12577 ( .A1(n12601), .A2(n12600), .ZN(n12639) );
  AND2_X1 U12578 ( .A1(n12598), .A2(n12640), .ZN(n12638) );
  OR2_X1 U12579 ( .A1(n12600), .A2(n12601), .ZN(n12640) );
  OR2_X1 U12580 ( .A1(n8191), .A2(n8133), .ZN(n12601) );
  OR2_X1 U12581 ( .A1(n12641), .A2(n12642), .ZN(n12600) );
  AND2_X1 U12582 ( .A1(n12597), .A2(n12596), .ZN(n12642) );
  AND2_X1 U12583 ( .A1(n12594), .A2(n12643), .ZN(n12641) );
  OR2_X1 U12584 ( .A1(n12596), .A2(n12597), .ZN(n12643) );
  OR2_X1 U12585 ( .A1(n8287), .A2(n8133), .ZN(n12597) );
  OR2_X1 U12586 ( .A1(n12644), .A2(n12645), .ZN(n12596) );
  AND2_X1 U12587 ( .A1(n12593), .A2(n12592), .ZN(n12645) );
  AND2_X1 U12588 ( .A1(n12590), .A2(n12646), .ZN(n12644) );
  OR2_X1 U12589 ( .A1(n12592), .A2(n12593), .ZN(n12646) );
  OR2_X1 U12590 ( .A1(n8608), .A2(n8133), .ZN(n12593) );
  OR2_X1 U12591 ( .A1(n12647), .A2(n12648), .ZN(n12592) );
  AND2_X1 U12592 ( .A1(n12587), .A2(n12589), .ZN(n12648) );
  AND2_X1 U12593 ( .A1(n12649), .A2(n12588), .ZN(n12647) );
  OR2_X1 U12594 ( .A1(n12587), .A2(n12589), .ZN(n12649) );
  OR2_X1 U12595 ( .A1(n12650), .A2(n12651), .ZN(n12589) );
  AND2_X1 U12596 ( .A1(n12585), .A2(n12584), .ZN(n12651) );
  AND2_X1 U12597 ( .A1(n12582), .A2(n12652), .ZN(n12650) );
  OR2_X1 U12598 ( .A1(n12584), .A2(n12585), .ZN(n12652) );
  OR2_X1 U12599 ( .A1(n8598), .A2(n8133), .ZN(n12585) );
  OR2_X1 U12600 ( .A1(n12653), .A2(n12654), .ZN(n12584) );
  AND2_X1 U12601 ( .A1(n12581), .A2(n12580), .ZN(n12654) );
  AND2_X1 U12602 ( .A1(n12578), .A2(n12655), .ZN(n12653) );
  OR2_X1 U12603 ( .A1(n12580), .A2(n12581), .ZN(n12655) );
  OR2_X1 U12604 ( .A1(n8593), .A2(n8133), .ZN(n12581) );
  OR2_X1 U12605 ( .A1(n12656), .A2(n12657), .ZN(n12580) );
  AND2_X1 U12606 ( .A1(n12577), .A2(n12576), .ZN(n12657) );
  AND2_X1 U12607 ( .A1(n12574), .A2(n12658), .ZN(n12656) );
  OR2_X1 U12608 ( .A1(n12576), .A2(n12577), .ZN(n12658) );
  OR2_X1 U12609 ( .A1(n8588), .A2(n8133), .ZN(n12577) );
  OR2_X1 U12610 ( .A1(n12659), .A2(n12660), .ZN(n12576) );
  AND2_X1 U12611 ( .A1(n12573), .A2(n12572), .ZN(n12660) );
  AND2_X1 U12612 ( .A1(n12570), .A2(n12661), .ZN(n12659) );
  OR2_X1 U12613 ( .A1(n12572), .A2(n12573), .ZN(n12661) );
  OR2_X1 U12614 ( .A1(n8583), .A2(n8133), .ZN(n12573) );
  OR2_X1 U12615 ( .A1(n12662), .A2(n12663), .ZN(n12572) );
  AND2_X1 U12616 ( .A1(n12569), .A2(n12568), .ZN(n12663) );
  AND2_X1 U12617 ( .A1(n12566), .A2(n12664), .ZN(n12662) );
  OR2_X1 U12618 ( .A1(n12568), .A2(n12569), .ZN(n12664) );
  OR2_X1 U12619 ( .A1(n8578), .A2(n8133), .ZN(n12569) );
  OR2_X1 U12620 ( .A1(n12665), .A2(n12666), .ZN(n12568) );
  AND2_X1 U12621 ( .A1(n12565), .A2(n12564), .ZN(n12666) );
  AND2_X1 U12622 ( .A1(n12562), .A2(n12667), .ZN(n12665) );
  OR2_X1 U12623 ( .A1(n12564), .A2(n12565), .ZN(n12667) );
  OR2_X1 U12624 ( .A1(n8573), .A2(n8133), .ZN(n12565) );
  OR2_X1 U12625 ( .A1(n12668), .A2(n12669), .ZN(n12564) );
  AND2_X1 U12626 ( .A1(n12561), .A2(n12560), .ZN(n12669) );
  AND2_X1 U12627 ( .A1(n12558), .A2(n12670), .ZN(n12668) );
  OR2_X1 U12628 ( .A1(n12560), .A2(n12561), .ZN(n12670) );
  OR2_X1 U12629 ( .A1(n8568), .A2(n8133), .ZN(n12561) );
  OR2_X1 U12630 ( .A1(n12671), .A2(n12672), .ZN(n12560) );
  AND2_X1 U12631 ( .A1(n12557), .A2(n12556), .ZN(n12672) );
  AND2_X1 U12632 ( .A1(n12554), .A2(n12673), .ZN(n12671) );
  OR2_X1 U12633 ( .A1(n12556), .A2(n12557), .ZN(n12673) );
  OR2_X1 U12634 ( .A1(n8563), .A2(n8133), .ZN(n12557) );
  OR2_X1 U12635 ( .A1(n12674), .A2(n12675), .ZN(n12556) );
  AND2_X1 U12636 ( .A1(n12553), .A2(n12552), .ZN(n12675) );
  AND2_X1 U12637 ( .A1(n12550), .A2(n12676), .ZN(n12674) );
  OR2_X1 U12638 ( .A1(n12552), .A2(n12553), .ZN(n12676) );
  OR2_X1 U12639 ( .A1(n8558), .A2(n8133), .ZN(n12553) );
  OR2_X1 U12640 ( .A1(n12677), .A2(n12678), .ZN(n12552) );
  AND2_X1 U12641 ( .A1(n12549), .A2(n12548), .ZN(n12678) );
  AND2_X1 U12642 ( .A1(n12546), .A2(n12679), .ZN(n12677) );
  OR2_X1 U12643 ( .A1(n12548), .A2(n12549), .ZN(n12679) );
  OR2_X1 U12644 ( .A1(n8553), .A2(n8133), .ZN(n12549) );
  OR2_X1 U12645 ( .A1(n12680), .A2(n12681), .ZN(n12548) );
  AND2_X1 U12646 ( .A1(n12545), .A2(n12544), .ZN(n12681) );
  AND2_X1 U12647 ( .A1(n12542), .A2(n12682), .ZN(n12680) );
  OR2_X1 U12648 ( .A1(n12544), .A2(n12545), .ZN(n12682) );
  OR2_X1 U12649 ( .A1(n8548), .A2(n8133), .ZN(n12545) );
  OR2_X1 U12650 ( .A1(n12683), .A2(n12684), .ZN(n12544) );
  AND2_X1 U12651 ( .A1(n12541), .A2(n12540), .ZN(n12684) );
  AND2_X1 U12652 ( .A1(n12538), .A2(n12685), .ZN(n12683) );
  OR2_X1 U12653 ( .A1(n12540), .A2(n12541), .ZN(n12685) );
  OR2_X1 U12654 ( .A1(n8543), .A2(n8133), .ZN(n12541) );
  OR2_X1 U12655 ( .A1(n12686), .A2(n12687), .ZN(n12540) );
  AND2_X1 U12656 ( .A1(n12537), .A2(n12536), .ZN(n12687) );
  AND2_X1 U12657 ( .A1(n12534), .A2(n12688), .ZN(n12686) );
  OR2_X1 U12658 ( .A1(n12536), .A2(n12537), .ZN(n12688) );
  OR2_X1 U12659 ( .A1(n8538), .A2(n8133), .ZN(n12537) );
  OR2_X1 U12660 ( .A1(n12689), .A2(n12690), .ZN(n12536) );
  AND2_X1 U12661 ( .A1(n12533), .A2(n12532), .ZN(n12690) );
  AND2_X1 U12662 ( .A1(n12530), .A2(n12691), .ZN(n12689) );
  OR2_X1 U12663 ( .A1(n12532), .A2(n12533), .ZN(n12691) );
  OR2_X1 U12664 ( .A1(n8533), .A2(n8133), .ZN(n12533) );
  OR2_X1 U12665 ( .A1(n12692), .A2(n12693), .ZN(n12532) );
  AND2_X1 U12666 ( .A1(n12529), .A2(n12528), .ZN(n12693) );
  AND2_X1 U12667 ( .A1(n12526), .A2(n12694), .ZN(n12692) );
  OR2_X1 U12668 ( .A1(n12528), .A2(n12529), .ZN(n12694) );
  OR2_X1 U12669 ( .A1(n8528), .A2(n8133), .ZN(n12529) );
  OR2_X1 U12670 ( .A1(n12695), .A2(n12696), .ZN(n12528) );
  AND2_X1 U12671 ( .A1(n12525), .A2(n12524), .ZN(n12696) );
  AND2_X1 U12672 ( .A1(n12522), .A2(n12697), .ZN(n12695) );
  OR2_X1 U12673 ( .A1(n12524), .A2(n12525), .ZN(n12697) );
  OR2_X1 U12674 ( .A1(n8523), .A2(n8133), .ZN(n12525) );
  OR2_X1 U12675 ( .A1(n12698), .A2(n12699), .ZN(n12524) );
  AND2_X1 U12676 ( .A1(n12519), .A2(n12520), .ZN(n12699) );
  AND2_X1 U12677 ( .A1(n12700), .A2(n12701), .ZN(n12698) );
  OR2_X1 U12678 ( .A1(n12520), .A2(n12519), .ZN(n12701) );
  OR2_X1 U12679 ( .A1(n8515), .A2(n8133), .ZN(n12519) );
  OR2_X1 U12680 ( .A1(n8133), .A2(n12702), .ZN(n12520) );
  OR2_X1 U12681 ( .A1(n8050), .A2(n8956), .ZN(n12702) );
  INV_X1 U12682 ( .A(n12521), .ZN(n12700) );
  OR2_X1 U12683 ( .A1(n12703), .A2(n12704), .ZN(n12521) );
  AND2_X1 U12684 ( .A1(b_11_), .A2(n12705), .ZN(n12704) );
  OR2_X1 U12685 ( .A1(n12706), .A2(n7343), .ZN(n12705) );
  AND2_X1 U12686 ( .A1(a_30_), .A2(n7981), .ZN(n12706) );
  AND2_X1 U12687 ( .A1(b_10_), .A2(n12707), .ZN(n12703) );
  OR2_X1 U12688 ( .A1(n12708), .A2(n7347), .ZN(n12707) );
  AND2_X1 U12689 ( .A1(a_31_), .A2(n8050), .ZN(n12708) );
  XOR2_X1 U12690 ( .A(n12709), .B(n12710), .Z(n12522) );
  XNOR2_X1 U12691 ( .A(n12711), .B(n12712), .ZN(n12709) );
  XOR2_X1 U12692 ( .A(n12713), .B(n12714), .Z(n12526) );
  XOR2_X1 U12693 ( .A(n12715), .B(n12716), .Z(n12714) );
  XOR2_X1 U12694 ( .A(n12717), .B(n12718), .Z(n12530) );
  XOR2_X1 U12695 ( .A(n12719), .B(n12720), .Z(n12718) );
  XOR2_X1 U12696 ( .A(n12721), .B(n12722), .Z(n12534) );
  XOR2_X1 U12697 ( .A(n12723), .B(n12724), .Z(n12722) );
  XOR2_X1 U12698 ( .A(n12725), .B(n12726), .Z(n12538) );
  XOR2_X1 U12699 ( .A(n12727), .B(n12728), .Z(n12726) );
  XOR2_X1 U12700 ( .A(n12729), .B(n12730), .Z(n12542) );
  XOR2_X1 U12701 ( .A(n12731), .B(n12732), .Z(n12730) );
  XOR2_X1 U12702 ( .A(n12733), .B(n12734), .Z(n12546) );
  XOR2_X1 U12703 ( .A(n12735), .B(n12736), .Z(n12734) );
  XOR2_X1 U12704 ( .A(n12737), .B(n12738), .Z(n12550) );
  XOR2_X1 U12705 ( .A(n12739), .B(n12740), .Z(n12738) );
  XOR2_X1 U12706 ( .A(n12741), .B(n12742), .Z(n12554) );
  XOR2_X1 U12707 ( .A(n12743), .B(n12744), .Z(n12742) );
  XOR2_X1 U12708 ( .A(n12745), .B(n12746), .Z(n12558) );
  XOR2_X1 U12709 ( .A(n12747), .B(n12748), .Z(n12746) );
  XOR2_X1 U12710 ( .A(n12749), .B(n12750), .Z(n12562) );
  XOR2_X1 U12711 ( .A(n12751), .B(n12752), .Z(n12750) );
  XOR2_X1 U12712 ( .A(n12753), .B(n12754), .Z(n12566) );
  XOR2_X1 U12713 ( .A(n12755), .B(n12756), .Z(n12754) );
  XOR2_X1 U12714 ( .A(n12757), .B(n12758), .Z(n12570) );
  XOR2_X1 U12715 ( .A(n12759), .B(n12760), .Z(n12758) );
  XOR2_X1 U12716 ( .A(n12761), .B(n12762), .Z(n12574) );
  XOR2_X1 U12717 ( .A(n12763), .B(n12764), .Z(n12762) );
  XOR2_X1 U12718 ( .A(n12765), .B(n12766), .Z(n12578) );
  XOR2_X1 U12719 ( .A(n12767), .B(n12768), .Z(n12766) );
  XOR2_X1 U12720 ( .A(n12769), .B(n12770), .Z(n12582) );
  XOR2_X1 U12721 ( .A(n12771), .B(n12772), .Z(n12770) );
  XOR2_X1 U12722 ( .A(n12773), .B(n12774), .Z(n12587) );
  XOR2_X1 U12723 ( .A(n12775), .B(n12776), .Z(n12774) );
  XOR2_X1 U12724 ( .A(n12777), .B(n12778), .Z(n12590) );
  XOR2_X1 U12725 ( .A(n12779), .B(n12780), .Z(n12778) );
  XNOR2_X1 U12726 ( .A(n12781), .B(n12782), .ZN(n12594) );
  XNOR2_X1 U12727 ( .A(n12783), .B(n12784), .ZN(n12781) );
  XOR2_X1 U12728 ( .A(n12785), .B(n12786), .Z(n12598) );
  XOR2_X1 U12729 ( .A(n12787), .B(n12788), .Z(n12786) );
  XOR2_X1 U12730 ( .A(n12789), .B(n12790), .Z(n12602) );
  XOR2_X1 U12731 ( .A(n12791), .B(n12792), .Z(n12790) );
  XOR2_X1 U12732 ( .A(n12793), .B(n12794), .Z(n12606) );
  XOR2_X1 U12733 ( .A(n12795), .B(n12796), .Z(n12794) );
  XOR2_X1 U12734 ( .A(n12797), .B(n12798), .Z(n12610) );
  XOR2_X1 U12735 ( .A(n12799), .B(n12800), .Z(n12798) );
  XOR2_X1 U12736 ( .A(n12801), .B(n12802), .Z(n12614) );
  XOR2_X1 U12737 ( .A(n12803), .B(n12804), .Z(n12802) );
  XOR2_X1 U12738 ( .A(n12805), .B(n12806), .Z(n12618) );
  XOR2_X1 U12739 ( .A(n12807), .B(n12808), .Z(n12806) );
  XOR2_X1 U12740 ( .A(n11744), .B(n12809), .Z(n11737) );
  XOR2_X1 U12741 ( .A(n11743), .B(n11742), .Z(n12809) );
  OR2_X1 U12742 ( .A1(n8050), .A2(n7828), .ZN(n11742) );
  OR2_X1 U12743 ( .A1(n12810), .A2(n12811), .ZN(n11743) );
  AND2_X1 U12744 ( .A1(n12808), .A2(n12807), .ZN(n12811) );
  AND2_X1 U12745 ( .A1(n12805), .A2(n12812), .ZN(n12810) );
  OR2_X1 U12746 ( .A1(n12808), .A2(n12807), .ZN(n12812) );
  OR2_X1 U12747 ( .A1(n12813), .A2(n12814), .ZN(n12807) );
  AND2_X1 U12748 ( .A1(n12804), .A2(n12803), .ZN(n12814) );
  AND2_X1 U12749 ( .A1(n12801), .A2(n12815), .ZN(n12813) );
  OR2_X1 U12750 ( .A1(n12804), .A2(n12803), .ZN(n12815) );
  OR2_X1 U12751 ( .A1(n12816), .A2(n12817), .ZN(n12803) );
  AND2_X1 U12752 ( .A1(n12800), .A2(n12799), .ZN(n12817) );
  AND2_X1 U12753 ( .A1(n12797), .A2(n12818), .ZN(n12816) );
  OR2_X1 U12754 ( .A1(n12800), .A2(n12799), .ZN(n12818) );
  OR2_X1 U12755 ( .A1(n12819), .A2(n12820), .ZN(n12799) );
  AND2_X1 U12756 ( .A1(n12796), .A2(n12795), .ZN(n12820) );
  AND2_X1 U12757 ( .A1(n12793), .A2(n12821), .ZN(n12819) );
  OR2_X1 U12758 ( .A1(n12796), .A2(n12795), .ZN(n12821) );
  OR2_X1 U12759 ( .A1(n12822), .A2(n12823), .ZN(n12795) );
  AND2_X1 U12760 ( .A1(n12792), .A2(n12791), .ZN(n12823) );
  AND2_X1 U12761 ( .A1(n12789), .A2(n12824), .ZN(n12822) );
  OR2_X1 U12762 ( .A1(n12792), .A2(n12791), .ZN(n12824) );
  OR2_X1 U12763 ( .A1(n12825), .A2(n12826), .ZN(n12791) );
  AND2_X1 U12764 ( .A1(n12788), .A2(n12787), .ZN(n12826) );
  AND2_X1 U12765 ( .A1(n12785), .A2(n12827), .ZN(n12825) );
  OR2_X1 U12766 ( .A1(n12788), .A2(n12787), .ZN(n12827) );
  OR2_X1 U12767 ( .A1(n12828), .A2(n12829), .ZN(n12787) );
  AND2_X1 U12768 ( .A1(n12782), .A2(n12784), .ZN(n12829) );
  AND2_X1 U12769 ( .A1(n12830), .A2(n12783), .ZN(n12828) );
  OR2_X1 U12770 ( .A1(n12782), .A2(n12784), .ZN(n12830) );
  OR2_X1 U12771 ( .A1(n12831), .A2(n12832), .ZN(n12784) );
  AND2_X1 U12772 ( .A1(n12780), .A2(n12779), .ZN(n12832) );
  AND2_X1 U12773 ( .A1(n12777), .A2(n12833), .ZN(n12831) );
  OR2_X1 U12774 ( .A1(n12780), .A2(n12779), .ZN(n12833) );
  OR2_X1 U12775 ( .A1(n12834), .A2(n12835), .ZN(n12779) );
  AND2_X1 U12776 ( .A1(n12776), .A2(n12775), .ZN(n12835) );
  AND2_X1 U12777 ( .A1(n12773), .A2(n12836), .ZN(n12834) );
  OR2_X1 U12778 ( .A1(n12776), .A2(n12775), .ZN(n12836) );
  OR2_X1 U12779 ( .A1(n12837), .A2(n12838), .ZN(n12775) );
  AND2_X1 U12780 ( .A1(n12772), .A2(n12771), .ZN(n12838) );
  AND2_X1 U12781 ( .A1(n12769), .A2(n12839), .ZN(n12837) );
  OR2_X1 U12782 ( .A1(n12772), .A2(n12771), .ZN(n12839) );
  OR2_X1 U12783 ( .A1(n12840), .A2(n12841), .ZN(n12771) );
  AND2_X1 U12784 ( .A1(n12768), .A2(n12767), .ZN(n12841) );
  AND2_X1 U12785 ( .A1(n12765), .A2(n12842), .ZN(n12840) );
  OR2_X1 U12786 ( .A1(n12768), .A2(n12767), .ZN(n12842) );
  OR2_X1 U12787 ( .A1(n12843), .A2(n12844), .ZN(n12767) );
  AND2_X1 U12788 ( .A1(n12764), .A2(n12763), .ZN(n12844) );
  AND2_X1 U12789 ( .A1(n12761), .A2(n12845), .ZN(n12843) );
  OR2_X1 U12790 ( .A1(n12764), .A2(n12763), .ZN(n12845) );
  OR2_X1 U12791 ( .A1(n12846), .A2(n12847), .ZN(n12763) );
  AND2_X1 U12792 ( .A1(n12760), .A2(n12759), .ZN(n12847) );
  AND2_X1 U12793 ( .A1(n12757), .A2(n12848), .ZN(n12846) );
  OR2_X1 U12794 ( .A1(n12760), .A2(n12759), .ZN(n12848) );
  OR2_X1 U12795 ( .A1(n12849), .A2(n12850), .ZN(n12759) );
  AND2_X1 U12796 ( .A1(n12756), .A2(n12755), .ZN(n12850) );
  AND2_X1 U12797 ( .A1(n12753), .A2(n12851), .ZN(n12849) );
  OR2_X1 U12798 ( .A1(n12756), .A2(n12755), .ZN(n12851) );
  OR2_X1 U12799 ( .A1(n12852), .A2(n12853), .ZN(n12755) );
  AND2_X1 U12800 ( .A1(n12752), .A2(n12751), .ZN(n12853) );
  AND2_X1 U12801 ( .A1(n12749), .A2(n12854), .ZN(n12852) );
  OR2_X1 U12802 ( .A1(n12752), .A2(n12751), .ZN(n12854) );
  OR2_X1 U12803 ( .A1(n12855), .A2(n12856), .ZN(n12751) );
  AND2_X1 U12804 ( .A1(n12748), .A2(n12747), .ZN(n12856) );
  AND2_X1 U12805 ( .A1(n12745), .A2(n12857), .ZN(n12855) );
  OR2_X1 U12806 ( .A1(n12748), .A2(n12747), .ZN(n12857) );
  OR2_X1 U12807 ( .A1(n12858), .A2(n12859), .ZN(n12747) );
  AND2_X1 U12808 ( .A1(n12744), .A2(n12743), .ZN(n12859) );
  AND2_X1 U12809 ( .A1(n12741), .A2(n12860), .ZN(n12858) );
  OR2_X1 U12810 ( .A1(n12744), .A2(n12743), .ZN(n12860) );
  OR2_X1 U12811 ( .A1(n12861), .A2(n12862), .ZN(n12743) );
  AND2_X1 U12812 ( .A1(n12740), .A2(n12739), .ZN(n12862) );
  AND2_X1 U12813 ( .A1(n12737), .A2(n12863), .ZN(n12861) );
  OR2_X1 U12814 ( .A1(n12740), .A2(n12739), .ZN(n12863) );
  OR2_X1 U12815 ( .A1(n12864), .A2(n12865), .ZN(n12739) );
  AND2_X1 U12816 ( .A1(n12736), .A2(n12735), .ZN(n12865) );
  AND2_X1 U12817 ( .A1(n12733), .A2(n12866), .ZN(n12864) );
  OR2_X1 U12818 ( .A1(n12736), .A2(n12735), .ZN(n12866) );
  OR2_X1 U12819 ( .A1(n12867), .A2(n12868), .ZN(n12735) );
  AND2_X1 U12820 ( .A1(n12732), .A2(n12731), .ZN(n12868) );
  AND2_X1 U12821 ( .A1(n12729), .A2(n12869), .ZN(n12867) );
  OR2_X1 U12822 ( .A1(n12732), .A2(n12731), .ZN(n12869) );
  OR2_X1 U12823 ( .A1(n12870), .A2(n12871), .ZN(n12731) );
  AND2_X1 U12824 ( .A1(n12728), .A2(n12727), .ZN(n12871) );
  AND2_X1 U12825 ( .A1(n12725), .A2(n12872), .ZN(n12870) );
  OR2_X1 U12826 ( .A1(n12728), .A2(n12727), .ZN(n12872) );
  OR2_X1 U12827 ( .A1(n12873), .A2(n12874), .ZN(n12727) );
  AND2_X1 U12828 ( .A1(n12724), .A2(n12723), .ZN(n12874) );
  AND2_X1 U12829 ( .A1(n12721), .A2(n12875), .ZN(n12873) );
  OR2_X1 U12830 ( .A1(n12724), .A2(n12723), .ZN(n12875) );
  OR2_X1 U12831 ( .A1(n12876), .A2(n12877), .ZN(n12723) );
  AND2_X1 U12832 ( .A1(n12720), .A2(n12719), .ZN(n12877) );
  AND2_X1 U12833 ( .A1(n12717), .A2(n12878), .ZN(n12876) );
  OR2_X1 U12834 ( .A1(n12720), .A2(n12719), .ZN(n12878) );
  OR2_X1 U12835 ( .A1(n12879), .A2(n12880), .ZN(n12719) );
  AND2_X1 U12836 ( .A1(n12716), .A2(n12715), .ZN(n12880) );
  AND2_X1 U12837 ( .A1(n12713), .A2(n12881), .ZN(n12879) );
  OR2_X1 U12838 ( .A1(n12716), .A2(n12715), .ZN(n12881) );
  OR2_X1 U12839 ( .A1(n12882), .A2(n12883), .ZN(n12715) );
  AND2_X1 U12840 ( .A1(n12710), .A2(n12711), .ZN(n12883) );
  AND2_X1 U12841 ( .A1(n12884), .A2(n12885), .ZN(n12882) );
  OR2_X1 U12842 ( .A1(n12710), .A2(n12711), .ZN(n12885) );
  OR2_X1 U12843 ( .A1(n8956), .A2(n12886), .ZN(n12711) );
  OR2_X1 U12844 ( .A1(n8050), .A2(n7981), .ZN(n12886) );
  OR2_X1 U12845 ( .A1(n8050), .A2(n8515), .ZN(n12710) );
  INV_X1 U12846 ( .A(n12712), .ZN(n12884) );
  OR2_X1 U12847 ( .A1(n12887), .A2(n12888), .ZN(n12712) );
  AND2_X1 U12848 ( .A1(b_9_), .A2(n12889), .ZN(n12888) );
  OR2_X1 U12849 ( .A1(n12890), .A2(n7347), .ZN(n12889) );
  AND2_X1 U12850 ( .A1(a_31_), .A2(n7981), .ZN(n12890) );
  AND2_X1 U12851 ( .A1(b_10_), .A2(n12891), .ZN(n12887) );
  OR2_X1 U12852 ( .A1(n12892), .A2(n7343), .ZN(n12891) );
  AND2_X1 U12853 ( .A1(a_30_), .A2(n7912), .ZN(n12892) );
  OR2_X1 U12854 ( .A1(n8050), .A2(n8523), .ZN(n12716) );
  XOR2_X1 U12855 ( .A(n12893), .B(n12894), .Z(n12713) );
  XNOR2_X1 U12856 ( .A(n12895), .B(n12896), .ZN(n12893) );
  OR2_X1 U12857 ( .A1(n8050), .A2(n8528), .ZN(n12720) );
  XOR2_X1 U12858 ( .A(n12897), .B(n12898), .Z(n12717) );
  XOR2_X1 U12859 ( .A(n12899), .B(n12900), .Z(n12898) );
  OR2_X1 U12860 ( .A1(n8050), .A2(n8533), .ZN(n12724) );
  XOR2_X1 U12861 ( .A(n12901), .B(n12902), .Z(n12721) );
  XOR2_X1 U12862 ( .A(n12903), .B(n12904), .Z(n12902) );
  OR2_X1 U12863 ( .A1(n8050), .A2(n8538), .ZN(n12728) );
  XOR2_X1 U12864 ( .A(n12905), .B(n12906), .Z(n12725) );
  XOR2_X1 U12865 ( .A(n12907), .B(n12908), .Z(n12906) );
  OR2_X1 U12866 ( .A1(n8050), .A2(n8543), .ZN(n12732) );
  XOR2_X1 U12867 ( .A(n12909), .B(n12910), .Z(n12729) );
  XOR2_X1 U12868 ( .A(n12911), .B(n12912), .Z(n12910) );
  OR2_X1 U12869 ( .A1(n8050), .A2(n8548), .ZN(n12736) );
  XOR2_X1 U12870 ( .A(n12913), .B(n12914), .Z(n12733) );
  XOR2_X1 U12871 ( .A(n12915), .B(n12916), .Z(n12914) );
  OR2_X1 U12872 ( .A1(n8050), .A2(n8553), .ZN(n12740) );
  XOR2_X1 U12873 ( .A(n12917), .B(n12918), .Z(n12737) );
  XOR2_X1 U12874 ( .A(n12919), .B(n12920), .Z(n12918) );
  OR2_X1 U12875 ( .A1(n8050), .A2(n8558), .ZN(n12744) );
  XOR2_X1 U12876 ( .A(n12921), .B(n12922), .Z(n12741) );
  XOR2_X1 U12877 ( .A(n12923), .B(n12924), .Z(n12922) );
  OR2_X1 U12878 ( .A1(n8050), .A2(n8563), .ZN(n12748) );
  XOR2_X1 U12879 ( .A(n12925), .B(n12926), .Z(n12745) );
  XOR2_X1 U12880 ( .A(n12927), .B(n12928), .Z(n12926) );
  OR2_X1 U12881 ( .A1(n8050), .A2(n8568), .ZN(n12752) );
  XOR2_X1 U12882 ( .A(n12929), .B(n12930), .Z(n12749) );
  XOR2_X1 U12883 ( .A(n12931), .B(n12932), .Z(n12930) );
  OR2_X1 U12884 ( .A1(n8050), .A2(n8573), .ZN(n12756) );
  XOR2_X1 U12885 ( .A(n12933), .B(n12934), .Z(n12753) );
  XOR2_X1 U12886 ( .A(n12935), .B(n12936), .Z(n12934) );
  OR2_X1 U12887 ( .A1(n8050), .A2(n8578), .ZN(n12760) );
  XOR2_X1 U12888 ( .A(n12937), .B(n12938), .Z(n12757) );
  XOR2_X1 U12889 ( .A(n12939), .B(n12940), .Z(n12938) );
  OR2_X1 U12890 ( .A1(n8050), .A2(n8583), .ZN(n12764) );
  XOR2_X1 U12891 ( .A(n12941), .B(n12942), .Z(n12761) );
  XOR2_X1 U12892 ( .A(n12943), .B(n12944), .Z(n12942) );
  OR2_X1 U12893 ( .A1(n8050), .A2(n8588), .ZN(n12768) );
  XOR2_X1 U12894 ( .A(n12945), .B(n12946), .Z(n12765) );
  XOR2_X1 U12895 ( .A(n12947), .B(n12948), .Z(n12946) );
  OR2_X1 U12896 ( .A1(n8050), .A2(n8593), .ZN(n12772) );
  XOR2_X1 U12897 ( .A(n12949), .B(n12950), .Z(n12769) );
  XOR2_X1 U12898 ( .A(n12951), .B(n12952), .Z(n12950) );
  OR2_X1 U12899 ( .A1(n8050), .A2(n8598), .ZN(n12776) );
  XOR2_X1 U12900 ( .A(n12953), .B(n12954), .Z(n12773) );
  XOR2_X1 U12901 ( .A(n12955), .B(n12956), .Z(n12954) );
  OR2_X1 U12902 ( .A1(n8050), .A2(n8603), .ZN(n12780) );
  XOR2_X1 U12903 ( .A(n12957), .B(n12958), .Z(n12777) );
  XOR2_X1 U12904 ( .A(n12959), .B(n12960), .Z(n12958) );
  XOR2_X1 U12905 ( .A(n12961), .B(n12962), .Z(n12782) );
  XOR2_X1 U12906 ( .A(n12963), .B(n12964), .Z(n12962) );
  OR2_X1 U12907 ( .A1(n8050), .A2(n8287), .ZN(n12788) );
  XOR2_X1 U12908 ( .A(n12965), .B(n12966), .Z(n12785) );
  XOR2_X1 U12909 ( .A(n12967), .B(n12968), .Z(n12966) );
  OR2_X1 U12910 ( .A1(n8050), .A2(n8191), .ZN(n12792) );
  XNOR2_X1 U12911 ( .A(n12969), .B(n12970), .ZN(n12789) );
  XNOR2_X1 U12912 ( .A(n12971), .B(n12972), .ZN(n12969) );
  OR2_X1 U12913 ( .A1(n8050), .A2(n8107), .ZN(n12796) );
  XOR2_X1 U12914 ( .A(n12973), .B(n12974), .Z(n12793) );
  XOR2_X1 U12915 ( .A(n12975), .B(n12976), .Z(n12974) );
  OR2_X1 U12916 ( .A1(n8050), .A2(n8025), .ZN(n12800) );
  XOR2_X1 U12917 ( .A(n12977), .B(n12978), .Z(n12797) );
  XOR2_X1 U12918 ( .A(n12979), .B(n12980), .Z(n12978) );
  OR2_X1 U12919 ( .A1(n8050), .A2(n7955), .ZN(n12804) );
  XOR2_X1 U12920 ( .A(n12981), .B(n12982), .Z(n12801) );
  XOR2_X1 U12921 ( .A(n12983), .B(n12984), .Z(n12982) );
  OR2_X1 U12922 ( .A1(n8050), .A2(n7887), .ZN(n12808) );
  XOR2_X1 U12923 ( .A(n12985), .B(n12986), .Z(n12805) );
  XOR2_X1 U12924 ( .A(n12987), .B(n12988), .Z(n12986) );
  XOR2_X1 U12925 ( .A(n11751), .B(n12989), .Z(n11744) );
  XOR2_X1 U12926 ( .A(n11750), .B(n11749), .Z(n12989) );
  OR2_X1 U12927 ( .A1(n7981), .A2(n7887), .ZN(n11749) );
  OR2_X1 U12928 ( .A1(n12990), .A2(n12991), .ZN(n11750) );
  AND2_X1 U12929 ( .A1(n12988), .A2(n12987), .ZN(n12991) );
  AND2_X1 U12930 ( .A1(n12985), .A2(n12992), .ZN(n12990) );
  OR2_X1 U12931 ( .A1(n12987), .A2(n12988), .ZN(n12992) );
  OR2_X1 U12932 ( .A1(n7981), .A2(n7955), .ZN(n12988) );
  OR2_X1 U12933 ( .A1(n12993), .A2(n12994), .ZN(n12987) );
  AND2_X1 U12934 ( .A1(n12984), .A2(n12983), .ZN(n12994) );
  AND2_X1 U12935 ( .A1(n12981), .A2(n12995), .ZN(n12993) );
  OR2_X1 U12936 ( .A1(n12983), .A2(n12984), .ZN(n12995) );
  OR2_X1 U12937 ( .A1(n7981), .A2(n8025), .ZN(n12984) );
  OR2_X1 U12938 ( .A1(n12996), .A2(n12997), .ZN(n12983) );
  AND2_X1 U12939 ( .A1(n12980), .A2(n12979), .ZN(n12997) );
  AND2_X1 U12940 ( .A1(n12977), .A2(n12998), .ZN(n12996) );
  OR2_X1 U12941 ( .A1(n12979), .A2(n12980), .ZN(n12998) );
  OR2_X1 U12942 ( .A1(n7981), .A2(n8107), .ZN(n12980) );
  OR2_X1 U12943 ( .A1(n12999), .A2(n13000), .ZN(n12979) );
  AND2_X1 U12944 ( .A1(n12976), .A2(n12975), .ZN(n13000) );
  AND2_X1 U12945 ( .A1(n12973), .A2(n13001), .ZN(n12999) );
  OR2_X1 U12946 ( .A1(n12975), .A2(n12976), .ZN(n13001) );
  OR2_X1 U12947 ( .A1(n7981), .A2(n8191), .ZN(n12976) );
  OR2_X1 U12948 ( .A1(n13002), .A2(n13003), .ZN(n12975) );
  AND2_X1 U12949 ( .A1(n12970), .A2(n12972), .ZN(n13003) );
  AND2_X1 U12950 ( .A1(n13004), .A2(n12971), .ZN(n13002) );
  OR2_X1 U12951 ( .A1(n12970), .A2(n12972), .ZN(n13004) );
  OR2_X1 U12952 ( .A1(n13005), .A2(n13006), .ZN(n12972) );
  AND2_X1 U12953 ( .A1(n12968), .A2(n12967), .ZN(n13006) );
  AND2_X1 U12954 ( .A1(n12965), .A2(n13007), .ZN(n13005) );
  OR2_X1 U12955 ( .A1(n12967), .A2(n12968), .ZN(n13007) );
  OR2_X1 U12956 ( .A1(n8608), .A2(n7981), .ZN(n12968) );
  OR2_X1 U12957 ( .A1(n13008), .A2(n13009), .ZN(n12967) );
  AND2_X1 U12958 ( .A1(n12964), .A2(n12963), .ZN(n13009) );
  AND2_X1 U12959 ( .A1(n12961), .A2(n13010), .ZN(n13008) );
  OR2_X1 U12960 ( .A1(n12963), .A2(n12964), .ZN(n13010) );
  OR2_X1 U12961 ( .A1(n7981), .A2(n8603), .ZN(n12964) );
  OR2_X1 U12962 ( .A1(n13011), .A2(n13012), .ZN(n12963) );
  AND2_X1 U12963 ( .A1(n12960), .A2(n12959), .ZN(n13012) );
  AND2_X1 U12964 ( .A1(n12957), .A2(n13013), .ZN(n13011) );
  OR2_X1 U12965 ( .A1(n12959), .A2(n12960), .ZN(n13013) );
  OR2_X1 U12966 ( .A1(n7981), .A2(n8598), .ZN(n12960) );
  OR2_X1 U12967 ( .A1(n13014), .A2(n13015), .ZN(n12959) );
  AND2_X1 U12968 ( .A1(n12956), .A2(n12955), .ZN(n13015) );
  AND2_X1 U12969 ( .A1(n12953), .A2(n13016), .ZN(n13014) );
  OR2_X1 U12970 ( .A1(n12955), .A2(n12956), .ZN(n13016) );
  OR2_X1 U12971 ( .A1(n7981), .A2(n8593), .ZN(n12956) );
  OR2_X1 U12972 ( .A1(n13017), .A2(n13018), .ZN(n12955) );
  AND2_X1 U12973 ( .A1(n12952), .A2(n12951), .ZN(n13018) );
  AND2_X1 U12974 ( .A1(n12949), .A2(n13019), .ZN(n13017) );
  OR2_X1 U12975 ( .A1(n12951), .A2(n12952), .ZN(n13019) );
  OR2_X1 U12976 ( .A1(n7981), .A2(n8588), .ZN(n12952) );
  OR2_X1 U12977 ( .A1(n13020), .A2(n13021), .ZN(n12951) );
  AND2_X1 U12978 ( .A1(n12948), .A2(n12947), .ZN(n13021) );
  AND2_X1 U12979 ( .A1(n12945), .A2(n13022), .ZN(n13020) );
  OR2_X1 U12980 ( .A1(n12947), .A2(n12948), .ZN(n13022) );
  OR2_X1 U12981 ( .A1(n7981), .A2(n8583), .ZN(n12948) );
  OR2_X1 U12982 ( .A1(n13023), .A2(n13024), .ZN(n12947) );
  AND2_X1 U12983 ( .A1(n12944), .A2(n12943), .ZN(n13024) );
  AND2_X1 U12984 ( .A1(n12941), .A2(n13025), .ZN(n13023) );
  OR2_X1 U12985 ( .A1(n12943), .A2(n12944), .ZN(n13025) );
  OR2_X1 U12986 ( .A1(n7981), .A2(n8578), .ZN(n12944) );
  OR2_X1 U12987 ( .A1(n13026), .A2(n13027), .ZN(n12943) );
  AND2_X1 U12988 ( .A1(n12940), .A2(n12939), .ZN(n13027) );
  AND2_X1 U12989 ( .A1(n12937), .A2(n13028), .ZN(n13026) );
  OR2_X1 U12990 ( .A1(n12939), .A2(n12940), .ZN(n13028) );
  OR2_X1 U12991 ( .A1(n7981), .A2(n8573), .ZN(n12940) );
  OR2_X1 U12992 ( .A1(n13029), .A2(n13030), .ZN(n12939) );
  AND2_X1 U12993 ( .A1(n12933), .A2(n12936), .ZN(n13030) );
  AND2_X1 U12994 ( .A1(n13031), .A2(n12935), .ZN(n13029) );
  OR2_X1 U12995 ( .A1(n13032), .A2(n13033), .ZN(n12935) );
  AND2_X1 U12996 ( .A1(n12932), .A2(n12931), .ZN(n13033) );
  AND2_X1 U12997 ( .A1(n12929), .A2(n13034), .ZN(n13032) );
  OR2_X1 U12998 ( .A1(n12931), .A2(n12932), .ZN(n13034) );
  OR2_X1 U12999 ( .A1(n7981), .A2(n8563), .ZN(n12932) );
  OR2_X1 U13000 ( .A1(n13035), .A2(n13036), .ZN(n12931) );
  AND2_X1 U13001 ( .A1(n12925), .A2(n12928), .ZN(n13036) );
  AND2_X1 U13002 ( .A1(n13037), .A2(n12927), .ZN(n13035) );
  OR2_X1 U13003 ( .A1(n13038), .A2(n13039), .ZN(n12927) );
  AND2_X1 U13004 ( .A1(n12921), .A2(n12924), .ZN(n13039) );
  AND2_X1 U13005 ( .A1(n13040), .A2(n12923), .ZN(n13038) );
  OR2_X1 U13006 ( .A1(n13041), .A2(n13042), .ZN(n12923) );
  AND2_X1 U13007 ( .A1(n12917), .A2(n12920), .ZN(n13042) );
  AND2_X1 U13008 ( .A1(n13043), .A2(n12919), .ZN(n13041) );
  OR2_X1 U13009 ( .A1(n13044), .A2(n13045), .ZN(n12919) );
  AND2_X1 U13010 ( .A1(n12913), .A2(n12916), .ZN(n13045) );
  AND2_X1 U13011 ( .A1(n13046), .A2(n12915), .ZN(n13044) );
  OR2_X1 U13012 ( .A1(n13047), .A2(n13048), .ZN(n12915) );
  AND2_X1 U13013 ( .A1(n12909), .A2(n12912), .ZN(n13048) );
  AND2_X1 U13014 ( .A1(n13049), .A2(n12911), .ZN(n13047) );
  OR2_X1 U13015 ( .A1(n13050), .A2(n13051), .ZN(n12911) );
  AND2_X1 U13016 ( .A1(n12905), .A2(n12908), .ZN(n13051) );
  AND2_X1 U13017 ( .A1(n13052), .A2(n12907), .ZN(n13050) );
  OR2_X1 U13018 ( .A1(n13053), .A2(n13054), .ZN(n12907) );
  AND2_X1 U13019 ( .A1(n12901), .A2(n12904), .ZN(n13054) );
  AND2_X1 U13020 ( .A1(n13055), .A2(n12903), .ZN(n13053) );
  OR2_X1 U13021 ( .A1(n13056), .A2(n13057), .ZN(n12903) );
  AND2_X1 U13022 ( .A1(n12897), .A2(n12900), .ZN(n13057) );
  AND2_X1 U13023 ( .A1(n13058), .A2(n12899), .ZN(n13056) );
  OR2_X1 U13024 ( .A1(n13059), .A2(n13060), .ZN(n12899) );
  AND2_X1 U13025 ( .A1(n12894), .A2(n12895), .ZN(n13060) );
  AND2_X1 U13026 ( .A1(n13061), .A2(n13062), .ZN(n13059) );
  OR2_X1 U13027 ( .A1(n12895), .A2(n12894), .ZN(n13062) );
  OR2_X1 U13028 ( .A1(n7981), .A2(n8515), .ZN(n12894) );
  OR2_X1 U13029 ( .A1(n8956), .A2(n13063), .ZN(n12895) );
  OR2_X1 U13030 ( .A1(n7981), .A2(n7912), .ZN(n13063) );
  INV_X1 U13031 ( .A(n12896), .ZN(n13061) );
  OR2_X1 U13032 ( .A1(n13064), .A2(n13065), .ZN(n12896) );
  AND2_X1 U13033 ( .A1(b_9_), .A2(n13066), .ZN(n13065) );
  OR2_X1 U13034 ( .A1(n13067), .A2(n7343), .ZN(n13066) );
  AND2_X1 U13035 ( .A1(a_30_), .A2(n7857), .ZN(n13067) );
  AND2_X1 U13036 ( .A1(b_8_), .A2(n13068), .ZN(n13064) );
  OR2_X1 U13037 ( .A1(n13069), .A2(n7347), .ZN(n13068) );
  AND2_X1 U13038 ( .A1(a_31_), .A2(n7912), .ZN(n13069) );
  OR2_X1 U13039 ( .A1(n12900), .A2(n12897), .ZN(n13058) );
  XOR2_X1 U13040 ( .A(n13070), .B(n13071), .Z(n12897) );
  XNOR2_X1 U13041 ( .A(n13072), .B(n13073), .ZN(n13070) );
  OR2_X1 U13042 ( .A1(n7981), .A2(n8523), .ZN(n12900) );
  OR2_X1 U13043 ( .A1(n12904), .A2(n12901), .ZN(n13055) );
  XOR2_X1 U13044 ( .A(n13074), .B(n13075), .Z(n12901) );
  XOR2_X1 U13045 ( .A(n13076), .B(n13077), .Z(n13075) );
  OR2_X1 U13046 ( .A1(n7981), .A2(n8528), .ZN(n12904) );
  OR2_X1 U13047 ( .A1(n12908), .A2(n12905), .ZN(n13052) );
  XOR2_X1 U13048 ( .A(n13078), .B(n13079), .Z(n12905) );
  XOR2_X1 U13049 ( .A(n13080), .B(n13081), .Z(n13079) );
  OR2_X1 U13050 ( .A1(n7981), .A2(n8533), .ZN(n12908) );
  OR2_X1 U13051 ( .A1(n12912), .A2(n12909), .ZN(n13049) );
  XOR2_X1 U13052 ( .A(n13082), .B(n13083), .Z(n12909) );
  XOR2_X1 U13053 ( .A(n13084), .B(n13085), .Z(n13083) );
  OR2_X1 U13054 ( .A1(n7981), .A2(n8538), .ZN(n12912) );
  OR2_X1 U13055 ( .A1(n12916), .A2(n12913), .ZN(n13046) );
  XOR2_X1 U13056 ( .A(n13086), .B(n13087), .Z(n12913) );
  XOR2_X1 U13057 ( .A(n13088), .B(n13089), .Z(n13087) );
  OR2_X1 U13058 ( .A1(n7981), .A2(n8543), .ZN(n12916) );
  OR2_X1 U13059 ( .A1(n12920), .A2(n12917), .ZN(n13043) );
  XOR2_X1 U13060 ( .A(n13090), .B(n13091), .Z(n12917) );
  XOR2_X1 U13061 ( .A(n13092), .B(n13093), .Z(n13091) );
  OR2_X1 U13062 ( .A1(n7981), .A2(n8548), .ZN(n12920) );
  OR2_X1 U13063 ( .A1(n12924), .A2(n12921), .ZN(n13040) );
  XOR2_X1 U13064 ( .A(n13094), .B(n13095), .Z(n12921) );
  XOR2_X1 U13065 ( .A(n13096), .B(n13097), .Z(n13095) );
  OR2_X1 U13066 ( .A1(n7981), .A2(n8553), .ZN(n12924) );
  OR2_X1 U13067 ( .A1(n12928), .A2(n12925), .ZN(n13037) );
  XOR2_X1 U13068 ( .A(n13098), .B(n13099), .Z(n12925) );
  XOR2_X1 U13069 ( .A(n13100), .B(n13101), .Z(n13099) );
  OR2_X1 U13070 ( .A1(n7981), .A2(n8558), .ZN(n12928) );
  XOR2_X1 U13071 ( .A(n13102), .B(n13103), .Z(n12929) );
  XOR2_X1 U13072 ( .A(n13104), .B(n13105), .Z(n13103) );
  OR2_X1 U13073 ( .A1(n12936), .A2(n12933), .ZN(n13031) );
  XOR2_X1 U13074 ( .A(n13106), .B(n13107), .Z(n12933) );
  XOR2_X1 U13075 ( .A(n13108), .B(n13109), .Z(n13107) );
  OR2_X1 U13076 ( .A1(n7981), .A2(n8568), .ZN(n12936) );
  XOR2_X1 U13077 ( .A(n13110), .B(n13111), .Z(n12937) );
  XOR2_X1 U13078 ( .A(n13112), .B(n13113), .Z(n13111) );
  XOR2_X1 U13079 ( .A(n13114), .B(n13115), .Z(n12941) );
  XOR2_X1 U13080 ( .A(n13116), .B(n13117), .Z(n13115) );
  XOR2_X1 U13081 ( .A(n13118), .B(n13119), .Z(n12945) );
  XOR2_X1 U13082 ( .A(n13120), .B(n13121), .Z(n13119) );
  XOR2_X1 U13083 ( .A(n13122), .B(n13123), .Z(n12949) );
  XOR2_X1 U13084 ( .A(n13124), .B(n13125), .Z(n13123) );
  XOR2_X1 U13085 ( .A(n13126), .B(n13127), .Z(n12953) );
  XOR2_X1 U13086 ( .A(n13128), .B(n13129), .Z(n13127) );
  XOR2_X1 U13087 ( .A(n13130), .B(n13131), .Z(n12957) );
  XOR2_X1 U13088 ( .A(n13132), .B(n13133), .Z(n13131) );
  XOR2_X1 U13089 ( .A(n13134), .B(n13135), .Z(n12961) );
  XOR2_X1 U13090 ( .A(n13136), .B(n13137), .Z(n13135) );
  XOR2_X1 U13091 ( .A(n13138), .B(n13139), .Z(n12965) );
  XOR2_X1 U13092 ( .A(n13140), .B(n13141), .Z(n13139) );
  XOR2_X1 U13093 ( .A(n13142), .B(n13143), .Z(n12970) );
  XOR2_X1 U13094 ( .A(n13144), .B(n13145), .Z(n13143) );
  XOR2_X1 U13095 ( .A(n13146), .B(n13147), .Z(n12973) );
  XOR2_X1 U13096 ( .A(n13148), .B(n13149), .Z(n13147) );
  XNOR2_X1 U13097 ( .A(n13150), .B(n13151), .ZN(n12977) );
  XNOR2_X1 U13098 ( .A(n13152), .B(n13153), .ZN(n13150) );
  XOR2_X1 U13099 ( .A(n13154), .B(n13155), .Z(n12981) );
  XOR2_X1 U13100 ( .A(n13156), .B(n13157), .Z(n13155) );
  XOR2_X1 U13101 ( .A(n13158), .B(n13159), .Z(n12985) );
  XOR2_X1 U13102 ( .A(n13160), .B(n13161), .Z(n13159) );
  XOR2_X1 U13103 ( .A(n11758), .B(n13162), .Z(n11751) );
  XOR2_X1 U13104 ( .A(n11757), .B(n11756), .Z(n13162) );
  OR2_X1 U13105 ( .A1(n7912), .A2(n7955), .ZN(n11756) );
  OR2_X1 U13106 ( .A1(n13163), .A2(n13164), .ZN(n11757) );
  AND2_X1 U13107 ( .A1(n13161), .A2(n13160), .ZN(n13164) );
  AND2_X1 U13108 ( .A1(n13158), .A2(n13165), .ZN(n13163) );
  OR2_X1 U13109 ( .A1(n13160), .A2(n13161), .ZN(n13165) );
  OR2_X1 U13110 ( .A1(n7912), .A2(n8025), .ZN(n13161) );
  OR2_X1 U13111 ( .A1(n13166), .A2(n13167), .ZN(n13160) );
  AND2_X1 U13112 ( .A1(n13157), .A2(n13156), .ZN(n13167) );
  AND2_X1 U13113 ( .A1(n13154), .A2(n13168), .ZN(n13166) );
  OR2_X1 U13114 ( .A1(n13156), .A2(n13157), .ZN(n13168) );
  OR2_X1 U13115 ( .A1(n7912), .A2(n8107), .ZN(n13157) );
  OR2_X1 U13116 ( .A1(n13169), .A2(n13170), .ZN(n13156) );
  AND2_X1 U13117 ( .A1(n13151), .A2(n13153), .ZN(n13170) );
  AND2_X1 U13118 ( .A1(n13171), .A2(n13152), .ZN(n13169) );
  OR2_X1 U13119 ( .A1(n13151), .A2(n13153), .ZN(n13171) );
  OR2_X1 U13120 ( .A1(n13172), .A2(n13173), .ZN(n13153) );
  AND2_X1 U13121 ( .A1(n13149), .A2(n13148), .ZN(n13173) );
  AND2_X1 U13122 ( .A1(n13146), .A2(n13174), .ZN(n13172) );
  OR2_X1 U13123 ( .A1(n13148), .A2(n13149), .ZN(n13174) );
  OR2_X1 U13124 ( .A1(n7912), .A2(n8287), .ZN(n13149) );
  OR2_X1 U13125 ( .A1(n13175), .A2(n13176), .ZN(n13148) );
  AND2_X1 U13126 ( .A1(n13145), .A2(n13144), .ZN(n13176) );
  AND2_X1 U13127 ( .A1(n13142), .A2(n13177), .ZN(n13175) );
  OR2_X1 U13128 ( .A1(n13144), .A2(n13145), .ZN(n13177) );
  OR2_X1 U13129 ( .A1(n8608), .A2(n7912), .ZN(n13145) );
  OR2_X1 U13130 ( .A1(n13178), .A2(n13179), .ZN(n13144) );
  AND2_X1 U13131 ( .A1(n13141), .A2(n13140), .ZN(n13179) );
  AND2_X1 U13132 ( .A1(n13138), .A2(n13180), .ZN(n13178) );
  OR2_X1 U13133 ( .A1(n13140), .A2(n13141), .ZN(n13180) );
  OR2_X1 U13134 ( .A1(n7912), .A2(n8603), .ZN(n13141) );
  OR2_X1 U13135 ( .A1(n13181), .A2(n13182), .ZN(n13140) );
  AND2_X1 U13136 ( .A1(n13137), .A2(n13136), .ZN(n13182) );
  AND2_X1 U13137 ( .A1(n13134), .A2(n13183), .ZN(n13181) );
  OR2_X1 U13138 ( .A1(n13136), .A2(n13137), .ZN(n13183) );
  OR2_X1 U13139 ( .A1(n7912), .A2(n8598), .ZN(n13137) );
  OR2_X1 U13140 ( .A1(n13184), .A2(n13185), .ZN(n13136) );
  AND2_X1 U13141 ( .A1(n13133), .A2(n13132), .ZN(n13185) );
  AND2_X1 U13142 ( .A1(n13130), .A2(n13186), .ZN(n13184) );
  OR2_X1 U13143 ( .A1(n13132), .A2(n13133), .ZN(n13186) );
  OR2_X1 U13144 ( .A1(n7912), .A2(n8593), .ZN(n13133) );
  OR2_X1 U13145 ( .A1(n13187), .A2(n13188), .ZN(n13132) );
  AND2_X1 U13146 ( .A1(n13129), .A2(n13128), .ZN(n13188) );
  AND2_X1 U13147 ( .A1(n13126), .A2(n13189), .ZN(n13187) );
  OR2_X1 U13148 ( .A1(n13128), .A2(n13129), .ZN(n13189) );
  OR2_X1 U13149 ( .A1(n7912), .A2(n8588), .ZN(n13129) );
  OR2_X1 U13150 ( .A1(n13190), .A2(n13191), .ZN(n13128) );
  AND2_X1 U13151 ( .A1(n13125), .A2(n13124), .ZN(n13191) );
  AND2_X1 U13152 ( .A1(n13122), .A2(n13192), .ZN(n13190) );
  OR2_X1 U13153 ( .A1(n13124), .A2(n13125), .ZN(n13192) );
  OR2_X1 U13154 ( .A1(n7912), .A2(n8583), .ZN(n13125) );
  OR2_X1 U13155 ( .A1(n13193), .A2(n13194), .ZN(n13124) );
  AND2_X1 U13156 ( .A1(n13121), .A2(n13120), .ZN(n13194) );
  AND2_X1 U13157 ( .A1(n13118), .A2(n13195), .ZN(n13193) );
  OR2_X1 U13158 ( .A1(n13120), .A2(n13121), .ZN(n13195) );
  OR2_X1 U13159 ( .A1(n7912), .A2(n8578), .ZN(n13121) );
  OR2_X1 U13160 ( .A1(n13196), .A2(n13197), .ZN(n13120) );
  AND2_X1 U13161 ( .A1(n13117), .A2(n13116), .ZN(n13197) );
  AND2_X1 U13162 ( .A1(n13114), .A2(n13198), .ZN(n13196) );
  OR2_X1 U13163 ( .A1(n13116), .A2(n13117), .ZN(n13198) );
  OR2_X1 U13164 ( .A1(n7912), .A2(n8573), .ZN(n13117) );
  OR2_X1 U13165 ( .A1(n13199), .A2(n13200), .ZN(n13116) );
  AND2_X1 U13166 ( .A1(n13113), .A2(n13112), .ZN(n13200) );
  AND2_X1 U13167 ( .A1(n13110), .A2(n13201), .ZN(n13199) );
  OR2_X1 U13168 ( .A1(n13112), .A2(n13113), .ZN(n13201) );
  OR2_X1 U13169 ( .A1(n7912), .A2(n8568), .ZN(n13113) );
  OR2_X1 U13170 ( .A1(n13202), .A2(n13203), .ZN(n13112) );
  AND2_X1 U13171 ( .A1(n13106), .A2(n13109), .ZN(n13203) );
  AND2_X1 U13172 ( .A1(n13204), .A2(n13108), .ZN(n13202) );
  OR2_X1 U13173 ( .A1(n13205), .A2(n13206), .ZN(n13108) );
  AND2_X1 U13174 ( .A1(n13105), .A2(n13104), .ZN(n13206) );
  AND2_X1 U13175 ( .A1(n13102), .A2(n13207), .ZN(n13205) );
  OR2_X1 U13176 ( .A1(n13104), .A2(n13105), .ZN(n13207) );
  OR2_X1 U13177 ( .A1(n7912), .A2(n8558), .ZN(n13105) );
  OR2_X1 U13178 ( .A1(n13208), .A2(n13209), .ZN(n13104) );
  AND2_X1 U13179 ( .A1(n13098), .A2(n13101), .ZN(n13209) );
  AND2_X1 U13180 ( .A1(n13210), .A2(n13100), .ZN(n13208) );
  OR2_X1 U13181 ( .A1(n13211), .A2(n13212), .ZN(n13100) );
  AND2_X1 U13182 ( .A1(n13094), .A2(n13097), .ZN(n13212) );
  AND2_X1 U13183 ( .A1(n13213), .A2(n13096), .ZN(n13211) );
  OR2_X1 U13184 ( .A1(n13214), .A2(n13215), .ZN(n13096) );
  AND2_X1 U13185 ( .A1(n13090), .A2(n13093), .ZN(n13215) );
  AND2_X1 U13186 ( .A1(n13216), .A2(n13092), .ZN(n13214) );
  OR2_X1 U13187 ( .A1(n13217), .A2(n13218), .ZN(n13092) );
  AND2_X1 U13188 ( .A1(n13086), .A2(n13089), .ZN(n13218) );
  AND2_X1 U13189 ( .A1(n13219), .A2(n13088), .ZN(n13217) );
  OR2_X1 U13190 ( .A1(n13220), .A2(n13221), .ZN(n13088) );
  AND2_X1 U13191 ( .A1(n13082), .A2(n13085), .ZN(n13221) );
  AND2_X1 U13192 ( .A1(n13222), .A2(n13084), .ZN(n13220) );
  OR2_X1 U13193 ( .A1(n13223), .A2(n13224), .ZN(n13084) );
  AND2_X1 U13194 ( .A1(n13078), .A2(n13081), .ZN(n13224) );
  AND2_X1 U13195 ( .A1(n13225), .A2(n13080), .ZN(n13223) );
  OR2_X1 U13196 ( .A1(n13226), .A2(n13227), .ZN(n13080) );
  AND2_X1 U13197 ( .A1(n13074), .A2(n13077), .ZN(n13227) );
  AND2_X1 U13198 ( .A1(n13228), .A2(n13076), .ZN(n13226) );
  OR2_X1 U13199 ( .A1(n13229), .A2(n13230), .ZN(n13076) );
  AND2_X1 U13200 ( .A1(n13071), .A2(n13072), .ZN(n13230) );
  AND2_X1 U13201 ( .A1(n13231), .A2(n13232), .ZN(n13229) );
  OR2_X1 U13202 ( .A1(n13072), .A2(n13071), .ZN(n13232) );
  OR2_X1 U13203 ( .A1(n7912), .A2(n8515), .ZN(n13071) );
  OR2_X1 U13204 ( .A1(n7857), .A2(n13233), .ZN(n13072) );
  OR2_X1 U13205 ( .A1(n7912), .A2(n8956), .ZN(n13233) );
  INV_X1 U13206 ( .A(n13073), .ZN(n13231) );
  OR2_X1 U13207 ( .A1(n13234), .A2(n13235), .ZN(n13073) );
  AND2_X1 U13208 ( .A1(b_8_), .A2(n13236), .ZN(n13235) );
  OR2_X1 U13209 ( .A1(n13237), .A2(n7343), .ZN(n13236) );
  AND2_X1 U13210 ( .A1(a_30_), .A2(n7798), .ZN(n13237) );
  AND2_X1 U13211 ( .A1(b_7_), .A2(n13238), .ZN(n13234) );
  OR2_X1 U13212 ( .A1(n13239), .A2(n7347), .ZN(n13238) );
  AND2_X1 U13213 ( .A1(a_31_), .A2(n7857), .ZN(n13239) );
  OR2_X1 U13214 ( .A1(n13077), .A2(n13074), .ZN(n13228) );
  XOR2_X1 U13215 ( .A(n13240), .B(n13241), .Z(n13074) );
  XNOR2_X1 U13216 ( .A(n13242), .B(n13243), .ZN(n13240) );
  OR2_X1 U13217 ( .A1(n7912), .A2(n8523), .ZN(n13077) );
  OR2_X1 U13218 ( .A1(n13081), .A2(n13078), .ZN(n13225) );
  XOR2_X1 U13219 ( .A(n13244), .B(n13245), .Z(n13078) );
  XOR2_X1 U13220 ( .A(n13246), .B(n13247), .Z(n13245) );
  OR2_X1 U13221 ( .A1(n7912), .A2(n8528), .ZN(n13081) );
  OR2_X1 U13222 ( .A1(n13085), .A2(n13082), .ZN(n13222) );
  XOR2_X1 U13223 ( .A(n13248), .B(n13249), .Z(n13082) );
  XOR2_X1 U13224 ( .A(n13250), .B(n13251), .Z(n13249) );
  OR2_X1 U13225 ( .A1(n7912), .A2(n8533), .ZN(n13085) );
  OR2_X1 U13226 ( .A1(n13089), .A2(n13086), .ZN(n13219) );
  XOR2_X1 U13227 ( .A(n13252), .B(n13253), .Z(n13086) );
  XOR2_X1 U13228 ( .A(n13254), .B(n13255), .Z(n13253) );
  OR2_X1 U13229 ( .A1(n7912), .A2(n8538), .ZN(n13089) );
  OR2_X1 U13230 ( .A1(n13093), .A2(n13090), .ZN(n13216) );
  XOR2_X1 U13231 ( .A(n13256), .B(n13257), .Z(n13090) );
  XOR2_X1 U13232 ( .A(n13258), .B(n13259), .Z(n13257) );
  OR2_X1 U13233 ( .A1(n7912), .A2(n8543), .ZN(n13093) );
  OR2_X1 U13234 ( .A1(n13097), .A2(n13094), .ZN(n13213) );
  XOR2_X1 U13235 ( .A(n13260), .B(n13261), .Z(n13094) );
  XOR2_X1 U13236 ( .A(n13262), .B(n13263), .Z(n13261) );
  OR2_X1 U13237 ( .A1(n7912), .A2(n8548), .ZN(n13097) );
  OR2_X1 U13238 ( .A1(n13101), .A2(n13098), .ZN(n13210) );
  XOR2_X1 U13239 ( .A(n13264), .B(n13265), .Z(n13098) );
  XOR2_X1 U13240 ( .A(n13266), .B(n13267), .Z(n13265) );
  OR2_X1 U13241 ( .A1(n7912), .A2(n8553), .ZN(n13101) );
  XOR2_X1 U13242 ( .A(n13268), .B(n13269), .Z(n13102) );
  XOR2_X1 U13243 ( .A(n13270), .B(n13271), .Z(n13269) );
  OR2_X1 U13244 ( .A1(n13109), .A2(n13106), .ZN(n13204) );
  XOR2_X1 U13245 ( .A(n13272), .B(n13273), .Z(n13106) );
  XOR2_X1 U13246 ( .A(n13274), .B(n13275), .Z(n13273) );
  OR2_X1 U13247 ( .A1(n7912), .A2(n8563), .ZN(n13109) );
  XOR2_X1 U13248 ( .A(n13276), .B(n13277), .Z(n13110) );
  XOR2_X1 U13249 ( .A(n13278), .B(n13279), .Z(n13277) );
  XOR2_X1 U13250 ( .A(n13280), .B(n13281), .Z(n13114) );
  XOR2_X1 U13251 ( .A(n13282), .B(n13283), .Z(n13281) );
  XOR2_X1 U13252 ( .A(n13284), .B(n13285), .Z(n13118) );
  XOR2_X1 U13253 ( .A(n13286), .B(n13287), .Z(n13285) );
  XOR2_X1 U13254 ( .A(n13288), .B(n13289), .Z(n13122) );
  XOR2_X1 U13255 ( .A(n13290), .B(n13291), .Z(n13289) );
  XOR2_X1 U13256 ( .A(n13292), .B(n13293), .Z(n13126) );
  XOR2_X1 U13257 ( .A(n13294), .B(n13295), .Z(n13293) );
  XOR2_X1 U13258 ( .A(n13296), .B(n13297), .Z(n13130) );
  XOR2_X1 U13259 ( .A(n13298), .B(n13299), .Z(n13297) );
  XOR2_X1 U13260 ( .A(n13300), .B(n13301), .Z(n13134) );
  XOR2_X1 U13261 ( .A(n13302), .B(n13303), .Z(n13301) );
  XOR2_X1 U13262 ( .A(n13304), .B(n13305), .Z(n13138) );
  XOR2_X1 U13263 ( .A(n13306), .B(n13307), .Z(n13305) );
  XOR2_X1 U13264 ( .A(n13308), .B(n13309), .Z(n13142) );
  XOR2_X1 U13265 ( .A(n13310), .B(n13311), .Z(n13309) );
  XOR2_X1 U13266 ( .A(n13312), .B(n13313), .Z(n13146) );
  XOR2_X1 U13267 ( .A(n13314), .B(n13315), .Z(n13313) );
  XOR2_X1 U13268 ( .A(n13316), .B(n13317), .Z(n13151) );
  XOR2_X1 U13269 ( .A(n13318), .B(n13319), .Z(n13317) );
  XOR2_X1 U13270 ( .A(n13320), .B(n13321), .Z(n13154) );
  XOR2_X1 U13271 ( .A(n13322), .B(n13323), .Z(n13321) );
  XNOR2_X1 U13272 ( .A(n13324), .B(n13325), .ZN(n13158) );
  XNOR2_X1 U13273 ( .A(n13326), .B(n13327), .ZN(n13324) );
  XOR2_X1 U13274 ( .A(n11765), .B(n13328), .Z(n11758) );
  XOR2_X1 U13275 ( .A(n11764), .B(n11763), .Z(n13328) );
  OR2_X1 U13276 ( .A1(n7857), .A2(n8025), .ZN(n11763) );
  OR2_X1 U13277 ( .A1(n13329), .A2(n13330), .ZN(n11764) );
  AND2_X1 U13278 ( .A1(n13325), .A2(n13327), .ZN(n13330) );
  AND2_X1 U13279 ( .A1(n13331), .A2(n13326), .ZN(n13329) );
  OR2_X1 U13280 ( .A1(n13325), .A2(n13327), .ZN(n13331) );
  OR2_X1 U13281 ( .A1(n13332), .A2(n13333), .ZN(n13327) );
  AND2_X1 U13282 ( .A1(n13323), .A2(n13322), .ZN(n13333) );
  AND2_X1 U13283 ( .A1(n13320), .A2(n13334), .ZN(n13332) );
  OR2_X1 U13284 ( .A1(n13322), .A2(n13323), .ZN(n13334) );
  OR2_X1 U13285 ( .A1(n7857), .A2(n8191), .ZN(n13323) );
  OR2_X1 U13286 ( .A1(n13335), .A2(n13336), .ZN(n13322) );
  AND2_X1 U13287 ( .A1(n13319), .A2(n13318), .ZN(n13336) );
  AND2_X1 U13288 ( .A1(n13316), .A2(n13337), .ZN(n13335) );
  OR2_X1 U13289 ( .A1(n13318), .A2(n13319), .ZN(n13337) );
  OR2_X1 U13290 ( .A1(n7857), .A2(n8287), .ZN(n13319) );
  OR2_X1 U13291 ( .A1(n13338), .A2(n13339), .ZN(n13318) );
  AND2_X1 U13292 ( .A1(n13315), .A2(n13314), .ZN(n13339) );
  AND2_X1 U13293 ( .A1(n13312), .A2(n13340), .ZN(n13338) );
  OR2_X1 U13294 ( .A1(n13314), .A2(n13315), .ZN(n13340) );
  OR2_X1 U13295 ( .A1(n8608), .A2(n7857), .ZN(n13315) );
  OR2_X1 U13296 ( .A1(n13341), .A2(n13342), .ZN(n13314) );
  AND2_X1 U13297 ( .A1(n13311), .A2(n13310), .ZN(n13342) );
  AND2_X1 U13298 ( .A1(n13308), .A2(n13343), .ZN(n13341) );
  OR2_X1 U13299 ( .A1(n13310), .A2(n13311), .ZN(n13343) );
  OR2_X1 U13300 ( .A1(n7857), .A2(n8603), .ZN(n13311) );
  OR2_X1 U13301 ( .A1(n13344), .A2(n13345), .ZN(n13310) );
  AND2_X1 U13302 ( .A1(n13307), .A2(n13306), .ZN(n13345) );
  AND2_X1 U13303 ( .A1(n13304), .A2(n13346), .ZN(n13344) );
  OR2_X1 U13304 ( .A1(n13306), .A2(n13307), .ZN(n13346) );
  OR2_X1 U13305 ( .A1(n7857), .A2(n8598), .ZN(n13307) );
  OR2_X1 U13306 ( .A1(n13347), .A2(n13348), .ZN(n13306) );
  AND2_X1 U13307 ( .A1(n13303), .A2(n13302), .ZN(n13348) );
  AND2_X1 U13308 ( .A1(n13300), .A2(n13349), .ZN(n13347) );
  OR2_X1 U13309 ( .A1(n13302), .A2(n13303), .ZN(n13349) );
  OR2_X1 U13310 ( .A1(n7857), .A2(n8593), .ZN(n13303) );
  OR2_X1 U13311 ( .A1(n13350), .A2(n13351), .ZN(n13302) );
  AND2_X1 U13312 ( .A1(n13299), .A2(n13298), .ZN(n13351) );
  AND2_X1 U13313 ( .A1(n13296), .A2(n13352), .ZN(n13350) );
  OR2_X1 U13314 ( .A1(n13298), .A2(n13299), .ZN(n13352) );
  OR2_X1 U13315 ( .A1(n7857), .A2(n8588), .ZN(n13299) );
  OR2_X1 U13316 ( .A1(n13353), .A2(n13354), .ZN(n13298) );
  AND2_X1 U13317 ( .A1(n13295), .A2(n13294), .ZN(n13354) );
  AND2_X1 U13318 ( .A1(n13292), .A2(n13355), .ZN(n13353) );
  OR2_X1 U13319 ( .A1(n13294), .A2(n13295), .ZN(n13355) );
  OR2_X1 U13320 ( .A1(n7857), .A2(n8583), .ZN(n13295) );
  OR2_X1 U13321 ( .A1(n13356), .A2(n13357), .ZN(n13294) );
  AND2_X1 U13322 ( .A1(n13291), .A2(n13290), .ZN(n13357) );
  AND2_X1 U13323 ( .A1(n13288), .A2(n13358), .ZN(n13356) );
  OR2_X1 U13324 ( .A1(n13290), .A2(n13291), .ZN(n13358) );
  OR2_X1 U13325 ( .A1(n7857), .A2(n8578), .ZN(n13291) );
  OR2_X1 U13326 ( .A1(n13359), .A2(n13360), .ZN(n13290) );
  AND2_X1 U13327 ( .A1(n13287), .A2(n13286), .ZN(n13360) );
  AND2_X1 U13328 ( .A1(n13284), .A2(n13361), .ZN(n13359) );
  OR2_X1 U13329 ( .A1(n13286), .A2(n13287), .ZN(n13361) );
  OR2_X1 U13330 ( .A1(n7857), .A2(n8573), .ZN(n13287) );
  OR2_X1 U13331 ( .A1(n13362), .A2(n13363), .ZN(n13286) );
  AND2_X1 U13332 ( .A1(n13283), .A2(n13282), .ZN(n13363) );
  AND2_X1 U13333 ( .A1(n13280), .A2(n13364), .ZN(n13362) );
  OR2_X1 U13334 ( .A1(n13282), .A2(n13283), .ZN(n13364) );
  OR2_X1 U13335 ( .A1(n7857), .A2(n8568), .ZN(n13283) );
  OR2_X1 U13336 ( .A1(n13365), .A2(n13366), .ZN(n13282) );
  AND2_X1 U13337 ( .A1(n13279), .A2(n13278), .ZN(n13366) );
  AND2_X1 U13338 ( .A1(n13276), .A2(n13367), .ZN(n13365) );
  OR2_X1 U13339 ( .A1(n13278), .A2(n13279), .ZN(n13367) );
  OR2_X1 U13340 ( .A1(n7857), .A2(n8563), .ZN(n13279) );
  OR2_X1 U13341 ( .A1(n13368), .A2(n13369), .ZN(n13278) );
  AND2_X1 U13342 ( .A1(n13272), .A2(n13275), .ZN(n13369) );
  AND2_X1 U13343 ( .A1(n13370), .A2(n13274), .ZN(n13368) );
  OR2_X1 U13344 ( .A1(n13371), .A2(n13372), .ZN(n13274) );
  AND2_X1 U13345 ( .A1(n13271), .A2(n13270), .ZN(n13372) );
  AND2_X1 U13346 ( .A1(n13268), .A2(n13373), .ZN(n13371) );
  OR2_X1 U13347 ( .A1(n13270), .A2(n13271), .ZN(n13373) );
  OR2_X1 U13348 ( .A1(n7857), .A2(n8553), .ZN(n13271) );
  OR2_X1 U13349 ( .A1(n13374), .A2(n13375), .ZN(n13270) );
  AND2_X1 U13350 ( .A1(n13264), .A2(n13267), .ZN(n13375) );
  AND2_X1 U13351 ( .A1(n13376), .A2(n13266), .ZN(n13374) );
  OR2_X1 U13352 ( .A1(n13377), .A2(n13378), .ZN(n13266) );
  AND2_X1 U13353 ( .A1(n13260), .A2(n13263), .ZN(n13378) );
  AND2_X1 U13354 ( .A1(n13379), .A2(n13262), .ZN(n13377) );
  OR2_X1 U13355 ( .A1(n13380), .A2(n13381), .ZN(n13262) );
  AND2_X1 U13356 ( .A1(n13256), .A2(n13259), .ZN(n13381) );
  AND2_X1 U13357 ( .A1(n13382), .A2(n13258), .ZN(n13380) );
  OR2_X1 U13358 ( .A1(n13383), .A2(n13384), .ZN(n13258) );
  AND2_X1 U13359 ( .A1(n13252), .A2(n13255), .ZN(n13384) );
  AND2_X1 U13360 ( .A1(n13385), .A2(n13254), .ZN(n13383) );
  OR2_X1 U13361 ( .A1(n13386), .A2(n13387), .ZN(n13254) );
  AND2_X1 U13362 ( .A1(n13248), .A2(n13251), .ZN(n13387) );
  AND2_X1 U13363 ( .A1(n13388), .A2(n13250), .ZN(n13386) );
  OR2_X1 U13364 ( .A1(n13389), .A2(n13390), .ZN(n13250) );
  AND2_X1 U13365 ( .A1(n13244), .A2(n13247), .ZN(n13390) );
  AND2_X1 U13366 ( .A1(n13391), .A2(n13246), .ZN(n13389) );
  OR2_X1 U13367 ( .A1(n13392), .A2(n13393), .ZN(n13246) );
  AND2_X1 U13368 ( .A1(n13241), .A2(n13242), .ZN(n13393) );
  AND2_X1 U13369 ( .A1(n13394), .A2(n13395), .ZN(n13392) );
  OR2_X1 U13370 ( .A1(n13242), .A2(n13241), .ZN(n13395) );
  OR2_X1 U13371 ( .A1(n8515), .A2(n7857), .ZN(n13241) );
  OR2_X1 U13372 ( .A1(n7798), .A2(n13396), .ZN(n13242) );
  OR2_X1 U13373 ( .A1(n8956), .A2(n7857), .ZN(n13396) );
  INV_X1 U13374 ( .A(n13243), .ZN(n13394) );
  OR2_X1 U13375 ( .A1(n13397), .A2(n13398), .ZN(n13243) );
  AND2_X1 U13376 ( .A1(b_7_), .A2(n13399), .ZN(n13398) );
  OR2_X1 U13377 ( .A1(n13400), .A2(n7343), .ZN(n13399) );
  AND2_X1 U13378 ( .A1(a_30_), .A2(n7759), .ZN(n13400) );
  AND2_X1 U13379 ( .A1(b_6_), .A2(n13401), .ZN(n13397) );
  OR2_X1 U13380 ( .A1(n13402), .A2(n7347), .ZN(n13401) );
  AND2_X1 U13381 ( .A1(a_31_), .A2(n7798), .ZN(n13402) );
  OR2_X1 U13382 ( .A1(n13247), .A2(n13244), .ZN(n13391) );
  XOR2_X1 U13383 ( .A(n13403), .B(n13404), .Z(n13244) );
  XNOR2_X1 U13384 ( .A(n13405), .B(n13406), .ZN(n13403) );
  OR2_X1 U13385 ( .A1(n8523), .A2(n7857), .ZN(n13247) );
  OR2_X1 U13386 ( .A1(n13251), .A2(n13248), .ZN(n13388) );
  XOR2_X1 U13387 ( .A(n13407), .B(n13408), .Z(n13248) );
  XOR2_X1 U13388 ( .A(n13409), .B(n13410), .Z(n13408) );
  OR2_X1 U13389 ( .A1(n7857), .A2(n8528), .ZN(n13251) );
  OR2_X1 U13390 ( .A1(n13255), .A2(n13252), .ZN(n13385) );
  XOR2_X1 U13391 ( .A(n13411), .B(n13412), .Z(n13252) );
  XOR2_X1 U13392 ( .A(n13413), .B(n13414), .Z(n13412) );
  OR2_X1 U13393 ( .A1(n7857), .A2(n8533), .ZN(n13255) );
  OR2_X1 U13394 ( .A1(n13259), .A2(n13256), .ZN(n13382) );
  XOR2_X1 U13395 ( .A(n13415), .B(n13416), .Z(n13256) );
  XOR2_X1 U13396 ( .A(n13417), .B(n13418), .Z(n13416) );
  OR2_X1 U13397 ( .A1(n7857), .A2(n8538), .ZN(n13259) );
  OR2_X1 U13398 ( .A1(n13263), .A2(n13260), .ZN(n13379) );
  XOR2_X1 U13399 ( .A(n13419), .B(n13420), .Z(n13260) );
  XOR2_X1 U13400 ( .A(n13421), .B(n13422), .Z(n13420) );
  OR2_X1 U13401 ( .A1(n7857), .A2(n8543), .ZN(n13263) );
  OR2_X1 U13402 ( .A1(n13267), .A2(n13264), .ZN(n13376) );
  XOR2_X1 U13403 ( .A(n13423), .B(n13424), .Z(n13264) );
  XOR2_X1 U13404 ( .A(n13425), .B(n13426), .Z(n13424) );
  OR2_X1 U13405 ( .A1(n7857), .A2(n8548), .ZN(n13267) );
  XOR2_X1 U13406 ( .A(n13427), .B(n13428), .Z(n13268) );
  XOR2_X1 U13407 ( .A(n13429), .B(n13430), .Z(n13428) );
  OR2_X1 U13408 ( .A1(n13275), .A2(n13272), .ZN(n13370) );
  XOR2_X1 U13409 ( .A(n13431), .B(n13432), .Z(n13272) );
  XOR2_X1 U13410 ( .A(n13433), .B(n13434), .Z(n13432) );
  OR2_X1 U13411 ( .A1(n7857), .A2(n8558), .ZN(n13275) );
  XOR2_X1 U13412 ( .A(n13435), .B(n13436), .Z(n13276) );
  XOR2_X1 U13413 ( .A(n13437), .B(n13438), .Z(n13436) );
  XOR2_X1 U13414 ( .A(n13439), .B(n13440), .Z(n13280) );
  XOR2_X1 U13415 ( .A(n13441), .B(n13442), .Z(n13440) );
  XOR2_X1 U13416 ( .A(n13443), .B(n13444), .Z(n13284) );
  XOR2_X1 U13417 ( .A(n13445), .B(n13446), .Z(n13444) );
  XOR2_X1 U13418 ( .A(n13447), .B(n13448), .Z(n13288) );
  XOR2_X1 U13419 ( .A(n13449), .B(n13450), .Z(n13448) );
  XOR2_X1 U13420 ( .A(n13451), .B(n13452), .Z(n13292) );
  XOR2_X1 U13421 ( .A(n13453), .B(n13454), .Z(n13452) );
  XOR2_X1 U13422 ( .A(n13455), .B(n13456), .Z(n13296) );
  XOR2_X1 U13423 ( .A(n13457), .B(n13458), .Z(n13456) );
  XOR2_X1 U13424 ( .A(n13459), .B(n13460), .Z(n13300) );
  XOR2_X1 U13425 ( .A(n13461), .B(n13462), .Z(n13460) );
  XOR2_X1 U13426 ( .A(n13463), .B(n13464), .Z(n13304) );
  XOR2_X1 U13427 ( .A(n13465), .B(n13466), .Z(n13464) );
  XOR2_X1 U13428 ( .A(n13467), .B(n13468), .Z(n13308) );
  XOR2_X1 U13429 ( .A(n13469), .B(n13470), .Z(n13468) );
  XOR2_X1 U13430 ( .A(n13471), .B(n13472), .Z(n13312) );
  XOR2_X1 U13431 ( .A(n13473), .B(n13474), .Z(n13472) );
  XOR2_X1 U13432 ( .A(n13475), .B(n13476), .Z(n13316) );
  XOR2_X1 U13433 ( .A(n13477), .B(n13478), .Z(n13476) );
  XOR2_X1 U13434 ( .A(n13479), .B(n13480), .Z(n13320) );
  XOR2_X1 U13435 ( .A(n13481), .B(n13482), .Z(n13480) );
  XOR2_X1 U13436 ( .A(n13483), .B(n13484), .Z(n13325) );
  XOR2_X1 U13437 ( .A(n13485), .B(n13486), .Z(n13484) );
  XOR2_X1 U13438 ( .A(n11804), .B(n13487), .Z(n11765) );
  XOR2_X1 U13439 ( .A(n11803), .B(n11802), .Z(n13487) );
  OR2_X1 U13440 ( .A1(n7798), .A2(n8107), .ZN(n11802) );
  OR2_X1 U13441 ( .A1(n13488), .A2(n13489), .ZN(n11803) );
  AND2_X1 U13442 ( .A1(n13486), .A2(n13485), .ZN(n13489) );
  AND2_X1 U13443 ( .A1(n13483), .A2(n13490), .ZN(n13488) );
  OR2_X1 U13444 ( .A1(n13485), .A2(n13486), .ZN(n13490) );
  OR2_X1 U13445 ( .A1(n7798), .A2(n8191), .ZN(n13486) );
  OR2_X1 U13446 ( .A1(n13491), .A2(n13492), .ZN(n13485) );
  AND2_X1 U13447 ( .A1(n13482), .A2(n13481), .ZN(n13492) );
  AND2_X1 U13448 ( .A1(n13479), .A2(n13493), .ZN(n13491) );
  OR2_X1 U13449 ( .A1(n13481), .A2(n13482), .ZN(n13493) );
  OR2_X1 U13450 ( .A1(n7798), .A2(n8287), .ZN(n13482) );
  OR2_X1 U13451 ( .A1(n13494), .A2(n13495), .ZN(n13481) );
  AND2_X1 U13452 ( .A1(n13478), .A2(n13477), .ZN(n13495) );
  AND2_X1 U13453 ( .A1(n13475), .A2(n13496), .ZN(n13494) );
  OR2_X1 U13454 ( .A1(n13477), .A2(n13478), .ZN(n13496) );
  OR2_X1 U13455 ( .A1(n8608), .A2(n7798), .ZN(n13478) );
  OR2_X1 U13456 ( .A1(n13497), .A2(n13498), .ZN(n13477) );
  AND2_X1 U13457 ( .A1(n13474), .A2(n13473), .ZN(n13498) );
  AND2_X1 U13458 ( .A1(n13471), .A2(n13499), .ZN(n13497) );
  OR2_X1 U13459 ( .A1(n13473), .A2(n13474), .ZN(n13499) );
  OR2_X1 U13460 ( .A1(n7798), .A2(n8603), .ZN(n13474) );
  OR2_X1 U13461 ( .A1(n13500), .A2(n13501), .ZN(n13473) );
  AND2_X1 U13462 ( .A1(n13470), .A2(n13469), .ZN(n13501) );
  AND2_X1 U13463 ( .A1(n13467), .A2(n13502), .ZN(n13500) );
  OR2_X1 U13464 ( .A1(n13469), .A2(n13470), .ZN(n13502) );
  OR2_X1 U13465 ( .A1(n7798), .A2(n8598), .ZN(n13470) );
  OR2_X1 U13466 ( .A1(n13503), .A2(n13504), .ZN(n13469) );
  AND2_X1 U13467 ( .A1(n13466), .A2(n13465), .ZN(n13504) );
  AND2_X1 U13468 ( .A1(n13463), .A2(n13505), .ZN(n13503) );
  OR2_X1 U13469 ( .A1(n13465), .A2(n13466), .ZN(n13505) );
  OR2_X1 U13470 ( .A1(n7798), .A2(n8593), .ZN(n13466) );
  OR2_X1 U13471 ( .A1(n13506), .A2(n13507), .ZN(n13465) );
  AND2_X1 U13472 ( .A1(n13462), .A2(n13461), .ZN(n13507) );
  AND2_X1 U13473 ( .A1(n13459), .A2(n13508), .ZN(n13506) );
  OR2_X1 U13474 ( .A1(n13461), .A2(n13462), .ZN(n13508) );
  OR2_X1 U13475 ( .A1(n7798), .A2(n8588), .ZN(n13462) );
  OR2_X1 U13476 ( .A1(n13509), .A2(n13510), .ZN(n13461) );
  AND2_X1 U13477 ( .A1(n13458), .A2(n13457), .ZN(n13510) );
  AND2_X1 U13478 ( .A1(n13455), .A2(n13511), .ZN(n13509) );
  OR2_X1 U13479 ( .A1(n13457), .A2(n13458), .ZN(n13511) );
  OR2_X1 U13480 ( .A1(n7798), .A2(n8583), .ZN(n13458) );
  OR2_X1 U13481 ( .A1(n13512), .A2(n13513), .ZN(n13457) );
  AND2_X1 U13482 ( .A1(n13454), .A2(n13453), .ZN(n13513) );
  AND2_X1 U13483 ( .A1(n13451), .A2(n13514), .ZN(n13512) );
  OR2_X1 U13484 ( .A1(n13453), .A2(n13454), .ZN(n13514) );
  OR2_X1 U13485 ( .A1(n7798), .A2(n8578), .ZN(n13454) );
  OR2_X1 U13486 ( .A1(n13515), .A2(n13516), .ZN(n13453) );
  AND2_X1 U13487 ( .A1(n13450), .A2(n13449), .ZN(n13516) );
  AND2_X1 U13488 ( .A1(n13447), .A2(n13517), .ZN(n13515) );
  OR2_X1 U13489 ( .A1(n13449), .A2(n13450), .ZN(n13517) );
  OR2_X1 U13490 ( .A1(n7798), .A2(n8573), .ZN(n13450) );
  OR2_X1 U13491 ( .A1(n13518), .A2(n13519), .ZN(n13449) );
  AND2_X1 U13492 ( .A1(n13446), .A2(n13445), .ZN(n13519) );
  AND2_X1 U13493 ( .A1(n13443), .A2(n13520), .ZN(n13518) );
  OR2_X1 U13494 ( .A1(n13445), .A2(n13446), .ZN(n13520) );
  OR2_X1 U13495 ( .A1(n7798), .A2(n8568), .ZN(n13446) );
  OR2_X1 U13496 ( .A1(n13521), .A2(n13522), .ZN(n13445) );
  AND2_X1 U13497 ( .A1(n13442), .A2(n13441), .ZN(n13522) );
  AND2_X1 U13498 ( .A1(n13439), .A2(n13523), .ZN(n13521) );
  OR2_X1 U13499 ( .A1(n13441), .A2(n13442), .ZN(n13523) );
  OR2_X1 U13500 ( .A1(n7798), .A2(n8563), .ZN(n13442) );
  OR2_X1 U13501 ( .A1(n13524), .A2(n13525), .ZN(n13441) );
  AND2_X1 U13502 ( .A1(n13438), .A2(n13437), .ZN(n13525) );
  AND2_X1 U13503 ( .A1(n13435), .A2(n13526), .ZN(n13524) );
  OR2_X1 U13504 ( .A1(n13437), .A2(n13438), .ZN(n13526) );
  OR2_X1 U13505 ( .A1(n7798), .A2(n8558), .ZN(n13438) );
  OR2_X1 U13506 ( .A1(n13527), .A2(n13528), .ZN(n13437) );
  AND2_X1 U13507 ( .A1(n13431), .A2(n13434), .ZN(n13528) );
  AND2_X1 U13508 ( .A1(n13529), .A2(n13433), .ZN(n13527) );
  OR2_X1 U13509 ( .A1(n13530), .A2(n13531), .ZN(n13433) );
  AND2_X1 U13510 ( .A1(n13430), .A2(n13429), .ZN(n13531) );
  AND2_X1 U13511 ( .A1(n13427), .A2(n13532), .ZN(n13530) );
  OR2_X1 U13512 ( .A1(n13429), .A2(n13430), .ZN(n13532) );
  OR2_X1 U13513 ( .A1(n7798), .A2(n8548), .ZN(n13430) );
  OR2_X1 U13514 ( .A1(n13533), .A2(n13534), .ZN(n13429) );
  AND2_X1 U13515 ( .A1(n13423), .A2(n13426), .ZN(n13534) );
  AND2_X1 U13516 ( .A1(n13535), .A2(n13425), .ZN(n13533) );
  OR2_X1 U13517 ( .A1(n13536), .A2(n13537), .ZN(n13425) );
  AND2_X1 U13518 ( .A1(n13419), .A2(n13422), .ZN(n13537) );
  AND2_X1 U13519 ( .A1(n13538), .A2(n13421), .ZN(n13536) );
  OR2_X1 U13520 ( .A1(n13539), .A2(n13540), .ZN(n13421) );
  AND2_X1 U13521 ( .A1(n13415), .A2(n13418), .ZN(n13540) );
  AND2_X1 U13522 ( .A1(n13541), .A2(n13417), .ZN(n13539) );
  OR2_X1 U13523 ( .A1(n13542), .A2(n13543), .ZN(n13417) );
  AND2_X1 U13524 ( .A1(n13411), .A2(n13414), .ZN(n13543) );
  AND2_X1 U13525 ( .A1(n13544), .A2(n13413), .ZN(n13542) );
  OR2_X1 U13526 ( .A1(n13545), .A2(n13546), .ZN(n13413) );
  AND2_X1 U13527 ( .A1(n13407), .A2(n13410), .ZN(n13546) );
  AND2_X1 U13528 ( .A1(n13547), .A2(n13409), .ZN(n13545) );
  OR2_X1 U13529 ( .A1(n13548), .A2(n13549), .ZN(n13409) );
  AND2_X1 U13530 ( .A1(n13404), .A2(n13405), .ZN(n13549) );
  AND2_X1 U13531 ( .A1(n13550), .A2(n13551), .ZN(n13548) );
  OR2_X1 U13532 ( .A1(n13405), .A2(n13404), .ZN(n13551) );
  OR2_X1 U13533 ( .A1(n8515), .A2(n7798), .ZN(n13404) );
  OR2_X1 U13534 ( .A1(n7759), .A2(n13552), .ZN(n13405) );
  OR2_X1 U13535 ( .A1(n8956), .A2(n7798), .ZN(n13552) );
  INV_X1 U13536 ( .A(n13406), .ZN(n13550) );
  OR2_X1 U13537 ( .A1(n13553), .A2(n13554), .ZN(n13406) );
  AND2_X1 U13538 ( .A1(b_6_), .A2(n13555), .ZN(n13554) );
  OR2_X1 U13539 ( .A1(n13556), .A2(n7343), .ZN(n13555) );
  AND2_X1 U13540 ( .A1(a_30_), .A2(n7715), .ZN(n13556) );
  AND2_X1 U13541 ( .A1(b_5_), .A2(n13557), .ZN(n13553) );
  OR2_X1 U13542 ( .A1(n13558), .A2(n7347), .ZN(n13557) );
  AND2_X1 U13543 ( .A1(a_31_), .A2(n7759), .ZN(n13558) );
  OR2_X1 U13544 ( .A1(n13410), .A2(n13407), .ZN(n13547) );
  XOR2_X1 U13545 ( .A(n13559), .B(n13560), .Z(n13407) );
  XNOR2_X1 U13546 ( .A(n13561), .B(n13562), .ZN(n13559) );
  OR2_X1 U13547 ( .A1(n8523), .A2(n7798), .ZN(n13410) );
  OR2_X1 U13548 ( .A1(n13414), .A2(n13411), .ZN(n13544) );
  XOR2_X1 U13549 ( .A(n13563), .B(n13564), .Z(n13411) );
  XOR2_X1 U13550 ( .A(n13565), .B(n13566), .Z(n13564) );
  OR2_X1 U13551 ( .A1(n8528), .A2(n7798), .ZN(n13414) );
  OR2_X1 U13552 ( .A1(n13418), .A2(n13415), .ZN(n13541) );
  XOR2_X1 U13553 ( .A(n13567), .B(n13568), .Z(n13415) );
  XOR2_X1 U13554 ( .A(n13569), .B(n13570), .Z(n13568) );
  OR2_X1 U13555 ( .A1(n7798), .A2(n8533), .ZN(n13418) );
  OR2_X1 U13556 ( .A1(n13422), .A2(n13419), .ZN(n13538) );
  XOR2_X1 U13557 ( .A(n13571), .B(n13572), .Z(n13419) );
  XOR2_X1 U13558 ( .A(n13573), .B(n13574), .Z(n13572) );
  OR2_X1 U13559 ( .A1(n7798), .A2(n8538), .ZN(n13422) );
  OR2_X1 U13560 ( .A1(n13426), .A2(n13423), .ZN(n13535) );
  XOR2_X1 U13561 ( .A(n13575), .B(n13576), .Z(n13423) );
  XOR2_X1 U13562 ( .A(n13577), .B(n13578), .Z(n13576) );
  OR2_X1 U13563 ( .A1(n7798), .A2(n8543), .ZN(n13426) );
  XOR2_X1 U13564 ( .A(n13579), .B(n13580), .Z(n13427) );
  XOR2_X1 U13565 ( .A(n13581), .B(n13582), .Z(n13580) );
  OR2_X1 U13566 ( .A1(n13434), .A2(n13431), .ZN(n13529) );
  XOR2_X1 U13567 ( .A(n13583), .B(n13584), .Z(n13431) );
  XOR2_X1 U13568 ( .A(n13585), .B(n13586), .Z(n13584) );
  OR2_X1 U13569 ( .A1(n7798), .A2(n8553), .ZN(n13434) );
  XOR2_X1 U13570 ( .A(n13587), .B(n13588), .Z(n13435) );
  XOR2_X1 U13571 ( .A(n13589), .B(n13590), .Z(n13588) );
  XOR2_X1 U13572 ( .A(n13591), .B(n13592), .Z(n13439) );
  XOR2_X1 U13573 ( .A(n13593), .B(n13594), .Z(n13592) );
  XOR2_X1 U13574 ( .A(n13595), .B(n13596), .Z(n13443) );
  XOR2_X1 U13575 ( .A(n13597), .B(n13598), .Z(n13596) );
  XOR2_X1 U13576 ( .A(n13599), .B(n13600), .Z(n13447) );
  XOR2_X1 U13577 ( .A(n13601), .B(n13602), .Z(n13600) );
  XOR2_X1 U13578 ( .A(n13603), .B(n13604), .Z(n13451) );
  XOR2_X1 U13579 ( .A(n13605), .B(n13606), .Z(n13604) );
  XOR2_X1 U13580 ( .A(n13607), .B(n13608), .Z(n13455) );
  XOR2_X1 U13581 ( .A(n13609), .B(n13610), .Z(n13608) );
  XOR2_X1 U13582 ( .A(n13611), .B(n13612), .Z(n13459) );
  XOR2_X1 U13583 ( .A(n13613), .B(n13614), .Z(n13612) );
  XOR2_X1 U13584 ( .A(n13615), .B(n13616), .Z(n13463) );
  XOR2_X1 U13585 ( .A(n13617), .B(n13618), .Z(n13616) );
  XOR2_X1 U13586 ( .A(n13619), .B(n13620), .Z(n13467) );
  XOR2_X1 U13587 ( .A(n13621), .B(n13622), .Z(n13620) );
  XOR2_X1 U13588 ( .A(n13623), .B(n13624), .Z(n13471) );
  XOR2_X1 U13589 ( .A(n13625), .B(n13626), .Z(n13624) );
  XOR2_X1 U13590 ( .A(n13627), .B(n13628), .Z(n13475) );
  XOR2_X1 U13591 ( .A(n13629), .B(n13630), .Z(n13628) );
  XOR2_X1 U13592 ( .A(n13631), .B(n13632), .Z(n13479) );
  XOR2_X1 U13593 ( .A(n13633), .B(n13634), .Z(n13632) );
  XOR2_X1 U13594 ( .A(n13635), .B(n13636), .Z(n13483) );
  XOR2_X1 U13595 ( .A(n13637), .B(n13638), .Z(n13636) );
  XOR2_X1 U13596 ( .A(n11773), .B(n13639), .Z(n11804) );
  XOR2_X1 U13597 ( .A(n11772), .B(n11771), .Z(n13639) );
  OR2_X1 U13598 ( .A1(n7759), .A2(n8191), .ZN(n11771) );
  OR2_X1 U13599 ( .A1(n13640), .A2(n13641), .ZN(n11772) );
  AND2_X1 U13600 ( .A1(n13638), .A2(n13637), .ZN(n13641) );
  AND2_X1 U13601 ( .A1(n13635), .A2(n13642), .ZN(n13640) );
  OR2_X1 U13602 ( .A1(n13637), .A2(n13638), .ZN(n13642) );
  OR2_X1 U13603 ( .A1(n7759), .A2(n8287), .ZN(n13638) );
  OR2_X1 U13604 ( .A1(n13643), .A2(n13644), .ZN(n13637) );
  AND2_X1 U13605 ( .A1(n13634), .A2(n13633), .ZN(n13644) );
  AND2_X1 U13606 ( .A1(n13631), .A2(n13645), .ZN(n13643) );
  OR2_X1 U13607 ( .A1(n13633), .A2(n13634), .ZN(n13645) );
  OR2_X1 U13608 ( .A1(n8608), .A2(n7759), .ZN(n13634) );
  OR2_X1 U13609 ( .A1(n13646), .A2(n13647), .ZN(n13633) );
  AND2_X1 U13610 ( .A1(n13630), .A2(n13629), .ZN(n13647) );
  AND2_X1 U13611 ( .A1(n13627), .A2(n13648), .ZN(n13646) );
  OR2_X1 U13612 ( .A1(n13629), .A2(n13630), .ZN(n13648) );
  OR2_X1 U13613 ( .A1(n7759), .A2(n8603), .ZN(n13630) );
  OR2_X1 U13614 ( .A1(n13649), .A2(n13650), .ZN(n13629) );
  AND2_X1 U13615 ( .A1(n13626), .A2(n13625), .ZN(n13650) );
  AND2_X1 U13616 ( .A1(n13623), .A2(n13651), .ZN(n13649) );
  OR2_X1 U13617 ( .A1(n13625), .A2(n13626), .ZN(n13651) );
  OR2_X1 U13618 ( .A1(n7759), .A2(n8598), .ZN(n13626) );
  OR2_X1 U13619 ( .A1(n13652), .A2(n13653), .ZN(n13625) );
  AND2_X1 U13620 ( .A1(n13622), .A2(n13621), .ZN(n13653) );
  AND2_X1 U13621 ( .A1(n13619), .A2(n13654), .ZN(n13652) );
  OR2_X1 U13622 ( .A1(n13621), .A2(n13622), .ZN(n13654) );
  OR2_X1 U13623 ( .A1(n7759), .A2(n8593), .ZN(n13622) );
  OR2_X1 U13624 ( .A1(n13655), .A2(n13656), .ZN(n13621) );
  AND2_X1 U13625 ( .A1(n13618), .A2(n13617), .ZN(n13656) );
  AND2_X1 U13626 ( .A1(n13615), .A2(n13657), .ZN(n13655) );
  OR2_X1 U13627 ( .A1(n13617), .A2(n13618), .ZN(n13657) );
  OR2_X1 U13628 ( .A1(n7759), .A2(n8588), .ZN(n13618) );
  OR2_X1 U13629 ( .A1(n13658), .A2(n13659), .ZN(n13617) );
  AND2_X1 U13630 ( .A1(n13614), .A2(n13613), .ZN(n13659) );
  AND2_X1 U13631 ( .A1(n13611), .A2(n13660), .ZN(n13658) );
  OR2_X1 U13632 ( .A1(n13613), .A2(n13614), .ZN(n13660) );
  OR2_X1 U13633 ( .A1(n7759), .A2(n8583), .ZN(n13614) );
  OR2_X1 U13634 ( .A1(n13661), .A2(n13662), .ZN(n13613) );
  AND2_X1 U13635 ( .A1(n13610), .A2(n13609), .ZN(n13662) );
  AND2_X1 U13636 ( .A1(n13607), .A2(n13663), .ZN(n13661) );
  OR2_X1 U13637 ( .A1(n13609), .A2(n13610), .ZN(n13663) );
  OR2_X1 U13638 ( .A1(n7759), .A2(n8578), .ZN(n13610) );
  OR2_X1 U13639 ( .A1(n13664), .A2(n13665), .ZN(n13609) );
  AND2_X1 U13640 ( .A1(n13606), .A2(n13605), .ZN(n13665) );
  AND2_X1 U13641 ( .A1(n13603), .A2(n13666), .ZN(n13664) );
  OR2_X1 U13642 ( .A1(n13605), .A2(n13606), .ZN(n13666) );
  OR2_X1 U13643 ( .A1(n7759), .A2(n8573), .ZN(n13606) );
  OR2_X1 U13644 ( .A1(n13667), .A2(n13668), .ZN(n13605) );
  AND2_X1 U13645 ( .A1(n13602), .A2(n13601), .ZN(n13668) );
  AND2_X1 U13646 ( .A1(n13599), .A2(n13669), .ZN(n13667) );
  OR2_X1 U13647 ( .A1(n13601), .A2(n13602), .ZN(n13669) );
  OR2_X1 U13648 ( .A1(n7759), .A2(n8568), .ZN(n13602) );
  OR2_X1 U13649 ( .A1(n13670), .A2(n13671), .ZN(n13601) );
  AND2_X1 U13650 ( .A1(n13598), .A2(n13597), .ZN(n13671) );
  AND2_X1 U13651 ( .A1(n13595), .A2(n13672), .ZN(n13670) );
  OR2_X1 U13652 ( .A1(n13597), .A2(n13598), .ZN(n13672) );
  OR2_X1 U13653 ( .A1(n7759), .A2(n8563), .ZN(n13598) );
  OR2_X1 U13654 ( .A1(n13673), .A2(n13674), .ZN(n13597) );
  AND2_X1 U13655 ( .A1(n13594), .A2(n13593), .ZN(n13674) );
  AND2_X1 U13656 ( .A1(n13591), .A2(n13675), .ZN(n13673) );
  OR2_X1 U13657 ( .A1(n13593), .A2(n13594), .ZN(n13675) );
  OR2_X1 U13658 ( .A1(n7759), .A2(n8558), .ZN(n13594) );
  OR2_X1 U13659 ( .A1(n13676), .A2(n13677), .ZN(n13593) );
  AND2_X1 U13660 ( .A1(n13590), .A2(n13589), .ZN(n13677) );
  AND2_X1 U13661 ( .A1(n13587), .A2(n13678), .ZN(n13676) );
  OR2_X1 U13662 ( .A1(n13589), .A2(n13590), .ZN(n13678) );
  OR2_X1 U13663 ( .A1(n7759), .A2(n8553), .ZN(n13590) );
  OR2_X1 U13664 ( .A1(n13679), .A2(n13680), .ZN(n13589) );
  AND2_X1 U13665 ( .A1(n13583), .A2(n13586), .ZN(n13680) );
  AND2_X1 U13666 ( .A1(n13681), .A2(n13585), .ZN(n13679) );
  OR2_X1 U13667 ( .A1(n13682), .A2(n13683), .ZN(n13585) );
  AND2_X1 U13668 ( .A1(n13582), .A2(n13581), .ZN(n13683) );
  AND2_X1 U13669 ( .A1(n13579), .A2(n13684), .ZN(n13682) );
  OR2_X1 U13670 ( .A1(n13581), .A2(n13582), .ZN(n13684) );
  OR2_X1 U13671 ( .A1(n7759), .A2(n8543), .ZN(n13582) );
  OR2_X1 U13672 ( .A1(n13685), .A2(n13686), .ZN(n13581) );
  AND2_X1 U13673 ( .A1(n13575), .A2(n13578), .ZN(n13686) );
  AND2_X1 U13674 ( .A1(n13687), .A2(n13577), .ZN(n13685) );
  OR2_X1 U13675 ( .A1(n13688), .A2(n13689), .ZN(n13577) );
  AND2_X1 U13676 ( .A1(n13571), .A2(n13574), .ZN(n13689) );
  AND2_X1 U13677 ( .A1(n13690), .A2(n13573), .ZN(n13688) );
  OR2_X1 U13678 ( .A1(n13691), .A2(n13692), .ZN(n13573) );
  AND2_X1 U13679 ( .A1(n13567), .A2(n13570), .ZN(n13692) );
  AND2_X1 U13680 ( .A1(n13693), .A2(n13569), .ZN(n13691) );
  OR2_X1 U13681 ( .A1(n13694), .A2(n13695), .ZN(n13569) );
  AND2_X1 U13682 ( .A1(n13563), .A2(n13566), .ZN(n13695) );
  AND2_X1 U13683 ( .A1(n13696), .A2(n13565), .ZN(n13694) );
  OR2_X1 U13684 ( .A1(n13697), .A2(n13698), .ZN(n13565) );
  AND2_X1 U13685 ( .A1(n13560), .A2(n13561), .ZN(n13698) );
  AND2_X1 U13686 ( .A1(n13699), .A2(n13700), .ZN(n13697) );
  OR2_X1 U13687 ( .A1(n13561), .A2(n13560), .ZN(n13700) );
  OR2_X1 U13688 ( .A1(n8515), .A2(n7759), .ZN(n13560) );
  OR2_X1 U13689 ( .A1(n7715), .A2(n13701), .ZN(n13561) );
  OR2_X1 U13690 ( .A1(n8956), .A2(n7759), .ZN(n13701) );
  INV_X1 U13691 ( .A(n13562), .ZN(n13699) );
  OR2_X1 U13692 ( .A1(n13702), .A2(n13703), .ZN(n13562) );
  AND2_X1 U13693 ( .A1(b_5_), .A2(n13704), .ZN(n13703) );
  OR2_X1 U13694 ( .A1(n13705), .A2(n7343), .ZN(n13704) );
  AND2_X1 U13695 ( .A1(a_30_), .A2(n7689), .ZN(n13705) );
  AND2_X1 U13696 ( .A1(b_4_), .A2(n13706), .ZN(n13702) );
  OR2_X1 U13697 ( .A1(n13707), .A2(n7347), .ZN(n13706) );
  AND2_X1 U13698 ( .A1(a_31_), .A2(n7715), .ZN(n13707) );
  OR2_X1 U13699 ( .A1(n13566), .A2(n13563), .ZN(n13696) );
  XOR2_X1 U13700 ( .A(n13708), .B(n13709), .Z(n13563) );
  XNOR2_X1 U13701 ( .A(n13710), .B(n13711), .ZN(n13708) );
  OR2_X1 U13702 ( .A1(n8523), .A2(n7759), .ZN(n13566) );
  OR2_X1 U13703 ( .A1(n13570), .A2(n13567), .ZN(n13693) );
  XOR2_X1 U13704 ( .A(n13712), .B(n13713), .Z(n13567) );
  XOR2_X1 U13705 ( .A(n13714), .B(n13715), .Z(n13713) );
  OR2_X1 U13706 ( .A1(n8528), .A2(n7759), .ZN(n13570) );
  OR2_X1 U13707 ( .A1(n13574), .A2(n13571), .ZN(n13690) );
  XOR2_X1 U13708 ( .A(n13716), .B(n13717), .Z(n13571) );
  XOR2_X1 U13709 ( .A(n13718), .B(n13719), .Z(n13717) );
  OR2_X1 U13710 ( .A1(n8533), .A2(n7759), .ZN(n13574) );
  OR2_X1 U13711 ( .A1(n13578), .A2(n13575), .ZN(n13687) );
  XOR2_X1 U13712 ( .A(n13720), .B(n13721), .Z(n13575) );
  XOR2_X1 U13713 ( .A(n13722), .B(n13723), .Z(n13721) );
  OR2_X1 U13714 ( .A1(n7759), .A2(n8538), .ZN(n13578) );
  XOR2_X1 U13715 ( .A(n13724), .B(n13725), .Z(n13579) );
  XOR2_X1 U13716 ( .A(n13726), .B(n13727), .Z(n13725) );
  OR2_X1 U13717 ( .A1(n13586), .A2(n13583), .ZN(n13681) );
  XOR2_X1 U13718 ( .A(n13728), .B(n13729), .Z(n13583) );
  XOR2_X1 U13719 ( .A(n13730), .B(n13731), .Z(n13729) );
  OR2_X1 U13720 ( .A1(n7759), .A2(n8548), .ZN(n13586) );
  XOR2_X1 U13721 ( .A(n13732), .B(n13733), .Z(n13587) );
  XOR2_X1 U13722 ( .A(n13734), .B(n13735), .Z(n13733) );
  XOR2_X1 U13723 ( .A(n13736), .B(n13737), .Z(n13591) );
  XOR2_X1 U13724 ( .A(n13738), .B(n13739), .Z(n13737) );
  XOR2_X1 U13725 ( .A(n13740), .B(n13741), .Z(n13595) );
  XOR2_X1 U13726 ( .A(n13742), .B(n13743), .Z(n13741) );
  XOR2_X1 U13727 ( .A(n13744), .B(n13745), .Z(n13599) );
  XOR2_X1 U13728 ( .A(n13746), .B(n13747), .Z(n13745) );
  XOR2_X1 U13729 ( .A(n13748), .B(n13749), .Z(n13603) );
  XOR2_X1 U13730 ( .A(n13750), .B(n13751), .Z(n13749) );
  XOR2_X1 U13731 ( .A(n13752), .B(n13753), .Z(n13607) );
  XOR2_X1 U13732 ( .A(n13754), .B(n13755), .Z(n13753) );
  XOR2_X1 U13733 ( .A(n13756), .B(n13757), .Z(n13611) );
  XOR2_X1 U13734 ( .A(n13758), .B(n13759), .Z(n13757) );
  XOR2_X1 U13735 ( .A(n13760), .B(n13761), .Z(n13615) );
  XOR2_X1 U13736 ( .A(n13762), .B(n13763), .Z(n13761) );
  XOR2_X1 U13737 ( .A(n13764), .B(n13765), .Z(n13619) );
  XOR2_X1 U13738 ( .A(n13766), .B(n13767), .Z(n13765) );
  XOR2_X1 U13739 ( .A(n13768), .B(n13769), .Z(n13623) );
  XOR2_X1 U13740 ( .A(n13770), .B(n13771), .Z(n13769) );
  XOR2_X1 U13741 ( .A(n13772), .B(n13773), .Z(n13627) );
  XOR2_X1 U13742 ( .A(n13774), .B(n13775), .Z(n13773) );
  XOR2_X1 U13743 ( .A(n13776), .B(n13777), .Z(n13631) );
  XOR2_X1 U13744 ( .A(n13778), .B(n13779), .Z(n13777) );
  XOR2_X1 U13745 ( .A(n13780), .B(n13781), .Z(n13635) );
  XOR2_X1 U13746 ( .A(n13782), .B(n13783), .Z(n13781) );
  XOR2_X1 U13747 ( .A(n11780), .B(n13784), .Z(n11773) );
  XOR2_X1 U13748 ( .A(n11779), .B(n11778), .Z(n13784) );
  OR2_X1 U13749 ( .A1(n7715), .A2(n8287), .ZN(n11778) );
  OR2_X1 U13750 ( .A1(n13785), .A2(n13786), .ZN(n11779) );
  AND2_X1 U13751 ( .A1(n13783), .A2(n13782), .ZN(n13786) );
  AND2_X1 U13752 ( .A1(n13780), .A2(n13787), .ZN(n13785) );
  OR2_X1 U13753 ( .A1(n13782), .A2(n13783), .ZN(n13787) );
  OR2_X1 U13754 ( .A1(n8608), .A2(n7715), .ZN(n13783) );
  OR2_X1 U13755 ( .A1(n13788), .A2(n13789), .ZN(n13782) );
  AND2_X1 U13756 ( .A1(n13779), .A2(n13778), .ZN(n13789) );
  AND2_X1 U13757 ( .A1(n13776), .A2(n13790), .ZN(n13788) );
  OR2_X1 U13758 ( .A1(n13778), .A2(n13779), .ZN(n13790) );
  OR2_X1 U13759 ( .A1(n7715), .A2(n8603), .ZN(n13779) );
  OR2_X1 U13760 ( .A1(n13791), .A2(n13792), .ZN(n13778) );
  AND2_X1 U13761 ( .A1(n13775), .A2(n13774), .ZN(n13792) );
  AND2_X1 U13762 ( .A1(n13772), .A2(n13793), .ZN(n13791) );
  OR2_X1 U13763 ( .A1(n13774), .A2(n13775), .ZN(n13793) );
  OR2_X1 U13764 ( .A1(n7715), .A2(n8598), .ZN(n13775) );
  OR2_X1 U13765 ( .A1(n13794), .A2(n13795), .ZN(n13774) );
  AND2_X1 U13766 ( .A1(n13771), .A2(n13770), .ZN(n13795) );
  AND2_X1 U13767 ( .A1(n13768), .A2(n13796), .ZN(n13794) );
  OR2_X1 U13768 ( .A1(n13770), .A2(n13771), .ZN(n13796) );
  OR2_X1 U13769 ( .A1(n7715), .A2(n8593), .ZN(n13771) );
  OR2_X1 U13770 ( .A1(n13797), .A2(n13798), .ZN(n13770) );
  AND2_X1 U13771 ( .A1(n13767), .A2(n13766), .ZN(n13798) );
  AND2_X1 U13772 ( .A1(n13764), .A2(n13799), .ZN(n13797) );
  OR2_X1 U13773 ( .A1(n13766), .A2(n13767), .ZN(n13799) );
  OR2_X1 U13774 ( .A1(n7715), .A2(n8588), .ZN(n13767) );
  OR2_X1 U13775 ( .A1(n13800), .A2(n13801), .ZN(n13766) );
  AND2_X1 U13776 ( .A1(n13763), .A2(n13762), .ZN(n13801) );
  AND2_X1 U13777 ( .A1(n13760), .A2(n13802), .ZN(n13800) );
  OR2_X1 U13778 ( .A1(n13762), .A2(n13763), .ZN(n13802) );
  OR2_X1 U13779 ( .A1(n7715), .A2(n8583), .ZN(n13763) );
  OR2_X1 U13780 ( .A1(n13803), .A2(n13804), .ZN(n13762) );
  AND2_X1 U13781 ( .A1(n13759), .A2(n13758), .ZN(n13804) );
  AND2_X1 U13782 ( .A1(n13756), .A2(n13805), .ZN(n13803) );
  OR2_X1 U13783 ( .A1(n13758), .A2(n13759), .ZN(n13805) );
  OR2_X1 U13784 ( .A1(n7715), .A2(n8578), .ZN(n13759) );
  OR2_X1 U13785 ( .A1(n13806), .A2(n13807), .ZN(n13758) );
  AND2_X1 U13786 ( .A1(n13755), .A2(n13754), .ZN(n13807) );
  AND2_X1 U13787 ( .A1(n13752), .A2(n13808), .ZN(n13806) );
  OR2_X1 U13788 ( .A1(n13754), .A2(n13755), .ZN(n13808) );
  OR2_X1 U13789 ( .A1(n7715), .A2(n8573), .ZN(n13755) );
  OR2_X1 U13790 ( .A1(n13809), .A2(n13810), .ZN(n13754) );
  AND2_X1 U13791 ( .A1(n13751), .A2(n13750), .ZN(n13810) );
  AND2_X1 U13792 ( .A1(n13748), .A2(n13811), .ZN(n13809) );
  OR2_X1 U13793 ( .A1(n13750), .A2(n13751), .ZN(n13811) );
  OR2_X1 U13794 ( .A1(n7715), .A2(n8568), .ZN(n13751) );
  OR2_X1 U13795 ( .A1(n13812), .A2(n13813), .ZN(n13750) );
  AND2_X1 U13796 ( .A1(n13747), .A2(n13746), .ZN(n13813) );
  AND2_X1 U13797 ( .A1(n13744), .A2(n13814), .ZN(n13812) );
  OR2_X1 U13798 ( .A1(n13746), .A2(n13747), .ZN(n13814) );
  OR2_X1 U13799 ( .A1(n7715), .A2(n8563), .ZN(n13747) );
  OR2_X1 U13800 ( .A1(n13815), .A2(n13816), .ZN(n13746) );
  AND2_X1 U13801 ( .A1(n13743), .A2(n13742), .ZN(n13816) );
  AND2_X1 U13802 ( .A1(n13740), .A2(n13817), .ZN(n13815) );
  OR2_X1 U13803 ( .A1(n13742), .A2(n13743), .ZN(n13817) );
  OR2_X1 U13804 ( .A1(n7715), .A2(n8558), .ZN(n13743) );
  OR2_X1 U13805 ( .A1(n13818), .A2(n13819), .ZN(n13742) );
  AND2_X1 U13806 ( .A1(n13739), .A2(n13738), .ZN(n13819) );
  AND2_X1 U13807 ( .A1(n13736), .A2(n13820), .ZN(n13818) );
  OR2_X1 U13808 ( .A1(n13738), .A2(n13739), .ZN(n13820) );
  OR2_X1 U13809 ( .A1(n7715), .A2(n8553), .ZN(n13739) );
  OR2_X1 U13810 ( .A1(n13821), .A2(n13822), .ZN(n13738) );
  AND2_X1 U13811 ( .A1(n13735), .A2(n13734), .ZN(n13822) );
  AND2_X1 U13812 ( .A1(n13732), .A2(n13823), .ZN(n13821) );
  OR2_X1 U13813 ( .A1(n13734), .A2(n13735), .ZN(n13823) );
  OR2_X1 U13814 ( .A1(n7715), .A2(n8548), .ZN(n13735) );
  OR2_X1 U13815 ( .A1(n13824), .A2(n13825), .ZN(n13734) );
  AND2_X1 U13816 ( .A1(n13728), .A2(n13731), .ZN(n13825) );
  AND2_X1 U13817 ( .A1(n13826), .A2(n13730), .ZN(n13824) );
  OR2_X1 U13818 ( .A1(n13827), .A2(n13828), .ZN(n13730) );
  AND2_X1 U13819 ( .A1(n13727), .A2(n13726), .ZN(n13828) );
  AND2_X1 U13820 ( .A1(n13724), .A2(n13829), .ZN(n13827) );
  OR2_X1 U13821 ( .A1(n13726), .A2(n13727), .ZN(n13829) );
  OR2_X1 U13822 ( .A1(n8538), .A2(n7715), .ZN(n13727) );
  OR2_X1 U13823 ( .A1(n13830), .A2(n13831), .ZN(n13726) );
  AND2_X1 U13824 ( .A1(n13720), .A2(n13723), .ZN(n13831) );
  AND2_X1 U13825 ( .A1(n13832), .A2(n13722), .ZN(n13830) );
  OR2_X1 U13826 ( .A1(n13833), .A2(n13834), .ZN(n13722) );
  AND2_X1 U13827 ( .A1(n13716), .A2(n13719), .ZN(n13834) );
  AND2_X1 U13828 ( .A1(n13835), .A2(n13718), .ZN(n13833) );
  OR2_X1 U13829 ( .A1(n13836), .A2(n13837), .ZN(n13718) );
  AND2_X1 U13830 ( .A1(n13712), .A2(n13715), .ZN(n13837) );
  AND2_X1 U13831 ( .A1(n13838), .A2(n13714), .ZN(n13836) );
  OR2_X1 U13832 ( .A1(n13839), .A2(n13840), .ZN(n13714) );
  AND2_X1 U13833 ( .A1(n13709), .A2(n13710), .ZN(n13840) );
  AND2_X1 U13834 ( .A1(n13841), .A2(n13842), .ZN(n13839) );
  OR2_X1 U13835 ( .A1(n13710), .A2(n13709), .ZN(n13842) );
  OR2_X1 U13836 ( .A1(n8515), .A2(n7715), .ZN(n13709) );
  OR2_X1 U13837 ( .A1(n7689), .A2(n13843), .ZN(n13710) );
  OR2_X1 U13838 ( .A1(n8956), .A2(n7715), .ZN(n13843) );
  INV_X1 U13839 ( .A(n13711), .ZN(n13841) );
  OR2_X1 U13840 ( .A1(n13844), .A2(n13845), .ZN(n13711) );
  AND2_X1 U13841 ( .A1(b_4_), .A2(n13846), .ZN(n13845) );
  OR2_X1 U13842 ( .A1(n13847), .A2(n7343), .ZN(n13846) );
  AND2_X1 U13843 ( .A1(a_30_), .A2(n7659), .ZN(n13847) );
  AND2_X1 U13844 ( .A1(b_3_), .A2(n13848), .ZN(n13844) );
  OR2_X1 U13845 ( .A1(n13849), .A2(n7347), .ZN(n13848) );
  AND2_X1 U13846 ( .A1(a_31_), .A2(n7689), .ZN(n13849) );
  OR2_X1 U13847 ( .A1(n13715), .A2(n13712), .ZN(n13838) );
  XOR2_X1 U13848 ( .A(n13850), .B(n13851), .Z(n13712) );
  XNOR2_X1 U13849 ( .A(n13852), .B(n13853), .ZN(n13850) );
  OR2_X1 U13850 ( .A1(n8523), .A2(n7715), .ZN(n13715) );
  OR2_X1 U13851 ( .A1(n13719), .A2(n13716), .ZN(n13835) );
  XOR2_X1 U13852 ( .A(n13854), .B(n13855), .Z(n13716) );
  XOR2_X1 U13853 ( .A(n13856), .B(n13857), .Z(n13855) );
  OR2_X1 U13854 ( .A1(n8528), .A2(n7715), .ZN(n13719) );
  OR2_X1 U13855 ( .A1(n13723), .A2(n13720), .ZN(n13832) );
  XOR2_X1 U13856 ( .A(n13858), .B(n13859), .Z(n13720) );
  XOR2_X1 U13857 ( .A(n13860), .B(n13861), .Z(n13859) );
  OR2_X1 U13858 ( .A1(n8533), .A2(n7715), .ZN(n13723) );
  XOR2_X1 U13859 ( .A(n13862), .B(n13863), .Z(n13724) );
  XOR2_X1 U13860 ( .A(n13864), .B(n13865), .Z(n13863) );
  OR2_X1 U13861 ( .A1(n13731), .A2(n13728), .ZN(n13826) );
  XOR2_X1 U13862 ( .A(n13866), .B(n13867), .Z(n13728) );
  XOR2_X1 U13863 ( .A(n13868), .B(n13869), .Z(n13867) );
  OR2_X1 U13864 ( .A1(n7715), .A2(n8543), .ZN(n13731) );
  XOR2_X1 U13865 ( .A(n13870), .B(n13871), .Z(n13732) );
  XOR2_X1 U13866 ( .A(n13872), .B(n13873), .Z(n13871) );
  XOR2_X1 U13867 ( .A(n13874), .B(n13875), .Z(n13736) );
  XOR2_X1 U13868 ( .A(n13876), .B(n13877), .Z(n13875) );
  XOR2_X1 U13869 ( .A(n13878), .B(n13879), .Z(n13740) );
  XOR2_X1 U13870 ( .A(n13880), .B(n13881), .Z(n13879) );
  XOR2_X1 U13871 ( .A(n13882), .B(n13883), .Z(n13744) );
  XOR2_X1 U13872 ( .A(n13884), .B(n13885), .Z(n13883) );
  XOR2_X1 U13873 ( .A(n13886), .B(n13887), .Z(n13748) );
  XOR2_X1 U13874 ( .A(n13888), .B(n13889), .Z(n13887) );
  XOR2_X1 U13875 ( .A(n13890), .B(n13891), .Z(n13752) );
  XOR2_X1 U13876 ( .A(n13892), .B(n13893), .Z(n13891) );
  XOR2_X1 U13877 ( .A(n13894), .B(n13895), .Z(n13756) );
  XOR2_X1 U13878 ( .A(n13896), .B(n13897), .Z(n13895) );
  XOR2_X1 U13879 ( .A(n13898), .B(n13899), .Z(n13760) );
  XOR2_X1 U13880 ( .A(n13900), .B(n13901), .Z(n13899) );
  XOR2_X1 U13881 ( .A(n13902), .B(n13903), .Z(n13764) );
  XOR2_X1 U13882 ( .A(n13904), .B(n13905), .Z(n13903) );
  XOR2_X1 U13883 ( .A(n13906), .B(n13907), .Z(n13768) );
  XOR2_X1 U13884 ( .A(n13908), .B(n13909), .Z(n13907) );
  XOR2_X1 U13885 ( .A(n13910), .B(n13911), .Z(n13772) );
  XOR2_X1 U13886 ( .A(n13912), .B(n13913), .Z(n13911) );
  XOR2_X1 U13887 ( .A(n13914), .B(n13915), .Z(n13776) );
  XOR2_X1 U13888 ( .A(n13916), .B(n13917), .Z(n13915) );
  XOR2_X1 U13889 ( .A(n13918), .B(n13919), .Z(n13780) );
  XOR2_X1 U13890 ( .A(n13920), .B(n13921), .Z(n13919) );
  XOR2_X1 U13891 ( .A(n11787), .B(n13922), .Z(n11780) );
  XOR2_X1 U13892 ( .A(n11786), .B(n11785), .Z(n13922) );
  OR2_X1 U13893 ( .A1(n8608), .A2(n7689), .ZN(n11785) );
  OR2_X1 U13894 ( .A1(n13923), .A2(n13924), .ZN(n11786) );
  AND2_X1 U13895 ( .A1(n13921), .A2(n13920), .ZN(n13924) );
  AND2_X1 U13896 ( .A1(n13918), .A2(n13925), .ZN(n13923) );
  OR2_X1 U13897 ( .A1(n13920), .A2(n13921), .ZN(n13925) );
  OR2_X1 U13898 ( .A1(n7689), .A2(n8603), .ZN(n13921) );
  OR2_X1 U13899 ( .A1(n13926), .A2(n13927), .ZN(n13920) );
  AND2_X1 U13900 ( .A1(n13917), .A2(n13916), .ZN(n13927) );
  AND2_X1 U13901 ( .A1(n13914), .A2(n13928), .ZN(n13926) );
  OR2_X1 U13902 ( .A1(n13916), .A2(n13917), .ZN(n13928) );
  OR2_X1 U13903 ( .A1(n7689), .A2(n8598), .ZN(n13917) );
  OR2_X1 U13904 ( .A1(n13929), .A2(n13930), .ZN(n13916) );
  AND2_X1 U13905 ( .A1(n13913), .A2(n13912), .ZN(n13930) );
  AND2_X1 U13906 ( .A1(n13910), .A2(n13931), .ZN(n13929) );
  OR2_X1 U13907 ( .A1(n13912), .A2(n13913), .ZN(n13931) );
  OR2_X1 U13908 ( .A1(n7689), .A2(n8593), .ZN(n13913) );
  OR2_X1 U13909 ( .A1(n13932), .A2(n13933), .ZN(n13912) );
  AND2_X1 U13910 ( .A1(n13909), .A2(n13908), .ZN(n13933) );
  AND2_X1 U13911 ( .A1(n13906), .A2(n13934), .ZN(n13932) );
  OR2_X1 U13912 ( .A1(n13908), .A2(n13909), .ZN(n13934) );
  OR2_X1 U13913 ( .A1(n7689), .A2(n8588), .ZN(n13909) );
  OR2_X1 U13914 ( .A1(n13935), .A2(n13936), .ZN(n13908) );
  AND2_X1 U13915 ( .A1(n13905), .A2(n13904), .ZN(n13936) );
  AND2_X1 U13916 ( .A1(n13902), .A2(n13937), .ZN(n13935) );
  OR2_X1 U13917 ( .A1(n13904), .A2(n13905), .ZN(n13937) );
  OR2_X1 U13918 ( .A1(n7689), .A2(n8583), .ZN(n13905) );
  OR2_X1 U13919 ( .A1(n13938), .A2(n13939), .ZN(n13904) );
  AND2_X1 U13920 ( .A1(n13901), .A2(n13900), .ZN(n13939) );
  AND2_X1 U13921 ( .A1(n13898), .A2(n13940), .ZN(n13938) );
  OR2_X1 U13922 ( .A1(n13900), .A2(n13901), .ZN(n13940) );
  OR2_X1 U13923 ( .A1(n7689), .A2(n8578), .ZN(n13901) );
  OR2_X1 U13924 ( .A1(n13941), .A2(n13942), .ZN(n13900) );
  AND2_X1 U13925 ( .A1(n13897), .A2(n13896), .ZN(n13942) );
  AND2_X1 U13926 ( .A1(n13894), .A2(n13943), .ZN(n13941) );
  OR2_X1 U13927 ( .A1(n13896), .A2(n13897), .ZN(n13943) );
  OR2_X1 U13928 ( .A1(n7689), .A2(n8573), .ZN(n13897) );
  OR2_X1 U13929 ( .A1(n13944), .A2(n13945), .ZN(n13896) );
  AND2_X1 U13930 ( .A1(n13893), .A2(n13892), .ZN(n13945) );
  AND2_X1 U13931 ( .A1(n13890), .A2(n13946), .ZN(n13944) );
  OR2_X1 U13932 ( .A1(n13892), .A2(n13893), .ZN(n13946) );
  OR2_X1 U13933 ( .A1(n7689), .A2(n8568), .ZN(n13893) );
  OR2_X1 U13934 ( .A1(n13947), .A2(n13948), .ZN(n13892) );
  AND2_X1 U13935 ( .A1(n13889), .A2(n13888), .ZN(n13948) );
  AND2_X1 U13936 ( .A1(n13886), .A2(n13949), .ZN(n13947) );
  OR2_X1 U13937 ( .A1(n13888), .A2(n13889), .ZN(n13949) );
  OR2_X1 U13938 ( .A1(n7689), .A2(n8563), .ZN(n13889) );
  OR2_X1 U13939 ( .A1(n13950), .A2(n13951), .ZN(n13888) );
  AND2_X1 U13940 ( .A1(n13885), .A2(n13884), .ZN(n13951) );
  AND2_X1 U13941 ( .A1(n13882), .A2(n13952), .ZN(n13950) );
  OR2_X1 U13942 ( .A1(n13884), .A2(n13885), .ZN(n13952) );
  OR2_X1 U13943 ( .A1(n7689), .A2(n8558), .ZN(n13885) );
  OR2_X1 U13944 ( .A1(n13953), .A2(n13954), .ZN(n13884) );
  AND2_X1 U13945 ( .A1(n13881), .A2(n13880), .ZN(n13954) );
  AND2_X1 U13946 ( .A1(n13878), .A2(n13955), .ZN(n13953) );
  OR2_X1 U13947 ( .A1(n13880), .A2(n13881), .ZN(n13955) );
  OR2_X1 U13948 ( .A1(n7689), .A2(n8553), .ZN(n13881) );
  OR2_X1 U13949 ( .A1(n13956), .A2(n13957), .ZN(n13880) );
  AND2_X1 U13950 ( .A1(n13877), .A2(n13876), .ZN(n13957) );
  AND2_X1 U13951 ( .A1(n13874), .A2(n13958), .ZN(n13956) );
  OR2_X1 U13952 ( .A1(n13876), .A2(n13877), .ZN(n13958) );
  OR2_X1 U13953 ( .A1(n7689), .A2(n8548), .ZN(n13877) );
  OR2_X1 U13954 ( .A1(n13959), .A2(n13960), .ZN(n13876) );
  AND2_X1 U13955 ( .A1(n13873), .A2(n13872), .ZN(n13960) );
  AND2_X1 U13956 ( .A1(n13870), .A2(n13961), .ZN(n13959) );
  OR2_X1 U13957 ( .A1(n13872), .A2(n13873), .ZN(n13961) );
  OR2_X1 U13958 ( .A1(n8543), .A2(n7689), .ZN(n13873) );
  OR2_X1 U13959 ( .A1(n13962), .A2(n13963), .ZN(n13872) );
  AND2_X1 U13960 ( .A1(n13866), .A2(n13869), .ZN(n13963) );
  AND2_X1 U13961 ( .A1(n13964), .A2(n13868), .ZN(n13962) );
  OR2_X1 U13962 ( .A1(n13965), .A2(n13966), .ZN(n13868) );
  AND2_X1 U13963 ( .A1(n13865), .A2(n13864), .ZN(n13966) );
  AND2_X1 U13964 ( .A1(n13862), .A2(n13967), .ZN(n13965) );
  OR2_X1 U13965 ( .A1(n13864), .A2(n13865), .ZN(n13967) );
  OR2_X1 U13966 ( .A1(n8533), .A2(n7689), .ZN(n13865) );
  OR2_X1 U13967 ( .A1(n13968), .A2(n13969), .ZN(n13864) );
  AND2_X1 U13968 ( .A1(n13858), .A2(n13861), .ZN(n13969) );
  AND2_X1 U13969 ( .A1(n13970), .A2(n13860), .ZN(n13968) );
  OR2_X1 U13970 ( .A1(n13971), .A2(n13972), .ZN(n13860) );
  AND2_X1 U13971 ( .A1(n13854), .A2(n13857), .ZN(n13972) );
  AND2_X1 U13972 ( .A1(n13973), .A2(n13856), .ZN(n13971) );
  OR2_X1 U13973 ( .A1(n13974), .A2(n13975), .ZN(n13856) );
  AND2_X1 U13974 ( .A1(n13851), .A2(n13852), .ZN(n13975) );
  AND2_X1 U13975 ( .A1(n13976), .A2(n13977), .ZN(n13974) );
  OR2_X1 U13976 ( .A1(n13852), .A2(n13851), .ZN(n13977) );
  OR2_X1 U13977 ( .A1(n8515), .A2(n7689), .ZN(n13851) );
  OR2_X1 U13978 ( .A1(n7659), .A2(n13978), .ZN(n13852) );
  OR2_X1 U13979 ( .A1(n8956), .A2(n7689), .ZN(n13978) );
  INV_X1 U13980 ( .A(n13853), .ZN(n13976) );
  OR2_X1 U13981 ( .A1(n13979), .A2(n13980), .ZN(n13853) );
  AND2_X1 U13982 ( .A1(b_3_), .A2(n13981), .ZN(n13980) );
  OR2_X1 U13983 ( .A1(n13982), .A2(n7343), .ZN(n13981) );
  AND2_X1 U13984 ( .A1(a_30_), .A2(n13983), .ZN(n13982) );
  AND2_X1 U13985 ( .A1(b_2_), .A2(n13984), .ZN(n13979) );
  OR2_X1 U13986 ( .A1(n13985), .A2(n7347), .ZN(n13984) );
  AND2_X1 U13987 ( .A1(a_31_), .A2(n7659), .ZN(n13985) );
  OR2_X1 U13988 ( .A1(n13857), .A2(n13854), .ZN(n13973) );
  XOR2_X1 U13989 ( .A(n13986), .B(n13987), .Z(n13854) );
  XNOR2_X1 U13990 ( .A(n13988), .B(n13989), .ZN(n13986) );
  OR2_X1 U13991 ( .A1(n8523), .A2(n7689), .ZN(n13857) );
  OR2_X1 U13992 ( .A1(n13861), .A2(n13858), .ZN(n13970) );
  XOR2_X1 U13993 ( .A(n13990), .B(n13991), .Z(n13858) );
  XOR2_X1 U13994 ( .A(n13992), .B(n13993), .Z(n13991) );
  OR2_X1 U13995 ( .A1(n8528), .A2(n7689), .ZN(n13861) );
  XOR2_X1 U13996 ( .A(n13994), .B(n13995), .Z(n13862) );
  XOR2_X1 U13997 ( .A(n13996), .B(n13997), .Z(n13995) );
  OR2_X1 U13998 ( .A1(n13869), .A2(n13866), .ZN(n13964) );
  XOR2_X1 U13999 ( .A(n13998), .B(n13999), .Z(n13866) );
  XOR2_X1 U14000 ( .A(n14000), .B(n14001), .Z(n13999) );
  OR2_X1 U14001 ( .A1(n8538), .A2(n7689), .ZN(n13869) );
  XOR2_X1 U14002 ( .A(n14002), .B(n14003), .Z(n13870) );
  XOR2_X1 U14003 ( .A(n14004), .B(n14005), .Z(n14003) );
  XOR2_X1 U14004 ( .A(n14006), .B(n14007), .Z(n13874) );
  XOR2_X1 U14005 ( .A(n14008), .B(n14009), .Z(n14007) );
  XOR2_X1 U14006 ( .A(n14010), .B(n14011), .Z(n13878) );
  XOR2_X1 U14007 ( .A(n14012), .B(n14013), .Z(n14011) );
  XOR2_X1 U14008 ( .A(n14014), .B(n14015), .Z(n13882) );
  XOR2_X1 U14009 ( .A(n14016), .B(n14017), .Z(n14015) );
  XOR2_X1 U14010 ( .A(n14018), .B(n14019), .Z(n13886) );
  XOR2_X1 U14011 ( .A(n14020), .B(n14021), .Z(n14019) );
  XOR2_X1 U14012 ( .A(n14022), .B(n14023), .Z(n13890) );
  XOR2_X1 U14013 ( .A(n14024), .B(n14025), .Z(n14023) );
  XOR2_X1 U14014 ( .A(n14026), .B(n14027), .Z(n13894) );
  XOR2_X1 U14015 ( .A(n14028), .B(n14029), .Z(n14027) );
  XOR2_X1 U14016 ( .A(n14030), .B(n14031), .Z(n13898) );
  XOR2_X1 U14017 ( .A(n14032), .B(n14033), .Z(n14031) );
  XOR2_X1 U14018 ( .A(n14034), .B(n14035), .Z(n13902) );
  XOR2_X1 U14019 ( .A(n14036), .B(n14037), .Z(n14035) );
  XOR2_X1 U14020 ( .A(n14038), .B(n14039), .Z(n13906) );
  XOR2_X1 U14021 ( .A(n14040), .B(n14041), .Z(n14039) );
  XOR2_X1 U14022 ( .A(n14042), .B(n14043), .Z(n13910) );
  XOR2_X1 U14023 ( .A(n14044), .B(n14045), .Z(n14043) );
  XOR2_X1 U14024 ( .A(n14046), .B(n14047), .Z(n13914) );
  XOR2_X1 U14025 ( .A(n14048), .B(n14049), .Z(n14047) );
  XOR2_X1 U14026 ( .A(n14050), .B(n14051), .Z(n13918) );
  XOR2_X1 U14027 ( .A(n14052), .B(n14053), .Z(n14051) );
  XOR2_X1 U14028 ( .A(n11794), .B(n14054), .Z(n11787) );
  XOR2_X1 U14029 ( .A(n11793), .B(n11792), .Z(n14054) );
  OR2_X1 U14030 ( .A1(n7659), .A2(n8603), .ZN(n11792) );
  OR2_X1 U14031 ( .A1(n14055), .A2(n14056), .ZN(n11793) );
  AND2_X1 U14032 ( .A1(n14053), .A2(n14052), .ZN(n14056) );
  AND2_X1 U14033 ( .A1(n14050), .A2(n14057), .ZN(n14055) );
  OR2_X1 U14034 ( .A1(n14052), .A2(n14053), .ZN(n14057) );
  OR2_X1 U14035 ( .A1(n7659), .A2(n8598), .ZN(n14053) );
  OR2_X1 U14036 ( .A1(n14058), .A2(n14059), .ZN(n14052) );
  AND2_X1 U14037 ( .A1(n14049), .A2(n14048), .ZN(n14059) );
  AND2_X1 U14038 ( .A1(n14046), .A2(n14060), .ZN(n14058) );
  OR2_X1 U14039 ( .A1(n14048), .A2(n14049), .ZN(n14060) );
  OR2_X1 U14040 ( .A1(n7659), .A2(n8593), .ZN(n14049) );
  OR2_X1 U14041 ( .A1(n14061), .A2(n14062), .ZN(n14048) );
  AND2_X1 U14042 ( .A1(n14045), .A2(n14044), .ZN(n14062) );
  AND2_X1 U14043 ( .A1(n14042), .A2(n14063), .ZN(n14061) );
  OR2_X1 U14044 ( .A1(n14044), .A2(n14045), .ZN(n14063) );
  OR2_X1 U14045 ( .A1(n7659), .A2(n8588), .ZN(n14045) );
  OR2_X1 U14046 ( .A1(n14064), .A2(n14065), .ZN(n14044) );
  AND2_X1 U14047 ( .A1(n14041), .A2(n14040), .ZN(n14065) );
  AND2_X1 U14048 ( .A1(n14038), .A2(n14066), .ZN(n14064) );
  OR2_X1 U14049 ( .A1(n14040), .A2(n14041), .ZN(n14066) );
  OR2_X1 U14050 ( .A1(n7659), .A2(n8583), .ZN(n14041) );
  OR2_X1 U14051 ( .A1(n14067), .A2(n14068), .ZN(n14040) );
  AND2_X1 U14052 ( .A1(n14037), .A2(n14036), .ZN(n14068) );
  AND2_X1 U14053 ( .A1(n14034), .A2(n14069), .ZN(n14067) );
  OR2_X1 U14054 ( .A1(n14036), .A2(n14037), .ZN(n14069) );
  OR2_X1 U14055 ( .A1(n7659), .A2(n8578), .ZN(n14037) );
  OR2_X1 U14056 ( .A1(n14070), .A2(n14071), .ZN(n14036) );
  AND2_X1 U14057 ( .A1(n14033), .A2(n14032), .ZN(n14071) );
  AND2_X1 U14058 ( .A1(n14030), .A2(n14072), .ZN(n14070) );
  OR2_X1 U14059 ( .A1(n14032), .A2(n14033), .ZN(n14072) );
  OR2_X1 U14060 ( .A1(n7659), .A2(n8573), .ZN(n14033) );
  OR2_X1 U14061 ( .A1(n14073), .A2(n14074), .ZN(n14032) );
  AND2_X1 U14062 ( .A1(n14029), .A2(n14028), .ZN(n14074) );
  AND2_X1 U14063 ( .A1(n14026), .A2(n14075), .ZN(n14073) );
  OR2_X1 U14064 ( .A1(n14028), .A2(n14029), .ZN(n14075) );
  OR2_X1 U14065 ( .A1(n7659), .A2(n8568), .ZN(n14029) );
  OR2_X1 U14066 ( .A1(n14076), .A2(n14077), .ZN(n14028) );
  AND2_X1 U14067 ( .A1(n14025), .A2(n14024), .ZN(n14077) );
  AND2_X1 U14068 ( .A1(n14022), .A2(n14078), .ZN(n14076) );
  OR2_X1 U14069 ( .A1(n14024), .A2(n14025), .ZN(n14078) );
  OR2_X1 U14070 ( .A1(n7659), .A2(n8563), .ZN(n14025) );
  OR2_X1 U14071 ( .A1(n14079), .A2(n14080), .ZN(n14024) );
  AND2_X1 U14072 ( .A1(n14021), .A2(n14020), .ZN(n14080) );
  AND2_X1 U14073 ( .A1(n14018), .A2(n14081), .ZN(n14079) );
  OR2_X1 U14074 ( .A1(n14020), .A2(n14021), .ZN(n14081) );
  OR2_X1 U14075 ( .A1(n7659), .A2(n8558), .ZN(n14021) );
  OR2_X1 U14076 ( .A1(n14082), .A2(n14083), .ZN(n14020) );
  AND2_X1 U14077 ( .A1(n14017), .A2(n14016), .ZN(n14083) );
  AND2_X1 U14078 ( .A1(n14014), .A2(n14084), .ZN(n14082) );
  OR2_X1 U14079 ( .A1(n14016), .A2(n14017), .ZN(n14084) );
  OR2_X1 U14080 ( .A1(n7659), .A2(n8553), .ZN(n14017) );
  OR2_X1 U14081 ( .A1(n14085), .A2(n14086), .ZN(n14016) );
  AND2_X1 U14082 ( .A1(n14013), .A2(n14012), .ZN(n14086) );
  AND2_X1 U14083 ( .A1(n14010), .A2(n14087), .ZN(n14085) );
  OR2_X1 U14084 ( .A1(n14012), .A2(n14013), .ZN(n14087) );
  OR2_X1 U14085 ( .A1(n8548), .A2(n7659), .ZN(n14013) );
  OR2_X1 U14086 ( .A1(n14088), .A2(n14089), .ZN(n14012) );
  AND2_X1 U14087 ( .A1(n14009), .A2(n14008), .ZN(n14089) );
  AND2_X1 U14088 ( .A1(n14006), .A2(n14090), .ZN(n14088) );
  OR2_X1 U14089 ( .A1(n14008), .A2(n14009), .ZN(n14090) );
  OR2_X1 U14090 ( .A1(n8543), .A2(n7659), .ZN(n14009) );
  OR2_X1 U14091 ( .A1(n14091), .A2(n14092), .ZN(n14008) );
  AND2_X1 U14092 ( .A1(n14005), .A2(n14004), .ZN(n14092) );
  AND2_X1 U14093 ( .A1(n14002), .A2(n14093), .ZN(n14091) );
  OR2_X1 U14094 ( .A1(n14004), .A2(n14005), .ZN(n14093) );
  OR2_X1 U14095 ( .A1(n8538), .A2(n7659), .ZN(n14005) );
  OR2_X1 U14096 ( .A1(n14094), .A2(n14095), .ZN(n14004) );
  AND2_X1 U14097 ( .A1(n13998), .A2(n14001), .ZN(n14095) );
  AND2_X1 U14098 ( .A1(n14096), .A2(n14000), .ZN(n14094) );
  OR2_X1 U14099 ( .A1(n14097), .A2(n14098), .ZN(n14000) );
  AND2_X1 U14100 ( .A1(n13997), .A2(n13996), .ZN(n14098) );
  AND2_X1 U14101 ( .A1(n13994), .A2(n14099), .ZN(n14097) );
  OR2_X1 U14102 ( .A1(n13996), .A2(n13997), .ZN(n14099) );
  OR2_X1 U14103 ( .A1(n8528), .A2(n7659), .ZN(n13997) );
  OR2_X1 U14104 ( .A1(n14100), .A2(n14101), .ZN(n13996) );
  AND2_X1 U14105 ( .A1(n13990), .A2(n13993), .ZN(n14101) );
  AND2_X1 U14106 ( .A1(n14102), .A2(n13992), .ZN(n14100) );
  OR2_X1 U14107 ( .A1(n14103), .A2(n14104), .ZN(n13992) );
  AND2_X1 U14108 ( .A1(n13987), .A2(n13988), .ZN(n14104) );
  AND2_X1 U14109 ( .A1(n14105), .A2(n14106), .ZN(n14103) );
  OR2_X1 U14110 ( .A1(n13988), .A2(n13987), .ZN(n14106) );
  OR2_X1 U14111 ( .A1(n8515), .A2(n7659), .ZN(n13987) );
  OR2_X1 U14112 ( .A1(n13983), .A2(n14107), .ZN(n13988) );
  OR2_X1 U14113 ( .A1(n8956), .A2(n7659), .ZN(n14107) );
  INV_X1 U14114 ( .A(n13989), .ZN(n14105) );
  OR2_X1 U14115 ( .A1(n14108), .A2(n14109), .ZN(n13989) );
  AND2_X1 U14116 ( .A1(b_2_), .A2(n14110), .ZN(n14109) );
  OR2_X1 U14117 ( .A1(n14111), .A2(n7343), .ZN(n14110) );
  AND2_X1 U14118 ( .A1(a_30_), .A2(n14112), .ZN(n14111) );
  AND2_X1 U14119 ( .A1(b_1_), .A2(n14113), .ZN(n14108) );
  OR2_X1 U14120 ( .A1(n14114), .A2(n7347), .ZN(n14113) );
  AND2_X1 U14121 ( .A1(a_31_), .A2(n13983), .ZN(n14114) );
  OR2_X1 U14122 ( .A1(n13993), .A2(n13990), .ZN(n14102) );
  XOR2_X1 U14123 ( .A(n14115), .B(n14116), .Z(n13990) );
  XNOR2_X1 U14124 ( .A(n14117), .B(n14118), .ZN(n14115) );
  OR2_X1 U14125 ( .A1(n8523), .A2(n7659), .ZN(n13993) );
  XOR2_X1 U14126 ( .A(n14119), .B(n14120), .Z(n13994) );
  XOR2_X1 U14127 ( .A(n14121), .B(n14122), .Z(n14120) );
  OR2_X1 U14128 ( .A1(n14001), .A2(n13998), .ZN(n14096) );
  XOR2_X1 U14129 ( .A(n14123), .B(n14124), .Z(n13998) );
  XOR2_X1 U14130 ( .A(n14125), .B(n14126), .Z(n14124) );
  OR2_X1 U14131 ( .A1(n8533), .A2(n7659), .ZN(n14001) );
  XOR2_X1 U14132 ( .A(n14127), .B(n14128), .Z(n14002) );
  XOR2_X1 U14133 ( .A(n14129), .B(n14130), .Z(n14128) );
  XOR2_X1 U14134 ( .A(n14131), .B(n14132), .Z(n14006) );
  XOR2_X1 U14135 ( .A(n14133), .B(n14134), .Z(n14132) );
  XOR2_X1 U14136 ( .A(n14135), .B(n14136), .Z(n14010) );
  XOR2_X1 U14137 ( .A(n14137), .B(n14138), .Z(n14136) );
  XOR2_X1 U14138 ( .A(n14139), .B(n14140), .Z(n14014) );
  XOR2_X1 U14139 ( .A(n14141), .B(n14142), .Z(n14140) );
  XOR2_X1 U14140 ( .A(n14143), .B(n14144), .Z(n14018) );
  XOR2_X1 U14141 ( .A(n14145), .B(n14146), .Z(n14144) );
  XOR2_X1 U14142 ( .A(n14147), .B(n14148), .Z(n14022) );
  XOR2_X1 U14143 ( .A(n14149), .B(n14150), .Z(n14148) );
  XOR2_X1 U14144 ( .A(n14151), .B(n14152), .Z(n14026) );
  XOR2_X1 U14145 ( .A(n14153), .B(n14154), .Z(n14152) );
  XOR2_X1 U14146 ( .A(n14155), .B(n14156), .Z(n14030) );
  XOR2_X1 U14147 ( .A(n14157), .B(n14158), .Z(n14156) );
  XOR2_X1 U14148 ( .A(n14159), .B(n14160), .Z(n14034) );
  XOR2_X1 U14149 ( .A(n14161), .B(n14162), .Z(n14160) );
  XOR2_X1 U14150 ( .A(n14163), .B(n14164), .Z(n14038) );
  XOR2_X1 U14151 ( .A(n14165), .B(n14166), .Z(n14164) );
  XOR2_X1 U14152 ( .A(n14167), .B(n14168), .Z(n14042) );
  XOR2_X1 U14153 ( .A(n14169), .B(n14170), .Z(n14168) );
  XOR2_X1 U14154 ( .A(n14171), .B(n14172), .Z(n14046) );
  XOR2_X1 U14155 ( .A(n14173), .B(n14174), .Z(n14172) );
  XOR2_X1 U14156 ( .A(n14175), .B(n14176), .Z(n14050) );
  XOR2_X1 U14157 ( .A(n14177), .B(n14178), .Z(n14176) );
  XOR2_X1 U14158 ( .A(n14179), .B(n14180), .Z(n11794) );
  XOR2_X1 U14159 ( .A(n14181), .B(n14182), .Z(n14180) );
  AND2_X1 U14160 ( .A1(n7548), .A2(n14183), .ZN(n7550) );
  AND2_X1 U14161 ( .A1(n7549), .A2(n7547), .ZN(n14183) );
  XOR2_X1 U14162 ( .A(n14184), .B(n14185), .Z(n7547) );
  OR2_X1 U14163 ( .A1(n14186), .A2(n7660), .ZN(n14184) );
  XNOR2_X1 U14164 ( .A(n14187), .B(n14188), .ZN(n7549) );
  XOR2_X1 U14165 ( .A(n14189), .B(n14190), .Z(n14188) );
  INV_X1 U14166 ( .A(n7630), .ZN(n7548) );
  OR2_X1 U14167 ( .A1(n14191), .A2(n14192), .ZN(n7630) );
  AND2_X1 U14168 ( .A1(n7651), .A2(n7650), .ZN(n14192) );
  AND2_X1 U14169 ( .A1(n7648), .A2(n14193), .ZN(n14191) );
  OR2_X1 U14170 ( .A1(n7650), .A2(n7651), .ZN(n14193) );
  OR2_X1 U14171 ( .A1(n13983), .A2(n7660), .ZN(n7651) );
  OR2_X1 U14172 ( .A1(n14194), .A2(n14195), .ZN(n7650) );
  AND2_X1 U14173 ( .A1(n7670), .A2(n7669), .ZN(n14195) );
  AND2_X1 U14174 ( .A1(n7667), .A2(n14196), .ZN(n14194) );
  OR2_X1 U14175 ( .A1(n7669), .A2(n7670), .ZN(n14196) );
  OR2_X1 U14176 ( .A1(n13983), .A2(n7697), .ZN(n7670) );
  OR2_X1 U14177 ( .A1(n14197), .A2(n14198), .ZN(n7669) );
  AND2_X1 U14178 ( .A1(n7705), .A2(n7707), .ZN(n14198) );
  AND2_X1 U14179 ( .A1(n14199), .A2(n7706), .ZN(n14197) );
  OR2_X1 U14180 ( .A1(n7705), .A2(n7707), .ZN(n14199) );
  OR2_X1 U14181 ( .A1(n14200), .A2(n14201), .ZN(n7707) );
  AND2_X1 U14182 ( .A1(n7740), .A2(n7739), .ZN(n14201) );
  AND2_X1 U14183 ( .A1(n7737), .A2(n14202), .ZN(n14200) );
  OR2_X1 U14184 ( .A1(n7739), .A2(n7740), .ZN(n14202) );
  OR2_X1 U14185 ( .A1(n13983), .A2(n7820), .ZN(n7740) );
  OR2_X1 U14186 ( .A1(n14203), .A2(n14204), .ZN(n7739) );
  AND2_X1 U14187 ( .A1(n7784), .A2(n7783), .ZN(n14204) );
  AND2_X1 U14188 ( .A1(n7781), .A2(n14205), .ZN(n14203) );
  OR2_X1 U14189 ( .A1(n7783), .A2(n7784), .ZN(n14205) );
  OR2_X1 U14190 ( .A1(n13983), .A2(n7828), .ZN(n7784) );
  OR2_X1 U14191 ( .A1(n14206), .A2(n14207), .ZN(n7783) );
  AND2_X1 U14192 ( .A1(n7838), .A2(n7837), .ZN(n14207) );
  AND2_X1 U14193 ( .A1(n7835), .A2(n14208), .ZN(n14206) );
  OR2_X1 U14194 ( .A1(n7837), .A2(n7838), .ZN(n14208) );
  OR2_X1 U14195 ( .A1(n13983), .A2(n7887), .ZN(n7838) );
  OR2_X1 U14196 ( .A1(n14209), .A2(n14210), .ZN(n7837) );
  AND2_X1 U14197 ( .A1(n7897), .A2(n7896), .ZN(n14210) );
  AND2_X1 U14198 ( .A1(n7894), .A2(n14211), .ZN(n14209) );
  OR2_X1 U14199 ( .A1(n7896), .A2(n7897), .ZN(n14211) );
  OR2_X1 U14200 ( .A1(n13983), .A2(n7955), .ZN(n7897) );
  OR2_X1 U14201 ( .A1(n14212), .A2(n14213), .ZN(n7896) );
  AND2_X1 U14202 ( .A1(n7965), .A2(n7964), .ZN(n14213) );
  AND2_X1 U14203 ( .A1(n7962), .A2(n14214), .ZN(n14212) );
  OR2_X1 U14204 ( .A1(n7964), .A2(n7965), .ZN(n14214) );
  OR2_X1 U14205 ( .A1(n13983), .A2(n8025), .ZN(n7965) );
  OR2_X1 U14206 ( .A1(n14215), .A2(n14216), .ZN(n7964) );
  AND2_X1 U14207 ( .A1(n8035), .A2(n8034), .ZN(n14216) );
  AND2_X1 U14208 ( .A1(n8032), .A2(n14217), .ZN(n14215) );
  OR2_X1 U14209 ( .A1(n8034), .A2(n8035), .ZN(n14217) );
  OR2_X1 U14210 ( .A1(n13983), .A2(n8107), .ZN(n8035) );
  OR2_X1 U14211 ( .A1(n14218), .A2(n14219), .ZN(n8034) );
  AND2_X1 U14212 ( .A1(n8117), .A2(n8116), .ZN(n14219) );
  AND2_X1 U14213 ( .A1(n8114), .A2(n14220), .ZN(n14218) );
  OR2_X1 U14214 ( .A1(n8116), .A2(n8117), .ZN(n14220) );
  OR2_X1 U14215 ( .A1(n13983), .A2(n8191), .ZN(n8117) );
  OR2_X1 U14216 ( .A1(n14221), .A2(n14222), .ZN(n8116) );
  AND2_X1 U14217 ( .A1(n8201), .A2(n8200), .ZN(n14222) );
  AND2_X1 U14218 ( .A1(n8198), .A2(n14223), .ZN(n14221) );
  OR2_X1 U14219 ( .A1(n8200), .A2(n8201), .ZN(n14223) );
  OR2_X1 U14220 ( .A1(n13983), .A2(n8287), .ZN(n8201) );
  OR2_X1 U14221 ( .A1(n14224), .A2(n14225), .ZN(n8200) );
  AND2_X1 U14222 ( .A1(n8297), .A2(n8296), .ZN(n14225) );
  AND2_X1 U14223 ( .A1(n8294), .A2(n14226), .ZN(n14224) );
  OR2_X1 U14224 ( .A1(n8296), .A2(n8297), .ZN(n14226) );
  OR2_X1 U14225 ( .A1(n8608), .A2(n13983), .ZN(n8297) );
  OR2_X1 U14226 ( .A1(n14227), .A2(n14228), .ZN(n8296) );
  AND2_X1 U14227 ( .A1(n11799), .A2(n11798), .ZN(n14228) );
  AND2_X1 U14228 ( .A1(n11796), .A2(n14229), .ZN(n14227) );
  OR2_X1 U14229 ( .A1(n11798), .A2(n11799), .ZN(n14229) );
  OR2_X1 U14230 ( .A1(n13983), .A2(n8603), .ZN(n11799) );
  OR2_X1 U14231 ( .A1(n14230), .A2(n14231), .ZN(n11798) );
  AND2_X1 U14232 ( .A1(n14182), .A2(n14181), .ZN(n14231) );
  AND2_X1 U14233 ( .A1(n14179), .A2(n14232), .ZN(n14230) );
  OR2_X1 U14234 ( .A1(n14181), .A2(n14182), .ZN(n14232) );
  OR2_X1 U14235 ( .A1(n13983), .A2(n8598), .ZN(n14182) );
  OR2_X1 U14236 ( .A1(n14233), .A2(n14234), .ZN(n14181) );
  AND2_X1 U14237 ( .A1(n14178), .A2(n14177), .ZN(n14234) );
  AND2_X1 U14238 ( .A1(n14175), .A2(n14235), .ZN(n14233) );
  OR2_X1 U14239 ( .A1(n14177), .A2(n14178), .ZN(n14235) );
  OR2_X1 U14240 ( .A1(n13983), .A2(n8593), .ZN(n14178) );
  OR2_X1 U14241 ( .A1(n14236), .A2(n14237), .ZN(n14177) );
  AND2_X1 U14242 ( .A1(n14174), .A2(n14173), .ZN(n14237) );
  AND2_X1 U14243 ( .A1(n14171), .A2(n14238), .ZN(n14236) );
  OR2_X1 U14244 ( .A1(n14173), .A2(n14174), .ZN(n14238) );
  OR2_X1 U14245 ( .A1(n13983), .A2(n8588), .ZN(n14174) );
  OR2_X1 U14246 ( .A1(n14239), .A2(n14240), .ZN(n14173) );
  AND2_X1 U14247 ( .A1(n14170), .A2(n14169), .ZN(n14240) );
  AND2_X1 U14248 ( .A1(n14167), .A2(n14241), .ZN(n14239) );
  OR2_X1 U14249 ( .A1(n14169), .A2(n14170), .ZN(n14241) );
  OR2_X1 U14250 ( .A1(n13983), .A2(n8583), .ZN(n14170) );
  OR2_X1 U14251 ( .A1(n14242), .A2(n14243), .ZN(n14169) );
  AND2_X1 U14252 ( .A1(n14166), .A2(n14165), .ZN(n14243) );
  AND2_X1 U14253 ( .A1(n14163), .A2(n14244), .ZN(n14242) );
  OR2_X1 U14254 ( .A1(n14165), .A2(n14166), .ZN(n14244) );
  OR2_X1 U14255 ( .A1(n13983), .A2(n8578), .ZN(n14166) );
  OR2_X1 U14256 ( .A1(n14245), .A2(n14246), .ZN(n14165) );
  AND2_X1 U14257 ( .A1(n14162), .A2(n14161), .ZN(n14246) );
  AND2_X1 U14258 ( .A1(n14159), .A2(n14247), .ZN(n14245) );
  OR2_X1 U14259 ( .A1(n14161), .A2(n14162), .ZN(n14247) );
  OR2_X1 U14260 ( .A1(n13983), .A2(n8573), .ZN(n14162) );
  OR2_X1 U14261 ( .A1(n14248), .A2(n14249), .ZN(n14161) );
  AND2_X1 U14262 ( .A1(n14158), .A2(n14157), .ZN(n14249) );
  AND2_X1 U14263 ( .A1(n14155), .A2(n14250), .ZN(n14248) );
  OR2_X1 U14264 ( .A1(n14157), .A2(n14158), .ZN(n14250) );
  OR2_X1 U14265 ( .A1(n13983), .A2(n8568), .ZN(n14158) );
  OR2_X1 U14266 ( .A1(n14251), .A2(n14252), .ZN(n14157) );
  AND2_X1 U14267 ( .A1(n14154), .A2(n14153), .ZN(n14252) );
  AND2_X1 U14268 ( .A1(n14151), .A2(n14253), .ZN(n14251) );
  OR2_X1 U14269 ( .A1(n14153), .A2(n14154), .ZN(n14253) );
  OR2_X1 U14270 ( .A1(n13983), .A2(n8563), .ZN(n14154) );
  OR2_X1 U14271 ( .A1(n14254), .A2(n14255), .ZN(n14153) );
  AND2_X1 U14272 ( .A1(n14150), .A2(n14149), .ZN(n14255) );
  AND2_X1 U14273 ( .A1(n14147), .A2(n14256), .ZN(n14254) );
  OR2_X1 U14274 ( .A1(n14149), .A2(n14150), .ZN(n14256) );
  OR2_X1 U14275 ( .A1(n13983), .A2(n8558), .ZN(n14150) );
  OR2_X1 U14276 ( .A1(n14257), .A2(n14258), .ZN(n14149) );
  AND2_X1 U14277 ( .A1(n14146), .A2(n14145), .ZN(n14258) );
  AND2_X1 U14278 ( .A1(n14143), .A2(n14259), .ZN(n14257) );
  OR2_X1 U14279 ( .A1(n14145), .A2(n14146), .ZN(n14259) );
  OR2_X1 U14280 ( .A1(n8553), .A2(n13983), .ZN(n14146) );
  OR2_X1 U14281 ( .A1(n14260), .A2(n14261), .ZN(n14145) );
  AND2_X1 U14282 ( .A1(n14142), .A2(n14141), .ZN(n14261) );
  AND2_X1 U14283 ( .A1(n14139), .A2(n14262), .ZN(n14260) );
  OR2_X1 U14284 ( .A1(n14141), .A2(n14142), .ZN(n14262) );
  OR2_X1 U14285 ( .A1(n8548), .A2(n13983), .ZN(n14142) );
  OR2_X1 U14286 ( .A1(n14263), .A2(n14264), .ZN(n14141) );
  AND2_X1 U14287 ( .A1(n14138), .A2(n14137), .ZN(n14264) );
  AND2_X1 U14288 ( .A1(n14135), .A2(n14265), .ZN(n14263) );
  OR2_X1 U14289 ( .A1(n14137), .A2(n14138), .ZN(n14265) );
  OR2_X1 U14290 ( .A1(n8543), .A2(n13983), .ZN(n14138) );
  OR2_X1 U14291 ( .A1(n14266), .A2(n14267), .ZN(n14137) );
  AND2_X1 U14292 ( .A1(n14134), .A2(n14133), .ZN(n14267) );
  AND2_X1 U14293 ( .A1(n14131), .A2(n14268), .ZN(n14266) );
  OR2_X1 U14294 ( .A1(n14133), .A2(n14134), .ZN(n14268) );
  OR2_X1 U14295 ( .A1(n8538), .A2(n13983), .ZN(n14134) );
  OR2_X1 U14296 ( .A1(n14269), .A2(n14270), .ZN(n14133) );
  AND2_X1 U14297 ( .A1(n14130), .A2(n14129), .ZN(n14270) );
  AND2_X1 U14298 ( .A1(n14127), .A2(n14271), .ZN(n14269) );
  OR2_X1 U14299 ( .A1(n14129), .A2(n14130), .ZN(n14271) );
  OR2_X1 U14300 ( .A1(n8533), .A2(n13983), .ZN(n14130) );
  OR2_X1 U14301 ( .A1(n14272), .A2(n14273), .ZN(n14129) );
  AND2_X1 U14302 ( .A1(n14123), .A2(n14126), .ZN(n14273) );
  AND2_X1 U14303 ( .A1(n14274), .A2(n14125), .ZN(n14272) );
  OR2_X1 U14304 ( .A1(n14275), .A2(n14276), .ZN(n14125) );
  AND2_X1 U14305 ( .A1(n14122), .A2(n14121), .ZN(n14276) );
  AND2_X1 U14306 ( .A1(n14119), .A2(n14277), .ZN(n14275) );
  OR2_X1 U14307 ( .A1(n14121), .A2(n14122), .ZN(n14277) );
  OR2_X1 U14308 ( .A1(n8523), .A2(n13983), .ZN(n14122) );
  OR2_X1 U14309 ( .A1(n14278), .A2(n14279), .ZN(n14121) );
  AND2_X1 U14310 ( .A1(n14116), .A2(n14117), .ZN(n14279) );
  AND2_X1 U14311 ( .A1(n14280), .A2(n14281), .ZN(n14278) );
  OR2_X1 U14312 ( .A1(n14117), .A2(n14116), .ZN(n14281) );
  OR2_X1 U14313 ( .A1(n8515), .A2(n13983), .ZN(n14116) );
  OR2_X1 U14314 ( .A1(n14112), .A2(n14282), .ZN(n14117) );
  OR2_X1 U14315 ( .A1(n8956), .A2(n13983), .ZN(n14282) );
  INV_X1 U14316 ( .A(n14118), .ZN(n14280) );
  OR2_X1 U14317 ( .A1(n14283), .A2(n14284), .ZN(n14118) );
  AND2_X1 U14318 ( .A1(b_1_), .A2(n14285), .ZN(n14284) );
  OR2_X1 U14319 ( .A1(n14286), .A2(n7343), .ZN(n14285) );
  AND2_X1 U14320 ( .A1(n14287), .A2(a_30_), .ZN(n7343) );
  AND2_X1 U14321 ( .A1(a_30_), .A2(n14186), .ZN(n14286) );
  AND2_X1 U14322 ( .A1(b_0_), .A2(n14288), .ZN(n14283) );
  OR2_X1 U14323 ( .A1(n14289), .A2(n7347), .ZN(n14288) );
  AND2_X1 U14324 ( .A1(n14290), .A2(a_31_), .ZN(n7347) );
  AND2_X1 U14325 ( .A1(a_31_), .A2(n14112), .ZN(n14289) );
  XOR2_X1 U14326 ( .A(n14291), .B(n14292), .Z(n14119) );
  XOR2_X1 U14327 ( .A(n14293), .B(n14294), .Z(n14291) );
  OR2_X1 U14328 ( .A1(n14126), .A2(n14123), .ZN(n14274) );
  XNOR2_X1 U14329 ( .A(n14295), .B(n14296), .ZN(n14123) );
  XNOR2_X1 U14330 ( .A(n14297), .B(n14298), .ZN(n14296) );
  OR2_X1 U14331 ( .A1(n8528), .A2(n13983), .ZN(n14126) );
  XNOR2_X1 U14332 ( .A(n14299), .B(n14300), .ZN(n14127) );
  XNOR2_X1 U14333 ( .A(n14301), .B(n14302), .ZN(n14299) );
  XNOR2_X1 U14334 ( .A(n14303), .B(n14304), .ZN(n14131) );
  XNOR2_X1 U14335 ( .A(n14305), .B(n14306), .ZN(n14303) );
  XNOR2_X1 U14336 ( .A(n14307), .B(n14308), .ZN(n14135) );
  XNOR2_X1 U14337 ( .A(n14309), .B(n14310), .ZN(n14307) );
  XNOR2_X1 U14338 ( .A(n14311), .B(n14312), .ZN(n14139) );
  XNOR2_X1 U14339 ( .A(n14313), .B(n14314), .ZN(n14311) );
  XNOR2_X1 U14340 ( .A(n14315), .B(n14316), .ZN(n14143) );
  XNOR2_X1 U14341 ( .A(n14317), .B(n14318), .ZN(n14315) );
  XNOR2_X1 U14342 ( .A(n14319), .B(n14320), .ZN(n14147) );
  XNOR2_X1 U14343 ( .A(n14321), .B(n14322), .ZN(n14319) );
  XNOR2_X1 U14344 ( .A(n14323), .B(n14324), .ZN(n14151) );
  XNOR2_X1 U14345 ( .A(n14325), .B(n14326), .ZN(n14323) );
  XNOR2_X1 U14346 ( .A(n14327), .B(n14328), .ZN(n14155) );
  XNOR2_X1 U14347 ( .A(n14329), .B(n14330), .ZN(n14327) );
  XNOR2_X1 U14348 ( .A(n14331), .B(n14332), .ZN(n14159) );
  XNOR2_X1 U14349 ( .A(n14333), .B(n14334), .ZN(n14331) );
  XNOR2_X1 U14350 ( .A(n14335), .B(n14336), .ZN(n14163) );
  XNOR2_X1 U14351 ( .A(n14337), .B(n14338), .ZN(n14335) );
  XNOR2_X1 U14352 ( .A(n14339), .B(n14340), .ZN(n14167) );
  XNOR2_X1 U14353 ( .A(n14341), .B(n14342), .ZN(n14339) );
  XNOR2_X1 U14354 ( .A(n14343), .B(n14344), .ZN(n14171) );
  XNOR2_X1 U14355 ( .A(n14345), .B(n14346), .ZN(n14343) );
  XNOR2_X1 U14356 ( .A(n14347), .B(n14348), .ZN(n14175) );
  XNOR2_X1 U14357 ( .A(n14349), .B(n14350), .ZN(n14347) );
  XNOR2_X1 U14358 ( .A(n14351), .B(n14352), .ZN(n14179) );
  XNOR2_X1 U14359 ( .A(n14353), .B(n14354), .ZN(n14351) );
  XNOR2_X1 U14360 ( .A(n14355), .B(n14356), .ZN(n11796) );
  XNOR2_X1 U14361 ( .A(n14357), .B(n14358), .ZN(n14355) );
  XNOR2_X1 U14362 ( .A(n14359), .B(n14360), .ZN(n8294) );
  XNOR2_X1 U14363 ( .A(n14361), .B(n14362), .ZN(n14359) );
  XNOR2_X1 U14364 ( .A(n14363), .B(n14364), .ZN(n8198) );
  XNOR2_X1 U14365 ( .A(n14365), .B(n14366), .ZN(n14363) );
  XNOR2_X1 U14366 ( .A(n14367), .B(n14368), .ZN(n8114) );
  XNOR2_X1 U14367 ( .A(n14369), .B(n14370), .ZN(n14367) );
  XNOR2_X1 U14368 ( .A(n14371), .B(n14372), .ZN(n8032) );
  XNOR2_X1 U14369 ( .A(n14373), .B(n14374), .ZN(n14371) );
  XOR2_X1 U14370 ( .A(n14375), .B(n14376), .Z(n7962) );
  XOR2_X1 U14371 ( .A(n14377), .B(n14378), .Z(n14376) );
  XOR2_X1 U14372 ( .A(n14379), .B(n14380), .Z(n7894) );
  XOR2_X1 U14373 ( .A(n14381), .B(n14382), .Z(n14380) );
  XOR2_X1 U14374 ( .A(n14383), .B(n14384), .Z(n7835) );
  XOR2_X1 U14375 ( .A(n14385), .B(n14386), .Z(n14384) );
  XOR2_X1 U14376 ( .A(n14387), .B(n14388), .Z(n7781) );
  XOR2_X1 U14377 ( .A(n14389), .B(n14390), .Z(n14388) );
  XOR2_X1 U14378 ( .A(n14391), .B(n14392), .Z(n7737) );
  XOR2_X1 U14379 ( .A(n14393), .B(n14394), .Z(n14392) );
  XOR2_X1 U14380 ( .A(n14395), .B(n14396), .Z(n7705) );
  XOR2_X1 U14381 ( .A(n14397), .B(n14398), .Z(n14396) );
  XOR2_X1 U14382 ( .A(n14399), .B(n14400), .Z(n7667) );
  XOR2_X1 U14383 ( .A(n14401), .B(n14402), .Z(n14400) );
  XOR2_X1 U14384 ( .A(n14403), .B(n14404), .Z(n7648) );
  XOR2_X1 U14385 ( .A(n14405), .B(n14406), .Z(n14404) );
  AND2_X1 U14386 ( .A1(n14407), .A2(a_0_), .ZN(n7627) );
  INV_X1 U14387 ( .A(n14185), .ZN(n14407) );
  OR2_X1 U14388 ( .A1(n14408), .A2(n14409), .ZN(n14185) );
  AND2_X1 U14389 ( .A1(n14187), .A2(n14189), .ZN(n14409) );
  AND2_X1 U14390 ( .A1(n14410), .A2(n14190), .ZN(n14408) );
  OR2_X1 U14391 ( .A1(n14112), .A2(n7660), .ZN(n14190) );
  INV_X1 U14392 ( .A(a_0_), .ZN(n7660) );
  OR2_X1 U14393 ( .A1(n14189), .A2(n14187), .ZN(n14410) );
  OR2_X1 U14394 ( .A1(n14186), .A2(n7697), .ZN(n14187) );
  OR2_X1 U14395 ( .A1(n14411), .A2(n14412), .ZN(n14189) );
  AND2_X1 U14396 ( .A1(n14403), .A2(n14405), .ZN(n14412) );
  AND2_X1 U14397 ( .A1(n14413), .A2(n14406), .ZN(n14411) );
  OR2_X1 U14398 ( .A1(n14405), .A2(n14403), .ZN(n14413) );
  OR2_X1 U14399 ( .A1(n14186), .A2(n7730), .ZN(n14403) );
  OR2_X1 U14400 ( .A1(n14414), .A2(n14415), .ZN(n14405) );
  AND2_X1 U14401 ( .A1(n14399), .A2(n14401), .ZN(n14415) );
  AND2_X1 U14402 ( .A1(n14416), .A2(n14402), .ZN(n14414) );
  OR2_X1 U14403 ( .A1(n14186), .A2(n7820), .ZN(n14402) );
  OR2_X1 U14404 ( .A1(n14401), .A2(n14399), .ZN(n14416) );
  OR2_X1 U14405 ( .A1(n14112), .A2(n7730), .ZN(n14399) );
  OR2_X1 U14406 ( .A1(n14417), .A2(n14418), .ZN(n14401) );
  AND2_X1 U14407 ( .A1(n14395), .A2(n14397), .ZN(n14418) );
  AND2_X1 U14408 ( .A1(n14419), .A2(n14398), .ZN(n14417) );
  OR2_X1 U14409 ( .A1(n14186), .A2(n7828), .ZN(n14398) );
  OR2_X1 U14410 ( .A1(n14397), .A2(n14395), .ZN(n14419) );
  OR2_X1 U14411 ( .A1(n14112), .A2(n7820), .ZN(n14395) );
  OR2_X1 U14412 ( .A1(n14420), .A2(n14421), .ZN(n14397) );
  AND2_X1 U14413 ( .A1(n14391), .A2(n14393), .ZN(n14421) );
  AND2_X1 U14414 ( .A1(n14422), .A2(n14394), .ZN(n14420) );
  OR2_X1 U14415 ( .A1(n14186), .A2(n7887), .ZN(n14394) );
  OR2_X1 U14416 ( .A1(n14393), .A2(n14391), .ZN(n14422) );
  OR2_X1 U14417 ( .A1(n14112), .A2(n7828), .ZN(n14391) );
  OR2_X1 U14418 ( .A1(n14423), .A2(n14424), .ZN(n14393) );
  AND2_X1 U14419 ( .A1(n14387), .A2(n14389), .ZN(n14424) );
  AND2_X1 U14420 ( .A1(n14425), .A2(n14390), .ZN(n14423) );
  OR2_X1 U14421 ( .A1(n14186), .A2(n7955), .ZN(n14390) );
  OR2_X1 U14422 ( .A1(n14389), .A2(n14387), .ZN(n14425) );
  OR2_X1 U14423 ( .A1(n14112), .A2(n7887), .ZN(n14387) );
  OR2_X1 U14424 ( .A1(n14426), .A2(n14427), .ZN(n14389) );
  AND2_X1 U14425 ( .A1(n14383), .A2(n14385), .ZN(n14427) );
  AND2_X1 U14426 ( .A1(n14428), .A2(n14386), .ZN(n14426) );
  OR2_X1 U14427 ( .A1(n14186), .A2(n8025), .ZN(n14386) );
  OR2_X1 U14428 ( .A1(n14385), .A2(n14383), .ZN(n14428) );
  OR2_X1 U14429 ( .A1(n14112), .A2(n7955), .ZN(n14383) );
  OR2_X1 U14430 ( .A1(n14429), .A2(n14430), .ZN(n14385) );
  AND2_X1 U14431 ( .A1(n14379), .A2(n14381), .ZN(n14430) );
  AND2_X1 U14432 ( .A1(n14431), .A2(n14382), .ZN(n14429) );
  OR2_X1 U14433 ( .A1(n14186), .A2(n8107), .ZN(n14382) );
  OR2_X1 U14434 ( .A1(n14381), .A2(n14379), .ZN(n14431) );
  OR2_X1 U14435 ( .A1(n14112), .A2(n8025), .ZN(n14379) );
  OR2_X1 U14436 ( .A1(n14432), .A2(n14433), .ZN(n14381) );
  AND2_X1 U14437 ( .A1(n14375), .A2(n14377), .ZN(n14433) );
  AND2_X1 U14438 ( .A1(n14434), .A2(n14378), .ZN(n14432) );
  OR2_X1 U14439 ( .A1(n14186), .A2(n8191), .ZN(n14378) );
  OR2_X1 U14440 ( .A1(n14377), .A2(n14375), .ZN(n14434) );
  OR2_X1 U14441 ( .A1(n14112), .A2(n8107), .ZN(n14375) );
  OR2_X1 U14442 ( .A1(n14435), .A2(n14436), .ZN(n14377) );
  AND2_X1 U14443 ( .A1(n14372), .A2(n14374), .ZN(n14436) );
  AND2_X1 U14444 ( .A1(n14437), .A2(n14373), .ZN(n14435) );
  OR2_X1 U14445 ( .A1(n14186), .A2(n8287), .ZN(n14373) );
  OR2_X1 U14446 ( .A1(n14374), .A2(n14372), .ZN(n14437) );
  OR2_X1 U14447 ( .A1(n14112), .A2(n8191), .ZN(n14372) );
  OR2_X1 U14448 ( .A1(n14438), .A2(n14439), .ZN(n14374) );
  AND2_X1 U14449 ( .A1(n14368), .A2(n14370), .ZN(n14439) );
  AND2_X1 U14450 ( .A1(n14440), .A2(n14369), .ZN(n14438) );
  OR2_X1 U14451 ( .A1(n8608), .A2(n14186), .ZN(n14369) );
  OR2_X1 U14452 ( .A1(n14370), .A2(n14368), .ZN(n14440) );
  OR2_X1 U14453 ( .A1(n14112), .A2(n8287), .ZN(n14368) );
  OR2_X1 U14454 ( .A1(n14441), .A2(n14442), .ZN(n14370) );
  AND2_X1 U14455 ( .A1(n14364), .A2(n14366), .ZN(n14442) );
  AND2_X1 U14456 ( .A1(n14443), .A2(n14365), .ZN(n14441) );
  OR2_X1 U14457 ( .A1(n14186), .A2(n8603), .ZN(n14365) );
  OR2_X1 U14458 ( .A1(n14366), .A2(n14364), .ZN(n14443) );
  OR2_X1 U14459 ( .A1(n8608), .A2(n14112), .ZN(n14364) );
  OR2_X1 U14460 ( .A1(n14444), .A2(n14445), .ZN(n14366) );
  AND2_X1 U14461 ( .A1(n14360), .A2(n14362), .ZN(n14445) );
  AND2_X1 U14462 ( .A1(n14446), .A2(n14361), .ZN(n14444) );
  OR2_X1 U14463 ( .A1(n14186), .A2(n8598), .ZN(n14361) );
  OR2_X1 U14464 ( .A1(n14362), .A2(n14360), .ZN(n14446) );
  OR2_X1 U14465 ( .A1(n14112), .A2(n8603), .ZN(n14360) );
  OR2_X1 U14466 ( .A1(n14447), .A2(n14448), .ZN(n14362) );
  AND2_X1 U14467 ( .A1(n14356), .A2(n14358), .ZN(n14448) );
  AND2_X1 U14468 ( .A1(n14449), .A2(n14357), .ZN(n14447) );
  OR2_X1 U14469 ( .A1(n14186), .A2(n8593), .ZN(n14357) );
  OR2_X1 U14470 ( .A1(n14358), .A2(n14356), .ZN(n14449) );
  OR2_X1 U14471 ( .A1(n14112), .A2(n8598), .ZN(n14356) );
  OR2_X1 U14472 ( .A1(n14450), .A2(n14451), .ZN(n14358) );
  AND2_X1 U14473 ( .A1(n14352), .A2(n14354), .ZN(n14451) );
  AND2_X1 U14474 ( .A1(n14452), .A2(n14353), .ZN(n14450) );
  OR2_X1 U14475 ( .A1(n14186), .A2(n8588), .ZN(n14353) );
  OR2_X1 U14476 ( .A1(n14354), .A2(n14352), .ZN(n14452) );
  OR2_X1 U14477 ( .A1(n14112), .A2(n8593), .ZN(n14352) );
  OR2_X1 U14478 ( .A1(n14453), .A2(n14454), .ZN(n14354) );
  AND2_X1 U14479 ( .A1(n14348), .A2(n14350), .ZN(n14454) );
  AND2_X1 U14480 ( .A1(n14455), .A2(n14349), .ZN(n14453) );
  OR2_X1 U14481 ( .A1(n14186), .A2(n8583), .ZN(n14349) );
  OR2_X1 U14482 ( .A1(n14350), .A2(n14348), .ZN(n14455) );
  OR2_X1 U14483 ( .A1(n14112), .A2(n8588), .ZN(n14348) );
  OR2_X1 U14484 ( .A1(n14456), .A2(n14457), .ZN(n14350) );
  AND2_X1 U14485 ( .A1(n14344), .A2(n14346), .ZN(n14457) );
  AND2_X1 U14486 ( .A1(n14458), .A2(n14345), .ZN(n14456) );
  OR2_X1 U14487 ( .A1(n14186), .A2(n8578), .ZN(n14345) );
  OR2_X1 U14488 ( .A1(n14346), .A2(n14344), .ZN(n14458) );
  OR2_X1 U14489 ( .A1(n14112), .A2(n8583), .ZN(n14344) );
  OR2_X1 U14490 ( .A1(n14459), .A2(n14460), .ZN(n14346) );
  AND2_X1 U14491 ( .A1(n14340), .A2(n14342), .ZN(n14460) );
  AND2_X1 U14492 ( .A1(n14461), .A2(n14341), .ZN(n14459) );
  OR2_X1 U14493 ( .A1(n14186), .A2(n8573), .ZN(n14341) );
  OR2_X1 U14494 ( .A1(n14342), .A2(n14340), .ZN(n14461) );
  OR2_X1 U14495 ( .A1(n14112), .A2(n8578), .ZN(n14340) );
  OR2_X1 U14496 ( .A1(n14462), .A2(n14463), .ZN(n14342) );
  AND2_X1 U14497 ( .A1(n14336), .A2(n14338), .ZN(n14463) );
  AND2_X1 U14498 ( .A1(n14464), .A2(n14337), .ZN(n14462) );
  OR2_X1 U14499 ( .A1(n14186), .A2(n8568), .ZN(n14337) );
  OR2_X1 U14500 ( .A1(n14338), .A2(n14336), .ZN(n14464) );
  OR2_X1 U14501 ( .A1(n14112), .A2(n8573), .ZN(n14336) );
  OR2_X1 U14502 ( .A1(n14465), .A2(n14466), .ZN(n14338) );
  AND2_X1 U14503 ( .A1(n14332), .A2(n14334), .ZN(n14466) );
  AND2_X1 U14504 ( .A1(n14467), .A2(n14333), .ZN(n14465) );
  OR2_X1 U14505 ( .A1(n8563), .A2(n14186), .ZN(n14333) );
  OR2_X1 U14506 ( .A1(n14334), .A2(n14332), .ZN(n14467) );
  OR2_X1 U14507 ( .A1(n14112), .A2(n8568), .ZN(n14332) );
  OR2_X1 U14508 ( .A1(n14468), .A2(n14469), .ZN(n14334) );
  AND2_X1 U14509 ( .A1(n14328), .A2(n14330), .ZN(n14469) );
  AND2_X1 U14510 ( .A1(n14470), .A2(n14329), .ZN(n14468) );
  OR2_X1 U14511 ( .A1(n8558), .A2(n14186), .ZN(n14329) );
  OR2_X1 U14512 ( .A1(n14330), .A2(n14328), .ZN(n14470) );
  OR2_X1 U14513 ( .A1(n14112), .A2(n8563), .ZN(n14328) );
  OR2_X1 U14514 ( .A1(n14471), .A2(n14472), .ZN(n14330) );
  AND2_X1 U14515 ( .A1(n14324), .A2(n14326), .ZN(n14472) );
  AND2_X1 U14516 ( .A1(n14473), .A2(n14325), .ZN(n14471) );
  OR2_X1 U14517 ( .A1(n8553), .A2(n14186), .ZN(n14325) );
  OR2_X1 U14518 ( .A1(n14326), .A2(n14324), .ZN(n14473) );
  OR2_X1 U14519 ( .A1(n8558), .A2(n14112), .ZN(n14324) );
  OR2_X1 U14520 ( .A1(n14474), .A2(n14475), .ZN(n14326) );
  AND2_X1 U14521 ( .A1(n14320), .A2(n14322), .ZN(n14475) );
  AND2_X1 U14522 ( .A1(n14476), .A2(n14321), .ZN(n14474) );
  OR2_X1 U14523 ( .A1(n8548), .A2(n14186), .ZN(n14321) );
  OR2_X1 U14524 ( .A1(n14322), .A2(n14320), .ZN(n14476) );
  OR2_X1 U14525 ( .A1(n8553), .A2(n14112), .ZN(n14320) );
  OR2_X1 U14526 ( .A1(n14477), .A2(n14478), .ZN(n14322) );
  AND2_X1 U14527 ( .A1(n14316), .A2(n14318), .ZN(n14478) );
  AND2_X1 U14528 ( .A1(n14479), .A2(n14317), .ZN(n14477) );
  OR2_X1 U14529 ( .A1(n8543), .A2(n14186), .ZN(n14317) );
  OR2_X1 U14530 ( .A1(n14318), .A2(n14316), .ZN(n14479) );
  OR2_X1 U14531 ( .A1(n8548), .A2(n14112), .ZN(n14316) );
  OR2_X1 U14532 ( .A1(n14480), .A2(n14481), .ZN(n14318) );
  AND2_X1 U14533 ( .A1(n14312), .A2(n14314), .ZN(n14481) );
  AND2_X1 U14534 ( .A1(n14482), .A2(n14313), .ZN(n14480) );
  OR2_X1 U14535 ( .A1(n8538), .A2(n14186), .ZN(n14313) );
  OR2_X1 U14536 ( .A1(n14314), .A2(n14312), .ZN(n14482) );
  OR2_X1 U14537 ( .A1(n8543), .A2(n14112), .ZN(n14312) );
  OR2_X1 U14538 ( .A1(n14483), .A2(n14484), .ZN(n14314) );
  AND2_X1 U14539 ( .A1(n14308), .A2(n14310), .ZN(n14484) );
  AND2_X1 U14540 ( .A1(n14485), .A2(n14309), .ZN(n14483) );
  OR2_X1 U14541 ( .A1(n8533), .A2(n14186), .ZN(n14309) );
  OR2_X1 U14542 ( .A1(n14310), .A2(n14308), .ZN(n14485) );
  OR2_X1 U14543 ( .A1(n8538), .A2(n14112), .ZN(n14308) );
  OR2_X1 U14544 ( .A1(n14486), .A2(n14487), .ZN(n14310) );
  AND2_X1 U14545 ( .A1(n14304), .A2(n14306), .ZN(n14487) );
  AND2_X1 U14546 ( .A1(n14488), .A2(n14305), .ZN(n14486) );
  OR2_X1 U14547 ( .A1(n8528), .A2(n14186), .ZN(n14305) );
  OR2_X1 U14548 ( .A1(n14306), .A2(n14304), .ZN(n14488) );
  OR2_X1 U14549 ( .A1(n8533), .A2(n14112), .ZN(n14304) );
  OR2_X1 U14550 ( .A1(n14489), .A2(n14490), .ZN(n14306) );
  AND2_X1 U14551 ( .A1(n14300), .A2(n14302), .ZN(n14490) );
  AND2_X1 U14552 ( .A1(n14491), .A2(n14301), .ZN(n14489) );
  OR2_X1 U14553 ( .A1(n8523), .A2(n14186), .ZN(n14301) );
  OR2_X1 U14554 ( .A1(n14302), .A2(n14300), .ZN(n14491) );
  OR2_X1 U14555 ( .A1(n8528), .A2(n14112), .ZN(n14300) );
  OR2_X1 U14556 ( .A1(n14492), .A2(n14493), .ZN(n14302) );
  AND2_X1 U14557 ( .A1(n14295), .A2(n14298), .ZN(n14493) );
  AND2_X1 U14558 ( .A1(n14297), .A2(n14494), .ZN(n14492) );
  OR2_X1 U14559 ( .A1(n14298), .A2(n14295), .ZN(n14494) );
  OR2_X1 U14560 ( .A1(n8523), .A2(n14112), .ZN(n14295) );
  OR2_X1 U14561 ( .A1(n8515), .A2(n14186), .ZN(n14298) );
  AND2_X1 U14562 ( .A1(n14495), .A2(n14294), .ZN(n14297) );
  OR2_X1 U14563 ( .A1(n14186), .A2(n14496), .ZN(n14294) );
  OR2_X1 U14564 ( .A1(n8956), .A2(n14112), .ZN(n14496) );
  OR2_X1 U14565 ( .A1(n14290), .A2(n14287), .ZN(n8956) );
  INV_X1 U14566 ( .A(a_31_), .ZN(n14287) );
  INV_X1 U14567 ( .A(b_0_), .ZN(n14186) );
  INV_X1 U14568 ( .A(n14497), .ZN(n14495) );
  AND2_X1 U14569 ( .A1(n14292), .A2(n14293), .ZN(n14497) );
  AND2_X1 U14570 ( .A1(a_29_), .A2(b_1_), .ZN(n14293) );
  AND2_X1 U14571 ( .A1(b_0_), .A2(a_30_), .ZN(n14292) );
  OR2_X1 U14572 ( .A1(n14498), .A2(n14499), .ZN(Result_add_9_) );
  OR2_X1 U14573 ( .A1(n14500), .A2(n14501), .ZN(n14499) );
  AND2_X1 U14574 ( .A1(n14502), .A2(n7912), .ZN(n14501) );
  XNOR2_X1 U14575 ( .A(a_9_), .B(n14503), .ZN(n14502) );
  AND2_X1 U14576 ( .A1(n14504), .A2(b_9_), .ZN(n14500) );
  AND2_X1 U14577 ( .A1(n14503), .A2(n8191), .ZN(n14504) );
  INV_X1 U14578 ( .A(n14505), .ZN(n14498) );
  OR2_X1 U14579 ( .A1(n14503), .A2(n13152), .ZN(n14505) );
  XOR2_X1 U14580 ( .A(n14506), .B(n14507), .Z(Result_add_8_) );
  OR2_X1 U14581 ( .A1(n14508), .A2(n14509), .ZN(n14507) );
  OR2_X1 U14582 ( .A1(n14510), .A2(n14511), .ZN(Result_add_7_) );
  OR2_X1 U14583 ( .A1(n14512), .A2(n14513), .ZN(n14511) );
  AND2_X1 U14584 ( .A1(n14514), .A2(n7798), .ZN(n14513) );
  XNOR2_X1 U14585 ( .A(a_7_), .B(n14515), .ZN(n14514) );
  AND2_X1 U14586 ( .A1(n14516), .A2(b_7_), .ZN(n14512) );
  AND2_X1 U14587 ( .A1(n14515), .A2(n8025), .ZN(n14516) );
  INV_X1 U14588 ( .A(n14517), .ZN(n14510) );
  OR2_X1 U14589 ( .A1(n14515), .A2(n8264), .ZN(n14517) );
  XOR2_X1 U14590 ( .A(n14518), .B(n14519), .Z(Result_add_6_) );
  OR2_X1 U14591 ( .A1(n14520), .A2(n14521), .ZN(n14519) );
  OR2_X1 U14592 ( .A1(n14522), .A2(n14523), .ZN(Result_add_5_) );
  OR2_X1 U14593 ( .A1(n14524), .A2(n14525), .ZN(n14523) );
  AND2_X1 U14594 ( .A1(n14526), .A2(n7715), .ZN(n14525) );
  XNOR2_X1 U14595 ( .A(a_5_), .B(n14527), .ZN(n14526) );
  AND2_X1 U14596 ( .A1(n14528), .A2(b_5_), .ZN(n14524) );
  AND2_X1 U14597 ( .A1(n14527), .A2(n7887), .ZN(n14528) );
  INV_X1 U14598 ( .A(n14529), .ZN(n14522) );
  OR2_X1 U14599 ( .A1(n14527), .A2(n7946), .ZN(n14529) );
  XOR2_X1 U14600 ( .A(n14530), .B(n14531), .Z(Result_add_4_) );
  OR2_X1 U14601 ( .A1(n14532), .A2(n14533), .ZN(n14531) );
  OR2_X1 U14602 ( .A1(n14534), .A2(n14535), .ZN(Result_add_3_) );
  OR2_X1 U14603 ( .A1(n14536), .A2(n14537), .ZN(n14535) );
  AND2_X1 U14604 ( .A1(n14538), .A2(n7659), .ZN(n14537) );
  XNOR2_X1 U14605 ( .A(a_3_), .B(n14539), .ZN(n14538) );
  AND2_X1 U14606 ( .A1(n14540), .A2(b_3_), .ZN(n14536) );
  AND2_X1 U14607 ( .A1(n14539), .A2(n7820), .ZN(n14540) );
  INV_X1 U14608 ( .A(n14541), .ZN(n14534) );
  OR2_X1 U14609 ( .A1(n14539), .A2(n7736), .ZN(n14541) );
  XNOR2_X1 U14610 ( .A(n7348), .B(a_31_), .ZN(Result_add_31_) );
  INV_X1 U14611 ( .A(b_31_), .ZN(n7348) );
  OR2_X1 U14612 ( .A1(n14542), .A2(n14543), .ZN(Result_add_30_) );
  OR2_X1 U14613 ( .A1(n14544), .A2(n14545), .ZN(n14543) );
  AND2_X1 U14614 ( .A1(n14546), .A2(b_30_), .ZN(n14545) );
  AND2_X1 U14615 ( .A1(n14547), .A2(n7344), .ZN(n14544) );
  XNOR2_X1 U14616 ( .A(n14290), .B(Result_mul_63_), .ZN(n14547) );
  INV_X1 U14617 ( .A(n7350), .ZN(n14542) );
  OR2_X1 U14618 ( .A1(n7344), .A2(n14548), .ZN(n7350) );
  XOR2_X1 U14619 ( .A(n14549), .B(n14550), .Z(Result_add_2_) );
  OR2_X1 U14620 ( .A1(n14551), .A2(n14552), .ZN(n14550) );
  OR2_X1 U14621 ( .A1(n14553), .A2(n14554), .ZN(Result_add_29_) );
  OR2_X1 U14622 ( .A1(n14555), .A2(n14556), .ZN(n14554) );
  AND2_X1 U14623 ( .A1(n14557), .A2(n8520), .ZN(n14556) );
  XNOR2_X1 U14624 ( .A(n8515), .B(n14558), .ZN(n14557) );
  AND2_X1 U14625 ( .A1(n14559), .A2(b_29_), .ZN(n14555) );
  AND2_X1 U14626 ( .A1(n14560), .A2(n8515), .ZN(n14559) );
  AND2_X1 U14627 ( .A1(n14558), .A2(n14561), .ZN(n14553) );
  INV_X1 U14628 ( .A(n14560), .ZN(n14558) );
  XNOR2_X1 U14629 ( .A(n14562), .B(n14563), .ZN(Result_add_28_) );
  AND2_X1 U14630 ( .A1(n8971), .A2(n14564), .ZN(n14563) );
  OR2_X1 U14631 ( .A1(n14565), .A2(n14566), .ZN(Result_add_27_) );
  OR2_X1 U14632 ( .A1(n14567), .A2(n14568), .ZN(n14566) );
  AND2_X1 U14633 ( .A1(n14569), .A2(n8962), .ZN(n14568) );
  XNOR2_X1 U14634 ( .A(n8528), .B(n14570), .ZN(n14569) );
  AND2_X1 U14635 ( .A1(n14571), .A2(b_27_), .ZN(n14567) );
  AND2_X1 U14636 ( .A1(n14572), .A2(n8528), .ZN(n14571) );
  AND2_X1 U14637 ( .A1(n14570), .A2(n14573), .ZN(n14565) );
  XNOR2_X1 U14638 ( .A(n14574), .B(n14575), .ZN(Result_add_26_) );
  AND2_X1 U14639 ( .A1(n9435), .A2(n14576), .ZN(n14575) );
  OR2_X1 U14640 ( .A1(n14577), .A2(n14578), .ZN(Result_add_25_) );
  OR2_X1 U14641 ( .A1(n14579), .A2(n14580), .ZN(n14578) );
  AND2_X1 U14642 ( .A1(n14581), .A2(n9311), .ZN(n14580) );
  XNOR2_X1 U14643 ( .A(n8538), .B(n14582), .ZN(n14581) );
  AND2_X1 U14644 ( .A1(n14583), .A2(b_25_), .ZN(n14579) );
  AND2_X1 U14645 ( .A1(n14584), .A2(n8538), .ZN(n14583) );
  AND2_X1 U14646 ( .A1(n14582), .A2(n14585), .ZN(n14577) );
  XNOR2_X1 U14647 ( .A(n14586), .B(n14587), .ZN(Result_add_24_) );
  AND2_X1 U14648 ( .A1(n9861), .A2(n14588), .ZN(n14587) );
  OR2_X1 U14649 ( .A1(n14589), .A2(n14590), .ZN(Result_add_23_) );
  OR2_X1 U14650 ( .A1(n14591), .A2(n14592), .ZN(n14590) );
  AND2_X1 U14651 ( .A1(n14593), .A2(n9836), .ZN(n14592) );
  XNOR2_X1 U14652 ( .A(n8548), .B(n14594), .ZN(n14593) );
  AND2_X1 U14653 ( .A1(n14595), .A2(b_23_), .ZN(n14591) );
  AND2_X1 U14654 ( .A1(n14596), .A2(n8548), .ZN(n14595) );
  AND2_X1 U14655 ( .A1(n14594), .A2(n14597), .ZN(n14589) );
  XNOR2_X1 U14656 ( .A(n14598), .B(n14599), .ZN(Result_add_22_) );
  AND2_X1 U14657 ( .A1(n10306), .A2(n14600), .ZN(n14599) );
  OR2_X1 U14658 ( .A1(n14601), .A2(n14602), .ZN(Result_add_21_) );
  OR2_X1 U14659 ( .A1(n14603), .A2(n14604), .ZN(n14602) );
  AND2_X1 U14660 ( .A1(n14605), .A2(n10273), .ZN(n14604) );
  XNOR2_X1 U14661 ( .A(n8558), .B(n14606), .ZN(n14605) );
  AND2_X1 U14662 ( .A1(n14607), .A2(b_21_), .ZN(n14603) );
  AND2_X1 U14663 ( .A1(n14608), .A2(n8558), .ZN(n14607) );
  AND2_X1 U14664 ( .A1(n14606), .A2(n14609), .ZN(n14601) );
  XNOR2_X1 U14665 ( .A(n14610), .B(n14611), .ZN(Result_add_20_) );
  AND2_X1 U14666 ( .A1(n10768), .A2(n14612), .ZN(n14611) );
  OR2_X1 U14667 ( .A1(n14613), .A2(n14614), .ZN(Result_add_1_) );
  OR2_X1 U14668 ( .A1(n14615), .A2(n14616), .ZN(n14614) );
  AND2_X1 U14669 ( .A1(n14617), .A2(n14112), .ZN(n14616) );
  XNOR2_X1 U14670 ( .A(a_1_), .B(n14618), .ZN(n14617) );
  AND2_X1 U14671 ( .A1(n14619), .A2(b_1_), .ZN(n14615) );
  AND2_X1 U14672 ( .A1(n14618), .A2(n7697), .ZN(n14619) );
  INV_X1 U14673 ( .A(n14620), .ZN(n14613) );
  OR2_X1 U14674 ( .A1(n14618), .A2(n14406), .ZN(n14620) );
  OR2_X1 U14675 ( .A1(n14621), .A2(n14622), .ZN(Result_add_19_) );
  OR2_X1 U14676 ( .A1(n14623), .A2(n14624), .ZN(n14622) );
  AND2_X1 U14677 ( .A1(n14625), .A2(n10727), .ZN(n14624) );
  XNOR2_X1 U14678 ( .A(n8568), .B(n14626), .ZN(n14625) );
  AND2_X1 U14679 ( .A1(n14627), .A2(b_19_), .ZN(n14623) );
  AND2_X1 U14680 ( .A1(n14628), .A2(n8568), .ZN(n14627) );
  AND2_X1 U14681 ( .A1(n14626), .A2(n14629), .ZN(n14621) );
  XNOR2_X1 U14682 ( .A(n14630), .B(n14631), .ZN(Result_add_18_) );
  AND2_X1 U14683 ( .A1(n11193), .A2(n14632), .ZN(n14631) );
  OR2_X1 U14684 ( .A1(n14633), .A2(n14634), .ZN(Result_add_17_) );
  OR2_X1 U14685 ( .A1(n14635), .A2(n14636), .ZN(n14634) );
  AND2_X1 U14686 ( .A1(n14637), .A2(n11144), .ZN(n14636) );
  XNOR2_X1 U14687 ( .A(n8578), .B(n14638), .ZN(n14637) );
  AND2_X1 U14688 ( .A1(n14639), .A2(b_17_), .ZN(n14635) );
  AND2_X1 U14689 ( .A1(n14640), .A2(n8578), .ZN(n14639) );
  AND2_X1 U14690 ( .A1(n14638), .A2(n14641), .ZN(n14633) );
  XNOR2_X1 U14691 ( .A(n14642), .B(n14643), .ZN(Result_add_16_) );
  AND2_X1 U14692 ( .A1(n11649), .A2(n14644), .ZN(n14643) );
  OR2_X1 U14693 ( .A1(n14645), .A2(n14646), .ZN(Result_add_15_) );
  OR2_X1 U14694 ( .A1(n14647), .A2(n14648), .ZN(n14646) );
  AND2_X1 U14695 ( .A1(n14649), .A2(n11592), .ZN(n14648) );
  XNOR2_X1 U14696 ( .A(n8588), .B(n14650), .ZN(n14649) );
  AND2_X1 U14697 ( .A1(n14651), .A2(b_15_), .ZN(n14647) );
  AND2_X1 U14698 ( .A1(n14652), .A2(n8588), .ZN(n14651) );
  AND2_X1 U14699 ( .A1(n14650), .A2(n14653), .ZN(n14645) );
  XNOR2_X1 U14700 ( .A(n14654), .B(n14655), .ZN(Result_add_14_) );
  AND2_X1 U14701 ( .A1(n12178), .A2(n14656), .ZN(n14655) );
  INV_X1 U14702 ( .A(n14657), .ZN(n14656) );
  OR2_X1 U14703 ( .A1(n14658), .A2(n14659), .ZN(Result_add_13_) );
  OR2_X1 U14704 ( .A1(n14660), .A2(n14661), .ZN(n14659) );
  AND2_X1 U14705 ( .A1(n14662), .A2(n8216), .ZN(n14661) );
  XNOR2_X1 U14706 ( .A(a_13_), .B(n14663), .ZN(n14662) );
  AND2_X1 U14707 ( .A1(n14664), .A2(b_13_), .ZN(n14660) );
  AND2_X1 U14708 ( .A1(n14663), .A2(n8598), .ZN(n14664) );
  INV_X1 U14709 ( .A(n14665), .ZN(n14658) );
  OR2_X1 U14710 ( .A1(n14663), .A2(n12387), .ZN(n14665) );
  XOR2_X1 U14711 ( .A(n14666), .B(n14667), .Z(Result_add_12_) );
  OR2_X1 U14712 ( .A1(n14668), .A2(n14669), .ZN(n14667) );
  OR2_X1 U14713 ( .A1(n14670), .A2(n14671), .ZN(Result_add_11_) );
  OR2_X1 U14714 ( .A1(n14672), .A2(n14673), .ZN(n14671) );
  AND2_X1 U14715 ( .A1(n14674), .A2(n8050), .ZN(n14673) );
  XNOR2_X1 U14716 ( .A(a_11_), .B(n14675), .ZN(n14674) );
  AND2_X1 U14717 ( .A1(n14676), .A2(b_11_), .ZN(n14672) );
  AND2_X1 U14718 ( .A1(n14675), .A2(n8608), .ZN(n14676) );
  INV_X1 U14719 ( .A(n14677), .ZN(n14670) );
  OR2_X1 U14720 ( .A1(n14675), .A2(n12783), .ZN(n14677) );
  XOR2_X1 U14721 ( .A(n14678), .B(n14679), .Z(Result_add_10_) );
  OR2_X1 U14722 ( .A1(n14680), .A2(n14681), .ZN(n14679) );
  XOR2_X1 U14723 ( .A(n14682), .B(n14683), .Z(Result_add_0_) );
  XNOR2_X1 U14724 ( .A(a_0_), .B(b_0_), .ZN(n14683) );
  OR2_X1 U14725 ( .A1(n14684), .A2(n14685), .ZN(n14682) );
  AND2_X1 U14726 ( .A1(n7697), .A2(n14112), .ZN(n14685) );
  AND2_X1 U14727 ( .A1(n14618), .A2(n14406), .ZN(n14684) );
  OR2_X1 U14728 ( .A1(n14112), .A2(n7697), .ZN(n14406) );
  INV_X1 U14729 ( .A(a_1_), .ZN(n7697) );
  INV_X1 U14730 ( .A(b_1_), .ZN(n14112) );
  OR2_X1 U14731 ( .A1(n14686), .A2(n14551), .ZN(n14618) );
  AND2_X1 U14732 ( .A1(n7730), .A2(n13983), .ZN(n14551) );
  INV_X1 U14733 ( .A(b_2_), .ZN(n13983) );
  INV_X1 U14734 ( .A(a_2_), .ZN(n7730) );
  AND2_X1 U14735 ( .A1(n14549), .A2(n7706), .ZN(n14686) );
  INV_X1 U14736 ( .A(n14552), .ZN(n7706) );
  AND2_X1 U14737 ( .A1(b_2_), .A2(a_2_), .ZN(n14552) );
  OR2_X1 U14738 ( .A1(n14687), .A2(n14688), .ZN(n14549) );
  AND2_X1 U14739 ( .A1(n7820), .A2(n7659), .ZN(n14688) );
  AND2_X1 U14740 ( .A1(n14539), .A2(n7736), .ZN(n14687) );
  OR2_X1 U14741 ( .A1(n7659), .A2(n7820), .ZN(n7736) );
  INV_X1 U14742 ( .A(a_3_), .ZN(n7820) );
  OR2_X1 U14743 ( .A1(n14689), .A2(n14532), .ZN(n14539) );
  AND2_X1 U14744 ( .A1(n7828), .A2(n7689), .ZN(n14532) );
  INV_X1 U14745 ( .A(b_4_), .ZN(n7689) );
  INV_X1 U14746 ( .A(a_4_), .ZN(n7828) );
  AND2_X1 U14747 ( .A1(n14530), .A2(n7826), .ZN(n14689) );
  INV_X1 U14748 ( .A(n14533), .ZN(n7826) );
  AND2_X1 U14749 ( .A1(b_4_), .A2(a_4_), .ZN(n14533) );
  OR2_X1 U14750 ( .A1(n14690), .A2(n14691), .ZN(n14530) );
  AND2_X1 U14751 ( .A1(n7887), .A2(n7715), .ZN(n14691) );
  AND2_X1 U14752 ( .A1(n14527), .A2(n7946), .ZN(n14690) );
  OR2_X1 U14753 ( .A1(n7715), .A2(n7887), .ZN(n7946) );
  INV_X1 U14754 ( .A(a_5_), .ZN(n7887) );
  OR2_X1 U14755 ( .A1(n14692), .A2(n14520), .ZN(n14527) );
  AND2_X1 U14756 ( .A1(n7955), .A2(n7759), .ZN(n14520) );
  INV_X1 U14757 ( .A(b_6_), .ZN(n7759) );
  INV_X1 U14758 ( .A(a_6_), .ZN(n7955) );
  AND2_X1 U14759 ( .A1(n14518), .A2(n8091), .ZN(n14692) );
  INV_X1 U14760 ( .A(n14521), .ZN(n8091) );
  AND2_X1 U14761 ( .A1(b_6_), .A2(a_6_), .ZN(n14521) );
  OR2_X1 U14762 ( .A1(n14693), .A2(n14694), .ZN(n14518) );
  AND2_X1 U14763 ( .A1(n8025), .A2(n7798), .ZN(n14694) );
  AND2_X1 U14764 ( .A1(n14515), .A2(n8264), .ZN(n14693) );
  OR2_X1 U14765 ( .A1(n7798), .A2(n8025), .ZN(n8264) );
  INV_X1 U14766 ( .A(a_7_), .ZN(n8025) );
  OR2_X1 U14767 ( .A1(n14695), .A2(n14508), .ZN(n14515) );
  AND2_X1 U14768 ( .A1(n8107), .A2(n7857), .ZN(n14508) );
  INV_X1 U14769 ( .A(b_8_), .ZN(n7857) );
  INV_X1 U14770 ( .A(a_8_), .ZN(n8107) );
  AND2_X1 U14771 ( .A1(n14506), .A2(n13326), .ZN(n14695) );
  INV_X1 U14772 ( .A(n14509), .ZN(n13326) );
  AND2_X1 U14773 ( .A1(b_8_), .A2(a_8_), .ZN(n14509) );
  OR2_X1 U14774 ( .A1(n14696), .A2(n14697), .ZN(n14506) );
  AND2_X1 U14775 ( .A1(n8191), .A2(n7912), .ZN(n14697) );
  AND2_X1 U14776 ( .A1(n14503), .A2(n13152), .ZN(n14696) );
  OR2_X1 U14777 ( .A1(n7912), .A2(n8191), .ZN(n13152) );
  INV_X1 U14778 ( .A(a_9_), .ZN(n8191) );
  OR2_X1 U14779 ( .A1(n14698), .A2(n14680), .ZN(n14503) );
  AND2_X1 U14780 ( .A1(n8287), .A2(n7981), .ZN(n14680) );
  INV_X1 U14781 ( .A(b_10_), .ZN(n7981) );
  INV_X1 U14782 ( .A(a_10_), .ZN(n8287) );
  AND2_X1 U14783 ( .A1(n14678), .A2(n12971), .ZN(n14698) );
  INV_X1 U14784 ( .A(n14681), .ZN(n12971) );
  AND2_X1 U14785 ( .A1(b_10_), .A2(a_10_), .ZN(n14681) );
  OR2_X1 U14786 ( .A1(n14699), .A2(n14700), .ZN(n14678) );
  AND2_X1 U14787 ( .A1(n8608), .A2(n8050), .ZN(n14700) );
  AND2_X1 U14788 ( .A1(n14675), .A2(n12783), .ZN(n14699) );
  OR2_X1 U14789 ( .A1(n8608), .A2(n8050), .ZN(n12783) );
  INV_X1 U14790 ( .A(a_11_), .ZN(n8608) );
  OR2_X1 U14791 ( .A1(n14701), .A2(n14668), .ZN(n14675) );
  AND2_X1 U14792 ( .A1(n8603), .A2(n8133), .ZN(n14668) );
  INV_X1 U14793 ( .A(b_12_), .ZN(n8133) );
  INV_X1 U14794 ( .A(a_12_), .ZN(n8603) );
  AND2_X1 U14795 ( .A1(n14666), .A2(n12588), .ZN(n14701) );
  INV_X1 U14796 ( .A(n14669), .ZN(n12588) );
  AND2_X1 U14797 ( .A1(a_12_), .A2(b_12_), .ZN(n14669) );
  OR2_X1 U14798 ( .A1(n14702), .A2(n14703), .ZN(n14666) );
  AND2_X1 U14799 ( .A1(n8598), .A2(n8216), .ZN(n14703) );
  AND2_X1 U14800 ( .A1(n14663), .A2(n12387), .ZN(n14702) );
  OR2_X1 U14801 ( .A1(n8598), .A2(n8216), .ZN(n12387) );
  INV_X1 U14802 ( .A(b_13_), .ZN(n8216) );
  INV_X1 U14803 ( .A(a_13_), .ZN(n8598) );
  OR2_X1 U14804 ( .A1(n14704), .A2(n14657), .ZN(n14663) );
  AND2_X1 U14805 ( .A1(n8593), .A2(n11718), .ZN(n14657) );
  AND2_X1 U14806 ( .A1(n14654), .A2(n12178), .ZN(n14704) );
  OR2_X1 U14807 ( .A1(n8593), .A2(n11718), .ZN(n12178) );
  INV_X1 U14808 ( .A(b_14_), .ZN(n11718) );
  INV_X1 U14809 ( .A(a_14_), .ZN(n8593) );
  OR2_X1 U14810 ( .A1(n14705), .A2(n14706), .ZN(n14654) );
  AND2_X1 U14811 ( .A1(n8588), .A2(n11592), .ZN(n14706) );
  INV_X1 U14812 ( .A(b_15_), .ZN(n11592) );
  INV_X1 U14813 ( .A(a_15_), .ZN(n8588) );
  AND2_X1 U14814 ( .A1(n14652), .A2(n11963), .ZN(n14705) );
  INV_X1 U14815 ( .A(n14653), .ZN(n11963) );
  AND2_X1 U14816 ( .A1(a_15_), .A2(b_15_), .ZN(n14653) );
  INV_X1 U14817 ( .A(n14650), .ZN(n14652) );
  AND2_X1 U14818 ( .A1(n14707), .A2(n14644), .ZN(n14650) );
  OR2_X1 U14819 ( .A1(a_16_), .A2(b_16_), .ZN(n14644) );
  INV_X1 U14820 ( .A(n14708), .ZN(n14707) );
  AND2_X1 U14821 ( .A1(n14642), .A2(n11649), .ZN(n14708) );
  OR2_X1 U14822 ( .A1(n8583), .A2(n11391), .ZN(n11649) );
  INV_X1 U14823 ( .A(b_16_), .ZN(n11391) );
  INV_X1 U14824 ( .A(a_16_), .ZN(n8583) );
  OR2_X1 U14825 ( .A1(n14709), .A2(n14710), .ZN(n14642) );
  AND2_X1 U14826 ( .A1(n8578), .A2(n11144), .ZN(n14710) );
  INV_X1 U14827 ( .A(b_17_), .ZN(n11144) );
  INV_X1 U14828 ( .A(a_17_), .ZN(n8578) );
  AND2_X1 U14829 ( .A1(n14640), .A2(n11440), .ZN(n14709) );
  INV_X1 U14830 ( .A(n14641), .ZN(n11440) );
  AND2_X1 U14831 ( .A1(a_17_), .A2(b_17_), .ZN(n14641) );
  INV_X1 U14832 ( .A(n14638), .ZN(n14640) );
  AND2_X1 U14833 ( .A1(n14711), .A2(n14632), .ZN(n14638) );
  OR2_X1 U14834 ( .A1(a_18_), .A2(b_18_), .ZN(n14632) );
  INV_X1 U14835 ( .A(n14712), .ZN(n14711) );
  AND2_X1 U14836 ( .A1(n14630), .A2(n11193), .ZN(n14712) );
  OR2_X1 U14837 ( .A1(n8573), .A2(n10933), .ZN(n11193) );
  INV_X1 U14838 ( .A(b_18_), .ZN(n10933) );
  INV_X1 U14839 ( .A(a_18_), .ZN(n8573) );
  OR2_X1 U14840 ( .A1(n14713), .A2(n14714), .ZN(n14630) );
  AND2_X1 U14841 ( .A1(n8568), .A2(n10727), .ZN(n14714) );
  INV_X1 U14842 ( .A(b_19_), .ZN(n10727) );
  INV_X1 U14843 ( .A(a_19_), .ZN(n8568) );
  AND2_X1 U14844 ( .A1(n14628), .A2(n10978), .ZN(n14713) );
  INV_X1 U14845 ( .A(n14629), .ZN(n10978) );
  AND2_X1 U14846 ( .A1(a_19_), .A2(b_19_), .ZN(n14629) );
  INV_X1 U14847 ( .A(n14626), .ZN(n14628) );
  AND2_X1 U14848 ( .A1(n14715), .A2(n14612), .ZN(n14626) );
  OR2_X1 U14849 ( .A1(a_20_), .A2(b_20_), .ZN(n14612) );
  INV_X1 U14850 ( .A(n14716), .ZN(n14715) );
  AND2_X1 U14851 ( .A1(n14610), .A2(n10768), .ZN(n14716) );
  OR2_X1 U14852 ( .A1(n8563), .A2(n10407), .ZN(n10768) );
  INV_X1 U14853 ( .A(b_20_), .ZN(n10407) );
  INV_X1 U14854 ( .A(a_20_), .ZN(n8563) );
  OR2_X1 U14855 ( .A1(n14717), .A2(n14718), .ZN(n14610) );
  AND2_X1 U14856 ( .A1(n8558), .A2(n10273), .ZN(n14718) );
  INV_X1 U14857 ( .A(b_21_), .ZN(n10273) );
  INV_X1 U14858 ( .A(a_21_), .ZN(n8558) );
  AND2_X1 U14859 ( .A1(n14608), .A2(n10551), .ZN(n14717) );
  INV_X1 U14860 ( .A(n14609), .ZN(n10551) );
  AND2_X1 U14861 ( .A1(a_21_), .A2(b_21_), .ZN(n14609) );
  INV_X1 U14862 ( .A(n14606), .ZN(n14608) );
  AND2_X1 U14863 ( .A1(n14719), .A2(n14600), .ZN(n14606) );
  OR2_X1 U14864 ( .A1(a_22_), .A2(b_22_), .ZN(n14600) );
  INV_X1 U14865 ( .A(n14720), .ZN(n14719) );
  AND2_X1 U14866 ( .A1(n14598), .A2(n10306), .ZN(n14720) );
  OR2_X1 U14867 ( .A1(n8553), .A2(n10057), .ZN(n10306) );
  INV_X1 U14868 ( .A(b_22_), .ZN(n10057) );
  INV_X1 U14869 ( .A(a_22_), .ZN(n8553) );
  OR2_X1 U14870 ( .A1(n14721), .A2(n14722), .ZN(n14598) );
  AND2_X1 U14871 ( .A1(n8548), .A2(n9836), .ZN(n14722) );
  INV_X1 U14872 ( .A(b_23_), .ZN(n9836) );
  INV_X1 U14873 ( .A(a_23_), .ZN(n8548) );
  AND2_X1 U14874 ( .A1(n14596), .A2(n10082), .ZN(n14721) );
  INV_X1 U14875 ( .A(n14597), .ZN(n10082) );
  AND2_X1 U14876 ( .A1(a_23_), .A2(b_23_), .ZN(n14597) );
  INV_X1 U14877 ( .A(n14594), .ZN(n14596) );
  AND2_X1 U14878 ( .A1(n14723), .A2(n14588), .ZN(n14594) );
  OR2_X1 U14879 ( .A1(a_24_), .A2(b_24_), .ZN(n14588) );
  INV_X1 U14880 ( .A(n14724), .ZN(n14723) );
  AND2_X1 U14881 ( .A1(n14586), .A2(n9861), .ZN(n14724) );
  OR2_X1 U14882 ( .A1(n8543), .A2(n9631), .ZN(n9861) );
  INV_X1 U14883 ( .A(b_24_), .ZN(n9631) );
  INV_X1 U14884 ( .A(a_24_), .ZN(n8543) );
  OR2_X1 U14885 ( .A1(n14725), .A2(n14726), .ZN(n14586) );
  AND2_X1 U14886 ( .A1(n8538), .A2(n9311), .ZN(n14726) );
  INV_X1 U14887 ( .A(b_25_), .ZN(n9311) );
  INV_X1 U14888 ( .A(a_25_), .ZN(n8538) );
  AND2_X1 U14889 ( .A1(n14584), .A2(n9652), .ZN(n14725) );
  INV_X1 U14890 ( .A(n14585), .ZN(n9652) );
  AND2_X1 U14891 ( .A1(a_25_), .A2(b_25_), .ZN(n14585) );
  INV_X1 U14892 ( .A(n14582), .ZN(n14584) );
  AND2_X1 U14893 ( .A1(n14727), .A2(n14576), .ZN(n14582) );
  OR2_X1 U14894 ( .A1(a_26_), .A2(b_26_), .ZN(n14576) );
  INV_X1 U14895 ( .A(n14728), .ZN(n14727) );
  AND2_X1 U14896 ( .A1(n14574), .A2(n9435), .ZN(n14728) );
  OR2_X1 U14897 ( .A1(n8533), .A2(n9185), .ZN(n9435) );
  INV_X1 U14898 ( .A(b_26_), .ZN(n9185) );
  INV_X1 U14899 ( .A(a_26_), .ZN(n8533) );
  OR2_X1 U14900 ( .A1(n14729), .A2(n14730), .ZN(n14574) );
  AND2_X1 U14901 ( .A1(n8528), .A2(n8962), .ZN(n14730) );
  INV_X1 U14902 ( .A(b_27_), .ZN(n8962) );
  INV_X1 U14903 ( .A(a_27_), .ZN(n8528) );
  AND2_X1 U14904 ( .A1(n14572), .A2(n9194), .ZN(n14729) );
  INV_X1 U14905 ( .A(n14573), .ZN(n9194) );
  AND2_X1 U14906 ( .A1(a_27_), .A2(b_27_), .ZN(n14573) );
  INV_X1 U14907 ( .A(n14570), .ZN(n14572) );
  AND2_X1 U14908 ( .A1(n14731), .A2(n14564), .ZN(n14570) );
  OR2_X1 U14909 ( .A1(a_28_), .A2(b_28_), .ZN(n14564) );
  INV_X1 U14910 ( .A(n14732), .ZN(n14731) );
  AND2_X1 U14911 ( .A1(n14562), .A2(n8971), .ZN(n14732) );
  OR2_X1 U14912 ( .A1(n8523), .A2(n8744), .ZN(n8971) );
  INV_X1 U14913 ( .A(b_28_), .ZN(n8744) );
  INV_X1 U14914 ( .A(a_28_), .ZN(n8523) );
  OR2_X1 U14915 ( .A1(n14733), .A2(n14734), .ZN(n14562) );
  AND2_X1 U14916 ( .A1(n8515), .A2(n8520), .ZN(n14734) );
  INV_X1 U14917 ( .A(b_29_), .ZN(n8520) );
  INV_X1 U14918 ( .A(a_29_), .ZN(n8515) );
  AND2_X1 U14919 ( .A1(n14560), .A2(n8749), .ZN(n14733) );
  INV_X1 U14920 ( .A(n14561), .ZN(n8749) );
  AND2_X1 U14921 ( .A1(a_29_), .A2(b_29_), .ZN(n14561) );
  OR2_X1 U14922 ( .A1(n14735), .A2(n14546), .ZN(n14560) );
  AND2_X1 U14923 ( .A1(n14736), .A2(n14290), .ZN(n14546) );
  AND2_X1 U14924 ( .A1(n14548), .A2(n7344), .ZN(n14735) );
  OR2_X1 U14925 ( .A1(n14290), .A2(n14736), .ZN(n14548) );
  INV_X1 U14926 ( .A(Result_mul_63_), .ZN(n14736) );
  AND2_X1 U14927 ( .A1(a_31_), .A2(b_31_), .ZN(Result_mul_63_) );
  INV_X1 U14928 ( .A(a_30_), .ZN(n14290) );
endmodule

