module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n1109_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n172_, keyIn_0_45 );
not g001 ( new_n173_, N102 );
and g002 ( new_n174_, new_n173_, keyIn_0_16 );
not g003 ( new_n175_, N108 );
not g004 ( new_n176_, keyIn_0_16 );
and g005 ( new_n177_, new_n176_, N102 );
or g006 ( new_n178_, new_n177_, new_n175_ );
or g007 ( new_n179_, new_n178_, new_n174_ );
not g008 ( new_n180_, new_n179_ );
and g009 ( new_n181_, new_n180_, keyIn_0_28 );
not g010 ( new_n182_, keyIn_0_28 );
and g011 ( new_n183_, new_n179_, new_n182_ );
or g012 ( new_n184_, new_n181_, new_n183_ );
or g013 ( new_n185_, keyIn_0_14, N89 );
not g014 ( new_n186_, N95 );
and g015 ( new_n187_, keyIn_0_14, N89 );
or g016 ( new_n188_, new_n187_, new_n186_ );
not g017 ( new_n189_, new_n188_ );
and g018 ( new_n190_, new_n189_, new_n185_ );
not g019 ( new_n191_, new_n190_ );
or g020 ( new_n192_, new_n191_, keyIn_0_27 );
not g021 ( new_n193_, keyIn_0_27 );
or g022 ( new_n194_, new_n190_, new_n193_ );
and g023 ( new_n195_, new_n192_, new_n194_ );
not g024 ( new_n196_, keyIn_0_26 );
not g025 ( new_n197_, N76 );
and g026 ( new_n198_, new_n197_, keyIn_0_12 );
not g027 ( new_n199_, new_n198_ );
or g028 ( new_n200_, new_n197_, keyIn_0_12 );
and g029 ( new_n201_, new_n200_, N82 );
and g030 ( new_n202_, new_n201_, new_n199_ );
not g031 ( new_n203_, new_n202_ );
or g032 ( new_n204_, new_n203_, new_n196_ );
or g033 ( new_n205_, new_n202_, keyIn_0_26 );
and g034 ( new_n206_, new_n204_, new_n205_ );
and g035 ( new_n207_, new_n195_, new_n206_ );
and g036 ( new_n208_, new_n207_, new_n184_ );
not g037 ( new_n209_, N1 );
and g038 ( new_n210_, new_n209_, keyIn_0_0 );
not g039 ( new_n211_, new_n210_ );
or g040 ( new_n212_, new_n209_, keyIn_0_0 );
and g041 ( new_n213_, new_n212_, N4 );
and g042 ( new_n214_, new_n213_, new_n211_ );
not g043 ( new_n215_, new_n214_ );
and g044 ( new_n216_, new_n215_, keyIn_0_18 );
not g045 ( new_n217_, keyIn_0_18 );
and g046 ( new_n218_, new_n214_, new_n217_ );
or g047 ( new_n219_, new_n216_, new_n218_ );
not g048 ( new_n220_, keyIn_0_21 );
not g049 ( new_n221_, N11 );
and g050 ( new_n222_, new_n221_, keyIn_0_2 );
not g051 ( new_n223_, new_n222_ );
or g052 ( new_n224_, new_n221_, keyIn_0_2 );
and g053 ( new_n225_, new_n224_, N17 );
and g054 ( new_n226_, new_n225_, new_n223_ );
not g055 ( new_n227_, new_n226_ );
and g056 ( new_n228_, new_n227_, new_n220_ );
and g057 ( new_n229_, new_n226_, keyIn_0_21 );
or g058 ( new_n230_, new_n228_, new_n229_ );
and g059 ( new_n231_, new_n219_, new_n230_ );
not g060 ( new_n232_, N50 );
and g061 ( new_n233_, new_n232_, keyIn_0_8 );
not g062 ( new_n234_, N56 );
not g063 ( new_n235_, keyIn_0_8 );
and g064 ( new_n236_, new_n235_, N50 );
or g065 ( new_n237_, new_n236_, new_n234_ );
or g066 ( new_n238_, new_n237_, new_n233_ );
and g067 ( new_n239_, new_n238_, keyIn_0_24 );
not g068 ( new_n240_, keyIn_0_24 );
not g069 ( new_n241_, new_n233_ );
or g070 ( new_n242_, new_n232_, keyIn_0_8 );
and g071 ( new_n243_, new_n242_, N56 );
and g072 ( new_n244_, new_n243_, new_n241_ );
and g073 ( new_n245_, new_n244_, new_n240_ );
or g074 ( new_n246_, new_n239_, new_n245_ );
not g075 ( new_n247_, keyIn_0_25 );
not g076 ( new_n248_, N63 );
and g077 ( new_n249_, new_n248_, keyIn_0_10 );
not g078 ( new_n250_, N69 );
not g079 ( new_n251_, keyIn_0_10 );
and g080 ( new_n252_, new_n251_, N63 );
or g081 ( new_n253_, new_n252_, new_n250_ );
or g082 ( new_n254_, new_n253_, new_n249_ );
or g083 ( new_n255_, new_n254_, new_n247_ );
not g084 ( new_n256_, new_n249_ );
or g085 ( new_n257_, new_n248_, keyIn_0_10 );
and g086 ( new_n258_, new_n257_, N69 );
and g087 ( new_n259_, new_n258_, new_n256_ );
or g088 ( new_n260_, new_n259_, keyIn_0_25 );
and g089 ( new_n261_, new_n255_, new_n260_ );
and g090 ( new_n262_, new_n246_, new_n261_ );
not g091 ( new_n263_, keyIn_0_23 );
and g092 ( new_n264_, keyIn_0_6, N37 );
not g093 ( new_n265_, keyIn_0_6 );
not g094 ( new_n266_, N37 );
and g095 ( new_n267_, new_n265_, new_n266_ );
or g096 ( new_n268_, new_n267_, new_n264_ );
and g097 ( new_n269_, new_n268_, N43 );
and g098 ( new_n270_, new_n269_, new_n263_ );
not g099 ( new_n271_, N43 );
not g100 ( new_n272_, new_n264_ );
or g101 ( new_n273_, keyIn_0_6, N37 );
and g102 ( new_n274_, new_n272_, new_n273_ );
or g103 ( new_n275_, new_n274_, new_n271_ );
and g104 ( new_n276_, new_n275_, keyIn_0_23 );
or g105 ( new_n277_, new_n270_, new_n276_ );
not g106 ( new_n278_, keyIn_0_22 );
not g107 ( new_n279_, N24 );
and g108 ( new_n280_, new_n279_, keyIn_0_4 );
not g109 ( new_n281_, N30 );
not g110 ( new_n282_, keyIn_0_4 );
and g111 ( new_n283_, new_n282_, N24 );
or g112 ( new_n284_, new_n283_, new_n281_ );
or g113 ( new_n285_, new_n284_, new_n280_ );
and g114 ( new_n286_, new_n285_, new_n278_ );
not g115 ( new_n287_, new_n280_ );
or g116 ( new_n288_, new_n279_, keyIn_0_4 );
and g117 ( new_n289_, new_n288_, N30 );
and g118 ( new_n290_, new_n289_, new_n287_ );
and g119 ( new_n291_, new_n290_, keyIn_0_22 );
or g120 ( new_n292_, new_n286_, new_n291_ );
and g121 ( new_n293_, new_n277_, new_n292_ );
and g122 ( new_n294_, new_n293_, new_n262_ );
and g123 ( new_n295_, new_n294_, new_n231_ );
and g124 ( new_n296_, new_n295_, new_n208_ );
and g125 ( new_n297_, new_n296_, new_n172_ );
not g126 ( new_n298_, new_n297_ );
or g127 ( new_n299_, new_n296_, new_n172_ );
and g128 ( N223, new_n298_, new_n299_ );
not g129 ( new_n301_, keyIn_0_76 );
not g130 ( new_n302_, keyIn_0_63 );
not g131 ( new_n303_, keyIn_0_52 );
not g132 ( new_n304_, keyIn_0_46 );
or g133 ( new_n305_, N223, new_n304_ );
not g134 ( new_n306_, new_n296_ );
and g135 ( new_n307_, new_n306_, keyIn_0_45 );
or g136 ( new_n308_, new_n307_, new_n297_ );
or g137 ( new_n309_, new_n308_, keyIn_0_46 );
and g138 ( new_n310_, new_n309_, new_n305_ );
and g139 ( new_n311_, new_n310_, new_n246_ );
not g140 ( new_n312_, new_n311_ );
or g141 ( new_n313_, new_n310_, new_n246_ );
and g142 ( new_n314_, new_n312_, new_n313_ );
and g143 ( new_n315_, new_n314_, new_n303_ );
not g144 ( new_n316_, new_n315_ );
or g145 ( new_n317_, new_n314_, new_n303_ );
and g146 ( new_n318_, new_n316_, new_n317_ );
not g147 ( new_n319_, new_n318_ );
not g148 ( new_n320_, N60 );
and g149 ( new_n321_, new_n234_, keyIn_0_9 );
not g150 ( new_n322_, new_n321_ );
or g151 ( new_n323_, new_n234_, keyIn_0_9 );
and g152 ( new_n324_, new_n322_, new_n323_ );
not g153 ( new_n325_, new_n324_ );
and g154 ( new_n326_, new_n325_, new_n320_ );
not g155 ( new_n327_, new_n326_ );
and g156 ( new_n328_, new_n327_, keyIn_0_35 );
not g157 ( new_n329_, new_n328_ );
or g158 ( new_n330_, new_n327_, keyIn_0_35 );
and g159 ( new_n331_, new_n329_, new_n330_ );
or g160 ( new_n332_, new_n319_, new_n331_ );
not g161 ( new_n333_, new_n332_ );
or g162 ( new_n334_, new_n333_, new_n302_ );
or g163 ( new_n335_, new_n332_, keyIn_0_63 );
and g164 ( new_n336_, new_n334_, new_n335_ );
not g165 ( new_n337_, keyIn_0_53 );
and g166 ( new_n338_, new_n310_, new_n261_ );
not g167 ( new_n339_, new_n338_ );
or g168 ( new_n340_, new_n310_, new_n261_ );
and g169 ( new_n341_, new_n339_, new_n340_ );
and g170 ( new_n342_, new_n341_, new_n337_ );
not g171 ( new_n343_, new_n342_ );
or g172 ( new_n344_, new_n341_, new_n337_ );
and g173 ( new_n345_, new_n343_, new_n344_ );
not g174 ( new_n346_, N73 );
and g175 ( new_n347_, keyIn_0_11, N69 );
not g176 ( new_n348_, new_n347_ );
or g177 ( new_n349_, keyIn_0_11, N69 );
and g178 ( new_n350_, new_n348_, new_n349_ );
and g179 ( new_n351_, new_n350_, new_n346_ );
not g180 ( new_n352_, new_n351_ );
and g181 ( new_n353_, new_n352_, keyIn_0_37 );
not g182 ( new_n354_, new_n353_ );
or g183 ( new_n355_, new_n352_, keyIn_0_37 );
and g184 ( new_n356_, new_n354_, new_n355_ );
not g185 ( new_n357_, new_n356_ );
and g186 ( new_n358_, new_n345_, new_n357_ );
not g187 ( new_n359_, new_n358_ );
or g188 ( new_n360_, new_n359_, keyIn_0_64 );
not g189 ( new_n361_, keyIn_0_64 );
or g190 ( new_n362_, new_n358_, new_n361_ );
and g191 ( new_n363_, new_n360_, new_n362_ );
not g192 ( new_n364_, keyIn_0_67 );
not g193 ( new_n365_, keyIn_0_56 );
not g194 ( new_n366_, new_n184_ );
and g195 ( new_n367_, new_n308_, keyIn_0_46 );
and g196 ( new_n368_, N223, new_n304_ );
or g197 ( new_n369_, new_n367_, new_n368_ );
and g198 ( new_n370_, new_n369_, new_n366_ );
and g199 ( new_n371_, new_n310_, new_n184_ );
or g200 ( new_n372_, new_n370_, new_n371_ );
and g201 ( new_n373_, new_n372_, new_n365_ );
not g202 ( new_n374_, new_n373_ );
or g203 ( new_n375_, new_n372_, new_n365_ );
and g204 ( new_n376_, new_n374_, new_n375_ );
not g205 ( new_n377_, N112 );
and g206 ( new_n378_, keyIn_0_17, N108 );
not g207 ( new_n379_, new_n378_ );
or g208 ( new_n380_, keyIn_0_17, N108 );
and g209 ( new_n381_, new_n379_, new_n380_ );
not g210 ( new_n382_, new_n381_ );
and g211 ( new_n383_, new_n382_, new_n377_ );
and g212 ( new_n384_, new_n383_, keyIn_0_43 );
not g213 ( new_n385_, new_n384_ );
or g214 ( new_n386_, new_n383_, keyIn_0_43 );
and g215 ( new_n387_, new_n385_, new_n386_ );
not g216 ( new_n388_, new_n387_ );
or g217 ( new_n389_, new_n376_, new_n388_ );
not g218 ( new_n390_, new_n389_ );
or g219 ( new_n391_, new_n390_, new_n364_ );
or g220 ( new_n392_, new_n389_, keyIn_0_67 );
and g221 ( new_n393_, new_n391_, new_n392_ );
and g222 ( new_n394_, new_n363_, new_n393_ );
and g223 ( new_n395_, new_n394_, new_n336_ );
not g224 ( new_n396_, keyIn_0_49 );
not g225 ( new_n397_, new_n230_ );
and g226 ( new_n398_, new_n369_, new_n397_ );
and g227 ( new_n399_, new_n310_, new_n230_ );
or g228 ( new_n400_, new_n398_, new_n399_ );
and g229 ( new_n401_, new_n400_, new_n396_ );
not g230 ( new_n402_, new_n401_ );
or g231 ( new_n403_, new_n400_, new_n396_ );
and g232 ( new_n404_, new_n402_, new_n403_ );
not g233 ( new_n405_, N21 );
and g234 ( new_n406_, keyIn_0_3, N17 );
not g235 ( new_n407_, new_n406_ );
or g236 ( new_n408_, keyIn_0_3, N17 );
and g237 ( new_n409_, new_n407_, new_n408_ );
not g238 ( new_n410_, new_n409_ );
and g239 ( new_n411_, new_n410_, new_n405_ );
not g240 ( new_n412_, new_n411_ );
and g241 ( new_n413_, new_n412_, keyIn_0_29 );
not g242 ( new_n414_, new_n413_ );
or g243 ( new_n415_, new_n412_, keyIn_0_29 );
and g244 ( new_n416_, new_n414_, new_n415_ );
not g245 ( new_n417_, new_n416_ );
and g246 ( new_n418_, new_n404_, new_n417_ );
not g247 ( new_n419_, new_n418_ );
or g248 ( new_n420_, new_n419_, keyIn_0_60 );
not g249 ( new_n421_, keyIn_0_60 );
or g250 ( new_n422_, new_n418_, new_n421_ );
and g251 ( new_n423_, new_n420_, new_n422_ );
not g252 ( new_n424_, new_n219_ );
and g253 ( new_n425_, new_n369_, new_n424_ );
and g254 ( new_n426_, new_n310_, new_n219_ );
or g255 ( new_n427_, new_n425_, new_n426_ );
and g256 ( new_n428_, new_n427_, keyIn_0_48 );
not g257 ( new_n429_, new_n428_ );
or g258 ( new_n430_, new_n427_, keyIn_0_48 );
and g259 ( new_n431_, new_n429_, new_n430_ );
not g260 ( new_n432_, N8 );
and g261 ( new_n433_, keyIn_0_1, N4 );
not g262 ( new_n434_, new_n433_ );
or g263 ( new_n435_, keyIn_0_1, N4 );
and g264 ( new_n436_, new_n434_, new_n435_ );
and g265 ( new_n437_, new_n436_, new_n432_ );
not g266 ( new_n438_, new_n437_ );
and g267 ( new_n439_, new_n438_, keyIn_0_19 );
not g268 ( new_n440_, new_n439_ );
or g269 ( new_n441_, new_n438_, keyIn_0_19 );
and g270 ( new_n442_, new_n440_, new_n441_ );
not g271 ( new_n443_, new_n442_ );
and g272 ( new_n444_, new_n431_, new_n443_ );
not g273 ( new_n445_, new_n444_ );
and g274 ( new_n446_, new_n445_, keyIn_0_58 );
not g275 ( new_n447_, keyIn_0_58 );
and g276 ( new_n448_, new_n444_, new_n447_ );
or g277 ( new_n449_, new_n446_, new_n448_ );
and g278 ( new_n450_, new_n423_, new_n449_ );
not g279 ( new_n451_, keyIn_0_61 );
not g280 ( new_n452_, keyIn_0_50 );
not g281 ( new_n453_, new_n292_ );
and g282 ( new_n454_, new_n369_, new_n453_ );
and g283 ( new_n455_, new_n310_, new_n292_ );
or g284 ( new_n456_, new_n454_, new_n455_ );
or g285 ( new_n457_, new_n456_, new_n452_ );
or g286 ( new_n458_, new_n310_, new_n292_ );
or g287 ( new_n459_, new_n369_, new_n453_ );
and g288 ( new_n460_, new_n459_, new_n458_ );
or g289 ( new_n461_, new_n460_, keyIn_0_50 );
and g290 ( new_n462_, new_n457_, new_n461_ );
and g291 ( new_n463_, keyIn_0_5, N30 );
not g292 ( new_n464_, new_n463_ );
not g293 ( new_n465_, N34 );
or g294 ( new_n466_, keyIn_0_5, N30 );
and g295 ( new_n467_, new_n466_, new_n465_ );
and g296 ( new_n468_, new_n467_, new_n464_ );
and g297 ( new_n469_, new_n468_, keyIn_0_31 );
not g298 ( new_n470_, new_n469_ );
or g299 ( new_n471_, new_n468_, keyIn_0_31 );
and g300 ( new_n472_, new_n470_, new_n471_ );
or g301 ( new_n473_, new_n462_, new_n472_ );
and g302 ( new_n474_, new_n473_, new_n451_ );
and g303 ( new_n475_, new_n460_, keyIn_0_50 );
and g304 ( new_n476_, new_n456_, new_n452_ );
or g305 ( new_n477_, new_n476_, new_n475_ );
not g306 ( new_n478_, new_n472_ );
and g307 ( new_n479_, new_n477_, new_n478_ );
and g308 ( new_n480_, new_n479_, keyIn_0_61 );
or g309 ( new_n481_, new_n474_, new_n480_ );
not g310 ( new_n482_, keyIn_0_62 );
not g311 ( new_n483_, keyIn_0_51 );
not g312 ( new_n484_, new_n277_ );
and g313 ( new_n485_, new_n369_, new_n484_ );
and g314 ( new_n486_, new_n310_, new_n277_ );
or g315 ( new_n487_, new_n485_, new_n486_ );
and g316 ( new_n488_, new_n487_, new_n483_ );
or g317 ( new_n489_, new_n310_, new_n277_ );
or g318 ( new_n490_, new_n369_, new_n484_ );
and g319 ( new_n491_, new_n490_, new_n489_ );
and g320 ( new_n492_, new_n491_, keyIn_0_51 );
or g321 ( new_n493_, new_n488_, new_n492_ );
not g322 ( new_n494_, keyIn_0_33 );
not g323 ( new_n495_, N47 );
and g324 ( new_n496_, keyIn_0_7, N43 );
not g325 ( new_n497_, new_n496_ );
or g326 ( new_n498_, keyIn_0_7, N43 );
and g327 ( new_n499_, new_n497_, new_n498_ );
not g328 ( new_n500_, new_n499_ );
and g329 ( new_n501_, new_n500_, new_n495_ );
not g330 ( new_n502_, new_n501_ );
and g331 ( new_n503_, new_n502_, new_n494_ );
and g332 ( new_n504_, new_n501_, keyIn_0_33 );
or g333 ( new_n505_, new_n503_, new_n504_ );
or g334 ( new_n506_, new_n493_, new_n505_ );
or g335 ( new_n507_, new_n506_, new_n482_ );
or g336 ( new_n508_, new_n491_, keyIn_0_51 );
or g337 ( new_n509_, new_n487_, new_n483_ );
and g338 ( new_n510_, new_n509_, new_n508_ );
not g339 ( new_n511_, new_n505_ );
and g340 ( new_n512_, new_n510_, new_n511_ );
or g341 ( new_n513_, new_n512_, keyIn_0_62 );
and g342 ( new_n514_, new_n507_, new_n513_ );
and g343 ( new_n515_, new_n481_, new_n514_ );
not g344 ( new_n516_, keyIn_0_66 );
not g345 ( new_n517_, new_n195_ );
and g346 ( new_n518_, new_n369_, new_n517_ );
and g347 ( new_n519_, new_n310_, new_n195_ );
or g348 ( new_n520_, new_n518_, new_n519_ );
and g349 ( new_n521_, new_n520_, keyIn_0_55 );
not g350 ( new_n522_, keyIn_0_55 );
or g351 ( new_n523_, new_n310_, new_n195_ );
or g352 ( new_n524_, new_n369_, new_n517_ );
and g353 ( new_n525_, new_n524_, new_n523_ );
and g354 ( new_n526_, new_n525_, new_n522_ );
or g355 ( new_n527_, new_n521_, new_n526_ );
not g356 ( new_n528_, keyIn_0_41 );
not g357 ( new_n529_, N99 );
and g358 ( new_n530_, keyIn_0_15, N95 );
not g359 ( new_n531_, new_n530_ );
or g360 ( new_n532_, keyIn_0_15, N95 );
and g361 ( new_n533_, new_n531_, new_n532_ );
not g362 ( new_n534_, new_n533_ );
and g363 ( new_n535_, new_n534_, new_n529_ );
not g364 ( new_n536_, new_n535_ );
and g365 ( new_n537_, new_n536_, new_n528_ );
and g366 ( new_n538_, new_n535_, keyIn_0_41 );
or g367 ( new_n539_, new_n537_, new_n538_ );
or g368 ( new_n540_, new_n527_, new_n539_ );
or g369 ( new_n541_, new_n540_, new_n516_ );
or g370 ( new_n542_, new_n525_, new_n522_ );
or g371 ( new_n543_, new_n520_, keyIn_0_55 );
and g372 ( new_n544_, new_n543_, new_n542_ );
not g373 ( new_n545_, new_n539_ );
and g374 ( new_n546_, new_n544_, new_n545_ );
or g375 ( new_n547_, new_n546_, keyIn_0_66 );
and g376 ( new_n548_, new_n541_, new_n547_ );
not g377 ( new_n549_, keyIn_0_54 );
not g378 ( new_n550_, new_n206_ );
and g379 ( new_n551_, new_n369_, new_n550_ );
and g380 ( new_n552_, new_n310_, new_n206_ );
or g381 ( new_n553_, new_n551_, new_n552_ );
and g382 ( new_n554_, new_n553_, new_n549_ );
or g383 ( new_n555_, new_n310_, new_n206_ );
or g384 ( new_n556_, new_n369_, new_n550_ );
and g385 ( new_n557_, new_n556_, new_n555_ );
and g386 ( new_n558_, new_n557_, keyIn_0_54 );
or g387 ( new_n559_, new_n554_, new_n558_ );
not g388 ( new_n560_, N86 );
and g389 ( new_n561_, keyIn_0_13, N82 );
not g390 ( new_n562_, new_n561_ );
or g391 ( new_n563_, keyIn_0_13, N82 );
and g392 ( new_n564_, new_n562_, new_n563_ );
and g393 ( new_n565_, new_n564_, new_n560_ );
not g394 ( new_n566_, new_n565_ );
and g395 ( new_n567_, new_n566_, keyIn_0_39 );
not g396 ( new_n568_, new_n567_ );
or g397 ( new_n569_, new_n566_, keyIn_0_39 );
and g398 ( new_n570_, new_n568_, new_n569_ );
or g399 ( new_n571_, new_n559_, new_n570_ );
or g400 ( new_n572_, new_n571_, keyIn_0_65 );
not g401 ( new_n573_, keyIn_0_65 );
or g402 ( new_n574_, new_n557_, keyIn_0_54 );
or g403 ( new_n575_, new_n553_, new_n549_ );
and g404 ( new_n576_, new_n575_, new_n574_ );
not g405 ( new_n577_, new_n570_ );
and g406 ( new_n578_, new_n576_, new_n577_ );
or g407 ( new_n579_, new_n578_, new_n573_ );
and g408 ( new_n580_, new_n572_, new_n579_ );
and g409 ( new_n581_, new_n548_, new_n580_ );
and g410 ( new_n582_, new_n515_, new_n581_ );
and g411 ( new_n583_, new_n582_, new_n450_ );
and g412 ( new_n584_, new_n583_, new_n395_ );
not g413 ( new_n585_, new_n584_ );
and g414 ( new_n586_, new_n585_, new_n301_ );
and g415 ( new_n587_, new_n584_, keyIn_0_76 );
or g416 ( N329, new_n586_, new_n587_ );
not g417 ( new_n589_, keyIn_0_107 );
not g418 ( new_n590_, keyIn_0_86 );
and g419 ( new_n591_, N329, new_n590_ );
or g420 ( new_n592_, new_n584_, keyIn_0_76 );
not g421 ( new_n593_, new_n587_ );
and g422 ( new_n594_, new_n593_, new_n592_ );
and g423 ( new_n595_, new_n594_, keyIn_0_86 );
or g424 ( new_n596_, new_n591_, new_n595_ );
and g425 ( new_n597_, new_n596_, new_n336_ );
not g426 ( new_n598_, new_n336_ );
or g427 ( new_n599_, new_n594_, keyIn_0_86 );
or g428 ( new_n600_, N329, new_n590_ );
and g429 ( new_n601_, new_n600_, new_n599_ );
and g430 ( new_n602_, new_n601_, new_n598_ );
or g431 ( new_n603_, new_n597_, new_n602_ );
not g432 ( new_n604_, new_n603_ );
and g433 ( new_n605_, new_n604_, keyIn_0_92 );
not g434 ( new_n606_, keyIn_0_92 );
and g435 ( new_n607_, new_n603_, new_n606_ );
not g436 ( new_n608_, N66 );
and g437 ( new_n609_, new_n325_, new_n608_ );
not g438 ( new_n610_, new_n609_ );
and g439 ( new_n611_, new_n610_, keyIn_0_36 );
not g440 ( new_n612_, new_n611_ );
or g441 ( new_n613_, new_n610_, keyIn_0_36 );
and g442 ( new_n614_, new_n612_, new_n613_ );
or g443 ( new_n615_, new_n319_, new_n614_ );
not g444 ( new_n616_, new_n615_ );
and g445 ( new_n617_, new_n616_, keyIn_0_71 );
not g446 ( new_n618_, new_n617_ );
or g447 ( new_n619_, new_n616_, keyIn_0_71 );
and g448 ( new_n620_, new_n618_, new_n619_ );
and g449 ( new_n621_, new_n620_, keyIn_0_81 );
not g450 ( new_n622_, new_n621_ );
or g451 ( new_n623_, new_n620_, keyIn_0_81 );
and g452 ( new_n624_, new_n622_, new_n623_ );
or g453 ( new_n625_, new_n607_, new_n624_ );
or g454 ( new_n626_, new_n625_, new_n605_ );
not g455 ( new_n627_, new_n626_ );
and g456 ( new_n628_, new_n627_, keyIn_0_102 );
not g457 ( new_n629_, keyIn_0_102 );
and g458 ( new_n630_, new_n626_, new_n629_ );
or g459 ( new_n631_, new_n628_, new_n630_ );
and g460 ( new_n632_, new_n596_, new_n449_ );
not g461 ( new_n633_, new_n632_ );
or g462 ( new_n634_, new_n596_, new_n449_ );
and g463 ( new_n635_, new_n633_, new_n634_ );
and g464 ( new_n636_, new_n635_, keyIn_0_88 );
not g465 ( new_n637_, new_n636_ );
or g466 ( new_n638_, new_n635_, keyIn_0_88 );
not g467 ( new_n639_, keyIn_0_77 );
not g468 ( new_n640_, keyIn_0_20 );
not g469 ( new_n641_, N14 );
and g470 ( new_n642_, new_n436_, new_n641_ );
and g471 ( new_n643_, new_n642_, new_n640_ );
not g472 ( new_n644_, new_n643_ );
or g473 ( new_n645_, new_n642_, new_n640_ );
and g474 ( new_n646_, new_n644_, new_n645_ );
and g475 ( new_n647_, new_n431_, new_n646_ );
and g476 ( new_n648_, new_n647_, keyIn_0_59 );
not g477 ( new_n649_, new_n648_ );
or g478 ( new_n650_, new_n647_, keyIn_0_59 );
and g479 ( new_n651_, new_n649_, new_n650_ );
and g480 ( new_n652_, new_n651_, new_n639_ );
not g481 ( new_n653_, new_n652_ );
or g482 ( new_n654_, new_n651_, new_n639_ );
and g483 ( new_n655_, new_n653_, new_n654_ );
and g484 ( new_n656_, new_n638_, new_n655_ );
and g485 ( new_n657_, new_n656_, new_n637_ );
not g486 ( new_n658_, new_n657_ );
and g487 ( new_n659_, new_n658_, keyIn_0_98 );
not g488 ( new_n660_, keyIn_0_98 );
and g489 ( new_n661_, new_n657_, new_n660_ );
or g490 ( new_n662_, new_n659_, new_n661_ );
not g491 ( new_n663_, keyIn_0_90 );
and g492 ( new_n664_, new_n596_, new_n481_ );
not g493 ( new_n665_, new_n664_ );
or g494 ( new_n666_, new_n596_, new_n481_ );
and g495 ( new_n667_, new_n665_, new_n666_ );
and g496 ( new_n668_, new_n667_, new_n663_ );
not g497 ( new_n669_, new_n668_ );
or g498 ( new_n670_, new_n667_, new_n663_ );
not g499 ( new_n671_, N40 );
and g500 ( new_n672_, new_n466_, new_n671_ );
and g501 ( new_n673_, new_n672_, new_n464_ );
and g502 ( new_n674_, new_n673_, keyIn_0_32 );
not g503 ( new_n675_, new_n674_ );
or g504 ( new_n676_, new_n673_, keyIn_0_32 );
and g505 ( new_n677_, new_n675_, new_n676_ );
or g506 ( new_n678_, new_n462_, new_n677_ );
and g507 ( new_n679_, new_n678_, keyIn_0_69 );
not g508 ( new_n680_, new_n679_ );
or g509 ( new_n681_, new_n678_, keyIn_0_69 );
and g510 ( new_n682_, new_n680_, new_n681_ );
and g511 ( new_n683_, new_n682_, keyIn_0_79 );
not g512 ( new_n684_, new_n683_ );
or g513 ( new_n685_, new_n682_, keyIn_0_79 );
and g514 ( new_n686_, new_n684_, new_n685_ );
and g515 ( new_n687_, new_n670_, new_n686_ );
and g516 ( new_n688_, new_n687_, new_n669_ );
not g517 ( new_n689_, new_n688_ );
and g518 ( new_n690_, new_n689_, keyIn_0_100 );
not g519 ( new_n691_, keyIn_0_100 );
and g520 ( new_n692_, new_n688_, new_n691_ );
or g521 ( new_n693_, new_n690_, new_n692_ );
and g522 ( new_n694_, new_n662_, new_n693_ );
and g523 ( new_n695_, new_n694_, new_n631_ );
not g524 ( new_n696_, keyIn_0_99 );
and g525 ( new_n697_, new_n596_, new_n423_ );
not g526 ( new_n698_, new_n697_ );
or g527 ( new_n699_, new_n596_, new_n423_ );
and g528 ( new_n700_, new_n698_, new_n699_ );
and g529 ( new_n701_, new_n700_, keyIn_0_89 );
not g530 ( new_n702_, new_n701_ );
or g531 ( new_n703_, new_n700_, keyIn_0_89 );
and g532 ( new_n704_, new_n702_, new_n703_ );
not g533 ( new_n705_, new_n704_ );
not g534 ( new_n706_, N27 );
and g535 ( new_n707_, new_n410_, new_n706_ );
not g536 ( new_n708_, new_n707_ );
and g537 ( new_n709_, new_n708_, keyIn_0_30 );
not g538 ( new_n710_, new_n709_ );
or g539 ( new_n711_, new_n708_, keyIn_0_30 );
and g540 ( new_n712_, new_n710_, new_n711_ );
and g541 ( new_n713_, new_n404_, new_n712_ );
and g542 ( new_n714_, new_n713_, keyIn_0_68 );
not g543 ( new_n715_, new_n714_ );
or g544 ( new_n716_, new_n713_, keyIn_0_68 );
and g545 ( new_n717_, new_n715_, new_n716_ );
and g546 ( new_n718_, new_n717_, keyIn_0_78 );
not g547 ( new_n719_, new_n718_ );
or g548 ( new_n720_, new_n717_, keyIn_0_78 );
and g549 ( new_n721_, new_n719_, new_n720_ );
not g550 ( new_n722_, new_n721_ );
and g551 ( new_n723_, new_n705_, new_n722_ );
or g552 ( new_n724_, new_n723_, new_n696_ );
not g553 ( new_n725_, keyIn_0_101 );
and g554 ( new_n726_, new_n596_, new_n514_ );
not g555 ( new_n727_, new_n726_ );
or g556 ( new_n728_, new_n596_, new_n514_ );
and g557 ( new_n729_, new_n727_, new_n728_ );
or g558 ( new_n730_, new_n729_, keyIn_0_91 );
not g559 ( new_n731_, new_n730_ );
and g560 ( new_n732_, new_n729_, keyIn_0_91 );
or g561 ( new_n733_, new_n731_, new_n732_ );
not g562 ( new_n734_, keyIn_0_70 );
not g563 ( new_n735_, N53 );
and g564 ( new_n736_, new_n500_, new_n735_ );
not g565 ( new_n737_, new_n736_ );
and g566 ( new_n738_, new_n737_, keyIn_0_34 );
not g567 ( new_n739_, new_n738_ );
or g568 ( new_n740_, new_n737_, keyIn_0_34 );
and g569 ( new_n741_, new_n739_, new_n740_ );
or g570 ( new_n742_, new_n493_, new_n741_ );
not g571 ( new_n743_, new_n742_ );
and g572 ( new_n744_, new_n743_, new_n734_ );
and g573 ( new_n745_, new_n742_, keyIn_0_70 );
or g574 ( new_n746_, new_n744_, new_n745_ );
not g575 ( new_n747_, new_n746_ );
and g576 ( new_n748_, new_n747_, keyIn_0_80 );
not g577 ( new_n749_, new_n748_ );
or g578 ( new_n750_, new_n747_, keyIn_0_80 );
and g579 ( new_n751_, new_n749_, new_n750_ );
not g580 ( new_n752_, new_n751_ );
and g581 ( new_n753_, new_n733_, new_n752_ );
or g582 ( new_n754_, new_n753_, new_n725_ );
and g583 ( new_n755_, new_n724_, new_n754_ );
or g584 ( new_n756_, new_n704_, new_n721_ );
or g585 ( new_n757_, new_n756_, keyIn_0_99 );
not g586 ( new_n758_, new_n732_ );
and g587 ( new_n759_, new_n758_, new_n730_ );
or g588 ( new_n760_, new_n759_, new_n751_ );
or g589 ( new_n761_, new_n760_, keyIn_0_101 );
and g590 ( new_n762_, new_n757_, new_n761_ );
and g591 ( new_n763_, new_n755_, new_n762_ );
not g592 ( new_n764_, new_n393_ );
or g593 ( new_n765_, new_n601_, new_n764_ );
or g594 ( new_n766_, new_n596_, new_n393_ );
and g595 ( new_n767_, new_n766_, new_n765_ );
and g596 ( new_n768_, new_n767_, keyIn_0_97 );
not g597 ( new_n769_, keyIn_0_97 );
and g598 ( new_n770_, new_n596_, new_n393_ );
and g599 ( new_n771_, new_n601_, new_n764_ );
or g600 ( new_n772_, new_n770_, new_n771_ );
and g601 ( new_n773_, new_n772_, new_n769_ );
not g602 ( new_n774_, N115 );
and g603 ( new_n775_, new_n382_, new_n774_ );
not g604 ( new_n776_, new_n775_ );
and g605 ( new_n777_, new_n776_, keyIn_0_44 );
not g606 ( new_n778_, new_n777_ );
or g607 ( new_n779_, new_n776_, keyIn_0_44 );
and g608 ( new_n780_, new_n778_, new_n779_ );
or g609 ( new_n781_, new_n376_, new_n780_ );
and g610 ( new_n782_, new_n781_, keyIn_0_75 );
not g611 ( new_n783_, new_n782_ );
or g612 ( new_n784_, new_n781_, keyIn_0_75 );
and g613 ( new_n785_, new_n783_, new_n784_ );
not g614 ( new_n786_, new_n785_ );
and g615 ( new_n787_, new_n786_, keyIn_0_85 );
not g616 ( new_n788_, new_n787_ );
or g617 ( new_n789_, new_n786_, keyIn_0_85 );
and g618 ( new_n790_, new_n788_, new_n789_ );
or g619 ( new_n791_, new_n773_, new_n790_ );
or g620 ( new_n792_, new_n791_, new_n768_ );
or g621 ( new_n793_, new_n792_, keyIn_0_106 );
not g622 ( new_n794_, keyIn_0_106 );
not g623 ( new_n795_, new_n768_ );
or g624 ( new_n796_, new_n767_, keyIn_0_97 );
not g625 ( new_n797_, new_n790_ );
and g626 ( new_n798_, new_n796_, new_n797_ );
and g627 ( new_n799_, new_n798_, new_n795_ );
or g628 ( new_n800_, new_n799_, new_n794_ );
and g629 ( new_n801_, new_n793_, new_n800_ );
and g630 ( new_n802_, new_n596_, new_n548_ );
not g631 ( new_n803_, new_n548_ );
and g632 ( new_n804_, new_n601_, new_n803_ );
or g633 ( new_n805_, new_n802_, new_n804_ );
or g634 ( new_n806_, new_n805_, keyIn_0_96 );
not g635 ( new_n807_, keyIn_0_96 );
or g636 ( new_n808_, new_n601_, new_n803_ );
or g637 ( new_n809_, new_n596_, new_n548_ );
and g638 ( new_n810_, new_n809_, new_n808_ );
or g639 ( new_n811_, new_n810_, new_n807_ );
and g640 ( new_n812_, new_n806_, new_n811_ );
not g641 ( new_n813_, keyIn_0_84 );
not g642 ( new_n814_, keyIn_0_74 );
not g643 ( new_n815_, N105 );
and g644 ( new_n816_, new_n534_, new_n815_ );
not g645 ( new_n817_, new_n816_ );
and g646 ( new_n818_, new_n817_, keyIn_0_42 );
not g647 ( new_n819_, new_n818_ );
or g648 ( new_n820_, new_n817_, keyIn_0_42 );
and g649 ( new_n821_, new_n819_, new_n820_ );
and g650 ( new_n822_, new_n544_, new_n821_ );
and g651 ( new_n823_, new_n822_, new_n814_ );
not g652 ( new_n824_, new_n823_ );
or g653 ( new_n825_, new_n822_, new_n814_ );
and g654 ( new_n826_, new_n824_, new_n825_ );
not g655 ( new_n827_, new_n826_ );
and g656 ( new_n828_, new_n827_, new_n813_ );
and g657 ( new_n829_, new_n826_, keyIn_0_84 );
or g658 ( new_n830_, new_n828_, new_n829_ );
or g659 ( new_n831_, new_n812_, new_n830_ );
or g660 ( new_n832_, new_n831_, keyIn_0_105 );
not g661 ( new_n833_, keyIn_0_105 );
and g662 ( new_n834_, new_n810_, new_n807_ );
and g663 ( new_n835_, new_n805_, keyIn_0_96 );
or g664 ( new_n836_, new_n835_, new_n834_ );
not g665 ( new_n837_, new_n830_ );
and g666 ( new_n838_, new_n836_, new_n837_ );
or g667 ( new_n839_, new_n838_, new_n833_ );
and g668 ( new_n840_, new_n832_, new_n839_ );
and g669 ( new_n841_, new_n801_, new_n840_ );
not g670 ( new_n842_, keyIn_0_103 );
not g671 ( new_n843_, keyIn_0_93 );
and g672 ( new_n844_, new_n596_, new_n363_ );
not g673 ( new_n845_, new_n363_ );
and g674 ( new_n846_, new_n601_, new_n845_ );
or g675 ( new_n847_, new_n844_, new_n846_ );
or g676 ( new_n848_, new_n847_, new_n843_ );
or g677 ( new_n849_, new_n601_, new_n845_ );
or g678 ( new_n850_, new_n596_, new_n363_ );
and g679 ( new_n851_, new_n850_, new_n849_ );
or g680 ( new_n852_, new_n851_, keyIn_0_93 );
and g681 ( new_n853_, new_n848_, new_n852_ );
not g682 ( new_n854_, keyIn_0_72 );
not g683 ( new_n855_, new_n344_ );
or g684 ( new_n856_, new_n855_, new_n342_ );
not g685 ( new_n857_, N79 );
and g686 ( new_n858_, new_n350_, new_n857_ );
not g687 ( new_n859_, new_n858_ );
and g688 ( new_n860_, new_n859_, keyIn_0_38 );
not g689 ( new_n861_, new_n860_ );
or g690 ( new_n862_, new_n859_, keyIn_0_38 );
and g691 ( new_n863_, new_n861_, new_n862_ );
or g692 ( new_n864_, new_n856_, new_n863_ );
not g693 ( new_n865_, new_n864_ );
and g694 ( new_n866_, new_n865_, new_n854_ );
and g695 ( new_n867_, new_n864_, keyIn_0_72 );
or g696 ( new_n868_, new_n866_, new_n867_ );
not g697 ( new_n869_, new_n868_ );
and g698 ( new_n870_, new_n869_, keyIn_0_82 );
not g699 ( new_n871_, new_n870_ );
or g700 ( new_n872_, new_n869_, keyIn_0_82 );
and g701 ( new_n873_, new_n871_, new_n872_ );
not g702 ( new_n874_, new_n873_ );
or g703 ( new_n875_, new_n853_, new_n874_ );
or g704 ( new_n876_, new_n875_, new_n842_ );
not g705 ( new_n877_, keyIn_0_104 );
not g706 ( new_n878_, keyIn_0_94 );
and g707 ( new_n879_, new_n596_, new_n580_ );
not g708 ( new_n880_, new_n580_ );
and g709 ( new_n881_, new_n601_, new_n880_ );
or g710 ( new_n882_, new_n879_, new_n881_ );
or g711 ( new_n883_, new_n882_, new_n878_ );
or g712 ( new_n884_, new_n601_, new_n880_ );
or g713 ( new_n885_, new_n596_, new_n580_ );
and g714 ( new_n886_, new_n885_, new_n884_ );
or g715 ( new_n887_, new_n886_, keyIn_0_94 );
and g716 ( new_n888_, new_n883_, new_n887_ );
not g717 ( new_n889_, keyIn_0_73 );
not g718 ( new_n890_, N92 );
and g719 ( new_n891_, new_n564_, new_n890_ );
not g720 ( new_n892_, new_n891_ );
and g721 ( new_n893_, new_n892_, keyIn_0_40 );
not g722 ( new_n894_, new_n893_ );
or g723 ( new_n895_, new_n892_, keyIn_0_40 );
and g724 ( new_n896_, new_n894_, new_n895_ );
or g725 ( new_n897_, new_n559_, new_n896_ );
not g726 ( new_n898_, new_n897_ );
and g727 ( new_n899_, new_n898_, new_n889_ );
and g728 ( new_n900_, new_n897_, keyIn_0_73 );
or g729 ( new_n901_, new_n899_, new_n900_ );
not g730 ( new_n902_, new_n901_ );
and g731 ( new_n903_, new_n902_, keyIn_0_83 );
not g732 ( new_n904_, new_n903_ );
or g733 ( new_n905_, new_n902_, keyIn_0_83 );
and g734 ( new_n906_, new_n904_, new_n905_ );
not g735 ( new_n907_, new_n906_ );
or g736 ( new_n908_, new_n888_, new_n907_ );
or g737 ( new_n909_, new_n908_, new_n877_ );
and g738 ( new_n910_, new_n876_, new_n909_ );
and g739 ( new_n911_, new_n851_, keyIn_0_93 );
and g740 ( new_n912_, new_n847_, new_n843_ );
or g741 ( new_n913_, new_n912_, new_n911_ );
and g742 ( new_n914_, new_n913_, new_n873_ );
or g743 ( new_n915_, new_n914_, keyIn_0_103 );
and g744 ( new_n916_, new_n886_, keyIn_0_94 );
and g745 ( new_n917_, new_n882_, new_n878_ );
or g746 ( new_n918_, new_n917_, new_n916_ );
and g747 ( new_n919_, new_n918_, new_n906_ );
or g748 ( new_n920_, new_n919_, keyIn_0_104 );
and g749 ( new_n921_, new_n915_, new_n920_ );
and g750 ( new_n922_, new_n910_, new_n921_ );
and g751 ( new_n923_, new_n841_, new_n922_ );
and g752 ( new_n924_, new_n923_, new_n763_ );
and g753 ( new_n925_, new_n924_, new_n695_ );
not g754 ( new_n926_, new_n925_ );
and g755 ( new_n927_, new_n926_, new_n589_ );
and g756 ( new_n928_, new_n925_, keyIn_0_107 );
or g757 ( N370, new_n927_, new_n928_ );
not g758 ( new_n930_, keyIn_0_120 );
not g759 ( new_n931_, keyIn_0_113 );
or g760 ( new_n932_, new_n925_, keyIn_0_107 );
not g761 ( new_n933_, new_n928_ );
and g762 ( new_n934_, new_n933_, new_n932_ );
or g763 ( new_n935_, new_n934_, keyIn_0_108 );
not g764 ( new_n936_, keyIn_0_108 );
or g765 ( new_n937_, N370, new_n936_ );
and g766 ( new_n938_, new_n937_, new_n935_ );
or g767 ( new_n939_, new_n938_, new_n735_ );
or g768 ( new_n940_, new_n939_, keyIn_0_109 );
not g769 ( new_n941_, keyIn_0_109 );
and g770 ( new_n942_, N370, new_n936_ );
and g771 ( new_n943_, new_n934_, keyIn_0_108 );
or g772 ( new_n944_, new_n942_, new_n943_ );
and g773 ( new_n945_, new_n944_, N53 );
or g774 ( new_n946_, new_n945_, new_n941_ );
and g775 ( new_n947_, new_n940_, new_n946_ );
and g776 ( new_n948_, N329, keyIn_0_87 );
not g777 ( new_n949_, new_n948_ );
or g778 ( new_n950_, N329, keyIn_0_87 );
and g779 ( new_n951_, new_n949_, new_n950_ );
not g780 ( new_n952_, new_n951_ );
and g781 ( new_n953_, new_n952_, N47 );
and g782 ( new_n954_, new_n953_, keyIn_0_95 );
not g783 ( new_n955_, new_n954_ );
or g784 ( new_n956_, new_n953_, keyIn_0_95 );
and g785 ( new_n957_, new_n955_, new_n956_ );
not g786 ( new_n958_, keyIn_0_57 );
and g787 ( new_n959_, N223, keyIn_0_47 );
not g788 ( new_n960_, new_n959_ );
or g789 ( new_n961_, N223, keyIn_0_47 );
and g790 ( new_n962_, new_n960_, new_n961_ );
and g791 ( new_n963_, new_n962_, N37 );
and g792 ( new_n964_, new_n963_, new_n958_ );
not g793 ( new_n965_, new_n964_ );
or g794 ( new_n966_, new_n963_, new_n958_ );
and g795 ( new_n967_, new_n965_, new_n966_ );
or g796 ( new_n968_, new_n967_, new_n271_ );
or g797 ( new_n969_, new_n957_, new_n968_ );
or g798 ( new_n970_, new_n947_, new_n969_ );
and g799 ( new_n971_, new_n970_, new_n931_ );
and g800 ( new_n972_, new_n945_, new_n941_ );
and g801 ( new_n973_, new_n939_, keyIn_0_109 );
or g802 ( new_n974_, new_n973_, new_n972_ );
not g803 ( new_n975_, new_n969_ );
and g804 ( new_n976_, new_n974_, new_n975_ );
and g805 ( new_n977_, new_n976_, keyIn_0_113 );
or g806 ( new_n978_, new_n971_, new_n977_ );
not g807 ( new_n979_, keyIn_0_114 );
and g808 ( new_n980_, new_n944_, N66 );
and g809 ( new_n981_, new_n952_, N60 );
and g810 ( new_n982_, new_n962_, N50 );
or g811 ( new_n983_, new_n982_, new_n234_ );
or g812 ( new_n984_, new_n981_, new_n983_ );
or g813 ( new_n985_, new_n980_, new_n984_ );
and g814 ( new_n986_, new_n985_, new_n979_ );
not g815 ( new_n987_, new_n986_ );
or g816 ( new_n988_, new_n985_, new_n979_ );
and g817 ( new_n989_, new_n987_, new_n988_ );
and g818 ( new_n990_, new_n978_, new_n989_ );
not g819 ( new_n991_, keyIn_0_111 );
and g820 ( new_n992_, new_n944_, N27 );
and g821 ( new_n993_, new_n952_, N21 );
not g822 ( new_n994_, N17 );
and g823 ( new_n995_, new_n962_, N11 );
or g824 ( new_n996_, new_n995_, new_n994_ );
or g825 ( new_n997_, new_n993_, new_n996_ );
or g826 ( new_n998_, new_n992_, new_n997_ );
and g827 ( new_n999_, new_n998_, new_n991_ );
not g828 ( new_n1000_, new_n999_ );
or g829 ( new_n1001_, new_n998_, new_n991_ );
and g830 ( new_n1002_, new_n1000_, new_n1001_ );
and g831 ( new_n1003_, new_n944_, N40 );
and g832 ( new_n1004_, new_n952_, N34 );
and g833 ( new_n1005_, new_n962_, N24 );
or g834 ( new_n1006_, new_n1005_, new_n281_ );
or g835 ( new_n1007_, new_n1004_, new_n1006_ );
or g836 ( new_n1008_, new_n1003_, new_n1007_ );
and g837 ( new_n1009_, new_n1008_, keyIn_0_112 );
not g838 ( new_n1010_, new_n1009_ );
or g839 ( new_n1011_, new_n1008_, keyIn_0_112 );
and g840 ( new_n1012_, new_n1010_, new_n1011_ );
and g841 ( new_n1013_, new_n1002_, new_n1012_ );
and g842 ( new_n1014_, new_n944_, N115 );
and g843 ( new_n1015_, new_n952_, N112 );
and g844 ( new_n1016_, new_n962_, N102 );
or g845 ( new_n1017_, new_n1016_, new_n175_ );
or g846 ( new_n1018_, new_n1015_, new_n1017_ );
or g847 ( new_n1019_, new_n1014_, new_n1018_ );
not g848 ( new_n1020_, new_n1019_ );
and g849 ( new_n1021_, new_n1020_, keyIn_0_118 );
not g850 ( new_n1022_, keyIn_0_118 );
and g851 ( new_n1023_, new_n1019_, new_n1022_ );
or g852 ( new_n1024_, new_n1021_, new_n1023_ );
and g853 ( new_n1025_, new_n944_, N105 );
and g854 ( new_n1026_, new_n952_, N99 );
and g855 ( new_n1027_, new_n962_, N89 );
or g856 ( new_n1028_, new_n1027_, new_n186_ );
or g857 ( new_n1029_, new_n1026_, new_n1028_ );
or g858 ( new_n1030_, new_n1025_, new_n1029_ );
not g859 ( new_n1031_, new_n1030_ );
and g860 ( new_n1032_, new_n1031_, keyIn_0_117 );
not g861 ( new_n1033_, keyIn_0_117 );
and g862 ( new_n1034_, new_n1030_, new_n1033_ );
or g863 ( new_n1035_, new_n1032_, new_n1034_ );
and g864 ( new_n1036_, new_n1024_, new_n1035_ );
not g865 ( new_n1037_, keyIn_0_115 );
and g866 ( new_n1038_, new_n944_, N79 );
and g867 ( new_n1039_, new_n952_, N73 );
and g868 ( new_n1040_, new_n962_, N63 );
or g869 ( new_n1041_, new_n1040_, new_n250_ );
or g870 ( new_n1042_, new_n1039_, new_n1041_ );
or g871 ( new_n1043_, new_n1038_, new_n1042_ );
not g872 ( new_n1044_, new_n1043_ );
or g873 ( new_n1045_, new_n1044_, new_n1037_ );
or g874 ( new_n1046_, new_n1043_, keyIn_0_115 );
and g875 ( new_n1047_, new_n1045_, new_n1046_ );
not g876 ( new_n1048_, keyIn_0_116 );
and g877 ( new_n1049_, new_n944_, N92 );
and g878 ( new_n1050_, new_n952_, N86 );
not g879 ( new_n1051_, N82 );
and g880 ( new_n1052_, new_n962_, N76 );
or g881 ( new_n1053_, new_n1052_, new_n1051_ );
or g882 ( new_n1054_, new_n1050_, new_n1053_ );
or g883 ( new_n1055_, new_n1049_, new_n1054_ );
not g884 ( new_n1056_, new_n1055_ );
or g885 ( new_n1057_, new_n1056_, new_n1048_ );
or g886 ( new_n1058_, new_n1055_, keyIn_0_116 );
and g887 ( new_n1059_, new_n1057_, new_n1058_ );
and g888 ( new_n1060_, new_n1047_, new_n1059_ );
and g889 ( new_n1061_, new_n1036_, new_n1060_ );
and g890 ( new_n1062_, new_n1061_, new_n1013_ );
and g891 ( new_n1063_, new_n1062_, new_n990_ );
and g892 ( new_n1064_, new_n1063_, keyIn_0_119 );
not g893 ( new_n1065_, new_n1064_ );
or g894 ( new_n1066_, new_n1063_, keyIn_0_119 );
not g895 ( new_n1067_, keyIn_0_110 );
and g896 ( new_n1068_, new_n944_, N14 );
and g897 ( new_n1069_, new_n952_, N8 );
not g898 ( new_n1070_, N4 );
and g899 ( new_n1071_, new_n962_, N1 );
or g900 ( new_n1072_, new_n1071_, new_n1070_ );
or g901 ( new_n1073_, new_n1069_, new_n1072_ );
or g902 ( new_n1074_, new_n1068_, new_n1073_ );
not g903 ( new_n1075_, new_n1074_ );
or g904 ( new_n1076_, new_n1075_, new_n1067_ );
or g905 ( new_n1077_, new_n1074_, keyIn_0_110 );
and g906 ( new_n1078_, new_n1076_, new_n1077_ );
and g907 ( new_n1079_, new_n1066_, new_n1078_ );
and g908 ( new_n1080_, new_n1079_, new_n1065_ );
and g909 ( new_n1081_, new_n1080_, new_n930_ );
not g910 ( new_n1082_, new_n1081_ );
or g911 ( new_n1083_, new_n1080_, new_n930_ );
and g912 ( N421, new_n1082_, new_n1083_ );
not g913 ( new_n1085_, keyIn_0_125 );
not g914 ( new_n1086_, keyIn_0_121 );
not g915 ( new_n1087_, new_n1012_ );
or g916 ( new_n1088_, new_n978_, new_n1087_ );
and g917 ( new_n1089_, new_n1088_, new_n1086_ );
or g918 ( new_n1090_, new_n976_, keyIn_0_113 );
or g919 ( new_n1091_, new_n970_, new_n931_ );
and g920 ( new_n1092_, new_n1091_, new_n1090_ );
and g921 ( new_n1093_, new_n1092_, new_n1012_ );
and g922 ( new_n1094_, new_n1093_, keyIn_0_121 );
or g923 ( new_n1095_, new_n1089_, new_n1094_ );
and g924 ( new_n1096_, new_n1013_, new_n989_ );
and g925 ( new_n1097_, new_n1095_, new_n1096_ );
not g926 ( new_n1098_, new_n1097_ );
and g927 ( new_n1099_, new_n1098_, new_n1085_ );
and g928 ( new_n1100_, new_n1097_, keyIn_0_125 );
or g929 ( N430, new_n1099_, new_n1100_ );
or g930 ( new_n1102_, new_n1092_, new_n1087_ );
not g931 ( new_n1103_, new_n989_ );
or g932 ( new_n1104_, new_n1103_, new_n1047_ );
or g933 ( new_n1105_, new_n1102_, new_n1104_ );
and g934 ( new_n1106_, new_n1105_, keyIn_0_122 );
not g935 ( new_n1107_, keyIn_0_122 );
and g936 ( new_n1108_, new_n978_, new_n1012_ );
not g937 ( new_n1109_, new_n1104_ );
and g938 ( new_n1110_, new_n1108_, new_n1109_ );
and g939 ( new_n1111_, new_n1110_, new_n1107_ );
or g940 ( new_n1112_, new_n1106_, new_n1111_ );
not g941 ( new_n1113_, new_n1013_ );
or g942 ( new_n1114_, new_n1092_, new_n1103_ );
or g943 ( new_n1115_, new_n1114_, new_n1059_ );
or g944 ( new_n1116_, new_n1115_, keyIn_0_123 );
not g945 ( new_n1117_, keyIn_0_123 );
not g946 ( new_n1118_, new_n1059_ );
and g947 ( new_n1119_, new_n990_, new_n1118_ );
or g948 ( new_n1120_, new_n1119_, new_n1117_ );
and g949 ( new_n1121_, new_n1116_, new_n1120_ );
or g950 ( new_n1122_, new_n1121_, new_n1113_ );
or g951 ( new_n1123_, new_n1122_, new_n1112_ );
or g952 ( new_n1124_, new_n1123_, keyIn_0_126 );
not g953 ( new_n1125_, keyIn_0_126 );
or g954 ( new_n1126_, new_n1110_, new_n1107_ );
not g955 ( new_n1127_, new_n1111_ );
and g956 ( new_n1128_, new_n1127_, new_n1126_ );
and g957 ( new_n1129_, new_n1119_, new_n1117_ );
and g958 ( new_n1130_, new_n1115_, keyIn_0_123 );
or g959 ( new_n1131_, new_n1130_, new_n1129_ );
and g960 ( new_n1132_, new_n1131_, new_n1013_ );
and g961 ( new_n1133_, new_n1132_, new_n1128_ );
or g962 ( new_n1134_, new_n1133_, new_n1125_ );
and g963 ( N431, new_n1124_, new_n1134_ );
not g964 ( new_n1136_, keyIn_0_127 );
or g965 ( new_n1137_, new_n1118_, new_n1035_ );
or g966 ( new_n1138_, new_n1102_, new_n1137_ );
and g967 ( new_n1139_, new_n1138_, keyIn_0_124 );
not g968 ( new_n1140_, new_n1139_ );
or g969 ( new_n1141_, new_n1138_, keyIn_0_124 );
and g970 ( new_n1142_, new_n1140_, new_n1141_ );
not g971 ( new_n1143_, new_n1002_ );
or g972 ( new_n1144_, new_n1093_, keyIn_0_121 );
or g973 ( new_n1145_, new_n1088_, new_n1086_ );
and g974 ( new_n1146_, new_n1145_, new_n1144_ );
or g975 ( new_n1147_, new_n1146_, new_n1143_ );
or g976 ( new_n1148_, new_n1147_, new_n1112_ );
or g977 ( new_n1149_, new_n1148_, new_n1142_ );
or g978 ( new_n1150_, new_n1149_, new_n1136_ );
not g979 ( new_n1151_, new_n1142_ );
and g980 ( new_n1152_, new_n1095_, new_n1002_ );
and g981 ( new_n1153_, new_n1128_, new_n1152_ );
and g982 ( new_n1154_, new_n1153_, new_n1151_ );
or g983 ( new_n1155_, new_n1154_, keyIn_0_127 );
and g984 ( N432, new_n1150_, new_n1155_ );
endmodule