module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n620_, new_n368_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n292_, new_n215_, new_n626_, new_n152_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n953_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n851_, new_n932_, new_n878_, new_n543_, new_n113_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n126_, new_n810_, new_n940_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n893_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n107_, new_n182_, new_n407_, new_n666_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n515_, new_n332_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n930_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n574_, new_n881_, new_n928_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n947_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n106_, keyIn_0_24 );
not g001 ( new_n107_, N65 );
or g002 ( new_n108_, new_n107_, N69 );
not g003 ( new_n109_, N69 );
or g004 ( new_n110_, new_n109_, N65 );
and g005 ( new_n111_, new_n108_, new_n110_ );
not g006 ( new_n112_, N77 );
and g007 ( new_n113_, new_n112_, N73 );
not g008 ( new_n114_, N73 );
and g009 ( new_n115_, new_n114_, N77 );
or g010 ( new_n116_, new_n113_, new_n115_ );
or g011 ( new_n117_, new_n116_, new_n111_ );
and g012 ( new_n118_, new_n109_, N65 );
and g013 ( new_n119_, new_n107_, N69 );
or g014 ( new_n120_, new_n118_, new_n119_ );
or g015 ( new_n121_, new_n114_, N77 );
or g016 ( new_n122_, new_n112_, N73 );
and g017 ( new_n123_, new_n121_, new_n122_ );
or g018 ( new_n124_, new_n120_, new_n123_ );
and g019 ( new_n125_, new_n117_, new_n124_ );
or g020 ( new_n126_, new_n125_, keyIn_0_4 );
not g021 ( new_n127_, keyIn_0_4 );
and g022 ( new_n128_, new_n120_, new_n123_ );
and g023 ( new_n129_, new_n116_, new_n111_ );
or g024 ( new_n130_, new_n128_, new_n129_ );
or g025 ( new_n131_, new_n130_, new_n127_ );
and g026 ( new_n132_, new_n131_, new_n126_ );
not g027 ( new_n133_, keyIn_0_5 );
not g028 ( new_n134_, N81 );
or g029 ( new_n135_, new_n134_, N85 );
not g030 ( new_n136_, N85 );
or g031 ( new_n137_, new_n136_, N81 );
and g032 ( new_n138_, new_n135_, new_n137_ );
not g033 ( new_n139_, N93 );
and g034 ( new_n140_, new_n139_, N89 );
not g035 ( new_n141_, N89 );
and g036 ( new_n142_, new_n141_, N93 );
or g037 ( new_n143_, new_n140_, new_n142_ );
or g038 ( new_n144_, new_n143_, new_n138_ );
and g039 ( new_n145_, new_n136_, N81 );
and g040 ( new_n146_, new_n134_, N85 );
or g041 ( new_n147_, new_n145_, new_n146_ );
or g042 ( new_n148_, new_n141_, N93 );
or g043 ( new_n149_, new_n139_, N89 );
and g044 ( new_n150_, new_n148_, new_n149_ );
or g045 ( new_n151_, new_n147_, new_n150_ );
and g046 ( new_n152_, new_n144_, new_n151_ );
and g047 ( new_n153_, new_n152_, new_n133_ );
and g048 ( new_n154_, new_n147_, new_n150_ );
and g049 ( new_n155_, new_n143_, new_n138_ );
or g050 ( new_n156_, new_n154_, new_n155_ );
and g051 ( new_n157_, new_n156_, keyIn_0_5 );
or g052 ( new_n158_, new_n157_, new_n153_ );
or g053 ( new_n159_, new_n158_, new_n132_ );
and g054 ( new_n160_, new_n130_, new_n127_ );
and g055 ( new_n161_, new_n125_, keyIn_0_4 );
or g056 ( new_n162_, new_n160_, new_n161_ );
or g057 ( new_n163_, new_n156_, keyIn_0_5 );
or g058 ( new_n164_, new_n152_, new_n133_ );
and g059 ( new_n165_, new_n163_, new_n164_ );
or g060 ( new_n166_, new_n162_, new_n165_ );
and g061 ( new_n167_, new_n159_, new_n166_ );
or g062 ( new_n168_, new_n167_, keyIn_0_20 );
not g063 ( new_n169_, keyIn_0_20 );
and g064 ( new_n170_, new_n162_, new_n165_ );
and g065 ( new_n171_, new_n158_, new_n132_ );
or g066 ( new_n172_, new_n170_, new_n171_ );
or g067 ( new_n173_, new_n172_, new_n169_ );
and g068 ( new_n174_, new_n173_, new_n168_ );
and g069 ( new_n175_, N129, N137 );
not g070 ( new_n176_, new_n175_ );
or g071 ( new_n177_, new_n174_, new_n176_ );
and g072 ( new_n178_, new_n172_, new_n169_ );
and g073 ( new_n179_, new_n167_, keyIn_0_20 );
or g074 ( new_n180_, new_n178_, new_n179_ );
or g075 ( new_n181_, new_n180_, new_n175_ );
and g076 ( new_n182_, new_n181_, new_n177_ );
or g077 ( new_n183_, new_n182_, new_n106_ );
and g078 ( new_n184_, new_n180_, new_n175_ );
and g079 ( new_n185_, new_n174_, new_n176_ );
or g080 ( new_n186_, new_n184_, new_n185_ );
or g081 ( new_n187_, new_n186_, keyIn_0_24 );
and g082 ( new_n188_, new_n187_, new_n183_ );
not g083 ( new_n189_, N49 );
and g084 ( new_n190_, new_n189_, N33 );
not g085 ( new_n191_, N33 );
and g086 ( new_n192_, new_n191_, N49 );
or g087 ( new_n193_, new_n190_, new_n192_ );
not g088 ( new_n194_, new_n193_ );
not g089 ( new_n195_, N17 );
and g090 ( new_n196_, new_n195_, N1 );
not g091 ( new_n197_, N1 );
and g092 ( new_n198_, new_n197_, N17 );
or g093 ( new_n199_, new_n196_, new_n198_ );
and g094 ( new_n200_, new_n194_, new_n199_ );
not g095 ( new_n201_, new_n200_ );
or g096 ( new_n202_, new_n194_, new_n199_ );
and g097 ( new_n203_, new_n201_, new_n202_ );
and g098 ( new_n204_, new_n203_, keyIn_0_8 );
not g099 ( new_n205_, new_n204_ );
or g100 ( new_n206_, new_n203_, keyIn_0_8 );
and g101 ( new_n207_, new_n205_, new_n206_ );
or g102 ( new_n208_, new_n188_, new_n207_ );
and g103 ( new_n209_, new_n186_, keyIn_0_24 );
and g104 ( new_n210_, new_n182_, new_n106_ );
or g105 ( new_n211_, new_n209_, new_n210_ );
not g106 ( new_n212_, new_n207_ );
or g107 ( new_n213_, new_n211_, new_n212_ );
and g108 ( new_n214_, new_n213_, new_n208_ );
and g109 ( new_n215_, new_n211_, new_n212_ );
and g110 ( new_n216_, new_n188_, new_n207_ );
or g111 ( new_n217_, new_n215_, new_n216_ );
not g112 ( new_n218_, keyIn_0_25 );
not g113 ( new_n219_, keyIn_0_21 );
not g114 ( new_n220_, N101 );
and g115 ( new_n221_, new_n220_, N97 );
not g116 ( new_n222_, N97 );
and g117 ( new_n223_, new_n222_, N101 );
or g118 ( new_n224_, new_n221_, new_n223_ );
not g119 ( new_n225_, N105 );
or g120 ( new_n226_, new_n225_, N109 );
not g121 ( new_n227_, N109 );
or g122 ( new_n228_, new_n227_, N105 );
and g123 ( new_n229_, new_n226_, new_n228_ );
and g124 ( new_n230_, new_n224_, new_n229_ );
or g125 ( new_n231_, new_n222_, N101 );
or g126 ( new_n232_, new_n220_, N97 );
and g127 ( new_n233_, new_n231_, new_n232_ );
and g128 ( new_n234_, new_n227_, N105 );
and g129 ( new_n235_, new_n225_, N109 );
or g130 ( new_n236_, new_n234_, new_n235_ );
and g131 ( new_n237_, new_n236_, new_n233_ );
or g132 ( new_n238_, new_n230_, new_n237_ );
and g133 ( new_n239_, new_n238_, keyIn_0_6 );
not g134 ( new_n240_, keyIn_0_6 );
or g135 ( new_n241_, new_n236_, new_n233_ );
or g136 ( new_n242_, new_n224_, new_n229_ );
and g137 ( new_n243_, new_n241_, new_n242_ );
and g138 ( new_n244_, new_n243_, new_n240_ );
or g139 ( new_n245_, new_n239_, new_n244_ );
not g140 ( new_n246_, keyIn_0_7 );
not g141 ( new_n247_, N117 );
and g142 ( new_n248_, new_n247_, N113 );
not g143 ( new_n249_, N113 );
and g144 ( new_n250_, new_n249_, N117 );
or g145 ( new_n251_, new_n248_, new_n250_ );
not g146 ( new_n252_, N121 );
or g147 ( new_n253_, new_n252_, N125 );
not g148 ( new_n254_, N125 );
or g149 ( new_n255_, new_n254_, N121 );
and g150 ( new_n256_, new_n253_, new_n255_ );
and g151 ( new_n257_, new_n251_, new_n256_ );
or g152 ( new_n258_, new_n249_, N117 );
or g153 ( new_n259_, new_n247_, N113 );
and g154 ( new_n260_, new_n258_, new_n259_ );
and g155 ( new_n261_, new_n254_, N121 );
and g156 ( new_n262_, new_n252_, N125 );
or g157 ( new_n263_, new_n261_, new_n262_ );
and g158 ( new_n264_, new_n263_, new_n260_ );
or g159 ( new_n265_, new_n257_, new_n264_ );
and g160 ( new_n266_, new_n265_, new_n246_ );
or g161 ( new_n267_, new_n263_, new_n260_ );
or g162 ( new_n268_, new_n251_, new_n256_ );
and g163 ( new_n269_, new_n267_, new_n268_ );
and g164 ( new_n270_, new_n269_, keyIn_0_7 );
or g165 ( new_n271_, new_n266_, new_n270_ );
or g166 ( new_n272_, new_n245_, new_n271_ );
or g167 ( new_n273_, new_n243_, new_n240_ );
or g168 ( new_n274_, new_n238_, keyIn_0_6 );
and g169 ( new_n275_, new_n274_, new_n273_ );
or g170 ( new_n276_, new_n269_, keyIn_0_7 );
or g171 ( new_n277_, new_n265_, new_n246_ );
and g172 ( new_n278_, new_n277_, new_n276_ );
or g173 ( new_n279_, new_n275_, new_n278_ );
and g174 ( new_n280_, new_n272_, new_n279_ );
and g175 ( new_n281_, new_n280_, new_n219_ );
and g176 ( new_n282_, new_n275_, new_n278_ );
and g177 ( new_n283_, new_n245_, new_n271_ );
or g178 ( new_n284_, new_n283_, new_n282_ );
and g179 ( new_n285_, new_n284_, keyIn_0_21 );
or g180 ( new_n286_, new_n281_, new_n285_ );
and g181 ( new_n287_, N130, N137 );
not g182 ( new_n288_, new_n287_ );
and g183 ( new_n289_, new_n286_, new_n288_ );
or g184 ( new_n290_, new_n284_, keyIn_0_21 );
or g185 ( new_n291_, new_n280_, new_n219_ );
and g186 ( new_n292_, new_n291_, new_n290_ );
and g187 ( new_n293_, new_n292_, new_n287_ );
or g188 ( new_n294_, new_n289_, new_n293_ );
and g189 ( new_n295_, new_n294_, new_n218_ );
or g190 ( new_n296_, new_n292_, new_n287_ );
or g191 ( new_n297_, new_n286_, new_n288_ );
and g192 ( new_n298_, new_n297_, new_n296_ );
and g193 ( new_n299_, new_n298_, keyIn_0_25 );
or g194 ( new_n300_, new_n295_, new_n299_ );
not g195 ( new_n301_, N53 );
and g196 ( new_n302_, new_n301_, N37 );
not g197 ( new_n303_, N37 );
and g198 ( new_n304_, new_n303_, N53 );
or g199 ( new_n305_, new_n302_, new_n304_ );
not g200 ( new_n306_, new_n305_ );
not g201 ( new_n307_, N21 );
and g202 ( new_n308_, new_n307_, N5 );
not g203 ( new_n309_, N5 );
and g204 ( new_n310_, new_n309_, N21 );
or g205 ( new_n311_, new_n308_, new_n310_ );
and g206 ( new_n312_, new_n306_, new_n311_ );
not g207 ( new_n313_, new_n312_ );
or g208 ( new_n314_, new_n306_, new_n311_ );
and g209 ( new_n315_, new_n313_, new_n314_ );
not g210 ( new_n316_, new_n315_ );
and g211 ( new_n317_, new_n316_, keyIn_0_9 );
not g212 ( new_n318_, new_n317_ );
or g213 ( new_n319_, new_n316_, keyIn_0_9 );
and g214 ( new_n320_, new_n318_, new_n319_ );
not g215 ( new_n321_, new_n320_ );
or g216 ( new_n322_, new_n300_, new_n321_ );
or g217 ( new_n323_, new_n298_, keyIn_0_25 );
or g218 ( new_n324_, new_n294_, new_n218_ );
and g219 ( new_n325_, new_n324_, new_n323_ );
or g220 ( new_n326_, new_n325_, new_n320_ );
and g221 ( new_n327_, new_n322_, new_n326_ );
or g222 ( new_n328_, new_n217_, new_n327_ );
not g223 ( new_n329_, keyIn_0_22 );
and g224 ( new_n330_, new_n162_, new_n245_ );
and g225 ( new_n331_, new_n132_, new_n275_ );
or g226 ( new_n332_, new_n330_, new_n331_ );
and g227 ( new_n333_, new_n332_, new_n329_ );
not g228 ( new_n334_, new_n333_ );
or g229 ( new_n335_, new_n332_, new_n329_ );
and g230 ( new_n336_, new_n334_, new_n335_ );
and g231 ( new_n337_, N131, N137 );
not g232 ( new_n338_, new_n337_ );
and g233 ( new_n339_, new_n336_, new_n338_ );
not g234 ( new_n340_, new_n339_ );
or g235 ( new_n341_, new_n336_, new_n338_ );
and g236 ( new_n342_, new_n340_, new_n341_ );
not g237 ( new_n343_, new_n342_ );
and g238 ( new_n344_, new_n343_, keyIn_0_26 );
not g239 ( new_n345_, keyIn_0_26 );
and g240 ( new_n346_, new_n342_, new_n345_ );
or g241 ( new_n347_, new_n344_, new_n346_ );
not g242 ( new_n348_, keyIn_0_10 );
not g243 ( new_n349_, N57 );
and g244 ( new_n350_, new_n349_, N41 );
not g245 ( new_n351_, N41 );
and g246 ( new_n352_, new_n351_, N57 );
or g247 ( new_n353_, new_n350_, new_n352_ );
not g248 ( new_n354_, new_n353_ );
not g249 ( new_n355_, N25 );
and g250 ( new_n356_, new_n355_, N9 );
not g251 ( new_n357_, N9 );
and g252 ( new_n358_, new_n357_, N25 );
or g253 ( new_n359_, new_n356_, new_n358_ );
and g254 ( new_n360_, new_n354_, new_n359_ );
not g255 ( new_n361_, new_n360_ );
or g256 ( new_n362_, new_n354_, new_n359_ );
and g257 ( new_n363_, new_n361_, new_n362_ );
not g258 ( new_n364_, new_n363_ );
and g259 ( new_n365_, new_n364_, new_n348_ );
and g260 ( new_n366_, new_n363_, keyIn_0_10 );
or g261 ( new_n367_, new_n365_, new_n366_ );
not g262 ( new_n368_, new_n367_ );
and g263 ( new_n369_, new_n347_, new_n368_ );
or g264 ( new_n370_, new_n342_, new_n345_ );
not g265 ( new_n371_, new_n346_ );
and g266 ( new_n372_, new_n371_, new_n370_ );
and g267 ( new_n373_, new_n372_, new_n367_ );
or g268 ( new_n374_, new_n369_, new_n373_ );
or g269 ( new_n375_, new_n328_, new_n374_ );
and g270 ( new_n376_, new_n325_, new_n320_ );
and g271 ( new_n377_, new_n300_, new_n321_ );
or g272 ( new_n378_, new_n377_, new_n376_ );
or g273 ( new_n379_, new_n378_, new_n214_ );
or g274 ( new_n380_, new_n379_, new_n374_ );
and g275 ( new_n381_, new_n375_, new_n380_ );
not g276 ( new_n382_, keyIn_0_27 );
and g277 ( new_n383_, new_n271_, new_n165_ );
and g278 ( new_n384_, new_n158_, new_n278_ );
or g279 ( new_n385_, new_n383_, new_n384_ );
and g280 ( new_n386_, new_n385_, keyIn_0_23 );
not g281 ( new_n387_, new_n386_ );
or g282 ( new_n388_, new_n385_, keyIn_0_23 );
and g283 ( new_n389_, new_n387_, new_n388_ );
and g284 ( new_n390_, N132, N137 );
and g285 ( new_n391_, new_n389_, new_n390_ );
not g286 ( new_n392_, new_n391_ );
or g287 ( new_n393_, new_n389_, new_n390_ );
and g288 ( new_n394_, new_n392_, new_n393_ );
not g289 ( new_n395_, new_n394_ );
and g290 ( new_n396_, new_n395_, new_n382_ );
and g291 ( new_n397_, new_n394_, keyIn_0_27 );
or g292 ( new_n398_, new_n396_, new_n397_ );
not g293 ( new_n399_, N61 );
and g294 ( new_n400_, new_n399_, N45 );
not g295 ( new_n401_, N45 );
and g296 ( new_n402_, new_n401_, N61 );
or g297 ( new_n403_, new_n400_, new_n402_ );
not g298 ( new_n404_, new_n403_ );
not g299 ( new_n405_, N29 );
and g300 ( new_n406_, new_n405_, N13 );
not g301 ( new_n407_, N13 );
and g302 ( new_n408_, new_n407_, N29 );
or g303 ( new_n409_, new_n406_, new_n408_ );
and g304 ( new_n410_, new_n404_, new_n409_ );
not g305 ( new_n411_, new_n410_ );
or g306 ( new_n412_, new_n404_, new_n409_ );
and g307 ( new_n413_, new_n411_, new_n412_ );
not g308 ( new_n414_, new_n413_ );
and g309 ( new_n415_, new_n414_, keyIn_0_11 );
not g310 ( new_n416_, new_n415_ );
or g311 ( new_n417_, new_n414_, keyIn_0_11 );
and g312 ( new_n418_, new_n416_, new_n417_ );
and g313 ( new_n419_, new_n398_, new_n418_ );
or g314 ( new_n420_, new_n394_, keyIn_0_27 );
not g315 ( new_n421_, new_n397_ );
and g316 ( new_n422_, new_n421_, new_n420_ );
not g317 ( new_n423_, new_n418_ );
and g318 ( new_n424_, new_n422_, new_n423_ );
or g319 ( new_n425_, new_n419_, new_n424_ );
or g320 ( new_n426_, new_n381_, new_n425_ );
or g321 ( new_n427_, new_n422_, new_n423_ );
or g322 ( new_n428_, new_n398_, new_n418_ );
and g323 ( new_n429_, new_n428_, new_n427_ );
or g324 ( new_n430_, new_n429_, new_n374_ );
or g325 ( new_n431_, new_n372_, new_n367_ );
or g326 ( new_n432_, new_n347_, new_n368_ );
and g327 ( new_n433_, new_n432_, new_n431_ );
or g328 ( new_n434_, new_n425_, new_n433_ );
and g329 ( new_n435_, new_n430_, new_n434_ );
and g330 ( new_n436_, new_n214_, new_n327_ );
not g331 ( new_n437_, new_n436_ );
or g332 ( new_n438_, new_n435_, new_n437_ );
and g333 ( new_n439_, new_n426_, new_n438_ );
or g334 ( new_n440_, new_n439_, new_n214_ );
not g335 ( new_n441_, keyIn_0_1 );
and g336 ( new_n442_, new_n307_, N17 );
and g337 ( new_n443_, new_n195_, N21 );
or g338 ( new_n444_, new_n442_, new_n443_ );
or g339 ( new_n445_, new_n355_, N29 );
or g340 ( new_n446_, new_n405_, N25 );
and g341 ( new_n447_, new_n445_, new_n446_ );
and g342 ( new_n448_, new_n444_, new_n447_ );
or g343 ( new_n449_, new_n195_, N21 );
or g344 ( new_n450_, new_n307_, N17 );
and g345 ( new_n451_, new_n449_, new_n450_ );
and g346 ( new_n452_, new_n405_, N25 );
and g347 ( new_n453_, new_n355_, N29 );
or g348 ( new_n454_, new_n452_, new_n453_ );
and g349 ( new_n455_, new_n454_, new_n451_ );
or g350 ( new_n456_, new_n448_, new_n455_ );
and g351 ( new_n457_, new_n456_, new_n441_ );
or g352 ( new_n458_, new_n454_, new_n451_ );
or g353 ( new_n459_, new_n444_, new_n447_ );
and g354 ( new_n460_, new_n458_, new_n459_ );
and g355 ( new_n461_, new_n460_, keyIn_0_1 );
or g356 ( new_n462_, new_n457_, new_n461_ );
and g357 ( new_n463_, new_n301_, N49 );
and g358 ( new_n464_, new_n189_, N53 );
or g359 ( new_n465_, new_n463_, new_n464_ );
or g360 ( new_n466_, new_n349_, N61 );
or g361 ( new_n467_, new_n399_, N57 );
and g362 ( new_n468_, new_n466_, new_n467_ );
and g363 ( new_n469_, new_n465_, new_n468_ );
or g364 ( new_n470_, new_n189_, N53 );
or g365 ( new_n471_, new_n301_, N49 );
and g366 ( new_n472_, new_n470_, new_n471_ );
and g367 ( new_n473_, new_n399_, N57 );
and g368 ( new_n474_, new_n349_, N61 );
or g369 ( new_n475_, new_n473_, new_n474_ );
and g370 ( new_n476_, new_n475_, new_n472_ );
or g371 ( new_n477_, new_n469_, new_n476_ );
or g372 ( new_n478_, new_n477_, keyIn_0_3 );
not g373 ( new_n479_, keyIn_0_3 );
or g374 ( new_n480_, new_n475_, new_n472_ );
or g375 ( new_n481_, new_n465_, new_n468_ );
and g376 ( new_n482_, new_n480_, new_n481_ );
or g377 ( new_n483_, new_n482_, new_n479_ );
and g378 ( new_n484_, new_n478_, new_n483_ );
and g379 ( new_n485_, new_n462_, new_n484_ );
or g380 ( new_n486_, new_n460_, keyIn_0_1 );
or g381 ( new_n487_, new_n456_, new_n441_ );
and g382 ( new_n488_, new_n487_, new_n486_ );
and g383 ( new_n489_, new_n482_, new_n479_ );
and g384 ( new_n490_, new_n477_, keyIn_0_3 );
or g385 ( new_n491_, new_n490_, new_n489_ );
and g386 ( new_n492_, new_n491_, new_n488_ );
or g387 ( new_n493_, new_n485_, new_n492_ );
and g388 ( new_n494_, new_n493_, keyIn_0_19 );
not g389 ( new_n495_, new_n494_ );
or g390 ( new_n496_, new_n493_, keyIn_0_19 );
and g391 ( new_n497_, new_n495_, new_n496_ );
and g392 ( new_n498_, N136, N137 );
and g393 ( new_n499_, new_n497_, new_n498_ );
not g394 ( new_n500_, new_n499_ );
or g395 ( new_n501_, new_n497_, new_n498_ );
and g396 ( new_n502_, new_n500_, new_n501_ );
not g397 ( new_n503_, new_n502_ );
and g398 ( new_n504_, new_n503_, keyIn_0_31 );
not g399 ( new_n505_, keyIn_0_31 );
and g400 ( new_n506_, new_n502_, new_n505_ );
or g401 ( new_n507_, new_n504_, new_n506_ );
not g402 ( new_n508_, keyIn_0_15 );
and g403 ( new_n509_, new_n254_, N109 );
and g404 ( new_n510_, new_n227_, N125 );
or g405 ( new_n511_, new_n509_, new_n510_ );
not g406 ( new_n512_, new_n511_ );
and g407 ( new_n513_, new_n139_, N77 );
and g408 ( new_n514_, new_n112_, N93 );
or g409 ( new_n515_, new_n513_, new_n514_ );
and g410 ( new_n516_, new_n512_, new_n515_ );
not g411 ( new_n517_, new_n516_ );
or g412 ( new_n518_, new_n512_, new_n515_ );
and g413 ( new_n519_, new_n517_, new_n518_ );
not g414 ( new_n520_, new_n519_ );
and g415 ( new_n521_, new_n520_, new_n508_ );
and g416 ( new_n522_, new_n519_, keyIn_0_15 );
or g417 ( new_n523_, new_n521_, new_n522_ );
not g418 ( new_n524_, new_n523_ );
or g419 ( new_n525_, new_n507_, new_n524_ );
or g420 ( new_n526_, new_n502_, new_n505_ );
not g421 ( new_n527_, new_n506_ );
and g422 ( new_n528_, new_n527_, new_n526_ );
or g423 ( new_n529_, new_n528_, new_n523_ );
and g424 ( new_n530_, new_n525_, new_n529_ );
not g425 ( new_n531_, keyIn_0_30 );
not g426 ( new_n532_, keyIn_0_2 );
and g427 ( new_n533_, new_n303_, N33 );
and g428 ( new_n534_, new_n191_, N37 );
or g429 ( new_n535_, new_n533_, new_n534_ );
or g430 ( new_n536_, new_n351_, N45 );
or g431 ( new_n537_, new_n401_, N41 );
and g432 ( new_n538_, new_n536_, new_n537_ );
and g433 ( new_n539_, new_n535_, new_n538_ );
or g434 ( new_n540_, new_n191_, N37 );
or g435 ( new_n541_, new_n303_, N33 );
and g436 ( new_n542_, new_n540_, new_n541_ );
and g437 ( new_n543_, new_n401_, N41 );
and g438 ( new_n544_, new_n351_, N45 );
or g439 ( new_n545_, new_n543_, new_n544_ );
and g440 ( new_n546_, new_n545_, new_n542_ );
or g441 ( new_n547_, new_n539_, new_n546_ );
and g442 ( new_n548_, new_n547_, new_n532_ );
or g443 ( new_n549_, new_n545_, new_n542_ );
or g444 ( new_n550_, new_n535_, new_n538_ );
and g445 ( new_n551_, new_n549_, new_n550_ );
and g446 ( new_n552_, new_n551_, keyIn_0_2 );
or g447 ( new_n553_, new_n548_, new_n552_ );
not g448 ( new_n554_, keyIn_0_0 );
and g449 ( new_n555_, new_n309_, N1 );
and g450 ( new_n556_, new_n197_, N5 );
or g451 ( new_n557_, new_n555_, new_n556_ );
or g452 ( new_n558_, new_n357_, N13 );
or g453 ( new_n559_, new_n407_, N9 );
and g454 ( new_n560_, new_n558_, new_n559_ );
and g455 ( new_n561_, new_n557_, new_n560_ );
or g456 ( new_n562_, new_n197_, N5 );
or g457 ( new_n563_, new_n309_, N1 );
and g458 ( new_n564_, new_n562_, new_n563_ );
and g459 ( new_n565_, new_n407_, N9 );
and g460 ( new_n566_, new_n357_, N13 );
or g461 ( new_n567_, new_n565_, new_n566_ );
and g462 ( new_n568_, new_n567_, new_n564_ );
or g463 ( new_n569_, new_n561_, new_n568_ );
or g464 ( new_n570_, new_n569_, new_n554_ );
or g465 ( new_n571_, new_n567_, new_n564_ );
or g466 ( new_n572_, new_n557_, new_n560_ );
and g467 ( new_n573_, new_n571_, new_n572_ );
or g468 ( new_n574_, new_n573_, keyIn_0_0 );
and g469 ( new_n575_, new_n570_, new_n574_ );
and g470 ( new_n576_, new_n553_, new_n575_ );
or g471 ( new_n577_, new_n551_, keyIn_0_2 );
or g472 ( new_n578_, new_n547_, new_n532_ );
and g473 ( new_n579_, new_n578_, new_n577_ );
and g474 ( new_n580_, new_n573_, keyIn_0_0 );
and g475 ( new_n581_, new_n569_, new_n554_ );
or g476 ( new_n582_, new_n581_, new_n580_ );
and g477 ( new_n583_, new_n582_, new_n579_ );
or g478 ( new_n584_, new_n576_, new_n583_ );
and g479 ( new_n585_, new_n584_, keyIn_0_18 );
not g480 ( new_n586_, new_n585_ );
or g481 ( new_n587_, new_n584_, keyIn_0_18 );
and g482 ( new_n588_, new_n586_, new_n587_ );
and g483 ( new_n589_, N135, N137 );
not g484 ( new_n590_, new_n589_ );
and g485 ( new_n591_, new_n588_, new_n590_ );
not g486 ( new_n592_, new_n591_ );
or g487 ( new_n593_, new_n588_, new_n590_ );
and g488 ( new_n594_, new_n592_, new_n593_ );
and g489 ( new_n595_, new_n594_, new_n531_ );
not g490 ( new_n596_, new_n595_ );
or g491 ( new_n597_, new_n594_, new_n531_ );
and g492 ( new_n598_, new_n596_, new_n597_ );
not g493 ( new_n599_, keyIn_0_14 );
and g494 ( new_n600_, new_n252_, N105 );
and g495 ( new_n601_, new_n225_, N121 );
or g496 ( new_n602_, new_n600_, new_n601_ );
not g497 ( new_n603_, new_n602_ );
and g498 ( new_n604_, new_n141_, N73 );
and g499 ( new_n605_, new_n114_, N89 );
or g500 ( new_n606_, new_n604_, new_n605_ );
and g501 ( new_n607_, new_n603_, new_n606_ );
not g502 ( new_n608_, new_n607_ );
or g503 ( new_n609_, new_n603_, new_n606_ );
and g504 ( new_n610_, new_n608_, new_n609_ );
not g505 ( new_n611_, new_n610_ );
and g506 ( new_n612_, new_n611_, new_n599_ );
and g507 ( new_n613_, new_n610_, keyIn_0_14 );
or g508 ( new_n614_, new_n612_, new_n613_ );
not g509 ( new_n615_, new_n614_ );
and g510 ( new_n616_, new_n598_, new_n615_ );
not g511 ( new_n617_, new_n593_ );
or g512 ( new_n618_, new_n617_, new_n591_ );
and g513 ( new_n619_, new_n618_, keyIn_0_30 );
or g514 ( new_n620_, new_n619_, new_n595_ );
and g515 ( new_n621_, new_n620_, new_n614_ );
or g516 ( new_n622_, new_n616_, new_n621_ );
and g517 ( new_n623_, new_n530_, new_n622_ );
or g518 ( new_n624_, new_n462_, new_n582_ );
or g519 ( new_n625_, new_n488_, new_n575_ );
and g520 ( new_n626_, new_n624_, new_n625_ );
and g521 ( new_n627_, new_n626_, keyIn_0_16 );
not g522 ( new_n628_, keyIn_0_16 );
and g523 ( new_n629_, new_n488_, new_n575_ );
and g524 ( new_n630_, new_n462_, new_n582_ );
or g525 ( new_n631_, new_n630_, new_n629_ );
and g526 ( new_n632_, new_n631_, new_n628_ );
or g527 ( new_n633_, new_n627_, new_n632_ );
and g528 ( new_n634_, N133, N137 );
and g529 ( new_n635_, new_n633_, new_n634_ );
or g530 ( new_n636_, new_n631_, new_n628_ );
or g531 ( new_n637_, new_n626_, keyIn_0_16 );
and g532 ( new_n638_, new_n637_, new_n636_ );
not g533 ( new_n639_, new_n634_ );
and g534 ( new_n640_, new_n638_, new_n639_ );
or g535 ( new_n641_, new_n635_, new_n640_ );
and g536 ( new_n642_, new_n641_, keyIn_0_28 );
not g537 ( new_n643_, keyIn_0_28 );
or g538 ( new_n644_, new_n638_, new_n639_ );
or g539 ( new_n645_, new_n633_, new_n634_ );
and g540 ( new_n646_, new_n645_, new_n644_ );
and g541 ( new_n647_, new_n646_, new_n643_ );
or g542 ( new_n648_, new_n642_, new_n647_ );
and g543 ( new_n649_, new_n249_, N97 );
and g544 ( new_n650_, new_n222_, N113 );
or g545 ( new_n651_, new_n649_, new_n650_ );
not g546 ( new_n652_, new_n651_ );
and g547 ( new_n653_, new_n134_, N65 );
and g548 ( new_n654_, new_n107_, N81 );
or g549 ( new_n655_, new_n653_, new_n654_ );
and g550 ( new_n656_, new_n652_, new_n655_ );
not g551 ( new_n657_, new_n656_ );
or g552 ( new_n658_, new_n652_, new_n655_ );
and g553 ( new_n659_, new_n657_, new_n658_ );
not g554 ( new_n660_, new_n659_ );
and g555 ( new_n661_, new_n660_, keyIn_0_12 );
not g556 ( new_n662_, new_n661_ );
or g557 ( new_n663_, new_n660_, keyIn_0_12 );
and g558 ( new_n664_, new_n662_, new_n663_ );
and g559 ( new_n665_, new_n648_, new_n664_ );
or g560 ( new_n666_, new_n646_, new_n643_ );
or g561 ( new_n667_, new_n641_, keyIn_0_28 );
and g562 ( new_n668_, new_n667_, new_n666_ );
not g563 ( new_n669_, new_n664_ );
and g564 ( new_n670_, new_n668_, new_n669_ );
or g565 ( new_n671_, new_n665_, new_n670_ );
not g566 ( new_n672_, keyIn_0_17 );
or g567 ( new_n673_, new_n491_, new_n553_ );
or g568 ( new_n674_, new_n484_, new_n579_ );
and g569 ( new_n675_, new_n673_, new_n674_ );
and g570 ( new_n676_, new_n675_, new_n672_ );
and g571 ( new_n677_, new_n484_, new_n579_ );
and g572 ( new_n678_, new_n491_, new_n553_ );
or g573 ( new_n679_, new_n678_, new_n677_ );
and g574 ( new_n680_, new_n679_, keyIn_0_17 );
or g575 ( new_n681_, new_n676_, new_n680_ );
and g576 ( new_n682_, N134, N137 );
not g577 ( new_n683_, new_n682_ );
and g578 ( new_n684_, new_n681_, new_n683_ );
or g579 ( new_n685_, new_n679_, keyIn_0_17 );
or g580 ( new_n686_, new_n675_, new_n672_ );
and g581 ( new_n687_, new_n686_, new_n685_ );
and g582 ( new_n688_, new_n687_, new_n682_ );
or g583 ( new_n689_, new_n684_, new_n688_ );
and g584 ( new_n690_, new_n689_, keyIn_0_29 );
not g585 ( new_n691_, keyIn_0_29 );
or g586 ( new_n692_, new_n687_, new_n682_ );
or g587 ( new_n693_, new_n681_, new_n683_ );
and g588 ( new_n694_, new_n693_, new_n692_ );
and g589 ( new_n695_, new_n694_, new_n691_ );
or g590 ( new_n696_, new_n690_, new_n695_ );
and g591 ( new_n697_, new_n247_, N101 );
and g592 ( new_n698_, new_n220_, N117 );
or g593 ( new_n699_, new_n697_, new_n698_ );
not g594 ( new_n700_, new_n699_ );
and g595 ( new_n701_, new_n136_, N69 );
and g596 ( new_n702_, new_n109_, N85 );
or g597 ( new_n703_, new_n701_, new_n702_ );
and g598 ( new_n704_, new_n700_, new_n703_ );
not g599 ( new_n705_, new_n704_ );
or g600 ( new_n706_, new_n700_, new_n703_ );
and g601 ( new_n707_, new_n705_, new_n706_ );
not g602 ( new_n708_, new_n707_ );
and g603 ( new_n709_, new_n708_, keyIn_0_13 );
not g604 ( new_n710_, new_n709_ );
or g605 ( new_n711_, new_n708_, keyIn_0_13 );
and g606 ( new_n712_, new_n710_, new_n711_ );
not g607 ( new_n713_, new_n712_ );
or g608 ( new_n714_, new_n696_, new_n713_ );
or g609 ( new_n715_, new_n694_, new_n691_ );
or g610 ( new_n716_, new_n689_, keyIn_0_29 );
and g611 ( new_n717_, new_n716_, new_n715_ );
or g612 ( new_n718_, new_n717_, new_n712_ );
and g613 ( new_n719_, new_n714_, new_n718_ );
and g614 ( new_n720_, new_n671_, new_n719_ );
and g615 ( new_n721_, new_n623_, new_n720_ );
not g616 ( new_n722_, new_n721_ );
or g617 ( new_n723_, new_n440_, new_n722_ );
and g618 ( new_n724_, new_n723_, N1 );
and g619 ( new_n725_, new_n378_, new_n214_ );
and g620 ( new_n726_, new_n725_, new_n433_ );
and g621 ( new_n727_, new_n217_, new_n327_ );
and g622 ( new_n728_, new_n727_, new_n433_ );
or g623 ( new_n729_, new_n726_, new_n728_ );
and g624 ( new_n730_, new_n729_, new_n429_ );
and g625 ( new_n731_, new_n425_, new_n433_ );
and g626 ( new_n732_, new_n429_, new_n374_ );
or g627 ( new_n733_, new_n732_, new_n731_ );
and g628 ( new_n734_, new_n733_, new_n436_ );
or g629 ( new_n735_, new_n730_, new_n734_ );
and g630 ( new_n736_, new_n735_, new_n217_ );
and g631 ( new_n737_, new_n736_, new_n721_ );
and g632 ( new_n738_, new_n737_, new_n197_ );
or g633 ( N724, new_n724_, new_n738_ );
or g634 ( new_n740_, new_n439_, new_n327_ );
or g635 ( new_n741_, new_n740_, new_n722_ );
and g636 ( new_n742_, new_n741_, N5 );
and g637 ( new_n743_, new_n735_, new_n378_ );
and g638 ( new_n744_, new_n743_, new_n721_ );
and g639 ( new_n745_, new_n744_, new_n309_ );
or g640 ( N725, new_n742_, new_n745_ );
or g641 ( new_n747_, new_n439_, new_n433_ );
or g642 ( new_n748_, new_n747_, new_n722_ );
and g643 ( new_n749_, new_n748_, N9 );
and g644 ( new_n750_, new_n735_, new_n374_ );
and g645 ( new_n751_, new_n750_, new_n721_ );
and g646 ( new_n752_, new_n751_, new_n357_ );
or g647 ( N726, new_n749_, new_n752_ );
or g648 ( new_n754_, new_n439_, new_n429_ );
or g649 ( new_n755_, new_n754_, new_n722_ );
and g650 ( new_n756_, new_n755_, N13 );
and g651 ( new_n757_, new_n735_, new_n425_ );
and g652 ( new_n758_, new_n757_, new_n721_ );
and g653 ( new_n759_, new_n758_, new_n407_ );
or g654 ( N727, new_n756_, new_n759_ );
and g655 ( new_n761_, new_n528_, new_n523_ );
and g656 ( new_n762_, new_n507_, new_n524_ );
or g657 ( new_n763_, new_n762_, new_n761_ );
or g658 ( new_n764_, new_n620_, new_n614_ );
or g659 ( new_n765_, new_n598_, new_n615_ );
and g660 ( new_n766_, new_n765_, new_n764_ );
and g661 ( new_n767_, new_n720_, new_n766_ );
and g662 ( new_n768_, new_n767_, new_n763_ );
not g663 ( new_n769_, new_n768_ );
or g664 ( new_n770_, new_n440_, new_n769_ );
and g665 ( new_n771_, new_n770_, N17 );
and g666 ( new_n772_, new_n736_, new_n768_ );
and g667 ( new_n773_, new_n772_, new_n195_ );
or g668 ( N728, new_n771_, new_n773_ );
or g669 ( new_n775_, new_n740_, new_n769_ );
and g670 ( new_n776_, new_n775_, N21 );
and g671 ( new_n777_, new_n743_, new_n768_ );
and g672 ( new_n778_, new_n777_, new_n307_ );
or g673 ( N729, new_n776_, new_n778_ );
or g674 ( new_n780_, new_n747_, new_n769_ );
and g675 ( new_n781_, new_n780_, N25 );
and g676 ( new_n782_, new_n750_, new_n768_ );
and g677 ( new_n783_, new_n782_, new_n355_ );
or g678 ( N730, new_n781_, new_n783_ );
or g679 ( new_n785_, new_n754_, new_n769_ );
and g680 ( new_n786_, new_n785_, N29 );
and g681 ( new_n787_, new_n757_, new_n768_ );
and g682 ( new_n788_, new_n787_, new_n405_ );
or g683 ( N731, new_n786_, new_n788_ );
or g684 ( new_n790_, new_n668_, new_n669_ );
or g685 ( new_n791_, new_n648_, new_n664_ );
and g686 ( new_n792_, new_n791_, new_n790_ );
and g687 ( new_n793_, new_n717_, new_n712_ );
and g688 ( new_n794_, new_n696_, new_n713_ );
or g689 ( new_n795_, new_n794_, new_n793_ );
and g690 ( new_n796_, new_n795_, new_n792_ );
and g691 ( new_n797_, new_n623_, new_n796_ );
not g692 ( new_n798_, new_n797_ );
or g693 ( new_n799_, new_n440_, new_n798_ );
and g694 ( new_n800_, new_n799_, N33 );
and g695 ( new_n801_, new_n736_, new_n797_ );
and g696 ( new_n802_, new_n801_, new_n191_ );
or g697 ( N732, new_n800_, new_n802_ );
or g698 ( new_n804_, new_n740_, new_n798_ );
and g699 ( new_n805_, new_n804_, N37 );
and g700 ( new_n806_, new_n743_, new_n797_ );
and g701 ( new_n807_, new_n806_, new_n303_ );
or g702 ( N733, new_n805_, new_n807_ );
or g703 ( new_n809_, new_n747_, new_n798_ );
and g704 ( new_n810_, new_n809_, N41 );
and g705 ( new_n811_, new_n750_, new_n797_ );
and g706 ( new_n812_, new_n811_, new_n351_ );
or g707 ( N734, new_n810_, new_n812_ );
or g708 ( new_n814_, new_n754_, new_n798_ );
and g709 ( new_n815_, new_n814_, N45 );
and g710 ( new_n816_, new_n757_, new_n797_ );
and g711 ( new_n817_, new_n816_, new_n401_ );
or g712 ( N735, new_n815_, new_n817_ );
and g713 ( new_n819_, new_n796_, new_n766_ );
and g714 ( new_n820_, new_n819_, new_n763_ );
not g715 ( new_n821_, new_n820_ );
or g716 ( new_n822_, new_n440_, new_n821_ );
and g717 ( new_n823_, new_n822_, N49 );
and g718 ( new_n824_, new_n736_, new_n820_ );
and g719 ( new_n825_, new_n824_, new_n189_ );
or g720 ( N736, new_n823_, new_n825_ );
or g721 ( new_n827_, new_n740_, new_n821_ );
and g722 ( new_n828_, new_n827_, N53 );
and g723 ( new_n829_, new_n743_, new_n820_ );
and g724 ( new_n830_, new_n829_, new_n301_ );
or g725 ( N737, new_n828_, new_n830_ );
or g726 ( new_n832_, new_n747_, new_n821_ );
and g727 ( new_n833_, new_n832_, N57 );
and g728 ( new_n834_, new_n750_, new_n820_ );
and g729 ( new_n835_, new_n834_, new_n349_ );
or g730 ( N738, new_n833_, new_n835_ );
or g731 ( new_n837_, new_n754_, new_n821_ );
and g732 ( new_n838_, new_n837_, N61 );
and g733 ( new_n839_, new_n757_, new_n820_ );
and g734 ( new_n840_, new_n839_, new_n399_ );
or g735 ( N739, new_n838_, new_n840_ );
or g736 ( new_n842_, new_n795_, new_n792_ );
or g737 ( new_n843_, new_n842_, new_n622_ );
or g738 ( new_n844_, new_n671_, new_n719_ );
or g739 ( new_n845_, new_n844_, new_n622_ );
and g740 ( new_n846_, new_n843_, new_n845_ );
or g741 ( new_n847_, new_n846_, new_n763_ );
or g742 ( new_n848_, new_n763_, new_n766_ );
or g743 ( new_n849_, new_n530_, new_n622_ );
and g744 ( new_n850_, new_n848_, new_n849_ );
and g745 ( new_n851_, new_n792_, new_n719_ );
not g746 ( new_n852_, new_n851_ );
or g747 ( new_n853_, new_n850_, new_n852_ );
and g748 ( new_n854_, new_n847_, new_n853_ );
or g749 ( new_n855_, new_n854_, new_n792_ );
and g750 ( new_n856_, new_n732_, new_n727_ );
not g751 ( new_n857_, new_n856_ );
or g752 ( new_n858_, new_n855_, new_n857_ );
and g753 ( new_n859_, new_n858_, N65 );
or g754 ( new_n860_, new_n767_, new_n819_ );
and g755 ( new_n861_, new_n860_, new_n530_ );
and g756 ( new_n862_, new_n763_, new_n766_ );
or g757 ( new_n863_, new_n862_, new_n623_ );
and g758 ( new_n864_, new_n863_, new_n851_ );
or g759 ( new_n865_, new_n861_, new_n864_ );
and g760 ( new_n866_, new_n865_, new_n671_ );
and g761 ( new_n867_, new_n866_, new_n856_ );
and g762 ( new_n868_, new_n867_, new_n107_ );
or g763 ( N740, new_n859_, new_n868_ );
or g764 ( new_n870_, new_n854_, new_n719_ );
or g765 ( new_n871_, new_n870_, new_n857_ );
and g766 ( new_n872_, new_n871_, N69 );
and g767 ( new_n873_, new_n865_, new_n795_ );
and g768 ( new_n874_, new_n873_, new_n856_ );
and g769 ( new_n875_, new_n874_, new_n109_ );
or g770 ( N741, new_n872_, new_n875_ );
or g771 ( new_n877_, new_n854_, new_n766_ );
or g772 ( new_n878_, new_n877_, new_n857_ );
and g773 ( new_n879_, new_n878_, N73 );
and g774 ( new_n880_, new_n865_, new_n622_ );
and g775 ( new_n881_, new_n880_, new_n856_ );
and g776 ( new_n882_, new_n881_, new_n114_ );
or g777 ( N742, new_n879_, new_n882_ );
or g778 ( new_n884_, new_n854_, new_n530_ );
or g779 ( new_n885_, new_n884_, new_n857_ );
and g780 ( new_n886_, new_n885_, N77 );
and g781 ( new_n887_, new_n865_, new_n763_ );
and g782 ( new_n888_, new_n887_, new_n856_ );
and g783 ( new_n889_, new_n888_, new_n112_ );
or g784 ( N743, new_n886_, new_n889_ );
and g785 ( new_n891_, new_n728_, new_n425_ );
not g786 ( new_n892_, new_n891_ );
or g787 ( new_n893_, new_n855_, new_n892_ );
and g788 ( new_n894_, new_n893_, N81 );
and g789 ( new_n895_, new_n866_, new_n891_ );
and g790 ( new_n896_, new_n895_, new_n134_ );
or g791 ( N744, new_n894_, new_n896_ );
or g792 ( new_n898_, new_n870_, new_n892_ );
and g793 ( new_n899_, new_n898_, N85 );
and g794 ( new_n900_, new_n873_, new_n891_ );
and g795 ( new_n901_, new_n900_, new_n136_ );
or g796 ( N745, new_n899_, new_n901_ );
or g797 ( new_n903_, new_n877_, new_n892_ );
and g798 ( new_n904_, new_n903_, N89 );
and g799 ( new_n905_, new_n880_, new_n891_ );
and g800 ( new_n906_, new_n905_, new_n141_ );
or g801 ( N746, new_n904_, new_n906_ );
or g802 ( new_n908_, new_n884_, new_n892_ );
and g803 ( new_n909_, new_n908_, N93 );
and g804 ( new_n910_, new_n887_, new_n891_ );
and g805 ( new_n911_, new_n910_, new_n139_ );
or g806 ( N747, new_n909_, new_n911_ );
and g807 ( new_n913_, new_n732_, new_n725_ );
not g808 ( new_n914_, new_n913_ );
or g809 ( new_n915_, new_n855_, new_n914_ );
and g810 ( new_n916_, new_n915_, N97 );
and g811 ( new_n917_, new_n866_, new_n913_ );
and g812 ( new_n918_, new_n917_, new_n222_ );
or g813 ( N748, new_n916_, new_n918_ );
or g814 ( new_n920_, new_n870_, new_n914_ );
and g815 ( new_n921_, new_n920_, N101 );
and g816 ( new_n922_, new_n873_, new_n913_ );
and g817 ( new_n923_, new_n922_, new_n220_ );
or g818 ( N749, new_n921_, new_n923_ );
or g819 ( new_n925_, new_n877_, new_n914_ );
and g820 ( new_n926_, new_n925_, N105 );
and g821 ( new_n927_, new_n880_, new_n913_ );
and g822 ( new_n928_, new_n927_, new_n225_ );
or g823 ( N750, new_n926_, new_n928_ );
or g824 ( new_n930_, new_n884_, new_n914_ );
and g825 ( new_n931_, new_n930_, N109 );
and g826 ( new_n932_, new_n887_, new_n913_ );
and g827 ( new_n933_, new_n932_, new_n227_ );
or g828 ( N751, new_n931_, new_n933_ );
and g829 ( new_n935_, new_n726_, new_n425_ );
not g830 ( new_n936_, new_n935_ );
or g831 ( new_n937_, new_n855_, new_n936_ );
and g832 ( new_n938_, new_n937_, N113 );
and g833 ( new_n939_, new_n866_, new_n935_ );
and g834 ( new_n940_, new_n939_, new_n249_ );
or g835 ( N752, new_n938_, new_n940_ );
or g836 ( new_n942_, new_n870_, new_n936_ );
and g837 ( new_n943_, new_n942_, N117 );
and g838 ( new_n944_, new_n873_, new_n935_ );
and g839 ( new_n945_, new_n944_, new_n247_ );
or g840 ( N753, new_n943_, new_n945_ );
or g841 ( new_n947_, new_n877_, new_n936_ );
and g842 ( new_n948_, new_n947_, N121 );
and g843 ( new_n949_, new_n880_, new_n935_ );
and g844 ( new_n950_, new_n949_, new_n252_ );
or g845 ( N754, new_n948_, new_n950_ );
or g846 ( new_n952_, new_n884_, new_n936_ );
and g847 ( new_n953_, new_n952_, N125 );
and g848 ( new_n954_, new_n887_, new_n935_ );
and g849 ( new_n955_, new_n954_, new_n254_ );
or g850 ( N755, new_n953_, new_n955_ );
endmodule