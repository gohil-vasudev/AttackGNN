module locked_c3540 (  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n137_, new_n138_, new_n140_, new_n141_, new_n142_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1108_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1133_, new_n1134_, new_n1135_;
  NOR2_X1 g000 ( .A1(G58), .A2(G68), .ZN(new_n137_) );
  INV_X1 g001 ( .A(new_n137_), .ZN(new_n138_) );
  NOR3_X1 g002 ( .A1(new_n138_), .A2(G50), .A3(G77), .ZN(G353) );
  INV_X1 g003 ( .A(G97), .ZN(new_n140_) );
  INV_X1 g004 ( .A(G107), .ZN(new_n141_) );
  NAND2_X1 g005 ( .A1(new_n140_), .A2(new_n141_), .ZN(new_n142_) );
  NAND2_X1 g006 ( .A1(new_n142_), .A2(G87), .ZN(G355) );
  INV_X1 g007 ( .A(KEYINPUT49), .ZN(new_n144_) );
  NAND2_X1 g008 ( .A1(G68), .A2(G238), .ZN(new_n145_) );
  NAND2_X1 g009 ( .A1(G77), .A2(G244), .ZN(new_n146_) );
  NAND2_X1 g010 ( .A1(G50), .A2(G226), .ZN(new_n147_) );
  NAND2_X1 g011 ( .A1(G58), .A2(G232), .ZN(new_n148_) );
  NAND4_X1 g012 ( .A1(new_n145_), .A2(new_n146_), .A3(new_n147_), .A4(new_n148_), .ZN(new_n149_) );
  NAND2_X1 g013 ( .A1(new_n149_), .A2(new_n144_), .ZN(new_n150_) );
  NOR2_X1 g014 ( .A1(new_n149_), .A2(new_n144_), .ZN(new_n151_) );
  NAND2_X1 g015 ( .A1(G87), .A2(G250), .ZN(new_n152_) );
  NAND2_X1 g016 ( .A1(G116), .A2(G270), .ZN(new_n153_) );
  NAND2_X1 g017 ( .A1(G97), .A2(G257), .ZN(new_n154_) );
  NAND3_X1 g018 ( .A1(new_n152_), .A2(new_n153_), .A3(new_n154_), .ZN(new_n155_) );
  NAND2_X1 g019 ( .A1(G107), .A2(G264), .ZN(new_n156_) );
  XOR2_X1 g020 ( .A(new_n156_), .B(KEYINPUT50), .Z(new_n157_) );
  NOR3_X1 g021 ( .A1(new_n157_), .A2(new_n151_), .A3(new_n155_), .ZN(new_n158_) );
  NAND2_X1 g022 ( .A1(new_n158_), .A2(new_n150_), .ZN(new_n159_) );
  NAND2_X1 g023 ( .A1(G1), .A2(G20), .ZN(new_n160_) );
  NAND2_X1 g024 ( .A1(new_n159_), .A2(new_n160_), .ZN(new_n161_) );
  INV_X1 g025 ( .A(KEYINPUT2), .ZN(new_n162_) );
  NAND2_X1 g026 ( .A1(G1), .A2(G13), .ZN(new_n163_) );
  NAND2_X1 g027 ( .A1(new_n163_), .A2(new_n162_), .ZN(new_n164_) );
  NAND3_X1 g028 ( .A1(G1), .A2(G13), .A3(KEYINPUT2), .ZN(new_n165_) );
  NAND2_X1 g029 ( .A1(new_n164_), .A2(new_n165_), .ZN(new_n166_) );
  NAND2_X1 g030 ( .A1(new_n166_), .A2(G20), .ZN(new_n167_) );
  INV_X1 g031 ( .A(new_n167_), .ZN(new_n168_) );
  INV_X1 g032 ( .A(G50), .ZN(new_n169_) );
  NOR2_X1 g033 ( .A1(new_n137_), .A2(new_n169_), .ZN(new_n170_) );
  NAND2_X1 g034 ( .A1(new_n168_), .A2(new_n170_), .ZN(new_n171_) );
  NOR2_X1 g035 ( .A1(new_n160_), .A2(G13), .ZN(new_n172_) );
  INV_X1 g036 ( .A(G257), .ZN(new_n173_) );
  INV_X1 g037 ( .A(G264), .ZN(new_n174_) );
  NAND2_X1 g038 ( .A1(new_n173_), .A2(new_n174_), .ZN(new_n175_) );
  NAND3_X1 g039 ( .A1(new_n172_), .A2(G250), .A3(new_n175_), .ZN(new_n176_) );
  NAND3_X1 g040 ( .A1(new_n161_), .A2(new_n171_), .A3(new_n176_), .ZN(new_n177_) );
  INV_X1 g041 ( .A(new_n177_), .ZN(G361) );
  XOR2_X1 g042 ( .A(G232), .B(G244), .Z(new_n179_) );
  XNOR2_X1 g043 ( .A(new_n179_), .B(G226), .ZN(new_n180_) );
  XNOR2_X1 g044 ( .A(new_n180_), .B(G238), .ZN(new_n181_) );
  XNOR2_X1 g045 ( .A(G264), .B(G270), .ZN(new_n182_) );
  XNOR2_X1 g046 ( .A(G250), .B(G257), .ZN(new_n183_) );
  XNOR2_X1 g047 ( .A(new_n182_), .B(new_n183_), .ZN(new_n184_) );
  XOR2_X1 g048 ( .A(new_n181_), .B(new_n184_), .Z(G358) );
  XOR2_X1 g049 ( .A(G97), .B(G107), .Z(new_n186_) );
  XNOR2_X1 g050 ( .A(new_n186_), .B(KEYINPUT51), .ZN(new_n187_) );
  XNOR2_X1 g051 ( .A(G87), .B(G116), .ZN(new_n188_) );
  XNOR2_X1 g052 ( .A(new_n187_), .B(new_n188_), .ZN(new_n189_) );
  XNOR2_X1 g053 ( .A(G50), .B(G77), .ZN(new_n190_) );
  XNOR2_X1 g054 ( .A(G58), .B(G68), .ZN(new_n191_) );
  XNOR2_X1 g055 ( .A(new_n190_), .B(new_n191_), .ZN(new_n192_) );
  XNOR2_X1 g056 ( .A(new_n189_), .B(new_n192_), .ZN(G351) );
  INV_X1 g057 ( .A(KEYINPUT4), .ZN(new_n194_) );
  XNOR2_X1 g058 ( .A(new_n163_), .B(KEYINPUT2), .ZN(new_n195_) );
  NAND4_X1 g059 ( .A1(G1), .A2(G20), .A3(G33), .A4(KEYINPUT3), .ZN(new_n196_) );
  INV_X1 g060 ( .A(KEYINPUT3), .ZN(new_n197_) );
  NAND3_X1 g061 ( .A1(G1), .A2(G20), .A3(G33), .ZN(new_n198_) );
  NAND2_X1 g062 ( .A1(new_n198_), .A2(new_n197_), .ZN(new_n199_) );
  NAND2_X1 g063 ( .A1(new_n199_), .A2(new_n196_), .ZN(new_n200_) );
  NAND2_X1 g064 ( .A1(new_n195_), .A2(new_n200_), .ZN(new_n201_) );
  NAND3_X1 g065 ( .A1(new_n201_), .A2(G20), .A3(new_n194_), .ZN(new_n202_) );
  NAND2_X1 g066 ( .A1(new_n201_), .A2(G20), .ZN(new_n203_) );
  NAND2_X1 g067 ( .A1(new_n203_), .A2(KEYINPUT4), .ZN(new_n204_) );
  NAND2_X1 g068 ( .A1(new_n204_), .A2(new_n202_), .ZN(new_n205_) );
  INV_X1 g069 ( .A(new_n205_), .ZN(new_n206_) );
  NAND2_X1 g070 ( .A1(new_n206_), .A2(new_n191_), .ZN(new_n207_) );
  INV_X1 g071 ( .A(new_n201_), .ZN(new_n208_) );
  INV_X1 g072 ( .A(G1), .ZN(new_n209_) );
  NAND2_X1 g073 ( .A1(new_n209_), .A2(G20), .ZN(new_n210_) );
  NAND2_X1 g074 ( .A1(new_n208_), .A2(new_n210_), .ZN(new_n211_) );
  INV_X1 g075 ( .A(new_n211_), .ZN(new_n212_) );
  NAND2_X1 g076 ( .A1(new_n212_), .A2(G58), .ZN(new_n213_) );
  INV_X1 g077 ( .A(G20), .ZN(new_n214_) );
  INV_X1 g078 ( .A(G33), .ZN(new_n215_) );
  NAND2_X1 g079 ( .A1(new_n166_), .A2(new_n215_), .ZN(new_n216_) );
  INV_X1 g080 ( .A(new_n216_), .ZN(new_n217_) );
  NAND2_X1 g081 ( .A1(new_n217_), .A2(new_n214_), .ZN(new_n218_) );
  INV_X1 g082 ( .A(new_n218_), .ZN(new_n219_) );
  NAND2_X1 g083 ( .A1(new_n219_), .A2(G159), .ZN(new_n220_) );
  NOR2_X1 g084 ( .A1(new_n215_), .A2(G20), .ZN(new_n221_) );
  NAND2_X1 g085 ( .A1(new_n166_), .A2(new_n221_), .ZN(new_n222_) );
  INV_X1 g086 ( .A(new_n222_), .ZN(new_n223_) );
  NAND2_X1 g087 ( .A1(new_n223_), .A2(G68), .ZN(new_n224_) );
  INV_X1 g088 ( .A(G58), .ZN(new_n225_) );
  NAND3_X1 g089 ( .A1(new_n209_), .A2(G13), .A3(G20), .ZN(new_n226_) );
  INV_X1 g090 ( .A(new_n226_), .ZN(new_n227_) );
  NAND2_X1 g091 ( .A1(new_n227_), .A2(new_n225_), .ZN(new_n228_) );
  NAND3_X1 g092 ( .A1(new_n220_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n229_) );
  INV_X1 g093 ( .A(new_n229_), .ZN(new_n230_) );
  NAND3_X1 g094 ( .A1(new_n230_), .A2(new_n207_), .A3(new_n213_), .ZN(new_n231_) );
  XOR2_X1 g095 ( .A(new_n231_), .B(KEYINPUT30), .Z(new_n232_) );
  INV_X1 g096 ( .A(new_n232_), .ZN(new_n233_) );
  INV_X1 g097 ( .A(KEYINPUT34), .ZN(new_n234_) );
  INV_X1 g098 ( .A(KEYINPUT32), .ZN(new_n235_) );
  NAND2_X1 g099 ( .A1(new_n217_), .A2(G1698), .ZN(new_n236_) );
  INV_X1 g100 ( .A(new_n236_), .ZN(new_n237_) );
  NAND2_X1 g101 ( .A1(new_n237_), .A2(G226), .ZN(new_n238_) );
  NAND2_X1 g102 ( .A1(new_n238_), .A2(new_n235_), .ZN(new_n239_) );
  NAND3_X1 g103 ( .A1(new_n237_), .A2(G226), .A3(KEYINPUT32), .ZN(new_n240_) );
  INV_X1 g104 ( .A(G1698), .ZN(new_n241_) );
  NAND3_X1 g105 ( .A1(new_n217_), .A2(G223), .A3(new_n241_), .ZN(new_n242_) );
  NAND4_X1 g106 ( .A1(new_n239_), .A2(KEYINPUT33), .A3(new_n240_), .A4(new_n242_), .ZN(new_n243_) );
  INV_X1 g107 ( .A(KEYINPUT33), .ZN(new_n244_) );
  NAND3_X1 g108 ( .A1(new_n239_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n245_) );
  NAND2_X1 g109 ( .A1(new_n245_), .A2(new_n244_), .ZN(new_n246_) );
  INV_X1 g110 ( .A(G41), .ZN(new_n247_) );
  INV_X1 g111 ( .A(G45), .ZN(new_n248_) );
  NAND2_X1 g112 ( .A1(new_n247_), .A2(new_n248_), .ZN(new_n249_) );
  NAND3_X1 g113 ( .A1(new_n249_), .A2(new_n209_), .A3(G274), .ZN(new_n250_) );
  NAND2_X1 g114 ( .A1(new_n249_), .A2(new_n209_), .ZN(new_n251_) );
  NAND2_X1 g115 ( .A1(G33), .A2(G41), .ZN(new_n252_) );
  NAND2_X1 g116 ( .A1(new_n166_), .A2(new_n252_), .ZN(new_n253_) );
  NAND2_X1 g117 ( .A1(new_n253_), .A2(new_n251_), .ZN(new_n254_) );
  INV_X1 g118 ( .A(new_n254_), .ZN(new_n255_) );
  NAND2_X1 g119 ( .A1(new_n255_), .A2(G232), .ZN(new_n256_) );
  NOR2_X1 g120 ( .A1(new_n215_), .A2(G41), .ZN(new_n257_) );
  NAND2_X1 g121 ( .A1(new_n166_), .A2(new_n257_), .ZN(new_n258_) );
  INV_X1 g122 ( .A(new_n258_), .ZN(new_n259_) );
  NAND2_X1 g123 ( .A1(new_n259_), .A2(G87), .ZN(new_n260_) );
  XOR2_X1 g124 ( .A(new_n260_), .B(KEYINPUT31), .Z(new_n261_) );
  NAND3_X1 g125 ( .A1(new_n261_), .A2(new_n250_), .A3(new_n256_), .ZN(new_n262_) );
  INV_X1 g126 ( .A(new_n262_), .ZN(new_n263_) );
  NAND3_X1 g127 ( .A1(new_n263_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n264_) );
  INV_X1 g128 ( .A(new_n264_), .ZN(new_n265_) );
  NAND2_X1 g129 ( .A1(new_n265_), .A2(G179), .ZN(new_n266_) );
  NAND2_X1 g130 ( .A1(new_n266_), .A2(new_n234_), .ZN(new_n267_) );
  NAND3_X1 g131 ( .A1(new_n265_), .A2(G179), .A3(KEYINPUT34), .ZN(new_n268_) );
  NAND2_X1 g132 ( .A1(new_n264_), .A2(G169), .ZN(new_n269_) );
  NAND3_X1 g133 ( .A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_) );
  NAND2_X1 g134 ( .A1(new_n270_), .A2(new_n233_), .ZN(new_n271_) );
  INV_X1 g135 ( .A(new_n271_), .ZN(new_n272_) );
  NAND2_X1 g136 ( .A1(new_n264_), .A2(G200), .ZN(new_n273_) );
  NAND2_X1 g137 ( .A1(new_n273_), .A2(KEYINPUT35), .ZN(new_n274_) );
  INV_X1 g138 ( .A(KEYINPUT35), .ZN(new_n275_) );
  NAND3_X1 g139 ( .A1(new_n264_), .A2(G200), .A3(new_n275_), .ZN(new_n276_) );
  NAND2_X1 g140 ( .A1(new_n265_), .A2(G190), .ZN(new_n277_) );
  NAND4_X1 g141 ( .A1(new_n274_), .A2(new_n232_), .A3(new_n277_), .A4(new_n276_), .ZN(new_n278_) );
  NAND3_X1 g142 ( .A1(new_n237_), .A2(G238), .A3(KEYINPUT6), .ZN(new_n279_) );
  INV_X1 g143 ( .A(KEYINPUT6), .ZN(new_n280_) );
  NAND3_X1 g144 ( .A1(new_n217_), .A2(G238), .A3(G1698), .ZN(new_n281_) );
  NAND2_X1 g145 ( .A1(new_n281_), .A2(new_n280_), .ZN(new_n282_) );
  NAND3_X1 g146 ( .A1(new_n217_), .A2(G232), .A3(new_n241_), .ZN(new_n283_) );
  NAND2_X1 g147 ( .A1(new_n259_), .A2(G107), .ZN(new_n284_) );
  NAND3_X1 g148 ( .A1(new_n283_), .A2(new_n250_), .A3(new_n284_), .ZN(new_n285_) );
  INV_X1 g149 ( .A(new_n285_), .ZN(new_n286_) );
  NAND4_X1 g150 ( .A1(new_n286_), .A2(new_n279_), .A3(KEYINPUT7), .A4(new_n282_), .ZN(new_n287_) );
  INV_X1 g151 ( .A(KEYINPUT7), .ZN(new_n288_) );
  NAND3_X1 g152 ( .A1(new_n286_), .A2(new_n279_), .A3(new_n282_), .ZN(new_n289_) );
  NAND2_X1 g153 ( .A1(new_n289_), .A2(new_n288_), .ZN(new_n290_) );
  NAND2_X1 g154 ( .A1(new_n255_), .A2(G244), .ZN(new_n291_) );
  NAND4_X1 g155 ( .A1(new_n290_), .A2(G179), .A3(new_n287_), .A4(new_n291_), .ZN(new_n292_) );
  NAND3_X1 g156 ( .A1(new_n290_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n293_) );
  NAND2_X1 g157 ( .A1(new_n293_), .A2(G169), .ZN(new_n294_) );
  NAND2_X1 g158 ( .A1(new_n294_), .A2(new_n292_), .ZN(new_n295_) );
  NAND2_X1 g159 ( .A1(new_n205_), .A2(new_n211_), .ZN(new_n296_) );
  NAND2_X1 g160 ( .A1(new_n296_), .A2(G77), .ZN(new_n297_) );
  NAND2_X1 g161 ( .A1(new_n219_), .A2(G58), .ZN(new_n298_) );
  NAND2_X1 g162 ( .A1(new_n223_), .A2(G87), .ZN(new_n299_) );
  INV_X1 g163 ( .A(G77), .ZN(new_n300_) );
  NAND2_X1 g164 ( .A1(new_n227_), .A2(new_n300_), .ZN(new_n301_) );
  NAND3_X1 g165 ( .A1(new_n298_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_) );
  INV_X1 g166 ( .A(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g167 ( .A1(new_n297_), .A2(new_n303_), .ZN(new_n304_) );
  NAND2_X1 g168 ( .A1(new_n295_), .A2(new_n304_), .ZN(new_n305_) );
  NAND4_X1 g169 ( .A1(new_n290_), .A2(G190), .A3(new_n287_), .A4(new_n291_), .ZN(new_n306_) );
  NAND2_X1 g170 ( .A1(new_n293_), .A2(G200), .ZN(new_n307_) );
  NAND4_X1 g171 ( .A1(new_n307_), .A2(new_n297_), .A3(new_n303_), .A4(new_n306_), .ZN(new_n308_) );
  NAND2_X1 g172 ( .A1(new_n305_), .A2(new_n308_), .ZN(new_n309_) );
  INV_X1 g173 ( .A(new_n309_), .ZN(new_n310_) );
  INV_X1 g174 ( .A(KEYINPUT37), .ZN(new_n311_) );
  NAND2_X1 g175 ( .A1(new_n296_), .A2(G50), .ZN(new_n312_) );
  NAND2_X1 g176 ( .A1(new_n206_), .A2(new_n138_), .ZN(new_n313_) );
  NAND2_X1 g177 ( .A1(new_n219_), .A2(G150), .ZN(new_n314_) );
  NAND2_X1 g178 ( .A1(new_n223_), .A2(G58), .ZN(new_n315_) );
  NAND2_X1 g179 ( .A1(new_n227_), .A2(new_n169_), .ZN(new_n316_) );
  NAND4_X1 g180 ( .A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_) );
  INV_X1 g181 ( .A(new_n317_), .ZN(new_n318_) );
  NAND2_X1 g182 ( .A1(new_n318_), .A2(new_n312_), .ZN(new_n319_) );
  INV_X1 g183 ( .A(G179), .ZN(new_n320_) );
  NAND2_X1 g184 ( .A1(new_n255_), .A2(G226), .ZN(new_n321_) );
  INV_X1 g185 ( .A(new_n321_), .ZN(new_n322_) );
  NAND3_X1 g186 ( .A1(new_n217_), .A2(G223), .A3(G1698), .ZN(new_n323_) );
  NAND2_X1 g187 ( .A1(new_n259_), .A2(G77), .ZN(new_n324_) );
  NAND3_X1 g188 ( .A1(new_n323_), .A2(new_n250_), .A3(new_n324_), .ZN(new_n325_) );
  INV_X1 g189 ( .A(KEYINPUT36), .ZN(new_n326_) );
  NAND3_X1 g190 ( .A1(new_n217_), .A2(G222), .A3(new_n241_), .ZN(new_n327_) );
  XNOR2_X1 g191 ( .A(new_n327_), .B(new_n326_), .ZN(new_n328_) );
  NOR3_X1 g192 ( .A1(new_n328_), .A2(new_n322_), .A3(new_n325_), .ZN(new_n329_) );
  NAND2_X1 g193 ( .A1(new_n329_), .A2(new_n320_), .ZN(new_n330_) );
  INV_X1 g194 ( .A(G169), .ZN(new_n331_) );
  INV_X1 g195 ( .A(new_n325_), .ZN(new_n332_) );
  XNOR2_X1 g196 ( .A(new_n327_), .B(KEYINPUT36), .ZN(new_n333_) );
  NAND3_X1 g197 ( .A1(new_n333_), .A2(new_n321_), .A3(new_n332_), .ZN(new_n334_) );
  NAND2_X1 g198 ( .A1(new_n334_), .A2(new_n331_), .ZN(new_n335_) );
  NAND2_X1 g199 ( .A1(new_n330_), .A2(new_n335_), .ZN(new_n336_) );
  INV_X1 g200 ( .A(new_n336_), .ZN(new_n337_) );
  NAND2_X1 g201 ( .A1(new_n337_), .A2(new_n319_), .ZN(new_n338_) );
  NAND2_X1 g202 ( .A1(new_n329_), .A2(G190), .ZN(new_n339_) );
  NAND2_X1 g203 ( .A1(new_n334_), .A2(G200), .ZN(new_n340_) );
  NAND4_X1 g204 ( .A1(new_n318_), .A2(new_n339_), .A3(new_n312_), .A4(new_n340_), .ZN(new_n341_) );
  NAND3_X1 g205 ( .A1(new_n338_), .A2(new_n311_), .A3(new_n341_), .ZN(new_n342_) );
  NAND2_X1 g206 ( .A1(new_n338_), .A2(new_n341_), .ZN(new_n343_) );
  NAND2_X1 g207 ( .A1(new_n343_), .A2(KEYINPUT37), .ZN(new_n344_) );
  NAND2_X1 g208 ( .A1(new_n344_), .A2(new_n342_), .ZN(new_n345_) );
  INV_X1 g209 ( .A(G68), .ZN(new_n346_) );
  NAND2_X1 g210 ( .A1(new_n205_), .A2(new_n226_), .ZN(new_n347_) );
  NAND2_X1 g211 ( .A1(new_n347_), .A2(new_n346_), .ZN(new_n348_) );
  NAND2_X1 g212 ( .A1(new_n212_), .A2(G68), .ZN(new_n349_) );
  INV_X1 g213 ( .A(new_n349_), .ZN(new_n350_) );
  NAND2_X1 g214 ( .A1(new_n219_), .A2(G50), .ZN(new_n351_) );
  NAND2_X1 g215 ( .A1(new_n223_), .A2(G77), .ZN(new_n352_) );
  NAND2_X1 g216 ( .A1(new_n351_), .A2(new_n352_), .ZN(new_n353_) );
  NOR2_X1 g217 ( .A1(new_n350_), .A2(new_n353_), .ZN(new_n354_) );
  NAND3_X1 g218 ( .A1(new_n217_), .A2(G226), .A3(new_n241_), .ZN(new_n355_) );
  NAND2_X1 g219 ( .A1(new_n259_), .A2(G97), .ZN(new_n356_) );
  NAND3_X1 g220 ( .A1(new_n355_), .A2(new_n250_), .A3(new_n356_), .ZN(new_n357_) );
  NAND2_X1 g221 ( .A1(new_n255_), .A2(G238), .ZN(new_n358_) );
  NAND3_X1 g222 ( .A1(new_n217_), .A2(G232), .A3(G1698), .ZN(new_n359_) );
  NAND2_X1 g223 ( .A1(new_n358_), .A2(new_n359_), .ZN(new_n360_) );
  NOR2_X1 g224 ( .A1(new_n360_), .A2(new_n357_), .ZN(new_n361_) );
  NAND2_X1 g225 ( .A1(new_n361_), .A2(G190), .ZN(new_n362_) );
  XNOR2_X1 g226 ( .A(new_n362_), .B(KEYINPUT28), .ZN(new_n363_) );
  INV_X1 g227 ( .A(G200), .ZN(new_n364_) );
  NOR2_X1 g228 ( .A1(new_n361_), .A2(new_n364_), .ZN(new_n365_) );
  XNOR2_X1 g229 ( .A(new_n365_), .B(KEYINPUT27), .ZN(new_n366_) );
  NAND4_X1 g230 ( .A1(new_n366_), .A2(new_n363_), .A3(new_n348_), .A4(new_n354_), .ZN(new_n367_) );
  INV_X1 g231 ( .A(new_n367_), .ZN(new_n368_) );
  NAND2_X1 g232 ( .A1(new_n354_), .A2(new_n348_), .ZN(new_n369_) );
  NOR3_X1 g233 ( .A1(new_n360_), .A2(new_n357_), .A3(G179), .ZN(new_n370_) );
  NOR2_X1 g234 ( .A1(new_n361_), .A2(G169), .ZN(new_n371_) );
  NOR2_X1 g235 ( .A1(new_n371_), .A2(new_n370_), .ZN(new_n372_) );
  NAND2_X1 g236 ( .A1(new_n372_), .A2(new_n369_), .ZN(new_n373_) );
  INV_X1 g237 ( .A(new_n373_), .ZN(new_n374_) );
  NOR2_X1 g238 ( .A1(new_n368_), .A2(new_n374_), .ZN(new_n375_) );
  NAND4_X1 g239 ( .A1(new_n345_), .A2(new_n278_), .A3(new_n310_), .A4(new_n375_), .ZN(new_n376_) );
  NOR2_X1 g240 ( .A1(new_n376_), .A2(new_n272_), .ZN(new_n377_) );
  INV_X1 g241 ( .A(new_n377_), .ZN(new_n378_) );
  NAND2_X1 g242 ( .A1(new_n347_), .A2(new_n141_), .ZN(new_n379_) );
  INV_X1 g243 ( .A(KEYINPUT17), .ZN(new_n380_) );
  NAND2_X1 g244 ( .A1(new_n209_), .A2(G33), .ZN(new_n381_) );
  NAND2_X1 g245 ( .A1(new_n226_), .A2(new_n381_), .ZN(new_n382_) );
  INV_X1 g246 ( .A(new_n382_), .ZN(new_n383_) );
  NAND4_X1 g247 ( .A1(new_n383_), .A2(new_n195_), .A3(G107), .A4(new_n200_), .ZN(new_n384_) );
  INV_X1 g248 ( .A(KEYINPUT16), .ZN(new_n385_) );
  NAND4_X1 g249 ( .A1(new_n166_), .A2(G116), .A3(new_n385_), .A4(new_n221_), .ZN(new_n386_) );
  NAND3_X1 g250 ( .A1(new_n166_), .A2(G116), .A3(new_n221_), .ZN(new_n387_) );
  NAND2_X1 g251 ( .A1(new_n387_), .A2(KEYINPUT16), .ZN(new_n388_) );
  NAND2_X1 g252 ( .A1(new_n388_), .A2(new_n386_), .ZN(new_n389_) );
  NAND3_X1 g253 ( .A1(new_n389_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n390_) );
  NAND2_X1 g254 ( .A1(new_n389_), .A2(new_n384_), .ZN(new_n391_) );
  NAND2_X1 g255 ( .A1(new_n391_), .A2(KEYINPUT17), .ZN(new_n392_) );
  NAND2_X1 g256 ( .A1(new_n392_), .A2(new_n390_), .ZN(new_n393_) );
  NAND2_X1 g257 ( .A1(new_n219_), .A2(G87), .ZN(new_n394_) );
  NAND3_X1 g258 ( .A1(new_n379_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_) );
  INV_X1 g259 ( .A(KEYINPUT15), .ZN(new_n396_) );
  INV_X1 g260 ( .A(KEYINPUT14), .ZN(new_n397_) );
  NAND3_X1 g261 ( .A1(new_n247_), .A2(G33), .A3(G294), .ZN(new_n398_) );
  INV_X1 g262 ( .A(new_n398_), .ZN(new_n399_) );
  NAND3_X1 g263 ( .A1(new_n166_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_) );
  NAND2_X1 g264 ( .A1(new_n166_), .A2(new_n399_), .ZN(new_n401_) );
  NAND2_X1 g265 ( .A1(new_n401_), .A2(KEYINPUT14), .ZN(new_n402_) );
  NAND2_X1 g266 ( .A1(new_n402_), .A2(new_n400_), .ZN(new_n403_) );
  NOR3_X1 g267 ( .A1(new_n248_), .A2(G1), .A3(G41), .ZN(new_n404_) );
  NAND2_X1 g268 ( .A1(new_n404_), .A2(G274), .ZN(new_n405_) );
  NOR2_X1 g269 ( .A1(new_n404_), .A2(new_n174_), .ZN(new_n406_) );
  NAND2_X1 g270 ( .A1(new_n253_), .A2(new_n406_), .ZN(new_n407_) );
  NAND4_X1 g271 ( .A1(new_n166_), .A2(new_n215_), .A3(G257), .A4(G1698), .ZN(new_n408_) );
  NAND4_X1 g272 ( .A1(new_n166_), .A2(new_n215_), .A3(G250), .A4(new_n241_), .ZN(new_n409_) );
  NAND2_X1 g273 ( .A1(new_n408_), .A2(new_n409_), .ZN(new_n410_) );
  INV_X1 g274 ( .A(new_n410_), .ZN(new_n411_) );
  NAND4_X1 g275 ( .A1(new_n411_), .A2(new_n403_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n412_) );
  INV_X1 g276 ( .A(new_n412_), .ZN(new_n413_) );
  NAND3_X1 g277 ( .A1(new_n413_), .A2(new_n320_), .A3(new_n396_), .ZN(new_n414_) );
  NAND2_X1 g278 ( .A1(new_n407_), .A2(new_n405_), .ZN(new_n415_) );
  INV_X1 g279 ( .A(new_n415_), .ZN(new_n416_) );
  NAND4_X1 g280 ( .A1(new_n416_), .A2(new_n320_), .A3(new_n403_), .A4(new_n411_), .ZN(new_n417_) );
  NAND2_X1 g281 ( .A1(new_n417_), .A2(KEYINPUT15), .ZN(new_n418_) );
  NAND2_X1 g282 ( .A1(new_n412_), .A2(new_n331_), .ZN(new_n419_) );
  NAND2_X1 g283 ( .A1(new_n418_), .A2(new_n419_), .ZN(new_n420_) );
  INV_X1 g284 ( .A(new_n420_), .ZN(new_n421_) );
  NAND3_X1 g285 ( .A1(new_n421_), .A2(new_n395_), .A3(new_n414_), .ZN(new_n422_) );
  NAND4_X1 g286 ( .A1(new_n416_), .A2(G190), .A3(new_n403_), .A4(new_n411_), .ZN(new_n423_) );
  NAND2_X1 g287 ( .A1(new_n412_), .A2(G200), .ZN(new_n424_) );
  NAND2_X1 g288 ( .A1(new_n424_), .A2(new_n423_), .ZN(new_n425_) );
  INV_X1 g289 ( .A(new_n425_), .ZN(new_n426_) );
  NAND4_X1 g290 ( .A1(new_n426_), .A2(new_n379_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n427_) );
  NAND3_X1 g291 ( .A1(new_n422_), .A2(new_n427_), .A3(KEYINPUT0), .ZN(new_n428_) );
  INV_X1 g292 ( .A(KEYINPUT0), .ZN(new_n429_) );
  NAND2_X1 g293 ( .A1(new_n422_), .A2(new_n427_), .ZN(new_n430_) );
  NAND2_X1 g294 ( .A1(new_n430_), .A2(new_n429_), .ZN(new_n431_) );
  NAND2_X1 g295 ( .A1(new_n431_), .A2(new_n428_), .ZN(new_n432_) );
  INV_X1 g296 ( .A(new_n432_), .ZN(new_n433_) );
  NAND3_X1 g297 ( .A1(new_n217_), .A2(G244), .A3(new_n241_), .ZN(new_n434_) );
  NAND3_X1 g298 ( .A1(new_n217_), .A2(G250), .A3(G1698), .ZN(new_n435_) );
  NAND2_X1 g299 ( .A1(new_n259_), .A2(G283), .ZN(new_n436_) );
  NAND4_X1 g300 ( .A1(new_n434_), .A2(new_n435_), .A3(new_n405_), .A4(new_n436_), .ZN(new_n437_) );
  NOR2_X1 g301 ( .A1(new_n437_), .A2(KEYINPUT12), .ZN(new_n438_) );
  INV_X1 g302 ( .A(new_n438_), .ZN(new_n439_) );
  NAND2_X1 g303 ( .A1(new_n437_), .A2(KEYINPUT12), .ZN(new_n440_) );
  INV_X1 g304 ( .A(new_n404_), .ZN(new_n441_) );
  NAND3_X1 g305 ( .A1(new_n253_), .A2(G257), .A3(new_n441_), .ZN(new_n442_) );
  NAND3_X1 g306 ( .A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n443_) );
  INV_X1 g307 ( .A(new_n443_), .ZN(new_n444_) );
  NAND2_X1 g308 ( .A1(new_n444_), .A2(new_n320_), .ZN(new_n445_) );
  NAND2_X1 g309 ( .A1(new_n443_), .A2(new_n331_), .ZN(new_n446_) );
  INV_X1 g310 ( .A(new_n186_), .ZN(new_n447_) );
  NAND2_X1 g311 ( .A1(new_n206_), .A2(new_n447_), .ZN(new_n448_) );
  NAND2_X1 g312 ( .A1(new_n223_), .A2(G107), .ZN(new_n449_) );
  NAND2_X1 g313 ( .A1(new_n227_), .A2(new_n140_), .ZN(new_n450_) );
  NAND3_X1 g314 ( .A1(new_n449_), .A2(KEYINPUT13), .A3(new_n450_), .ZN(new_n451_) );
  NAND2_X1 g315 ( .A1(new_n219_), .A2(G77), .ZN(new_n452_) );
  NAND2_X1 g316 ( .A1(new_n452_), .A2(new_n451_), .ZN(new_n453_) );
  INV_X1 g317 ( .A(KEYINPUT13), .ZN(new_n454_) );
  NAND2_X1 g318 ( .A1(new_n449_), .A2(new_n450_), .ZN(new_n455_) );
  NAND2_X1 g319 ( .A1(new_n455_), .A2(new_n454_), .ZN(new_n456_) );
  NOR2_X1 g320 ( .A1(new_n201_), .A2(new_n382_), .ZN(new_n457_) );
  NAND2_X1 g321 ( .A1(new_n457_), .A2(G97), .ZN(new_n458_) );
  NAND2_X1 g322 ( .A1(new_n456_), .A2(new_n458_), .ZN(new_n459_) );
  NOR2_X1 g323 ( .A1(new_n459_), .A2(new_n453_), .ZN(new_n460_) );
  NAND2_X1 g324 ( .A1(new_n460_), .A2(new_n448_), .ZN(new_n461_) );
  NAND3_X1 g325 ( .A1(new_n445_), .A2(new_n446_), .A3(new_n461_), .ZN(new_n462_) );
  NAND2_X1 g326 ( .A1(new_n444_), .A2(G190), .ZN(new_n463_) );
  NAND2_X1 g327 ( .A1(new_n443_), .A2(G200), .ZN(new_n464_) );
  NAND4_X1 g328 ( .A1(new_n463_), .A2(new_n464_), .A3(new_n448_), .A4(new_n460_), .ZN(new_n465_) );
  NAND2_X1 g329 ( .A1(new_n465_), .A2(new_n462_), .ZN(new_n466_) );
  INV_X1 g330 ( .A(new_n466_), .ZN(new_n467_) );
  INV_X1 g331 ( .A(KEYINPUT11), .ZN(new_n468_) );
  INV_X1 g332 ( .A(new_n457_), .ZN(new_n469_) );
  NAND2_X1 g333 ( .A1(new_n205_), .A2(new_n469_), .ZN(new_n470_) );
  NAND2_X1 g334 ( .A1(new_n470_), .A2(G116), .ZN(new_n471_) );
  NAND2_X1 g335 ( .A1(new_n219_), .A2(G97), .ZN(new_n472_) );
  NAND2_X1 g336 ( .A1(new_n223_), .A2(G283), .ZN(new_n473_) );
  INV_X1 g337 ( .A(G116), .ZN(new_n474_) );
  NAND2_X1 g338 ( .A1(new_n227_), .A2(new_n474_), .ZN(new_n475_) );
  NAND3_X1 g339 ( .A1(new_n472_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_) );
  INV_X1 g340 ( .A(new_n476_), .ZN(new_n477_) );
  NAND2_X1 g341 ( .A1(new_n471_), .A2(new_n477_), .ZN(new_n478_) );
  NAND4_X1 g342 ( .A1(new_n166_), .A2(new_n215_), .A3(G257), .A4(new_n241_), .ZN(new_n479_) );
  NAND3_X1 g343 ( .A1(new_n166_), .A2(G303), .A3(new_n257_), .ZN(new_n480_) );
  NAND3_X1 g344 ( .A1(new_n479_), .A2(new_n405_), .A3(new_n480_), .ZN(new_n481_) );
  INV_X1 g345 ( .A(new_n481_), .ZN(new_n482_) );
  NAND4_X1 g346 ( .A1(new_n253_), .A2(G270), .A3(KEYINPUT10), .A4(new_n441_), .ZN(new_n483_) );
  NAND3_X1 g347 ( .A1(new_n217_), .A2(G264), .A3(G1698), .ZN(new_n484_) );
  INV_X1 g348 ( .A(KEYINPUT10), .ZN(new_n485_) );
  NAND3_X1 g349 ( .A1(new_n253_), .A2(G270), .A3(new_n441_), .ZN(new_n486_) );
  NAND2_X1 g350 ( .A1(new_n486_), .A2(new_n485_), .ZN(new_n487_) );
  NAND4_X1 g351 ( .A1(new_n482_), .A2(new_n487_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n488_) );
  NAND2_X1 g352 ( .A1(new_n488_), .A2(G169), .ZN(new_n489_) );
  NAND2_X1 g353 ( .A1(new_n487_), .A2(new_n484_), .ZN(new_n490_) );
  INV_X1 g354 ( .A(new_n490_), .ZN(new_n491_) );
  NAND4_X1 g355 ( .A1(new_n491_), .A2(G179), .A3(new_n482_), .A4(new_n483_), .ZN(new_n492_) );
  NAND2_X1 g356 ( .A1(new_n492_), .A2(new_n489_), .ZN(new_n493_) );
  NAND2_X1 g357 ( .A1(new_n478_), .A2(new_n493_), .ZN(new_n494_) );
  NAND2_X1 g358 ( .A1(new_n488_), .A2(G200), .ZN(new_n495_) );
  NAND4_X1 g359 ( .A1(new_n491_), .A2(G190), .A3(new_n482_), .A4(new_n483_), .ZN(new_n496_) );
  NAND4_X1 g360 ( .A1(new_n471_), .A2(new_n477_), .A3(new_n496_), .A4(new_n495_), .ZN(new_n497_) );
  NAND2_X1 g361 ( .A1(new_n494_), .A2(new_n497_), .ZN(new_n498_) );
  XNOR2_X1 g362 ( .A(new_n498_), .B(new_n468_), .ZN(new_n499_) );
  INV_X1 g363 ( .A(KEYINPUT9), .ZN(new_n500_) );
  NAND2_X1 g364 ( .A1(new_n457_), .A2(G87), .ZN(new_n501_) );
  NAND2_X1 g365 ( .A1(new_n205_), .A2(new_n501_), .ZN(new_n502_) );
  INV_X1 g366 ( .A(G87), .ZN(new_n503_) );
  NAND3_X1 g367 ( .A1(new_n503_), .A2(new_n140_), .A3(new_n141_), .ZN(new_n504_) );
  NAND3_X1 g368 ( .A1(new_n502_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_) );
  NAND2_X1 g369 ( .A1(new_n502_), .A2(new_n504_), .ZN(new_n506_) );
  NAND2_X1 g370 ( .A1(new_n506_), .A2(KEYINPUT9), .ZN(new_n507_) );
  NAND2_X1 g371 ( .A1(new_n219_), .A2(G68), .ZN(new_n508_) );
  NAND2_X1 g372 ( .A1(new_n223_), .A2(G97), .ZN(new_n509_) );
  NAND2_X1 g373 ( .A1(new_n227_), .A2(new_n503_), .ZN(new_n510_) );
  NAND3_X1 g374 ( .A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_) );
  INV_X1 g375 ( .A(new_n511_), .ZN(new_n512_) );
  NAND3_X1 g376 ( .A1(new_n507_), .A2(new_n505_), .A3(new_n512_), .ZN(new_n513_) );
  INV_X1 g377 ( .A(new_n513_), .ZN(new_n514_) );
  NAND3_X1 g378 ( .A1(new_n217_), .A2(G244), .A3(G1698), .ZN(new_n515_) );
  NAND4_X1 g379 ( .A1(new_n166_), .A2(new_n215_), .A3(G238), .A4(new_n241_), .ZN(new_n516_) );
  NAND2_X1 g380 ( .A1(new_n515_), .A2(new_n516_), .ZN(new_n517_) );
  NAND2_X1 g381 ( .A1(new_n517_), .A2(KEYINPUT8), .ZN(new_n518_) );
  INV_X1 g382 ( .A(KEYINPUT8), .ZN(new_n519_) );
  NAND3_X1 g383 ( .A1(new_n515_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_) );
  NAND2_X1 g384 ( .A1(new_n209_), .A2(G45), .ZN(new_n521_) );
  NAND3_X1 g385 ( .A1(new_n253_), .A2(G250), .A3(new_n521_), .ZN(new_n522_) );
  INV_X1 g386 ( .A(new_n522_), .ZN(new_n523_) );
  NAND2_X1 g387 ( .A1(new_n259_), .A2(G116), .ZN(new_n524_) );
  NAND3_X1 g388 ( .A1(new_n209_), .A2(G45), .A3(G274), .ZN(new_n525_) );
  NAND2_X1 g389 ( .A1(new_n524_), .A2(new_n525_), .ZN(new_n526_) );
  NOR2_X1 g390 ( .A1(new_n526_), .A2(new_n523_), .ZN(new_n527_) );
  NAND3_X1 g391 ( .A1(new_n518_), .A2(new_n527_), .A3(new_n520_), .ZN(new_n528_) );
  NAND2_X1 g392 ( .A1(new_n528_), .A2(G200), .ZN(new_n529_) );
  INV_X1 g393 ( .A(new_n528_), .ZN(new_n530_) );
  NAND2_X1 g394 ( .A1(new_n530_), .A2(G190), .ZN(new_n531_) );
  NAND3_X1 g395 ( .A1(new_n514_), .A2(new_n529_), .A3(new_n531_), .ZN(new_n532_) );
  NAND2_X1 g396 ( .A1(new_n528_), .A2(G169), .ZN(new_n533_) );
  NAND2_X1 g397 ( .A1(new_n530_), .A2(G179), .ZN(new_n534_) );
  NAND2_X1 g398 ( .A1(new_n534_), .A2(new_n533_), .ZN(new_n535_) );
  NAND2_X1 g399 ( .A1(new_n535_), .A2(new_n513_), .ZN(new_n536_) );
  NAND2_X1 g400 ( .A1(new_n532_), .A2(new_n536_), .ZN(new_n537_) );
  NOR2_X1 g401 ( .A1(new_n499_), .A2(new_n537_), .ZN(new_n538_) );
  NAND2_X1 g402 ( .A1(new_n538_), .A2(new_n467_), .ZN(new_n539_) );
  NOR3_X1 g403 ( .A1(new_n378_), .A2(new_n433_), .A3(new_n539_), .ZN(G372) );
  INV_X1 g404 ( .A(new_n494_), .ZN(new_n541_) );
  NAND2_X1 g405 ( .A1(new_n432_), .A2(new_n541_), .ZN(new_n542_) );
  NAND2_X1 g406 ( .A1(new_n542_), .A2(new_n422_), .ZN(new_n543_) );
  NAND2_X1 g407 ( .A1(new_n543_), .A2(new_n467_), .ZN(new_n544_) );
  NAND3_X1 g408 ( .A1(new_n544_), .A2(new_n462_), .A3(new_n536_), .ZN(new_n545_) );
  NAND2_X1 g409 ( .A1(new_n545_), .A2(new_n532_), .ZN(new_n546_) );
  INV_X1 g410 ( .A(new_n546_), .ZN(new_n547_) );
  NAND2_X1 g411 ( .A1(new_n547_), .A2(new_n377_), .ZN(new_n548_) );
  NAND4_X1 g412 ( .A1(new_n367_), .A2(new_n295_), .A3(new_n304_), .A4(new_n373_), .ZN(new_n549_) );
  NAND2_X1 g413 ( .A1(new_n549_), .A2(new_n373_), .ZN(new_n550_) );
  NAND2_X1 g414 ( .A1(new_n550_), .A2(new_n278_), .ZN(new_n551_) );
  NAND2_X1 g415 ( .A1(new_n551_), .A2(new_n271_), .ZN(new_n552_) );
  NAND2_X1 g416 ( .A1(new_n552_), .A2(new_n345_), .ZN(new_n553_) );
  NAND2_X1 g417 ( .A1(new_n553_), .A2(new_n338_), .ZN(new_n554_) );
  INV_X1 g418 ( .A(new_n554_), .ZN(new_n555_) );
  NAND2_X1 g419 ( .A1(new_n548_), .A2(new_n555_), .ZN(G369) );
  INV_X1 g420 ( .A(new_n499_), .ZN(new_n557_) );
  INV_X1 g421 ( .A(G343), .ZN(new_n558_) );
  NAND4_X1 g422 ( .A1(new_n209_), .A2(new_n214_), .A3(G13), .A4(G213), .ZN(new_n559_) );
  NOR2_X1 g423 ( .A1(new_n559_), .A2(new_n558_), .ZN(new_n560_) );
  NAND2_X1 g424 ( .A1(new_n478_), .A2(new_n560_), .ZN(new_n561_) );
  NAND2_X1 g425 ( .A1(new_n557_), .A2(new_n561_), .ZN(new_n562_) );
  NAND2_X1 g426 ( .A1(new_n541_), .A2(new_n560_), .ZN(new_n563_) );
  NAND2_X1 g427 ( .A1(new_n562_), .A2(new_n563_), .ZN(new_n564_) );
  NAND2_X1 g428 ( .A1(new_n395_), .A2(new_n560_), .ZN(new_n565_) );
  NAND2_X1 g429 ( .A1(new_n432_), .A2(new_n565_), .ZN(new_n566_) );
  NAND4_X1 g430 ( .A1(new_n421_), .A2(new_n395_), .A3(new_n414_), .A4(new_n560_), .ZN(new_n567_) );
  NAND2_X1 g431 ( .A1(new_n566_), .A2(new_n567_), .ZN(new_n568_) );
  NAND3_X1 g432 ( .A1(new_n564_), .A2(new_n568_), .A3(G330), .ZN(new_n569_) );
  INV_X1 g433 ( .A(new_n560_), .ZN(new_n570_) );
  NAND2_X1 g434 ( .A1(new_n543_), .A2(new_n570_), .ZN(new_n571_) );
  NAND2_X1 g435 ( .A1(new_n569_), .A2(new_n571_), .ZN(G399) );
  NAND2_X1 g436 ( .A1(new_n547_), .A2(new_n570_), .ZN(new_n573_) );
  NAND4_X1 g437 ( .A1(new_n538_), .A2(new_n432_), .A3(new_n467_), .A4(new_n570_), .ZN(new_n574_) );
  INV_X1 g438 ( .A(KEYINPUT18), .ZN(new_n575_) );
  NAND3_X1 g439 ( .A1(new_n444_), .A2(new_n575_), .A3(new_n530_), .ZN(new_n576_) );
  NAND2_X1 g440 ( .A1(new_n444_), .A2(new_n530_), .ZN(new_n577_) );
  NAND2_X1 g441 ( .A1(new_n577_), .A2(KEYINPUT18), .ZN(new_n578_) );
  NOR2_X1 g442 ( .A1(new_n492_), .A2(new_n412_), .ZN(new_n579_) );
  NAND3_X1 g443 ( .A1(new_n578_), .A2(new_n576_), .A3(new_n579_), .ZN(new_n580_) );
  NOR2_X1 g444 ( .A1(new_n413_), .A2(G179), .ZN(new_n581_) );
  NAND4_X1 g445 ( .A1(new_n443_), .A2(new_n488_), .A3(new_n528_), .A4(new_n581_), .ZN(new_n582_) );
  NAND2_X1 g446 ( .A1(new_n580_), .A2(new_n582_), .ZN(new_n583_) );
  NAND2_X1 g447 ( .A1(new_n583_), .A2(new_n560_), .ZN(new_n584_) );
  NAND2_X1 g448 ( .A1(new_n574_), .A2(new_n584_), .ZN(new_n585_) );
  NAND2_X1 g449 ( .A1(new_n585_), .A2(G330), .ZN(new_n586_) );
  NAND2_X1 g450 ( .A1(new_n573_), .A2(new_n586_), .ZN(new_n587_) );
  NAND2_X1 g451 ( .A1(new_n587_), .A2(new_n209_), .ZN(new_n588_) );
  NOR2_X1 g452 ( .A1(new_n504_), .A2(G116), .ZN(new_n589_) );
  INV_X1 g453 ( .A(new_n172_), .ZN(new_n590_) );
  NOR2_X1 g454 ( .A1(new_n590_), .A2(G41), .ZN(new_n591_) );
  INV_X1 g455 ( .A(new_n591_), .ZN(new_n592_) );
  NAND3_X1 g456 ( .A1(new_n592_), .A2(G1), .A3(new_n589_), .ZN(new_n593_) );
  NAND2_X1 g457 ( .A1(new_n591_), .A2(new_n170_), .ZN(new_n594_) );
  NAND3_X1 g458 ( .A1(new_n588_), .A2(new_n593_), .A3(new_n594_), .ZN(G364) );
  INV_X1 g459 ( .A(new_n564_), .ZN(new_n596_) );
  NOR2_X1 g460 ( .A1(G13), .A2(G33), .ZN(new_n597_) );
  INV_X1 g461 ( .A(new_n597_), .ZN(new_n598_) );
  NOR2_X1 g462 ( .A1(new_n598_), .A2(G20), .ZN(new_n599_) );
  NAND3_X1 g463 ( .A1(new_n596_), .A2(KEYINPUT62), .A3(new_n599_), .ZN(new_n600_) );
  INV_X1 g464 ( .A(KEYINPUT62), .ZN(new_n601_) );
  NAND2_X1 g465 ( .A1(new_n596_), .A2(new_n599_), .ZN(new_n602_) );
  NAND2_X1 g466 ( .A1(new_n602_), .A2(new_n601_), .ZN(new_n603_) );
  NAND2_X1 g467 ( .A1(new_n172_), .A2(G33), .ZN(new_n604_) );
  XOR2_X1 g468 ( .A(new_n604_), .B(KEYINPUT24), .Z(new_n605_) );
  NAND2_X1 g469 ( .A1(new_n192_), .A2(G45), .ZN(new_n606_) );
  NAND2_X1 g470 ( .A1(new_n170_), .A2(new_n248_), .ZN(new_n607_) );
  NAND3_X1 g471 ( .A1(new_n606_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_) );
  NAND3_X1 g472 ( .A1(new_n590_), .A2(new_n474_), .A3(KEYINPUT60), .ZN(new_n609_) );
  NAND2_X1 g473 ( .A1(G355), .A2(new_n597_), .ZN(new_n610_) );
  INV_X1 g474 ( .A(KEYINPUT60), .ZN(new_n611_) );
  NAND2_X1 g475 ( .A1(new_n590_), .A2(new_n474_), .ZN(new_n612_) );
  NAND2_X1 g476 ( .A1(new_n612_), .A2(new_n611_), .ZN(new_n613_) );
  NAND4_X1 g477 ( .A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .A4(new_n613_), .ZN(new_n614_) );
  INV_X1 g478 ( .A(new_n599_), .ZN(new_n615_) );
  NAND2_X1 g479 ( .A1(new_n331_), .A2(G20), .ZN(new_n616_) );
  NAND2_X1 g480 ( .A1(new_n166_), .A2(new_n616_), .ZN(new_n617_) );
  NAND2_X1 g481 ( .A1(new_n615_), .A2(new_n617_), .ZN(new_n618_) );
  INV_X1 g482 ( .A(new_n618_), .ZN(new_n619_) );
  NAND2_X1 g483 ( .A1(new_n614_), .A2(new_n619_), .ZN(new_n620_) );
  INV_X1 g484 ( .A(new_n620_), .ZN(new_n621_) );
  NAND3_X1 g485 ( .A1(new_n320_), .A2(new_n364_), .A3(G190), .ZN(new_n622_) );
  NAND2_X1 g486 ( .A1(new_n622_), .A2(G20), .ZN(new_n623_) );
  INV_X1 g487 ( .A(new_n623_), .ZN(new_n624_) );
  NOR2_X1 g488 ( .A1(new_n624_), .A2(new_n140_), .ZN(new_n625_) );
  NAND2_X1 g489 ( .A1(G20), .A2(G179), .ZN(new_n626_) );
  NOR3_X1 g490 ( .A1(new_n626_), .A2(G190), .A3(G200), .ZN(new_n627_) );
  INV_X1 g491 ( .A(new_n627_), .ZN(new_n628_) );
  NOR2_X1 g492 ( .A1(new_n628_), .A2(new_n300_), .ZN(new_n629_) );
  INV_X1 g493 ( .A(G159), .ZN(new_n630_) );
  INV_X1 g494 ( .A(G190), .ZN(new_n631_) );
  NOR2_X1 g495 ( .A1(new_n214_), .A2(G179), .ZN(new_n632_) );
  NAND3_X1 g496 ( .A1(new_n632_), .A2(new_n631_), .A3(new_n364_), .ZN(new_n633_) );
  NOR2_X1 g497 ( .A1(new_n633_), .A2(new_n630_), .ZN(new_n634_) );
  NOR3_X1 g498 ( .A1(new_n626_), .A2(new_n364_), .A3(G190), .ZN(new_n635_) );
  INV_X1 g499 ( .A(new_n635_), .ZN(new_n636_) );
  NOR2_X1 g500 ( .A1(new_n636_), .A2(new_n346_), .ZN(new_n637_) );
  NOR4_X1 g501 ( .A1(new_n625_), .A2(new_n629_), .A3(new_n637_), .A4(new_n634_), .ZN(new_n638_) );
  NAND2_X1 g502 ( .A1(new_n638_), .A2(KEYINPUT61), .ZN(new_n639_) );
  INV_X1 g503 ( .A(KEYINPUT61), .ZN(new_n640_) );
  INV_X1 g504 ( .A(new_n638_), .ZN(new_n641_) );
  NAND2_X1 g505 ( .A1(new_n641_), .A2(new_n640_), .ZN(new_n642_) );
  INV_X1 g506 ( .A(new_n617_), .ZN(new_n643_) );
  NAND2_X1 g507 ( .A1(new_n643_), .A2(new_n215_), .ZN(new_n644_) );
  NAND3_X1 g508 ( .A1(new_n632_), .A2(new_n631_), .A3(G200), .ZN(new_n645_) );
  NOR2_X1 g509 ( .A1(new_n645_), .A2(new_n141_), .ZN(new_n646_) );
  NAND2_X1 g510 ( .A1(G190), .A2(G200), .ZN(new_n647_) );
  NOR2_X1 g511 ( .A1(new_n626_), .A2(new_n647_), .ZN(new_n648_) );
  NAND2_X1 g512 ( .A1(new_n648_), .A2(G50), .ZN(new_n649_) );
  NOR3_X1 g513 ( .A1(new_n626_), .A2(new_n631_), .A3(G200), .ZN(new_n650_) );
  NAND2_X1 g514 ( .A1(new_n650_), .A2(G58), .ZN(new_n651_) );
  NOR3_X1 g515 ( .A1(new_n647_), .A2(new_n214_), .A3(G179), .ZN(new_n652_) );
  NAND2_X1 g516 ( .A1(new_n652_), .A2(G87), .ZN(new_n653_) );
  NAND3_X1 g517 ( .A1(new_n651_), .A2(new_n653_), .A3(new_n649_), .ZN(new_n654_) );
  NOR3_X1 g518 ( .A1(new_n644_), .A2(new_n646_), .A3(new_n654_), .ZN(new_n655_) );
  NAND3_X1 g519 ( .A1(new_n642_), .A2(new_n639_), .A3(new_n655_), .ZN(new_n656_) );
  INV_X1 g520 ( .A(new_n645_), .ZN(new_n657_) );
  NAND2_X1 g521 ( .A1(new_n657_), .A2(G283), .ZN(new_n658_) );
  INV_X1 g522 ( .A(new_n633_), .ZN(new_n659_) );
  NAND2_X1 g523 ( .A1(new_n659_), .A2(G329), .ZN(new_n660_) );
  NAND2_X1 g524 ( .A1(new_n627_), .A2(G311), .ZN(new_n661_) );
  NAND2_X1 g525 ( .A1(new_n643_), .A2(G33), .ZN(new_n662_) );
  INV_X1 g526 ( .A(G322), .ZN(new_n663_) );
  INV_X1 g527 ( .A(new_n650_), .ZN(new_n664_) );
  NOR2_X1 g528 ( .A1(new_n664_), .A2(new_n663_), .ZN(new_n665_) );
  NAND2_X1 g529 ( .A1(new_n652_), .A2(G303), .ZN(new_n666_) );
  NAND2_X1 g530 ( .A1(new_n648_), .A2(G326), .ZN(new_n667_) );
  NAND2_X1 g531 ( .A1(new_n666_), .A2(new_n667_), .ZN(new_n668_) );
  NAND2_X1 g532 ( .A1(new_n623_), .A2(G294), .ZN(new_n669_) );
  NAND2_X1 g533 ( .A1(new_n635_), .A2(G317), .ZN(new_n670_) );
  NAND2_X1 g534 ( .A1(new_n669_), .A2(new_n670_), .ZN(new_n671_) );
  NOR4_X1 g535 ( .A1(new_n662_), .A2(new_n671_), .A3(new_n665_), .A4(new_n668_), .ZN(new_n672_) );
  NAND4_X1 g536 ( .A1(new_n672_), .A2(new_n658_), .A3(new_n660_), .A4(new_n661_), .ZN(new_n673_) );
  NAND3_X1 g537 ( .A1(new_n214_), .A2(G13), .A3(G45), .ZN(new_n674_) );
  NAND2_X1 g538 ( .A1(new_n674_), .A2(G1), .ZN(new_n675_) );
  XOR2_X1 g539 ( .A(new_n675_), .B(KEYINPUT1), .Z(new_n676_) );
  INV_X1 g540 ( .A(new_n676_), .ZN(new_n677_) );
  NAND2_X1 g541 ( .A1(new_n677_), .A2(new_n592_), .ZN(new_n678_) );
  INV_X1 g542 ( .A(new_n678_), .ZN(new_n679_) );
  NAND3_X1 g543 ( .A1(new_n656_), .A2(new_n673_), .A3(new_n679_), .ZN(new_n680_) );
  NOR2_X1 g544 ( .A1(new_n680_), .A2(new_n621_), .ZN(new_n681_) );
  NAND3_X1 g545 ( .A1(new_n603_), .A2(new_n600_), .A3(new_n681_), .ZN(new_n682_) );
  NAND2_X1 g546 ( .A1(new_n564_), .A2(G330), .ZN(new_n683_) );
  INV_X1 g547 ( .A(G330), .ZN(new_n684_) );
  NAND2_X1 g548 ( .A1(new_n596_), .A2(new_n684_), .ZN(new_n685_) );
  NAND3_X1 g549 ( .A1(new_n685_), .A2(new_n683_), .A3(new_n678_), .ZN(new_n686_) );
  NAND2_X1 g550 ( .A1(new_n682_), .A2(new_n686_), .ZN(G396) );
  INV_X1 g551 ( .A(new_n587_), .ZN(new_n688_) );
  NAND2_X1 g552 ( .A1(new_n304_), .A2(new_n560_), .ZN(new_n689_) );
  XOR2_X1 g553 ( .A(new_n689_), .B(KEYINPUT5), .Z(new_n690_) );
  NAND2_X1 g554 ( .A1(new_n310_), .A2(new_n690_), .ZN(new_n691_) );
  INV_X1 g555 ( .A(new_n690_), .ZN(new_n692_) );
  NAND2_X1 g556 ( .A1(new_n692_), .A2(new_n295_), .ZN(new_n693_) );
  NAND2_X1 g557 ( .A1(new_n691_), .A2(new_n693_), .ZN(new_n694_) );
  INV_X1 g558 ( .A(new_n694_), .ZN(new_n695_) );
  NAND2_X1 g559 ( .A1(new_n688_), .A2(new_n695_), .ZN(new_n696_) );
  NAND2_X1 g560 ( .A1(new_n587_), .A2(new_n694_), .ZN(new_n697_) );
  NAND3_X1 g561 ( .A1(new_n696_), .A2(new_n678_), .A3(new_n697_), .ZN(new_n698_) );
  NAND2_X1 g562 ( .A1(new_n695_), .A2(new_n597_), .ZN(new_n699_) );
  NAND2_X1 g563 ( .A1(new_n635_), .A2(G150), .ZN(new_n700_) );
  NAND2_X1 g564 ( .A1(new_n657_), .A2(G68), .ZN(new_n701_) );
  NAND2_X1 g565 ( .A1(new_n650_), .A2(G143), .ZN(new_n702_) );
  NAND3_X1 g566 ( .A1(new_n701_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_) );
  INV_X1 g567 ( .A(new_n703_), .ZN(new_n704_) );
  NAND2_X1 g568 ( .A1(new_n659_), .A2(G132), .ZN(new_n705_) );
  NAND2_X1 g569 ( .A1(new_n705_), .A2(KEYINPUT19), .ZN(new_n706_) );
  NOR2_X1 g570 ( .A1(new_n705_), .A2(KEYINPUT19), .ZN(new_n707_) );
  NOR2_X1 g571 ( .A1(new_n707_), .A2(new_n644_), .ZN(new_n708_) );
  NAND2_X1 g572 ( .A1(new_n627_), .A2(G159), .ZN(new_n709_) );
  NAND2_X1 g573 ( .A1(new_n623_), .A2(G58), .ZN(new_n710_) );
  NAND2_X1 g574 ( .A1(new_n652_), .A2(G50), .ZN(new_n711_) );
  NAND2_X1 g575 ( .A1(new_n648_), .A2(G137), .ZN(new_n712_) );
  NAND4_X1 g576 ( .A1(new_n710_), .A2(new_n709_), .A3(new_n711_), .A4(new_n712_), .ZN(new_n713_) );
  XOR2_X1 g577 ( .A(new_n713_), .B(KEYINPUT20), .Z(new_n714_) );
  NAND4_X1 g578 ( .A1(new_n714_), .A2(new_n704_), .A3(new_n706_), .A4(new_n708_), .ZN(new_n715_) );
  NAND2_X1 g579 ( .A1(new_n627_), .A2(G116), .ZN(new_n716_) );
  NAND2_X1 g580 ( .A1(new_n716_), .A2(KEYINPUT21), .ZN(new_n717_) );
  NOR2_X1 g581 ( .A1(new_n716_), .A2(KEYINPUT21), .ZN(new_n718_) );
  NAND2_X1 g582 ( .A1(new_n650_), .A2(G294), .ZN(new_n719_) );
  NAND2_X1 g583 ( .A1(new_n652_), .A2(G107), .ZN(new_n720_) );
  NAND2_X1 g584 ( .A1(new_n648_), .A2(G303), .ZN(new_n721_) );
  NAND4_X1 g585 ( .A1(new_n719_), .A2(new_n720_), .A3(G33), .A4(new_n721_), .ZN(new_n722_) );
  NOR2_X1 g586 ( .A1(new_n722_), .A2(new_n718_), .ZN(new_n723_) );
  NAND2_X1 g587 ( .A1(new_n657_), .A2(G87), .ZN(new_n724_) );
  XNOR2_X1 g588 ( .A(new_n724_), .B(KEYINPUT22), .ZN(new_n725_) );
  INV_X1 g589 ( .A(G311), .ZN(new_n726_) );
  NOR2_X1 g590 ( .A1(new_n633_), .A2(new_n726_), .ZN(new_n727_) );
  INV_X1 g591 ( .A(G283), .ZN(new_n728_) );
  NOR2_X1 g592 ( .A1(new_n636_), .A2(new_n728_), .ZN(new_n729_) );
  NOR4_X1 g593 ( .A1(new_n625_), .A2(new_n729_), .A3(new_n727_), .A4(new_n617_), .ZN(new_n730_) );
  NAND4_X1 g594 ( .A1(new_n725_), .A2(new_n730_), .A3(new_n717_), .A4(new_n723_), .ZN(new_n731_) );
  NAND2_X1 g595 ( .A1(new_n617_), .A2(new_n598_), .ZN(new_n732_) );
  INV_X1 g596 ( .A(new_n732_), .ZN(new_n733_) );
  NAND2_X1 g597 ( .A1(new_n733_), .A2(new_n300_), .ZN(new_n734_) );
  NAND2_X1 g598 ( .A1(new_n679_), .A2(new_n734_), .ZN(new_n735_) );
  INV_X1 g599 ( .A(new_n735_), .ZN(new_n736_) );
  NAND4_X1 g600 ( .A1(new_n699_), .A2(new_n715_), .A3(new_n731_), .A4(new_n736_), .ZN(new_n737_) );
  NAND2_X1 g601 ( .A1(new_n698_), .A2(new_n737_), .ZN(G384) );
  NAND2_X1 g602 ( .A1(new_n272_), .A2(new_n559_), .ZN(new_n739_) );
  NAND3_X1 g603 ( .A1(new_n545_), .A2(new_n308_), .A3(new_n532_), .ZN(new_n740_) );
  NAND2_X1 g604 ( .A1(new_n740_), .A2(new_n305_), .ZN(new_n741_) );
  INV_X1 g605 ( .A(KEYINPUT29), .ZN(new_n742_) );
  NAND2_X1 g606 ( .A1(new_n369_), .A2(new_n560_), .ZN(new_n743_) );
  NAND3_X1 g607 ( .A1(new_n367_), .A2(new_n373_), .A3(new_n743_), .ZN(new_n744_) );
  NAND2_X1 g608 ( .A1(new_n374_), .A2(new_n560_), .ZN(new_n745_) );
  NAND2_X1 g609 ( .A1(new_n744_), .A2(new_n745_), .ZN(new_n746_) );
  XNOR2_X1 g610 ( .A(new_n746_), .B(new_n742_), .ZN(new_n747_) );
  NAND3_X1 g611 ( .A1(new_n741_), .A2(new_n570_), .A3(new_n747_), .ZN(new_n748_) );
  NAND2_X1 g612 ( .A1(new_n374_), .A2(new_n570_), .ZN(new_n749_) );
  NAND2_X1 g613 ( .A1(new_n748_), .A2(new_n749_), .ZN(new_n750_) );
  INV_X1 g614 ( .A(new_n559_), .ZN(new_n751_) );
  NAND2_X1 g615 ( .A1(new_n233_), .A2(new_n751_), .ZN(new_n752_) );
  NAND2_X1 g616 ( .A1(new_n278_), .A2(new_n752_), .ZN(new_n753_) );
  NAND2_X1 g617 ( .A1(new_n271_), .A2(new_n753_), .ZN(new_n754_) );
  NAND3_X1 g618 ( .A1(new_n750_), .A2(new_n739_), .A3(new_n754_), .ZN(new_n755_) );
  NAND2_X1 g619 ( .A1(new_n755_), .A2(new_n739_), .ZN(new_n756_) );
  NAND4_X1 g620 ( .A1(new_n377_), .A2(new_n545_), .A3(new_n532_), .A4(new_n570_), .ZN(new_n757_) );
  NAND2_X1 g621 ( .A1(new_n555_), .A2(new_n757_), .ZN(new_n758_) );
  XNOR2_X1 g622 ( .A(new_n756_), .B(new_n758_), .ZN(new_n759_) );
  INV_X1 g623 ( .A(new_n747_), .ZN(new_n760_) );
  NAND2_X1 g624 ( .A1(new_n739_), .A2(new_n754_), .ZN(new_n761_) );
  NOR4_X1 g625 ( .A1(new_n378_), .A2(new_n761_), .A3(new_n760_), .A4(new_n695_), .ZN(new_n762_) );
  NOR3_X1 g626 ( .A1(new_n761_), .A2(new_n760_), .A3(new_n695_), .ZN(new_n763_) );
  NOR2_X1 g627 ( .A1(new_n763_), .A2(new_n377_), .ZN(new_n764_) );
  NOR3_X1 g628 ( .A1(new_n764_), .A2(new_n762_), .A3(new_n586_), .ZN(new_n765_) );
  XNOR2_X1 g629 ( .A(new_n759_), .B(new_n765_), .ZN(new_n766_) );
  NAND2_X1 g630 ( .A1(new_n766_), .A2(new_n167_), .ZN(new_n767_) );
  INV_X1 g631 ( .A(G13), .ZN(new_n768_) );
  NAND2_X1 g632 ( .A1(new_n768_), .A2(G1), .ZN(new_n769_) );
  NAND2_X1 g633 ( .A1(new_n767_), .A2(new_n769_), .ZN(new_n770_) );
  NAND2_X1 g634 ( .A1(G50), .A2(G58), .ZN(new_n771_) );
  XNOR2_X1 g635 ( .A(new_n771_), .B(G68), .ZN(new_n772_) );
  NAND2_X1 g636 ( .A1(new_n300_), .A2(G50), .ZN(new_n773_) );
  NAND2_X1 g637 ( .A1(new_n772_), .A2(new_n773_), .ZN(new_n774_) );
  NAND3_X1 g638 ( .A1(new_n774_), .A2(G1), .A3(new_n768_), .ZN(new_n775_) );
  NAND2_X1 g639 ( .A1(new_n770_), .A2(new_n775_), .ZN(new_n776_) );
  NAND3_X1 g640 ( .A1(new_n168_), .A2(G116), .A3(new_n186_), .ZN(new_n777_) );
  NAND2_X1 g641 ( .A1(new_n776_), .A2(new_n777_), .ZN(G367) );
  INV_X1 g642 ( .A(KEYINPUT55), .ZN(new_n779_) );
  INV_X1 g643 ( .A(KEYINPUT52), .ZN(new_n780_) );
  NAND2_X1 g644 ( .A1(new_n461_), .A2(new_n560_), .ZN(new_n781_) );
  NAND2_X1 g645 ( .A1(new_n571_), .A2(new_n781_), .ZN(new_n782_) );
  XNOR2_X1 g646 ( .A(new_n782_), .B(new_n467_), .ZN(new_n783_) );
  NAND2_X1 g647 ( .A1(new_n783_), .A2(new_n569_), .ZN(new_n784_) );
  INV_X1 g648 ( .A(new_n569_), .ZN(new_n785_) );
  XNOR2_X1 g649 ( .A(new_n782_), .B(new_n466_), .ZN(new_n786_) );
  NAND2_X1 g650 ( .A1(new_n786_), .A2(new_n785_), .ZN(new_n787_) );
  NAND2_X1 g651 ( .A1(new_n541_), .A2(new_n570_), .ZN(new_n788_) );
  NAND2_X1 g652 ( .A1(new_n788_), .A2(new_n565_), .ZN(new_n789_) );
  XOR2_X1 g653 ( .A(new_n432_), .B(new_n789_), .Z(new_n790_) );
  XNOR2_X1 g654 ( .A(new_n683_), .B(new_n790_), .ZN(new_n791_) );
  NAND3_X1 g655 ( .A1(new_n784_), .A2(new_n787_), .A3(new_n791_), .ZN(new_n792_) );
  NAND2_X1 g656 ( .A1(new_n792_), .A2(new_n780_), .ZN(new_n793_) );
  XNOR2_X1 g657 ( .A(new_n786_), .B(new_n569_), .ZN(new_n794_) );
  NAND3_X1 g658 ( .A1(new_n794_), .A2(KEYINPUT52), .A3(new_n791_), .ZN(new_n795_) );
  NAND3_X1 g659 ( .A1(new_n573_), .A2(new_n586_), .A3(new_n677_), .ZN(new_n796_) );
  INV_X1 g660 ( .A(new_n796_), .ZN(new_n797_) );
  NAND3_X1 g661 ( .A1(new_n795_), .A2(new_n793_), .A3(new_n797_), .ZN(new_n798_) );
  INV_X1 g662 ( .A(KEYINPUT53), .ZN(new_n799_) );
  INV_X1 g663 ( .A(new_n537_), .ZN(new_n800_) );
  NAND2_X1 g664 ( .A1(new_n544_), .A2(new_n462_), .ZN(new_n801_) );
  NAND2_X1 g665 ( .A1(new_n801_), .A2(new_n800_), .ZN(new_n802_) );
  NAND3_X1 g666 ( .A1(new_n544_), .A2(new_n462_), .A3(new_n537_), .ZN(new_n803_) );
  NAND3_X1 g667 ( .A1(new_n802_), .A2(new_n570_), .A3(new_n803_), .ZN(new_n804_) );
  NAND2_X1 g668 ( .A1(new_n532_), .A2(new_n560_), .ZN(new_n805_) );
  NAND3_X1 g669 ( .A1(new_n804_), .A2(new_n799_), .A3(new_n805_), .ZN(new_n806_) );
  NAND2_X1 g670 ( .A1(new_n804_), .A2(new_n805_), .ZN(new_n807_) );
  NAND2_X1 g671 ( .A1(new_n807_), .A2(KEYINPUT53), .ZN(new_n808_) );
  NAND4_X1 g672 ( .A1(new_n513_), .A2(new_n533_), .A3(new_n534_), .A4(new_n560_), .ZN(new_n809_) );
  NAND3_X1 g673 ( .A1(new_n808_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_) );
  NAND2_X1 g674 ( .A1(new_n467_), .A2(new_n781_), .ZN(new_n811_) );
  NAND4_X1 g675 ( .A1(new_n445_), .A2(new_n446_), .A3(new_n461_), .A4(new_n560_), .ZN(new_n812_) );
  NAND2_X1 g676 ( .A1(new_n811_), .A2(new_n812_), .ZN(new_n813_) );
  NAND2_X1 g677 ( .A1(new_n785_), .A2(new_n813_), .ZN(new_n814_) );
  NAND2_X1 g678 ( .A1(new_n810_), .A2(new_n814_), .ZN(new_n815_) );
  INV_X1 g679 ( .A(new_n810_), .ZN(new_n816_) );
  NAND3_X1 g680 ( .A1(new_n816_), .A2(new_n785_), .A3(new_n813_), .ZN(new_n817_) );
  NAND4_X1 g681 ( .A1(new_n798_), .A2(new_n817_), .A3(new_n678_), .A4(new_n815_), .ZN(new_n818_) );
  NAND2_X1 g682 ( .A1(new_n537_), .A2(new_n599_), .ZN(new_n819_) );
  NAND2_X1 g683 ( .A1(new_n627_), .A2(G50), .ZN(new_n820_) );
  NOR2_X1 g684 ( .A1(new_n624_), .A2(new_n346_), .ZN(new_n821_) );
  INV_X1 g685 ( .A(new_n821_), .ZN(new_n822_) );
  NAND2_X1 g686 ( .A1(new_n657_), .A2(G77), .ZN(new_n823_) );
  NAND2_X1 g687 ( .A1(new_n650_), .A2(G150), .ZN(new_n824_) );
  NAND2_X1 g688 ( .A1(new_n652_), .A2(G58), .ZN(new_n825_) );
  NAND2_X1 g689 ( .A1(new_n648_), .A2(G143), .ZN(new_n826_) );
  NAND3_X1 g690 ( .A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_) );
  NAND2_X1 g691 ( .A1(new_n659_), .A2(G137), .ZN(new_n828_) );
  NAND2_X1 g692 ( .A1(new_n635_), .A2(G159), .ZN(new_n829_) );
  NAND2_X1 g693 ( .A1(new_n828_), .A2(new_n829_), .ZN(new_n830_) );
  NOR3_X1 g694 ( .A1(new_n830_), .A2(new_n644_), .A3(new_n827_), .ZN(new_n831_) );
  NAND4_X1 g695 ( .A1(new_n831_), .A2(new_n820_), .A3(new_n822_), .A4(new_n823_), .ZN(new_n832_) );
  NOR2_X1 g696 ( .A1(new_n645_), .A2(new_n140_), .ZN(new_n833_) );
  INV_X1 g697 ( .A(new_n833_), .ZN(new_n834_) );
  NAND2_X1 g698 ( .A1(new_n659_), .A2(G317), .ZN(new_n835_) );
  NAND2_X1 g699 ( .A1(new_n834_), .A2(new_n835_), .ZN(new_n836_) );
  INV_X1 g700 ( .A(G294), .ZN(new_n837_) );
  NOR2_X1 g701 ( .A1(new_n636_), .A2(new_n837_), .ZN(new_n838_) );
  NOR2_X1 g702 ( .A1(new_n628_), .A2(new_n728_), .ZN(new_n839_) );
  INV_X1 g703 ( .A(new_n662_), .ZN(new_n840_) );
  NOR2_X1 g704 ( .A1(new_n624_), .A2(new_n141_), .ZN(new_n841_) );
  INV_X1 g705 ( .A(new_n652_), .ZN(new_n842_) );
  NOR2_X1 g706 ( .A1(new_n842_), .A2(new_n474_), .ZN(new_n843_) );
  INV_X1 g707 ( .A(G303), .ZN(new_n844_) );
  NOR2_X1 g708 ( .A1(new_n664_), .A2(new_n844_), .ZN(new_n845_) );
  NOR3_X1 g709 ( .A1(new_n841_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_) );
  NAND2_X1 g710 ( .A1(new_n648_), .A2(G311), .ZN(new_n847_) );
  XNOR2_X1 g711 ( .A(new_n847_), .B(KEYINPUT54), .ZN(new_n848_) );
  NAND3_X1 g712 ( .A1(new_n846_), .A2(new_n840_), .A3(new_n848_), .ZN(new_n849_) );
  NOR4_X1 g713 ( .A1(new_n849_), .A2(new_n836_), .A3(new_n838_), .A4(new_n839_), .ZN(new_n850_) );
  NAND2_X1 g714 ( .A1(new_n605_), .A2(new_n184_), .ZN(new_n851_) );
  NAND2_X1 g715 ( .A1(new_n590_), .A2(G87), .ZN(new_n852_) );
  NAND3_X1 g716 ( .A1(new_n851_), .A2(new_n619_), .A3(new_n852_), .ZN(new_n853_) );
  INV_X1 g717 ( .A(new_n853_), .ZN(new_n854_) );
  NOR3_X1 g718 ( .A1(new_n850_), .A2(new_n678_), .A3(new_n854_), .ZN(new_n855_) );
  NAND3_X1 g719 ( .A1(new_n819_), .A2(new_n832_), .A3(new_n855_), .ZN(new_n856_) );
  NAND3_X1 g720 ( .A1(new_n818_), .A2(new_n779_), .A3(new_n856_), .ZN(new_n857_) );
  NAND2_X1 g721 ( .A1(new_n818_), .A2(new_n856_), .ZN(new_n858_) );
  NAND2_X1 g722 ( .A1(new_n858_), .A2(KEYINPUT55), .ZN(new_n859_) );
  NAND2_X1 g723 ( .A1(new_n859_), .A2(new_n857_), .ZN(new_n860_) );
  INV_X1 g724 ( .A(new_n860_), .ZN(G387) );
  NAND3_X1 g725 ( .A1(new_n796_), .A2(new_n678_), .A3(new_n791_), .ZN(new_n862_) );
  INV_X1 g726 ( .A(new_n791_), .ZN(new_n863_) );
  NAND3_X1 g727 ( .A1(new_n688_), .A2(new_n591_), .A3(new_n863_), .ZN(new_n864_) );
  NAND3_X1 g728 ( .A1(new_n566_), .A2(new_n567_), .A3(new_n599_), .ZN(new_n865_) );
  NAND2_X1 g729 ( .A1(new_n181_), .A2(G45), .ZN(new_n866_) );
  NAND2_X1 g730 ( .A1(G68), .A2(G77), .ZN(new_n867_) );
  NAND4_X1 g731 ( .A1(new_n589_), .A2(new_n169_), .A3(G58), .A4(new_n867_), .ZN(new_n868_) );
  NAND2_X1 g732 ( .A1(new_n868_), .A2(new_n248_), .ZN(new_n869_) );
  XOR2_X1 g733 ( .A(new_n869_), .B(KEYINPUT23), .Z(new_n870_) );
  NAND2_X1 g734 ( .A1(new_n866_), .A2(new_n870_), .ZN(new_n871_) );
  NAND2_X1 g735 ( .A1(new_n871_), .A2(new_n605_), .ZN(new_n872_) );
  INV_X1 g736 ( .A(new_n589_), .ZN(new_n873_) );
  NAND2_X1 g737 ( .A1(new_n873_), .A2(new_n597_), .ZN(new_n874_) );
  NAND2_X1 g738 ( .A1(new_n590_), .A2(new_n141_), .ZN(new_n875_) );
  NAND3_X1 g739 ( .A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_) );
  NAND2_X1 g740 ( .A1(new_n876_), .A2(new_n619_), .ZN(new_n877_) );
  NAND2_X1 g741 ( .A1(new_n623_), .A2(G87), .ZN(new_n878_) );
  NAND2_X1 g742 ( .A1(new_n659_), .A2(G150), .ZN(new_n879_) );
  NAND2_X1 g743 ( .A1(new_n635_), .A2(G58), .ZN(new_n880_) );
  NAND3_X1 g744 ( .A1(new_n879_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_) );
  NOR2_X1 g745 ( .A1(new_n664_), .A2(new_n169_), .ZN(new_n882_) );
  NOR2_X1 g746 ( .A1(new_n842_), .A2(new_n300_), .ZN(new_n883_) );
  INV_X1 g747 ( .A(new_n648_), .ZN(new_n884_) );
  NOR2_X1 g748 ( .A1(new_n884_), .A2(new_n630_), .ZN(new_n885_) );
  NOR3_X1 g749 ( .A1(new_n882_), .A2(new_n883_), .A3(new_n885_), .ZN(new_n886_) );
  NAND2_X1 g750 ( .A1(new_n627_), .A2(G68), .ZN(new_n887_) );
  NAND3_X1 g751 ( .A1(new_n886_), .A2(new_n834_), .A3(new_n887_), .ZN(new_n888_) );
  NOR3_X1 g752 ( .A1(new_n888_), .A2(new_n644_), .A3(new_n881_), .ZN(new_n889_) );
  NAND2_X1 g753 ( .A1(new_n652_), .A2(G294), .ZN(new_n890_) );
  NAND2_X1 g754 ( .A1(new_n648_), .A2(G322), .ZN(new_n891_) );
  NAND2_X1 g755 ( .A1(new_n890_), .A2(new_n891_), .ZN(new_n892_) );
  XNOR2_X1 g756 ( .A(new_n892_), .B(KEYINPUT26), .ZN(new_n893_) );
  NAND2_X1 g757 ( .A1(new_n657_), .A2(G116), .ZN(new_n894_) );
  XNOR2_X1 g758 ( .A(new_n894_), .B(KEYINPUT25), .ZN(new_n895_) );
  NAND2_X1 g759 ( .A1(new_n635_), .A2(G311), .ZN(new_n896_) );
  NAND2_X1 g760 ( .A1(new_n623_), .A2(G283), .ZN(new_n897_) );
  NAND2_X1 g761 ( .A1(new_n659_), .A2(G326), .ZN(new_n898_) );
  NAND3_X1 g762 ( .A1(new_n898_), .A2(new_n897_), .A3(new_n896_), .ZN(new_n899_) );
  NAND2_X1 g763 ( .A1(new_n627_), .A2(G303), .ZN(new_n900_) );
  NAND2_X1 g764 ( .A1(new_n650_), .A2(G317), .ZN(new_n901_) );
  NAND3_X1 g765 ( .A1(new_n840_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_) );
  NOR4_X1 g766 ( .A1(new_n902_), .A2(new_n895_), .A3(new_n893_), .A4(new_n899_), .ZN(new_n903_) );
  NOR3_X1 g767 ( .A1(new_n903_), .A2(new_n678_), .A3(new_n889_), .ZN(new_n904_) );
  NAND3_X1 g768 ( .A1(new_n865_), .A2(new_n877_), .A3(new_n904_), .ZN(new_n905_) );
  NAND3_X1 g769 ( .A1(new_n864_), .A2(new_n862_), .A3(new_n905_), .ZN(G393) );
  NAND2_X1 g770 ( .A1(new_n784_), .A2(new_n787_), .ZN(new_n907_) );
  NAND3_X1 g771 ( .A1(new_n573_), .A2(new_n586_), .A3(new_n791_), .ZN(new_n908_) );
  NAND2_X1 g772 ( .A1(new_n907_), .A2(new_n908_), .ZN(new_n909_) );
  NAND4_X1 g773 ( .A1(new_n795_), .A2(new_n909_), .A3(new_n591_), .A4(new_n793_), .ZN(new_n910_) );
  NAND3_X1 g774 ( .A1(new_n794_), .A2(new_n678_), .A3(new_n796_), .ZN(new_n911_) );
  NAND3_X1 g775 ( .A1(new_n811_), .A2(new_n599_), .A3(new_n812_), .ZN(new_n912_) );
  INV_X1 g776 ( .A(KEYINPUT58), .ZN(new_n913_) );
  NOR2_X1 g777 ( .A1(new_n664_), .A2(new_n726_), .ZN(new_n914_) );
  NAND2_X1 g778 ( .A1(new_n623_), .A2(G116), .ZN(new_n915_) );
  NAND2_X1 g779 ( .A1(new_n659_), .A2(G322), .ZN(new_n916_) );
  NAND2_X1 g780 ( .A1(new_n627_), .A2(G294), .ZN(new_n917_) );
  NAND2_X1 g781 ( .A1(new_n635_), .A2(G303), .ZN(new_n918_) );
  NAND4_X1 g782 ( .A1(new_n916_), .A2(new_n915_), .A3(new_n917_), .A4(new_n918_), .ZN(new_n919_) );
  NOR4_X1 g783 ( .A1(new_n919_), .A2(new_n215_), .A3(new_n646_), .A4(new_n914_), .ZN(new_n920_) );
  NAND2_X1 g784 ( .A1(new_n920_), .A2(new_n913_), .ZN(new_n921_) );
  INV_X1 g785 ( .A(new_n920_), .ZN(new_n922_) );
  NAND2_X1 g786 ( .A1(new_n922_), .A2(KEYINPUT58), .ZN(new_n923_) );
  NAND2_X1 g787 ( .A1(new_n652_), .A2(G283), .ZN(new_n924_) );
  NAND2_X1 g788 ( .A1(new_n648_), .A2(G317), .ZN(new_n925_) );
  NAND2_X1 g789 ( .A1(new_n924_), .A2(new_n925_), .ZN(new_n926_) );
  XNOR2_X1 g790 ( .A(new_n926_), .B(KEYINPUT59), .ZN(new_n927_) );
  NAND3_X1 g791 ( .A1(new_n923_), .A2(new_n921_), .A3(new_n927_), .ZN(new_n928_) );
  NOR2_X1 g792 ( .A1(new_n624_), .A2(new_n300_), .ZN(new_n929_) );
  NOR2_X1 g793 ( .A1(new_n664_), .A2(new_n630_), .ZN(new_n930_) );
  NAND2_X1 g794 ( .A1(new_n635_), .A2(G50), .ZN(new_n931_) );
  NAND2_X1 g795 ( .A1(new_n627_), .A2(G58), .ZN(new_n932_) );
  NAND2_X1 g796 ( .A1(new_n659_), .A2(G143), .ZN(new_n933_) );
  NAND3_X1 g797 ( .A1(new_n933_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n934_) );
  NOR4_X1 g798 ( .A1(new_n934_), .A2(new_n929_), .A3(G33), .A4(new_n930_), .ZN(new_n935_) );
  NAND3_X1 g799 ( .A1(new_n648_), .A2(G150), .A3(KEYINPUT56), .ZN(new_n936_) );
  INV_X1 g800 ( .A(KEYINPUT56), .ZN(new_n937_) );
  NAND2_X1 g801 ( .A1(new_n648_), .A2(G150), .ZN(new_n938_) );
  NAND2_X1 g802 ( .A1(new_n938_), .A2(new_n937_), .ZN(new_n939_) );
  NAND2_X1 g803 ( .A1(new_n652_), .A2(G68), .ZN(new_n940_) );
  NAND3_X1 g804 ( .A1(new_n939_), .A2(new_n936_), .A3(new_n940_), .ZN(new_n941_) );
  XNOR2_X1 g805 ( .A(new_n941_), .B(KEYINPUT57), .ZN(new_n942_) );
  NAND3_X1 g806 ( .A1(new_n942_), .A2(new_n935_), .A3(new_n725_), .ZN(new_n943_) );
  NAND2_X1 g807 ( .A1(new_n928_), .A2(new_n943_), .ZN(new_n944_) );
  NAND2_X1 g808 ( .A1(new_n944_), .A2(new_n643_), .ZN(new_n945_) );
  NAND2_X1 g809 ( .A1(new_n189_), .A2(new_n605_), .ZN(new_n946_) );
  NAND2_X1 g810 ( .A1(new_n590_), .A2(G97), .ZN(new_n947_) );
  NAND3_X1 g811 ( .A1(new_n946_), .A2(new_n619_), .A3(new_n947_), .ZN(new_n948_) );
  NAND4_X1 g812 ( .A1(new_n912_), .A2(new_n679_), .A3(new_n945_), .A4(new_n948_), .ZN(new_n949_) );
  NAND2_X1 g813 ( .A1(new_n911_), .A2(new_n949_), .ZN(new_n950_) );
  INV_X1 g814 ( .A(new_n950_), .ZN(new_n951_) );
  NAND2_X1 g815 ( .A1(new_n951_), .A2(new_n910_), .ZN(G390) );
  NAND2_X1 g816 ( .A1(new_n741_), .A2(new_n570_), .ZN(new_n953_) );
  INV_X1 g817 ( .A(new_n586_), .ZN(new_n954_) );
  NAND2_X1 g818 ( .A1(new_n954_), .A2(new_n694_), .ZN(new_n955_) );
  NAND2_X1 g819 ( .A1(new_n953_), .A2(new_n955_), .ZN(new_n956_) );
  NAND2_X1 g820 ( .A1(new_n956_), .A2(new_n760_), .ZN(new_n957_) );
  NAND3_X1 g821 ( .A1(new_n953_), .A2(new_n747_), .A3(new_n955_), .ZN(new_n958_) );
  NAND2_X1 g822 ( .A1(new_n957_), .A2(new_n958_), .ZN(new_n959_) );
  INV_X1 g823 ( .A(KEYINPUT38), .ZN(new_n960_) );
  NAND3_X1 g824 ( .A1(new_n377_), .A2(G330), .A3(new_n585_), .ZN(new_n961_) );
  NAND3_X1 g825 ( .A1(new_n555_), .A2(new_n757_), .A3(new_n961_), .ZN(new_n962_) );
  XNOR2_X1 g826 ( .A(new_n962_), .B(new_n960_), .ZN(new_n963_) );
  INV_X1 g827 ( .A(KEYINPUT39), .ZN(new_n964_) );
  NAND4_X1 g828 ( .A1(new_n747_), .A2(new_n585_), .A3(G330), .A4(new_n694_), .ZN(new_n965_) );
  XNOR2_X1 g829 ( .A(new_n965_), .B(new_n964_), .ZN(new_n966_) );
  XNOR2_X1 g830 ( .A(new_n761_), .B(KEYINPUT40), .ZN(new_n967_) );
  NAND4_X1 g831 ( .A1(new_n966_), .A2(new_n748_), .A3(new_n749_), .A4(new_n967_), .ZN(new_n968_) );
  NAND3_X1 g832 ( .A1(new_n966_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n969_) );
  INV_X1 g833 ( .A(new_n967_), .ZN(new_n970_) );
  NAND2_X1 g834 ( .A1(new_n969_), .A2(new_n970_), .ZN(new_n971_) );
  NAND2_X1 g835 ( .A1(new_n971_), .A2(new_n968_), .ZN(new_n972_) );
  INV_X1 g836 ( .A(new_n972_), .ZN(new_n973_) );
  NAND3_X1 g837 ( .A1(new_n973_), .A2(new_n959_), .A3(new_n963_), .ZN(new_n974_) );
  NAND2_X1 g838 ( .A1(new_n959_), .A2(new_n963_), .ZN(new_n975_) );
  NAND2_X1 g839 ( .A1(new_n975_), .A2(new_n972_), .ZN(new_n976_) );
  NAND3_X1 g840 ( .A1(new_n974_), .A2(new_n591_), .A3(new_n976_), .ZN(new_n977_) );
  NAND2_X1 g841 ( .A1(new_n973_), .A2(new_n676_), .ZN(new_n978_) );
  NAND2_X1 g842 ( .A1(new_n761_), .A2(new_n597_), .ZN(new_n979_) );
  NAND2_X1 g843 ( .A1(new_n623_), .A2(G159), .ZN(new_n980_) );
  NAND2_X1 g844 ( .A1(new_n659_), .A2(G125), .ZN(new_n981_) );
  NAND2_X1 g845 ( .A1(new_n635_), .A2(G137), .ZN(new_n982_) );
  NAND2_X1 g846 ( .A1(new_n650_), .A2(G132), .ZN(new_n983_) );
  NAND2_X1 g847 ( .A1(new_n652_), .A2(G150), .ZN(new_n984_) );
  NAND2_X1 g848 ( .A1(new_n648_), .A2(G128), .ZN(new_n985_) );
  NAND3_X1 g849 ( .A1(new_n983_), .A2(new_n984_), .A3(new_n985_), .ZN(new_n986_) );
  NOR2_X1 g850 ( .A1(new_n645_), .A2(new_n169_), .ZN(new_n987_) );
  INV_X1 g851 ( .A(G143), .ZN(new_n988_) );
  NOR2_X1 g852 ( .A1(new_n628_), .A2(new_n988_), .ZN(new_n989_) );
  NOR4_X1 g853 ( .A1(new_n644_), .A2(new_n986_), .A3(new_n987_), .A4(new_n989_), .ZN(new_n990_) );
  NAND4_X1 g854 ( .A1(new_n990_), .A2(new_n980_), .A3(new_n981_), .A4(new_n982_), .ZN(new_n991_) );
  NOR2_X1 g855 ( .A1(new_n633_), .A2(new_n837_), .ZN(new_n992_) );
  NOR2_X1 g856 ( .A1(new_n628_), .A2(new_n140_), .ZN(new_n993_) );
  NOR2_X1 g857 ( .A1(new_n993_), .A2(new_n992_), .ZN(new_n994_) );
  XNOR2_X1 g858 ( .A(new_n994_), .B(KEYINPUT48), .ZN(new_n995_) );
  NAND2_X1 g859 ( .A1(new_n650_), .A2(G116), .ZN(new_n996_) );
  NOR2_X1 g860 ( .A1(new_n996_), .A2(KEYINPUT47), .ZN(new_n997_) );
  NAND2_X1 g861 ( .A1(new_n996_), .A2(KEYINPUT47), .ZN(new_n998_) );
  NAND2_X1 g862 ( .A1(new_n635_), .A2(G107), .ZN(new_n999_) );
  NAND2_X1 g863 ( .A1(new_n998_), .A2(new_n999_), .ZN(new_n1000_) );
  NAND2_X1 g864 ( .A1(new_n648_), .A2(G283), .ZN(new_n1001_) );
  NAND4_X1 g865 ( .A1(new_n840_), .A2(new_n653_), .A3(new_n701_), .A4(new_n1001_), .ZN(new_n1002_) );
  NOR4_X1 g866 ( .A1(new_n1002_), .A2(new_n929_), .A3(new_n997_), .A4(new_n1000_), .ZN(new_n1003_) );
  NAND2_X1 g867 ( .A1(new_n1003_), .A2(new_n995_), .ZN(new_n1004_) );
  NAND2_X1 g868 ( .A1(new_n733_), .A2(new_n225_), .ZN(new_n1005_) );
  NAND3_X1 g869 ( .A1(new_n1004_), .A2(new_n679_), .A3(new_n1005_), .ZN(new_n1006_) );
  INV_X1 g870 ( .A(new_n1006_), .ZN(new_n1007_) );
  NAND3_X1 g871 ( .A1(new_n979_), .A2(new_n991_), .A3(new_n1007_), .ZN(new_n1008_) );
  NAND2_X1 g872 ( .A1(new_n978_), .A2(new_n1008_), .ZN(new_n1009_) );
  INV_X1 g873 ( .A(new_n1009_), .ZN(new_n1010_) );
  NAND2_X1 g874 ( .A1(new_n1010_), .A2(new_n977_), .ZN(G378) );
  NAND4_X1 g875 ( .A1(new_n959_), .A2(new_n971_), .A3(KEYINPUT41), .A4(new_n968_), .ZN(new_n1012_) );
  INV_X1 g876 ( .A(KEYINPUT41), .ZN(new_n1013_) );
  NAND3_X1 g877 ( .A1(new_n959_), .A2(new_n971_), .A3(new_n968_), .ZN(new_n1014_) );
  NAND2_X1 g878 ( .A1(new_n1014_), .A2(new_n1013_), .ZN(new_n1015_) );
  NAND2_X1 g879 ( .A1(new_n1015_), .A2(new_n1012_), .ZN(new_n1016_) );
  NAND3_X1 g880 ( .A1(new_n1016_), .A2(new_n677_), .A3(new_n963_), .ZN(new_n1017_) );
  NAND2_X1 g881 ( .A1(new_n763_), .A2(new_n954_), .ZN(new_n1018_) );
  NAND3_X1 g882 ( .A1(new_n755_), .A2(new_n739_), .A3(new_n1018_), .ZN(new_n1019_) );
  NAND2_X1 g883 ( .A1(new_n319_), .A2(new_n751_), .ZN(new_n1020_) );
  NAND2_X1 g884 ( .A1(new_n345_), .A2(new_n1020_), .ZN(new_n1021_) );
  NAND3_X1 g885 ( .A1(new_n337_), .A2(new_n319_), .A3(new_n751_), .ZN(new_n1022_) );
  NAND2_X1 g886 ( .A1(new_n1021_), .A2(new_n1022_), .ZN(new_n1023_) );
  NAND2_X1 g887 ( .A1(new_n1019_), .A2(new_n1023_), .ZN(new_n1024_) );
  INV_X1 g888 ( .A(new_n1024_), .ZN(new_n1025_) );
  INV_X1 g889 ( .A(new_n1023_), .ZN(new_n1026_) );
  NAND4_X1 g890 ( .A1(new_n755_), .A2(new_n739_), .A3(new_n1018_), .A4(new_n1026_), .ZN(new_n1027_) );
  INV_X1 g891 ( .A(new_n1027_), .ZN(new_n1028_) );
  NOR3_X1 g892 ( .A1(new_n1025_), .A2(new_n679_), .A3(new_n1028_), .ZN(new_n1029_) );
  NAND2_X1 g893 ( .A1(new_n1017_), .A2(new_n1029_), .ZN(new_n1030_) );
  NAND2_X1 g894 ( .A1(new_n1026_), .A2(new_n597_), .ZN(new_n1031_) );
  NAND2_X1 g895 ( .A1(new_n657_), .A2(G159), .ZN(new_n1032_) );
  NAND2_X1 g896 ( .A1(new_n635_), .A2(G132), .ZN(new_n1033_) );
  NAND2_X1 g897 ( .A1(new_n1032_), .A2(new_n1033_), .ZN(new_n1034_) );
  NOR2_X1 g898 ( .A1(new_n1034_), .A2(KEYINPUT44), .ZN(new_n1035_) );
  NAND2_X1 g899 ( .A1(new_n652_), .A2(G143), .ZN(new_n1036_) );
  NAND2_X1 g900 ( .A1(new_n650_), .A2(G128), .ZN(new_n1037_) );
  NAND2_X1 g901 ( .A1(new_n648_), .A2(G125), .ZN(new_n1038_) );
  NAND3_X1 g902 ( .A1(new_n1036_), .A2(new_n1037_), .A3(new_n1038_), .ZN(new_n1039_) );
  NAND2_X1 g903 ( .A1(new_n623_), .A2(G150), .ZN(new_n1040_) );
  NAND2_X1 g904 ( .A1(new_n659_), .A2(G124), .ZN(new_n1041_) );
  NAND2_X1 g905 ( .A1(new_n1041_), .A2(new_n1040_), .ZN(new_n1042_) );
  NOR3_X1 g906 ( .A1(new_n1035_), .A2(new_n1039_), .A3(new_n1042_), .ZN(new_n1043_) );
  NAND2_X1 g907 ( .A1(new_n1034_), .A2(KEYINPUT44), .ZN(new_n1044_) );
  NAND2_X1 g908 ( .A1(new_n627_), .A2(G137), .ZN(new_n1045_) );
  XOR2_X1 g909 ( .A(new_n1045_), .B(KEYINPUT43), .Z(new_n1046_) );
  NAND3_X1 g910 ( .A1(new_n1043_), .A2(new_n1044_), .A3(new_n1046_), .ZN(new_n1047_) );
  NAND2_X1 g911 ( .A1(new_n1047_), .A2(new_n215_), .ZN(new_n1048_) );
  NOR2_X1 g912 ( .A1(new_n645_), .A2(new_n225_), .ZN(new_n1049_) );
  NOR2_X1 g913 ( .A1(new_n628_), .A2(new_n503_), .ZN(new_n1050_) );
  NAND2_X1 g914 ( .A1(new_n650_), .A2(G107), .ZN(new_n1051_) );
  XOR2_X1 g915 ( .A(new_n1051_), .B(KEYINPUT42), .Z(new_n1052_) );
  NOR3_X1 g916 ( .A1(new_n1052_), .A2(new_n1049_), .A3(new_n1050_), .ZN(new_n1053_) );
  NOR2_X1 g917 ( .A1(new_n884_), .A2(new_n474_), .ZN(new_n1054_) );
  NOR3_X1 g918 ( .A1(new_n821_), .A2(new_n883_), .A3(new_n1054_), .ZN(new_n1055_) );
  NAND2_X1 g919 ( .A1(new_n659_), .A2(G283), .ZN(new_n1056_) );
  NAND2_X1 g920 ( .A1(new_n635_), .A2(G97), .ZN(new_n1057_) );
  NAND4_X1 g921 ( .A1(new_n1053_), .A2(new_n1055_), .A3(new_n1056_), .A4(new_n1057_), .ZN(new_n1058_) );
  NAND2_X1 g922 ( .A1(new_n1058_), .A2(G33), .ZN(new_n1059_) );
  NAND4_X1 g923 ( .A1(new_n1048_), .A2(new_n1059_), .A3(new_n247_), .A4(new_n643_), .ZN(new_n1060_) );
  NAND2_X1 g924 ( .A1(new_n643_), .A2(new_n247_), .ZN(new_n1061_) );
  NAND3_X1 g925 ( .A1(new_n1061_), .A2(new_n169_), .A3(new_n598_), .ZN(new_n1062_) );
  NAND4_X1 g926 ( .A1(new_n1031_), .A2(new_n679_), .A3(new_n1060_), .A4(new_n1062_), .ZN(new_n1063_) );
  NAND2_X1 g927 ( .A1(new_n1030_), .A2(new_n1063_), .ZN(G375) );
  XNOR2_X1 g928 ( .A(new_n962_), .B(KEYINPUT38), .ZN(new_n1065_) );
  NAND3_X1 g929 ( .A1(new_n1065_), .A2(new_n957_), .A3(new_n958_), .ZN(new_n1066_) );
  NAND3_X1 g930 ( .A1(new_n975_), .A2(new_n1066_), .A3(KEYINPUT46), .ZN(new_n1067_) );
  INV_X1 g931 ( .A(KEYINPUT46), .ZN(new_n1068_) );
  NAND2_X1 g932 ( .A1(new_n975_), .A2(new_n1066_), .ZN(new_n1069_) );
  NAND2_X1 g933 ( .A1(new_n1069_), .A2(new_n1068_), .ZN(new_n1070_) );
  NAND2_X1 g934 ( .A1(new_n1070_), .A2(new_n1067_), .ZN(new_n1071_) );
  NAND2_X1 g935 ( .A1(new_n1071_), .A2(new_n591_), .ZN(new_n1072_) );
  NAND2_X1 g936 ( .A1(new_n959_), .A2(new_n676_), .ZN(new_n1073_) );
  NAND2_X1 g937 ( .A1(new_n760_), .A2(new_n597_), .ZN(new_n1074_) );
  NAND2_X1 g938 ( .A1(new_n623_), .A2(G50), .ZN(new_n1075_) );
  NAND2_X1 g939 ( .A1(new_n659_), .A2(G128), .ZN(new_n1076_) );
  NAND2_X1 g940 ( .A1(new_n627_), .A2(G150), .ZN(new_n1077_) );
  NAND2_X1 g941 ( .A1(new_n650_), .A2(G137), .ZN(new_n1078_) );
  NAND2_X1 g942 ( .A1(new_n652_), .A2(G159), .ZN(new_n1079_) );
  NAND2_X1 g943 ( .A1(new_n648_), .A2(G132), .ZN(new_n1080_) );
  NAND3_X1 g944 ( .A1(new_n1078_), .A2(new_n1079_), .A3(new_n1080_), .ZN(new_n1081_) );
  NOR2_X1 g945 ( .A1(new_n636_), .A2(new_n988_), .ZN(new_n1082_) );
  NOR4_X1 g946 ( .A1(new_n644_), .A2(new_n1081_), .A3(new_n1049_), .A4(new_n1082_), .ZN(new_n1083_) );
  NAND4_X1 g947 ( .A1(new_n1083_), .A2(new_n1075_), .A3(new_n1076_), .A4(new_n1077_), .ZN(new_n1084_) );
  NOR2_X1 g948 ( .A1(new_n636_), .A2(new_n474_), .ZN(new_n1085_) );
  NOR2_X1 g949 ( .A1(new_n633_), .A2(new_n844_), .ZN(new_n1086_) );
  NOR2_X1 g950 ( .A1(new_n628_), .A2(new_n141_), .ZN(new_n1087_) );
  NOR3_X1 g951 ( .A1(new_n1085_), .A2(new_n1087_), .A3(new_n1086_), .ZN(new_n1088_) );
  NOR2_X1 g952 ( .A1(new_n664_), .A2(new_n728_), .ZN(new_n1089_) );
  NOR2_X1 g953 ( .A1(new_n842_), .A2(new_n140_), .ZN(new_n1090_) );
  NOR2_X1 g954 ( .A1(new_n884_), .A2(new_n837_), .ZN(new_n1091_) );
  NAND2_X1 g955 ( .A1(new_n823_), .A2(new_n878_), .ZN(new_n1092_) );
  NOR4_X1 g956 ( .A1(new_n1092_), .A2(new_n1089_), .A3(new_n1090_), .A4(new_n1091_), .ZN(new_n1093_) );
  NAND3_X1 g957 ( .A1(new_n1093_), .A2(new_n840_), .A3(new_n1088_), .ZN(new_n1094_) );
  NAND2_X1 g958 ( .A1(new_n733_), .A2(new_n346_), .ZN(new_n1095_) );
  NAND4_X1 g959 ( .A1(new_n1084_), .A2(new_n1094_), .A3(new_n679_), .A4(new_n1095_), .ZN(new_n1096_) );
  XNOR2_X1 g960 ( .A(new_n1096_), .B(KEYINPUT45), .ZN(new_n1097_) );
  NAND2_X1 g961 ( .A1(new_n1074_), .A2(new_n1097_), .ZN(new_n1098_) );
  NAND2_X1 g962 ( .A1(new_n1073_), .A2(new_n1098_), .ZN(new_n1099_) );
  INV_X1 g963 ( .A(new_n1099_), .ZN(new_n1100_) );
  NAND2_X1 g964 ( .A1(new_n1072_), .A2(new_n1100_), .ZN(G381) );
  INV_X1 g965 ( .A(G381), .ZN(new_n1102_) );
  INV_X1 g966 ( .A(G378), .ZN(new_n1103_) );
  NAND3_X1 g967 ( .A1(new_n1103_), .A2(new_n1030_), .A3(new_n1063_), .ZN(new_n1104_) );
  INV_X1 g968 ( .A(new_n1104_), .ZN(new_n1105_) );
  NOR4_X1 g969 ( .A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1106_) );
  NAND4_X1 g970 ( .A1(new_n1105_), .A2(new_n860_), .A3(new_n1102_), .A4(new_n1106_), .ZN(G407) );
  NAND2_X1 g971 ( .A1(new_n1105_), .A2(new_n558_), .ZN(new_n1108_) );
  NAND3_X1 g972 ( .A1(G407), .A2(new_n1108_), .A3(G213), .ZN(G409) );
  NAND2_X1 g973 ( .A1(G375), .A2(G378), .ZN(new_n1110_) );
  NAND2_X1 g974 ( .A1(new_n558_), .A2(G213), .ZN(new_n1111_) );
  NAND3_X1 g975 ( .A1(new_n1110_), .A2(new_n1104_), .A3(new_n1111_), .ZN(new_n1112_) );
  NAND3_X1 g976 ( .A1(new_n558_), .A2(G213), .A3(G2897), .ZN(new_n1113_) );
  XOR2_X1 g977 ( .A(new_n1113_), .B(KEYINPUT63), .Z(new_n1114_) );
  XNOR2_X1 g978 ( .A(G390), .B(G396), .ZN(new_n1115_) );
  NAND2_X1 g979 ( .A1(G381), .A2(new_n1115_), .ZN(new_n1116_) );
  INV_X1 g980 ( .A(G396), .ZN(new_n1117_) );
  XNOR2_X1 g981 ( .A(G390), .B(new_n1117_), .ZN(new_n1118_) );
  NAND3_X1 g982 ( .A1(new_n1118_), .A2(new_n1072_), .A3(new_n1100_), .ZN(new_n1119_) );
  NAND2_X1 g983 ( .A1(new_n1116_), .A2(new_n1119_), .ZN(new_n1120_) );
  XNOR2_X1 g984 ( .A(G384), .B(G393), .ZN(new_n1121_) );
  NAND3_X1 g985 ( .A1(new_n859_), .A2(new_n857_), .A3(new_n1121_), .ZN(new_n1122_) );
  INV_X1 g986 ( .A(new_n1121_), .ZN(new_n1123_) );
  NAND2_X1 g987 ( .A1(new_n860_), .A2(new_n1123_), .ZN(new_n1124_) );
  NAND2_X1 g988 ( .A1(new_n1124_), .A2(new_n1122_), .ZN(new_n1125_) );
  NAND2_X1 g989 ( .A1(new_n1120_), .A2(new_n1125_), .ZN(new_n1126_) );
  NAND4_X1 g990 ( .A1(new_n1116_), .A2(new_n1119_), .A3(new_n1124_), .A4(new_n1122_), .ZN(new_n1127_) );
  NAND2_X1 g991 ( .A1(new_n1126_), .A2(new_n1127_), .ZN(new_n1128_) );
  NAND3_X1 g992 ( .A1(new_n1128_), .A2(new_n1112_), .A3(new_n1114_), .ZN(new_n1129_) );
  NAND2_X1 g993 ( .A1(new_n1112_), .A2(new_n1114_), .ZN(new_n1130_) );
  NAND3_X1 g994 ( .A1(new_n1130_), .A2(new_n1126_), .A3(new_n1127_), .ZN(new_n1131_) );
  NAND2_X1 g995 ( .A1(new_n1129_), .A2(new_n1131_), .ZN(G405) );
  NAND2_X1 g996 ( .A1(new_n1110_), .A2(new_n1104_), .ZN(new_n1133_) );
  NAND2_X1 g997 ( .A1(new_n1128_), .A2(new_n1133_), .ZN(new_n1134_) );
  NAND4_X1 g998 ( .A1(new_n1126_), .A2(new_n1104_), .A3(new_n1110_), .A4(new_n1127_), .ZN(new_n1135_) );
  NAND2_X1 g999 ( .A1(new_n1134_), .A2(new_n1135_), .ZN(G402) );
endmodule


