module add_mul_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, 
        b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, operation, Result_0_, 
        Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, 
        Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, 
        Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959;

  NAND2_X1 U464 ( .A1(n448), .A2(n449), .ZN(Result_9_) );
  NAND2_X1 U465 ( .A1(n450), .A2(n451), .ZN(n449) );
  NAND2_X1 U466 ( .A1(n452), .A2(n453), .ZN(n450) );
  NAND2_X1 U467 ( .A1(n454), .A2(n455), .ZN(n453) );
  OR2_X1 U468 ( .A1(n456), .A2(n457), .ZN(n454) );
  NAND2_X1 U469 ( .A1(n458), .A2(n459), .ZN(n452) );
  XOR2_X1 U470 ( .A(b_1_), .B(a_1_), .Z(n458) );
  NAND2_X1 U471 ( .A1(n460), .A2(operation), .ZN(n448) );
  XOR2_X1 U472 ( .A(n461), .B(n462), .Z(n460) );
  XOR2_X1 U473 ( .A(n463), .B(n464), .Z(n462) );
  NOR2_X1 U474 ( .A1(n465), .A2(n466), .ZN(n464) );
  NAND2_X1 U475 ( .A1(n467), .A2(n468), .ZN(Result_8_) );
  NAND2_X1 U476 ( .A1(n469), .A2(n451), .ZN(n468) );
  XOR2_X1 U477 ( .A(n470), .B(n471), .Z(n469) );
  NOR2_X1 U478 ( .A1(n472), .A2(n473), .ZN(n471) );
  INV_X1 U479 ( .A(n474), .ZN(n473) );
  NOR2_X1 U480 ( .A1(b_0_), .A2(a_0_), .ZN(n472) );
  NOR2_X1 U481 ( .A1(n457), .A2(n475), .ZN(n470) );
  NOR2_X1 U482 ( .A1(n456), .A2(n455), .ZN(n475) );
  INV_X1 U483 ( .A(n459), .ZN(n455) );
  NOR2_X1 U484 ( .A1(n476), .A2(n477), .ZN(n459) );
  NOR2_X1 U485 ( .A1(n478), .A2(n479), .ZN(n477) );
  NOR2_X1 U486 ( .A1(b_1_), .A2(a_1_), .ZN(n457) );
  NAND2_X1 U487 ( .A1(n480), .A2(operation), .ZN(n467) );
  XNOR2_X1 U488 ( .A(n481), .B(n482), .ZN(n480) );
  NAND2_X1 U489 ( .A1(n483), .A2(n484), .ZN(n481) );
  NOR2_X1 U490 ( .A1(n485), .A2(n451), .ZN(Result_7_) );
  XNOR2_X1 U491 ( .A(n486), .B(n487), .ZN(n485) );
  NOR2_X1 U492 ( .A1(n451), .A2(n488), .ZN(Result_6_) );
  NAND2_X1 U493 ( .A1(n489), .A2(n490), .ZN(n488) );
  NAND2_X1 U494 ( .A1(n491), .A2(n492), .ZN(n489) );
  NOR2_X1 U495 ( .A1(n493), .A2(n451), .ZN(Result_5_) );
  XOR2_X1 U496 ( .A(n490), .B(n494), .Z(n493) );
  NOR2_X1 U497 ( .A1(n495), .A2(n496), .ZN(n494) );
  NOR2_X1 U498 ( .A1(n497), .A2(n498), .ZN(n496) );
  INV_X1 U499 ( .A(n499), .ZN(n490) );
  NOR2_X1 U500 ( .A1(n500), .A2(n451), .ZN(Result_4_) );
  XNOR2_X1 U501 ( .A(n501), .B(n502), .ZN(n500) );
  NOR2_X1 U502 ( .A1(n503), .A2(n451), .ZN(Result_3_) );
  XOR2_X1 U503 ( .A(n504), .B(n505), .Z(n503) );
  NAND2_X1 U504 ( .A1(n506), .A2(n507), .ZN(n504) );
  NOR2_X1 U505 ( .A1(n451), .A2(n508), .ZN(Result_2_) );
  XOR2_X1 U506 ( .A(n509), .B(n510), .Z(n508) );
  NAND2_X1 U507 ( .A1(n511), .A2(n512), .ZN(n510) );
  NOR2_X1 U508 ( .A1(n451), .A2(n513), .ZN(Result_1_) );
  XOR2_X1 U509 ( .A(n514), .B(n515), .Z(n513) );
  NAND2_X1 U510 ( .A1(n516), .A2(n517), .ZN(n515) );
  NAND2_X1 U511 ( .A1(n518), .A2(n519), .ZN(Result_15_) );
  NAND2_X1 U512 ( .A1(n520), .A2(n451), .ZN(n519) );
  XOR2_X1 U513 ( .A(b_7_), .B(a_7_), .Z(n520) );
  NAND2_X1 U514 ( .A1(operation), .A2(n521), .ZN(n518) );
  NAND2_X1 U515 ( .A1(n522), .A2(n523), .ZN(Result_14_) );
  NAND2_X1 U516 ( .A1(n524), .A2(n451), .ZN(n523) );
  NAND2_X1 U517 ( .A1(n525), .A2(n526), .ZN(n524) );
  NOR2_X1 U518 ( .A1(n527), .A2(n528), .ZN(n525) );
  NOR2_X1 U519 ( .A1(n529), .A2(n530), .ZN(n528) );
  NAND2_X1 U520 ( .A1(n531), .A2(n532), .ZN(n530) );
  NOR2_X1 U521 ( .A1(b_6_), .A2(n533), .ZN(n527) );
  XOR2_X1 U522 ( .A(n531), .B(a_6_), .Z(n533) );
  NAND2_X1 U523 ( .A1(n534), .A2(operation), .ZN(n522) );
  XOR2_X1 U524 ( .A(n535), .B(n536), .Z(n534) );
  NAND2_X1 U525 ( .A1(b_7_), .A2(a_6_), .ZN(n536) );
  NAND2_X1 U526 ( .A1(n537), .A2(n538), .ZN(Result_13_) );
  NAND2_X1 U527 ( .A1(n539), .A2(n451), .ZN(n538) );
  NAND2_X1 U528 ( .A1(n540), .A2(n541), .ZN(n539) );
  NAND2_X1 U529 ( .A1(n542), .A2(n543), .ZN(n541) );
  NOR2_X1 U530 ( .A1(n544), .A2(n545), .ZN(n540) );
  NOR2_X1 U531 ( .A1(b_5_), .A2(n546), .ZN(n545) );
  XOR2_X1 U532 ( .A(a_5_), .B(n547), .Z(n546) );
  NOR2_X1 U533 ( .A1(n548), .A2(n549), .ZN(n544) );
  NAND2_X1 U534 ( .A1(n547), .A2(n550), .ZN(n549) );
  INV_X1 U535 ( .A(n543), .ZN(n547) );
  NAND2_X1 U536 ( .A1(n551), .A2(operation), .ZN(n537) );
  XNOR2_X1 U537 ( .A(n552), .B(n553), .ZN(n551) );
  XOR2_X1 U538 ( .A(n554), .B(n555), .Z(n553) );
  NAND2_X1 U539 ( .A1(b_7_), .A2(a_5_), .ZN(n554) );
  NAND2_X1 U540 ( .A1(n556), .A2(n557), .ZN(Result_12_) );
  NAND2_X1 U541 ( .A1(n558), .A2(n451), .ZN(n557) );
  XNOR2_X1 U542 ( .A(n559), .B(n560), .ZN(n558) );
  NAND2_X1 U543 ( .A1(n561), .A2(n562), .ZN(n559) );
  NAND2_X1 U544 ( .A1(n563), .A2(operation), .ZN(n556) );
  XNOR2_X1 U545 ( .A(n564), .B(n565), .ZN(n563) );
  NAND2_X1 U546 ( .A1(n566), .A2(n567), .ZN(n564) );
  NAND2_X1 U547 ( .A1(n568), .A2(n569), .ZN(Result_11_) );
  NAND2_X1 U548 ( .A1(n570), .A2(n451), .ZN(n569) );
  NAND2_X1 U549 ( .A1(n571), .A2(n572), .ZN(n570) );
  NAND2_X1 U550 ( .A1(n573), .A2(n574), .ZN(n572) );
  NOR2_X1 U551 ( .A1(n575), .A2(n576), .ZN(n571) );
  NOR2_X1 U552 ( .A1(b_3_), .A2(n577), .ZN(n576) );
  XOR2_X1 U553 ( .A(n578), .B(n574), .Z(n577) );
  NOR2_X1 U554 ( .A1(n579), .A2(n580), .ZN(n575) );
  OR2_X1 U555 ( .A1(n574), .A2(a_3_), .ZN(n580) );
  NAND2_X1 U556 ( .A1(n581), .A2(operation), .ZN(n568) );
  XOR2_X1 U557 ( .A(n582), .B(n583), .Z(n581) );
  XNOR2_X1 U558 ( .A(n584), .B(n585), .ZN(n583) );
  NAND2_X1 U559 ( .A1(b_7_), .A2(a_3_), .ZN(n584) );
  NAND2_X1 U560 ( .A1(n586), .A2(n587), .ZN(Result_10_) );
  NAND2_X1 U561 ( .A1(n588), .A2(n451), .ZN(n587) );
  XNOR2_X1 U562 ( .A(n479), .B(n589), .ZN(n588) );
  NOR2_X1 U563 ( .A1(n478), .A2(n476), .ZN(n589) );
  NOR2_X1 U564 ( .A1(b_2_), .A2(a_2_), .ZN(n478) );
  AND2_X1 U565 ( .A1(n590), .A2(n591), .ZN(n479) );
  NAND2_X1 U566 ( .A1(n592), .A2(n574), .ZN(n591) );
  NAND2_X1 U567 ( .A1(n561), .A2(n593), .ZN(n574) );
  NAND2_X1 U568 ( .A1(n562), .A2(n560), .ZN(n593) );
  OR2_X1 U569 ( .A1(n542), .A2(n594), .ZN(n560) );
  AND2_X1 U570 ( .A1(n595), .A2(n543), .ZN(n594) );
  NAND2_X1 U571 ( .A1(n596), .A2(n597), .ZN(n543) );
  NAND2_X1 U572 ( .A1(n521), .A2(n598), .ZN(n597) );
  NAND2_X1 U573 ( .A1(n529), .A2(n532), .ZN(n598) );
  NAND2_X1 U574 ( .A1(n548), .A2(n550), .ZN(n595) );
  NAND2_X1 U575 ( .A1(n599), .A2(n600), .ZN(n562) );
  NAND2_X1 U576 ( .A1(n579), .A2(n578), .ZN(n592) );
  NAND2_X1 U577 ( .A1(n601), .A2(operation), .ZN(n586) );
  XOR2_X1 U578 ( .A(n602), .B(n603), .Z(n601) );
  XOR2_X1 U579 ( .A(n604), .B(n605), .Z(n603) );
  NOR2_X1 U580 ( .A1(n606), .A2(n451), .ZN(Result_0_) );
  INV_X1 U581 ( .A(operation), .ZN(n451) );
  NOR2_X1 U582 ( .A1(n607), .A2(n608), .ZN(n606) );
  NAND2_X1 U583 ( .A1(n609), .A2(n517), .ZN(n608) );
  NAND2_X1 U584 ( .A1(n610), .A2(n611), .ZN(n517) );
  NOR2_X1 U585 ( .A1(n612), .A2(n613), .ZN(n611) );
  NOR2_X1 U586 ( .A1(n614), .A2(n474), .ZN(n610) );
  NAND2_X1 U587 ( .A1(n516), .A2(n514), .ZN(n609) );
  NAND2_X1 U588 ( .A1(n511), .A2(n615), .ZN(n514) );
  NAND2_X1 U589 ( .A1(n512), .A2(n509), .ZN(n615) );
  NAND2_X1 U590 ( .A1(n506), .A2(n616), .ZN(n509) );
  NAND2_X1 U591 ( .A1(n505), .A2(n507), .ZN(n616) );
  NAND2_X1 U592 ( .A1(n617), .A2(n618), .ZN(n507) );
  NAND2_X1 U593 ( .A1(n619), .A2(n620), .ZN(n618) );
  XOR2_X1 U594 ( .A(n621), .B(n622), .Z(n617) );
  AND2_X1 U595 ( .A1(n501), .A2(n502), .ZN(n505) );
  NAND2_X1 U596 ( .A1(n623), .A2(n624), .ZN(n502) );
  NAND2_X1 U597 ( .A1(n499), .A2(n498), .ZN(n624) );
  NOR2_X1 U598 ( .A1(n492), .A2(n491), .ZN(n499) );
  XNOR2_X1 U599 ( .A(n625), .B(n626), .ZN(n491) );
  OR2_X1 U600 ( .A1(n487), .A2(n486), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n627), .B(n628), .ZN(n486) );
  XOR2_X1 U602 ( .A(n629), .B(n630), .Z(n627) );
  AND2_X1 U603 ( .A1(n483), .A2(n631), .ZN(n487) );
  NAND2_X1 U604 ( .A1(n482), .A2(n484), .ZN(n631) );
  NAND2_X1 U605 ( .A1(n632), .A2(n633), .ZN(n484) );
  NAND2_X1 U606 ( .A1(a_0_), .A2(b_7_), .ZN(n633) );
  INV_X1 U607 ( .A(n634), .ZN(n632) );
  XOR2_X1 U608 ( .A(n635), .B(n636), .Z(n482) );
  XOR2_X1 U609 ( .A(n637), .B(n638), .Z(n635) );
  NAND2_X1 U610 ( .A1(a_0_), .A2(n634), .ZN(n483) );
  NAND2_X1 U611 ( .A1(n639), .A2(n640), .ZN(n634) );
  NAND2_X1 U612 ( .A1(n641), .A2(a_1_), .ZN(n640) );
  NOR2_X1 U613 ( .A1(n642), .A2(n465), .ZN(n641) );
  NOR2_X1 U614 ( .A1(n461), .A2(n463), .ZN(n642) );
  NAND2_X1 U615 ( .A1(n461), .A2(n463), .ZN(n639) );
  NAND2_X1 U616 ( .A1(n643), .A2(n644), .ZN(n463) );
  NAND2_X1 U617 ( .A1(n605), .A2(n645), .ZN(n644) );
  NAND2_X1 U618 ( .A1(n604), .A2(n602), .ZN(n645) );
  NOR2_X1 U619 ( .A1(n465), .A2(n646), .ZN(n605) );
  INV_X1 U620 ( .A(b_7_), .ZN(n465) );
  OR2_X1 U621 ( .A1(n602), .A2(n604), .ZN(n643) );
  AND2_X1 U622 ( .A1(n647), .A2(n648), .ZN(n604) );
  NAND2_X1 U623 ( .A1(n649), .A2(b_7_), .ZN(n648) );
  NOR2_X1 U624 ( .A1(n650), .A2(n578), .ZN(n649) );
  NOR2_X1 U625 ( .A1(n582), .A2(n585), .ZN(n650) );
  NAND2_X1 U626 ( .A1(n582), .A2(n585), .ZN(n647) );
  NAND2_X1 U627 ( .A1(n566), .A2(n651), .ZN(n585) );
  NAND2_X1 U628 ( .A1(n565), .A2(n567), .ZN(n651) );
  NAND2_X1 U629 ( .A1(n652), .A2(n653), .ZN(n567) );
  NAND2_X1 U630 ( .A1(b_7_), .A2(a_4_), .ZN(n653) );
  INV_X1 U631 ( .A(n654), .ZN(n652) );
  XNOR2_X1 U632 ( .A(n655), .B(n656), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n657), .A2(n658), .ZN(n655) );
  NAND2_X1 U634 ( .A1(a_4_), .A2(n654), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n659), .A2(n660), .ZN(n654) );
  NAND2_X1 U636 ( .A1(n661), .A2(b_7_), .ZN(n660) );
  NOR2_X1 U637 ( .A1(n662), .A2(n550), .ZN(n661) );
  NOR2_X1 U638 ( .A1(n555), .A2(n552), .ZN(n662) );
  NAND2_X1 U639 ( .A1(n555), .A2(n552), .ZN(n659) );
  XNOR2_X1 U640 ( .A(n596), .B(n663), .ZN(n552) );
  NOR2_X1 U641 ( .A1(n664), .A2(n548), .ZN(n663) );
  INV_X1 U642 ( .A(n526), .ZN(n555) );
  NAND2_X1 U643 ( .A1(n665), .A2(n521), .ZN(n526) );
  INV_X1 U644 ( .A(n531), .ZN(n521) );
  NAND2_X1 U645 ( .A1(b_7_), .A2(a_7_), .ZN(n531) );
  INV_X1 U646 ( .A(n596), .ZN(n665) );
  NAND2_X1 U647 ( .A1(b_6_), .A2(a_6_), .ZN(n596) );
  XNOR2_X1 U648 ( .A(n666), .B(n667), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n668), .B(n669), .ZN(n667) );
  XNOR2_X1 U650 ( .A(n670), .B(n671), .ZN(n602) );
  XOR2_X1 U651 ( .A(n672), .B(n673), .Z(n670) );
  NOR2_X1 U652 ( .A1(n578), .A2(n529), .ZN(n673) );
  XOR2_X1 U653 ( .A(n674), .B(n675), .Z(n461) );
  XOR2_X1 U654 ( .A(n676), .B(n677), .Z(n674) );
  NOR2_X1 U655 ( .A1(n678), .A2(n495), .ZN(n623) );
  AND2_X1 U656 ( .A1(n497), .A2(n498), .ZN(n495) );
  AND2_X1 U657 ( .A1(n679), .A2(n680), .ZN(n498) );
  NAND2_X1 U658 ( .A1(n681), .A2(n682), .ZN(n679) );
  INV_X1 U659 ( .A(n683), .ZN(n682) );
  XOR2_X1 U660 ( .A(n684), .B(n685), .Z(n681) );
  NOR2_X1 U661 ( .A1(n625), .A2(n626), .ZN(n497) );
  XOR2_X1 U662 ( .A(n686), .B(n687), .Z(n626) );
  NAND2_X1 U663 ( .A1(n688), .A2(n689), .ZN(n686) );
  AND2_X1 U664 ( .A1(n690), .A2(n691), .ZN(n625) );
  NAND2_X1 U665 ( .A1(n629), .A2(n692), .ZN(n691) );
  OR2_X1 U666 ( .A1(n628), .A2(n630), .ZN(n692) );
  NOR2_X1 U667 ( .A1(n693), .A2(n529), .ZN(n629) );
  NAND2_X1 U668 ( .A1(n628), .A2(n630), .ZN(n690) );
  NAND2_X1 U669 ( .A1(n694), .A2(n695), .ZN(n630) );
  NAND2_X1 U670 ( .A1(n638), .A2(n696), .ZN(n695) );
  OR2_X1 U671 ( .A1(n637), .A2(n636), .ZN(n696) );
  NOR2_X1 U672 ( .A1(n466), .A2(n529), .ZN(n638) );
  NAND2_X1 U673 ( .A1(n636), .A2(n637), .ZN(n694) );
  NAND2_X1 U674 ( .A1(n697), .A2(n698), .ZN(n637) );
  NAND2_X1 U675 ( .A1(n677), .A2(n699), .ZN(n698) );
  OR2_X1 U676 ( .A1(n675), .A2(n676), .ZN(n699) );
  NOR2_X1 U677 ( .A1(n646), .A2(n529), .ZN(n677) );
  NAND2_X1 U678 ( .A1(n675), .A2(n676), .ZN(n697) );
  NAND2_X1 U679 ( .A1(n700), .A2(n701), .ZN(n676) );
  NAND2_X1 U680 ( .A1(n702), .A2(b_6_), .ZN(n701) );
  NOR2_X1 U681 ( .A1(n703), .A2(n578), .ZN(n702) );
  NOR2_X1 U682 ( .A1(n671), .A2(n672), .ZN(n703) );
  NAND2_X1 U683 ( .A1(n671), .A2(n672), .ZN(n700) );
  NAND2_X1 U684 ( .A1(n704), .A2(n705), .ZN(n672) );
  NAND2_X1 U685 ( .A1(n669), .A2(n706), .ZN(n705) );
  OR2_X1 U686 ( .A1(n668), .A2(n666), .ZN(n706) );
  NOR2_X1 U687 ( .A1(n529), .A2(n600), .ZN(n669) );
  INV_X1 U688 ( .A(b_6_), .ZN(n529) );
  NAND2_X1 U689 ( .A1(n666), .A2(n668), .ZN(n704) );
  NAND2_X1 U690 ( .A1(n657), .A2(n707), .ZN(n668) );
  NAND2_X1 U691 ( .A1(n656), .A2(n658), .ZN(n707) );
  NAND2_X1 U692 ( .A1(n708), .A2(n709), .ZN(n658) );
  INV_X1 U693 ( .A(n710), .ZN(n709) );
  NAND2_X1 U694 ( .A1(b_6_), .A2(a_5_), .ZN(n708) );
  XNOR2_X1 U695 ( .A(n711), .B(n712), .ZN(n656) );
  NOR2_X1 U696 ( .A1(n664), .A2(n599), .ZN(n712) );
  NAND2_X1 U697 ( .A1(n710), .A2(a_5_), .ZN(n657) );
  NOR2_X1 U698 ( .A1(n535), .A2(n711), .ZN(n710) );
  NAND2_X1 U699 ( .A1(b_6_), .A2(a_7_), .ZN(n535) );
  XNOR2_X1 U700 ( .A(n713), .B(n714), .ZN(n666) );
  XNOR2_X1 U701 ( .A(n542), .B(n715), .ZN(n713) );
  XNOR2_X1 U702 ( .A(n716), .B(n717), .ZN(n671) );
  NAND2_X1 U703 ( .A1(n718), .A2(n719), .ZN(n716) );
  XOR2_X1 U704 ( .A(n720), .B(n721), .Z(n675) );
  XOR2_X1 U705 ( .A(n722), .B(n723), .Z(n720) );
  NOR2_X1 U706 ( .A1(n548), .A2(n578), .ZN(n723) );
  XNOR2_X1 U707 ( .A(n724), .B(n725), .ZN(n636) );
  XOR2_X1 U708 ( .A(n726), .B(n727), .Z(n725) );
  NAND2_X1 U709 ( .A1(a_2_), .A2(b_5_), .ZN(n727) );
  XOR2_X1 U710 ( .A(n728), .B(n729), .Z(n628) );
  XOR2_X1 U711 ( .A(n730), .B(n731), .Z(n729) );
  INV_X1 U712 ( .A(n680), .ZN(n678) );
  NAND2_X1 U713 ( .A1(n732), .A2(n683), .ZN(n680) );
  NAND2_X1 U714 ( .A1(n688), .A2(n733), .ZN(n683) );
  NAND2_X1 U715 ( .A1(n687), .A2(n689), .ZN(n733) );
  NAND2_X1 U716 ( .A1(n734), .A2(n735), .ZN(n689) );
  NAND2_X1 U717 ( .A1(a_0_), .A2(b_5_), .ZN(n735) );
  INV_X1 U718 ( .A(n736), .ZN(n734) );
  XNOR2_X1 U719 ( .A(n737), .B(n738), .ZN(n687) );
  NAND2_X1 U720 ( .A1(n739), .A2(n740), .ZN(n737) );
  NAND2_X1 U721 ( .A1(a_0_), .A2(n736), .ZN(n688) );
  NAND2_X1 U722 ( .A1(n741), .A2(n742), .ZN(n736) );
  NAND2_X1 U723 ( .A1(n731), .A2(n743), .ZN(n742) );
  NAND2_X1 U724 ( .A1(n730), .A2(n728), .ZN(n743) );
  NOR2_X1 U725 ( .A1(n466), .A2(n548), .ZN(n731) );
  OR2_X1 U726 ( .A1(n728), .A2(n730), .ZN(n741) );
  AND2_X1 U727 ( .A1(n744), .A2(n745), .ZN(n730) );
  NAND2_X1 U728 ( .A1(n746), .A2(a_2_), .ZN(n745) );
  NOR2_X1 U729 ( .A1(n747), .A2(n548), .ZN(n746) );
  NOR2_X1 U730 ( .A1(n726), .A2(n724), .ZN(n747) );
  NAND2_X1 U731 ( .A1(n724), .A2(n726), .ZN(n744) );
  NAND2_X1 U732 ( .A1(n748), .A2(n749), .ZN(n726) );
  NAND2_X1 U733 ( .A1(n750), .A2(a_3_), .ZN(n749) );
  NOR2_X1 U734 ( .A1(n751), .A2(n548), .ZN(n750) );
  NOR2_X1 U735 ( .A1(n721), .A2(n722), .ZN(n751) );
  NAND2_X1 U736 ( .A1(n721), .A2(n722), .ZN(n748) );
  NAND2_X1 U737 ( .A1(n718), .A2(n752), .ZN(n722) );
  NAND2_X1 U738 ( .A1(n717), .A2(n719), .ZN(n752) );
  NAND2_X1 U739 ( .A1(n753), .A2(n754), .ZN(n719) );
  NAND2_X1 U740 ( .A1(b_5_), .A2(a_4_), .ZN(n754) );
  INV_X1 U741 ( .A(n755), .ZN(n753) );
  XOR2_X1 U742 ( .A(n756), .B(n757), .Z(n717) );
  NOR2_X1 U743 ( .A1(n758), .A2(n759), .ZN(n757) );
  NOR2_X1 U744 ( .A1(n760), .A2(n761), .ZN(n758) );
  NOR2_X1 U745 ( .A1(n550), .A2(n599), .ZN(n761) );
  INV_X1 U746 ( .A(n762), .ZN(n760) );
  NAND2_X1 U747 ( .A1(a_4_), .A2(n755), .ZN(n718) );
  NAND2_X1 U748 ( .A1(n763), .A2(n764), .ZN(n755) );
  NAND2_X1 U749 ( .A1(n715), .A2(n765), .ZN(n764) );
  OR2_X1 U750 ( .A1(n714), .A2(n542), .ZN(n765) );
  NOR2_X1 U751 ( .A1(n766), .A2(n711), .ZN(n715) );
  NAND2_X1 U752 ( .A1(b_5_), .A2(a_6_), .ZN(n711) );
  NAND2_X1 U753 ( .A1(a_7_), .A2(b_4_), .ZN(n766) );
  NAND2_X1 U754 ( .A1(n542), .A2(n714), .ZN(n763) );
  XOR2_X1 U755 ( .A(n767), .B(n768), .Z(n714) );
  NOR2_X1 U756 ( .A1(n548), .A2(n550), .ZN(n542) );
  INV_X1 U757 ( .A(b_5_), .ZN(n548) );
  XNOR2_X1 U758 ( .A(n769), .B(n770), .ZN(n721) );
  XOR2_X1 U759 ( .A(n561), .B(n771), .Z(n769) );
  XNOR2_X1 U760 ( .A(n772), .B(n773), .ZN(n724) );
  XOR2_X1 U761 ( .A(n774), .B(n775), .Z(n773) );
  XOR2_X1 U762 ( .A(n776), .B(n777), .Z(n728) );
  NAND2_X1 U763 ( .A1(n778), .A2(n779), .ZN(n776) );
  XNOR2_X1 U764 ( .A(n684), .B(n685), .ZN(n732) );
  XNOR2_X1 U765 ( .A(n780), .B(n781), .ZN(n684) );
  NOR2_X1 U766 ( .A1(n599), .A2(n693), .ZN(n781) );
  XOR2_X1 U767 ( .A(n620), .B(n619), .Z(n501) );
  NAND2_X1 U768 ( .A1(n782), .A2(n783), .ZN(n506) );
  XOR2_X1 U769 ( .A(n622), .B(n784), .Z(n783) );
  INV_X1 U770 ( .A(n621), .ZN(n784) );
  AND2_X1 U771 ( .A1(n620), .A2(n619), .ZN(n782) );
  XOR2_X1 U772 ( .A(n785), .B(n786), .Z(n619) );
  XNOR2_X1 U773 ( .A(n787), .B(n788), .ZN(n786) );
  NAND2_X1 U774 ( .A1(a_0_), .A2(b_3_), .ZN(n788) );
  NAND2_X1 U775 ( .A1(n789), .A2(n790), .ZN(n620) );
  NAND2_X1 U776 ( .A1(n791), .A2(a_0_), .ZN(n790) );
  NOR2_X1 U777 ( .A1(n792), .A2(n599), .ZN(n791) );
  NOR2_X1 U778 ( .A1(n685), .A2(n780), .ZN(n792) );
  NAND2_X1 U779 ( .A1(n685), .A2(n780), .ZN(n789) );
  NAND2_X1 U780 ( .A1(n739), .A2(n793), .ZN(n780) );
  NAND2_X1 U781 ( .A1(n738), .A2(n740), .ZN(n793) );
  NAND2_X1 U782 ( .A1(n794), .A2(n795), .ZN(n740) );
  NAND2_X1 U783 ( .A1(a_1_), .A2(b_4_), .ZN(n795) );
  INV_X1 U784 ( .A(n796), .ZN(n794) );
  XNOR2_X1 U785 ( .A(n797), .B(n798), .ZN(n738) );
  XOR2_X1 U786 ( .A(n799), .B(n800), .Z(n797) );
  NAND2_X1 U787 ( .A1(a_2_), .A2(b_3_), .ZN(n799) );
  NAND2_X1 U788 ( .A1(a_1_), .A2(n796), .ZN(n739) );
  NAND2_X1 U789 ( .A1(n778), .A2(n801), .ZN(n796) );
  NAND2_X1 U790 ( .A1(n777), .A2(n779), .ZN(n801) );
  NAND2_X1 U791 ( .A1(n802), .A2(n803), .ZN(n779) );
  NAND2_X1 U792 ( .A1(a_2_), .A2(b_4_), .ZN(n803) );
  XNOR2_X1 U793 ( .A(n804), .B(n805), .ZN(n777) );
  XOR2_X1 U794 ( .A(n590), .B(n806), .Z(n805) );
  OR2_X1 U795 ( .A1(n802), .A2(n646), .ZN(n778) );
  NAND2_X1 U796 ( .A1(n807), .A2(n808), .ZN(n802) );
  NAND2_X1 U797 ( .A1(n772), .A2(n809), .ZN(n808) );
  OR2_X1 U798 ( .A1(n775), .A2(n774), .ZN(n809) );
  XOR2_X1 U799 ( .A(n810), .B(n811), .Z(n772) );
  NAND2_X1 U800 ( .A1(n812), .A2(n813), .ZN(n810) );
  NAND2_X1 U801 ( .A1(n775), .A2(n774), .ZN(n807) );
  NAND2_X1 U802 ( .A1(n814), .A2(n815), .ZN(n774) );
  NAND2_X1 U803 ( .A1(n770), .A2(n816), .ZN(n815) );
  OR2_X1 U804 ( .A1(n561), .A2(n771), .ZN(n816) );
  XNOR2_X1 U805 ( .A(n817), .B(n818), .ZN(n770) );
  NOR2_X1 U806 ( .A1(n819), .A2(n820), .ZN(n818) );
  NOR2_X1 U807 ( .A1(n821), .A2(n822), .ZN(n819) );
  NOR2_X1 U808 ( .A1(n579), .A2(n550), .ZN(n822) );
  INV_X1 U809 ( .A(n823), .ZN(n821) );
  NAND2_X1 U810 ( .A1(n771), .A2(n561), .ZN(n814) );
  NAND2_X1 U811 ( .A1(b_4_), .A2(a_4_), .ZN(n561) );
  NOR2_X1 U812 ( .A1(n759), .A2(n824), .ZN(n771) );
  AND2_X1 U813 ( .A1(n756), .A2(n825), .ZN(n824) );
  NAND2_X1 U814 ( .A1(n762), .A2(n826), .ZN(n825) );
  NAND2_X1 U815 ( .A1(b_4_), .A2(a_5_), .ZN(n826) );
  AND2_X1 U816 ( .A1(n823), .A2(n827), .ZN(n756) );
  NAND2_X1 U817 ( .A1(n828), .A2(n829), .ZN(n827) );
  NAND2_X1 U818 ( .A1(b_3_), .A2(a_6_), .ZN(n828) );
  NOR2_X1 U819 ( .A1(n762), .A2(n550), .ZN(n759) );
  NAND2_X1 U820 ( .A1(n767), .A2(n768), .ZN(n762) );
  NOR2_X1 U821 ( .A1(n599), .A2(n532), .ZN(n768) );
  INV_X1 U822 ( .A(b_4_), .ZN(n599) );
  NOR2_X1 U823 ( .A1(n579), .A2(n664), .ZN(n767) );
  NAND2_X1 U824 ( .A1(a_3_), .A2(b_4_), .ZN(n775) );
  XNOR2_X1 U825 ( .A(n830), .B(n831), .ZN(n685) );
  XOR2_X1 U826 ( .A(n832), .B(n833), .Z(n831) );
  NAND2_X1 U827 ( .A1(n834), .A2(n835), .ZN(n512) );
  NAND2_X1 U828 ( .A1(n621), .A2(n836), .ZN(n835) );
  NAND2_X1 U829 ( .A1(n837), .A2(n621), .ZN(n511) );
  XNOR2_X1 U830 ( .A(n838), .B(n839), .ZN(n621) );
  NAND2_X1 U831 ( .A1(n840), .A2(n841), .ZN(n838) );
  NOR2_X1 U832 ( .A1(n622), .A2(n834), .ZN(n837) );
  XNOR2_X1 U833 ( .A(n612), .B(n613), .ZN(n834) );
  INV_X1 U834 ( .A(n836), .ZN(n622) );
  NAND2_X1 U835 ( .A1(n842), .A2(n843), .ZN(n836) );
  NAND2_X1 U836 ( .A1(n844), .A2(a_0_), .ZN(n843) );
  NOR2_X1 U837 ( .A1(n845), .A2(n579), .ZN(n844) );
  NOR2_X1 U838 ( .A1(n787), .A2(n785), .ZN(n845) );
  NAND2_X1 U839 ( .A1(n787), .A2(n785), .ZN(n842) );
  XOR2_X1 U840 ( .A(n846), .B(n847), .Z(n785) );
  XOR2_X1 U841 ( .A(n848), .B(n849), .Z(n846) );
  AND2_X1 U842 ( .A1(n850), .A2(n851), .ZN(n787) );
  NAND2_X1 U843 ( .A1(n832), .A2(n852), .ZN(n851) );
  NAND2_X1 U844 ( .A1(n833), .A2(n830), .ZN(n852) );
  AND2_X1 U845 ( .A1(n853), .A2(n854), .ZN(n832) );
  NAND2_X1 U846 ( .A1(n855), .A2(a_2_), .ZN(n854) );
  NOR2_X1 U847 ( .A1(n856), .A2(n579), .ZN(n855) );
  NOR2_X1 U848 ( .A1(n800), .A2(n798), .ZN(n856) );
  NAND2_X1 U849 ( .A1(n800), .A2(n798), .ZN(n853) );
  XOR2_X1 U850 ( .A(n857), .B(n858), .Z(n798) );
  XNOR2_X1 U851 ( .A(n859), .B(n860), .ZN(n857) );
  NAND2_X1 U852 ( .A1(a_3_), .A2(b_2_), .ZN(n859) );
  AND2_X1 U853 ( .A1(n861), .A2(n862), .ZN(n800) );
  NAND2_X1 U854 ( .A1(n863), .A2(n864), .ZN(n862) );
  NAND2_X1 U855 ( .A1(n573), .A2(n804), .ZN(n864) );
  INV_X1 U856 ( .A(n806), .ZN(n863) );
  NAND2_X1 U857 ( .A1(n812), .A2(n865), .ZN(n806) );
  NAND2_X1 U858 ( .A1(n811), .A2(n813), .ZN(n865) );
  NAND2_X1 U859 ( .A1(n866), .A2(n867), .ZN(n813) );
  NAND2_X1 U860 ( .A1(a_4_), .A2(b_3_), .ZN(n867) );
  XNOR2_X1 U861 ( .A(n868), .B(n869), .ZN(n811) );
  NAND2_X1 U862 ( .A1(n870), .A2(n871), .ZN(n868) );
  OR2_X1 U863 ( .A1(n600), .A2(n866), .ZN(n812) );
  NOR2_X1 U864 ( .A1(n820), .A2(n872), .ZN(n866) );
  AND2_X1 U865 ( .A1(n817), .A2(n873), .ZN(n872) );
  NAND2_X1 U866 ( .A1(n823), .A2(n874), .ZN(n873) );
  NAND2_X1 U867 ( .A1(a_5_), .A2(b_3_), .ZN(n874) );
  XOR2_X1 U868 ( .A(n875), .B(n876), .Z(n817) );
  NOR2_X1 U869 ( .A1(n823), .A2(n550), .ZN(n820) );
  NAND2_X1 U870 ( .A1(n877), .A2(b_3_), .ZN(n823) );
  NOR2_X1 U871 ( .A1(n829), .A2(n532), .ZN(n877) );
  NAND2_X1 U872 ( .A1(b_2_), .A2(a_7_), .ZN(n829) );
  OR2_X1 U873 ( .A1(n804), .A2(n573), .ZN(n861) );
  INV_X1 U874 ( .A(n590), .ZN(n573) );
  NAND2_X1 U875 ( .A1(a_3_), .A2(b_3_), .ZN(n590) );
  XNOR2_X1 U876 ( .A(n878), .B(n879), .ZN(n804) );
  NAND2_X1 U877 ( .A1(n880), .A2(n881), .ZN(n878) );
  OR2_X1 U878 ( .A1(n830), .A2(n833), .ZN(n850) );
  NOR2_X1 U879 ( .A1(n466), .A2(n579), .ZN(n833) );
  INV_X1 U880 ( .A(b_3_), .ZN(n579) );
  XOR2_X1 U881 ( .A(n882), .B(n883), .Z(n830) );
  XOR2_X1 U882 ( .A(n884), .B(n476), .Z(n882) );
  NAND2_X1 U883 ( .A1(n885), .A2(n886), .ZN(n516) );
  OR2_X1 U884 ( .A1(n613), .A2(n612), .ZN(n886) );
  AND2_X1 U885 ( .A1(n840), .A2(n887), .ZN(n612) );
  NAND2_X1 U886 ( .A1(n839), .A2(n841), .ZN(n887) );
  NAND2_X1 U887 ( .A1(n888), .A2(n889), .ZN(n841) );
  NAND2_X1 U888 ( .A1(a_0_), .A2(b_2_), .ZN(n889) );
  INV_X1 U889 ( .A(n890), .ZN(n888) );
  XOR2_X1 U890 ( .A(n891), .B(n892), .Z(n839) );
  XNOR2_X1 U891 ( .A(n456), .B(n893), .ZN(n892) );
  NAND2_X1 U892 ( .A1(b_0_), .A2(a_2_), .ZN(n891) );
  NAND2_X1 U893 ( .A1(a_0_), .A2(n890), .ZN(n840) );
  NAND2_X1 U894 ( .A1(n894), .A2(n895), .ZN(n890) );
  NAND2_X1 U895 ( .A1(n849), .A2(n896), .ZN(n895) );
  OR2_X1 U896 ( .A1(n848), .A2(n847), .ZN(n896) );
  NOR2_X1 U897 ( .A1(n466), .A2(n897), .ZN(n849) );
  NAND2_X1 U898 ( .A1(n847), .A2(n848), .ZN(n894) );
  NAND2_X1 U899 ( .A1(n898), .A2(n899), .ZN(n848) );
  NAND2_X1 U900 ( .A1(n476), .A2(n900), .ZN(n899) );
  OR2_X1 U901 ( .A1(n884), .A2(n883), .ZN(n900) );
  NOR2_X1 U902 ( .A1(n646), .A2(n897), .ZN(n476) );
  NAND2_X1 U903 ( .A1(n883), .A2(n884), .ZN(n898) );
  NAND2_X1 U904 ( .A1(n901), .A2(n902), .ZN(n884) );
  NAND2_X1 U905 ( .A1(n903), .A2(a_3_), .ZN(n902) );
  NOR2_X1 U906 ( .A1(n904), .A2(n897), .ZN(n903) );
  NOR2_X1 U907 ( .A1(n858), .A2(n860), .ZN(n904) );
  NAND2_X1 U908 ( .A1(n858), .A2(n860), .ZN(n901) );
  NAND2_X1 U909 ( .A1(n880), .A2(n905), .ZN(n860) );
  NAND2_X1 U910 ( .A1(n879), .A2(n881), .ZN(n905) );
  NAND2_X1 U911 ( .A1(n906), .A2(n907), .ZN(n881) );
  NAND2_X1 U912 ( .A1(a_4_), .A2(b_2_), .ZN(n907) );
  INV_X1 U913 ( .A(n908), .ZN(n906) );
  XOR2_X1 U914 ( .A(n909), .B(n910), .Z(n879) );
  AND2_X1 U915 ( .A1(n911), .A2(n912), .ZN(n910) );
  NAND2_X1 U916 ( .A1(a_4_), .A2(n908), .ZN(n880) );
  NAND2_X1 U917 ( .A1(n870), .A2(n913), .ZN(n908) );
  NAND2_X1 U918 ( .A1(n869), .A2(n871), .ZN(n913) );
  NAND2_X1 U919 ( .A1(n914), .A2(n915), .ZN(n871) );
  NAND2_X1 U920 ( .A1(a_5_), .A2(b_2_), .ZN(n915) );
  AND2_X1 U921 ( .A1(n911), .A2(n916), .ZN(n869) );
  NAND2_X1 U922 ( .A1(n917), .A2(n918), .ZN(n916) );
  NAND2_X1 U923 ( .A1(b_0_), .A2(a_7_), .ZN(n918) );
  NAND2_X1 U924 ( .A1(b_1_), .A2(a_6_), .ZN(n917) );
  OR2_X1 U925 ( .A1(n914), .A2(n550), .ZN(n870) );
  NAND2_X1 U926 ( .A1(n875), .A2(n876), .ZN(n914) );
  NOR2_X1 U927 ( .A1(n532), .A2(n897), .ZN(n875) );
  INV_X1 U928 ( .A(b_2_), .ZN(n897) );
  INV_X1 U929 ( .A(a_6_), .ZN(n532) );
  XOR2_X1 U930 ( .A(n919), .B(n920), .Z(n858) );
  XOR2_X1 U931 ( .A(n921), .B(n922), .Z(n919) );
  XOR2_X1 U932 ( .A(n923), .B(n924), .Z(n883) );
  XNOR2_X1 U933 ( .A(n925), .B(n926), .ZN(n924) );
  NAND2_X1 U934 ( .A1(b_0_), .A2(a_4_), .ZN(n923) );
  XOR2_X1 U935 ( .A(n927), .B(n928), .Z(n847) );
  NOR2_X1 U936 ( .A1(n929), .A2(n930), .ZN(n928) );
  INV_X1 U937 ( .A(n931), .ZN(n930) );
  NOR2_X1 U938 ( .A1(n932), .A2(n933), .ZN(n929) );
  XNOR2_X1 U939 ( .A(n934), .B(n935), .ZN(n613) );
  NOR2_X1 U940 ( .A1(n936), .A2(n937), .ZN(n935) );
  INV_X1 U941 ( .A(n938), .ZN(n937) );
  NOR2_X1 U942 ( .A1(n939), .A2(n940), .ZN(n936) );
  XOR2_X1 U943 ( .A(n474), .B(n614), .Z(n885) );
  NAND2_X1 U944 ( .A1(b_0_), .A2(a_0_), .ZN(n474) );
  AND2_X1 U945 ( .A1(n614), .A2(a_0_), .ZN(n607) );
  NAND2_X1 U946 ( .A1(n938), .A2(n941), .ZN(n614) );
  NAND2_X1 U947 ( .A1(n942), .A2(n934), .ZN(n941) );
  NAND2_X1 U948 ( .A1(n943), .A2(n944), .ZN(n934) );
  NAND2_X1 U949 ( .A1(n945), .A2(b_0_), .ZN(n944) );
  NOR2_X1 U950 ( .A1(n946), .A2(n646), .ZN(n945) );
  NOR2_X1 U951 ( .A1(n456), .A2(n893), .ZN(n946) );
  NAND2_X1 U952 ( .A1(n456), .A2(n893), .ZN(n943) );
  NAND2_X1 U953 ( .A1(n931), .A2(n947), .ZN(n893) );
  NAND2_X1 U954 ( .A1(n948), .A2(n927), .ZN(n947) );
  NAND2_X1 U955 ( .A1(n949), .A2(n950), .ZN(n927) );
  NAND2_X1 U956 ( .A1(n951), .A2(b_0_), .ZN(n950) );
  NOR2_X1 U957 ( .A1(n952), .A2(n600), .ZN(n951) );
  NOR2_X1 U958 ( .A1(n926), .A2(n925), .ZN(n952) );
  NAND2_X1 U959 ( .A1(n926), .A2(n925), .ZN(n949) );
  NAND2_X1 U960 ( .A1(n953), .A2(n954), .ZN(n925) );
  NAND2_X1 U961 ( .A1(n920), .A2(n955), .ZN(n954) );
  OR2_X1 U962 ( .A1(n922), .A2(n921), .ZN(n955) );
  AND2_X1 U963 ( .A1(b_0_), .A2(a_5_), .ZN(n920) );
  NAND2_X1 U964 ( .A1(n921), .A2(n922), .ZN(n953) );
  NAND2_X1 U965 ( .A1(n956), .A2(n911), .ZN(n922) );
  NAND2_X1 U966 ( .A1(n912), .A2(n876), .ZN(n911) );
  NOR2_X1 U967 ( .A1(n957), .A2(n664), .ZN(n876) );
  INV_X1 U968 ( .A(a_7_), .ZN(n664) );
  NAND2_X1 U969 ( .A1(n909), .A2(n912), .ZN(n956) );
  AND2_X1 U970 ( .A1(b_0_), .A2(a_6_), .ZN(n912) );
  NOR2_X1 U971 ( .A1(n957), .A2(n550), .ZN(n909) );
  INV_X1 U972 ( .A(a_5_), .ZN(n550) );
  NOR2_X1 U973 ( .A1(n600), .A2(n957), .ZN(n921) );
  INV_X1 U974 ( .A(a_4_), .ZN(n600) );
  NOR2_X1 U975 ( .A1(n578), .A2(n957), .ZN(n926) );
  INV_X1 U976 ( .A(a_3_), .ZN(n578) );
  NAND2_X1 U977 ( .A1(n958), .A2(n646), .ZN(n948) );
  NAND2_X1 U978 ( .A1(n933), .A2(n932), .ZN(n931) );
  INV_X1 U979 ( .A(n958), .ZN(n932) );
  NAND2_X1 U980 ( .A1(b_0_), .A2(a_3_), .ZN(n958) );
  NOR2_X1 U981 ( .A1(n957), .A2(n646), .ZN(n933) );
  INV_X1 U982 ( .A(a_2_), .ZN(n646) );
  NOR2_X1 U983 ( .A1(n466), .A2(n957), .ZN(n456) );
  INV_X1 U984 ( .A(a_1_), .ZN(n466) );
  NAND2_X1 U985 ( .A1(n959), .A2(n693), .ZN(n942) );
  NAND2_X1 U986 ( .A1(n940), .A2(n939), .ZN(n938) );
  INV_X1 U987 ( .A(n959), .ZN(n939) );
  NAND2_X1 U988 ( .A1(b_0_), .A2(a_1_), .ZN(n959) );
  NOR2_X1 U989 ( .A1(n957), .A2(n693), .ZN(n940) );
  INV_X1 U990 ( .A(a_0_), .ZN(n693) );
  INV_X1 U991 ( .A(b_1_), .ZN(n957) );
endmodule

