module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n614_, new_n445_, new_n236_, new_n238_, new_n479_, new_n608_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n601_, new_n556_, new_n456_, new_n246_, new_n170_, new_n266_, new_n367_, new_n542_, new_n173_, new_n220_, new_n419_, new_n534_, new_n214_, new_n451_, new_n489_, new_n602_, new_n188_, new_n240_, new_n413_, new_n526_, new_n211_, new_n552_, new_n342_, new_n462_, new_n603_, new_n564_, new_n500_, new_n317_, new_n344_, new_n287_, new_n504_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n257_, new_n481_, new_n212_, new_n449_, new_n364_, new_n580_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n315_, new_n326_, new_n554_, new_n164_, new_n230_, new_n281_, new_n430_, new_n482_, new_n606_, new_n589_, new_n248_, new_n350_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n565_, new_n150_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n491_, new_n549_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n206_, new_n254_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n587_, new_n465_, new_n263_, new_n334_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n524_, new_n277_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n528_, new_n179_, new_n572_, new_n436_, new_n397_, new_n399_, new_n596_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n166_, new_n162_, new_n457_, new_n161_, new_n553_, new_n333_, new_n290_, new_n369_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n308_, new_n232_, new_n258_, new_n176_, new_n156_, new_n306_, new_n494_, new_n291_, new_n261_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n604_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n460_, new_n505_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n485_, new_n525_, new_n562_, new_n578_, new_n177_, new_n493_, new_n547_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n570_, new_n598_, new_n143_, new_n520_, new_n145_, new_n253_, new_n237_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n507_, new_n605_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n592_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n522_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n569_, new_n555_, new_n174_, new_n468_, new_n354_, new_n392_, new_n444_, new_n518_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n203_, new_n316_, new_n590_, new_n417_, new_n515_, new_n332_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n440_, new_n531_, new_n593_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n242_, new_n503_, new_n527_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n435_, new_n265_, new_n370_, new_n278_, new_n304_, new_n523_, new_n217_, new_n269_, new_n512_, new_n599_, new_n412_, new_n327_, new_n594_, new_n561_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n336_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n567_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n322_, new_n228_, new_n545_, new_n611_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n284_, new_n293_, new_n551_, new_n168_, new_n279_, new_n455_, new_n618_, new_n521_, new_n356_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n405_;

not g000 ( new_n138_, keyIn_0_41 );
xnor g001 ( new_n139_, N89, N93 );
xnor g002 ( new_n140_, N81, N85 );
xor g003 ( new_n141_, new_n139_, new_n140_ );
not g004 ( new_n142_, new_n141_ );
xnor g005 ( new_n143_, N73, N77 );
xnor g006 ( new_n144_, new_n143_, keyIn_0_6 );
xnor g007 ( new_n145_, N65, N69 );
nand g008 ( new_n146_, new_n145_, keyIn_0_5 );
or g009 ( new_n147_, new_n145_, keyIn_0_5 );
nand g010 ( new_n148_, new_n144_, new_n146_, new_n147_ );
not g011 ( new_n149_, keyIn_0_6 );
xnor g012 ( new_n150_, new_n143_, new_n149_ );
xnor g013 ( new_n151_, new_n145_, keyIn_0_5 );
nand g014 ( new_n152_, new_n150_, new_n151_ );
nand g015 ( new_n153_, new_n148_, new_n152_ );
nand g016 ( new_n154_, new_n153_, new_n142_ );
nand g017 ( new_n155_, new_n148_, new_n152_, new_n141_ );
nand g018 ( new_n156_, new_n154_, new_n155_ );
nand g019 ( new_n157_, N129, N137 );
nand g020 ( new_n158_, new_n156_, new_n157_ );
nand g021 ( new_n159_, new_n154_, N129, N137, new_n155_ );
nand g022 ( new_n160_, new_n158_, new_n159_ );
xnor g023 ( new_n161_, N33, N49 );
xnor g024 ( new_n162_, N1, N17 );
xnor g025 ( new_n163_, new_n161_, new_n162_ );
xnor g026 ( new_n164_, new_n160_, new_n163_ );
not g027 ( new_n165_, keyIn_0_36 );
xnor g028 ( new_n166_, N121, N125 );
or g029 ( new_n167_, new_n166_, keyIn_0_7 );
nand g030 ( new_n168_, new_n166_, keyIn_0_7 );
xnor g031 ( new_n169_, N113, N117 );
nand g032 ( new_n170_, new_n167_, new_n168_, new_n169_ );
xnor g033 ( new_n171_, new_n166_, keyIn_0_7 );
not g034 ( new_n172_, new_n169_ );
nand g035 ( new_n173_, new_n171_, new_n172_ );
nand g036 ( new_n174_, new_n173_, new_n170_ );
nand g037 ( new_n175_, new_n174_, keyIn_0_19 );
not g038 ( new_n176_, keyIn_0_19 );
nand g039 ( new_n177_, new_n173_, new_n176_, new_n170_ );
nand g040 ( new_n178_, new_n175_, new_n177_ );
not g041 ( new_n179_, keyIn_0_18 );
xor g042 ( new_n180_, N97, N101 );
xnor g043 ( new_n181_, N105, N109 );
nand g044 ( new_n182_, new_n180_, new_n181_ );
xnor g045 ( new_n183_, N97, N101 );
xor g046 ( new_n184_, N105, N109 );
nand g047 ( new_n185_, new_n184_, new_n183_ );
nand g048 ( new_n186_, new_n182_, new_n185_, new_n179_ );
nand g049 ( new_n187_, new_n182_, new_n185_ );
nand g050 ( new_n188_, new_n187_, keyIn_0_18 );
nand g051 ( new_n189_, new_n188_, new_n186_ );
nand g052 ( new_n190_, new_n178_, new_n189_ );
nand g053 ( new_n191_, new_n175_, new_n177_, new_n186_, new_n188_ );
nand g054 ( new_n192_, new_n190_, new_n191_ );
nand g055 ( new_n193_, new_n192_, keyIn_0_22 );
not g056 ( new_n194_, keyIn_0_22 );
nand g057 ( new_n195_, new_n190_, new_n194_, new_n191_ );
nand g058 ( new_n196_, new_n193_, new_n195_ );
nand g059 ( new_n197_, N130, N137 );
xor g060 ( new_n198_, new_n197_, keyIn_0_8 );
not g061 ( new_n199_, new_n198_ );
nand g062 ( new_n200_, new_n196_, new_n199_ );
nand g063 ( new_n201_, new_n193_, new_n195_, new_n198_ );
xor g064 ( new_n202_, N5, N21 );
xnor g065 ( new_n203_, new_n202_, keyIn_0_12 );
xor g066 ( new_n204_, N37, N53 );
xnor g067 ( new_n205_, new_n204_, keyIn_0_13 );
xor g068 ( new_n206_, new_n203_, new_n205_ );
nand g069 ( new_n207_, new_n200_, new_n201_, new_n206_ );
nand g070 ( new_n208_, new_n200_, new_n201_ );
not g071 ( new_n209_, new_n206_ );
nand g072 ( new_n210_, new_n208_, new_n209_ );
nand g073 ( new_n211_, new_n210_, new_n164_, new_n207_ );
not g074 ( new_n212_, keyIn_0_23 );
nand g075 ( new_n213_, new_n175_, new_n141_, new_n177_ );
nand g076 ( new_n214_, new_n178_, new_n142_ );
nand g077 ( new_n215_, N132, N137 );
xnor g078 ( new_n216_, new_n215_, keyIn_0_9 );
nand g079 ( new_n217_, new_n214_, new_n213_, new_n216_ );
nand g080 ( new_n218_, new_n214_, new_n213_ );
not g081 ( new_n219_, new_n216_ );
nand g082 ( new_n220_, new_n218_, new_n219_ );
nand g083 ( new_n221_, new_n220_, new_n217_ );
nand g084 ( new_n222_, new_n221_, new_n212_ );
nand g085 ( new_n223_, new_n220_, keyIn_0_23, new_n217_ );
xor g086 ( new_n224_, N13, N29 );
xnor g087 ( new_n225_, new_n224_, keyIn_0_14 );
xnor g088 ( new_n226_, N45, N61 );
xnor g089 ( new_n227_, new_n225_, new_n226_ );
nand g090 ( new_n228_, new_n222_, new_n223_, new_n227_ );
nand g091 ( new_n229_, new_n222_, new_n223_ );
not g092 ( new_n230_, new_n227_ );
nand g093 ( new_n231_, new_n229_, new_n230_ );
not g094 ( new_n232_, keyIn_0_26 );
nand g095 ( new_n233_, new_n148_, new_n152_, new_n188_, new_n186_ );
nand g096 ( new_n234_, new_n153_, new_n189_ );
nand g097 ( new_n235_, new_n234_, N131, N137, new_n233_ );
nand g098 ( new_n236_, new_n234_, new_n233_ );
nand g099 ( new_n237_, N131, N137 );
nand g100 ( new_n238_, new_n236_, new_n237_ );
nand g101 ( new_n239_, new_n238_, new_n235_ );
xnor g102 ( new_n240_, N41, N57 );
xnor g103 ( new_n241_, N9, N25 );
xor g104 ( new_n242_, new_n240_, new_n241_ );
not g105 ( new_n243_, new_n242_ );
nand g106 ( new_n244_, new_n239_, new_n243_ );
nand g107 ( new_n245_, new_n238_, new_n235_, new_n242_ );
nand g108 ( new_n246_, new_n244_, new_n245_ );
nand g109 ( new_n247_, new_n246_, keyIn_0_24 );
not g110 ( new_n248_, keyIn_0_24 );
nand g111 ( new_n249_, new_n244_, new_n248_, new_n245_ );
nand g112 ( new_n250_, new_n247_, new_n232_, new_n249_ );
nand g113 ( new_n251_, new_n247_, new_n249_ );
nand g114 ( new_n252_, new_n251_, keyIn_0_26 );
nand g115 ( new_n253_, new_n252_, new_n231_, new_n228_, new_n250_ );
nor g116 ( new_n254_, new_n253_, new_n211_ );
xnor g117 ( new_n255_, new_n254_, new_n165_ );
and g118 ( new_n256_, new_n231_, new_n228_ );
not g119 ( new_n257_, new_n164_ );
nand g120 ( new_n258_, new_n210_, new_n207_ );
nand g121 ( new_n259_, new_n258_, new_n257_, new_n251_ );
not g122 ( new_n260_, new_n251_ );
xnor g123 ( new_n261_, new_n164_, keyIn_0_25 );
nand g124 ( new_n262_, new_n261_, new_n207_, new_n210_, new_n260_ );
nand g125 ( new_n263_, new_n259_, new_n262_ );
nand g126 ( new_n264_, new_n263_, new_n256_ );
not g127 ( new_n265_, new_n258_ );
not g128 ( new_n266_, new_n256_ );
nand g129 ( new_n267_, new_n266_, new_n257_, new_n265_, new_n251_ );
nand g130 ( new_n268_, new_n264_, new_n267_ );
nor g131 ( new_n269_, new_n255_, new_n268_ );
not g132 ( new_n270_, keyIn_0_21 );
not g133 ( new_n271_, N37 );
not g134 ( new_n272_, N33 );
nand g135 ( new_n273_, new_n272_, keyIn_0_2 );
not g136 ( new_n274_, keyIn_0_2 );
nand g137 ( new_n275_, new_n274_, N33 );
nand g138 ( new_n276_, new_n273_, new_n275_ );
nand g139 ( new_n277_, new_n276_, new_n271_ );
nand g140 ( new_n278_, new_n273_, new_n275_, N37 );
nand g141 ( new_n279_, new_n277_, new_n278_ );
not g142 ( new_n280_, keyIn_0_3 );
xnor g143 ( new_n281_, N41, N45 );
nand g144 ( new_n282_, new_n281_, new_n280_ );
or g145 ( new_n283_, N41, N45 );
nand g146 ( new_n284_, N41, N45 );
nand g147 ( new_n285_, new_n283_, keyIn_0_3, new_n284_ );
nand g148 ( new_n286_, new_n282_, new_n285_ );
nand g149 ( new_n287_, new_n279_, new_n286_ );
nand g150 ( new_n288_, new_n277_, new_n282_, new_n278_, new_n285_ );
nand g151 ( new_n289_, new_n287_, new_n288_ );
nand g152 ( new_n290_, new_n289_, keyIn_0_17 );
not g153 ( new_n291_, keyIn_0_17 );
nand g154 ( new_n292_, new_n287_, new_n291_, new_n288_ );
nand g155 ( new_n293_, new_n290_, new_n292_ );
xnor g156 ( new_n294_, N1, N5 );
or g157 ( new_n295_, N9, N13 );
nand g158 ( new_n296_, N9, N13 );
nand g159 ( new_n297_, new_n294_, new_n295_, new_n296_ );
xor g160 ( new_n298_, N1, N5 );
nand g161 ( new_n299_, new_n295_, new_n296_ );
nand g162 ( new_n300_, new_n298_, new_n299_ );
nand g163 ( new_n301_, new_n300_, new_n297_ );
nand g164 ( new_n302_, new_n301_, keyIn_0_16 );
not g165 ( new_n303_, keyIn_0_16 );
nand g166 ( new_n304_, new_n300_, new_n303_, new_n297_ );
nand g167 ( new_n305_, new_n302_, new_n304_ );
not g168 ( new_n306_, new_n305_ );
nand g169 ( new_n307_, new_n293_, new_n306_ );
nand g170 ( new_n308_, new_n290_, new_n292_, new_n305_ );
nand g171 ( new_n309_, new_n307_, new_n308_ );
nand g172 ( new_n310_, new_n309_, new_n270_ );
nand g173 ( new_n311_, new_n307_, keyIn_0_21, new_n308_ );
nand g174 ( new_n312_, new_n310_, new_n311_ );
nand g175 ( new_n313_, N135, N137 );
xor g176 ( new_n314_, new_n313_, keyIn_0_10 );
not g177 ( new_n315_, new_n314_ );
nand g178 ( new_n316_, new_n312_, new_n315_ );
nand g179 ( new_n317_, new_n310_, new_n311_, new_n314_ );
nand g180 ( new_n318_, new_n316_, new_n317_ );
xor g181 ( new_n319_, N105, N121 );
xnor g182 ( new_n320_, N73, N89 );
xnor g183 ( new_n321_, new_n319_, new_n320_ );
xnor g184 ( new_n322_, new_n321_, keyIn_0_20 );
not g185 ( new_n323_, new_n322_ );
nand g186 ( new_n324_, new_n318_, new_n323_ );
nand g187 ( new_n325_, new_n316_, new_n317_, new_n322_ );
nand g188 ( new_n326_, new_n324_, new_n325_ );
not g189 ( new_n327_, new_n326_ );
nor g190 ( new_n328_, new_n269_, new_n327_ );
not g191 ( new_n329_, keyIn_0_4 );
xnor g192 ( new_n330_, N57, N61 );
xnor g193 ( new_n331_, new_n330_, new_n329_ );
xnor g194 ( new_n332_, N49, N53 );
nor g195 ( new_n333_, new_n331_, new_n332_ );
and g196 ( new_n334_, new_n331_, new_n332_ );
nor g197 ( new_n335_, new_n334_, new_n333_ );
nand g198 ( new_n336_, new_n293_, new_n335_ );
xnor g199 ( new_n337_, new_n331_, new_n332_ );
nand g200 ( new_n338_, new_n337_, new_n290_, new_n292_ );
nand g201 ( new_n339_, new_n336_, new_n338_ );
nand g202 ( new_n340_, N134, N137 );
nand g203 ( new_n341_, new_n339_, new_n340_ );
nand g204 ( new_n342_, new_n336_, N134, N137, new_n338_ );
nand g205 ( new_n343_, new_n341_, new_n342_ );
xnor g206 ( new_n344_, N101, N117 );
xnor g207 ( new_n345_, N69, N85 );
xor g208 ( new_n346_, new_n344_, new_n345_ );
not g209 ( new_n347_, new_n346_ );
nand g210 ( new_n348_, new_n343_, new_n347_ );
nand g211 ( new_n349_, new_n341_, new_n342_, new_n346_ );
not g212 ( new_n350_, keyIn_0_0 );
or g213 ( new_n351_, N17, N21 );
nand g214 ( new_n352_, N17, N21 );
nand g215 ( new_n353_, new_n351_, new_n350_, new_n352_ );
nand g216 ( new_n354_, new_n351_, new_n352_ );
nand g217 ( new_n355_, new_n354_, keyIn_0_0 );
not g218 ( new_n356_, keyIn_0_1 );
or g219 ( new_n357_, N25, N29 );
nand g220 ( new_n358_, N25, N29 );
nand g221 ( new_n359_, new_n357_, new_n356_, new_n358_ );
nand g222 ( new_n360_, new_n357_, new_n358_ );
nand g223 ( new_n361_, new_n360_, keyIn_0_1 );
nand g224 ( new_n362_, new_n355_, new_n361_, new_n353_, new_n359_ );
nand g225 ( new_n363_, new_n355_, new_n353_ );
nand g226 ( new_n364_, new_n361_, new_n359_ );
nand g227 ( new_n365_, new_n363_, new_n364_ );
nand g228 ( new_n366_, new_n305_, new_n362_, new_n365_ );
nand g229 ( new_n367_, new_n365_, new_n362_ );
nand g230 ( new_n368_, new_n367_, new_n302_, new_n304_ );
nand g231 ( new_n369_, new_n366_, new_n368_ );
nand g232 ( new_n370_, N133, N137 );
not g233 ( new_n371_, new_n370_ );
nand g234 ( new_n372_, new_n369_, new_n371_ );
nand g235 ( new_n373_, new_n366_, new_n368_, new_n370_ );
xnor g236 ( new_n374_, N97, N113 );
xnor g237 ( new_n375_, new_n374_, keyIn_0_15 );
xor g238 ( new_n376_, N65, N81 );
xnor g239 ( new_n377_, new_n375_, new_n376_ );
not g240 ( new_n378_, new_n377_ );
nand g241 ( new_n379_, new_n372_, new_n373_, new_n378_ );
nand g242 ( new_n380_, new_n372_, new_n373_ );
nand g243 ( new_n381_, new_n380_, new_n377_ );
nand g244 ( new_n382_, new_n381_, new_n379_ );
nand g245 ( new_n383_, new_n348_, new_n349_, new_n382_ );
nand g246 ( new_n384_, new_n337_, new_n362_, new_n365_ );
nand g247 ( new_n385_, new_n335_, new_n367_ );
nand g248 ( new_n386_, new_n384_, new_n385_ );
nand g249 ( new_n387_, N136, N137 );
xnor g250 ( new_n388_, new_n387_, keyIn_0_11 );
nand g251 ( new_n389_, new_n386_, new_n388_ );
not g252 ( new_n390_, new_n388_ );
nand g253 ( new_n391_, new_n384_, new_n385_, new_n390_ );
xnor g254 ( new_n392_, N109, N125 );
xnor g255 ( new_n393_, N77, N93 );
xor g256 ( new_n394_, new_n392_, new_n393_ );
not g257 ( new_n395_, new_n394_ );
nand g258 ( new_n396_, new_n389_, new_n391_, new_n395_ );
nand g259 ( new_n397_, new_n389_, new_n391_ );
nand g260 ( new_n398_, new_n397_, new_n394_ );
nand g261 ( new_n399_, new_n398_, new_n396_ );
nor g262 ( new_n400_, new_n383_, new_n399_ );
nand g263 ( new_n401_, new_n328_, new_n164_, new_n400_ );
xnor g264 ( new_n402_, new_n401_, new_n138_ );
xnor g265 ( N724, new_n402_, N1 );
nand g266 ( new_n404_, new_n328_, new_n258_, new_n400_ );
xnor g267 ( new_n405_, new_n404_, keyIn_0_42 );
xnor g268 ( N725, new_n405_, N5 );
and g269 ( new_n407_, new_n328_, new_n400_ );
nand g270 ( new_n408_, new_n407_, new_n260_ );
xnor g271 ( N726, new_n408_, N9 );
nand g272 ( new_n410_, new_n407_, new_n266_ );
xnor g273 ( N727, new_n410_, N13 );
and g274 ( new_n412_, new_n210_, new_n164_, new_n207_ );
and g275 ( new_n413_, new_n252_, new_n250_ );
nand g276 ( new_n414_, new_n413_, new_n412_, new_n256_ );
nand g277 ( new_n415_, new_n414_, new_n165_ );
nand g278 ( new_n416_, new_n254_, keyIn_0_36 );
nand g279 ( new_n417_, new_n415_, new_n416_ );
nand g280 ( new_n418_, new_n417_, new_n264_, new_n267_ );
not g281 ( new_n419_, new_n399_ );
nor g282 ( new_n420_, new_n326_, new_n383_, new_n419_ );
and g283 ( new_n421_, new_n418_, new_n420_ );
nand g284 ( new_n422_, new_n421_, new_n164_ );
xnor g285 ( new_n423_, new_n422_, N17 );
xnor g286 ( N728, new_n423_, keyIn_0_54 );
nand g287 ( new_n425_, new_n421_, new_n258_ );
xnor g288 ( new_n426_, new_n425_, N21 );
xnor g289 ( N729, new_n426_, keyIn_0_55 );
nand g290 ( new_n428_, new_n421_, new_n260_ );
xnor g291 ( N730, new_n428_, N25 );
not g292 ( new_n430_, keyIn_0_43 );
nand g293 ( new_n431_, new_n421_, new_n266_ );
xnor g294 ( new_n432_, new_n431_, new_n430_ );
xnor g295 ( N731, new_n432_, N29 );
nand g296 ( new_n434_, new_n348_, new_n349_ );
not g297 ( new_n435_, new_n434_ );
nor g298 ( new_n436_, new_n435_, new_n382_, new_n399_ );
nand g299 ( new_n437_, new_n328_, new_n164_, new_n436_ );
xnor g300 ( new_n438_, new_n437_, N33 );
xnor g301 ( N732, new_n438_, keyIn_0_56 );
nand g302 ( new_n440_, new_n328_, new_n258_, new_n436_ );
xnor g303 ( new_n441_, new_n440_, new_n271_ );
xnor g304 ( N733, new_n441_, keyIn_0_57 );
not g305 ( new_n443_, keyIn_0_44 );
nand g306 ( new_n444_, new_n328_, new_n260_, new_n436_ );
xnor g307 ( new_n445_, new_n444_, new_n443_ );
xnor g308 ( N734, new_n445_, N41 );
nand g309 ( new_n447_, new_n328_, keyIn_0_45, new_n266_, new_n436_ );
not g310 ( new_n448_, keyIn_0_45 );
nand g311 ( new_n449_, new_n418_, new_n266_, new_n326_, new_n436_ );
nand g312 ( new_n450_, new_n449_, new_n448_ );
nand g313 ( new_n451_, new_n447_, new_n450_ );
nand g314 ( new_n452_, new_n451_, N45 );
not g315 ( new_n453_, N45 );
nand g316 ( new_n454_, new_n447_, new_n453_, new_n450_ );
nand g317 ( new_n455_, new_n452_, new_n454_ );
nand g318 ( new_n456_, new_n455_, keyIn_0_58 );
not g319 ( new_n457_, keyIn_0_58 );
nand g320 ( new_n458_, new_n452_, new_n457_, new_n454_ );
nand g321 ( N735, new_n456_, new_n458_ );
not g322 ( new_n460_, keyIn_0_39 );
xor g323 ( new_n461_, new_n326_, keyIn_0_27 );
nor g324 ( new_n462_, new_n461_, new_n435_, new_n382_, new_n419_ );
nand g325 ( new_n463_, new_n418_, new_n462_ );
nand g326 ( new_n464_, new_n463_, new_n460_ );
nand g327 ( new_n465_, new_n418_, keyIn_0_39, new_n462_ );
nand g328 ( new_n466_, new_n464_, new_n465_ );
nand g329 ( new_n467_, new_n466_, new_n164_ );
nand g330 ( new_n468_, new_n467_, N49 );
not g331 ( new_n469_, N49 );
nand g332 ( new_n470_, new_n466_, new_n469_, new_n164_ );
nand g333 ( new_n471_, new_n468_, new_n470_ );
nand g334 ( new_n472_, new_n471_, keyIn_0_59 );
not g335 ( new_n473_, keyIn_0_59 );
nand g336 ( new_n474_, new_n468_, new_n473_, new_n470_ );
nand g337 ( N736, new_n472_, new_n474_ );
nand g338 ( new_n476_, new_n466_, new_n258_ );
nand g339 ( new_n477_, new_n476_, keyIn_0_46 );
not g340 ( new_n478_, keyIn_0_46 );
nand g341 ( new_n479_, new_n466_, new_n478_, new_n258_ );
nand g342 ( new_n480_, new_n477_, new_n479_ );
nand g343 ( new_n481_, new_n480_, N53 );
not g344 ( new_n482_, N53 );
nand g345 ( new_n483_, new_n477_, new_n482_, new_n479_ );
nand g346 ( N737, new_n481_, new_n483_ );
nand g347 ( new_n485_, new_n466_, new_n260_ );
xnor g348 ( N738, new_n485_, N57 );
nand g349 ( new_n487_, new_n466_, new_n266_ );
xnor g350 ( N739, new_n487_, N61 );
not g351 ( new_n489_, N65 );
not g352 ( new_n490_, keyIn_0_37 );
not g353 ( new_n491_, keyIn_0_31 );
nand g354 ( new_n492_, new_n324_, new_n491_, new_n325_ );
nand g355 ( new_n493_, new_n326_, keyIn_0_31 );
nand g356 ( new_n494_, new_n493_, new_n490_, new_n436_, new_n492_ );
nand g357 ( new_n495_, new_n493_, new_n436_, new_n492_ );
nand g358 ( new_n496_, new_n495_, keyIn_0_37 );
not g359 ( new_n497_, keyIn_0_32 );
nand g360 ( new_n498_, new_n324_, new_n497_, new_n325_ );
nand g361 ( new_n499_, new_n326_, keyIn_0_32 );
not g362 ( new_n500_, keyIn_0_33 );
nand g363 ( new_n501_, new_n399_, new_n500_ );
nand g364 ( new_n502_, new_n398_, keyIn_0_33, new_n396_ );
nand g365 ( new_n503_, new_n501_, new_n502_ );
nor g366 ( new_n504_, new_n503_, new_n383_ );
nand g367 ( new_n505_, new_n499_, new_n498_, new_n504_ );
nand g368 ( new_n506_, new_n434_, keyIn_0_28 );
not g369 ( new_n507_, keyIn_0_28 );
nand g370 ( new_n508_, new_n348_, new_n507_, new_n349_ );
nand g371 ( new_n509_, new_n506_, new_n508_ );
nor g372 ( new_n510_, new_n419_, new_n382_ );
nand g373 ( new_n511_, new_n509_, new_n324_, new_n325_, new_n510_ );
not g374 ( new_n512_, keyIn_0_30 );
xnor g375 ( new_n513_, new_n399_, new_n512_ );
nand g376 ( new_n514_, new_n382_, keyIn_0_29 );
not g377 ( new_n515_, keyIn_0_29 );
nand g378 ( new_n516_, new_n381_, new_n515_, new_n379_ );
and g379 ( new_n517_, new_n348_, new_n514_, new_n349_, new_n516_ );
nand g380 ( new_n518_, new_n326_, new_n513_, new_n517_ );
and g381 ( new_n519_, new_n511_, new_n518_ );
nand g382 ( new_n520_, new_n496_, new_n519_, new_n494_, new_n505_ );
nand g383 ( new_n521_, new_n520_, keyIn_0_38 );
not g384 ( new_n522_, keyIn_0_38 );
and g385 ( new_n523_, new_n505_, new_n511_, new_n518_ );
nand g386 ( new_n524_, new_n523_, new_n522_, new_n494_, new_n496_ );
nand g387 ( new_n525_, new_n256_, new_n260_ );
nor g388 ( new_n526_, new_n525_, new_n211_ );
nand g389 ( new_n527_, new_n521_, new_n524_, new_n526_ );
nand g390 ( new_n528_, new_n527_, keyIn_0_40 );
not g391 ( new_n529_, keyIn_0_40 );
nand g392 ( new_n530_, new_n521_, new_n524_, new_n529_, new_n526_ );
nand g393 ( new_n531_, new_n528_, new_n530_ );
nand g394 ( new_n532_, new_n531_, new_n382_ );
nand g395 ( new_n533_, new_n532_, keyIn_0_47 );
not g396 ( new_n534_, keyIn_0_47 );
nand g397 ( new_n535_, new_n531_, new_n534_, new_n382_ );
nand g398 ( new_n536_, new_n533_, new_n535_ );
nand g399 ( new_n537_, new_n536_, new_n489_ );
nand g400 ( new_n538_, new_n533_, N65, new_n535_ );
nand g401 ( N740, new_n537_, new_n538_ );
not g402 ( new_n540_, N69 );
nand g403 ( new_n541_, new_n531_, new_n434_ );
nand g404 ( new_n542_, new_n541_, keyIn_0_48 );
not g405 ( new_n543_, keyIn_0_48 );
nand g406 ( new_n544_, new_n531_, new_n543_, new_n434_ );
nand g407 ( new_n545_, new_n542_, new_n544_ );
nand g408 ( new_n546_, new_n545_, new_n540_ );
nand g409 ( new_n547_, new_n542_, N69, new_n544_ );
nand g410 ( N741, new_n546_, new_n547_ );
nand g411 ( new_n549_, new_n531_, new_n326_ );
xnor g412 ( N742, new_n549_, N73 );
nand g413 ( new_n551_, new_n531_, new_n399_ );
nand g414 ( new_n552_, new_n551_, N77 );
not g415 ( new_n553_, N77 );
nand g416 ( new_n554_, new_n531_, new_n553_, new_n399_ );
nand g417 ( new_n555_, new_n552_, new_n554_ );
nand g418 ( new_n556_, new_n555_, keyIn_0_60 );
not g419 ( new_n557_, keyIn_0_60 );
nand g420 ( new_n558_, new_n552_, new_n557_, new_n554_ );
nand g421 ( N743, new_n556_, new_n558_ );
not g422 ( new_n560_, new_n382_ );
and g423 ( new_n561_, new_n521_, new_n524_ );
nor g424 ( new_n562_, new_n258_, keyIn_0_34 );
and g425 ( new_n563_, new_n258_, keyIn_0_34 );
nand g426 ( new_n564_, new_n251_, new_n164_ );
nor g427 ( new_n565_, new_n563_, new_n562_, new_n256_, new_n564_ );
nand g428 ( new_n566_, new_n561_, new_n565_ );
nor g429 ( new_n567_, new_n566_, new_n560_ );
xor g430 ( N744, new_n567_, N81 );
nand g431 ( new_n569_, new_n561_, new_n434_, new_n565_ );
xnor g432 ( new_n570_, new_n569_, keyIn_0_49 );
xnor g433 ( N745, new_n570_, N85 );
nand g434 ( new_n572_, new_n561_, new_n326_, new_n565_ );
xnor g435 ( new_n573_, new_n572_, N89 );
xnor g436 ( N746, new_n573_, keyIn_0_61 );
nor g437 ( new_n575_, new_n566_, new_n419_ );
xor g438 ( N747, new_n575_, N93 );
xor g439 ( new_n577_, new_n164_, keyIn_0_35 );
nor g440 ( new_n578_, new_n525_, new_n265_, new_n577_ );
nand g441 ( new_n579_, new_n561_, new_n578_ );
nor g442 ( new_n580_, new_n579_, new_n560_ );
xor g443 ( N748, new_n580_, N97 );
nand g444 ( new_n582_, new_n561_, new_n434_, new_n578_ );
xnor g445 ( new_n583_, new_n582_, keyIn_0_50 );
xnor g446 ( N749, new_n583_, N101 );
nor g447 ( new_n585_, new_n579_, new_n327_ );
xor g448 ( N750, new_n585_, N105 );
nor g449 ( new_n587_, new_n579_, new_n419_ );
xor g450 ( N751, new_n587_, N109 );
nor g451 ( new_n589_, new_n259_, new_n256_ );
nand g452 ( new_n590_, new_n561_, new_n382_, new_n589_ );
xnor g453 ( N752, new_n590_, N113 );
not g454 ( new_n592_, N117 );
nand g455 ( new_n593_, new_n561_, new_n434_, new_n589_ );
xnor g456 ( new_n594_, new_n593_, keyIn_0_51 );
xnor g457 ( N753, new_n594_, new_n592_ );
not g458 ( new_n596_, keyIn_0_62 );
not g459 ( new_n597_, N121 );
nand g460 ( new_n598_, new_n521_, new_n524_, new_n326_, new_n589_ );
or g461 ( new_n599_, new_n598_, keyIn_0_52 );
nand g462 ( new_n600_, new_n598_, keyIn_0_52 );
nand g463 ( new_n601_, new_n599_, new_n600_ );
nand g464 ( new_n602_, new_n601_, new_n597_ );
nand g465 ( new_n603_, new_n599_, N121, new_n600_ );
nand g466 ( new_n604_, new_n602_, new_n603_ );
nand g467 ( new_n605_, new_n604_, new_n596_ );
nand g468 ( new_n606_, new_n602_, keyIn_0_62, new_n603_ );
nand g469 ( N754, new_n605_, new_n606_ );
not g470 ( new_n608_, keyIn_0_63 );
nand g471 ( new_n609_, new_n521_, new_n524_, new_n399_, new_n589_ );
or g472 ( new_n610_, new_n609_, keyIn_0_53 );
nand g473 ( new_n611_, new_n609_, keyIn_0_53 );
nand g474 ( new_n612_, new_n610_, new_n611_ );
nand g475 ( new_n613_, new_n612_, N125 );
not g476 ( new_n614_, N125 );
nand g477 ( new_n615_, new_n610_, new_n614_, new_n611_ );
nand g478 ( new_n616_, new_n613_, new_n615_ );
nand g479 ( new_n617_, new_n616_, new_n608_ );
nand g480 ( new_n618_, new_n613_, keyIn_0_63, new_n615_ );
nand g481 ( N755, new_n617_, new_n618_ );
endmodule