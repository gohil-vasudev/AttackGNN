module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n691_, new_n456_, new_n1024_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n1124_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n1109_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n861_, new_n1091_, new_n310_, new_n144_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n1096_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n802_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n138_, N69 );
and g001 ( new_n139_, new_n138_, N65 );
not g002 ( new_n140_, N65 );
and g003 ( new_n141_, new_n140_, N69 );
or g004 ( new_n142_, new_n139_, new_n141_ );
not g005 ( new_n143_, N73 );
not g006 ( new_n144_, N77 );
and g007 ( new_n145_, new_n143_, new_n144_ );
and g008 ( new_n146_, N73, N77 );
or g009 ( new_n147_, new_n145_, new_n146_ );
and g010 ( new_n148_, new_n142_, new_n147_ );
not g011 ( new_n149_, new_n148_ );
or g012 ( new_n150_, new_n142_, new_n147_ );
and g013 ( new_n151_, new_n149_, new_n150_ );
not g014 ( new_n152_, new_n151_ );
not g015 ( new_n153_, N85 );
and g016 ( new_n154_, new_n153_, N81 );
not g017 ( new_n155_, N81 );
and g018 ( new_n156_, new_n155_, N85 );
or g019 ( new_n157_, new_n154_, new_n156_ );
not g020 ( new_n158_, N89 );
not g021 ( new_n159_, N93 );
and g022 ( new_n160_, new_n158_, new_n159_ );
and g023 ( new_n161_, N89, N93 );
or g024 ( new_n162_, new_n160_, new_n161_ );
and g025 ( new_n163_, new_n157_, new_n162_ );
not g026 ( new_n164_, new_n163_ );
or g027 ( new_n165_, new_n157_, new_n162_ );
and g028 ( new_n166_, new_n164_, new_n165_ );
and g029 ( new_n167_, new_n152_, new_n166_ );
not g030 ( new_n168_, new_n166_ );
and g031 ( new_n169_, new_n168_, new_n151_ );
or g032 ( new_n170_, new_n167_, new_n169_ );
and g033 ( new_n171_, N129, N137 );
not g034 ( new_n172_, new_n171_ );
and g035 ( new_n173_, new_n170_, new_n172_ );
not g036 ( new_n174_, new_n173_ );
or g037 ( new_n175_, new_n170_, new_n172_ );
and g038 ( new_n176_, new_n174_, new_n175_ );
not g039 ( new_n177_, new_n176_ );
not g040 ( new_n178_, N17 );
and g041 ( new_n179_, new_n178_, N1 );
not g042 ( new_n180_, N1 );
and g043 ( new_n181_, new_n180_, N17 );
or g044 ( new_n182_, new_n179_, new_n181_ );
not g045 ( new_n183_, N33 );
not g046 ( new_n184_, N49 );
and g047 ( new_n185_, new_n183_, new_n184_ );
and g048 ( new_n186_, N33, N49 );
or g049 ( new_n187_, new_n185_, new_n186_ );
and g050 ( new_n188_, new_n182_, new_n187_ );
not g051 ( new_n189_, new_n188_ );
or g052 ( new_n190_, new_n182_, new_n187_ );
and g053 ( new_n191_, new_n189_, new_n190_ );
not g054 ( new_n192_, new_n191_ );
and g055 ( new_n193_, new_n177_, new_n192_ );
and g056 ( new_n194_, new_n176_, new_n191_ );
or g057 ( new_n195_, new_n193_, new_n194_ );
not g058 ( new_n196_, new_n195_ );
not g059 ( new_n197_, keyIn_0_22 );
not g060 ( new_n198_, keyIn_0_13 );
not g061 ( new_n199_, N21 );
and g062 ( new_n200_, new_n178_, new_n199_ );
and g063 ( new_n201_, N17, N21 );
or g064 ( new_n202_, new_n200_, new_n201_ );
and g065 ( new_n203_, new_n202_, keyIn_0_2 );
not g066 ( new_n204_, keyIn_0_2 );
or g067 ( new_n205_, N17, N21 );
not g068 ( new_n206_, new_n201_ );
and g069 ( new_n207_, new_n206_, new_n205_ );
and g070 ( new_n208_, new_n207_, new_n204_ );
or g071 ( new_n209_, new_n203_, new_n208_ );
not g072 ( new_n210_, N25 );
not g073 ( new_n211_, N29 );
and g074 ( new_n212_, new_n210_, new_n211_ );
and g075 ( new_n213_, N25, N29 );
or g076 ( new_n214_, new_n212_, new_n213_ );
and g077 ( new_n215_, new_n214_, keyIn_0_3 );
not g078 ( new_n216_, keyIn_0_3 );
or g079 ( new_n217_, N25, N29 );
not g080 ( new_n218_, new_n213_ );
and g081 ( new_n219_, new_n218_, new_n217_ );
and g082 ( new_n220_, new_n219_, new_n216_ );
or g083 ( new_n221_, new_n215_, new_n220_ );
or g084 ( new_n222_, new_n209_, new_n221_ );
or g085 ( new_n223_, new_n207_, new_n204_ );
or g086 ( new_n224_, new_n202_, keyIn_0_2 );
and g087 ( new_n225_, new_n224_, new_n223_ );
or g088 ( new_n226_, new_n219_, new_n216_ );
or g089 ( new_n227_, new_n214_, keyIn_0_3 );
and g090 ( new_n228_, new_n227_, new_n226_ );
or g091 ( new_n229_, new_n225_, new_n228_ );
and g092 ( new_n230_, new_n222_, new_n229_ );
and g093 ( new_n231_, new_n230_, new_n198_ );
and g094 ( new_n232_, new_n225_, new_n228_ );
and g095 ( new_n233_, new_n209_, new_n221_ );
or g096 ( new_n234_, new_n233_, new_n232_ );
and g097 ( new_n235_, new_n234_, keyIn_0_13 );
or g098 ( new_n236_, new_n231_, new_n235_ );
not g099 ( new_n237_, N9 );
not g100 ( new_n238_, N13 );
and g101 ( new_n239_, new_n237_, new_n238_ );
and g102 ( new_n240_, N9, N13 );
or g103 ( new_n241_, new_n239_, new_n240_ );
and g104 ( new_n242_, new_n241_, keyIn_0_1 );
not g105 ( new_n243_, keyIn_0_1 );
or g106 ( new_n244_, N9, N13 );
not g107 ( new_n245_, new_n240_ );
and g108 ( new_n246_, new_n245_, new_n244_ );
and g109 ( new_n247_, new_n246_, new_n243_ );
or g110 ( new_n248_, new_n242_, new_n247_ );
not g111 ( new_n249_, keyIn_0_0 );
not g112 ( new_n250_, N5 );
and g113 ( new_n251_, new_n180_, new_n250_ );
and g114 ( new_n252_, N1, N5 );
or g115 ( new_n253_, new_n251_, new_n252_ );
or g116 ( new_n254_, new_n253_, new_n249_ );
or g117 ( new_n255_, N1, N5 );
not g118 ( new_n256_, new_n252_ );
and g119 ( new_n257_, new_n256_, new_n255_ );
or g120 ( new_n258_, new_n257_, keyIn_0_0 );
and g121 ( new_n259_, new_n254_, new_n258_ );
or g122 ( new_n260_, new_n248_, new_n259_ );
or g123 ( new_n261_, new_n246_, new_n243_ );
or g124 ( new_n262_, new_n241_, keyIn_0_1 );
and g125 ( new_n263_, new_n262_, new_n261_ );
and g126 ( new_n264_, new_n257_, keyIn_0_0 );
and g127 ( new_n265_, new_n253_, new_n249_ );
or g128 ( new_n266_, new_n265_, new_n264_ );
or g129 ( new_n267_, new_n266_, new_n263_ );
and g130 ( new_n268_, new_n260_, new_n267_ );
or g131 ( new_n269_, new_n268_, keyIn_0_12 );
not g132 ( new_n270_, keyIn_0_12 );
and g133 ( new_n271_, new_n266_, new_n263_ );
and g134 ( new_n272_, new_n248_, new_n259_ );
or g135 ( new_n273_, new_n271_, new_n272_ );
or g136 ( new_n274_, new_n273_, new_n270_ );
and g137 ( new_n275_, new_n269_, new_n274_ );
and g138 ( new_n276_, new_n236_, new_n275_ );
or g139 ( new_n277_, new_n234_, keyIn_0_13 );
or g140 ( new_n278_, new_n230_, new_n198_ );
and g141 ( new_n279_, new_n277_, new_n278_ );
and g142 ( new_n280_, new_n273_, new_n270_ );
and g143 ( new_n281_, new_n268_, keyIn_0_12 );
or g144 ( new_n282_, new_n280_, new_n281_ );
and g145 ( new_n283_, new_n282_, new_n279_ );
or g146 ( new_n284_, new_n276_, new_n283_ );
and g147 ( new_n285_, new_n284_, keyIn_0_18 );
not g148 ( new_n286_, keyIn_0_18 );
or g149 ( new_n287_, new_n282_, new_n279_ );
or g150 ( new_n288_, new_n236_, new_n275_ );
and g151 ( new_n289_, new_n287_, new_n288_ );
and g152 ( new_n290_, new_n289_, new_n286_ );
or g153 ( new_n291_, new_n285_, new_n290_ );
and g154 ( new_n292_, N133, N137 );
and g155 ( new_n293_, new_n292_, keyIn_0_6 );
not g156 ( new_n294_, new_n293_ );
or g157 ( new_n295_, new_n292_, keyIn_0_6 );
and g158 ( new_n296_, new_n294_, new_n295_ );
not g159 ( new_n297_, new_n296_ );
and g160 ( new_n298_, new_n291_, new_n297_ );
or g161 ( new_n299_, new_n289_, new_n286_ );
or g162 ( new_n300_, new_n284_, keyIn_0_18 );
and g163 ( new_n301_, new_n300_, new_n299_ );
and g164 ( new_n302_, new_n301_, new_n296_ );
or g165 ( new_n303_, new_n298_, new_n302_ );
and g166 ( new_n304_, new_n303_, keyIn_0_20 );
not g167 ( new_n305_, keyIn_0_20 );
or g168 ( new_n306_, new_n301_, new_n296_ );
or g169 ( new_n307_, new_n291_, new_n297_ );
and g170 ( new_n308_, new_n307_, new_n306_ );
and g171 ( new_n309_, new_n308_, new_n305_ );
or g172 ( new_n310_, new_n304_, new_n309_ );
and g173 ( new_n311_, new_n155_, N65 );
and g174 ( new_n312_, new_n140_, N81 );
or g175 ( new_n313_, new_n311_, new_n312_ );
and g176 ( new_n314_, new_n313_, keyIn_0_8 );
not g177 ( new_n315_, new_n314_ );
or g178 ( new_n316_, new_n313_, keyIn_0_8 );
and g179 ( new_n317_, new_n315_, new_n316_ );
not g180 ( new_n318_, new_n317_ );
not g181 ( new_n319_, N97 );
not g182 ( new_n320_, N113 );
and g183 ( new_n321_, new_n319_, new_n320_ );
and g184 ( new_n322_, N97, N113 );
or g185 ( new_n323_, new_n321_, new_n322_ );
and g186 ( new_n324_, new_n323_, keyIn_0_9 );
not g187 ( new_n325_, new_n324_ );
or g188 ( new_n326_, new_n323_, keyIn_0_9 );
and g189 ( new_n327_, new_n325_, new_n326_ );
not g190 ( new_n328_, new_n327_ );
and g191 ( new_n329_, new_n318_, new_n328_ );
and g192 ( new_n330_, new_n317_, new_n327_ );
or g193 ( new_n331_, new_n329_, new_n330_ );
and g194 ( new_n332_, new_n331_, keyIn_0_16 );
not g195 ( new_n333_, new_n332_ );
or g196 ( new_n334_, new_n331_, keyIn_0_16 );
and g197 ( new_n335_, new_n333_, new_n334_ );
not g198 ( new_n336_, new_n335_ );
and g199 ( new_n337_, new_n310_, new_n336_ );
or g200 ( new_n338_, new_n308_, new_n305_ );
or g201 ( new_n339_, new_n303_, keyIn_0_20 );
and g202 ( new_n340_, new_n339_, new_n338_ );
and g203 ( new_n341_, new_n340_, new_n335_ );
or g204 ( new_n342_, new_n337_, new_n341_ );
or g205 ( new_n343_, new_n342_, new_n197_ );
or g206 ( new_n344_, new_n340_, new_n335_ );
or g207 ( new_n345_, new_n310_, new_n336_ );
and g208 ( new_n346_, new_n345_, new_n344_ );
or g209 ( new_n347_, new_n346_, keyIn_0_22 );
and g210 ( new_n348_, new_n343_, new_n347_ );
not g211 ( new_n349_, keyIn_0_14 );
not g212 ( new_n350_, N41 );
not g213 ( new_n351_, N45 );
and g214 ( new_n352_, new_n350_, new_n351_ );
and g215 ( new_n353_, N41, N45 );
or g216 ( new_n354_, new_n352_, new_n353_ );
and g217 ( new_n355_, new_n354_, keyIn_0_5 );
not g218 ( new_n356_, keyIn_0_5 );
or g219 ( new_n357_, N41, N45 );
not g220 ( new_n358_, new_n353_ );
and g221 ( new_n359_, new_n358_, new_n357_ );
and g222 ( new_n360_, new_n359_, new_n356_ );
or g223 ( new_n361_, new_n355_, new_n360_ );
not g224 ( new_n362_, N37 );
and g225 ( new_n363_, new_n183_, new_n362_ );
and g226 ( new_n364_, N33, N37 );
or g227 ( new_n365_, new_n363_, new_n364_ );
and g228 ( new_n366_, new_n365_, keyIn_0_4 );
not g229 ( new_n367_, keyIn_0_4 );
or g230 ( new_n368_, N33, N37 );
not g231 ( new_n369_, new_n364_ );
and g232 ( new_n370_, new_n369_, new_n368_ );
and g233 ( new_n371_, new_n370_, new_n367_ );
or g234 ( new_n372_, new_n366_, new_n371_ );
and g235 ( new_n373_, new_n361_, new_n372_ );
or g236 ( new_n374_, new_n359_, new_n356_ );
or g237 ( new_n375_, new_n354_, keyIn_0_5 );
and g238 ( new_n376_, new_n375_, new_n374_ );
or g239 ( new_n377_, new_n370_, new_n367_ );
or g240 ( new_n378_, new_n365_, keyIn_0_4 );
and g241 ( new_n379_, new_n378_, new_n377_ );
and g242 ( new_n380_, new_n376_, new_n379_ );
or g243 ( new_n381_, new_n373_, new_n380_ );
and g244 ( new_n382_, new_n381_, new_n349_ );
or g245 ( new_n383_, new_n376_, new_n379_ );
or g246 ( new_n384_, new_n361_, new_n372_ );
and g247 ( new_n385_, new_n384_, new_n383_ );
and g248 ( new_n386_, new_n385_, keyIn_0_14 );
or g249 ( new_n387_, new_n382_, new_n386_ );
not g250 ( new_n388_, N53 );
and g251 ( new_n389_, new_n184_, new_n388_ );
and g252 ( new_n390_, N49, N53 );
or g253 ( new_n391_, new_n389_, new_n390_ );
not g254 ( new_n392_, N57 );
not g255 ( new_n393_, N61 );
and g256 ( new_n394_, new_n392_, new_n393_ );
and g257 ( new_n395_, N57, N61 );
or g258 ( new_n396_, new_n394_, new_n395_ );
and g259 ( new_n397_, new_n391_, new_n396_ );
not g260 ( new_n398_, new_n397_ );
or g261 ( new_n399_, new_n391_, new_n396_ );
and g262 ( new_n400_, new_n398_, new_n399_ );
not g263 ( new_n401_, new_n400_ );
and g264 ( new_n402_, new_n387_, new_n401_ );
or g265 ( new_n403_, new_n385_, keyIn_0_14 );
or g266 ( new_n404_, new_n381_, new_n349_ );
and g267 ( new_n405_, new_n403_, new_n404_ );
and g268 ( new_n406_, new_n405_, new_n400_ );
or g269 ( new_n407_, new_n402_, new_n406_ );
and g270 ( new_n408_, N134, N137 );
not g271 ( new_n409_, new_n408_ );
and g272 ( new_n410_, new_n407_, new_n409_ );
not g273 ( new_n411_, new_n410_ );
or g274 ( new_n412_, new_n407_, new_n409_ );
and g275 ( new_n413_, new_n411_, new_n412_ );
not g276 ( new_n414_, new_n413_ );
and g277 ( new_n415_, new_n153_, N69 );
and g278 ( new_n416_, new_n138_, N85 );
or g279 ( new_n417_, new_n415_, new_n416_ );
not g280 ( new_n418_, N101 );
not g281 ( new_n419_, N117 );
and g282 ( new_n420_, new_n418_, new_n419_ );
and g283 ( new_n421_, N101, N117 );
or g284 ( new_n422_, new_n420_, new_n421_ );
and g285 ( new_n423_, new_n417_, new_n422_ );
not g286 ( new_n424_, new_n423_ );
or g287 ( new_n425_, new_n417_, new_n422_ );
and g288 ( new_n426_, new_n424_, new_n425_ );
not g289 ( new_n427_, new_n426_ );
and g290 ( new_n428_, new_n414_, new_n427_ );
and g291 ( new_n429_, new_n413_, new_n426_ );
or g292 ( new_n430_, new_n428_, new_n429_ );
and g293 ( new_n431_, new_n348_, new_n430_ );
not g294 ( new_n432_, keyIn_0_19 );
or g295 ( new_n433_, new_n282_, new_n387_ );
or g296 ( new_n434_, new_n275_, new_n405_ );
and g297 ( new_n435_, new_n433_, new_n434_ );
and g298 ( new_n436_, new_n435_, new_n432_ );
and g299 ( new_n437_, new_n275_, new_n405_ );
and g300 ( new_n438_, new_n282_, new_n387_ );
or g301 ( new_n439_, new_n438_, new_n437_ );
and g302 ( new_n440_, new_n439_, keyIn_0_19 );
or g303 ( new_n441_, new_n436_, new_n440_ );
and g304 ( new_n442_, N135, N137 );
and g305 ( new_n443_, new_n442_, keyIn_0_7 );
not g306 ( new_n444_, new_n443_ );
or g307 ( new_n445_, new_n442_, keyIn_0_7 );
and g308 ( new_n446_, new_n444_, new_n445_ );
not g309 ( new_n447_, new_n446_ );
and g310 ( new_n448_, new_n441_, new_n447_ );
or g311 ( new_n449_, new_n439_, keyIn_0_19 );
or g312 ( new_n450_, new_n435_, new_n432_ );
and g313 ( new_n451_, new_n450_, new_n449_ );
and g314 ( new_n452_, new_n451_, new_n446_ );
or g315 ( new_n453_, new_n448_, new_n452_ );
and g316 ( new_n454_, new_n453_, keyIn_0_21 );
not g317 ( new_n455_, keyIn_0_21 );
or g318 ( new_n456_, new_n451_, new_n446_ );
or g319 ( new_n457_, new_n441_, new_n447_ );
and g320 ( new_n458_, new_n457_, new_n456_ );
and g321 ( new_n459_, new_n458_, new_n455_ );
or g322 ( new_n460_, new_n454_, new_n459_ );
not g323 ( new_n461_, keyIn_0_17 );
and g324 ( new_n462_, new_n158_, N73 );
and g325 ( new_n463_, new_n143_, N89 );
or g326 ( new_n464_, new_n462_, new_n463_ );
and g327 ( new_n465_, new_n464_, keyIn_0_10 );
not g328 ( new_n466_, new_n465_ );
or g329 ( new_n467_, new_n464_, keyIn_0_10 );
and g330 ( new_n468_, new_n466_, new_n467_ );
not g331 ( new_n469_, new_n468_ );
not g332 ( new_n470_, N121 );
and g333 ( new_n471_, new_n470_, N105 );
not g334 ( new_n472_, N105 );
and g335 ( new_n473_, new_n472_, N121 );
or g336 ( new_n474_, new_n471_, new_n473_ );
and g337 ( new_n475_, new_n474_, keyIn_0_11 );
not g338 ( new_n476_, new_n475_ );
or g339 ( new_n477_, new_n474_, keyIn_0_11 );
and g340 ( new_n478_, new_n476_, new_n477_ );
not g341 ( new_n479_, new_n478_ );
and g342 ( new_n480_, new_n469_, new_n479_ );
and g343 ( new_n481_, new_n468_, new_n478_ );
or g344 ( new_n482_, new_n480_, new_n481_ );
and g345 ( new_n483_, new_n482_, new_n461_ );
not g346 ( new_n484_, new_n483_ );
or g347 ( new_n485_, new_n482_, new_n461_ );
and g348 ( new_n486_, new_n484_, new_n485_ );
and g349 ( new_n487_, new_n460_, new_n486_ );
or g350 ( new_n488_, new_n458_, new_n455_ );
or g351 ( new_n489_, new_n453_, keyIn_0_21 );
and g352 ( new_n490_, new_n489_, new_n488_ );
not g353 ( new_n491_, new_n486_ );
and g354 ( new_n492_, new_n490_, new_n491_ );
or g355 ( new_n493_, new_n487_, new_n492_ );
or g356 ( new_n494_, new_n493_, keyIn_0_23 );
not g357 ( new_n495_, keyIn_0_23 );
or g358 ( new_n496_, new_n490_, new_n491_ );
or g359 ( new_n497_, new_n460_, new_n486_ );
and g360 ( new_n498_, new_n497_, new_n496_ );
or g361 ( new_n499_, new_n498_, new_n495_ );
and g362 ( new_n500_, new_n494_, new_n499_ );
not g363 ( new_n501_, keyIn_0_24 );
and g364 ( new_n502_, new_n195_, new_n501_ );
not g365 ( new_n503_, new_n502_ );
and g366 ( new_n504_, new_n196_, keyIn_0_24 );
not g367 ( new_n505_, new_n504_ );
and g368 ( new_n506_, new_n418_, N97 );
and g369 ( new_n507_, new_n319_, N101 );
or g370 ( new_n508_, new_n506_, new_n507_ );
not g371 ( new_n509_, N109 );
and g372 ( new_n510_, new_n472_, new_n509_ );
and g373 ( new_n511_, N105, N109 );
or g374 ( new_n512_, new_n510_, new_n511_ );
and g375 ( new_n513_, new_n508_, new_n512_ );
not g376 ( new_n514_, new_n513_ );
or g377 ( new_n515_, new_n508_, new_n512_ );
and g378 ( new_n516_, new_n514_, new_n515_ );
and g379 ( new_n517_, new_n152_, new_n516_ );
not g380 ( new_n518_, new_n516_ );
and g381 ( new_n519_, new_n518_, new_n151_ );
or g382 ( new_n520_, new_n517_, new_n519_ );
and g383 ( new_n521_, N131, N137 );
not g384 ( new_n522_, new_n521_ );
and g385 ( new_n523_, new_n520_, new_n522_ );
not g386 ( new_n524_, new_n523_ );
or g387 ( new_n525_, new_n520_, new_n522_ );
and g388 ( new_n526_, new_n524_, new_n525_ );
not g389 ( new_n527_, new_n526_ );
and g390 ( new_n528_, new_n210_, N9 );
and g391 ( new_n529_, new_n237_, N25 );
or g392 ( new_n530_, new_n528_, new_n529_ );
and g393 ( new_n531_, new_n350_, new_n392_ );
and g394 ( new_n532_, N41, N57 );
or g395 ( new_n533_, new_n531_, new_n532_ );
and g396 ( new_n534_, new_n530_, new_n533_ );
not g397 ( new_n535_, new_n534_ );
or g398 ( new_n536_, new_n530_, new_n533_ );
and g399 ( new_n537_, new_n535_, new_n536_ );
not g400 ( new_n538_, new_n537_ );
and g401 ( new_n539_, new_n527_, new_n538_ );
and g402 ( new_n540_, new_n526_, new_n537_ );
or g403 ( new_n541_, new_n539_, new_n540_ );
not g404 ( new_n542_, new_n541_ );
and g405 ( new_n543_, new_n419_, N113 );
and g406 ( new_n544_, new_n320_, N117 );
or g407 ( new_n545_, new_n543_, new_n544_ );
not g408 ( new_n546_, N125 );
and g409 ( new_n547_, new_n470_, new_n546_ );
and g410 ( new_n548_, N121, N125 );
or g411 ( new_n549_, new_n547_, new_n548_ );
and g412 ( new_n550_, new_n545_, new_n549_ );
not g413 ( new_n551_, new_n550_ );
or g414 ( new_n552_, new_n545_, new_n549_ );
and g415 ( new_n553_, new_n551_, new_n552_ );
not g416 ( new_n554_, new_n553_ );
and g417 ( new_n555_, new_n554_, new_n516_ );
and g418 ( new_n556_, new_n518_, new_n553_ );
or g419 ( new_n557_, new_n555_, new_n556_ );
and g420 ( new_n558_, N130, N137 );
not g421 ( new_n559_, new_n558_ );
and g422 ( new_n560_, new_n557_, new_n559_ );
not g423 ( new_n561_, new_n560_ );
or g424 ( new_n562_, new_n557_, new_n559_ );
and g425 ( new_n563_, new_n561_, new_n562_ );
not g426 ( new_n564_, new_n563_ );
and g427 ( new_n565_, new_n199_, N5 );
and g428 ( new_n566_, new_n250_, N21 );
or g429 ( new_n567_, new_n565_, new_n566_ );
and g430 ( new_n568_, new_n362_, new_n388_ );
and g431 ( new_n569_, N37, N53 );
or g432 ( new_n570_, new_n568_, new_n569_ );
and g433 ( new_n571_, new_n567_, new_n570_ );
not g434 ( new_n572_, new_n571_ );
or g435 ( new_n573_, new_n567_, new_n570_ );
and g436 ( new_n574_, new_n572_, new_n573_ );
not g437 ( new_n575_, new_n574_ );
and g438 ( new_n576_, new_n564_, new_n575_ );
and g439 ( new_n577_, new_n563_, new_n574_ );
or g440 ( new_n578_, new_n576_, new_n577_ );
and g441 ( new_n579_, new_n542_, new_n578_ );
and g442 ( new_n580_, new_n505_, new_n579_ );
and g443 ( new_n581_, new_n580_, new_n503_ );
not g444 ( new_n582_, new_n581_ );
and g445 ( new_n583_, new_n196_, new_n578_ );
and g446 ( new_n584_, new_n583_, new_n541_ );
not g447 ( new_n585_, new_n584_ );
not g448 ( new_n586_, new_n578_ );
and g449 ( new_n587_, new_n586_, new_n195_ );
and g450 ( new_n588_, new_n587_, new_n541_ );
not g451 ( new_n589_, new_n588_ );
and g452 ( new_n590_, new_n585_, new_n589_ );
and g453 ( new_n591_, new_n582_, new_n590_ );
and g454 ( new_n592_, new_n168_, new_n553_ );
and g455 ( new_n593_, new_n554_, new_n166_ );
or g456 ( new_n594_, new_n592_, new_n593_ );
and g457 ( new_n595_, N132, N137 );
not g458 ( new_n596_, new_n595_ );
and g459 ( new_n597_, new_n594_, new_n596_ );
not g460 ( new_n598_, new_n597_ );
or g461 ( new_n599_, new_n594_, new_n596_ );
and g462 ( new_n600_, new_n598_, new_n599_ );
not g463 ( new_n601_, new_n600_ );
and g464 ( new_n602_, new_n211_, N13 );
and g465 ( new_n603_, new_n238_, N29 );
or g466 ( new_n604_, new_n602_, new_n603_ );
and g467 ( new_n605_, new_n351_, new_n393_ );
and g468 ( new_n606_, N45, N61 );
or g469 ( new_n607_, new_n605_, new_n606_ );
and g470 ( new_n608_, new_n604_, new_n607_ );
not g471 ( new_n609_, new_n608_ );
or g472 ( new_n610_, new_n604_, new_n607_ );
and g473 ( new_n611_, new_n609_, new_n610_ );
not g474 ( new_n612_, new_n611_ );
and g475 ( new_n613_, new_n612_, keyIn_0_15 );
not g476 ( new_n614_, new_n613_ );
or g477 ( new_n615_, new_n612_, keyIn_0_15 );
and g478 ( new_n616_, new_n614_, new_n615_ );
not g479 ( new_n617_, new_n616_ );
and g480 ( new_n618_, new_n601_, new_n617_ );
and g481 ( new_n619_, new_n600_, new_n616_ );
or g482 ( new_n620_, new_n618_, new_n619_ );
not g483 ( new_n621_, new_n620_ );
or g484 ( new_n622_, new_n591_, new_n621_ );
and g485 ( new_n623_, new_n195_, new_n541_ );
and g486 ( new_n624_, new_n621_, new_n578_ );
and g487 ( new_n625_, new_n624_, new_n623_ );
not g488 ( new_n626_, new_n625_ );
and g489 ( new_n627_, new_n622_, new_n626_ );
not g490 ( new_n628_, new_n627_ );
and g491 ( new_n629_, new_n236_, new_n401_ );
and g492 ( new_n630_, new_n279_, new_n400_ );
or g493 ( new_n631_, new_n629_, new_n630_ );
and g494 ( new_n632_, N136, N137 );
not g495 ( new_n633_, new_n632_ );
and g496 ( new_n634_, new_n631_, new_n633_ );
not g497 ( new_n635_, new_n634_ );
or g498 ( new_n636_, new_n631_, new_n633_ );
and g499 ( new_n637_, new_n635_, new_n636_ );
not g500 ( new_n638_, new_n637_ );
and g501 ( new_n639_, new_n159_, N77 );
and g502 ( new_n640_, new_n144_, N93 );
or g503 ( new_n641_, new_n639_, new_n640_ );
and g504 ( new_n642_, new_n509_, new_n546_ );
and g505 ( new_n643_, N109, N125 );
or g506 ( new_n644_, new_n642_, new_n643_ );
and g507 ( new_n645_, new_n641_, new_n644_ );
not g508 ( new_n646_, new_n645_ );
or g509 ( new_n647_, new_n641_, new_n644_ );
and g510 ( new_n648_, new_n646_, new_n647_ );
not g511 ( new_n649_, new_n648_ );
and g512 ( new_n650_, new_n638_, new_n649_ );
and g513 ( new_n651_, new_n637_, new_n648_ );
or g514 ( new_n652_, new_n650_, new_n651_ );
and g515 ( new_n653_, new_n628_, new_n652_ );
and g516 ( new_n654_, new_n500_, new_n653_ );
and g517 ( new_n655_, new_n431_, new_n654_ );
and g518 ( new_n656_, new_n655_, new_n196_ );
not g519 ( new_n657_, new_n656_ );
and g520 ( new_n658_, new_n657_, N1 );
and g521 ( new_n659_, new_n656_, new_n180_ );
or g522 ( N724, new_n658_, new_n659_ );
and g523 ( new_n661_, new_n655_, new_n586_ );
not g524 ( new_n662_, new_n661_ );
and g525 ( new_n663_, new_n662_, N5 );
and g526 ( new_n664_, new_n661_, new_n250_ );
or g527 ( N725, new_n663_, new_n664_ );
and g528 ( new_n666_, new_n655_, new_n542_ );
not g529 ( new_n667_, new_n666_ );
and g530 ( new_n668_, new_n667_, N9 );
and g531 ( new_n669_, new_n666_, new_n237_ );
or g532 ( N726, new_n668_, new_n669_ );
and g533 ( new_n671_, new_n655_, new_n621_ );
not g534 ( new_n672_, new_n671_ );
and g535 ( new_n673_, new_n672_, N13 );
and g536 ( new_n674_, new_n671_, new_n238_ );
or g537 ( N727, new_n673_, new_n674_ );
and g538 ( new_n676_, new_n498_, new_n495_ );
and g539 ( new_n677_, new_n493_, keyIn_0_23 );
or g540 ( new_n678_, new_n677_, new_n676_ );
not g541 ( new_n679_, new_n652_ );
and g542 ( new_n680_, new_n628_, new_n679_ );
and g543 ( new_n681_, new_n678_, new_n680_ );
and g544 ( new_n682_, new_n681_, new_n431_ );
and g545 ( new_n683_, new_n682_, new_n196_ );
not g546 ( new_n684_, new_n683_ );
and g547 ( new_n685_, new_n684_, N17 );
and g548 ( new_n686_, new_n683_, new_n178_ );
or g549 ( N728, new_n685_, new_n686_ );
and g550 ( new_n688_, new_n682_, new_n586_ );
not g551 ( new_n689_, new_n688_ );
and g552 ( new_n690_, new_n689_, N21 );
and g553 ( new_n691_, new_n688_, new_n199_ );
or g554 ( N729, new_n690_, new_n691_ );
and g555 ( new_n693_, new_n682_, new_n542_ );
not g556 ( new_n694_, new_n693_ );
and g557 ( new_n695_, new_n694_, N25 );
and g558 ( new_n696_, new_n693_, new_n210_ );
or g559 ( N730, new_n695_, new_n696_ );
and g560 ( new_n698_, new_n682_, new_n621_ );
not g561 ( new_n699_, new_n698_ );
and g562 ( new_n700_, new_n699_, N29 );
and g563 ( new_n701_, new_n698_, new_n211_ );
or g564 ( N731, new_n700_, new_n701_ );
and g565 ( new_n703_, new_n346_, keyIn_0_22 );
and g566 ( new_n704_, new_n342_, new_n197_ );
or g567 ( new_n705_, new_n704_, new_n703_ );
not g568 ( new_n706_, new_n430_ );
and g569 ( new_n707_, new_n705_, new_n706_ );
and g570 ( new_n708_, new_n707_, new_n654_ );
and g571 ( new_n709_, new_n708_, new_n196_ );
not g572 ( new_n710_, new_n709_ );
and g573 ( new_n711_, new_n710_, N33 );
and g574 ( new_n712_, new_n709_, new_n183_ );
or g575 ( N732, new_n711_, new_n712_ );
and g576 ( new_n714_, new_n708_, new_n586_ );
not g577 ( new_n715_, new_n714_ );
and g578 ( new_n716_, new_n715_, N37 );
and g579 ( new_n717_, new_n714_, new_n362_ );
or g580 ( N733, new_n716_, new_n717_ );
and g581 ( new_n719_, new_n708_, new_n542_ );
not g582 ( new_n720_, new_n719_ );
and g583 ( new_n721_, new_n720_, N41 );
and g584 ( new_n722_, new_n719_, new_n350_ );
or g585 ( N734, new_n721_, new_n722_ );
and g586 ( new_n724_, new_n708_, new_n621_ );
not g587 ( new_n725_, new_n724_ );
and g588 ( new_n726_, new_n725_, N45 );
and g589 ( new_n727_, new_n724_, new_n351_ );
or g590 ( N735, new_n726_, new_n727_ );
and g591 ( new_n729_, new_n681_, new_n707_ );
and g592 ( new_n730_, new_n729_, new_n196_ );
not g593 ( new_n731_, new_n730_ );
and g594 ( new_n732_, new_n731_, N49 );
and g595 ( new_n733_, new_n730_, new_n184_ );
or g596 ( N736, new_n732_, new_n733_ );
and g597 ( new_n735_, new_n729_, new_n586_ );
not g598 ( new_n736_, new_n735_ );
and g599 ( new_n737_, new_n736_, N53 );
and g600 ( new_n738_, new_n735_, new_n388_ );
or g601 ( N737, new_n737_, new_n738_ );
and g602 ( new_n740_, new_n729_, new_n542_ );
not g603 ( new_n741_, new_n740_ );
and g604 ( new_n742_, new_n741_, N57 );
and g605 ( new_n743_, new_n740_, new_n392_ );
or g606 ( N738, new_n742_, new_n743_ );
and g607 ( new_n745_, new_n729_, new_n621_ );
not g608 ( new_n746_, new_n745_ );
and g609 ( new_n747_, new_n746_, N61 );
and g610 ( new_n748_, new_n745_, new_n393_ );
or g611 ( N739, new_n747_, new_n748_ );
not g612 ( new_n750_, keyIn_0_52 );
not g613 ( new_n751_, keyIn_0_36 );
and g614 ( new_n752_, new_n500_, keyIn_0_27 );
not g615 ( new_n753_, new_n752_ );
or g616 ( new_n754_, new_n500_, keyIn_0_27 );
and g617 ( new_n755_, new_n753_, new_n754_ );
not g618 ( new_n756_, keyIn_0_25 );
and g619 ( new_n757_, new_n348_, new_n756_ );
and g620 ( new_n758_, new_n705_, keyIn_0_25 );
not g621 ( new_n759_, keyIn_0_26 );
and g622 ( new_n760_, new_n430_, new_n759_ );
and g623 ( new_n761_, new_n706_, keyIn_0_26 );
or g624 ( new_n762_, new_n761_, new_n652_ );
or g625 ( new_n763_, new_n762_, new_n760_ );
or g626 ( new_n764_, new_n758_, new_n763_ );
or g627 ( new_n765_, new_n764_, new_n757_ );
or g628 ( new_n766_, new_n765_, new_n755_ );
and g629 ( new_n767_, new_n766_, keyIn_0_32 );
not g630 ( new_n768_, new_n767_ );
or g631 ( new_n769_, new_n766_, keyIn_0_32 );
and g632 ( new_n770_, new_n768_, new_n769_ );
not g633 ( new_n771_, new_n770_ );
or g634 ( new_n772_, new_n678_, keyIn_0_31 );
not g635 ( new_n773_, keyIn_0_31 );
or g636 ( new_n774_, new_n500_, new_n773_ );
and g637 ( new_n775_, new_n772_, new_n774_ );
or g638 ( new_n776_, new_n705_, new_n706_ );
or g639 ( new_n777_, new_n776_, new_n679_ );
or g640 ( new_n778_, new_n777_, new_n775_ );
and g641 ( new_n779_, new_n778_, keyIn_0_35 );
not g642 ( new_n780_, keyIn_0_35 );
and g643 ( new_n781_, new_n500_, new_n773_ );
and g644 ( new_n782_, new_n678_, keyIn_0_31 );
or g645 ( new_n783_, new_n782_, new_n781_ );
and g646 ( new_n784_, new_n431_, new_n652_ );
and g647 ( new_n785_, new_n783_, new_n784_ );
and g648 ( new_n786_, new_n785_, new_n780_ );
or g649 ( new_n787_, new_n779_, new_n786_ );
not g650 ( new_n788_, keyIn_0_33 );
not g651 ( new_n789_, keyIn_0_28 );
and g652 ( new_n790_, new_n705_, new_n789_ );
and g653 ( new_n791_, new_n348_, keyIn_0_28 );
and g654 ( new_n792_, new_n430_, new_n652_ );
not g655 ( new_n793_, new_n792_ );
or g656 ( new_n794_, new_n678_, new_n793_ );
or g657 ( new_n795_, new_n794_, new_n791_ );
or g658 ( new_n796_, new_n795_, new_n790_ );
and g659 ( new_n797_, new_n796_, new_n788_ );
not g660 ( new_n798_, new_n790_ );
or g661 ( new_n799_, new_n705_, new_n789_ );
and g662 ( new_n800_, new_n500_, new_n792_ );
and g663 ( new_n801_, new_n799_, new_n800_ );
and g664 ( new_n802_, new_n801_, new_n798_ );
and g665 ( new_n803_, new_n802_, keyIn_0_33 );
or g666 ( new_n804_, new_n797_, new_n803_ );
and g667 ( new_n805_, new_n787_, new_n804_ );
not g668 ( new_n806_, keyIn_0_34 );
and g669 ( new_n807_, new_n705_, keyIn_0_29 );
not g670 ( new_n808_, new_n807_ );
or g671 ( new_n809_, new_n705_, keyIn_0_29 );
and g672 ( new_n810_, new_n808_, new_n809_ );
not g673 ( new_n811_, keyIn_0_30 );
and g674 ( new_n812_, new_n678_, new_n811_ );
and g675 ( new_n813_, new_n500_, keyIn_0_30 );
and g676 ( new_n814_, new_n706_, new_n652_ );
not g677 ( new_n815_, new_n814_ );
or g678 ( new_n816_, new_n813_, new_n815_ );
or g679 ( new_n817_, new_n816_, new_n812_ );
or g680 ( new_n818_, new_n817_, new_n810_ );
or g681 ( new_n819_, new_n818_, new_n806_ );
not g682 ( new_n820_, new_n810_ );
not g683 ( new_n821_, new_n812_ );
or g684 ( new_n822_, new_n678_, new_n811_ );
and g685 ( new_n823_, new_n822_, new_n814_ );
and g686 ( new_n824_, new_n823_, new_n821_ );
and g687 ( new_n825_, new_n824_, new_n820_ );
or g688 ( new_n826_, new_n825_, keyIn_0_34 );
and g689 ( new_n827_, new_n819_, new_n826_ );
and g690 ( new_n828_, new_n805_, new_n827_ );
and g691 ( new_n829_, new_n828_, new_n771_ );
and g692 ( new_n830_, new_n829_, new_n751_ );
not g693 ( new_n831_, new_n830_ );
or g694 ( new_n832_, new_n829_, new_n751_ );
and g695 ( new_n833_, new_n831_, new_n832_ );
and g696 ( new_n834_, new_n542_, new_n620_ );
and g697 ( new_n835_, new_n583_, new_n834_ );
not g698 ( new_n836_, new_n835_ );
or g699 ( new_n837_, new_n833_, new_n836_ );
or g700 ( new_n838_, new_n837_, keyIn_0_37 );
not g701 ( new_n839_, keyIn_0_37 );
or g702 ( new_n840_, new_n785_, new_n780_ );
or g703 ( new_n841_, new_n778_, keyIn_0_35 );
and g704 ( new_n842_, new_n841_, new_n840_ );
or g705 ( new_n843_, new_n802_, keyIn_0_33 );
or g706 ( new_n844_, new_n796_, new_n788_ );
and g707 ( new_n845_, new_n844_, new_n843_ );
or g708 ( new_n846_, new_n842_, new_n845_ );
and g709 ( new_n847_, new_n825_, keyIn_0_34 );
and g710 ( new_n848_, new_n818_, new_n806_ );
or g711 ( new_n849_, new_n848_, new_n847_ );
or g712 ( new_n850_, new_n846_, new_n849_ );
or g713 ( new_n851_, new_n850_, new_n770_ );
and g714 ( new_n852_, new_n851_, keyIn_0_36 );
or g715 ( new_n853_, new_n852_, new_n830_ );
and g716 ( new_n854_, new_n853_, new_n835_ );
or g717 ( new_n855_, new_n854_, new_n839_ );
and g718 ( new_n856_, new_n838_, new_n855_ );
or g719 ( new_n857_, new_n856_, new_n705_ );
and g720 ( new_n858_, new_n857_, keyIn_0_40 );
not g721 ( new_n859_, keyIn_0_40 );
and g722 ( new_n860_, new_n854_, new_n839_ );
and g723 ( new_n861_, new_n837_, keyIn_0_37 );
or g724 ( new_n862_, new_n861_, new_n860_ );
and g725 ( new_n863_, new_n862_, new_n348_ );
and g726 ( new_n864_, new_n863_, new_n859_ );
or g727 ( new_n865_, new_n858_, new_n864_ );
and g728 ( new_n866_, new_n865_, N65 );
or g729 ( new_n867_, new_n863_, new_n859_ );
or g730 ( new_n868_, new_n857_, keyIn_0_40 );
and g731 ( new_n869_, new_n868_, new_n867_ );
and g732 ( new_n870_, new_n869_, new_n140_ );
or g733 ( new_n871_, new_n866_, new_n870_ );
and g734 ( new_n872_, new_n871_, new_n750_ );
or g735 ( new_n873_, new_n869_, new_n140_ );
or g736 ( new_n874_, new_n865_, N65 );
and g737 ( new_n875_, new_n874_, new_n873_ );
and g738 ( new_n876_, new_n875_, keyIn_0_52 );
or g739 ( N740, new_n872_, new_n876_ );
not g740 ( new_n878_, keyIn_0_53 );
not g741 ( new_n879_, keyIn_0_41 );
or g742 ( new_n880_, new_n856_, new_n430_ );
and g743 ( new_n881_, new_n880_, new_n879_ );
and g744 ( new_n882_, new_n862_, new_n706_ );
and g745 ( new_n883_, new_n882_, keyIn_0_41 );
or g746 ( new_n884_, new_n881_, new_n883_ );
and g747 ( new_n885_, new_n884_, new_n138_ );
or g748 ( new_n886_, new_n882_, keyIn_0_41 );
or g749 ( new_n887_, new_n880_, new_n879_ );
and g750 ( new_n888_, new_n887_, new_n886_ );
and g751 ( new_n889_, new_n888_, N69 );
or g752 ( new_n890_, new_n885_, new_n889_ );
and g753 ( new_n891_, new_n890_, new_n878_ );
or g754 ( new_n892_, new_n888_, N69 );
or g755 ( new_n893_, new_n884_, new_n138_ );
and g756 ( new_n894_, new_n893_, new_n892_ );
and g757 ( new_n895_, new_n894_, keyIn_0_53 );
or g758 ( N741, new_n891_, new_n895_ );
or g759 ( new_n897_, new_n856_, new_n678_ );
and g760 ( new_n898_, new_n897_, keyIn_0_42 );
not g761 ( new_n899_, keyIn_0_42 );
and g762 ( new_n900_, new_n862_, new_n500_ );
and g763 ( new_n901_, new_n900_, new_n899_ );
or g764 ( new_n902_, new_n898_, new_n901_ );
and g765 ( new_n903_, new_n902_, new_n143_ );
or g766 ( new_n904_, new_n900_, new_n899_ );
or g767 ( new_n905_, new_n897_, keyIn_0_42 );
and g768 ( new_n906_, new_n905_, new_n904_ );
and g769 ( new_n907_, new_n906_, N73 );
or g770 ( new_n908_, new_n903_, new_n907_ );
and g771 ( new_n909_, new_n908_, keyIn_0_54 );
not g772 ( new_n910_, keyIn_0_54 );
or g773 ( new_n911_, new_n906_, N73 );
or g774 ( new_n912_, new_n902_, new_n143_ );
and g775 ( new_n913_, new_n912_, new_n911_ );
and g776 ( new_n914_, new_n913_, new_n910_ );
or g777 ( N742, new_n909_, new_n914_ );
not g778 ( new_n916_, keyIn_0_55 );
or g779 ( new_n917_, new_n856_, new_n652_ );
and g780 ( new_n918_, new_n917_, keyIn_0_43 );
not g781 ( new_n919_, keyIn_0_43 );
and g782 ( new_n920_, new_n862_, new_n679_ );
and g783 ( new_n921_, new_n920_, new_n919_ );
or g784 ( new_n922_, new_n918_, new_n921_ );
and g785 ( new_n923_, new_n922_, N77 );
or g786 ( new_n924_, new_n920_, new_n919_ );
or g787 ( new_n925_, new_n917_, keyIn_0_43 );
and g788 ( new_n926_, new_n925_, new_n924_ );
and g789 ( new_n927_, new_n926_, new_n144_ );
or g790 ( new_n928_, new_n923_, new_n927_ );
and g791 ( new_n929_, new_n928_, new_n916_ );
or g792 ( new_n930_, new_n926_, new_n144_ );
or g793 ( new_n931_, new_n922_, N77 );
and g794 ( new_n932_, new_n931_, new_n930_ );
and g795 ( new_n933_, new_n932_, keyIn_0_55 );
or g796 ( N743, new_n929_, new_n933_ );
not g797 ( new_n935_, keyIn_0_44 );
and g798 ( new_n936_, new_n584_, new_n621_ );
not g799 ( new_n937_, new_n936_ );
or g800 ( new_n938_, new_n833_, new_n937_ );
and g801 ( new_n939_, new_n938_, keyIn_0_38 );
not g802 ( new_n940_, keyIn_0_38 );
and g803 ( new_n941_, new_n853_, new_n936_ );
and g804 ( new_n942_, new_n941_, new_n940_ );
or g805 ( new_n943_, new_n939_, new_n942_ );
or g806 ( new_n944_, new_n943_, new_n705_ );
and g807 ( new_n945_, new_n944_, new_n935_ );
or g808 ( new_n946_, new_n941_, new_n940_ );
or g809 ( new_n947_, new_n938_, keyIn_0_38 );
and g810 ( new_n948_, new_n947_, new_n946_ );
and g811 ( new_n949_, new_n948_, new_n348_ );
and g812 ( new_n950_, new_n949_, keyIn_0_44 );
or g813 ( new_n951_, new_n945_, new_n950_ );
and g814 ( new_n952_, new_n951_, new_n155_ );
or g815 ( new_n953_, new_n949_, keyIn_0_44 );
or g816 ( new_n954_, new_n944_, new_n935_ );
and g817 ( new_n955_, new_n954_, new_n953_ );
and g818 ( new_n956_, new_n955_, N81 );
or g819 ( new_n957_, new_n952_, new_n956_ );
and g820 ( new_n958_, new_n957_, keyIn_0_56 );
not g821 ( new_n959_, keyIn_0_56 );
or g822 ( new_n960_, new_n955_, N81 );
or g823 ( new_n961_, new_n951_, new_n155_ );
and g824 ( new_n962_, new_n960_, new_n961_ );
and g825 ( new_n963_, new_n962_, new_n959_ );
or g826 ( N744, new_n958_, new_n963_ );
not g827 ( new_n965_, keyIn_0_57 );
or g828 ( new_n966_, new_n943_, new_n430_ );
and g829 ( new_n967_, new_n966_, keyIn_0_45 );
not g830 ( new_n968_, keyIn_0_45 );
and g831 ( new_n969_, new_n948_, new_n706_ );
and g832 ( new_n970_, new_n969_, new_n968_ );
or g833 ( new_n971_, new_n967_, new_n970_ );
and g834 ( new_n972_, new_n971_, N85 );
or g835 ( new_n973_, new_n969_, new_n968_ );
or g836 ( new_n974_, new_n966_, keyIn_0_45 );
and g837 ( new_n975_, new_n974_, new_n973_ );
and g838 ( new_n976_, new_n975_, new_n153_ );
or g839 ( new_n977_, new_n972_, new_n976_ );
and g840 ( new_n978_, new_n977_, new_n965_ );
or g841 ( new_n979_, new_n975_, new_n153_ );
or g842 ( new_n980_, new_n971_, N85 );
and g843 ( new_n981_, new_n979_, new_n980_ );
and g844 ( new_n982_, new_n981_, keyIn_0_57 );
or g845 ( N745, new_n978_, new_n982_ );
or g846 ( new_n984_, new_n943_, new_n678_ );
and g847 ( new_n985_, new_n984_, keyIn_0_46 );
not g848 ( new_n986_, keyIn_0_46 );
and g849 ( new_n987_, new_n948_, new_n500_ );
and g850 ( new_n988_, new_n987_, new_n986_ );
or g851 ( new_n989_, new_n985_, new_n988_ );
and g852 ( new_n990_, new_n989_, N89 );
or g853 ( new_n991_, new_n987_, new_n986_ );
or g854 ( new_n992_, new_n984_, keyIn_0_46 );
and g855 ( new_n993_, new_n992_, new_n991_ );
and g856 ( new_n994_, new_n993_, new_n158_ );
or g857 ( new_n995_, new_n990_, new_n994_ );
and g858 ( new_n996_, new_n995_, keyIn_0_58 );
not g859 ( new_n997_, keyIn_0_58 );
or g860 ( new_n998_, new_n993_, new_n158_ );
or g861 ( new_n999_, new_n989_, N89 );
and g862 ( new_n1000_, new_n998_, new_n999_ );
and g863 ( new_n1001_, new_n1000_, new_n997_ );
or g864 ( N746, new_n996_, new_n1001_ );
not g865 ( new_n1003_, keyIn_0_59 );
or g866 ( new_n1004_, new_n943_, new_n652_ );
and g867 ( new_n1005_, new_n1004_, keyIn_0_47 );
not g868 ( new_n1006_, keyIn_0_47 );
and g869 ( new_n1007_, new_n948_, new_n679_ );
and g870 ( new_n1008_, new_n1007_, new_n1006_ );
or g871 ( new_n1009_, new_n1005_, new_n1008_ );
and g872 ( new_n1010_, new_n1009_, N93 );
or g873 ( new_n1011_, new_n1007_, new_n1006_ );
or g874 ( new_n1012_, new_n1004_, keyIn_0_47 );
and g875 ( new_n1013_, new_n1012_, new_n1011_ );
and g876 ( new_n1014_, new_n1013_, new_n159_ );
or g877 ( new_n1015_, new_n1010_, new_n1014_ );
and g878 ( new_n1016_, new_n1015_, new_n1003_ );
or g879 ( new_n1017_, new_n1013_, new_n159_ );
or g880 ( new_n1018_, new_n1009_, N93 );
and g881 ( new_n1019_, new_n1017_, new_n1018_ );
and g882 ( new_n1020_, new_n1019_, keyIn_0_59 );
or g883 ( N747, new_n1016_, new_n1020_ );
and g884 ( new_n1022_, new_n587_, new_n834_ );
not g885 ( new_n1023_, new_n1022_ );
or g886 ( new_n1024_, new_n833_, new_n1023_ );
or g887 ( new_n1025_, new_n1024_, keyIn_0_39 );
not g888 ( new_n1026_, keyIn_0_39 );
and g889 ( new_n1027_, new_n853_, new_n1022_ );
or g890 ( new_n1028_, new_n1027_, new_n1026_ );
and g891 ( new_n1029_, new_n1025_, new_n1028_ );
or g892 ( new_n1030_, new_n1029_, new_n705_ );
and g893 ( new_n1031_, new_n1030_, keyIn_0_48 );
not g894 ( new_n1032_, keyIn_0_48 );
and g895 ( new_n1033_, new_n1027_, new_n1026_ );
and g896 ( new_n1034_, new_n1024_, keyIn_0_39 );
or g897 ( new_n1035_, new_n1034_, new_n1033_ );
and g898 ( new_n1036_, new_n1035_, new_n348_ );
and g899 ( new_n1037_, new_n1036_, new_n1032_ );
or g900 ( new_n1038_, new_n1031_, new_n1037_ );
and g901 ( new_n1039_, new_n1038_, N97 );
or g902 ( new_n1040_, new_n1036_, new_n1032_ );
or g903 ( new_n1041_, new_n1030_, keyIn_0_48 );
and g904 ( new_n1042_, new_n1041_, new_n1040_ );
and g905 ( new_n1043_, new_n1042_, new_n319_ );
or g906 ( new_n1044_, new_n1039_, new_n1043_ );
and g907 ( new_n1045_, new_n1044_, keyIn_0_60 );
not g908 ( new_n1046_, keyIn_0_60 );
or g909 ( new_n1047_, new_n1042_, new_n319_ );
or g910 ( new_n1048_, new_n1038_, N97 );
and g911 ( new_n1049_, new_n1048_, new_n1047_ );
and g912 ( new_n1050_, new_n1049_, new_n1046_ );
or g913 ( N748, new_n1045_, new_n1050_ );
not g914 ( new_n1052_, keyIn_0_49 );
or g915 ( new_n1053_, new_n1029_, new_n430_ );
and g916 ( new_n1054_, new_n1053_, new_n1052_ );
and g917 ( new_n1055_, new_n1035_, new_n706_ );
and g918 ( new_n1056_, new_n1055_, keyIn_0_49 );
or g919 ( new_n1057_, new_n1054_, new_n1056_ );
and g920 ( new_n1058_, new_n1057_, new_n418_ );
or g921 ( new_n1059_, new_n1055_, keyIn_0_49 );
or g922 ( new_n1060_, new_n1053_, new_n1052_ );
and g923 ( new_n1061_, new_n1060_, new_n1059_ );
and g924 ( new_n1062_, new_n1061_, N101 );
or g925 ( new_n1063_, new_n1058_, new_n1062_ );
and g926 ( new_n1064_, new_n1063_, keyIn_0_61 );
not g927 ( new_n1065_, keyIn_0_61 );
or g928 ( new_n1066_, new_n1061_, N101 );
or g929 ( new_n1067_, new_n1057_, new_n418_ );
and g930 ( new_n1068_, new_n1067_, new_n1066_ );
and g931 ( new_n1069_, new_n1068_, new_n1065_ );
or g932 ( N749, new_n1064_, new_n1069_ );
not g933 ( new_n1071_, keyIn_0_50 );
or g934 ( new_n1072_, new_n1029_, new_n678_ );
and g935 ( new_n1073_, new_n1072_, new_n1071_ );
and g936 ( new_n1074_, new_n1035_, new_n500_ );
and g937 ( new_n1075_, new_n1074_, keyIn_0_50 );
or g938 ( new_n1076_, new_n1073_, new_n1075_ );
and g939 ( new_n1077_, new_n1076_, new_n472_ );
or g940 ( new_n1078_, new_n1074_, keyIn_0_50 );
or g941 ( new_n1079_, new_n1072_, new_n1071_ );
and g942 ( new_n1080_, new_n1079_, new_n1078_ );
and g943 ( new_n1081_, new_n1080_, N105 );
or g944 ( new_n1082_, new_n1077_, new_n1081_ );
and g945 ( new_n1083_, new_n1082_, keyIn_0_62 );
not g946 ( new_n1084_, keyIn_0_62 );
or g947 ( new_n1085_, new_n1080_, N105 );
or g948 ( new_n1086_, new_n1076_, new_n472_ );
and g949 ( new_n1087_, new_n1086_, new_n1085_ );
and g950 ( new_n1088_, new_n1087_, new_n1084_ );
or g951 ( N750, new_n1083_, new_n1088_ );
not g952 ( new_n1090_, keyIn_0_63 );
or g953 ( new_n1091_, new_n1029_, new_n652_ );
and g954 ( new_n1092_, new_n1091_, keyIn_0_51 );
not g955 ( new_n1093_, keyIn_0_51 );
and g956 ( new_n1094_, new_n1035_, new_n679_ );
and g957 ( new_n1095_, new_n1094_, new_n1093_ );
or g958 ( new_n1096_, new_n1092_, new_n1095_ );
and g959 ( new_n1097_, new_n1096_, new_n509_ );
or g960 ( new_n1098_, new_n1094_, new_n1093_ );
or g961 ( new_n1099_, new_n1091_, keyIn_0_51 );
and g962 ( new_n1100_, new_n1099_, new_n1098_ );
and g963 ( new_n1101_, new_n1100_, N109 );
or g964 ( new_n1102_, new_n1097_, new_n1101_ );
and g965 ( new_n1103_, new_n1102_, new_n1090_ );
or g966 ( new_n1104_, new_n1100_, N109 );
or g967 ( new_n1105_, new_n1096_, new_n509_ );
and g968 ( new_n1106_, new_n1105_, new_n1104_ );
and g969 ( new_n1107_, new_n1106_, keyIn_0_63 );
or g970 ( N751, new_n1103_, new_n1107_ );
and g971 ( new_n1109_, new_n588_, new_n621_ );
and g972 ( new_n1110_, new_n853_, new_n1109_ );
and g973 ( new_n1111_, new_n1110_, new_n348_ );
not g974 ( new_n1112_, new_n1111_ );
and g975 ( new_n1113_, new_n1112_, N113 );
and g976 ( new_n1114_, new_n1111_, new_n320_ );
or g977 ( N752, new_n1113_, new_n1114_ );
and g978 ( new_n1116_, new_n1110_, new_n706_ );
not g979 ( new_n1117_, new_n1116_ );
and g980 ( new_n1118_, new_n1117_, N117 );
and g981 ( new_n1119_, new_n1116_, new_n419_ );
or g982 ( N753, new_n1118_, new_n1119_ );
and g983 ( new_n1121_, new_n1110_, new_n500_ );
not g984 ( new_n1122_, new_n1121_ );
and g985 ( new_n1123_, new_n1122_, N121 );
and g986 ( new_n1124_, new_n1121_, new_n470_ );
or g987 ( N754, new_n1123_, new_n1124_ );
and g988 ( new_n1126_, new_n1110_, new_n679_ );
not g989 ( new_n1127_, new_n1126_ );
and g990 ( new_n1128_, new_n1127_, N125 );
and g991 ( new_n1129_, new_n1126_, new_n546_ );
or g992 ( N755, new_n1128_, new_n1129_ );
endmodule