module add_mul_sub_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, operation_0_, operation_1_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, 
        Result_20_, Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, 
        Result_26_, Result_27_, Result_28_, Result_29_, Result_30_, Result_31_
 );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_,
         operation_0_, operation_1_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343;

  OR2_X1 U2155 ( .A1(n2123), .A2(n2124), .ZN(Result_9_) );
  AND2_X1 U2156 ( .A1(n2125), .A2(n2126), .ZN(n2123) );
  XOR2_X1 U2157 ( .A(n2127), .B(n2128), .Z(n2125) );
  OR2_X1 U2158 ( .A1(n2129), .A2(n2124), .ZN(Result_8_) );
  AND2_X1 U2159 ( .A1(n2126), .A2(n2130), .ZN(n2129) );
  XOR2_X1 U2160 ( .A(n2131), .B(n2132), .Z(n2130) );
  OR2_X1 U2161 ( .A1(n2133), .A2(n2124), .ZN(Result_7_) );
  AND2_X1 U2162 ( .A1(n2126), .A2(n2134), .ZN(n2133) );
  XOR2_X1 U2163 ( .A(n2135), .B(n2136), .Z(n2134) );
  OR2_X1 U2164 ( .A1(n2137), .A2(n2124), .ZN(Result_6_) );
  AND2_X1 U2165 ( .A1(n2126), .A2(n2138), .ZN(n2137) );
  XOR2_X1 U2166 ( .A(n2139), .B(n2140), .Z(n2138) );
  OR2_X1 U2167 ( .A1(n2141), .A2(n2124), .ZN(Result_5_) );
  AND2_X1 U2168 ( .A1(n2126), .A2(n2142), .ZN(n2141) );
  XOR2_X1 U2169 ( .A(n2143), .B(n2144), .Z(n2142) );
  OR2_X1 U2170 ( .A1(n2145), .A2(n2124), .ZN(Result_4_) );
  AND2_X1 U2171 ( .A1(n2126), .A2(n2146), .ZN(n2145) );
  XOR2_X1 U2172 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR2_X1 U2173 ( .A1(n2149), .A2(n2124), .ZN(Result_3_) );
  AND2_X1 U2174 ( .A1(n2126), .A2(n2150), .ZN(n2149) );
  XOR2_X1 U2175 ( .A(n2151), .B(n2152), .Z(n2150) );
  OR2_X1 U2176 ( .A1(n2153), .A2(n2154), .ZN(Result_31_) );
  AND2_X1 U2177 ( .A1(n2155), .A2(n2126), .ZN(n2154) );
  AND2_X1 U2178 ( .A1(n2156), .A2(n2157), .ZN(n2153) );
  OR3_X1 U2179 ( .A1(n2158), .A2(n2159), .A3(n2160), .ZN(n2157) );
  OR2_X1 U2180 ( .A1(n2161), .A2(n2162), .ZN(n2156) );
  OR3_X1 U2181 ( .A1(n2163), .A2(n2164), .A3(n2165), .ZN(Result_30_) );
  AND3_X1 U2182 ( .A1(n2162), .A2(a_14_), .A3(n2126), .ZN(n2165) );
  AND2_X1 U2183 ( .A1(n2166), .A2(n2167), .ZN(n2164) );
  OR2_X1 U2184 ( .A1(n2168), .A2(n2169), .ZN(n2166) );
  AND2_X1 U2185 ( .A1(a_14_), .A2(n2170), .ZN(n2169) );
  OR2_X1 U2186 ( .A1(n2171), .A2(n2172), .ZN(n2170) );
  AND2_X1 U2187 ( .A1(n2126), .A2(b_15_), .ZN(n2171) );
  AND2_X1 U2188 ( .A1(n2173), .A2(n2174), .ZN(n2168) );
  AND2_X1 U2189 ( .A1(b_14_), .A2(n2175), .ZN(n2163) );
  OR3_X1 U2190 ( .A1(n2176), .A2(n2177), .A3(n2178), .ZN(n2175) );
  AND2_X1 U2191 ( .A1(n2126), .A2(n2179), .ZN(n2178) );
  OR2_X1 U2192 ( .A1(n2161), .A2(n2180), .ZN(n2179) );
  AND2_X1 U2193 ( .A1(n2172), .A2(n2174), .ZN(n2177) );
  OR3_X1 U2194 ( .A1(n2181), .A2(n2182), .A3(n2183), .ZN(n2172) );
  AND2_X1 U2195 ( .A1(n2158), .A2(n2184), .ZN(n2183) );
  AND2_X1 U2196 ( .A1(n2159), .A2(n2185), .ZN(n2182) );
  AND2_X1 U2197 ( .A1(n2160), .A2(n2186), .ZN(n2181) );
  AND2_X1 U2198 ( .A1(a_14_), .A2(n2173), .ZN(n2176) );
  OR3_X1 U2199 ( .A1(n2187), .A2(n2188), .A3(n2189), .ZN(n2173) );
  AND2_X1 U2200 ( .A1(n2158), .A2(n2162), .ZN(n2189) );
  AND2_X1 U2201 ( .A1(n2159), .A2(n2161), .ZN(n2188) );
  AND2_X1 U2202 ( .A1(n2160), .A2(n2155), .ZN(n2187) );
  INV_X1 U2203 ( .A(n2186), .ZN(n2155) );
  OR2_X1 U2204 ( .A1(n2190), .A2(n2124), .ZN(Result_2_) );
  AND2_X1 U2205 ( .A1(n2126), .A2(n2191), .ZN(n2190) );
  XOR2_X1 U2206 ( .A(n2192), .B(n2193), .Z(n2191) );
  OR3_X1 U2207 ( .A1(n2194), .A2(n2195), .A3(n2196), .ZN(Result_29_) );
  AND2_X1 U2208 ( .A1(n2197), .A2(n2126), .ZN(n2196) );
  XOR2_X1 U2209 ( .A(n2198), .B(n2199), .Z(n2197) );
  XOR2_X1 U2210 ( .A(n2200), .B(n2201), .Z(n2199) );
  AND2_X1 U2211 ( .A1(n2202), .A2(n2203), .ZN(n2195) );
  OR3_X1 U2212 ( .A1(n2204), .A2(n2205), .A3(n2206), .ZN(n2203) );
  AND2_X1 U2213 ( .A1(n2158), .A2(n2207), .ZN(n2206) );
  AND2_X1 U2214 ( .A1(n2159), .A2(n2208), .ZN(n2205) );
  AND2_X1 U2215 ( .A1(n2160), .A2(n2209), .ZN(n2204) );
  INV_X1 U2216 ( .A(n2210), .ZN(n2209) );
  INV_X1 U2217 ( .A(n2211), .ZN(n2202) );
  AND2_X1 U2218 ( .A1(n2211), .A2(n2212), .ZN(n2194) );
  OR3_X1 U2219 ( .A1(n2213), .A2(n2214), .A3(n2215), .ZN(n2212) );
  AND2_X1 U2220 ( .A1(n2158), .A2(n2216), .ZN(n2215) );
  INV_X1 U2221 ( .A(n2207), .ZN(n2216) );
  AND2_X1 U2222 ( .A1(n2159), .A2(n2217), .ZN(n2214) );
  INV_X1 U2223 ( .A(n2208), .ZN(n2217) );
  AND2_X1 U2224 ( .A1(n2210), .A2(n2160), .ZN(n2213) );
  XNOR2_X1 U2225 ( .A(n2218), .B(b_13_), .ZN(n2211) );
  OR3_X1 U2226 ( .A1(n2219), .A2(n2220), .A3(n2221), .ZN(Result_28_) );
  AND2_X1 U2227 ( .A1(n2222), .A2(n2126), .ZN(n2221) );
  XNOR2_X1 U2228 ( .A(n2223), .B(n2224), .ZN(n2222) );
  XOR2_X1 U2229 ( .A(n2225), .B(n2226), .Z(n2224) );
  AND2_X1 U2230 ( .A1(n2227), .A2(n2228), .ZN(n2220) );
  OR3_X1 U2231 ( .A1(n2229), .A2(n2230), .A3(n2231), .ZN(n2228) );
  AND2_X1 U2232 ( .A1(n2158), .A2(n2232), .ZN(n2231) );
  AND2_X1 U2233 ( .A1(n2159), .A2(n2233), .ZN(n2230) );
  AND2_X1 U2234 ( .A1(n2234), .A2(n2160), .ZN(n2229) );
  INV_X1 U2235 ( .A(n2235), .ZN(n2234) );
  INV_X1 U2236 ( .A(n2236), .ZN(n2227) );
  AND2_X1 U2237 ( .A1(n2236), .A2(n2237), .ZN(n2219) );
  OR3_X1 U2238 ( .A1(n2238), .A2(n2239), .A3(n2240), .ZN(n2237) );
  AND2_X1 U2239 ( .A1(n2158), .A2(n2241), .ZN(n2240) );
  INV_X1 U2240 ( .A(n2232), .ZN(n2241) );
  AND2_X1 U2241 ( .A1(n2159), .A2(n2242), .ZN(n2239) );
  INV_X1 U2242 ( .A(n2233), .ZN(n2242) );
  AND2_X1 U2243 ( .A1(n2160), .A2(n2235), .ZN(n2238) );
  XNOR2_X1 U2244 ( .A(n2243), .B(b_12_), .ZN(n2236) );
  OR3_X1 U2245 ( .A1(n2244), .A2(n2245), .A3(n2246), .ZN(Result_27_) );
  AND2_X1 U2246 ( .A1(n2247), .A2(n2126), .ZN(n2246) );
  XNOR2_X1 U2247 ( .A(n2248), .B(n2249), .ZN(n2247) );
  XOR2_X1 U2248 ( .A(n2250), .B(n2251), .Z(n2249) );
  AND2_X1 U2249 ( .A1(n2252), .A2(n2253), .ZN(n2245) );
  OR3_X1 U2250 ( .A1(n2254), .A2(n2255), .A3(n2256), .ZN(n2253) );
  AND2_X1 U2251 ( .A1(n2158), .A2(n2257), .ZN(n2256) );
  AND2_X1 U2252 ( .A1(n2159), .A2(n2258), .ZN(n2255) );
  AND2_X1 U2253 ( .A1(n2259), .A2(n2160), .ZN(n2254) );
  INV_X1 U2254 ( .A(n2260), .ZN(n2259) );
  INV_X1 U2255 ( .A(n2261), .ZN(n2252) );
  AND2_X1 U2256 ( .A1(n2261), .A2(n2262), .ZN(n2244) );
  OR3_X1 U2257 ( .A1(n2263), .A2(n2264), .A3(n2265), .ZN(n2262) );
  AND2_X1 U2258 ( .A1(n2158), .A2(n2266), .ZN(n2265) );
  INV_X1 U2259 ( .A(n2257), .ZN(n2266) );
  AND2_X1 U2260 ( .A1(n2159), .A2(n2267), .ZN(n2264) );
  INV_X1 U2261 ( .A(n2258), .ZN(n2267) );
  AND2_X1 U2262 ( .A1(n2160), .A2(n2260), .ZN(n2263) );
  XNOR2_X1 U2263 ( .A(n2268), .B(b_11_), .ZN(n2261) );
  OR3_X1 U2264 ( .A1(n2269), .A2(n2270), .A3(n2271), .ZN(Result_26_) );
  AND2_X1 U2265 ( .A1(n2272), .A2(n2126), .ZN(n2271) );
  XNOR2_X1 U2266 ( .A(n2273), .B(n2274), .ZN(n2272) );
  XOR2_X1 U2267 ( .A(n2275), .B(n2276), .Z(n2274) );
  AND2_X1 U2268 ( .A1(n2277), .A2(n2278), .ZN(n2270) );
  OR3_X1 U2269 ( .A1(n2279), .A2(n2280), .A3(n2281), .ZN(n2278) );
  AND2_X1 U2270 ( .A1(n2158), .A2(n2282), .ZN(n2281) );
  AND2_X1 U2271 ( .A1(n2159), .A2(n2283), .ZN(n2280) );
  AND2_X1 U2272 ( .A1(n2284), .A2(n2160), .ZN(n2279) );
  INV_X1 U2273 ( .A(n2285), .ZN(n2284) );
  INV_X1 U2274 ( .A(n2286), .ZN(n2277) );
  AND2_X1 U2275 ( .A1(n2286), .A2(n2287), .ZN(n2269) );
  OR3_X1 U2276 ( .A1(n2288), .A2(n2289), .A3(n2290), .ZN(n2287) );
  AND2_X1 U2277 ( .A1(n2158), .A2(n2291), .ZN(n2290) );
  INV_X1 U2278 ( .A(n2282), .ZN(n2291) );
  AND2_X1 U2279 ( .A1(n2159), .A2(n2292), .ZN(n2289) );
  INV_X1 U2280 ( .A(n2283), .ZN(n2292) );
  AND2_X1 U2281 ( .A1(n2160), .A2(n2285), .ZN(n2288) );
  XNOR2_X1 U2282 ( .A(n2293), .B(b_10_), .ZN(n2286) );
  OR3_X1 U2283 ( .A1(n2294), .A2(n2295), .A3(n2296), .ZN(Result_25_) );
  AND2_X1 U2284 ( .A1(n2297), .A2(n2126), .ZN(n2296) );
  XNOR2_X1 U2285 ( .A(n2298), .B(n2299), .ZN(n2297) );
  XOR2_X1 U2286 ( .A(n2300), .B(n2301), .Z(n2299) );
  AND2_X1 U2287 ( .A1(n2302), .A2(n2303), .ZN(n2295) );
  OR3_X1 U2288 ( .A1(n2304), .A2(n2305), .A3(n2306), .ZN(n2303) );
  AND2_X1 U2289 ( .A1(n2158), .A2(n2307), .ZN(n2306) );
  AND2_X1 U2290 ( .A1(n2159), .A2(n2308), .ZN(n2305) );
  AND2_X1 U2291 ( .A1(n2309), .A2(n2160), .ZN(n2304) );
  INV_X1 U2292 ( .A(n2310), .ZN(n2309) );
  INV_X1 U2293 ( .A(n2311), .ZN(n2302) );
  AND2_X1 U2294 ( .A1(n2311), .A2(n2312), .ZN(n2294) );
  OR3_X1 U2295 ( .A1(n2313), .A2(n2314), .A3(n2315), .ZN(n2312) );
  AND2_X1 U2296 ( .A1(n2158), .A2(n2316), .ZN(n2315) );
  INV_X1 U2297 ( .A(n2307), .ZN(n2316) );
  AND2_X1 U2298 ( .A1(n2159), .A2(n2317), .ZN(n2314) );
  INV_X1 U2299 ( .A(n2308), .ZN(n2317) );
  AND2_X1 U2300 ( .A1(n2160), .A2(n2310), .ZN(n2313) );
  XNOR2_X1 U2301 ( .A(n2318), .B(b_9_), .ZN(n2311) );
  OR3_X1 U2302 ( .A1(n2319), .A2(n2320), .A3(n2321), .ZN(Result_24_) );
  AND2_X1 U2303 ( .A1(n2322), .A2(n2126), .ZN(n2321) );
  XNOR2_X1 U2304 ( .A(n2323), .B(n2324), .ZN(n2322) );
  XOR2_X1 U2305 ( .A(n2325), .B(n2326), .Z(n2324) );
  AND2_X1 U2306 ( .A1(n2327), .A2(n2328), .ZN(n2320) );
  OR3_X1 U2307 ( .A1(n2329), .A2(n2330), .A3(n2331), .ZN(n2328) );
  AND2_X1 U2308 ( .A1(n2158), .A2(n2332), .ZN(n2331) );
  INV_X1 U2309 ( .A(n2333), .ZN(n2332) );
  AND2_X1 U2310 ( .A1(n2159), .A2(n2334), .ZN(n2330) );
  INV_X1 U2311 ( .A(n2335), .ZN(n2334) );
  AND2_X1 U2312 ( .A1(n2160), .A2(n2336), .ZN(n2329) );
  AND2_X1 U2313 ( .A1(n2337), .A2(n2338), .ZN(n2319) );
  INV_X1 U2314 ( .A(n2327), .ZN(n2338) );
  AND2_X1 U2315 ( .A1(n2339), .A2(n2340), .ZN(n2327) );
  OR2_X1 U2316 ( .A1(a_8_), .A2(b_8_), .ZN(n2339) );
  OR3_X1 U2317 ( .A1(n2341), .A2(n2342), .A3(n2343), .ZN(n2337) );
  AND2_X1 U2318 ( .A1(n2158), .A2(n2333), .ZN(n2343) );
  AND2_X1 U2319 ( .A1(n2159), .A2(n2335), .ZN(n2342) );
  AND2_X1 U2320 ( .A1(n2344), .A2(n2160), .ZN(n2341) );
  INV_X1 U2321 ( .A(n2336), .ZN(n2344) );
  OR3_X1 U2322 ( .A1(n2345), .A2(n2346), .A3(n2347), .ZN(Result_23_) );
  AND2_X1 U2323 ( .A1(n2348), .A2(n2126), .ZN(n2347) );
  XNOR2_X1 U2324 ( .A(n2349), .B(n2350), .ZN(n2348) );
  XOR2_X1 U2325 ( .A(n2351), .B(n2352), .Z(n2350) );
  AND2_X1 U2326 ( .A1(n2353), .A2(n2354), .ZN(n2346) );
  OR3_X1 U2327 ( .A1(n2355), .A2(n2356), .A3(n2357), .ZN(n2354) );
  AND2_X1 U2328 ( .A1(n2158), .A2(n2358), .ZN(n2357) );
  INV_X1 U2329 ( .A(n2359), .ZN(n2358) );
  AND2_X1 U2330 ( .A1(n2159), .A2(n2360), .ZN(n2356) );
  INV_X1 U2331 ( .A(n2361), .ZN(n2360) );
  AND2_X1 U2332 ( .A1(n2160), .A2(n2362), .ZN(n2355) );
  AND2_X1 U2333 ( .A1(n2363), .A2(n2364), .ZN(n2345) );
  INV_X1 U2334 ( .A(n2353), .ZN(n2364) );
  AND2_X1 U2335 ( .A1(n2365), .A2(n2366), .ZN(n2353) );
  OR2_X1 U2336 ( .A1(a_7_), .A2(b_7_), .ZN(n2365) );
  OR3_X1 U2337 ( .A1(n2367), .A2(n2368), .A3(n2369), .ZN(n2363) );
  AND2_X1 U2338 ( .A1(n2158), .A2(n2359), .ZN(n2369) );
  AND2_X1 U2339 ( .A1(n2159), .A2(n2361), .ZN(n2368) );
  AND2_X1 U2340 ( .A1(n2370), .A2(n2160), .ZN(n2367) );
  INV_X1 U2341 ( .A(n2362), .ZN(n2370) );
  OR3_X1 U2342 ( .A1(n2371), .A2(n2372), .A3(n2373), .ZN(Result_22_) );
  AND2_X1 U2343 ( .A1(n2374), .A2(n2126), .ZN(n2373) );
  XNOR2_X1 U2344 ( .A(n2375), .B(n2376), .ZN(n2374) );
  XOR2_X1 U2345 ( .A(n2377), .B(n2378), .Z(n2376) );
  AND2_X1 U2346 ( .A1(n2379), .A2(n2380), .ZN(n2372) );
  OR3_X1 U2347 ( .A1(n2381), .A2(n2382), .A3(n2383), .ZN(n2380) );
  AND2_X1 U2348 ( .A1(n2158), .A2(n2384), .ZN(n2383) );
  INV_X1 U2349 ( .A(n2385), .ZN(n2384) );
  AND2_X1 U2350 ( .A1(n2159), .A2(n2386), .ZN(n2382) );
  INV_X1 U2351 ( .A(n2387), .ZN(n2386) );
  AND2_X1 U2352 ( .A1(n2160), .A2(n2388), .ZN(n2381) );
  AND2_X1 U2353 ( .A1(n2389), .A2(n2390), .ZN(n2371) );
  INV_X1 U2354 ( .A(n2379), .ZN(n2390) );
  AND2_X1 U2355 ( .A1(n2391), .A2(n2392), .ZN(n2379) );
  OR2_X1 U2356 ( .A1(a_6_), .A2(b_6_), .ZN(n2391) );
  OR3_X1 U2357 ( .A1(n2393), .A2(n2394), .A3(n2395), .ZN(n2389) );
  AND2_X1 U2358 ( .A1(n2158), .A2(n2385), .ZN(n2395) );
  AND2_X1 U2359 ( .A1(n2159), .A2(n2387), .ZN(n2394) );
  AND2_X1 U2360 ( .A1(n2396), .A2(n2160), .ZN(n2393) );
  INV_X1 U2361 ( .A(n2388), .ZN(n2396) );
  OR3_X1 U2362 ( .A1(n2397), .A2(n2398), .A3(n2399), .ZN(Result_21_) );
  AND2_X1 U2363 ( .A1(n2400), .A2(n2126), .ZN(n2399) );
  XNOR2_X1 U2364 ( .A(n2401), .B(n2402), .ZN(n2400) );
  XOR2_X1 U2365 ( .A(n2403), .B(n2404), .Z(n2402) );
  AND2_X1 U2366 ( .A1(n2405), .A2(n2406), .ZN(n2398) );
  OR3_X1 U2367 ( .A1(n2407), .A2(n2408), .A3(n2409), .ZN(n2406) );
  AND2_X1 U2368 ( .A1(n2158), .A2(n2410), .ZN(n2409) );
  INV_X1 U2369 ( .A(n2411), .ZN(n2410) );
  AND2_X1 U2370 ( .A1(n2159), .A2(n2412), .ZN(n2408) );
  INV_X1 U2371 ( .A(n2413), .ZN(n2412) );
  AND2_X1 U2372 ( .A1(n2160), .A2(n2414), .ZN(n2407) );
  AND2_X1 U2373 ( .A1(n2415), .A2(n2416), .ZN(n2397) );
  INV_X1 U2374 ( .A(n2405), .ZN(n2416) );
  AND2_X1 U2375 ( .A1(n2417), .A2(n2418), .ZN(n2405) );
  OR2_X1 U2376 ( .A1(a_5_), .A2(b_5_), .ZN(n2417) );
  OR3_X1 U2377 ( .A1(n2419), .A2(n2420), .A3(n2421), .ZN(n2415) );
  AND2_X1 U2378 ( .A1(n2158), .A2(n2411), .ZN(n2421) );
  AND2_X1 U2379 ( .A1(n2159), .A2(n2413), .ZN(n2420) );
  AND2_X1 U2380 ( .A1(n2422), .A2(n2160), .ZN(n2419) );
  INV_X1 U2381 ( .A(n2414), .ZN(n2422) );
  OR3_X1 U2382 ( .A1(n2423), .A2(n2424), .A3(n2425), .ZN(Result_20_) );
  AND2_X1 U2383 ( .A1(n2426), .A2(n2126), .ZN(n2425) );
  XNOR2_X1 U2384 ( .A(n2427), .B(n2428), .ZN(n2426) );
  XOR2_X1 U2385 ( .A(n2429), .B(n2430), .Z(n2428) );
  AND2_X1 U2386 ( .A1(n2431), .A2(n2432), .ZN(n2424) );
  OR3_X1 U2387 ( .A1(n2433), .A2(n2434), .A3(n2435), .ZN(n2432) );
  AND2_X1 U2388 ( .A1(n2158), .A2(n2436), .ZN(n2435) );
  INV_X1 U2389 ( .A(n2437), .ZN(n2436) );
  AND2_X1 U2390 ( .A1(n2159), .A2(n2438), .ZN(n2434) );
  INV_X1 U2391 ( .A(n2439), .ZN(n2438) );
  AND2_X1 U2392 ( .A1(n2160), .A2(n2440), .ZN(n2433) );
  AND2_X1 U2393 ( .A1(n2441), .A2(n2442), .ZN(n2423) );
  INV_X1 U2394 ( .A(n2431), .ZN(n2442) );
  AND2_X1 U2395 ( .A1(n2443), .A2(n2444), .ZN(n2431) );
  OR2_X1 U2396 ( .A1(a_4_), .A2(b_4_), .ZN(n2443) );
  OR3_X1 U2397 ( .A1(n2445), .A2(n2446), .A3(n2447), .ZN(n2441) );
  AND2_X1 U2398 ( .A1(n2158), .A2(n2437), .ZN(n2447) );
  AND2_X1 U2399 ( .A1(n2159), .A2(n2439), .ZN(n2446) );
  AND2_X1 U2400 ( .A1(n2448), .A2(n2160), .ZN(n2445) );
  INV_X1 U2401 ( .A(n2440), .ZN(n2448) );
  OR2_X1 U2402 ( .A1(n2449), .A2(n2124), .ZN(Result_1_) );
  AND2_X1 U2403 ( .A1(n2126), .A2(n2450), .ZN(n2449) );
  XOR2_X1 U2404 ( .A(n2451), .B(n2452), .Z(n2450) );
  AND2_X1 U2405 ( .A1(n2453), .A2(n2454), .ZN(n2452) );
  OR2_X1 U2406 ( .A1(n2455), .A2(n2456), .ZN(n2454) );
  AND2_X1 U2407 ( .A1(n2457), .A2(n2458), .ZN(n2455) );
  INV_X1 U2408 ( .A(n2459), .ZN(n2453) );
  OR3_X1 U2409 ( .A1(n2460), .A2(n2461), .A3(n2462), .ZN(Result_19_) );
  AND2_X1 U2410 ( .A1(n2463), .A2(n2126), .ZN(n2462) );
  XNOR2_X1 U2411 ( .A(n2464), .B(n2465), .ZN(n2463) );
  XOR2_X1 U2412 ( .A(n2466), .B(n2467), .Z(n2465) );
  AND2_X1 U2413 ( .A1(n2468), .A2(n2469), .ZN(n2461) );
  OR3_X1 U2414 ( .A1(n2470), .A2(n2471), .A3(n2472), .ZN(n2469) );
  AND2_X1 U2415 ( .A1(n2158), .A2(n2473), .ZN(n2472) );
  INV_X1 U2416 ( .A(n2474), .ZN(n2473) );
  AND2_X1 U2417 ( .A1(n2159), .A2(n2475), .ZN(n2471) );
  INV_X1 U2418 ( .A(n2476), .ZN(n2475) );
  AND2_X1 U2419 ( .A1(n2160), .A2(n2477), .ZN(n2470) );
  AND2_X1 U2420 ( .A1(n2478), .A2(n2479), .ZN(n2460) );
  INV_X1 U2421 ( .A(n2468), .ZN(n2479) );
  AND2_X1 U2422 ( .A1(n2480), .A2(n2481), .ZN(n2468) );
  OR2_X1 U2423 ( .A1(a_3_), .A2(b_3_), .ZN(n2480) );
  OR3_X1 U2424 ( .A1(n2482), .A2(n2483), .A3(n2484), .ZN(n2478) );
  AND2_X1 U2425 ( .A1(n2158), .A2(n2474), .ZN(n2484) );
  AND2_X1 U2426 ( .A1(n2159), .A2(n2476), .ZN(n2483) );
  AND2_X1 U2427 ( .A1(n2485), .A2(n2160), .ZN(n2482) );
  INV_X1 U2428 ( .A(n2477), .ZN(n2485) );
  OR3_X1 U2429 ( .A1(n2486), .A2(n2487), .A3(n2488), .ZN(Result_18_) );
  AND2_X1 U2430 ( .A1(n2489), .A2(n2126), .ZN(n2488) );
  XNOR2_X1 U2431 ( .A(n2490), .B(n2491), .ZN(n2489) );
  XOR2_X1 U2432 ( .A(n2492), .B(n2493), .Z(n2491) );
  AND2_X1 U2433 ( .A1(n2494), .A2(n2495), .ZN(n2487) );
  OR3_X1 U2434 ( .A1(n2496), .A2(n2497), .A3(n2498), .ZN(n2495) );
  AND2_X1 U2435 ( .A1(n2158), .A2(n2499), .ZN(n2498) );
  INV_X1 U2436 ( .A(n2500), .ZN(n2499) );
  AND2_X1 U2437 ( .A1(n2159), .A2(n2501), .ZN(n2497) );
  INV_X1 U2438 ( .A(n2502), .ZN(n2501) );
  AND2_X1 U2439 ( .A1(n2160), .A2(n2503), .ZN(n2496) );
  AND2_X1 U2440 ( .A1(n2504), .A2(n2505), .ZN(n2486) );
  INV_X1 U2441 ( .A(n2494), .ZN(n2505) );
  AND2_X1 U2442 ( .A1(n2506), .A2(n2507), .ZN(n2494) );
  OR2_X1 U2443 ( .A1(a_2_), .A2(b_2_), .ZN(n2506) );
  OR3_X1 U2444 ( .A1(n2508), .A2(n2509), .A3(n2510), .ZN(n2504) );
  AND2_X1 U2445 ( .A1(n2158), .A2(n2500), .ZN(n2510) );
  AND2_X1 U2446 ( .A1(n2159), .A2(n2502), .ZN(n2509) );
  AND2_X1 U2447 ( .A1(n2511), .A2(n2160), .ZN(n2508) );
  INV_X1 U2448 ( .A(n2503), .ZN(n2511) );
  OR3_X1 U2449 ( .A1(n2512), .A2(n2513), .A3(n2514), .ZN(Result_17_) );
  AND2_X1 U2450 ( .A1(n2515), .A2(n2126), .ZN(n2514) );
  XNOR2_X1 U2451 ( .A(n2516), .B(n2517), .ZN(n2515) );
  XOR2_X1 U2452 ( .A(n2518), .B(n2519), .Z(n2517) );
  AND2_X1 U2453 ( .A1(n2520), .A2(n2521), .ZN(n2513) );
  OR3_X1 U2454 ( .A1(n2522), .A2(n2523), .A3(n2524), .ZN(n2521) );
  AND2_X1 U2455 ( .A1(n2158), .A2(n2525), .ZN(n2524) );
  INV_X1 U2456 ( .A(n2526), .ZN(n2525) );
  AND2_X1 U2457 ( .A1(n2159), .A2(n2527), .ZN(n2523) );
  INV_X1 U2458 ( .A(n2528), .ZN(n2527) );
  AND2_X1 U2459 ( .A1(n2160), .A2(n2529), .ZN(n2522) );
  AND2_X1 U2460 ( .A1(n2530), .A2(n2531), .ZN(n2512) );
  INV_X1 U2461 ( .A(n2520), .ZN(n2531) );
  AND2_X1 U2462 ( .A1(n2532), .A2(n2533), .ZN(n2520) );
  OR2_X1 U2463 ( .A1(a_1_), .A2(b_1_), .ZN(n2532) );
  OR3_X1 U2464 ( .A1(n2534), .A2(n2535), .A3(n2536), .ZN(n2530) );
  AND2_X1 U2465 ( .A1(n2158), .A2(n2526), .ZN(n2536) );
  AND2_X1 U2466 ( .A1(n2159), .A2(n2528), .ZN(n2535) );
  AND2_X1 U2467 ( .A1(n2537), .A2(n2160), .ZN(n2534) );
  INV_X1 U2468 ( .A(n2529), .ZN(n2537) );
  OR3_X1 U2469 ( .A1(n2538), .A2(n2539), .A3(n2540), .ZN(Result_16_) );
  AND2_X1 U2470 ( .A1(n2541), .A2(n2126), .ZN(n2540) );
  XNOR2_X1 U2471 ( .A(n2542), .B(n2543), .ZN(n2541) );
  XOR2_X1 U2472 ( .A(n2544), .B(n2545), .Z(n2543) );
  AND2_X1 U2473 ( .A1(n2546), .A2(n2547), .ZN(n2539) );
  OR3_X1 U2474 ( .A1(n2548), .A2(n2549), .A3(n2550), .ZN(n2546) );
  AND2_X1 U2475 ( .A1(n2551), .A2(n2158), .ZN(n2550) );
  AND2_X1 U2476 ( .A1(n2159), .A2(n2552), .ZN(n2549) );
  INV_X1 U2477 ( .A(n2553), .ZN(n2552) );
  AND2_X1 U2478 ( .A1(n2160), .A2(n2554), .ZN(n2548) );
  AND2_X1 U2479 ( .A1(n2555), .A2(n2556), .ZN(n2538) );
  OR3_X1 U2480 ( .A1(n2557), .A2(n2558), .A3(n2559), .ZN(n2556) );
  AND2_X1 U2481 ( .A1(n2158), .A2(n2560), .ZN(n2559) );
  AND2_X1 U2482 ( .A1(n2159), .A2(n2553), .ZN(n2558) );
  AND2_X1 U2483 ( .A1(n2561), .A2(n2160), .ZN(n2557) );
  AND2_X1 U2484 ( .A1(n2562), .A2(n2563), .ZN(n2160) );
  INV_X1 U2485 ( .A(n2554), .ZN(n2561) );
  OR2_X1 U2486 ( .A1(n2564), .A2(n2565), .ZN(n2554) );
  AND2_X1 U2487 ( .A1(n2566), .A2(n2567), .ZN(n2565) );
  AND2_X1 U2488 ( .A1(n2529), .A2(n2533), .ZN(n2564) );
  OR2_X1 U2489 ( .A1(n2568), .A2(n2569), .ZN(n2529) );
  AND2_X1 U2490 ( .A1(n2570), .A2(n2571), .ZN(n2569) );
  AND2_X1 U2491 ( .A1(n2503), .A2(n2507), .ZN(n2568) );
  OR2_X1 U2492 ( .A1(n2572), .A2(n2573), .ZN(n2503) );
  AND2_X1 U2493 ( .A1(n2574), .A2(n2575), .ZN(n2573) );
  AND2_X1 U2494 ( .A1(n2477), .A2(n2481), .ZN(n2572) );
  OR2_X1 U2495 ( .A1(n2576), .A2(n2577), .ZN(n2477) );
  AND2_X1 U2496 ( .A1(n2578), .A2(n2579), .ZN(n2577) );
  AND2_X1 U2497 ( .A1(n2440), .A2(n2444), .ZN(n2576) );
  OR2_X1 U2498 ( .A1(n2580), .A2(n2581), .ZN(n2440) );
  AND2_X1 U2499 ( .A1(n2582), .A2(n2583), .ZN(n2581) );
  AND2_X1 U2500 ( .A1(n2414), .A2(n2418), .ZN(n2580) );
  OR2_X1 U2501 ( .A1(n2584), .A2(n2585), .ZN(n2414) );
  AND2_X1 U2502 ( .A1(n2586), .A2(n2587), .ZN(n2585) );
  AND2_X1 U2503 ( .A1(n2388), .A2(n2392), .ZN(n2584) );
  OR2_X1 U2504 ( .A1(n2588), .A2(n2589), .ZN(n2388) );
  AND2_X1 U2505 ( .A1(n2590), .A2(n2591), .ZN(n2589) );
  AND2_X1 U2506 ( .A1(n2362), .A2(n2366), .ZN(n2588) );
  OR2_X1 U2507 ( .A1(n2592), .A2(n2593), .ZN(n2362) );
  AND2_X1 U2508 ( .A1(n2594), .A2(n2595), .ZN(n2593) );
  AND2_X1 U2509 ( .A1(n2336), .A2(n2340), .ZN(n2592) );
  OR2_X1 U2510 ( .A1(n2596), .A2(n2597), .ZN(n2336) );
  AND2_X1 U2511 ( .A1(n2318), .A2(n2598), .ZN(n2597) );
  AND2_X1 U2512 ( .A1(n2310), .A2(n2599), .ZN(n2596) );
  OR2_X1 U2513 ( .A1(n2600), .A2(n2601), .ZN(n2310) );
  AND2_X1 U2514 ( .A1(n2293), .A2(n2602), .ZN(n2601) );
  AND2_X1 U2515 ( .A1(n2285), .A2(n2603), .ZN(n2600) );
  OR2_X1 U2516 ( .A1(n2604), .A2(n2605), .ZN(n2285) );
  AND2_X1 U2517 ( .A1(n2268), .A2(n2606), .ZN(n2605) );
  AND2_X1 U2518 ( .A1(n2260), .A2(n2607), .ZN(n2604) );
  OR2_X1 U2519 ( .A1(n2608), .A2(n2609), .ZN(n2260) );
  AND2_X1 U2520 ( .A1(n2243), .A2(n2610), .ZN(n2609) );
  AND2_X1 U2521 ( .A1(n2235), .A2(n2611), .ZN(n2608) );
  OR2_X1 U2522 ( .A1(n2612), .A2(n2613), .ZN(n2235) );
  AND2_X1 U2523 ( .A1(n2218), .A2(n2614), .ZN(n2613) );
  AND2_X1 U2524 ( .A1(n2210), .A2(n2615), .ZN(n2612) );
  AND2_X1 U2525 ( .A1(n2616), .A2(n2617), .ZN(n2210) );
  OR2_X1 U2526 ( .A1(n2167), .A2(n2618), .ZN(n2617) );
  AND2_X1 U2527 ( .A1(n2174), .A2(n2186), .ZN(n2618) );
  OR2_X1 U2528 ( .A1(n2619), .A2(n2620), .ZN(n2186) );
  INV_X1 U2529 ( .A(n2547), .ZN(n2555) );
  OR2_X1 U2530 ( .A1(n2621), .A2(n2622), .ZN(n2547) );
  INV_X1 U2531 ( .A(n2623), .ZN(n2621) );
  OR2_X1 U2532 ( .A1(n2624), .A2(n2124), .ZN(Result_15_) );
  AND2_X1 U2533 ( .A1(n2126), .A2(n2625), .ZN(n2624) );
  XOR2_X1 U2534 ( .A(n2626), .B(n2627), .Z(n2625) );
  OR2_X1 U2535 ( .A1(n2628), .A2(n2124), .ZN(Result_14_) );
  AND3_X1 U2536 ( .A1(n2629), .A2(n2630), .A3(n2126), .ZN(n2628) );
  OR2_X1 U2537 ( .A1(n2631), .A2(n2632), .ZN(n2629) );
  AND2_X1 U2538 ( .A1(n2626), .A2(n2627), .ZN(n2631) );
  OR2_X1 U2539 ( .A1(n2633), .A2(n2124), .ZN(Result_13_) );
  AND2_X1 U2540 ( .A1(n2126), .A2(n2634), .ZN(n2633) );
  XOR2_X1 U2541 ( .A(n2630), .B(n2635), .Z(n2634) );
  OR2_X1 U2542 ( .A1(n2636), .A2(n2637), .ZN(n2635) );
  AND2_X1 U2543 ( .A1(n2638), .A2(n2639), .ZN(n2636) );
  OR2_X1 U2544 ( .A1(n2640), .A2(n2641), .ZN(n2638) );
  INV_X1 U2545 ( .A(n2642), .ZN(n2630) );
  OR2_X1 U2546 ( .A1(n2643), .A2(n2124), .ZN(Result_12_) );
  AND2_X1 U2547 ( .A1(n2644), .A2(n2126), .ZN(n2643) );
  XOR2_X1 U2548 ( .A(n2645), .B(n2646), .Z(n2644) );
  AND2_X1 U2549 ( .A1(n2647), .A2(n2648), .ZN(n2646) );
  OR2_X1 U2550 ( .A1(n2649), .A2(n2650), .ZN(n2648) );
  INV_X1 U2551 ( .A(n2651), .ZN(n2647) );
  OR2_X1 U2552 ( .A1(n2652), .A2(n2124), .ZN(Result_11_) );
  AND2_X1 U2553 ( .A1(n2653), .A2(n2126), .ZN(n2652) );
  XOR2_X1 U2554 ( .A(n2654), .B(n2655), .Z(n2653) );
  AND2_X1 U2555 ( .A1(n2656), .A2(n2657), .ZN(n2655) );
  OR2_X1 U2556 ( .A1(n2658), .A2(n2659), .ZN(n2657) );
  AND2_X1 U2557 ( .A1(n2660), .A2(n2661), .ZN(n2658) );
  INV_X1 U2558 ( .A(n2662), .ZN(n2656) );
  OR2_X1 U2559 ( .A1(n2663), .A2(n2124), .ZN(Result_10_) );
  AND2_X1 U2560 ( .A1(n2664), .A2(n2126), .ZN(n2663) );
  XOR2_X1 U2561 ( .A(n2665), .B(n2666), .Z(n2664) );
  AND2_X1 U2562 ( .A1(n2667), .A2(n2668), .ZN(n2666) );
  OR2_X1 U2563 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  AND2_X1 U2564 ( .A1(n2671), .A2(n2672), .ZN(n2670) );
  INV_X1 U2565 ( .A(n2673), .ZN(n2667) );
  OR2_X1 U2566 ( .A1(n2674), .A2(n2124), .ZN(Result_0_) );
  OR2_X1 U2567 ( .A1(n2675), .A2(n2676), .ZN(n2124) );
  AND2_X1 U2568 ( .A1(n2158), .A2(n2677), .ZN(n2676) );
  INV_X1 U2569 ( .A(n2678), .ZN(n2677) );
  AND2_X1 U2570 ( .A1(n2679), .A2(n2623), .ZN(n2678) );
  OR2_X1 U2571 ( .A1(n2551), .A2(n2622), .ZN(n2679) );
  INV_X1 U2572 ( .A(n2560), .ZN(n2551) );
  OR2_X1 U2573 ( .A1(n2680), .A2(n2681), .ZN(n2560) );
  AND2_X1 U2574 ( .A1(n2526), .A2(n2566), .ZN(n2681) );
  AND2_X1 U2575 ( .A1(b_1_), .A2(n2682), .ZN(n2680) );
  OR2_X1 U2576 ( .A1(n2566), .A2(n2526), .ZN(n2682) );
  OR2_X1 U2577 ( .A1(n2683), .A2(n2684), .ZN(n2526) );
  AND2_X1 U2578 ( .A1(n2500), .A2(n2570), .ZN(n2684) );
  AND2_X1 U2579 ( .A1(b_2_), .A2(n2685), .ZN(n2683) );
  OR2_X1 U2580 ( .A1(n2570), .A2(n2500), .ZN(n2685) );
  OR2_X1 U2581 ( .A1(n2686), .A2(n2687), .ZN(n2500) );
  AND2_X1 U2582 ( .A1(n2474), .A2(n2574), .ZN(n2687) );
  AND2_X1 U2583 ( .A1(b_3_), .A2(n2688), .ZN(n2686) );
  OR2_X1 U2584 ( .A1(n2574), .A2(n2474), .ZN(n2688) );
  OR2_X1 U2585 ( .A1(n2689), .A2(n2690), .ZN(n2474) );
  AND2_X1 U2586 ( .A1(n2437), .A2(n2578), .ZN(n2690) );
  AND2_X1 U2587 ( .A1(b_4_), .A2(n2691), .ZN(n2689) );
  OR2_X1 U2588 ( .A1(n2578), .A2(n2437), .ZN(n2691) );
  OR2_X1 U2589 ( .A1(n2692), .A2(n2693), .ZN(n2437) );
  AND2_X1 U2590 ( .A1(n2411), .A2(n2582), .ZN(n2693) );
  AND2_X1 U2591 ( .A1(b_5_), .A2(n2694), .ZN(n2692) );
  OR2_X1 U2592 ( .A1(n2582), .A2(n2411), .ZN(n2694) );
  OR2_X1 U2593 ( .A1(n2695), .A2(n2696), .ZN(n2411) );
  AND2_X1 U2594 ( .A1(n2385), .A2(n2586), .ZN(n2696) );
  AND2_X1 U2595 ( .A1(b_6_), .A2(n2697), .ZN(n2695) );
  OR2_X1 U2596 ( .A1(n2586), .A2(n2385), .ZN(n2697) );
  OR2_X1 U2597 ( .A1(n2698), .A2(n2699), .ZN(n2385) );
  AND2_X1 U2598 ( .A1(n2359), .A2(n2590), .ZN(n2699) );
  AND2_X1 U2599 ( .A1(b_7_), .A2(n2700), .ZN(n2698) );
  OR2_X1 U2600 ( .A1(n2590), .A2(n2359), .ZN(n2700) );
  OR2_X1 U2601 ( .A1(n2701), .A2(n2702), .ZN(n2359) );
  AND2_X1 U2602 ( .A1(n2333), .A2(n2594), .ZN(n2702) );
  AND2_X1 U2603 ( .A1(b_8_), .A2(n2703), .ZN(n2701) );
  OR2_X1 U2604 ( .A1(n2594), .A2(n2333), .ZN(n2703) );
  OR2_X1 U2605 ( .A1(n2704), .A2(n2705), .ZN(n2333) );
  AND2_X1 U2606 ( .A1(n2307), .A2(n2318), .ZN(n2705) );
  AND2_X1 U2607 ( .A1(b_9_), .A2(n2706), .ZN(n2704) );
  OR2_X1 U2608 ( .A1(n2318), .A2(n2307), .ZN(n2706) );
  OR2_X1 U2609 ( .A1(n2707), .A2(n2708), .ZN(n2307) );
  AND2_X1 U2610 ( .A1(n2282), .A2(n2293), .ZN(n2708) );
  AND2_X1 U2611 ( .A1(b_10_), .A2(n2709), .ZN(n2707) );
  OR2_X1 U2612 ( .A1(n2293), .A2(n2282), .ZN(n2709) );
  OR2_X1 U2613 ( .A1(n2710), .A2(n2711), .ZN(n2282) );
  AND2_X1 U2614 ( .A1(n2257), .A2(n2268), .ZN(n2711) );
  AND2_X1 U2615 ( .A1(b_11_), .A2(n2712), .ZN(n2710) );
  OR2_X1 U2616 ( .A1(n2268), .A2(n2257), .ZN(n2712) );
  OR2_X1 U2617 ( .A1(n2713), .A2(n2714), .ZN(n2257) );
  AND2_X1 U2618 ( .A1(n2232), .A2(n2243), .ZN(n2714) );
  AND2_X1 U2619 ( .A1(b_12_), .A2(n2715), .ZN(n2713) );
  OR2_X1 U2620 ( .A1(n2243), .A2(n2232), .ZN(n2715) );
  OR2_X1 U2621 ( .A1(n2716), .A2(n2717), .ZN(n2232) );
  AND2_X1 U2622 ( .A1(n2207), .A2(n2218), .ZN(n2717) );
  AND2_X1 U2623 ( .A1(b_13_), .A2(n2718), .ZN(n2716) );
  OR2_X1 U2624 ( .A1(n2218), .A2(n2207), .ZN(n2718) );
  OR2_X1 U2625 ( .A1(n2719), .A2(n2720), .ZN(n2207) );
  AND2_X1 U2626 ( .A1(n2162), .A2(n2174), .ZN(n2720) );
  AND2_X1 U2627 ( .A1(b_14_), .A2(n2721), .ZN(n2719) );
  OR2_X1 U2628 ( .A1(n2162), .A2(n2174), .ZN(n2721) );
  INV_X1 U2629 ( .A(n2184), .ZN(n2162) );
  OR2_X1 U2630 ( .A1(a_15_), .A2(n2620), .ZN(n2184) );
  AND2_X1 U2631 ( .A1(n2563), .A2(operation_1_), .ZN(n2158) );
  INV_X1 U2632 ( .A(operation_0_), .ZN(n2563) );
  AND3_X1 U2633 ( .A1(n2722), .A2(n2623), .A3(n2159), .ZN(n2675) );
  AND2_X1 U2634 ( .A1(n2562), .A2(operation_0_), .ZN(n2159) );
  INV_X1 U2635 ( .A(operation_1_), .ZN(n2562) );
  OR2_X1 U2636 ( .A1(a_0_), .A2(n2723), .ZN(n2623) );
  OR2_X1 U2637 ( .A1(n2622), .A2(n2553), .ZN(n2722) );
  OR2_X1 U2638 ( .A1(n2724), .A2(n2725), .ZN(n2553) );
  AND2_X1 U2639 ( .A1(a_1_), .A2(n2528), .ZN(n2725) );
  AND2_X1 U2640 ( .A1(n2726), .A2(n2567), .ZN(n2724) );
  OR2_X1 U2641 ( .A1(a_1_), .A2(n2528), .ZN(n2726) );
  OR2_X1 U2642 ( .A1(n2727), .A2(n2728), .ZN(n2528) );
  AND2_X1 U2643 ( .A1(a_2_), .A2(n2502), .ZN(n2728) );
  AND2_X1 U2644 ( .A1(n2729), .A2(n2571), .ZN(n2727) );
  OR2_X1 U2645 ( .A1(a_2_), .A2(n2502), .ZN(n2729) );
  OR2_X1 U2646 ( .A1(n2730), .A2(n2731), .ZN(n2502) );
  AND2_X1 U2647 ( .A1(a_3_), .A2(n2476), .ZN(n2731) );
  AND2_X1 U2648 ( .A1(n2732), .A2(n2575), .ZN(n2730) );
  OR2_X1 U2649 ( .A1(a_3_), .A2(n2476), .ZN(n2732) );
  OR2_X1 U2650 ( .A1(n2733), .A2(n2734), .ZN(n2476) );
  AND2_X1 U2651 ( .A1(a_4_), .A2(n2439), .ZN(n2734) );
  AND2_X1 U2652 ( .A1(n2735), .A2(n2579), .ZN(n2733) );
  OR2_X1 U2653 ( .A1(a_4_), .A2(n2439), .ZN(n2735) );
  OR2_X1 U2654 ( .A1(n2736), .A2(n2737), .ZN(n2439) );
  AND2_X1 U2655 ( .A1(a_5_), .A2(n2413), .ZN(n2737) );
  AND2_X1 U2656 ( .A1(n2738), .A2(n2583), .ZN(n2736) );
  OR2_X1 U2657 ( .A1(a_5_), .A2(n2413), .ZN(n2738) );
  OR2_X1 U2658 ( .A1(n2739), .A2(n2740), .ZN(n2413) );
  AND2_X1 U2659 ( .A1(a_6_), .A2(n2387), .ZN(n2740) );
  AND2_X1 U2660 ( .A1(n2741), .A2(n2587), .ZN(n2739) );
  OR2_X1 U2661 ( .A1(a_6_), .A2(n2387), .ZN(n2741) );
  OR2_X1 U2662 ( .A1(n2742), .A2(n2743), .ZN(n2387) );
  AND2_X1 U2663 ( .A1(a_7_), .A2(n2361), .ZN(n2743) );
  AND2_X1 U2664 ( .A1(n2744), .A2(n2591), .ZN(n2742) );
  OR2_X1 U2665 ( .A1(a_7_), .A2(n2361), .ZN(n2744) );
  OR2_X1 U2666 ( .A1(n2745), .A2(n2746), .ZN(n2361) );
  AND2_X1 U2667 ( .A1(a_8_), .A2(n2335), .ZN(n2746) );
  AND2_X1 U2668 ( .A1(n2747), .A2(n2595), .ZN(n2745) );
  OR2_X1 U2669 ( .A1(a_8_), .A2(n2335), .ZN(n2747) );
  OR2_X1 U2670 ( .A1(n2748), .A2(n2749), .ZN(n2335) );
  AND2_X1 U2671 ( .A1(a_9_), .A2(n2308), .ZN(n2749) );
  AND2_X1 U2672 ( .A1(n2750), .A2(n2598), .ZN(n2748) );
  OR2_X1 U2673 ( .A1(a_9_), .A2(n2308), .ZN(n2750) );
  OR2_X1 U2674 ( .A1(n2751), .A2(n2752), .ZN(n2308) );
  AND2_X1 U2675 ( .A1(a_10_), .A2(n2283), .ZN(n2752) );
  AND2_X1 U2676 ( .A1(n2753), .A2(n2602), .ZN(n2751) );
  OR2_X1 U2677 ( .A1(a_10_), .A2(n2283), .ZN(n2753) );
  OR2_X1 U2678 ( .A1(n2754), .A2(n2755), .ZN(n2283) );
  AND2_X1 U2679 ( .A1(a_11_), .A2(n2258), .ZN(n2755) );
  AND2_X1 U2680 ( .A1(n2756), .A2(n2606), .ZN(n2754) );
  OR2_X1 U2681 ( .A1(a_11_), .A2(n2258), .ZN(n2756) );
  OR2_X1 U2682 ( .A1(n2757), .A2(n2758), .ZN(n2258) );
  AND2_X1 U2683 ( .A1(a_12_), .A2(n2233), .ZN(n2758) );
  AND2_X1 U2684 ( .A1(n2759), .A2(n2610), .ZN(n2757) );
  OR2_X1 U2685 ( .A1(a_12_), .A2(n2233), .ZN(n2759) );
  OR2_X1 U2686 ( .A1(n2760), .A2(n2761), .ZN(n2233) );
  AND2_X1 U2687 ( .A1(a_13_), .A2(n2208), .ZN(n2761) );
  AND2_X1 U2688 ( .A1(n2762), .A2(n2614), .ZN(n2760) );
  OR2_X1 U2689 ( .A1(a_13_), .A2(n2208), .ZN(n2762) );
  OR2_X1 U2690 ( .A1(n2763), .A2(n2764), .ZN(n2208) );
  AND2_X1 U2691 ( .A1(a_14_), .A2(n2161), .ZN(n2764) );
  AND2_X1 U2692 ( .A1(n2765), .A2(n2167), .ZN(n2763) );
  OR2_X1 U2693 ( .A1(n2161), .A2(a_14_), .ZN(n2765) );
  INV_X1 U2694 ( .A(n2185), .ZN(n2161) );
  OR2_X1 U2695 ( .A1(b_15_), .A2(n2619), .ZN(n2185) );
  AND2_X1 U2696 ( .A1(n2723), .A2(a_0_), .ZN(n2622) );
  AND2_X1 U2697 ( .A1(n2126), .A2(n2766), .ZN(n2674) );
  OR3_X1 U2698 ( .A1(n2459), .A2(n2767), .A3(n2768), .ZN(n2766) );
  AND2_X1 U2699 ( .A1(n2769), .A2(a_0_), .ZN(n2768) );
  INV_X1 U2700 ( .A(n2770), .ZN(n2769) );
  AND2_X1 U2701 ( .A1(n2451), .A2(n2456), .ZN(n2767) );
  AND2_X1 U2702 ( .A1(n2192), .A2(n2193), .ZN(n2451) );
  XOR2_X1 U2703 ( .A(n2458), .B(n2457), .Z(n2193) );
  OR2_X1 U2704 ( .A1(n2771), .A2(n2772), .ZN(n2192) );
  AND2_X1 U2705 ( .A1(n2151), .A2(n2152), .ZN(n2772) );
  INV_X1 U2706 ( .A(n2773), .ZN(n2152) );
  OR2_X1 U2707 ( .A1(n2774), .A2(n2771), .ZN(n2773) );
  AND2_X1 U2708 ( .A1(n2775), .A2(n2776), .ZN(n2774) );
  OR2_X1 U2709 ( .A1(n2777), .A2(n2778), .ZN(n2151) );
  AND2_X1 U2710 ( .A1(n2147), .A2(n2148), .ZN(n2777) );
  INV_X1 U2711 ( .A(n2779), .ZN(n2148) );
  OR2_X1 U2712 ( .A1(n2780), .A2(n2778), .ZN(n2779) );
  INV_X1 U2713 ( .A(n2781), .ZN(n2778) );
  OR2_X1 U2714 ( .A1(n2782), .A2(n2783), .ZN(n2781) );
  AND2_X1 U2715 ( .A1(n2782), .A2(n2783), .ZN(n2780) );
  OR2_X1 U2716 ( .A1(n2784), .A2(n2785), .ZN(n2783) );
  AND2_X1 U2717 ( .A1(n2786), .A2(n2787), .ZN(n2785) );
  AND2_X1 U2718 ( .A1(n2788), .A2(n2789), .ZN(n2784) );
  OR2_X1 U2719 ( .A1(n2787), .A2(n2786), .ZN(n2789) );
  XOR2_X1 U2720 ( .A(n2790), .B(n2791), .Z(n2782) );
  XOR2_X1 U2721 ( .A(n2792), .B(n2793), .Z(n2791) );
  OR2_X1 U2722 ( .A1(n2794), .A2(n2795), .ZN(n2147) );
  AND2_X1 U2723 ( .A1(n2143), .A2(n2144), .ZN(n2795) );
  INV_X1 U2724 ( .A(n2796), .ZN(n2144) );
  OR2_X1 U2725 ( .A1(n2797), .A2(n2794), .ZN(n2796) );
  AND2_X1 U2726 ( .A1(n2798), .A2(n2799), .ZN(n2797) );
  OR2_X1 U2727 ( .A1(n2800), .A2(n2801), .ZN(n2143) );
  AND2_X1 U2728 ( .A1(n2139), .A2(n2140), .ZN(n2800) );
  INV_X1 U2729 ( .A(n2802), .ZN(n2140) );
  OR2_X1 U2730 ( .A1(n2803), .A2(n2801), .ZN(n2802) );
  INV_X1 U2731 ( .A(n2804), .ZN(n2801) );
  OR2_X1 U2732 ( .A1(n2805), .A2(n2806), .ZN(n2804) );
  AND2_X1 U2733 ( .A1(n2805), .A2(n2806), .ZN(n2803) );
  OR2_X1 U2734 ( .A1(n2807), .A2(n2808), .ZN(n2806) );
  AND2_X1 U2735 ( .A1(n2809), .A2(n2810), .ZN(n2808) );
  AND2_X1 U2736 ( .A1(n2811), .A2(n2812), .ZN(n2807) );
  OR2_X1 U2737 ( .A1(n2810), .A2(n2809), .ZN(n2812) );
  XOR2_X1 U2738 ( .A(n2813), .B(n2814), .Z(n2805) );
  XOR2_X1 U2739 ( .A(n2815), .B(n2816), .Z(n2814) );
  OR2_X1 U2740 ( .A1(n2817), .A2(n2818), .ZN(n2139) );
  AND2_X1 U2741 ( .A1(n2135), .A2(n2136), .ZN(n2818) );
  INV_X1 U2742 ( .A(n2819), .ZN(n2136) );
  OR2_X1 U2743 ( .A1(n2820), .A2(n2817), .ZN(n2819) );
  AND2_X1 U2744 ( .A1(n2821), .A2(n2822), .ZN(n2820) );
  OR2_X1 U2745 ( .A1(n2823), .A2(n2824), .ZN(n2135) );
  AND2_X1 U2746 ( .A1(n2131), .A2(n2132), .ZN(n2823) );
  INV_X1 U2747 ( .A(n2825), .ZN(n2132) );
  OR2_X1 U2748 ( .A1(n2826), .A2(n2824), .ZN(n2825) );
  INV_X1 U2749 ( .A(n2827), .ZN(n2824) );
  OR2_X1 U2750 ( .A1(n2828), .A2(n2829), .ZN(n2827) );
  AND2_X1 U2751 ( .A1(n2828), .A2(n2829), .ZN(n2826) );
  OR2_X1 U2752 ( .A1(n2830), .A2(n2831), .ZN(n2829) );
  AND2_X1 U2753 ( .A1(n2832), .A2(n2833), .ZN(n2831) );
  AND2_X1 U2754 ( .A1(n2834), .A2(n2835), .ZN(n2830) );
  OR2_X1 U2755 ( .A1(n2833), .A2(n2832), .ZN(n2835) );
  XOR2_X1 U2756 ( .A(n2836), .B(n2837), .Z(n2828) );
  XOR2_X1 U2757 ( .A(n2838), .B(n2839), .Z(n2837) );
  OR2_X1 U2758 ( .A1(n2840), .A2(n2841), .ZN(n2131) );
  AND2_X1 U2759 ( .A1(n2127), .A2(n2128), .ZN(n2841) );
  INV_X1 U2760 ( .A(n2842), .ZN(n2128) );
  OR2_X1 U2761 ( .A1(n2843), .A2(n2840), .ZN(n2842) );
  AND2_X1 U2762 ( .A1(n2844), .A2(n2845), .ZN(n2843) );
  OR2_X1 U2763 ( .A1(n2846), .A2(n2847), .ZN(n2127) );
  INV_X1 U2764 ( .A(n2848), .ZN(n2847) );
  OR2_X1 U2765 ( .A1(n2849), .A2(n2673), .ZN(n2846) );
  AND3_X1 U2766 ( .A1(n2672), .A2(n2671), .A3(n2669), .ZN(n2673) );
  AND2_X1 U2767 ( .A1(n2669), .A2(n2665), .ZN(n2849) );
  OR2_X1 U2768 ( .A1(n2850), .A2(n2662), .ZN(n2665) );
  AND3_X1 U2769 ( .A1(n2661), .A2(n2659), .A3(n2660), .ZN(n2662) );
  AND2_X1 U2770 ( .A1(n2659), .A2(n2654), .ZN(n2850) );
  OR2_X1 U2771 ( .A1(n2851), .A2(n2651), .ZN(n2654) );
  AND2_X1 U2772 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  AND2_X1 U2773 ( .A1(n2650), .A2(n2645), .ZN(n2851) );
  OR2_X1 U2774 ( .A1(n2852), .A2(n2637), .ZN(n2645) );
  INV_X1 U2775 ( .A(n2853), .ZN(n2637) );
  OR3_X1 U2776 ( .A1(n2641), .A2(n2640), .A3(n2639), .ZN(n2853) );
  AND2_X1 U2777 ( .A1(n2642), .A2(n2854), .ZN(n2852) );
  INV_X1 U2778 ( .A(n2639), .ZN(n2854) );
  OR2_X1 U2779 ( .A1(n2855), .A2(n2649), .ZN(n2639) );
  INV_X1 U2780 ( .A(n2856), .ZN(n2649) );
  OR2_X1 U2781 ( .A1(n2857), .A2(n2858), .ZN(n2856) );
  AND2_X1 U2782 ( .A1(n2857), .A2(n2858), .ZN(n2855) );
  OR2_X1 U2783 ( .A1(n2859), .A2(n2860), .ZN(n2858) );
  AND2_X1 U2784 ( .A1(n2861), .A2(n2862), .ZN(n2860) );
  AND2_X1 U2785 ( .A1(n2863), .A2(n2864), .ZN(n2859) );
  OR2_X1 U2786 ( .A1(n2862), .A2(n2861), .ZN(n2864) );
  XOR2_X1 U2787 ( .A(n2865), .B(n2866), .Z(n2857) );
  XOR2_X1 U2788 ( .A(n2867), .B(n2868), .Z(n2866) );
  AND3_X1 U2789 ( .A1(n2627), .A2(n2632), .A3(n2626), .ZN(n2642) );
  INV_X1 U2790 ( .A(n2869), .ZN(n2626) );
  OR2_X1 U2791 ( .A1(n2870), .A2(n2871), .ZN(n2869) );
  AND2_X1 U2792 ( .A1(n2545), .A2(n2544), .ZN(n2871) );
  AND2_X1 U2793 ( .A1(n2542), .A2(n2872), .ZN(n2870) );
  OR2_X1 U2794 ( .A1(n2545), .A2(n2544), .ZN(n2872) );
  OR2_X1 U2795 ( .A1(n2873), .A2(n2874), .ZN(n2544) );
  AND2_X1 U2796 ( .A1(n2519), .A2(n2518), .ZN(n2874) );
  AND2_X1 U2797 ( .A1(n2516), .A2(n2875), .ZN(n2873) );
  OR2_X1 U2798 ( .A1(n2519), .A2(n2518), .ZN(n2875) );
  OR2_X1 U2799 ( .A1(n2876), .A2(n2877), .ZN(n2518) );
  AND2_X1 U2800 ( .A1(n2493), .A2(n2492), .ZN(n2877) );
  AND2_X1 U2801 ( .A1(n2490), .A2(n2878), .ZN(n2876) );
  OR2_X1 U2802 ( .A1(n2493), .A2(n2492), .ZN(n2878) );
  OR2_X1 U2803 ( .A1(n2879), .A2(n2880), .ZN(n2492) );
  AND2_X1 U2804 ( .A1(n2467), .A2(n2466), .ZN(n2880) );
  AND2_X1 U2805 ( .A1(n2464), .A2(n2881), .ZN(n2879) );
  OR2_X1 U2806 ( .A1(n2467), .A2(n2466), .ZN(n2881) );
  OR2_X1 U2807 ( .A1(n2882), .A2(n2883), .ZN(n2466) );
  AND2_X1 U2808 ( .A1(n2430), .A2(n2429), .ZN(n2883) );
  AND2_X1 U2809 ( .A1(n2427), .A2(n2884), .ZN(n2882) );
  OR2_X1 U2810 ( .A1(n2430), .A2(n2429), .ZN(n2884) );
  OR2_X1 U2811 ( .A1(n2885), .A2(n2886), .ZN(n2429) );
  AND2_X1 U2812 ( .A1(n2404), .A2(n2403), .ZN(n2886) );
  AND2_X1 U2813 ( .A1(n2401), .A2(n2887), .ZN(n2885) );
  OR2_X1 U2814 ( .A1(n2404), .A2(n2403), .ZN(n2887) );
  OR2_X1 U2815 ( .A1(n2888), .A2(n2889), .ZN(n2403) );
  AND2_X1 U2816 ( .A1(n2378), .A2(n2377), .ZN(n2889) );
  AND2_X1 U2817 ( .A1(n2375), .A2(n2890), .ZN(n2888) );
  OR2_X1 U2818 ( .A1(n2378), .A2(n2377), .ZN(n2890) );
  OR2_X1 U2819 ( .A1(n2891), .A2(n2892), .ZN(n2377) );
  AND2_X1 U2820 ( .A1(n2352), .A2(n2351), .ZN(n2892) );
  AND2_X1 U2821 ( .A1(n2349), .A2(n2893), .ZN(n2891) );
  OR2_X1 U2822 ( .A1(n2352), .A2(n2351), .ZN(n2893) );
  OR2_X1 U2823 ( .A1(n2894), .A2(n2895), .ZN(n2351) );
  AND2_X1 U2824 ( .A1(n2326), .A2(n2325), .ZN(n2895) );
  AND2_X1 U2825 ( .A1(n2323), .A2(n2896), .ZN(n2894) );
  OR2_X1 U2826 ( .A1(n2326), .A2(n2325), .ZN(n2896) );
  OR2_X1 U2827 ( .A1(n2897), .A2(n2898), .ZN(n2325) );
  AND2_X1 U2828 ( .A1(n2301), .A2(n2300), .ZN(n2898) );
  AND2_X1 U2829 ( .A1(n2298), .A2(n2899), .ZN(n2897) );
  OR2_X1 U2830 ( .A1(n2301), .A2(n2300), .ZN(n2899) );
  OR2_X1 U2831 ( .A1(n2900), .A2(n2901), .ZN(n2300) );
  AND2_X1 U2832 ( .A1(n2276), .A2(n2275), .ZN(n2901) );
  AND2_X1 U2833 ( .A1(n2273), .A2(n2902), .ZN(n2900) );
  OR2_X1 U2834 ( .A1(n2276), .A2(n2275), .ZN(n2902) );
  OR2_X1 U2835 ( .A1(n2903), .A2(n2904), .ZN(n2275) );
  AND2_X1 U2836 ( .A1(n2251), .A2(n2250), .ZN(n2904) );
  AND2_X1 U2837 ( .A1(n2248), .A2(n2905), .ZN(n2903) );
  OR2_X1 U2838 ( .A1(n2251), .A2(n2250), .ZN(n2905) );
  OR2_X1 U2839 ( .A1(n2906), .A2(n2907), .ZN(n2250) );
  AND2_X1 U2840 ( .A1(n2226), .A2(n2225), .ZN(n2907) );
  AND2_X1 U2841 ( .A1(n2223), .A2(n2908), .ZN(n2906) );
  OR2_X1 U2842 ( .A1(n2226), .A2(n2225), .ZN(n2908) );
  OR2_X1 U2843 ( .A1(n2909), .A2(n2910), .ZN(n2225) );
  AND2_X1 U2844 ( .A1(n2198), .A2(n2201), .ZN(n2910) );
  AND2_X1 U2845 ( .A1(n2911), .A2(n2912), .ZN(n2909) );
  OR2_X1 U2846 ( .A1(n2198), .A2(n2201), .ZN(n2912) );
  OR2_X1 U2847 ( .A1(n2218), .A2(n2620), .ZN(n2201) );
  OR2_X1 U2848 ( .A1(n2167), .A2(n2616), .ZN(n2198) );
  OR2_X1 U2849 ( .A1(n2620), .A2(n2913), .ZN(n2616) );
  INV_X1 U2850 ( .A(n2200), .ZN(n2911) );
  OR2_X1 U2851 ( .A1(n2914), .A2(n2915), .ZN(n2200) );
  AND2_X1 U2852 ( .A1(b_14_), .A2(n2916), .ZN(n2915) );
  OR2_X1 U2853 ( .A1(n2917), .A2(n2918), .ZN(n2916) );
  AND2_X1 U2854 ( .A1(a_14_), .A2(n2614), .ZN(n2917) );
  AND2_X1 U2855 ( .A1(b_13_), .A2(n2919), .ZN(n2914) );
  OR2_X1 U2856 ( .A1(n2920), .A2(n2180), .ZN(n2919) );
  AND2_X1 U2857 ( .A1(a_15_), .A2(n2167), .ZN(n2920) );
  OR2_X1 U2858 ( .A1(n2243), .A2(n2620), .ZN(n2226) );
  XNOR2_X1 U2859 ( .A(n2921), .B(n2922), .ZN(n2223) );
  XOR2_X1 U2860 ( .A(n2923), .B(n2924), .Z(n2922) );
  OR2_X1 U2861 ( .A1(n2268), .A2(n2620), .ZN(n2251) );
  XOR2_X1 U2862 ( .A(n2925), .B(n2926), .Z(n2248) );
  XOR2_X1 U2863 ( .A(n2927), .B(n2928), .Z(n2926) );
  OR2_X1 U2864 ( .A1(n2293), .A2(n2620), .ZN(n2276) );
  XOR2_X1 U2865 ( .A(n2929), .B(n2930), .Z(n2273) );
  XOR2_X1 U2866 ( .A(n2931), .B(n2932), .Z(n2930) );
  OR2_X1 U2867 ( .A1(n2318), .A2(n2620), .ZN(n2301) );
  XOR2_X1 U2868 ( .A(n2933), .B(n2934), .Z(n2298) );
  XOR2_X1 U2869 ( .A(n2935), .B(n2936), .Z(n2934) );
  OR2_X1 U2870 ( .A1(n2594), .A2(n2620), .ZN(n2326) );
  XOR2_X1 U2871 ( .A(n2937), .B(n2938), .Z(n2323) );
  XOR2_X1 U2872 ( .A(n2939), .B(n2940), .Z(n2938) );
  OR2_X1 U2873 ( .A1(n2590), .A2(n2620), .ZN(n2352) );
  XOR2_X1 U2874 ( .A(n2941), .B(n2942), .Z(n2349) );
  XOR2_X1 U2875 ( .A(n2943), .B(n2944), .Z(n2942) );
  OR2_X1 U2876 ( .A1(n2586), .A2(n2620), .ZN(n2378) );
  XOR2_X1 U2877 ( .A(n2945), .B(n2946), .Z(n2375) );
  XOR2_X1 U2878 ( .A(n2947), .B(n2948), .Z(n2946) );
  OR2_X1 U2879 ( .A1(n2582), .A2(n2620), .ZN(n2404) );
  XOR2_X1 U2880 ( .A(n2949), .B(n2950), .Z(n2401) );
  XOR2_X1 U2881 ( .A(n2951), .B(n2952), .Z(n2950) );
  OR2_X1 U2882 ( .A1(n2578), .A2(n2620), .ZN(n2430) );
  XOR2_X1 U2883 ( .A(n2953), .B(n2954), .Z(n2427) );
  XOR2_X1 U2884 ( .A(n2955), .B(n2956), .Z(n2954) );
  OR2_X1 U2885 ( .A1(n2574), .A2(n2620), .ZN(n2467) );
  XOR2_X1 U2886 ( .A(n2957), .B(n2958), .Z(n2464) );
  XOR2_X1 U2887 ( .A(n2959), .B(n2960), .Z(n2958) );
  OR2_X1 U2888 ( .A1(n2570), .A2(n2620), .ZN(n2493) );
  XOR2_X1 U2889 ( .A(n2961), .B(n2962), .Z(n2490) );
  XOR2_X1 U2890 ( .A(n2963), .B(n2964), .Z(n2962) );
  OR2_X1 U2891 ( .A1(n2566), .A2(n2620), .ZN(n2519) );
  XOR2_X1 U2892 ( .A(n2965), .B(n2966), .Z(n2516) );
  XOR2_X1 U2893 ( .A(n2967), .B(n2968), .Z(n2966) );
  OR2_X1 U2894 ( .A1(n2969), .A2(n2620), .ZN(n2545) );
  INV_X1 U2895 ( .A(b_15_), .ZN(n2620) );
  XOR2_X1 U2896 ( .A(n2970), .B(n2971), .Z(n2542) );
  XOR2_X1 U2897 ( .A(n2972), .B(n2973), .Z(n2971) );
  XOR2_X1 U2898 ( .A(n2640), .B(n2641), .Z(n2632) );
  OR2_X1 U2899 ( .A1(n2974), .A2(n2975), .ZN(n2641) );
  AND2_X1 U2900 ( .A1(n2976), .A2(n2977), .ZN(n2975) );
  AND2_X1 U2901 ( .A1(n2978), .A2(n2979), .ZN(n2974) );
  OR2_X1 U2902 ( .A1(n2976), .A2(n2977), .ZN(n2979) );
  XOR2_X1 U2903 ( .A(n2863), .B(n2980), .Z(n2640) );
  XOR2_X1 U2904 ( .A(n2862), .B(n2861), .Z(n2980) );
  OR2_X1 U2905 ( .A1(n2969), .A2(n2614), .ZN(n2861) );
  OR2_X1 U2906 ( .A1(n2981), .A2(n2982), .ZN(n2862) );
  AND2_X1 U2907 ( .A1(n2983), .A2(n2984), .ZN(n2982) );
  AND2_X1 U2908 ( .A1(n2985), .A2(n2986), .ZN(n2981) );
  OR2_X1 U2909 ( .A1(n2984), .A2(n2983), .ZN(n2986) );
  XOR2_X1 U2910 ( .A(n2987), .B(n2988), .Z(n2863) );
  XOR2_X1 U2911 ( .A(n2989), .B(n2990), .Z(n2988) );
  XNOR2_X1 U2912 ( .A(n2978), .B(n2991), .ZN(n2627) );
  XOR2_X1 U2913 ( .A(n2977), .B(n2976), .Z(n2991) );
  OR2_X1 U2914 ( .A1(n2969), .A2(n2167), .ZN(n2976) );
  OR2_X1 U2915 ( .A1(n2992), .A2(n2993), .ZN(n2977) );
  AND2_X1 U2916 ( .A1(n2973), .A2(n2972), .ZN(n2993) );
  AND2_X1 U2917 ( .A1(n2970), .A2(n2994), .ZN(n2992) );
  OR2_X1 U2918 ( .A1(n2972), .A2(n2973), .ZN(n2994) );
  OR2_X1 U2919 ( .A1(n2566), .A2(n2167), .ZN(n2973) );
  OR2_X1 U2920 ( .A1(n2995), .A2(n2996), .ZN(n2972) );
  AND2_X1 U2921 ( .A1(n2968), .A2(n2967), .ZN(n2996) );
  AND2_X1 U2922 ( .A1(n2965), .A2(n2997), .ZN(n2995) );
  OR2_X1 U2923 ( .A1(n2967), .A2(n2968), .ZN(n2997) );
  OR2_X1 U2924 ( .A1(n2570), .A2(n2167), .ZN(n2968) );
  OR2_X1 U2925 ( .A1(n2998), .A2(n2999), .ZN(n2967) );
  AND2_X1 U2926 ( .A1(n2964), .A2(n2963), .ZN(n2999) );
  AND2_X1 U2927 ( .A1(n2961), .A2(n3000), .ZN(n2998) );
  OR2_X1 U2928 ( .A1(n2963), .A2(n2964), .ZN(n3000) );
  OR2_X1 U2929 ( .A1(n2574), .A2(n2167), .ZN(n2964) );
  OR2_X1 U2930 ( .A1(n3001), .A2(n3002), .ZN(n2963) );
  AND2_X1 U2931 ( .A1(n2960), .A2(n2959), .ZN(n3002) );
  AND2_X1 U2932 ( .A1(n2957), .A2(n3003), .ZN(n3001) );
  OR2_X1 U2933 ( .A1(n2959), .A2(n2960), .ZN(n3003) );
  OR2_X1 U2934 ( .A1(n2578), .A2(n2167), .ZN(n2960) );
  OR2_X1 U2935 ( .A1(n3004), .A2(n3005), .ZN(n2959) );
  AND2_X1 U2936 ( .A1(n2956), .A2(n2955), .ZN(n3005) );
  AND2_X1 U2937 ( .A1(n2953), .A2(n3006), .ZN(n3004) );
  OR2_X1 U2938 ( .A1(n2955), .A2(n2956), .ZN(n3006) );
  OR2_X1 U2939 ( .A1(n2582), .A2(n2167), .ZN(n2956) );
  OR2_X1 U2940 ( .A1(n3007), .A2(n3008), .ZN(n2955) );
  AND2_X1 U2941 ( .A1(n2952), .A2(n2951), .ZN(n3008) );
  AND2_X1 U2942 ( .A1(n2949), .A2(n3009), .ZN(n3007) );
  OR2_X1 U2943 ( .A1(n2951), .A2(n2952), .ZN(n3009) );
  OR2_X1 U2944 ( .A1(n2586), .A2(n2167), .ZN(n2952) );
  OR2_X1 U2945 ( .A1(n3010), .A2(n3011), .ZN(n2951) );
  AND2_X1 U2946 ( .A1(n2948), .A2(n2947), .ZN(n3011) );
  AND2_X1 U2947 ( .A1(n2945), .A2(n3012), .ZN(n3010) );
  OR2_X1 U2948 ( .A1(n2947), .A2(n2948), .ZN(n3012) );
  OR2_X1 U2949 ( .A1(n2590), .A2(n2167), .ZN(n2948) );
  OR2_X1 U2950 ( .A1(n3013), .A2(n3014), .ZN(n2947) );
  AND2_X1 U2951 ( .A1(n2944), .A2(n2943), .ZN(n3014) );
  AND2_X1 U2952 ( .A1(n2941), .A2(n3015), .ZN(n3013) );
  OR2_X1 U2953 ( .A1(n2943), .A2(n2944), .ZN(n3015) );
  OR2_X1 U2954 ( .A1(n2594), .A2(n2167), .ZN(n2944) );
  OR2_X1 U2955 ( .A1(n3016), .A2(n3017), .ZN(n2943) );
  AND2_X1 U2956 ( .A1(n2940), .A2(n2939), .ZN(n3017) );
  AND2_X1 U2957 ( .A1(n2937), .A2(n3018), .ZN(n3016) );
  OR2_X1 U2958 ( .A1(n2939), .A2(n2940), .ZN(n3018) );
  OR2_X1 U2959 ( .A1(n2318), .A2(n2167), .ZN(n2940) );
  OR2_X1 U2960 ( .A1(n3019), .A2(n3020), .ZN(n2939) );
  AND2_X1 U2961 ( .A1(n2936), .A2(n2935), .ZN(n3020) );
  AND2_X1 U2962 ( .A1(n2933), .A2(n3021), .ZN(n3019) );
  OR2_X1 U2963 ( .A1(n2935), .A2(n2936), .ZN(n3021) );
  OR2_X1 U2964 ( .A1(n2293), .A2(n2167), .ZN(n2936) );
  OR2_X1 U2965 ( .A1(n3022), .A2(n3023), .ZN(n2935) );
  AND2_X1 U2966 ( .A1(n2932), .A2(n2931), .ZN(n3023) );
  AND2_X1 U2967 ( .A1(n2929), .A2(n3024), .ZN(n3022) );
  OR2_X1 U2968 ( .A1(n2931), .A2(n2932), .ZN(n3024) );
  OR2_X1 U2969 ( .A1(n2268), .A2(n2167), .ZN(n2932) );
  OR2_X1 U2970 ( .A1(n3025), .A2(n3026), .ZN(n2931) );
  AND2_X1 U2971 ( .A1(n2928), .A2(n2927), .ZN(n3026) );
  AND2_X1 U2972 ( .A1(n2925), .A2(n3027), .ZN(n3025) );
  OR2_X1 U2973 ( .A1(n2927), .A2(n2928), .ZN(n3027) );
  OR2_X1 U2974 ( .A1(n2243), .A2(n2167), .ZN(n2928) );
  OR2_X1 U2975 ( .A1(n3028), .A2(n3029), .ZN(n2927) );
  AND2_X1 U2976 ( .A1(n2921), .A2(n2924), .ZN(n3029) );
  AND2_X1 U2977 ( .A1(n3030), .A2(n3031), .ZN(n3028) );
  OR2_X1 U2978 ( .A1(n2924), .A2(n2921), .ZN(n3031) );
  OR2_X1 U2979 ( .A1(n2218), .A2(n2167), .ZN(n2921) );
  OR3_X1 U2980 ( .A1(n2167), .A2(n2614), .A3(n2913), .ZN(n2924) );
  INV_X1 U2981 ( .A(b_14_), .ZN(n2167) );
  INV_X1 U2982 ( .A(n2923), .ZN(n3030) );
  OR2_X1 U2983 ( .A1(n3032), .A2(n3033), .ZN(n2923) );
  AND2_X1 U2984 ( .A1(b_13_), .A2(n3034), .ZN(n3033) );
  OR2_X1 U2985 ( .A1(n3035), .A2(n2918), .ZN(n3034) );
  AND2_X1 U2986 ( .A1(a_14_), .A2(n2610), .ZN(n3035) );
  AND2_X1 U2987 ( .A1(b_12_), .A2(n3036), .ZN(n3032) );
  OR2_X1 U2988 ( .A1(n3037), .A2(n2180), .ZN(n3036) );
  AND2_X1 U2989 ( .A1(a_15_), .A2(n2614), .ZN(n3037) );
  XNOR2_X1 U2990 ( .A(n2615), .B(n3038), .ZN(n2925) );
  XOR2_X1 U2991 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR2_X1 U2992 ( .A(n3041), .B(n3042), .Z(n2929) );
  XOR2_X1 U2993 ( .A(n3043), .B(n3044), .Z(n3042) );
  XOR2_X1 U2994 ( .A(n3045), .B(n3046), .Z(n2933) );
  XOR2_X1 U2995 ( .A(n3047), .B(n3048), .Z(n3046) );
  XOR2_X1 U2996 ( .A(n3049), .B(n3050), .Z(n2937) );
  XOR2_X1 U2997 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR2_X1 U2998 ( .A(n3053), .B(n3054), .Z(n2941) );
  XOR2_X1 U2999 ( .A(n3055), .B(n3056), .Z(n3054) );
  XOR2_X1 U3000 ( .A(n3057), .B(n3058), .Z(n2945) );
  XOR2_X1 U3001 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR2_X1 U3002 ( .A(n3061), .B(n3062), .Z(n2949) );
  XOR2_X1 U3003 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR2_X1 U3004 ( .A(n3065), .B(n3066), .Z(n2953) );
  XOR2_X1 U3005 ( .A(n3067), .B(n3068), .Z(n3066) );
  XOR2_X1 U3006 ( .A(n3069), .B(n3070), .Z(n2957) );
  XOR2_X1 U3007 ( .A(n3071), .B(n3072), .Z(n3070) );
  XOR2_X1 U3008 ( .A(n3073), .B(n3074), .Z(n2961) );
  XOR2_X1 U3009 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR2_X1 U3010 ( .A(n3077), .B(n3078), .Z(n2965) );
  XOR2_X1 U3011 ( .A(n3079), .B(n3080), .Z(n3078) );
  XOR2_X1 U3012 ( .A(n3081), .B(n3082), .Z(n2970) );
  XOR2_X1 U3013 ( .A(n3083), .B(n3084), .Z(n3082) );
  XOR2_X1 U3014 ( .A(n2985), .B(n3085), .Z(n2978) );
  XOR2_X1 U3015 ( .A(n2984), .B(n2983), .Z(n3085) );
  OR2_X1 U3016 ( .A1(n2566), .A2(n2614), .ZN(n2983) );
  OR2_X1 U3017 ( .A1(n3086), .A2(n3087), .ZN(n2984) );
  AND2_X1 U3018 ( .A1(n3084), .A2(n3083), .ZN(n3087) );
  AND2_X1 U3019 ( .A1(n3081), .A2(n3088), .ZN(n3086) );
  OR2_X1 U3020 ( .A1(n3083), .A2(n3084), .ZN(n3088) );
  OR2_X1 U3021 ( .A1(n2570), .A2(n2614), .ZN(n3084) );
  OR2_X1 U3022 ( .A1(n3089), .A2(n3090), .ZN(n3083) );
  AND2_X1 U3023 ( .A1(n3080), .A2(n3079), .ZN(n3090) );
  AND2_X1 U3024 ( .A1(n3077), .A2(n3091), .ZN(n3089) );
  OR2_X1 U3025 ( .A1(n3079), .A2(n3080), .ZN(n3091) );
  OR2_X1 U3026 ( .A1(n2574), .A2(n2614), .ZN(n3080) );
  OR2_X1 U3027 ( .A1(n3092), .A2(n3093), .ZN(n3079) );
  AND2_X1 U3028 ( .A1(n3076), .A2(n3075), .ZN(n3093) );
  AND2_X1 U3029 ( .A1(n3073), .A2(n3094), .ZN(n3092) );
  OR2_X1 U3030 ( .A1(n3075), .A2(n3076), .ZN(n3094) );
  OR2_X1 U3031 ( .A1(n2578), .A2(n2614), .ZN(n3076) );
  OR2_X1 U3032 ( .A1(n3095), .A2(n3096), .ZN(n3075) );
  AND2_X1 U3033 ( .A1(n3072), .A2(n3071), .ZN(n3096) );
  AND2_X1 U3034 ( .A1(n3069), .A2(n3097), .ZN(n3095) );
  OR2_X1 U3035 ( .A1(n3071), .A2(n3072), .ZN(n3097) );
  OR2_X1 U3036 ( .A1(n2582), .A2(n2614), .ZN(n3072) );
  OR2_X1 U3037 ( .A1(n3098), .A2(n3099), .ZN(n3071) );
  AND2_X1 U3038 ( .A1(n3068), .A2(n3067), .ZN(n3099) );
  AND2_X1 U3039 ( .A1(n3065), .A2(n3100), .ZN(n3098) );
  OR2_X1 U3040 ( .A1(n3067), .A2(n3068), .ZN(n3100) );
  OR2_X1 U3041 ( .A1(n2586), .A2(n2614), .ZN(n3068) );
  OR2_X1 U3042 ( .A1(n3101), .A2(n3102), .ZN(n3067) );
  AND2_X1 U3043 ( .A1(n3064), .A2(n3063), .ZN(n3102) );
  AND2_X1 U3044 ( .A1(n3061), .A2(n3103), .ZN(n3101) );
  OR2_X1 U3045 ( .A1(n3063), .A2(n3064), .ZN(n3103) );
  OR2_X1 U3046 ( .A1(n2590), .A2(n2614), .ZN(n3064) );
  OR2_X1 U3047 ( .A1(n3104), .A2(n3105), .ZN(n3063) );
  AND2_X1 U3048 ( .A1(n3060), .A2(n3059), .ZN(n3105) );
  AND2_X1 U3049 ( .A1(n3057), .A2(n3106), .ZN(n3104) );
  OR2_X1 U3050 ( .A1(n3059), .A2(n3060), .ZN(n3106) );
  OR2_X1 U3051 ( .A1(n2594), .A2(n2614), .ZN(n3060) );
  OR2_X1 U3052 ( .A1(n3107), .A2(n3108), .ZN(n3059) );
  AND2_X1 U3053 ( .A1(n3056), .A2(n3055), .ZN(n3108) );
  AND2_X1 U3054 ( .A1(n3053), .A2(n3109), .ZN(n3107) );
  OR2_X1 U3055 ( .A1(n3055), .A2(n3056), .ZN(n3109) );
  OR2_X1 U3056 ( .A1(n2318), .A2(n2614), .ZN(n3056) );
  OR2_X1 U3057 ( .A1(n3110), .A2(n3111), .ZN(n3055) );
  AND2_X1 U3058 ( .A1(n3052), .A2(n3051), .ZN(n3111) );
  AND2_X1 U3059 ( .A1(n3049), .A2(n3112), .ZN(n3110) );
  OR2_X1 U3060 ( .A1(n3051), .A2(n3052), .ZN(n3112) );
  OR2_X1 U3061 ( .A1(n2293), .A2(n2614), .ZN(n3052) );
  OR2_X1 U3062 ( .A1(n3113), .A2(n3114), .ZN(n3051) );
  AND2_X1 U3063 ( .A1(n3048), .A2(n3047), .ZN(n3114) );
  AND2_X1 U3064 ( .A1(n3045), .A2(n3115), .ZN(n3113) );
  OR2_X1 U3065 ( .A1(n3047), .A2(n3048), .ZN(n3115) );
  OR2_X1 U3066 ( .A1(n2268), .A2(n2614), .ZN(n3048) );
  OR2_X1 U3067 ( .A1(n3116), .A2(n3117), .ZN(n3047) );
  AND2_X1 U3068 ( .A1(n3044), .A2(n3043), .ZN(n3117) );
  AND2_X1 U3069 ( .A1(n3041), .A2(n3118), .ZN(n3116) );
  OR2_X1 U3070 ( .A1(n3043), .A2(n3044), .ZN(n3118) );
  OR2_X1 U3071 ( .A1(n2243), .A2(n2614), .ZN(n3044) );
  OR2_X1 U3072 ( .A1(n3119), .A2(n3120), .ZN(n3043) );
  AND2_X1 U3073 ( .A1(n2615), .A2(n3040), .ZN(n3120) );
  AND2_X1 U3074 ( .A1(n3121), .A2(n3122), .ZN(n3119) );
  OR2_X1 U3075 ( .A1(n3040), .A2(n2615), .ZN(n3122) );
  OR2_X1 U3076 ( .A1(n2218), .A2(n2614), .ZN(n2615) );
  OR3_X1 U3077 ( .A1(n2614), .A2(n2610), .A3(n2913), .ZN(n3040) );
  INV_X1 U3078 ( .A(b_13_), .ZN(n2614) );
  INV_X1 U3079 ( .A(n3039), .ZN(n3121) );
  OR2_X1 U3080 ( .A1(n3123), .A2(n3124), .ZN(n3039) );
  AND2_X1 U3081 ( .A1(b_12_), .A2(n3125), .ZN(n3124) );
  OR2_X1 U3082 ( .A1(n3126), .A2(n2918), .ZN(n3125) );
  AND2_X1 U3083 ( .A1(a_14_), .A2(n2606), .ZN(n3126) );
  AND2_X1 U3084 ( .A1(b_11_), .A2(n3127), .ZN(n3123) );
  OR2_X1 U3085 ( .A1(n3128), .A2(n2180), .ZN(n3127) );
  AND2_X1 U3086 ( .A1(a_15_), .A2(n2610), .ZN(n3128) );
  XNOR2_X1 U3087 ( .A(n3129), .B(n3130), .ZN(n3041) );
  XOR2_X1 U3088 ( .A(n3131), .B(n3132), .Z(n3130) );
  XOR2_X1 U3089 ( .A(n3133), .B(n3134), .Z(n3045) );
  XOR2_X1 U3090 ( .A(n3135), .B(n2611), .Z(n3134) );
  XOR2_X1 U3091 ( .A(n3136), .B(n3137), .Z(n3049) );
  XOR2_X1 U3092 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR2_X1 U3093 ( .A(n3140), .B(n3141), .Z(n3053) );
  XOR2_X1 U3094 ( .A(n3142), .B(n3143), .Z(n3141) );
  XOR2_X1 U3095 ( .A(n3144), .B(n3145), .Z(n3057) );
  XOR2_X1 U3096 ( .A(n3146), .B(n3147), .Z(n3145) );
  XOR2_X1 U3097 ( .A(n3148), .B(n3149), .Z(n3061) );
  XOR2_X1 U3098 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR2_X1 U3099 ( .A(n3152), .B(n3153), .Z(n3065) );
  XOR2_X1 U3100 ( .A(n3154), .B(n3155), .Z(n3153) );
  XOR2_X1 U3101 ( .A(n3156), .B(n3157), .Z(n3069) );
  XOR2_X1 U3102 ( .A(n3158), .B(n3159), .Z(n3157) );
  XOR2_X1 U3103 ( .A(n3160), .B(n3161), .Z(n3073) );
  XOR2_X1 U3104 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR2_X1 U3105 ( .A(n3164), .B(n3165), .Z(n3077) );
  XOR2_X1 U3106 ( .A(n3166), .B(n3167), .Z(n3165) );
  XOR2_X1 U3107 ( .A(n3168), .B(n3169), .Z(n3081) );
  XOR2_X1 U3108 ( .A(n3170), .B(n3171), .Z(n3169) );
  XOR2_X1 U3109 ( .A(n3172), .B(n3173), .Z(n2985) );
  XOR2_X1 U3110 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR2_X1 U3111 ( .A(n2661), .B(n2660), .Z(n2650) );
  INV_X1 U3112 ( .A(n3176), .ZN(n2660) );
  OR2_X1 U3113 ( .A1(n3177), .A2(n3178), .ZN(n3176) );
  AND2_X1 U3114 ( .A1(n2868), .A2(n2867), .ZN(n3178) );
  AND2_X1 U3115 ( .A1(n2865), .A2(n3179), .ZN(n3177) );
  OR2_X1 U3116 ( .A1(n2867), .A2(n2868), .ZN(n3179) );
  OR2_X1 U3117 ( .A1(n2969), .A2(n2610), .ZN(n2868) );
  OR2_X1 U3118 ( .A1(n3180), .A2(n3181), .ZN(n2867) );
  AND2_X1 U3119 ( .A1(n2990), .A2(n2989), .ZN(n3181) );
  AND2_X1 U3120 ( .A1(n2987), .A2(n3182), .ZN(n3180) );
  OR2_X1 U3121 ( .A1(n2989), .A2(n2990), .ZN(n3182) );
  OR2_X1 U3122 ( .A1(n2566), .A2(n2610), .ZN(n2990) );
  OR2_X1 U3123 ( .A1(n3183), .A2(n3184), .ZN(n2989) );
  AND2_X1 U3124 ( .A1(n3175), .A2(n3174), .ZN(n3184) );
  AND2_X1 U3125 ( .A1(n3172), .A2(n3185), .ZN(n3183) );
  OR2_X1 U3126 ( .A1(n3174), .A2(n3175), .ZN(n3185) );
  OR2_X1 U3127 ( .A1(n2570), .A2(n2610), .ZN(n3175) );
  OR2_X1 U3128 ( .A1(n3186), .A2(n3187), .ZN(n3174) );
  AND2_X1 U3129 ( .A1(n3171), .A2(n3170), .ZN(n3187) );
  AND2_X1 U3130 ( .A1(n3168), .A2(n3188), .ZN(n3186) );
  OR2_X1 U3131 ( .A1(n3170), .A2(n3171), .ZN(n3188) );
  OR2_X1 U3132 ( .A1(n2574), .A2(n2610), .ZN(n3171) );
  OR2_X1 U3133 ( .A1(n3189), .A2(n3190), .ZN(n3170) );
  AND2_X1 U3134 ( .A1(n3167), .A2(n3166), .ZN(n3190) );
  AND2_X1 U3135 ( .A1(n3164), .A2(n3191), .ZN(n3189) );
  OR2_X1 U3136 ( .A1(n3166), .A2(n3167), .ZN(n3191) );
  OR2_X1 U3137 ( .A1(n2578), .A2(n2610), .ZN(n3167) );
  OR2_X1 U3138 ( .A1(n3192), .A2(n3193), .ZN(n3166) );
  AND2_X1 U3139 ( .A1(n3163), .A2(n3162), .ZN(n3193) );
  AND2_X1 U3140 ( .A1(n3160), .A2(n3194), .ZN(n3192) );
  OR2_X1 U3141 ( .A1(n3162), .A2(n3163), .ZN(n3194) );
  OR2_X1 U3142 ( .A1(n2582), .A2(n2610), .ZN(n3163) );
  OR2_X1 U3143 ( .A1(n3195), .A2(n3196), .ZN(n3162) );
  AND2_X1 U3144 ( .A1(n3159), .A2(n3158), .ZN(n3196) );
  AND2_X1 U3145 ( .A1(n3156), .A2(n3197), .ZN(n3195) );
  OR2_X1 U3146 ( .A1(n3158), .A2(n3159), .ZN(n3197) );
  OR2_X1 U3147 ( .A1(n2586), .A2(n2610), .ZN(n3159) );
  OR2_X1 U3148 ( .A1(n3198), .A2(n3199), .ZN(n3158) );
  AND2_X1 U3149 ( .A1(n3155), .A2(n3154), .ZN(n3199) );
  AND2_X1 U3150 ( .A1(n3152), .A2(n3200), .ZN(n3198) );
  OR2_X1 U3151 ( .A1(n3154), .A2(n3155), .ZN(n3200) );
  OR2_X1 U3152 ( .A1(n2590), .A2(n2610), .ZN(n3155) );
  OR2_X1 U3153 ( .A1(n3201), .A2(n3202), .ZN(n3154) );
  AND2_X1 U3154 ( .A1(n3151), .A2(n3150), .ZN(n3202) );
  AND2_X1 U3155 ( .A1(n3148), .A2(n3203), .ZN(n3201) );
  OR2_X1 U3156 ( .A1(n3150), .A2(n3151), .ZN(n3203) );
  OR2_X1 U3157 ( .A1(n2594), .A2(n2610), .ZN(n3151) );
  OR2_X1 U3158 ( .A1(n3204), .A2(n3205), .ZN(n3150) );
  AND2_X1 U3159 ( .A1(n3147), .A2(n3146), .ZN(n3205) );
  AND2_X1 U3160 ( .A1(n3144), .A2(n3206), .ZN(n3204) );
  OR2_X1 U3161 ( .A1(n3146), .A2(n3147), .ZN(n3206) );
  OR2_X1 U3162 ( .A1(n2318), .A2(n2610), .ZN(n3147) );
  OR2_X1 U3163 ( .A1(n3207), .A2(n3208), .ZN(n3146) );
  AND2_X1 U3164 ( .A1(n3143), .A2(n3142), .ZN(n3208) );
  AND2_X1 U3165 ( .A1(n3140), .A2(n3209), .ZN(n3207) );
  OR2_X1 U3166 ( .A1(n3142), .A2(n3143), .ZN(n3209) );
  OR2_X1 U3167 ( .A1(n2293), .A2(n2610), .ZN(n3143) );
  OR2_X1 U3168 ( .A1(n3210), .A2(n3211), .ZN(n3142) );
  AND2_X1 U3169 ( .A1(n3139), .A2(n3138), .ZN(n3211) );
  AND2_X1 U3170 ( .A1(n3136), .A2(n3212), .ZN(n3210) );
  OR2_X1 U3171 ( .A1(n3138), .A2(n3139), .ZN(n3212) );
  OR2_X1 U3172 ( .A1(n2268), .A2(n2610), .ZN(n3139) );
  OR2_X1 U3173 ( .A1(n3213), .A2(n3214), .ZN(n3138) );
  AND2_X1 U3174 ( .A1(n2611), .A2(n3135), .ZN(n3214) );
  AND2_X1 U3175 ( .A1(n3133), .A2(n3215), .ZN(n3213) );
  OR2_X1 U3176 ( .A1(n3135), .A2(n2611), .ZN(n3215) );
  OR2_X1 U3177 ( .A1(n2243), .A2(n2610), .ZN(n2611) );
  OR2_X1 U3178 ( .A1(n3216), .A2(n3217), .ZN(n3135) );
  AND2_X1 U3179 ( .A1(n3129), .A2(n3132), .ZN(n3217) );
  AND2_X1 U3180 ( .A1(n3218), .A2(n3219), .ZN(n3216) );
  OR2_X1 U3181 ( .A1(n3132), .A2(n3129), .ZN(n3219) );
  OR2_X1 U3182 ( .A1(n2218), .A2(n2610), .ZN(n3129) );
  OR3_X1 U3183 ( .A1(n2610), .A2(n2606), .A3(n2913), .ZN(n3132) );
  INV_X1 U3184 ( .A(b_12_), .ZN(n2610) );
  INV_X1 U3185 ( .A(n3131), .ZN(n3218) );
  OR2_X1 U3186 ( .A1(n3220), .A2(n3221), .ZN(n3131) );
  AND2_X1 U3187 ( .A1(b_11_), .A2(n3222), .ZN(n3221) );
  OR2_X1 U3188 ( .A1(n3223), .A2(n2918), .ZN(n3222) );
  AND2_X1 U3189 ( .A1(a_14_), .A2(n2602), .ZN(n3223) );
  AND2_X1 U3190 ( .A1(b_10_), .A2(n3224), .ZN(n3220) );
  OR2_X1 U3191 ( .A1(n3225), .A2(n2180), .ZN(n3224) );
  AND2_X1 U3192 ( .A1(a_15_), .A2(n2606), .ZN(n3225) );
  XNOR2_X1 U3193 ( .A(n3226), .B(n3227), .ZN(n3133) );
  XOR2_X1 U3194 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR2_X1 U3195 ( .A(n3230), .B(n3231), .Z(n3136) );
  XOR2_X1 U3196 ( .A(n3232), .B(n3233), .Z(n3231) );
  XOR2_X1 U3197 ( .A(n3234), .B(n3235), .Z(n3140) );
  XOR2_X1 U3198 ( .A(n3236), .B(n2607), .Z(n3235) );
  XOR2_X1 U3199 ( .A(n3237), .B(n3238), .Z(n3144) );
  XOR2_X1 U3200 ( .A(n3239), .B(n3240), .Z(n3238) );
  XOR2_X1 U3201 ( .A(n3241), .B(n3242), .Z(n3148) );
  XOR2_X1 U3202 ( .A(n3243), .B(n3244), .Z(n3242) );
  XOR2_X1 U3203 ( .A(n3245), .B(n3246), .Z(n3152) );
  XOR2_X1 U3204 ( .A(n3247), .B(n3248), .Z(n3246) );
  XOR2_X1 U3205 ( .A(n3249), .B(n3250), .Z(n3156) );
  XOR2_X1 U3206 ( .A(n3251), .B(n3252), .Z(n3250) );
  XOR2_X1 U3207 ( .A(n3253), .B(n3254), .Z(n3160) );
  XOR2_X1 U3208 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR2_X1 U3209 ( .A(n3257), .B(n3258), .Z(n3164) );
  XOR2_X1 U3210 ( .A(n3259), .B(n3260), .Z(n3258) );
  XOR2_X1 U3211 ( .A(n3261), .B(n3262), .Z(n3168) );
  XOR2_X1 U3212 ( .A(n3263), .B(n3264), .Z(n3262) );
  XOR2_X1 U3213 ( .A(n3265), .B(n3266), .Z(n3172) );
  XOR2_X1 U3214 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR2_X1 U3215 ( .A(n3269), .B(n3270), .Z(n2987) );
  XOR2_X1 U3216 ( .A(n3271), .B(n3272), .Z(n3270) );
  XOR2_X1 U3217 ( .A(n3273), .B(n3274), .Z(n2865) );
  XOR2_X1 U3218 ( .A(n3275), .B(n3276), .Z(n3274) );
  XNOR2_X1 U3219 ( .A(n3277), .B(n3278), .ZN(n2661) );
  XOR2_X1 U3220 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR2_X1 U3221 ( .A(n2672), .B(n2671), .Z(n2659) );
  INV_X1 U3222 ( .A(n3281), .ZN(n2671) );
  OR2_X1 U3223 ( .A1(n3282), .A2(n3283), .ZN(n3281) );
  AND2_X1 U3224 ( .A1(n3280), .A2(n3279), .ZN(n3283) );
  AND2_X1 U3225 ( .A1(n3277), .A2(n3284), .ZN(n3282) );
  OR2_X1 U3226 ( .A1(n3279), .A2(n3280), .ZN(n3284) );
  OR2_X1 U3227 ( .A1(n2969), .A2(n2606), .ZN(n3280) );
  OR2_X1 U3228 ( .A1(n3285), .A2(n3286), .ZN(n3279) );
  AND2_X1 U3229 ( .A1(n3276), .A2(n3275), .ZN(n3286) );
  AND2_X1 U3230 ( .A1(n3273), .A2(n3287), .ZN(n3285) );
  OR2_X1 U3231 ( .A1(n3275), .A2(n3276), .ZN(n3287) );
  OR2_X1 U3232 ( .A1(n2566), .A2(n2606), .ZN(n3276) );
  OR2_X1 U3233 ( .A1(n3288), .A2(n3289), .ZN(n3275) );
  AND2_X1 U3234 ( .A1(n3272), .A2(n3271), .ZN(n3289) );
  AND2_X1 U3235 ( .A1(n3269), .A2(n3290), .ZN(n3288) );
  OR2_X1 U3236 ( .A1(n3271), .A2(n3272), .ZN(n3290) );
  OR2_X1 U3237 ( .A1(n2570), .A2(n2606), .ZN(n3272) );
  OR2_X1 U3238 ( .A1(n3291), .A2(n3292), .ZN(n3271) );
  AND2_X1 U3239 ( .A1(n3268), .A2(n3267), .ZN(n3292) );
  AND2_X1 U3240 ( .A1(n3265), .A2(n3293), .ZN(n3291) );
  OR2_X1 U3241 ( .A1(n3267), .A2(n3268), .ZN(n3293) );
  OR2_X1 U3242 ( .A1(n2574), .A2(n2606), .ZN(n3268) );
  OR2_X1 U3243 ( .A1(n3294), .A2(n3295), .ZN(n3267) );
  AND2_X1 U3244 ( .A1(n3264), .A2(n3263), .ZN(n3295) );
  AND2_X1 U3245 ( .A1(n3261), .A2(n3296), .ZN(n3294) );
  OR2_X1 U3246 ( .A1(n3263), .A2(n3264), .ZN(n3296) );
  OR2_X1 U3247 ( .A1(n2578), .A2(n2606), .ZN(n3264) );
  OR2_X1 U3248 ( .A1(n3297), .A2(n3298), .ZN(n3263) );
  AND2_X1 U3249 ( .A1(n3260), .A2(n3259), .ZN(n3298) );
  AND2_X1 U3250 ( .A1(n3257), .A2(n3299), .ZN(n3297) );
  OR2_X1 U3251 ( .A1(n3259), .A2(n3260), .ZN(n3299) );
  OR2_X1 U3252 ( .A1(n2582), .A2(n2606), .ZN(n3260) );
  OR2_X1 U3253 ( .A1(n3300), .A2(n3301), .ZN(n3259) );
  AND2_X1 U3254 ( .A1(n3256), .A2(n3255), .ZN(n3301) );
  AND2_X1 U3255 ( .A1(n3253), .A2(n3302), .ZN(n3300) );
  OR2_X1 U3256 ( .A1(n3255), .A2(n3256), .ZN(n3302) );
  OR2_X1 U3257 ( .A1(n2586), .A2(n2606), .ZN(n3256) );
  OR2_X1 U3258 ( .A1(n3303), .A2(n3304), .ZN(n3255) );
  AND2_X1 U3259 ( .A1(n3252), .A2(n3251), .ZN(n3304) );
  AND2_X1 U3260 ( .A1(n3249), .A2(n3305), .ZN(n3303) );
  OR2_X1 U3261 ( .A1(n3251), .A2(n3252), .ZN(n3305) );
  OR2_X1 U3262 ( .A1(n2590), .A2(n2606), .ZN(n3252) );
  OR2_X1 U3263 ( .A1(n3306), .A2(n3307), .ZN(n3251) );
  AND2_X1 U3264 ( .A1(n3248), .A2(n3247), .ZN(n3307) );
  AND2_X1 U3265 ( .A1(n3245), .A2(n3308), .ZN(n3306) );
  OR2_X1 U3266 ( .A1(n3247), .A2(n3248), .ZN(n3308) );
  OR2_X1 U3267 ( .A1(n2594), .A2(n2606), .ZN(n3248) );
  OR2_X1 U3268 ( .A1(n3309), .A2(n3310), .ZN(n3247) );
  AND2_X1 U3269 ( .A1(n3244), .A2(n3243), .ZN(n3310) );
  AND2_X1 U3270 ( .A1(n3241), .A2(n3311), .ZN(n3309) );
  OR2_X1 U3271 ( .A1(n3243), .A2(n3244), .ZN(n3311) );
  OR2_X1 U3272 ( .A1(n2318), .A2(n2606), .ZN(n3244) );
  OR2_X1 U3273 ( .A1(n3312), .A2(n3313), .ZN(n3243) );
  AND2_X1 U3274 ( .A1(n3240), .A2(n3239), .ZN(n3313) );
  AND2_X1 U3275 ( .A1(n3237), .A2(n3314), .ZN(n3312) );
  OR2_X1 U3276 ( .A1(n3239), .A2(n3240), .ZN(n3314) );
  OR2_X1 U3277 ( .A1(n2293), .A2(n2606), .ZN(n3240) );
  OR2_X1 U3278 ( .A1(n3315), .A2(n3316), .ZN(n3239) );
  AND2_X1 U3279 ( .A1(n2607), .A2(n3236), .ZN(n3316) );
  AND2_X1 U3280 ( .A1(n3234), .A2(n3317), .ZN(n3315) );
  OR2_X1 U3281 ( .A1(n3236), .A2(n2607), .ZN(n3317) );
  OR2_X1 U3282 ( .A1(n2268), .A2(n2606), .ZN(n2607) );
  OR2_X1 U3283 ( .A1(n3318), .A2(n3319), .ZN(n3236) );
  AND2_X1 U3284 ( .A1(n3233), .A2(n3232), .ZN(n3319) );
  AND2_X1 U3285 ( .A1(n3230), .A2(n3320), .ZN(n3318) );
  OR2_X1 U3286 ( .A1(n3232), .A2(n3233), .ZN(n3320) );
  OR2_X1 U3287 ( .A1(n2243), .A2(n2606), .ZN(n3233) );
  OR2_X1 U3288 ( .A1(n3321), .A2(n3322), .ZN(n3232) );
  AND2_X1 U3289 ( .A1(n3226), .A2(n3229), .ZN(n3322) );
  AND2_X1 U3290 ( .A1(n3323), .A2(n3324), .ZN(n3321) );
  OR2_X1 U3291 ( .A1(n3229), .A2(n3226), .ZN(n3324) );
  OR2_X1 U3292 ( .A1(n2218), .A2(n2606), .ZN(n3226) );
  OR3_X1 U3293 ( .A1(n2606), .A2(n2602), .A3(n2913), .ZN(n3229) );
  INV_X1 U3294 ( .A(b_11_), .ZN(n2606) );
  INV_X1 U3295 ( .A(n3228), .ZN(n3323) );
  OR2_X1 U3296 ( .A1(n3325), .A2(n3326), .ZN(n3228) );
  AND2_X1 U3297 ( .A1(b_9_), .A2(n3327), .ZN(n3326) );
  OR2_X1 U3298 ( .A1(n3328), .A2(n2180), .ZN(n3327) );
  AND2_X1 U3299 ( .A1(a_15_), .A2(n2602), .ZN(n3328) );
  AND2_X1 U3300 ( .A1(b_10_), .A2(n3329), .ZN(n3325) );
  OR2_X1 U3301 ( .A1(n3330), .A2(n2918), .ZN(n3329) );
  AND2_X1 U3302 ( .A1(a_14_), .A2(n2598), .ZN(n3330) );
  XNOR2_X1 U3303 ( .A(n3331), .B(n3332), .ZN(n3230) );
  XOR2_X1 U3304 ( .A(n3333), .B(n3334), .Z(n3332) );
  XOR2_X1 U3305 ( .A(n3335), .B(n3336), .Z(n3234) );
  XOR2_X1 U3306 ( .A(n3337), .B(n3338), .Z(n3336) );
  XOR2_X1 U3307 ( .A(n3339), .B(n3340), .Z(n3237) );
  XOR2_X1 U3308 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR2_X1 U3309 ( .A(n3343), .B(n3344), .Z(n3241) );
  XOR2_X1 U3310 ( .A(n3345), .B(n2603), .Z(n3344) );
  XOR2_X1 U3311 ( .A(n3346), .B(n3347), .Z(n3245) );
  XOR2_X1 U3312 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR2_X1 U3313 ( .A(n3350), .B(n3351), .Z(n3249) );
  XOR2_X1 U3314 ( .A(n3352), .B(n3353), .Z(n3351) );
  XOR2_X1 U3315 ( .A(n3354), .B(n3355), .Z(n3253) );
  XOR2_X1 U3316 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR2_X1 U3317 ( .A(n3358), .B(n3359), .Z(n3257) );
  XOR2_X1 U3318 ( .A(n3360), .B(n3361), .Z(n3359) );
  XOR2_X1 U3319 ( .A(n3362), .B(n3363), .Z(n3261) );
  XOR2_X1 U3320 ( .A(n3364), .B(n3365), .Z(n3363) );
  XOR2_X1 U3321 ( .A(n3366), .B(n3367), .Z(n3265) );
  XOR2_X1 U3322 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR2_X1 U3323 ( .A(n3370), .B(n3371), .Z(n3269) );
  XOR2_X1 U3324 ( .A(n3372), .B(n3373), .Z(n3371) );
  XOR2_X1 U3325 ( .A(n3374), .B(n3375), .Z(n3273) );
  XOR2_X1 U3326 ( .A(n3376), .B(n3377), .Z(n3375) );
  XOR2_X1 U3327 ( .A(n3378), .B(n3379), .Z(n3277) );
  XOR2_X1 U3328 ( .A(n3380), .B(n3381), .Z(n3379) );
  XNOR2_X1 U3329 ( .A(n3382), .B(n3383), .ZN(n2672) );
  XOR2_X1 U3330 ( .A(n3384), .B(n3385), .Z(n3383) );
  AND2_X1 U3331 ( .A1(n3386), .A2(n2848), .ZN(n2669) );
  OR2_X1 U3332 ( .A1(n3387), .A2(n3388), .ZN(n2848) );
  INV_X1 U3333 ( .A(n3389), .ZN(n3386) );
  AND2_X1 U3334 ( .A1(n3387), .A2(n3388), .ZN(n3389) );
  OR2_X1 U3335 ( .A1(n3390), .A2(n3391), .ZN(n3388) );
  AND2_X1 U3336 ( .A1(n3385), .A2(n3384), .ZN(n3391) );
  AND2_X1 U3337 ( .A1(n3382), .A2(n3392), .ZN(n3390) );
  OR2_X1 U3338 ( .A1(n3385), .A2(n3384), .ZN(n3392) );
  OR2_X1 U3339 ( .A1(n3393), .A2(n3394), .ZN(n3384) );
  AND2_X1 U3340 ( .A1(n3381), .A2(n3380), .ZN(n3394) );
  AND2_X1 U3341 ( .A1(n3378), .A2(n3395), .ZN(n3393) );
  OR2_X1 U3342 ( .A1(n3381), .A2(n3380), .ZN(n3395) );
  OR2_X1 U3343 ( .A1(n3396), .A2(n3397), .ZN(n3380) );
  AND2_X1 U3344 ( .A1(n3377), .A2(n3376), .ZN(n3397) );
  AND2_X1 U3345 ( .A1(n3374), .A2(n3398), .ZN(n3396) );
  OR2_X1 U3346 ( .A1(n3377), .A2(n3376), .ZN(n3398) );
  OR2_X1 U3347 ( .A1(n3399), .A2(n3400), .ZN(n3376) );
  AND2_X1 U3348 ( .A1(n3370), .A2(n3373), .ZN(n3400) );
  AND2_X1 U3349 ( .A1(n3401), .A2(n3372), .ZN(n3399) );
  OR2_X1 U3350 ( .A1(n3402), .A2(n3403), .ZN(n3372) );
  AND2_X1 U3351 ( .A1(n3369), .A2(n3368), .ZN(n3403) );
  AND2_X1 U3352 ( .A1(n3366), .A2(n3404), .ZN(n3402) );
  OR2_X1 U3353 ( .A1(n3369), .A2(n3368), .ZN(n3404) );
  OR2_X1 U3354 ( .A1(n3405), .A2(n3406), .ZN(n3368) );
  AND2_X1 U3355 ( .A1(n3362), .A2(n3365), .ZN(n3406) );
  AND2_X1 U3356 ( .A1(n3407), .A2(n3364), .ZN(n3405) );
  OR2_X1 U3357 ( .A1(n3408), .A2(n3409), .ZN(n3364) );
  AND2_X1 U3358 ( .A1(n3358), .A2(n3361), .ZN(n3409) );
  AND2_X1 U3359 ( .A1(n3410), .A2(n3360), .ZN(n3408) );
  OR2_X1 U3360 ( .A1(n3411), .A2(n3412), .ZN(n3360) );
  AND2_X1 U3361 ( .A1(n3354), .A2(n3357), .ZN(n3412) );
  AND2_X1 U3362 ( .A1(n3413), .A2(n3356), .ZN(n3411) );
  OR2_X1 U3363 ( .A1(n3414), .A2(n3415), .ZN(n3356) );
  AND2_X1 U3364 ( .A1(n3350), .A2(n3353), .ZN(n3415) );
  AND2_X1 U3365 ( .A1(n3416), .A2(n3352), .ZN(n3414) );
  OR2_X1 U3366 ( .A1(n3417), .A2(n3418), .ZN(n3352) );
  AND2_X1 U3367 ( .A1(n3346), .A2(n3349), .ZN(n3418) );
  AND2_X1 U3368 ( .A1(n3419), .A2(n3348), .ZN(n3417) );
  OR2_X1 U3369 ( .A1(n3420), .A2(n3421), .ZN(n3348) );
  AND2_X1 U3370 ( .A1(n3343), .A2(n2603), .ZN(n3421) );
  AND2_X1 U3371 ( .A1(n3422), .A2(n3345), .ZN(n3420) );
  OR2_X1 U3372 ( .A1(n3423), .A2(n3424), .ZN(n3345) );
  AND2_X1 U3373 ( .A1(n3339), .A2(n3342), .ZN(n3424) );
  AND2_X1 U3374 ( .A1(n3425), .A2(n3341), .ZN(n3423) );
  OR2_X1 U3375 ( .A1(n3426), .A2(n3427), .ZN(n3341) );
  AND2_X1 U3376 ( .A1(n3335), .A2(n3338), .ZN(n3427) );
  AND2_X1 U3377 ( .A1(n3428), .A2(n3337), .ZN(n3426) );
  OR2_X1 U3378 ( .A1(n3429), .A2(n3430), .ZN(n3337) );
  AND2_X1 U3379 ( .A1(n3331), .A2(n3334), .ZN(n3430) );
  AND2_X1 U3380 ( .A1(n3431), .A2(n3432), .ZN(n3429) );
  OR2_X1 U3381 ( .A1(n3331), .A2(n3334), .ZN(n3432) );
  OR3_X1 U3382 ( .A1(n2602), .A2(n2598), .A3(n2913), .ZN(n3334) );
  OR2_X1 U3383 ( .A1(n2218), .A2(n2602), .ZN(n3331) );
  INV_X1 U3384 ( .A(n3333), .ZN(n3431) );
  OR2_X1 U3385 ( .A1(n3433), .A2(n3434), .ZN(n3333) );
  AND2_X1 U3386 ( .A1(b_9_), .A2(n3435), .ZN(n3434) );
  OR2_X1 U3387 ( .A1(n3436), .A2(n2918), .ZN(n3435) );
  AND2_X1 U3388 ( .A1(a_14_), .A2(n2595), .ZN(n3436) );
  AND2_X1 U3389 ( .A1(b_8_), .A2(n3437), .ZN(n3433) );
  OR2_X1 U3390 ( .A1(n3438), .A2(n2180), .ZN(n3437) );
  AND2_X1 U3391 ( .A1(a_15_), .A2(n2598), .ZN(n3438) );
  OR2_X1 U3392 ( .A1(n3335), .A2(n3338), .ZN(n3428) );
  OR2_X1 U3393 ( .A1(n2243), .A2(n2602), .ZN(n3338) );
  XNOR2_X1 U3394 ( .A(n3439), .B(n3440), .ZN(n3335) );
  XOR2_X1 U3395 ( .A(n3441), .B(n3442), .Z(n3440) );
  OR2_X1 U3396 ( .A1(n3339), .A2(n3342), .ZN(n3425) );
  OR2_X1 U3397 ( .A1(n2268), .A2(n2602), .ZN(n3342) );
  XOR2_X1 U3398 ( .A(n3443), .B(n3444), .Z(n3339) );
  XOR2_X1 U3399 ( .A(n3445), .B(n3446), .Z(n3444) );
  OR2_X1 U3400 ( .A1(n3343), .A2(n2603), .ZN(n3422) );
  OR2_X1 U3401 ( .A1(n2293), .A2(n2602), .ZN(n2603) );
  XOR2_X1 U3402 ( .A(n3447), .B(n3448), .Z(n3343) );
  XOR2_X1 U3403 ( .A(n3449), .B(n3450), .Z(n3448) );
  OR2_X1 U3404 ( .A1(n3346), .A2(n3349), .ZN(n3419) );
  OR2_X1 U3405 ( .A1(n2318), .A2(n2602), .ZN(n3349) );
  XOR2_X1 U3406 ( .A(n3451), .B(n3452), .Z(n3346) );
  XOR2_X1 U3407 ( .A(n3453), .B(n3454), .Z(n3452) );
  OR2_X1 U3408 ( .A1(n3350), .A2(n3353), .ZN(n3416) );
  OR2_X1 U3409 ( .A1(n2594), .A2(n2602), .ZN(n3353) );
  XOR2_X1 U3410 ( .A(n3455), .B(n3456), .Z(n3350) );
  XOR2_X1 U3411 ( .A(n3457), .B(n2599), .Z(n3456) );
  OR2_X1 U3412 ( .A1(n3354), .A2(n3357), .ZN(n3413) );
  OR2_X1 U3413 ( .A1(n2590), .A2(n2602), .ZN(n3357) );
  XOR2_X1 U3414 ( .A(n3458), .B(n3459), .Z(n3354) );
  XOR2_X1 U3415 ( .A(n3460), .B(n3461), .Z(n3459) );
  OR2_X1 U3416 ( .A1(n3358), .A2(n3361), .ZN(n3410) );
  OR2_X1 U3417 ( .A1(n2586), .A2(n2602), .ZN(n3361) );
  XOR2_X1 U3418 ( .A(n3462), .B(n3463), .Z(n3358) );
  XOR2_X1 U3419 ( .A(n3464), .B(n3465), .Z(n3463) );
  OR2_X1 U3420 ( .A1(n3362), .A2(n3365), .ZN(n3407) );
  OR2_X1 U3421 ( .A1(n2582), .A2(n2602), .ZN(n3365) );
  XOR2_X1 U3422 ( .A(n3466), .B(n3467), .Z(n3362) );
  XOR2_X1 U3423 ( .A(n3468), .B(n3469), .Z(n3467) );
  OR2_X1 U3424 ( .A1(n2578), .A2(n2602), .ZN(n3369) );
  XOR2_X1 U3425 ( .A(n3470), .B(n3471), .Z(n3366) );
  XOR2_X1 U3426 ( .A(n3472), .B(n3473), .Z(n3471) );
  OR2_X1 U3427 ( .A1(n3370), .A2(n3373), .ZN(n3401) );
  OR2_X1 U3428 ( .A1(n2574), .A2(n2602), .ZN(n3373) );
  XOR2_X1 U3429 ( .A(n3474), .B(n3475), .Z(n3370) );
  XOR2_X1 U3430 ( .A(n3476), .B(n3477), .Z(n3475) );
  OR2_X1 U3431 ( .A1(n2570), .A2(n2602), .ZN(n3377) );
  XOR2_X1 U3432 ( .A(n3478), .B(n3479), .Z(n3374) );
  XOR2_X1 U3433 ( .A(n3480), .B(n3481), .Z(n3479) );
  OR2_X1 U3434 ( .A1(n2566), .A2(n2602), .ZN(n3381) );
  XOR2_X1 U3435 ( .A(n3482), .B(n3483), .Z(n3378) );
  XOR2_X1 U3436 ( .A(n3484), .B(n3485), .Z(n3483) );
  OR2_X1 U3437 ( .A1(n2969), .A2(n2602), .ZN(n3385) );
  INV_X1 U3438 ( .A(b_10_), .ZN(n2602) );
  XOR2_X1 U3439 ( .A(n3486), .B(n3487), .Z(n3382) );
  XOR2_X1 U3440 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR2_X1 U3441 ( .A(n3490), .B(n3491), .Z(n3387) );
  XOR2_X1 U3442 ( .A(n3492), .B(n3493), .Z(n3491) );
  INV_X1 U3443 ( .A(n3494), .ZN(n2840) );
  OR2_X1 U3444 ( .A1(n2844), .A2(n2845), .ZN(n3494) );
  OR2_X1 U3445 ( .A1(n3495), .A2(n3496), .ZN(n2845) );
  AND2_X1 U3446 ( .A1(n3493), .A2(n3492), .ZN(n3496) );
  AND2_X1 U3447 ( .A1(n3490), .A2(n3497), .ZN(n3495) );
  OR2_X1 U3448 ( .A1(n3493), .A2(n3492), .ZN(n3497) );
  OR2_X1 U3449 ( .A1(n3498), .A2(n3499), .ZN(n3492) );
  AND2_X1 U3450 ( .A1(n3489), .A2(n3488), .ZN(n3499) );
  AND2_X1 U3451 ( .A1(n3486), .A2(n3500), .ZN(n3498) );
  OR2_X1 U3452 ( .A1(n3489), .A2(n3488), .ZN(n3500) );
  OR2_X1 U3453 ( .A1(n3501), .A2(n3502), .ZN(n3488) );
  AND2_X1 U3454 ( .A1(n3485), .A2(n3484), .ZN(n3502) );
  AND2_X1 U3455 ( .A1(n3482), .A2(n3503), .ZN(n3501) );
  OR2_X1 U3456 ( .A1(n3485), .A2(n3484), .ZN(n3503) );
  OR2_X1 U3457 ( .A1(n3504), .A2(n3505), .ZN(n3484) );
  AND2_X1 U3458 ( .A1(n3481), .A2(n3480), .ZN(n3505) );
  AND2_X1 U3459 ( .A1(n3478), .A2(n3506), .ZN(n3504) );
  OR2_X1 U3460 ( .A1(n3481), .A2(n3480), .ZN(n3506) );
  OR2_X1 U3461 ( .A1(n3507), .A2(n3508), .ZN(n3480) );
  AND2_X1 U3462 ( .A1(n3474), .A2(n3477), .ZN(n3508) );
  AND2_X1 U3463 ( .A1(n3509), .A2(n3476), .ZN(n3507) );
  OR2_X1 U3464 ( .A1(n3510), .A2(n3511), .ZN(n3476) );
  AND2_X1 U3465 ( .A1(n3473), .A2(n3472), .ZN(n3511) );
  AND2_X1 U3466 ( .A1(n3470), .A2(n3512), .ZN(n3510) );
  OR2_X1 U3467 ( .A1(n3473), .A2(n3472), .ZN(n3512) );
  OR2_X1 U3468 ( .A1(n3513), .A2(n3514), .ZN(n3472) );
  AND2_X1 U3469 ( .A1(n3466), .A2(n3469), .ZN(n3514) );
  AND2_X1 U3470 ( .A1(n3515), .A2(n3468), .ZN(n3513) );
  OR2_X1 U3471 ( .A1(n3516), .A2(n3517), .ZN(n3468) );
  AND2_X1 U3472 ( .A1(n3462), .A2(n3465), .ZN(n3517) );
  AND2_X1 U3473 ( .A1(n3518), .A2(n3464), .ZN(n3516) );
  OR2_X1 U3474 ( .A1(n3519), .A2(n3520), .ZN(n3464) );
  AND2_X1 U3475 ( .A1(n3458), .A2(n3461), .ZN(n3520) );
  AND2_X1 U3476 ( .A1(n3521), .A2(n3460), .ZN(n3519) );
  OR2_X1 U3477 ( .A1(n3522), .A2(n3523), .ZN(n3460) );
  AND2_X1 U3478 ( .A1(n3455), .A2(n2599), .ZN(n3523) );
  AND2_X1 U3479 ( .A1(n3524), .A2(n3457), .ZN(n3522) );
  OR2_X1 U3480 ( .A1(n3525), .A2(n3526), .ZN(n3457) );
  AND2_X1 U3481 ( .A1(n3451), .A2(n3454), .ZN(n3526) );
  AND2_X1 U3482 ( .A1(n3527), .A2(n3453), .ZN(n3525) );
  OR2_X1 U3483 ( .A1(n3528), .A2(n3529), .ZN(n3453) );
  AND2_X1 U3484 ( .A1(n3447), .A2(n3450), .ZN(n3529) );
  AND2_X1 U3485 ( .A1(n3530), .A2(n3449), .ZN(n3528) );
  OR2_X1 U3486 ( .A1(n3531), .A2(n3532), .ZN(n3449) );
  AND2_X1 U3487 ( .A1(n3443), .A2(n3446), .ZN(n3532) );
  AND2_X1 U3488 ( .A1(n3533), .A2(n3445), .ZN(n3531) );
  OR2_X1 U3489 ( .A1(n3534), .A2(n3535), .ZN(n3445) );
  AND2_X1 U3490 ( .A1(n3439), .A2(n3442), .ZN(n3535) );
  AND2_X1 U3491 ( .A1(n3536), .A2(n3537), .ZN(n3534) );
  OR2_X1 U3492 ( .A1(n3439), .A2(n3442), .ZN(n3537) );
  OR3_X1 U3493 ( .A1(n2598), .A2(n2595), .A3(n2913), .ZN(n3442) );
  OR2_X1 U3494 ( .A1(n2218), .A2(n2598), .ZN(n3439) );
  INV_X1 U3495 ( .A(n3441), .ZN(n3536) );
  OR2_X1 U3496 ( .A1(n3538), .A2(n3539), .ZN(n3441) );
  AND2_X1 U3497 ( .A1(b_8_), .A2(n3540), .ZN(n3539) );
  OR2_X1 U3498 ( .A1(n3541), .A2(n2918), .ZN(n3540) );
  AND2_X1 U3499 ( .A1(a_14_), .A2(n2591), .ZN(n3541) );
  AND2_X1 U3500 ( .A1(b_7_), .A2(n3542), .ZN(n3538) );
  OR2_X1 U3501 ( .A1(n3543), .A2(n2180), .ZN(n3542) );
  AND2_X1 U3502 ( .A1(a_15_), .A2(n2595), .ZN(n3543) );
  OR2_X1 U3503 ( .A1(n3443), .A2(n3446), .ZN(n3533) );
  OR2_X1 U3504 ( .A1(n2243), .A2(n2598), .ZN(n3446) );
  XNOR2_X1 U3505 ( .A(n3544), .B(n3545), .ZN(n3443) );
  XOR2_X1 U3506 ( .A(n3546), .B(n3547), .Z(n3545) );
  OR2_X1 U3507 ( .A1(n3447), .A2(n3450), .ZN(n3530) );
  OR2_X1 U3508 ( .A1(n2268), .A2(n2598), .ZN(n3450) );
  XOR2_X1 U3509 ( .A(n3548), .B(n3549), .Z(n3447) );
  XOR2_X1 U3510 ( .A(n3550), .B(n3551), .Z(n3549) );
  OR2_X1 U3511 ( .A1(n3451), .A2(n3454), .ZN(n3527) );
  OR2_X1 U3512 ( .A1(n2293), .A2(n2598), .ZN(n3454) );
  XOR2_X1 U3513 ( .A(n3552), .B(n3553), .Z(n3451) );
  XOR2_X1 U3514 ( .A(n3554), .B(n3555), .Z(n3553) );
  OR2_X1 U3515 ( .A1(n3455), .A2(n2599), .ZN(n3524) );
  OR2_X1 U3516 ( .A1(n2318), .A2(n2598), .ZN(n2599) );
  XOR2_X1 U3517 ( .A(n3556), .B(n3557), .Z(n3455) );
  XOR2_X1 U3518 ( .A(n3558), .B(n3559), .Z(n3557) );
  OR2_X1 U3519 ( .A1(n3458), .A2(n3461), .ZN(n3521) );
  OR2_X1 U3520 ( .A1(n2594), .A2(n2598), .ZN(n3461) );
  XOR2_X1 U3521 ( .A(n3560), .B(n3561), .Z(n3458) );
  XOR2_X1 U3522 ( .A(n3562), .B(n3563), .Z(n3561) );
  OR2_X1 U3523 ( .A1(n3462), .A2(n3465), .ZN(n3518) );
  OR2_X1 U3524 ( .A1(n2590), .A2(n2598), .ZN(n3465) );
  XOR2_X1 U3525 ( .A(n3564), .B(n3565), .Z(n3462) );
  XOR2_X1 U3526 ( .A(n3566), .B(n2340), .Z(n3565) );
  OR2_X1 U3527 ( .A1(n3466), .A2(n3469), .ZN(n3515) );
  OR2_X1 U3528 ( .A1(n2586), .A2(n2598), .ZN(n3469) );
  XOR2_X1 U3529 ( .A(n3567), .B(n3568), .Z(n3466) );
  XOR2_X1 U3530 ( .A(n3569), .B(n3570), .Z(n3568) );
  OR2_X1 U3531 ( .A1(n2582), .A2(n2598), .ZN(n3473) );
  XOR2_X1 U3532 ( .A(n3571), .B(n3572), .Z(n3470) );
  XOR2_X1 U3533 ( .A(n3573), .B(n3574), .Z(n3572) );
  OR2_X1 U3534 ( .A1(n3474), .A2(n3477), .ZN(n3509) );
  OR2_X1 U3535 ( .A1(n2578), .A2(n2598), .ZN(n3477) );
  XOR2_X1 U3536 ( .A(n3575), .B(n3576), .Z(n3474) );
  XOR2_X1 U3537 ( .A(n3577), .B(n3578), .Z(n3576) );
  OR2_X1 U3538 ( .A1(n2574), .A2(n2598), .ZN(n3481) );
  XOR2_X1 U3539 ( .A(n3579), .B(n3580), .Z(n3478) );
  XOR2_X1 U3540 ( .A(n3581), .B(n3582), .Z(n3580) );
  OR2_X1 U3541 ( .A1(n2570), .A2(n2598), .ZN(n3485) );
  XOR2_X1 U3542 ( .A(n3583), .B(n3584), .Z(n3482) );
  XOR2_X1 U3543 ( .A(n3585), .B(n3586), .Z(n3584) );
  OR2_X1 U3544 ( .A1(n2566), .A2(n2598), .ZN(n3489) );
  XOR2_X1 U3545 ( .A(n3587), .B(n3588), .Z(n3486) );
  XOR2_X1 U3546 ( .A(n3589), .B(n3590), .Z(n3588) );
  OR2_X1 U3547 ( .A1(n2969), .A2(n2598), .ZN(n3493) );
  INV_X1 U3548 ( .A(b_9_), .ZN(n2598) );
  XOR2_X1 U3549 ( .A(n3591), .B(n3592), .Z(n3490) );
  XOR2_X1 U3550 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR2_X1 U3551 ( .A(n2834), .B(n3595), .Z(n2844) );
  XOR2_X1 U3552 ( .A(n2833), .B(n2832), .Z(n3595) );
  OR2_X1 U3553 ( .A1(n2969), .A2(n2595), .ZN(n2832) );
  OR2_X1 U3554 ( .A1(n3596), .A2(n3597), .ZN(n2833) );
  AND2_X1 U3555 ( .A1(n3594), .A2(n3593), .ZN(n3597) );
  AND2_X1 U3556 ( .A1(n3591), .A2(n3598), .ZN(n3596) );
  OR2_X1 U3557 ( .A1(n3593), .A2(n3594), .ZN(n3598) );
  OR2_X1 U3558 ( .A1(n2566), .A2(n2595), .ZN(n3594) );
  OR2_X1 U3559 ( .A1(n3599), .A2(n3600), .ZN(n3593) );
  AND2_X1 U3560 ( .A1(n3590), .A2(n3589), .ZN(n3600) );
  AND2_X1 U3561 ( .A1(n3587), .A2(n3601), .ZN(n3599) );
  OR2_X1 U3562 ( .A1(n3589), .A2(n3590), .ZN(n3601) );
  OR2_X1 U3563 ( .A1(n2570), .A2(n2595), .ZN(n3590) );
  OR2_X1 U3564 ( .A1(n3602), .A2(n3603), .ZN(n3589) );
  AND2_X1 U3565 ( .A1(n3586), .A2(n3585), .ZN(n3603) );
  AND2_X1 U3566 ( .A1(n3583), .A2(n3604), .ZN(n3602) );
  OR2_X1 U3567 ( .A1(n3585), .A2(n3586), .ZN(n3604) );
  OR2_X1 U3568 ( .A1(n2574), .A2(n2595), .ZN(n3586) );
  OR2_X1 U3569 ( .A1(n3605), .A2(n3606), .ZN(n3585) );
  AND2_X1 U3570 ( .A1(n3582), .A2(n3581), .ZN(n3606) );
  AND2_X1 U3571 ( .A1(n3579), .A2(n3607), .ZN(n3605) );
  OR2_X1 U3572 ( .A1(n3581), .A2(n3582), .ZN(n3607) );
  OR2_X1 U3573 ( .A1(n2578), .A2(n2595), .ZN(n3582) );
  OR2_X1 U3574 ( .A1(n3608), .A2(n3609), .ZN(n3581) );
  AND2_X1 U3575 ( .A1(n3575), .A2(n3578), .ZN(n3609) );
  AND2_X1 U3576 ( .A1(n3610), .A2(n3577), .ZN(n3608) );
  OR2_X1 U3577 ( .A1(n3611), .A2(n3612), .ZN(n3577) );
  AND2_X1 U3578 ( .A1(n3574), .A2(n3573), .ZN(n3612) );
  AND2_X1 U3579 ( .A1(n3571), .A2(n3613), .ZN(n3611) );
  OR2_X1 U3580 ( .A1(n3573), .A2(n3574), .ZN(n3613) );
  OR2_X1 U3581 ( .A1(n2586), .A2(n2595), .ZN(n3574) );
  OR2_X1 U3582 ( .A1(n3614), .A2(n3615), .ZN(n3573) );
  AND2_X1 U3583 ( .A1(n3567), .A2(n3570), .ZN(n3615) );
  AND2_X1 U3584 ( .A1(n3616), .A2(n3569), .ZN(n3614) );
  OR2_X1 U3585 ( .A1(n3617), .A2(n3618), .ZN(n3569) );
  AND2_X1 U3586 ( .A1(n3564), .A2(n2340), .ZN(n3618) );
  AND2_X1 U3587 ( .A1(n3619), .A2(n3566), .ZN(n3617) );
  OR2_X1 U3588 ( .A1(n3620), .A2(n3621), .ZN(n3566) );
  AND2_X1 U3589 ( .A1(n3560), .A2(n3563), .ZN(n3621) );
  AND2_X1 U3590 ( .A1(n3622), .A2(n3562), .ZN(n3620) );
  OR2_X1 U3591 ( .A1(n3623), .A2(n3624), .ZN(n3562) );
  AND2_X1 U3592 ( .A1(n3556), .A2(n3559), .ZN(n3624) );
  AND2_X1 U3593 ( .A1(n3625), .A2(n3558), .ZN(n3623) );
  OR2_X1 U3594 ( .A1(n3626), .A2(n3627), .ZN(n3558) );
  AND2_X1 U3595 ( .A1(n3552), .A2(n3555), .ZN(n3627) );
  AND2_X1 U3596 ( .A1(n3628), .A2(n3554), .ZN(n3626) );
  OR2_X1 U3597 ( .A1(n3629), .A2(n3630), .ZN(n3554) );
  AND2_X1 U3598 ( .A1(n3548), .A2(n3551), .ZN(n3630) );
  AND2_X1 U3599 ( .A1(n3631), .A2(n3550), .ZN(n3629) );
  OR2_X1 U3600 ( .A1(n3632), .A2(n3633), .ZN(n3550) );
  AND2_X1 U3601 ( .A1(n3544), .A2(n3547), .ZN(n3633) );
  AND2_X1 U3602 ( .A1(n3634), .A2(n3635), .ZN(n3632) );
  OR2_X1 U3603 ( .A1(n3547), .A2(n3544), .ZN(n3635) );
  OR2_X1 U3604 ( .A1(n2218), .A2(n2595), .ZN(n3544) );
  OR3_X1 U3605 ( .A1(n2595), .A2(n2591), .A3(n2913), .ZN(n3547) );
  INV_X1 U3606 ( .A(n3546), .ZN(n3634) );
  OR2_X1 U3607 ( .A1(n3636), .A2(n3637), .ZN(n3546) );
  AND2_X1 U3608 ( .A1(b_7_), .A2(n3638), .ZN(n3637) );
  OR2_X1 U3609 ( .A1(n3639), .A2(n2918), .ZN(n3638) );
  AND2_X1 U3610 ( .A1(a_14_), .A2(n2587), .ZN(n3639) );
  AND2_X1 U3611 ( .A1(b_6_), .A2(n3640), .ZN(n3636) );
  OR2_X1 U3612 ( .A1(n3641), .A2(n2180), .ZN(n3640) );
  AND2_X1 U3613 ( .A1(a_15_), .A2(n2591), .ZN(n3641) );
  OR2_X1 U3614 ( .A1(n3551), .A2(n3548), .ZN(n3631) );
  XNOR2_X1 U3615 ( .A(n3642), .B(n3643), .ZN(n3548) );
  XOR2_X1 U3616 ( .A(n3644), .B(n3645), .Z(n3643) );
  OR2_X1 U3617 ( .A1(n2243), .A2(n2595), .ZN(n3551) );
  OR2_X1 U3618 ( .A1(n3555), .A2(n3552), .ZN(n3628) );
  XOR2_X1 U3619 ( .A(n3646), .B(n3647), .Z(n3552) );
  XOR2_X1 U3620 ( .A(n3648), .B(n3649), .Z(n3647) );
  OR2_X1 U3621 ( .A1(n2268), .A2(n2595), .ZN(n3555) );
  OR2_X1 U3622 ( .A1(n3559), .A2(n3556), .ZN(n3625) );
  XOR2_X1 U3623 ( .A(n3650), .B(n3651), .Z(n3556) );
  XOR2_X1 U3624 ( .A(n3652), .B(n3653), .Z(n3651) );
  OR2_X1 U3625 ( .A1(n2293), .A2(n2595), .ZN(n3559) );
  OR2_X1 U3626 ( .A1(n3563), .A2(n3560), .ZN(n3622) );
  XOR2_X1 U3627 ( .A(n3654), .B(n3655), .Z(n3560) );
  XOR2_X1 U3628 ( .A(n3656), .B(n3657), .Z(n3655) );
  OR2_X1 U3629 ( .A1(n2318), .A2(n2595), .ZN(n3563) );
  OR2_X1 U3630 ( .A1(n2340), .A2(n3564), .ZN(n3619) );
  XOR2_X1 U3631 ( .A(n3658), .B(n3659), .Z(n3564) );
  XOR2_X1 U3632 ( .A(n3660), .B(n3661), .Z(n3659) );
  OR2_X1 U3633 ( .A1(n2594), .A2(n2595), .ZN(n2340) );
  OR2_X1 U3634 ( .A1(n3570), .A2(n3567), .ZN(n3616) );
  XOR2_X1 U3635 ( .A(n3662), .B(n3663), .Z(n3567) );
  XOR2_X1 U3636 ( .A(n3664), .B(n3665), .Z(n3663) );
  OR2_X1 U3637 ( .A1(n2590), .A2(n2595), .ZN(n3570) );
  XOR2_X1 U3638 ( .A(n3666), .B(n3667), .Z(n3571) );
  XOR2_X1 U3639 ( .A(n3668), .B(n2366), .Z(n3667) );
  OR2_X1 U3640 ( .A1(n3578), .A2(n3575), .ZN(n3610) );
  XOR2_X1 U3641 ( .A(n3669), .B(n3670), .Z(n3575) );
  XOR2_X1 U3642 ( .A(n3671), .B(n3672), .Z(n3670) );
  OR2_X1 U3643 ( .A1(n2582), .A2(n2595), .ZN(n3578) );
  INV_X1 U3644 ( .A(b_8_), .ZN(n2595) );
  XOR2_X1 U3645 ( .A(n3673), .B(n3674), .Z(n3579) );
  XOR2_X1 U3646 ( .A(n3675), .B(n3676), .Z(n3674) );
  XOR2_X1 U3647 ( .A(n3677), .B(n3678), .Z(n3583) );
  XOR2_X1 U3648 ( .A(n3679), .B(n3680), .Z(n3678) );
  XOR2_X1 U3649 ( .A(n3681), .B(n3682), .Z(n3587) );
  XOR2_X1 U3650 ( .A(n3683), .B(n3684), .Z(n3682) );
  XOR2_X1 U3651 ( .A(n3685), .B(n3686), .Z(n3591) );
  XOR2_X1 U3652 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR2_X1 U3653 ( .A(n3689), .B(n3690), .Z(n2834) );
  XOR2_X1 U3654 ( .A(n3691), .B(n3692), .Z(n3690) );
  INV_X1 U3655 ( .A(n3693), .ZN(n2817) );
  OR2_X1 U3656 ( .A1(n2821), .A2(n2822), .ZN(n3693) );
  OR2_X1 U3657 ( .A1(n3694), .A2(n3695), .ZN(n2822) );
  AND2_X1 U3658 ( .A1(n2839), .A2(n2838), .ZN(n3695) );
  AND2_X1 U3659 ( .A1(n2836), .A2(n3696), .ZN(n3694) );
  OR2_X1 U3660 ( .A1(n2838), .A2(n2839), .ZN(n3696) );
  OR2_X1 U3661 ( .A1(n2969), .A2(n2591), .ZN(n2839) );
  OR2_X1 U3662 ( .A1(n3697), .A2(n3698), .ZN(n2838) );
  AND2_X1 U3663 ( .A1(n3692), .A2(n3691), .ZN(n3698) );
  AND2_X1 U3664 ( .A1(n3689), .A2(n3699), .ZN(n3697) );
  OR2_X1 U3665 ( .A1(n3691), .A2(n3692), .ZN(n3699) );
  OR2_X1 U3666 ( .A1(n2566), .A2(n2591), .ZN(n3692) );
  OR2_X1 U3667 ( .A1(n3700), .A2(n3701), .ZN(n3691) );
  AND2_X1 U3668 ( .A1(n3688), .A2(n3687), .ZN(n3701) );
  AND2_X1 U3669 ( .A1(n3685), .A2(n3702), .ZN(n3700) );
  OR2_X1 U3670 ( .A1(n3687), .A2(n3688), .ZN(n3702) );
  OR2_X1 U3671 ( .A1(n2570), .A2(n2591), .ZN(n3688) );
  OR2_X1 U3672 ( .A1(n3703), .A2(n3704), .ZN(n3687) );
  AND2_X1 U3673 ( .A1(n3684), .A2(n3683), .ZN(n3704) );
  AND2_X1 U3674 ( .A1(n3681), .A2(n3705), .ZN(n3703) );
  OR2_X1 U3675 ( .A1(n3683), .A2(n3684), .ZN(n3705) );
  OR2_X1 U3676 ( .A1(n2574), .A2(n2591), .ZN(n3684) );
  OR2_X1 U3677 ( .A1(n3706), .A2(n3707), .ZN(n3683) );
  AND2_X1 U3678 ( .A1(n3680), .A2(n3679), .ZN(n3707) );
  AND2_X1 U3679 ( .A1(n3677), .A2(n3708), .ZN(n3706) );
  OR2_X1 U3680 ( .A1(n3679), .A2(n3680), .ZN(n3708) );
  OR2_X1 U3681 ( .A1(n2578), .A2(n2591), .ZN(n3680) );
  OR2_X1 U3682 ( .A1(n3709), .A2(n3710), .ZN(n3679) );
  AND2_X1 U3683 ( .A1(n3676), .A2(n3675), .ZN(n3710) );
  AND2_X1 U3684 ( .A1(n3673), .A2(n3711), .ZN(n3709) );
  OR2_X1 U3685 ( .A1(n3675), .A2(n3676), .ZN(n3711) );
  OR2_X1 U3686 ( .A1(n2582), .A2(n2591), .ZN(n3676) );
  OR2_X1 U3687 ( .A1(n3712), .A2(n3713), .ZN(n3675) );
  AND2_X1 U3688 ( .A1(n3669), .A2(n3672), .ZN(n3713) );
  AND2_X1 U3689 ( .A1(n3714), .A2(n3671), .ZN(n3712) );
  OR2_X1 U3690 ( .A1(n3715), .A2(n3716), .ZN(n3671) );
  AND2_X1 U3691 ( .A1(n2366), .A2(n3668), .ZN(n3716) );
  AND2_X1 U3692 ( .A1(n3666), .A2(n3717), .ZN(n3715) );
  OR2_X1 U3693 ( .A1(n3668), .A2(n2366), .ZN(n3717) );
  OR2_X1 U3694 ( .A1(n2590), .A2(n2591), .ZN(n2366) );
  OR2_X1 U3695 ( .A1(n3718), .A2(n3719), .ZN(n3668) );
  AND2_X1 U3696 ( .A1(n3662), .A2(n3665), .ZN(n3719) );
  AND2_X1 U3697 ( .A1(n3720), .A2(n3664), .ZN(n3718) );
  OR2_X1 U3698 ( .A1(n3721), .A2(n3722), .ZN(n3664) );
  AND2_X1 U3699 ( .A1(n3658), .A2(n3661), .ZN(n3722) );
  AND2_X1 U3700 ( .A1(n3723), .A2(n3660), .ZN(n3721) );
  OR2_X1 U3701 ( .A1(n3724), .A2(n3725), .ZN(n3660) );
  AND2_X1 U3702 ( .A1(n3654), .A2(n3657), .ZN(n3725) );
  AND2_X1 U3703 ( .A1(n3726), .A2(n3656), .ZN(n3724) );
  OR2_X1 U3704 ( .A1(n3727), .A2(n3728), .ZN(n3656) );
  AND2_X1 U3705 ( .A1(n3650), .A2(n3653), .ZN(n3728) );
  AND2_X1 U3706 ( .A1(n3729), .A2(n3652), .ZN(n3727) );
  OR2_X1 U3707 ( .A1(n3730), .A2(n3731), .ZN(n3652) );
  AND2_X1 U3708 ( .A1(n3646), .A2(n3649), .ZN(n3731) );
  AND2_X1 U3709 ( .A1(n3732), .A2(n3648), .ZN(n3730) );
  OR2_X1 U3710 ( .A1(n3733), .A2(n3734), .ZN(n3648) );
  AND2_X1 U3711 ( .A1(n3642), .A2(n3645), .ZN(n3734) );
  AND2_X1 U3712 ( .A1(n3735), .A2(n3736), .ZN(n3733) );
  OR2_X1 U3713 ( .A1(n3645), .A2(n3642), .ZN(n3736) );
  OR2_X1 U3714 ( .A1(n2218), .A2(n2591), .ZN(n3642) );
  OR3_X1 U3715 ( .A1(n2591), .A2(n2587), .A3(n2913), .ZN(n3645) );
  INV_X1 U3716 ( .A(n3644), .ZN(n3735) );
  OR2_X1 U3717 ( .A1(n3737), .A2(n3738), .ZN(n3644) );
  AND2_X1 U3718 ( .A1(b_6_), .A2(n3739), .ZN(n3738) );
  OR2_X1 U3719 ( .A1(n3740), .A2(n2918), .ZN(n3739) );
  AND2_X1 U3720 ( .A1(a_14_), .A2(n2583), .ZN(n3740) );
  AND2_X1 U3721 ( .A1(b_5_), .A2(n3741), .ZN(n3737) );
  OR2_X1 U3722 ( .A1(n3742), .A2(n2180), .ZN(n3741) );
  AND2_X1 U3723 ( .A1(a_15_), .A2(n2587), .ZN(n3742) );
  OR2_X1 U3724 ( .A1(n3649), .A2(n3646), .ZN(n3732) );
  XNOR2_X1 U3725 ( .A(n3743), .B(n3744), .ZN(n3646) );
  XOR2_X1 U3726 ( .A(n3745), .B(n3746), .Z(n3744) );
  OR2_X1 U3727 ( .A1(n2243), .A2(n2591), .ZN(n3649) );
  OR2_X1 U3728 ( .A1(n3653), .A2(n3650), .ZN(n3729) );
  XOR2_X1 U3729 ( .A(n3747), .B(n3748), .Z(n3650) );
  XOR2_X1 U3730 ( .A(n3749), .B(n3750), .Z(n3748) );
  OR2_X1 U3731 ( .A1(n2268), .A2(n2591), .ZN(n3653) );
  OR2_X1 U3732 ( .A1(n3657), .A2(n3654), .ZN(n3726) );
  XOR2_X1 U3733 ( .A(n3751), .B(n3752), .Z(n3654) );
  XOR2_X1 U3734 ( .A(n3753), .B(n3754), .Z(n3752) );
  OR2_X1 U3735 ( .A1(n2293), .A2(n2591), .ZN(n3657) );
  OR2_X1 U3736 ( .A1(n3661), .A2(n3658), .ZN(n3723) );
  XOR2_X1 U3737 ( .A(n3755), .B(n3756), .Z(n3658) );
  XOR2_X1 U3738 ( .A(n3757), .B(n3758), .Z(n3756) );
  OR2_X1 U3739 ( .A1(n2318), .A2(n2591), .ZN(n3661) );
  OR2_X1 U3740 ( .A1(n3665), .A2(n3662), .ZN(n3720) );
  XOR2_X1 U3741 ( .A(n3759), .B(n3760), .Z(n3662) );
  XOR2_X1 U3742 ( .A(n3761), .B(n3762), .Z(n3760) );
  OR2_X1 U3743 ( .A1(n2594), .A2(n2591), .ZN(n3665) );
  XOR2_X1 U3744 ( .A(n3763), .B(n3764), .Z(n3666) );
  XOR2_X1 U3745 ( .A(n3765), .B(n3766), .Z(n3764) );
  OR2_X1 U3746 ( .A1(n3672), .A2(n3669), .ZN(n3714) );
  XOR2_X1 U3747 ( .A(n3767), .B(n3768), .Z(n3669) );
  XOR2_X1 U3748 ( .A(n3769), .B(n3770), .Z(n3768) );
  OR2_X1 U3749 ( .A1(n2586), .A2(n2591), .ZN(n3672) );
  INV_X1 U3750 ( .A(b_7_), .ZN(n2591) );
  XOR2_X1 U3751 ( .A(n3771), .B(n3772), .Z(n3673) );
  XOR2_X1 U3752 ( .A(n3773), .B(n2392), .Z(n3772) );
  XOR2_X1 U3753 ( .A(n3774), .B(n3775), .Z(n3677) );
  XOR2_X1 U3754 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR2_X1 U3755 ( .A(n3778), .B(n3779), .Z(n3681) );
  XOR2_X1 U3756 ( .A(n3780), .B(n3781), .Z(n3779) );
  XOR2_X1 U3757 ( .A(n3782), .B(n3783), .Z(n3685) );
  XOR2_X1 U3758 ( .A(n3784), .B(n3785), .Z(n3783) );
  XOR2_X1 U3759 ( .A(n3786), .B(n3787), .Z(n3689) );
  XOR2_X1 U3760 ( .A(n3788), .B(n3789), .Z(n3787) );
  XOR2_X1 U3761 ( .A(n3790), .B(n3791), .Z(n2836) );
  XOR2_X1 U3762 ( .A(n3792), .B(n3793), .Z(n3791) );
  XOR2_X1 U3763 ( .A(n2811), .B(n3794), .Z(n2821) );
  XOR2_X1 U3764 ( .A(n2810), .B(n2809), .Z(n3794) );
  OR2_X1 U3765 ( .A1(n2969), .A2(n2587), .ZN(n2809) );
  OR2_X1 U3766 ( .A1(n3795), .A2(n3796), .ZN(n2810) );
  AND2_X1 U3767 ( .A1(n3793), .A2(n3792), .ZN(n3796) );
  AND2_X1 U3768 ( .A1(n3790), .A2(n3797), .ZN(n3795) );
  OR2_X1 U3769 ( .A1(n3792), .A2(n3793), .ZN(n3797) );
  OR2_X1 U3770 ( .A1(n2566), .A2(n2587), .ZN(n3793) );
  OR2_X1 U3771 ( .A1(n3798), .A2(n3799), .ZN(n3792) );
  AND2_X1 U3772 ( .A1(n3789), .A2(n3788), .ZN(n3799) );
  AND2_X1 U3773 ( .A1(n3786), .A2(n3800), .ZN(n3798) );
  OR2_X1 U3774 ( .A1(n3788), .A2(n3789), .ZN(n3800) );
  OR2_X1 U3775 ( .A1(n2570), .A2(n2587), .ZN(n3789) );
  OR2_X1 U3776 ( .A1(n3801), .A2(n3802), .ZN(n3788) );
  AND2_X1 U3777 ( .A1(n3785), .A2(n3784), .ZN(n3802) );
  AND2_X1 U3778 ( .A1(n3782), .A2(n3803), .ZN(n3801) );
  OR2_X1 U3779 ( .A1(n3784), .A2(n3785), .ZN(n3803) );
  OR2_X1 U3780 ( .A1(n2574), .A2(n2587), .ZN(n3785) );
  OR2_X1 U3781 ( .A1(n3804), .A2(n3805), .ZN(n3784) );
  AND2_X1 U3782 ( .A1(n3781), .A2(n3780), .ZN(n3805) );
  AND2_X1 U3783 ( .A1(n3778), .A2(n3806), .ZN(n3804) );
  OR2_X1 U3784 ( .A1(n3780), .A2(n3781), .ZN(n3806) );
  OR2_X1 U3785 ( .A1(n2578), .A2(n2587), .ZN(n3781) );
  OR2_X1 U3786 ( .A1(n3807), .A2(n3808), .ZN(n3780) );
  AND2_X1 U3787 ( .A1(n3777), .A2(n3776), .ZN(n3808) );
  AND2_X1 U3788 ( .A1(n3774), .A2(n3809), .ZN(n3807) );
  OR2_X1 U3789 ( .A1(n3776), .A2(n3777), .ZN(n3809) );
  OR2_X1 U3790 ( .A1(n2582), .A2(n2587), .ZN(n3777) );
  OR2_X1 U3791 ( .A1(n3810), .A2(n3811), .ZN(n3776) );
  AND2_X1 U3792 ( .A1(n2392), .A2(n3773), .ZN(n3811) );
  AND2_X1 U3793 ( .A1(n3771), .A2(n3812), .ZN(n3810) );
  OR2_X1 U3794 ( .A1(n3773), .A2(n2392), .ZN(n3812) );
  OR2_X1 U3795 ( .A1(n2586), .A2(n2587), .ZN(n2392) );
  OR2_X1 U3796 ( .A1(n3813), .A2(n3814), .ZN(n3773) );
  AND2_X1 U3797 ( .A1(n3767), .A2(n3770), .ZN(n3814) );
  AND2_X1 U3798 ( .A1(n3815), .A2(n3769), .ZN(n3813) );
  OR2_X1 U3799 ( .A1(n3816), .A2(n3817), .ZN(n3769) );
  AND2_X1 U3800 ( .A1(n3766), .A2(n3765), .ZN(n3817) );
  AND2_X1 U3801 ( .A1(n3763), .A2(n3818), .ZN(n3816) );
  OR2_X1 U3802 ( .A1(n3765), .A2(n3766), .ZN(n3818) );
  OR2_X1 U3803 ( .A1(n2594), .A2(n2587), .ZN(n3766) );
  OR2_X1 U3804 ( .A1(n3819), .A2(n3820), .ZN(n3765) );
  AND2_X1 U3805 ( .A1(n3759), .A2(n3762), .ZN(n3820) );
  AND2_X1 U3806 ( .A1(n3821), .A2(n3761), .ZN(n3819) );
  OR2_X1 U3807 ( .A1(n3822), .A2(n3823), .ZN(n3761) );
  AND2_X1 U3808 ( .A1(n3755), .A2(n3758), .ZN(n3823) );
  AND2_X1 U3809 ( .A1(n3824), .A2(n3757), .ZN(n3822) );
  OR2_X1 U3810 ( .A1(n3825), .A2(n3826), .ZN(n3757) );
  AND2_X1 U3811 ( .A1(n3751), .A2(n3754), .ZN(n3826) );
  AND2_X1 U3812 ( .A1(n3827), .A2(n3753), .ZN(n3825) );
  OR2_X1 U3813 ( .A1(n3828), .A2(n3829), .ZN(n3753) );
  AND2_X1 U3814 ( .A1(n3747), .A2(n3750), .ZN(n3829) );
  AND2_X1 U3815 ( .A1(n3830), .A2(n3749), .ZN(n3828) );
  OR2_X1 U3816 ( .A1(n3831), .A2(n3832), .ZN(n3749) );
  AND2_X1 U3817 ( .A1(n3743), .A2(n3746), .ZN(n3832) );
  AND2_X1 U3818 ( .A1(n3833), .A2(n3834), .ZN(n3831) );
  OR2_X1 U3819 ( .A1(n3746), .A2(n3743), .ZN(n3834) );
  OR2_X1 U3820 ( .A1(n2218), .A2(n2587), .ZN(n3743) );
  OR3_X1 U3821 ( .A1(n2587), .A2(n2583), .A3(n2913), .ZN(n3746) );
  INV_X1 U3822 ( .A(n3745), .ZN(n3833) );
  OR2_X1 U3823 ( .A1(n3835), .A2(n3836), .ZN(n3745) );
  AND2_X1 U3824 ( .A1(b_5_), .A2(n3837), .ZN(n3836) );
  OR2_X1 U3825 ( .A1(n3838), .A2(n2918), .ZN(n3837) );
  AND2_X1 U3826 ( .A1(a_14_), .A2(n2579), .ZN(n3838) );
  AND2_X1 U3827 ( .A1(b_4_), .A2(n3839), .ZN(n3835) );
  OR2_X1 U3828 ( .A1(n3840), .A2(n2180), .ZN(n3839) );
  AND2_X1 U3829 ( .A1(a_15_), .A2(n2583), .ZN(n3840) );
  OR2_X1 U3830 ( .A1(n3750), .A2(n3747), .ZN(n3830) );
  XNOR2_X1 U3831 ( .A(n3841), .B(n3842), .ZN(n3747) );
  XOR2_X1 U3832 ( .A(n3843), .B(n3844), .Z(n3842) );
  OR2_X1 U3833 ( .A1(n2243), .A2(n2587), .ZN(n3750) );
  OR2_X1 U3834 ( .A1(n3754), .A2(n3751), .ZN(n3827) );
  XOR2_X1 U3835 ( .A(n3845), .B(n3846), .Z(n3751) );
  XOR2_X1 U3836 ( .A(n3847), .B(n3848), .Z(n3846) );
  OR2_X1 U3837 ( .A1(n2268), .A2(n2587), .ZN(n3754) );
  OR2_X1 U3838 ( .A1(n3758), .A2(n3755), .ZN(n3824) );
  XOR2_X1 U3839 ( .A(n3849), .B(n3850), .Z(n3755) );
  XOR2_X1 U3840 ( .A(n3851), .B(n3852), .Z(n3850) );
  OR2_X1 U3841 ( .A1(n2293), .A2(n2587), .ZN(n3758) );
  OR2_X1 U3842 ( .A1(n3762), .A2(n3759), .ZN(n3821) );
  XOR2_X1 U3843 ( .A(n3853), .B(n3854), .Z(n3759) );
  XOR2_X1 U3844 ( .A(n3855), .B(n3856), .Z(n3854) );
  OR2_X1 U3845 ( .A1(n2318), .A2(n2587), .ZN(n3762) );
  XOR2_X1 U3846 ( .A(n3857), .B(n3858), .Z(n3763) );
  XOR2_X1 U3847 ( .A(n3859), .B(n3860), .Z(n3858) );
  OR2_X1 U3848 ( .A1(n3770), .A2(n3767), .ZN(n3815) );
  XOR2_X1 U3849 ( .A(n3861), .B(n3862), .Z(n3767) );
  XOR2_X1 U3850 ( .A(n3863), .B(n3864), .Z(n3862) );
  OR2_X1 U3851 ( .A1(n2590), .A2(n2587), .ZN(n3770) );
  INV_X1 U3852 ( .A(b_6_), .ZN(n2587) );
  XOR2_X1 U3853 ( .A(n3865), .B(n3866), .Z(n3771) );
  XOR2_X1 U3854 ( .A(n3867), .B(n3868), .Z(n3866) );
  XOR2_X1 U3855 ( .A(n3869), .B(n3870), .Z(n3774) );
  XOR2_X1 U3856 ( .A(n3871), .B(n3872), .Z(n3870) );
  XOR2_X1 U3857 ( .A(n3873), .B(n3874), .Z(n3778) );
  XOR2_X1 U3858 ( .A(n3875), .B(n2418), .Z(n3874) );
  XOR2_X1 U3859 ( .A(n3876), .B(n3877), .Z(n3782) );
  XOR2_X1 U3860 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR2_X1 U3861 ( .A(n3880), .B(n3881), .Z(n3786) );
  XOR2_X1 U3862 ( .A(n3882), .B(n3883), .Z(n3881) );
  XOR2_X1 U3863 ( .A(n3884), .B(n3885), .Z(n3790) );
  XOR2_X1 U3864 ( .A(n3886), .B(n3887), .Z(n3885) );
  XOR2_X1 U3865 ( .A(n3888), .B(n3889), .Z(n2811) );
  XOR2_X1 U3866 ( .A(n3890), .B(n3891), .Z(n3889) );
  INV_X1 U3867 ( .A(n3892), .ZN(n2794) );
  OR2_X1 U3868 ( .A1(n2798), .A2(n2799), .ZN(n3892) );
  OR2_X1 U3869 ( .A1(n3893), .A2(n3894), .ZN(n2799) );
  AND2_X1 U3870 ( .A1(n2816), .A2(n2815), .ZN(n3894) );
  AND2_X1 U3871 ( .A1(n2813), .A2(n3895), .ZN(n3893) );
  OR2_X1 U3872 ( .A1(n2815), .A2(n2816), .ZN(n3895) );
  OR2_X1 U3873 ( .A1(n2969), .A2(n2583), .ZN(n2816) );
  OR2_X1 U3874 ( .A1(n3896), .A2(n3897), .ZN(n2815) );
  AND2_X1 U3875 ( .A1(n3891), .A2(n3890), .ZN(n3897) );
  AND2_X1 U3876 ( .A1(n3888), .A2(n3898), .ZN(n3896) );
  OR2_X1 U3877 ( .A1(n3890), .A2(n3891), .ZN(n3898) );
  OR2_X1 U3878 ( .A1(n2566), .A2(n2583), .ZN(n3891) );
  OR2_X1 U3879 ( .A1(n3899), .A2(n3900), .ZN(n3890) );
  AND2_X1 U3880 ( .A1(n3887), .A2(n3886), .ZN(n3900) );
  AND2_X1 U3881 ( .A1(n3884), .A2(n3901), .ZN(n3899) );
  OR2_X1 U3882 ( .A1(n3886), .A2(n3887), .ZN(n3901) );
  OR2_X1 U3883 ( .A1(n2570), .A2(n2583), .ZN(n3887) );
  OR2_X1 U3884 ( .A1(n3902), .A2(n3903), .ZN(n3886) );
  AND2_X1 U3885 ( .A1(n3883), .A2(n3882), .ZN(n3903) );
  AND2_X1 U3886 ( .A1(n3880), .A2(n3904), .ZN(n3902) );
  OR2_X1 U3887 ( .A1(n3882), .A2(n3883), .ZN(n3904) );
  OR2_X1 U3888 ( .A1(n2574), .A2(n2583), .ZN(n3883) );
  OR2_X1 U3889 ( .A1(n3905), .A2(n3906), .ZN(n3882) );
  AND2_X1 U3890 ( .A1(n3879), .A2(n3878), .ZN(n3906) );
  AND2_X1 U3891 ( .A1(n3876), .A2(n3907), .ZN(n3905) );
  OR2_X1 U3892 ( .A1(n3878), .A2(n3879), .ZN(n3907) );
  OR2_X1 U3893 ( .A1(n2578), .A2(n2583), .ZN(n3879) );
  OR2_X1 U3894 ( .A1(n3908), .A2(n3909), .ZN(n3878) );
  AND2_X1 U3895 ( .A1(n2418), .A2(n3875), .ZN(n3909) );
  AND2_X1 U3896 ( .A1(n3873), .A2(n3910), .ZN(n3908) );
  OR2_X1 U3897 ( .A1(n3875), .A2(n2418), .ZN(n3910) );
  OR2_X1 U3898 ( .A1(n2582), .A2(n2583), .ZN(n2418) );
  OR2_X1 U3899 ( .A1(n3911), .A2(n3912), .ZN(n3875) );
  AND2_X1 U3900 ( .A1(n3872), .A2(n3871), .ZN(n3912) );
  AND2_X1 U3901 ( .A1(n3869), .A2(n3913), .ZN(n3911) );
  OR2_X1 U3902 ( .A1(n3871), .A2(n3872), .ZN(n3913) );
  OR2_X1 U3903 ( .A1(n2586), .A2(n2583), .ZN(n3872) );
  OR2_X1 U3904 ( .A1(n3914), .A2(n3915), .ZN(n3871) );
  AND2_X1 U3905 ( .A1(n3868), .A2(n3867), .ZN(n3915) );
  AND2_X1 U3906 ( .A1(n3865), .A2(n3916), .ZN(n3914) );
  OR2_X1 U3907 ( .A1(n3867), .A2(n3868), .ZN(n3916) );
  OR2_X1 U3908 ( .A1(n2590), .A2(n2583), .ZN(n3868) );
  OR2_X1 U3909 ( .A1(n3917), .A2(n3918), .ZN(n3867) );
  AND2_X1 U3910 ( .A1(n3861), .A2(n3864), .ZN(n3918) );
  AND2_X1 U3911 ( .A1(n3919), .A2(n3863), .ZN(n3917) );
  OR2_X1 U3912 ( .A1(n3920), .A2(n3921), .ZN(n3863) );
  AND2_X1 U3913 ( .A1(n3860), .A2(n3859), .ZN(n3921) );
  AND2_X1 U3914 ( .A1(n3857), .A2(n3922), .ZN(n3920) );
  OR2_X1 U3915 ( .A1(n3859), .A2(n3860), .ZN(n3922) );
  OR2_X1 U3916 ( .A1(n2318), .A2(n2583), .ZN(n3860) );
  OR2_X1 U3917 ( .A1(n3923), .A2(n3924), .ZN(n3859) );
  AND2_X1 U3918 ( .A1(n3853), .A2(n3856), .ZN(n3924) );
  AND2_X1 U3919 ( .A1(n3925), .A2(n3855), .ZN(n3923) );
  OR2_X1 U3920 ( .A1(n3926), .A2(n3927), .ZN(n3855) );
  AND2_X1 U3921 ( .A1(n3849), .A2(n3852), .ZN(n3927) );
  AND2_X1 U3922 ( .A1(n3928), .A2(n3851), .ZN(n3926) );
  OR2_X1 U3923 ( .A1(n3929), .A2(n3930), .ZN(n3851) );
  AND2_X1 U3924 ( .A1(n3845), .A2(n3848), .ZN(n3930) );
  AND2_X1 U3925 ( .A1(n3931), .A2(n3847), .ZN(n3929) );
  OR2_X1 U3926 ( .A1(n3932), .A2(n3933), .ZN(n3847) );
  AND2_X1 U3927 ( .A1(n3841), .A2(n3844), .ZN(n3933) );
  AND2_X1 U3928 ( .A1(n3934), .A2(n3935), .ZN(n3932) );
  OR2_X1 U3929 ( .A1(n3844), .A2(n3841), .ZN(n3935) );
  OR2_X1 U3930 ( .A1(n2218), .A2(n2583), .ZN(n3841) );
  OR3_X1 U3931 ( .A1(n2583), .A2(n2579), .A3(n2913), .ZN(n3844) );
  INV_X1 U3932 ( .A(n3843), .ZN(n3934) );
  OR2_X1 U3933 ( .A1(n3936), .A2(n3937), .ZN(n3843) );
  AND2_X1 U3934 ( .A1(b_4_), .A2(n3938), .ZN(n3937) );
  OR2_X1 U3935 ( .A1(n3939), .A2(n2918), .ZN(n3938) );
  AND2_X1 U3936 ( .A1(a_14_), .A2(n2575), .ZN(n3939) );
  AND2_X1 U3937 ( .A1(b_3_), .A2(n3940), .ZN(n3936) );
  OR2_X1 U3938 ( .A1(n3941), .A2(n2180), .ZN(n3940) );
  AND2_X1 U3939 ( .A1(a_15_), .A2(n2579), .ZN(n3941) );
  OR2_X1 U3940 ( .A1(n3848), .A2(n3845), .ZN(n3931) );
  XNOR2_X1 U3941 ( .A(n3942), .B(n3943), .ZN(n3845) );
  XOR2_X1 U3942 ( .A(n3944), .B(n3945), .Z(n3943) );
  OR2_X1 U3943 ( .A1(n2243), .A2(n2583), .ZN(n3848) );
  OR2_X1 U3944 ( .A1(n3852), .A2(n3849), .ZN(n3928) );
  XOR2_X1 U3945 ( .A(n3946), .B(n3947), .Z(n3849) );
  XOR2_X1 U3946 ( .A(n3948), .B(n3949), .Z(n3947) );
  OR2_X1 U3947 ( .A1(n2268), .A2(n2583), .ZN(n3852) );
  OR2_X1 U3948 ( .A1(n3856), .A2(n3853), .ZN(n3925) );
  XOR2_X1 U3949 ( .A(n3950), .B(n3951), .Z(n3853) );
  XOR2_X1 U3950 ( .A(n3952), .B(n3953), .Z(n3951) );
  OR2_X1 U3951 ( .A1(n2293), .A2(n2583), .ZN(n3856) );
  XOR2_X1 U3952 ( .A(n3954), .B(n3955), .Z(n3857) );
  XOR2_X1 U3953 ( .A(n3956), .B(n3957), .Z(n3955) );
  OR2_X1 U3954 ( .A1(n3864), .A2(n3861), .ZN(n3919) );
  XOR2_X1 U3955 ( .A(n3958), .B(n3959), .Z(n3861) );
  XOR2_X1 U3956 ( .A(n3960), .B(n3961), .Z(n3959) );
  OR2_X1 U3957 ( .A1(n2594), .A2(n2583), .ZN(n3864) );
  INV_X1 U3958 ( .A(b_5_), .ZN(n2583) );
  XOR2_X1 U3959 ( .A(n3962), .B(n3963), .Z(n3865) );
  XOR2_X1 U3960 ( .A(n3964), .B(n3965), .Z(n3963) );
  XOR2_X1 U3961 ( .A(n3966), .B(n3967), .Z(n3869) );
  XOR2_X1 U3962 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR2_X1 U3963 ( .A(n3970), .B(n3971), .Z(n3873) );
  XOR2_X1 U3964 ( .A(n3972), .B(n3973), .Z(n3971) );
  XOR2_X1 U3965 ( .A(n3974), .B(n3975), .Z(n3876) );
  XOR2_X1 U3966 ( .A(n3976), .B(n3977), .Z(n3975) );
  XOR2_X1 U3967 ( .A(n3978), .B(n3979), .Z(n3880) );
  XOR2_X1 U3968 ( .A(n3980), .B(n2444), .Z(n3979) );
  XOR2_X1 U3969 ( .A(n3981), .B(n3982), .Z(n3884) );
  XOR2_X1 U3970 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR2_X1 U3971 ( .A(n3985), .B(n3986), .Z(n3888) );
  XOR2_X1 U3972 ( .A(n3987), .B(n3988), .Z(n3986) );
  XOR2_X1 U3973 ( .A(n3989), .B(n3990), .Z(n2813) );
  XOR2_X1 U3974 ( .A(n3991), .B(n3992), .Z(n3990) );
  XOR2_X1 U3975 ( .A(n2788), .B(n3993), .Z(n2798) );
  XOR2_X1 U3976 ( .A(n2787), .B(n2786), .Z(n3993) );
  OR2_X1 U3977 ( .A1(n2969), .A2(n2579), .ZN(n2786) );
  OR2_X1 U3978 ( .A1(n3994), .A2(n3995), .ZN(n2787) );
  AND2_X1 U3979 ( .A1(n3992), .A2(n3991), .ZN(n3995) );
  AND2_X1 U3980 ( .A1(n3989), .A2(n3996), .ZN(n3994) );
  OR2_X1 U3981 ( .A1(n3991), .A2(n3992), .ZN(n3996) );
  OR2_X1 U3982 ( .A1(n2566), .A2(n2579), .ZN(n3992) );
  OR2_X1 U3983 ( .A1(n3997), .A2(n3998), .ZN(n3991) );
  AND2_X1 U3984 ( .A1(n3988), .A2(n3987), .ZN(n3998) );
  AND2_X1 U3985 ( .A1(n3985), .A2(n3999), .ZN(n3997) );
  OR2_X1 U3986 ( .A1(n3987), .A2(n3988), .ZN(n3999) );
  OR2_X1 U3987 ( .A1(n2570), .A2(n2579), .ZN(n3988) );
  OR2_X1 U3988 ( .A1(n4000), .A2(n4001), .ZN(n3987) );
  AND2_X1 U3989 ( .A1(n3984), .A2(n3983), .ZN(n4001) );
  AND2_X1 U3990 ( .A1(n3981), .A2(n4002), .ZN(n4000) );
  OR2_X1 U3991 ( .A1(n3983), .A2(n3984), .ZN(n4002) );
  OR2_X1 U3992 ( .A1(n2574), .A2(n2579), .ZN(n3984) );
  OR2_X1 U3993 ( .A1(n4003), .A2(n4004), .ZN(n3983) );
  AND2_X1 U3994 ( .A1(n2444), .A2(n3980), .ZN(n4004) );
  AND2_X1 U3995 ( .A1(n3978), .A2(n4005), .ZN(n4003) );
  OR2_X1 U3996 ( .A1(n3980), .A2(n2444), .ZN(n4005) );
  OR2_X1 U3997 ( .A1(n2578), .A2(n2579), .ZN(n2444) );
  OR2_X1 U3998 ( .A1(n4006), .A2(n4007), .ZN(n3980) );
  AND2_X1 U3999 ( .A1(n3977), .A2(n3976), .ZN(n4007) );
  AND2_X1 U4000 ( .A1(n3974), .A2(n4008), .ZN(n4006) );
  OR2_X1 U4001 ( .A1(n3976), .A2(n3977), .ZN(n4008) );
  OR2_X1 U4002 ( .A1(n2582), .A2(n2579), .ZN(n3977) );
  OR2_X1 U4003 ( .A1(n4009), .A2(n4010), .ZN(n3976) );
  AND2_X1 U4004 ( .A1(n3973), .A2(n3972), .ZN(n4010) );
  AND2_X1 U4005 ( .A1(n3970), .A2(n4011), .ZN(n4009) );
  OR2_X1 U4006 ( .A1(n3972), .A2(n3973), .ZN(n4011) );
  OR2_X1 U4007 ( .A1(n2586), .A2(n2579), .ZN(n3973) );
  OR2_X1 U4008 ( .A1(n4012), .A2(n4013), .ZN(n3972) );
  AND2_X1 U4009 ( .A1(n3969), .A2(n3968), .ZN(n4013) );
  AND2_X1 U4010 ( .A1(n3966), .A2(n4014), .ZN(n4012) );
  OR2_X1 U4011 ( .A1(n3968), .A2(n3969), .ZN(n4014) );
  OR2_X1 U4012 ( .A1(n2590), .A2(n2579), .ZN(n3969) );
  OR2_X1 U4013 ( .A1(n4015), .A2(n4016), .ZN(n3968) );
  AND2_X1 U4014 ( .A1(n3965), .A2(n3964), .ZN(n4016) );
  AND2_X1 U4015 ( .A1(n3962), .A2(n4017), .ZN(n4015) );
  OR2_X1 U4016 ( .A1(n3964), .A2(n3965), .ZN(n4017) );
  OR2_X1 U4017 ( .A1(n2594), .A2(n2579), .ZN(n3965) );
  OR2_X1 U4018 ( .A1(n4018), .A2(n4019), .ZN(n3964) );
  AND2_X1 U4019 ( .A1(n3958), .A2(n3961), .ZN(n4019) );
  AND2_X1 U4020 ( .A1(n4020), .A2(n3960), .ZN(n4018) );
  OR2_X1 U4021 ( .A1(n4021), .A2(n4022), .ZN(n3960) );
  AND2_X1 U4022 ( .A1(n3957), .A2(n3956), .ZN(n4022) );
  AND2_X1 U4023 ( .A1(n3954), .A2(n4023), .ZN(n4021) );
  OR2_X1 U4024 ( .A1(n3956), .A2(n3957), .ZN(n4023) );
  OR2_X1 U4025 ( .A1(n2293), .A2(n2579), .ZN(n3957) );
  OR2_X1 U4026 ( .A1(n4024), .A2(n4025), .ZN(n3956) );
  AND2_X1 U4027 ( .A1(n3950), .A2(n3953), .ZN(n4025) );
  AND2_X1 U4028 ( .A1(n4026), .A2(n3952), .ZN(n4024) );
  OR2_X1 U4029 ( .A1(n4027), .A2(n4028), .ZN(n3952) );
  AND2_X1 U4030 ( .A1(n3946), .A2(n3949), .ZN(n4028) );
  AND2_X1 U4031 ( .A1(n4029), .A2(n3948), .ZN(n4027) );
  OR2_X1 U4032 ( .A1(n4030), .A2(n4031), .ZN(n3948) );
  AND2_X1 U4033 ( .A1(n3942), .A2(n3945), .ZN(n4031) );
  AND2_X1 U4034 ( .A1(n4032), .A2(n4033), .ZN(n4030) );
  OR2_X1 U4035 ( .A1(n3945), .A2(n3942), .ZN(n4033) );
  OR2_X1 U4036 ( .A1(n2218), .A2(n2579), .ZN(n3942) );
  OR3_X1 U4037 ( .A1(n2579), .A2(n2575), .A3(n2913), .ZN(n3945) );
  INV_X1 U4038 ( .A(n3944), .ZN(n4032) );
  OR2_X1 U4039 ( .A1(n4034), .A2(n4035), .ZN(n3944) );
  AND2_X1 U4040 ( .A1(b_3_), .A2(n4036), .ZN(n4035) );
  OR2_X1 U4041 ( .A1(n4037), .A2(n2918), .ZN(n4036) );
  AND2_X1 U4042 ( .A1(a_14_), .A2(n2571), .ZN(n4037) );
  AND2_X1 U4043 ( .A1(b_2_), .A2(n4038), .ZN(n4034) );
  OR2_X1 U4044 ( .A1(n4039), .A2(n2180), .ZN(n4038) );
  AND2_X1 U4045 ( .A1(a_15_), .A2(n2575), .ZN(n4039) );
  OR2_X1 U4046 ( .A1(n3949), .A2(n3946), .ZN(n4029) );
  XNOR2_X1 U4047 ( .A(n4040), .B(n4041), .ZN(n3946) );
  XOR2_X1 U4048 ( .A(n4042), .B(n4043), .Z(n4041) );
  OR2_X1 U4049 ( .A1(n2243), .A2(n2579), .ZN(n3949) );
  OR2_X1 U4050 ( .A1(n3953), .A2(n3950), .ZN(n4026) );
  XOR2_X1 U4051 ( .A(n4044), .B(n4045), .Z(n3950) );
  XOR2_X1 U4052 ( .A(n4046), .B(n4047), .Z(n4045) );
  OR2_X1 U4053 ( .A1(n2268), .A2(n2579), .ZN(n3953) );
  XOR2_X1 U4054 ( .A(n4048), .B(n4049), .Z(n3954) );
  XOR2_X1 U4055 ( .A(n4050), .B(n4051), .Z(n4049) );
  OR2_X1 U4056 ( .A1(n3961), .A2(n3958), .ZN(n4020) );
  XOR2_X1 U4057 ( .A(n4052), .B(n4053), .Z(n3958) );
  XOR2_X1 U4058 ( .A(n4054), .B(n4055), .Z(n4053) );
  OR2_X1 U4059 ( .A1(n2318), .A2(n2579), .ZN(n3961) );
  INV_X1 U4060 ( .A(b_4_), .ZN(n2579) );
  XOR2_X1 U4061 ( .A(n4056), .B(n4057), .Z(n3962) );
  XOR2_X1 U4062 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR2_X1 U4063 ( .A(n4060), .B(n4061), .Z(n3966) );
  XOR2_X1 U4064 ( .A(n4062), .B(n4063), .Z(n4061) );
  XOR2_X1 U4065 ( .A(n4064), .B(n4065), .Z(n3970) );
  XOR2_X1 U4066 ( .A(n4066), .B(n4067), .Z(n4065) );
  XOR2_X1 U4067 ( .A(n4068), .B(n4069), .Z(n3974) );
  XOR2_X1 U4068 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR2_X1 U4069 ( .A(n4072), .B(n4073), .Z(n3978) );
  XOR2_X1 U4070 ( .A(n4074), .B(n4075), .Z(n4073) );
  XOR2_X1 U4071 ( .A(n4076), .B(n4077), .Z(n3981) );
  XOR2_X1 U4072 ( .A(n4078), .B(n4079), .Z(n4077) );
  XOR2_X1 U4073 ( .A(n4080), .B(n4081), .Z(n3985) );
  XOR2_X1 U4074 ( .A(n4082), .B(n2481), .Z(n4081) );
  XOR2_X1 U4075 ( .A(n4083), .B(n4084), .Z(n3989) );
  XOR2_X1 U4076 ( .A(n4085), .B(n4086), .Z(n4084) );
  XOR2_X1 U4077 ( .A(n4087), .B(n4088), .Z(n2788) );
  XOR2_X1 U4078 ( .A(n4089), .B(n4090), .Z(n4088) );
  INV_X1 U4079 ( .A(n4091), .ZN(n2771) );
  OR2_X1 U4080 ( .A1(n2775), .A2(n2776), .ZN(n4091) );
  OR2_X1 U4081 ( .A1(n4092), .A2(n4093), .ZN(n2776) );
  AND2_X1 U4082 ( .A1(n2793), .A2(n2792), .ZN(n4093) );
  AND2_X1 U4083 ( .A1(n2790), .A2(n4094), .ZN(n4092) );
  OR2_X1 U4084 ( .A1(n2792), .A2(n2793), .ZN(n4094) );
  OR2_X1 U4085 ( .A1(n2969), .A2(n2575), .ZN(n2793) );
  OR2_X1 U4086 ( .A1(n4095), .A2(n4096), .ZN(n2792) );
  AND2_X1 U4087 ( .A1(n4090), .A2(n4089), .ZN(n4096) );
  AND2_X1 U4088 ( .A1(n4087), .A2(n4097), .ZN(n4095) );
  OR2_X1 U4089 ( .A1(n4089), .A2(n4090), .ZN(n4097) );
  OR2_X1 U4090 ( .A1(n2566), .A2(n2575), .ZN(n4090) );
  OR2_X1 U4091 ( .A1(n4098), .A2(n4099), .ZN(n4089) );
  AND2_X1 U4092 ( .A1(n4086), .A2(n4085), .ZN(n4099) );
  AND2_X1 U4093 ( .A1(n4083), .A2(n4100), .ZN(n4098) );
  OR2_X1 U4094 ( .A1(n4085), .A2(n4086), .ZN(n4100) );
  OR2_X1 U4095 ( .A1(n2570), .A2(n2575), .ZN(n4086) );
  OR2_X1 U4096 ( .A1(n4101), .A2(n4102), .ZN(n4085) );
  AND2_X1 U4097 ( .A1(n2481), .A2(n4082), .ZN(n4102) );
  AND2_X1 U4098 ( .A1(n4080), .A2(n4103), .ZN(n4101) );
  OR2_X1 U4099 ( .A1(n4082), .A2(n2481), .ZN(n4103) );
  OR2_X1 U4100 ( .A1(n2574), .A2(n2575), .ZN(n2481) );
  OR2_X1 U4101 ( .A1(n4104), .A2(n4105), .ZN(n4082) );
  AND2_X1 U4102 ( .A1(n4079), .A2(n4078), .ZN(n4105) );
  AND2_X1 U4103 ( .A1(n4076), .A2(n4106), .ZN(n4104) );
  OR2_X1 U4104 ( .A1(n4078), .A2(n4079), .ZN(n4106) );
  OR2_X1 U4105 ( .A1(n2578), .A2(n2575), .ZN(n4079) );
  OR2_X1 U4106 ( .A1(n4107), .A2(n4108), .ZN(n4078) );
  AND2_X1 U4107 ( .A1(n4075), .A2(n4074), .ZN(n4108) );
  AND2_X1 U4108 ( .A1(n4072), .A2(n4109), .ZN(n4107) );
  OR2_X1 U4109 ( .A1(n4074), .A2(n4075), .ZN(n4109) );
  OR2_X1 U4110 ( .A1(n2582), .A2(n2575), .ZN(n4075) );
  OR2_X1 U4111 ( .A1(n4110), .A2(n4111), .ZN(n4074) );
  AND2_X1 U4112 ( .A1(n4071), .A2(n4070), .ZN(n4111) );
  AND2_X1 U4113 ( .A1(n4068), .A2(n4112), .ZN(n4110) );
  OR2_X1 U4114 ( .A1(n4070), .A2(n4071), .ZN(n4112) );
  OR2_X1 U4115 ( .A1(n2586), .A2(n2575), .ZN(n4071) );
  OR2_X1 U4116 ( .A1(n4113), .A2(n4114), .ZN(n4070) );
  AND2_X1 U4117 ( .A1(n4067), .A2(n4066), .ZN(n4114) );
  AND2_X1 U4118 ( .A1(n4064), .A2(n4115), .ZN(n4113) );
  OR2_X1 U4119 ( .A1(n4066), .A2(n4067), .ZN(n4115) );
  OR2_X1 U4120 ( .A1(n2590), .A2(n2575), .ZN(n4067) );
  OR2_X1 U4121 ( .A1(n4116), .A2(n4117), .ZN(n4066) );
  AND2_X1 U4122 ( .A1(n4063), .A2(n4062), .ZN(n4117) );
  AND2_X1 U4123 ( .A1(n4060), .A2(n4118), .ZN(n4116) );
  OR2_X1 U4124 ( .A1(n4062), .A2(n4063), .ZN(n4118) );
  OR2_X1 U4125 ( .A1(n2594), .A2(n2575), .ZN(n4063) );
  OR2_X1 U4126 ( .A1(n4119), .A2(n4120), .ZN(n4062) );
  AND2_X1 U4127 ( .A1(n4059), .A2(n4058), .ZN(n4120) );
  AND2_X1 U4128 ( .A1(n4056), .A2(n4121), .ZN(n4119) );
  OR2_X1 U4129 ( .A1(n4058), .A2(n4059), .ZN(n4121) );
  OR2_X1 U4130 ( .A1(n2318), .A2(n2575), .ZN(n4059) );
  OR2_X1 U4131 ( .A1(n4122), .A2(n4123), .ZN(n4058) );
  AND2_X1 U4132 ( .A1(n4052), .A2(n4055), .ZN(n4123) );
  AND2_X1 U4133 ( .A1(n4124), .A2(n4054), .ZN(n4122) );
  OR2_X1 U4134 ( .A1(n4125), .A2(n4126), .ZN(n4054) );
  AND2_X1 U4135 ( .A1(n4051), .A2(n4050), .ZN(n4126) );
  AND2_X1 U4136 ( .A1(n4048), .A2(n4127), .ZN(n4125) );
  OR2_X1 U4137 ( .A1(n4050), .A2(n4051), .ZN(n4127) );
  OR2_X1 U4138 ( .A1(n2268), .A2(n2575), .ZN(n4051) );
  OR2_X1 U4139 ( .A1(n4128), .A2(n4129), .ZN(n4050) );
  AND2_X1 U4140 ( .A1(n4044), .A2(n4047), .ZN(n4129) );
  AND2_X1 U4141 ( .A1(n4130), .A2(n4046), .ZN(n4128) );
  OR2_X1 U4142 ( .A1(n4131), .A2(n4132), .ZN(n4046) );
  AND2_X1 U4143 ( .A1(n4040), .A2(n4043), .ZN(n4132) );
  AND2_X1 U4144 ( .A1(n4133), .A2(n4134), .ZN(n4131) );
  OR2_X1 U4145 ( .A1(n4043), .A2(n4040), .ZN(n4134) );
  OR2_X1 U4146 ( .A1(n2218), .A2(n2575), .ZN(n4040) );
  OR3_X1 U4147 ( .A1(n2575), .A2(n2571), .A3(n2913), .ZN(n4043) );
  INV_X1 U4148 ( .A(n4042), .ZN(n4133) );
  OR2_X1 U4149 ( .A1(n4135), .A2(n4136), .ZN(n4042) );
  AND2_X1 U4150 ( .A1(b_2_), .A2(n4137), .ZN(n4136) );
  OR2_X1 U4151 ( .A1(n4138), .A2(n2918), .ZN(n4137) );
  AND2_X1 U4152 ( .A1(a_14_), .A2(n2567), .ZN(n4138) );
  AND2_X1 U4153 ( .A1(b_1_), .A2(n4139), .ZN(n4135) );
  OR2_X1 U4154 ( .A1(n4140), .A2(n2180), .ZN(n4139) );
  AND2_X1 U4155 ( .A1(a_15_), .A2(n2571), .ZN(n4140) );
  OR2_X1 U4156 ( .A1(n4047), .A2(n4044), .ZN(n4130) );
  XNOR2_X1 U4157 ( .A(n4141), .B(n4142), .ZN(n4044) );
  XOR2_X1 U4158 ( .A(n4143), .B(n4144), .Z(n4142) );
  OR2_X1 U4159 ( .A1(n2243), .A2(n2575), .ZN(n4047) );
  XOR2_X1 U4160 ( .A(n4145), .B(n4146), .Z(n4048) );
  XOR2_X1 U4161 ( .A(n4147), .B(n4148), .Z(n4146) );
  OR2_X1 U4162 ( .A1(n4055), .A2(n4052), .ZN(n4124) );
  XOR2_X1 U4163 ( .A(n4149), .B(n4150), .Z(n4052) );
  XOR2_X1 U4164 ( .A(n4151), .B(n4152), .Z(n4150) );
  OR2_X1 U4165 ( .A1(n2293), .A2(n2575), .ZN(n4055) );
  INV_X1 U4166 ( .A(b_3_), .ZN(n2575) );
  XOR2_X1 U4167 ( .A(n4153), .B(n4154), .Z(n4056) );
  XOR2_X1 U4168 ( .A(n4155), .B(n4156), .Z(n4154) );
  XOR2_X1 U4169 ( .A(n4157), .B(n4158), .Z(n4060) );
  XOR2_X1 U4170 ( .A(n4159), .B(n4160), .Z(n4158) );
  XOR2_X1 U4171 ( .A(n4161), .B(n4162), .Z(n4064) );
  XOR2_X1 U4172 ( .A(n4163), .B(n4164), .Z(n4162) );
  XOR2_X1 U4173 ( .A(n4165), .B(n4166), .Z(n4068) );
  XOR2_X1 U4174 ( .A(n4167), .B(n4168), .Z(n4166) );
  XOR2_X1 U4175 ( .A(n4169), .B(n4170), .Z(n4072) );
  XOR2_X1 U4176 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR2_X1 U4177 ( .A(n4173), .B(n4174), .Z(n4076) );
  XOR2_X1 U4178 ( .A(n4175), .B(n4176), .Z(n4174) );
  XOR2_X1 U4179 ( .A(n4177), .B(n4178), .Z(n4080) );
  XOR2_X1 U4180 ( .A(n4179), .B(n4180), .Z(n4178) );
  XOR2_X1 U4181 ( .A(n4181), .B(n4182), .Z(n4083) );
  XOR2_X1 U4182 ( .A(n4183), .B(n4184), .Z(n4182) );
  XOR2_X1 U4183 ( .A(n4185), .B(n4186), .Z(n4087) );
  XOR2_X1 U4184 ( .A(n4187), .B(n2507), .Z(n4186) );
  XOR2_X1 U4185 ( .A(n4188), .B(n4189), .Z(n2790) );
  XOR2_X1 U4186 ( .A(n4190), .B(n4191), .Z(n4189) );
  XOR2_X1 U4187 ( .A(n4192), .B(n4193), .Z(n2775) );
  XOR2_X1 U4188 ( .A(n4194), .B(n4195), .Z(n4193) );
  AND3_X1 U4189 ( .A1(n2458), .A2(n2456), .A3(n2457), .ZN(n2459) );
  INV_X1 U4190 ( .A(n4196), .ZN(n2457) );
  OR2_X1 U4191 ( .A1(n4197), .A2(n4198), .ZN(n4196) );
  AND2_X1 U4192 ( .A1(n4195), .A2(n4194), .ZN(n4198) );
  AND2_X1 U4193 ( .A1(n4192), .A2(n4199), .ZN(n4197) );
  OR2_X1 U4194 ( .A1(n4194), .A2(n4195), .ZN(n4199) );
  OR2_X1 U4195 ( .A1(n2969), .A2(n2571), .ZN(n4195) );
  OR2_X1 U4196 ( .A1(n4200), .A2(n4201), .ZN(n4194) );
  AND2_X1 U4197 ( .A1(n4191), .A2(n4190), .ZN(n4201) );
  AND2_X1 U4198 ( .A1(n4188), .A2(n4202), .ZN(n4200) );
  OR2_X1 U4199 ( .A1(n4190), .A2(n4191), .ZN(n4202) );
  OR2_X1 U4200 ( .A1(n2566), .A2(n2571), .ZN(n4191) );
  OR2_X1 U4201 ( .A1(n4203), .A2(n4204), .ZN(n4190) );
  AND2_X1 U4202 ( .A1(n2507), .A2(n4187), .ZN(n4204) );
  AND2_X1 U4203 ( .A1(n4185), .A2(n4205), .ZN(n4203) );
  OR2_X1 U4204 ( .A1(n4187), .A2(n2507), .ZN(n4205) );
  OR2_X1 U4205 ( .A1(n2570), .A2(n2571), .ZN(n2507) );
  OR2_X1 U4206 ( .A1(n4206), .A2(n4207), .ZN(n4187) );
  AND2_X1 U4207 ( .A1(n4184), .A2(n4183), .ZN(n4207) );
  AND2_X1 U4208 ( .A1(n4181), .A2(n4208), .ZN(n4206) );
  OR2_X1 U4209 ( .A1(n4183), .A2(n4184), .ZN(n4208) );
  OR2_X1 U4210 ( .A1(n2574), .A2(n2571), .ZN(n4184) );
  OR2_X1 U4211 ( .A1(n4209), .A2(n4210), .ZN(n4183) );
  AND2_X1 U4212 ( .A1(n4180), .A2(n4179), .ZN(n4210) );
  AND2_X1 U4213 ( .A1(n4177), .A2(n4211), .ZN(n4209) );
  OR2_X1 U4214 ( .A1(n4179), .A2(n4180), .ZN(n4211) );
  OR2_X1 U4215 ( .A1(n2578), .A2(n2571), .ZN(n4180) );
  OR2_X1 U4216 ( .A1(n4212), .A2(n4213), .ZN(n4179) );
  AND2_X1 U4217 ( .A1(n4176), .A2(n4175), .ZN(n4213) );
  AND2_X1 U4218 ( .A1(n4173), .A2(n4214), .ZN(n4212) );
  OR2_X1 U4219 ( .A1(n4175), .A2(n4176), .ZN(n4214) );
  OR2_X1 U4220 ( .A1(n2582), .A2(n2571), .ZN(n4176) );
  OR2_X1 U4221 ( .A1(n4215), .A2(n4216), .ZN(n4175) );
  AND2_X1 U4222 ( .A1(n4172), .A2(n4171), .ZN(n4216) );
  AND2_X1 U4223 ( .A1(n4169), .A2(n4217), .ZN(n4215) );
  OR2_X1 U4224 ( .A1(n4171), .A2(n4172), .ZN(n4217) );
  OR2_X1 U4225 ( .A1(n2586), .A2(n2571), .ZN(n4172) );
  OR2_X1 U4226 ( .A1(n4218), .A2(n4219), .ZN(n4171) );
  AND2_X1 U4227 ( .A1(n4168), .A2(n4167), .ZN(n4219) );
  AND2_X1 U4228 ( .A1(n4165), .A2(n4220), .ZN(n4218) );
  OR2_X1 U4229 ( .A1(n4167), .A2(n4168), .ZN(n4220) );
  OR2_X1 U4230 ( .A1(n2590), .A2(n2571), .ZN(n4168) );
  OR2_X1 U4231 ( .A1(n4221), .A2(n4222), .ZN(n4167) );
  AND2_X1 U4232 ( .A1(n4164), .A2(n4163), .ZN(n4222) );
  AND2_X1 U4233 ( .A1(n4161), .A2(n4223), .ZN(n4221) );
  OR2_X1 U4234 ( .A1(n4163), .A2(n4164), .ZN(n4223) );
  OR2_X1 U4235 ( .A1(n2594), .A2(n2571), .ZN(n4164) );
  OR2_X1 U4236 ( .A1(n4224), .A2(n4225), .ZN(n4163) );
  AND2_X1 U4237 ( .A1(n4160), .A2(n4159), .ZN(n4225) );
  AND2_X1 U4238 ( .A1(n4157), .A2(n4226), .ZN(n4224) );
  OR2_X1 U4239 ( .A1(n4159), .A2(n4160), .ZN(n4226) );
  OR2_X1 U4240 ( .A1(n2318), .A2(n2571), .ZN(n4160) );
  OR2_X1 U4241 ( .A1(n4227), .A2(n4228), .ZN(n4159) );
  AND2_X1 U4242 ( .A1(n4156), .A2(n4155), .ZN(n4228) );
  AND2_X1 U4243 ( .A1(n4153), .A2(n4229), .ZN(n4227) );
  OR2_X1 U4244 ( .A1(n4155), .A2(n4156), .ZN(n4229) );
  OR2_X1 U4245 ( .A1(n2293), .A2(n2571), .ZN(n4156) );
  OR2_X1 U4246 ( .A1(n4230), .A2(n4231), .ZN(n4155) );
  AND2_X1 U4247 ( .A1(n4149), .A2(n4152), .ZN(n4231) );
  AND2_X1 U4248 ( .A1(n4232), .A2(n4151), .ZN(n4230) );
  OR2_X1 U4249 ( .A1(n4233), .A2(n4234), .ZN(n4151) );
  AND2_X1 U4250 ( .A1(n4148), .A2(n4147), .ZN(n4234) );
  AND2_X1 U4251 ( .A1(n4145), .A2(n4235), .ZN(n4233) );
  OR2_X1 U4252 ( .A1(n4147), .A2(n4148), .ZN(n4235) );
  OR2_X1 U4253 ( .A1(n2243), .A2(n2571), .ZN(n4148) );
  OR2_X1 U4254 ( .A1(n4236), .A2(n4237), .ZN(n4147) );
  AND2_X1 U4255 ( .A1(n4141), .A2(n4144), .ZN(n4237) );
  AND2_X1 U4256 ( .A1(n4238), .A2(n4239), .ZN(n4236) );
  OR2_X1 U4257 ( .A1(n4144), .A2(n4141), .ZN(n4239) );
  OR2_X1 U4258 ( .A1(n2218), .A2(n2571), .ZN(n4141) );
  OR3_X1 U4259 ( .A1(n2571), .A2(n2567), .A3(n2913), .ZN(n4144) );
  INV_X1 U4260 ( .A(n4143), .ZN(n4238) );
  OR2_X1 U4261 ( .A1(n4240), .A2(n4241), .ZN(n4143) );
  AND2_X1 U4262 ( .A1(b_1_), .A2(n4242), .ZN(n4241) );
  OR2_X1 U4263 ( .A1(n4243), .A2(n2918), .ZN(n4242) );
  AND2_X1 U4264 ( .A1(n2619), .A2(a_14_), .ZN(n2918) );
  AND2_X1 U4265 ( .A1(a_14_), .A2(n2723), .ZN(n4243) );
  AND2_X1 U4266 ( .A1(b_0_), .A2(n4244), .ZN(n4240) );
  OR2_X1 U4267 ( .A1(n4245), .A2(n2180), .ZN(n4244) );
  AND2_X1 U4268 ( .A1(n2174), .A2(a_15_), .ZN(n2180) );
  AND2_X1 U4269 ( .A1(a_15_), .A2(n2567), .ZN(n4245) );
  XNOR2_X1 U4270 ( .A(n4246), .B(n4247), .ZN(n4145) );
  OR2_X1 U4271 ( .A1(n4248), .A2(n4249), .ZN(n4246) );
  INV_X1 U4272 ( .A(n4250), .ZN(n4249) );
  AND2_X1 U4273 ( .A1(n4251), .A2(n4252), .ZN(n4248) );
  OR2_X1 U4274 ( .A1(n2723), .A2(n2174), .ZN(n4251) );
  OR2_X1 U4275 ( .A1(n4152), .A2(n4149), .ZN(n4232) );
  XOR2_X1 U4276 ( .A(n4253), .B(n4254), .Z(n4149) );
  XOR2_X1 U4277 ( .A(n4255), .B(n4256), .Z(n4253) );
  OR2_X1 U4278 ( .A1(n2268), .A2(n2571), .ZN(n4152) );
  INV_X1 U4279 ( .A(b_2_), .ZN(n2571) );
  XNOR2_X1 U4280 ( .A(n4257), .B(n4258), .ZN(n4153) );
  XNOR2_X1 U4281 ( .A(n4259), .B(n4260), .ZN(n4257) );
  XNOR2_X1 U4282 ( .A(n4261), .B(n4262), .ZN(n4157) );
  XNOR2_X1 U4283 ( .A(n4263), .B(n4264), .ZN(n4261) );
  XNOR2_X1 U4284 ( .A(n4265), .B(n4266), .ZN(n4161) );
  XNOR2_X1 U4285 ( .A(n4267), .B(n4268), .ZN(n4265) );
  XOR2_X1 U4286 ( .A(n4269), .B(n4270), .Z(n4165) );
  XOR2_X1 U4287 ( .A(n4271), .B(n4272), .Z(n4270) );
  XOR2_X1 U4288 ( .A(n4273), .B(n4274), .Z(n4169) );
  XOR2_X1 U4289 ( .A(n4275), .B(n4276), .Z(n4274) );
  XOR2_X1 U4290 ( .A(n4277), .B(n4278), .Z(n4173) );
  XOR2_X1 U4291 ( .A(n4279), .B(n4280), .Z(n4278) );
  XOR2_X1 U4292 ( .A(n4281), .B(n4282), .Z(n4177) );
  XOR2_X1 U4293 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR2_X1 U4294 ( .A(n4285), .B(n4286), .Z(n4181) );
  XOR2_X1 U4295 ( .A(n4287), .B(n4288), .Z(n4286) );
  XOR2_X1 U4296 ( .A(n4289), .B(n4290), .Z(n4185) );
  XOR2_X1 U4297 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR2_X1 U4298 ( .A(n4293), .B(n4294), .Z(n4188) );
  XOR2_X1 U4299 ( .A(n4295), .B(n4296), .Z(n4294) );
  XOR2_X1 U4300 ( .A(n4297), .B(n4298), .Z(n4192) );
  XOR2_X1 U4301 ( .A(n4299), .B(n2533), .Z(n4298) );
  XOR2_X1 U4302 ( .A(n4300), .B(n2770), .Z(n2456) );
  OR2_X1 U4303 ( .A1(n4301), .A2(n4302), .ZN(n2770) );
  AND2_X1 U4304 ( .A1(n4303), .A2(n4304), .ZN(n4302) );
  AND2_X1 U4305 ( .A1(n4305), .A2(n4306), .ZN(n4301) );
  OR2_X1 U4306 ( .A1(n4304), .A2(n4303), .ZN(n4305) );
  OR2_X1 U4307 ( .A1(n2723), .A2(n2969), .ZN(n4300) );
  XNOR2_X1 U4308 ( .A(n4303), .B(n4307), .ZN(n2458) );
  XOR2_X1 U4309 ( .A(n4304), .B(n4306), .Z(n4307) );
  OR2_X1 U4310 ( .A1(n2969), .A2(n2567), .ZN(n4306) );
  INV_X1 U4311 ( .A(a_0_), .ZN(n2969) );
  OR2_X1 U4312 ( .A1(n4308), .A2(n4309), .ZN(n4304) );
  AND2_X1 U4313 ( .A1(n4297), .A2(n4299), .ZN(n4309) );
  AND2_X1 U4314 ( .A1(n4310), .A2(n2533), .ZN(n4308) );
  OR2_X1 U4315 ( .A1(n2566), .A2(n2567), .ZN(n2533) );
  OR2_X1 U4316 ( .A1(n4299), .A2(n4297), .ZN(n4310) );
  OR2_X1 U4317 ( .A1(n2723), .A2(n2570), .ZN(n4297) );
  OR2_X1 U4318 ( .A1(n4311), .A2(n4312), .ZN(n4299) );
  AND2_X1 U4319 ( .A1(n4293), .A2(n4295), .ZN(n4312) );
  AND2_X1 U4320 ( .A1(n4313), .A2(n4296), .ZN(n4311) );
  OR2_X1 U4321 ( .A1(n2723), .A2(n2574), .ZN(n4296) );
  OR2_X1 U4322 ( .A1(n4295), .A2(n4293), .ZN(n4313) );
  OR2_X1 U4323 ( .A1(n2570), .A2(n2567), .ZN(n4293) );
  INV_X1 U4324 ( .A(a_2_), .ZN(n2570) );
  OR2_X1 U4325 ( .A1(n4314), .A2(n4315), .ZN(n4295) );
  AND2_X1 U4326 ( .A1(n4289), .A2(n4291), .ZN(n4315) );
  AND2_X1 U4327 ( .A1(n4316), .A2(n4292), .ZN(n4314) );
  OR2_X1 U4328 ( .A1(n2723), .A2(n2578), .ZN(n4292) );
  OR2_X1 U4329 ( .A1(n4291), .A2(n4289), .ZN(n4316) );
  OR2_X1 U4330 ( .A1(n2574), .A2(n2567), .ZN(n4289) );
  INV_X1 U4331 ( .A(a_3_), .ZN(n2574) );
  OR2_X1 U4332 ( .A1(n4317), .A2(n4318), .ZN(n4291) );
  AND2_X1 U4333 ( .A1(n4285), .A2(n4287), .ZN(n4318) );
  AND2_X1 U4334 ( .A1(n4319), .A2(n4288), .ZN(n4317) );
  OR2_X1 U4335 ( .A1(n2723), .A2(n2582), .ZN(n4288) );
  OR2_X1 U4336 ( .A1(n4287), .A2(n4285), .ZN(n4319) );
  OR2_X1 U4337 ( .A1(n2578), .A2(n2567), .ZN(n4285) );
  INV_X1 U4338 ( .A(a_4_), .ZN(n2578) );
  OR2_X1 U4339 ( .A1(n4320), .A2(n4321), .ZN(n4287) );
  AND2_X1 U4340 ( .A1(n4281), .A2(n4283), .ZN(n4321) );
  AND2_X1 U4341 ( .A1(n4322), .A2(n4284), .ZN(n4320) );
  OR2_X1 U4342 ( .A1(n2723), .A2(n2586), .ZN(n4284) );
  OR2_X1 U4343 ( .A1(n4283), .A2(n4281), .ZN(n4322) );
  OR2_X1 U4344 ( .A1(n2582), .A2(n2567), .ZN(n4281) );
  INV_X1 U4345 ( .A(a_5_), .ZN(n2582) );
  OR2_X1 U4346 ( .A1(n4323), .A2(n4324), .ZN(n4283) );
  AND2_X1 U4347 ( .A1(n4277), .A2(n4279), .ZN(n4324) );
  AND2_X1 U4348 ( .A1(n4325), .A2(n4280), .ZN(n4323) );
  OR2_X1 U4349 ( .A1(n2723), .A2(n2590), .ZN(n4280) );
  OR2_X1 U4350 ( .A1(n4279), .A2(n4277), .ZN(n4325) );
  OR2_X1 U4351 ( .A1(n2586), .A2(n2567), .ZN(n4277) );
  INV_X1 U4352 ( .A(a_6_), .ZN(n2586) );
  OR2_X1 U4353 ( .A1(n4326), .A2(n4327), .ZN(n4279) );
  AND2_X1 U4354 ( .A1(n4273), .A2(n4275), .ZN(n4327) );
  AND2_X1 U4355 ( .A1(n4328), .A2(n4276), .ZN(n4326) );
  OR2_X1 U4356 ( .A1(n2723), .A2(n2594), .ZN(n4276) );
  OR2_X1 U4357 ( .A1(n4275), .A2(n4273), .ZN(n4328) );
  OR2_X1 U4358 ( .A1(n2590), .A2(n2567), .ZN(n4273) );
  INV_X1 U4359 ( .A(a_7_), .ZN(n2590) );
  OR2_X1 U4360 ( .A1(n4329), .A2(n4330), .ZN(n4275) );
  AND2_X1 U4361 ( .A1(n4269), .A2(n4271), .ZN(n4330) );
  AND2_X1 U4362 ( .A1(n4331), .A2(n4272), .ZN(n4329) );
  OR2_X1 U4363 ( .A1(n2723), .A2(n2318), .ZN(n4272) );
  OR2_X1 U4364 ( .A1(n4271), .A2(n4269), .ZN(n4331) );
  OR2_X1 U4365 ( .A1(n2594), .A2(n2567), .ZN(n4269) );
  INV_X1 U4366 ( .A(a_8_), .ZN(n2594) );
  OR2_X1 U4367 ( .A1(n4332), .A2(n4333), .ZN(n4271) );
  AND2_X1 U4368 ( .A1(n4266), .A2(n4268), .ZN(n4333) );
  AND2_X1 U4369 ( .A1(n4334), .A2(n4267), .ZN(n4332) );
  OR2_X1 U4370 ( .A1(n2723), .A2(n2293), .ZN(n4267) );
  OR2_X1 U4371 ( .A1(n4268), .A2(n4266), .ZN(n4334) );
  OR2_X1 U4372 ( .A1(n2318), .A2(n2567), .ZN(n4266) );
  INV_X1 U4373 ( .A(a_9_), .ZN(n2318) );
  OR2_X1 U4374 ( .A1(n4335), .A2(n4336), .ZN(n4268) );
  AND2_X1 U4375 ( .A1(n4262), .A2(n4264), .ZN(n4336) );
  AND2_X1 U4376 ( .A1(n4337), .A2(n4263), .ZN(n4335) );
  OR2_X1 U4377 ( .A1(n2723), .A2(n2268), .ZN(n4263) );
  OR2_X1 U4378 ( .A1(n4264), .A2(n4262), .ZN(n4337) );
  OR2_X1 U4379 ( .A1(n2293), .A2(n2567), .ZN(n4262) );
  INV_X1 U4380 ( .A(a_10_), .ZN(n2293) );
  OR2_X1 U4381 ( .A1(n4338), .A2(n4339), .ZN(n4264) );
  AND2_X1 U4382 ( .A1(n4258), .A2(n4260), .ZN(n4339) );
  AND2_X1 U4383 ( .A1(n4340), .A2(n4259), .ZN(n4338) );
  OR2_X1 U4384 ( .A1(n2723), .A2(n2243), .ZN(n4259) );
  OR2_X1 U4385 ( .A1(n4260), .A2(n4258), .ZN(n4340) );
  OR2_X1 U4386 ( .A1(n2268), .A2(n2567), .ZN(n4258) );
  INV_X1 U4387 ( .A(a_11_), .ZN(n2268) );
  OR2_X1 U4388 ( .A1(n4341), .A2(n4342), .ZN(n4260) );
  AND2_X1 U4389 ( .A1(n4254), .A2(n4256), .ZN(n4342) );
  AND2_X1 U4390 ( .A1(n4255), .A2(n4343), .ZN(n4341) );
  OR2_X1 U4391 ( .A1(n4256), .A2(n4254), .ZN(n4343) );
  OR2_X1 U4392 ( .A1(n2243), .A2(n2567), .ZN(n4254) );
  INV_X1 U4393 ( .A(a_12_), .ZN(n2243) );
  OR2_X1 U4394 ( .A1(n2723), .A2(n2218), .ZN(n4256) );
  AND2_X1 U4395 ( .A1(n4250), .A2(n4247), .ZN(n4255) );
  OR3_X1 U4396 ( .A1(n2723), .A2(n2567), .A3(n2913), .ZN(n4247) );
  OR2_X1 U4397 ( .A1(n2619), .A2(n2174), .ZN(n2913) );
  INV_X1 U4398 ( .A(a_15_), .ZN(n2619) );
  OR3_X1 U4399 ( .A1(n2723), .A2(n2174), .A3(n4252), .ZN(n4250) );
  OR2_X1 U4400 ( .A1(n2218), .A2(n2567), .ZN(n4252) );
  INV_X1 U4401 ( .A(b_1_), .ZN(n2567) );
  INV_X1 U4402 ( .A(a_13_), .ZN(n2218) );
  INV_X1 U4403 ( .A(a_14_), .ZN(n2174) );
  OR2_X1 U4404 ( .A1(n2723), .A2(n2566), .ZN(n4303) );
  INV_X1 U4405 ( .A(a_1_), .ZN(n2566) );
  INV_X1 U4406 ( .A(b_0_), .ZN(n2723) );
  AND2_X1 U4407 ( .A1(operation_0_), .A2(operation_1_), .ZN(n2126) );
endmodule

