module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n1009_, new_n238_, new_n479_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n158_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n144_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1074_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n1022_, new_n968_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n837_, new_n801_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n1096_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n994_, new_n982_, new_n422_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n138_, N81 );
not g001 ( new_n139_, N85 );
and g002 ( new_n140_, new_n138_, new_n139_ );
and g003 ( new_n141_, N81, N85 );
or g004 ( new_n142_, new_n140_, new_n141_ );
not g005 ( new_n143_, new_n142_ );
not g006 ( new_n144_, N89 );
not g007 ( new_n145_, N93 );
and g008 ( new_n146_, new_n144_, new_n145_ );
and g009 ( new_n147_, N89, N93 );
or g010 ( new_n148_, new_n146_, new_n147_ );
not g011 ( new_n149_, new_n148_ );
and g012 ( new_n150_, new_n143_, new_n149_ );
and g013 ( new_n151_, new_n142_, new_n148_ );
or g014 ( new_n152_, new_n150_, new_n151_ );
and g015 ( new_n153_, N65, N69 );
not g016 ( new_n154_, N65 );
not g017 ( new_n155_, N69 );
and g018 ( new_n156_, new_n154_, new_n155_ );
or g019 ( new_n157_, new_n156_, new_n153_ );
and g020 ( new_n158_, new_n157_, keyIn_0_5 );
or g021 ( new_n159_, new_n153_, keyIn_0_5 );
or g022 ( new_n160_, new_n159_, new_n156_ );
not g023 ( new_n161_, new_n160_ );
or g024 ( new_n162_, new_n161_, new_n158_ );
not g025 ( new_n163_, new_n162_ );
and g026 ( new_n164_, N73, N77 );
not g027 ( new_n165_, N73 );
not g028 ( new_n166_, N77 );
and g029 ( new_n167_, new_n165_, new_n166_ );
or g030 ( new_n168_, new_n167_, new_n164_ );
and g031 ( new_n169_, new_n168_, keyIn_0_6 );
not g032 ( new_n170_, new_n169_ );
or g033 ( new_n171_, new_n168_, keyIn_0_6 );
and g034 ( new_n172_, new_n170_, new_n171_ );
and g035 ( new_n173_, new_n163_, new_n172_ );
not g036 ( new_n174_, new_n173_ );
or g037 ( new_n175_, new_n163_, new_n172_ );
and g038 ( new_n176_, new_n174_, new_n175_ );
and g039 ( new_n177_, new_n176_, new_n152_ );
not g040 ( new_n178_, new_n152_ );
not g041 ( new_n179_, new_n176_ );
and g042 ( new_n180_, new_n179_, new_n178_ );
or g043 ( new_n181_, new_n180_, new_n177_ );
and g044 ( new_n182_, N129, N137 );
not g045 ( new_n183_, new_n182_ );
and g046 ( new_n184_, new_n181_, new_n183_ );
not g047 ( new_n185_, new_n184_ );
or g048 ( new_n186_, new_n181_, new_n183_ );
and g049 ( new_n187_, new_n185_, new_n186_ );
not g050 ( new_n188_, N17 );
and g051 ( new_n189_, new_n188_, N1 );
not g052 ( new_n190_, N1 );
and g053 ( new_n191_, new_n190_, N17 );
or g054 ( new_n192_, new_n189_, new_n191_ );
not g055 ( new_n193_, new_n192_ );
not g056 ( new_n194_, N33 );
not g057 ( new_n195_, N49 );
and g058 ( new_n196_, new_n194_, new_n195_ );
and g059 ( new_n197_, N33, N49 );
or g060 ( new_n198_, new_n196_, new_n197_ );
not g061 ( new_n199_, new_n198_ );
and g062 ( new_n200_, new_n193_, new_n199_ );
and g063 ( new_n201_, new_n192_, new_n198_ );
or g064 ( new_n202_, new_n200_, new_n201_ );
and g065 ( new_n203_, new_n187_, new_n202_ );
not g066 ( new_n204_, new_n203_ );
or g067 ( new_n205_, new_n187_, new_n202_ );
and g068 ( new_n206_, new_n204_, new_n205_ );
not g069 ( new_n207_, new_n206_ );
not g070 ( new_n208_, keyIn_0_18 );
not g071 ( new_n209_, N101 );
and g072 ( new_n210_, new_n209_, N97 );
not g073 ( new_n211_, N97 );
and g074 ( new_n212_, new_n211_, N101 );
or g075 ( new_n213_, new_n210_, new_n212_ );
and g076 ( new_n214_, N105, N109 );
not g077 ( new_n215_, N105 );
not g078 ( new_n216_, N109 );
and g079 ( new_n217_, new_n215_, new_n216_ );
or g080 ( new_n218_, new_n217_, new_n214_ );
and g081 ( new_n219_, new_n213_, new_n218_ );
not g082 ( new_n220_, new_n219_ );
or g083 ( new_n221_, new_n213_, new_n218_ );
and g084 ( new_n222_, new_n220_, new_n221_ );
and g085 ( new_n223_, new_n222_, new_n208_ );
not g086 ( new_n224_, new_n223_ );
or g087 ( new_n225_, new_n222_, new_n208_ );
and g088 ( new_n226_, new_n224_, new_n225_ );
and g089 ( new_n227_, N121, N125 );
not g090 ( new_n228_, N121 );
not g091 ( new_n229_, N125 );
and g092 ( new_n230_, new_n228_, new_n229_ );
or g093 ( new_n231_, new_n230_, new_n227_ );
or g094 ( new_n232_, new_n231_, keyIn_0_7 );
and g095 ( new_n233_, new_n231_, keyIn_0_7 );
not g096 ( new_n234_, new_n233_ );
and g097 ( new_n235_, new_n234_, new_n232_ );
not g098 ( new_n236_, N117 );
and g099 ( new_n237_, new_n236_, N113 );
not g100 ( new_n238_, N113 );
and g101 ( new_n239_, new_n238_, N117 );
or g102 ( new_n240_, new_n237_, new_n239_ );
not g103 ( new_n241_, new_n240_ );
and g104 ( new_n242_, new_n235_, new_n241_ );
not g105 ( new_n243_, new_n242_ );
or g106 ( new_n244_, new_n235_, new_n241_ );
and g107 ( new_n245_, new_n243_, new_n244_ );
not g108 ( new_n246_, new_n245_ );
and g109 ( new_n247_, new_n246_, keyIn_0_19 );
not g110 ( new_n248_, new_n247_ );
or g111 ( new_n249_, new_n246_, keyIn_0_19 );
and g112 ( new_n250_, new_n248_, new_n249_ );
or g113 ( new_n251_, new_n250_, new_n226_ );
not g114 ( new_n252_, new_n251_ );
and g115 ( new_n253_, new_n250_, new_n226_ );
or g116 ( new_n254_, new_n252_, new_n253_ );
and g117 ( new_n255_, new_n254_, keyIn_0_22 );
not g118 ( new_n256_, keyIn_0_22 );
not g119 ( new_n257_, new_n253_ );
and g120 ( new_n258_, new_n257_, new_n251_ );
and g121 ( new_n259_, new_n258_, new_n256_ );
or g122 ( new_n260_, new_n255_, new_n259_ );
not g123 ( new_n261_, keyIn_0_8 );
and g124 ( new_n262_, N130, N137 );
and g125 ( new_n263_, new_n262_, new_n261_ );
not g126 ( new_n264_, new_n263_ );
or g127 ( new_n265_, new_n262_, new_n261_ );
and g128 ( new_n266_, new_n264_, new_n265_ );
not g129 ( new_n267_, new_n266_ );
and g130 ( new_n268_, new_n260_, new_n267_ );
or g131 ( new_n269_, new_n258_, new_n256_ );
or g132 ( new_n270_, new_n254_, keyIn_0_22 );
and g133 ( new_n271_, new_n270_, new_n269_ );
and g134 ( new_n272_, new_n271_, new_n266_ );
or g135 ( new_n273_, new_n268_, new_n272_ );
not g136 ( new_n274_, N21 );
and g137 ( new_n275_, new_n274_, N5 );
not g138 ( new_n276_, N5 );
and g139 ( new_n277_, new_n276_, N21 );
or g140 ( new_n278_, new_n275_, new_n277_ );
and g141 ( new_n279_, new_n278_, keyIn_0_12 );
not g142 ( new_n280_, new_n279_ );
or g143 ( new_n281_, new_n278_, keyIn_0_12 );
and g144 ( new_n282_, new_n280_, new_n281_ );
not g145 ( new_n283_, N53 );
and g146 ( new_n284_, new_n283_, N37 );
not g147 ( new_n285_, N37 );
and g148 ( new_n286_, new_n285_, N53 );
or g149 ( new_n287_, new_n284_, new_n286_ );
and g150 ( new_n288_, new_n287_, keyIn_0_13 );
not g151 ( new_n289_, new_n288_ );
or g152 ( new_n290_, new_n287_, keyIn_0_13 );
and g153 ( new_n291_, new_n289_, new_n290_ );
and g154 ( new_n292_, new_n282_, new_n291_ );
not g155 ( new_n293_, new_n292_ );
or g156 ( new_n294_, new_n282_, new_n291_ );
and g157 ( new_n295_, new_n293_, new_n294_ );
not g158 ( new_n296_, new_n295_ );
or g159 ( new_n297_, new_n273_, new_n296_ );
or g160 ( new_n298_, new_n271_, new_n266_ );
or g161 ( new_n299_, new_n260_, new_n267_ );
and g162 ( new_n300_, new_n299_, new_n298_ );
or g163 ( new_n301_, new_n300_, new_n295_ );
and g164 ( new_n302_, new_n297_, new_n301_ );
and g165 ( new_n303_, new_n302_, new_n207_ );
not g166 ( new_n304_, keyIn_0_23 );
or g167 ( new_n305_, new_n250_, new_n178_ );
not g168 ( new_n306_, new_n305_ );
and g169 ( new_n307_, new_n250_, new_n178_ );
or g170 ( new_n308_, new_n306_, new_n307_ );
and g171 ( new_n309_, N132, N137 );
and g172 ( new_n310_, new_n309_, keyIn_0_9 );
not g173 ( new_n311_, new_n310_ );
or g174 ( new_n312_, new_n309_, keyIn_0_9 );
and g175 ( new_n313_, new_n311_, new_n312_ );
not g176 ( new_n314_, new_n313_ );
and g177 ( new_n315_, new_n308_, new_n314_ );
not g178 ( new_n316_, new_n307_ );
and g179 ( new_n317_, new_n316_, new_n305_ );
and g180 ( new_n318_, new_n317_, new_n313_ );
or g181 ( new_n319_, new_n315_, new_n318_ );
or g182 ( new_n320_, new_n319_, new_n304_ );
or g183 ( new_n321_, new_n317_, new_n313_ );
or g184 ( new_n322_, new_n308_, new_n314_ );
and g185 ( new_n323_, new_n322_, new_n321_ );
or g186 ( new_n324_, new_n323_, keyIn_0_23 );
and g187 ( new_n325_, new_n320_, new_n324_ );
not g188 ( new_n326_, N29 );
and g189 ( new_n327_, new_n326_, N13 );
not g190 ( new_n328_, N13 );
and g191 ( new_n329_, new_n328_, N29 );
or g192 ( new_n330_, new_n327_, new_n329_ );
and g193 ( new_n331_, new_n330_, keyIn_0_14 );
not g194 ( new_n332_, new_n331_ );
or g195 ( new_n333_, new_n330_, keyIn_0_14 );
and g196 ( new_n334_, new_n332_, new_n333_ );
not g197 ( new_n335_, new_n334_ );
not g198 ( new_n336_, N61 );
and g199 ( new_n337_, new_n336_, N45 );
not g200 ( new_n338_, N45 );
and g201 ( new_n339_, new_n338_, N61 );
or g202 ( new_n340_, new_n337_, new_n339_ );
and g203 ( new_n341_, new_n335_, new_n340_ );
not g204 ( new_n342_, new_n341_ );
or g205 ( new_n343_, new_n335_, new_n340_ );
and g206 ( new_n344_, new_n342_, new_n343_ );
and g207 ( new_n345_, new_n325_, new_n344_ );
not g208 ( new_n346_, new_n345_ );
and g209 ( new_n347_, new_n323_, keyIn_0_23 );
and g210 ( new_n348_, new_n319_, new_n304_ );
or g211 ( new_n349_, new_n348_, new_n347_ );
not g212 ( new_n350_, new_n344_ );
and g213 ( new_n351_, new_n349_, new_n350_ );
not g214 ( new_n352_, new_n351_ );
and g215 ( new_n353_, new_n352_, new_n346_ );
and g216 ( new_n354_, new_n179_, new_n226_ );
not g217 ( new_n355_, new_n354_ );
or g218 ( new_n356_, new_n179_, new_n226_ );
and g219 ( new_n357_, new_n355_, new_n356_ );
and g220 ( new_n358_, N131, N137 );
and g221 ( new_n359_, new_n357_, new_n358_ );
not g222 ( new_n360_, new_n357_ );
not g223 ( new_n361_, new_n358_ );
and g224 ( new_n362_, new_n360_, new_n361_ );
or g225 ( new_n363_, new_n362_, new_n359_ );
not g226 ( new_n364_, N9 );
not g227 ( new_n365_, N25 );
and g228 ( new_n366_, new_n364_, new_n365_ );
and g229 ( new_n367_, N9, N25 );
or g230 ( new_n368_, new_n366_, new_n367_ );
not g231 ( new_n369_, new_n368_ );
not g232 ( new_n370_, N41 );
not g233 ( new_n371_, N57 );
and g234 ( new_n372_, new_n370_, new_n371_ );
and g235 ( new_n373_, N41, N57 );
or g236 ( new_n374_, new_n372_, new_n373_ );
not g237 ( new_n375_, new_n374_ );
and g238 ( new_n376_, new_n369_, new_n375_ );
and g239 ( new_n377_, new_n368_, new_n374_ );
or g240 ( new_n378_, new_n376_, new_n377_ );
and g241 ( new_n379_, new_n363_, new_n378_ );
not g242 ( new_n380_, new_n359_ );
or g243 ( new_n381_, new_n357_, new_n358_ );
and g244 ( new_n382_, new_n380_, new_n381_ );
not g245 ( new_n383_, new_n378_ );
and g246 ( new_n384_, new_n382_, new_n383_ );
or g247 ( new_n385_, new_n379_, new_n384_ );
and g248 ( new_n386_, new_n385_, keyIn_0_24 );
not g249 ( new_n387_, keyIn_0_24 );
or g250 ( new_n388_, new_n382_, new_n383_ );
or g251 ( new_n389_, new_n363_, new_n378_ );
and g252 ( new_n390_, new_n389_, new_n388_ );
and g253 ( new_n391_, new_n390_, new_n387_ );
or g254 ( new_n392_, new_n386_, new_n391_ );
or g255 ( new_n393_, new_n392_, keyIn_0_26 );
not g256 ( new_n394_, keyIn_0_26 );
or g257 ( new_n395_, new_n390_, new_n387_ );
or g258 ( new_n396_, new_n385_, keyIn_0_24 );
and g259 ( new_n397_, new_n396_, new_n395_ );
or g260 ( new_n398_, new_n397_, new_n394_ );
and g261 ( new_n399_, new_n393_, new_n398_ );
and g262 ( new_n400_, new_n353_, new_n399_ );
and g263 ( new_n401_, new_n400_, new_n303_ );
or g264 ( new_n402_, new_n401_, keyIn_0_36 );
not g265 ( new_n403_, keyIn_0_36 );
and g266 ( new_n404_, new_n300_, new_n295_ );
and g267 ( new_n405_, new_n273_, new_n296_ );
or g268 ( new_n406_, new_n405_, new_n404_ );
or g269 ( new_n407_, new_n406_, new_n206_ );
or g270 ( new_n408_, new_n351_, new_n345_ );
and g271 ( new_n409_, new_n397_, new_n394_ );
and g272 ( new_n410_, new_n392_, keyIn_0_26 );
or g273 ( new_n411_, new_n410_, new_n409_ );
or g274 ( new_n412_, new_n411_, new_n408_ );
or g275 ( new_n413_, new_n412_, new_n407_ );
or g276 ( new_n414_, new_n413_, new_n403_ );
and g277 ( new_n415_, new_n414_, new_n402_ );
and g278 ( new_n416_, new_n392_, new_n206_ );
and g279 ( new_n417_, new_n408_, new_n416_ );
and g280 ( new_n418_, new_n417_, new_n302_ );
and g281 ( new_n419_, new_n406_, new_n416_ );
or g282 ( new_n420_, new_n206_, keyIn_0_25 );
and g283 ( new_n421_, new_n206_, keyIn_0_25 );
not g284 ( new_n422_, new_n421_ );
and g285 ( new_n423_, new_n422_, new_n420_ );
and g286 ( new_n424_, new_n423_, new_n397_ );
and g287 ( new_n425_, new_n302_, new_n424_ );
or g288 ( new_n426_, new_n419_, new_n425_ );
and g289 ( new_n427_, new_n426_, new_n353_ );
or g290 ( new_n428_, new_n427_, new_n418_ );
or g291 ( new_n429_, new_n415_, new_n428_ );
not g292 ( new_n430_, keyIn_0_21 );
and g293 ( new_n431_, new_n194_, keyIn_0_2 );
not g294 ( new_n432_, keyIn_0_2 );
and g295 ( new_n433_, new_n432_, N33 );
or g296 ( new_n434_, new_n431_, new_n433_ );
and g297 ( new_n435_, new_n434_, new_n285_ );
or g298 ( new_n436_, new_n432_, N33 );
or g299 ( new_n437_, new_n194_, keyIn_0_2 );
and g300 ( new_n438_, new_n436_, new_n437_ );
and g301 ( new_n439_, new_n438_, N37 );
or g302 ( new_n440_, new_n435_, new_n439_ );
not g303 ( new_n441_, keyIn_0_3 );
and g304 ( new_n442_, new_n370_, new_n338_ );
and g305 ( new_n443_, N41, N45 );
or g306 ( new_n444_, new_n442_, new_n443_ );
and g307 ( new_n445_, new_n444_, new_n441_ );
not g308 ( new_n446_, new_n443_ );
or g309 ( new_n447_, N41, N45 );
and g310 ( new_n448_, new_n447_, keyIn_0_3 );
and g311 ( new_n449_, new_n448_, new_n446_ );
or g312 ( new_n450_, new_n445_, new_n449_ );
and g313 ( new_n451_, new_n440_, new_n450_ );
or g314 ( new_n452_, new_n438_, N37 );
or g315 ( new_n453_, new_n434_, new_n285_ );
and g316 ( new_n454_, new_n453_, new_n452_ );
and g317 ( new_n455_, new_n446_, new_n447_ );
or g318 ( new_n456_, new_n455_, keyIn_0_3 );
not g319 ( new_n457_, new_n449_ );
and g320 ( new_n458_, new_n457_, new_n456_ );
and g321 ( new_n459_, new_n454_, new_n458_ );
or g322 ( new_n460_, new_n451_, new_n459_ );
and g323 ( new_n461_, new_n460_, keyIn_0_17 );
not g324 ( new_n462_, keyIn_0_17 );
or g325 ( new_n463_, new_n454_, new_n458_ );
or g326 ( new_n464_, new_n440_, new_n450_ );
and g327 ( new_n465_, new_n464_, new_n463_ );
and g328 ( new_n466_, new_n465_, new_n462_ );
or g329 ( new_n467_, new_n461_, new_n466_ );
and g330 ( new_n468_, new_n276_, N1 );
and g331 ( new_n469_, new_n190_, N5 );
or g332 ( new_n470_, new_n468_, new_n469_ );
not g333 ( new_n471_, new_n470_ );
and g334 ( new_n472_, new_n364_, new_n328_ );
and g335 ( new_n473_, N9, N13 );
or g336 ( new_n474_, new_n472_, new_n473_ );
not g337 ( new_n475_, new_n474_ );
and g338 ( new_n476_, new_n471_, new_n475_ );
and g339 ( new_n477_, new_n470_, new_n474_ );
or g340 ( new_n478_, new_n476_, new_n477_ );
and g341 ( new_n479_, new_n478_, keyIn_0_16 );
not g342 ( new_n480_, new_n479_ );
or g343 ( new_n481_, new_n478_, keyIn_0_16 );
and g344 ( new_n482_, new_n480_, new_n481_ );
and g345 ( new_n483_, new_n467_, new_n482_ );
or g346 ( new_n484_, new_n465_, new_n462_ );
or g347 ( new_n485_, new_n460_, keyIn_0_17 );
and g348 ( new_n486_, new_n485_, new_n484_ );
not g349 ( new_n487_, keyIn_0_16 );
not g350 ( new_n488_, new_n478_ );
and g351 ( new_n489_, new_n488_, new_n487_ );
or g352 ( new_n490_, new_n489_, new_n479_ );
and g353 ( new_n491_, new_n486_, new_n490_ );
or g354 ( new_n492_, new_n483_, new_n491_ );
and g355 ( new_n493_, new_n492_, new_n430_ );
or g356 ( new_n494_, new_n486_, new_n490_ );
or g357 ( new_n495_, new_n467_, new_n482_ );
and g358 ( new_n496_, new_n495_, new_n494_ );
and g359 ( new_n497_, new_n496_, keyIn_0_21 );
or g360 ( new_n498_, new_n493_, new_n497_ );
not g361 ( new_n499_, keyIn_0_10 );
and g362 ( new_n500_, N135, N137 );
and g363 ( new_n501_, new_n500_, new_n499_ );
not g364 ( new_n502_, new_n501_ );
or g365 ( new_n503_, new_n500_, new_n499_ );
and g366 ( new_n504_, new_n502_, new_n503_ );
not g367 ( new_n505_, new_n504_ );
and g368 ( new_n506_, new_n498_, new_n505_ );
or g369 ( new_n507_, new_n496_, keyIn_0_21 );
or g370 ( new_n508_, new_n492_, new_n430_ );
and g371 ( new_n509_, new_n508_, new_n507_ );
and g372 ( new_n510_, new_n509_, new_n504_ );
or g373 ( new_n511_, new_n506_, new_n510_ );
not g374 ( new_n512_, keyIn_0_20 );
and g375 ( new_n513_, new_n144_, N73 );
and g376 ( new_n514_, new_n165_, N89 );
or g377 ( new_n515_, new_n513_, new_n514_ );
not g378 ( new_n516_, new_n515_ );
and g379 ( new_n517_, new_n215_, new_n228_ );
and g380 ( new_n518_, N105, N121 );
or g381 ( new_n519_, new_n517_, new_n518_ );
not g382 ( new_n520_, new_n519_ );
and g383 ( new_n521_, new_n516_, new_n520_ );
and g384 ( new_n522_, new_n515_, new_n519_ );
or g385 ( new_n523_, new_n521_, new_n522_ );
and g386 ( new_n524_, new_n523_, new_n512_ );
not g387 ( new_n525_, new_n524_ );
or g388 ( new_n526_, new_n523_, new_n512_ );
and g389 ( new_n527_, new_n525_, new_n526_ );
not g390 ( new_n528_, new_n527_ );
and g391 ( new_n529_, new_n511_, new_n528_ );
or g392 ( new_n530_, new_n509_, new_n504_ );
or g393 ( new_n531_, new_n498_, new_n505_ );
and g394 ( new_n532_, new_n531_, new_n530_ );
and g395 ( new_n533_, new_n532_, new_n527_ );
or g396 ( new_n534_, new_n529_, new_n533_ );
and g397 ( new_n535_, new_n429_, new_n534_ );
not g398 ( new_n536_, keyIn_0_4 );
and g399 ( new_n537_, N57, N61 );
and g400 ( new_n538_, new_n371_, new_n336_ );
or g401 ( new_n539_, new_n538_, new_n537_ );
or g402 ( new_n540_, new_n539_, new_n536_ );
and g403 ( new_n541_, new_n539_, new_n536_ );
not g404 ( new_n542_, new_n541_ );
and g405 ( new_n543_, new_n542_, new_n540_ );
not g406 ( new_n544_, new_n543_ );
and g407 ( new_n545_, new_n195_, new_n283_ );
and g408 ( new_n546_, N49, N53 );
or g409 ( new_n547_, new_n545_, new_n546_ );
and g410 ( new_n548_, new_n544_, new_n547_ );
not g411 ( new_n549_, new_n548_ );
or g412 ( new_n550_, new_n544_, new_n547_ );
and g413 ( new_n551_, new_n549_, new_n550_ );
and g414 ( new_n552_, new_n188_, new_n274_ );
and g415 ( new_n553_, N17, N21 );
or g416 ( new_n554_, new_n552_, new_n553_ );
and g417 ( new_n555_, new_n554_, keyIn_0_0 );
not g418 ( new_n556_, new_n555_ );
or g419 ( new_n557_, new_n554_, keyIn_0_0 );
and g420 ( new_n558_, new_n556_, new_n557_ );
and g421 ( new_n559_, new_n365_, new_n326_ );
and g422 ( new_n560_, N25, N29 );
or g423 ( new_n561_, new_n559_, new_n560_ );
and g424 ( new_n562_, new_n561_, keyIn_0_1 );
not g425 ( new_n563_, new_n562_ );
or g426 ( new_n564_, new_n561_, keyIn_0_1 );
and g427 ( new_n565_, new_n563_, new_n564_ );
or g428 ( new_n566_, new_n558_, new_n565_ );
not g429 ( new_n567_, new_n566_ );
and g430 ( new_n568_, new_n558_, new_n565_ );
or g431 ( new_n569_, new_n567_, new_n568_ );
and g432 ( new_n570_, new_n551_, new_n569_ );
not g433 ( new_n571_, new_n570_ );
or g434 ( new_n572_, new_n551_, new_n569_ );
and g435 ( new_n573_, new_n571_, new_n572_ );
and g436 ( new_n574_, N136, N137 );
and g437 ( new_n575_, new_n574_, keyIn_0_11 );
not g438 ( new_n576_, new_n575_ );
or g439 ( new_n577_, new_n574_, keyIn_0_11 );
and g440 ( new_n578_, new_n576_, new_n577_ );
and g441 ( new_n579_, new_n573_, new_n578_ );
not g442 ( new_n580_, new_n572_ );
or g443 ( new_n581_, new_n580_, new_n570_ );
not g444 ( new_n582_, new_n578_ );
and g445 ( new_n583_, new_n581_, new_n582_ );
or g446 ( new_n584_, new_n583_, new_n579_ );
and g447 ( new_n585_, new_n166_, new_n145_ );
and g448 ( new_n586_, N77, N93 );
or g449 ( new_n587_, new_n585_, new_n586_ );
not g450 ( new_n588_, new_n587_ );
and g451 ( new_n589_, new_n216_, new_n229_ );
and g452 ( new_n590_, N109, N125 );
or g453 ( new_n591_, new_n589_, new_n590_ );
not g454 ( new_n592_, new_n591_ );
and g455 ( new_n593_, new_n588_, new_n592_ );
and g456 ( new_n594_, new_n587_, new_n591_ );
or g457 ( new_n595_, new_n593_, new_n594_ );
or g458 ( new_n596_, new_n584_, new_n595_ );
not g459 ( new_n597_, new_n579_ );
or g460 ( new_n598_, new_n573_, new_n578_ );
and g461 ( new_n599_, new_n597_, new_n598_ );
not g462 ( new_n600_, new_n595_ );
or g463 ( new_n601_, new_n599_, new_n600_ );
and g464 ( new_n602_, new_n601_, new_n596_ );
and g465 ( new_n603_, new_n467_, new_n551_ );
not g466 ( new_n604_, new_n603_ );
or g467 ( new_n605_, new_n467_, new_n551_ );
and g468 ( new_n606_, new_n604_, new_n605_ );
and g469 ( new_n607_, N134, N137 );
or g470 ( new_n608_, new_n606_, new_n607_ );
and g471 ( new_n609_, new_n606_, new_n607_ );
not g472 ( new_n610_, new_n609_ );
and g473 ( new_n611_, new_n610_, new_n608_ );
and g474 ( new_n612_, new_n155_, new_n139_ );
and g475 ( new_n613_, N69, N85 );
or g476 ( new_n614_, new_n612_, new_n613_ );
not g477 ( new_n615_, new_n614_ );
and g478 ( new_n616_, new_n209_, new_n236_ );
and g479 ( new_n617_, N101, N117 );
or g480 ( new_n618_, new_n616_, new_n617_ );
not g481 ( new_n619_, new_n618_ );
and g482 ( new_n620_, new_n615_, new_n619_ );
and g483 ( new_n621_, new_n614_, new_n618_ );
or g484 ( new_n622_, new_n620_, new_n621_ );
not g485 ( new_n623_, new_n622_ );
or g486 ( new_n624_, new_n611_, new_n623_ );
not g487 ( new_n625_, new_n608_ );
or g488 ( new_n626_, new_n625_, new_n609_ );
or g489 ( new_n627_, new_n626_, new_n622_ );
and g490 ( new_n628_, new_n627_, new_n624_ );
not g491 ( new_n629_, new_n568_ );
and g492 ( new_n630_, new_n629_, new_n566_ );
or g493 ( new_n631_, new_n490_, new_n630_ );
or g494 ( new_n632_, new_n569_, new_n482_ );
and g495 ( new_n633_, new_n632_, new_n631_ );
and g496 ( new_n634_, N133, N137 );
or g497 ( new_n635_, new_n633_, new_n634_ );
and g498 ( new_n636_, new_n569_, new_n482_ );
and g499 ( new_n637_, new_n490_, new_n630_ );
or g500 ( new_n638_, new_n636_, new_n637_ );
not g501 ( new_n639_, new_n634_ );
or g502 ( new_n640_, new_n638_, new_n639_ );
and g503 ( new_n641_, new_n640_, new_n635_ );
and g504 ( new_n642_, new_n211_, new_n238_ );
and g505 ( new_n643_, N97, N113 );
or g506 ( new_n644_, new_n642_, new_n643_ );
and g507 ( new_n645_, new_n644_, keyIn_0_15 );
not g508 ( new_n646_, new_n645_ );
or g509 ( new_n647_, new_n644_, keyIn_0_15 );
and g510 ( new_n648_, new_n646_, new_n647_ );
not g511 ( new_n649_, new_n648_ );
and g512 ( new_n650_, new_n154_, new_n138_ );
and g513 ( new_n651_, N65, N81 );
or g514 ( new_n652_, new_n650_, new_n651_ );
and g515 ( new_n653_, new_n649_, new_n652_ );
not g516 ( new_n654_, new_n653_ );
or g517 ( new_n655_, new_n649_, new_n652_ );
and g518 ( new_n656_, new_n654_, new_n655_ );
and g519 ( new_n657_, new_n641_, new_n656_ );
and g520 ( new_n658_, new_n638_, new_n639_ );
and g521 ( new_n659_, new_n633_, new_n634_ );
or g522 ( new_n660_, new_n658_, new_n659_ );
not g523 ( new_n661_, new_n656_ );
and g524 ( new_n662_, new_n660_, new_n661_ );
or g525 ( new_n663_, new_n662_, new_n657_ );
and g526 ( new_n664_, new_n628_, new_n663_ );
and g527 ( new_n665_, new_n664_, new_n602_ );
and g528 ( new_n666_, new_n535_, new_n665_ );
and g529 ( new_n667_, new_n666_, new_n207_ );
and g530 ( new_n668_, new_n667_, keyIn_0_41 );
not g531 ( new_n669_, new_n668_ );
or g532 ( new_n670_, new_n667_, keyIn_0_41 );
and g533 ( new_n671_, new_n669_, new_n670_ );
not g534 ( new_n672_, new_n671_ );
and g535 ( new_n673_, new_n672_, N1 );
and g536 ( new_n674_, new_n671_, new_n190_ );
or g537 ( N724, new_n673_, new_n674_ );
and g538 ( new_n676_, new_n666_, new_n406_ );
and g539 ( new_n677_, new_n676_, keyIn_0_42 );
not g540 ( new_n678_, new_n677_ );
or g541 ( new_n679_, new_n676_, keyIn_0_42 );
and g542 ( new_n680_, new_n678_, new_n679_ );
not g543 ( new_n681_, new_n680_ );
and g544 ( new_n682_, new_n681_, new_n276_ );
and g545 ( new_n683_, new_n680_, N5 );
or g546 ( N725, new_n682_, new_n683_ );
and g547 ( new_n685_, new_n666_, new_n397_ );
not g548 ( new_n686_, new_n685_ );
and g549 ( new_n687_, new_n686_, N9 );
and g550 ( new_n688_, new_n685_, new_n364_ );
or g551 ( N726, new_n687_, new_n688_ );
and g552 ( new_n690_, new_n666_, new_n408_ );
not g553 ( new_n691_, new_n690_ );
and g554 ( new_n692_, new_n691_, N13 );
and g555 ( new_n693_, new_n690_, new_n328_ );
or g556 ( N727, new_n692_, new_n693_ );
or g557 ( new_n695_, new_n532_, new_n527_ );
or g558 ( new_n696_, new_n511_, new_n528_ );
and g559 ( new_n697_, new_n696_, new_n695_ );
and g560 ( new_n698_, new_n599_, new_n600_ );
and g561 ( new_n699_, new_n584_, new_n595_ );
or g562 ( new_n700_, new_n698_, new_n699_ );
and g563 ( new_n701_, new_n664_, new_n700_ );
and g564 ( new_n702_, new_n701_, new_n697_ );
and g565 ( new_n703_, new_n429_, new_n702_ );
and g566 ( new_n704_, new_n703_, new_n207_ );
and g567 ( new_n705_, new_n704_, new_n188_ );
not g568 ( new_n706_, new_n705_ );
or g569 ( new_n707_, new_n704_, new_n188_ );
and g570 ( new_n708_, new_n706_, new_n707_ );
not g571 ( new_n709_, new_n708_ );
and g572 ( new_n710_, new_n709_, keyIn_0_54 );
not g573 ( new_n711_, keyIn_0_54 );
and g574 ( new_n712_, new_n708_, new_n711_ );
or g575 ( N728, new_n710_, new_n712_ );
and g576 ( new_n714_, new_n703_, new_n406_ );
and g577 ( new_n715_, new_n714_, new_n274_ );
not g578 ( new_n716_, new_n715_ );
or g579 ( new_n717_, new_n714_, new_n274_ );
and g580 ( new_n718_, new_n716_, new_n717_ );
not g581 ( new_n719_, new_n718_ );
and g582 ( new_n720_, new_n719_, keyIn_0_55 );
not g583 ( new_n721_, keyIn_0_55 );
and g584 ( new_n722_, new_n718_, new_n721_ );
or g585 ( N729, new_n720_, new_n722_ );
and g586 ( new_n724_, new_n703_, new_n397_ );
not g587 ( new_n725_, new_n724_ );
and g588 ( new_n726_, new_n725_, N25 );
and g589 ( new_n727_, new_n724_, new_n365_ );
or g590 ( N730, new_n726_, new_n727_ );
and g591 ( new_n729_, new_n703_, new_n408_ );
and g592 ( new_n730_, new_n729_, keyIn_0_43 );
not g593 ( new_n731_, new_n730_ );
or g594 ( new_n732_, new_n729_, keyIn_0_43 );
and g595 ( new_n733_, new_n731_, new_n732_ );
not g596 ( new_n734_, new_n733_ );
and g597 ( new_n735_, new_n734_, N29 );
and g598 ( new_n736_, new_n733_, new_n326_ );
or g599 ( N731, new_n735_, new_n736_ );
or g600 ( new_n738_, new_n628_, new_n663_ );
not g601 ( new_n739_, new_n738_ );
and g602 ( new_n740_, new_n739_, new_n602_ );
and g603 ( new_n741_, new_n535_, new_n740_ );
and g604 ( new_n742_, new_n741_, new_n207_ );
and g605 ( new_n743_, new_n742_, new_n194_ );
not g606 ( new_n744_, new_n743_ );
or g607 ( new_n745_, new_n742_, new_n194_ );
and g608 ( new_n746_, new_n744_, new_n745_ );
not g609 ( new_n747_, new_n746_ );
and g610 ( new_n748_, new_n747_, keyIn_0_56 );
not g611 ( new_n749_, keyIn_0_56 );
and g612 ( new_n750_, new_n746_, new_n749_ );
or g613 ( N732, new_n748_, new_n750_ );
and g614 ( new_n752_, new_n741_, new_n406_ );
and g615 ( new_n753_, new_n752_, N37 );
not g616 ( new_n754_, new_n753_ );
or g617 ( new_n755_, new_n752_, N37 );
and g618 ( new_n756_, new_n754_, new_n755_ );
not g619 ( new_n757_, new_n756_ );
and g620 ( new_n758_, new_n757_, keyIn_0_57 );
not g621 ( new_n759_, keyIn_0_57 );
and g622 ( new_n760_, new_n756_, new_n759_ );
or g623 ( N733, new_n758_, new_n760_ );
and g624 ( new_n762_, new_n741_, new_n397_ );
and g625 ( new_n763_, new_n762_, keyIn_0_44 );
not g626 ( new_n764_, new_n763_ );
or g627 ( new_n765_, new_n762_, keyIn_0_44 );
and g628 ( new_n766_, new_n764_, new_n765_ );
not g629 ( new_n767_, new_n766_ );
and g630 ( new_n768_, new_n767_, N41 );
and g631 ( new_n769_, new_n766_, new_n370_ );
or g632 ( N734, new_n768_, new_n769_ );
and g633 ( new_n771_, new_n741_, new_n408_ );
and g634 ( new_n772_, new_n771_, keyIn_0_45 );
not g635 ( new_n773_, keyIn_0_45 );
and g636 ( new_n774_, new_n413_, new_n403_ );
and g637 ( new_n775_, new_n401_, keyIn_0_36 );
or g638 ( new_n776_, new_n774_, new_n775_ );
not g639 ( new_n777_, new_n418_ );
not g640 ( new_n778_, new_n416_ );
or g641 ( new_n779_, new_n302_, new_n778_ );
not g642 ( new_n780_, new_n425_ );
and g643 ( new_n781_, new_n780_, new_n779_ );
or g644 ( new_n782_, new_n781_, new_n408_ );
and g645 ( new_n783_, new_n782_, new_n777_ );
and g646 ( new_n784_, new_n776_, new_n783_ );
or g647 ( new_n785_, new_n784_, new_n697_ );
or g648 ( new_n786_, new_n738_, new_n700_ );
or g649 ( new_n787_, new_n785_, new_n786_ );
or g650 ( new_n788_, new_n787_, new_n353_ );
and g651 ( new_n789_, new_n788_, new_n773_ );
or g652 ( new_n790_, new_n789_, new_n772_ );
and g653 ( new_n791_, new_n790_, N45 );
not g654 ( new_n792_, new_n772_ );
or g655 ( new_n793_, new_n771_, keyIn_0_45 );
and g656 ( new_n794_, new_n792_, new_n793_ );
and g657 ( new_n795_, new_n794_, new_n338_ );
or g658 ( new_n796_, new_n795_, new_n791_ );
and g659 ( new_n797_, new_n796_, keyIn_0_58 );
not g660 ( new_n798_, keyIn_0_58 );
or g661 ( new_n799_, new_n794_, new_n338_ );
or g662 ( new_n800_, new_n790_, N45 );
and g663 ( new_n801_, new_n799_, new_n800_ );
and g664 ( new_n802_, new_n801_, new_n798_ );
or g665 ( N735, new_n797_, new_n802_ );
not g666 ( new_n804_, keyIn_0_39 );
and g667 ( new_n805_, new_n534_, keyIn_0_27 );
not g668 ( new_n806_, new_n805_ );
or g669 ( new_n807_, new_n534_, keyIn_0_27 );
and g670 ( new_n808_, new_n806_, new_n807_ );
not g671 ( new_n809_, new_n808_ );
and g672 ( new_n810_, new_n739_, new_n700_ );
and g673 ( new_n811_, new_n809_, new_n810_ );
and g674 ( new_n812_, new_n429_, new_n811_ );
not g675 ( new_n813_, new_n812_ );
and g676 ( new_n814_, new_n813_, new_n804_ );
and g677 ( new_n815_, new_n812_, keyIn_0_39 );
or g678 ( new_n816_, new_n814_, new_n815_ );
and g679 ( new_n817_, new_n816_, new_n207_ );
or g680 ( new_n818_, new_n817_, new_n195_ );
and g681 ( new_n819_, new_n817_, new_n195_ );
not g682 ( new_n820_, new_n819_ );
and g683 ( new_n821_, new_n820_, new_n818_ );
not g684 ( new_n822_, new_n821_ );
and g685 ( new_n823_, new_n822_, keyIn_0_59 );
not g686 ( new_n824_, keyIn_0_59 );
and g687 ( new_n825_, new_n821_, new_n824_ );
or g688 ( N736, new_n823_, new_n825_ );
not g689 ( new_n827_, keyIn_0_46 );
and g690 ( new_n828_, new_n816_, new_n406_ );
or g691 ( new_n829_, new_n828_, new_n827_ );
and g692 ( new_n830_, new_n828_, new_n827_ );
not g693 ( new_n831_, new_n830_ );
and g694 ( new_n832_, new_n831_, new_n829_ );
not g695 ( new_n833_, new_n832_ );
and g696 ( new_n834_, new_n833_, N53 );
and g697 ( new_n835_, new_n832_, new_n283_ );
or g698 ( N737, new_n834_, new_n835_ );
and g699 ( new_n837_, new_n816_, new_n397_ );
not g700 ( new_n838_, new_n837_ );
and g701 ( new_n839_, new_n838_, N57 );
and g702 ( new_n840_, new_n837_, new_n371_ );
or g703 ( N738, new_n839_, new_n840_ );
and g704 ( new_n842_, new_n816_, new_n408_ );
not g705 ( new_n843_, new_n842_ );
and g706 ( new_n844_, new_n843_, N61 );
and g707 ( new_n845_, new_n842_, new_n336_ );
or g708 ( N739, new_n844_, new_n845_ );
or g709 ( new_n847_, new_n660_, new_n661_ );
or g710 ( new_n848_, new_n641_, new_n656_ );
and g711 ( new_n849_, new_n847_, new_n848_ );
not g712 ( new_n850_, keyIn_0_40 );
not g713 ( new_n851_, keyIn_0_38 );
not g714 ( new_n852_, keyIn_0_37 );
not g715 ( new_n853_, keyIn_0_31 );
and g716 ( new_n854_, new_n697_, new_n853_ );
not g717 ( new_n855_, new_n854_ );
or g718 ( new_n856_, new_n697_, new_n853_ );
and g719 ( new_n857_, new_n740_, new_n856_ );
and g720 ( new_n858_, new_n857_, new_n855_ );
and g721 ( new_n859_, new_n858_, new_n852_ );
not g722 ( new_n860_, new_n859_ );
or g723 ( new_n861_, new_n858_, new_n852_ );
not g724 ( new_n862_, keyIn_0_32 );
and g725 ( new_n863_, new_n697_, new_n862_ );
and g726 ( new_n864_, new_n534_, keyIn_0_32 );
and g727 ( new_n865_, new_n626_, new_n622_ );
and g728 ( new_n866_, new_n611_, new_n623_ );
or g729 ( new_n867_, new_n865_, new_n866_ );
or g730 ( new_n868_, new_n867_, new_n849_ );
and g731 ( new_n869_, new_n602_, keyIn_0_33 );
not g732 ( new_n870_, keyIn_0_33 );
and g733 ( new_n871_, new_n700_, new_n870_ );
or g734 ( new_n872_, new_n871_, new_n869_ );
or g735 ( new_n873_, new_n868_, new_n872_ );
or g736 ( new_n874_, new_n864_, new_n873_ );
or g737 ( new_n875_, new_n874_, new_n863_ );
and g738 ( new_n876_, new_n867_, keyIn_0_28 );
not g739 ( new_n877_, new_n876_ );
not g740 ( new_n878_, keyIn_0_28 );
and g741 ( new_n879_, new_n628_, new_n878_ );
not g742 ( new_n880_, new_n879_ );
and g743 ( new_n881_, new_n880_, new_n877_ );
and g744 ( new_n882_, new_n700_, new_n849_ );
not g745 ( new_n883_, new_n882_ );
or g746 ( new_n884_, new_n534_, new_n883_ );
or g747 ( new_n885_, new_n881_, new_n884_ );
and g748 ( new_n886_, new_n602_, keyIn_0_30 );
not g749 ( new_n887_, keyIn_0_30 );
and g750 ( new_n888_, new_n700_, new_n887_ );
or g751 ( new_n889_, new_n888_, new_n886_ );
not g752 ( new_n890_, keyIn_0_29 );
or g753 ( new_n891_, new_n849_, new_n890_ );
or g754 ( new_n892_, new_n663_, keyIn_0_29 );
and g755 ( new_n893_, new_n892_, new_n891_ );
and g756 ( new_n894_, new_n893_, new_n628_ );
and g757 ( new_n895_, new_n894_, new_n889_ );
and g758 ( new_n896_, new_n895_, new_n534_ );
not g759 ( new_n897_, new_n896_ );
and g760 ( new_n898_, new_n885_, new_n897_ );
and g761 ( new_n899_, new_n898_, new_n875_ );
and g762 ( new_n900_, new_n899_, new_n861_ );
and g763 ( new_n901_, new_n900_, new_n860_ );
or g764 ( new_n902_, new_n901_, new_n851_ );
and g765 ( new_n903_, new_n534_, keyIn_0_31 );
or g766 ( new_n904_, new_n903_, new_n786_ );
or g767 ( new_n905_, new_n904_, new_n854_ );
and g768 ( new_n906_, new_n905_, keyIn_0_37 );
not g769 ( new_n907_, new_n863_ );
or g770 ( new_n908_, new_n697_, new_n862_ );
not g771 ( new_n909_, new_n872_ );
and g772 ( new_n910_, new_n909_, new_n664_ );
and g773 ( new_n911_, new_n908_, new_n910_ );
and g774 ( new_n912_, new_n911_, new_n907_ );
or g775 ( new_n913_, new_n876_, new_n879_ );
and g776 ( new_n914_, new_n697_, new_n882_ );
and g777 ( new_n915_, new_n914_, new_n913_ );
or g778 ( new_n916_, new_n915_, new_n896_ );
or g779 ( new_n917_, new_n912_, new_n916_ );
or g780 ( new_n918_, new_n917_, new_n906_ );
or g781 ( new_n919_, new_n918_, new_n859_ );
or g782 ( new_n920_, new_n919_, keyIn_0_38 );
and g783 ( new_n921_, new_n920_, new_n902_ );
and g784 ( new_n922_, new_n353_, new_n397_ );
and g785 ( new_n923_, new_n922_, new_n303_ );
and g786 ( new_n924_, new_n921_, new_n923_ );
or g787 ( new_n925_, new_n924_, new_n850_ );
and g788 ( new_n926_, new_n919_, keyIn_0_38 );
and g789 ( new_n927_, new_n901_, new_n851_ );
or g790 ( new_n928_, new_n926_, new_n927_ );
not g791 ( new_n929_, new_n923_ );
or g792 ( new_n930_, new_n928_, new_n929_ );
or g793 ( new_n931_, new_n930_, keyIn_0_40 );
and g794 ( new_n932_, new_n931_, new_n925_ );
or g795 ( new_n933_, new_n932_, new_n849_ );
and g796 ( new_n934_, new_n933_, keyIn_0_47 );
not g797 ( new_n935_, keyIn_0_47 );
and g798 ( new_n936_, new_n930_, keyIn_0_40 );
and g799 ( new_n937_, new_n924_, new_n850_ );
or g800 ( new_n938_, new_n936_, new_n937_ );
and g801 ( new_n939_, new_n938_, new_n663_ );
and g802 ( new_n940_, new_n939_, new_n935_ );
or g803 ( new_n941_, new_n934_, new_n940_ );
and g804 ( new_n942_, new_n941_, new_n154_ );
or g805 ( new_n943_, new_n939_, new_n935_ );
or g806 ( new_n944_, new_n933_, keyIn_0_47 );
and g807 ( new_n945_, new_n944_, new_n943_ );
and g808 ( new_n946_, new_n945_, N65 );
or g809 ( N740, new_n942_, new_n946_ );
or g810 ( new_n948_, new_n932_, new_n628_ );
and g811 ( new_n949_, new_n948_, keyIn_0_48 );
not g812 ( new_n950_, keyIn_0_48 );
and g813 ( new_n951_, new_n938_, new_n867_ );
and g814 ( new_n952_, new_n951_, new_n950_ );
or g815 ( new_n953_, new_n949_, new_n952_ );
and g816 ( new_n954_, new_n953_, new_n155_ );
or g817 ( new_n955_, new_n951_, new_n950_ );
or g818 ( new_n956_, new_n948_, keyIn_0_48 );
and g819 ( new_n957_, new_n956_, new_n955_ );
and g820 ( new_n958_, new_n957_, N69 );
or g821 ( N741, new_n954_, new_n958_ );
and g822 ( new_n960_, new_n938_, new_n534_ );
not g823 ( new_n961_, new_n960_ );
and g824 ( new_n962_, new_n961_, N73 );
and g825 ( new_n963_, new_n960_, new_n165_ );
or g826 ( N742, new_n962_, new_n963_ );
or g827 ( new_n965_, new_n932_, new_n602_ );
and g828 ( new_n966_, new_n965_, N77 );
and g829 ( new_n967_, new_n938_, new_n700_ );
and g830 ( new_n968_, new_n967_, new_n166_ );
or g831 ( new_n969_, new_n966_, new_n968_ );
and g832 ( new_n970_, new_n969_, keyIn_0_60 );
not g833 ( new_n971_, keyIn_0_60 );
or g834 ( new_n972_, new_n967_, new_n166_ );
or g835 ( new_n973_, new_n965_, N77 );
and g836 ( new_n974_, new_n973_, new_n972_ );
and g837 ( new_n975_, new_n974_, new_n971_ );
or g838 ( N743, new_n970_, new_n975_ );
not g839 ( new_n977_, keyIn_0_34 );
and g840 ( new_n978_, new_n302_, new_n977_ );
not g841 ( new_n979_, new_n978_ );
and g842 ( new_n980_, new_n406_, keyIn_0_34 );
not g843 ( new_n981_, new_n980_ );
and g844 ( new_n982_, new_n392_, new_n207_ );
and g845 ( new_n983_, new_n408_, new_n982_ );
and g846 ( new_n984_, new_n981_, new_n983_ );
and g847 ( new_n985_, new_n984_, new_n979_ );
and g848 ( new_n986_, new_n921_, new_n985_ );
and g849 ( new_n987_, new_n986_, new_n663_ );
not g850 ( new_n988_, new_n987_ );
and g851 ( new_n989_, new_n988_, N81 );
and g852 ( new_n990_, new_n987_, new_n138_ );
or g853 ( N744, new_n989_, new_n990_ );
and g854 ( new_n992_, new_n986_, new_n867_ );
not g855 ( new_n993_, new_n992_ );
and g856 ( new_n994_, new_n993_, keyIn_0_49 );
not g857 ( new_n995_, keyIn_0_49 );
and g858 ( new_n996_, new_n992_, new_n995_ );
or g859 ( new_n997_, new_n994_, new_n996_ );
and g860 ( new_n998_, new_n997_, N85 );
not g861 ( new_n999_, new_n997_ );
and g862 ( new_n1000_, new_n999_, new_n139_ );
or g863 ( N745, new_n1000_, new_n998_ );
and g864 ( new_n1002_, new_n986_, new_n534_ );
not g865 ( new_n1003_, new_n1002_ );
and g866 ( new_n1004_, new_n1003_, N89 );
and g867 ( new_n1005_, new_n1002_, new_n144_ );
or g868 ( new_n1006_, new_n1004_, new_n1005_ );
and g869 ( new_n1007_, new_n1006_, keyIn_0_61 );
not g870 ( new_n1008_, keyIn_0_61 );
not g871 ( new_n1009_, new_n1006_ );
and g872 ( new_n1010_, new_n1009_, new_n1008_ );
or g873 ( N746, new_n1010_, new_n1007_ );
and g874 ( new_n1012_, new_n986_, new_n700_ );
not g875 ( new_n1013_, new_n1012_ );
and g876 ( new_n1014_, new_n1013_, N93 );
and g877 ( new_n1015_, new_n1012_, new_n145_ );
or g878 ( N747, new_n1014_, new_n1015_ );
and g879 ( new_n1017_, new_n206_, keyIn_0_35 );
not g880 ( new_n1018_, new_n1017_ );
or g881 ( new_n1019_, new_n206_, keyIn_0_35 );
and g882 ( new_n1020_, new_n1018_, new_n1019_ );
and g883 ( new_n1021_, new_n406_, new_n1020_ );
and g884 ( new_n1022_, new_n922_, new_n1021_ );
and g885 ( new_n1023_, new_n921_, new_n1022_ );
and g886 ( new_n1024_, new_n1023_, new_n663_ );
not g887 ( new_n1025_, new_n1024_ );
and g888 ( new_n1026_, new_n1025_, N97 );
and g889 ( new_n1027_, new_n1024_, new_n211_ );
or g890 ( N748, new_n1026_, new_n1027_ );
and g891 ( new_n1029_, new_n1023_, new_n867_ );
not g892 ( new_n1030_, new_n1029_ );
and g893 ( new_n1031_, new_n1030_, keyIn_0_50 );
not g894 ( new_n1032_, keyIn_0_50 );
and g895 ( new_n1033_, new_n1029_, new_n1032_ );
or g896 ( new_n1034_, new_n1031_, new_n1033_ );
and g897 ( new_n1035_, new_n1034_, N101 );
not g898 ( new_n1036_, new_n1034_ );
and g899 ( new_n1037_, new_n1036_, new_n209_ );
or g900 ( N749, new_n1037_, new_n1035_ );
and g901 ( new_n1039_, new_n1023_, new_n534_ );
not g902 ( new_n1040_, new_n1039_ );
and g903 ( new_n1041_, new_n1040_, N105 );
and g904 ( new_n1042_, new_n1039_, new_n215_ );
or g905 ( N750, new_n1041_, new_n1042_ );
and g906 ( new_n1044_, new_n1023_, new_n700_ );
not g907 ( new_n1045_, new_n1044_ );
and g908 ( new_n1046_, new_n1045_, N109 );
and g909 ( new_n1047_, new_n1044_, new_n216_ );
or g910 ( N751, new_n1046_, new_n1047_ );
and g911 ( new_n1049_, new_n419_, new_n408_ );
and g912 ( new_n1050_, new_n921_, new_n1049_ );
and g913 ( new_n1051_, new_n1050_, new_n663_ );
not g914 ( new_n1052_, new_n1051_ );
and g915 ( new_n1053_, new_n1052_, N113 );
and g916 ( new_n1054_, new_n1051_, new_n238_ );
or g917 ( N752, new_n1053_, new_n1054_ );
and g918 ( new_n1056_, new_n1050_, new_n867_ );
not g919 ( new_n1057_, new_n1056_ );
and g920 ( new_n1058_, new_n1057_, keyIn_0_51 );
not g921 ( new_n1059_, keyIn_0_51 );
and g922 ( new_n1060_, new_n1056_, new_n1059_ );
or g923 ( new_n1061_, new_n1058_, new_n1060_ );
and g924 ( new_n1062_, new_n1061_, new_n236_ );
not g925 ( new_n1063_, new_n1061_ );
and g926 ( new_n1064_, new_n1063_, N117 );
or g927 ( N753, new_n1064_, new_n1062_ );
not g928 ( new_n1066_, keyIn_0_62 );
not g929 ( new_n1067_, keyIn_0_52 );
and g930 ( new_n1068_, new_n1050_, new_n534_ );
and g931 ( new_n1069_, new_n1068_, new_n1067_ );
not g932 ( new_n1070_, new_n1049_ );
or g933 ( new_n1071_, new_n928_, new_n1070_ );
or g934 ( new_n1072_, new_n1071_, new_n697_ );
and g935 ( new_n1073_, new_n1072_, keyIn_0_52 );
or g936 ( new_n1074_, new_n1073_, new_n1069_ );
and g937 ( new_n1075_, new_n1074_, new_n228_ );
or g938 ( new_n1076_, new_n1072_, keyIn_0_52 );
or g939 ( new_n1077_, new_n1068_, new_n1067_ );
and g940 ( new_n1078_, new_n1076_, new_n1077_ );
and g941 ( new_n1079_, new_n1078_, N121 );
or g942 ( new_n1080_, new_n1075_, new_n1079_ );
and g943 ( new_n1081_, new_n1080_, new_n1066_ );
or g944 ( new_n1082_, new_n1078_, N121 );
or g945 ( new_n1083_, new_n1074_, new_n228_ );
and g946 ( new_n1084_, new_n1082_, new_n1083_ );
and g947 ( new_n1085_, new_n1084_, keyIn_0_62 );
or g948 ( N754, new_n1081_, new_n1085_ );
not g949 ( new_n1087_, keyIn_0_63 );
not g950 ( new_n1088_, keyIn_0_53 );
and g951 ( new_n1089_, new_n1050_, new_n700_ );
and g952 ( new_n1090_, new_n1089_, new_n1088_ );
or g953 ( new_n1091_, new_n1071_, new_n602_ );
and g954 ( new_n1092_, new_n1091_, keyIn_0_53 );
or g955 ( new_n1093_, new_n1092_, new_n1090_ );
and g956 ( new_n1094_, new_n1093_, N125 );
or g957 ( new_n1095_, new_n1091_, keyIn_0_53 );
or g958 ( new_n1096_, new_n1089_, new_n1088_ );
and g959 ( new_n1097_, new_n1095_, new_n1096_ );
and g960 ( new_n1098_, new_n1097_, new_n229_ );
or g961 ( new_n1099_, new_n1094_, new_n1098_ );
and g962 ( new_n1100_, new_n1099_, new_n1087_ );
or g963 ( new_n1101_, new_n1097_, new_n229_ );
or g964 ( new_n1102_, new_n1093_, N125 );
and g965 ( new_n1103_, new_n1101_, new_n1102_ );
and g966 ( new_n1104_, new_n1103_, keyIn_0_63 );
or g967 ( N755, new_n1100_, new_n1104_ );
endmodule