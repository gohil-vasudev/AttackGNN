module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n246_, new_n682_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n840_, new_n735_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n953_, new_n257_, new_n481_, new_n212_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n903_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n385_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n650_, new_n708_, new_n750_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n394_, new_n299_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n426_, new_n235_, new_n398_, new_n301_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n668_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n276_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n860_, new_n306_, new_n494_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n749_, new_n861_, new_n310_, new_n275_, new_n998_, new_n352_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n824_, new_n520_, new_n1001_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n231_, new_n219_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n285_, new_n692_, new_n502_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n252_, new_n585_, new_n751_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n712_, new_n1017_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n434_, new_n200_, new_n947_, new_n994_, new_n422_, new_n964_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n172_, keyIn_0_21 );
or g001 ( new_n173_, keyIn_0_12, N102 );
and g002 ( new_n174_, keyIn_0_12, N102 );
not g003 ( new_n175_, new_n174_ );
and g004 ( new_n176_, new_n175_, N108, new_n173_ );
or g005 ( new_n177_, new_n176_, new_n172_ );
not g006 ( new_n178_, N108 );
not g007 ( new_n179_, new_n173_ );
or g008 ( new_n180_, new_n179_, new_n174_, keyIn_0_21, new_n178_ );
and g009 ( new_n181_, new_n177_, new_n180_ );
not g010 ( new_n182_, N95 );
not g011 ( new_n183_, keyIn_0_11 );
or g012 ( new_n184_, new_n183_, N89 );
not g013 ( new_n185_, N89 );
or g014 ( new_n186_, new_n185_, keyIn_0_11 );
and g015 ( new_n187_, new_n184_, new_n186_ );
or g016 ( new_n188_, new_n187_, keyIn_0_20, new_n182_ );
not g017 ( new_n189_, keyIn_0_20 );
and g018 ( new_n190_, new_n185_, keyIn_0_11 );
and g019 ( new_n191_, new_n183_, N89 );
or g020 ( new_n192_, new_n190_, new_n191_ );
and g021 ( new_n193_, new_n192_, N95 );
or g022 ( new_n194_, new_n193_, new_n189_ );
or g023 ( new_n195_, keyIn_0_7, N50 );
and g024 ( new_n196_, keyIn_0_7, N50 );
not g025 ( new_n197_, new_n196_ );
and g026 ( new_n198_, new_n197_, keyIn_0_19, N56, new_n195_ );
not g027 ( new_n199_, keyIn_0_19 );
not g028 ( new_n200_, N56 );
not g029 ( new_n201_, keyIn_0_7 );
not g030 ( new_n202_, N50 );
and g031 ( new_n203_, new_n201_, new_n202_ );
or g032 ( new_n204_, new_n203_, new_n200_, new_n196_ );
and g033 ( new_n205_, new_n204_, new_n199_ );
or g034 ( new_n206_, new_n205_, new_n198_ );
and g035 ( new_n207_, new_n206_, new_n181_, new_n188_, new_n194_ );
not g036 ( new_n208_, keyIn_0_18 );
not g037 ( new_n209_, N43 );
not g038 ( new_n210_, keyIn_0_6 );
or g039 ( new_n211_, new_n210_, N37 );
not g040 ( new_n212_, N37 );
or g041 ( new_n213_, new_n212_, keyIn_0_6 );
and g042 ( new_n214_, new_n211_, new_n213_ );
or g043 ( new_n215_, new_n214_, new_n209_ );
and g044 ( new_n216_, new_n215_, new_n208_ );
not g045 ( new_n217_, new_n214_ );
and g046 ( new_n218_, new_n217_, keyIn_0_18, N43 );
or g047 ( new_n219_, new_n216_, new_n218_ );
not g048 ( new_n220_, N82 );
not g049 ( new_n221_, keyIn_0_9 );
and g050 ( new_n222_, new_n221_, N76 );
not g051 ( new_n223_, N76 );
and g052 ( new_n224_, new_n223_, keyIn_0_9 );
or g053 ( new_n225_, new_n222_, new_n224_, new_n220_ );
not g054 ( new_n226_, N17 );
and g055 ( new_n227_, keyIn_0_2, N11 );
not g056 ( new_n228_, new_n227_ );
or g057 ( new_n229_, keyIn_0_2, N11 );
and g058 ( new_n230_, new_n228_, new_n229_ );
or g059 ( new_n231_, new_n230_, new_n226_ );
not g060 ( new_n232_, N63 );
and g061 ( new_n233_, new_n232_, N69 );
not g062 ( new_n234_, new_n233_ );
and g063 ( new_n235_, new_n231_, new_n225_, new_n234_ );
not g064 ( new_n236_, keyIn_0_14 );
or g065 ( new_n237_, keyIn_0_0, N1 );
not g066 ( new_n238_, new_n237_ );
and g067 ( new_n239_, keyIn_0_0, N1 );
or g068 ( new_n240_, new_n238_, new_n239_ );
and g069 ( new_n241_, new_n240_, N4 );
or g070 ( new_n242_, new_n241_, new_n236_ );
not g071 ( new_n243_, N4 );
not g072 ( new_n244_, new_n240_ );
or g073 ( new_n245_, new_n244_, keyIn_0_14, new_n243_ );
not g074 ( new_n246_, keyIn_0_17 );
not g075 ( new_n247_, N30 );
not g076 ( new_n248_, keyIn_0_4 );
not g077 ( new_n249_, N24 );
and g078 ( new_n250_, new_n248_, new_n249_ );
and g079 ( new_n251_, keyIn_0_4, N24 );
or g080 ( new_n252_, new_n250_, new_n247_, new_n251_ );
and g081 ( new_n253_, new_n252_, new_n246_ );
not g082 ( new_n254_, new_n250_ );
not g083 ( new_n255_, new_n251_ );
and g084 ( new_n256_, new_n254_, keyIn_0_17, N30, new_n255_ );
or g085 ( new_n257_, new_n253_, new_n256_ );
and g086 ( new_n258_, new_n257_, new_n242_, new_n245_ );
and g087 ( new_n259_, new_n207_, new_n258_, new_n219_, new_n235_ );
not g088 ( new_n260_, new_n259_ );
and g089 ( new_n261_, new_n260_, keyIn_0_38 );
not g090 ( new_n262_, keyIn_0_38 );
and g091 ( new_n263_, new_n259_, new_n262_ );
or g092 ( N223, new_n261_, new_n263_ );
not g093 ( new_n265_, keyIn_0_80 );
not g094 ( new_n266_, keyIn_0_59 );
not g095 ( new_n267_, keyIn_0_43 );
not g096 ( new_n268_, keyIn_0_37 );
or g097 ( new_n269_, new_n259_, new_n268_ );
and g098 ( new_n270_, new_n219_, new_n235_ );
and g099 ( new_n271_, new_n270_, new_n268_, new_n207_, new_n258_ );
not g100 ( new_n272_, new_n271_ );
and g101 ( new_n273_, new_n269_, new_n272_ );
or g102 ( new_n274_, new_n273_, new_n233_ );
and g103 ( new_n275_, new_n269_, new_n233_, new_n272_ );
not g104 ( new_n276_, new_n275_ );
and g105 ( new_n277_, new_n274_, new_n276_ );
or g106 ( new_n278_, new_n277_, new_n267_ );
and g107 ( new_n279_, new_n274_, new_n267_, new_n276_ );
not g108 ( new_n280_, new_n279_ );
and g109 ( new_n281_, new_n278_, new_n280_ );
not g110 ( new_n282_, N73 );
and g111 ( new_n283_, new_n282_, N69 );
and g112 ( new_n284_, new_n283_, keyIn_0_29 );
not g113 ( new_n285_, new_n284_ );
or g114 ( new_n286_, new_n283_, keyIn_0_29 );
and g115 ( new_n287_, new_n285_, new_n286_ );
or g116 ( new_n288_, new_n281_, new_n287_ );
and g117 ( new_n289_, new_n288_, new_n266_ );
not g118 ( new_n290_, new_n281_ );
not g119 ( new_n291_, new_n287_ );
and g120 ( new_n292_, new_n290_, keyIn_0_59, new_n291_ );
or g121 ( new_n293_, new_n289_, new_n292_ );
not g122 ( new_n294_, keyIn_0_41 );
not g123 ( new_n295_, new_n219_ );
or g124 ( new_n296_, new_n273_, new_n295_ );
and g125 ( new_n297_, new_n273_, new_n295_ );
not g126 ( new_n298_, new_n297_ );
and g127 ( new_n299_, new_n298_, new_n296_ );
or g128 ( new_n300_, new_n299_, new_n294_ );
and g129 ( new_n301_, new_n299_, new_n294_ );
not g130 ( new_n302_, new_n301_ );
not g131 ( new_n303_, keyIn_0_25 );
not g132 ( new_n304_, N47 );
and g133 ( new_n305_, new_n304_, N43 );
or g134 ( new_n306_, new_n305_, new_n303_ );
or g135 ( new_n307_, new_n209_, keyIn_0_25, N47 );
and g136 ( new_n308_, new_n306_, new_n307_ );
and g137 ( new_n309_, new_n302_, new_n300_, new_n308_ );
or g138 ( new_n310_, new_n309_, keyIn_0_58 );
and g139 ( new_n311_, new_n302_, keyIn_0_58, new_n300_, new_n308_ );
not g140 ( new_n312_, new_n311_ );
and g141 ( new_n313_, new_n310_, new_n312_ );
not g142 ( new_n314_, keyIn_0_62 );
not g143 ( new_n315_, new_n181_ );
or g144 ( new_n316_, new_n273_, new_n315_ );
not g145 ( new_n317_, new_n269_ );
or g146 ( new_n318_, new_n317_, new_n181_, new_n271_ );
and g147 ( new_n319_, new_n316_, keyIn_0_47, new_n318_ );
not g148 ( new_n320_, new_n319_ );
and g149 ( new_n321_, new_n316_, new_n318_ );
or g150 ( new_n322_, new_n321_, keyIn_0_47 );
and g151 ( new_n323_, new_n322_, new_n320_ );
not g152 ( new_n324_, new_n323_ );
not g153 ( new_n325_, keyIn_0_35 );
not g154 ( new_n326_, N112 );
and g155 ( new_n327_, keyIn_0_13, N108 );
not g156 ( new_n328_, new_n327_ );
or g157 ( new_n329_, keyIn_0_13, N108 );
and g158 ( new_n330_, new_n328_, new_n329_ );
not g159 ( new_n331_, new_n330_ );
and g160 ( new_n332_, new_n331_, new_n326_ );
not g161 ( new_n333_, new_n332_ );
and g162 ( new_n334_, new_n333_, new_n325_ );
and g163 ( new_n335_, new_n332_, keyIn_0_35 );
or g164 ( new_n336_, new_n334_, new_n335_ );
and g165 ( new_n337_, new_n324_, new_n314_, new_n336_ );
not g166 ( new_n338_, new_n336_ );
or g167 ( new_n339_, new_n323_, new_n338_ );
and g168 ( new_n340_, new_n339_, keyIn_0_62 );
or g169 ( new_n341_, new_n340_, new_n337_ );
and g170 ( new_n342_, new_n293_, new_n341_, new_n313_ );
not g171 ( new_n343_, keyIn_0_45 );
and g172 ( new_n344_, new_n194_, new_n188_ );
not g173 ( new_n345_, new_n344_ );
or g174 ( new_n346_, new_n273_, new_n345_ );
and g175 ( new_n347_, new_n345_, new_n268_ );
not g176 ( new_n348_, new_n347_ );
and g177 ( new_n349_, new_n346_, new_n343_, new_n348_ );
not g178 ( new_n350_, new_n349_ );
and g179 ( new_n351_, new_n346_, new_n348_ );
or g180 ( new_n352_, new_n351_, new_n343_ );
and g181 ( new_n353_, new_n352_, new_n350_ );
not g182 ( new_n354_, new_n353_ );
not g183 ( new_n355_, keyIn_0_33 );
not g184 ( new_n356_, N99 );
and g185 ( new_n357_, new_n356_, N95 );
and g186 ( new_n358_, new_n357_, new_n355_ );
not g187 ( new_n359_, new_n358_ );
or g188 ( new_n360_, new_n357_, new_n355_ );
and g189 ( new_n361_, new_n359_, new_n360_ );
not g190 ( new_n362_, new_n361_ );
and g191 ( new_n363_, new_n354_, keyIn_0_61, new_n362_ );
not g192 ( new_n364_, keyIn_0_61 );
or g193 ( new_n365_, new_n353_, new_n361_ );
and g194 ( new_n366_, new_n365_, new_n364_ );
or g195 ( new_n367_, new_n366_, new_n363_ );
not g196 ( new_n368_, keyIn_0_60 );
not g197 ( new_n369_, new_n273_ );
and g198 ( new_n370_, new_n369_, new_n225_ );
not g199 ( new_n371_, new_n225_ );
and g200 ( new_n372_, new_n273_, new_n371_ );
or g201 ( new_n373_, new_n370_, new_n372_ );
not g202 ( new_n374_, keyIn_0_31 );
not g203 ( new_n375_, N86 );
and g204 ( new_n376_, keyIn_0_10, N82 );
not g205 ( new_n377_, new_n376_ );
or g206 ( new_n378_, keyIn_0_10, N82 );
and g207 ( new_n379_, new_n377_, new_n378_ );
not g208 ( new_n380_, new_n379_ );
and g209 ( new_n381_, new_n380_, new_n375_ );
not g210 ( new_n382_, new_n381_ );
and g211 ( new_n383_, new_n382_, new_n374_ );
and g212 ( new_n384_, new_n381_, keyIn_0_31 );
or g213 ( new_n385_, new_n383_, new_n384_ );
and g214 ( new_n386_, new_n373_, new_n385_ );
not g215 ( new_n387_, new_n386_ );
or g216 ( new_n388_, new_n387_, new_n368_ );
or g217 ( new_n389_, new_n386_, keyIn_0_60 );
and g218 ( new_n390_, new_n388_, new_n389_ );
not g219 ( new_n391_, keyIn_0_54 );
and g220 ( new_n392_, new_n242_, new_n245_ );
not g221 ( new_n393_, new_n392_ );
and g222 ( new_n394_, new_n273_, new_n393_ );
and g223 ( new_n395_, new_n369_, new_n392_ );
or g224 ( new_n396_, new_n395_, new_n394_ );
not g225 ( new_n397_, N8 );
and g226 ( new_n398_, keyIn_0_1, N4 );
not g227 ( new_n399_, new_n398_ );
or g228 ( new_n400_, keyIn_0_1, N4 );
and g229 ( new_n401_, new_n399_, new_n400_ );
not g230 ( new_n402_, new_n401_ );
and g231 ( new_n403_, new_n402_, new_n397_ );
not g232 ( new_n404_, new_n403_ );
and g233 ( new_n405_, new_n404_, keyIn_0_15 );
not g234 ( new_n406_, new_n405_ );
or g235 ( new_n407_, new_n404_, keyIn_0_15 );
and g236 ( new_n408_, new_n406_, new_n407_ );
not g237 ( new_n409_, new_n408_ );
and g238 ( new_n410_, new_n396_, new_n409_ );
or g239 ( new_n411_, new_n410_, new_n391_ );
not g240 ( new_n412_, new_n396_ );
or g241 ( new_n413_, new_n412_, keyIn_0_54, new_n408_ );
and g242 ( new_n414_, new_n411_, new_n413_ );
not g243 ( new_n415_, keyIn_0_42 );
not g244 ( new_n416_, new_n206_ );
or g245 ( new_n417_, new_n273_, new_n416_ );
and g246 ( new_n418_, new_n273_, new_n416_ );
not g247 ( new_n419_, new_n418_ );
and g248 ( new_n420_, new_n419_, new_n417_ );
or g249 ( new_n421_, new_n420_, new_n415_ );
and g250 ( new_n422_, new_n420_, new_n415_ );
not g251 ( new_n423_, new_n422_ );
and g252 ( new_n424_, new_n423_, new_n421_ );
not g253 ( new_n425_, N60 );
and g254 ( new_n426_, keyIn_0_8, N56 );
not g255 ( new_n427_, new_n426_ );
or g256 ( new_n428_, keyIn_0_8, N56 );
and g257 ( new_n429_, new_n427_, new_n428_ );
not g258 ( new_n430_, new_n429_ );
and g259 ( new_n431_, new_n430_, new_n425_ );
not g260 ( new_n432_, new_n431_ );
and g261 ( new_n433_, new_n432_, keyIn_0_27 );
not g262 ( new_n434_, new_n433_ );
or g263 ( new_n435_, new_n432_, keyIn_0_27 );
and g264 ( new_n436_, new_n434_, new_n435_ );
or g265 ( new_n437_, new_n424_, new_n436_ );
and g266 ( new_n438_, new_n390_, new_n414_, new_n437_ );
and g267 ( new_n439_, new_n367_, new_n438_ );
not g268 ( new_n440_, keyIn_0_56 );
not g269 ( new_n441_, new_n231_ );
or g270 ( new_n442_, new_n273_, new_n441_ );
and g271 ( new_n443_, new_n269_, new_n272_, new_n441_ );
not g272 ( new_n444_, new_n443_ );
and g273 ( new_n445_, new_n442_, keyIn_0_39, new_n444_ );
not g274 ( new_n446_, new_n445_ );
and g275 ( new_n447_, new_n442_, new_n444_ );
or g276 ( new_n448_, new_n447_, keyIn_0_39 );
and g277 ( new_n449_, new_n448_, new_n446_ );
not g278 ( new_n450_, new_n449_ );
not g279 ( new_n451_, N21 );
and g280 ( new_n452_, new_n226_, keyIn_0_3 );
not g281 ( new_n453_, new_n452_ );
or g282 ( new_n454_, new_n226_, keyIn_0_3 );
and g283 ( new_n455_, new_n453_, new_n454_ );
not g284 ( new_n456_, new_n455_ );
and g285 ( new_n457_, new_n456_, new_n451_ );
not g286 ( new_n458_, new_n457_ );
and g287 ( new_n459_, new_n458_, keyIn_0_22 );
not g288 ( new_n460_, new_n459_ );
or g289 ( new_n461_, new_n458_, keyIn_0_22 );
and g290 ( new_n462_, new_n460_, new_n461_ );
not g291 ( new_n463_, new_n462_ );
and g292 ( new_n464_, new_n450_, new_n440_, new_n463_ );
or g293 ( new_n465_, new_n449_, new_n462_ );
and g294 ( new_n466_, new_n465_, keyIn_0_56 );
or g295 ( new_n467_, new_n466_, new_n464_ );
not g296 ( new_n468_, keyIn_0_40 );
not g297 ( new_n469_, new_n257_ );
or g298 ( new_n470_, new_n273_, new_n469_ );
or g299 ( new_n471_, new_n257_, keyIn_0_37 );
and g300 ( new_n472_, new_n470_, new_n471_ );
or g301 ( new_n473_, new_n472_, new_n468_ );
and g302 ( new_n474_, new_n472_, new_n468_ );
not g303 ( new_n475_, new_n474_ );
not g304 ( new_n476_, N34 );
and g305 ( new_n477_, new_n247_, keyIn_0_5 );
not g306 ( new_n478_, new_n477_ );
or g307 ( new_n479_, new_n247_, keyIn_0_5 );
and g308 ( new_n480_, new_n478_, new_n479_ );
not g309 ( new_n481_, new_n480_ );
and g310 ( new_n482_, new_n481_, new_n476_ );
not g311 ( new_n483_, new_n482_ );
and g312 ( new_n484_, new_n483_, keyIn_0_23 );
not g313 ( new_n485_, keyIn_0_23 );
and g314 ( new_n486_, new_n482_, new_n485_ );
or g315 ( new_n487_, new_n484_, new_n486_ );
and g316 ( new_n488_, new_n475_, new_n473_, new_n487_ );
and g317 ( new_n489_, new_n488_, keyIn_0_57 );
not g318 ( new_n490_, keyIn_0_57 );
not g319 ( new_n491_, new_n488_ );
and g320 ( new_n492_, new_n491_, new_n490_ );
or g321 ( new_n493_, new_n492_, new_n489_ );
and g322 ( new_n494_, new_n467_, new_n493_ );
and g323 ( new_n495_, new_n342_, new_n439_, new_n494_ );
or g324 ( new_n496_, new_n495_, keyIn_0_71 );
and g325 ( new_n497_, new_n342_, keyIn_0_71, new_n439_, new_n494_ );
not g326 ( new_n498_, new_n497_ );
and g327 ( new_n499_, new_n496_, new_n498_ );
not g328 ( new_n500_, new_n499_ );
and g329 ( new_n501_, new_n500_, new_n265_ );
and g330 ( new_n502_, new_n499_, keyIn_0_80 );
or g331 ( N329, new_n501_, new_n502_ );
not g332 ( new_n504_, keyIn_0_95 );
not g333 ( new_n505_, new_n493_ );
not g334 ( new_n506_, keyIn_0_78 );
or g335 ( new_n507_, new_n499_, new_n506_ );
and g336 ( new_n508_, new_n496_, new_n506_, new_n498_ );
not g337 ( new_n509_, new_n508_ );
and g338 ( new_n510_, new_n507_, new_n509_ );
or g339 ( new_n511_, new_n510_, new_n505_ );
and g340 ( new_n512_, new_n507_, new_n505_, new_n509_ );
not g341 ( new_n513_, new_n512_ );
and g342 ( new_n514_, new_n511_, new_n513_ );
not g343 ( new_n515_, keyIn_0_73 );
not g344 ( new_n516_, keyIn_0_64 );
not g345 ( new_n517_, keyIn_0_24 );
or g346 ( new_n518_, new_n480_, N40 );
not g347 ( new_n519_, new_n518_ );
and g348 ( new_n520_, new_n519_, new_n517_ );
and g349 ( new_n521_, new_n518_, keyIn_0_24 );
or g350 ( new_n522_, new_n520_, new_n521_ );
and g351 ( new_n523_, new_n475_, new_n473_, new_n522_ );
and g352 ( new_n524_, new_n523_, new_n516_ );
not g353 ( new_n525_, new_n524_ );
or g354 ( new_n526_, new_n523_, new_n516_ );
and g355 ( new_n527_, new_n525_, new_n526_ );
and g356 ( new_n528_, new_n527_, new_n515_ );
not g357 ( new_n529_, new_n528_ );
or g358 ( new_n530_, new_n527_, new_n515_ );
and g359 ( new_n531_, new_n529_, new_n530_ );
or g360 ( new_n532_, new_n514_, new_n531_ );
and g361 ( new_n533_, new_n532_, new_n504_ );
not g362 ( new_n534_, new_n514_ );
not g363 ( new_n535_, new_n531_ );
and g364 ( new_n536_, new_n534_, keyIn_0_95, new_n535_ );
or g365 ( new_n537_, new_n533_, new_n536_ );
not g366 ( new_n538_, new_n313_ );
or g367 ( new_n539_, new_n510_, new_n538_ );
and g368 ( new_n540_, new_n507_, new_n538_, new_n509_ );
not g369 ( new_n541_, new_n540_ );
and g370 ( new_n542_, new_n539_, new_n541_ );
not g371 ( new_n543_, keyIn_0_65 );
not g372 ( new_n544_, N53 );
and g373 ( new_n545_, new_n544_, N43 );
or g374 ( new_n546_, new_n545_, keyIn_0_26 );
not g375 ( new_n547_, keyIn_0_26 );
or g376 ( new_n548_, new_n547_, new_n209_, N53 );
and g377 ( new_n549_, new_n302_, new_n300_, new_n546_, new_n548_ );
and g378 ( new_n550_, new_n549_, new_n543_ );
not g379 ( new_n551_, new_n550_ );
or g380 ( new_n552_, new_n549_, new_n543_ );
and g381 ( new_n553_, new_n551_, new_n552_ );
or g382 ( new_n554_, new_n542_, new_n553_ );
and g383 ( new_n555_, new_n554_, keyIn_0_96 );
not g384 ( new_n556_, keyIn_0_96 );
not g385 ( new_n557_, new_n542_ );
not g386 ( new_n558_, new_n553_ );
and g387 ( new_n559_, new_n557_, new_n556_, new_n558_ );
or g388 ( new_n560_, new_n555_, new_n559_ );
and g389 ( new_n561_, new_n537_, new_n560_ );
not g390 ( new_n562_, keyIn_0_86 );
not g391 ( new_n563_, new_n390_ );
or g392 ( new_n564_, new_n510_, new_n563_ );
and g393 ( new_n565_, new_n507_, new_n563_, new_n509_ );
not g394 ( new_n566_, new_n565_ );
and g395 ( new_n567_, new_n564_, new_n566_ );
or g396 ( new_n568_, new_n567_, new_n562_ );
and g397 ( new_n569_, new_n564_, new_n562_, new_n566_ );
not g398 ( new_n570_, new_n569_ );
and g399 ( new_n571_, new_n568_, new_n570_ );
not g400 ( new_n572_, new_n373_ );
not g401 ( new_n573_, keyIn_0_32 );
or g402 ( new_n574_, new_n379_, N92 );
and g403 ( new_n575_, new_n574_, new_n573_ );
not g404 ( new_n576_, new_n575_ );
or g405 ( new_n577_, new_n574_, new_n573_ );
and g406 ( new_n578_, new_n576_, new_n577_ );
or g407 ( new_n579_, new_n572_, new_n578_ );
and g408 ( new_n580_, new_n579_, keyIn_0_68 );
not g409 ( new_n581_, new_n580_ );
or g410 ( new_n582_, new_n579_, keyIn_0_68 );
and g411 ( new_n583_, new_n581_, new_n582_ );
not g412 ( new_n584_, new_n583_ );
or g413 ( new_n585_, new_n584_, keyIn_0_75 );
not g414 ( new_n586_, keyIn_0_75 );
or g415 ( new_n587_, new_n583_, new_n586_ );
and g416 ( new_n588_, new_n585_, new_n587_ );
or g417 ( new_n589_, new_n571_, new_n588_ );
not g418 ( new_n590_, new_n437_ );
or g419 ( new_n591_, new_n510_, new_n590_ );
and g420 ( new_n592_, new_n507_, new_n590_, new_n509_ );
not g421 ( new_n593_, new_n592_ );
and g422 ( new_n594_, new_n591_, new_n593_ );
or g423 ( new_n595_, new_n594_, keyIn_0_83 );
and g424 ( new_n596_, new_n591_, keyIn_0_83, new_n593_ );
not g425 ( new_n597_, new_n596_ );
and g426 ( new_n598_, new_n595_, new_n597_ );
not g427 ( new_n599_, keyIn_0_28 );
or g428 ( new_n600_, new_n429_, N66 );
and g429 ( new_n601_, new_n600_, new_n599_ );
not g430 ( new_n602_, new_n601_ );
or g431 ( new_n603_, new_n600_, new_n599_ );
and g432 ( new_n604_, new_n602_, new_n603_ );
or g433 ( new_n605_, new_n424_, new_n604_ );
not g434 ( new_n606_, new_n605_ );
or g435 ( new_n607_, new_n606_, keyIn_0_66 );
not g436 ( new_n608_, keyIn_0_66 );
or g437 ( new_n609_, new_n605_, new_n608_ );
and g438 ( new_n610_, new_n607_, new_n609_ );
or g439 ( new_n611_, new_n598_, new_n610_ );
and g440 ( new_n612_, new_n589_, new_n611_ );
not g441 ( new_n613_, new_n467_ );
or g442 ( new_n614_, new_n510_, new_n613_ );
and g443 ( new_n615_, new_n510_, new_n613_ );
not g444 ( new_n616_, new_n615_ );
and g445 ( new_n617_, new_n616_, new_n614_ );
or g446 ( new_n618_, new_n617_, keyIn_0_82 );
and g447 ( new_n619_, new_n617_, keyIn_0_82 );
not g448 ( new_n620_, new_n619_ );
or g449 ( new_n621_, new_n449_, N27, new_n455_ );
not g450 ( new_n622_, new_n621_ );
and g451 ( new_n623_, new_n622_, keyIn_0_63 );
not g452 ( new_n624_, new_n623_ );
or g453 ( new_n625_, new_n622_, keyIn_0_63 );
and g454 ( new_n626_, new_n624_, new_n625_ );
not g455 ( new_n627_, new_n626_ );
and g456 ( new_n628_, new_n620_, new_n618_, new_n627_ );
or g457 ( new_n629_, new_n628_, keyIn_0_94 );
not g458 ( new_n630_, keyIn_0_94 );
not g459 ( new_n631_, new_n618_ );
or g460 ( new_n632_, new_n631_, new_n619_, new_n630_, new_n626_ );
and g461 ( new_n633_, new_n561_, new_n612_, new_n629_, new_n632_ );
not g462 ( new_n634_, new_n414_ );
and g463 ( new_n635_, new_n507_, new_n634_, new_n509_ );
not g464 ( new_n636_, new_n635_ );
or g465 ( new_n637_, new_n510_, new_n634_ );
and g466 ( new_n638_, new_n637_, keyIn_0_81, new_n636_ );
not g467 ( new_n639_, new_n638_ );
and g468 ( new_n640_, new_n637_, new_n636_ );
or g469 ( new_n641_, new_n640_, keyIn_0_81 );
or g470 ( new_n642_, new_n401_, N14 );
and g471 ( new_n643_, new_n642_, keyIn_0_16 );
not g472 ( new_n644_, new_n643_ );
or g473 ( new_n645_, new_n642_, keyIn_0_16 );
and g474 ( new_n646_, new_n644_, new_n645_ );
or g475 ( new_n647_, new_n412_, new_n646_ );
and g476 ( new_n648_, new_n647_, keyIn_0_55 );
not g477 ( new_n649_, new_n648_ );
or g478 ( new_n650_, new_n647_, keyIn_0_55 );
and g479 ( new_n651_, new_n649_, new_n650_ );
not g480 ( new_n652_, new_n651_ );
and g481 ( new_n653_, new_n652_, keyIn_0_72 );
not g482 ( new_n654_, keyIn_0_72 );
and g483 ( new_n655_, new_n651_, new_n654_ );
or g484 ( new_n656_, new_n653_, new_n655_ );
and g485 ( new_n657_, new_n641_, new_n639_, new_n656_ );
and g486 ( new_n658_, new_n657_, keyIn_0_93 );
not g487 ( new_n659_, keyIn_0_93 );
not g488 ( new_n660_, new_n657_ );
and g489 ( new_n661_, new_n660_, new_n659_ );
or g490 ( new_n662_, new_n661_, new_n658_ );
not g491 ( new_n663_, keyIn_0_97 );
not g492 ( new_n664_, new_n293_ );
or g493 ( new_n665_, new_n510_, new_n664_ );
and g494 ( new_n666_, new_n507_, new_n664_, new_n509_ );
not g495 ( new_n667_, new_n666_ );
and g496 ( new_n668_, new_n665_, keyIn_0_85, new_n667_ );
not g497 ( new_n669_, new_n668_ );
and g498 ( new_n670_, new_n665_, new_n667_ );
or g499 ( new_n671_, new_n670_, keyIn_0_85 );
not g500 ( new_n672_, keyIn_0_67 );
not g501 ( new_n673_, N79 );
and g502 ( new_n674_, new_n673_, N69 );
and g503 ( new_n675_, new_n674_, keyIn_0_30 );
not g504 ( new_n676_, new_n675_ );
or g505 ( new_n677_, new_n674_, keyIn_0_30 );
and g506 ( new_n678_, new_n676_, new_n677_ );
or g507 ( new_n679_, new_n281_, new_n678_ );
and g508 ( new_n680_, new_n679_, new_n672_ );
not g509 ( new_n681_, new_n680_ );
or g510 ( new_n682_, new_n679_, new_n672_ );
and g511 ( new_n683_, new_n681_, new_n682_ );
not g512 ( new_n684_, new_n683_ );
and g513 ( new_n685_, new_n684_, keyIn_0_74 );
not g514 ( new_n686_, keyIn_0_74 );
and g515 ( new_n687_, new_n683_, new_n686_ );
or g516 ( new_n688_, new_n685_, new_n687_ );
and g517 ( new_n689_, new_n671_, new_n669_, new_n688_ );
and g518 ( new_n690_, new_n689_, new_n663_ );
not g519 ( new_n691_, new_n689_ );
and g520 ( new_n692_, new_n691_, keyIn_0_97 );
or g521 ( new_n693_, new_n692_, new_n690_ );
and g522 ( new_n694_, new_n662_, new_n693_ );
not g523 ( new_n695_, keyIn_0_88 );
not g524 ( new_n696_, new_n367_ );
or g525 ( new_n697_, new_n510_, new_n696_ );
and g526 ( new_n698_, new_n507_, new_n696_, new_n509_ );
not g527 ( new_n699_, new_n698_ );
and g528 ( new_n700_, new_n697_, new_n695_, new_n699_ );
not g529 ( new_n701_, new_n700_ );
and g530 ( new_n702_, new_n697_, new_n699_ );
or g531 ( new_n703_, new_n702_, new_n695_ );
and g532 ( new_n704_, new_n703_, new_n701_ );
not g533 ( new_n705_, new_n704_ );
not g534 ( new_n706_, N105 );
and g535 ( new_n707_, new_n706_, N95 );
and g536 ( new_n708_, new_n707_, keyIn_0_34 );
not g537 ( new_n709_, new_n708_ );
or g538 ( new_n710_, new_n707_, keyIn_0_34 );
and g539 ( new_n711_, new_n709_, new_n710_ );
or g540 ( new_n712_, new_n353_, new_n711_ );
and g541 ( new_n713_, new_n712_, keyIn_0_69 );
not g542 ( new_n714_, new_n713_ );
or g543 ( new_n715_, new_n712_, keyIn_0_69 );
and g544 ( new_n716_, new_n714_, new_n715_ );
not g545 ( new_n717_, new_n716_ );
and g546 ( new_n718_, new_n717_, keyIn_0_76 );
not g547 ( new_n719_, new_n718_ );
or g548 ( new_n720_, new_n717_, keyIn_0_76 );
and g549 ( new_n721_, new_n719_, new_n720_ );
not g550 ( new_n722_, new_n721_ );
and g551 ( new_n723_, new_n705_, keyIn_0_98, new_n722_ );
not g552 ( new_n724_, keyIn_0_98 );
or g553 ( new_n725_, new_n704_, new_n721_ );
and g554 ( new_n726_, new_n725_, new_n724_ );
or g555 ( new_n727_, new_n726_, new_n723_ );
not g556 ( new_n728_, keyIn_0_99 );
not g557 ( new_n729_, new_n341_ );
or g558 ( new_n730_, new_n510_, new_n729_ );
and g559 ( new_n731_, new_n507_, new_n729_, new_n509_ );
not g560 ( new_n732_, new_n731_ );
and g561 ( new_n733_, new_n730_, keyIn_0_90, new_n732_ );
not g562 ( new_n734_, new_n733_ );
and g563 ( new_n735_, new_n730_, new_n732_ );
or g564 ( new_n736_, new_n735_, keyIn_0_90 );
and g565 ( new_n737_, new_n736_, new_n734_ );
not g566 ( new_n738_, new_n737_ );
not g567 ( new_n739_, keyIn_0_70 );
or g568 ( new_n740_, new_n330_, N115 );
and g569 ( new_n741_, new_n740_, keyIn_0_36 );
not g570 ( new_n742_, new_n741_ );
or g571 ( new_n743_, new_n740_, keyIn_0_36 );
and g572 ( new_n744_, new_n742_, new_n743_ );
or g573 ( new_n745_, new_n323_, new_n744_ );
and g574 ( new_n746_, new_n745_, new_n739_ );
not g575 ( new_n747_, new_n746_ );
or g576 ( new_n748_, new_n745_, new_n739_ );
and g577 ( new_n749_, new_n747_, new_n748_ );
not g578 ( new_n750_, new_n749_ );
and g579 ( new_n751_, new_n750_, keyIn_0_77 );
not g580 ( new_n752_, new_n751_ );
or g581 ( new_n753_, new_n750_, keyIn_0_77 );
and g582 ( new_n754_, new_n752_, new_n753_ );
not g583 ( new_n755_, new_n754_ );
and g584 ( new_n756_, new_n738_, new_n728_, new_n755_ );
or g585 ( new_n757_, new_n737_, new_n754_ );
and g586 ( new_n758_, new_n757_, keyIn_0_99 );
or g587 ( new_n759_, new_n758_, new_n756_ );
and g588 ( new_n760_, new_n694_, new_n633_, new_n727_, new_n759_ );
not g589 ( N370, new_n760_ );
not g590 ( new_n762_, keyIn_0_115 );
not g591 ( new_n763_, keyIn_0_114 );
not g592 ( new_n764_, keyIn_0_107 );
not g593 ( new_n765_, keyIn_0_100 );
and g594 ( new_n766_, new_n727_, new_n759_ );
and g595 ( new_n767_, new_n766_, new_n765_, new_n633_, new_n694_ );
not g596 ( new_n768_, new_n767_ );
or g597 ( new_n769_, new_n760_, new_n765_ );
and g598 ( new_n770_, new_n769_, new_n768_, new_n764_, N92 );
not g599 ( new_n771_, new_n770_ );
and g600 ( new_n772_, new_n769_, N92, new_n768_ );
or g601 ( new_n773_, new_n772_, new_n764_ );
and g602 ( new_n774_, new_n773_, new_n771_ );
and g603 ( new_n775_, new_n500_, keyIn_0_79 );
not g604 ( new_n776_, keyIn_0_79 );
and g605 ( new_n777_, new_n499_, new_n776_ );
or g606 ( new_n778_, new_n775_, new_n777_ );
and g607 ( new_n779_, new_n778_, N86 );
and g608 ( new_n780_, new_n260_, N76 );
not g609 ( new_n781_, new_n780_ );
and g610 ( new_n782_, new_n781_, keyIn_0_51 );
not g611 ( new_n783_, new_n782_ );
or g612 ( new_n784_, new_n781_, keyIn_0_51 );
and g613 ( new_n785_, new_n783_, new_n784_ );
or g614 ( new_n786_, new_n779_, new_n220_, new_n785_ );
or g615 ( new_n787_, new_n774_, new_n786_ );
and g616 ( new_n788_, new_n787_, new_n763_ );
not g617 ( new_n789_, new_n774_ );
not g618 ( new_n790_, new_n786_ );
and g619 ( new_n791_, new_n789_, keyIn_0_114, new_n790_ );
or g620 ( new_n792_, new_n788_, new_n791_ );
and g621 ( new_n793_, new_n769_, new_n768_, keyIn_0_106, N79 );
not g622 ( new_n794_, new_n793_ );
and g623 ( new_n795_, new_n769_, N79, new_n768_ );
or g624 ( new_n796_, new_n795_, keyIn_0_106 );
and g625 ( new_n797_, new_n796_, new_n794_ );
not g626 ( new_n798_, N69 );
and g627 ( new_n799_, new_n778_, N73 );
not g628 ( new_n800_, new_n799_ );
and g629 ( new_n801_, new_n800_, keyIn_0_91 );
not g630 ( new_n802_, new_n801_ );
or g631 ( new_n803_, new_n800_, keyIn_0_91 );
and g632 ( new_n804_, new_n802_, new_n803_ );
and g633 ( new_n805_, new_n260_, N63 );
not g634 ( new_n806_, new_n805_ );
and g635 ( new_n807_, new_n806_, keyIn_0_50 );
not g636 ( new_n808_, new_n807_ );
or g637 ( new_n809_, new_n806_, keyIn_0_50 );
and g638 ( new_n810_, new_n808_, new_n809_ );
or g639 ( new_n811_, new_n804_, new_n798_, new_n810_ );
or g640 ( new_n812_, new_n797_, new_n811_ );
and g641 ( new_n813_, new_n812_, keyIn_0_113 );
not g642 ( new_n814_, new_n813_ );
not g643 ( new_n815_, keyIn_0_113 );
not g644 ( new_n816_, new_n797_ );
not g645 ( new_n817_, new_n811_ );
and g646 ( new_n818_, new_n816_, new_n815_, new_n817_ );
not g647 ( new_n819_, new_n818_ );
and g648 ( new_n820_, new_n769_, N105, new_n768_ );
and g649 ( new_n821_, new_n820_, keyIn_0_108 );
not g650 ( new_n822_, new_n821_ );
or g651 ( new_n823_, new_n820_, keyIn_0_108 );
and g652 ( new_n824_, new_n822_, new_n823_ );
not g653 ( new_n825_, keyIn_0_92 );
and g654 ( new_n826_, new_n778_, N99 );
not g655 ( new_n827_, new_n826_ );
and g656 ( new_n828_, new_n827_, new_n825_ );
and g657 ( new_n829_, new_n826_, keyIn_0_92 );
not g658 ( new_n830_, keyIn_0_52 );
and g659 ( new_n831_, new_n260_, N89 );
not g660 ( new_n832_, new_n831_ );
and g661 ( new_n833_, new_n832_, new_n830_ );
and g662 ( new_n834_, new_n831_, keyIn_0_52 );
or g663 ( new_n835_, new_n833_, new_n834_ );
not g664 ( new_n836_, new_n835_ );
or g665 ( new_n837_, new_n828_, new_n829_, new_n182_, new_n836_ );
or g666 ( new_n838_, new_n824_, new_n837_ );
and g667 ( new_n839_, new_n769_, new_n768_ );
and g668 ( new_n840_, new_n839_, N115 );
and g669 ( new_n841_, new_n778_, N112 );
not g670 ( new_n842_, keyIn_0_53 );
and g671 ( new_n843_, new_n260_, N102 );
not g672 ( new_n844_, new_n843_ );
and g673 ( new_n845_, new_n844_, new_n842_ );
and g674 ( new_n846_, new_n843_, keyIn_0_53 );
or g675 ( new_n847_, new_n845_, new_n846_ );
not g676 ( new_n848_, new_n847_ );
or g677 ( new_n849_, new_n840_, new_n178_, new_n841_, new_n848_ );
and g678 ( new_n850_, new_n838_, new_n849_ );
and g679 ( new_n851_, new_n792_, new_n814_, new_n819_, new_n850_ );
not g680 ( new_n852_, keyIn_0_105 );
and g681 ( new_n853_, new_n769_, N66, new_n768_ );
or g682 ( new_n854_, new_n853_, new_n852_ );
not g683 ( new_n855_, new_n854_ );
and g684 ( new_n856_, new_n853_, new_n852_ );
and g685 ( new_n857_, new_n778_, N60 );
not g686 ( new_n858_, new_n857_ );
and g687 ( new_n859_, new_n858_, keyIn_0_89 );
not g688 ( new_n860_, new_n859_ );
or g689 ( new_n861_, new_n858_, keyIn_0_89 );
and g690 ( new_n862_, new_n860_, new_n861_ );
and g691 ( new_n863_, new_n260_, N50 );
and g692 ( new_n864_, new_n863_, keyIn_0_49 );
or g693 ( new_n865_, new_n863_, keyIn_0_49 );
not g694 ( new_n866_, new_n865_ );
or g695 ( new_n867_, new_n862_, new_n200_, new_n864_, new_n866_ );
or g696 ( new_n868_, new_n855_, new_n856_, keyIn_0_112, new_n867_ );
not g697 ( new_n869_, keyIn_0_112 );
not g698 ( new_n870_, new_n856_ );
not g699 ( new_n871_, new_n867_ );
and g700 ( new_n872_, new_n870_, new_n854_, new_n871_ );
or g701 ( new_n873_, new_n872_, new_n869_ );
and g702 ( new_n874_, new_n873_, new_n868_ );
and g703 ( new_n875_, new_n769_, N53, new_n768_ );
and g704 ( new_n876_, new_n875_, keyIn_0_104 );
not g705 ( new_n877_, new_n876_ );
or g706 ( new_n878_, new_n875_, keyIn_0_104 );
and g707 ( new_n879_, new_n877_, new_n878_ );
not g708 ( new_n880_, keyIn_0_87 );
and g709 ( new_n881_, new_n778_, N47 );
not g710 ( new_n882_, new_n881_ );
and g711 ( new_n883_, new_n882_, new_n880_ );
and g712 ( new_n884_, new_n881_, keyIn_0_87 );
not g713 ( new_n885_, keyIn_0_48 );
and g714 ( new_n886_, new_n260_, N37 );
and g715 ( new_n887_, new_n886_, new_n885_ );
not g716 ( new_n888_, new_n887_ );
or g717 ( new_n889_, new_n886_, new_n885_ );
and g718 ( new_n890_, new_n888_, N43, new_n889_ );
not g719 ( new_n891_, new_n890_ );
or g720 ( new_n892_, new_n883_, new_n884_, new_n891_ );
or g721 ( new_n893_, new_n879_, new_n892_ );
not g722 ( new_n894_, new_n893_ );
or g723 ( new_n895_, new_n874_, new_n894_ );
not g724 ( new_n896_, new_n895_ );
not g725 ( new_n897_, keyIn_0_110 );
not g726 ( new_n898_, keyIn_0_102 );
and g727 ( new_n899_, new_n839_, N27 );
and g728 ( new_n900_, new_n899_, new_n898_ );
not g729 ( new_n901_, new_n900_ );
or g730 ( new_n902_, new_n899_, new_n898_ );
and g731 ( new_n903_, new_n901_, new_n902_ );
not g732 ( new_n904_, keyIn_0_84 );
and g733 ( new_n905_, new_n778_, N21 );
and g734 ( new_n906_, new_n905_, new_n904_ );
or g735 ( new_n907_, new_n905_, new_n904_ );
not g736 ( new_n908_, new_n907_ );
and g737 ( new_n909_, new_n260_, N11 );
or g738 ( new_n910_, new_n908_, new_n226_, new_n906_, new_n909_ );
or g739 ( new_n911_, new_n903_, new_n910_ );
and g740 ( new_n912_, new_n911_, new_n897_ );
not g741 ( new_n913_, new_n912_ );
not g742 ( new_n914_, new_n903_ );
not g743 ( new_n915_, new_n910_ );
and g744 ( new_n916_, new_n914_, keyIn_0_110, new_n915_ );
not g745 ( new_n917_, new_n916_ );
not g746 ( new_n918_, keyIn_0_103 );
and g747 ( new_n919_, new_n769_, new_n768_, new_n918_, N40 );
not g748 ( new_n920_, new_n919_ );
and g749 ( new_n921_, new_n769_, N40, new_n768_ );
or g750 ( new_n922_, new_n921_, new_n918_ );
and g751 ( new_n923_, new_n922_, new_n920_ );
and g752 ( new_n924_, new_n778_, N34 );
not g753 ( new_n925_, keyIn_0_46 );
and g754 ( new_n926_, new_n260_, N24 );
and g755 ( new_n927_, new_n926_, new_n925_ );
or g756 ( new_n928_, new_n926_, new_n925_ );
not g757 ( new_n929_, new_n928_ );
or g758 ( new_n930_, new_n924_, new_n247_, new_n927_, new_n929_ );
or g759 ( new_n931_, new_n923_, new_n930_ );
and g760 ( new_n932_, new_n931_, keyIn_0_111 );
not g761 ( new_n933_, keyIn_0_111 );
not g762 ( new_n934_, new_n923_ );
not g763 ( new_n935_, new_n930_ );
and g764 ( new_n936_, new_n934_, new_n933_, new_n935_ );
or g765 ( new_n937_, new_n932_, new_n936_ );
not g766 ( new_n938_, new_n937_ );
and g767 ( new_n939_, new_n913_, new_n938_, new_n917_ );
and g768 ( new_n940_, new_n939_, new_n762_, new_n851_, new_n896_ );
not g769 ( new_n941_, new_n940_ );
and g770 ( new_n942_, new_n939_, new_n851_, new_n896_ );
or g771 ( new_n943_, new_n942_, new_n762_ );
and g772 ( new_n944_, new_n943_, new_n941_ );
not g773 ( new_n945_, keyIn_0_109 );
and g774 ( new_n946_, new_n839_, N14 );
or g775 ( new_n947_, new_n946_, keyIn_0_101 );
not g776 ( new_n948_, new_n947_ );
and g777 ( new_n949_, new_n946_, keyIn_0_101 );
and g778 ( new_n950_, new_n778_, N8 );
and g779 ( new_n951_, new_n260_, N1 );
and g780 ( new_n952_, new_n951_, keyIn_0_44 );
or g781 ( new_n953_, new_n951_, keyIn_0_44 );
not g782 ( new_n954_, new_n953_ );
or g783 ( new_n955_, new_n950_, new_n243_, new_n952_, new_n954_ );
or g784 ( new_n956_, new_n948_, new_n949_, new_n955_ );
not g785 ( new_n957_, new_n956_ );
and g786 ( new_n958_, new_n957_, new_n945_ );
and g787 ( new_n959_, new_n956_, keyIn_0_109 );
or g788 ( new_n960_, new_n958_, new_n959_ );
not g789 ( new_n961_, new_n960_ );
or g790 ( new_n962_, new_n944_, new_n961_ );
and g791 ( new_n963_, new_n962_, keyIn_0_120 );
not g792 ( new_n964_, keyIn_0_120 );
not g793 ( new_n965_, new_n944_ );
and g794 ( new_n966_, new_n965_, new_n964_, new_n960_ );
or g795 ( N421, new_n963_, new_n966_ );
not g796 ( new_n968_, keyIn_0_125 );
not g797 ( new_n969_, new_n874_ );
not g798 ( new_n970_, keyIn_0_121 );
not g799 ( new_n971_, keyIn_0_116 );
and g800 ( new_n972_, new_n894_, new_n971_ );
and g801 ( new_n973_, new_n893_, keyIn_0_116 );
or g802 ( new_n974_, new_n937_, new_n972_, new_n973_ );
or g803 ( new_n975_, new_n974_, new_n970_ );
not g804 ( new_n976_, new_n974_ );
or g805 ( new_n977_, new_n976_, keyIn_0_121 );
and g806 ( new_n978_, new_n977_, new_n975_, new_n969_, new_n939_ );
not g807 ( new_n979_, new_n978_ );
and g808 ( new_n980_, new_n979_, new_n968_ );
and g809 ( new_n981_, new_n978_, keyIn_0_125 );
or g810 ( N430, new_n980_, new_n981_ );
not g811 ( new_n983_, keyIn_0_123 );
not g812 ( new_n984_, new_n788_ );
not g813 ( new_n985_, new_n791_ );
and g814 ( new_n986_, new_n984_, keyIn_0_118, new_n985_ );
not g815 ( new_n987_, keyIn_0_118 );
and g816 ( new_n988_, new_n792_, new_n987_ );
or g817 ( new_n989_, new_n988_, new_n895_, new_n986_ );
and g818 ( new_n990_, new_n989_, new_n983_ );
not g819 ( new_n991_, new_n986_ );
not g820 ( new_n992_, new_n988_ );
and g821 ( new_n993_, new_n992_, keyIn_0_123, new_n896_, new_n991_ );
or g822 ( new_n994_, new_n990_, new_n993_ );
not g823 ( new_n995_, keyIn_0_122 );
and g824 ( new_n996_, new_n814_, keyIn_0_117, new_n819_ );
not g825 ( new_n997_, keyIn_0_117 );
or g826 ( new_n998_, new_n813_, new_n818_ );
and g827 ( new_n999_, new_n998_, new_n997_ );
or g828 ( new_n1000_, new_n999_, new_n996_ );
or g829 ( new_n1001_, new_n932_, new_n894_, new_n936_ );
not g830 ( new_n1002_, new_n1001_ );
and g831 ( new_n1003_, new_n1002_, new_n969_ );
and g832 ( new_n1004_, new_n1000_, new_n995_, new_n1003_ );
not g833 ( new_n1005_, new_n1004_ );
and g834 ( new_n1006_, new_n1000_, new_n1003_ );
or g835 ( new_n1007_, new_n1006_, new_n995_ );
and g836 ( new_n1008_, new_n994_, new_n939_, new_n1005_, new_n1007_ );
not g837 ( new_n1009_, new_n1008_ );
and g838 ( new_n1010_, new_n1009_, keyIn_0_126 );
not g839 ( new_n1011_, keyIn_0_126 );
and g840 ( new_n1012_, new_n1008_, new_n1011_ );
or g841 ( N431, new_n1010_, new_n1012_ );
not g842 ( new_n1014_, keyIn_0_127 );
and g843 ( new_n1015_, new_n977_, new_n975_, new_n913_, new_n917_ );
not g844 ( new_n1016_, keyIn_0_119 );
and g845 ( new_n1017_, new_n838_, new_n1016_ );
not g846 ( new_n1018_, new_n1017_ );
or g847 ( new_n1019_, new_n838_, new_n1016_ );
and g848 ( new_n1020_, new_n1018_, new_n1019_ );
not g849 ( new_n1021_, new_n1020_ );
and g850 ( new_n1022_, new_n1021_, keyIn_0_124, new_n792_, new_n1002_ );
not g851 ( new_n1023_, keyIn_0_124 );
not g852 ( new_n1024_, new_n792_ );
or g853 ( new_n1025_, new_n1020_, new_n1024_, new_n1001_ );
and g854 ( new_n1026_, new_n1025_, new_n1023_ );
or g855 ( new_n1027_, new_n1026_, new_n1022_ );
and g856 ( new_n1028_, new_n1015_, new_n1027_, new_n1007_, new_n1005_ );
and g857 ( new_n1029_, new_n1028_, new_n1014_ );
not g858 ( new_n1030_, new_n1028_ );
and g859 ( new_n1031_, new_n1030_, keyIn_0_127 );
or g860 ( N432, new_n1031_, new_n1029_ );
endmodule