module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n266_, new_n667_, new_n367_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n761_, new_n564_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n629_, new_n702_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n363_, new_n165_, new_n441_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n543_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n273_, new_n224_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n237_, new_n858_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n826_, new_n837_, new_n801_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n531_, new_n593_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n769_, new_n651_, new_n433_, new_n435_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n412_, new_n607_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n627_, new_n704_, new_n195_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n138_, N1 );
not g001 ( new_n139_, keyIn_0_17 );
not g002 ( new_n140_, keyIn_0_2 );
not g003 ( new_n141_, N33 );
not g004 ( new_n142_, N37 );
nand g005 ( new_n143_, new_n141_, new_n142_ );
nand g006 ( new_n144_, N33, N37 );
nand g007 ( new_n145_, new_n143_, new_n144_ );
nand g008 ( new_n146_, new_n145_, new_n140_ );
nand g009 ( new_n147_, new_n143_, keyIn_0_2, new_n144_ );
nand g010 ( new_n148_, new_n146_, new_n147_ );
not g011 ( new_n149_, N41 );
not g012 ( new_n150_, N45 );
nand g013 ( new_n151_, new_n149_, new_n150_ );
nand g014 ( new_n152_, N41, N45 );
nand g015 ( new_n153_, new_n151_, new_n152_ );
nand g016 ( new_n154_, new_n153_, keyIn_0_3 );
not g017 ( new_n155_, keyIn_0_3 );
nand g018 ( new_n156_, new_n151_, new_n155_, new_n152_ );
nand g019 ( new_n157_, new_n154_, new_n156_ );
nand g020 ( new_n158_, new_n148_, new_n157_ );
nand g021 ( new_n159_, new_n146_, new_n154_, new_n147_, new_n156_ );
nand g022 ( new_n160_, new_n158_, new_n159_ );
nand g023 ( new_n161_, new_n160_, new_n139_ );
nand g024 ( new_n162_, new_n158_, keyIn_0_17, new_n159_ );
nand g025 ( new_n163_, new_n161_, new_n162_ );
not g026 ( new_n164_, N49 );
not g027 ( new_n165_, N53 );
nand g028 ( new_n166_, new_n164_, new_n165_ );
nand g029 ( new_n167_, N49, N53 );
nand g030 ( new_n168_, new_n166_, new_n167_ );
nand g031 ( new_n169_, new_n168_, keyIn_0_4 );
not g032 ( new_n170_, keyIn_0_4 );
nand g033 ( new_n171_, new_n166_, new_n170_, new_n167_ );
nand g034 ( new_n172_, new_n169_, new_n171_ );
not g035 ( new_n173_, N57 );
not g036 ( new_n174_, N61 );
nand g037 ( new_n175_, new_n173_, new_n174_ );
nand g038 ( new_n176_, N57, N61 );
nand g039 ( new_n177_, new_n175_, new_n176_ );
nand g040 ( new_n178_, new_n172_, new_n177_ );
nand g041 ( new_n179_, new_n169_, new_n171_, new_n175_, new_n176_ );
nand g042 ( new_n180_, new_n178_, new_n179_ );
nand g043 ( new_n181_, new_n163_, new_n180_ );
nand g044 ( new_n182_, new_n161_, new_n162_, new_n178_, new_n179_ );
nand g045 ( new_n183_, new_n181_, new_n182_ );
nand g046 ( new_n184_, N134, N137 );
nand g047 ( new_n185_, new_n183_, new_n184_ );
nand g048 ( new_n186_, new_n181_, N134, N137, new_n182_ );
nand g049 ( new_n187_, new_n185_, new_n186_ );
not g050 ( new_n188_, N69 );
not g051 ( new_n189_, N85 );
nand g052 ( new_n190_, new_n188_, new_n189_ );
nand g053 ( new_n191_, N69, N85 );
nand g054 ( new_n192_, new_n190_, new_n191_ );
not g055 ( new_n193_, N101 );
not g056 ( new_n194_, N117 );
nand g057 ( new_n195_, new_n193_, new_n194_ );
nand g058 ( new_n196_, N101, N117 );
nand g059 ( new_n197_, new_n195_, new_n196_ );
nand g060 ( new_n198_, new_n192_, new_n197_ );
nand g061 ( new_n199_, new_n190_, new_n195_, new_n191_, new_n196_ );
nand g062 ( new_n200_, new_n198_, new_n199_ );
nand g063 ( new_n201_, new_n187_, new_n200_ );
nand g064 ( new_n202_, new_n185_, new_n186_, new_n198_, new_n199_ );
nand g065 ( new_n203_, new_n201_, new_n202_ );
not g066 ( new_n204_, N5 );
nand g067 ( new_n205_, new_n138_, new_n204_ );
nand g068 ( new_n206_, N1, N5 );
nand g069 ( new_n207_, new_n205_, new_n206_ );
not g070 ( new_n208_, N9 );
not g071 ( new_n209_, N13 );
nand g072 ( new_n210_, new_n208_, new_n209_ );
nand g073 ( new_n211_, N9, N13 );
nand g074 ( new_n212_, new_n210_, new_n211_ );
nand g075 ( new_n213_, new_n207_, new_n212_ );
nand g076 ( new_n214_, new_n205_, new_n210_, new_n206_, new_n211_ );
nand g077 ( new_n215_, new_n213_, new_n214_ );
nand g078 ( new_n216_, new_n215_, keyIn_0_16 );
not g079 ( new_n217_, keyIn_0_16 );
nand g080 ( new_n218_, new_n213_, new_n217_, new_n214_ );
nand g081 ( new_n219_, new_n216_, new_n218_ );
not g082 ( new_n220_, N25 );
not g083 ( new_n221_, N29 );
nand g084 ( new_n222_, new_n220_, new_n221_ );
nand g085 ( new_n223_, N25, N29 );
nand g086 ( new_n224_, new_n222_, new_n223_ );
nand g087 ( new_n225_, new_n224_, keyIn_0_1 );
not g088 ( new_n226_, keyIn_0_1 );
nand g089 ( new_n227_, new_n222_, new_n226_, new_n223_ );
nand g090 ( new_n228_, new_n225_, new_n227_ );
not g091 ( new_n229_, N21 );
nand g092 ( new_n230_, new_n229_, N17 );
not g093 ( new_n231_, N17 );
nand g094 ( new_n232_, new_n231_, N21 );
nand g095 ( new_n233_, new_n230_, new_n232_ );
nand g096 ( new_n234_, new_n233_, keyIn_0_0 );
not g097 ( new_n235_, keyIn_0_0 );
nand g098 ( new_n236_, new_n230_, new_n232_, new_n235_ );
nand g099 ( new_n237_, new_n234_, new_n236_ );
nand g100 ( new_n238_, new_n228_, new_n237_ );
nand g101 ( new_n239_, new_n225_, new_n234_, new_n227_, new_n236_ );
nand g102 ( new_n240_, new_n238_, new_n239_ );
nand g103 ( new_n241_, new_n219_, new_n240_ );
not g104 ( new_n242_, new_n219_ );
nand g105 ( new_n243_, new_n242_, new_n238_, new_n239_ );
nand g106 ( new_n244_, new_n243_, new_n241_ );
nand g107 ( new_n245_, N133, N137 );
nand g108 ( new_n246_, new_n244_, new_n245_ );
nand g109 ( new_n247_, new_n243_, N133, N137, new_n241_ );
nand g110 ( new_n248_, new_n246_, new_n247_ );
not g111 ( new_n249_, N113 );
nand g112 ( new_n250_, new_n249_, N97 );
not g113 ( new_n251_, N97 );
nand g114 ( new_n252_, new_n251_, N113 );
nand g115 ( new_n253_, new_n250_, new_n252_ );
nand g116 ( new_n254_, new_n253_, keyIn_0_15 );
not g117 ( new_n255_, keyIn_0_15 );
nand g118 ( new_n256_, new_n250_, new_n252_, new_n255_ );
nand g119 ( new_n257_, new_n254_, new_n256_ );
nand g120 ( new_n258_, N65, N81 );
not g121 ( new_n259_, new_n258_ );
nor g122 ( new_n260_, N65, N81 );
nor g123 ( new_n261_, new_n259_, new_n260_ );
nand g124 ( new_n262_, new_n257_, new_n261_ );
not g125 ( new_n263_, new_n261_ );
nand g126 ( new_n264_, new_n254_, new_n263_, new_n256_ );
nand g127 ( new_n265_, new_n262_, new_n264_ );
nand g128 ( new_n266_, new_n248_, new_n265_ );
nand g129 ( new_n267_, new_n246_, new_n247_, new_n262_, new_n264_ );
nand g130 ( new_n268_, new_n266_, new_n267_ );
not g131 ( new_n269_, new_n268_ );
nand g132 ( new_n270_, new_n203_, new_n269_ );
not g133 ( new_n271_, new_n270_ );
nand g134 ( new_n272_, new_n240_, new_n180_ );
nand g135 ( new_n273_, new_n238_, new_n178_, new_n179_, new_n239_ );
nand g136 ( new_n274_, new_n272_, new_n273_ );
nand g137 ( new_n275_, new_n274_, keyIn_0_11 );
not g138 ( new_n276_, keyIn_0_11 );
nand g139 ( new_n277_, new_n272_, new_n276_, new_n273_ );
nand g140 ( new_n278_, new_n275_, new_n277_ );
nand g141 ( new_n279_, N136, N137 );
nand g142 ( new_n280_, new_n278_, new_n279_ );
nand g143 ( new_n281_, new_n275_, N136, N137, new_n277_ );
nand g144 ( new_n282_, new_n280_, new_n281_ );
not g145 ( new_n283_, N77 );
not g146 ( new_n284_, N93 );
nand g147 ( new_n285_, new_n283_, new_n284_ );
nand g148 ( new_n286_, N77, N93 );
nand g149 ( new_n287_, new_n285_, new_n286_ );
not g150 ( new_n288_, N109 );
not g151 ( new_n289_, N125 );
nand g152 ( new_n290_, new_n288_, new_n289_ );
nand g153 ( new_n291_, N109, N125 );
nand g154 ( new_n292_, new_n290_, new_n291_ );
nand g155 ( new_n293_, new_n287_, new_n292_ );
nand g156 ( new_n294_, new_n285_, new_n290_, new_n286_, new_n291_ );
nand g157 ( new_n295_, new_n293_, new_n294_ );
not g158 ( new_n296_, new_n295_ );
nand g159 ( new_n297_, new_n282_, new_n296_ );
nand g160 ( new_n298_, new_n280_, new_n281_, new_n295_ );
nand g161 ( new_n299_, new_n297_, new_n298_ );
nand g162 ( new_n300_, new_n271_, new_n299_ );
not g163 ( new_n301_, new_n300_ );
not g164 ( new_n302_, N65 );
nand g165 ( new_n303_, new_n302_, new_n188_ );
nand g166 ( new_n304_, N65, N69 );
nand g167 ( new_n305_, new_n303_, new_n304_ );
nand g168 ( new_n306_, new_n305_, keyIn_0_5 );
not g169 ( new_n307_, keyIn_0_5 );
nand g170 ( new_n308_, new_n303_, new_n307_, new_n304_ );
nand g171 ( new_n309_, new_n306_, new_n308_ );
nand g172 ( new_n310_, new_n309_, keyIn_0_6 );
not g173 ( new_n311_, keyIn_0_6 );
nand g174 ( new_n312_, new_n306_, new_n311_, new_n308_ );
nand g175 ( new_n313_, new_n310_, new_n312_ );
nand g176 ( new_n314_, N73, N77 );
not g177 ( new_n315_, new_n314_ );
nor g178 ( new_n316_, N73, N77 );
nor g179 ( new_n317_, new_n315_, new_n316_ );
not g180 ( new_n318_, new_n317_ );
nand g181 ( new_n319_, new_n313_, new_n318_ );
nand g182 ( new_n320_, new_n310_, new_n312_, new_n317_ );
nand g183 ( new_n321_, new_n319_, new_n320_ );
not g184 ( new_n322_, N81 );
nand g185 ( new_n323_, new_n322_, new_n189_ );
nand g186 ( new_n324_, N81, N85 );
nand g187 ( new_n325_, new_n323_, new_n324_ );
not g188 ( new_n326_, N89 );
nand g189 ( new_n327_, new_n326_, new_n284_ );
nand g190 ( new_n328_, N89, N93 );
nand g191 ( new_n329_, new_n327_, new_n328_ );
nand g192 ( new_n330_, new_n325_, new_n329_ );
nand g193 ( new_n331_, new_n323_, new_n327_, new_n324_, new_n328_ );
nand g194 ( new_n332_, new_n330_, new_n331_ );
not g195 ( new_n333_, new_n332_ );
nand g196 ( new_n334_, new_n321_, new_n333_ );
nand g197 ( new_n335_, new_n319_, new_n320_, new_n332_ );
nand g198 ( new_n336_, N129, N137 );
nand g199 ( new_n337_, new_n334_, new_n335_, new_n336_ );
nand g200 ( new_n338_, new_n334_, new_n335_ );
nand g201 ( new_n339_, new_n338_, N129, N137 );
nand g202 ( new_n340_, new_n339_, new_n337_ );
nand g203 ( new_n341_, new_n138_, new_n231_ );
nand g204 ( new_n342_, N1, N17 );
nand g205 ( new_n343_, new_n341_, new_n342_ );
nand g206 ( new_n344_, new_n141_, new_n164_ );
nand g207 ( new_n345_, N33, N49 );
nand g208 ( new_n346_, new_n344_, new_n345_ );
nand g209 ( new_n347_, new_n343_, new_n346_ );
nand g210 ( new_n348_, new_n341_, new_n344_, new_n342_, new_n345_ );
nand g211 ( new_n349_, new_n347_, new_n348_ );
nand g212 ( new_n350_, new_n340_, new_n349_ );
nand g213 ( new_n351_, new_n339_, new_n337_, new_n347_, new_n348_ );
nand g214 ( new_n352_, new_n350_, new_n351_ );
not g215 ( new_n353_, new_n352_ );
not g216 ( new_n354_, keyIn_0_23 );
not g217 ( new_n355_, N121 );
nand g218 ( new_n356_, new_n355_, new_n289_ );
nand g219 ( new_n357_, N121, N125 );
nand g220 ( new_n358_, new_n356_, new_n357_ );
nand g221 ( new_n359_, new_n358_, keyIn_0_7 );
not g222 ( new_n360_, keyIn_0_7 );
nand g223 ( new_n361_, new_n356_, new_n360_, new_n357_ );
nand g224 ( new_n362_, new_n359_, new_n361_ );
nand g225 ( new_n363_, new_n249_, new_n194_ );
nand g226 ( new_n364_, N113, N117 );
nand g227 ( new_n365_, new_n363_, new_n364_ );
nand g228 ( new_n366_, new_n362_, new_n365_ );
nand g229 ( new_n367_, new_n359_, new_n361_, new_n363_, new_n364_ );
nand g230 ( new_n368_, new_n366_, new_n367_ );
nand g231 ( new_n369_, new_n368_, keyIn_0_19 );
not g232 ( new_n370_, keyIn_0_19 );
nand g233 ( new_n371_, new_n366_, new_n370_, new_n367_ );
nand g234 ( new_n372_, new_n369_, new_n371_ );
nand g235 ( new_n373_, new_n372_, new_n333_ );
nand g236 ( new_n374_, new_n369_, new_n332_, new_n371_ );
nand g237 ( new_n375_, new_n373_, new_n374_ );
nand g238 ( new_n376_, N132, N137 );
nand g239 ( new_n377_, new_n376_, keyIn_0_9 );
not g240 ( new_n378_, keyIn_0_9 );
nand g241 ( new_n379_, new_n378_, N132, N137 );
nand g242 ( new_n380_, new_n377_, new_n379_ );
nand g243 ( new_n381_, new_n375_, new_n380_ );
nand g244 ( new_n382_, new_n373_, new_n374_, new_n377_, new_n379_ );
nand g245 ( new_n383_, new_n381_, new_n382_ );
nand g246 ( new_n384_, new_n383_, new_n354_ );
nand g247 ( new_n385_, new_n381_, keyIn_0_23, new_n382_ );
nand g248 ( new_n386_, new_n384_, new_n385_ );
nor g249 ( new_n387_, N13, N29 );
not g250 ( new_n388_, new_n387_ );
nand g251 ( new_n389_, N13, N29 );
nand g252 ( new_n390_, new_n388_, new_n389_ );
nand g253 ( new_n391_, new_n390_, keyIn_0_14 );
not g254 ( new_n392_, new_n391_ );
nor g255 ( new_n393_, new_n390_, keyIn_0_14 );
nor g256 ( new_n394_, new_n392_, new_n393_ );
not g257 ( new_n395_, new_n394_ );
nand g258 ( new_n396_, N45, N61 );
not g259 ( new_n397_, new_n396_ );
nor g260 ( new_n398_, N45, N61 );
nor g261 ( new_n399_, new_n397_, new_n398_ );
not g262 ( new_n400_, new_n399_ );
nand g263 ( new_n401_, new_n395_, new_n400_ );
nand g264 ( new_n402_, new_n394_, new_n399_ );
nand g265 ( new_n403_, new_n401_, new_n402_ );
nand g266 ( new_n404_, new_n386_, new_n403_ );
nand g267 ( new_n405_, new_n384_, new_n385_, new_n401_, new_n402_ );
nand g268 ( new_n406_, new_n404_, new_n405_ );
nand g269 ( new_n407_, new_n193_, N97 );
nand g270 ( new_n408_, new_n251_, N101 );
nand g271 ( new_n409_, new_n407_, new_n408_ );
not g272 ( new_n410_, N105 );
nand g273 ( new_n411_, new_n410_, new_n288_ );
nand g274 ( new_n412_, N105, N109 );
nand g275 ( new_n413_, new_n411_, new_n412_ );
nand g276 ( new_n414_, new_n409_, new_n413_ );
nand g277 ( new_n415_, new_n411_, new_n407_, new_n408_, new_n412_ );
nand g278 ( new_n416_, new_n414_, new_n415_ );
nand g279 ( new_n417_, new_n416_, keyIn_0_18 );
not g280 ( new_n418_, keyIn_0_18 );
nand g281 ( new_n419_, new_n414_, new_n418_, new_n415_ );
nand g282 ( new_n420_, new_n417_, new_n419_ );
nand g283 ( new_n421_, new_n372_, new_n420_ );
not g284 ( new_n422_, new_n420_ );
nand g285 ( new_n423_, new_n369_, new_n422_, new_n371_ );
nand g286 ( new_n424_, new_n421_, new_n423_ );
nand g287 ( new_n425_, new_n424_, keyIn_0_22 );
not g288 ( new_n426_, keyIn_0_22 );
nand g289 ( new_n427_, new_n421_, new_n426_, new_n423_ );
nand g290 ( new_n428_, new_n425_, new_n427_ );
nand g291 ( new_n429_, new_n428_, keyIn_0_8 );
not g292 ( new_n430_, keyIn_0_8 );
nand g293 ( new_n431_, new_n425_, new_n430_, new_n427_ );
nand g294 ( new_n432_, new_n429_, new_n431_ );
nand g295 ( new_n433_, N130, N137 );
nand g296 ( new_n434_, new_n432_, new_n433_ );
nand g297 ( new_n435_, new_n429_, N130, N137, new_n431_ );
nand g298 ( new_n436_, new_n434_, new_n435_ );
nor g299 ( new_n437_, N5, N21 );
not g300 ( new_n438_, new_n437_ );
nand g301 ( new_n439_, N5, N21 );
nand g302 ( new_n440_, new_n438_, new_n439_ );
nand g303 ( new_n441_, new_n440_, keyIn_0_12 );
not g304 ( new_n442_, new_n441_ );
nor g305 ( new_n443_, new_n440_, keyIn_0_12 );
nor g306 ( new_n444_, new_n442_, new_n443_ );
not g307 ( new_n445_, new_n444_ );
nor g308 ( new_n446_, N37, N53 );
not g309 ( new_n447_, new_n446_ );
nand g310 ( new_n448_, N37, N53 );
nand g311 ( new_n449_, new_n447_, new_n448_ );
nand g312 ( new_n450_, new_n449_, keyIn_0_13 );
not g313 ( new_n451_, new_n450_ );
nor g314 ( new_n452_, new_n449_, keyIn_0_13 );
nor g315 ( new_n453_, new_n451_, new_n452_ );
not g316 ( new_n454_, new_n453_ );
nand g317 ( new_n455_, new_n445_, new_n454_ );
nand g318 ( new_n456_, new_n444_, new_n453_ );
nand g319 ( new_n457_, new_n455_, new_n456_ );
nand g320 ( new_n458_, new_n436_, new_n457_ );
nand g321 ( new_n459_, new_n434_, new_n435_, new_n455_, new_n456_ );
nand g322 ( new_n460_, new_n458_, new_n459_ );
not g323 ( new_n461_, new_n460_ );
nand g324 ( new_n462_, new_n321_, new_n420_ );
nand g325 ( new_n463_, new_n319_, new_n422_, new_n320_ );
nand g326 ( new_n464_, N131, N137 );
nand g327 ( new_n465_, new_n462_, new_n463_, new_n464_ );
nand g328 ( new_n466_, new_n462_, new_n463_ );
nand g329 ( new_n467_, new_n466_, N131, N137 );
nand g330 ( new_n468_, new_n467_, new_n465_ );
nand g331 ( new_n469_, new_n220_, N9 );
nand g332 ( new_n470_, new_n208_, N25 );
nand g333 ( new_n471_, new_n469_, new_n470_ );
nand g334 ( new_n472_, new_n149_, new_n173_ );
nand g335 ( new_n473_, N41, N57 );
nand g336 ( new_n474_, new_n472_, new_n473_ );
nand g337 ( new_n475_, new_n471_, new_n474_ );
nand g338 ( new_n476_, new_n472_, new_n469_, new_n470_, new_n473_ );
nand g339 ( new_n477_, new_n475_, new_n476_ );
nand g340 ( new_n478_, new_n468_, new_n477_ );
nand g341 ( new_n479_, new_n467_, new_n465_, new_n475_, new_n476_ );
nand g342 ( new_n480_, new_n478_, new_n479_ );
nand g343 ( new_n481_, new_n480_, keyIn_0_24 );
not g344 ( new_n482_, keyIn_0_24 );
nand g345 ( new_n483_, new_n478_, new_n482_, new_n479_ );
nand g346 ( new_n484_, new_n481_, new_n483_ );
not g347 ( new_n485_, new_n484_ );
nand g348 ( new_n486_, new_n461_, new_n352_, new_n485_ );
nand g349 ( new_n487_, new_n352_, keyIn_0_25 );
not g350 ( new_n488_, keyIn_0_25 );
nand g351 ( new_n489_, new_n353_, new_n488_ );
nand g352 ( new_n490_, new_n460_, new_n484_, new_n487_, new_n489_ );
nand g353 ( new_n491_, new_n486_, new_n490_ );
nand g354 ( new_n492_, new_n491_, new_n406_ );
not g355 ( new_n493_, new_n406_ );
nand g356 ( new_n494_, new_n460_, new_n352_, new_n493_, new_n485_ );
not g357 ( new_n495_, keyIn_0_36 );
not g358 ( new_n496_, keyIn_0_26 );
nand g359 ( new_n497_, new_n485_, new_n496_ );
nand g360 ( new_n498_, new_n484_, keyIn_0_26 );
nand g361 ( new_n499_, new_n497_, new_n498_ );
nand g362 ( new_n500_, new_n406_, new_n353_ );
not g363 ( new_n501_, new_n500_ );
nand g364 ( new_n502_, new_n499_, new_n460_, new_n501_ );
nand g365 ( new_n503_, new_n502_, new_n495_ );
nand g366 ( new_n504_, new_n499_, keyIn_0_36, new_n460_, new_n501_ );
nand g367 ( new_n505_, new_n503_, new_n504_ );
nand g368 ( new_n506_, new_n505_, new_n492_, new_n494_ );
not g369 ( new_n507_, keyIn_0_21 );
nand g370 ( new_n508_, new_n163_, new_n219_ );
nand g371 ( new_n509_, new_n161_, new_n162_, new_n242_ );
nand g372 ( new_n510_, new_n508_, new_n509_ );
nand g373 ( new_n511_, new_n510_, new_n507_ );
nand g374 ( new_n512_, new_n508_, keyIn_0_21, new_n509_ );
nand g375 ( new_n513_, new_n511_, new_n512_ );
nand g376 ( new_n514_, new_n513_, keyIn_0_10 );
not g377 ( new_n515_, keyIn_0_10 );
nand g378 ( new_n516_, new_n511_, new_n515_, new_n512_ );
nand g379 ( new_n517_, new_n514_, new_n516_ );
nand g380 ( new_n518_, N135, N137 );
nand g381 ( new_n519_, new_n517_, new_n518_ );
nand g382 ( new_n520_, new_n514_, N135, N137, new_n516_ );
nand g383 ( new_n521_, new_n519_, new_n520_ );
not g384 ( new_n522_, N73 );
nand g385 ( new_n523_, new_n522_, new_n326_ );
nand g386 ( new_n524_, N73, N89 );
nand g387 ( new_n525_, new_n523_, new_n524_ );
nand g388 ( new_n526_, new_n410_, new_n355_ );
nand g389 ( new_n527_, N105, N121 );
nand g390 ( new_n528_, new_n526_, new_n527_ );
nand g391 ( new_n529_, new_n525_, new_n528_ );
nand g392 ( new_n530_, new_n523_, new_n526_, new_n524_, new_n527_ );
nand g393 ( new_n531_, new_n529_, new_n530_ );
nand g394 ( new_n532_, new_n531_, keyIn_0_20 );
not g395 ( new_n533_, keyIn_0_20 );
nand g396 ( new_n534_, new_n529_, new_n533_, new_n530_ );
nand g397 ( new_n535_, new_n532_, new_n534_ );
not g398 ( new_n536_, new_n535_ );
nand g399 ( new_n537_, new_n521_, new_n536_ );
nand g400 ( new_n538_, new_n519_, new_n520_, new_n535_ );
nand g401 ( new_n539_, new_n537_, new_n538_ );
nand g402 ( new_n540_, new_n506_, new_n539_ );
not g403 ( new_n541_, new_n540_ );
nand g404 ( new_n542_, new_n541_, new_n301_, new_n353_ );
nand g405 ( new_n543_, new_n542_, keyIn_0_41 );
not g406 ( new_n544_, keyIn_0_41 );
nand g407 ( new_n545_, new_n541_, new_n544_, new_n301_, new_n353_ );
nand g408 ( new_n546_, new_n543_, new_n545_ );
nand g409 ( new_n547_, new_n546_, new_n138_ );
nand g410 ( new_n548_, new_n543_, N1, new_n545_ );
nand g411 ( N724, new_n547_, new_n548_ );
nand g412 ( new_n550_, new_n541_, new_n301_, new_n461_ );
nand g413 ( new_n551_, new_n550_, keyIn_0_42 );
not g414 ( new_n552_, keyIn_0_42 );
nand g415 ( new_n553_, new_n541_, new_n552_, new_n301_, new_n461_ );
nand g416 ( new_n554_, new_n551_, new_n553_ );
nand g417 ( new_n555_, new_n554_, N5 );
nand g418 ( new_n556_, new_n551_, new_n204_, new_n553_ );
nand g419 ( N725, new_n555_, new_n556_ );
nand g420 ( new_n558_, new_n541_, new_n301_ );
not g421 ( new_n559_, new_n558_ );
nand g422 ( new_n560_, new_n559_, new_n484_ );
nand g423 ( new_n561_, new_n560_, N9 );
nand g424 ( new_n562_, new_n559_, new_n208_, new_n484_ );
nand g425 ( N726, new_n561_, new_n562_ );
nand g426 ( new_n564_, new_n559_, new_n493_ );
nand g427 ( new_n565_, new_n564_, N13 );
nand g428 ( new_n566_, new_n559_, new_n209_, new_n493_ );
nand g429 ( N727, new_n565_, new_n566_ );
not g430 ( new_n568_, new_n299_ );
nand g431 ( new_n569_, new_n506_, new_n568_ );
not g432 ( new_n570_, new_n569_ );
not g433 ( new_n571_, new_n539_ );
nand g434 ( new_n572_, new_n571_, new_n271_ );
not g435 ( new_n573_, new_n572_ );
nand g436 ( new_n574_, new_n570_, new_n573_ );
not g437 ( new_n575_, new_n574_ );
nand g438 ( new_n576_, new_n575_, new_n353_ );
nand g439 ( new_n577_, new_n576_, N17 );
nand g440 ( new_n578_, new_n575_, new_n231_, new_n353_ );
nand g441 ( new_n579_, new_n577_, new_n578_ );
nand g442 ( new_n580_, new_n579_, keyIn_0_54 );
not g443 ( new_n581_, keyIn_0_54 );
nand g444 ( new_n582_, new_n577_, new_n581_, new_n578_ );
nand g445 ( N728, new_n580_, new_n582_ );
nand g446 ( new_n584_, new_n575_, new_n461_ );
nand g447 ( new_n585_, new_n584_, N21 );
nand g448 ( new_n586_, new_n575_, new_n229_, new_n461_ );
nand g449 ( new_n587_, new_n585_, new_n586_ );
nand g450 ( new_n588_, new_n587_, keyIn_0_55 );
not g451 ( new_n589_, keyIn_0_55 );
nand g452 ( new_n590_, new_n585_, new_n589_, new_n586_ );
nand g453 ( N729, new_n588_, new_n590_ );
nand g454 ( new_n592_, new_n575_, new_n484_ );
nand g455 ( new_n593_, new_n592_, N25 );
nand g456 ( new_n594_, new_n575_, new_n220_, new_n484_ );
nand g457 ( N730, new_n593_, new_n594_ );
not g458 ( new_n596_, keyIn_0_43 );
nand g459 ( new_n597_, new_n575_, new_n493_ );
nand g460 ( new_n598_, new_n597_, new_n596_ );
nand g461 ( new_n599_, new_n575_, keyIn_0_43, new_n493_ );
nand g462 ( new_n600_, new_n598_, new_n599_ );
nand g463 ( new_n601_, new_n600_, N29 );
nand g464 ( new_n602_, new_n598_, new_n221_, new_n599_ );
nand g465 ( N731, new_n601_, new_n602_ );
not g466 ( new_n604_, new_n203_ );
nand g467 ( new_n605_, new_n604_, new_n268_ );
nor g468 ( new_n606_, new_n605_, new_n568_ );
nand g469 ( new_n607_, new_n541_, new_n353_, new_n606_ );
nand g470 ( new_n608_, new_n607_, N33 );
nand g471 ( new_n609_, new_n541_, new_n141_, new_n353_, new_n606_ );
nand g472 ( new_n610_, new_n608_, new_n609_ );
nand g473 ( new_n611_, new_n610_, keyIn_0_56 );
not g474 ( new_n612_, keyIn_0_56 );
nand g475 ( new_n613_, new_n608_, new_n612_, new_n609_ );
nand g476 ( N732, new_n611_, new_n613_ );
nand g477 ( new_n615_, new_n541_, new_n461_, new_n606_ );
nand g478 ( new_n616_, new_n615_, new_n142_ );
nand g479 ( new_n617_, new_n541_, N37, new_n461_, new_n606_ );
nand g480 ( new_n618_, new_n616_, new_n617_ );
nand g481 ( new_n619_, new_n618_, keyIn_0_57 );
not g482 ( new_n620_, keyIn_0_57 );
nand g483 ( new_n621_, new_n616_, new_n620_, new_n617_ );
nand g484 ( N733, new_n619_, new_n621_ );
not g485 ( new_n623_, keyIn_0_44 );
nand g486 ( new_n624_, new_n606_, new_n484_ );
not g487 ( new_n625_, new_n624_ );
nand g488 ( new_n626_, new_n541_, new_n625_ );
nand g489 ( new_n627_, new_n626_, new_n623_ );
nand g490 ( new_n628_, new_n541_, keyIn_0_44, new_n625_ );
nand g491 ( new_n629_, new_n627_, new_n628_ );
nand g492 ( new_n630_, new_n629_, N41 );
nand g493 ( new_n631_, new_n627_, new_n149_, new_n628_ );
nand g494 ( N734, new_n630_, new_n631_ );
nor g495 ( new_n633_, new_n406_, new_n605_, new_n568_ );
nand g496 ( new_n634_, new_n541_, new_n633_ );
nand g497 ( new_n635_, new_n634_, keyIn_0_45 );
not g498 ( new_n636_, keyIn_0_45 );
nand g499 ( new_n637_, new_n541_, new_n636_, new_n633_ );
nand g500 ( new_n638_, new_n635_, new_n637_ );
nand g501 ( new_n639_, new_n638_, new_n150_ );
nand g502 ( new_n640_, new_n635_, N45, new_n637_ );
nand g503 ( new_n641_, new_n639_, new_n640_ );
nand g504 ( new_n642_, new_n641_, keyIn_0_58 );
not g505 ( new_n643_, keyIn_0_58 );
nand g506 ( new_n644_, new_n639_, new_n643_, new_n640_ );
nand g507 ( N735, new_n642_, new_n644_ );
not g508 ( new_n646_, keyIn_0_59 );
not g509 ( new_n647_, keyIn_0_39 );
nand g510 ( new_n648_, new_n571_, keyIn_0_27 );
not g511 ( new_n649_, keyIn_0_27 );
nand g512 ( new_n650_, new_n539_, new_n649_ );
nand g513 ( new_n651_, new_n648_, new_n604_, new_n268_, new_n650_ );
not g514 ( new_n652_, new_n651_ );
nand g515 ( new_n653_, new_n506_, new_n568_, new_n652_ );
nand g516 ( new_n654_, new_n653_, new_n647_ );
nand g517 ( new_n655_, new_n506_, keyIn_0_39, new_n568_, new_n652_ );
nand g518 ( new_n656_, new_n654_, new_n655_ );
nand g519 ( new_n657_, new_n656_, new_n353_ );
nand g520 ( new_n658_, new_n657_, new_n164_ );
nand g521 ( new_n659_, new_n656_, N49, new_n353_ );
nand g522 ( new_n660_, new_n658_, new_n659_ );
nand g523 ( new_n661_, new_n660_, new_n646_ );
nand g524 ( new_n662_, new_n658_, keyIn_0_59, new_n659_ );
nand g525 ( N736, new_n661_, new_n662_ );
not g526 ( new_n664_, keyIn_0_46 );
nand g527 ( new_n665_, new_n656_, new_n461_ );
nand g528 ( new_n666_, new_n665_, new_n664_ );
nand g529 ( new_n667_, new_n656_, keyIn_0_46, new_n461_ );
nand g530 ( new_n668_, new_n666_, new_n667_ );
nand g531 ( new_n669_, new_n668_, new_n165_ );
nand g532 ( new_n670_, new_n666_, N53, new_n667_ );
nand g533 ( N737, new_n669_, new_n670_ );
nand g534 ( new_n672_, new_n656_, new_n484_ );
nand g535 ( new_n673_, new_n672_, N57 );
nand g536 ( new_n674_, new_n656_, new_n173_, new_n484_ );
nand g537 ( N738, new_n673_, new_n674_ );
nand g538 ( new_n676_, new_n656_, new_n493_ );
nand g539 ( new_n677_, new_n676_, N61 );
nand g540 ( new_n678_, new_n656_, new_n174_, new_n493_ );
nand g541 ( N739, new_n677_, new_n678_ );
not g542 ( new_n680_, keyIn_0_47 );
not g543 ( new_n681_, keyIn_0_37 );
not g544 ( new_n682_, keyIn_0_31 );
nand g545 ( new_n683_, new_n537_, new_n682_, new_n538_ );
nand g546 ( new_n684_, new_n539_, keyIn_0_31 );
nand g547 ( new_n685_, new_n684_, new_n681_, new_n606_, new_n683_ );
not g548 ( new_n686_, keyIn_0_32 );
nand g549 ( new_n687_, new_n539_, new_n686_ );
nand g550 ( new_n688_, new_n537_, keyIn_0_32, new_n538_ );
nand g551 ( new_n689_, new_n687_, new_n688_ );
not g552 ( new_n690_, keyIn_0_33 );
nand g553 ( new_n691_, new_n568_, new_n690_ );
nand g554 ( new_n692_, new_n299_, keyIn_0_33 );
nand g555 ( new_n693_, new_n271_, new_n691_, new_n692_ );
not g556 ( new_n694_, new_n693_ );
nand g557 ( new_n695_, new_n689_, new_n694_ );
nand g558 ( new_n696_, new_n299_, keyIn_0_30 );
not g559 ( new_n697_, keyIn_0_30 );
nand g560 ( new_n698_, new_n297_, new_n697_, new_n298_ );
nand g561 ( new_n699_, new_n696_, new_n698_ );
not g562 ( new_n700_, keyIn_0_29 );
nand g563 ( new_n701_, new_n268_, new_n700_ );
nand g564 ( new_n702_, new_n266_, keyIn_0_29, new_n267_ );
nand g565 ( new_n703_, new_n701_, new_n702_ );
not g566 ( new_n704_, new_n703_ );
nand g567 ( new_n705_, new_n699_, new_n203_, new_n704_ );
not g568 ( new_n706_, new_n705_ );
nand g569 ( new_n707_, new_n706_, new_n539_ );
nand g570 ( new_n708_, new_n604_, keyIn_0_28 );
not g571 ( new_n709_, keyIn_0_28 );
nand g572 ( new_n710_, new_n203_, new_n709_ );
nand g573 ( new_n711_, new_n708_, new_n710_ );
nand g574 ( new_n712_, new_n568_, new_n268_ );
not g575 ( new_n713_, new_n712_ );
nand g576 ( new_n714_, new_n537_, new_n711_, new_n538_, new_n713_ );
nand g577 ( new_n715_, new_n707_, new_n714_ );
not g578 ( new_n716_, new_n715_ );
nand g579 ( new_n717_, new_n695_, new_n716_, new_n685_ );
not g580 ( new_n718_, new_n717_ );
not g581 ( new_n719_, keyIn_0_38 );
nand g582 ( new_n720_, new_n684_, new_n606_, new_n683_ );
nand g583 ( new_n721_, new_n720_, keyIn_0_37 );
nand g584 ( new_n722_, new_n721_, new_n719_ );
not g585 ( new_n723_, new_n722_ );
nand g586 ( new_n724_, new_n718_, new_n723_ );
nand g587 ( new_n725_, new_n721_, new_n695_, new_n685_, new_n716_ );
nand g588 ( new_n726_, new_n725_, keyIn_0_38 );
nand g589 ( new_n727_, new_n460_, new_n484_, new_n501_ );
not g590 ( new_n728_, new_n727_ );
nand g591 ( new_n729_, new_n724_, new_n726_, new_n728_ );
nand g592 ( new_n730_, new_n729_, keyIn_0_40 );
not g593 ( new_n731_, keyIn_0_40 );
nand g594 ( new_n732_, new_n724_, new_n731_, new_n726_, new_n728_ );
nand g595 ( new_n733_, new_n730_, new_n732_ );
nand g596 ( new_n734_, new_n733_, new_n269_ );
nand g597 ( new_n735_, new_n734_, new_n680_ );
nand g598 ( new_n736_, new_n733_, keyIn_0_47, new_n269_ );
nand g599 ( new_n737_, new_n735_, new_n736_ );
nand g600 ( new_n738_, new_n737_, N65 );
nand g601 ( new_n739_, new_n735_, new_n302_, new_n736_ );
nand g602 ( N740, new_n738_, new_n739_ );
not g603 ( new_n741_, keyIn_0_48 );
nand g604 ( new_n742_, new_n733_, new_n604_ );
nand g605 ( new_n743_, new_n742_, new_n741_ );
nand g606 ( new_n744_, new_n733_, keyIn_0_48, new_n604_ );
nand g607 ( new_n745_, new_n743_, new_n744_ );
nand g608 ( new_n746_, new_n745_, N69 );
nand g609 ( new_n747_, new_n743_, new_n188_, new_n744_ );
nand g610 ( N741, new_n746_, new_n747_ );
nand g611 ( new_n749_, new_n733_, new_n539_ );
nand g612 ( new_n750_, new_n749_, N73 );
nand g613 ( new_n751_, new_n733_, new_n522_, new_n539_ );
nand g614 ( N742, new_n750_, new_n751_ );
not g615 ( new_n753_, keyIn_0_60 );
nand g616 ( new_n754_, new_n733_, new_n568_ );
nand g617 ( new_n755_, new_n754_, new_n283_ );
nand g618 ( new_n756_, new_n733_, N77, new_n568_ );
nand g619 ( new_n757_, new_n755_, new_n756_ );
nand g620 ( new_n758_, new_n757_, new_n753_ );
nand g621 ( new_n759_, new_n755_, keyIn_0_60, new_n756_ );
nand g622 ( N743, new_n758_, new_n759_ );
nor g623 ( new_n761_, new_n717_, new_n722_ );
not g624 ( new_n762_, new_n726_ );
nor g625 ( new_n763_, new_n762_, new_n761_ );
not g626 ( new_n764_, keyIn_0_34 );
nand g627 ( new_n765_, new_n461_, new_n764_ );
nand g628 ( new_n766_, new_n460_, keyIn_0_34 );
nand g629 ( new_n767_, new_n765_, new_n766_ );
nand g630 ( new_n768_, new_n767_, new_n353_, new_n493_, new_n485_ );
not g631 ( new_n769_, new_n768_ );
nand g632 ( new_n770_, new_n763_, new_n769_ );
not g633 ( new_n771_, new_n770_ );
nand g634 ( new_n772_, new_n771_, new_n269_ );
nand g635 ( new_n773_, new_n772_, N81 );
nand g636 ( new_n774_, new_n771_, new_n322_, new_n269_ );
nand g637 ( N744, new_n773_, new_n774_ );
not g638 ( new_n776_, keyIn_0_49 );
nand g639 ( new_n777_, new_n763_, new_n604_, new_n769_ );
nand g640 ( new_n778_, new_n777_, new_n776_ );
nand g641 ( new_n779_, new_n763_, new_n604_ );
not g642 ( new_n780_, new_n779_ );
nand g643 ( new_n781_, new_n780_, keyIn_0_49, new_n769_ );
nand g644 ( new_n782_, new_n781_, new_n778_ );
nand g645 ( new_n783_, new_n782_, new_n189_ );
nand g646 ( new_n784_, new_n781_, N85, new_n778_ );
nand g647 ( N745, new_n783_, new_n784_ );
not g648 ( new_n786_, keyIn_0_61 );
nand g649 ( new_n787_, new_n763_, new_n539_, new_n769_ );
nand g650 ( new_n788_, new_n787_, new_n326_ );
nand g651 ( new_n789_, new_n763_, N89, new_n539_, new_n769_ );
nand g652 ( new_n790_, new_n788_, new_n789_ );
nand g653 ( new_n791_, new_n790_, new_n786_ );
nand g654 ( new_n792_, new_n788_, keyIn_0_61, new_n789_ );
nand g655 ( N746, new_n791_, new_n792_ );
nand g656 ( new_n794_, new_n771_, new_n568_ );
nand g657 ( new_n795_, new_n794_, N93 );
nand g658 ( new_n796_, new_n771_, new_n284_, new_n568_ );
nand g659 ( N747, new_n795_, new_n796_ );
nand g660 ( new_n798_, new_n353_, keyIn_0_35 );
not g661 ( new_n799_, keyIn_0_35 );
nand g662 ( new_n800_, new_n352_, new_n799_ );
nand g663 ( new_n801_, new_n798_, new_n800_ );
nand g664 ( new_n802_, new_n801_, new_n406_, new_n484_ );
nor g665 ( new_n803_, new_n802_, new_n460_ );
nand g666 ( new_n804_, new_n763_, new_n803_ );
not g667 ( new_n805_, new_n804_ );
nand g668 ( new_n806_, new_n805_, new_n269_ );
nand g669 ( new_n807_, new_n806_, N97 );
nand g670 ( new_n808_, new_n805_, new_n251_, new_n269_ );
nand g671 ( N748, new_n807_, new_n808_ );
nand g672 ( new_n810_, new_n763_, new_n604_, new_n803_ );
nand g673 ( new_n811_, new_n810_, keyIn_0_50 );
not g674 ( new_n812_, keyIn_0_50 );
nand g675 ( new_n813_, new_n780_, new_n812_, new_n803_ );
nand g676 ( new_n814_, new_n813_, new_n811_ );
nand g677 ( new_n815_, new_n814_, N101 );
nand g678 ( new_n816_, new_n813_, new_n193_, new_n811_ );
nand g679 ( N749, new_n815_, new_n816_ );
nand g680 ( new_n818_, new_n805_, new_n539_ );
nand g681 ( new_n819_, new_n818_, N105 );
nand g682 ( new_n820_, new_n805_, new_n410_, new_n539_ );
nand g683 ( N750, new_n819_, new_n820_ );
nand g684 ( new_n822_, new_n805_, new_n568_ );
nand g685 ( new_n823_, new_n822_, N109 );
nand g686 ( new_n824_, new_n805_, new_n288_, new_n568_ );
nand g687 ( N751, new_n823_, new_n824_ );
nand g688 ( new_n826_, new_n461_, new_n352_, new_n493_, new_n485_ );
not g689 ( new_n827_, new_n826_ );
nand g690 ( new_n828_, new_n763_, new_n827_ );
not g691 ( new_n829_, new_n828_ );
nand g692 ( new_n830_, new_n829_, new_n269_ );
nand g693 ( new_n831_, new_n830_, N113 );
nand g694 ( new_n832_, new_n829_, new_n249_, new_n269_ );
nand g695 ( N752, new_n831_, new_n832_ );
not g696 ( new_n834_, keyIn_0_51 );
nand g697 ( new_n835_, new_n763_, new_n604_, new_n827_ );
nand g698 ( new_n836_, new_n835_, new_n834_ );
nand g699 ( new_n837_, new_n780_, keyIn_0_51, new_n827_ );
nand g700 ( new_n838_, new_n837_, new_n836_ );
nand g701 ( new_n839_, new_n838_, N117 );
nand g702 ( new_n840_, new_n837_, new_n194_, new_n836_ );
nand g703 ( N753, new_n839_, new_n840_ );
nand g704 ( new_n842_, new_n724_, new_n539_, new_n726_, new_n827_ );
nand g705 ( new_n843_, new_n842_, keyIn_0_52 );
not g706 ( new_n844_, keyIn_0_52 );
nand g707 ( new_n845_, new_n763_, new_n844_, new_n539_, new_n827_ );
nand g708 ( new_n846_, new_n845_, new_n843_ );
nand g709 ( new_n847_, new_n846_, N121 );
nand g710 ( new_n848_, new_n845_, new_n355_, new_n843_ );
nand g711 ( new_n849_, new_n847_, new_n848_ );
nand g712 ( new_n850_, new_n849_, keyIn_0_62 );
not g713 ( new_n851_, keyIn_0_62 );
nand g714 ( new_n852_, new_n847_, new_n851_, new_n848_ );
nand g715 ( N754, new_n850_, new_n852_ );
not g716 ( new_n854_, keyIn_0_53 );
nand g717 ( new_n855_, new_n724_, new_n568_, new_n726_, new_n827_ );
nand g718 ( new_n856_, new_n855_, new_n854_ );
nand g719 ( new_n857_, new_n763_, keyIn_0_53, new_n568_, new_n827_ );
nand g720 ( new_n858_, new_n857_, new_n856_ );
nand g721 ( new_n859_, new_n858_, N125 );
nand g722 ( new_n860_, new_n857_, new_n289_, new_n856_ );
nand g723 ( new_n861_, new_n859_, new_n860_ );
nand g724 ( new_n862_, new_n861_, keyIn_0_63 );
not g725 ( new_n863_, keyIn_0_63 );
nand g726 ( new_n864_, new_n859_, new_n863_, new_n860_ );
nand g727 ( N755, new_n862_, new_n864_ );
endmodule