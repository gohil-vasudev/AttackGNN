module add_mul_combine_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_mul_0_, Result_mul_1_, 
        Result_mul_2_, Result_mul_3_, Result_mul_4_, Result_mul_5_, 
        Result_mul_6_, Result_mul_7_, Result_mul_8_, Result_mul_9_, 
        Result_mul_10_, Result_mul_11_, Result_mul_12_, Result_mul_13_, 
        Result_mul_14_, Result_mul_15_, Result_mul_16_, Result_mul_17_, 
        Result_mul_18_, Result_mul_19_, Result_mul_20_, Result_mul_21_, 
        Result_mul_22_, Result_mul_23_, Result_mul_24_, Result_mul_25_, 
        Result_mul_26_, Result_mul_27_, Result_mul_28_, Result_mul_29_, 
        Result_mul_30_, Result_mul_31_, Result_mul_32_, Result_mul_33_, 
        Result_mul_34_, Result_mul_35_, Result_mul_36_, Result_mul_37_, 
        Result_mul_38_, Result_mul_39_, Result_mul_40_, Result_mul_41_, 
        Result_mul_42_, Result_mul_43_, Result_mul_44_, Result_mul_45_, 
        Result_mul_46_, Result_mul_47_, Result_mul_48_, Result_mul_49_, 
        Result_mul_50_, Result_mul_51_, Result_mul_52_, Result_mul_53_, 
        Result_mul_54_, Result_mul_55_, Result_mul_56_, Result_mul_57_, 
        Result_mul_58_, Result_mul_59_, Result_mul_60_, Result_mul_61_, 
        Result_mul_62_, Result_mul_63_, Result_add_0_, Result_add_1_, 
        Result_add_2_, Result_add_3_, Result_add_4_, Result_add_5_, 
        Result_add_6_, Result_add_7_, Result_add_8_, Result_add_9_, 
        Result_add_10_, Result_add_11_, Result_add_12_, Result_add_13_, 
        Result_add_14_, Result_add_15_, Result_add_16_, Result_add_17_, 
        Result_add_18_, Result_add_19_, Result_add_20_, Result_add_21_, 
        Result_add_22_, Result_add_23_, Result_add_24_, Result_add_25_, 
        Result_add_26_, Result_add_27_, Result_add_28_, Result_add_29_, 
        Result_add_30_, Result_add_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_mul_0_, Result_mul_1_, Result_mul_2_, Result_mul_3_,
         Result_mul_4_, Result_mul_5_, Result_mul_6_, Result_mul_7_,
         Result_mul_8_, Result_mul_9_, Result_mul_10_, Result_mul_11_,
         Result_mul_12_, Result_mul_13_, Result_mul_14_, Result_mul_15_,
         Result_mul_16_, Result_mul_17_, Result_mul_18_, Result_mul_19_,
         Result_mul_20_, Result_mul_21_, Result_mul_22_, Result_mul_23_,
         Result_mul_24_, Result_mul_25_, Result_mul_26_, Result_mul_27_,
         Result_mul_28_, Result_mul_29_, Result_mul_30_, Result_mul_31_,
         Result_mul_32_, Result_mul_33_, Result_mul_34_, Result_mul_35_,
         Result_mul_36_, Result_mul_37_, Result_mul_38_, Result_mul_39_,
         Result_mul_40_, Result_mul_41_, Result_mul_42_, Result_mul_43_,
         Result_mul_44_, Result_mul_45_, Result_mul_46_, Result_mul_47_,
         Result_mul_48_, Result_mul_49_, Result_mul_50_, Result_mul_51_,
         Result_mul_52_, Result_mul_53_, Result_mul_54_, Result_mul_55_,
         Result_mul_56_, Result_mul_57_, Result_mul_58_, Result_mul_59_,
         Result_mul_60_, Result_mul_61_, Result_mul_62_, Result_mul_63_,
         Result_add_0_, Result_add_1_, Result_add_2_, Result_add_3_,
         Result_add_4_, Result_add_5_, Result_add_6_, Result_add_7_,
         Result_add_8_, Result_add_9_, Result_add_10_, Result_add_11_,
         Result_add_12_, Result_add_13_, Result_add_14_, Result_add_15_,
         Result_add_16_, Result_add_17_, Result_add_18_, Result_add_19_,
         Result_add_20_, Result_add_21_, Result_add_22_, Result_add_23_,
         Result_add_24_, Result_add_25_, Result_add_26_, Result_add_27_,
         Result_add_28_, Result_add_29_, Result_add_30_, Result_add_31_;
  wire   n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666;

  INV_X2 U7345 ( .A(b_27_), .ZN(n8183) );
  INV_X2 U7346 ( .A(b_7_), .ZN(n12673) );
  INV_X2 U7347 ( .A(b_16_), .ZN(n10683) );
  INV_X2 U7348 ( .A(b_22_), .ZN(n9312) );
  INV_X2 U7349 ( .A(b_30_), .ZN(n7274) );
  NAND2_X2 U7350 ( .A1(a_30_), .A2(n14290), .ZN(n7272) );
  NAND2_X2 U7351 ( .A1(a_31_), .A2(n14287), .ZN(n7268) );
  INV_X2 U7352 ( .A(a_15_), .ZN(n7346) );
  INV_X2 U7353 ( .A(a_9_), .ZN(n7870) );
  INV_X2 U7354 ( .A(a_20_), .ZN(n7987) );
  INV_X2 U7355 ( .A(a_25_), .ZN(n7923) );
  INV_X2 U7356 ( .A(a_18_), .ZN(n7764) );
  INV_X2 U7357 ( .A(a_24_), .ZN(n7691) );
  INV_X2 U7358 ( .A(a_23_), .ZN(n7916) );
  INV_X2 U7359 ( .A(a_17_), .ZN(n7337) );
  INV_X2 U7360 ( .A(a_21_), .ZN(n7909) );
  INV_X2 U7361 ( .A(a_29_), .ZN(n7946) );
  NOR2_X2 U7362 ( .A1(n14290), .A2(n14287), .ZN(n7954) );
  XOR2_X1 U7363 ( .A(n7249), .B(n7250), .Z(Result_mul_9_) );
  AND2_X1 U7364 ( .A1(n7251), .A2(n7252), .ZN(n7250) );
  XOR2_X1 U7365 ( .A(n7253), .B(n7254), .Z(Result_mul_8_) );
  AND2_X1 U7366 ( .A1(n7255), .A2(n7256), .ZN(n7254) );
  XOR2_X1 U7367 ( .A(n7257), .B(n7258), .Z(Result_mul_7_) );
  AND2_X1 U7368 ( .A1(n7259), .A2(n7260), .ZN(n7258) );
  XOR2_X1 U7369 ( .A(n7261), .B(n7262), .Z(Result_mul_6_) );
  AND2_X1 U7370 ( .A1(n7263), .A2(n7264), .ZN(n7262) );
  NAND2_X1 U7371 ( .A1(n7265), .A2(n7266), .ZN(Result_mul_62_) );
  NAND2_X1 U7372 ( .A1(b_30_), .A2(n7267), .ZN(n7266) );
  NAND2_X1 U7373 ( .A1(n7268), .A2(n7269), .ZN(n7267) );
  NAND2_X1 U7374 ( .A1(a_31_), .A2(n7270), .ZN(n7269) );
  NAND2_X1 U7375 ( .A1(b_31_), .A2(n7271), .ZN(n7265) );
  NAND2_X1 U7376 ( .A1(n7272), .A2(n7273), .ZN(n7271) );
  NAND2_X1 U7377 ( .A1(a_30_), .A2(n7274), .ZN(n7273) );
  XOR2_X1 U7378 ( .A(n7275), .B(n7276), .Z(Result_mul_61_) );
  XOR2_X1 U7379 ( .A(n7277), .B(n7278), .Z(n7276) );
  NAND2_X1 U7380 ( .A1(b_31_), .A2(a_29_), .ZN(n7275) );
  XOR2_X1 U7381 ( .A(n7279), .B(n7280), .Z(Result_mul_60_) );
  XNOR2_X1 U7382 ( .A(n7281), .B(n7282), .ZN(n7280) );
  NAND2_X1 U7383 ( .A1(b_31_), .A2(a_28_), .ZN(n7282) );
  XOR2_X1 U7384 ( .A(n7283), .B(n7284), .Z(Result_mul_5_) );
  AND2_X1 U7385 ( .A1(n7285), .A2(n7286), .ZN(n7284) );
  XNOR2_X1 U7386 ( .A(n7287), .B(n7288), .ZN(Result_mul_59_) );
  NAND2_X1 U7387 ( .A1(n7289), .A2(n7290), .ZN(n7287) );
  XOR2_X1 U7388 ( .A(n7291), .B(n7292), .Z(Result_mul_58_) );
  XOR2_X1 U7389 ( .A(n7293), .B(n7294), .Z(n7291) );
  NOR2_X1 U7390 ( .A1(n7295), .A2(n7270), .ZN(n7294) );
  XNOR2_X1 U7391 ( .A(n7296), .B(n7297), .ZN(Result_mul_57_) );
  NAND2_X1 U7392 ( .A1(n7298), .A2(n7299), .ZN(n7296) );
  XOR2_X1 U7393 ( .A(n7300), .B(n7301), .Z(Result_mul_56_) );
  XNOR2_X1 U7394 ( .A(n7302), .B(n7303), .ZN(n7301) );
  NAND2_X1 U7395 ( .A1(b_31_), .A2(a_24_), .ZN(n7302) );
  XNOR2_X1 U7396 ( .A(n7304), .B(n7305), .ZN(Result_mul_55_) );
  NAND2_X1 U7397 ( .A1(n7306), .A2(n7307), .ZN(n7304) );
  XOR2_X1 U7398 ( .A(n7308), .B(n7309), .Z(Result_mul_54_) );
  XOR2_X1 U7399 ( .A(n7310), .B(n7311), .Z(n7309) );
  NOR2_X1 U7400 ( .A1(n7312), .A2(n7270), .ZN(n7311) );
  XOR2_X1 U7401 ( .A(n7313), .B(n7314), .Z(Result_mul_53_) );
  XNOR2_X1 U7402 ( .A(n7315), .B(n7316), .ZN(n7314) );
  NAND2_X1 U7403 ( .A1(b_31_), .A2(a_21_), .ZN(n7316) );
  XOR2_X1 U7404 ( .A(n7317), .B(n7318), .Z(Result_mul_52_) );
  XNOR2_X1 U7405 ( .A(n7319), .B(n7320), .ZN(n7318) );
  NAND2_X1 U7406 ( .A1(b_31_), .A2(a_20_), .ZN(n7320) );
  XNOR2_X1 U7407 ( .A(n7321), .B(n7322), .ZN(Result_mul_51_) );
  XOR2_X1 U7408 ( .A(n7323), .B(n7324), .Z(n7322) );
  NAND2_X1 U7409 ( .A1(b_31_), .A2(a_19_), .ZN(n7324) );
  XOR2_X1 U7410 ( .A(n7325), .B(n7326), .Z(Result_mul_50_) );
  XNOR2_X1 U7411 ( .A(n7327), .B(n7328), .ZN(n7326) );
  NAND2_X1 U7412 ( .A1(b_31_), .A2(a_18_), .ZN(n7328) );
  XOR2_X1 U7413 ( .A(n7329), .B(n7330), .Z(Result_mul_4_) );
  AND2_X1 U7414 ( .A1(n7331), .A2(n7332), .ZN(n7330) );
  XOR2_X1 U7415 ( .A(n7333), .B(n7334), .Z(Result_mul_49_) );
  XOR2_X1 U7416 ( .A(n7335), .B(n7336), .Z(n7333) );
  NOR2_X1 U7417 ( .A1(n7337), .A2(n7270), .ZN(n7336) );
  XOR2_X1 U7418 ( .A(n7338), .B(n7339), .Z(Result_mul_48_) );
  XNOR2_X1 U7419 ( .A(n7340), .B(n7341), .ZN(n7339) );
  NAND2_X1 U7420 ( .A1(b_31_), .A2(a_16_), .ZN(n7341) );
  XOR2_X1 U7421 ( .A(n7342), .B(n7343), .Z(Result_mul_47_) );
  XOR2_X1 U7422 ( .A(n7344), .B(n7345), .Z(n7342) );
  NOR2_X1 U7423 ( .A1(n7346), .A2(n7270), .ZN(n7345) );
  XOR2_X1 U7424 ( .A(n7347), .B(n7348), .Z(Result_mul_46_) );
  XNOR2_X1 U7425 ( .A(n7349), .B(n7350), .ZN(n7348) );
  NAND2_X1 U7426 ( .A1(b_31_), .A2(a_14_), .ZN(n7350) );
  XOR2_X1 U7427 ( .A(n7351), .B(n7352), .Z(Result_mul_45_) );
  XOR2_X1 U7428 ( .A(n7353), .B(n7354), .Z(n7351) );
  NOR2_X1 U7429 ( .A1(n7355), .A2(n7270), .ZN(n7354) );
  XOR2_X1 U7430 ( .A(n7356), .B(n7357), .Z(Result_mul_44_) );
  XNOR2_X1 U7431 ( .A(n7358), .B(n7359), .ZN(n7357) );
  NAND2_X1 U7432 ( .A1(b_31_), .A2(a_12_), .ZN(n7359) );
  XNOR2_X1 U7433 ( .A(n7360), .B(n7361), .ZN(Result_mul_43_) );
  XOR2_X1 U7434 ( .A(n7362), .B(n7363), .Z(n7361) );
  NAND2_X1 U7435 ( .A1(b_31_), .A2(a_11_), .ZN(n7363) );
  XOR2_X1 U7436 ( .A(n7364), .B(n7365), .Z(Result_mul_42_) );
  XNOR2_X1 U7437 ( .A(n7366), .B(n7367), .ZN(n7365) );
  NAND2_X1 U7438 ( .A1(b_31_), .A2(a_10_), .ZN(n7367) );
  XOR2_X1 U7439 ( .A(n7368), .B(n7369), .Z(Result_mul_41_) );
  XNOR2_X1 U7440 ( .A(n7370), .B(n7371), .ZN(n7369) );
  NAND2_X1 U7441 ( .A1(b_31_), .A2(a_9_), .ZN(n7371) );
  XOR2_X1 U7442 ( .A(n7372), .B(n7373), .Z(Result_mul_40_) );
  XNOR2_X1 U7443 ( .A(n7374), .B(n7375), .ZN(n7373) );
  NAND2_X1 U7444 ( .A1(b_31_), .A2(a_8_), .ZN(n7375) );
  XOR2_X1 U7445 ( .A(n7376), .B(n7377), .Z(Result_mul_3_) );
  AND2_X1 U7446 ( .A1(n7378), .A2(n7379), .ZN(n7377) );
  XNOR2_X1 U7447 ( .A(n7380), .B(n7381), .ZN(Result_mul_39_) );
  XOR2_X1 U7448 ( .A(n7382), .B(n7383), .Z(n7381) );
  NAND2_X1 U7449 ( .A1(b_31_), .A2(a_7_), .ZN(n7383) );
  XOR2_X1 U7450 ( .A(n7384), .B(n7385), .Z(Result_mul_38_) );
  XOR2_X1 U7451 ( .A(n7386), .B(n7387), .Z(n7384) );
  NOR2_X1 U7452 ( .A1(n7388), .A2(n7270), .ZN(n7387) );
  XOR2_X1 U7453 ( .A(n7389), .B(n7390), .Z(Result_mul_37_) );
  XOR2_X1 U7454 ( .A(n7391), .B(n7392), .Z(n7389) );
  NOR2_X1 U7455 ( .A1(n7393), .A2(n7270), .ZN(n7392) );
  XOR2_X1 U7456 ( .A(n7394), .B(n7395), .Z(Result_mul_36_) );
  XOR2_X1 U7457 ( .A(n7396), .B(n7397), .Z(n7394) );
  NOR2_X1 U7458 ( .A1(n7398), .A2(n7270), .ZN(n7397) );
  XNOR2_X1 U7459 ( .A(n7399), .B(n7400), .ZN(Result_mul_35_) );
  XOR2_X1 U7460 ( .A(n7401), .B(n7402), .Z(n7400) );
  NAND2_X1 U7461 ( .A1(b_31_), .A2(a_3_), .ZN(n7402) );
  XOR2_X1 U7462 ( .A(n7403), .B(n7404), .Z(Result_mul_34_) );
  XNOR2_X1 U7463 ( .A(n7405), .B(n7406), .ZN(n7404) );
  NAND2_X1 U7464 ( .A1(b_31_), .A2(a_2_), .ZN(n7406) );
  XOR2_X1 U7465 ( .A(n7407), .B(n7408), .Z(Result_mul_33_) );
  XOR2_X1 U7466 ( .A(n7409), .B(n7410), .Z(n7407) );
  NOR2_X1 U7467 ( .A1(n7411), .A2(n7270), .ZN(n7410) );
  INV_X1 U7468 ( .A(b_31_), .ZN(n7270) );
  XOR2_X1 U7469 ( .A(n7412), .B(n7413), .Z(Result_mul_32_) );
  XNOR2_X1 U7470 ( .A(n7414), .B(n7415), .ZN(n7413) );
  NAND2_X1 U7471 ( .A1(b_31_), .A2(a_0_), .ZN(n7415) );
  XOR2_X1 U7472 ( .A(n7416), .B(n7417), .Z(Result_mul_31_) );
  NOR2_X1 U7473 ( .A1(n7418), .A2(n7419), .ZN(Result_mul_30_) );
  NOR2_X1 U7474 ( .A1(n7420), .A2(n7421), .ZN(n7419) );
  AND2_X1 U7475 ( .A1(n7417), .A2(n7416), .ZN(n7420) );
  XOR2_X1 U7476 ( .A(n7422), .B(n7423), .Z(Result_mul_2_) );
  AND2_X1 U7477 ( .A1(n7424), .A2(n7425), .ZN(n7423) );
  XNOR2_X1 U7478 ( .A(n7418), .B(n7426), .ZN(Result_mul_29_) );
  NAND2_X1 U7479 ( .A1(n7427), .A2(n7428), .ZN(n7426) );
  XNOR2_X1 U7480 ( .A(n7429), .B(n7430), .ZN(Result_mul_28_) );
  NAND2_X1 U7481 ( .A1(n7431), .A2(n7432), .ZN(n7429) );
  XNOR2_X1 U7482 ( .A(n7433), .B(n7434), .ZN(Result_mul_27_) );
  NAND2_X1 U7483 ( .A1(n7435), .A2(n7436), .ZN(n7433) );
  XOR2_X1 U7484 ( .A(n7437), .B(n7438), .Z(Result_mul_26_) );
  AND2_X1 U7485 ( .A1(n7439), .A2(n7440), .ZN(n7438) );
  XOR2_X1 U7486 ( .A(n7441), .B(n7442), .Z(Result_mul_25_) );
  AND2_X1 U7487 ( .A1(n7443), .A2(n7444), .ZN(n7442) );
  XOR2_X1 U7488 ( .A(n7445), .B(n7446), .Z(Result_mul_24_) );
  AND2_X1 U7489 ( .A1(n7447), .A2(n7448), .ZN(n7446) );
  XOR2_X1 U7490 ( .A(n7449), .B(n7450), .Z(Result_mul_23_) );
  AND2_X1 U7491 ( .A1(n7451), .A2(n7452), .ZN(n7450) );
  XOR2_X1 U7492 ( .A(n7453), .B(n7454), .Z(Result_mul_22_) );
  AND2_X1 U7493 ( .A1(n7455), .A2(n7456), .ZN(n7454) );
  XOR2_X1 U7494 ( .A(n7457), .B(n7458), .Z(Result_mul_21_) );
  AND2_X1 U7495 ( .A1(n7459), .A2(n7460), .ZN(n7458) );
  XOR2_X1 U7496 ( .A(n7461), .B(n7462), .Z(Result_mul_20_) );
  AND2_X1 U7497 ( .A1(n7463), .A2(n7464), .ZN(n7462) );
  XOR2_X1 U7498 ( .A(n7465), .B(n7466), .Z(Result_mul_1_) );
  AND2_X1 U7499 ( .A1(n7467), .A2(n7468), .ZN(n7466) );
  XOR2_X1 U7500 ( .A(n7469), .B(n7470), .Z(Result_mul_19_) );
  AND2_X1 U7501 ( .A1(n7471), .A2(n7472), .ZN(n7470) );
  XOR2_X1 U7502 ( .A(n7473), .B(n7474), .Z(Result_mul_18_) );
  AND2_X1 U7503 ( .A1(n7475), .A2(n7476), .ZN(n7474) );
  XOR2_X1 U7504 ( .A(n7477), .B(n7478), .Z(Result_mul_17_) );
  AND2_X1 U7505 ( .A1(n7479), .A2(n7480), .ZN(n7478) );
  XOR2_X1 U7506 ( .A(n7481), .B(n7482), .Z(Result_mul_16_) );
  AND2_X1 U7507 ( .A1(n7483), .A2(n7484), .ZN(n7482) );
  XOR2_X1 U7508 ( .A(n7485), .B(n7486), .Z(Result_mul_15_) );
  AND2_X1 U7509 ( .A1(n7487), .A2(n7488), .ZN(n7486) );
  XOR2_X1 U7510 ( .A(n7489), .B(n7490), .Z(Result_mul_14_) );
  AND2_X1 U7511 ( .A1(n7491), .A2(n7492), .ZN(n7490) );
  XOR2_X1 U7512 ( .A(n7493), .B(n7494), .Z(Result_mul_13_) );
  AND2_X1 U7513 ( .A1(n7495), .A2(n7496), .ZN(n7494) );
  XOR2_X1 U7514 ( .A(n7497), .B(n7498), .Z(Result_mul_12_) );
  AND2_X1 U7515 ( .A1(n7499), .A2(n7500), .ZN(n7498) );
  XOR2_X1 U7516 ( .A(n7501), .B(n7502), .Z(Result_mul_11_) );
  AND2_X1 U7517 ( .A1(n7503), .A2(n7504), .ZN(n7502) );
  XOR2_X1 U7518 ( .A(n7505), .B(n7506), .Z(Result_mul_10_) );
  AND2_X1 U7519 ( .A1(n7507), .A2(n7508), .ZN(n7506) );
  NAND3_X1 U7520 ( .A1(n7509), .A2(n7468), .A3(n7510), .ZN(Result_mul_0_) );
  NAND2_X1 U7521 ( .A1(a_0_), .A2(n7511), .ZN(n7510) );
  OR4_X1 U7522 ( .A1(n7511), .A2(n7512), .A3(n7513), .A4(n7514), .ZN(n7468) );
  NAND2_X1 U7523 ( .A1(n7467), .A2(n7465), .ZN(n7509) );
  NAND2_X1 U7524 ( .A1(n7425), .A2(n7515), .ZN(n7465) );
  NAND2_X1 U7525 ( .A1(n7424), .A2(n7422), .ZN(n7515) );
  NAND2_X1 U7526 ( .A1(n7379), .A2(n7516), .ZN(n7422) );
  NAND2_X1 U7527 ( .A1(n7378), .A2(n7376), .ZN(n7516) );
  NAND2_X1 U7528 ( .A1(n7332), .A2(n7517), .ZN(n7376) );
  NAND2_X1 U7529 ( .A1(n7331), .A2(n7329), .ZN(n7517) );
  NAND2_X1 U7530 ( .A1(n7286), .A2(n7518), .ZN(n7329) );
  NAND2_X1 U7531 ( .A1(n7285), .A2(n7283), .ZN(n7518) );
  NAND2_X1 U7532 ( .A1(n7264), .A2(n7519), .ZN(n7283) );
  NAND2_X1 U7533 ( .A1(n7263), .A2(n7261), .ZN(n7519) );
  NAND2_X1 U7534 ( .A1(n7260), .A2(n7520), .ZN(n7261) );
  NAND2_X1 U7535 ( .A1(n7259), .A2(n7257), .ZN(n7520) );
  NAND2_X1 U7536 ( .A1(n7256), .A2(n7521), .ZN(n7257) );
  NAND2_X1 U7537 ( .A1(n7255), .A2(n7253), .ZN(n7521) );
  NAND2_X1 U7538 ( .A1(n7252), .A2(n7522), .ZN(n7253) );
  NAND2_X1 U7539 ( .A1(n7251), .A2(n7249), .ZN(n7522) );
  NAND2_X1 U7540 ( .A1(n7508), .A2(n7523), .ZN(n7249) );
  NAND2_X1 U7541 ( .A1(n7505), .A2(n7507), .ZN(n7523) );
  NAND2_X1 U7542 ( .A1(n7524), .A2(n7525), .ZN(n7507) );
  NAND2_X1 U7543 ( .A1(n7504), .A2(n7526), .ZN(n7505) );
  NAND2_X1 U7544 ( .A1(n7501), .A2(n7503), .ZN(n7526) );
  NAND2_X1 U7545 ( .A1(n7527), .A2(n7528), .ZN(n7503) );
  NAND2_X1 U7546 ( .A1(n7529), .A2(n7525), .ZN(n7528) );
  NAND2_X1 U7547 ( .A1(n7530), .A2(n7531), .ZN(n7527) );
  NAND2_X1 U7548 ( .A1(n7500), .A2(n7532), .ZN(n7501) );
  NAND2_X1 U7549 ( .A1(n7497), .A2(n7499), .ZN(n7532) );
  NAND2_X1 U7550 ( .A1(n7533), .A2(n7534), .ZN(n7499) );
  XNOR2_X1 U7551 ( .A(n7530), .B(n7531), .ZN(n7533) );
  NAND2_X1 U7552 ( .A1(n7496), .A2(n7535), .ZN(n7497) );
  NAND2_X1 U7553 ( .A1(n7493), .A2(n7495), .ZN(n7535) );
  NAND2_X1 U7554 ( .A1(n7536), .A2(n7537), .ZN(n7495) );
  NAND2_X1 U7555 ( .A1(n7538), .A2(n7534), .ZN(n7537) );
  NAND2_X1 U7556 ( .A1(n7539), .A2(n7540), .ZN(n7536) );
  NAND2_X1 U7557 ( .A1(n7492), .A2(n7541), .ZN(n7493) );
  NAND2_X1 U7558 ( .A1(n7491), .A2(n7489), .ZN(n7541) );
  NAND2_X1 U7559 ( .A1(n7488), .A2(n7542), .ZN(n7489) );
  NAND2_X1 U7560 ( .A1(n7487), .A2(n7485), .ZN(n7542) );
  NAND2_X1 U7561 ( .A1(n7484), .A2(n7543), .ZN(n7485) );
  NAND2_X1 U7562 ( .A1(n7481), .A2(n7483), .ZN(n7543) );
  NAND2_X1 U7563 ( .A1(n7544), .A2(n7545), .ZN(n7483) );
  NAND2_X1 U7564 ( .A1(n7546), .A2(n7547), .ZN(n7545) );
  XNOR2_X1 U7565 ( .A(n7548), .B(n7549), .ZN(n7544) );
  NAND2_X1 U7566 ( .A1(n7480), .A2(n7550), .ZN(n7481) );
  NAND2_X1 U7567 ( .A1(n7479), .A2(n7477), .ZN(n7550) );
  NAND2_X1 U7568 ( .A1(n7475), .A2(n7551), .ZN(n7477) );
  NAND2_X1 U7569 ( .A1(n7473), .A2(n7476), .ZN(n7551) );
  NAND2_X1 U7570 ( .A1(n7552), .A2(n7553), .ZN(n7476) );
  NAND2_X1 U7571 ( .A1(n7554), .A2(n7555), .ZN(n7553) );
  XNOR2_X1 U7572 ( .A(n7556), .B(n7557), .ZN(n7552) );
  NAND2_X1 U7573 ( .A1(n7472), .A2(n7558), .ZN(n7473) );
  NAND2_X1 U7574 ( .A1(n7469), .A2(n7471), .ZN(n7558) );
  NAND2_X1 U7575 ( .A1(n7559), .A2(n7560), .ZN(n7471) );
  NAND2_X1 U7576 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  XNOR2_X1 U7577 ( .A(n7554), .B(n7555), .ZN(n7559) );
  NAND2_X1 U7578 ( .A1(n7463), .A2(n7563), .ZN(n7469) );
  NAND2_X1 U7579 ( .A1(n7461), .A2(n7464), .ZN(n7563) );
  NAND2_X1 U7580 ( .A1(n7564), .A2(n7565), .ZN(n7464) );
  XOR2_X1 U7581 ( .A(n7562), .B(n7566), .Z(n7564) );
  NAND2_X1 U7582 ( .A1(n7459), .A2(n7567), .ZN(n7461) );
  NAND2_X1 U7583 ( .A1(n7457), .A2(n7460), .ZN(n7567) );
  NAND2_X1 U7584 ( .A1(n7568), .A2(n7569), .ZN(n7460) );
  NAND2_X1 U7585 ( .A1(n7570), .A2(n7565), .ZN(n7569) );
  NAND2_X1 U7586 ( .A1(n7571), .A2(n7572), .ZN(n7568) );
  NAND2_X1 U7587 ( .A1(n7455), .A2(n7573), .ZN(n7457) );
  NAND2_X1 U7588 ( .A1(n7453), .A2(n7456), .ZN(n7573) );
  NAND2_X1 U7589 ( .A1(n7574), .A2(n7575), .ZN(n7456) );
  NAND2_X1 U7590 ( .A1(n7576), .A2(n7577), .ZN(n7575) );
  XNOR2_X1 U7591 ( .A(n7572), .B(n7571), .ZN(n7574) );
  NAND2_X1 U7592 ( .A1(n7452), .A2(n7578), .ZN(n7453) );
  NAND2_X1 U7593 ( .A1(n7449), .A2(n7451), .ZN(n7578) );
  NAND2_X1 U7594 ( .A1(n7579), .A2(n7580), .ZN(n7451) );
  NAND2_X1 U7595 ( .A1(n7581), .A2(n7582), .ZN(n7580) );
  XNOR2_X1 U7596 ( .A(n7577), .B(n7576), .ZN(n7579) );
  NAND2_X1 U7597 ( .A1(n7447), .A2(n7583), .ZN(n7449) );
  NAND2_X1 U7598 ( .A1(n7445), .A2(n7448), .ZN(n7583) );
  NAND2_X1 U7599 ( .A1(n7584), .A2(n7585), .ZN(n7448) );
  XOR2_X1 U7600 ( .A(n7582), .B(n7586), .Z(n7584) );
  NAND2_X1 U7601 ( .A1(n7443), .A2(n7587), .ZN(n7445) );
  NAND2_X1 U7602 ( .A1(n7441), .A2(n7444), .ZN(n7587) );
  NAND2_X1 U7603 ( .A1(n7588), .A2(n7589), .ZN(n7444) );
  NAND2_X1 U7604 ( .A1(n7590), .A2(n7585), .ZN(n7589) );
  NAND2_X1 U7605 ( .A1(n7591), .A2(n7592), .ZN(n7588) );
  NAND2_X1 U7606 ( .A1(n7440), .A2(n7593), .ZN(n7441) );
  NAND2_X1 U7607 ( .A1(n7439), .A2(n7437), .ZN(n7593) );
  NAND2_X1 U7608 ( .A1(n7594), .A2(n7435), .ZN(n7437) );
  OR2_X1 U7609 ( .A1(n7595), .A2(n7596), .ZN(n7435) );
  NAND2_X1 U7610 ( .A1(n7436), .A2(n7434), .ZN(n7594) );
  NAND2_X1 U7611 ( .A1(n7597), .A2(n7432), .ZN(n7434) );
  NAND4_X1 U7612 ( .A1(n7598), .A2(n7599), .A3(n7600), .A4(n7596), .ZN(n7432)
         );
  NAND2_X1 U7613 ( .A1(n7601), .A2(n7602), .ZN(n7599) );
  NAND2_X1 U7614 ( .A1(n7431), .A2(n7430), .ZN(n7597) );
  NAND2_X1 U7615 ( .A1(n7428), .A2(n7603), .ZN(n7430) );
  NAND2_X1 U7616 ( .A1(n7418), .A2(n7427), .ZN(n7603) );
  NAND2_X1 U7617 ( .A1(n7604), .A2(n7605), .ZN(n7427) );
  NAND2_X1 U7618 ( .A1(n7606), .A2(n7607), .ZN(n7605) );
  XOR2_X1 U7619 ( .A(n7600), .B(n7608), .Z(n7604) );
  AND3_X1 U7620 ( .A1(n7421), .A2(n7417), .A3(n7416), .ZN(n7418) );
  XNOR2_X1 U7621 ( .A(n7609), .B(n7610), .ZN(n7416) );
  XNOR2_X1 U7622 ( .A(n7611), .B(n7612), .ZN(n7609) );
  NOR2_X1 U7623 ( .A1(n7613), .A2(n7274), .ZN(n7612) );
  NAND2_X1 U7624 ( .A1(n7614), .A2(n7615), .ZN(n7417) );
  NAND3_X1 U7625 ( .A1(a_0_), .A2(n7616), .A3(b_31_), .ZN(n7615) );
  NAND2_X1 U7626 ( .A1(n7414), .A2(n7412), .ZN(n7616) );
  OR2_X1 U7627 ( .A1(n7412), .A2(n7414), .ZN(n7614) );
  AND2_X1 U7628 ( .A1(n7617), .A2(n7618), .ZN(n7414) );
  NAND3_X1 U7629 ( .A1(a_1_), .A2(n7619), .A3(b_31_), .ZN(n7618) );
  OR2_X1 U7630 ( .A1(n7409), .A2(n7408), .ZN(n7619) );
  NAND2_X1 U7631 ( .A1(n7408), .A2(n7409), .ZN(n7617) );
  NAND2_X1 U7632 ( .A1(n7620), .A2(n7621), .ZN(n7409) );
  NAND3_X1 U7633 ( .A1(a_2_), .A2(n7622), .A3(b_31_), .ZN(n7621) );
  NAND2_X1 U7634 ( .A1(n7405), .A2(n7403), .ZN(n7622) );
  OR2_X1 U7635 ( .A1(n7403), .A2(n7405), .ZN(n7620) );
  AND2_X1 U7636 ( .A1(n7623), .A2(n7624), .ZN(n7405) );
  NAND3_X1 U7637 ( .A1(a_3_), .A2(n7625), .A3(b_31_), .ZN(n7624) );
  OR2_X1 U7638 ( .A1(n7401), .A2(n7399), .ZN(n7625) );
  NAND2_X1 U7639 ( .A1(n7399), .A2(n7401), .ZN(n7623) );
  NAND2_X1 U7640 ( .A1(n7626), .A2(n7627), .ZN(n7401) );
  NAND3_X1 U7641 ( .A1(a_4_), .A2(n7628), .A3(b_31_), .ZN(n7627) );
  OR2_X1 U7642 ( .A1(n7396), .A2(n7395), .ZN(n7628) );
  NAND2_X1 U7643 ( .A1(n7395), .A2(n7396), .ZN(n7626) );
  NAND2_X1 U7644 ( .A1(n7629), .A2(n7630), .ZN(n7396) );
  NAND3_X1 U7645 ( .A1(a_5_), .A2(n7631), .A3(b_31_), .ZN(n7630) );
  OR2_X1 U7646 ( .A1(n7391), .A2(n7390), .ZN(n7631) );
  NAND2_X1 U7647 ( .A1(n7390), .A2(n7391), .ZN(n7629) );
  NAND2_X1 U7648 ( .A1(n7632), .A2(n7633), .ZN(n7391) );
  NAND3_X1 U7649 ( .A1(a_6_), .A2(n7634), .A3(b_31_), .ZN(n7633) );
  OR2_X1 U7650 ( .A1(n7386), .A2(n7385), .ZN(n7634) );
  NAND2_X1 U7651 ( .A1(n7385), .A2(n7386), .ZN(n7632) );
  NAND2_X1 U7652 ( .A1(n7635), .A2(n7636), .ZN(n7386) );
  NAND3_X1 U7653 ( .A1(a_7_), .A2(n7637), .A3(b_31_), .ZN(n7636) );
  OR2_X1 U7654 ( .A1(n7382), .A2(n7380), .ZN(n7637) );
  NAND2_X1 U7655 ( .A1(n7380), .A2(n7382), .ZN(n7635) );
  NAND2_X1 U7656 ( .A1(n7638), .A2(n7639), .ZN(n7382) );
  NAND3_X1 U7657 ( .A1(a_8_), .A2(n7640), .A3(b_31_), .ZN(n7639) );
  NAND2_X1 U7658 ( .A1(n7374), .A2(n7372), .ZN(n7640) );
  OR2_X1 U7659 ( .A1(n7372), .A2(n7374), .ZN(n7638) );
  AND2_X1 U7660 ( .A1(n7641), .A2(n7642), .ZN(n7374) );
  NAND3_X1 U7661 ( .A1(a_9_), .A2(n7643), .A3(b_31_), .ZN(n7642) );
  NAND2_X1 U7662 ( .A1(n7370), .A2(n7368), .ZN(n7643) );
  OR2_X1 U7663 ( .A1(n7368), .A2(n7370), .ZN(n7641) );
  AND2_X1 U7664 ( .A1(n7644), .A2(n7645), .ZN(n7370) );
  NAND3_X1 U7665 ( .A1(a_10_), .A2(n7646), .A3(b_31_), .ZN(n7645) );
  NAND2_X1 U7666 ( .A1(n7366), .A2(n7364), .ZN(n7646) );
  OR2_X1 U7667 ( .A1(n7364), .A2(n7366), .ZN(n7644) );
  AND2_X1 U7668 ( .A1(n7647), .A2(n7648), .ZN(n7366) );
  NAND3_X1 U7669 ( .A1(a_11_), .A2(n7649), .A3(b_31_), .ZN(n7648) );
  OR2_X1 U7670 ( .A1(n7362), .A2(n7360), .ZN(n7649) );
  NAND2_X1 U7671 ( .A1(n7360), .A2(n7362), .ZN(n7647) );
  NAND2_X1 U7672 ( .A1(n7650), .A2(n7651), .ZN(n7362) );
  NAND3_X1 U7673 ( .A1(a_12_), .A2(n7652), .A3(b_31_), .ZN(n7651) );
  NAND2_X1 U7674 ( .A1(n7358), .A2(n7356), .ZN(n7652) );
  OR2_X1 U7675 ( .A1(n7356), .A2(n7358), .ZN(n7650) );
  AND2_X1 U7676 ( .A1(n7653), .A2(n7654), .ZN(n7358) );
  NAND3_X1 U7677 ( .A1(a_13_), .A2(n7655), .A3(b_31_), .ZN(n7654) );
  OR2_X1 U7678 ( .A1(n7353), .A2(n7352), .ZN(n7655) );
  NAND2_X1 U7679 ( .A1(n7352), .A2(n7353), .ZN(n7653) );
  NAND2_X1 U7680 ( .A1(n7656), .A2(n7657), .ZN(n7353) );
  NAND3_X1 U7681 ( .A1(a_14_), .A2(n7658), .A3(b_31_), .ZN(n7657) );
  NAND2_X1 U7682 ( .A1(n7349), .A2(n7347), .ZN(n7658) );
  OR2_X1 U7683 ( .A1(n7347), .A2(n7349), .ZN(n7656) );
  AND2_X1 U7684 ( .A1(n7659), .A2(n7660), .ZN(n7349) );
  NAND3_X1 U7685 ( .A1(a_15_), .A2(n7661), .A3(b_31_), .ZN(n7660) );
  OR2_X1 U7686 ( .A1(n7344), .A2(n7343), .ZN(n7661) );
  NAND2_X1 U7687 ( .A1(n7343), .A2(n7344), .ZN(n7659) );
  NAND2_X1 U7688 ( .A1(n7662), .A2(n7663), .ZN(n7344) );
  NAND3_X1 U7689 ( .A1(a_16_), .A2(n7664), .A3(b_31_), .ZN(n7663) );
  NAND2_X1 U7690 ( .A1(n7340), .A2(n7338), .ZN(n7664) );
  OR2_X1 U7691 ( .A1(n7338), .A2(n7340), .ZN(n7662) );
  AND2_X1 U7692 ( .A1(n7665), .A2(n7666), .ZN(n7340) );
  NAND3_X1 U7693 ( .A1(a_17_), .A2(n7667), .A3(b_31_), .ZN(n7666) );
  OR2_X1 U7694 ( .A1(n7335), .A2(n7334), .ZN(n7667) );
  NAND2_X1 U7695 ( .A1(n7334), .A2(n7335), .ZN(n7665) );
  NAND2_X1 U7696 ( .A1(n7668), .A2(n7669), .ZN(n7335) );
  NAND3_X1 U7697 ( .A1(a_18_), .A2(n7670), .A3(b_31_), .ZN(n7669) );
  NAND2_X1 U7698 ( .A1(n7327), .A2(n7325), .ZN(n7670) );
  OR2_X1 U7699 ( .A1(n7325), .A2(n7327), .ZN(n7668) );
  AND2_X1 U7700 ( .A1(n7671), .A2(n7672), .ZN(n7327) );
  NAND3_X1 U7701 ( .A1(a_19_), .A2(n7673), .A3(b_31_), .ZN(n7672) );
  OR2_X1 U7702 ( .A1(n7323), .A2(n7321), .ZN(n7673) );
  NAND2_X1 U7703 ( .A1(n7321), .A2(n7323), .ZN(n7671) );
  NAND2_X1 U7704 ( .A1(n7674), .A2(n7675), .ZN(n7323) );
  NAND3_X1 U7705 ( .A1(a_20_), .A2(n7676), .A3(b_31_), .ZN(n7675) );
  NAND2_X1 U7706 ( .A1(n7319), .A2(n7317), .ZN(n7676) );
  OR2_X1 U7707 ( .A1(n7317), .A2(n7319), .ZN(n7674) );
  AND2_X1 U7708 ( .A1(n7677), .A2(n7678), .ZN(n7319) );
  NAND3_X1 U7709 ( .A1(a_21_), .A2(n7679), .A3(b_31_), .ZN(n7678) );
  NAND2_X1 U7710 ( .A1(n7315), .A2(n7313), .ZN(n7679) );
  OR2_X1 U7711 ( .A1(n7313), .A2(n7315), .ZN(n7677) );
  AND2_X1 U7712 ( .A1(n7680), .A2(n7681), .ZN(n7315) );
  NAND3_X1 U7713 ( .A1(a_22_), .A2(n7682), .A3(b_31_), .ZN(n7681) );
  NAND2_X1 U7714 ( .A1(n7310), .A2(n7308), .ZN(n7682) );
  OR2_X1 U7715 ( .A1(n7308), .A2(n7310), .ZN(n7680) );
  AND2_X1 U7716 ( .A1(n7306), .A2(n7683), .ZN(n7310) );
  NAND2_X1 U7717 ( .A1(n7305), .A2(n7307), .ZN(n7683) );
  NAND2_X1 U7718 ( .A1(n7684), .A2(n7685), .ZN(n7307) );
  NAND2_X1 U7719 ( .A1(b_31_), .A2(a_23_), .ZN(n7685) );
  INV_X1 U7720 ( .A(n7686), .ZN(n7684) );
  XOR2_X1 U7721 ( .A(n7687), .B(n7688), .Z(n7305) );
  XOR2_X1 U7722 ( .A(n7689), .B(n7690), .Z(n7687) );
  NOR2_X1 U7723 ( .A1(n7691), .A2(n7274), .ZN(n7690) );
  NAND2_X1 U7724 ( .A1(a_23_), .A2(n7686), .ZN(n7306) );
  NAND2_X1 U7725 ( .A1(n7692), .A2(n7693), .ZN(n7686) );
  NAND3_X1 U7726 ( .A1(a_24_), .A2(n7694), .A3(b_31_), .ZN(n7693) );
  OR2_X1 U7727 ( .A1(n7303), .A2(n7300), .ZN(n7694) );
  NAND2_X1 U7728 ( .A1(n7300), .A2(n7303), .ZN(n7692) );
  NAND2_X1 U7729 ( .A1(n7298), .A2(n7695), .ZN(n7303) );
  NAND2_X1 U7730 ( .A1(n7297), .A2(n7299), .ZN(n7695) );
  NAND2_X1 U7731 ( .A1(n7696), .A2(n7697), .ZN(n7299) );
  NAND2_X1 U7732 ( .A1(b_31_), .A2(a_25_), .ZN(n7697) );
  INV_X1 U7733 ( .A(n7698), .ZN(n7696) );
  XNOR2_X1 U7734 ( .A(n7699), .B(n7700), .ZN(n7297) );
  NAND2_X1 U7735 ( .A1(n7701), .A2(n7702), .ZN(n7699) );
  NAND2_X1 U7736 ( .A1(a_25_), .A2(n7698), .ZN(n7298) );
  NAND2_X1 U7737 ( .A1(n7703), .A2(n7704), .ZN(n7698) );
  NAND3_X1 U7738 ( .A1(a_26_), .A2(n7705), .A3(b_31_), .ZN(n7704) );
  OR2_X1 U7739 ( .A1(n7293), .A2(n7292), .ZN(n7705) );
  NAND2_X1 U7740 ( .A1(n7292), .A2(n7293), .ZN(n7703) );
  NAND2_X1 U7741 ( .A1(n7289), .A2(n7706), .ZN(n7293) );
  NAND2_X1 U7742 ( .A1(n7288), .A2(n7290), .ZN(n7706) );
  NAND2_X1 U7743 ( .A1(n7707), .A2(n7708), .ZN(n7290) );
  NAND2_X1 U7744 ( .A1(b_31_), .A2(a_27_), .ZN(n7708) );
  INV_X1 U7745 ( .A(n7709), .ZN(n7707) );
  XNOR2_X1 U7746 ( .A(n7710), .B(n7711), .ZN(n7288) );
  XOR2_X1 U7747 ( .A(n7712), .B(n7713), .Z(n7710) );
  NAND2_X1 U7748 ( .A1(b_30_), .A2(a_28_), .ZN(n7712) );
  NAND2_X1 U7749 ( .A1(a_27_), .A2(n7709), .ZN(n7289) );
  NAND2_X1 U7750 ( .A1(n7714), .A2(n7715), .ZN(n7709) );
  NAND3_X1 U7751 ( .A1(a_28_), .A2(n7716), .A3(b_31_), .ZN(n7715) );
  NAND2_X1 U7752 ( .A1(n7281), .A2(n7279), .ZN(n7716) );
  OR2_X1 U7753 ( .A1(n7279), .A2(n7281), .ZN(n7714) );
  AND2_X1 U7754 ( .A1(n7717), .A2(n7718), .ZN(n7281) );
  NAND3_X1 U7755 ( .A1(a_29_), .A2(n7719), .A3(b_31_), .ZN(n7718) );
  OR2_X1 U7756 ( .A1(n7278), .A2(n7720), .ZN(n7719) );
  NAND2_X1 U7757 ( .A1(n7720), .A2(n7278), .ZN(n7717) );
  NAND3_X1 U7758 ( .A1(n7721), .A2(n7722), .A3(n7723), .ZN(n7278) );
  OR2_X1 U7759 ( .A1(n7272), .A2(n7274), .ZN(n7723) );
  NAND2_X1 U7760 ( .A1(n7724), .A2(n7725), .ZN(n7722) );
  NAND2_X1 U7761 ( .A1(b_29_), .A2(n7726), .ZN(n7721) );
  NAND2_X1 U7762 ( .A1(n7268), .A2(n7727), .ZN(n7726) );
  NAND2_X1 U7763 ( .A1(a_31_), .A2(n7274), .ZN(n7727) );
  INV_X1 U7764 ( .A(n7277), .ZN(n7720) );
  XNOR2_X1 U7765 ( .A(n7728), .B(n7729), .ZN(n7279) );
  XOR2_X1 U7766 ( .A(n7730), .B(n7731), .Z(n7728) );
  XNOR2_X1 U7767 ( .A(n7732), .B(n7733), .ZN(n7292) );
  NAND2_X1 U7768 ( .A1(n7734), .A2(n7735), .ZN(n7732) );
  XOR2_X1 U7769 ( .A(n7736), .B(n7737), .Z(n7300) );
  XOR2_X1 U7770 ( .A(n7738), .B(n7739), .Z(n7736) );
  XNOR2_X1 U7771 ( .A(n7740), .B(n7741), .ZN(n7308) );
  XOR2_X1 U7772 ( .A(n7742), .B(n7743), .Z(n7740) );
  XNOR2_X1 U7773 ( .A(n7744), .B(n7745), .ZN(n7313) );
  XOR2_X1 U7774 ( .A(n7746), .B(n7747), .Z(n7744) );
  NOR2_X1 U7775 ( .A1(n7312), .A2(n7274), .ZN(n7747) );
  XNOR2_X1 U7776 ( .A(n7748), .B(n7749), .ZN(n7317) );
  XOR2_X1 U7777 ( .A(n7750), .B(n7751), .Z(n7748) );
  XNOR2_X1 U7778 ( .A(n7752), .B(n7753), .ZN(n7321) );
  XOR2_X1 U7779 ( .A(n7754), .B(n7755), .Z(n7753) );
  NAND2_X1 U7780 ( .A1(b_30_), .A2(a_20_), .ZN(n7755) );
  XOR2_X1 U7781 ( .A(n7756), .B(n7757), .Z(n7325) );
  XNOR2_X1 U7782 ( .A(n7758), .B(n7759), .ZN(n7757) );
  XNOR2_X1 U7783 ( .A(n7760), .B(n7761), .ZN(n7334) );
  XNOR2_X1 U7784 ( .A(n7762), .B(n7763), .ZN(n7760) );
  NOR2_X1 U7785 ( .A1(n7764), .A2(n7274), .ZN(n7763) );
  XOR2_X1 U7786 ( .A(n7765), .B(n7766), .Z(n7338) );
  XNOR2_X1 U7787 ( .A(n7767), .B(n7768), .ZN(n7766) );
  XNOR2_X1 U7788 ( .A(n7769), .B(n7770), .ZN(n7343) );
  XNOR2_X1 U7789 ( .A(n7771), .B(n7772), .ZN(n7769) );
  NOR2_X1 U7790 ( .A1(n7773), .A2(n7274), .ZN(n7772) );
  XOR2_X1 U7791 ( .A(n7774), .B(n7775), .Z(n7347) );
  XNOR2_X1 U7792 ( .A(n7776), .B(n7777), .ZN(n7775) );
  XNOR2_X1 U7793 ( .A(n7778), .B(n7779), .ZN(n7352) );
  XNOR2_X1 U7794 ( .A(n7780), .B(n7781), .ZN(n7778) );
  NOR2_X1 U7795 ( .A1(n7782), .A2(n7274), .ZN(n7781) );
  XNOR2_X1 U7796 ( .A(n7783), .B(n7784), .ZN(n7356) );
  XOR2_X1 U7797 ( .A(n7785), .B(n7786), .Z(n7783) );
  XNOR2_X1 U7798 ( .A(n7787), .B(n7788), .ZN(n7360) );
  XOR2_X1 U7799 ( .A(n7789), .B(n7790), .Z(n7788) );
  NAND2_X1 U7800 ( .A1(b_30_), .A2(a_12_), .ZN(n7790) );
  XOR2_X1 U7801 ( .A(n7791), .B(n7792), .Z(n7364) );
  XNOR2_X1 U7802 ( .A(n7793), .B(n7794), .ZN(n7792) );
  XNOR2_X1 U7803 ( .A(n7795), .B(n7796), .ZN(n7368) );
  XOR2_X1 U7804 ( .A(n7797), .B(n7798), .Z(n7795) );
  NOR2_X1 U7805 ( .A1(n7799), .A2(n7274), .ZN(n7798) );
  XNOR2_X1 U7806 ( .A(n7800), .B(n7801), .ZN(n7372) );
  XOR2_X1 U7807 ( .A(n7802), .B(n7803), .Z(n7800) );
  XNOR2_X1 U7808 ( .A(n7804), .B(n7805), .ZN(n7380) );
  XOR2_X1 U7809 ( .A(n7806), .B(n7807), .Z(n7805) );
  NAND2_X1 U7810 ( .A1(b_30_), .A2(a_8_), .ZN(n7807) );
  XNOR2_X1 U7811 ( .A(n7808), .B(n7809), .ZN(n7385) );
  XNOR2_X1 U7812 ( .A(n7810), .B(n7811), .ZN(n7809) );
  XNOR2_X1 U7813 ( .A(n7812), .B(n7813), .ZN(n7390) );
  XNOR2_X1 U7814 ( .A(n7814), .B(n7815), .ZN(n7812) );
  NOR2_X1 U7815 ( .A1(n7388), .A2(n7274), .ZN(n7815) );
  XNOR2_X1 U7816 ( .A(n7816), .B(n7817), .ZN(n7395) );
  XNOR2_X1 U7817 ( .A(n7818), .B(n7819), .ZN(n7816) );
  XNOR2_X1 U7818 ( .A(n7820), .B(n7821), .ZN(n7399) );
  XNOR2_X1 U7819 ( .A(n7822), .B(n7823), .ZN(n7820) );
  NOR2_X1 U7820 ( .A1(n7398), .A2(n7274), .ZN(n7823) );
  XOR2_X1 U7821 ( .A(n7824), .B(n7825), .Z(n7403) );
  XNOR2_X1 U7822 ( .A(n7826), .B(n7827), .ZN(n7825) );
  XNOR2_X1 U7823 ( .A(n7828), .B(n7829), .ZN(n7408) );
  XNOR2_X1 U7824 ( .A(n7830), .B(n7831), .ZN(n7828) );
  NOR2_X1 U7825 ( .A1(n7832), .A2(n7274), .ZN(n7831) );
  XOR2_X1 U7826 ( .A(n7833), .B(n7834), .Z(n7412) );
  XOR2_X1 U7827 ( .A(n7835), .B(n7836), .Z(n7834) );
  NAND2_X1 U7828 ( .A1(b_30_), .A2(a_1_), .ZN(n7836) );
  XOR2_X1 U7829 ( .A(n7607), .B(n7606), .Z(n7421) );
  NAND3_X1 U7830 ( .A1(n7606), .A2(n7607), .A3(n7837), .ZN(n7428) );
  XOR2_X1 U7831 ( .A(n7598), .B(n7600), .Z(n7837) );
  NAND2_X1 U7832 ( .A1(n7838), .A2(n7839), .ZN(n7607) );
  NAND3_X1 U7833 ( .A1(a_0_), .A2(n7840), .A3(b_30_), .ZN(n7839) );
  NAND2_X1 U7834 ( .A1(n7611), .A2(n7610), .ZN(n7840) );
  OR2_X1 U7835 ( .A1(n7610), .A2(n7611), .ZN(n7838) );
  AND2_X1 U7836 ( .A1(n7841), .A2(n7842), .ZN(n7611) );
  NAND3_X1 U7837 ( .A1(a_1_), .A2(n7843), .A3(b_30_), .ZN(n7842) );
  OR2_X1 U7838 ( .A1(n7833), .A2(n7835), .ZN(n7843) );
  NAND2_X1 U7839 ( .A1(n7833), .A2(n7835), .ZN(n7841) );
  NAND2_X1 U7840 ( .A1(n7844), .A2(n7845), .ZN(n7835) );
  NAND3_X1 U7841 ( .A1(a_2_), .A2(n7846), .A3(b_30_), .ZN(n7845) );
  NAND2_X1 U7842 ( .A1(n7830), .A2(n7829), .ZN(n7846) );
  OR2_X1 U7843 ( .A1(n7829), .A2(n7830), .ZN(n7844) );
  AND2_X1 U7844 ( .A1(n7847), .A2(n7848), .ZN(n7830) );
  NAND2_X1 U7845 ( .A1(n7827), .A2(n7849), .ZN(n7848) );
  OR2_X1 U7846 ( .A1(n7824), .A2(n7826), .ZN(n7849) );
  NOR2_X1 U7847 ( .A1(n7274), .A2(n7850), .ZN(n7827) );
  NAND2_X1 U7848 ( .A1(n7824), .A2(n7826), .ZN(n7847) );
  NAND2_X1 U7849 ( .A1(n7851), .A2(n7852), .ZN(n7826) );
  NAND3_X1 U7850 ( .A1(a_4_), .A2(n7853), .A3(b_30_), .ZN(n7852) );
  NAND2_X1 U7851 ( .A1(n7822), .A2(n7821), .ZN(n7853) );
  OR2_X1 U7852 ( .A1(n7821), .A2(n7822), .ZN(n7851) );
  AND2_X1 U7853 ( .A1(n7854), .A2(n7855), .ZN(n7822) );
  NAND2_X1 U7854 ( .A1(n7819), .A2(n7856), .ZN(n7855) );
  NAND2_X1 U7855 ( .A1(n7818), .A2(n7817), .ZN(n7856) );
  NOR2_X1 U7856 ( .A1(n7274), .A2(n7393), .ZN(n7819) );
  OR2_X1 U7857 ( .A1(n7817), .A2(n7818), .ZN(n7854) );
  AND2_X1 U7858 ( .A1(n7857), .A2(n7858), .ZN(n7818) );
  NAND3_X1 U7859 ( .A1(a_6_), .A2(n7859), .A3(b_30_), .ZN(n7858) );
  NAND2_X1 U7860 ( .A1(n7814), .A2(n7813), .ZN(n7859) );
  OR2_X1 U7861 ( .A1(n7813), .A2(n7814), .ZN(n7857) );
  AND2_X1 U7862 ( .A1(n7860), .A2(n7861), .ZN(n7814) );
  NAND2_X1 U7863 ( .A1(n7811), .A2(n7862), .ZN(n7861) );
  OR2_X1 U7864 ( .A1(n7810), .A2(n7808), .ZN(n7862) );
  NOR2_X1 U7865 ( .A1(n7274), .A2(n7863), .ZN(n7811) );
  NAND2_X1 U7866 ( .A1(n7808), .A2(n7810), .ZN(n7860) );
  NAND2_X1 U7867 ( .A1(n7864), .A2(n7865), .ZN(n7810) );
  NAND3_X1 U7868 ( .A1(a_8_), .A2(n7866), .A3(b_30_), .ZN(n7865) );
  OR2_X1 U7869 ( .A1(n7806), .A2(n7804), .ZN(n7866) );
  NAND2_X1 U7870 ( .A1(n7804), .A2(n7806), .ZN(n7864) );
  NAND2_X1 U7871 ( .A1(n7867), .A2(n7868), .ZN(n7806) );
  NAND2_X1 U7872 ( .A1(n7803), .A2(n7869), .ZN(n7868) );
  OR2_X1 U7873 ( .A1(n7801), .A2(n7802), .ZN(n7869) );
  NOR2_X1 U7874 ( .A1(n7274), .A2(n7870), .ZN(n7803) );
  NAND2_X1 U7875 ( .A1(n7801), .A2(n7802), .ZN(n7867) );
  NAND2_X1 U7876 ( .A1(n7871), .A2(n7872), .ZN(n7802) );
  NAND3_X1 U7877 ( .A1(a_10_), .A2(n7873), .A3(b_30_), .ZN(n7872) );
  OR2_X1 U7878 ( .A1(n7796), .A2(n7797), .ZN(n7873) );
  NAND2_X1 U7879 ( .A1(n7796), .A2(n7797), .ZN(n7871) );
  NAND2_X1 U7880 ( .A1(n7874), .A2(n7875), .ZN(n7797) );
  NAND2_X1 U7881 ( .A1(n7794), .A2(n7876), .ZN(n7875) );
  OR2_X1 U7882 ( .A1(n7791), .A2(n7793), .ZN(n7876) );
  NOR2_X1 U7883 ( .A1(n7274), .A2(n7877), .ZN(n7794) );
  NAND2_X1 U7884 ( .A1(n7791), .A2(n7793), .ZN(n7874) );
  NAND2_X1 U7885 ( .A1(n7878), .A2(n7879), .ZN(n7793) );
  NAND3_X1 U7886 ( .A1(a_12_), .A2(n7880), .A3(b_30_), .ZN(n7879) );
  OR2_X1 U7887 ( .A1(n7789), .A2(n7787), .ZN(n7880) );
  NAND2_X1 U7888 ( .A1(n7787), .A2(n7789), .ZN(n7878) );
  NAND2_X1 U7889 ( .A1(n7881), .A2(n7882), .ZN(n7789) );
  NAND2_X1 U7890 ( .A1(n7786), .A2(n7883), .ZN(n7882) );
  OR2_X1 U7891 ( .A1(n7784), .A2(n7785), .ZN(n7883) );
  NOR2_X1 U7892 ( .A1(n7274), .A2(n7355), .ZN(n7786) );
  NAND2_X1 U7893 ( .A1(n7784), .A2(n7785), .ZN(n7881) );
  NAND2_X1 U7894 ( .A1(n7884), .A2(n7885), .ZN(n7785) );
  NAND3_X1 U7895 ( .A1(a_14_), .A2(n7886), .A3(b_30_), .ZN(n7885) );
  NAND2_X1 U7896 ( .A1(n7780), .A2(n7779), .ZN(n7886) );
  OR2_X1 U7897 ( .A1(n7779), .A2(n7780), .ZN(n7884) );
  AND2_X1 U7898 ( .A1(n7887), .A2(n7888), .ZN(n7780) );
  NAND2_X1 U7899 ( .A1(n7777), .A2(n7889), .ZN(n7888) );
  OR2_X1 U7900 ( .A1(n7774), .A2(n7776), .ZN(n7889) );
  NOR2_X1 U7901 ( .A1(n7274), .A2(n7346), .ZN(n7777) );
  NAND2_X1 U7902 ( .A1(n7774), .A2(n7776), .ZN(n7887) );
  NAND2_X1 U7903 ( .A1(n7890), .A2(n7891), .ZN(n7776) );
  NAND3_X1 U7904 ( .A1(a_16_), .A2(n7892), .A3(b_30_), .ZN(n7891) );
  NAND2_X1 U7905 ( .A1(n7771), .A2(n7770), .ZN(n7892) );
  OR2_X1 U7906 ( .A1(n7770), .A2(n7771), .ZN(n7890) );
  AND2_X1 U7907 ( .A1(n7893), .A2(n7894), .ZN(n7771) );
  NAND2_X1 U7908 ( .A1(n7768), .A2(n7895), .ZN(n7894) );
  OR2_X1 U7909 ( .A1(n7765), .A2(n7767), .ZN(n7895) );
  NOR2_X1 U7910 ( .A1(n7274), .A2(n7337), .ZN(n7768) );
  NAND2_X1 U7911 ( .A1(n7765), .A2(n7767), .ZN(n7893) );
  NAND2_X1 U7912 ( .A1(n7896), .A2(n7897), .ZN(n7767) );
  NAND3_X1 U7913 ( .A1(a_18_), .A2(n7898), .A3(b_30_), .ZN(n7897) );
  NAND2_X1 U7914 ( .A1(n7762), .A2(n7761), .ZN(n7898) );
  OR2_X1 U7915 ( .A1(n7761), .A2(n7762), .ZN(n7896) );
  AND2_X1 U7916 ( .A1(n7899), .A2(n7900), .ZN(n7762) );
  NAND2_X1 U7917 ( .A1(n7759), .A2(n7901), .ZN(n7900) );
  OR2_X1 U7918 ( .A1(n7756), .A2(n7758), .ZN(n7901) );
  NOR2_X1 U7919 ( .A1(n7274), .A2(n7902), .ZN(n7759) );
  NAND2_X1 U7920 ( .A1(n7756), .A2(n7758), .ZN(n7899) );
  NAND2_X1 U7921 ( .A1(n7903), .A2(n7904), .ZN(n7758) );
  NAND3_X1 U7922 ( .A1(a_20_), .A2(n7905), .A3(b_30_), .ZN(n7904) );
  OR2_X1 U7923 ( .A1(n7754), .A2(n7752), .ZN(n7905) );
  NAND2_X1 U7924 ( .A1(n7752), .A2(n7754), .ZN(n7903) );
  NAND2_X1 U7925 ( .A1(n7906), .A2(n7907), .ZN(n7754) );
  NAND2_X1 U7926 ( .A1(n7751), .A2(n7908), .ZN(n7907) );
  OR2_X1 U7927 ( .A1(n7749), .A2(n7750), .ZN(n7908) );
  NOR2_X1 U7928 ( .A1(n7274), .A2(n7909), .ZN(n7751) );
  NAND2_X1 U7929 ( .A1(n7749), .A2(n7750), .ZN(n7906) );
  NAND2_X1 U7930 ( .A1(n7910), .A2(n7911), .ZN(n7750) );
  NAND3_X1 U7931 ( .A1(a_22_), .A2(n7912), .A3(b_30_), .ZN(n7911) );
  OR2_X1 U7932 ( .A1(n7745), .A2(n7746), .ZN(n7912) );
  NAND2_X1 U7933 ( .A1(n7745), .A2(n7746), .ZN(n7910) );
  NAND2_X1 U7934 ( .A1(n7913), .A2(n7914), .ZN(n7746) );
  NAND2_X1 U7935 ( .A1(n7743), .A2(n7915), .ZN(n7914) );
  OR2_X1 U7936 ( .A1(n7741), .A2(n7742), .ZN(n7915) );
  NOR2_X1 U7937 ( .A1(n7274), .A2(n7916), .ZN(n7743) );
  NAND2_X1 U7938 ( .A1(n7741), .A2(n7742), .ZN(n7913) );
  NAND2_X1 U7939 ( .A1(n7917), .A2(n7918), .ZN(n7742) );
  NAND3_X1 U7940 ( .A1(a_24_), .A2(n7919), .A3(b_30_), .ZN(n7918) );
  OR2_X1 U7941 ( .A1(n7688), .A2(n7689), .ZN(n7919) );
  NAND2_X1 U7942 ( .A1(n7688), .A2(n7689), .ZN(n7917) );
  NAND2_X1 U7943 ( .A1(n7920), .A2(n7921), .ZN(n7689) );
  NAND2_X1 U7944 ( .A1(n7739), .A2(n7922), .ZN(n7921) );
  OR2_X1 U7945 ( .A1(n7737), .A2(n7738), .ZN(n7922) );
  NOR2_X1 U7946 ( .A1(n7274), .A2(n7923), .ZN(n7739) );
  NAND2_X1 U7947 ( .A1(n7737), .A2(n7738), .ZN(n7920) );
  NAND2_X1 U7948 ( .A1(n7701), .A2(n7924), .ZN(n7738) );
  NAND2_X1 U7949 ( .A1(n7700), .A2(n7702), .ZN(n7924) );
  NAND2_X1 U7950 ( .A1(n7925), .A2(n7926), .ZN(n7702) );
  NAND2_X1 U7951 ( .A1(b_30_), .A2(a_26_), .ZN(n7926) );
  INV_X1 U7952 ( .A(n7927), .ZN(n7925) );
  XNOR2_X1 U7953 ( .A(n7928), .B(n7929), .ZN(n7700) );
  NAND2_X1 U7954 ( .A1(n7930), .A2(n7931), .ZN(n7928) );
  NAND2_X1 U7955 ( .A1(a_26_), .A2(n7927), .ZN(n7701) );
  NAND2_X1 U7956 ( .A1(n7734), .A2(n7932), .ZN(n7927) );
  NAND2_X1 U7957 ( .A1(n7733), .A2(n7735), .ZN(n7932) );
  NAND2_X1 U7958 ( .A1(n7933), .A2(n7934), .ZN(n7735) );
  NAND2_X1 U7959 ( .A1(b_30_), .A2(a_27_), .ZN(n7934) );
  INV_X1 U7960 ( .A(n7935), .ZN(n7933) );
  XNOR2_X1 U7961 ( .A(n7936), .B(n7937), .ZN(n7733) );
  XOR2_X1 U7962 ( .A(n7938), .B(n7939), .Z(n7936) );
  NAND2_X1 U7963 ( .A1(b_29_), .A2(a_28_), .ZN(n7938) );
  NAND2_X1 U7964 ( .A1(a_27_), .A2(n7935), .ZN(n7734) );
  NAND2_X1 U7965 ( .A1(n7940), .A2(n7941), .ZN(n7935) );
  NAND3_X1 U7966 ( .A1(a_28_), .A2(n7942), .A3(b_30_), .ZN(n7941) );
  NAND2_X1 U7967 ( .A1(n7713), .A2(n7711), .ZN(n7942) );
  OR2_X1 U7968 ( .A1(n7711), .A2(n7713), .ZN(n7940) );
  AND2_X1 U7969 ( .A1(n7943), .A2(n7944), .ZN(n7713) );
  NAND2_X1 U7970 ( .A1(n7729), .A2(n7945), .ZN(n7944) );
  OR2_X1 U7971 ( .A1(n7730), .A2(n7731), .ZN(n7945) );
  NOR2_X1 U7972 ( .A1(n7274), .A2(n7946), .ZN(n7729) );
  NAND2_X1 U7973 ( .A1(n7731), .A2(n7730), .ZN(n7943) );
  NAND2_X1 U7974 ( .A1(n7947), .A2(n7948), .ZN(n7730) );
  NAND2_X1 U7975 ( .A1(b_28_), .A2(n7949), .ZN(n7948) );
  NAND2_X1 U7976 ( .A1(n7268), .A2(n7950), .ZN(n7949) );
  NAND2_X1 U7977 ( .A1(a_31_), .A2(n7725), .ZN(n7950) );
  NAND2_X1 U7978 ( .A1(b_29_), .A2(n7951), .ZN(n7947) );
  NAND2_X1 U7979 ( .A1(n7272), .A2(n7952), .ZN(n7951) );
  NAND2_X1 U7980 ( .A1(a_30_), .A2(n7953), .ZN(n7952) );
  AND3_X1 U7981 ( .A1(b_29_), .A2(n7954), .A3(b_30_), .ZN(n7731) );
  XNOR2_X1 U7982 ( .A(n7955), .B(n7956), .ZN(n7711) );
  XOR2_X1 U7983 ( .A(n7957), .B(n7958), .Z(n7955) );
  XNOR2_X1 U7984 ( .A(n7959), .B(n7960), .ZN(n7737) );
  NAND2_X1 U7985 ( .A1(n7961), .A2(n7962), .ZN(n7959) );
  XNOR2_X1 U7986 ( .A(n7963), .B(n7964), .ZN(n7688) );
  XNOR2_X1 U7987 ( .A(n7965), .B(n7966), .ZN(n7963) );
  XNOR2_X1 U7988 ( .A(n7967), .B(n7968), .ZN(n7741) );
  XNOR2_X1 U7989 ( .A(n7969), .B(n7970), .ZN(n7967) );
  NOR2_X1 U7990 ( .A1(n7691), .A2(n7725), .ZN(n7970) );
  XNOR2_X1 U7991 ( .A(n7971), .B(n7972), .ZN(n7745) );
  XNOR2_X1 U7992 ( .A(n7973), .B(n7974), .ZN(n7972) );
  XNOR2_X1 U7993 ( .A(n7975), .B(n7976), .ZN(n7749) );
  XOR2_X1 U7994 ( .A(n7977), .B(n7978), .Z(n7976) );
  NAND2_X1 U7995 ( .A1(b_29_), .A2(a_22_), .ZN(n7978) );
  XOR2_X1 U7996 ( .A(n7979), .B(n7980), .Z(n7752) );
  XOR2_X1 U7997 ( .A(n7981), .B(n7982), .Z(n7979) );
  XNOR2_X1 U7998 ( .A(n7983), .B(n7984), .ZN(n7756) );
  XNOR2_X1 U7999 ( .A(n7985), .B(n7986), .ZN(n7983) );
  NOR2_X1 U8000 ( .A1(n7987), .A2(n7725), .ZN(n7986) );
  XNOR2_X1 U8001 ( .A(n7988), .B(n7989), .ZN(n7761) );
  XOR2_X1 U8002 ( .A(n7990), .B(n7991), .Z(n7988) );
  XNOR2_X1 U8003 ( .A(n7992), .B(n7993), .ZN(n7765) );
  XNOR2_X1 U8004 ( .A(n7994), .B(n7995), .ZN(n7992) );
  NOR2_X1 U8005 ( .A1(n7764), .A2(n7725), .ZN(n7995) );
  XNOR2_X1 U8006 ( .A(n7996), .B(n7997), .ZN(n7770) );
  XOR2_X1 U8007 ( .A(n7998), .B(n7999), .Z(n7996) );
  XNOR2_X1 U8008 ( .A(n8000), .B(n8001), .ZN(n7774) );
  XOR2_X1 U8009 ( .A(n8002), .B(n8003), .Z(n8001) );
  NAND2_X1 U8010 ( .A1(b_29_), .A2(a_16_), .ZN(n8003) );
  XOR2_X1 U8011 ( .A(n8004), .B(n8005), .Z(n7779) );
  XNOR2_X1 U8012 ( .A(n8006), .B(n8007), .ZN(n8005) );
  XNOR2_X1 U8013 ( .A(n8008), .B(n8009), .ZN(n7784) );
  XNOR2_X1 U8014 ( .A(n8010), .B(n8011), .ZN(n8008) );
  NOR2_X1 U8015 ( .A1(n7782), .A2(n7725), .ZN(n8011) );
  XOR2_X1 U8016 ( .A(n8012), .B(n8013), .Z(n7787) );
  XOR2_X1 U8017 ( .A(n8014), .B(n8015), .Z(n8012) );
  XNOR2_X1 U8018 ( .A(n8016), .B(n8017), .ZN(n7791) );
  XNOR2_X1 U8019 ( .A(n8018), .B(n8019), .ZN(n8016) );
  NOR2_X1 U8020 ( .A1(n8020), .A2(n7725), .ZN(n8019) );
  XNOR2_X1 U8021 ( .A(n8021), .B(n8022), .ZN(n7796) );
  XNOR2_X1 U8022 ( .A(n8023), .B(n8024), .ZN(n8022) );
  XNOR2_X1 U8023 ( .A(n8025), .B(n8026), .ZN(n7801) );
  XNOR2_X1 U8024 ( .A(n8027), .B(n8028), .ZN(n8025) );
  NOR2_X1 U8025 ( .A1(n7799), .A2(n7725), .ZN(n8028) );
  XOR2_X1 U8026 ( .A(n8029), .B(n8030), .Z(n7804) );
  XOR2_X1 U8027 ( .A(n8031), .B(n8032), .Z(n8029) );
  XOR2_X1 U8028 ( .A(n8033), .B(n8034), .Z(n7808) );
  XOR2_X1 U8029 ( .A(n8035), .B(n8036), .Z(n8033) );
  NOR2_X1 U8030 ( .A1(n8037), .A2(n7725), .ZN(n8036) );
  XOR2_X1 U8031 ( .A(n8038), .B(n8039), .Z(n7813) );
  XNOR2_X1 U8032 ( .A(n8040), .B(n8041), .ZN(n8039) );
  XNOR2_X1 U8033 ( .A(n8042), .B(n8043), .ZN(n7817) );
  XNOR2_X1 U8034 ( .A(n8044), .B(n8045), .ZN(n8042) );
  NAND2_X1 U8035 ( .A1(b_29_), .A2(a_6_), .ZN(n8044) );
  XNOR2_X1 U8036 ( .A(n8046), .B(n8047), .ZN(n7821) );
  XOR2_X1 U8037 ( .A(n8048), .B(n8049), .Z(n8046) );
  XNOR2_X1 U8038 ( .A(n8050), .B(n8051), .ZN(n7824) );
  XNOR2_X1 U8039 ( .A(n8052), .B(n8053), .ZN(n8050) );
  NOR2_X1 U8040 ( .A1(n7398), .A2(n7725), .ZN(n8053) );
  XOR2_X1 U8041 ( .A(n8054), .B(n8055), .Z(n7829) );
  XOR2_X1 U8042 ( .A(n8056), .B(n8057), .Z(n8055) );
  NAND2_X1 U8043 ( .A1(b_29_), .A2(a_3_), .ZN(n8057) );
  XNOR2_X1 U8044 ( .A(n8058), .B(n8059), .ZN(n7833) );
  XNOR2_X1 U8045 ( .A(n8060), .B(n8061), .ZN(n8058) );
  XNOR2_X1 U8046 ( .A(n8062), .B(n8063), .ZN(n7610) );
  XOR2_X1 U8047 ( .A(n8064), .B(n8065), .Z(n8062) );
  NOR2_X1 U8048 ( .A1(n7411), .A2(n7725), .ZN(n8065) );
  XNOR2_X1 U8049 ( .A(n8066), .B(n8067), .ZN(n7606) );
  NAND2_X1 U8050 ( .A1(n8068), .A2(n8069), .ZN(n8066) );
  NAND2_X1 U8051 ( .A1(n8070), .A2(n8071), .ZN(n7431) );
  NAND2_X1 U8052 ( .A1(n7598), .A2(n7600), .ZN(n8071) );
  NAND2_X1 U8053 ( .A1(n8068), .A2(n8072), .ZN(n7600) );
  NAND2_X1 U8054 ( .A1(n8067), .A2(n8069), .ZN(n8072) );
  NAND2_X1 U8055 ( .A1(n8073), .A2(n8074), .ZN(n8069) );
  NAND2_X1 U8056 ( .A1(b_29_), .A2(a_0_), .ZN(n8074) );
  INV_X1 U8057 ( .A(n8075), .ZN(n8073) );
  XOR2_X1 U8058 ( .A(n8076), .B(n8077), .Z(n8067) );
  XOR2_X1 U8059 ( .A(n8078), .B(n8079), .Z(n8076) );
  NAND2_X1 U8060 ( .A1(a_0_), .A2(n8075), .ZN(n8068) );
  NAND2_X1 U8061 ( .A1(n8080), .A2(n8081), .ZN(n8075) );
  NAND3_X1 U8062 ( .A1(a_1_), .A2(n8082), .A3(b_29_), .ZN(n8081) );
  OR2_X1 U8063 ( .A1(n8064), .A2(n8063), .ZN(n8082) );
  NAND2_X1 U8064 ( .A1(n8063), .A2(n8064), .ZN(n8080) );
  NAND2_X1 U8065 ( .A1(n8083), .A2(n8084), .ZN(n8064) );
  NAND2_X1 U8066 ( .A1(n8060), .A2(n8085), .ZN(n8084) );
  NAND2_X1 U8067 ( .A1(n8059), .A2(n8061), .ZN(n8085) );
  NAND2_X1 U8068 ( .A1(n8086), .A2(n8087), .ZN(n8060) );
  NAND3_X1 U8069 ( .A1(a_3_), .A2(n8088), .A3(b_29_), .ZN(n8087) );
  OR2_X1 U8070 ( .A1(n8056), .A2(n8054), .ZN(n8088) );
  NAND2_X1 U8071 ( .A1(n8054), .A2(n8056), .ZN(n8086) );
  NAND2_X1 U8072 ( .A1(n8089), .A2(n8090), .ZN(n8056) );
  NAND3_X1 U8073 ( .A1(a_4_), .A2(n8091), .A3(b_29_), .ZN(n8090) );
  NAND2_X1 U8074 ( .A1(n8052), .A2(n8051), .ZN(n8091) );
  OR2_X1 U8075 ( .A1(n8051), .A2(n8052), .ZN(n8089) );
  AND2_X1 U8076 ( .A1(n8092), .A2(n8093), .ZN(n8052) );
  NAND2_X1 U8077 ( .A1(n8049), .A2(n8094), .ZN(n8093) );
  OR2_X1 U8078 ( .A1(n8048), .A2(n8047), .ZN(n8094) );
  NOR2_X1 U8079 ( .A1(n7725), .A2(n7393), .ZN(n8049) );
  NAND2_X1 U8080 ( .A1(n8047), .A2(n8048), .ZN(n8092) );
  NAND2_X1 U8081 ( .A1(n8095), .A2(n8096), .ZN(n8048) );
  NAND3_X1 U8082 ( .A1(a_6_), .A2(n8097), .A3(b_29_), .ZN(n8096) );
  OR2_X1 U8083 ( .A1(n8045), .A2(n8043), .ZN(n8097) );
  NAND2_X1 U8084 ( .A1(n8043), .A2(n8045), .ZN(n8095) );
  NAND2_X1 U8085 ( .A1(n8098), .A2(n8099), .ZN(n8045) );
  NAND2_X1 U8086 ( .A1(n8041), .A2(n8100), .ZN(n8099) );
  OR2_X1 U8087 ( .A1(n8040), .A2(n8038), .ZN(n8100) );
  NOR2_X1 U8088 ( .A1(n7725), .A2(n7863), .ZN(n8041) );
  NAND2_X1 U8089 ( .A1(n8038), .A2(n8040), .ZN(n8098) );
  NAND2_X1 U8090 ( .A1(n8101), .A2(n8102), .ZN(n8040) );
  NAND3_X1 U8091 ( .A1(a_8_), .A2(n8103), .A3(b_29_), .ZN(n8102) );
  OR2_X1 U8092 ( .A1(n8035), .A2(n8034), .ZN(n8103) );
  NAND2_X1 U8093 ( .A1(n8034), .A2(n8035), .ZN(n8101) );
  NAND2_X1 U8094 ( .A1(n8104), .A2(n8105), .ZN(n8035) );
  NAND2_X1 U8095 ( .A1(n8032), .A2(n8106), .ZN(n8105) );
  OR2_X1 U8096 ( .A1(n8031), .A2(n8030), .ZN(n8106) );
  NOR2_X1 U8097 ( .A1(n7725), .A2(n7870), .ZN(n8032) );
  NAND2_X1 U8098 ( .A1(n8030), .A2(n8031), .ZN(n8104) );
  NAND2_X1 U8099 ( .A1(n8107), .A2(n8108), .ZN(n8031) );
  NAND3_X1 U8100 ( .A1(a_10_), .A2(n8109), .A3(b_29_), .ZN(n8108) );
  NAND2_X1 U8101 ( .A1(n8027), .A2(n8026), .ZN(n8109) );
  OR2_X1 U8102 ( .A1(n8026), .A2(n8027), .ZN(n8107) );
  AND2_X1 U8103 ( .A1(n8110), .A2(n8111), .ZN(n8027) );
  NAND2_X1 U8104 ( .A1(n8024), .A2(n8112), .ZN(n8111) );
  OR2_X1 U8105 ( .A1(n8023), .A2(n8021), .ZN(n8112) );
  NOR2_X1 U8106 ( .A1(n7725), .A2(n7877), .ZN(n8024) );
  NAND2_X1 U8107 ( .A1(n8021), .A2(n8023), .ZN(n8110) );
  NAND2_X1 U8108 ( .A1(n8113), .A2(n8114), .ZN(n8023) );
  NAND3_X1 U8109 ( .A1(a_12_), .A2(n8115), .A3(b_29_), .ZN(n8114) );
  NAND2_X1 U8110 ( .A1(n8018), .A2(n8017), .ZN(n8115) );
  OR2_X1 U8111 ( .A1(n8017), .A2(n8018), .ZN(n8113) );
  AND2_X1 U8112 ( .A1(n8116), .A2(n8117), .ZN(n8018) );
  NAND2_X1 U8113 ( .A1(n8015), .A2(n8118), .ZN(n8117) );
  OR2_X1 U8114 ( .A1(n8014), .A2(n8013), .ZN(n8118) );
  NOR2_X1 U8115 ( .A1(n7725), .A2(n7355), .ZN(n8015) );
  NAND2_X1 U8116 ( .A1(n8013), .A2(n8014), .ZN(n8116) );
  NAND2_X1 U8117 ( .A1(n8119), .A2(n8120), .ZN(n8014) );
  NAND3_X1 U8118 ( .A1(a_14_), .A2(n8121), .A3(b_29_), .ZN(n8120) );
  NAND2_X1 U8119 ( .A1(n8010), .A2(n8009), .ZN(n8121) );
  OR2_X1 U8120 ( .A1(n8009), .A2(n8010), .ZN(n8119) );
  AND2_X1 U8121 ( .A1(n8122), .A2(n8123), .ZN(n8010) );
  NAND2_X1 U8122 ( .A1(n8007), .A2(n8124), .ZN(n8123) );
  OR2_X1 U8123 ( .A1(n8006), .A2(n8004), .ZN(n8124) );
  NOR2_X1 U8124 ( .A1(n7725), .A2(n7346), .ZN(n8007) );
  NAND2_X1 U8125 ( .A1(n8004), .A2(n8006), .ZN(n8122) );
  NAND2_X1 U8126 ( .A1(n8125), .A2(n8126), .ZN(n8006) );
  NAND3_X1 U8127 ( .A1(a_16_), .A2(n8127), .A3(b_29_), .ZN(n8126) );
  OR2_X1 U8128 ( .A1(n8002), .A2(n8000), .ZN(n8127) );
  NAND2_X1 U8129 ( .A1(n8000), .A2(n8002), .ZN(n8125) );
  NAND2_X1 U8130 ( .A1(n8128), .A2(n8129), .ZN(n8002) );
  NAND2_X1 U8131 ( .A1(n7999), .A2(n8130), .ZN(n8129) );
  OR2_X1 U8132 ( .A1(n7998), .A2(n7997), .ZN(n8130) );
  NOR2_X1 U8133 ( .A1(n7725), .A2(n7337), .ZN(n7999) );
  NAND2_X1 U8134 ( .A1(n7997), .A2(n7998), .ZN(n8128) );
  NAND2_X1 U8135 ( .A1(n8131), .A2(n8132), .ZN(n7998) );
  NAND3_X1 U8136 ( .A1(a_18_), .A2(n8133), .A3(b_29_), .ZN(n8132) );
  NAND2_X1 U8137 ( .A1(n7994), .A2(n7993), .ZN(n8133) );
  OR2_X1 U8138 ( .A1(n7993), .A2(n7994), .ZN(n8131) );
  AND2_X1 U8139 ( .A1(n8134), .A2(n8135), .ZN(n7994) );
  NAND2_X1 U8140 ( .A1(n7991), .A2(n8136), .ZN(n8135) );
  OR2_X1 U8141 ( .A1(n7990), .A2(n7989), .ZN(n8136) );
  NOR2_X1 U8142 ( .A1(n7725), .A2(n7902), .ZN(n7991) );
  NAND2_X1 U8143 ( .A1(n7989), .A2(n7990), .ZN(n8134) );
  NAND2_X1 U8144 ( .A1(n8137), .A2(n8138), .ZN(n7990) );
  NAND3_X1 U8145 ( .A1(a_20_), .A2(n8139), .A3(b_29_), .ZN(n8138) );
  NAND2_X1 U8146 ( .A1(n7985), .A2(n7984), .ZN(n8139) );
  OR2_X1 U8147 ( .A1(n7984), .A2(n7985), .ZN(n8137) );
  AND2_X1 U8148 ( .A1(n8140), .A2(n8141), .ZN(n7985) );
  NAND2_X1 U8149 ( .A1(n7982), .A2(n8142), .ZN(n8141) );
  OR2_X1 U8150 ( .A1(n7981), .A2(n7980), .ZN(n8142) );
  NOR2_X1 U8151 ( .A1(n7725), .A2(n7909), .ZN(n7982) );
  NAND2_X1 U8152 ( .A1(n7980), .A2(n7981), .ZN(n8140) );
  NAND2_X1 U8153 ( .A1(n8143), .A2(n8144), .ZN(n7981) );
  NAND3_X1 U8154 ( .A1(a_22_), .A2(n8145), .A3(b_29_), .ZN(n8144) );
  OR2_X1 U8155 ( .A1(n7977), .A2(n7975), .ZN(n8145) );
  NAND2_X1 U8156 ( .A1(n7975), .A2(n7977), .ZN(n8143) );
  NAND2_X1 U8157 ( .A1(n8146), .A2(n8147), .ZN(n7977) );
  NAND2_X1 U8158 ( .A1(n7974), .A2(n8148), .ZN(n8147) );
  OR2_X1 U8159 ( .A1(n7973), .A2(n7971), .ZN(n8148) );
  NOR2_X1 U8160 ( .A1(n7725), .A2(n7916), .ZN(n7974) );
  NAND2_X1 U8161 ( .A1(n7971), .A2(n7973), .ZN(n8146) );
  NAND2_X1 U8162 ( .A1(n8149), .A2(n8150), .ZN(n7973) );
  NAND3_X1 U8163 ( .A1(a_24_), .A2(n8151), .A3(b_29_), .ZN(n8150) );
  NAND2_X1 U8164 ( .A1(n7969), .A2(n7968), .ZN(n8151) );
  OR2_X1 U8165 ( .A1(n7968), .A2(n7969), .ZN(n8149) );
  AND2_X1 U8166 ( .A1(n8152), .A2(n8153), .ZN(n7969) );
  NAND2_X1 U8167 ( .A1(n7966), .A2(n8154), .ZN(n8153) );
  NAND2_X1 U8168 ( .A1(n7965), .A2(n7964), .ZN(n8154) );
  NOR2_X1 U8169 ( .A1(n7725), .A2(n7923), .ZN(n7966) );
  OR2_X1 U8170 ( .A1(n7964), .A2(n7965), .ZN(n8152) );
  AND2_X1 U8171 ( .A1(n7961), .A2(n8155), .ZN(n7965) );
  NAND2_X1 U8172 ( .A1(n7960), .A2(n7962), .ZN(n8155) );
  NAND2_X1 U8173 ( .A1(n8156), .A2(n8157), .ZN(n7962) );
  NAND2_X1 U8174 ( .A1(b_29_), .A2(a_26_), .ZN(n8157) );
  INV_X1 U8175 ( .A(n8158), .ZN(n8156) );
  XNOR2_X1 U8176 ( .A(n8159), .B(n8160), .ZN(n7960) );
  NAND2_X1 U8177 ( .A1(n8161), .A2(n8162), .ZN(n8159) );
  NAND2_X1 U8178 ( .A1(a_26_), .A2(n8158), .ZN(n7961) );
  NAND2_X1 U8179 ( .A1(n7930), .A2(n8163), .ZN(n8158) );
  NAND2_X1 U8180 ( .A1(n7929), .A2(n7931), .ZN(n8163) );
  NAND2_X1 U8181 ( .A1(n8164), .A2(n8165), .ZN(n7931) );
  NAND2_X1 U8182 ( .A1(b_29_), .A2(a_27_), .ZN(n8165) );
  INV_X1 U8183 ( .A(n8166), .ZN(n8164) );
  XNOR2_X1 U8184 ( .A(n8167), .B(n8168), .ZN(n7929) );
  XOR2_X1 U8185 ( .A(n8169), .B(n8170), .Z(n8167) );
  NAND2_X1 U8186 ( .A1(a_27_), .A2(n8166), .ZN(n7930) );
  NAND2_X1 U8187 ( .A1(n8171), .A2(n8172), .ZN(n8166) );
  NAND3_X1 U8188 ( .A1(a_28_), .A2(n8173), .A3(b_29_), .ZN(n8172) );
  NAND2_X1 U8189 ( .A1(n7939), .A2(n7937), .ZN(n8173) );
  OR2_X1 U8190 ( .A1(n7937), .A2(n7939), .ZN(n8171) );
  AND2_X1 U8191 ( .A1(n8174), .A2(n8175), .ZN(n7939) );
  NAND2_X1 U8192 ( .A1(n7956), .A2(n8176), .ZN(n8175) );
  OR2_X1 U8193 ( .A1(n7957), .A2(n7958), .ZN(n8176) );
  NAND2_X1 U8194 ( .A1(n7958), .A2(n7957), .ZN(n8174) );
  NAND2_X1 U8195 ( .A1(n8177), .A2(n8178), .ZN(n7957) );
  NAND2_X1 U8196 ( .A1(b_27_), .A2(n8179), .ZN(n8178) );
  NAND2_X1 U8197 ( .A1(n7268), .A2(n8180), .ZN(n8179) );
  NAND2_X1 U8198 ( .A1(a_31_), .A2(n7953), .ZN(n8180) );
  NAND2_X1 U8199 ( .A1(b_28_), .A2(n8181), .ZN(n8177) );
  NAND2_X1 U8200 ( .A1(n7272), .A2(n8182), .ZN(n8181) );
  NAND2_X1 U8201 ( .A1(a_30_), .A2(n8183), .ZN(n8182) );
  AND3_X1 U8202 ( .A1(b_28_), .A2(n7954), .A3(b_29_), .ZN(n7958) );
  XNOR2_X1 U8203 ( .A(n8184), .B(n8185), .ZN(n7937) );
  XOR2_X1 U8204 ( .A(n8186), .B(n8187), .Z(n8184) );
  XOR2_X1 U8205 ( .A(n8188), .B(n8189), .Z(n7964) );
  NAND2_X1 U8206 ( .A1(n8190), .A2(n8191), .ZN(n8188) );
  XNOR2_X1 U8207 ( .A(n8192), .B(n8193), .ZN(n7968) );
  XOR2_X1 U8208 ( .A(n8194), .B(n8195), .Z(n8192) );
  XOR2_X1 U8209 ( .A(n8196), .B(n8197), .Z(n7971) );
  XOR2_X1 U8210 ( .A(n8198), .B(n8199), .Z(n8196) );
  NOR2_X1 U8211 ( .A1(n7691), .A2(n7953), .ZN(n8199) );
  XNOR2_X1 U8212 ( .A(n8200), .B(n8201), .ZN(n7975) );
  XNOR2_X1 U8213 ( .A(n8202), .B(n8203), .ZN(n8201) );
  XNOR2_X1 U8214 ( .A(n8204), .B(n8205), .ZN(n7980) );
  XNOR2_X1 U8215 ( .A(n8206), .B(n8207), .ZN(n8204) );
  NOR2_X1 U8216 ( .A1(n7312), .A2(n7953), .ZN(n8207) );
  XOR2_X1 U8217 ( .A(n8208), .B(n8209), .Z(n7984) );
  XNOR2_X1 U8218 ( .A(n8210), .B(n8211), .ZN(n8209) );
  XNOR2_X1 U8219 ( .A(n8212), .B(n8213), .ZN(n7989) );
  XNOR2_X1 U8220 ( .A(n8214), .B(n8215), .ZN(n8212) );
  NOR2_X1 U8221 ( .A1(n7987), .A2(n7953), .ZN(n8215) );
  XOR2_X1 U8222 ( .A(n8216), .B(n8217), .Z(n7993) );
  XNOR2_X1 U8223 ( .A(n8218), .B(n8219), .ZN(n8217) );
  XNOR2_X1 U8224 ( .A(n8220), .B(n8221), .ZN(n7997) );
  XNOR2_X1 U8225 ( .A(n8222), .B(n8223), .ZN(n8220) );
  NOR2_X1 U8226 ( .A1(n7764), .A2(n7953), .ZN(n8223) );
  XOR2_X1 U8227 ( .A(n8224), .B(n8225), .Z(n8000) );
  XOR2_X1 U8228 ( .A(n8226), .B(n8227), .Z(n8224) );
  XNOR2_X1 U8229 ( .A(n8228), .B(n8229), .ZN(n8004) );
  XOR2_X1 U8230 ( .A(n8230), .B(n8231), .Z(n8229) );
  NAND2_X1 U8231 ( .A1(b_28_), .A2(a_16_), .ZN(n8231) );
  XOR2_X1 U8232 ( .A(n8232), .B(n8233), .Z(n8009) );
  XNOR2_X1 U8233 ( .A(n8234), .B(n8235), .ZN(n8233) );
  XNOR2_X1 U8234 ( .A(n8236), .B(n8237), .ZN(n8013) );
  XNOR2_X1 U8235 ( .A(n8238), .B(n8239), .ZN(n8236) );
  NOR2_X1 U8236 ( .A1(n7782), .A2(n7953), .ZN(n8239) );
  XNOR2_X1 U8237 ( .A(n8240), .B(n8241), .ZN(n8017) );
  XOR2_X1 U8238 ( .A(n8242), .B(n8243), .Z(n8240) );
  XNOR2_X1 U8239 ( .A(n8244), .B(n8245), .ZN(n8021) );
  XOR2_X1 U8240 ( .A(n8246), .B(n8247), .Z(n8245) );
  NAND2_X1 U8241 ( .A1(b_28_), .A2(a_12_), .ZN(n8247) );
  XOR2_X1 U8242 ( .A(n8248), .B(n8249), .Z(n8026) );
  XNOR2_X1 U8243 ( .A(n8250), .B(n8251), .ZN(n8249) );
  XNOR2_X1 U8244 ( .A(n8252), .B(n8253), .ZN(n8030) );
  XOR2_X1 U8245 ( .A(n8254), .B(n8255), .Z(n8252) );
  NAND2_X1 U8246 ( .A1(b_28_), .A2(a_10_), .ZN(n8254) );
  XNOR2_X1 U8247 ( .A(n8256), .B(n8257), .ZN(n8034) );
  XNOR2_X1 U8248 ( .A(n8258), .B(n8259), .ZN(n8256) );
  XNOR2_X1 U8249 ( .A(n8260), .B(n8261), .ZN(n8038) );
  XOR2_X1 U8250 ( .A(n8262), .B(n8263), .Z(n8261) );
  NAND2_X1 U8251 ( .A1(b_28_), .A2(a_8_), .ZN(n8263) );
  XNOR2_X1 U8252 ( .A(n8264), .B(n8265), .ZN(n8043) );
  XNOR2_X1 U8253 ( .A(n8266), .B(n8267), .ZN(n8265) );
  XNOR2_X1 U8254 ( .A(n8268), .B(n8269), .ZN(n8047) );
  XNOR2_X1 U8255 ( .A(n8270), .B(n8271), .ZN(n8268) );
  NOR2_X1 U8256 ( .A1(n7388), .A2(n7953), .ZN(n8271) );
  XOR2_X1 U8257 ( .A(n8272), .B(n8273), .Z(n8051) );
  XNOR2_X1 U8258 ( .A(n8274), .B(n8275), .ZN(n8273) );
  XNOR2_X1 U8259 ( .A(n8276), .B(n8277), .ZN(n8054) );
  XNOR2_X1 U8260 ( .A(n8278), .B(n8279), .ZN(n8276) );
  NOR2_X1 U8261 ( .A1(n7398), .A2(n7953), .ZN(n8279) );
  OR2_X1 U8262 ( .A1(n8061), .A2(n8059), .ZN(n8083) );
  XOR2_X1 U8263 ( .A(n8280), .B(n8281), .Z(n8059) );
  XOR2_X1 U8264 ( .A(n8282), .B(n8283), .Z(n8281) );
  NAND2_X1 U8265 ( .A1(b_28_), .A2(a_3_), .ZN(n8283) );
  NAND2_X1 U8266 ( .A1(b_29_), .A2(a_2_), .ZN(n8061) );
  XNOR2_X1 U8267 ( .A(n8284), .B(n8285), .ZN(n8063) );
  XNOR2_X1 U8268 ( .A(n8286), .B(n8287), .ZN(n8284) );
  INV_X1 U8269 ( .A(n7608), .ZN(n7598) );
  XOR2_X1 U8270 ( .A(n8288), .B(n8289), .Z(n7608) );
  XNOR2_X1 U8271 ( .A(n8290), .B(n8291), .ZN(n8288) );
  NOR2_X1 U8272 ( .A1(n7613), .A2(n7953), .ZN(n8291) );
  XNOR2_X1 U8273 ( .A(n7602), .B(n7601), .ZN(n8070) );
  NAND2_X1 U8274 ( .A1(n7596), .A2(n7595), .ZN(n7436) );
  NAND2_X1 U8275 ( .A1(n8292), .A2(n8293), .ZN(n7595) );
  NAND2_X1 U8276 ( .A1(n8294), .A2(n8295), .ZN(n8292) );
  OR2_X1 U8277 ( .A1(n7602), .A2(n7601), .ZN(n7596) );
  AND2_X1 U8278 ( .A1(n8296), .A2(n8297), .ZN(n7601) );
  NAND3_X1 U8279 ( .A1(a_0_), .A2(n8298), .A3(b_28_), .ZN(n8297) );
  NAND2_X1 U8280 ( .A1(n8290), .A2(n8289), .ZN(n8298) );
  OR2_X1 U8281 ( .A1(n8289), .A2(n8290), .ZN(n8296) );
  AND2_X1 U8282 ( .A1(n8299), .A2(n8300), .ZN(n8290) );
  NAND2_X1 U8283 ( .A1(n8079), .A2(n8301), .ZN(n8300) );
  OR2_X1 U8284 ( .A1(n8078), .A2(n8077), .ZN(n8301) );
  NOR2_X1 U8285 ( .A1(n7953), .A2(n7411), .ZN(n8079) );
  NAND2_X1 U8286 ( .A1(n8077), .A2(n8078), .ZN(n8299) );
  NAND2_X1 U8287 ( .A1(n8302), .A2(n8303), .ZN(n8078) );
  NAND2_X1 U8288 ( .A1(n8286), .A2(n8304), .ZN(n8303) );
  NAND2_X1 U8289 ( .A1(n8285), .A2(n8287), .ZN(n8304) );
  NAND2_X1 U8290 ( .A1(n8305), .A2(n8306), .ZN(n8286) );
  NAND3_X1 U8291 ( .A1(a_3_), .A2(n8307), .A3(b_28_), .ZN(n8306) );
  OR2_X1 U8292 ( .A1(n8282), .A2(n8280), .ZN(n8307) );
  NAND2_X1 U8293 ( .A1(n8280), .A2(n8282), .ZN(n8305) );
  NAND2_X1 U8294 ( .A1(n8308), .A2(n8309), .ZN(n8282) );
  NAND3_X1 U8295 ( .A1(a_4_), .A2(n8310), .A3(b_28_), .ZN(n8309) );
  NAND2_X1 U8296 ( .A1(n8278), .A2(n8277), .ZN(n8310) );
  OR2_X1 U8297 ( .A1(n8277), .A2(n8278), .ZN(n8308) );
  AND2_X1 U8298 ( .A1(n8311), .A2(n8312), .ZN(n8278) );
  NAND2_X1 U8299 ( .A1(n8275), .A2(n8313), .ZN(n8312) );
  OR2_X1 U8300 ( .A1(n8274), .A2(n8272), .ZN(n8313) );
  NOR2_X1 U8301 ( .A1(n7953), .A2(n7393), .ZN(n8275) );
  NAND2_X1 U8302 ( .A1(n8272), .A2(n8274), .ZN(n8311) );
  NAND2_X1 U8303 ( .A1(n8314), .A2(n8315), .ZN(n8274) );
  NAND3_X1 U8304 ( .A1(a_6_), .A2(n8316), .A3(b_28_), .ZN(n8315) );
  NAND2_X1 U8305 ( .A1(n8270), .A2(n8269), .ZN(n8316) );
  OR2_X1 U8306 ( .A1(n8269), .A2(n8270), .ZN(n8314) );
  AND2_X1 U8307 ( .A1(n8317), .A2(n8318), .ZN(n8270) );
  NAND2_X1 U8308 ( .A1(n8267), .A2(n8319), .ZN(n8318) );
  OR2_X1 U8309 ( .A1(n8266), .A2(n8264), .ZN(n8319) );
  NOR2_X1 U8310 ( .A1(n7953), .A2(n7863), .ZN(n8267) );
  NAND2_X1 U8311 ( .A1(n8264), .A2(n8266), .ZN(n8317) );
  NAND2_X1 U8312 ( .A1(n8320), .A2(n8321), .ZN(n8266) );
  NAND3_X1 U8313 ( .A1(a_8_), .A2(n8322), .A3(b_28_), .ZN(n8321) );
  OR2_X1 U8314 ( .A1(n8262), .A2(n8260), .ZN(n8322) );
  NAND2_X1 U8315 ( .A1(n8260), .A2(n8262), .ZN(n8320) );
  NAND2_X1 U8316 ( .A1(n8323), .A2(n8324), .ZN(n8262) );
  NAND2_X1 U8317 ( .A1(n8259), .A2(n8325), .ZN(n8324) );
  NAND2_X1 U8318 ( .A1(n8258), .A2(n8257), .ZN(n8325) );
  NOR2_X1 U8319 ( .A1(n7953), .A2(n7870), .ZN(n8259) );
  OR2_X1 U8320 ( .A1(n8257), .A2(n8258), .ZN(n8323) );
  AND2_X1 U8321 ( .A1(n8326), .A2(n8327), .ZN(n8258) );
  NAND3_X1 U8322 ( .A1(a_10_), .A2(n8328), .A3(b_28_), .ZN(n8327) );
  NAND2_X1 U8323 ( .A1(n8255), .A2(n8253), .ZN(n8328) );
  OR2_X1 U8324 ( .A1(n8253), .A2(n8255), .ZN(n8326) );
  AND2_X1 U8325 ( .A1(n8329), .A2(n8330), .ZN(n8255) );
  NAND2_X1 U8326 ( .A1(n8251), .A2(n8331), .ZN(n8330) );
  OR2_X1 U8327 ( .A1(n8250), .A2(n8248), .ZN(n8331) );
  NOR2_X1 U8328 ( .A1(n7953), .A2(n7877), .ZN(n8251) );
  NAND2_X1 U8329 ( .A1(n8248), .A2(n8250), .ZN(n8329) );
  NAND2_X1 U8330 ( .A1(n8332), .A2(n8333), .ZN(n8250) );
  NAND3_X1 U8331 ( .A1(a_12_), .A2(n8334), .A3(b_28_), .ZN(n8333) );
  OR2_X1 U8332 ( .A1(n8246), .A2(n8244), .ZN(n8334) );
  NAND2_X1 U8333 ( .A1(n8244), .A2(n8246), .ZN(n8332) );
  NAND2_X1 U8334 ( .A1(n8335), .A2(n8336), .ZN(n8246) );
  NAND2_X1 U8335 ( .A1(n8243), .A2(n8337), .ZN(n8336) );
  OR2_X1 U8336 ( .A1(n8242), .A2(n8241), .ZN(n8337) );
  NOR2_X1 U8337 ( .A1(n7953), .A2(n7355), .ZN(n8243) );
  NAND2_X1 U8338 ( .A1(n8241), .A2(n8242), .ZN(n8335) );
  NAND2_X1 U8339 ( .A1(n8338), .A2(n8339), .ZN(n8242) );
  NAND3_X1 U8340 ( .A1(a_14_), .A2(n8340), .A3(b_28_), .ZN(n8339) );
  NAND2_X1 U8341 ( .A1(n8238), .A2(n8237), .ZN(n8340) );
  OR2_X1 U8342 ( .A1(n8237), .A2(n8238), .ZN(n8338) );
  AND2_X1 U8343 ( .A1(n8341), .A2(n8342), .ZN(n8238) );
  NAND2_X1 U8344 ( .A1(n8235), .A2(n8343), .ZN(n8342) );
  OR2_X1 U8345 ( .A1(n8234), .A2(n8232), .ZN(n8343) );
  NOR2_X1 U8346 ( .A1(n7953), .A2(n7346), .ZN(n8235) );
  NAND2_X1 U8347 ( .A1(n8232), .A2(n8234), .ZN(n8341) );
  NAND2_X1 U8348 ( .A1(n8344), .A2(n8345), .ZN(n8234) );
  NAND3_X1 U8349 ( .A1(a_16_), .A2(n8346), .A3(b_28_), .ZN(n8345) );
  OR2_X1 U8350 ( .A1(n8230), .A2(n8228), .ZN(n8346) );
  NAND2_X1 U8351 ( .A1(n8228), .A2(n8230), .ZN(n8344) );
  NAND2_X1 U8352 ( .A1(n8347), .A2(n8348), .ZN(n8230) );
  NAND2_X1 U8353 ( .A1(n8227), .A2(n8349), .ZN(n8348) );
  OR2_X1 U8354 ( .A1(n8226), .A2(n8225), .ZN(n8349) );
  NOR2_X1 U8355 ( .A1(n7953), .A2(n7337), .ZN(n8227) );
  NAND2_X1 U8356 ( .A1(n8225), .A2(n8226), .ZN(n8347) );
  NAND2_X1 U8357 ( .A1(n8350), .A2(n8351), .ZN(n8226) );
  NAND3_X1 U8358 ( .A1(a_18_), .A2(n8352), .A3(b_28_), .ZN(n8351) );
  NAND2_X1 U8359 ( .A1(n8222), .A2(n8221), .ZN(n8352) );
  OR2_X1 U8360 ( .A1(n8221), .A2(n8222), .ZN(n8350) );
  AND2_X1 U8361 ( .A1(n8353), .A2(n8354), .ZN(n8222) );
  NAND2_X1 U8362 ( .A1(n8219), .A2(n8355), .ZN(n8354) );
  OR2_X1 U8363 ( .A1(n8218), .A2(n8216), .ZN(n8355) );
  NOR2_X1 U8364 ( .A1(n7953), .A2(n7902), .ZN(n8219) );
  NAND2_X1 U8365 ( .A1(n8216), .A2(n8218), .ZN(n8353) );
  NAND2_X1 U8366 ( .A1(n8356), .A2(n8357), .ZN(n8218) );
  NAND3_X1 U8367 ( .A1(a_20_), .A2(n8358), .A3(b_28_), .ZN(n8357) );
  NAND2_X1 U8368 ( .A1(n8214), .A2(n8213), .ZN(n8358) );
  OR2_X1 U8369 ( .A1(n8213), .A2(n8214), .ZN(n8356) );
  AND2_X1 U8370 ( .A1(n8359), .A2(n8360), .ZN(n8214) );
  NAND2_X1 U8371 ( .A1(n8211), .A2(n8361), .ZN(n8360) );
  OR2_X1 U8372 ( .A1(n8210), .A2(n8208), .ZN(n8361) );
  NOR2_X1 U8373 ( .A1(n7953), .A2(n7909), .ZN(n8211) );
  NAND2_X1 U8374 ( .A1(n8208), .A2(n8210), .ZN(n8359) );
  NAND2_X1 U8375 ( .A1(n8362), .A2(n8363), .ZN(n8210) );
  NAND3_X1 U8376 ( .A1(a_22_), .A2(n8364), .A3(b_28_), .ZN(n8363) );
  NAND2_X1 U8377 ( .A1(n8206), .A2(n8205), .ZN(n8364) );
  OR2_X1 U8378 ( .A1(n8205), .A2(n8206), .ZN(n8362) );
  AND2_X1 U8379 ( .A1(n8365), .A2(n8366), .ZN(n8206) );
  NAND2_X1 U8380 ( .A1(n8203), .A2(n8367), .ZN(n8366) );
  OR2_X1 U8381 ( .A1(n8202), .A2(n8200), .ZN(n8367) );
  NOR2_X1 U8382 ( .A1(n7953), .A2(n7916), .ZN(n8203) );
  NAND2_X1 U8383 ( .A1(n8200), .A2(n8202), .ZN(n8365) );
  NAND2_X1 U8384 ( .A1(n8368), .A2(n8369), .ZN(n8202) );
  NAND3_X1 U8385 ( .A1(a_24_), .A2(n8370), .A3(b_28_), .ZN(n8369) );
  OR2_X1 U8386 ( .A1(n8198), .A2(n8197), .ZN(n8370) );
  NAND2_X1 U8387 ( .A1(n8197), .A2(n8198), .ZN(n8368) );
  NAND2_X1 U8388 ( .A1(n8371), .A2(n8372), .ZN(n8198) );
  NAND2_X1 U8389 ( .A1(n8195), .A2(n8373), .ZN(n8372) );
  OR2_X1 U8390 ( .A1(n8194), .A2(n8193), .ZN(n8373) );
  NOR2_X1 U8391 ( .A1(n7953), .A2(n7923), .ZN(n8195) );
  NAND2_X1 U8392 ( .A1(n8193), .A2(n8194), .ZN(n8371) );
  NAND2_X1 U8393 ( .A1(n8190), .A2(n8374), .ZN(n8194) );
  NAND2_X1 U8394 ( .A1(n8189), .A2(n8191), .ZN(n8374) );
  NAND2_X1 U8395 ( .A1(n8375), .A2(n8376), .ZN(n8191) );
  NAND2_X1 U8396 ( .A1(b_28_), .A2(a_26_), .ZN(n8376) );
  INV_X1 U8397 ( .A(n8377), .ZN(n8375) );
  XOR2_X1 U8398 ( .A(n8378), .B(n8379), .Z(n8189) );
  XOR2_X1 U8399 ( .A(n8380), .B(n8381), .Z(n8378) );
  NAND2_X1 U8400 ( .A1(a_26_), .A2(n8377), .ZN(n8190) );
  NAND2_X1 U8401 ( .A1(n8161), .A2(n8382), .ZN(n8377) );
  NAND2_X1 U8402 ( .A1(n8160), .A2(n8162), .ZN(n8382) );
  NAND2_X1 U8403 ( .A1(n8383), .A2(n8384), .ZN(n8162) );
  NAND2_X1 U8404 ( .A1(b_28_), .A2(a_27_), .ZN(n8384) );
  INV_X1 U8405 ( .A(n8385), .ZN(n8383) );
  XNOR2_X1 U8406 ( .A(n8386), .B(n8387), .ZN(n8160) );
  XOR2_X1 U8407 ( .A(n8388), .B(n8389), .Z(n8386) );
  NAND2_X1 U8408 ( .A1(b_27_), .A2(a_28_), .ZN(n8388) );
  NAND2_X1 U8409 ( .A1(a_27_), .A2(n8385), .ZN(n8161) );
  NAND2_X1 U8410 ( .A1(n8390), .A2(n8391), .ZN(n8385) );
  NAND2_X1 U8411 ( .A1(n8392), .A2(n8393), .ZN(n8391) );
  NAND2_X1 U8412 ( .A1(n8170), .A2(n8168), .ZN(n8393) );
  INV_X1 U8413 ( .A(n8169), .ZN(n8392) );
  OR2_X1 U8414 ( .A1(n8168), .A2(n8170), .ZN(n8390) );
  AND2_X1 U8415 ( .A1(n8394), .A2(n8395), .ZN(n8170) );
  NAND2_X1 U8416 ( .A1(n8185), .A2(n8396), .ZN(n8395) );
  OR2_X1 U8417 ( .A1(n8186), .A2(n8187), .ZN(n8396) );
  NOR2_X1 U8418 ( .A1(n7953), .A2(n7946), .ZN(n8185) );
  NAND2_X1 U8419 ( .A1(n8187), .A2(n8186), .ZN(n8394) );
  NAND2_X1 U8420 ( .A1(n8397), .A2(n8398), .ZN(n8186) );
  NAND2_X1 U8421 ( .A1(b_26_), .A2(n8399), .ZN(n8398) );
  NAND2_X1 U8422 ( .A1(n7268), .A2(n8400), .ZN(n8399) );
  NAND2_X1 U8423 ( .A1(a_31_), .A2(n8183), .ZN(n8400) );
  NAND2_X1 U8424 ( .A1(b_27_), .A2(n8401), .ZN(n8397) );
  NAND2_X1 U8425 ( .A1(n7272), .A2(n8402), .ZN(n8401) );
  NAND2_X1 U8426 ( .A1(a_30_), .A2(n8403), .ZN(n8402) );
  AND3_X1 U8427 ( .A1(b_27_), .A2(n7954), .A3(b_28_), .ZN(n8187) );
  XNOR2_X1 U8428 ( .A(n8404), .B(n8405), .ZN(n8168) );
  XOR2_X1 U8429 ( .A(n8406), .B(n8407), .Z(n8404) );
  XNOR2_X1 U8430 ( .A(n8408), .B(n8409), .ZN(n8193) );
  NAND2_X1 U8431 ( .A1(n8410), .A2(n8411), .ZN(n8408) );
  XNOR2_X1 U8432 ( .A(n8412), .B(n8413), .ZN(n8197) );
  XNOR2_X1 U8433 ( .A(n8414), .B(n8415), .ZN(n8412) );
  XNOR2_X1 U8434 ( .A(n8416), .B(n8417), .ZN(n8200) );
  XOR2_X1 U8435 ( .A(n8418), .B(n8419), .Z(n8417) );
  NAND2_X1 U8436 ( .A1(b_27_), .A2(a_24_), .ZN(n8419) );
  XNOR2_X1 U8437 ( .A(n8420), .B(n8421), .ZN(n8205) );
  XOR2_X1 U8438 ( .A(n8422), .B(n8423), .Z(n8420) );
  XNOR2_X1 U8439 ( .A(n8424), .B(n8425), .ZN(n8208) );
  XNOR2_X1 U8440 ( .A(n8426), .B(n8427), .ZN(n8424) );
  NOR2_X1 U8441 ( .A1(n7312), .A2(n8183), .ZN(n8427) );
  XNOR2_X1 U8442 ( .A(n8428), .B(n8429), .ZN(n8213) );
  XOR2_X1 U8443 ( .A(n8430), .B(n8431), .Z(n8428) );
  XNOR2_X1 U8444 ( .A(n8432), .B(n8433), .ZN(n8216) );
  XNOR2_X1 U8445 ( .A(n8434), .B(n8435), .ZN(n8432) );
  NOR2_X1 U8446 ( .A1(n7987), .A2(n8183), .ZN(n8435) );
  XOR2_X1 U8447 ( .A(n8436), .B(n8437), .Z(n8221) );
  XNOR2_X1 U8448 ( .A(n8438), .B(n8439), .ZN(n8437) );
  XNOR2_X1 U8449 ( .A(n8440), .B(n8441), .ZN(n8225) );
  XNOR2_X1 U8450 ( .A(n8442), .B(n8443), .ZN(n8440) );
  NOR2_X1 U8451 ( .A1(n7764), .A2(n8183), .ZN(n8443) );
  XOR2_X1 U8452 ( .A(n8444), .B(n8445), .Z(n8228) );
  XOR2_X1 U8453 ( .A(n8446), .B(n8447), .Z(n8444) );
  XNOR2_X1 U8454 ( .A(n8448), .B(n8449), .ZN(n8232) );
  XNOR2_X1 U8455 ( .A(n8450), .B(n8451), .ZN(n8448) );
  NOR2_X1 U8456 ( .A1(n7773), .A2(n8183), .ZN(n8451) );
  XOR2_X1 U8457 ( .A(n8452), .B(n8453), .Z(n8237) );
  XNOR2_X1 U8458 ( .A(n8454), .B(n8455), .ZN(n8453) );
  XNOR2_X1 U8459 ( .A(n8456), .B(n8457), .ZN(n8241) );
  XNOR2_X1 U8460 ( .A(n8458), .B(n8459), .ZN(n8456) );
  NOR2_X1 U8461 ( .A1(n7782), .A2(n8183), .ZN(n8459) );
  XNOR2_X1 U8462 ( .A(n8460), .B(n8461), .ZN(n8244) );
  XNOR2_X1 U8463 ( .A(n8462), .B(n8463), .ZN(n8460) );
  XNOR2_X1 U8464 ( .A(n8464), .B(n8465), .ZN(n8248) );
  XOR2_X1 U8465 ( .A(n8466), .B(n8467), .Z(n8465) );
  NAND2_X1 U8466 ( .A1(b_27_), .A2(a_12_), .ZN(n8467) );
  XOR2_X1 U8467 ( .A(n8468), .B(n8469), .Z(n8253) );
  XNOR2_X1 U8468 ( .A(n8470), .B(n8471), .ZN(n8469) );
  XNOR2_X1 U8469 ( .A(n8472), .B(n8473), .ZN(n8257) );
  XOR2_X1 U8470 ( .A(n8474), .B(n8475), .Z(n8472) );
  NOR2_X1 U8471 ( .A1(n7799), .A2(n8183), .ZN(n8475) );
  XOR2_X1 U8472 ( .A(n8476), .B(n8477), .Z(n8260) );
  XOR2_X1 U8473 ( .A(n8478), .B(n8479), .Z(n8476) );
  XOR2_X1 U8474 ( .A(n8480), .B(n8481), .Z(n8264) );
  XOR2_X1 U8475 ( .A(n8482), .B(n8483), .Z(n8480) );
  NOR2_X1 U8476 ( .A1(n8037), .A2(n8183), .ZN(n8483) );
  XOR2_X1 U8477 ( .A(n8484), .B(n8485), .Z(n8269) );
  XOR2_X1 U8478 ( .A(n8486), .B(n8487), .Z(n8485) );
  NAND2_X1 U8479 ( .A1(b_27_), .A2(a_7_), .ZN(n8487) );
  XNOR2_X1 U8480 ( .A(n8488), .B(n8489), .ZN(n8272) );
  XNOR2_X1 U8481 ( .A(n8490), .B(n8491), .ZN(n8488) );
  NOR2_X1 U8482 ( .A1(n7388), .A2(n8183), .ZN(n8491) );
  XNOR2_X1 U8483 ( .A(n8492), .B(n8493), .ZN(n8277) );
  XOR2_X1 U8484 ( .A(n8494), .B(n8495), .Z(n8492) );
  XNOR2_X1 U8485 ( .A(n8496), .B(n8497), .ZN(n8280) );
  XNOR2_X1 U8486 ( .A(n8498), .B(n8499), .ZN(n8496) );
  NOR2_X1 U8487 ( .A1(n7398), .A2(n8183), .ZN(n8499) );
  OR2_X1 U8488 ( .A1(n8287), .A2(n8285), .ZN(n8302) );
  XOR2_X1 U8489 ( .A(n8500), .B(n8501), .Z(n8285) );
  NAND2_X1 U8490 ( .A1(n8502), .A2(n8503), .ZN(n8500) );
  NAND2_X1 U8491 ( .A1(b_28_), .A2(a_2_), .ZN(n8287) );
  XNOR2_X1 U8492 ( .A(n8504), .B(n8505), .ZN(n8077) );
  NAND2_X1 U8493 ( .A1(n8506), .A2(n8507), .ZN(n8504) );
  XNOR2_X1 U8494 ( .A(n8508), .B(n8509), .ZN(n8289) );
  XOR2_X1 U8495 ( .A(n8510), .B(n8511), .Z(n8508) );
  NOR2_X1 U8496 ( .A1(n7411), .A2(n8183), .ZN(n8511) );
  XNOR2_X1 U8497 ( .A(n8512), .B(n8513), .ZN(n7602) );
  XNOR2_X1 U8498 ( .A(n8514), .B(n8515), .ZN(n8513) );
  NAND2_X1 U8499 ( .A1(n8516), .A2(n8293), .ZN(n7439) );
  INV_X1 U8500 ( .A(n8517), .ZN(n8293) );
  XOR2_X1 U8501 ( .A(n7592), .B(n8518), .Z(n8516) );
  NAND2_X1 U8502 ( .A1(n8519), .A2(n8517), .ZN(n7440) );
  NOR2_X1 U8503 ( .A1(n8295), .A2(n8294), .ZN(n8517) );
  XOR2_X1 U8504 ( .A(n8520), .B(n8521), .Z(n8294) );
  XOR2_X1 U8505 ( .A(n8522), .B(n8523), .Z(n8521) );
  NAND2_X1 U8506 ( .A1(b_26_), .A2(a_0_), .ZN(n8523) );
  NAND2_X1 U8507 ( .A1(n8524), .A2(n8525), .ZN(n8295) );
  NAND2_X1 U8508 ( .A1(n8514), .A2(n8526), .ZN(n8525) );
  OR2_X1 U8509 ( .A1(n8515), .A2(n8512), .ZN(n8526) );
  AND2_X1 U8510 ( .A1(n8527), .A2(n8528), .ZN(n8514) );
  NAND3_X1 U8511 ( .A1(a_1_), .A2(n8529), .A3(b_27_), .ZN(n8528) );
  OR2_X1 U8512 ( .A1(n8510), .A2(n8509), .ZN(n8529) );
  NAND2_X1 U8513 ( .A1(n8509), .A2(n8510), .ZN(n8527) );
  NAND2_X1 U8514 ( .A1(n8506), .A2(n8530), .ZN(n8510) );
  NAND2_X1 U8515 ( .A1(n8505), .A2(n8507), .ZN(n8530) );
  NAND2_X1 U8516 ( .A1(n8531), .A2(n8532), .ZN(n8507) );
  NAND2_X1 U8517 ( .A1(b_27_), .A2(a_2_), .ZN(n8532) );
  INV_X1 U8518 ( .A(n8533), .ZN(n8531) );
  XNOR2_X1 U8519 ( .A(n8534), .B(n8535), .ZN(n8505) );
  XNOR2_X1 U8520 ( .A(n8536), .B(n8537), .ZN(n8534) );
  NOR2_X1 U8521 ( .A1(n7850), .A2(n8403), .ZN(n8537) );
  NAND2_X1 U8522 ( .A1(a_2_), .A2(n8533), .ZN(n8506) );
  NAND2_X1 U8523 ( .A1(n8502), .A2(n8538), .ZN(n8533) );
  NAND2_X1 U8524 ( .A1(n8501), .A2(n8503), .ZN(n8538) );
  NAND2_X1 U8525 ( .A1(n8539), .A2(n8540), .ZN(n8503) );
  NAND2_X1 U8526 ( .A1(b_27_), .A2(a_3_), .ZN(n8540) );
  INV_X1 U8527 ( .A(n8541), .ZN(n8539) );
  XNOR2_X1 U8528 ( .A(n8542), .B(n8543), .ZN(n8501) );
  XNOR2_X1 U8529 ( .A(n8544), .B(n8545), .ZN(n8543) );
  NAND2_X1 U8530 ( .A1(a_3_), .A2(n8541), .ZN(n8502) );
  NAND2_X1 U8531 ( .A1(n8546), .A2(n8547), .ZN(n8541) );
  NAND3_X1 U8532 ( .A1(a_4_), .A2(n8548), .A3(b_27_), .ZN(n8547) );
  NAND2_X1 U8533 ( .A1(n8498), .A2(n8497), .ZN(n8548) );
  OR2_X1 U8534 ( .A1(n8497), .A2(n8498), .ZN(n8546) );
  AND2_X1 U8535 ( .A1(n8549), .A2(n8550), .ZN(n8498) );
  NAND2_X1 U8536 ( .A1(n8495), .A2(n8551), .ZN(n8550) );
  OR2_X1 U8537 ( .A1(n8494), .A2(n8493), .ZN(n8551) );
  NOR2_X1 U8538 ( .A1(n8183), .A2(n7393), .ZN(n8495) );
  NAND2_X1 U8539 ( .A1(n8493), .A2(n8494), .ZN(n8549) );
  NAND2_X1 U8540 ( .A1(n8552), .A2(n8553), .ZN(n8494) );
  NAND3_X1 U8541 ( .A1(a_6_), .A2(n8554), .A3(b_27_), .ZN(n8553) );
  NAND2_X1 U8542 ( .A1(n8490), .A2(n8489), .ZN(n8554) );
  OR2_X1 U8543 ( .A1(n8489), .A2(n8490), .ZN(n8552) );
  AND2_X1 U8544 ( .A1(n8555), .A2(n8556), .ZN(n8490) );
  NAND3_X1 U8545 ( .A1(a_7_), .A2(n8557), .A3(b_27_), .ZN(n8556) );
  OR2_X1 U8546 ( .A1(n8486), .A2(n8484), .ZN(n8557) );
  NAND2_X1 U8547 ( .A1(n8484), .A2(n8486), .ZN(n8555) );
  NAND2_X1 U8548 ( .A1(n8558), .A2(n8559), .ZN(n8486) );
  NAND3_X1 U8549 ( .A1(a_8_), .A2(n8560), .A3(b_27_), .ZN(n8559) );
  OR2_X1 U8550 ( .A1(n8482), .A2(n8481), .ZN(n8560) );
  NAND2_X1 U8551 ( .A1(n8481), .A2(n8482), .ZN(n8558) );
  NAND2_X1 U8552 ( .A1(n8561), .A2(n8562), .ZN(n8482) );
  NAND2_X1 U8553 ( .A1(n8479), .A2(n8563), .ZN(n8562) );
  OR2_X1 U8554 ( .A1(n8478), .A2(n8477), .ZN(n8563) );
  NOR2_X1 U8555 ( .A1(n8183), .A2(n7870), .ZN(n8479) );
  NAND2_X1 U8556 ( .A1(n8477), .A2(n8478), .ZN(n8561) );
  NAND2_X1 U8557 ( .A1(n8564), .A2(n8565), .ZN(n8478) );
  NAND3_X1 U8558 ( .A1(a_10_), .A2(n8566), .A3(b_27_), .ZN(n8565) );
  OR2_X1 U8559 ( .A1(n8474), .A2(n8473), .ZN(n8566) );
  NAND2_X1 U8560 ( .A1(n8473), .A2(n8474), .ZN(n8564) );
  NAND2_X1 U8561 ( .A1(n8567), .A2(n8568), .ZN(n8474) );
  NAND2_X1 U8562 ( .A1(n8471), .A2(n8569), .ZN(n8568) );
  OR2_X1 U8563 ( .A1(n8470), .A2(n8468), .ZN(n8569) );
  NOR2_X1 U8564 ( .A1(n8183), .A2(n7877), .ZN(n8471) );
  NAND2_X1 U8565 ( .A1(n8468), .A2(n8470), .ZN(n8567) );
  NAND2_X1 U8566 ( .A1(n8570), .A2(n8571), .ZN(n8470) );
  NAND3_X1 U8567 ( .A1(a_12_), .A2(n8572), .A3(b_27_), .ZN(n8571) );
  OR2_X1 U8568 ( .A1(n8466), .A2(n8464), .ZN(n8572) );
  NAND2_X1 U8569 ( .A1(n8464), .A2(n8466), .ZN(n8570) );
  NAND2_X1 U8570 ( .A1(n8573), .A2(n8574), .ZN(n8466) );
  NAND2_X1 U8571 ( .A1(n8463), .A2(n8575), .ZN(n8574) );
  NAND2_X1 U8572 ( .A1(n8462), .A2(n8461), .ZN(n8575) );
  NOR2_X1 U8573 ( .A1(n8183), .A2(n7355), .ZN(n8463) );
  OR2_X1 U8574 ( .A1(n8461), .A2(n8462), .ZN(n8573) );
  AND2_X1 U8575 ( .A1(n8576), .A2(n8577), .ZN(n8462) );
  NAND3_X1 U8576 ( .A1(a_14_), .A2(n8578), .A3(b_27_), .ZN(n8577) );
  NAND2_X1 U8577 ( .A1(n8458), .A2(n8457), .ZN(n8578) );
  OR2_X1 U8578 ( .A1(n8457), .A2(n8458), .ZN(n8576) );
  AND2_X1 U8579 ( .A1(n8579), .A2(n8580), .ZN(n8458) );
  NAND2_X1 U8580 ( .A1(n8455), .A2(n8581), .ZN(n8580) );
  OR2_X1 U8581 ( .A1(n8454), .A2(n8452), .ZN(n8581) );
  NOR2_X1 U8582 ( .A1(n8183), .A2(n7346), .ZN(n8455) );
  NAND2_X1 U8583 ( .A1(n8452), .A2(n8454), .ZN(n8579) );
  NAND2_X1 U8584 ( .A1(n8582), .A2(n8583), .ZN(n8454) );
  NAND3_X1 U8585 ( .A1(a_16_), .A2(n8584), .A3(b_27_), .ZN(n8583) );
  NAND2_X1 U8586 ( .A1(n8450), .A2(n8449), .ZN(n8584) );
  OR2_X1 U8587 ( .A1(n8449), .A2(n8450), .ZN(n8582) );
  AND2_X1 U8588 ( .A1(n8585), .A2(n8586), .ZN(n8450) );
  NAND2_X1 U8589 ( .A1(n8447), .A2(n8587), .ZN(n8586) );
  OR2_X1 U8590 ( .A1(n8446), .A2(n8445), .ZN(n8587) );
  NOR2_X1 U8591 ( .A1(n8183), .A2(n7337), .ZN(n8447) );
  NAND2_X1 U8592 ( .A1(n8445), .A2(n8446), .ZN(n8585) );
  NAND2_X1 U8593 ( .A1(n8588), .A2(n8589), .ZN(n8446) );
  NAND3_X1 U8594 ( .A1(a_18_), .A2(n8590), .A3(b_27_), .ZN(n8589) );
  NAND2_X1 U8595 ( .A1(n8442), .A2(n8441), .ZN(n8590) );
  OR2_X1 U8596 ( .A1(n8441), .A2(n8442), .ZN(n8588) );
  AND2_X1 U8597 ( .A1(n8591), .A2(n8592), .ZN(n8442) );
  NAND2_X1 U8598 ( .A1(n8439), .A2(n8593), .ZN(n8592) );
  OR2_X1 U8599 ( .A1(n8438), .A2(n8436), .ZN(n8593) );
  NOR2_X1 U8600 ( .A1(n8183), .A2(n7902), .ZN(n8439) );
  NAND2_X1 U8601 ( .A1(n8436), .A2(n8438), .ZN(n8591) );
  NAND2_X1 U8602 ( .A1(n8594), .A2(n8595), .ZN(n8438) );
  NAND3_X1 U8603 ( .A1(a_20_), .A2(n8596), .A3(b_27_), .ZN(n8595) );
  NAND2_X1 U8604 ( .A1(n8434), .A2(n8433), .ZN(n8596) );
  OR2_X1 U8605 ( .A1(n8433), .A2(n8434), .ZN(n8594) );
  AND2_X1 U8606 ( .A1(n8597), .A2(n8598), .ZN(n8434) );
  NAND2_X1 U8607 ( .A1(n8431), .A2(n8599), .ZN(n8598) );
  OR2_X1 U8608 ( .A1(n8430), .A2(n8429), .ZN(n8599) );
  NOR2_X1 U8609 ( .A1(n8183), .A2(n7909), .ZN(n8431) );
  NAND2_X1 U8610 ( .A1(n8429), .A2(n8430), .ZN(n8597) );
  NAND2_X1 U8611 ( .A1(n8600), .A2(n8601), .ZN(n8430) );
  NAND3_X1 U8612 ( .A1(a_22_), .A2(n8602), .A3(b_27_), .ZN(n8601) );
  NAND2_X1 U8613 ( .A1(n8426), .A2(n8425), .ZN(n8602) );
  OR2_X1 U8614 ( .A1(n8425), .A2(n8426), .ZN(n8600) );
  AND2_X1 U8615 ( .A1(n8603), .A2(n8604), .ZN(n8426) );
  NAND2_X1 U8616 ( .A1(n8423), .A2(n8605), .ZN(n8604) );
  OR2_X1 U8617 ( .A1(n8422), .A2(n8421), .ZN(n8605) );
  NOR2_X1 U8618 ( .A1(n8183), .A2(n7916), .ZN(n8423) );
  NAND2_X1 U8619 ( .A1(n8421), .A2(n8422), .ZN(n8603) );
  NAND2_X1 U8620 ( .A1(n8606), .A2(n8607), .ZN(n8422) );
  NAND3_X1 U8621 ( .A1(a_24_), .A2(n8608), .A3(b_27_), .ZN(n8607) );
  OR2_X1 U8622 ( .A1(n8418), .A2(n8416), .ZN(n8608) );
  NAND2_X1 U8623 ( .A1(n8416), .A2(n8418), .ZN(n8606) );
  NAND2_X1 U8624 ( .A1(n8609), .A2(n8610), .ZN(n8418) );
  NAND2_X1 U8625 ( .A1(n8415), .A2(n8611), .ZN(n8610) );
  NAND2_X1 U8626 ( .A1(n8414), .A2(n8413), .ZN(n8611) );
  NOR2_X1 U8627 ( .A1(n8183), .A2(n7923), .ZN(n8415) );
  OR2_X1 U8628 ( .A1(n8413), .A2(n8414), .ZN(n8609) );
  AND2_X1 U8629 ( .A1(n8410), .A2(n8612), .ZN(n8414) );
  NAND2_X1 U8630 ( .A1(n8409), .A2(n8411), .ZN(n8612) );
  NAND2_X1 U8631 ( .A1(n8613), .A2(n8614), .ZN(n8411) );
  NAND2_X1 U8632 ( .A1(b_27_), .A2(a_26_), .ZN(n8614) );
  INV_X1 U8633 ( .A(n8615), .ZN(n8613) );
  XNOR2_X1 U8634 ( .A(n8616), .B(n8617), .ZN(n8409) );
  NAND2_X1 U8635 ( .A1(n8618), .A2(n8619), .ZN(n8616) );
  NAND2_X1 U8636 ( .A1(a_26_), .A2(n8615), .ZN(n8410) );
  NAND2_X1 U8637 ( .A1(n8620), .A2(n8621), .ZN(n8615) );
  NAND2_X1 U8638 ( .A1(n8379), .A2(n8622), .ZN(n8621) );
  OR2_X1 U8639 ( .A1(n8380), .A2(n8381), .ZN(n8622) );
  XNOR2_X1 U8640 ( .A(n8623), .B(n8624), .ZN(n8379) );
  XOR2_X1 U8641 ( .A(n8625), .B(n8626), .Z(n8623) );
  NAND2_X1 U8642 ( .A1(b_26_), .A2(a_28_), .ZN(n8625) );
  NAND2_X1 U8643 ( .A1(n8381), .A2(n8380), .ZN(n8620) );
  NAND2_X1 U8644 ( .A1(n8627), .A2(n8628), .ZN(n8380) );
  NAND3_X1 U8645 ( .A1(a_28_), .A2(n8629), .A3(b_27_), .ZN(n8628) );
  NAND2_X1 U8646 ( .A1(n8389), .A2(n8387), .ZN(n8629) );
  OR2_X1 U8647 ( .A1(n8387), .A2(n8389), .ZN(n8627) );
  AND2_X1 U8648 ( .A1(n8630), .A2(n8631), .ZN(n8389) );
  NAND2_X1 U8649 ( .A1(n8405), .A2(n8632), .ZN(n8631) );
  OR2_X1 U8650 ( .A1(n8406), .A2(n8407), .ZN(n8632) );
  NOR2_X1 U8651 ( .A1(n8183), .A2(n7946), .ZN(n8405) );
  NAND2_X1 U8652 ( .A1(n8407), .A2(n8406), .ZN(n8630) );
  NAND2_X1 U8653 ( .A1(n8633), .A2(n8634), .ZN(n8406) );
  NAND2_X1 U8654 ( .A1(b_25_), .A2(n8635), .ZN(n8634) );
  NAND2_X1 U8655 ( .A1(n7268), .A2(n8636), .ZN(n8635) );
  NAND2_X1 U8656 ( .A1(a_31_), .A2(n8403), .ZN(n8636) );
  NAND2_X1 U8657 ( .A1(b_26_), .A2(n8637), .ZN(n8633) );
  NAND2_X1 U8658 ( .A1(n7272), .A2(n8638), .ZN(n8637) );
  NAND2_X1 U8659 ( .A1(a_30_), .A2(n8639), .ZN(n8638) );
  AND3_X1 U8660 ( .A1(b_26_), .A2(n7954), .A3(b_27_), .ZN(n8407) );
  XNOR2_X1 U8661 ( .A(n8640), .B(n8641), .ZN(n8387) );
  XOR2_X1 U8662 ( .A(n8642), .B(n8643), .Z(n8640) );
  XNOR2_X1 U8663 ( .A(n8644), .B(n8645), .ZN(n8413) );
  XOR2_X1 U8664 ( .A(n8646), .B(n8647), .Z(n8644) );
  XNOR2_X1 U8665 ( .A(n8648), .B(n8649), .ZN(n8416) );
  XNOR2_X1 U8666 ( .A(n8650), .B(n8651), .ZN(n8649) );
  XNOR2_X1 U8667 ( .A(n8652), .B(n8653), .ZN(n8421) );
  XNOR2_X1 U8668 ( .A(n8654), .B(n8655), .ZN(n8652) );
  NOR2_X1 U8669 ( .A1(n7691), .A2(n8403), .ZN(n8655) );
  XOR2_X1 U8670 ( .A(n8656), .B(n8657), .Z(n8425) );
  XNOR2_X1 U8671 ( .A(n8658), .B(n8659), .ZN(n8657) );
  XNOR2_X1 U8672 ( .A(n8660), .B(n8661), .ZN(n8429) );
  XOR2_X1 U8673 ( .A(n8662), .B(n8663), .Z(n8661) );
  NAND2_X1 U8674 ( .A1(b_26_), .A2(a_22_), .ZN(n8663) );
  XNOR2_X1 U8675 ( .A(n8664), .B(n8665), .ZN(n8433) );
  XOR2_X1 U8676 ( .A(n8666), .B(n8667), .Z(n8664) );
  XNOR2_X1 U8677 ( .A(n8668), .B(n8669), .ZN(n8436) );
  XNOR2_X1 U8678 ( .A(n8670), .B(n8671), .ZN(n8668) );
  NOR2_X1 U8679 ( .A1(n7987), .A2(n8403), .ZN(n8671) );
  XOR2_X1 U8680 ( .A(n8672), .B(n8673), .Z(n8441) );
  XNOR2_X1 U8681 ( .A(n8674), .B(n8675), .ZN(n8673) );
  XNOR2_X1 U8682 ( .A(n8676), .B(n8677), .ZN(n8445) );
  XNOR2_X1 U8683 ( .A(n8678), .B(n8679), .ZN(n8676) );
  NOR2_X1 U8684 ( .A1(n7764), .A2(n8403), .ZN(n8679) );
  XNOR2_X1 U8685 ( .A(n8680), .B(n8681), .ZN(n8449) );
  XOR2_X1 U8686 ( .A(n8682), .B(n8683), .Z(n8680) );
  XNOR2_X1 U8687 ( .A(n8684), .B(n8685), .ZN(n8452) );
  XOR2_X1 U8688 ( .A(n8686), .B(n8687), .Z(n8685) );
  NAND2_X1 U8689 ( .A1(b_26_), .A2(a_16_), .ZN(n8687) );
  XOR2_X1 U8690 ( .A(n8688), .B(n8689), .Z(n8457) );
  XNOR2_X1 U8691 ( .A(n8690), .B(n8691), .ZN(n8689) );
  XNOR2_X1 U8692 ( .A(n8692), .B(n8693), .ZN(n8461) );
  XOR2_X1 U8693 ( .A(n8694), .B(n8695), .Z(n8692) );
  NOR2_X1 U8694 ( .A1(n7782), .A2(n8403), .ZN(n8695) );
  XOR2_X1 U8695 ( .A(n8696), .B(n8697), .Z(n8464) );
  XOR2_X1 U8696 ( .A(n8698), .B(n8699), .Z(n8696) );
  XNOR2_X1 U8697 ( .A(n8700), .B(n8701), .ZN(n8468) );
  XNOR2_X1 U8698 ( .A(n8702), .B(n8703), .ZN(n8700) );
  NOR2_X1 U8699 ( .A1(n8020), .A2(n8403), .ZN(n8703) );
  XNOR2_X1 U8700 ( .A(n8704), .B(n8705), .ZN(n8473) );
  XNOR2_X1 U8701 ( .A(n8706), .B(n8707), .ZN(n8705) );
  XNOR2_X1 U8702 ( .A(n8708), .B(n8709), .ZN(n8477) );
  XNOR2_X1 U8703 ( .A(n8710), .B(n8711), .ZN(n8708) );
  NOR2_X1 U8704 ( .A1(n7799), .A2(n8403), .ZN(n8711) );
  XNOR2_X1 U8705 ( .A(n8712), .B(n8713), .ZN(n8481) );
  XNOR2_X1 U8706 ( .A(n8714), .B(n8715), .ZN(n8712) );
  XNOR2_X1 U8707 ( .A(n8716), .B(n8717), .ZN(n8484) );
  XOR2_X1 U8708 ( .A(n8718), .B(n8719), .Z(n8717) );
  NAND2_X1 U8709 ( .A1(b_26_), .A2(a_8_), .ZN(n8719) );
  XOR2_X1 U8710 ( .A(n8720), .B(n8721), .Z(n8489) );
  NAND2_X1 U8711 ( .A1(n8722), .A2(n8723), .ZN(n8720) );
  XNOR2_X1 U8712 ( .A(n8724), .B(n8725), .ZN(n8493) );
  XOR2_X1 U8713 ( .A(n8726), .B(n8727), .Z(n8724) );
  NAND2_X1 U8714 ( .A1(b_26_), .A2(a_6_), .ZN(n8726) );
  XOR2_X1 U8715 ( .A(n8728), .B(n8729), .Z(n8497) );
  XOR2_X1 U8716 ( .A(n8730), .B(n8731), .Z(n8729) );
  NAND2_X1 U8717 ( .A1(b_26_), .A2(a_5_), .ZN(n8731) );
  XNOR2_X1 U8718 ( .A(n8732), .B(n8733), .ZN(n8509) );
  XNOR2_X1 U8719 ( .A(n8734), .B(n8735), .ZN(n8733) );
  NAND2_X1 U8720 ( .A1(n8512), .A2(n8515), .ZN(n8524) );
  NAND2_X1 U8721 ( .A1(b_27_), .A2(a_0_), .ZN(n8515) );
  XOR2_X1 U8722 ( .A(n8736), .B(n8737), .Z(n8512) );
  XNOR2_X1 U8723 ( .A(n8738), .B(n8739), .ZN(n8736) );
  XOR2_X1 U8724 ( .A(n7592), .B(n7591), .Z(n8519) );
  NAND4_X1 U8725 ( .A1(n7591), .A2(n7590), .A3(n7592), .A4(n7585), .ZN(n7443)
         );
  INV_X1 U8726 ( .A(n8740), .ZN(n7585) );
  NAND2_X1 U8727 ( .A1(n8741), .A2(n8742), .ZN(n7592) );
  NAND3_X1 U8728 ( .A1(a_0_), .A2(n8743), .A3(b_26_), .ZN(n8742) );
  OR2_X1 U8729 ( .A1(n8522), .A2(n8520), .ZN(n8743) );
  NAND2_X1 U8730 ( .A1(n8520), .A2(n8522), .ZN(n8741) );
  NAND2_X1 U8731 ( .A1(n8744), .A2(n8745), .ZN(n8522) );
  NAND2_X1 U8732 ( .A1(n8739), .A2(n8746), .ZN(n8745) );
  NAND2_X1 U8733 ( .A1(n8738), .A2(n8737), .ZN(n8746) );
  NOR2_X1 U8734 ( .A1(n8403), .A2(n7411), .ZN(n8739) );
  OR2_X1 U8735 ( .A1(n8737), .A2(n8738), .ZN(n8744) );
  AND2_X1 U8736 ( .A1(n8747), .A2(n8748), .ZN(n8738) );
  NAND2_X1 U8737 ( .A1(n8735), .A2(n8749), .ZN(n8748) );
  OR2_X1 U8738 ( .A1(n8734), .A2(n8732), .ZN(n8749) );
  NOR2_X1 U8739 ( .A1(n8403), .A2(n7832), .ZN(n8735) );
  NAND2_X1 U8740 ( .A1(n8732), .A2(n8734), .ZN(n8747) );
  NAND2_X1 U8741 ( .A1(n8750), .A2(n8751), .ZN(n8734) );
  NAND3_X1 U8742 ( .A1(a_3_), .A2(n8752), .A3(b_26_), .ZN(n8751) );
  NAND2_X1 U8743 ( .A1(n8536), .A2(n8535), .ZN(n8752) );
  OR2_X1 U8744 ( .A1(n8535), .A2(n8536), .ZN(n8750) );
  AND2_X1 U8745 ( .A1(n8753), .A2(n8754), .ZN(n8536) );
  NAND2_X1 U8746 ( .A1(n8545), .A2(n8755), .ZN(n8754) );
  OR2_X1 U8747 ( .A1(n8544), .A2(n8542), .ZN(n8755) );
  NOR2_X1 U8748 ( .A1(n8403), .A2(n7398), .ZN(n8545) );
  NAND2_X1 U8749 ( .A1(n8542), .A2(n8544), .ZN(n8753) );
  NAND2_X1 U8750 ( .A1(n8756), .A2(n8757), .ZN(n8544) );
  NAND3_X1 U8751 ( .A1(a_5_), .A2(n8758), .A3(b_26_), .ZN(n8757) );
  OR2_X1 U8752 ( .A1(n8730), .A2(n8728), .ZN(n8758) );
  NAND2_X1 U8753 ( .A1(n8728), .A2(n8730), .ZN(n8756) );
  NAND2_X1 U8754 ( .A1(n8759), .A2(n8760), .ZN(n8730) );
  NAND3_X1 U8755 ( .A1(a_6_), .A2(n8761), .A3(b_26_), .ZN(n8760) );
  NAND2_X1 U8756 ( .A1(n8727), .A2(n8725), .ZN(n8761) );
  OR2_X1 U8757 ( .A1(n8725), .A2(n8727), .ZN(n8759) );
  AND2_X1 U8758 ( .A1(n8722), .A2(n8762), .ZN(n8727) );
  NAND2_X1 U8759 ( .A1(n8721), .A2(n8723), .ZN(n8762) );
  NAND2_X1 U8760 ( .A1(n8763), .A2(n8764), .ZN(n8723) );
  NAND2_X1 U8761 ( .A1(b_26_), .A2(a_7_), .ZN(n8764) );
  INV_X1 U8762 ( .A(n8765), .ZN(n8763) );
  XOR2_X1 U8763 ( .A(n8766), .B(n8767), .Z(n8721) );
  XOR2_X1 U8764 ( .A(n8768), .B(n8769), .Z(n8766) );
  NOR2_X1 U8765 ( .A1(n8037), .A2(n8639), .ZN(n8769) );
  NAND2_X1 U8766 ( .A1(a_7_), .A2(n8765), .ZN(n8722) );
  NAND2_X1 U8767 ( .A1(n8770), .A2(n8771), .ZN(n8765) );
  NAND3_X1 U8768 ( .A1(a_8_), .A2(n8772), .A3(b_26_), .ZN(n8771) );
  OR2_X1 U8769 ( .A1(n8718), .A2(n8716), .ZN(n8772) );
  NAND2_X1 U8770 ( .A1(n8716), .A2(n8718), .ZN(n8770) );
  NAND2_X1 U8771 ( .A1(n8773), .A2(n8774), .ZN(n8718) );
  NAND2_X1 U8772 ( .A1(n8715), .A2(n8775), .ZN(n8774) );
  NAND2_X1 U8773 ( .A1(n8714), .A2(n8713), .ZN(n8775) );
  NOR2_X1 U8774 ( .A1(n8403), .A2(n7870), .ZN(n8715) );
  OR2_X1 U8775 ( .A1(n8713), .A2(n8714), .ZN(n8773) );
  AND2_X1 U8776 ( .A1(n8776), .A2(n8777), .ZN(n8714) );
  NAND3_X1 U8777 ( .A1(a_10_), .A2(n8778), .A3(b_26_), .ZN(n8777) );
  NAND2_X1 U8778 ( .A1(n8710), .A2(n8709), .ZN(n8778) );
  OR2_X1 U8779 ( .A1(n8709), .A2(n8710), .ZN(n8776) );
  AND2_X1 U8780 ( .A1(n8779), .A2(n8780), .ZN(n8710) );
  NAND2_X1 U8781 ( .A1(n8707), .A2(n8781), .ZN(n8780) );
  OR2_X1 U8782 ( .A1(n8706), .A2(n8704), .ZN(n8781) );
  NOR2_X1 U8783 ( .A1(n8403), .A2(n7877), .ZN(n8707) );
  NAND2_X1 U8784 ( .A1(n8704), .A2(n8706), .ZN(n8779) );
  NAND2_X1 U8785 ( .A1(n8782), .A2(n8783), .ZN(n8706) );
  NAND3_X1 U8786 ( .A1(a_12_), .A2(n8784), .A3(b_26_), .ZN(n8783) );
  NAND2_X1 U8787 ( .A1(n8702), .A2(n8701), .ZN(n8784) );
  OR2_X1 U8788 ( .A1(n8701), .A2(n8702), .ZN(n8782) );
  AND2_X1 U8789 ( .A1(n8785), .A2(n8786), .ZN(n8702) );
  NAND2_X1 U8790 ( .A1(n8699), .A2(n8787), .ZN(n8786) );
  OR2_X1 U8791 ( .A1(n8698), .A2(n8697), .ZN(n8787) );
  NOR2_X1 U8792 ( .A1(n8403), .A2(n7355), .ZN(n8699) );
  NAND2_X1 U8793 ( .A1(n8697), .A2(n8698), .ZN(n8785) );
  NAND2_X1 U8794 ( .A1(n8788), .A2(n8789), .ZN(n8698) );
  NAND3_X1 U8795 ( .A1(a_14_), .A2(n8790), .A3(b_26_), .ZN(n8789) );
  OR2_X1 U8796 ( .A1(n8694), .A2(n8693), .ZN(n8790) );
  NAND2_X1 U8797 ( .A1(n8693), .A2(n8694), .ZN(n8788) );
  NAND2_X1 U8798 ( .A1(n8791), .A2(n8792), .ZN(n8694) );
  NAND2_X1 U8799 ( .A1(n8691), .A2(n8793), .ZN(n8792) );
  OR2_X1 U8800 ( .A1(n8690), .A2(n8688), .ZN(n8793) );
  NOR2_X1 U8801 ( .A1(n8403), .A2(n7346), .ZN(n8691) );
  NAND2_X1 U8802 ( .A1(n8688), .A2(n8690), .ZN(n8791) );
  NAND2_X1 U8803 ( .A1(n8794), .A2(n8795), .ZN(n8690) );
  NAND3_X1 U8804 ( .A1(a_16_), .A2(n8796), .A3(b_26_), .ZN(n8795) );
  OR2_X1 U8805 ( .A1(n8686), .A2(n8684), .ZN(n8796) );
  NAND2_X1 U8806 ( .A1(n8684), .A2(n8686), .ZN(n8794) );
  NAND2_X1 U8807 ( .A1(n8797), .A2(n8798), .ZN(n8686) );
  NAND2_X1 U8808 ( .A1(n8683), .A2(n8799), .ZN(n8798) );
  OR2_X1 U8809 ( .A1(n8682), .A2(n8681), .ZN(n8799) );
  NOR2_X1 U8810 ( .A1(n8403), .A2(n7337), .ZN(n8683) );
  NAND2_X1 U8811 ( .A1(n8681), .A2(n8682), .ZN(n8797) );
  NAND2_X1 U8812 ( .A1(n8800), .A2(n8801), .ZN(n8682) );
  NAND3_X1 U8813 ( .A1(a_18_), .A2(n8802), .A3(b_26_), .ZN(n8801) );
  NAND2_X1 U8814 ( .A1(n8678), .A2(n8677), .ZN(n8802) );
  OR2_X1 U8815 ( .A1(n8677), .A2(n8678), .ZN(n8800) );
  AND2_X1 U8816 ( .A1(n8803), .A2(n8804), .ZN(n8678) );
  NAND2_X1 U8817 ( .A1(n8675), .A2(n8805), .ZN(n8804) );
  OR2_X1 U8818 ( .A1(n8674), .A2(n8672), .ZN(n8805) );
  NOR2_X1 U8819 ( .A1(n8403), .A2(n7902), .ZN(n8675) );
  NAND2_X1 U8820 ( .A1(n8672), .A2(n8674), .ZN(n8803) );
  NAND2_X1 U8821 ( .A1(n8806), .A2(n8807), .ZN(n8674) );
  NAND3_X1 U8822 ( .A1(a_20_), .A2(n8808), .A3(b_26_), .ZN(n8807) );
  NAND2_X1 U8823 ( .A1(n8670), .A2(n8669), .ZN(n8808) );
  OR2_X1 U8824 ( .A1(n8669), .A2(n8670), .ZN(n8806) );
  AND2_X1 U8825 ( .A1(n8809), .A2(n8810), .ZN(n8670) );
  NAND2_X1 U8826 ( .A1(n8667), .A2(n8811), .ZN(n8810) );
  OR2_X1 U8827 ( .A1(n8666), .A2(n8665), .ZN(n8811) );
  NOR2_X1 U8828 ( .A1(n8403), .A2(n7909), .ZN(n8667) );
  NAND2_X1 U8829 ( .A1(n8665), .A2(n8666), .ZN(n8809) );
  NAND2_X1 U8830 ( .A1(n8812), .A2(n8813), .ZN(n8666) );
  NAND3_X1 U8831 ( .A1(a_22_), .A2(n8814), .A3(b_26_), .ZN(n8813) );
  OR2_X1 U8832 ( .A1(n8662), .A2(n8660), .ZN(n8814) );
  NAND2_X1 U8833 ( .A1(n8660), .A2(n8662), .ZN(n8812) );
  NAND2_X1 U8834 ( .A1(n8815), .A2(n8816), .ZN(n8662) );
  NAND2_X1 U8835 ( .A1(n8659), .A2(n8817), .ZN(n8816) );
  OR2_X1 U8836 ( .A1(n8658), .A2(n8656), .ZN(n8817) );
  NOR2_X1 U8837 ( .A1(n8403), .A2(n7916), .ZN(n8659) );
  NAND2_X1 U8838 ( .A1(n8656), .A2(n8658), .ZN(n8815) );
  NAND2_X1 U8839 ( .A1(n8818), .A2(n8819), .ZN(n8658) );
  NAND3_X1 U8840 ( .A1(a_24_), .A2(n8820), .A3(b_26_), .ZN(n8819) );
  NAND2_X1 U8841 ( .A1(n8654), .A2(n8653), .ZN(n8820) );
  OR2_X1 U8842 ( .A1(n8653), .A2(n8654), .ZN(n8818) );
  AND2_X1 U8843 ( .A1(n8821), .A2(n8822), .ZN(n8654) );
  NAND2_X1 U8844 ( .A1(n8651), .A2(n8823), .ZN(n8822) );
  OR2_X1 U8845 ( .A1(n8650), .A2(n8648), .ZN(n8823) );
  NOR2_X1 U8846 ( .A1(n8403), .A2(n7923), .ZN(n8651) );
  NAND2_X1 U8847 ( .A1(n8648), .A2(n8650), .ZN(n8821) );
  NAND2_X1 U8848 ( .A1(n8824), .A2(n8825), .ZN(n8650) );
  NAND2_X1 U8849 ( .A1(n8647), .A2(n8826), .ZN(n8825) );
  OR2_X1 U8850 ( .A1(n8646), .A2(n8645), .ZN(n8826) );
  INV_X1 U8851 ( .A(n8827), .ZN(n8647) );
  NAND2_X1 U8852 ( .A1(n8645), .A2(n8646), .ZN(n8824) );
  NAND2_X1 U8853 ( .A1(n8618), .A2(n8828), .ZN(n8646) );
  NAND2_X1 U8854 ( .A1(n8617), .A2(n8619), .ZN(n8828) );
  NAND2_X1 U8855 ( .A1(n8829), .A2(n8830), .ZN(n8619) );
  NAND2_X1 U8856 ( .A1(b_26_), .A2(a_27_), .ZN(n8830) );
  INV_X1 U8857 ( .A(n8831), .ZN(n8829) );
  XNOR2_X1 U8858 ( .A(n8832), .B(n8833), .ZN(n8617) );
  XOR2_X1 U8859 ( .A(n8834), .B(n8835), .Z(n8832) );
  NAND2_X1 U8860 ( .A1(b_25_), .A2(a_28_), .ZN(n8834) );
  NAND2_X1 U8861 ( .A1(a_27_), .A2(n8831), .ZN(n8618) );
  NAND2_X1 U8862 ( .A1(n8836), .A2(n8837), .ZN(n8831) );
  NAND3_X1 U8863 ( .A1(a_28_), .A2(n8838), .A3(b_26_), .ZN(n8837) );
  NAND2_X1 U8864 ( .A1(n8626), .A2(n8624), .ZN(n8838) );
  OR2_X1 U8865 ( .A1(n8624), .A2(n8626), .ZN(n8836) );
  AND2_X1 U8866 ( .A1(n8839), .A2(n8840), .ZN(n8626) );
  NAND2_X1 U8867 ( .A1(n8641), .A2(n8841), .ZN(n8840) );
  OR2_X1 U8868 ( .A1(n8642), .A2(n8643), .ZN(n8841) );
  NOR2_X1 U8869 ( .A1(n8403), .A2(n7946), .ZN(n8641) );
  NAND2_X1 U8870 ( .A1(n8643), .A2(n8642), .ZN(n8839) );
  NAND2_X1 U8871 ( .A1(n8842), .A2(n8843), .ZN(n8642) );
  NAND2_X1 U8872 ( .A1(b_24_), .A2(n8844), .ZN(n8843) );
  NAND2_X1 U8873 ( .A1(n7268), .A2(n8845), .ZN(n8844) );
  NAND2_X1 U8874 ( .A1(a_31_), .A2(n8639), .ZN(n8845) );
  NAND2_X1 U8875 ( .A1(b_25_), .A2(n8846), .ZN(n8842) );
  NAND2_X1 U8876 ( .A1(n7272), .A2(n8847), .ZN(n8846) );
  NAND2_X1 U8877 ( .A1(a_30_), .A2(n8848), .ZN(n8847) );
  AND3_X1 U8878 ( .A1(b_25_), .A2(n7954), .A3(b_26_), .ZN(n8643) );
  XNOR2_X1 U8879 ( .A(n8849), .B(n8850), .ZN(n8624) );
  XOR2_X1 U8880 ( .A(n8851), .B(n8852), .Z(n8849) );
  XNOR2_X1 U8881 ( .A(n8853), .B(n8854), .ZN(n8645) );
  NAND2_X1 U8882 ( .A1(n8855), .A2(n8856), .ZN(n8853) );
  XNOR2_X1 U8883 ( .A(n8857), .B(n8858), .ZN(n8648) );
  NAND2_X1 U8884 ( .A1(n8859), .A2(n8860), .ZN(n8857) );
  XNOR2_X1 U8885 ( .A(n8861), .B(n8862), .ZN(n8653) );
  XOR2_X1 U8886 ( .A(n8863), .B(n8864), .Z(n8861) );
  XNOR2_X1 U8887 ( .A(n8865), .B(n8866), .ZN(n8656) );
  XNOR2_X1 U8888 ( .A(n8867), .B(n8868), .ZN(n8865) );
  NOR2_X1 U8889 ( .A1(n7691), .A2(n8639), .ZN(n8868) );
  XNOR2_X1 U8890 ( .A(n8869), .B(n8870), .ZN(n8660) );
  XNOR2_X1 U8891 ( .A(n8871), .B(n8872), .ZN(n8870) );
  XNOR2_X1 U8892 ( .A(n8873), .B(n8874), .ZN(n8665) );
  XOR2_X1 U8893 ( .A(n8875), .B(n8876), .Z(n8874) );
  NAND2_X1 U8894 ( .A1(b_25_), .A2(a_22_), .ZN(n8876) );
  XNOR2_X1 U8895 ( .A(n8877), .B(n8878), .ZN(n8669) );
  XOR2_X1 U8896 ( .A(n8879), .B(n8880), .Z(n8877) );
  XNOR2_X1 U8897 ( .A(n8881), .B(n8882), .ZN(n8672) );
  XNOR2_X1 U8898 ( .A(n8883), .B(n8884), .ZN(n8881) );
  NOR2_X1 U8899 ( .A1(n7987), .A2(n8639), .ZN(n8884) );
  XOR2_X1 U8900 ( .A(n8885), .B(n8886), .Z(n8677) );
  XNOR2_X1 U8901 ( .A(n8887), .B(n8888), .ZN(n8886) );
  XNOR2_X1 U8902 ( .A(n8889), .B(n8890), .ZN(n8681) );
  XNOR2_X1 U8903 ( .A(n8891), .B(n8892), .ZN(n8889) );
  NOR2_X1 U8904 ( .A1(n7764), .A2(n8639), .ZN(n8892) );
  XOR2_X1 U8905 ( .A(n8893), .B(n8894), .Z(n8684) );
  XOR2_X1 U8906 ( .A(n8895), .B(n8896), .Z(n8893) );
  XNOR2_X1 U8907 ( .A(n8897), .B(n8898), .ZN(n8688) );
  XOR2_X1 U8908 ( .A(n8899), .B(n8900), .Z(n8898) );
  NAND2_X1 U8909 ( .A1(b_25_), .A2(a_16_), .ZN(n8900) );
  XNOR2_X1 U8910 ( .A(n8901), .B(n8902), .ZN(n8693) );
  XNOR2_X1 U8911 ( .A(n8903), .B(n8904), .ZN(n8902) );
  XNOR2_X1 U8912 ( .A(n8905), .B(n8906), .ZN(n8697) );
  XOR2_X1 U8913 ( .A(n8907), .B(n8908), .Z(n8905) );
  NAND2_X1 U8914 ( .A1(b_25_), .A2(a_14_), .ZN(n8907) );
  XNOR2_X1 U8915 ( .A(n8909), .B(n8910), .ZN(n8701) );
  XOR2_X1 U8916 ( .A(n8911), .B(n8912), .Z(n8909) );
  XOR2_X1 U8917 ( .A(n8913), .B(n8914), .Z(n8704) );
  XOR2_X1 U8918 ( .A(n8915), .B(n8916), .Z(n8913) );
  NOR2_X1 U8919 ( .A1(n8020), .A2(n8639), .ZN(n8916) );
  XOR2_X1 U8920 ( .A(n8917), .B(n8918), .Z(n8709) );
  XOR2_X1 U8921 ( .A(n8919), .B(n8920), .Z(n8918) );
  NAND2_X1 U8922 ( .A1(b_25_), .A2(a_11_), .ZN(n8920) );
  XNOR2_X1 U8923 ( .A(n8921), .B(n8922), .ZN(n8713) );
  XOR2_X1 U8924 ( .A(n8923), .B(n8924), .Z(n8921) );
  NOR2_X1 U8925 ( .A1(n7799), .A2(n8639), .ZN(n8924) );
  XOR2_X1 U8926 ( .A(n8925), .B(n8926), .Z(n8716) );
  XOR2_X1 U8927 ( .A(n8927), .B(n8928), .Z(n8925) );
  XNOR2_X1 U8928 ( .A(n8929), .B(n8930), .ZN(n8725) );
  XOR2_X1 U8929 ( .A(n8931), .B(n8932), .Z(n8929) );
  NOR2_X1 U8930 ( .A1(n7863), .A2(n8639), .ZN(n8932) );
  XNOR2_X1 U8931 ( .A(n8933), .B(n8934), .ZN(n8728) );
  XOR2_X1 U8932 ( .A(n8935), .B(n8936), .Z(n8934) );
  XNOR2_X1 U8933 ( .A(n8937), .B(n8938), .ZN(n8542) );
  XNOR2_X1 U8934 ( .A(n8939), .B(n8940), .ZN(n8937) );
  NOR2_X1 U8935 ( .A1(n7393), .A2(n8639), .ZN(n8940) );
  XOR2_X1 U8936 ( .A(n8941), .B(n8942), .Z(n8535) );
  XOR2_X1 U8937 ( .A(n8943), .B(n8944), .Z(n8942) );
  NAND2_X1 U8938 ( .A1(b_25_), .A2(a_4_), .ZN(n8944) );
  XNOR2_X1 U8939 ( .A(n8945), .B(n8946), .ZN(n8732) );
  XOR2_X1 U8940 ( .A(n8947), .B(n8948), .Z(n8946) );
  NAND2_X1 U8941 ( .A1(b_25_), .A2(a_3_), .ZN(n8948) );
  XNOR2_X1 U8942 ( .A(n8949), .B(n8950), .ZN(n8737) );
  XOR2_X1 U8943 ( .A(n8951), .B(n8952), .Z(n8949) );
  NOR2_X1 U8944 ( .A1(n7832), .A2(n8639), .ZN(n8952) );
  XOR2_X1 U8945 ( .A(n8953), .B(n8954), .Z(n8520) );
  XOR2_X1 U8946 ( .A(n8955), .B(n8956), .Z(n8953) );
  NOR2_X1 U8947 ( .A1(n7411), .A2(n8639), .ZN(n8956) );
  NAND2_X1 U8948 ( .A1(n8957), .A2(n8958), .ZN(n7590) );
  INV_X1 U8949 ( .A(n8518), .ZN(n7591) );
  XOR2_X1 U8950 ( .A(n8959), .B(n8960), .Z(n8518) );
  XNOR2_X1 U8951 ( .A(n8961), .B(n8962), .ZN(n8960) );
  NAND2_X1 U8952 ( .A1(n8963), .A2(n8740), .ZN(n7447) );
  NOR2_X1 U8953 ( .A1(n8958), .A2(n8957), .ZN(n8740) );
  AND2_X1 U8954 ( .A1(n8964), .A2(n8965), .ZN(n8957) );
  NAND2_X1 U8955 ( .A1(n8962), .A2(n8966), .ZN(n8965) );
  OR2_X1 U8956 ( .A1(n8961), .A2(n8959), .ZN(n8966) );
  NOR2_X1 U8957 ( .A1(n8639), .A2(n7613), .ZN(n8962) );
  NAND2_X1 U8958 ( .A1(n8959), .A2(n8961), .ZN(n8964) );
  NAND2_X1 U8959 ( .A1(n8967), .A2(n8968), .ZN(n8961) );
  NAND3_X1 U8960 ( .A1(a_1_), .A2(n8969), .A3(b_25_), .ZN(n8968) );
  OR2_X1 U8961 ( .A1(n8955), .A2(n8954), .ZN(n8969) );
  NAND2_X1 U8962 ( .A1(n8954), .A2(n8955), .ZN(n8967) );
  NAND2_X1 U8963 ( .A1(n8970), .A2(n8971), .ZN(n8955) );
  NAND3_X1 U8964 ( .A1(a_2_), .A2(n8972), .A3(b_25_), .ZN(n8971) );
  OR2_X1 U8965 ( .A1(n8951), .A2(n8950), .ZN(n8972) );
  NAND2_X1 U8966 ( .A1(n8950), .A2(n8951), .ZN(n8970) );
  NAND2_X1 U8967 ( .A1(n8973), .A2(n8974), .ZN(n8951) );
  NAND3_X1 U8968 ( .A1(a_3_), .A2(n8975), .A3(b_25_), .ZN(n8974) );
  OR2_X1 U8969 ( .A1(n8947), .A2(n8945), .ZN(n8975) );
  NAND2_X1 U8970 ( .A1(n8945), .A2(n8947), .ZN(n8973) );
  NAND2_X1 U8971 ( .A1(n8976), .A2(n8977), .ZN(n8947) );
  NAND3_X1 U8972 ( .A1(a_4_), .A2(n8978), .A3(b_25_), .ZN(n8977) );
  OR2_X1 U8973 ( .A1(n8943), .A2(n8941), .ZN(n8978) );
  NAND2_X1 U8974 ( .A1(n8941), .A2(n8943), .ZN(n8976) );
  NAND2_X1 U8975 ( .A1(n8979), .A2(n8980), .ZN(n8943) );
  NAND3_X1 U8976 ( .A1(a_5_), .A2(n8981), .A3(b_25_), .ZN(n8980) );
  NAND2_X1 U8977 ( .A1(n8939), .A2(n8938), .ZN(n8981) );
  OR2_X1 U8978 ( .A1(n8938), .A2(n8939), .ZN(n8979) );
  AND2_X1 U8979 ( .A1(n8982), .A2(n8983), .ZN(n8939) );
  NAND2_X1 U8980 ( .A1(n8935), .A2(n8984), .ZN(n8983) );
  NAND2_X1 U8981 ( .A1(n8985), .A2(n8936), .ZN(n8984) );
  INV_X1 U8982 ( .A(n8933), .ZN(n8985) );
  NAND2_X1 U8983 ( .A1(n8986), .A2(n8987), .ZN(n8935) );
  NAND3_X1 U8984 ( .A1(a_7_), .A2(n8988), .A3(b_25_), .ZN(n8987) );
  OR2_X1 U8985 ( .A1(n8931), .A2(n8930), .ZN(n8988) );
  NAND2_X1 U8986 ( .A1(n8930), .A2(n8931), .ZN(n8986) );
  NAND2_X1 U8987 ( .A1(n8989), .A2(n8990), .ZN(n8931) );
  NAND3_X1 U8988 ( .A1(a_8_), .A2(n8991), .A3(b_25_), .ZN(n8990) );
  OR2_X1 U8989 ( .A1(n8768), .A2(n8767), .ZN(n8991) );
  NAND2_X1 U8990 ( .A1(n8767), .A2(n8768), .ZN(n8989) );
  NAND2_X1 U8991 ( .A1(n8992), .A2(n8993), .ZN(n8768) );
  NAND2_X1 U8992 ( .A1(n8928), .A2(n8994), .ZN(n8993) );
  OR2_X1 U8993 ( .A1(n8927), .A2(n8926), .ZN(n8994) );
  NOR2_X1 U8994 ( .A1(n8639), .A2(n7870), .ZN(n8928) );
  NAND2_X1 U8995 ( .A1(n8926), .A2(n8927), .ZN(n8992) );
  NAND2_X1 U8996 ( .A1(n8995), .A2(n8996), .ZN(n8927) );
  NAND3_X1 U8997 ( .A1(a_10_), .A2(n8997), .A3(b_25_), .ZN(n8996) );
  OR2_X1 U8998 ( .A1(n8923), .A2(n8922), .ZN(n8997) );
  NAND2_X1 U8999 ( .A1(n8922), .A2(n8923), .ZN(n8995) );
  NAND2_X1 U9000 ( .A1(n8998), .A2(n8999), .ZN(n8923) );
  NAND3_X1 U9001 ( .A1(a_11_), .A2(n9000), .A3(b_25_), .ZN(n8999) );
  OR2_X1 U9002 ( .A1(n8919), .A2(n8917), .ZN(n9000) );
  NAND2_X1 U9003 ( .A1(n8917), .A2(n8919), .ZN(n8998) );
  NAND2_X1 U9004 ( .A1(n9001), .A2(n9002), .ZN(n8919) );
  NAND3_X1 U9005 ( .A1(a_12_), .A2(n9003), .A3(b_25_), .ZN(n9002) );
  OR2_X1 U9006 ( .A1(n8915), .A2(n8914), .ZN(n9003) );
  NAND2_X1 U9007 ( .A1(n8914), .A2(n8915), .ZN(n9001) );
  NAND2_X1 U9008 ( .A1(n9004), .A2(n9005), .ZN(n8915) );
  NAND2_X1 U9009 ( .A1(n8912), .A2(n9006), .ZN(n9005) );
  OR2_X1 U9010 ( .A1(n8911), .A2(n8910), .ZN(n9006) );
  NOR2_X1 U9011 ( .A1(n8639), .A2(n7355), .ZN(n8912) );
  NAND2_X1 U9012 ( .A1(n8910), .A2(n8911), .ZN(n9004) );
  NAND2_X1 U9013 ( .A1(n9007), .A2(n9008), .ZN(n8911) );
  NAND3_X1 U9014 ( .A1(a_14_), .A2(n9009), .A3(b_25_), .ZN(n9008) );
  NAND2_X1 U9015 ( .A1(n8908), .A2(n8906), .ZN(n9009) );
  OR2_X1 U9016 ( .A1(n8906), .A2(n8908), .ZN(n9007) );
  AND2_X1 U9017 ( .A1(n9010), .A2(n9011), .ZN(n8908) );
  NAND2_X1 U9018 ( .A1(n8904), .A2(n9012), .ZN(n9011) );
  OR2_X1 U9019 ( .A1(n8903), .A2(n8901), .ZN(n9012) );
  NOR2_X1 U9020 ( .A1(n8639), .A2(n7346), .ZN(n8904) );
  NAND2_X1 U9021 ( .A1(n8901), .A2(n8903), .ZN(n9010) );
  NAND2_X1 U9022 ( .A1(n9013), .A2(n9014), .ZN(n8903) );
  NAND3_X1 U9023 ( .A1(a_16_), .A2(n9015), .A3(b_25_), .ZN(n9014) );
  OR2_X1 U9024 ( .A1(n8899), .A2(n8897), .ZN(n9015) );
  NAND2_X1 U9025 ( .A1(n8897), .A2(n8899), .ZN(n9013) );
  NAND2_X1 U9026 ( .A1(n9016), .A2(n9017), .ZN(n8899) );
  NAND2_X1 U9027 ( .A1(n8896), .A2(n9018), .ZN(n9017) );
  OR2_X1 U9028 ( .A1(n8895), .A2(n8894), .ZN(n9018) );
  NOR2_X1 U9029 ( .A1(n8639), .A2(n7337), .ZN(n8896) );
  NAND2_X1 U9030 ( .A1(n8894), .A2(n8895), .ZN(n9016) );
  NAND2_X1 U9031 ( .A1(n9019), .A2(n9020), .ZN(n8895) );
  NAND3_X1 U9032 ( .A1(a_18_), .A2(n9021), .A3(b_25_), .ZN(n9020) );
  NAND2_X1 U9033 ( .A1(n8891), .A2(n8890), .ZN(n9021) );
  OR2_X1 U9034 ( .A1(n8890), .A2(n8891), .ZN(n9019) );
  AND2_X1 U9035 ( .A1(n9022), .A2(n9023), .ZN(n8891) );
  NAND2_X1 U9036 ( .A1(n8888), .A2(n9024), .ZN(n9023) );
  OR2_X1 U9037 ( .A1(n8887), .A2(n8885), .ZN(n9024) );
  NOR2_X1 U9038 ( .A1(n8639), .A2(n7902), .ZN(n8888) );
  NAND2_X1 U9039 ( .A1(n8885), .A2(n8887), .ZN(n9022) );
  NAND2_X1 U9040 ( .A1(n9025), .A2(n9026), .ZN(n8887) );
  NAND3_X1 U9041 ( .A1(a_20_), .A2(n9027), .A3(b_25_), .ZN(n9026) );
  NAND2_X1 U9042 ( .A1(n8883), .A2(n8882), .ZN(n9027) );
  OR2_X1 U9043 ( .A1(n8882), .A2(n8883), .ZN(n9025) );
  AND2_X1 U9044 ( .A1(n9028), .A2(n9029), .ZN(n8883) );
  NAND2_X1 U9045 ( .A1(n8880), .A2(n9030), .ZN(n9029) );
  OR2_X1 U9046 ( .A1(n8879), .A2(n8878), .ZN(n9030) );
  NOR2_X1 U9047 ( .A1(n8639), .A2(n7909), .ZN(n8880) );
  NAND2_X1 U9048 ( .A1(n8878), .A2(n8879), .ZN(n9028) );
  NAND2_X1 U9049 ( .A1(n9031), .A2(n9032), .ZN(n8879) );
  NAND3_X1 U9050 ( .A1(a_22_), .A2(n9033), .A3(b_25_), .ZN(n9032) );
  OR2_X1 U9051 ( .A1(n8875), .A2(n8873), .ZN(n9033) );
  NAND2_X1 U9052 ( .A1(n8873), .A2(n8875), .ZN(n9031) );
  NAND2_X1 U9053 ( .A1(n9034), .A2(n9035), .ZN(n8875) );
  NAND2_X1 U9054 ( .A1(n8872), .A2(n9036), .ZN(n9035) );
  OR2_X1 U9055 ( .A1(n8871), .A2(n8869), .ZN(n9036) );
  NOR2_X1 U9056 ( .A1(n8639), .A2(n7916), .ZN(n8872) );
  NAND2_X1 U9057 ( .A1(n8869), .A2(n8871), .ZN(n9034) );
  NAND2_X1 U9058 ( .A1(n9037), .A2(n9038), .ZN(n8871) );
  NAND3_X1 U9059 ( .A1(a_24_), .A2(n9039), .A3(b_25_), .ZN(n9038) );
  NAND2_X1 U9060 ( .A1(n8867), .A2(n8866), .ZN(n9039) );
  OR2_X1 U9061 ( .A1(n8866), .A2(n8867), .ZN(n9037) );
  AND2_X1 U9062 ( .A1(n9040), .A2(n9041), .ZN(n8867) );
  NAND2_X1 U9063 ( .A1(n8864), .A2(n9042), .ZN(n9041) );
  OR2_X1 U9064 ( .A1(n8863), .A2(n8862), .ZN(n9042) );
  NAND2_X1 U9065 ( .A1(n8862), .A2(n8863), .ZN(n9040) );
  NAND2_X1 U9066 ( .A1(n8859), .A2(n9043), .ZN(n8863) );
  NAND2_X1 U9067 ( .A1(n8858), .A2(n8860), .ZN(n9043) );
  NAND2_X1 U9068 ( .A1(n9044), .A2(n9045), .ZN(n8860) );
  NAND2_X1 U9069 ( .A1(b_25_), .A2(a_26_), .ZN(n9045) );
  INV_X1 U9070 ( .A(n9046), .ZN(n9044) );
  XNOR2_X1 U9071 ( .A(n9047), .B(n9048), .ZN(n8858) );
  NAND2_X1 U9072 ( .A1(n9049), .A2(n9050), .ZN(n9047) );
  NAND2_X1 U9073 ( .A1(a_26_), .A2(n9046), .ZN(n8859) );
  NAND2_X1 U9074 ( .A1(n8855), .A2(n9051), .ZN(n9046) );
  NAND2_X1 U9075 ( .A1(n8854), .A2(n8856), .ZN(n9051) );
  NAND2_X1 U9076 ( .A1(n9052), .A2(n9053), .ZN(n8856) );
  NAND2_X1 U9077 ( .A1(b_25_), .A2(a_27_), .ZN(n9053) );
  INV_X1 U9078 ( .A(n9054), .ZN(n9052) );
  XNOR2_X1 U9079 ( .A(n9055), .B(n9056), .ZN(n8854) );
  XOR2_X1 U9080 ( .A(n9057), .B(n9058), .Z(n9055) );
  NAND2_X1 U9081 ( .A1(b_24_), .A2(a_28_), .ZN(n9057) );
  NAND2_X1 U9082 ( .A1(a_27_), .A2(n9054), .ZN(n8855) );
  NAND2_X1 U9083 ( .A1(n9059), .A2(n9060), .ZN(n9054) );
  NAND3_X1 U9084 ( .A1(a_28_), .A2(n9061), .A3(b_25_), .ZN(n9060) );
  NAND2_X1 U9085 ( .A1(n8835), .A2(n8833), .ZN(n9061) );
  OR2_X1 U9086 ( .A1(n8833), .A2(n8835), .ZN(n9059) );
  AND2_X1 U9087 ( .A1(n9062), .A2(n9063), .ZN(n8835) );
  NAND2_X1 U9088 ( .A1(n8850), .A2(n9064), .ZN(n9063) );
  OR2_X1 U9089 ( .A1(n8851), .A2(n8852), .ZN(n9064) );
  NOR2_X1 U9090 ( .A1(n8639), .A2(n7946), .ZN(n8850) );
  NAND2_X1 U9091 ( .A1(n8852), .A2(n8851), .ZN(n9062) );
  NAND2_X1 U9092 ( .A1(n9065), .A2(n9066), .ZN(n8851) );
  NAND2_X1 U9093 ( .A1(b_23_), .A2(n9067), .ZN(n9066) );
  NAND2_X1 U9094 ( .A1(n7268), .A2(n9068), .ZN(n9067) );
  NAND2_X1 U9095 ( .A1(a_31_), .A2(n8848), .ZN(n9068) );
  NAND2_X1 U9096 ( .A1(b_24_), .A2(n9069), .ZN(n9065) );
  NAND2_X1 U9097 ( .A1(n7272), .A2(n9070), .ZN(n9069) );
  NAND2_X1 U9098 ( .A1(a_30_), .A2(n9071), .ZN(n9070) );
  AND3_X1 U9099 ( .A1(b_24_), .A2(n7954), .A3(b_25_), .ZN(n8852) );
  XNOR2_X1 U9100 ( .A(n9072), .B(n9073), .ZN(n8833) );
  XOR2_X1 U9101 ( .A(n9074), .B(n9075), .Z(n9072) );
  XNOR2_X1 U9102 ( .A(n9076), .B(n9077), .ZN(n8862) );
  NAND2_X1 U9103 ( .A1(n9078), .A2(n9079), .ZN(n9076) );
  XNOR2_X1 U9104 ( .A(n9080), .B(n9081), .ZN(n8866) );
  XOR2_X1 U9105 ( .A(n9082), .B(n9083), .Z(n9080) );
  XNOR2_X1 U9106 ( .A(n9084), .B(n9085), .ZN(n8869) );
  XNOR2_X1 U9107 ( .A(n9086), .B(n9087), .ZN(n9084) );
  XNOR2_X1 U9108 ( .A(n9088), .B(n9089), .ZN(n8873) );
  XNOR2_X1 U9109 ( .A(n9090), .B(n9091), .ZN(n9089) );
  XNOR2_X1 U9110 ( .A(n9092), .B(n9093), .ZN(n8878) );
  XOR2_X1 U9111 ( .A(n9094), .B(n9095), .Z(n9093) );
  NAND2_X1 U9112 ( .A1(b_24_), .A2(a_22_), .ZN(n9095) );
  XNOR2_X1 U9113 ( .A(n9096), .B(n9097), .ZN(n8882) );
  XOR2_X1 U9114 ( .A(n9098), .B(n9099), .Z(n9096) );
  XNOR2_X1 U9115 ( .A(n9100), .B(n9101), .ZN(n8885) );
  XNOR2_X1 U9116 ( .A(n9102), .B(n9103), .ZN(n9100) );
  NOR2_X1 U9117 ( .A1(n7987), .A2(n8848), .ZN(n9103) );
  XOR2_X1 U9118 ( .A(n9104), .B(n9105), .Z(n8890) );
  XNOR2_X1 U9119 ( .A(n9106), .B(n9107), .ZN(n9105) );
  XNOR2_X1 U9120 ( .A(n9108), .B(n9109), .ZN(n8894) );
  XNOR2_X1 U9121 ( .A(n9110), .B(n9111), .ZN(n9108) );
  NOR2_X1 U9122 ( .A1(n7764), .A2(n8848), .ZN(n9111) );
  XOR2_X1 U9123 ( .A(n9112), .B(n9113), .Z(n8897) );
  XOR2_X1 U9124 ( .A(n9114), .B(n9115), .Z(n9112) );
  XNOR2_X1 U9125 ( .A(n9116), .B(n9117), .ZN(n8901) );
  XOR2_X1 U9126 ( .A(n9118), .B(n9119), .Z(n9117) );
  NAND2_X1 U9127 ( .A1(b_24_), .A2(a_16_), .ZN(n9119) );
  XOR2_X1 U9128 ( .A(n9120), .B(n9121), .Z(n8906) );
  XNOR2_X1 U9129 ( .A(n9122), .B(n9123), .ZN(n9121) );
  XNOR2_X1 U9130 ( .A(n9124), .B(n9125), .ZN(n8910) );
  XOR2_X1 U9131 ( .A(n9126), .B(n9127), .Z(n9124) );
  NAND2_X1 U9132 ( .A1(b_24_), .A2(a_14_), .ZN(n9126) );
  XNOR2_X1 U9133 ( .A(n9128), .B(n9129), .ZN(n8914) );
  XNOR2_X1 U9134 ( .A(n9130), .B(n9131), .ZN(n9128) );
  XNOR2_X1 U9135 ( .A(n9132), .B(n9133), .ZN(n8917) );
  XOR2_X1 U9136 ( .A(n9134), .B(n9135), .Z(n9133) );
  NAND2_X1 U9137 ( .A1(b_24_), .A2(a_12_), .ZN(n9135) );
  XNOR2_X1 U9138 ( .A(n9136), .B(n9137), .ZN(n8922) );
  NAND2_X1 U9139 ( .A1(n9138), .A2(n9139), .ZN(n9136) );
  XNOR2_X1 U9140 ( .A(n9140), .B(n9141), .ZN(n8926) );
  XNOR2_X1 U9141 ( .A(n9142), .B(n9143), .ZN(n9141) );
  NOR2_X1 U9142 ( .A1(n7799), .A2(n8848), .ZN(n9143) );
  XNOR2_X1 U9143 ( .A(n9144), .B(n9145), .ZN(n8767) );
  XNOR2_X1 U9144 ( .A(n9146), .B(n9147), .ZN(n9145) );
  XNOR2_X1 U9145 ( .A(n9148), .B(n9149), .ZN(n8930) );
  XOR2_X1 U9146 ( .A(n9150), .B(n9151), .Z(n9148) );
  NAND2_X1 U9147 ( .A1(b_24_), .A2(a_8_), .ZN(n9150) );
  NAND2_X1 U9148 ( .A1(n9152), .A2(n8933), .ZN(n8982) );
  XNOR2_X1 U9149 ( .A(n9153), .B(n9154), .ZN(n8933) );
  NAND2_X1 U9150 ( .A1(n9155), .A2(n9156), .ZN(n9153) );
  INV_X1 U9151 ( .A(n8936), .ZN(n9152) );
  NAND2_X1 U9152 ( .A1(b_25_), .A2(a_6_), .ZN(n8936) );
  XNOR2_X1 U9153 ( .A(n9157), .B(n9158), .ZN(n8938) );
  XOR2_X1 U9154 ( .A(n9159), .B(n9160), .Z(n9157) );
  XNOR2_X1 U9155 ( .A(n9161), .B(n9162), .ZN(n8941) );
  XNOR2_X1 U9156 ( .A(n9163), .B(n9164), .ZN(n9161) );
  XNOR2_X1 U9157 ( .A(n9165), .B(n9166), .ZN(n8945) );
  XNOR2_X1 U9158 ( .A(n9167), .B(n9168), .ZN(n9165) );
  NOR2_X1 U9159 ( .A1(n7398), .A2(n8848), .ZN(n9168) );
  XNOR2_X1 U9160 ( .A(n9169), .B(n9170), .ZN(n8950) );
  NAND2_X1 U9161 ( .A1(n9171), .A2(n9172), .ZN(n9169) );
  XNOR2_X1 U9162 ( .A(n9173), .B(n9174), .ZN(n8954) );
  NAND2_X1 U9163 ( .A1(n9175), .A2(n9176), .ZN(n9173) );
  XOR2_X1 U9164 ( .A(n9177), .B(n9178), .Z(n8959) );
  XOR2_X1 U9165 ( .A(n9179), .B(n9180), .Z(n9178) );
  XNOR2_X1 U9166 ( .A(n9181), .B(n9182), .ZN(n8958) );
  XOR2_X1 U9167 ( .A(n9183), .B(n9184), .Z(n9181) );
  NOR2_X1 U9168 ( .A1(n7613), .A2(n8848), .ZN(n9184) );
  XOR2_X1 U9169 ( .A(n7582), .B(n7581), .Z(n8963) );
  NAND3_X1 U9170 ( .A1(n7581), .A2(n7582), .A3(n9185), .ZN(n7452) );
  XOR2_X1 U9171 ( .A(n7577), .B(n7576), .Z(n9185) );
  NAND2_X1 U9172 ( .A1(n9186), .A2(n9187), .ZN(n7582) );
  NAND3_X1 U9173 ( .A1(a_0_), .A2(n9188), .A3(b_24_), .ZN(n9187) );
  OR2_X1 U9174 ( .A1(n9183), .A2(n9182), .ZN(n9188) );
  NAND2_X1 U9175 ( .A1(n9182), .A2(n9183), .ZN(n9186) );
  NAND2_X1 U9176 ( .A1(n9189), .A2(n9190), .ZN(n9183) );
  NAND2_X1 U9177 ( .A1(n9179), .A2(n9191), .ZN(n9190) );
  NAND2_X1 U9178 ( .A1(n9177), .A2(n9180), .ZN(n9191) );
  NAND2_X1 U9179 ( .A1(n9175), .A2(n9192), .ZN(n9179) );
  NAND2_X1 U9180 ( .A1(n9174), .A2(n9176), .ZN(n9192) );
  NAND2_X1 U9181 ( .A1(n9193), .A2(n9194), .ZN(n9176) );
  NAND2_X1 U9182 ( .A1(b_24_), .A2(a_2_), .ZN(n9194) );
  INV_X1 U9183 ( .A(n9195), .ZN(n9193) );
  XNOR2_X1 U9184 ( .A(n9196), .B(n9197), .ZN(n9174) );
  XOR2_X1 U9185 ( .A(n9198), .B(n9199), .Z(n9197) );
  NAND2_X1 U9186 ( .A1(b_23_), .A2(a_3_), .ZN(n9199) );
  NAND2_X1 U9187 ( .A1(a_2_), .A2(n9195), .ZN(n9175) );
  NAND2_X1 U9188 ( .A1(n9171), .A2(n9200), .ZN(n9195) );
  NAND2_X1 U9189 ( .A1(n9170), .A2(n9172), .ZN(n9200) );
  NAND2_X1 U9190 ( .A1(n9201), .A2(n9202), .ZN(n9172) );
  NAND2_X1 U9191 ( .A1(b_24_), .A2(a_3_), .ZN(n9202) );
  INV_X1 U9192 ( .A(n9203), .ZN(n9201) );
  XNOR2_X1 U9193 ( .A(n9204), .B(n9205), .ZN(n9170) );
  XOR2_X1 U9194 ( .A(n9206), .B(n9207), .Z(n9205) );
  NAND2_X1 U9195 ( .A1(b_23_), .A2(a_4_), .ZN(n9207) );
  NAND2_X1 U9196 ( .A1(a_3_), .A2(n9203), .ZN(n9171) );
  NAND2_X1 U9197 ( .A1(n9208), .A2(n9209), .ZN(n9203) );
  NAND3_X1 U9198 ( .A1(a_4_), .A2(n9210), .A3(b_24_), .ZN(n9209) );
  NAND2_X1 U9199 ( .A1(n9167), .A2(n9166), .ZN(n9210) );
  OR2_X1 U9200 ( .A1(n9166), .A2(n9167), .ZN(n9208) );
  AND2_X1 U9201 ( .A1(n9211), .A2(n9212), .ZN(n9167) );
  NAND2_X1 U9202 ( .A1(n9164), .A2(n9213), .ZN(n9212) );
  NAND2_X1 U9203 ( .A1(n9163), .A2(n9162), .ZN(n9213) );
  NOR2_X1 U9204 ( .A1(n8848), .A2(n7393), .ZN(n9164) );
  OR2_X1 U9205 ( .A1(n9162), .A2(n9163), .ZN(n9211) );
  AND2_X1 U9206 ( .A1(n9214), .A2(n9215), .ZN(n9163) );
  NAND2_X1 U9207 ( .A1(n9160), .A2(n9216), .ZN(n9215) );
  OR2_X1 U9208 ( .A1(n9158), .A2(n9159), .ZN(n9216) );
  NAND2_X1 U9209 ( .A1(n9155), .A2(n9217), .ZN(n9160) );
  NAND2_X1 U9210 ( .A1(n9154), .A2(n9156), .ZN(n9217) );
  NAND2_X1 U9211 ( .A1(n9218), .A2(n9219), .ZN(n9156) );
  NAND2_X1 U9212 ( .A1(b_24_), .A2(a_7_), .ZN(n9219) );
  INV_X1 U9213 ( .A(n9220), .ZN(n9218) );
  XNOR2_X1 U9214 ( .A(n9221), .B(n9222), .ZN(n9154) );
  XNOR2_X1 U9215 ( .A(n9223), .B(n9224), .ZN(n9222) );
  NAND2_X1 U9216 ( .A1(a_7_), .A2(n9220), .ZN(n9155) );
  NAND2_X1 U9217 ( .A1(n9225), .A2(n9226), .ZN(n9220) );
  NAND3_X1 U9218 ( .A1(a_8_), .A2(n9227), .A3(b_24_), .ZN(n9226) );
  NAND2_X1 U9219 ( .A1(n9151), .A2(n9149), .ZN(n9227) );
  OR2_X1 U9220 ( .A1(n9149), .A2(n9151), .ZN(n9225) );
  AND2_X1 U9221 ( .A1(n9228), .A2(n9229), .ZN(n9151) );
  NAND2_X1 U9222 ( .A1(n9147), .A2(n9230), .ZN(n9229) );
  OR2_X1 U9223 ( .A1(n9146), .A2(n9144), .ZN(n9230) );
  NOR2_X1 U9224 ( .A1(n8848), .A2(n7870), .ZN(n9147) );
  NAND2_X1 U9225 ( .A1(n9144), .A2(n9146), .ZN(n9228) );
  NAND2_X1 U9226 ( .A1(n9231), .A2(n9232), .ZN(n9146) );
  NAND3_X1 U9227 ( .A1(a_10_), .A2(n9233), .A3(b_24_), .ZN(n9232) );
  OR2_X1 U9228 ( .A1(n9142), .A2(n9140), .ZN(n9233) );
  NAND2_X1 U9229 ( .A1(n9140), .A2(n9142), .ZN(n9231) );
  NAND2_X1 U9230 ( .A1(n9138), .A2(n9234), .ZN(n9142) );
  NAND2_X1 U9231 ( .A1(n9137), .A2(n9139), .ZN(n9234) );
  NAND2_X1 U9232 ( .A1(n9235), .A2(n9236), .ZN(n9139) );
  NAND2_X1 U9233 ( .A1(b_24_), .A2(a_11_), .ZN(n9236) );
  INV_X1 U9234 ( .A(n9237), .ZN(n9235) );
  XNOR2_X1 U9235 ( .A(n9238), .B(n9239), .ZN(n9137) );
  XNOR2_X1 U9236 ( .A(n9240), .B(n9241), .ZN(n9238) );
  NOR2_X1 U9237 ( .A1(n8020), .A2(n9071), .ZN(n9241) );
  NAND2_X1 U9238 ( .A1(a_11_), .A2(n9237), .ZN(n9138) );
  NAND2_X1 U9239 ( .A1(n9242), .A2(n9243), .ZN(n9237) );
  NAND3_X1 U9240 ( .A1(a_12_), .A2(n9244), .A3(b_24_), .ZN(n9243) );
  OR2_X1 U9241 ( .A1(n9134), .A2(n9132), .ZN(n9244) );
  NAND2_X1 U9242 ( .A1(n9132), .A2(n9134), .ZN(n9242) );
  NAND2_X1 U9243 ( .A1(n9245), .A2(n9246), .ZN(n9134) );
  NAND2_X1 U9244 ( .A1(n9131), .A2(n9247), .ZN(n9246) );
  NAND2_X1 U9245 ( .A1(n9130), .A2(n9129), .ZN(n9247) );
  NOR2_X1 U9246 ( .A1(n8848), .A2(n7355), .ZN(n9131) );
  OR2_X1 U9247 ( .A1(n9129), .A2(n9130), .ZN(n9245) );
  AND2_X1 U9248 ( .A1(n9248), .A2(n9249), .ZN(n9130) );
  NAND3_X1 U9249 ( .A1(a_14_), .A2(n9250), .A3(b_24_), .ZN(n9249) );
  NAND2_X1 U9250 ( .A1(n9127), .A2(n9125), .ZN(n9250) );
  OR2_X1 U9251 ( .A1(n9125), .A2(n9127), .ZN(n9248) );
  AND2_X1 U9252 ( .A1(n9251), .A2(n9252), .ZN(n9127) );
  NAND2_X1 U9253 ( .A1(n9123), .A2(n9253), .ZN(n9252) );
  OR2_X1 U9254 ( .A1(n9122), .A2(n9120), .ZN(n9253) );
  NOR2_X1 U9255 ( .A1(n8848), .A2(n7346), .ZN(n9123) );
  NAND2_X1 U9256 ( .A1(n9120), .A2(n9122), .ZN(n9251) );
  NAND2_X1 U9257 ( .A1(n9254), .A2(n9255), .ZN(n9122) );
  NAND3_X1 U9258 ( .A1(a_16_), .A2(n9256), .A3(b_24_), .ZN(n9255) );
  OR2_X1 U9259 ( .A1(n9118), .A2(n9116), .ZN(n9256) );
  NAND2_X1 U9260 ( .A1(n9116), .A2(n9118), .ZN(n9254) );
  NAND2_X1 U9261 ( .A1(n9257), .A2(n9258), .ZN(n9118) );
  NAND2_X1 U9262 ( .A1(n9115), .A2(n9259), .ZN(n9258) );
  OR2_X1 U9263 ( .A1(n9114), .A2(n9113), .ZN(n9259) );
  NOR2_X1 U9264 ( .A1(n8848), .A2(n7337), .ZN(n9115) );
  NAND2_X1 U9265 ( .A1(n9113), .A2(n9114), .ZN(n9257) );
  NAND2_X1 U9266 ( .A1(n9260), .A2(n9261), .ZN(n9114) );
  NAND3_X1 U9267 ( .A1(a_18_), .A2(n9262), .A3(b_24_), .ZN(n9261) );
  NAND2_X1 U9268 ( .A1(n9110), .A2(n9109), .ZN(n9262) );
  OR2_X1 U9269 ( .A1(n9109), .A2(n9110), .ZN(n9260) );
  AND2_X1 U9270 ( .A1(n9263), .A2(n9264), .ZN(n9110) );
  NAND2_X1 U9271 ( .A1(n9107), .A2(n9265), .ZN(n9264) );
  OR2_X1 U9272 ( .A1(n9106), .A2(n9104), .ZN(n9265) );
  NOR2_X1 U9273 ( .A1(n8848), .A2(n7902), .ZN(n9107) );
  NAND2_X1 U9274 ( .A1(n9104), .A2(n9106), .ZN(n9263) );
  NAND2_X1 U9275 ( .A1(n9266), .A2(n9267), .ZN(n9106) );
  NAND3_X1 U9276 ( .A1(a_20_), .A2(n9268), .A3(b_24_), .ZN(n9267) );
  NAND2_X1 U9277 ( .A1(n9102), .A2(n9101), .ZN(n9268) );
  OR2_X1 U9278 ( .A1(n9101), .A2(n9102), .ZN(n9266) );
  AND2_X1 U9279 ( .A1(n9269), .A2(n9270), .ZN(n9102) );
  NAND2_X1 U9280 ( .A1(n9099), .A2(n9271), .ZN(n9270) );
  OR2_X1 U9281 ( .A1(n9098), .A2(n9097), .ZN(n9271) );
  NOR2_X1 U9282 ( .A1(n8848), .A2(n7909), .ZN(n9099) );
  NAND2_X1 U9283 ( .A1(n9097), .A2(n9098), .ZN(n9269) );
  NAND2_X1 U9284 ( .A1(n9272), .A2(n9273), .ZN(n9098) );
  NAND3_X1 U9285 ( .A1(a_22_), .A2(n9274), .A3(b_24_), .ZN(n9273) );
  OR2_X1 U9286 ( .A1(n9094), .A2(n9092), .ZN(n9274) );
  NAND2_X1 U9287 ( .A1(n9092), .A2(n9094), .ZN(n9272) );
  NAND2_X1 U9288 ( .A1(n9275), .A2(n9276), .ZN(n9094) );
  NAND2_X1 U9289 ( .A1(n9091), .A2(n9277), .ZN(n9276) );
  OR2_X1 U9290 ( .A1(n9090), .A2(n9088), .ZN(n9277) );
  NOR2_X1 U9291 ( .A1(n8848), .A2(n7916), .ZN(n9091) );
  NAND2_X1 U9292 ( .A1(n9088), .A2(n9090), .ZN(n9275) );
  NAND2_X1 U9293 ( .A1(n9278), .A2(n9279), .ZN(n9090) );
  NAND2_X1 U9294 ( .A1(n9087), .A2(n9280), .ZN(n9279) );
  NAND2_X1 U9295 ( .A1(n9086), .A2(n9085), .ZN(n9280) );
  OR2_X1 U9296 ( .A1(n9085), .A2(n9086), .ZN(n9278) );
  AND2_X1 U9297 ( .A1(n9281), .A2(n9282), .ZN(n9086) );
  NAND2_X1 U9298 ( .A1(n9083), .A2(n9283), .ZN(n9282) );
  OR2_X1 U9299 ( .A1(n9082), .A2(n9081), .ZN(n9283) );
  NOR2_X1 U9300 ( .A1(n8848), .A2(n7923), .ZN(n9083) );
  NAND2_X1 U9301 ( .A1(n9081), .A2(n9082), .ZN(n9281) );
  NAND2_X1 U9302 ( .A1(n9078), .A2(n9284), .ZN(n9082) );
  NAND2_X1 U9303 ( .A1(n9077), .A2(n9079), .ZN(n9284) );
  NAND2_X1 U9304 ( .A1(n9285), .A2(n9286), .ZN(n9079) );
  NAND2_X1 U9305 ( .A1(b_24_), .A2(a_26_), .ZN(n9286) );
  INV_X1 U9306 ( .A(n9287), .ZN(n9285) );
  XNOR2_X1 U9307 ( .A(n9288), .B(n9289), .ZN(n9077) );
  NAND2_X1 U9308 ( .A1(n9290), .A2(n9291), .ZN(n9288) );
  NAND2_X1 U9309 ( .A1(a_26_), .A2(n9287), .ZN(n9078) );
  NAND2_X1 U9310 ( .A1(n9049), .A2(n9292), .ZN(n9287) );
  NAND2_X1 U9311 ( .A1(n9048), .A2(n9050), .ZN(n9292) );
  NAND2_X1 U9312 ( .A1(n9293), .A2(n9294), .ZN(n9050) );
  NAND2_X1 U9313 ( .A1(b_24_), .A2(a_27_), .ZN(n9294) );
  INV_X1 U9314 ( .A(n9295), .ZN(n9293) );
  XNOR2_X1 U9315 ( .A(n9296), .B(n9297), .ZN(n9048) );
  XOR2_X1 U9316 ( .A(n9298), .B(n9299), .Z(n9296) );
  NAND2_X1 U9317 ( .A1(b_23_), .A2(a_28_), .ZN(n9298) );
  NAND2_X1 U9318 ( .A1(a_27_), .A2(n9295), .ZN(n9049) );
  NAND2_X1 U9319 ( .A1(n9300), .A2(n9301), .ZN(n9295) );
  NAND3_X1 U9320 ( .A1(a_28_), .A2(n9302), .A3(b_24_), .ZN(n9301) );
  NAND2_X1 U9321 ( .A1(n9058), .A2(n9056), .ZN(n9302) );
  OR2_X1 U9322 ( .A1(n9056), .A2(n9058), .ZN(n9300) );
  AND2_X1 U9323 ( .A1(n9303), .A2(n9304), .ZN(n9058) );
  NAND2_X1 U9324 ( .A1(n9073), .A2(n9305), .ZN(n9304) );
  OR2_X1 U9325 ( .A1(n9074), .A2(n9075), .ZN(n9305) );
  NOR2_X1 U9326 ( .A1(n8848), .A2(n7946), .ZN(n9073) );
  NAND2_X1 U9327 ( .A1(n9075), .A2(n9074), .ZN(n9303) );
  NAND2_X1 U9328 ( .A1(n9306), .A2(n9307), .ZN(n9074) );
  NAND2_X1 U9329 ( .A1(b_22_), .A2(n9308), .ZN(n9307) );
  NAND2_X1 U9330 ( .A1(n7268), .A2(n9309), .ZN(n9308) );
  NAND2_X1 U9331 ( .A1(a_31_), .A2(n9071), .ZN(n9309) );
  NAND2_X1 U9332 ( .A1(b_23_), .A2(n9310), .ZN(n9306) );
  NAND2_X1 U9333 ( .A1(n7272), .A2(n9311), .ZN(n9310) );
  NAND2_X1 U9334 ( .A1(a_30_), .A2(n9312), .ZN(n9311) );
  AND3_X1 U9335 ( .A1(b_23_), .A2(n7954), .A3(b_24_), .ZN(n9075) );
  XNOR2_X1 U9336 ( .A(n9313), .B(n9314), .ZN(n9056) );
  XOR2_X1 U9337 ( .A(n9315), .B(n9316), .Z(n9313) );
  XNOR2_X1 U9338 ( .A(n9317), .B(n9318), .ZN(n9081) );
  NAND2_X1 U9339 ( .A1(n9319), .A2(n9320), .ZN(n9317) );
  XNOR2_X1 U9340 ( .A(n9321), .B(n9322), .ZN(n9085) );
  XOR2_X1 U9341 ( .A(n9323), .B(n9324), .Z(n9321) );
  XNOR2_X1 U9342 ( .A(n9325), .B(n9326), .ZN(n9088) );
  XNOR2_X1 U9343 ( .A(n9327), .B(n9328), .ZN(n9325) );
  NOR2_X1 U9344 ( .A1(n7691), .A2(n9071), .ZN(n9328) );
  XNOR2_X1 U9345 ( .A(n9329), .B(n9330), .ZN(n9092) );
  XNOR2_X1 U9346 ( .A(n9331), .B(n9332), .ZN(n9330) );
  XNOR2_X1 U9347 ( .A(n9333), .B(n9334), .ZN(n9097) );
  XOR2_X1 U9348 ( .A(n9335), .B(n9336), .Z(n9334) );
  NAND2_X1 U9349 ( .A1(b_23_), .A2(a_22_), .ZN(n9336) );
  XNOR2_X1 U9350 ( .A(n9337), .B(n9338), .ZN(n9101) );
  XOR2_X1 U9351 ( .A(n9339), .B(n9340), .Z(n9337) );
  XNOR2_X1 U9352 ( .A(n9341), .B(n9342), .ZN(n9104) );
  XNOR2_X1 U9353 ( .A(n9343), .B(n9344), .ZN(n9341) );
  NOR2_X1 U9354 ( .A1(n7987), .A2(n9071), .ZN(n9344) );
  XOR2_X1 U9355 ( .A(n9345), .B(n9346), .Z(n9109) );
  XNOR2_X1 U9356 ( .A(n9347), .B(n9348), .ZN(n9346) );
  XNOR2_X1 U9357 ( .A(n9349), .B(n9350), .ZN(n9113) );
  XNOR2_X1 U9358 ( .A(n9351), .B(n9352), .ZN(n9349) );
  NOR2_X1 U9359 ( .A1(n7764), .A2(n9071), .ZN(n9352) );
  XNOR2_X1 U9360 ( .A(n9353), .B(n9354), .ZN(n9116) );
  XNOR2_X1 U9361 ( .A(n9355), .B(n9356), .ZN(n9353) );
  XNOR2_X1 U9362 ( .A(n9357), .B(n9358), .ZN(n9120) );
  XOR2_X1 U9363 ( .A(n9359), .B(n9360), .Z(n9358) );
  NAND2_X1 U9364 ( .A1(b_23_), .A2(a_16_), .ZN(n9360) );
  XOR2_X1 U9365 ( .A(n9361), .B(n9362), .Z(n9125) );
  XOR2_X1 U9366 ( .A(n9363), .B(n9364), .Z(n9362) );
  NAND2_X1 U9367 ( .A1(b_23_), .A2(a_15_), .ZN(n9364) );
  XOR2_X1 U9368 ( .A(n9365), .B(n9366), .Z(n9129) );
  NAND2_X1 U9369 ( .A1(n9367), .A2(n9368), .ZN(n9365) );
  XOR2_X1 U9370 ( .A(n9369), .B(n9370), .Z(n9132) );
  XOR2_X1 U9371 ( .A(n9371), .B(n9372), .Z(n9369) );
  XOR2_X1 U9372 ( .A(n9373), .B(n9374), .Z(n9140) );
  XOR2_X1 U9373 ( .A(n9375), .B(n9376), .Z(n9373) );
  NOR2_X1 U9374 ( .A1(n7877), .A2(n9071), .ZN(n9376) );
  XNOR2_X1 U9375 ( .A(n9377), .B(n9378), .ZN(n9144) );
  NAND2_X1 U9376 ( .A1(n9379), .A2(n9380), .ZN(n9377) );
  XOR2_X1 U9377 ( .A(n9381), .B(n9382), .Z(n9149) );
  XNOR2_X1 U9378 ( .A(n9383), .B(n9384), .ZN(n9382) );
  NAND2_X1 U9379 ( .A1(n9159), .A2(n9158), .ZN(n9214) );
  XNOR2_X1 U9380 ( .A(n9385), .B(n9386), .ZN(n9158) );
  XOR2_X1 U9381 ( .A(n9387), .B(n9388), .Z(n9386) );
  NAND2_X1 U9382 ( .A1(b_23_), .A2(a_7_), .ZN(n9388) );
  NOR2_X1 U9383 ( .A1(n8848), .A2(n7388), .ZN(n9159) );
  XOR2_X1 U9384 ( .A(n9389), .B(n9390), .Z(n9162) );
  NAND2_X1 U9385 ( .A1(n9391), .A2(n9392), .ZN(n9389) );
  XNOR2_X1 U9386 ( .A(n9393), .B(n9394), .ZN(n9166) );
  XOR2_X1 U9387 ( .A(n9395), .B(n9396), .Z(n9393) );
  NOR2_X1 U9388 ( .A1(n7393), .A2(n9071), .ZN(n9396) );
  NAND2_X1 U9389 ( .A1(n9397), .A2(n9398), .ZN(n9189) );
  INV_X1 U9390 ( .A(n9177), .ZN(n9398) );
  XOR2_X1 U9391 ( .A(n9399), .B(n9400), .Z(n9177) );
  XOR2_X1 U9392 ( .A(n9401), .B(n9402), .Z(n9400) );
  NAND2_X1 U9393 ( .A1(b_23_), .A2(a_2_), .ZN(n9402) );
  INV_X1 U9394 ( .A(n9180), .ZN(n9397) );
  NAND2_X1 U9395 ( .A1(b_24_), .A2(a_1_), .ZN(n9180) );
  XNOR2_X1 U9396 ( .A(n9403), .B(n9404), .ZN(n9182) );
  XOR2_X1 U9397 ( .A(n9405), .B(n9406), .Z(n9404) );
  NAND2_X1 U9398 ( .A1(b_23_), .A2(a_1_), .ZN(n9406) );
  INV_X1 U9399 ( .A(n7586), .ZN(n7581) );
  XOR2_X1 U9400 ( .A(n9407), .B(n9408), .Z(n7586) );
  XOR2_X1 U9401 ( .A(n9409), .B(n9410), .Z(n9408) );
  NAND2_X1 U9402 ( .A1(b_23_), .A2(a_0_), .ZN(n9410) );
  NAND3_X1 U9403 ( .A1(n9411), .A2(n7577), .A3(n7576), .ZN(n7455) );
  XNOR2_X1 U9404 ( .A(n9412), .B(n9413), .ZN(n7576) );
  NAND2_X1 U9405 ( .A1(n9414), .A2(n9415), .ZN(n9412) );
  NAND2_X1 U9406 ( .A1(n9416), .A2(n9417), .ZN(n7577) );
  NAND3_X1 U9407 ( .A1(a_0_), .A2(n9418), .A3(b_23_), .ZN(n9417) );
  OR2_X1 U9408 ( .A1(n9409), .A2(n9407), .ZN(n9418) );
  NAND2_X1 U9409 ( .A1(n9407), .A2(n9409), .ZN(n9416) );
  NAND2_X1 U9410 ( .A1(n9419), .A2(n9420), .ZN(n9409) );
  NAND3_X1 U9411 ( .A1(a_1_), .A2(n9421), .A3(b_23_), .ZN(n9420) );
  OR2_X1 U9412 ( .A1(n9405), .A2(n9403), .ZN(n9421) );
  NAND2_X1 U9413 ( .A1(n9403), .A2(n9405), .ZN(n9419) );
  NAND2_X1 U9414 ( .A1(n9422), .A2(n9423), .ZN(n9405) );
  NAND3_X1 U9415 ( .A1(a_2_), .A2(n9424), .A3(b_23_), .ZN(n9423) );
  OR2_X1 U9416 ( .A1(n9401), .A2(n9399), .ZN(n9424) );
  NAND2_X1 U9417 ( .A1(n9399), .A2(n9401), .ZN(n9422) );
  NAND2_X1 U9418 ( .A1(n9425), .A2(n9426), .ZN(n9401) );
  NAND3_X1 U9419 ( .A1(a_3_), .A2(n9427), .A3(b_23_), .ZN(n9426) );
  OR2_X1 U9420 ( .A1(n9198), .A2(n9196), .ZN(n9427) );
  NAND2_X1 U9421 ( .A1(n9196), .A2(n9198), .ZN(n9425) );
  NAND2_X1 U9422 ( .A1(n9428), .A2(n9429), .ZN(n9198) );
  NAND3_X1 U9423 ( .A1(a_4_), .A2(n9430), .A3(b_23_), .ZN(n9429) );
  OR2_X1 U9424 ( .A1(n9206), .A2(n9204), .ZN(n9430) );
  NAND2_X1 U9425 ( .A1(n9204), .A2(n9206), .ZN(n9428) );
  NAND2_X1 U9426 ( .A1(n9431), .A2(n9432), .ZN(n9206) );
  NAND3_X1 U9427 ( .A1(a_5_), .A2(n9433), .A3(b_23_), .ZN(n9432) );
  OR2_X1 U9428 ( .A1(n9395), .A2(n9394), .ZN(n9433) );
  NAND2_X1 U9429 ( .A1(n9394), .A2(n9395), .ZN(n9431) );
  NAND2_X1 U9430 ( .A1(n9391), .A2(n9434), .ZN(n9395) );
  NAND2_X1 U9431 ( .A1(n9390), .A2(n9392), .ZN(n9434) );
  NAND2_X1 U9432 ( .A1(n9435), .A2(n9436), .ZN(n9392) );
  NAND2_X1 U9433 ( .A1(b_23_), .A2(a_6_), .ZN(n9436) );
  INV_X1 U9434 ( .A(n9437), .ZN(n9435) );
  XNOR2_X1 U9435 ( .A(n9438), .B(n9439), .ZN(n9390) );
  XNOR2_X1 U9436 ( .A(n9440), .B(n9441), .ZN(n9439) );
  NAND2_X1 U9437 ( .A1(a_6_), .A2(n9437), .ZN(n9391) );
  NAND2_X1 U9438 ( .A1(n9442), .A2(n9443), .ZN(n9437) );
  NAND3_X1 U9439 ( .A1(a_7_), .A2(n9444), .A3(b_23_), .ZN(n9443) );
  OR2_X1 U9440 ( .A1(n9387), .A2(n9385), .ZN(n9444) );
  NAND2_X1 U9441 ( .A1(n9385), .A2(n9387), .ZN(n9442) );
  NAND2_X1 U9442 ( .A1(n9445), .A2(n9446), .ZN(n9387) );
  NAND2_X1 U9443 ( .A1(n9224), .A2(n9447), .ZN(n9446) );
  OR2_X1 U9444 ( .A1(n9223), .A2(n9221), .ZN(n9447) );
  NOR2_X1 U9445 ( .A1(n9071), .A2(n8037), .ZN(n9224) );
  NAND2_X1 U9446 ( .A1(n9221), .A2(n9223), .ZN(n9445) );
  NAND2_X1 U9447 ( .A1(n9448), .A2(n9449), .ZN(n9223) );
  NAND2_X1 U9448 ( .A1(n9384), .A2(n9450), .ZN(n9449) );
  OR2_X1 U9449 ( .A1(n9383), .A2(n9381), .ZN(n9450) );
  NOR2_X1 U9450 ( .A1(n9071), .A2(n7870), .ZN(n9384) );
  NAND2_X1 U9451 ( .A1(n9381), .A2(n9383), .ZN(n9448) );
  NAND2_X1 U9452 ( .A1(n9379), .A2(n9451), .ZN(n9383) );
  NAND2_X1 U9453 ( .A1(n9378), .A2(n9380), .ZN(n9451) );
  NAND2_X1 U9454 ( .A1(n9452), .A2(n9453), .ZN(n9380) );
  NAND2_X1 U9455 ( .A1(b_23_), .A2(a_10_), .ZN(n9453) );
  INV_X1 U9456 ( .A(n9454), .ZN(n9452) );
  XNOR2_X1 U9457 ( .A(n9455), .B(n9456), .ZN(n9378) );
  XNOR2_X1 U9458 ( .A(n9457), .B(n9458), .ZN(n9456) );
  NAND2_X1 U9459 ( .A1(a_10_), .A2(n9454), .ZN(n9379) );
  NAND2_X1 U9460 ( .A1(n9459), .A2(n9460), .ZN(n9454) );
  NAND3_X1 U9461 ( .A1(a_11_), .A2(n9461), .A3(b_23_), .ZN(n9460) );
  OR2_X1 U9462 ( .A1(n9375), .A2(n9374), .ZN(n9461) );
  NAND2_X1 U9463 ( .A1(n9374), .A2(n9375), .ZN(n9459) );
  NAND2_X1 U9464 ( .A1(n9462), .A2(n9463), .ZN(n9375) );
  NAND3_X1 U9465 ( .A1(a_12_), .A2(n9464), .A3(b_23_), .ZN(n9463) );
  NAND2_X1 U9466 ( .A1(n9240), .A2(n9239), .ZN(n9464) );
  OR2_X1 U9467 ( .A1(n9239), .A2(n9240), .ZN(n9462) );
  AND2_X1 U9468 ( .A1(n9465), .A2(n9466), .ZN(n9240) );
  NAND2_X1 U9469 ( .A1(n9372), .A2(n9467), .ZN(n9466) );
  OR2_X1 U9470 ( .A1(n9371), .A2(n9370), .ZN(n9467) );
  NOR2_X1 U9471 ( .A1(n9071), .A2(n7355), .ZN(n9372) );
  NAND2_X1 U9472 ( .A1(n9370), .A2(n9371), .ZN(n9465) );
  NAND2_X1 U9473 ( .A1(n9367), .A2(n9468), .ZN(n9371) );
  NAND2_X1 U9474 ( .A1(n9366), .A2(n9368), .ZN(n9468) );
  NAND2_X1 U9475 ( .A1(n9469), .A2(n9470), .ZN(n9368) );
  NAND2_X1 U9476 ( .A1(b_23_), .A2(a_14_), .ZN(n9470) );
  INV_X1 U9477 ( .A(n9471), .ZN(n9469) );
  XNOR2_X1 U9478 ( .A(n9472), .B(n9473), .ZN(n9366) );
  XNOR2_X1 U9479 ( .A(n9474), .B(n9475), .ZN(n9473) );
  NAND2_X1 U9480 ( .A1(a_14_), .A2(n9471), .ZN(n9367) );
  NAND2_X1 U9481 ( .A1(n9476), .A2(n9477), .ZN(n9471) );
  NAND3_X1 U9482 ( .A1(a_15_), .A2(n9478), .A3(b_23_), .ZN(n9477) );
  OR2_X1 U9483 ( .A1(n9363), .A2(n9361), .ZN(n9478) );
  NAND2_X1 U9484 ( .A1(n9361), .A2(n9363), .ZN(n9476) );
  NAND2_X1 U9485 ( .A1(n9479), .A2(n9480), .ZN(n9363) );
  NAND3_X1 U9486 ( .A1(a_16_), .A2(n9481), .A3(b_23_), .ZN(n9480) );
  OR2_X1 U9487 ( .A1(n9359), .A2(n9357), .ZN(n9481) );
  NAND2_X1 U9488 ( .A1(n9357), .A2(n9359), .ZN(n9479) );
  NAND2_X1 U9489 ( .A1(n9482), .A2(n9483), .ZN(n9359) );
  NAND2_X1 U9490 ( .A1(n9356), .A2(n9484), .ZN(n9483) );
  NAND2_X1 U9491 ( .A1(n9355), .A2(n9354), .ZN(n9484) );
  NOR2_X1 U9492 ( .A1(n9071), .A2(n7337), .ZN(n9356) );
  OR2_X1 U9493 ( .A1(n9354), .A2(n9355), .ZN(n9482) );
  AND2_X1 U9494 ( .A1(n9485), .A2(n9486), .ZN(n9355) );
  NAND3_X1 U9495 ( .A1(a_18_), .A2(n9487), .A3(b_23_), .ZN(n9486) );
  NAND2_X1 U9496 ( .A1(n9351), .A2(n9350), .ZN(n9487) );
  OR2_X1 U9497 ( .A1(n9350), .A2(n9351), .ZN(n9485) );
  AND2_X1 U9498 ( .A1(n9488), .A2(n9489), .ZN(n9351) );
  NAND2_X1 U9499 ( .A1(n9348), .A2(n9490), .ZN(n9489) );
  OR2_X1 U9500 ( .A1(n9347), .A2(n9345), .ZN(n9490) );
  NOR2_X1 U9501 ( .A1(n9071), .A2(n7902), .ZN(n9348) );
  NAND2_X1 U9502 ( .A1(n9345), .A2(n9347), .ZN(n9488) );
  NAND2_X1 U9503 ( .A1(n9491), .A2(n9492), .ZN(n9347) );
  NAND3_X1 U9504 ( .A1(a_20_), .A2(n9493), .A3(b_23_), .ZN(n9492) );
  NAND2_X1 U9505 ( .A1(n9343), .A2(n9342), .ZN(n9493) );
  OR2_X1 U9506 ( .A1(n9342), .A2(n9343), .ZN(n9491) );
  AND2_X1 U9507 ( .A1(n9494), .A2(n9495), .ZN(n9343) );
  NAND2_X1 U9508 ( .A1(n9340), .A2(n9496), .ZN(n9495) );
  OR2_X1 U9509 ( .A1(n9339), .A2(n9338), .ZN(n9496) );
  NOR2_X1 U9510 ( .A1(n9071), .A2(n7909), .ZN(n9340) );
  NAND2_X1 U9511 ( .A1(n9338), .A2(n9339), .ZN(n9494) );
  NAND2_X1 U9512 ( .A1(n9497), .A2(n9498), .ZN(n9339) );
  NAND3_X1 U9513 ( .A1(a_22_), .A2(n9499), .A3(b_23_), .ZN(n9498) );
  OR2_X1 U9514 ( .A1(n9335), .A2(n9333), .ZN(n9499) );
  NAND2_X1 U9515 ( .A1(n9333), .A2(n9335), .ZN(n9497) );
  NAND2_X1 U9516 ( .A1(n9500), .A2(n9501), .ZN(n9335) );
  NAND2_X1 U9517 ( .A1(n9332), .A2(n9502), .ZN(n9501) );
  OR2_X1 U9518 ( .A1(n9331), .A2(n9329), .ZN(n9502) );
  NAND2_X1 U9519 ( .A1(n9329), .A2(n9331), .ZN(n9500) );
  NAND2_X1 U9520 ( .A1(n9503), .A2(n9504), .ZN(n9331) );
  NAND3_X1 U9521 ( .A1(a_24_), .A2(n9505), .A3(b_23_), .ZN(n9504) );
  NAND2_X1 U9522 ( .A1(n9327), .A2(n9326), .ZN(n9505) );
  OR2_X1 U9523 ( .A1(n9326), .A2(n9327), .ZN(n9503) );
  AND2_X1 U9524 ( .A1(n9506), .A2(n9507), .ZN(n9327) );
  NAND2_X1 U9525 ( .A1(n9324), .A2(n9508), .ZN(n9507) );
  OR2_X1 U9526 ( .A1(n9323), .A2(n9322), .ZN(n9508) );
  NOR2_X1 U9527 ( .A1(n9071), .A2(n7923), .ZN(n9324) );
  NAND2_X1 U9528 ( .A1(n9322), .A2(n9323), .ZN(n9506) );
  NAND2_X1 U9529 ( .A1(n9319), .A2(n9509), .ZN(n9323) );
  NAND2_X1 U9530 ( .A1(n9318), .A2(n9320), .ZN(n9509) );
  NAND2_X1 U9531 ( .A1(n9510), .A2(n9511), .ZN(n9320) );
  NAND2_X1 U9532 ( .A1(b_23_), .A2(a_26_), .ZN(n9511) );
  INV_X1 U9533 ( .A(n9512), .ZN(n9510) );
  XNOR2_X1 U9534 ( .A(n9513), .B(n9514), .ZN(n9318) );
  NAND2_X1 U9535 ( .A1(n9515), .A2(n9516), .ZN(n9513) );
  NAND2_X1 U9536 ( .A1(a_26_), .A2(n9512), .ZN(n9319) );
  NAND2_X1 U9537 ( .A1(n9290), .A2(n9517), .ZN(n9512) );
  NAND2_X1 U9538 ( .A1(n9289), .A2(n9291), .ZN(n9517) );
  NAND2_X1 U9539 ( .A1(n9518), .A2(n9519), .ZN(n9291) );
  NAND2_X1 U9540 ( .A1(b_23_), .A2(a_27_), .ZN(n9519) );
  INV_X1 U9541 ( .A(n9520), .ZN(n9518) );
  XNOR2_X1 U9542 ( .A(n9521), .B(n9522), .ZN(n9289) );
  XOR2_X1 U9543 ( .A(n9523), .B(n9524), .Z(n9521) );
  NAND2_X1 U9544 ( .A1(b_22_), .A2(a_28_), .ZN(n9523) );
  NAND2_X1 U9545 ( .A1(a_27_), .A2(n9520), .ZN(n9290) );
  NAND2_X1 U9546 ( .A1(n9525), .A2(n9526), .ZN(n9520) );
  NAND3_X1 U9547 ( .A1(a_28_), .A2(n9527), .A3(b_23_), .ZN(n9526) );
  NAND2_X1 U9548 ( .A1(n9299), .A2(n9297), .ZN(n9527) );
  OR2_X1 U9549 ( .A1(n9297), .A2(n9299), .ZN(n9525) );
  AND2_X1 U9550 ( .A1(n9528), .A2(n9529), .ZN(n9299) );
  NAND2_X1 U9551 ( .A1(n9314), .A2(n9530), .ZN(n9529) );
  OR2_X1 U9552 ( .A1(n9315), .A2(n9316), .ZN(n9530) );
  NOR2_X1 U9553 ( .A1(n9071), .A2(n7946), .ZN(n9314) );
  NAND2_X1 U9554 ( .A1(n9316), .A2(n9315), .ZN(n9528) );
  NAND2_X1 U9555 ( .A1(n9531), .A2(n9532), .ZN(n9315) );
  NAND2_X1 U9556 ( .A1(b_21_), .A2(n9533), .ZN(n9532) );
  NAND2_X1 U9557 ( .A1(n7268), .A2(n9534), .ZN(n9533) );
  NAND2_X1 U9558 ( .A1(a_31_), .A2(n9312), .ZN(n9534) );
  NAND2_X1 U9559 ( .A1(b_22_), .A2(n9535), .ZN(n9531) );
  NAND2_X1 U9560 ( .A1(n7272), .A2(n9536), .ZN(n9535) );
  NAND2_X1 U9561 ( .A1(a_30_), .A2(n9537), .ZN(n9536) );
  AND3_X1 U9562 ( .A1(b_22_), .A2(n7954), .A3(b_23_), .ZN(n9316) );
  XNOR2_X1 U9563 ( .A(n9538), .B(n9539), .ZN(n9297) );
  XOR2_X1 U9564 ( .A(n9540), .B(n9541), .Z(n9538) );
  XNOR2_X1 U9565 ( .A(n9542), .B(n9543), .ZN(n9322) );
  NAND2_X1 U9566 ( .A1(n9544), .A2(n9545), .ZN(n9542) );
  XNOR2_X1 U9567 ( .A(n9546), .B(n9547), .ZN(n9326) );
  XOR2_X1 U9568 ( .A(n9548), .B(n9549), .Z(n9546) );
  XNOR2_X1 U9569 ( .A(n9550), .B(n9551), .ZN(n9329) );
  XNOR2_X1 U9570 ( .A(n9552), .B(n9553), .ZN(n9550) );
  NOR2_X1 U9571 ( .A1(n7691), .A2(n9312), .ZN(n9553) );
  XNOR2_X1 U9572 ( .A(n9554), .B(n9555), .ZN(n9333) );
  XNOR2_X1 U9573 ( .A(n9556), .B(n9557), .ZN(n9555) );
  XNOR2_X1 U9574 ( .A(n9558), .B(n9559), .ZN(n9338) );
  XNOR2_X1 U9575 ( .A(n9560), .B(n9561), .ZN(n9558) );
  XNOR2_X1 U9576 ( .A(n9562), .B(n9563), .ZN(n9342) );
  XOR2_X1 U9577 ( .A(n9564), .B(n9565), .Z(n9562) );
  XNOR2_X1 U9578 ( .A(n9566), .B(n9567), .ZN(n9345) );
  XNOR2_X1 U9579 ( .A(n9568), .B(n9569), .ZN(n9566) );
  NOR2_X1 U9580 ( .A1(n7987), .A2(n9312), .ZN(n9569) );
  XOR2_X1 U9581 ( .A(n9570), .B(n9571), .Z(n9350) );
  XNOR2_X1 U9582 ( .A(n9572), .B(n9573), .ZN(n9571) );
  XNOR2_X1 U9583 ( .A(n9574), .B(n9575), .ZN(n9354) );
  XOR2_X1 U9584 ( .A(n9576), .B(n9577), .Z(n9574) );
  NOR2_X1 U9585 ( .A1(n7764), .A2(n9312), .ZN(n9577) );
  XOR2_X1 U9586 ( .A(n9578), .B(n9579), .Z(n9357) );
  XOR2_X1 U9587 ( .A(n9580), .B(n9581), .Z(n9578) );
  XNOR2_X1 U9588 ( .A(n9582), .B(n9583), .ZN(n9361) );
  XOR2_X1 U9589 ( .A(n9584), .B(n9585), .Z(n9583) );
  NAND2_X1 U9590 ( .A1(b_22_), .A2(a_16_), .ZN(n9585) );
  XNOR2_X1 U9591 ( .A(n9586), .B(n9587), .ZN(n9370) );
  XNOR2_X1 U9592 ( .A(n9588), .B(n9589), .ZN(n9586) );
  NOR2_X1 U9593 ( .A1(n7782), .A2(n9312), .ZN(n9589) );
  XOR2_X1 U9594 ( .A(n9590), .B(n9591), .Z(n9239) );
  XNOR2_X1 U9595 ( .A(n9592), .B(n9593), .ZN(n9591) );
  XNOR2_X1 U9596 ( .A(n9594), .B(n9595), .ZN(n9374) );
  XNOR2_X1 U9597 ( .A(n9596), .B(n9597), .ZN(n9594) );
  NOR2_X1 U9598 ( .A1(n8020), .A2(n9312), .ZN(n9597) );
  XNOR2_X1 U9599 ( .A(n9598), .B(n9599), .ZN(n9381) );
  XNOR2_X1 U9600 ( .A(n9600), .B(n9601), .ZN(n9598) );
  NOR2_X1 U9601 ( .A1(n7799), .A2(n9312), .ZN(n9601) );
  XNOR2_X1 U9602 ( .A(n9602), .B(n9603), .ZN(n9221) );
  XNOR2_X1 U9603 ( .A(n9604), .B(n9605), .ZN(n9602) );
  NOR2_X1 U9604 ( .A1(n7870), .A2(n9312), .ZN(n9605) );
  XNOR2_X1 U9605 ( .A(n9606), .B(n9607), .ZN(n9385) );
  XNOR2_X1 U9606 ( .A(n9608), .B(n9609), .ZN(n9607) );
  XNOR2_X1 U9607 ( .A(n9610), .B(n9611), .ZN(n9394) );
  XNOR2_X1 U9608 ( .A(n9612), .B(n9613), .ZN(n9610) );
  XOR2_X1 U9609 ( .A(n9614), .B(n9615), .Z(n9204) );
  XOR2_X1 U9610 ( .A(n9616), .B(n9617), .Z(n9614) );
  NOR2_X1 U9611 ( .A1(n7393), .A2(n9312), .ZN(n9617) );
  XNOR2_X1 U9612 ( .A(n9618), .B(n9619), .ZN(n9196) );
  XNOR2_X1 U9613 ( .A(n9620), .B(n9621), .ZN(n9619) );
  XOR2_X1 U9614 ( .A(n9622), .B(n9623), .Z(n9399) );
  XOR2_X1 U9615 ( .A(n9624), .B(n9625), .Z(n9622) );
  XOR2_X1 U9616 ( .A(n9626), .B(n9627), .Z(n9403) );
  XOR2_X1 U9617 ( .A(n9628), .B(n9629), .Z(n9626) );
  XOR2_X1 U9618 ( .A(n9630), .B(n9631), .Z(n9407) );
  XOR2_X1 U9619 ( .A(n9632), .B(n9633), .Z(n9630) );
  NOR2_X1 U9620 ( .A1(n7411), .A2(n9312), .ZN(n9633) );
  XOR2_X1 U9621 ( .A(n7572), .B(n7571), .Z(n9411) );
  NAND4_X1 U9622 ( .A1(n7571), .A2(n7570), .A3(n7572), .A4(n7565), .ZN(n7459)
         );
  INV_X1 U9623 ( .A(n9634), .ZN(n7565) );
  NAND2_X1 U9624 ( .A1(n9414), .A2(n9635), .ZN(n7572) );
  NAND2_X1 U9625 ( .A1(n9413), .A2(n9415), .ZN(n9635) );
  NAND2_X1 U9626 ( .A1(n9636), .A2(n9637), .ZN(n9415) );
  NAND2_X1 U9627 ( .A1(b_22_), .A2(a_0_), .ZN(n9637) );
  INV_X1 U9628 ( .A(n9638), .ZN(n9636) );
  XOR2_X1 U9629 ( .A(n9639), .B(n9640), .Z(n9413) );
  XOR2_X1 U9630 ( .A(n9641), .B(n9642), .Z(n9639) );
  NOR2_X1 U9631 ( .A1(n7411), .A2(n9537), .ZN(n9642) );
  NAND2_X1 U9632 ( .A1(a_0_), .A2(n9638), .ZN(n9414) );
  NAND2_X1 U9633 ( .A1(n9643), .A2(n9644), .ZN(n9638) );
  NAND3_X1 U9634 ( .A1(a_1_), .A2(n9645), .A3(b_22_), .ZN(n9644) );
  OR2_X1 U9635 ( .A1(n9632), .A2(n9631), .ZN(n9645) );
  NAND2_X1 U9636 ( .A1(n9631), .A2(n9632), .ZN(n9643) );
  NAND2_X1 U9637 ( .A1(n9646), .A2(n9647), .ZN(n9632) );
  NAND2_X1 U9638 ( .A1(n9629), .A2(n9648), .ZN(n9647) );
  OR2_X1 U9639 ( .A1(n9628), .A2(n9627), .ZN(n9648) );
  NOR2_X1 U9640 ( .A1(n9312), .A2(n7832), .ZN(n9629) );
  NAND2_X1 U9641 ( .A1(n9627), .A2(n9628), .ZN(n9646) );
  NAND2_X1 U9642 ( .A1(n9649), .A2(n9650), .ZN(n9628) );
  NAND2_X1 U9643 ( .A1(n9625), .A2(n9651), .ZN(n9650) );
  OR2_X1 U9644 ( .A1(n9624), .A2(n9623), .ZN(n9651) );
  NOR2_X1 U9645 ( .A1(n9312), .A2(n7850), .ZN(n9625) );
  NAND2_X1 U9646 ( .A1(n9623), .A2(n9624), .ZN(n9649) );
  NAND2_X1 U9647 ( .A1(n9652), .A2(n9653), .ZN(n9624) );
  NAND2_X1 U9648 ( .A1(n9621), .A2(n9654), .ZN(n9653) );
  OR2_X1 U9649 ( .A1(n9620), .A2(n9618), .ZN(n9654) );
  NOR2_X1 U9650 ( .A1(n9312), .A2(n7398), .ZN(n9621) );
  NAND2_X1 U9651 ( .A1(n9618), .A2(n9620), .ZN(n9652) );
  NAND2_X1 U9652 ( .A1(n9655), .A2(n9656), .ZN(n9620) );
  NAND3_X1 U9653 ( .A1(a_5_), .A2(n9657), .A3(b_22_), .ZN(n9656) );
  OR2_X1 U9654 ( .A1(n9616), .A2(n9615), .ZN(n9657) );
  NAND2_X1 U9655 ( .A1(n9615), .A2(n9616), .ZN(n9655) );
  NAND2_X1 U9656 ( .A1(n9658), .A2(n9659), .ZN(n9616) );
  NAND2_X1 U9657 ( .A1(n9613), .A2(n9660), .ZN(n9659) );
  NAND2_X1 U9658 ( .A1(n9612), .A2(n9611), .ZN(n9660) );
  NOR2_X1 U9659 ( .A1(n9312), .A2(n7388), .ZN(n9613) );
  OR2_X1 U9660 ( .A1(n9611), .A2(n9612), .ZN(n9658) );
  AND2_X1 U9661 ( .A1(n9661), .A2(n9662), .ZN(n9612) );
  NAND2_X1 U9662 ( .A1(n9441), .A2(n9663), .ZN(n9662) );
  OR2_X1 U9663 ( .A1(n9440), .A2(n9438), .ZN(n9663) );
  NOR2_X1 U9664 ( .A1(n9312), .A2(n7863), .ZN(n9441) );
  NAND2_X1 U9665 ( .A1(n9438), .A2(n9440), .ZN(n9661) );
  NAND2_X1 U9666 ( .A1(n9664), .A2(n9665), .ZN(n9440) );
  NAND2_X1 U9667 ( .A1(n9609), .A2(n9666), .ZN(n9665) );
  OR2_X1 U9668 ( .A1(n9608), .A2(n9606), .ZN(n9666) );
  NOR2_X1 U9669 ( .A1(n9312), .A2(n8037), .ZN(n9609) );
  NAND2_X1 U9670 ( .A1(n9606), .A2(n9608), .ZN(n9664) );
  NAND2_X1 U9671 ( .A1(n9667), .A2(n9668), .ZN(n9608) );
  NAND3_X1 U9672 ( .A1(a_9_), .A2(n9669), .A3(b_22_), .ZN(n9668) );
  NAND2_X1 U9673 ( .A1(n9604), .A2(n9603), .ZN(n9669) );
  OR2_X1 U9674 ( .A1(n9603), .A2(n9604), .ZN(n9667) );
  AND2_X1 U9675 ( .A1(n9670), .A2(n9671), .ZN(n9604) );
  NAND3_X1 U9676 ( .A1(a_10_), .A2(n9672), .A3(b_22_), .ZN(n9671) );
  NAND2_X1 U9677 ( .A1(n9600), .A2(n9599), .ZN(n9672) );
  OR2_X1 U9678 ( .A1(n9599), .A2(n9600), .ZN(n9670) );
  AND2_X1 U9679 ( .A1(n9673), .A2(n9674), .ZN(n9600) );
  NAND2_X1 U9680 ( .A1(n9458), .A2(n9675), .ZN(n9674) );
  OR2_X1 U9681 ( .A1(n9457), .A2(n9455), .ZN(n9675) );
  NOR2_X1 U9682 ( .A1(n9312), .A2(n7877), .ZN(n9458) );
  NAND2_X1 U9683 ( .A1(n9455), .A2(n9457), .ZN(n9673) );
  NAND2_X1 U9684 ( .A1(n9676), .A2(n9677), .ZN(n9457) );
  NAND3_X1 U9685 ( .A1(a_12_), .A2(n9678), .A3(b_22_), .ZN(n9677) );
  NAND2_X1 U9686 ( .A1(n9596), .A2(n9595), .ZN(n9678) );
  OR2_X1 U9687 ( .A1(n9595), .A2(n9596), .ZN(n9676) );
  AND2_X1 U9688 ( .A1(n9679), .A2(n9680), .ZN(n9596) );
  NAND2_X1 U9689 ( .A1(n9593), .A2(n9681), .ZN(n9680) );
  OR2_X1 U9690 ( .A1(n9592), .A2(n9590), .ZN(n9681) );
  NOR2_X1 U9691 ( .A1(n9312), .A2(n7355), .ZN(n9593) );
  NAND2_X1 U9692 ( .A1(n9590), .A2(n9592), .ZN(n9679) );
  NAND2_X1 U9693 ( .A1(n9682), .A2(n9683), .ZN(n9592) );
  NAND3_X1 U9694 ( .A1(a_14_), .A2(n9684), .A3(b_22_), .ZN(n9683) );
  NAND2_X1 U9695 ( .A1(n9588), .A2(n9587), .ZN(n9684) );
  OR2_X1 U9696 ( .A1(n9587), .A2(n9588), .ZN(n9682) );
  AND2_X1 U9697 ( .A1(n9685), .A2(n9686), .ZN(n9588) );
  NAND2_X1 U9698 ( .A1(n9475), .A2(n9687), .ZN(n9686) );
  OR2_X1 U9699 ( .A1(n9474), .A2(n9472), .ZN(n9687) );
  NOR2_X1 U9700 ( .A1(n9312), .A2(n7346), .ZN(n9475) );
  NAND2_X1 U9701 ( .A1(n9472), .A2(n9474), .ZN(n9685) );
  NAND2_X1 U9702 ( .A1(n9688), .A2(n9689), .ZN(n9474) );
  NAND3_X1 U9703 ( .A1(a_16_), .A2(n9690), .A3(b_22_), .ZN(n9689) );
  OR2_X1 U9704 ( .A1(n9584), .A2(n9582), .ZN(n9690) );
  NAND2_X1 U9705 ( .A1(n9582), .A2(n9584), .ZN(n9688) );
  NAND2_X1 U9706 ( .A1(n9691), .A2(n9692), .ZN(n9584) );
  NAND2_X1 U9707 ( .A1(n9581), .A2(n9693), .ZN(n9692) );
  OR2_X1 U9708 ( .A1(n9580), .A2(n9579), .ZN(n9693) );
  NOR2_X1 U9709 ( .A1(n9312), .A2(n7337), .ZN(n9581) );
  NAND2_X1 U9710 ( .A1(n9579), .A2(n9580), .ZN(n9691) );
  NAND2_X1 U9711 ( .A1(n9694), .A2(n9695), .ZN(n9580) );
  NAND3_X1 U9712 ( .A1(a_18_), .A2(n9696), .A3(b_22_), .ZN(n9695) );
  OR2_X1 U9713 ( .A1(n9576), .A2(n9575), .ZN(n9696) );
  NAND2_X1 U9714 ( .A1(n9575), .A2(n9576), .ZN(n9694) );
  NAND2_X1 U9715 ( .A1(n9697), .A2(n9698), .ZN(n9576) );
  NAND2_X1 U9716 ( .A1(n9573), .A2(n9699), .ZN(n9698) );
  OR2_X1 U9717 ( .A1(n9572), .A2(n9570), .ZN(n9699) );
  NOR2_X1 U9718 ( .A1(n9312), .A2(n7902), .ZN(n9573) );
  NAND2_X1 U9719 ( .A1(n9570), .A2(n9572), .ZN(n9697) );
  NAND2_X1 U9720 ( .A1(n9700), .A2(n9701), .ZN(n9572) );
  NAND3_X1 U9721 ( .A1(a_20_), .A2(n9702), .A3(b_22_), .ZN(n9701) );
  NAND2_X1 U9722 ( .A1(n9568), .A2(n9567), .ZN(n9702) );
  OR2_X1 U9723 ( .A1(n9567), .A2(n9568), .ZN(n9700) );
  AND2_X1 U9724 ( .A1(n9703), .A2(n9704), .ZN(n9568) );
  NAND2_X1 U9725 ( .A1(n9565), .A2(n9705), .ZN(n9704) );
  OR2_X1 U9726 ( .A1(n9564), .A2(n9563), .ZN(n9705) );
  NOR2_X1 U9727 ( .A1(n9312), .A2(n7909), .ZN(n9565) );
  NAND2_X1 U9728 ( .A1(n9563), .A2(n9564), .ZN(n9703) );
  NAND2_X1 U9729 ( .A1(n9706), .A2(n9707), .ZN(n9564) );
  NAND2_X1 U9730 ( .A1(n9561), .A2(n9708), .ZN(n9707) );
  NAND2_X1 U9731 ( .A1(n9560), .A2(n9559), .ZN(n9708) );
  OR2_X1 U9732 ( .A1(n9559), .A2(n9560), .ZN(n9706) );
  AND2_X1 U9733 ( .A1(n9709), .A2(n9710), .ZN(n9560) );
  NAND2_X1 U9734 ( .A1(n9557), .A2(n9711), .ZN(n9710) );
  OR2_X1 U9735 ( .A1(n9556), .A2(n9554), .ZN(n9711) );
  NOR2_X1 U9736 ( .A1(n9312), .A2(n7916), .ZN(n9557) );
  NAND2_X1 U9737 ( .A1(n9554), .A2(n9556), .ZN(n9709) );
  NAND2_X1 U9738 ( .A1(n9712), .A2(n9713), .ZN(n9556) );
  NAND3_X1 U9739 ( .A1(a_24_), .A2(n9714), .A3(b_22_), .ZN(n9713) );
  NAND2_X1 U9740 ( .A1(n9552), .A2(n9551), .ZN(n9714) );
  OR2_X1 U9741 ( .A1(n9551), .A2(n9552), .ZN(n9712) );
  AND2_X1 U9742 ( .A1(n9715), .A2(n9716), .ZN(n9552) );
  NAND2_X1 U9743 ( .A1(n9549), .A2(n9717), .ZN(n9716) );
  OR2_X1 U9744 ( .A1(n9548), .A2(n9547), .ZN(n9717) );
  NOR2_X1 U9745 ( .A1(n9312), .A2(n7923), .ZN(n9549) );
  NAND2_X1 U9746 ( .A1(n9547), .A2(n9548), .ZN(n9715) );
  NAND2_X1 U9747 ( .A1(n9544), .A2(n9718), .ZN(n9548) );
  NAND2_X1 U9748 ( .A1(n9543), .A2(n9545), .ZN(n9718) );
  NAND2_X1 U9749 ( .A1(n9719), .A2(n9720), .ZN(n9545) );
  NAND2_X1 U9750 ( .A1(b_22_), .A2(a_26_), .ZN(n9720) );
  INV_X1 U9751 ( .A(n9721), .ZN(n9719) );
  XNOR2_X1 U9752 ( .A(n9722), .B(n9723), .ZN(n9543) );
  NAND2_X1 U9753 ( .A1(n9724), .A2(n9725), .ZN(n9722) );
  NAND2_X1 U9754 ( .A1(a_26_), .A2(n9721), .ZN(n9544) );
  NAND2_X1 U9755 ( .A1(n9515), .A2(n9726), .ZN(n9721) );
  NAND2_X1 U9756 ( .A1(n9514), .A2(n9516), .ZN(n9726) );
  NAND2_X1 U9757 ( .A1(n9727), .A2(n9728), .ZN(n9516) );
  NAND2_X1 U9758 ( .A1(b_22_), .A2(a_27_), .ZN(n9728) );
  INV_X1 U9759 ( .A(n9729), .ZN(n9727) );
  XNOR2_X1 U9760 ( .A(n9730), .B(n9731), .ZN(n9514) );
  XOR2_X1 U9761 ( .A(n9732), .B(n9733), .Z(n9730) );
  NAND2_X1 U9762 ( .A1(b_21_), .A2(a_28_), .ZN(n9732) );
  NAND2_X1 U9763 ( .A1(a_27_), .A2(n9729), .ZN(n9515) );
  NAND2_X1 U9764 ( .A1(n9734), .A2(n9735), .ZN(n9729) );
  NAND3_X1 U9765 ( .A1(a_28_), .A2(n9736), .A3(b_22_), .ZN(n9735) );
  NAND2_X1 U9766 ( .A1(n9524), .A2(n9522), .ZN(n9736) );
  OR2_X1 U9767 ( .A1(n9522), .A2(n9524), .ZN(n9734) );
  AND2_X1 U9768 ( .A1(n9737), .A2(n9738), .ZN(n9524) );
  NAND2_X1 U9769 ( .A1(n9539), .A2(n9739), .ZN(n9738) );
  OR2_X1 U9770 ( .A1(n9540), .A2(n9541), .ZN(n9739) );
  NOR2_X1 U9771 ( .A1(n9312), .A2(n7946), .ZN(n9539) );
  NAND2_X1 U9772 ( .A1(n9541), .A2(n9540), .ZN(n9737) );
  NAND2_X1 U9773 ( .A1(n9740), .A2(n9741), .ZN(n9540) );
  NAND2_X1 U9774 ( .A1(b_20_), .A2(n9742), .ZN(n9741) );
  NAND2_X1 U9775 ( .A1(n7268), .A2(n9743), .ZN(n9742) );
  NAND2_X1 U9776 ( .A1(a_31_), .A2(n9537), .ZN(n9743) );
  NAND2_X1 U9777 ( .A1(b_21_), .A2(n9744), .ZN(n9740) );
  NAND2_X1 U9778 ( .A1(n7272), .A2(n9745), .ZN(n9744) );
  NAND2_X1 U9779 ( .A1(a_30_), .A2(n9746), .ZN(n9745) );
  AND3_X1 U9780 ( .A1(b_21_), .A2(n7954), .A3(b_22_), .ZN(n9541) );
  XNOR2_X1 U9781 ( .A(n9747), .B(n9748), .ZN(n9522) );
  XOR2_X1 U9782 ( .A(n9749), .B(n9750), .Z(n9747) );
  XNOR2_X1 U9783 ( .A(n9751), .B(n9752), .ZN(n9547) );
  NAND2_X1 U9784 ( .A1(n9753), .A2(n9754), .ZN(n9751) );
  XNOR2_X1 U9785 ( .A(n9755), .B(n9756), .ZN(n9551) );
  XOR2_X1 U9786 ( .A(n9757), .B(n9758), .Z(n9755) );
  XNOR2_X1 U9787 ( .A(n9759), .B(n9760), .ZN(n9554) );
  XNOR2_X1 U9788 ( .A(n9761), .B(n9762), .ZN(n9759) );
  NOR2_X1 U9789 ( .A1(n7691), .A2(n9537), .ZN(n9762) );
  XOR2_X1 U9790 ( .A(n9763), .B(n9764), .Z(n9559) );
  XNOR2_X1 U9791 ( .A(n9765), .B(n9766), .ZN(n9764) );
  XNOR2_X1 U9792 ( .A(n9767), .B(n9768), .ZN(n9563) );
  XOR2_X1 U9793 ( .A(n9769), .B(n9770), .Z(n9768) );
  NAND2_X1 U9794 ( .A1(b_21_), .A2(a_22_), .ZN(n9770) );
  XNOR2_X1 U9795 ( .A(n9771), .B(n9772), .ZN(n9567) );
  XOR2_X1 U9796 ( .A(n9773), .B(n9774), .Z(n9771) );
  XNOR2_X1 U9797 ( .A(n9775), .B(n9776), .ZN(n9570) );
  XNOR2_X1 U9798 ( .A(n9777), .B(n9778), .ZN(n9775) );
  NOR2_X1 U9799 ( .A1(n7987), .A2(n9537), .ZN(n9778) );
  XNOR2_X1 U9800 ( .A(n9779), .B(n9780), .ZN(n9575) );
  XNOR2_X1 U9801 ( .A(n9781), .B(n9782), .ZN(n9780) );
  XNOR2_X1 U9802 ( .A(n9783), .B(n9784), .ZN(n9579) );
  XNOR2_X1 U9803 ( .A(n9785), .B(n9786), .ZN(n9783) );
  NOR2_X1 U9804 ( .A1(n7764), .A2(n9537), .ZN(n9786) );
  XNOR2_X1 U9805 ( .A(n9787), .B(n9788), .ZN(n9582) );
  XNOR2_X1 U9806 ( .A(n9789), .B(n9790), .ZN(n9788) );
  XNOR2_X1 U9807 ( .A(n9791), .B(n9792), .ZN(n9472) );
  XNOR2_X1 U9808 ( .A(n9793), .B(n9794), .ZN(n9791) );
  NOR2_X1 U9809 ( .A1(n7773), .A2(n9537), .ZN(n9794) );
  XNOR2_X1 U9810 ( .A(n9795), .B(n9796), .ZN(n9587) );
  XOR2_X1 U9811 ( .A(n9797), .B(n9798), .Z(n9795) );
  XNOR2_X1 U9812 ( .A(n9799), .B(n9800), .ZN(n9590) );
  XNOR2_X1 U9813 ( .A(n9801), .B(n9802), .ZN(n9799) );
  NOR2_X1 U9814 ( .A1(n7782), .A2(n9537), .ZN(n9802) );
  XNOR2_X1 U9815 ( .A(n9803), .B(n9804), .ZN(n9595) );
  XOR2_X1 U9816 ( .A(n9805), .B(n9806), .Z(n9803) );
  XNOR2_X1 U9817 ( .A(n9807), .B(n9808), .ZN(n9455) );
  XOR2_X1 U9818 ( .A(n9809), .B(n9810), .Z(n9808) );
  NAND2_X1 U9819 ( .A1(b_21_), .A2(a_12_), .ZN(n9810) );
  XOR2_X1 U9820 ( .A(n9811), .B(n9812), .Z(n9599) );
  XNOR2_X1 U9821 ( .A(n9813), .B(n9814), .ZN(n9812) );
  XNOR2_X1 U9822 ( .A(n9815), .B(n9816), .ZN(n9603) );
  XOR2_X1 U9823 ( .A(n9817), .B(n9818), .Z(n9815) );
  XNOR2_X1 U9824 ( .A(n9819), .B(n9820), .ZN(n9606) );
  XNOR2_X1 U9825 ( .A(n9821), .B(n9822), .ZN(n9819) );
  NOR2_X1 U9826 ( .A1(n7870), .A2(n9537), .ZN(n9822) );
  XNOR2_X1 U9827 ( .A(n9823), .B(n9824), .ZN(n9438) );
  XOR2_X1 U9828 ( .A(n9825), .B(n9826), .Z(n9824) );
  NAND2_X1 U9829 ( .A1(b_21_), .A2(a_8_), .ZN(n9826) );
  XOR2_X1 U9830 ( .A(n9827), .B(n9828), .Z(n9611) );
  XOR2_X1 U9831 ( .A(n9829), .B(n9830), .Z(n9828) );
  NAND2_X1 U9832 ( .A1(b_21_), .A2(a_7_), .ZN(n9830) );
  XNOR2_X1 U9833 ( .A(n9831), .B(n9832), .ZN(n9615) );
  XOR2_X1 U9834 ( .A(n9833), .B(n9834), .Z(n9832) );
  NAND2_X1 U9835 ( .A1(b_21_), .A2(a_6_), .ZN(n9834) );
  XNOR2_X1 U9836 ( .A(n9835), .B(n9836), .ZN(n9618) );
  XNOR2_X1 U9837 ( .A(n9837), .B(n9838), .ZN(n9835) );
  NOR2_X1 U9838 ( .A1(n7393), .A2(n9537), .ZN(n9838) );
  XNOR2_X1 U9839 ( .A(n9839), .B(n9840), .ZN(n9623) );
  XOR2_X1 U9840 ( .A(n9841), .B(n9842), .Z(n9840) );
  NAND2_X1 U9841 ( .A1(b_21_), .A2(a_4_), .ZN(n9842) );
  XNOR2_X1 U9842 ( .A(n9843), .B(n9844), .ZN(n9627) );
  XOR2_X1 U9843 ( .A(n9845), .B(n9846), .Z(n9844) );
  NAND2_X1 U9844 ( .A1(b_21_), .A2(a_3_), .ZN(n9846) );
  XNOR2_X1 U9845 ( .A(n9847), .B(n9848), .ZN(n9631) );
  XOR2_X1 U9846 ( .A(n9849), .B(n9850), .Z(n9848) );
  NAND2_X1 U9847 ( .A1(b_21_), .A2(a_2_), .ZN(n9850) );
  NAND2_X1 U9848 ( .A1(n9851), .A2(n9852), .ZN(n7570) );
  XNOR2_X1 U9849 ( .A(n9853), .B(n9854), .ZN(n7571) );
  XNOR2_X1 U9850 ( .A(n9855), .B(n9856), .ZN(n9854) );
  NAND2_X1 U9851 ( .A1(n9857), .A2(n9634), .ZN(n7463) );
  NOR2_X1 U9852 ( .A1(n9852), .A2(n9851), .ZN(n9634) );
  AND2_X1 U9853 ( .A1(n9858), .A2(n9859), .ZN(n9851) );
  NAND2_X1 U9854 ( .A1(n9856), .A2(n9860), .ZN(n9859) );
  OR2_X1 U9855 ( .A1(n9855), .A2(n9853), .ZN(n9860) );
  NOR2_X1 U9856 ( .A1(n9537), .A2(n7613), .ZN(n9856) );
  NAND2_X1 U9857 ( .A1(n9853), .A2(n9855), .ZN(n9858) );
  NAND2_X1 U9858 ( .A1(n9861), .A2(n9862), .ZN(n9855) );
  NAND3_X1 U9859 ( .A1(a_1_), .A2(n9863), .A3(b_21_), .ZN(n9862) );
  OR2_X1 U9860 ( .A1(n9641), .A2(n9640), .ZN(n9863) );
  NAND2_X1 U9861 ( .A1(n9640), .A2(n9641), .ZN(n9861) );
  NAND2_X1 U9862 ( .A1(n9864), .A2(n9865), .ZN(n9641) );
  NAND3_X1 U9863 ( .A1(a_2_), .A2(n9866), .A3(b_21_), .ZN(n9865) );
  OR2_X1 U9864 ( .A1(n9849), .A2(n9847), .ZN(n9866) );
  NAND2_X1 U9865 ( .A1(n9847), .A2(n9849), .ZN(n9864) );
  NAND2_X1 U9866 ( .A1(n9867), .A2(n9868), .ZN(n9849) );
  NAND3_X1 U9867 ( .A1(a_3_), .A2(n9869), .A3(b_21_), .ZN(n9868) );
  OR2_X1 U9868 ( .A1(n9845), .A2(n9843), .ZN(n9869) );
  NAND2_X1 U9869 ( .A1(n9843), .A2(n9845), .ZN(n9867) );
  NAND2_X1 U9870 ( .A1(n9870), .A2(n9871), .ZN(n9845) );
  NAND3_X1 U9871 ( .A1(a_4_), .A2(n9872), .A3(b_21_), .ZN(n9871) );
  OR2_X1 U9872 ( .A1(n9841), .A2(n9839), .ZN(n9872) );
  NAND2_X1 U9873 ( .A1(n9839), .A2(n9841), .ZN(n9870) );
  NAND2_X1 U9874 ( .A1(n9873), .A2(n9874), .ZN(n9841) );
  NAND3_X1 U9875 ( .A1(a_5_), .A2(n9875), .A3(b_21_), .ZN(n9874) );
  NAND2_X1 U9876 ( .A1(n9837), .A2(n9836), .ZN(n9875) );
  OR2_X1 U9877 ( .A1(n9836), .A2(n9837), .ZN(n9873) );
  AND2_X1 U9878 ( .A1(n9876), .A2(n9877), .ZN(n9837) );
  NAND3_X1 U9879 ( .A1(a_6_), .A2(n9878), .A3(b_21_), .ZN(n9877) );
  OR2_X1 U9880 ( .A1(n9833), .A2(n9831), .ZN(n9878) );
  NAND2_X1 U9881 ( .A1(n9831), .A2(n9833), .ZN(n9876) );
  NAND2_X1 U9882 ( .A1(n9879), .A2(n9880), .ZN(n9833) );
  NAND3_X1 U9883 ( .A1(a_7_), .A2(n9881), .A3(b_21_), .ZN(n9880) );
  OR2_X1 U9884 ( .A1(n9829), .A2(n9827), .ZN(n9881) );
  NAND2_X1 U9885 ( .A1(n9827), .A2(n9829), .ZN(n9879) );
  NAND2_X1 U9886 ( .A1(n9882), .A2(n9883), .ZN(n9829) );
  NAND3_X1 U9887 ( .A1(a_8_), .A2(n9884), .A3(b_21_), .ZN(n9883) );
  OR2_X1 U9888 ( .A1(n9825), .A2(n9823), .ZN(n9884) );
  NAND2_X1 U9889 ( .A1(n9823), .A2(n9825), .ZN(n9882) );
  NAND2_X1 U9890 ( .A1(n9885), .A2(n9886), .ZN(n9825) );
  NAND3_X1 U9891 ( .A1(a_9_), .A2(n9887), .A3(b_21_), .ZN(n9886) );
  NAND2_X1 U9892 ( .A1(n9821), .A2(n9820), .ZN(n9887) );
  OR2_X1 U9893 ( .A1(n9820), .A2(n9821), .ZN(n9885) );
  AND2_X1 U9894 ( .A1(n9888), .A2(n9889), .ZN(n9821) );
  NAND2_X1 U9895 ( .A1(n9818), .A2(n9890), .ZN(n9889) );
  OR2_X1 U9896 ( .A1(n9817), .A2(n9816), .ZN(n9890) );
  NOR2_X1 U9897 ( .A1(n9537), .A2(n7799), .ZN(n9818) );
  NAND2_X1 U9898 ( .A1(n9816), .A2(n9817), .ZN(n9888) );
  NAND2_X1 U9899 ( .A1(n9891), .A2(n9892), .ZN(n9817) );
  NAND2_X1 U9900 ( .A1(n9814), .A2(n9893), .ZN(n9892) );
  OR2_X1 U9901 ( .A1(n9813), .A2(n9811), .ZN(n9893) );
  NOR2_X1 U9902 ( .A1(n9537), .A2(n7877), .ZN(n9814) );
  NAND2_X1 U9903 ( .A1(n9811), .A2(n9813), .ZN(n9891) );
  NAND2_X1 U9904 ( .A1(n9894), .A2(n9895), .ZN(n9813) );
  NAND3_X1 U9905 ( .A1(a_12_), .A2(n9896), .A3(b_21_), .ZN(n9895) );
  OR2_X1 U9906 ( .A1(n9809), .A2(n9807), .ZN(n9896) );
  NAND2_X1 U9907 ( .A1(n9807), .A2(n9809), .ZN(n9894) );
  NAND2_X1 U9908 ( .A1(n9897), .A2(n9898), .ZN(n9809) );
  NAND2_X1 U9909 ( .A1(n9806), .A2(n9899), .ZN(n9898) );
  OR2_X1 U9910 ( .A1(n9805), .A2(n9804), .ZN(n9899) );
  NOR2_X1 U9911 ( .A1(n9537), .A2(n7355), .ZN(n9806) );
  NAND2_X1 U9912 ( .A1(n9804), .A2(n9805), .ZN(n9897) );
  NAND2_X1 U9913 ( .A1(n9900), .A2(n9901), .ZN(n9805) );
  NAND3_X1 U9914 ( .A1(a_14_), .A2(n9902), .A3(b_21_), .ZN(n9901) );
  NAND2_X1 U9915 ( .A1(n9801), .A2(n9800), .ZN(n9902) );
  OR2_X1 U9916 ( .A1(n9800), .A2(n9801), .ZN(n9900) );
  AND2_X1 U9917 ( .A1(n9903), .A2(n9904), .ZN(n9801) );
  NAND2_X1 U9918 ( .A1(n9798), .A2(n9905), .ZN(n9904) );
  OR2_X1 U9919 ( .A1(n9797), .A2(n9796), .ZN(n9905) );
  NOR2_X1 U9920 ( .A1(n9537), .A2(n7346), .ZN(n9798) );
  NAND2_X1 U9921 ( .A1(n9796), .A2(n9797), .ZN(n9903) );
  NAND2_X1 U9922 ( .A1(n9906), .A2(n9907), .ZN(n9797) );
  NAND3_X1 U9923 ( .A1(a_16_), .A2(n9908), .A3(b_21_), .ZN(n9907) );
  NAND2_X1 U9924 ( .A1(n9793), .A2(n9792), .ZN(n9908) );
  OR2_X1 U9925 ( .A1(n9792), .A2(n9793), .ZN(n9906) );
  AND2_X1 U9926 ( .A1(n9909), .A2(n9910), .ZN(n9793) );
  NAND2_X1 U9927 ( .A1(n9790), .A2(n9911), .ZN(n9910) );
  OR2_X1 U9928 ( .A1(n9789), .A2(n9787), .ZN(n9911) );
  NOR2_X1 U9929 ( .A1(n9537), .A2(n7337), .ZN(n9790) );
  NAND2_X1 U9930 ( .A1(n9787), .A2(n9789), .ZN(n9909) );
  NAND2_X1 U9931 ( .A1(n9912), .A2(n9913), .ZN(n9789) );
  NAND3_X1 U9932 ( .A1(a_18_), .A2(n9914), .A3(b_21_), .ZN(n9913) );
  NAND2_X1 U9933 ( .A1(n9785), .A2(n9784), .ZN(n9914) );
  OR2_X1 U9934 ( .A1(n9784), .A2(n9785), .ZN(n9912) );
  AND2_X1 U9935 ( .A1(n9915), .A2(n9916), .ZN(n9785) );
  NAND2_X1 U9936 ( .A1(n9782), .A2(n9917), .ZN(n9916) );
  OR2_X1 U9937 ( .A1(n9781), .A2(n9779), .ZN(n9917) );
  NOR2_X1 U9938 ( .A1(n9537), .A2(n7902), .ZN(n9782) );
  NAND2_X1 U9939 ( .A1(n9779), .A2(n9781), .ZN(n9915) );
  NAND2_X1 U9940 ( .A1(n9918), .A2(n9919), .ZN(n9781) );
  NAND3_X1 U9941 ( .A1(a_20_), .A2(n9920), .A3(b_21_), .ZN(n9919) );
  NAND2_X1 U9942 ( .A1(n9777), .A2(n9776), .ZN(n9920) );
  OR2_X1 U9943 ( .A1(n9776), .A2(n9777), .ZN(n9918) );
  AND2_X1 U9944 ( .A1(n9921), .A2(n9922), .ZN(n9777) );
  NAND2_X1 U9945 ( .A1(n9774), .A2(n9923), .ZN(n9922) );
  OR2_X1 U9946 ( .A1(n9773), .A2(n9772), .ZN(n9923) );
  NAND2_X1 U9947 ( .A1(n9772), .A2(n9773), .ZN(n9921) );
  NAND2_X1 U9948 ( .A1(n9924), .A2(n9925), .ZN(n9773) );
  NAND3_X1 U9949 ( .A1(a_22_), .A2(n9926), .A3(b_21_), .ZN(n9925) );
  OR2_X1 U9950 ( .A1(n9769), .A2(n9767), .ZN(n9926) );
  NAND2_X1 U9951 ( .A1(n9767), .A2(n9769), .ZN(n9924) );
  NAND2_X1 U9952 ( .A1(n9927), .A2(n9928), .ZN(n9769) );
  NAND2_X1 U9953 ( .A1(n9766), .A2(n9929), .ZN(n9928) );
  OR2_X1 U9954 ( .A1(n9765), .A2(n9763), .ZN(n9929) );
  NOR2_X1 U9955 ( .A1(n9537), .A2(n7916), .ZN(n9766) );
  NAND2_X1 U9956 ( .A1(n9763), .A2(n9765), .ZN(n9927) );
  NAND2_X1 U9957 ( .A1(n9930), .A2(n9931), .ZN(n9765) );
  NAND3_X1 U9958 ( .A1(a_24_), .A2(n9932), .A3(b_21_), .ZN(n9931) );
  NAND2_X1 U9959 ( .A1(n9761), .A2(n9760), .ZN(n9932) );
  OR2_X1 U9960 ( .A1(n9760), .A2(n9761), .ZN(n9930) );
  AND2_X1 U9961 ( .A1(n9933), .A2(n9934), .ZN(n9761) );
  NAND2_X1 U9962 ( .A1(n9758), .A2(n9935), .ZN(n9934) );
  OR2_X1 U9963 ( .A1(n9757), .A2(n9756), .ZN(n9935) );
  NOR2_X1 U9964 ( .A1(n9537), .A2(n7923), .ZN(n9758) );
  NAND2_X1 U9965 ( .A1(n9756), .A2(n9757), .ZN(n9933) );
  NAND2_X1 U9966 ( .A1(n9753), .A2(n9936), .ZN(n9757) );
  NAND2_X1 U9967 ( .A1(n9752), .A2(n9754), .ZN(n9936) );
  NAND2_X1 U9968 ( .A1(n9937), .A2(n9938), .ZN(n9754) );
  NAND2_X1 U9969 ( .A1(b_21_), .A2(a_26_), .ZN(n9938) );
  INV_X1 U9970 ( .A(n9939), .ZN(n9937) );
  XNOR2_X1 U9971 ( .A(n9940), .B(n9941), .ZN(n9752) );
  NAND2_X1 U9972 ( .A1(n9942), .A2(n9943), .ZN(n9940) );
  NAND2_X1 U9973 ( .A1(a_26_), .A2(n9939), .ZN(n9753) );
  NAND2_X1 U9974 ( .A1(n9724), .A2(n9944), .ZN(n9939) );
  NAND2_X1 U9975 ( .A1(n9723), .A2(n9725), .ZN(n9944) );
  NAND2_X1 U9976 ( .A1(n9945), .A2(n9946), .ZN(n9725) );
  NAND2_X1 U9977 ( .A1(b_21_), .A2(a_27_), .ZN(n9946) );
  INV_X1 U9978 ( .A(n9947), .ZN(n9945) );
  XNOR2_X1 U9979 ( .A(n9948), .B(n9949), .ZN(n9723) );
  XOR2_X1 U9980 ( .A(n9950), .B(n9951), .Z(n9948) );
  NAND2_X1 U9981 ( .A1(b_20_), .A2(a_28_), .ZN(n9950) );
  NAND2_X1 U9982 ( .A1(a_27_), .A2(n9947), .ZN(n9724) );
  NAND2_X1 U9983 ( .A1(n9952), .A2(n9953), .ZN(n9947) );
  NAND3_X1 U9984 ( .A1(a_28_), .A2(n9954), .A3(b_21_), .ZN(n9953) );
  NAND2_X1 U9985 ( .A1(n9733), .A2(n9731), .ZN(n9954) );
  OR2_X1 U9986 ( .A1(n9731), .A2(n9733), .ZN(n9952) );
  AND2_X1 U9987 ( .A1(n9955), .A2(n9956), .ZN(n9733) );
  NAND2_X1 U9988 ( .A1(n9748), .A2(n9957), .ZN(n9956) );
  OR2_X1 U9989 ( .A1(n9749), .A2(n9750), .ZN(n9957) );
  NOR2_X1 U9990 ( .A1(n9537), .A2(n7946), .ZN(n9748) );
  NAND2_X1 U9991 ( .A1(n9750), .A2(n9749), .ZN(n9955) );
  NAND2_X1 U9992 ( .A1(n9958), .A2(n9959), .ZN(n9749) );
  NAND2_X1 U9993 ( .A1(b_19_), .A2(n9960), .ZN(n9959) );
  NAND2_X1 U9994 ( .A1(n7268), .A2(n9961), .ZN(n9960) );
  NAND2_X1 U9995 ( .A1(a_31_), .A2(n9746), .ZN(n9961) );
  NAND2_X1 U9996 ( .A1(b_20_), .A2(n9962), .ZN(n9958) );
  NAND2_X1 U9997 ( .A1(n7272), .A2(n9963), .ZN(n9962) );
  NAND2_X1 U9998 ( .A1(a_30_), .A2(n9964), .ZN(n9963) );
  AND3_X1 U9999 ( .A1(b_20_), .A2(n7954), .A3(b_21_), .ZN(n9750) );
  XNOR2_X1 U10000 ( .A(n9965), .B(n9966), .ZN(n9731) );
  XOR2_X1 U10001 ( .A(n9967), .B(n9968), .Z(n9965) );
  XNOR2_X1 U10002 ( .A(n9969), .B(n9970), .ZN(n9756) );
  NAND2_X1 U10003 ( .A1(n9971), .A2(n9972), .ZN(n9969) );
  XNOR2_X1 U10004 ( .A(n9973), .B(n9974), .ZN(n9760) );
  XOR2_X1 U10005 ( .A(n9975), .B(n9976), .Z(n9973) );
  XNOR2_X1 U10006 ( .A(n9977), .B(n9978), .ZN(n9763) );
  XNOR2_X1 U10007 ( .A(n9979), .B(n9980), .ZN(n9977) );
  NOR2_X1 U10008 ( .A1(n7691), .A2(n9746), .ZN(n9980) );
  XNOR2_X1 U10009 ( .A(n9981), .B(n9982), .ZN(n9767) );
  XNOR2_X1 U10010 ( .A(n9983), .B(n9984), .ZN(n9982) );
  XNOR2_X1 U10011 ( .A(n9985), .B(n9986), .ZN(n9772) );
  XOR2_X1 U10012 ( .A(n9987), .B(n9988), .Z(n9986) );
  NAND2_X1 U10013 ( .A1(b_20_), .A2(a_22_), .ZN(n9988) );
  XNOR2_X1 U10014 ( .A(n9989), .B(n9990), .ZN(n9776) );
  XOR2_X1 U10015 ( .A(n9991), .B(n9992), .Z(n9989) );
  XOR2_X1 U10016 ( .A(n9993), .B(n9994), .Z(n9779) );
  XOR2_X1 U10017 ( .A(n9995), .B(n9996), .Z(n9993) );
  XOR2_X1 U10018 ( .A(n9997), .B(n9998), .Z(n9784) );
  XNOR2_X1 U10019 ( .A(n9999), .B(n10000), .ZN(n9998) );
  XNOR2_X1 U10020 ( .A(n10001), .B(n10002), .ZN(n9787) );
  XNOR2_X1 U10021 ( .A(n10003), .B(n10004), .ZN(n10001) );
  NOR2_X1 U10022 ( .A1(n7764), .A2(n9746), .ZN(n10004) );
  XOR2_X1 U10023 ( .A(n10005), .B(n10006), .Z(n9792) );
  XNOR2_X1 U10024 ( .A(n10007), .B(n10008), .ZN(n10006) );
  XNOR2_X1 U10025 ( .A(n10009), .B(n10010), .ZN(n9796) );
  XNOR2_X1 U10026 ( .A(n10011), .B(n10012), .ZN(n10009) );
  NOR2_X1 U10027 ( .A1(n7773), .A2(n9746), .ZN(n10012) );
  XOR2_X1 U10028 ( .A(n10013), .B(n10014), .Z(n9800) );
  XNOR2_X1 U10029 ( .A(n10015), .B(n10016), .ZN(n10014) );
  XNOR2_X1 U10030 ( .A(n10017), .B(n10018), .ZN(n9804) );
  XNOR2_X1 U10031 ( .A(n10019), .B(n10020), .ZN(n10017) );
  NOR2_X1 U10032 ( .A1(n7782), .A2(n9746), .ZN(n10020) );
  XOR2_X1 U10033 ( .A(n10021), .B(n10022), .Z(n9807) );
  XOR2_X1 U10034 ( .A(n10023), .B(n10024), .Z(n10021) );
  XNOR2_X1 U10035 ( .A(n10025), .B(n10026), .ZN(n9811) );
  XNOR2_X1 U10036 ( .A(n10027), .B(n10028), .ZN(n10025) );
  NOR2_X1 U10037 ( .A1(n8020), .A2(n9746), .ZN(n10028) );
  XNOR2_X1 U10038 ( .A(n10029), .B(n10030), .ZN(n9816) );
  XOR2_X1 U10039 ( .A(n10031), .B(n10032), .Z(n10030) );
  NAND2_X1 U10040 ( .A1(b_20_), .A2(a_11_), .ZN(n10032) );
  XNOR2_X1 U10041 ( .A(n10033), .B(n10034), .ZN(n9820) );
  XOR2_X1 U10042 ( .A(n10035), .B(n10036), .Z(n10033) );
  XOR2_X1 U10043 ( .A(n10037), .B(n10038), .Z(n9823) );
  XOR2_X1 U10044 ( .A(n10039), .B(n10040), .Z(n10037) );
  XNOR2_X1 U10045 ( .A(n10041), .B(n10042), .ZN(n9827) );
  XNOR2_X1 U10046 ( .A(n10043), .B(n10044), .ZN(n10041) );
  NOR2_X1 U10047 ( .A1(n8037), .A2(n9746), .ZN(n10044) );
  XNOR2_X1 U10048 ( .A(n10045), .B(n10046), .ZN(n9831) );
  NAND2_X1 U10049 ( .A1(n10047), .A2(n10048), .ZN(n10045) );
  XNOR2_X1 U10050 ( .A(n10049), .B(n10050), .ZN(n9836) );
  NOR2_X1 U10051 ( .A1(n10051), .A2(n10052), .ZN(n10050) );
  NOR2_X1 U10052 ( .A1(n10053), .A2(n10054), .ZN(n10051) );
  NOR2_X1 U10053 ( .A1(n7388), .A2(n9746), .ZN(n10053) );
  XOR2_X1 U10054 ( .A(n10055), .B(n10056), .Z(n9839) );
  XOR2_X1 U10055 ( .A(n10057), .B(n10058), .Z(n10055) );
  XOR2_X1 U10056 ( .A(n10059), .B(n10060), .Z(n9843) );
  XOR2_X1 U10057 ( .A(n10061), .B(n10062), .Z(n10059) );
  NOR2_X1 U10058 ( .A1(n7398), .A2(n9746), .ZN(n10062) );
  XNOR2_X1 U10059 ( .A(n10063), .B(n10064), .ZN(n9847) );
  NAND2_X1 U10060 ( .A1(n10065), .A2(n10066), .ZN(n10063) );
  XNOR2_X1 U10061 ( .A(n10067), .B(n10068), .ZN(n9640) );
  NAND2_X1 U10062 ( .A1(n10069), .A2(n10070), .ZN(n10067) );
  XNOR2_X1 U10063 ( .A(n10071), .B(n10072), .ZN(n9853) );
  XNOR2_X1 U10064 ( .A(n10073), .B(n10074), .ZN(n10071) );
  XNOR2_X1 U10065 ( .A(n10075), .B(n10076), .ZN(n9852) );
  XOR2_X1 U10066 ( .A(n10077), .B(n10078), .Z(n10075) );
  NOR2_X1 U10067 ( .A1(n7613), .A2(n9746), .ZN(n10078) );
  XOR2_X1 U10068 ( .A(n7562), .B(n7561), .Z(n9857) );
  NAND3_X1 U10069 ( .A1(n7561), .A2(n7562), .A3(n10079), .ZN(n7472) );
  XOR2_X1 U10070 ( .A(n7555), .B(n7554), .Z(n10079) );
  NAND2_X1 U10071 ( .A1(n10080), .A2(n10081), .ZN(n7562) );
  NAND3_X1 U10072 ( .A1(a_0_), .A2(n10082), .A3(b_20_), .ZN(n10081) );
  OR2_X1 U10073 ( .A1(n10077), .A2(n10076), .ZN(n10082) );
  NAND2_X1 U10074 ( .A1(n10076), .A2(n10077), .ZN(n10080) );
  NAND2_X1 U10075 ( .A1(n10083), .A2(n10084), .ZN(n10077) );
  NAND2_X1 U10076 ( .A1(n10074), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U10077 ( .A1(n10073), .A2(n10072), .ZN(n10085) );
  NOR2_X1 U10078 ( .A1(n9746), .A2(n7411), .ZN(n10074) );
  OR2_X1 U10079 ( .A1(n10072), .A2(n10073), .ZN(n10083) );
  AND2_X1 U10080 ( .A1(n10069), .A2(n10086), .ZN(n10073) );
  NAND2_X1 U10081 ( .A1(n10068), .A2(n10070), .ZN(n10086) );
  NAND2_X1 U10082 ( .A1(n10087), .A2(n10088), .ZN(n10070) );
  NAND2_X1 U10083 ( .A1(b_20_), .A2(a_2_), .ZN(n10088) );
  INV_X1 U10084 ( .A(n10089), .ZN(n10087) );
  XNOR2_X1 U10085 ( .A(n10090), .B(n10091), .ZN(n10068) );
  XOR2_X1 U10086 ( .A(n10092), .B(n10093), .Z(n10091) );
  NAND2_X1 U10087 ( .A1(b_19_), .A2(a_3_), .ZN(n10093) );
  NAND2_X1 U10088 ( .A1(a_2_), .A2(n10089), .ZN(n10069) );
  NAND2_X1 U10089 ( .A1(n10065), .A2(n10094), .ZN(n10089) );
  NAND2_X1 U10090 ( .A1(n10064), .A2(n10066), .ZN(n10094) );
  NAND2_X1 U10091 ( .A1(n10095), .A2(n10096), .ZN(n10066) );
  NAND2_X1 U10092 ( .A1(b_20_), .A2(a_3_), .ZN(n10096) );
  INV_X1 U10093 ( .A(n10097), .ZN(n10095) );
  XOR2_X1 U10094 ( .A(n10098), .B(n10099), .Z(n10064) );
  XOR2_X1 U10095 ( .A(n10100), .B(n10101), .Z(n10098) );
  NOR2_X1 U10096 ( .A1(n7398), .A2(n9964), .ZN(n10101) );
  NAND2_X1 U10097 ( .A1(a_3_), .A2(n10097), .ZN(n10065) );
  NAND2_X1 U10098 ( .A1(n10102), .A2(n10103), .ZN(n10097) );
  NAND3_X1 U10099 ( .A1(a_4_), .A2(n10104), .A3(b_20_), .ZN(n10103) );
  OR2_X1 U10100 ( .A1(n10061), .A2(n10060), .ZN(n10104) );
  NAND2_X1 U10101 ( .A1(n10060), .A2(n10061), .ZN(n10102) );
  NAND2_X1 U10102 ( .A1(n10105), .A2(n10106), .ZN(n10061) );
  NAND2_X1 U10103 ( .A1(n10058), .A2(n10107), .ZN(n10106) );
  OR2_X1 U10104 ( .A1(n10057), .A2(n10056), .ZN(n10107) );
  NOR2_X1 U10105 ( .A1(n9746), .A2(n7393), .ZN(n10058) );
  NAND2_X1 U10106 ( .A1(n10056), .A2(n10057), .ZN(n10105) );
  OR2_X1 U10107 ( .A1(n10052), .A2(n10108), .ZN(n10057) );
  AND2_X1 U10108 ( .A1(n10049), .A2(n10109), .ZN(n10108) );
  NAND2_X1 U10109 ( .A1(n10110), .A2(n10111), .ZN(n10109) );
  NAND2_X1 U10110 ( .A1(b_20_), .A2(a_6_), .ZN(n10111) );
  XNOR2_X1 U10111 ( .A(n10112), .B(n10113), .ZN(n10049) );
  XOR2_X1 U10112 ( .A(n10114), .B(n10115), .Z(n10113) );
  NAND2_X1 U10113 ( .A1(b_19_), .A2(a_7_), .ZN(n10115) );
  NOR2_X1 U10114 ( .A1(n7388), .A2(n10110), .ZN(n10052) );
  INV_X1 U10115 ( .A(n10054), .ZN(n10110) );
  NAND2_X1 U10116 ( .A1(n10047), .A2(n10116), .ZN(n10054) );
  NAND2_X1 U10117 ( .A1(n10046), .A2(n10048), .ZN(n10116) );
  NAND2_X1 U10118 ( .A1(n10117), .A2(n10118), .ZN(n10048) );
  NAND2_X1 U10119 ( .A1(b_20_), .A2(a_7_), .ZN(n10118) );
  INV_X1 U10120 ( .A(n10119), .ZN(n10117) );
  XNOR2_X1 U10121 ( .A(n10120), .B(n10121), .ZN(n10046) );
  XOR2_X1 U10122 ( .A(n10122), .B(n10123), .Z(n10121) );
  NAND2_X1 U10123 ( .A1(b_19_), .A2(a_8_), .ZN(n10123) );
  NAND2_X1 U10124 ( .A1(a_7_), .A2(n10119), .ZN(n10047) );
  NAND2_X1 U10125 ( .A1(n10124), .A2(n10125), .ZN(n10119) );
  NAND3_X1 U10126 ( .A1(a_8_), .A2(n10126), .A3(b_20_), .ZN(n10125) );
  NAND2_X1 U10127 ( .A1(n10043), .A2(n10042), .ZN(n10126) );
  OR2_X1 U10128 ( .A1(n10042), .A2(n10043), .ZN(n10124) );
  AND2_X1 U10129 ( .A1(n10127), .A2(n10128), .ZN(n10043) );
  NAND2_X1 U10130 ( .A1(n10040), .A2(n10129), .ZN(n10128) );
  OR2_X1 U10131 ( .A1(n10039), .A2(n10038), .ZN(n10129) );
  NOR2_X1 U10132 ( .A1(n9746), .A2(n7870), .ZN(n10040) );
  NAND2_X1 U10133 ( .A1(n10038), .A2(n10039), .ZN(n10127) );
  NAND2_X1 U10134 ( .A1(n10130), .A2(n10131), .ZN(n10039) );
  NAND2_X1 U10135 ( .A1(n10036), .A2(n10132), .ZN(n10131) );
  OR2_X1 U10136 ( .A1(n10035), .A2(n10034), .ZN(n10132) );
  NOR2_X1 U10137 ( .A1(n9746), .A2(n7799), .ZN(n10036) );
  NAND2_X1 U10138 ( .A1(n10034), .A2(n10035), .ZN(n10130) );
  NAND2_X1 U10139 ( .A1(n10133), .A2(n10134), .ZN(n10035) );
  NAND3_X1 U10140 ( .A1(a_11_), .A2(n10135), .A3(b_20_), .ZN(n10134) );
  OR2_X1 U10141 ( .A1(n10031), .A2(n10029), .ZN(n10135) );
  NAND2_X1 U10142 ( .A1(n10029), .A2(n10031), .ZN(n10133) );
  NAND2_X1 U10143 ( .A1(n10136), .A2(n10137), .ZN(n10031) );
  NAND3_X1 U10144 ( .A1(a_12_), .A2(n10138), .A3(b_20_), .ZN(n10137) );
  NAND2_X1 U10145 ( .A1(n10027), .A2(n10026), .ZN(n10138) );
  OR2_X1 U10146 ( .A1(n10026), .A2(n10027), .ZN(n10136) );
  AND2_X1 U10147 ( .A1(n10139), .A2(n10140), .ZN(n10027) );
  NAND2_X1 U10148 ( .A1(n10024), .A2(n10141), .ZN(n10140) );
  OR2_X1 U10149 ( .A1(n10023), .A2(n10022), .ZN(n10141) );
  NOR2_X1 U10150 ( .A1(n9746), .A2(n7355), .ZN(n10024) );
  NAND2_X1 U10151 ( .A1(n10022), .A2(n10023), .ZN(n10139) );
  NAND2_X1 U10152 ( .A1(n10142), .A2(n10143), .ZN(n10023) );
  NAND3_X1 U10153 ( .A1(a_14_), .A2(n10144), .A3(b_20_), .ZN(n10143) );
  NAND2_X1 U10154 ( .A1(n10019), .A2(n10018), .ZN(n10144) );
  OR2_X1 U10155 ( .A1(n10018), .A2(n10019), .ZN(n10142) );
  AND2_X1 U10156 ( .A1(n10145), .A2(n10146), .ZN(n10019) );
  NAND2_X1 U10157 ( .A1(n10016), .A2(n10147), .ZN(n10146) );
  OR2_X1 U10158 ( .A1(n10015), .A2(n10013), .ZN(n10147) );
  NOR2_X1 U10159 ( .A1(n9746), .A2(n7346), .ZN(n10016) );
  NAND2_X1 U10160 ( .A1(n10013), .A2(n10015), .ZN(n10145) );
  NAND2_X1 U10161 ( .A1(n10148), .A2(n10149), .ZN(n10015) );
  NAND3_X1 U10162 ( .A1(a_16_), .A2(n10150), .A3(b_20_), .ZN(n10149) );
  NAND2_X1 U10163 ( .A1(n10011), .A2(n10010), .ZN(n10150) );
  OR2_X1 U10164 ( .A1(n10010), .A2(n10011), .ZN(n10148) );
  AND2_X1 U10165 ( .A1(n10151), .A2(n10152), .ZN(n10011) );
  NAND2_X1 U10166 ( .A1(n10008), .A2(n10153), .ZN(n10152) );
  OR2_X1 U10167 ( .A1(n10007), .A2(n10005), .ZN(n10153) );
  NOR2_X1 U10168 ( .A1(n9746), .A2(n7337), .ZN(n10008) );
  NAND2_X1 U10169 ( .A1(n10005), .A2(n10007), .ZN(n10151) );
  NAND2_X1 U10170 ( .A1(n10154), .A2(n10155), .ZN(n10007) );
  NAND3_X1 U10171 ( .A1(a_18_), .A2(n10156), .A3(b_20_), .ZN(n10155) );
  NAND2_X1 U10172 ( .A1(n10003), .A2(n10002), .ZN(n10156) );
  OR2_X1 U10173 ( .A1(n10002), .A2(n10003), .ZN(n10154) );
  AND2_X1 U10174 ( .A1(n10157), .A2(n10158), .ZN(n10003) );
  NAND2_X1 U10175 ( .A1(n10000), .A2(n10159), .ZN(n10158) );
  OR2_X1 U10176 ( .A1(n9999), .A2(n9997), .ZN(n10159) );
  NOR2_X1 U10177 ( .A1(n9746), .A2(n7902), .ZN(n10000) );
  NAND2_X1 U10178 ( .A1(n9997), .A2(n9999), .ZN(n10157) );
  NAND2_X1 U10179 ( .A1(n10160), .A2(n10161), .ZN(n9999) );
  NAND2_X1 U10180 ( .A1(n9996), .A2(n10162), .ZN(n10161) );
  OR2_X1 U10181 ( .A1(n9995), .A2(n9994), .ZN(n10162) );
  INV_X1 U10182 ( .A(n10163), .ZN(n9996) );
  NAND2_X1 U10183 ( .A1(n9994), .A2(n9995), .ZN(n10160) );
  NAND2_X1 U10184 ( .A1(n10164), .A2(n10165), .ZN(n9995) );
  NAND2_X1 U10185 ( .A1(n9992), .A2(n10166), .ZN(n10165) );
  OR2_X1 U10186 ( .A1(n9991), .A2(n9990), .ZN(n10166) );
  NOR2_X1 U10187 ( .A1(n9746), .A2(n7909), .ZN(n9992) );
  NAND2_X1 U10188 ( .A1(n9990), .A2(n9991), .ZN(n10164) );
  NAND2_X1 U10189 ( .A1(n10167), .A2(n10168), .ZN(n9991) );
  NAND3_X1 U10190 ( .A1(a_22_), .A2(n10169), .A3(b_20_), .ZN(n10168) );
  OR2_X1 U10191 ( .A1(n9987), .A2(n9985), .ZN(n10169) );
  NAND2_X1 U10192 ( .A1(n9985), .A2(n9987), .ZN(n10167) );
  NAND2_X1 U10193 ( .A1(n10170), .A2(n10171), .ZN(n9987) );
  NAND2_X1 U10194 ( .A1(n9984), .A2(n10172), .ZN(n10171) );
  OR2_X1 U10195 ( .A1(n9983), .A2(n9981), .ZN(n10172) );
  NOR2_X1 U10196 ( .A1(n9746), .A2(n7916), .ZN(n9984) );
  NAND2_X1 U10197 ( .A1(n9981), .A2(n9983), .ZN(n10170) );
  NAND2_X1 U10198 ( .A1(n10173), .A2(n10174), .ZN(n9983) );
  NAND3_X1 U10199 ( .A1(a_24_), .A2(n10175), .A3(b_20_), .ZN(n10174) );
  NAND2_X1 U10200 ( .A1(n9979), .A2(n9978), .ZN(n10175) );
  OR2_X1 U10201 ( .A1(n9978), .A2(n9979), .ZN(n10173) );
  AND2_X1 U10202 ( .A1(n10176), .A2(n10177), .ZN(n9979) );
  NAND2_X1 U10203 ( .A1(n9976), .A2(n10178), .ZN(n10177) );
  OR2_X1 U10204 ( .A1(n9975), .A2(n9974), .ZN(n10178) );
  NOR2_X1 U10205 ( .A1(n9746), .A2(n7923), .ZN(n9976) );
  NAND2_X1 U10206 ( .A1(n9974), .A2(n9975), .ZN(n10176) );
  NAND2_X1 U10207 ( .A1(n9971), .A2(n10179), .ZN(n9975) );
  NAND2_X1 U10208 ( .A1(n9970), .A2(n9972), .ZN(n10179) );
  NAND2_X1 U10209 ( .A1(n10180), .A2(n10181), .ZN(n9972) );
  NAND2_X1 U10210 ( .A1(b_20_), .A2(a_26_), .ZN(n10181) );
  INV_X1 U10211 ( .A(n10182), .ZN(n10180) );
  XNOR2_X1 U10212 ( .A(n10183), .B(n10184), .ZN(n9970) );
  NAND2_X1 U10213 ( .A1(n10185), .A2(n10186), .ZN(n10183) );
  NAND2_X1 U10214 ( .A1(a_26_), .A2(n10182), .ZN(n9971) );
  NAND2_X1 U10215 ( .A1(n9942), .A2(n10187), .ZN(n10182) );
  NAND2_X1 U10216 ( .A1(n9941), .A2(n9943), .ZN(n10187) );
  NAND2_X1 U10217 ( .A1(n10188), .A2(n10189), .ZN(n9943) );
  NAND2_X1 U10218 ( .A1(b_20_), .A2(a_27_), .ZN(n10189) );
  INV_X1 U10219 ( .A(n10190), .ZN(n10188) );
  XNOR2_X1 U10220 ( .A(n10191), .B(n10192), .ZN(n9941) );
  XOR2_X1 U10221 ( .A(n10193), .B(n10194), .Z(n10191) );
  NAND2_X1 U10222 ( .A1(b_19_), .A2(a_28_), .ZN(n10193) );
  NAND2_X1 U10223 ( .A1(a_27_), .A2(n10190), .ZN(n9942) );
  NAND2_X1 U10224 ( .A1(n10195), .A2(n10196), .ZN(n10190) );
  NAND3_X1 U10225 ( .A1(a_28_), .A2(n10197), .A3(b_20_), .ZN(n10196) );
  NAND2_X1 U10226 ( .A1(n9951), .A2(n9949), .ZN(n10197) );
  OR2_X1 U10227 ( .A1(n9949), .A2(n9951), .ZN(n10195) );
  AND2_X1 U10228 ( .A1(n10198), .A2(n10199), .ZN(n9951) );
  NAND2_X1 U10229 ( .A1(n9966), .A2(n10200), .ZN(n10199) );
  OR2_X1 U10230 ( .A1(n9967), .A2(n9968), .ZN(n10200) );
  NOR2_X1 U10231 ( .A1(n9746), .A2(n7946), .ZN(n9966) );
  NAND2_X1 U10232 ( .A1(n9968), .A2(n9967), .ZN(n10198) );
  NAND2_X1 U10233 ( .A1(n10201), .A2(n10202), .ZN(n9967) );
  NAND2_X1 U10234 ( .A1(b_18_), .A2(n10203), .ZN(n10202) );
  NAND2_X1 U10235 ( .A1(n7268), .A2(n10204), .ZN(n10203) );
  NAND2_X1 U10236 ( .A1(a_31_), .A2(n9964), .ZN(n10204) );
  NAND2_X1 U10237 ( .A1(b_19_), .A2(n10205), .ZN(n10201) );
  NAND2_X1 U10238 ( .A1(n7272), .A2(n10206), .ZN(n10205) );
  NAND2_X1 U10239 ( .A1(a_30_), .A2(n10207), .ZN(n10206) );
  AND3_X1 U10240 ( .A1(b_19_), .A2(n7954), .A3(b_20_), .ZN(n9968) );
  XNOR2_X1 U10241 ( .A(n10208), .B(n10209), .ZN(n9949) );
  XOR2_X1 U10242 ( .A(n10210), .B(n10211), .Z(n10208) );
  XNOR2_X1 U10243 ( .A(n10212), .B(n10213), .ZN(n9974) );
  NAND2_X1 U10244 ( .A1(n10214), .A2(n10215), .ZN(n10212) );
  XNOR2_X1 U10245 ( .A(n10216), .B(n10217), .ZN(n9978) );
  XOR2_X1 U10246 ( .A(n10218), .B(n10219), .Z(n10216) );
  XNOR2_X1 U10247 ( .A(n10220), .B(n10221), .ZN(n9981) );
  XNOR2_X1 U10248 ( .A(n10222), .B(n10223), .ZN(n10220) );
  NOR2_X1 U10249 ( .A1(n7691), .A2(n9964), .ZN(n10223) );
  XNOR2_X1 U10250 ( .A(n10224), .B(n10225), .ZN(n9985) );
  XNOR2_X1 U10251 ( .A(n10226), .B(n10227), .ZN(n10225) );
  XNOR2_X1 U10252 ( .A(n10228), .B(n10229), .ZN(n9990) );
  XOR2_X1 U10253 ( .A(n10230), .B(n10231), .Z(n10229) );
  NAND2_X1 U10254 ( .A1(b_19_), .A2(a_22_), .ZN(n10231) );
  XNOR2_X1 U10255 ( .A(n10232), .B(n10233), .ZN(n9994) );
  XNOR2_X1 U10256 ( .A(n10234), .B(n10235), .ZN(n10232) );
  XNOR2_X1 U10257 ( .A(n10236), .B(n10237), .ZN(n9997) );
  XOR2_X1 U10258 ( .A(n10238), .B(n10239), .Z(n10236) );
  NAND2_X1 U10259 ( .A1(b_19_), .A2(a_20_), .ZN(n10238) );
  XNOR2_X1 U10260 ( .A(n10240), .B(n10241), .ZN(n10002) );
  XOR2_X1 U10261 ( .A(n10242), .B(n10243), .Z(n10240) );
  XNOR2_X1 U10262 ( .A(n10244), .B(n10245), .ZN(n10005) );
  XNOR2_X1 U10263 ( .A(n10246), .B(n10247), .ZN(n10244) );
  NOR2_X1 U10264 ( .A1(n7764), .A2(n9964), .ZN(n10247) );
  XNOR2_X1 U10265 ( .A(n10248), .B(n10249), .ZN(n10010) );
  XOR2_X1 U10266 ( .A(n10250), .B(n10251), .Z(n10248) );
  XNOR2_X1 U10267 ( .A(n10252), .B(n10253), .ZN(n10013) );
  XOR2_X1 U10268 ( .A(n10254), .B(n10255), .Z(n10253) );
  NAND2_X1 U10269 ( .A1(b_19_), .A2(a_16_), .ZN(n10255) );
  XOR2_X1 U10270 ( .A(n10256), .B(n10257), .Z(n10018) );
  XNOR2_X1 U10271 ( .A(n10258), .B(n10259), .ZN(n10257) );
  XNOR2_X1 U10272 ( .A(n10260), .B(n10261), .ZN(n10022) );
  XOR2_X1 U10273 ( .A(n10262), .B(n10263), .Z(n10260) );
  NAND2_X1 U10274 ( .A1(b_19_), .A2(a_14_), .ZN(n10262) );
  XNOR2_X1 U10275 ( .A(n10264), .B(n10265), .ZN(n10026) );
  XOR2_X1 U10276 ( .A(n10266), .B(n10267), .Z(n10264) );
  XOR2_X1 U10277 ( .A(n10268), .B(n10269), .Z(n10029) );
  XOR2_X1 U10278 ( .A(n10270), .B(n10271), .Z(n10268) );
  XNOR2_X1 U10279 ( .A(n10272), .B(n10273), .ZN(n10034) );
  XOR2_X1 U10280 ( .A(n10274), .B(n10275), .Z(n10273) );
  NAND2_X1 U10281 ( .A1(b_19_), .A2(a_11_), .ZN(n10275) );
  XNOR2_X1 U10282 ( .A(n10276), .B(n10277), .ZN(n10038) );
  NAND2_X1 U10283 ( .A1(n10278), .A2(n10279), .ZN(n10276) );
  XNOR2_X1 U10284 ( .A(n10280), .B(n10281), .ZN(n10042) );
  XOR2_X1 U10285 ( .A(n10282), .B(n10283), .Z(n10280) );
  NOR2_X1 U10286 ( .A1(n7870), .A2(n9964), .ZN(n10283) );
  XNOR2_X1 U10287 ( .A(n10284), .B(n10285), .ZN(n10056) );
  XNOR2_X1 U10288 ( .A(n10286), .B(n10287), .ZN(n10284) );
  NOR2_X1 U10289 ( .A1(n7388), .A2(n9964), .ZN(n10287) );
  XNOR2_X1 U10290 ( .A(n10288), .B(n10289), .ZN(n10060) );
  XNOR2_X1 U10291 ( .A(n10290), .B(n10291), .ZN(n10288) );
  NOR2_X1 U10292 ( .A1(n7393), .A2(n9964), .ZN(n10291) );
  XOR2_X1 U10293 ( .A(n10292), .B(n10293), .Z(n10072) );
  XOR2_X1 U10294 ( .A(n10294), .B(n10295), .Z(n10293) );
  NAND2_X1 U10295 ( .A1(b_19_), .A2(a_2_), .ZN(n10295) );
  XNOR2_X1 U10296 ( .A(n10296), .B(n10297), .ZN(n10076) );
  XNOR2_X1 U10297 ( .A(n10298), .B(n10299), .ZN(n10296) );
  NOR2_X1 U10298 ( .A1(n7411), .A2(n9964), .ZN(n10299) );
  INV_X1 U10299 ( .A(n7566), .ZN(n7561) );
  XOR2_X1 U10300 ( .A(n10300), .B(n10301), .Z(n7566) );
  XOR2_X1 U10301 ( .A(n10302), .B(n10303), .Z(n10301) );
  NAND2_X1 U10302 ( .A1(b_19_), .A2(a_0_), .ZN(n10303) );
  NAND3_X1 U10303 ( .A1(n10304), .A2(n7555), .A3(n7554), .ZN(n7475) );
  XOR2_X1 U10304 ( .A(n10305), .B(n10306), .Z(n7554) );
  XOR2_X1 U10305 ( .A(n10307), .B(n10308), .Z(n10305) );
  NOR2_X1 U10306 ( .A1(n7613), .A2(n10207), .ZN(n10308) );
  NAND2_X1 U10307 ( .A1(n10309), .A2(n10310), .ZN(n7555) );
  NAND3_X1 U10308 ( .A1(a_0_), .A2(n10311), .A3(b_19_), .ZN(n10310) );
  OR2_X1 U10309 ( .A1(n10302), .A2(n10300), .ZN(n10311) );
  NAND2_X1 U10310 ( .A1(n10300), .A2(n10302), .ZN(n10309) );
  NAND2_X1 U10311 ( .A1(n10312), .A2(n10313), .ZN(n10302) );
  NAND3_X1 U10312 ( .A1(a_1_), .A2(n10314), .A3(b_19_), .ZN(n10313) );
  NAND2_X1 U10313 ( .A1(n10298), .A2(n10297), .ZN(n10314) );
  OR2_X1 U10314 ( .A1(n10297), .A2(n10298), .ZN(n10312) );
  AND2_X1 U10315 ( .A1(n10315), .A2(n10316), .ZN(n10298) );
  NAND3_X1 U10316 ( .A1(a_2_), .A2(n10317), .A3(b_19_), .ZN(n10316) );
  OR2_X1 U10317 ( .A1(n10294), .A2(n10292), .ZN(n10317) );
  NAND2_X1 U10318 ( .A1(n10292), .A2(n10294), .ZN(n10315) );
  NAND2_X1 U10319 ( .A1(n10318), .A2(n10319), .ZN(n10294) );
  NAND3_X1 U10320 ( .A1(a_3_), .A2(n10320), .A3(b_19_), .ZN(n10319) );
  OR2_X1 U10321 ( .A1(n10092), .A2(n10090), .ZN(n10320) );
  NAND2_X1 U10322 ( .A1(n10090), .A2(n10092), .ZN(n10318) );
  NAND2_X1 U10323 ( .A1(n10321), .A2(n10322), .ZN(n10092) );
  NAND3_X1 U10324 ( .A1(a_4_), .A2(n10323), .A3(b_19_), .ZN(n10322) );
  OR2_X1 U10325 ( .A1(n10100), .A2(n10099), .ZN(n10323) );
  NAND2_X1 U10326 ( .A1(n10099), .A2(n10100), .ZN(n10321) );
  NAND2_X1 U10327 ( .A1(n10324), .A2(n10325), .ZN(n10100) );
  NAND3_X1 U10328 ( .A1(a_5_), .A2(n10326), .A3(b_19_), .ZN(n10325) );
  NAND2_X1 U10329 ( .A1(n10290), .A2(n10289), .ZN(n10326) );
  OR2_X1 U10330 ( .A1(n10289), .A2(n10290), .ZN(n10324) );
  AND2_X1 U10331 ( .A1(n10327), .A2(n10328), .ZN(n10290) );
  NAND3_X1 U10332 ( .A1(a_6_), .A2(n10329), .A3(b_19_), .ZN(n10328) );
  NAND2_X1 U10333 ( .A1(n10286), .A2(n10285), .ZN(n10329) );
  OR2_X1 U10334 ( .A1(n10285), .A2(n10286), .ZN(n10327) );
  AND2_X1 U10335 ( .A1(n10330), .A2(n10331), .ZN(n10286) );
  NAND3_X1 U10336 ( .A1(a_7_), .A2(n10332), .A3(b_19_), .ZN(n10331) );
  OR2_X1 U10337 ( .A1(n10114), .A2(n10112), .ZN(n10332) );
  NAND2_X1 U10338 ( .A1(n10112), .A2(n10114), .ZN(n10330) );
  NAND2_X1 U10339 ( .A1(n10333), .A2(n10334), .ZN(n10114) );
  NAND3_X1 U10340 ( .A1(a_8_), .A2(n10335), .A3(b_19_), .ZN(n10334) );
  OR2_X1 U10341 ( .A1(n10122), .A2(n10120), .ZN(n10335) );
  NAND2_X1 U10342 ( .A1(n10120), .A2(n10122), .ZN(n10333) );
  NAND2_X1 U10343 ( .A1(n10336), .A2(n10337), .ZN(n10122) );
  NAND3_X1 U10344 ( .A1(a_9_), .A2(n10338), .A3(b_19_), .ZN(n10337) );
  OR2_X1 U10345 ( .A1(n10282), .A2(n10281), .ZN(n10338) );
  NAND2_X1 U10346 ( .A1(n10281), .A2(n10282), .ZN(n10336) );
  NAND2_X1 U10347 ( .A1(n10278), .A2(n10339), .ZN(n10282) );
  NAND2_X1 U10348 ( .A1(n10277), .A2(n10279), .ZN(n10339) );
  NAND2_X1 U10349 ( .A1(n10340), .A2(n10341), .ZN(n10279) );
  NAND2_X1 U10350 ( .A1(b_19_), .A2(a_10_), .ZN(n10341) );
  INV_X1 U10351 ( .A(n10342), .ZN(n10340) );
  XNOR2_X1 U10352 ( .A(n10343), .B(n10344), .ZN(n10277) );
  XNOR2_X1 U10353 ( .A(n10345), .B(n10346), .ZN(n10343) );
  NAND2_X1 U10354 ( .A1(a_10_), .A2(n10342), .ZN(n10278) );
  NAND2_X1 U10355 ( .A1(n10347), .A2(n10348), .ZN(n10342) );
  NAND3_X1 U10356 ( .A1(a_11_), .A2(n10349), .A3(b_19_), .ZN(n10348) );
  OR2_X1 U10357 ( .A1(n10274), .A2(n10272), .ZN(n10349) );
  NAND2_X1 U10358 ( .A1(n10272), .A2(n10274), .ZN(n10347) );
  NAND2_X1 U10359 ( .A1(n10350), .A2(n10351), .ZN(n10274) );
  NAND2_X1 U10360 ( .A1(n10271), .A2(n10352), .ZN(n10351) );
  OR2_X1 U10361 ( .A1(n10270), .A2(n10269), .ZN(n10352) );
  NOR2_X1 U10362 ( .A1(n9964), .A2(n8020), .ZN(n10271) );
  NAND2_X1 U10363 ( .A1(n10269), .A2(n10270), .ZN(n10350) );
  NAND2_X1 U10364 ( .A1(n10353), .A2(n10354), .ZN(n10270) );
  NAND2_X1 U10365 ( .A1(n10267), .A2(n10355), .ZN(n10354) );
  OR2_X1 U10366 ( .A1(n10266), .A2(n10265), .ZN(n10355) );
  NOR2_X1 U10367 ( .A1(n9964), .A2(n7355), .ZN(n10267) );
  NAND2_X1 U10368 ( .A1(n10265), .A2(n10266), .ZN(n10353) );
  NAND2_X1 U10369 ( .A1(n10356), .A2(n10357), .ZN(n10266) );
  NAND3_X1 U10370 ( .A1(a_14_), .A2(n10358), .A3(b_19_), .ZN(n10357) );
  NAND2_X1 U10371 ( .A1(n10263), .A2(n10261), .ZN(n10358) );
  OR2_X1 U10372 ( .A1(n10261), .A2(n10263), .ZN(n10356) );
  AND2_X1 U10373 ( .A1(n10359), .A2(n10360), .ZN(n10263) );
  NAND2_X1 U10374 ( .A1(n10259), .A2(n10361), .ZN(n10360) );
  OR2_X1 U10375 ( .A1(n10258), .A2(n10256), .ZN(n10361) );
  NOR2_X1 U10376 ( .A1(n9964), .A2(n7346), .ZN(n10259) );
  NAND2_X1 U10377 ( .A1(n10256), .A2(n10258), .ZN(n10359) );
  NAND2_X1 U10378 ( .A1(n10362), .A2(n10363), .ZN(n10258) );
  NAND3_X1 U10379 ( .A1(a_16_), .A2(n10364), .A3(b_19_), .ZN(n10363) );
  OR2_X1 U10380 ( .A1(n10254), .A2(n10252), .ZN(n10364) );
  NAND2_X1 U10381 ( .A1(n10252), .A2(n10254), .ZN(n10362) );
  NAND2_X1 U10382 ( .A1(n10365), .A2(n10366), .ZN(n10254) );
  NAND2_X1 U10383 ( .A1(n10251), .A2(n10367), .ZN(n10366) );
  OR2_X1 U10384 ( .A1(n10250), .A2(n10249), .ZN(n10367) );
  NOR2_X1 U10385 ( .A1(n9964), .A2(n7337), .ZN(n10251) );
  NAND2_X1 U10386 ( .A1(n10249), .A2(n10250), .ZN(n10365) );
  NAND2_X1 U10387 ( .A1(n10368), .A2(n10369), .ZN(n10250) );
  NAND3_X1 U10388 ( .A1(a_18_), .A2(n10370), .A3(b_19_), .ZN(n10369) );
  NAND2_X1 U10389 ( .A1(n10246), .A2(n10245), .ZN(n10370) );
  OR2_X1 U10390 ( .A1(n10245), .A2(n10246), .ZN(n10368) );
  AND2_X1 U10391 ( .A1(n10371), .A2(n10372), .ZN(n10246) );
  NAND2_X1 U10392 ( .A1(n10243), .A2(n10373), .ZN(n10372) );
  OR2_X1 U10393 ( .A1(n10242), .A2(n10241), .ZN(n10373) );
  NAND2_X1 U10394 ( .A1(n10241), .A2(n10242), .ZN(n10371) );
  NAND2_X1 U10395 ( .A1(n10374), .A2(n10375), .ZN(n10242) );
  NAND3_X1 U10396 ( .A1(a_20_), .A2(n10376), .A3(b_19_), .ZN(n10375) );
  NAND2_X1 U10397 ( .A1(n10239), .A2(n10237), .ZN(n10376) );
  OR2_X1 U10398 ( .A1(n10237), .A2(n10239), .ZN(n10374) );
  AND2_X1 U10399 ( .A1(n10377), .A2(n10378), .ZN(n10239) );
  NAND2_X1 U10400 ( .A1(n10235), .A2(n10379), .ZN(n10378) );
  NAND2_X1 U10401 ( .A1(n10234), .A2(n10233), .ZN(n10379) );
  NOR2_X1 U10402 ( .A1(n9964), .A2(n7909), .ZN(n10235) );
  OR2_X1 U10403 ( .A1(n10233), .A2(n10234), .ZN(n10377) );
  AND2_X1 U10404 ( .A1(n10380), .A2(n10381), .ZN(n10234) );
  NAND3_X1 U10405 ( .A1(a_22_), .A2(n10382), .A3(b_19_), .ZN(n10381) );
  OR2_X1 U10406 ( .A1(n10230), .A2(n10228), .ZN(n10382) );
  NAND2_X1 U10407 ( .A1(n10228), .A2(n10230), .ZN(n10380) );
  NAND2_X1 U10408 ( .A1(n10383), .A2(n10384), .ZN(n10230) );
  NAND2_X1 U10409 ( .A1(n10227), .A2(n10385), .ZN(n10384) );
  OR2_X1 U10410 ( .A1(n10226), .A2(n10224), .ZN(n10385) );
  NOR2_X1 U10411 ( .A1(n9964), .A2(n7916), .ZN(n10227) );
  NAND2_X1 U10412 ( .A1(n10224), .A2(n10226), .ZN(n10383) );
  NAND2_X1 U10413 ( .A1(n10386), .A2(n10387), .ZN(n10226) );
  NAND3_X1 U10414 ( .A1(a_24_), .A2(n10388), .A3(b_19_), .ZN(n10387) );
  NAND2_X1 U10415 ( .A1(n10222), .A2(n10221), .ZN(n10388) );
  OR2_X1 U10416 ( .A1(n10221), .A2(n10222), .ZN(n10386) );
  AND2_X1 U10417 ( .A1(n10389), .A2(n10390), .ZN(n10222) );
  NAND2_X1 U10418 ( .A1(n10219), .A2(n10391), .ZN(n10390) );
  OR2_X1 U10419 ( .A1(n10218), .A2(n10217), .ZN(n10391) );
  NOR2_X1 U10420 ( .A1(n9964), .A2(n7923), .ZN(n10219) );
  NAND2_X1 U10421 ( .A1(n10217), .A2(n10218), .ZN(n10389) );
  NAND2_X1 U10422 ( .A1(n10214), .A2(n10392), .ZN(n10218) );
  NAND2_X1 U10423 ( .A1(n10213), .A2(n10215), .ZN(n10392) );
  NAND2_X1 U10424 ( .A1(n10393), .A2(n10394), .ZN(n10215) );
  NAND2_X1 U10425 ( .A1(b_19_), .A2(a_26_), .ZN(n10394) );
  INV_X1 U10426 ( .A(n10395), .ZN(n10393) );
  XNOR2_X1 U10427 ( .A(n10396), .B(n10397), .ZN(n10213) );
  NAND2_X1 U10428 ( .A1(n10398), .A2(n10399), .ZN(n10396) );
  NAND2_X1 U10429 ( .A1(a_26_), .A2(n10395), .ZN(n10214) );
  NAND2_X1 U10430 ( .A1(n10185), .A2(n10400), .ZN(n10395) );
  NAND2_X1 U10431 ( .A1(n10184), .A2(n10186), .ZN(n10400) );
  NAND2_X1 U10432 ( .A1(n10401), .A2(n10402), .ZN(n10186) );
  NAND2_X1 U10433 ( .A1(b_19_), .A2(a_27_), .ZN(n10402) );
  INV_X1 U10434 ( .A(n10403), .ZN(n10401) );
  XNOR2_X1 U10435 ( .A(n10404), .B(n10405), .ZN(n10184) );
  XOR2_X1 U10436 ( .A(n10406), .B(n10407), .Z(n10404) );
  NAND2_X1 U10437 ( .A1(b_18_), .A2(a_28_), .ZN(n10406) );
  NAND2_X1 U10438 ( .A1(a_27_), .A2(n10403), .ZN(n10185) );
  NAND2_X1 U10439 ( .A1(n10408), .A2(n10409), .ZN(n10403) );
  NAND3_X1 U10440 ( .A1(a_28_), .A2(n10410), .A3(b_19_), .ZN(n10409) );
  NAND2_X1 U10441 ( .A1(n10194), .A2(n10192), .ZN(n10410) );
  OR2_X1 U10442 ( .A1(n10192), .A2(n10194), .ZN(n10408) );
  AND2_X1 U10443 ( .A1(n10411), .A2(n10412), .ZN(n10194) );
  NAND2_X1 U10444 ( .A1(n10209), .A2(n10413), .ZN(n10412) );
  OR2_X1 U10445 ( .A1(n10210), .A2(n10211), .ZN(n10413) );
  NOR2_X1 U10446 ( .A1(n9964), .A2(n7946), .ZN(n10209) );
  NAND2_X1 U10447 ( .A1(n10211), .A2(n10210), .ZN(n10411) );
  NAND2_X1 U10448 ( .A1(n10414), .A2(n10415), .ZN(n10210) );
  NAND2_X1 U10449 ( .A1(b_17_), .A2(n10416), .ZN(n10415) );
  NAND2_X1 U10450 ( .A1(n7268), .A2(n10417), .ZN(n10416) );
  NAND2_X1 U10451 ( .A1(a_31_), .A2(n10207), .ZN(n10417) );
  NAND2_X1 U10452 ( .A1(b_18_), .A2(n10418), .ZN(n10414) );
  NAND2_X1 U10453 ( .A1(n7272), .A2(n10419), .ZN(n10418) );
  NAND2_X1 U10454 ( .A1(a_30_), .A2(n10420), .ZN(n10419) );
  AND3_X1 U10455 ( .A1(b_19_), .A2(n7954), .A3(b_18_), .ZN(n10211) );
  XNOR2_X1 U10456 ( .A(n10421), .B(n10422), .ZN(n10192) );
  XOR2_X1 U10457 ( .A(n10423), .B(n10424), .Z(n10421) );
  XNOR2_X1 U10458 ( .A(n10425), .B(n10426), .ZN(n10217) );
  NAND2_X1 U10459 ( .A1(n10427), .A2(n10428), .ZN(n10425) );
  XNOR2_X1 U10460 ( .A(n10429), .B(n10430), .ZN(n10221) );
  XOR2_X1 U10461 ( .A(n10431), .B(n10432), .Z(n10429) );
  XNOR2_X1 U10462 ( .A(n10433), .B(n10434), .ZN(n10224) );
  XNOR2_X1 U10463 ( .A(n10435), .B(n10436), .ZN(n10433) );
  NOR2_X1 U10464 ( .A1(n7691), .A2(n10207), .ZN(n10436) );
  XNOR2_X1 U10465 ( .A(n10437), .B(n10438), .ZN(n10228) );
  XOR2_X1 U10466 ( .A(n10439), .B(n10440), .Z(n10438) );
  NAND2_X1 U10467 ( .A1(b_18_), .A2(a_23_), .ZN(n10440) );
  XOR2_X1 U10468 ( .A(n10441), .B(n10442), .Z(n10233) );
  NAND2_X1 U10469 ( .A1(n10443), .A2(n10444), .ZN(n10441) );
  XNOR2_X1 U10470 ( .A(n10445), .B(n10446), .ZN(n10237) );
  XOR2_X1 U10471 ( .A(n10447), .B(n10448), .Z(n10445) );
  XNOR2_X1 U10472 ( .A(n10449), .B(n10450), .ZN(n10241) );
  XNOR2_X1 U10473 ( .A(n10451), .B(n10452), .ZN(n10449) );
  NOR2_X1 U10474 ( .A1(n7987), .A2(n10207), .ZN(n10452) );
  XOR2_X1 U10475 ( .A(n10453), .B(n10454), .Z(n10245) );
  XNOR2_X1 U10476 ( .A(n10455), .B(n10456), .ZN(n10454) );
  XNOR2_X1 U10477 ( .A(n10457), .B(n10458), .ZN(n10249) );
  XNOR2_X1 U10478 ( .A(n10459), .B(n10460), .ZN(n10457) );
  XOR2_X1 U10479 ( .A(n10461), .B(n10462), .Z(n10252) );
  XOR2_X1 U10480 ( .A(n10463), .B(n10464), .Z(n10461) );
  XNOR2_X1 U10481 ( .A(n10465), .B(n10466), .ZN(n10256) );
  XOR2_X1 U10482 ( .A(n10467), .B(n10468), .Z(n10466) );
  NAND2_X1 U10483 ( .A1(b_18_), .A2(a_16_), .ZN(n10468) );
  XOR2_X1 U10484 ( .A(n10469), .B(n10470), .Z(n10261) );
  XNOR2_X1 U10485 ( .A(n10471), .B(n10472), .ZN(n10470) );
  XNOR2_X1 U10486 ( .A(n10473), .B(n10474), .ZN(n10265) );
  XNOR2_X1 U10487 ( .A(n10475), .B(n10476), .ZN(n10473) );
  NOR2_X1 U10488 ( .A1(n7782), .A2(n10207), .ZN(n10476) );
  XNOR2_X1 U10489 ( .A(n10477), .B(n10478), .ZN(n10269) );
  XNOR2_X1 U10490 ( .A(n10479), .B(n10480), .ZN(n10477) );
  NOR2_X1 U10491 ( .A1(n7355), .A2(n10207), .ZN(n10480) );
  XNOR2_X1 U10492 ( .A(n10481), .B(n10482), .ZN(n10272) );
  XNOR2_X1 U10493 ( .A(n10483), .B(n10484), .ZN(n10482) );
  XNOR2_X1 U10494 ( .A(n10485), .B(n10486), .ZN(n10281) );
  XNOR2_X1 U10495 ( .A(n10487), .B(n10488), .ZN(n10485) );
  NOR2_X1 U10496 ( .A1(n7799), .A2(n10207), .ZN(n10488) );
  XNOR2_X1 U10497 ( .A(n10489), .B(n10490), .ZN(n10120) );
  NAND2_X1 U10498 ( .A1(n10491), .A2(n10492), .ZN(n10489) );
  XNOR2_X1 U10499 ( .A(n10493), .B(n10494), .ZN(n10112) );
  NAND2_X1 U10500 ( .A1(n10495), .A2(n10496), .ZN(n10493) );
  XOR2_X1 U10501 ( .A(n10497), .B(n10498), .Z(n10285) );
  NAND2_X1 U10502 ( .A1(n10499), .A2(n10500), .ZN(n10497) );
  XOR2_X1 U10503 ( .A(n10501), .B(n10502), .Z(n10289) );
  NAND2_X1 U10504 ( .A1(n10503), .A2(n10504), .ZN(n10501) );
  XNOR2_X1 U10505 ( .A(n10505), .B(n10506), .ZN(n10099) );
  NAND2_X1 U10506 ( .A1(n10507), .A2(n10508), .ZN(n10505) );
  XNOR2_X1 U10507 ( .A(n10509), .B(n10510), .ZN(n10090) );
  NAND2_X1 U10508 ( .A1(n10511), .A2(n10512), .ZN(n10509) );
  XNOR2_X1 U10509 ( .A(n10513), .B(n10514), .ZN(n10292) );
  NAND2_X1 U10510 ( .A1(n10515), .A2(n10516), .ZN(n10513) );
  XOR2_X1 U10511 ( .A(n10517), .B(n10518), .Z(n10297) );
  NAND2_X1 U10512 ( .A1(n10519), .A2(n10520), .ZN(n10517) );
  XNOR2_X1 U10513 ( .A(n10521), .B(n10522), .ZN(n10300) );
  XNOR2_X1 U10514 ( .A(n10523), .B(n10524), .ZN(n10522) );
  XOR2_X1 U10515 ( .A(n7556), .B(n7557), .Z(n10304) );
  NAND2_X1 U10516 ( .A1(n10525), .A2(n10526), .ZN(n7479) );
  NAND2_X1 U10517 ( .A1(n7557), .A2(n7556), .ZN(n10526) );
  XNOR2_X1 U10518 ( .A(n7547), .B(n7546), .ZN(n10525) );
  NAND3_X1 U10519 ( .A1(n10527), .A2(n7556), .A3(n7557), .ZN(n7480) );
  XNOR2_X1 U10520 ( .A(n10528), .B(n10529), .ZN(n7557) );
  XOR2_X1 U10521 ( .A(n10530), .B(n10531), .Z(n10529) );
  NAND2_X1 U10522 ( .A1(b_17_), .A2(a_0_), .ZN(n10531) );
  NAND2_X1 U10523 ( .A1(n10532), .A2(n10533), .ZN(n7556) );
  NAND3_X1 U10524 ( .A1(a_0_), .A2(n10534), .A3(b_18_), .ZN(n10533) );
  OR2_X1 U10525 ( .A1(n10306), .A2(n10307), .ZN(n10534) );
  NAND2_X1 U10526 ( .A1(n10306), .A2(n10307), .ZN(n10532) );
  NAND2_X1 U10527 ( .A1(n10535), .A2(n10536), .ZN(n10307) );
  NAND2_X1 U10528 ( .A1(n10524), .A2(n10537), .ZN(n10536) );
  OR2_X1 U10529 ( .A1(n10521), .A2(n10523), .ZN(n10537) );
  NOR2_X1 U10530 ( .A1(n10207), .A2(n7411), .ZN(n10524) );
  NAND2_X1 U10531 ( .A1(n10521), .A2(n10523), .ZN(n10535) );
  NAND2_X1 U10532 ( .A1(n10519), .A2(n10538), .ZN(n10523) );
  NAND2_X1 U10533 ( .A1(n10518), .A2(n10520), .ZN(n10538) );
  NAND2_X1 U10534 ( .A1(n10539), .A2(n10540), .ZN(n10520) );
  NAND2_X1 U10535 ( .A1(b_18_), .A2(a_2_), .ZN(n10540) );
  INV_X1 U10536 ( .A(n10541), .ZN(n10539) );
  XOR2_X1 U10537 ( .A(n10542), .B(n10543), .Z(n10518) );
  XOR2_X1 U10538 ( .A(n10544), .B(n10545), .Z(n10542) );
  NOR2_X1 U10539 ( .A1(n7850), .A2(n10420), .ZN(n10545) );
  NAND2_X1 U10540 ( .A1(a_2_), .A2(n10541), .ZN(n10519) );
  NAND2_X1 U10541 ( .A1(n10515), .A2(n10546), .ZN(n10541) );
  NAND2_X1 U10542 ( .A1(n10514), .A2(n10516), .ZN(n10546) );
  NAND2_X1 U10543 ( .A1(n10547), .A2(n10548), .ZN(n10516) );
  NAND2_X1 U10544 ( .A1(b_18_), .A2(a_3_), .ZN(n10548) );
  INV_X1 U10545 ( .A(n10549), .ZN(n10547) );
  XNOR2_X1 U10546 ( .A(n10550), .B(n10551), .ZN(n10514) );
  XOR2_X1 U10547 ( .A(n10552), .B(n10553), .Z(n10551) );
  NAND2_X1 U10548 ( .A1(b_17_), .A2(a_4_), .ZN(n10553) );
  NAND2_X1 U10549 ( .A1(a_3_), .A2(n10549), .ZN(n10515) );
  NAND2_X1 U10550 ( .A1(n10511), .A2(n10554), .ZN(n10549) );
  NAND2_X1 U10551 ( .A1(n10510), .A2(n10512), .ZN(n10554) );
  NAND2_X1 U10552 ( .A1(n10555), .A2(n10556), .ZN(n10512) );
  NAND2_X1 U10553 ( .A1(b_18_), .A2(a_4_), .ZN(n10556) );
  INV_X1 U10554 ( .A(n10557), .ZN(n10555) );
  XOR2_X1 U10555 ( .A(n10558), .B(n10559), .Z(n10510) );
  XOR2_X1 U10556 ( .A(n10560), .B(n10561), .Z(n10558) );
  NOR2_X1 U10557 ( .A1(n7393), .A2(n10420), .ZN(n10561) );
  NAND2_X1 U10558 ( .A1(a_4_), .A2(n10557), .ZN(n10511) );
  NAND2_X1 U10559 ( .A1(n10507), .A2(n10562), .ZN(n10557) );
  NAND2_X1 U10560 ( .A1(n10506), .A2(n10508), .ZN(n10562) );
  NAND2_X1 U10561 ( .A1(n10563), .A2(n10564), .ZN(n10508) );
  NAND2_X1 U10562 ( .A1(b_18_), .A2(a_5_), .ZN(n10564) );
  INV_X1 U10563 ( .A(n10565), .ZN(n10563) );
  XNOR2_X1 U10564 ( .A(n10566), .B(n10567), .ZN(n10506) );
  XOR2_X1 U10565 ( .A(n10568), .B(n10569), .Z(n10567) );
  NAND2_X1 U10566 ( .A1(b_17_), .A2(a_6_), .ZN(n10569) );
  NAND2_X1 U10567 ( .A1(a_5_), .A2(n10565), .ZN(n10507) );
  NAND2_X1 U10568 ( .A1(n10503), .A2(n10570), .ZN(n10565) );
  NAND2_X1 U10569 ( .A1(n10502), .A2(n10504), .ZN(n10570) );
  NAND2_X1 U10570 ( .A1(n10571), .A2(n10572), .ZN(n10504) );
  NAND2_X1 U10571 ( .A1(b_18_), .A2(a_6_), .ZN(n10572) );
  INV_X1 U10572 ( .A(n10573), .ZN(n10571) );
  XNOR2_X1 U10573 ( .A(n10574), .B(n10575), .ZN(n10502) );
  XOR2_X1 U10574 ( .A(n10576), .B(n10577), .Z(n10575) );
  NAND2_X1 U10575 ( .A1(b_17_), .A2(a_7_), .ZN(n10577) );
  NAND2_X1 U10576 ( .A1(a_6_), .A2(n10573), .ZN(n10503) );
  NAND2_X1 U10577 ( .A1(n10499), .A2(n10578), .ZN(n10573) );
  NAND2_X1 U10578 ( .A1(n10498), .A2(n10500), .ZN(n10578) );
  NAND2_X1 U10579 ( .A1(n10579), .A2(n10580), .ZN(n10500) );
  NAND2_X1 U10580 ( .A1(b_18_), .A2(a_7_), .ZN(n10580) );
  INV_X1 U10581 ( .A(n10581), .ZN(n10579) );
  XNOR2_X1 U10582 ( .A(n10582), .B(n10583), .ZN(n10498) );
  XOR2_X1 U10583 ( .A(n10584), .B(n10585), .Z(n10583) );
  NAND2_X1 U10584 ( .A1(b_17_), .A2(a_8_), .ZN(n10585) );
  NAND2_X1 U10585 ( .A1(a_7_), .A2(n10581), .ZN(n10499) );
  NAND2_X1 U10586 ( .A1(n10495), .A2(n10586), .ZN(n10581) );
  NAND2_X1 U10587 ( .A1(n10494), .A2(n10496), .ZN(n10586) );
  NAND2_X1 U10588 ( .A1(n10587), .A2(n10588), .ZN(n10496) );
  NAND2_X1 U10589 ( .A1(b_18_), .A2(a_8_), .ZN(n10588) );
  INV_X1 U10590 ( .A(n10589), .ZN(n10587) );
  XNOR2_X1 U10591 ( .A(n10590), .B(n10591), .ZN(n10494) );
  XNOR2_X1 U10592 ( .A(n10592), .B(n10593), .ZN(n10590) );
  NOR2_X1 U10593 ( .A1(n7870), .A2(n10420), .ZN(n10593) );
  NAND2_X1 U10594 ( .A1(a_8_), .A2(n10589), .ZN(n10495) );
  NAND2_X1 U10595 ( .A1(n10491), .A2(n10594), .ZN(n10589) );
  NAND2_X1 U10596 ( .A1(n10490), .A2(n10492), .ZN(n10594) );
  NAND2_X1 U10597 ( .A1(n10595), .A2(n10596), .ZN(n10492) );
  NAND2_X1 U10598 ( .A1(b_18_), .A2(a_9_), .ZN(n10596) );
  INV_X1 U10599 ( .A(n10597), .ZN(n10595) );
  XNOR2_X1 U10600 ( .A(n10598), .B(n10599), .ZN(n10490) );
  XNOR2_X1 U10601 ( .A(n10600), .B(n10601), .ZN(n10598) );
  NOR2_X1 U10602 ( .A1(n7799), .A2(n10420), .ZN(n10601) );
  NAND2_X1 U10603 ( .A1(a_9_), .A2(n10597), .ZN(n10491) );
  NAND2_X1 U10604 ( .A1(n10602), .A2(n10603), .ZN(n10597) );
  NAND3_X1 U10605 ( .A1(a_10_), .A2(n10604), .A3(b_18_), .ZN(n10603) );
  NAND2_X1 U10606 ( .A1(n10487), .A2(n10486), .ZN(n10604) );
  OR2_X1 U10607 ( .A1(n10486), .A2(n10487), .ZN(n10602) );
  AND2_X1 U10608 ( .A1(n10605), .A2(n10606), .ZN(n10487) );
  NAND2_X1 U10609 ( .A1(n10346), .A2(n10607), .ZN(n10606) );
  NAND2_X1 U10610 ( .A1(n10345), .A2(n10344), .ZN(n10607) );
  NOR2_X1 U10611 ( .A1(n10207), .A2(n7877), .ZN(n10346) );
  OR2_X1 U10612 ( .A1(n10344), .A2(n10345), .ZN(n10605) );
  AND2_X1 U10613 ( .A1(n10608), .A2(n10609), .ZN(n10345) );
  NAND2_X1 U10614 ( .A1(n10484), .A2(n10610), .ZN(n10609) );
  OR2_X1 U10615 ( .A1(n10481), .A2(n10483), .ZN(n10610) );
  NOR2_X1 U10616 ( .A1(n10207), .A2(n8020), .ZN(n10484) );
  NAND2_X1 U10617 ( .A1(n10481), .A2(n10483), .ZN(n10608) );
  NAND2_X1 U10618 ( .A1(n10611), .A2(n10612), .ZN(n10483) );
  NAND3_X1 U10619 ( .A1(a_13_), .A2(n10613), .A3(b_18_), .ZN(n10612) );
  NAND2_X1 U10620 ( .A1(n10479), .A2(n10478), .ZN(n10613) );
  OR2_X1 U10621 ( .A1(n10478), .A2(n10479), .ZN(n10611) );
  AND2_X1 U10622 ( .A1(n10614), .A2(n10615), .ZN(n10479) );
  NAND3_X1 U10623 ( .A1(a_14_), .A2(n10616), .A3(b_18_), .ZN(n10615) );
  NAND2_X1 U10624 ( .A1(n10475), .A2(n10474), .ZN(n10616) );
  OR2_X1 U10625 ( .A1(n10474), .A2(n10475), .ZN(n10614) );
  AND2_X1 U10626 ( .A1(n10617), .A2(n10618), .ZN(n10475) );
  NAND2_X1 U10627 ( .A1(n10472), .A2(n10619), .ZN(n10618) );
  OR2_X1 U10628 ( .A1(n10469), .A2(n10471), .ZN(n10619) );
  NOR2_X1 U10629 ( .A1(n10207), .A2(n7346), .ZN(n10472) );
  NAND2_X1 U10630 ( .A1(n10469), .A2(n10471), .ZN(n10617) );
  NAND2_X1 U10631 ( .A1(n10620), .A2(n10621), .ZN(n10471) );
  NAND3_X1 U10632 ( .A1(a_16_), .A2(n10622), .A3(b_18_), .ZN(n10621) );
  OR2_X1 U10633 ( .A1(n10467), .A2(n10465), .ZN(n10622) );
  NAND2_X1 U10634 ( .A1(n10465), .A2(n10467), .ZN(n10620) );
  NAND2_X1 U10635 ( .A1(n10623), .A2(n10624), .ZN(n10467) );
  NAND2_X1 U10636 ( .A1(n10464), .A2(n10625), .ZN(n10624) );
  OR2_X1 U10637 ( .A1(n10462), .A2(n10463), .ZN(n10625) );
  NOR2_X1 U10638 ( .A1(n10207), .A2(n7337), .ZN(n10464) );
  NAND2_X1 U10639 ( .A1(n10462), .A2(n10463), .ZN(n10623) );
  NAND2_X1 U10640 ( .A1(n10626), .A2(n10627), .ZN(n10463) );
  NAND2_X1 U10641 ( .A1(n10460), .A2(n10628), .ZN(n10627) );
  NAND2_X1 U10642 ( .A1(n10459), .A2(n10458), .ZN(n10628) );
  OR2_X1 U10643 ( .A1(n10458), .A2(n10459), .ZN(n10626) );
  AND2_X1 U10644 ( .A1(n10629), .A2(n10630), .ZN(n10459) );
  NAND2_X1 U10645 ( .A1(n10456), .A2(n10631), .ZN(n10630) );
  OR2_X1 U10646 ( .A1(n10453), .A2(n10455), .ZN(n10631) );
  NOR2_X1 U10647 ( .A1(n10207), .A2(n7902), .ZN(n10456) );
  NAND2_X1 U10648 ( .A1(n10453), .A2(n10455), .ZN(n10629) );
  NAND2_X1 U10649 ( .A1(n10632), .A2(n10633), .ZN(n10455) );
  NAND3_X1 U10650 ( .A1(a_20_), .A2(n10634), .A3(b_18_), .ZN(n10633) );
  NAND2_X1 U10651 ( .A1(n10451), .A2(n10450), .ZN(n10634) );
  OR2_X1 U10652 ( .A1(n10450), .A2(n10451), .ZN(n10632) );
  AND2_X1 U10653 ( .A1(n10635), .A2(n10636), .ZN(n10451) );
  NAND2_X1 U10654 ( .A1(n10447), .A2(n10637), .ZN(n10636) );
  OR2_X1 U10655 ( .A1(n10446), .A2(n10448), .ZN(n10637) );
  NOR2_X1 U10656 ( .A1(n10207), .A2(n7909), .ZN(n10447) );
  NAND2_X1 U10657 ( .A1(n10446), .A2(n10448), .ZN(n10635) );
  NAND2_X1 U10658 ( .A1(n10443), .A2(n10638), .ZN(n10448) );
  NAND2_X1 U10659 ( .A1(n10442), .A2(n10444), .ZN(n10638) );
  NAND2_X1 U10660 ( .A1(n10639), .A2(n10640), .ZN(n10444) );
  NAND2_X1 U10661 ( .A1(b_18_), .A2(a_22_), .ZN(n10640) );
  INV_X1 U10662 ( .A(n10641), .ZN(n10639) );
  XNOR2_X1 U10663 ( .A(n10642), .B(n10643), .ZN(n10442) );
  XNOR2_X1 U10664 ( .A(n10644), .B(n10645), .ZN(n10643) );
  NAND2_X1 U10665 ( .A1(a_22_), .A2(n10641), .ZN(n10443) );
  NAND2_X1 U10666 ( .A1(n10646), .A2(n10647), .ZN(n10641) );
  NAND3_X1 U10667 ( .A1(a_23_), .A2(n10648), .A3(b_18_), .ZN(n10647) );
  OR2_X1 U10668 ( .A1(n10437), .A2(n10439), .ZN(n10648) );
  NAND2_X1 U10669 ( .A1(n10437), .A2(n10439), .ZN(n10646) );
  NAND2_X1 U10670 ( .A1(n10649), .A2(n10650), .ZN(n10439) );
  NAND3_X1 U10671 ( .A1(a_24_), .A2(n10651), .A3(b_18_), .ZN(n10650) );
  NAND2_X1 U10672 ( .A1(n10435), .A2(n10434), .ZN(n10651) );
  OR2_X1 U10673 ( .A1(n10434), .A2(n10435), .ZN(n10649) );
  AND2_X1 U10674 ( .A1(n10652), .A2(n10653), .ZN(n10435) );
  NAND2_X1 U10675 ( .A1(n10432), .A2(n10654), .ZN(n10653) );
  OR2_X1 U10676 ( .A1(n10430), .A2(n10431), .ZN(n10654) );
  NOR2_X1 U10677 ( .A1(n10207), .A2(n7923), .ZN(n10432) );
  NAND2_X1 U10678 ( .A1(n10430), .A2(n10431), .ZN(n10652) );
  NAND2_X1 U10679 ( .A1(n10427), .A2(n10655), .ZN(n10431) );
  NAND2_X1 U10680 ( .A1(n10426), .A2(n10428), .ZN(n10655) );
  NAND2_X1 U10681 ( .A1(n10656), .A2(n10657), .ZN(n10428) );
  NAND2_X1 U10682 ( .A1(b_18_), .A2(a_26_), .ZN(n10657) );
  INV_X1 U10683 ( .A(n10658), .ZN(n10656) );
  XNOR2_X1 U10684 ( .A(n10659), .B(n10660), .ZN(n10426) );
  NAND2_X1 U10685 ( .A1(n10661), .A2(n10662), .ZN(n10659) );
  NAND2_X1 U10686 ( .A1(a_26_), .A2(n10658), .ZN(n10427) );
  NAND2_X1 U10687 ( .A1(n10398), .A2(n10663), .ZN(n10658) );
  NAND2_X1 U10688 ( .A1(n10397), .A2(n10399), .ZN(n10663) );
  NAND2_X1 U10689 ( .A1(n10664), .A2(n10665), .ZN(n10399) );
  NAND2_X1 U10690 ( .A1(b_18_), .A2(a_27_), .ZN(n10665) );
  INV_X1 U10691 ( .A(n10666), .ZN(n10664) );
  XNOR2_X1 U10692 ( .A(n10667), .B(n10668), .ZN(n10397) );
  XOR2_X1 U10693 ( .A(n10669), .B(n10670), .Z(n10667) );
  NAND2_X1 U10694 ( .A1(b_17_), .A2(a_28_), .ZN(n10669) );
  NAND2_X1 U10695 ( .A1(a_27_), .A2(n10666), .ZN(n10398) );
  NAND2_X1 U10696 ( .A1(n10671), .A2(n10672), .ZN(n10666) );
  NAND3_X1 U10697 ( .A1(a_28_), .A2(n10673), .A3(b_18_), .ZN(n10672) );
  NAND2_X1 U10698 ( .A1(n10407), .A2(n10405), .ZN(n10673) );
  OR2_X1 U10699 ( .A1(n10405), .A2(n10407), .ZN(n10671) );
  AND2_X1 U10700 ( .A1(n10674), .A2(n10675), .ZN(n10407) );
  NAND2_X1 U10701 ( .A1(n10422), .A2(n10676), .ZN(n10675) );
  OR2_X1 U10702 ( .A1(n10423), .A2(n10424), .ZN(n10676) );
  NOR2_X1 U10703 ( .A1(n10207), .A2(n7946), .ZN(n10422) );
  NAND2_X1 U10704 ( .A1(n10424), .A2(n10423), .ZN(n10674) );
  NAND2_X1 U10705 ( .A1(n10677), .A2(n10678), .ZN(n10423) );
  NAND2_X1 U10706 ( .A1(b_16_), .A2(n10679), .ZN(n10678) );
  NAND2_X1 U10707 ( .A1(n7268), .A2(n10680), .ZN(n10679) );
  NAND2_X1 U10708 ( .A1(a_31_), .A2(n10420), .ZN(n10680) );
  NAND2_X1 U10709 ( .A1(b_17_), .A2(n10681), .ZN(n10677) );
  NAND2_X1 U10710 ( .A1(n7272), .A2(n10682), .ZN(n10681) );
  NAND2_X1 U10711 ( .A1(a_30_), .A2(n10683), .ZN(n10682) );
  AND3_X1 U10712 ( .A1(b_17_), .A2(n7954), .A3(b_18_), .ZN(n10424) );
  XNOR2_X1 U10713 ( .A(n10684), .B(n10685), .ZN(n10405) );
  XOR2_X1 U10714 ( .A(n10686), .B(n10687), .Z(n10684) );
  XNOR2_X1 U10715 ( .A(n10688), .B(n10689), .ZN(n10430) );
  NAND2_X1 U10716 ( .A1(n10690), .A2(n10691), .ZN(n10688) );
  XNOR2_X1 U10717 ( .A(n10692), .B(n10693), .ZN(n10434) );
  XOR2_X1 U10718 ( .A(n10694), .B(n10695), .Z(n10692) );
  XNOR2_X1 U10719 ( .A(n10696), .B(n10697), .ZN(n10437) );
  XNOR2_X1 U10720 ( .A(n10698), .B(n10699), .ZN(n10696) );
  NOR2_X1 U10721 ( .A1(n7691), .A2(n10420), .ZN(n10699) );
  XNOR2_X1 U10722 ( .A(n10700), .B(n10701), .ZN(n10446) );
  XOR2_X1 U10723 ( .A(n10702), .B(n10703), .Z(n10701) );
  NAND2_X1 U10724 ( .A1(b_17_), .A2(a_22_), .ZN(n10703) );
  XNOR2_X1 U10725 ( .A(n10704), .B(n10705), .ZN(n10450) );
  XOR2_X1 U10726 ( .A(n10706), .B(n10707), .Z(n10704) );
  XNOR2_X1 U10727 ( .A(n10708), .B(n10709), .ZN(n10453) );
  XNOR2_X1 U10728 ( .A(n10710), .B(n10711), .ZN(n10708) );
  NOR2_X1 U10729 ( .A1(n7987), .A2(n10420), .ZN(n10711) );
  XOR2_X1 U10730 ( .A(n10712), .B(n10713), .Z(n10458) );
  XNOR2_X1 U10731 ( .A(n10714), .B(n10715), .ZN(n10713) );
  XNOR2_X1 U10732 ( .A(n10716), .B(n10717), .ZN(n10462) );
  XNOR2_X1 U10733 ( .A(n10718), .B(n10719), .ZN(n10716) );
  NOR2_X1 U10734 ( .A1(n7764), .A2(n10420), .ZN(n10719) );
  XOR2_X1 U10735 ( .A(n10720), .B(n10721), .Z(n10465) );
  XOR2_X1 U10736 ( .A(n10722), .B(n10723), .Z(n10720) );
  XNOR2_X1 U10737 ( .A(n10724), .B(n10725), .ZN(n10469) );
  XOR2_X1 U10738 ( .A(n10726), .B(n10727), .Z(n10725) );
  NAND2_X1 U10739 ( .A1(b_17_), .A2(a_16_), .ZN(n10727) );
  XOR2_X1 U10740 ( .A(n10728), .B(n10729), .Z(n10474) );
  XNOR2_X1 U10741 ( .A(n10730), .B(n10731), .ZN(n10729) );
  XNOR2_X1 U10742 ( .A(n10732), .B(n10733), .ZN(n10478) );
  XOR2_X1 U10743 ( .A(n10734), .B(n10735), .Z(n10732) );
  XNOR2_X1 U10744 ( .A(n10736), .B(n10737), .ZN(n10481) );
  XOR2_X1 U10745 ( .A(n10738), .B(n10739), .Z(n10736) );
  NAND2_X1 U10746 ( .A1(b_17_), .A2(a_13_), .ZN(n10738) );
  XOR2_X1 U10747 ( .A(n10740), .B(n10741), .Z(n10344) );
  XOR2_X1 U10748 ( .A(n10742), .B(n10743), .Z(n10741) );
  NAND2_X1 U10749 ( .A1(b_17_), .A2(a_12_), .ZN(n10743) );
  XOR2_X1 U10750 ( .A(n10744), .B(n10745), .Z(n10486) );
  XOR2_X1 U10751 ( .A(n10746), .B(n10747), .Z(n10745) );
  NAND2_X1 U10752 ( .A1(b_17_), .A2(a_11_), .ZN(n10747) );
  XNOR2_X1 U10753 ( .A(n10748), .B(n10749), .ZN(n10521) );
  XOR2_X1 U10754 ( .A(n10750), .B(n10751), .Z(n10749) );
  NAND2_X1 U10755 ( .A1(b_17_), .A2(a_2_), .ZN(n10751) );
  XNOR2_X1 U10756 ( .A(n10752), .B(n10753), .ZN(n10306) );
  XOR2_X1 U10757 ( .A(n10754), .B(n10755), .Z(n10753) );
  NAND2_X1 U10758 ( .A1(b_17_), .A2(a_1_), .ZN(n10755) );
  XOR2_X1 U10759 ( .A(n7547), .B(n7546), .Z(n10527) );
  NAND3_X1 U10760 ( .A1(n7546), .A2(n7547), .A3(n10756), .ZN(n7484) );
  XOR2_X1 U10761 ( .A(n7549), .B(n7548), .Z(n10756) );
  NAND2_X1 U10762 ( .A1(n10757), .A2(n10758), .ZN(n7547) );
  NAND3_X1 U10763 ( .A1(a_0_), .A2(n10759), .A3(b_17_), .ZN(n10758) );
  OR2_X1 U10764 ( .A1(n10530), .A2(n10528), .ZN(n10759) );
  NAND2_X1 U10765 ( .A1(n10528), .A2(n10530), .ZN(n10757) );
  NAND2_X1 U10766 ( .A1(n10760), .A2(n10761), .ZN(n10530) );
  NAND3_X1 U10767 ( .A1(a_1_), .A2(n10762), .A3(b_17_), .ZN(n10761) );
  OR2_X1 U10768 ( .A1(n10754), .A2(n10752), .ZN(n10762) );
  NAND2_X1 U10769 ( .A1(n10752), .A2(n10754), .ZN(n10760) );
  NAND2_X1 U10770 ( .A1(n10763), .A2(n10764), .ZN(n10754) );
  NAND3_X1 U10771 ( .A1(a_2_), .A2(n10765), .A3(b_17_), .ZN(n10764) );
  OR2_X1 U10772 ( .A1(n10750), .A2(n10748), .ZN(n10765) );
  NAND2_X1 U10773 ( .A1(n10748), .A2(n10750), .ZN(n10763) );
  NAND2_X1 U10774 ( .A1(n10766), .A2(n10767), .ZN(n10750) );
  NAND3_X1 U10775 ( .A1(a_3_), .A2(n10768), .A3(b_17_), .ZN(n10767) );
  OR2_X1 U10776 ( .A1(n10544), .A2(n10543), .ZN(n10768) );
  NAND2_X1 U10777 ( .A1(n10543), .A2(n10544), .ZN(n10766) );
  NAND2_X1 U10778 ( .A1(n10769), .A2(n10770), .ZN(n10544) );
  NAND3_X1 U10779 ( .A1(a_4_), .A2(n10771), .A3(b_17_), .ZN(n10770) );
  OR2_X1 U10780 ( .A1(n10552), .A2(n10550), .ZN(n10771) );
  NAND2_X1 U10781 ( .A1(n10550), .A2(n10552), .ZN(n10769) );
  NAND2_X1 U10782 ( .A1(n10772), .A2(n10773), .ZN(n10552) );
  NAND3_X1 U10783 ( .A1(a_5_), .A2(n10774), .A3(b_17_), .ZN(n10773) );
  OR2_X1 U10784 ( .A1(n10560), .A2(n10559), .ZN(n10774) );
  NAND2_X1 U10785 ( .A1(n10559), .A2(n10560), .ZN(n10772) );
  NAND2_X1 U10786 ( .A1(n10775), .A2(n10776), .ZN(n10560) );
  NAND3_X1 U10787 ( .A1(a_6_), .A2(n10777), .A3(b_17_), .ZN(n10776) );
  OR2_X1 U10788 ( .A1(n10568), .A2(n10566), .ZN(n10777) );
  NAND2_X1 U10789 ( .A1(n10566), .A2(n10568), .ZN(n10775) );
  NAND2_X1 U10790 ( .A1(n10778), .A2(n10779), .ZN(n10568) );
  NAND3_X1 U10791 ( .A1(a_7_), .A2(n10780), .A3(b_17_), .ZN(n10779) );
  OR2_X1 U10792 ( .A1(n10576), .A2(n10574), .ZN(n10780) );
  NAND2_X1 U10793 ( .A1(n10574), .A2(n10576), .ZN(n10778) );
  NAND2_X1 U10794 ( .A1(n10781), .A2(n10782), .ZN(n10576) );
  NAND3_X1 U10795 ( .A1(a_8_), .A2(n10783), .A3(b_17_), .ZN(n10782) );
  OR2_X1 U10796 ( .A1(n10584), .A2(n10582), .ZN(n10783) );
  NAND2_X1 U10797 ( .A1(n10582), .A2(n10584), .ZN(n10781) );
  NAND2_X1 U10798 ( .A1(n10784), .A2(n10785), .ZN(n10584) );
  NAND3_X1 U10799 ( .A1(a_9_), .A2(n10786), .A3(b_17_), .ZN(n10785) );
  NAND2_X1 U10800 ( .A1(n10592), .A2(n10591), .ZN(n10786) );
  OR2_X1 U10801 ( .A1(n10591), .A2(n10592), .ZN(n10784) );
  AND2_X1 U10802 ( .A1(n10787), .A2(n10788), .ZN(n10592) );
  NAND3_X1 U10803 ( .A1(a_10_), .A2(n10789), .A3(b_17_), .ZN(n10788) );
  NAND2_X1 U10804 ( .A1(n10600), .A2(n10599), .ZN(n10789) );
  OR2_X1 U10805 ( .A1(n10599), .A2(n10600), .ZN(n10787) );
  AND2_X1 U10806 ( .A1(n10790), .A2(n10791), .ZN(n10600) );
  NAND3_X1 U10807 ( .A1(a_11_), .A2(n10792), .A3(b_17_), .ZN(n10791) );
  OR2_X1 U10808 ( .A1(n10746), .A2(n10744), .ZN(n10792) );
  NAND2_X1 U10809 ( .A1(n10744), .A2(n10746), .ZN(n10790) );
  NAND2_X1 U10810 ( .A1(n10793), .A2(n10794), .ZN(n10746) );
  NAND3_X1 U10811 ( .A1(a_12_), .A2(n10795), .A3(b_17_), .ZN(n10794) );
  OR2_X1 U10812 ( .A1(n10742), .A2(n10740), .ZN(n10795) );
  NAND2_X1 U10813 ( .A1(n10740), .A2(n10742), .ZN(n10793) );
  NAND2_X1 U10814 ( .A1(n10796), .A2(n10797), .ZN(n10742) );
  NAND3_X1 U10815 ( .A1(a_13_), .A2(n10798), .A3(b_17_), .ZN(n10797) );
  NAND2_X1 U10816 ( .A1(n10739), .A2(n10737), .ZN(n10798) );
  OR2_X1 U10817 ( .A1(n10737), .A2(n10739), .ZN(n10796) );
  AND2_X1 U10818 ( .A1(n10799), .A2(n10800), .ZN(n10739) );
  NAND2_X1 U10819 ( .A1(n10735), .A2(n10801), .ZN(n10800) );
  OR2_X1 U10820 ( .A1(n10734), .A2(n10733), .ZN(n10801) );
  NOR2_X1 U10821 ( .A1(n10420), .A2(n7782), .ZN(n10735) );
  NAND2_X1 U10822 ( .A1(n10733), .A2(n10734), .ZN(n10799) );
  NAND2_X1 U10823 ( .A1(n10802), .A2(n10803), .ZN(n10734) );
  NAND2_X1 U10824 ( .A1(n10731), .A2(n10804), .ZN(n10803) );
  OR2_X1 U10825 ( .A1(n10730), .A2(n10728), .ZN(n10804) );
  NOR2_X1 U10826 ( .A1(n10420), .A2(n7346), .ZN(n10731) );
  NAND2_X1 U10827 ( .A1(n10728), .A2(n10730), .ZN(n10802) );
  NAND2_X1 U10828 ( .A1(n10805), .A2(n10806), .ZN(n10730) );
  NAND3_X1 U10829 ( .A1(a_16_), .A2(n10807), .A3(b_17_), .ZN(n10806) );
  OR2_X1 U10830 ( .A1(n10726), .A2(n10724), .ZN(n10807) );
  NAND2_X1 U10831 ( .A1(n10724), .A2(n10726), .ZN(n10805) );
  NAND2_X1 U10832 ( .A1(n10808), .A2(n10809), .ZN(n10726) );
  NAND2_X1 U10833 ( .A1(n10723), .A2(n10810), .ZN(n10809) );
  OR2_X1 U10834 ( .A1(n10722), .A2(n10721), .ZN(n10810) );
  NAND2_X1 U10835 ( .A1(n10721), .A2(n10722), .ZN(n10808) );
  NAND2_X1 U10836 ( .A1(n10811), .A2(n10812), .ZN(n10722) );
  NAND3_X1 U10837 ( .A1(a_18_), .A2(n10813), .A3(b_17_), .ZN(n10812) );
  NAND2_X1 U10838 ( .A1(n10718), .A2(n10717), .ZN(n10813) );
  OR2_X1 U10839 ( .A1(n10717), .A2(n10718), .ZN(n10811) );
  AND2_X1 U10840 ( .A1(n10814), .A2(n10815), .ZN(n10718) );
  NAND2_X1 U10841 ( .A1(n10715), .A2(n10816), .ZN(n10815) );
  OR2_X1 U10842 ( .A1(n10714), .A2(n10712), .ZN(n10816) );
  NOR2_X1 U10843 ( .A1(n10420), .A2(n7902), .ZN(n10715) );
  NAND2_X1 U10844 ( .A1(n10712), .A2(n10714), .ZN(n10814) );
  NAND2_X1 U10845 ( .A1(n10817), .A2(n10818), .ZN(n10714) );
  NAND3_X1 U10846 ( .A1(a_20_), .A2(n10819), .A3(b_17_), .ZN(n10818) );
  NAND2_X1 U10847 ( .A1(n10710), .A2(n10709), .ZN(n10819) );
  OR2_X1 U10848 ( .A1(n10709), .A2(n10710), .ZN(n10817) );
  AND2_X1 U10849 ( .A1(n10820), .A2(n10821), .ZN(n10710) );
  NAND2_X1 U10850 ( .A1(n10707), .A2(n10822), .ZN(n10821) );
  OR2_X1 U10851 ( .A1(n10706), .A2(n10705), .ZN(n10822) );
  NOR2_X1 U10852 ( .A1(n10420), .A2(n7909), .ZN(n10707) );
  NAND2_X1 U10853 ( .A1(n10705), .A2(n10706), .ZN(n10820) );
  NAND2_X1 U10854 ( .A1(n10823), .A2(n10824), .ZN(n10706) );
  NAND3_X1 U10855 ( .A1(a_22_), .A2(n10825), .A3(b_17_), .ZN(n10824) );
  OR2_X1 U10856 ( .A1(n10702), .A2(n10700), .ZN(n10825) );
  NAND2_X1 U10857 ( .A1(n10700), .A2(n10702), .ZN(n10823) );
  NAND2_X1 U10858 ( .A1(n10826), .A2(n10827), .ZN(n10702) );
  NAND2_X1 U10859 ( .A1(n10645), .A2(n10828), .ZN(n10827) );
  OR2_X1 U10860 ( .A1(n10644), .A2(n10642), .ZN(n10828) );
  NOR2_X1 U10861 ( .A1(n10420), .A2(n7916), .ZN(n10645) );
  NAND2_X1 U10862 ( .A1(n10642), .A2(n10644), .ZN(n10826) );
  NAND2_X1 U10863 ( .A1(n10829), .A2(n10830), .ZN(n10644) );
  NAND3_X1 U10864 ( .A1(a_24_), .A2(n10831), .A3(b_17_), .ZN(n10830) );
  NAND2_X1 U10865 ( .A1(n10698), .A2(n10697), .ZN(n10831) );
  OR2_X1 U10866 ( .A1(n10697), .A2(n10698), .ZN(n10829) );
  AND2_X1 U10867 ( .A1(n10832), .A2(n10833), .ZN(n10698) );
  NAND2_X1 U10868 ( .A1(n10695), .A2(n10834), .ZN(n10833) );
  OR2_X1 U10869 ( .A1(n10694), .A2(n10693), .ZN(n10834) );
  NOR2_X1 U10870 ( .A1(n10420), .A2(n7923), .ZN(n10695) );
  NAND2_X1 U10871 ( .A1(n10693), .A2(n10694), .ZN(n10832) );
  NAND2_X1 U10872 ( .A1(n10690), .A2(n10835), .ZN(n10694) );
  NAND2_X1 U10873 ( .A1(n10689), .A2(n10691), .ZN(n10835) );
  NAND2_X1 U10874 ( .A1(n10836), .A2(n10837), .ZN(n10691) );
  NAND2_X1 U10875 ( .A1(b_17_), .A2(a_26_), .ZN(n10837) );
  INV_X1 U10876 ( .A(n10838), .ZN(n10836) );
  XNOR2_X1 U10877 ( .A(n10839), .B(n10840), .ZN(n10689) );
  NAND2_X1 U10878 ( .A1(n10841), .A2(n10842), .ZN(n10839) );
  NAND2_X1 U10879 ( .A1(a_26_), .A2(n10838), .ZN(n10690) );
  NAND2_X1 U10880 ( .A1(n10661), .A2(n10843), .ZN(n10838) );
  NAND2_X1 U10881 ( .A1(n10660), .A2(n10662), .ZN(n10843) );
  NAND2_X1 U10882 ( .A1(n10844), .A2(n10845), .ZN(n10662) );
  NAND2_X1 U10883 ( .A1(b_17_), .A2(a_27_), .ZN(n10845) );
  INV_X1 U10884 ( .A(n10846), .ZN(n10844) );
  XNOR2_X1 U10885 ( .A(n10847), .B(n10848), .ZN(n10660) );
  XOR2_X1 U10886 ( .A(n10849), .B(n10850), .Z(n10847) );
  NAND2_X1 U10887 ( .A1(b_16_), .A2(a_28_), .ZN(n10849) );
  NAND2_X1 U10888 ( .A1(a_27_), .A2(n10846), .ZN(n10661) );
  NAND2_X1 U10889 ( .A1(n10851), .A2(n10852), .ZN(n10846) );
  NAND3_X1 U10890 ( .A1(a_28_), .A2(n10853), .A3(b_17_), .ZN(n10852) );
  NAND2_X1 U10891 ( .A1(n10670), .A2(n10668), .ZN(n10853) );
  OR2_X1 U10892 ( .A1(n10668), .A2(n10670), .ZN(n10851) );
  AND2_X1 U10893 ( .A1(n10854), .A2(n10855), .ZN(n10670) );
  NAND2_X1 U10894 ( .A1(n10685), .A2(n10856), .ZN(n10855) );
  OR2_X1 U10895 ( .A1(n10686), .A2(n10687), .ZN(n10856) );
  NOR2_X1 U10896 ( .A1(n10420), .A2(n7946), .ZN(n10685) );
  NAND2_X1 U10897 ( .A1(n10687), .A2(n10686), .ZN(n10854) );
  NAND2_X1 U10898 ( .A1(n10857), .A2(n10858), .ZN(n10686) );
  NAND2_X1 U10899 ( .A1(b_15_), .A2(n10859), .ZN(n10858) );
  NAND2_X1 U10900 ( .A1(n7268), .A2(n10860), .ZN(n10859) );
  NAND2_X1 U10901 ( .A1(a_31_), .A2(n10683), .ZN(n10860) );
  NAND2_X1 U10902 ( .A1(b_16_), .A2(n10861), .ZN(n10857) );
  NAND2_X1 U10903 ( .A1(n7272), .A2(n10862), .ZN(n10861) );
  NAND2_X1 U10904 ( .A1(a_30_), .A2(n10863), .ZN(n10862) );
  AND3_X1 U10905 ( .A1(b_17_), .A2(n7954), .A3(b_16_), .ZN(n10687) );
  XNOR2_X1 U10906 ( .A(n10864), .B(n10865), .ZN(n10668) );
  XOR2_X1 U10907 ( .A(n10866), .B(n10867), .Z(n10864) );
  XNOR2_X1 U10908 ( .A(n10868), .B(n10869), .ZN(n10693) );
  NAND2_X1 U10909 ( .A1(n10870), .A2(n10871), .ZN(n10868) );
  XNOR2_X1 U10910 ( .A(n10872), .B(n10873), .ZN(n10697) );
  XOR2_X1 U10911 ( .A(n10874), .B(n10875), .Z(n10872) );
  XNOR2_X1 U10912 ( .A(n10876), .B(n10877), .ZN(n10642) );
  XNOR2_X1 U10913 ( .A(n10878), .B(n10879), .ZN(n10876) );
  NOR2_X1 U10914 ( .A1(n7691), .A2(n10683), .ZN(n10879) );
  XNOR2_X1 U10915 ( .A(n10880), .B(n10881), .ZN(n10700) );
  XNOR2_X1 U10916 ( .A(n10882), .B(n10883), .ZN(n10881) );
  XNOR2_X1 U10917 ( .A(n10884), .B(n10885), .ZN(n10705) );
  XNOR2_X1 U10918 ( .A(n10886), .B(n10887), .ZN(n10884) );
  NOR2_X1 U10919 ( .A1(n7312), .A2(n10683), .ZN(n10887) );
  XNOR2_X1 U10920 ( .A(n10888), .B(n10889), .ZN(n10709) );
  XOR2_X1 U10921 ( .A(n10890), .B(n10891), .Z(n10888) );
  XNOR2_X1 U10922 ( .A(n10892), .B(n10893), .ZN(n10712) );
  XNOR2_X1 U10923 ( .A(n10894), .B(n10895), .ZN(n10892) );
  NOR2_X1 U10924 ( .A1(n7987), .A2(n10683), .ZN(n10895) );
  XOR2_X1 U10925 ( .A(n10896), .B(n10897), .Z(n10717) );
  XNOR2_X1 U10926 ( .A(n10898), .B(n10899), .ZN(n10897) );
  XNOR2_X1 U10927 ( .A(n10900), .B(n10901), .ZN(n10721) );
  XNOR2_X1 U10928 ( .A(n10902), .B(n10903), .ZN(n10900) );
  NOR2_X1 U10929 ( .A1(n7764), .A2(n10683), .ZN(n10903) );
  XOR2_X1 U10930 ( .A(n10904), .B(n10905), .Z(n10724) );
  XOR2_X1 U10931 ( .A(n10906), .B(n10907), .Z(n10904) );
  XNOR2_X1 U10932 ( .A(n10908), .B(n10909), .ZN(n10728) );
  XNOR2_X1 U10933 ( .A(n10910), .B(n10911), .ZN(n10909) );
  XNOR2_X1 U10934 ( .A(n10912), .B(n10913), .ZN(n10733) );
  NAND2_X1 U10935 ( .A1(n10914), .A2(n10915), .ZN(n10912) );
  XNOR2_X1 U10936 ( .A(n10916), .B(n10917), .ZN(n10737) );
  XOR2_X1 U10937 ( .A(n10918), .B(n10919), .Z(n10916) );
  XNOR2_X1 U10938 ( .A(n10920), .B(n10921), .ZN(n10740) );
  XNOR2_X1 U10939 ( .A(n10922), .B(n10923), .ZN(n10920) );
  XNOR2_X1 U10940 ( .A(n10924), .B(n10925), .ZN(n10744) );
  XNOR2_X1 U10941 ( .A(n10926), .B(n10927), .ZN(n10924) );
  XNOR2_X1 U10942 ( .A(n10928), .B(n10929), .ZN(n10599) );
  XOR2_X1 U10943 ( .A(n10930), .B(n10931), .Z(n10928) );
  XNOR2_X1 U10944 ( .A(n10932), .B(n10933), .ZN(n10591) );
  XOR2_X1 U10945 ( .A(n10934), .B(n10935), .Z(n10932) );
  XNOR2_X1 U10946 ( .A(n10936), .B(n10937), .ZN(n10582) );
  XNOR2_X1 U10947 ( .A(n10938), .B(n10939), .ZN(n10937) );
  XNOR2_X1 U10948 ( .A(n10940), .B(n10941), .ZN(n10574) );
  XNOR2_X1 U10949 ( .A(n10942), .B(n10943), .ZN(n10940) );
  NOR2_X1 U10950 ( .A1(n8037), .A2(n10683), .ZN(n10943) );
  XNOR2_X1 U10951 ( .A(n10944), .B(n10945), .ZN(n10566) );
  XNOR2_X1 U10952 ( .A(n10946), .B(n10947), .ZN(n10945) );
  XNOR2_X1 U10953 ( .A(n10948), .B(n10949), .ZN(n10559) );
  XNOR2_X1 U10954 ( .A(n10950), .B(n10951), .ZN(n10948) );
  NOR2_X1 U10955 ( .A1(n7388), .A2(n10683), .ZN(n10951) );
  XNOR2_X1 U10956 ( .A(n10952), .B(n10953), .ZN(n10550) );
  NAND2_X1 U10957 ( .A1(n10954), .A2(n10955), .ZN(n10952) );
  XNOR2_X1 U10958 ( .A(n10956), .B(n10957), .ZN(n10543) );
  XNOR2_X1 U10959 ( .A(n10958), .B(n10959), .ZN(n10956) );
  XOR2_X1 U10960 ( .A(n10960), .B(n10961), .Z(n10748) );
  XOR2_X1 U10961 ( .A(n10962), .B(n10963), .Z(n10960) );
  XOR2_X1 U10962 ( .A(n10964), .B(n10965), .Z(n10752) );
  XOR2_X1 U10963 ( .A(n10966), .B(n10967), .Z(n10964) );
  XNOR2_X1 U10964 ( .A(n10968), .B(n10969), .ZN(n10528) );
  XNOR2_X1 U10965 ( .A(n10970), .B(n10971), .ZN(n10968) );
  NOR2_X1 U10966 ( .A1(n7411), .A2(n10683), .ZN(n10971) );
  XNOR2_X1 U10967 ( .A(n10972), .B(n10973), .ZN(n7546) );
  NAND2_X1 U10968 ( .A1(n10974), .A2(n10975), .ZN(n10972) );
  NAND2_X1 U10969 ( .A1(n10976), .A2(n10977), .ZN(n7487) );
  NAND2_X1 U10970 ( .A1(n7549), .A2(n7548), .ZN(n10977) );
  XOR2_X1 U10971 ( .A(n10978), .B(n10979), .Z(n10976) );
  NAND3_X1 U10972 ( .A1(n7549), .A2(n7548), .A3(n10980), .ZN(n7488) );
  XOR2_X1 U10973 ( .A(n10981), .B(n10978), .Z(n10980) );
  NAND2_X1 U10974 ( .A1(n10974), .A2(n10982), .ZN(n7548) );
  NAND2_X1 U10975 ( .A1(n10973), .A2(n10975), .ZN(n10982) );
  NAND2_X1 U10976 ( .A1(n10983), .A2(n10984), .ZN(n10975) );
  NAND2_X1 U10977 ( .A1(b_16_), .A2(a_0_), .ZN(n10984) );
  INV_X1 U10978 ( .A(n10985), .ZN(n10983) );
  XOR2_X1 U10979 ( .A(n10986), .B(n10987), .Z(n10973) );
  XOR2_X1 U10980 ( .A(n10988), .B(n10989), .Z(n10986) );
  NOR2_X1 U10981 ( .A1(n7411), .A2(n10863), .ZN(n10989) );
  NAND2_X1 U10982 ( .A1(a_0_), .A2(n10985), .ZN(n10974) );
  NAND2_X1 U10983 ( .A1(n10990), .A2(n10991), .ZN(n10985) );
  NAND3_X1 U10984 ( .A1(a_1_), .A2(n10992), .A3(b_16_), .ZN(n10991) );
  NAND2_X1 U10985 ( .A1(n10970), .A2(n10969), .ZN(n10992) );
  OR2_X1 U10986 ( .A1(n10969), .A2(n10970), .ZN(n10990) );
  AND2_X1 U10987 ( .A1(n10993), .A2(n10994), .ZN(n10970) );
  NAND2_X1 U10988 ( .A1(n10967), .A2(n10995), .ZN(n10994) );
  OR2_X1 U10989 ( .A1(n10965), .A2(n10966), .ZN(n10995) );
  NOR2_X1 U10990 ( .A1(n10683), .A2(n7832), .ZN(n10967) );
  NAND2_X1 U10991 ( .A1(n10965), .A2(n10966), .ZN(n10993) );
  NAND2_X1 U10992 ( .A1(n10996), .A2(n10997), .ZN(n10966) );
  NAND2_X1 U10993 ( .A1(n10963), .A2(n10998), .ZN(n10997) );
  OR2_X1 U10994 ( .A1(n10961), .A2(n10962), .ZN(n10998) );
  NOR2_X1 U10995 ( .A1(n10683), .A2(n7850), .ZN(n10963) );
  NAND2_X1 U10996 ( .A1(n10961), .A2(n10962), .ZN(n10996) );
  NAND2_X1 U10997 ( .A1(n10999), .A2(n11000), .ZN(n10962) );
  NAND2_X1 U10998 ( .A1(n10959), .A2(n11001), .ZN(n11000) );
  NAND2_X1 U10999 ( .A1(n10958), .A2(n10957), .ZN(n11001) );
  NOR2_X1 U11000 ( .A1(n10683), .A2(n7398), .ZN(n10959) );
  OR2_X1 U11001 ( .A1(n10957), .A2(n10958), .ZN(n10999) );
  AND2_X1 U11002 ( .A1(n10954), .A2(n11002), .ZN(n10958) );
  NAND2_X1 U11003 ( .A1(n10953), .A2(n10955), .ZN(n11002) );
  NAND2_X1 U11004 ( .A1(n11003), .A2(n11004), .ZN(n10955) );
  NAND2_X1 U11005 ( .A1(b_16_), .A2(a_5_), .ZN(n11004) );
  INV_X1 U11006 ( .A(n11005), .ZN(n11003) );
  XOR2_X1 U11007 ( .A(n11006), .B(n11007), .Z(n10953) );
  XOR2_X1 U11008 ( .A(n11008), .B(n11009), .Z(n11006) );
  NOR2_X1 U11009 ( .A1(n7388), .A2(n10863), .ZN(n11009) );
  NAND2_X1 U11010 ( .A1(a_5_), .A2(n11005), .ZN(n10954) );
  NAND2_X1 U11011 ( .A1(n11010), .A2(n11011), .ZN(n11005) );
  NAND3_X1 U11012 ( .A1(a_6_), .A2(n11012), .A3(b_16_), .ZN(n11011) );
  NAND2_X1 U11013 ( .A1(n10950), .A2(n10949), .ZN(n11012) );
  OR2_X1 U11014 ( .A1(n10949), .A2(n10950), .ZN(n11010) );
  AND2_X1 U11015 ( .A1(n11013), .A2(n11014), .ZN(n10950) );
  NAND2_X1 U11016 ( .A1(n10947), .A2(n11015), .ZN(n11014) );
  OR2_X1 U11017 ( .A1(n10944), .A2(n10946), .ZN(n11015) );
  NOR2_X1 U11018 ( .A1(n10683), .A2(n7863), .ZN(n10947) );
  NAND2_X1 U11019 ( .A1(n10944), .A2(n10946), .ZN(n11013) );
  NAND2_X1 U11020 ( .A1(n11016), .A2(n11017), .ZN(n10946) );
  NAND3_X1 U11021 ( .A1(a_8_), .A2(n11018), .A3(b_16_), .ZN(n11017) );
  NAND2_X1 U11022 ( .A1(n10942), .A2(n10941), .ZN(n11018) );
  OR2_X1 U11023 ( .A1(n10941), .A2(n10942), .ZN(n11016) );
  AND2_X1 U11024 ( .A1(n11019), .A2(n11020), .ZN(n10942) );
  NAND2_X1 U11025 ( .A1(n10939), .A2(n11021), .ZN(n11020) );
  OR2_X1 U11026 ( .A1(n10938), .A2(n10936), .ZN(n11021) );
  NOR2_X1 U11027 ( .A1(n10683), .A2(n7870), .ZN(n10939) );
  NAND2_X1 U11028 ( .A1(n10936), .A2(n10938), .ZN(n11019) );
  NAND2_X1 U11029 ( .A1(n11022), .A2(n11023), .ZN(n10938) );
  NAND2_X1 U11030 ( .A1(n10935), .A2(n11024), .ZN(n11023) );
  OR2_X1 U11031 ( .A1(n10933), .A2(n10934), .ZN(n11024) );
  NOR2_X1 U11032 ( .A1(n10683), .A2(n7799), .ZN(n10935) );
  NAND2_X1 U11033 ( .A1(n10933), .A2(n10934), .ZN(n11022) );
  NAND2_X1 U11034 ( .A1(n11025), .A2(n11026), .ZN(n10934) );
  NAND2_X1 U11035 ( .A1(n10931), .A2(n11027), .ZN(n11026) );
  OR2_X1 U11036 ( .A1(n10929), .A2(n10930), .ZN(n11027) );
  NOR2_X1 U11037 ( .A1(n10683), .A2(n7877), .ZN(n10931) );
  NAND2_X1 U11038 ( .A1(n10929), .A2(n10930), .ZN(n11025) );
  NAND2_X1 U11039 ( .A1(n11028), .A2(n11029), .ZN(n10930) );
  NAND2_X1 U11040 ( .A1(n10927), .A2(n11030), .ZN(n11029) );
  NAND2_X1 U11041 ( .A1(n10926), .A2(n10925), .ZN(n11030) );
  NOR2_X1 U11042 ( .A1(n10683), .A2(n8020), .ZN(n10927) );
  OR2_X1 U11043 ( .A1(n10925), .A2(n10926), .ZN(n11028) );
  AND2_X1 U11044 ( .A1(n11031), .A2(n11032), .ZN(n10926) );
  NAND2_X1 U11045 ( .A1(n10923), .A2(n11033), .ZN(n11032) );
  NAND2_X1 U11046 ( .A1(n10922), .A2(n10921), .ZN(n11033) );
  NOR2_X1 U11047 ( .A1(n10683), .A2(n7355), .ZN(n10923) );
  OR2_X1 U11048 ( .A1(n10921), .A2(n10922), .ZN(n11031) );
  AND2_X1 U11049 ( .A1(n11034), .A2(n11035), .ZN(n10922) );
  NAND2_X1 U11050 ( .A1(n10918), .A2(n11036), .ZN(n11035) );
  OR2_X1 U11051 ( .A1(n10917), .A2(n10919), .ZN(n11036) );
  NOR2_X1 U11052 ( .A1(n10683), .A2(n7782), .ZN(n10918) );
  NAND2_X1 U11053 ( .A1(n10917), .A2(n10919), .ZN(n11034) );
  NAND2_X1 U11054 ( .A1(n10914), .A2(n11037), .ZN(n10919) );
  NAND2_X1 U11055 ( .A1(n10913), .A2(n10915), .ZN(n11037) );
  NAND2_X1 U11056 ( .A1(n11038), .A2(n11039), .ZN(n10915) );
  NAND2_X1 U11057 ( .A1(b_16_), .A2(a_15_), .ZN(n11039) );
  INV_X1 U11058 ( .A(n11040), .ZN(n11038) );
  XNOR2_X1 U11059 ( .A(n11041), .B(n11042), .ZN(n10913) );
  XOR2_X1 U11060 ( .A(n11043), .B(n11044), .Z(n11042) );
  NAND2_X1 U11061 ( .A1(b_15_), .A2(a_16_), .ZN(n11044) );
  NAND2_X1 U11062 ( .A1(a_15_), .A2(n11040), .ZN(n10914) );
  NAND2_X1 U11063 ( .A1(n11045), .A2(n11046), .ZN(n11040) );
  NAND2_X1 U11064 ( .A1(n10910), .A2(n11047), .ZN(n11046) );
  OR2_X1 U11065 ( .A1(n10911), .A2(n10908), .ZN(n11047) );
  NAND2_X1 U11066 ( .A1(n10908), .A2(n10911), .ZN(n11045) );
  NAND2_X1 U11067 ( .A1(n11048), .A2(n11049), .ZN(n10911) );
  NAND2_X1 U11068 ( .A1(n10907), .A2(n11050), .ZN(n11049) );
  OR2_X1 U11069 ( .A1(n10905), .A2(n10906), .ZN(n11050) );
  NOR2_X1 U11070 ( .A1(n10683), .A2(n7337), .ZN(n10907) );
  NAND2_X1 U11071 ( .A1(n10905), .A2(n10906), .ZN(n11048) );
  NAND2_X1 U11072 ( .A1(n11051), .A2(n11052), .ZN(n10906) );
  NAND3_X1 U11073 ( .A1(a_18_), .A2(n11053), .A3(b_16_), .ZN(n11052) );
  NAND2_X1 U11074 ( .A1(n10902), .A2(n10901), .ZN(n11053) );
  OR2_X1 U11075 ( .A1(n10901), .A2(n10902), .ZN(n11051) );
  AND2_X1 U11076 ( .A1(n11054), .A2(n11055), .ZN(n10902) );
  NAND2_X1 U11077 ( .A1(n10899), .A2(n11056), .ZN(n11055) );
  OR2_X1 U11078 ( .A1(n10896), .A2(n10898), .ZN(n11056) );
  NOR2_X1 U11079 ( .A1(n10683), .A2(n7902), .ZN(n10899) );
  NAND2_X1 U11080 ( .A1(n10896), .A2(n10898), .ZN(n11054) );
  NAND2_X1 U11081 ( .A1(n11057), .A2(n11058), .ZN(n10898) );
  NAND3_X1 U11082 ( .A1(a_20_), .A2(n11059), .A3(b_16_), .ZN(n11058) );
  NAND2_X1 U11083 ( .A1(n10894), .A2(n10893), .ZN(n11059) );
  OR2_X1 U11084 ( .A1(n10893), .A2(n10894), .ZN(n11057) );
  AND2_X1 U11085 ( .A1(n11060), .A2(n11061), .ZN(n10894) );
  NAND2_X1 U11086 ( .A1(n10891), .A2(n11062), .ZN(n11061) );
  OR2_X1 U11087 ( .A1(n10889), .A2(n10890), .ZN(n11062) );
  NOR2_X1 U11088 ( .A1(n10683), .A2(n7909), .ZN(n10891) );
  NAND2_X1 U11089 ( .A1(n10889), .A2(n10890), .ZN(n11060) );
  NAND2_X1 U11090 ( .A1(n11063), .A2(n11064), .ZN(n10890) );
  NAND3_X1 U11091 ( .A1(a_22_), .A2(n11065), .A3(b_16_), .ZN(n11064) );
  NAND2_X1 U11092 ( .A1(n10886), .A2(n10885), .ZN(n11065) );
  OR2_X1 U11093 ( .A1(n10885), .A2(n10886), .ZN(n11063) );
  AND2_X1 U11094 ( .A1(n11066), .A2(n11067), .ZN(n10886) );
  NAND2_X1 U11095 ( .A1(n10883), .A2(n11068), .ZN(n11067) );
  OR2_X1 U11096 ( .A1(n10880), .A2(n10882), .ZN(n11068) );
  NOR2_X1 U11097 ( .A1(n10683), .A2(n7916), .ZN(n10883) );
  NAND2_X1 U11098 ( .A1(n10880), .A2(n10882), .ZN(n11066) );
  NAND2_X1 U11099 ( .A1(n11069), .A2(n11070), .ZN(n10882) );
  NAND3_X1 U11100 ( .A1(a_24_), .A2(n11071), .A3(b_16_), .ZN(n11070) );
  NAND2_X1 U11101 ( .A1(n10878), .A2(n10877), .ZN(n11071) );
  OR2_X1 U11102 ( .A1(n10877), .A2(n10878), .ZN(n11069) );
  AND2_X1 U11103 ( .A1(n11072), .A2(n11073), .ZN(n10878) );
  NAND2_X1 U11104 ( .A1(n10875), .A2(n11074), .ZN(n11073) );
  OR2_X1 U11105 ( .A1(n10873), .A2(n10874), .ZN(n11074) );
  NOR2_X1 U11106 ( .A1(n10683), .A2(n7923), .ZN(n10875) );
  NAND2_X1 U11107 ( .A1(n10873), .A2(n10874), .ZN(n11072) );
  NAND2_X1 U11108 ( .A1(n10870), .A2(n11075), .ZN(n10874) );
  NAND2_X1 U11109 ( .A1(n10869), .A2(n10871), .ZN(n11075) );
  NAND2_X1 U11110 ( .A1(n11076), .A2(n11077), .ZN(n10871) );
  NAND2_X1 U11111 ( .A1(b_16_), .A2(a_26_), .ZN(n11077) );
  INV_X1 U11112 ( .A(n11078), .ZN(n11076) );
  XNOR2_X1 U11113 ( .A(n11079), .B(n11080), .ZN(n10869) );
  NAND2_X1 U11114 ( .A1(n11081), .A2(n11082), .ZN(n11079) );
  NAND2_X1 U11115 ( .A1(a_26_), .A2(n11078), .ZN(n10870) );
  NAND2_X1 U11116 ( .A1(n10841), .A2(n11083), .ZN(n11078) );
  NAND2_X1 U11117 ( .A1(n10840), .A2(n10842), .ZN(n11083) );
  NAND2_X1 U11118 ( .A1(n11084), .A2(n11085), .ZN(n10842) );
  NAND2_X1 U11119 ( .A1(b_16_), .A2(a_27_), .ZN(n11085) );
  INV_X1 U11120 ( .A(n11086), .ZN(n11084) );
  XNOR2_X1 U11121 ( .A(n11087), .B(n11088), .ZN(n10840) );
  XOR2_X1 U11122 ( .A(n11089), .B(n11090), .Z(n11087) );
  NAND2_X1 U11123 ( .A1(b_15_), .A2(a_28_), .ZN(n11089) );
  NAND2_X1 U11124 ( .A1(a_27_), .A2(n11086), .ZN(n10841) );
  NAND2_X1 U11125 ( .A1(n11091), .A2(n11092), .ZN(n11086) );
  NAND3_X1 U11126 ( .A1(a_28_), .A2(n11093), .A3(b_16_), .ZN(n11092) );
  NAND2_X1 U11127 ( .A1(n10850), .A2(n10848), .ZN(n11093) );
  OR2_X1 U11128 ( .A1(n10848), .A2(n10850), .ZN(n11091) );
  AND2_X1 U11129 ( .A1(n11094), .A2(n11095), .ZN(n10850) );
  NAND2_X1 U11130 ( .A1(n10865), .A2(n11096), .ZN(n11095) );
  OR2_X1 U11131 ( .A1(n10866), .A2(n10867), .ZN(n11096) );
  NOR2_X1 U11132 ( .A1(n10683), .A2(n7946), .ZN(n10865) );
  NAND2_X1 U11133 ( .A1(n10867), .A2(n10866), .ZN(n11094) );
  NAND2_X1 U11134 ( .A1(n11097), .A2(n11098), .ZN(n10866) );
  NAND2_X1 U11135 ( .A1(b_14_), .A2(n11099), .ZN(n11098) );
  NAND2_X1 U11136 ( .A1(n7268), .A2(n11100), .ZN(n11099) );
  NAND2_X1 U11137 ( .A1(a_31_), .A2(n10863), .ZN(n11100) );
  NAND2_X1 U11138 ( .A1(b_15_), .A2(n11101), .ZN(n11097) );
  NAND2_X1 U11139 ( .A1(n7272), .A2(n11102), .ZN(n11101) );
  NAND2_X1 U11140 ( .A1(a_30_), .A2(n11103), .ZN(n11102) );
  AND3_X1 U11141 ( .A1(b_16_), .A2(n7954), .A3(b_15_), .ZN(n10867) );
  XNOR2_X1 U11142 ( .A(n11104), .B(n11105), .ZN(n10848) );
  XOR2_X1 U11143 ( .A(n11106), .B(n11107), .Z(n11104) );
  XNOR2_X1 U11144 ( .A(n11108), .B(n11109), .ZN(n10873) );
  NAND2_X1 U11145 ( .A1(n11110), .A2(n11111), .ZN(n11108) );
  XNOR2_X1 U11146 ( .A(n11112), .B(n11113), .ZN(n10877) );
  XOR2_X1 U11147 ( .A(n11114), .B(n11115), .Z(n11112) );
  XNOR2_X1 U11148 ( .A(n11116), .B(n11117), .ZN(n10880) );
  XNOR2_X1 U11149 ( .A(n11118), .B(n11119), .ZN(n11116) );
  NOR2_X1 U11150 ( .A1(n7691), .A2(n10863), .ZN(n11119) );
  XOR2_X1 U11151 ( .A(n11120), .B(n11121), .Z(n10885) );
  XNOR2_X1 U11152 ( .A(n11122), .B(n11123), .ZN(n11121) );
  XNOR2_X1 U11153 ( .A(n11124), .B(n11125), .ZN(n10889) );
  XNOR2_X1 U11154 ( .A(n11126), .B(n11127), .ZN(n11124) );
  NOR2_X1 U11155 ( .A1(n7312), .A2(n10863), .ZN(n11127) );
  XNOR2_X1 U11156 ( .A(n11128), .B(n11129), .ZN(n10893) );
  XOR2_X1 U11157 ( .A(n11130), .B(n11131), .Z(n11128) );
  XNOR2_X1 U11158 ( .A(n11132), .B(n11133), .ZN(n10896) );
  XNOR2_X1 U11159 ( .A(n11134), .B(n11135), .ZN(n11132) );
  NOR2_X1 U11160 ( .A1(n7987), .A2(n10863), .ZN(n11135) );
  XOR2_X1 U11161 ( .A(n11136), .B(n11137), .Z(n10901) );
  XNOR2_X1 U11162 ( .A(n11138), .B(n11139), .ZN(n11137) );
  XNOR2_X1 U11163 ( .A(n11140), .B(n11141), .ZN(n10905) );
  XNOR2_X1 U11164 ( .A(n11142), .B(n11143), .ZN(n11140) );
  NOR2_X1 U11165 ( .A1(n7764), .A2(n10863), .ZN(n11143) );
  XOR2_X1 U11166 ( .A(n11144), .B(n11145), .Z(n10908) );
  XOR2_X1 U11167 ( .A(n11146), .B(n11147), .Z(n11144) );
  XNOR2_X1 U11168 ( .A(n11148), .B(n11149), .ZN(n10917) );
  XNOR2_X1 U11169 ( .A(n11150), .B(n11151), .ZN(n11149) );
  XOR2_X1 U11170 ( .A(n11152), .B(n11153), .Z(n10921) );
  NAND2_X1 U11171 ( .A1(n11154), .A2(n11155), .ZN(n11152) );
  XOR2_X1 U11172 ( .A(n11156), .B(n11157), .Z(n10925) );
  XOR2_X1 U11173 ( .A(n11158), .B(n11159), .Z(n11157) );
  NAND2_X1 U11174 ( .A1(b_15_), .A2(a_13_), .ZN(n11159) );
  XNOR2_X1 U11175 ( .A(n11160), .B(n11161), .ZN(n10929) );
  XOR2_X1 U11176 ( .A(n11162), .B(n11163), .Z(n11161) );
  NAND2_X1 U11177 ( .A1(b_15_), .A2(a_12_), .ZN(n11163) );
  XNOR2_X1 U11178 ( .A(n11164), .B(n11165), .ZN(n10933) );
  XNOR2_X1 U11179 ( .A(n11166), .B(n11167), .ZN(n11164) );
  NOR2_X1 U11180 ( .A1(n7877), .A2(n10863), .ZN(n11167) );
  XNOR2_X1 U11181 ( .A(n11168), .B(n11169), .ZN(n10936) );
  XOR2_X1 U11182 ( .A(n11170), .B(n11171), .Z(n11169) );
  NAND2_X1 U11183 ( .A1(b_15_), .A2(a_10_), .ZN(n11171) );
  XNOR2_X1 U11184 ( .A(n11172), .B(n11173), .ZN(n10941) );
  XOR2_X1 U11185 ( .A(n11174), .B(n11175), .Z(n11172) );
  NOR2_X1 U11186 ( .A1(n7870), .A2(n10863), .ZN(n11175) );
  XNOR2_X1 U11187 ( .A(n11176), .B(n11177), .ZN(n10944) );
  XNOR2_X1 U11188 ( .A(n11178), .B(n11179), .ZN(n11176) );
  NOR2_X1 U11189 ( .A1(n8037), .A2(n10863), .ZN(n11179) );
  XOR2_X1 U11190 ( .A(n11180), .B(n11181), .Z(n10949) );
  XOR2_X1 U11191 ( .A(n11182), .B(n11183), .Z(n11181) );
  NAND2_X1 U11192 ( .A1(b_15_), .A2(a_7_), .ZN(n11183) );
  XNOR2_X1 U11193 ( .A(n11184), .B(n11185), .ZN(n10957) );
  XNOR2_X1 U11194 ( .A(n11186), .B(n11187), .ZN(n11184) );
  NAND2_X1 U11195 ( .A1(b_15_), .A2(a_5_), .ZN(n11186) );
  XNOR2_X1 U11196 ( .A(n11188), .B(n11189), .ZN(n10961) );
  XNOR2_X1 U11197 ( .A(n11190), .B(n11191), .ZN(n11188) );
  NOR2_X1 U11198 ( .A1(n7398), .A2(n10863), .ZN(n11191) );
  XNOR2_X1 U11199 ( .A(n11192), .B(n11193), .ZN(n10965) );
  XOR2_X1 U11200 ( .A(n11194), .B(n11195), .Z(n11193) );
  NAND2_X1 U11201 ( .A1(b_15_), .A2(a_3_), .ZN(n11195) );
  XOR2_X1 U11202 ( .A(n11196), .B(n11197), .Z(n10969) );
  XOR2_X1 U11203 ( .A(n11198), .B(n11199), .Z(n11197) );
  NAND2_X1 U11204 ( .A1(b_15_), .A2(a_2_), .ZN(n11199) );
  XNOR2_X1 U11205 ( .A(n11200), .B(n11201), .ZN(n7549) );
  XOR2_X1 U11206 ( .A(n11202), .B(n11203), .Z(n11201) );
  NAND2_X1 U11207 ( .A1(b_15_), .A2(a_0_), .ZN(n11203) );
  NAND2_X1 U11208 ( .A1(n11204), .A2(n11205), .ZN(n7491) );
  NAND2_X1 U11209 ( .A1(n10981), .A2(n10978), .ZN(n11205) );
  XNOR2_X1 U11210 ( .A(n7540), .B(n7539), .ZN(n11204) );
  NAND3_X1 U11211 ( .A1(n10981), .A2(n10978), .A3(n11206), .ZN(n7492) );
  XOR2_X1 U11212 ( .A(n7540), .B(n7539), .Z(n11206) );
  NAND2_X1 U11213 ( .A1(n11207), .A2(n11208), .ZN(n10978) );
  NAND3_X1 U11214 ( .A1(a_0_), .A2(n11209), .A3(b_15_), .ZN(n11208) );
  OR2_X1 U11215 ( .A1(n11202), .A2(n11200), .ZN(n11209) );
  NAND2_X1 U11216 ( .A1(n11200), .A2(n11202), .ZN(n11207) );
  NAND2_X1 U11217 ( .A1(n11210), .A2(n11211), .ZN(n11202) );
  NAND3_X1 U11218 ( .A1(a_1_), .A2(n11212), .A3(b_15_), .ZN(n11211) );
  OR2_X1 U11219 ( .A1(n10987), .A2(n10988), .ZN(n11212) );
  NAND2_X1 U11220 ( .A1(n10987), .A2(n10988), .ZN(n11210) );
  NAND2_X1 U11221 ( .A1(n11213), .A2(n11214), .ZN(n10988) );
  NAND3_X1 U11222 ( .A1(a_2_), .A2(n11215), .A3(b_15_), .ZN(n11214) );
  OR2_X1 U11223 ( .A1(n11196), .A2(n11198), .ZN(n11215) );
  NAND2_X1 U11224 ( .A1(n11196), .A2(n11198), .ZN(n11213) );
  NAND2_X1 U11225 ( .A1(n11216), .A2(n11217), .ZN(n11198) );
  NAND3_X1 U11226 ( .A1(a_3_), .A2(n11218), .A3(b_15_), .ZN(n11217) );
  OR2_X1 U11227 ( .A1(n11194), .A2(n11192), .ZN(n11218) );
  NAND2_X1 U11228 ( .A1(n11192), .A2(n11194), .ZN(n11216) );
  NAND2_X1 U11229 ( .A1(n11219), .A2(n11220), .ZN(n11194) );
  NAND3_X1 U11230 ( .A1(a_4_), .A2(n11221), .A3(b_15_), .ZN(n11220) );
  NAND2_X1 U11231 ( .A1(n11190), .A2(n11189), .ZN(n11221) );
  OR2_X1 U11232 ( .A1(n11189), .A2(n11190), .ZN(n11219) );
  AND2_X1 U11233 ( .A1(n11222), .A2(n11223), .ZN(n11190) );
  NAND3_X1 U11234 ( .A1(a_5_), .A2(n11224), .A3(b_15_), .ZN(n11223) );
  OR2_X1 U11235 ( .A1(n11185), .A2(n11187), .ZN(n11224) );
  NAND2_X1 U11236 ( .A1(n11185), .A2(n11187), .ZN(n11222) );
  NAND2_X1 U11237 ( .A1(n11225), .A2(n11226), .ZN(n11187) );
  NAND3_X1 U11238 ( .A1(a_6_), .A2(n11227), .A3(b_15_), .ZN(n11226) );
  OR2_X1 U11239 ( .A1(n11007), .A2(n11008), .ZN(n11227) );
  NAND2_X1 U11240 ( .A1(n11007), .A2(n11008), .ZN(n11225) );
  NAND2_X1 U11241 ( .A1(n11228), .A2(n11229), .ZN(n11008) );
  NAND3_X1 U11242 ( .A1(a_7_), .A2(n11230), .A3(b_15_), .ZN(n11229) );
  OR2_X1 U11243 ( .A1(n11180), .A2(n11182), .ZN(n11230) );
  NAND2_X1 U11244 ( .A1(n11180), .A2(n11182), .ZN(n11228) );
  NAND2_X1 U11245 ( .A1(n11231), .A2(n11232), .ZN(n11182) );
  NAND3_X1 U11246 ( .A1(a_8_), .A2(n11233), .A3(b_15_), .ZN(n11232) );
  NAND2_X1 U11247 ( .A1(n11178), .A2(n11177), .ZN(n11233) );
  OR2_X1 U11248 ( .A1(n11177), .A2(n11178), .ZN(n11231) );
  AND2_X1 U11249 ( .A1(n11234), .A2(n11235), .ZN(n11178) );
  NAND3_X1 U11250 ( .A1(a_9_), .A2(n11236), .A3(b_15_), .ZN(n11235) );
  OR2_X1 U11251 ( .A1(n11173), .A2(n11174), .ZN(n11236) );
  NAND2_X1 U11252 ( .A1(n11173), .A2(n11174), .ZN(n11234) );
  NAND2_X1 U11253 ( .A1(n11237), .A2(n11238), .ZN(n11174) );
  NAND3_X1 U11254 ( .A1(a_10_), .A2(n11239), .A3(b_15_), .ZN(n11238) );
  OR2_X1 U11255 ( .A1(n11168), .A2(n11170), .ZN(n11239) );
  NAND2_X1 U11256 ( .A1(n11168), .A2(n11170), .ZN(n11237) );
  NAND2_X1 U11257 ( .A1(n11240), .A2(n11241), .ZN(n11170) );
  NAND3_X1 U11258 ( .A1(a_11_), .A2(n11242), .A3(b_15_), .ZN(n11241) );
  NAND2_X1 U11259 ( .A1(n11166), .A2(n11165), .ZN(n11242) );
  OR2_X1 U11260 ( .A1(n11165), .A2(n11166), .ZN(n11240) );
  AND2_X1 U11261 ( .A1(n11243), .A2(n11244), .ZN(n11166) );
  NAND3_X1 U11262 ( .A1(a_12_), .A2(n11245), .A3(b_15_), .ZN(n11244) );
  OR2_X1 U11263 ( .A1(n11162), .A2(n11160), .ZN(n11245) );
  NAND2_X1 U11264 ( .A1(n11160), .A2(n11162), .ZN(n11243) );
  NAND2_X1 U11265 ( .A1(n11246), .A2(n11247), .ZN(n11162) );
  NAND3_X1 U11266 ( .A1(a_13_), .A2(n11248), .A3(b_15_), .ZN(n11247) );
  OR2_X1 U11267 ( .A1(n11156), .A2(n11158), .ZN(n11248) );
  NAND2_X1 U11268 ( .A1(n11156), .A2(n11158), .ZN(n11246) );
  NAND2_X1 U11269 ( .A1(n11154), .A2(n11249), .ZN(n11158) );
  NAND2_X1 U11270 ( .A1(n11153), .A2(n11155), .ZN(n11249) );
  NAND2_X1 U11271 ( .A1(n11250), .A2(n11251), .ZN(n11155) );
  NAND2_X1 U11272 ( .A1(b_15_), .A2(a_14_), .ZN(n11251) );
  INV_X1 U11273 ( .A(n11252), .ZN(n11250) );
  XOR2_X1 U11274 ( .A(n11253), .B(n11254), .Z(n11153) );
  XOR2_X1 U11275 ( .A(n11255), .B(n11256), .Z(n11253) );
  NAND2_X1 U11276 ( .A1(a_14_), .A2(n11252), .ZN(n11154) );
  NAND2_X1 U11277 ( .A1(n11257), .A2(n11258), .ZN(n11252) );
  NAND2_X1 U11278 ( .A1(n11148), .A2(n11259), .ZN(n11258) );
  OR2_X1 U11279 ( .A1(n11151), .A2(n11150), .ZN(n11259) );
  XNOR2_X1 U11280 ( .A(n11260), .B(n11261), .ZN(n11148) );
  XNOR2_X1 U11281 ( .A(n11262), .B(n11263), .ZN(n11261) );
  NAND2_X1 U11282 ( .A1(n11150), .A2(n11151), .ZN(n11257) );
  NAND2_X1 U11283 ( .A1(n11264), .A2(n11265), .ZN(n11151) );
  NAND3_X1 U11284 ( .A1(a_16_), .A2(n11266), .A3(b_15_), .ZN(n11265) );
  OR2_X1 U11285 ( .A1(n11043), .A2(n11041), .ZN(n11266) );
  NAND2_X1 U11286 ( .A1(n11041), .A2(n11043), .ZN(n11264) );
  NAND2_X1 U11287 ( .A1(n11267), .A2(n11268), .ZN(n11043) );
  NAND2_X1 U11288 ( .A1(n11147), .A2(n11269), .ZN(n11268) );
  OR2_X1 U11289 ( .A1(n11145), .A2(n11146), .ZN(n11269) );
  NOR2_X1 U11290 ( .A1(n10863), .A2(n7337), .ZN(n11147) );
  NAND2_X1 U11291 ( .A1(n11145), .A2(n11146), .ZN(n11267) );
  NAND2_X1 U11292 ( .A1(n11270), .A2(n11271), .ZN(n11146) );
  NAND3_X1 U11293 ( .A1(a_18_), .A2(n11272), .A3(b_15_), .ZN(n11271) );
  NAND2_X1 U11294 ( .A1(n11142), .A2(n11141), .ZN(n11272) );
  OR2_X1 U11295 ( .A1(n11141), .A2(n11142), .ZN(n11270) );
  AND2_X1 U11296 ( .A1(n11273), .A2(n11274), .ZN(n11142) );
  NAND2_X1 U11297 ( .A1(n11139), .A2(n11275), .ZN(n11274) );
  OR2_X1 U11298 ( .A1(n11136), .A2(n11138), .ZN(n11275) );
  NOR2_X1 U11299 ( .A1(n10863), .A2(n7902), .ZN(n11139) );
  NAND2_X1 U11300 ( .A1(n11136), .A2(n11138), .ZN(n11273) );
  NAND2_X1 U11301 ( .A1(n11276), .A2(n11277), .ZN(n11138) );
  NAND3_X1 U11302 ( .A1(a_20_), .A2(n11278), .A3(b_15_), .ZN(n11277) );
  NAND2_X1 U11303 ( .A1(n11134), .A2(n11133), .ZN(n11278) );
  OR2_X1 U11304 ( .A1(n11133), .A2(n11134), .ZN(n11276) );
  AND2_X1 U11305 ( .A1(n11279), .A2(n11280), .ZN(n11134) );
  NAND2_X1 U11306 ( .A1(n11131), .A2(n11281), .ZN(n11280) );
  OR2_X1 U11307 ( .A1(n11129), .A2(n11130), .ZN(n11281) );
  NOR2_X1 U11308 ( .A1(n10863), .A2(n7909), .ZN(n11131) );
  NAND2_X1 U11309 ( .A1(n11129), .A2(n11130), .ZN(n11279) );
  NAND2_X1 U11310 ( .A1(n11282), .A2(n11283), .ZN(n11130) );
  NAND3_X1 U11311 ( .A1(a_22_), .A2(n11284), .A3(b_15_), .ZN(n11283) );
  NAND2_X1 U11312 ( .A1(n11126), .A2(n11125), .ZN(n11284) );
  OR2_X1 U11313 ( .A1(n11125), .A2(n11126), .ZN(n11282) );
  AND2_X1 U11314 ( .A1(n11285), .A2(n11286), .ZN(n11126) );
  NAND2_X1 U11315 ( .A1(n11123), .A2(n11287), .ZN(n11286) );
  OR2_X1 U11316 ( .A1(n11120), .A2(n11122), .ZN(n11287) );
  NOR2_X1 U11317 ( .A1(n10863), .A2(n7916), .ZN(n11123) );
  NAND2_X1 U11318 ( .A1(n11120), .A2(n11122), .ZN(n11285) );
  NAND2_X1 U11319 ( .A1(n11288), .A2(n11289), .ZN(n11122) );
  NAND3_X1 U11320 ( .A1(a_24_), .A2(n11290), .A3(b_15_), .ZN(n11289) );
  NAND2_X1 U11321 ( .A1(n11118), .A2(n11117), .ZN(n11290) );
  OR2_X1 U11322 ( .A1(n11117), .A2(n11118), .ZN(n11288) );
  AND2_X1 U11323 ( .A1(n11291), .A2(n11292), .ZN(n11118) );
  NAND2_X1 U11324 ( .A1(n11115), .A2(n11293), .ZN(n11292) );
  OR2_X1 U11325 ( .A1(n11113), .A2(n11114), .ZN(n11293) );
  NOR2_X1 U11326 ( .A1(n10863), .A2(n7923), .ZN(n11115) );
  NAND2_X1 U11327 ( .A1(n11113), .A2(n11114), .ZN(n11291) );
  NAND2_X1 U11328 ( .A1(n11110), .A2(n11294), .ZN(n11114) );
  NAND2_X1 U11329 ( .A1(n11109), .A2(n11111), .ZN(n11294) );
  NAND2_X1 U11330 ( .A1(n11295), .A2(n11296), .ZN(n11111) );
  NAND2_X1 U11331 ( .A1(b_15_), .A2(a_26_), .ZN(n11296) );
  INV_X1 U11332 ( .A(n11297), .ZN(n11295) );
  XNOR2_X1 U11333 ( .A(n11298), .B(n11299), .ZN(n11109) );
  NAND2_X1 U11334 ( .A1(n11300), .A2(n11301), .ZN(n11298) );
  NAND2_X1 U11335 ( .A1(a_26_), .A2(n11297), .ZN(n11110) );
  NAND2_X1 U11336 ( .A1(n11081), .A2(n11302), .ZN(n11297) );
  NAND2_X1 U11337 ( .A1(n11080), .A2(n11082), .ZN(n11302) );
  NAND2_X1 U11338 ( .A1(n11303), .A2(n11304), .ZN(n11082) );
  NAND2_X1 U11339 ( .A1(b_15_), .A2(a_27_), .ZN(n11304) );
  INV_X1 U11340 ( .A(n11305), .ZN(n11303) );
  XNOR2_X1 U11341 ( .A(n11306), .B(n11307), .ZN(n11080) );
  XOR2_X1 U11342 ( .A(n11308), .B(n11309), .Z(n11306) );
  NAND2_X1 U11343 ( .A1(b_14_), .A2(a_28_), .ZN(n11308) );
  NAND2_X1 U11344 ( .A1(a_27_), .A2(n11305), .ZN(n11081) );
  NAND2_X1 U11345 ( .A1(n11310), .A2(n11311), .ZN(n11305) );
  NAND3_X1 U11346 ( .A1(a_28_), .A2(n11312), .A3(b_15_), .ZN(n11311) );
  NAND2_X1 U11347 ( .A1(n11090), .A2(n11088), .ZN(n11312) );
  OR2_X1 U11348 ( .A1(n11088), .A2(n11090), .ZN(n11310) );
  AND2_X1 U11349 ( .A1(n11313), .A2(n11314), .ZN(n11090) );
  NAND2_X1 U11350 ( .A1(n11105), .A2(n11315), .ZN(n11314) );
  OR2_X1 U11351 ( .A1(n11106), .A2(n11107), .ZN(n11315) );
  NOR2_X1 U11352 ( .A1(n10863), .A2(n7946), .ZN(n11105) );
  NAND2_X1 U11353 ( .A1(n11107), .A2(n11106), .ZN(n11313) );
  NAND2_X1 U11354 ( .A1(n11316), .A2(n11317), .ZN(n11106) );
  NAND2_X1 U11355 ( .A1(b_13_), .A2(n11318), .ZN(n11317) );
  NAND2_X1 U11356 ( .A1(n7268), .A2(n11319), .ZN(n11318) );
  NAND2_X1 U11357 ( .A1(a_31_), .A2(n11103), .ZN(n11319) );
  NAND2_X1 U11358 ( .A1(b_14_), .A2(n11320), .ZN(n11316) );
  NAND2_X1 U11359 ( .A1(n7272), .A2(n11321), .ZN(n11320) );
  NAND2_X1 U11360 ( .A1(a_30_), .A2(n11322), .ZN(n11321) );
  AND3_X1 U11361 ( .A1(b_14_), .A2(n7954), .A3(b_15_), .ZN(n11107) );
  XNOR2_X1 U11362 ( .A(n11323), .B(n11324), .ZN(n11088) );
  XOR2_X1 U11363 ( .A(n11325), .B(n11326), .Z(n11323) );
  XNOR2_X1 U11364 ( .A(n11327), .B(n11328), .ZN(n11113) );
  NAND2_X1 U11365 ( .A1(n11329), .A2(n11330), .ZN(n11327) );
  XNOR2_X1 U11366 ( .A(n11331), .B(n11332), .ZN(n11117) );
  XOR2_X1 U11367 ( .A(n11333), .B(n11334), .Z(n11331) );
  XNOR2_X1 U11368 ( .A(n11335), .B(n11336), .ZN(n11120) );
  XNOR2_X1 U11369 ( .A(n11337), .B(n11338), .ZN(n11335) );
  NOR2_X1 U11370 ( .A1(n7691), .A2(n11103), .ZN(n11338) );
  XOR2_X1 U11371 ( .A(n11339), .B(n11340), .Z(n11125) );
  XNOR2_X1 U11372 ( .A(n11341), .B(n11342), .ZN(n11340) );
  XNOR2_X1 U11373 ( .A(n11343), .B(n11344), .ZN(n11129) );
  XOR2_X1 U11374 ( .A(n11345), .B(n11346), .Z(n11344) );
  NAND2_X1 U11375 ( .A1(b_14_), .A2(a_22_), .ZN(n11346) );
  XNOR2_X1 U11376 ( .A(n11347), .B(n11348), .ZN(n11133) );
  XOR2_X1 U11377 ( .A(n11349), .B(n11350), .Z(n11347) );
  XNOR2_X1 U11378 ( .A(n11351), .B(n11352), .ZN(n11136) );
  XNOR2_X1 U11379 ( .A(n11353), .B(n11354), .ZN(n11351) );
  NOR2_X1 U11380 ( .A1(n7987), .A2(n11103), .ZN(n11354) );
  XOR2_X1 U11381 ( .A(n11355), .B(n11356), .Z(n11141) );
  XNOR2_X1 U11382 ( .A(n11357), .B(n11358), .ZN(n11356) );
  XNOR2_X1 U11383 ( .A(n11359), .B(n11360), .ZN(n11145) );
  XNOR2_X1 U11384 ( .A(n11361), .B(n11362), .ZN(n11359) );
  NOR2_X1 U11385 ( .A1(n7764), .A2(n11103), .ZN(n11362) );
  XOR2_X1 U11386 ( .A(n11363), .B(n11364), .Z(n11041) );
  XOR2_X1 U11387 ( .A(n11365), .B(n11366), .Z(n11363) );
  NOR2_X1 U11388 ( .A1(n7337), .A2(n11103), .ZN(n11366) );
  XNOR2_X1 U11389 ( .A(n11367), .B(n11368), .ZN(n11156) );
  XNOR2_X1 U11390 ( .A(n11369), .B(n11370), .ZN(n11367) );
  XNOR2_X1 U11391 ( .A(n11371), .B(n11372), .ZN(n11160) );
  NAND2_X1 U11392 ( .A1(n11373), .A2(n11374), .ZN(n11371) );
  XNOR2_X1 U11393 ( .A(n11375), .B(n11376), .ZN(n11165) );
  XOR2_X1 U11394 ( .A(n11377), .B(n11378), .Z(n11375) );
  XNOR2_X1 U11395 ( .A(n11379), .B(n11380), .ZN(n11168) );
  XNOR2_X1 U11396 ( .A(n11381), .B(n11382), .ZN(n11379) );
  NOR2_X1 U11397 ( .A1(n7877), .A2(n11103), .ZN(n11382) );
  XNOR2_X1 U11398 ( .A(n11383), .B(n11384), .ZN(n11173) );
  XNOR2_X1 U11399 ( .A(n11385), .B(n11386), .ZN(n11383) );
  XNOR2_X1 U11400 ( .A(n11387), .B(n11388), .ZN(n11177) );
  XOR2_X1 U11401 ( .A(n11389), .B(n11390), .Z(n11387) );
  NOR2_X1 U11402 ( .A1(n7870), .A2(n11103), .ZN(n11390) );
  XNOR2_X1 U11403 ( .A(n11391), .B(n11392), .ZN(n11180) );
  NAND2_X1 U11404 ( .A1(n11393), .A2(n11394), .ZN(n11391) );
  XNOR2_X1 U11405 ( .A(n11395), .B(n11396), .ZN(n11007) );
  NAND2_X1 U11406 ( .A1(n11397), .A2(n11398), .ZN(n11395) );
  XNOR2_X1 U11407 ( .A(n11399), .B(n11400), .ZN(n11185) );
  NAND2_X1 U11408 ( .A1(n11401), .A2(n11402), .ZN(n11399) );
  XOR2_X1 U11409 ( .A(n11403), .B(n11404), .Z(n11189) );
  NAND2_X1 U11410 ( .A1(n11405), .A2(n11406), .ZN(n11403) );
  XNOR2_X1 U11411 ( .A(n11407), .B(n11408), .ZN(n11192) );
  XNOR2_X1 U11412 ( .A(n11409), .B(n11410), .ZN(n11408) );
  XNOR2_X1 U11413 ( .A(n11411), .B(n11412), .ZN(n11196) );
  XNOR2_X1 U11414 ( .A(n11413), .B(n11414), .ZN(n11412) );
  XNOR2_X1 U11415 ( .A(n11415), .B(n11416), .ZN(n10987) );
  XNOR2_X1 U11416 ( .A(n11417), .B(n11418), .ZN(n11415) );
  NOR2_X1 U11417 ( .A1(n7832), .A2(n11103), .ZN(n11418) );
  XNOR2_X1 U11418 ( .A(n11419), .B(n11420), .ZN(n11200) );
  XNOR2_X1 U11419 ( .A(n11421), .B(n11422), .ZN(n11420) );
  INV_X1 U11420 ( .A(n10979), .ZN(n10981) );
  XOR2_X1 U11421 ( .A(n11423), .B(n11424), .Z(n10979) );
  XNOR2_X1 U11422 ( .A(n11425), .B(n11426), .ZN(n11423) );
  NOR2_X1 U11423 ( .A1(n7613), .A2(n11103), .ZN(n11426) );
  NAND4_X1 U11424 ( .A1(n7539), .A2(n7538), .A3(n7540), .A4(n7534), .ZN(n7496)
         );
  INV_X1 U11425 ( .A(n11427), .ZN(n7534) );
  NAND2_X1 U11426 ( .A1(n11428), .A2(n11429), .ZN(n7540) );
  NAND3_X1 U11427 ( .A1(a_0_), .A2(n11430), .A3(b_14_), .ZN(n11429) );
  NAND2_X1 U11428 ( .A1(n11425), .A2(n11424), .ZN(n11430) );
  OR2_X1 U11429 ( .A1(n11424), .A2(n11425), .ZN(n11428) );
  AND2_X1 U11430 ( .A1(n11431), .A2(n11432), .ZN(n11425) );
  NAND2_X1 U11431 ( .A1(n11422), .A2(n11433), .ZN(n11432) );
  OR2_X1 U11432 ( .A1(n11421), .A2(n11419), .ZN(n11433) );
  NOR2_X1 U11433 ( .A1(n11103), .A2(n7411), .ZN(n11422) );
  NAND2_X1 U11434 ( .A1(n11419), .A2(n11421), .ZN(n11431) );
  NAND2_X1 U11435 ( .A1(n11434), .A2(n11435), .ZN(n11421) );
  NAND3_X1 U11436 ( .A1(a_2_), .A2(n11436), .A3(b_14_), .ZN(n11435) );
  NAND2_X1 U11437 ( .A1(n11417), .A2(n11416), .ZN(n11436) );
  OR2_X1 U11438 ( .A1(n11416), .A2(n11417), .ZN(n11434) );
  AND2_X1 U11439 ( .A1(n11437), .A2(n11438), .ZN(n11417) );
  NAND2_X1 U11440 ( .A1(n11414), .A2(n11439), .ZN(n11438) );
  OR2_X1 U11441 ( .A1(n11413), .A2(n11411), .ZN(n11439) );
  NOR2_X1 U11442 ( .A1(n11103), .A2(n7850), .ZN(n11414) );
  NAND2_X1 U11443 ( .A1(n11411), .A2(n11413), .ZN(n11437) );
  NAND2_X1 U11444 ( .A1(n11440), .A2(n11441), .ZN(n11413) );
  NAND2_X1 U11445 ( .A1(n11410), .A2(n11442), .ZN(n11441) );
  OR2_X1 U11446 ( .A1(n11409), .A2(n11407), .ZN(n11442) );
  NOR2_X1 U11447 ( .A1(n11103), .A2(n7398), .ZN(n11410) );
  NAND2_X1 U11448 ( .A1(n11407), .A2(n11409), .ZN(n11440) );
  NAND2_X1 U11449 ( .A1(n11405), .A2(n11443), .ZN(n11409) );
  NAND2_X1 U11450 ( .A1(n11404), .A2(n11406), .ZN(n11443) );
  NAND2_X1 U11451 ( .A1(n11444), .A2(n11445), .ZN(n11406) );
  NAND2_X1 U11452 ( .A1(b_14_), .A2(a_5_), .ZN(n11445) );
  INV_X1 U11453 ( .A(n11446), .ZN(n11444) );
  XNOR2_X1 U11454 ( .A(n11447), .B(n11448), .ZN(n11404) );
  XOR2_X1 U11455 ( .A(n11449), .B(n11450), .Z(n11448) );
  NAND2_X1 U11456 ( .A1(b_13_), .A2(a_6_), .ZN(n11450) );
  NAND2_X1 U11457 ( .A1(a_5_), .A2(n11446), .ZN(n11405) );
  NAND2_X1 U11458 ( .A1(n11401), .A2(n11451), .ZN(n11446) );
  NAND2_X1 U11459 ( .A1(n11400), .A2(n11402), .ZN(n11451) );
  NAND2_X1 U11460 ( .A1(n11452), .A2(n11453), .ZN(n11402) );
  NAND2_X1 U11461 ( .A1(b_14_), .A2(a_6_), .ZN(n11453) );
  INV_X1 U11462 ( .A(n11454), .ZN(n11452) );
  XNOR2_X1 U11463 ( .A(n11455), .B(n11456), .ZN(n11400) );
  XOR2_X1 U11464 ( .A(n11457), .B(n11458), .Z(n11456) );
  NAND2_X1 U11465 ( .A1(b_13_), .A2(a_7_), .ZN(n11458) );
  NAND2_X1 U11466 ( .A1(a_6_), .A2(n11454), .ZN(n11401) );
  NAND2_X1 U11467 ( .A1(n11397), .A2(n11459), .ZN(n11454) );
  NAND2_X1 U11468 ( .A1(n11396), .A2(n11398), .ZN(n11459) );
  NAND2_X1 U11469 ( .A1(n11460), .A2(n11461), .ZN(n11398) );
  NAND2_X1 U11470 ( .A1(b_14_), .A2(a_7_), .ZN(n11461) );
  INV_X1 U11471 ( .A(n11462), .ZN(n11460) );
  XNOR2_X1 U11472 ( .A(n11463), .B(n11464), .ZN(n11396) );
  XOR2_X1 U11473 ( .A(n11465), .B(n11466), .Z(n11464) );
  NAND2_X1 U11474 ( .A1(b_13_), .A2(a_8_), .ZN(n11466) );
  NAND2_X1 U11475 ( .A1(a_7_), .A2(n11462), .ZN(n11397) );
  NAND2_X1 U11476 ( .A1(n11393), .A2(n11467), .ZN(n11462) );
  NAND2_X1 U11477 ( .A1(n11392), .A2(n11394), .ZN(n11467) );
  NAND2_X1 U11478 ( .A1(n11468), .A2(n11469), .ZN(n11394) );
  NAND2_X1 U11479 ( .A1(b_14_), .A2(a_8_), .ZN(n11469) );
  INV_X1 U11480 ( .A(n11470), .ZN(n11468) );
  XNOR2_X1 U11481 ( .A(n11471), .B(n11472), .ZN(n11392) );
  XNOR2_X1 U11482 ( .A(n11473), .B(n11474), .ZN(n11471) );
  NOR2_X1 U11483 ( .A1(n7870), .A2(n11322), .ZN(n11474) );
  NAND2_X1 U11484 ( .A1(a_8_), .A2(n11470), .ZN(n11393) );
  NAND2_X1 U11485 ( .A1(n11475), .A2(n11476), .ZN(n11470) );
  NAND3_X1 U11486 ( .A1(a_9_), .A2(n11477), .A3(b_14_), .ZN(n11476) );
  OR2_X1 U11487 ( .A1(n11389), .A2(n11388), .ZN(n11477) );
  NAND2_X1 U11488 ( .A1(n11388), .A2(n11389), .ZN(n11475) );
  NAND2_X1 U11489 ( .A1(n11478), .A2(n11479), .ZN(n11389) );
  NAND2_X1 U11490 ( .A1(n11386), .A2(n11480), .ZN(n11479) );
  NAND2_X1 U11491 ( .A1(n11385), .A2(n11384), .ZN(n11480) );
  NOR2_X1 U11492 ( .A1(n11103), .A2(n7799), .ZN(n11386) );
  OR2_X1 U11493 ( .A1(n11384), .A2(n11385), .ZN(n11478) );
  AND2_X1 U11494 ( .A1(n11481), .A2(n11482), .ZN(n11385) );
  NAND3_X1 U11495 ( .A1(a_11_), .A2(n11483), .A3(b_14_), .ZN(n11482) );
  NAND2_X1 U11496 ( .A1(n11381), .A2(n11380), .ZN(n11483) );
  OR2_X1 U11497 ( .A1(n11380), .A2(n11381), .ZN(n11481) );
  AND2_X1 U11498 ( .A1(n11484), .A2(n11485), .ZN(n11381) );
  NAND2_X1 U11499 ( .A1(n11378), .A2(n11486), .ZN(n11485) );
  OR2_X1 U11500 ( .A1(n11377), .A2(n11376), .ZN(n11486) );
  NOR2_X1 U11501 ( .A1(n11103), .A2(n8020), .ZN(n11378) );
  NAND2_X1 U11502 ( .A1(n11376), .A2(n11377), .ZN(n11484) );
  NAND2_X1 U11503 ( .A1(n11373), .A2(n11487), .ZN(n11377) );
  NAND2_X1 U11504 ( .A1(n11372), .A2(n11374), .ZN(n11487) );
  NAND2_X1 U11505 ( .A1(n11488), .A2(n11489), .ZN(n11374) );
  NAND2_X1 U11506 ( .A1(b_14_), .A2(a_13_), .ZN(n11489) );
  INV_X1 U11507 ( .A(n11490), .ZN(n11488) );
  XOR2_X1 U11508 ( .A(n11491), .B(n11492), .Z(n11372) );
  XOR2_X1 U11509 ( .A(n11493), .B(n11494), .Z(n11491) );
  NOR2_X1 U11510 ( .A1(n7782), .A2(n11322), .ZN(n11494) );
  NAND2_X1 U11511 ( .A1(a_13_), .A2(n11490), .ZN(n11373) );
  NAND2_X1 U11512 ( .A1(n11495), .A2(n11496), .ZN(n11490) );
  NAND2_X1 U11513 ( .A1(n11370), .A2(n11497), .ZN(n11496) );
  NAND2_X1 U11514 ( .A1(n11369), .A2(n11368), .ZN(n11497) );
  OR2_X1 U11515 ( .A1(n11368), .A2(n11369), .ZN(n11495) );
  AND2_X1 U11516 ( .A1(n11498), .A2(n11499), .ZN(n11369) );
  NAND2_X1 U11517 ( .A1(n11256), .A2(n11500), .ZN(n11499) );
  OR2_X1 U11518 ( .A1(n11255), .A2(n11254), .ZN(n11500) );
  NOR2_X1 U11519 ( .A1(n11103), .A2(n7346), .ZN(n11256) );
  NAND2_X1 U11520 ( .A1(n11254), .A2(n11255), .ZN(n11498) );
  NAND2_X1 U11521 ( .A1(n11501), .A2(n11502), .ZN(n11255) );
  NAND2_X1 U11522 ( .A1(n11263), .A2(n11503), .ZN(n11502) );
  OR2_X1 U11523 ( .A1(n11262), .A2(n11260), .ZN(n11503) );
  NOR2_X1 U11524 ( .A1(n11103), .A2(n7773), .ZN(n11263) );
  NAND2_X1 U11525 ( .A1(n11260), .A2(n11262), .ZN(n11501) );
  NAND2_X1 U11526 ( .A1(n11504), .A2(n11505), .ZN(n11262) );
  NAND3_X1 U11527 ( .A1(a_17_), .A2(n11506), .A3(b_14_), .ZN(n11505) );
  OR2_X1 U11528 ( .A1(n11365), .A2(n11364), .ZN(n11506) );
  NAND2_X1 U11529 ( .A1(n11364), .A2(n11365), .ZN(n11504) );
  NAND2_X1 U11530 ( .A1(n11507), .A2(n11508), .ZN(n11365) );
  NAND3_X1 U11531 ( .A1(a_18_), .A2(n11509), .A3(b_14_), .ZN(n11508) );
  NAND2_X1 U11532 ( .A1(n11361), .A2(n11360), .ZN(n11509) );
  OR2_X1 U11533 ( .A1(n11360), .A2(n11361), .ZN(n11507) );
  AND2_X1 U11534 ( .A1(n11510), .A2(n11511), .ZN(n11361) );
  NAND2_X1 U11535 ( .A1(n11358), .A2(n11512), .ZN(n11511) );
  OR2_X1 U11536 ( .A1(n11357), .A2(n11355), .ZN(n11512) );
  NOR2_X1 U11537 ( .A1(n11103), .A2(n7902), .ZN(n11358) );
  NAND2_X1 U11538 ( .A1(n11355), .A2(n11357), .ZN(n11510) );
  NAND2_X1 U11539 ( .A1(n11513), .A2(n11514), .ZN(n11357) );
  NAND3_X1 U11540 ( .A1(a_20_), .A2(n11515), .A3(b_14_), .ZN(n11514) );
  NAND2_X1 U11541 ( .A1(n11353), .A2(n11352), .ZN(n11515) );
  OR2_X1 U11542 ( .A1(n11352), .A2(n11353), .ZN(n11513) );
  AND2_X1 U11543 ( .A1(n11516), .A2(n11517), .ZN(n11353) );
  NAND2_X1 U11544 ( .A1(n11350), .A2(n11518), .ZN(n11517) );
  OR2_X1 U11545 ( .A1(n11349), .A2(n11348), .ZN(n11518) );
  NOR2_X1 U11546 ( .A1(n11103), .A2(n7909), .ZN(n11350) );
  NAND2_X1 U11547 ( .A1(n11348), .A2(n11349), .ZN(n11516) );
  NAND2_X1 U11548 ( .A1(n11519), .A2(n11520), .ZN(n11349) );
  NAND3_X1 U11549 ( .A1(a_22_), .A2(n11521), .A3(b_14_), .ZN(n11520) );
  OR2_X1 U11550 ( .A1(n11345), .A2(n11343), .ZN(n11521) );
  NAND2_X1 U11551 ( .A1(n11343), .A2(n11345), .ZN(n11519) );
  NAND2_X1 U11552 ( .A1(n11522), .A2(n11523), .ZN(n11345) );
  NAND2_X1 U11553 ( .A1(n11342), .A2(n11524), .ZN(n11523) );
  OR2_X1 U11554 ( .A1(n11341), .A2(n11339), .ZN(n11524) );
  NOR2_X1 U11555 ( .A1(n11103), .A2(n7916), .ZN(n11342) );
  NAND2_X1 U11556 ( .A1(n11339), .A2(n11341), .ZN(n11522) );
  NAND2_X1 U11557 ( .A1(n11525), .A2(n11526), .ZN(n11341) );
  NAND3_X1 U11558 ( .A1(a_24_), .A2(n11527), .A3(b_14_), .ZN(n11526) );
  NAND2_X1 U11559 ( .A1(n11337), .A2(n11336), .ZN(n11527) );
  OR2_X1 U11560 ( .A1(n11336), .A2(n11337), .ZN(n11525) );
  AND2_X1 U11561 ( .A1(n11528), .A2(n11529), .ZN(n11337) );
  NAND2_X1 U11562 ( .A1(n11334), .A2(n11530), .ZN(n11529) );
  OR2_X1 U11563 ( .A1(n11333), .A2(n11332), .ZN(n11530) );
  NOR2_X1 U11564 ( .A1(n11103), .A2(n7923), .ZN(n11334) );
  NAND2_X1 U11565 ( .A1(n11332), .A2(n11333), .ZN(n11528) );
  NAND2_X1 U11566 ( .A1(n11329), .A2(n11531), .ZN(n11333) );
  NAND2_X1 U11567 ( .A1(n11328), .A2(n11330), .ZN(n11531) );
  NAND2_X1 U11568 ( .A1(n11532), .A2(n11533), .ZN(n11330) );
  NAND2_X1 U11569 ( .A1(b_14_), .A2(a_26_), .ZN(n11533) );
  INV_X1 U11570 ( .A(n11534), .ZN(n11532) );
  XNOR2_X1 U11571 ( .A(n11535), .B(n11536), .ZN(n11328) );
  NAND2_X1 U11572 ( .A1(n11537), .A2(n11538), .ZN(n11535) );
  NAND2_X1 U11573 ( .A1(a_26_), .A2(n11534), .ZN(n11329) );
  NAND2_X1 U11574 ( .A1(n11300), .A2(n11539), .ZN(n11534) );
  NAND2_X1 U11575 ( .A1(n11299), .A2(n11301), .ZN(n11539) );
  NAND2_X1 U11576 ( .A1(n11540), .A2(n11541), .ZN(n11301) );
  NAND2_X1 U11577 ( .A1(b_14_), .A2(a_27_), .ZN(n11541) );
  INV_X1 U11578 ( .A(n11542), .ZN(n11540) );
  XNOR2_X1 U11579 ( .A(n11543), .B(n11544), .ZN(n11299) );
  XOR2_X1 U11580 ( .A(n11545), .B(n11546), .Z(n11543) );
  NAND2_X1 U11581 ( .A1(b_13_), .A2(a_28_), .ZN(n11545) );
  NAND2_X1 U11582 ( .A1(a_27_), .A2(n11542), .ZN(n11300) );
  NAND2_X1 U11583 ( .A1(n11547), .A2(n11548), .ZN(n11542) );
  NAND3_X1 U11584 ( .A1(a_28_), .A2(n11549), .A3(b_14_), .ZN(n11548) );
  NAND2_X1 U11585 ( .A1(n11309), .A2(n11307), .ZN(n11549) );
  OR2_X1 U11586 ( .A1(n11307), .A2(n11309), .ZN(n11547) );
  AND2_X1 U11587 ( .A1(n11550), .A2(n11551), .ZN(n11309) );
  NAND2_X1 U11588 ( .A1(n11324), .A2(n11552), .ZN(n11551) );
  OR2_X1 U11589 ( .A1(n11325), .A2(n11326), .ZN(n11552) );
  NOR2_X1 U11590 ( .A1(n11103), .A2(n7946), .ZN(n11324) );
  NAND2_X1 U11591 ( .A1(n11326), .A2(n11325), .ZN(n11550) );
  NAND2_X1 U11592 ( .A1(n11553), .A2(n11554), .ZN(n11325) );
  NAND2_X1 U11593 ( .A1(b_12_), .A2(n11555), .ZN(n11554) );
  NAND2_X1 U11594 ( .A1(n7268), .A2(n11556), .ZN(n11555) );
  NAND2_X1 U11595 ( .A1(a_31_), .A2(n11322), .ZN(n11556) );
  NAND2_X1 U11596 ( .A1(b_13_), .A2(n11557), .ZN(n11553) );
  NAND2_X1 U11597 ( .A1(n7272), .A2(n11558), .ZN(n11557) );
  NAND2_X1 U11598 ( .A1(a_30_), .A2(n11559), .ZN(n11558) );
  AND3_X1 U11599 ( .A1(b_13_), .A2(n7954), .A3(b_14_), .ZN(n11326) );
  XNOR2_X1 U11600 ( .A(n11560), .B(n11561), .ZN(n11307) );
  XOR2_X1 U11601 ( .A(n11562), .B(n11563), .Z(n11560) );
  XNOR2_X1 U11602 ( .A(n11564), .B(n11565), .ZN(n11332) );
  NAND2_X1 U11603 ( .A1(n11566), .A2(n11567), .ZN(n11564) );
  XNOR2_X1 U11604 ( .A(n11568), .B(n11569), .ZN(n11336) );
  XOR2_X1 U11605 ( .A(n11570), .B(n11571), .Z(n11568) );
  XNOR2_X1 U11606 ( .A(n11572), .B(n11573), .ZN(n11339) );
  XNOR2_X1 U11607 ( .A(n11574), .B(n11575), .ZN(n11572) );
  NOR2_X1 U11608 ( .A1(n7691), .A2(n11322), .ZN(n11575) );
  XNOR2_X1 U11609 ( .A(n11576), .B(n11577), .ZN(n11343) );
  XNOR2_X1 U11610 ( .A(n11578), .B(n11579), .ZN(n11577) );
  XNOR2_X1 U11611 ( .A(n11580), .B(n11581), .ZN(n11348) );
  XOR2_X1 U11612 ( .A(n11582), .B(n11583), .Z(n11581) );
  NAND2_X1 U11613 ( .A1(b_13_), .A2(a_22_), .ZN(n11583) );
  XNOR2_X1 U11614 ( .A(n11584), .B(n11585), .ZN(n11352) );
  XOR2_X1 U11615 ( .A(n11586), .B(n11587), .Z(n11584) );
  XNOR2_X1 U11616 ( .A(n11588), .B(n11589), .ZN(n11355) );
  XNOR2_X1 U11617 ( .A(n11590), .B(n11591), .ZN(n11588) );
  NOR2_X1 U11618 ( .A1(n7987), .A2(n11322), .ZN(n11591) );
  XOR2_X1 U11619 ( .A(n11592), .B(n11593), .Z(n11360) );
  XNOR2_X1 U11620 ( .A(n11594), .B(n11595), .ZN(n11593) );
  XNOR2_X1 U11621 ( .A(n11596), .B(n11597), .ZN(n11364) );
  XNOR2_X1 U11622 ( .A(n11598), .B(n11599), .ZN(n11596) );
  XNOR2_X1 U11623 ( .A(n11600), .B(n11601), .ZN(n11260) );
  XOR2_X1 U11624 ( .A(n11602), .B(n11603), .Z(n11600) );
  NAND2_X1 U11625 ( .A1(b_13_), .A2(a_17_), .ZN(n11602) );
  XNOR2_X1 U11626 ( .A(n11604), .B(n11605), .ZN(n11254) );
  XNOR2_X1 U11627 ( .A(n11606), .B(n11607), .ZN(n11604) );
  NOR2_X1 U11628 ( .A1(n7773), .A2(n11322), .ZN(n11607) );
  XOR2_X1 U11629 ( .A(n11608), .B(n11609), .Z(n11368) );
  XOR2_X1 U11630 ( .A(n11610), .B(n11611), .Z(n11609) );
  NAND2_X1 U11631 ( .A1(b_13_), .A2(a_15_), .ZN(n11611) );
  XOR2_X1 U11632 ( .A(n11612), .B(n11613), .Z(n11376) );
  XOR2_X1 U11633 ( .A(n11614), .B(n11615), .Z(n11612) );
  XNOR2_X1 U11634 ( .A(n11616), .B(n11617), .ZN(n11380) );
  XNOR2_X1 U11635 ( .A(n11618), .B(n11619), .ZN(n11616) );
  NAND2_X1 U11636 ( .A1(b_13_), .A2(a_12_), .ZN(n11618) );
  XOR2_X1 U11637 ( .A(n11620), .B(n11621), .Z(n11384) );
  XOR2_X1 U11638 ( .A(n11622), .B(n11623), .Z(n11621) );
  NAND2_X1 U11639 ( .A1(b_13_), .A2(a_11_), .ZN(n11623) );
  XNOR2_X1 U11640 ( .A(n11624), .B(n11625), .ZN(n11388) );
  XOR2_X1 U11641 ( .A(n11626), .B(n11627), .Z(n11625) );
  NAND2_X1 U11642 ( .A1(b_13_), .A2(a_10_), .ZN(n11627) );
  XNOR2_X1 U11643 ( .A(n11628), .B(n11629), .ZN(n11407) );
  XNOR2_X1 U11644 ( .A(n11630), .B(n11631), .ZN(n11628) );
  NOR2_X1 U11645 ( .A1(n7393), .A2(n11322), .ZN(n11631) );
  XNOR2_X1 U11646 ( .A(n11632), .B(n11633), .ZN(n11411) );
  XOR2_X1 U11647 ( .A(n11634), .B(n11635), .Z(n11633) );
  NAND2_X1 U11648 ( .A1(b_13_), .A2(a_4_), .ZN(n11635) );
  XNOR2_X1 U11649 ( .A(n11636), .B(n11637), .ZN(n11416) );
  XOR2_X1 U11650 ( .A(n11638), .B(n11639), .Z(n11636) );
  NOR2_X1 U11651 ( .A1(n7850), .A2(n11322), .ZN(n11639) );
  XNOR2_X1 U11652 ( .A(n11640), .B(n11641), .ZN(n11419) );
  XOR2_X1 U11653 ( .A(n11642), .B(n11643), .Z(n11641) );
  NAND2_X1 U11654 ( .A1(b_13_), .A2(a_2_), .ZN(n11643) );
  XNOR2_X1 U11655 ( .A(n11644), .B(n11645), .ZN(n11424) );
  XOR2_X1 U11656 ( .A(n11646), .B(n11647), .Z(n11644) );
  NOR2_X1 U11657 ( .A1(n7411), .A2(n11322), .ZN(n11647) );
  NAND2_X1 U11658 ( .A1(n11648), .A2(n11649), .ZN(n7538) );
  XNOR2_X1 U11659 ( .A(n11650), .B(n11651), .ZN(n7539) );
  XNOR2_X1 U11660 ( .A(n11652), .B(n11653), .ZN(n11651) );
  NAND2_X1 U11661 ( .A1(n11427), .A2(n11654), .ZN(n7500) );
  XOR2_X1 U11662 ( .A(n7531), .B(n7530), .Z(n11654) );
  NOR2_X1 U11663 ( .A1(n11649), .A2(n11648), .ZN(n11427) );
  AND2_X1 U11664 ( .A1(n11655), .A2(n11656), .ZN(n11648) );
  NAND2_X1 U11665 ( .A1(n11653), .A2(n11657), .ZN(n11656) );
  OR2_X1 U11666 ( .A1(n11652), .A2(n11650), .ZN(n11657) );
  NOR2_X1 U11667 ( .A1(n11322), .A2(n7613), .ZN(n11653) );
  NAND2_X1 U11668 ( .A1(n11650), .A2(n11652), .ZN(n11655) );
  NAND2_X1 U11669 ( .A1(n11658), .A2(n11659), .ZN(n11652) );
  NAND3_X1 U11670 ( .A1(a_1_), .A2(n11660), .A3(b_13_), .ZN(n11659) );
  OR2_X1 U11671 ( .A1(n11646), .A2(n11645), .ZN(n11660) );
  NAND2_X1 U11672 ( .A1(n11645), .A2(n11646), .ZN(n11658) );
  NAND2_X1 U11673 ( .A1(n11661), .A2(n11662), .ZN(n11646) );
  NAND3_X1 U11674 ( .A1(a_2_), .A2(n11663), .A3(b_13_), .ZN(n11662) );
  OR2_X1 U11675 ( .A1(n11642), .A2(n11640), .ZN(n11663) );
  NAND2_X1 U11676 ( .A1(n11640), .A2(n11642), .ZN(n11661) );
  NAND2_X1 U11677 ( .A1(n11664), .A2(n11665), .ZN(n11642) );
  NAND3_X1 U11678 ( .A1(a_3_), .A2(n11666), .A3(b_13_), .ZN(n11665) );
  OR2_X1 U11679 ( .A1(n11638), .A2(n11637), .ZN(n11666) );
  NAND2_X1 U11680 ( .A1(n11637), .A2(n11638), .ZN(n11664) );
  NAND2_X1 U11681 ( .A1(n11667), .A2(n11668), .ZN(n11638) );
  NAND3_X1 U11682 ( .A1(a_4_), .A2(n11669), .A3(b_13_), .ZN(n11668) );
  OR2_X1 U11683 ( .A1(n11634), .A2(n11632), .ZN(n11669) );
  NAND2_X1 U11684 ( .A1(n11632), .A2(n11634), .ZN(n11667) );
  NAND2_X1 U11685 ( .A1(n11670), .A2(n11671), .ZN(n11634) );
  NAND3_X1 U11686 ( .A1(a_5_), .A2(n11672), .A3(b_13_), .ZN(n11671) );
  NAND2_X1 U11687 ( .A1(n11630), .A2(n11629), .ZN(n11672) );
  OR2_X1 U11688 ( .A1(n11629), .A2(n11630), .ZN(n11670) );
  AND2_X1 U11689 ( .A1(n11673), .A2(n11674), .ZN(n11630) );
  NAND3_X1 U11690 ( .A1(a_6_), .A2(n11675), .A3(b_13_), .ZN(n11674) );
  OR2_X1 U11691 ( .A1(n11449), .A2(n11447), .ZN(n11675) );
  NAND2_X1 U11692 ( .A1(n11447), .A2(n11449), .ZN(n11673) );
  NAND2_X1 U11693 ( .A1(n11676), .A2(n11677), .ZN(n11449) );
  NAND3_X1 U11694 ( .A1(a_7_), .A2(n11678), .A3(b_13_), .ZN(n11677) );
  OR2_X1 U11695 ( .A1(n11457), .A2(n11455), .ZN(n11678) );
  NAND2_X1 U11696 ( .A1(n11455), .A2(n11457), .ZN(n11676) );
  NAND2_X1 U11697 ( .A1(n11679), .A2(n11680), .ZN(n11457) );
  NAND3_X1 U11698 ( .A1(a_8_), .A2(n11681), .A3(b_13_), .ZN(n11680) );
  OR2_X1 U11699 ( .A1(n11465), .A2(n11463), .ZN(n11681) );
  NAND2_X1 U11700 ( .A1(n11463), .A2(n11465), .ZN(n11679) );
  NAND2_X1 U11701 ( .A1(n11682), .A2(n11683), .ZN(n11465) );
  NAND3_X1 U11702 ( .A1(a_9_), .A2(n11684), .A3(b_13_), .ZN(n11683) );
  NAND2_X1 U11703 ( .A1(n11473), .A2(n11472), .ZN(n11684) );
  OR2_X1 U11704 ( .A1(n11472), .A2(n11473), .ZN(n11682) );
  AND2_X1 U11705 ( .A1(n11685), .A2(n11686), .ZN(n11473) );
  NAND3_X1 U11706 ( .A1(a_10_), .A2(n11687), .A3(b_13_), .ZN(n11686) );
  OR2_X1 U11707 ( .A1(n11626), .A2(n11624), .ZN(n11687) );
  NAND2_X1 U11708 ( .A1(n11624), .A2(n11626), .ZN(n11685) );
  NAND2_X1 U11709 ( .A1(n11688), .A2(n11689), .ZN(n11626) );
  NAND3_X1 U11710 ( .A1(a_11_), .A2(n11690), .A3(b_13_), .ZN(n11689) );
  OR2_X1 U11711 ( .A1(n11622), .A2(n11620), .ZN(n11690) );
  NAND2_X1 U11712 ( .A1(n11620), .A2(n11622), .ZN(n11688) );
  NAND2_X1 U11713 ( .A1(n11691), .A2(n11692), .ZN(n11622) );
  NAND3_X1 U11714 ( .A1(a_12_), .A2(n11693), .A3(b_13_), .ZN(n11692) );
  OR2_X1 U11715 ( .A1(n11619), .A2(n11617), .ZN(n11693) );
  NAND2_X1 U11716 ( .A1(n11617), .A2(n11619), .ZN(n11691) );
  NAND2_X1 U11717 ( .A1(n11694), .A2(n11695), .ZN(n11619) );
  NAND2_X1 U11718 ( .A1(n11613), .A2(n11696), .ZN(n11695) );
  OR2_X1 U11719 ( .A1(n11614), .A2(n11615), .ZN(n11696) );
  XNOR2_X1 U11720 ( .A(n11697), .B(n11698), .ZN(n11613) );
  NAND2_X1 U11721 ( .A1(n11699), .A2(n11700), .ZN(n11697) );
  NAND2_X1 U11722 ( .A1(n11615), .A2(n11614), .ZN(n11694) );
  NAND2_X1 U11723 ( .A1(n11701), .A2(n11702), .ZN(n11614) );
  NAND3_X1 U11724 ( .A1(a_14_), .A2(n11703), .A3(b_13_), .ZN(n11702) );
  OR2_X1 U11725 ( .A1(n11493), .A2(n11492), .ZN(n11703) );
  NAND2_X1 U11726 ( .A1(n11492), .A2(n11493), .ZN(n11701) );
  NAND2_X1 U11727 ( .A1(n11704), .A2(n11705), .ZN(n11493) );
  NAND3_X1 U11728 ( .A1(a_15_), .A2(n11706), .A3(b_13_), .ZN(n11705) );
  OR2_X1 U11729 ( .A1(n11610), .A2(n11608), .ZN(n11706) );
  NAND2_X1 U11730 ( .A1(n11608), .A2(n11610), .ZN(n11704) );
  NAND2_X1 U11731 ( .A1(n11707), .A2(n11708), .ZN(n11610) );
  NAND3_X1 U11732 ( .A1(a_16_), .A2(n11709), .A3(b_13_), .ZN(n11708) );
  NAND2_X1 U11733 ( .A1(n11606), .A2(n11605), .ZN(n11709) );
  OR2_X1 U11734 ( .A1(n11605), .A2(n11606), .ZN(n11707) );
  AND2_X1 U11735 ( .A1(n11710), .A2(n11711), .ZN(n11606) );
  NAND3_X1 U11736 ( .A1(a_17_), .A2(n11712), .A3(b_13_), .ZN(n11711) );
  NAND2_X1 U11737 ( .A1(n11603), .A2(n11601), .ZN(n11712) );
  OR2_X1 U11738 ( .A1(n11601), .A2(n11603), .ZN(n11710) );
  AND2_X1 U11739 ( .A1(n11713), .A2(n11714), .ZN(n11603) );
  NAND2_X1 U11740 ( .A1(n11599), .A2(n11715), .ZN(n11714) );
  NAND2_X1 U11741 ( .A1(n11598), .A2(n11597), .ZN(n11715) );
  NOR2_X1 U11742 ( .A1(n11322), .A2(n7764), .ZN(n11599) );
  OR2_X1 U11743 ( .A1(n11597), .A2(n11598), .ZN(n11713) );
  AND2_X1 U11744 ( .A1(n11716), .A2(n11717), .ZN(n11598) );
  NAND2_X1 U11745 ( .A1(n11595), .A2(n11718), .ZN(n11717) );
  OR2_X1 U11746 ( .A1(n11594), .A2(n11592), .ZN(n11718) );
  NOR2_X1 U11747 ( .A1(n11322), .A2(n7902), .ZN(n11595) );
  NAND2_X1 U11748 ( .A1(n11592), .A2(n11594), .ZN(n11716) );
  NAND2_X1 U11749 ( .A1(n11719), .A2(n11720), .ZN(n11594) );
  NAND3_X1 U11750 ( .A1(a_20_), .A2(n11721), .A3(b_13_), .ZN(n11720) );
  NAND2_X1 U11751 ( .A1(n11590), .A2(n11589), .ZN(n11721) );
  OR2_X1 U11752 ( .A1(n11589), .A2(n11590), .ZN(n11719) );
  AND2_X1 U11753 ( .A1(n11722), .A2(n11723), .ZN(n11590) );
  NAND2_X1 U11754 ( .A1(n11587), .A2(n11724), .ZN(n11723) );
  OR2_X1 U11755 ( .A1(n11586), .A2(n11585), .ZN(n11724) );
  NOR2_X1 U11756 ( .A1(n11322), .A2(n7909), .ZN(n11587) );
  NAND2_X1 U11757 ( .A1(n11585), .A2(n11586), .ZN(n11722) );
  NAND2_X1 U11758 ( .A1(n11725), .A2(n11726), .ZN(n11586) );
  NAND3_X1 U11759 ( .A1(a_22_), .A2(n11727), .A3(b_13_), .ZN(n11726) );
  OR2_X1 U11760 ( .A1(n11582), .A2(n11580), .ZN(n11727) );
  NAND2_X1 U11761 ( .A1(n11580), .A2(n11582), .ZN(n11725) );
  NAND2_X1 U11762 ( .A1(n11728), .A2(n11729), .ZN(n11582) );
  NAND2_X1 U11763 ( .A1(n11579), .A2(n11730), .ZN(n11729) );
  OR2_X1 U11764 ( .A1(n11578), .A2(n11576), .ZN(n11730) );
  NOR2_X1 U11765 ( .A1(n11322), .A2(n7916), .ZN(n11579) );
  NAND2_X1 U11766 ( .A1(n11576), .A2(n11578), .ZN(n11728) );
  NAND2_X1 U11767 ( .A1(n11731), .A2(n11732), .ZN(n11578) );
  NAND3_X1 U11768 ( .A1(a_24_), .A2(n11733), .A3(b_13_), .ZN(n11732) );
  NAND2_X1 U11769 ( .A1(n11574), .A2(n11573), .ZN(n11733) );
  OR2_X1 U11770 ( .A1(n11573), .A2(n11574), .ZN(n11731) );
  AND2_X1 U11771 ( .A1(n11734), .A2(n11735), .ZN(n11574) );
  NAND2_X1 U11772 ( .A1(n11571), .A2(n11736), .ZN(n11735) );
  OR2_X1 U11773 ( .A1(n11570), .A2(n11569), .ZN(n11736) );
  NOR2_X1 U11774 ( .A1(n11322), .A2(n7923), .ZN(n11571) );
  NAND2_X1 U11775 ( .A1(n11569), .A2(n11570), .ZN(n11734) );
  NAND2_X1 U11776 ( .A1(n11566), .A2(n11737), .ZN(n11570) );
  NAND2_X1 U11777 ( .A1(n11565), .A2(n11567), .ZN(n11737) );
  NAND2_X1 U11778 ( .A1(n11738), .A2(n11739), .ZN(n11567) );
  NAND2_X1 U11779 ( .A1(b_13_), .A2(a_26_), .ZN(n11739) );
  INV_X1 U11780 ( .A(n11740), .ZN(n11738) );
  XNOR2_X1 U11781 ( .A(n11741), .B(n11742), .ZN(n11565) );
  NAND2_X1 U11782 ( .A1(n11743), .A2(n11744), .ZN(n11741) );
  NAND2_X1 U11783 ( .A1(a_26_), .A2(n11740), .ZN(n11566) );
  NAND2_X1 U11784 ( .A1(n11537), .A2(n11745), .ZN(n11740) );
  NAND2_X1 U11785 ( .A1(n11536), .A2(n11538), .ZN(n11745) );
  NAND2_X1 U11786 ( .A1(n11746), .A2(n11747), .ZN(n11538) );
  NAND2_X1 U11787 ( .A1(b_13_), .A2(a_27_), .ZN(n11747) );
  INV_X1 U11788 ( .A(n11748), .ZN(n11746) );
  XNOR2_X1 U11789 ( .A(n11749), .B(n11750), .ZN(n11536) );
  XOR2_X1 U11790 ( .A(n11751), .B(n11752), .Z(n11749) );
  NAND2_X1 U11791 ( .A1(b_12_), .A2(a_28_), .ZN(n11751) );
  NAND2_X1 U11792 ( .A1(a_27_), .A2(n11748), .ZN(n11537) );
  NAND2_X1 U11793 ( .A1(n11753), .A2(n11754), .ZN(n11748) );
  NAND3_X1 U11794 ( .A1(a_28_), .A2(n11755), .A3(b_13_), .ZN(n11754) );
  NAND2_X1 U11795 ( .A1(n11546), .A2(n11544), .ZN(n11755) );
  OR2_X1 U11796 ( .A1(n11544), .A2(n11546), .ZN(n11753) );
  AND2_X1 U11797 ( .A1(n11756), .A2(n11757), .ZN(n11546) );
  NAND2_X1 U11798 ( .A1(n11561), .A2(n11758), .ZN(n11757) );
  OR2_X1 U11799 ( .A1(n11562), .A2(n11563), .ZN(n11758) );
  NOR2_X1 U11800 ( .A1(n11322), .A2(n7946), .ZN(n11561) );
  NAND2_X1 U11801 ( .A1(n11563), .A2(n11562), .ZN(n11756) );
  NAND2_X1 U11802 ( .A1(n11759), .A2(n11760), .ZN(n11562) );
  NAND2_X1 U11803 ( .A1(b_11_), .A2(n11761), .ZN(n11760) );
  NAND2_X1 U11804 ( .A1(n7268), .A2(n11762), .ZN(n11761) );
  NAND2_X1 U11805 ( .A1(a_31_), .A2(n11559), .ZN(n11762) );
  NAND2_X1 U11806 ( .A1(b_12_), .A2(n11763), .ZN(n11759) );
  NAND2_X1 U11807 ( .A1(n7272), .A2(n11764), .ZN(n11763) );
  NAND2_X1 U11808 ( .A1(a_30_), .A2(n11765), .ZN(n11764) );
  AND3_X1 U11809 ( .A1(b_12_), .A2(n7954), .A3(b_13_), .ZN(n11563) );
  XNOR2_X1 U11810 ( .A(n11766), .B(n11767), .ZN(n11544) );
  XOR2_X1 U11811 ( .A(n11768), .B(n11769), .Z(n11766) );
  XNOR2_X1 U11812 ( .A(n11770), .B(n11771), .ZN(n11569) );
  NAND2_X1 U11813 ( .A1(n11772), .A2(n11773), .ZN(n11770) );
  XNOR2_X1 U11814 ( .A(n11774), .B(n11775), .ZN(n11573) );
  XOR2_X1 U11815 ( .A(n11776), .B(n11777), .Z(n11774) );
  XNOR2_X1 U11816 ( .A(n11778), .B(n11779), .ZN(n11576) );
  XNOR2_X1 U11817 ( .A(n11780), .B(n11781), .ZN(n11778) );
  NOR2_X1 U11818 ( .A1(n7691), .A2(n11559), .ZN(n11781) );
  XNOR2_X1 U11819 ( .A(n11782), .B(n11783), .ZN(n11580) );
  XNOR2_X1 U11820 ( .A(n11784), .B(n11785), .ZN(n11783) );
  XNOR2_X1 U11821 ( .A(n11786), .B(n11787), .ZN(n11585) );
  XOR2_X1 U11822 ( .A(n11788), .B(n11789), .Z(n11787) );
  NAND2_X1 U11823 ( .A1(b_12_), .A2(a_22_), .ZN(n11789) );
  XNOR2_X1 U11824 ( .A(n11790), .B(n11791), .ZN(n11589) );
  XOR2_X1 U11825 ( .A(n11792), .B(n11793), .Z(n11790) );
  XNOR2_X1 U11826 ( .A(n11794), .B(n11795), .ZN(n11592) );
  XNOR2_X1 U11827 ( .A(n11796), .B(n11797), .ZN(n11794) );
  NOR2_X1 U11828 ( .A1(n7987), .A2(n11559), .ZN(n11797) );
  XOR2_X1 U11829 ( .A(n11798), .B(n11799), .Z(n11597) );
  NAND2_X1 U11830 ( .A1(n11800), .A2(n11801), .ZN(n11798) );
  XNOR2_X1 U11831 ( .A(n11802), .B(n11803), .ZN(n11601) );
  XOR2_X1 U11832 ( .A(n11804), .B(n11805), .Z(n11802) );
  XNOR2_X1 U11833 ( .A(n11806), .B(n11807), .ZN(n11605) );
  XOR2_X1 U11834 ( .A(n11808), .B(n11809), .Z(n11806) );
  XNOR2_X1 U11835 ( .A(n11810), .B(n11811), .ZN(n11608) );
  XNOR2_X1 U11836 ( .A(n11812), .B(n11813), .ZN(n11810) );
  NOR2_X1 U11837 ( .A1(n7773), .A2(n11559), .ZN(n11813) );
  XNOR2_X1 U11838 ( .A(n11814), .B(n11815), .ZN(n11492) );
  NAND2_X1 U11839 ( .A1(n11816), .A2(n11817), .ZN(n11814) );
  XNOR2_X1 U11840 ( .A(n11818), .B(n11819), .ZN(n11617) );
  XNOR2_X1 U11841 ( .A(n11820), .B(n11821), .ZN(n11819) );
  XNOR2_X1 U11842 ( .A(n11822), .B(n11823), .ZN(n11620) );
  XNOR2_X1 U11843 ( .A(n11824), .B(n11825), .ZN(n11823) );
  XNOR2_X1 U11844 ( .A(n11826), .B(n11827), .ZN(n11624) );
  NAND2_X1 U11845 ( .A1(n11828), .A2(n11829), .ZN(n11826) );
  XOR2_X1 U11846 ( .A(n11830), .B(n11831), .Z(n11472) );
  NAND2_X1 U11847 ( .A1(n11832), .A2(n11833), .ZN(n11830) );
  XNOR2_X1 U11848 ( .A(n11834), .B(n11835), .ZN(n11463) );
  XNOR2_X1 U11849 ( .A(n11836), .B(n11837), .ZN(n11835) );
  XOR2_X1 U11850 ( .A(n11838), .B(n11839), .Z(n11455) );
  XOR2_X1 U11851 ( .A(n11840), .B(n11841), .Z(n11838) );
  NOR2_X1 U11852 ( .A1(n8037), .A2(n11559), .ZN(n11841) );
  XNOR2_X1 U11853 ( .A(n11842), .B(n11843), .ZN(n11447) );
  NAND2_X1 U11854 ( .A1(n11844), .A2(n11845), .ZN(n11842) );
  XNOR2_X1 U11855 ( .A(n11846), .B(n11847), .ZN(n11629) );
  XOR2_X1 U11856 ( .A(n11848), .B(n11849), .Z(n11846) );
  XNOR2_X1 U11857 ( .A(n11850), .B(n11851), .ZN(n11632) );
  XOR2_X1 U11858 ( .A(n11852), .B(n11853), .Z(n11851) );
  NAND2_X1 U11859 ( .A1(b_12_), .A2(a_5_), .ZN(n11853) );
  XNOR2_X1 U11860 ( .A(n11854), .B(n11855), .ZN(n11637) );
  XNOR2_X1 U11861 ( .A(n11856), .B(n11857), .ZN(n11854) );
  XOR2_X1 U11862 ( .A(n11858), .B(n11859), .Z(n11640) );
  XOR2_X1 U11863 ( .A(n11860), .B(n11861), .Z(n11858) );
  NOR2_X1 U11864 ( .A1(n7850), .A2(n11559), .ZN(n11861) );
  XNOR2_X1 U11865 ( .A(n11862), .B(n11863), .ZN(n11645) );
  XNOR2_X1 U11866 ( .A(n11864), .B(n11865), .ZN(n11863) );
  XNOR2_X1 U11867 ( .A(n11866), .B(n11867), .ZN(n11650) );
  XNOR2_X1 U11868 ( .A(n11868), .B(n11869), .ZN(n11866) );
  XOR2_X1 U11869 ( .A(n11870), .B(n11871), .Z(n11649) );
  XNOR2_X1 U11870 ( .A(n11872), .B(n11873), .ZN(n11870) );
  NAND4_X1 U11871 ( .A1(n7530), .A2(n7529), .A3(n7525), .A4(n7531), .ZN(n7504)
         );
  NAND2_X1 U11872 ( .A1(n11874), .A2(n11875), .ZN(n7531) );
  NAND2_X1 U11873 ( .A1(n11873), .A2(n11876), .ZN(n11875) );
  NAND2_X1 U11874 ( .A1(n11872), .A2(n11871), .ZN(n11876) );
  NOR2_X1 U11875 ( .A1(n11559), .A2(n7613), .ZN(n11873) );
  OR2_X1 U11876 ( .A1(n11871), .A2(n11872), .ZN(n11874) );
  AND2_X1 U11877 ( .A1(n11877), .A2(n11878), .ZN(n11872) );
  NAND2_X1 U11878 ( .A1(n11869), .A2(n11879), .ZN(n11878) );
  NAND2_X1 U11879 ( .A1(n11868), .A2(n11867), .ZN(n11879) );
  NOR2_X1 U11880 ( .A1(n11559), .A2(n7411), .ZN(n11869) );
  OR2_X1 U11881 ( .A1(n11867), .A2(n11868), .ZN(n11877) );
  AND2_X1 U11882 ( .A1(n11880), .A2(n11881), .ZN(n11868) );
  NAND2_X1 U11883 ( .A1(n11865), .A2(n11882), .ZN(n11881) );
  OR2_X1 U11884 ( .A1(n11864), .A2(n11862), .ZN(n11882) );
  NOR2_X1 U11885 ( .A1(n11559), .A2(n7832), .ZN(n11865) );
  NAND2_X1 U11886 ( .A1(n11862), .A2(n11864), .ZN(n11880) );
  NAND2_X1 U11887 ( .A1(n11883), .A2(n11884), .ZN(n11864) );
  NAND3_X1 U11888 ( .A1(a_3_), .A2(n11885), .A3(b_12_), .ZN(n11884) );
  OR2_X1 U11889 ( .A1(n11860), .A2(n11859), .ZN(n11885) );
  NAND2_X1 U11890 ( .A1(n11859), .A2(n11860), .ZN(n11883) );
  NAND2_X1 U11891 ( .A1(n11886), .A2(n11887), .ZN(n11860) );
  NAND2_X1 U11892 ( .A1(n11857), .A2(n11888), .ZN(n11887) );
  NAND2_X1 U11893 ( .A1(n11856), .A2(n11855), .ZN(n11888) );
  NOR2_X1 U11894 ( .A1(n11559), .A2(n7398), .ZN(n11857) );
  OR2_X1 U11895 ( .A1(n11855), .A2(n11856), .ZN(n11886) );
  AND2_X1 U11896 ( .A1(n11889), .A2(n11890), .ZN(n11856) );
  NAND3_X1 U11897 ( .A1(a_5_), .A2(n11891), .A3(b_12_), .ZN(n11890) );
  OR2_X1 U11898 ( .A1(n11852), .A2(n11850), .ZN(n11891) );
  NAND2_X1 U11899 ( .A1(n11850), .A2(n11852), .ZN(n11889) );
  NAND2_X1 U11900 ( .A1(n11892), .A2(n11893), .ZN(n11852) );
  NAND2_X1 U11901 ( .A1(n11848), .A2(n11894), .ZN(n11893) );
  OR2_X1 U11902 ( .A1(n11849), .A2(n11847), .ZN(n11894) );
  NOR2_X1 U11903 ( .A1(n11559), .A2(n7388), .ZN(n11848) );
  NAND2_X1 U11904 ( .A1(n11847), .A2(n11849), .ZN(n11892) );
  NAND2_X1 U11905 ( .A1(n11844), .A2(n11895), .ZN(n11849) );
  NAND2_X1 U11906 ( .A1(n11843), .A2(n11845), .ZN(n11895) );
  NAND2_X1 U11907 ( .A1(n11896), .A2(n11897), .ZN(n11845) );
  NAND2_X1 U11908 ( .A1(b_12_), .A2(a_7_), .ZN(n11897) );
  INV_X1 U11909 ( .A(n11898), .ZN(n11896) );
  XNOR2_X1 U11910 ( .A(n11899), .B(n11900), .ZN(n11843) );
  XOR2_X1 U11911 ( .A(n11901), .B(n11902), .Z(n11900) );
  NAND2_X1 U11912 ( .A1(b_11_), .A2(a_8_), .ZN(n11902) );
  NAND2_X1 U11913 ( .A1(a_7_), .A2(n11898), .ZN(n11844) );
  NAND2_X1 U11914 ( .A1(n11903), .A2(n11904), .ZN(n11898) );
  NAND3_X1 U11915 ( .A1(a_8_), .A2(n11905), .A3(b_12_), .ZN(n11904) );
  OR2_X1 U11916 ( .A1(n11840), .A2(n11839), .ZN(n11905) );
  NAND2_X1 U11917 ( .A1(n11839), .A2(n11840), .ZN(n11903) );
  NAND2_X1 U11918 ( .A1(n11906), .A2(n11907), .ZN(n11840) );
  NAND2_X1 U11919 ( .A1(n11837), .A2(n11908), .ZN(n11907) );
  OR2_X1 U11920 ( .A1(n11836), .A2(n11834), .ZN(n11908) );
  NOR2_X1 U11921 ( .A1(n11559), .A2(n7870), .ZN(n11837) );
  NAND2_X1 U11922 ( .A1(n11834), .A2(n11836), .ZN(n11906) );
  NAND2_X1 U11923 ( .A1(n11832), .A2(n11909), .ZN(n11836) );
  NAND2_X1 U11924 ( .A1(n11831), .A2(n11833), .ZN(n11909) );
  NAND2_X1 U11925 ( .A1(n11910), .A2(n11911), .ZN(n11833) );
  NAND2_X1 U11926 ( .A1(b_12_), .A2(a_10_), .ZN(n11911) );
  INV_X1 U11927 ( .A(n11912), .ZN(n11910) );
  XOR2_X1 U11928 ( .A(n11913), .B(n11914), .Z(n11831) );
  XOR2_X1 U11929 ( .A(n11915), .B(n11916), .Z(n11913) );
  NAND2_X1 U11930 ( .A1(a_10_), .A2(n11912), .ZN(n11832) );
  NAND2_X1 U11931 ( .A1(n11828), .A2(n11917), .ZN(n11912) );
  NAND2_X1 U11932 ( .A1(n11827), .A2(n11829), .ZN(n11917) );
  NAND2_X1 U11933 ( .A1(n11918), .A2(n11919), .ZN(n11829) );
  NAND2_X1 U11934 ( .A1(b_12_), .A2(a_11_), .ZN(n11919) );
  INV_X1 U11935 ( .A(n11920), .ZN(n11918) );
  XOR2_X1 U11936 ( .A(n11921), .B(n11922), .Z(n11827) );
  XOR2_X1 U11937 ( .A(n11923), .B(n11924), .Z(n11921) );
  NOR2_X1 U11938 ( .A1(n8020), .A2(n11765), .ZN(n11924) );
  NAND2_X1 U11939 ( .A1(a_11_), .A2(n11920), .ZN(n11828) );
  NAND2_X1 U11940 ( .A1(n11925), .A2(n11926), .ZN(n11920) );
  NAND2_X1 U11941 ( .A1(n11824), .A2(n11927), .ZN(n11926) );
  OR2_X1 U11942 ( .A1(n11825), .A2(n11822), .ZN(n11927) );
  NAND2_X1 U11943 ( .A1(n11822), .A2(n11825), .ZN(n11925) );
  NAND2_X1 U11944 ( .A1(n11928), .A2(n11929), .ZN(n11825) );
  NAND2_X1 U11945 ( .A1(n11821), .A2(n11930), .ZN(n11929) );
  OR2_X1 U11946 ( .A1(n11820), .A2(n11818), .ZN(n11930) );
  NOR2_X1 U11947 ( .A1(n11559), .A2(n7355), .ZN(n11821) );
  NAND2_X1 U11948 ( .A1(n11818), .A2(n11820), .ZN(n11928) );
  NAND2_X1 U11949 ( .A1(n11699), .A2(n11931), .ZN(n11820) );
  NAND2_X1 U11950 ( .A1(n11698), .A2(n11700), .ZN(n11931) );
  NAND2_X1 U11951 ( .A1(n11932), .A2(n11933), .ZN(n11700) );
  NAND2_X1 U11952 ( .A1(b_12_), .A2(a_14_), .ZN(n11933) );
  INV_X1 U11953 ( .A(n11934), .ZN(n11932) );
  XNOR2_X1 U11954 ( .A(n11935), .B(n11936), .ZN(n11698) );
  XOR2_X1 U11955 ( .A(n11937), .B(n11938), .Z(n11936) );
  NAND2_X1 U11956 ( .A1(b_11_), .A2(a_15_), .ZN(n11938) );
  NAND2_X1 U11957 ( .A1(a_14_), .A2(n11934), .ZN(n11699) );
  NAND2_X1 U11958 ( .A1(n11816), .A2(n11939), .ZN(n11934) );
  NAND2_X1 U11959 ( .A1(n11815), .A2(n11817), .ZN(n11939) );
  NAND2_X1 U11960 ( .A1(n11940), .A2(n11941), .ZN(n11817) );
  NAND2_X1 U11961 ( .A1(b_12_), .A2(a_15_), .ZN(n11941) );
  INV_X1 U11962 ( .A(n11942), .ZN(n11940) );
  XNOR2_X1 U11963 ( .A(n11943), .B(n11944), .ZN(n11815) );
  XNOR2_X1 U11964 ( .A(n11945), .B(n11946), .ZN(n11943) );
  NOR2_X1 U11965 ( .A1(n7773), .A2(n11765), .ZN(n11946) );
  NAND2_X1 U11966 ( .A1(a_15_), .A2(n11942), .ZN(n11816) );
  NAND2_X1 U11967 ( .A1(n11947), .A2(n11948), .ZN(n11942) );
  NAND3_X1 U11968 ( .A1(a_16_), .A2(n11949), .A3(b_12_), .ZN(n11948) );
  NAND2_X1 U11969 ( .A1(n11812), .A2(n11811), .ZN(n11949) );
  OR2_X1 U11970 ( .A1(n11811), .A2(n11812), .ZN(n11947) );
  AND2_X1 U11971 ( .A1(n11950), .A2(n11951), .ZN(n11812) );
  NAND2_X1 U11972 ( .A1(n11808), .A2(n11952), .ZN(n11951) );
  OR2_X1 U11973 ( .A1(n11809), .A2(n11807), .ZN(n11952) );
  NOR2_X1 U11974 ( .A1(n11559), .A2(n7337), .ZN(n11808) );
  NAND2_X1 U11975 ( .A1(n11807), .A2(n11809), .ZN(n11950) );
  NAND2_X1 U11976 ( .A1(n11953), .A2(n11954), .ZN(n11809) );
  NAND2_X1 U11977 ( .A1(n11804), .A2(n11955), .ZN(n11954) );
  OR2_X1 U11978 ( .A1(n11805), .A2(n11803), .ZN(n11955) );
  NOR2_X1 U11979 ( .A1(n11559), .A2(n7764), .ZN(n11804) );
  NAND2_X1 U11980 ( .A1(n11803), .A2(n11805), .ZN(n11953) );
  NAND2_X1 U11981 ( .A1(n11800), .A2(n11956), .ZN(n11805) );
  NAND2_X1 U11982 ( .A1(n11799), .A2(n11801), .ZN(n11956) );
  NAND2_X1 U11983 ( .A1(n11957), .A2(n11958), .ZN(n11801) );
  NAND2_X1 U11984 ( .A1(b_12_), .A2(a_19_), .ZN(n11958) );
  INV_X1 U11985 ( .A(n11959), .ZN(n11957) );
  XOR2_X1 U11986 ( .A(n11960), .B(n11961), .Z(n11799) );
  XOR2_X1 U11987 ( .A(n11962), .B(n11963), .Z(n11960) );
  NOR2_X1 U11988 ( .A1(n7987), .A2(n11765), .ZN(n11963) );
  NAND2_X1 U11989 ( .A1(a_19_), .A2(n11959), .ZN(n11800) );
  NAND2_X1 U11990 ( .A1(n11964), .A2(n11965), .ZN(n11959) );
  NAND3_X1 U11991 ( .A1(a_20_), .A2(n11966), .A3(b_12_), .ZN(n11965) );
  NAND2_X1 U11992 ( .A1(n11796), .A2(n11795), .ZN(n11966) );
  OR2_X1 U11993 ( .A1(n11795), .A2(n11796), .ZN(n11964) );
  AND2_X1 U11994 ( .A1(n11967), .A2(n11968), .ZN(n11796) );
  NAND2_X1 U11995 ( .A1(n11793), .A2(n11969), .ZN(n11968) );
  OR2_X1 U11996 ( .A1(n11792), .A2(n11791), .ZN(n11969) );
  NOR2_X1 U11997 ( .A1(n11559), .A2(n7909), .ZN(n11793) );
  NAND2_X1 U11998 ( .A1(n11791), .A2(n11792), .ZN(n11967) );
  NAND2_X1 U11999 ( .A1(n11970), .A2(n11971), .ZN(n11792) );
  NAND3_X1 U12000 ( .A1(a_22_), .A2(n11972), .A3(b_12_), .ZN(n11971) );
  OR2_X1 U12001 ( .A1(n11788), .A2(n11786), .ZN(n11972) );
  NAND2_X1 U12002 ( .A1(n11786), .A2(n11788), .ZN(n11970) );
  NAND2_X1 U12003 ( .A1(n11973), .A2(n11974), .ZN(n11788) );
  NAND2_X1 U12004 ( .A1(n11785), .A2(n11975), .ZN(n11974) );
  OR2_X1 U12005 ( .A1(n11784), .A2(n11782), .ZN(n11975) );
  NOR2_X1 U12006 ( .A1(n11559), .A2(n7916), .ZN(n11785) );
  NAND2_X1 U12007 ( .A1(n11782), .A2(n11784), .ZN(n11973) );
  NAND2_X1 U12008 ( .A1(n11976), .A2(n11977), .ZN(n11784) );
  NAND3_X1 U12009 ( .A1(a_24_), .A2(n11978), .A3(b_12_), .ZN(n11977) );
  NAND2_X1 U12010 ( .A1(n11780), .A2(n11779), .ZN(n11978) );
  OR2_X1 U12011 ( .A1(n11779), .A2(n11780), .ZN(n11976) );
  AND2_X1 U12012 ( .A1(n11979), .A2(n11980), .ZN(n11780) );
  NAND2_X1 U12013 ( .A1(n11777), .A2(n11981), .ZN(n11980) );
  OR2_X1 U12014 ( .A1(n11776), .A2(n11775), .ZN(n11981) );
  NOR2_X1 U12015 ( .A1(n11559), .A2(n7923), .ZN(n11777) );
  NAND2_X1 U12016 ( .A1(n11775), .A2(n11776), .ZN(n11979) );
  NAND2_X1 U12017 ( .A1(n11772), .A2(n11982), .ZN(n11776) );
  NAND2_X1 U12018 ( .A1(n11771), .A2(n11773), .ZN(n11982) );
  NAND2_X1 U12019 ( .A1(n11983), .A2(n11984), .ZN(n11773) );
  NAND2_X1 U12020 ( .A1(b_12_), .A2(a_26_), .ZN(n11984) );
  INV_X1 U12021 ( .A(n11985), .ZN(n11983) );
  XNOR2_X1 U12022 ( .A(n11986), .B(n11987), .ZN(n11771) );
  NAND2_X1 U12023 ( .A1(n11988), .A2(n11989), .ZN(n11986) );
  NAND2_X1 U12024 ( .A1(a_26_), .A2(n11985), .ZN(n11772) );
  NAND2_X1 U12025 ( .A1(n11743), .A2(n11990), .ZN(n11985) );
  NAND2_X1 U12026 ( .A1(n11742), .A2(n11744), .ZN(n11990) );
  NAND2_X1 U12027 ( .A1(n11991), .A2(n11992), .ZN(n11744) );
  NAND2_X1 U12028 ( .A1(b_12_), .A2(a_27_), .ZN(n11992) );
  INV_X1 U12029 ( .A(n11993), .ZN(n11991) );
  XNOR2_X1 U12030 ( .A(n11994), .B(n11995), .ZN(n11742) );
  XOR2_X1 U12031 ( .A(n11996), .B(n11997), .Z(n11994) );
  NAND2_X1 U12032 ( .A1(b_11_), .A2(a_28_), .ZN(n11996) );
  NAND2_X1 U12033 ( .A1(a_27_), .A2(n11993), .ZN(n11743) );
  NAND2_X1 U12034 ( .A1(n11998), .A2(n11999), .ZN(n11993) );
  NAND3_X1 U12035 ( .A1(a_28_), .A2(n12000), .A3(b_12_), .ZN(n11999) );
  NAND2_X1 U12036 ( .A1(n11752), .A2(n11750), .ZN(n12000) );
  OR2_X1 U12037 ( .A1(n11750), .A2(n11752), .ZN(n11998) );
  AND2_X1 U12038 ( .A1(n12001), .A2(n12002), .ZN(n11752) );
  NAND2_X1 U12039 ( .A1(n11767), .A2(n12003), .ZN(n12002) );
  OR2_X1 U12040 ( .A1(n11768), .A2(n11769), .ZN(n12003) );
  NOR2_X1 U12041 ( .A1(n11559), .A2(n7946), .ZN(n11767) );
  NAND2_X1 U12042 ( .A1(n11769), .A2(n11768), .ZN(n12001) );
  NAND2_X1 U12043 ( .A1(n12004), .A2(n12005), .ZN(n11768) );
  NAND2_X1 U12044 ( .A1(b_10_), .A2(n12006), .ZN(n12005) );
  NAND2_X1 U12045 ( .A1(n7268), .A2(n12007), .ZN(n12006) );
  NAND2_X1 U12046 ( .A1(a_31_), .A2(n11765), .ZN(n12007) );
  NAND2_X1 U12047 ( .A1(b_11_), .A2(n12008), .ZN(n12004) );
  NAND2_X1 U12048 ( .A1(n7272), .A2(n12009), .ZN(n12008) );
  NAND2_X1 U12049 ( .A1(a_30_), .A2(n12010), .ZN(n12009) );
  AND3_X1 U12050 ( .A1(b_11_), .A2(n7954), .A3(b_12_), .ZN(n11769) );
  XNOR2_X1 U12051 ( .A(n12011), .B(n12012), .ZN(n11750) );
  XOR2_X1 U12052 ( .A(n12013), .B(n12014), .Z(n12011) );
  XNOR2_X1 U12053 ( .A(n12015), .B(n12016), .ZN(n11775) );
  NAND2_X1 U12054 ( .A1(n12017), .A2(n12018), .ZN(n12015) );
  XNOR2_X1 U12055 ( .A(n12019), .B(n12020), .ZN(n11779) );
  XOR2_X1 U12056 ( .A(n12021), .B(n12022), .Z(n12019) );
  XNOR2_X1 U12057 ( .A(n12023), .B(n12024), .ZN(n11782) );
  XNOR2_X1 U12058 ( .A(n12025), .B(n12026), .ZN(n12023) );
  NOR2_X1 U12059 ( .A1(n7691), .A2(n11765), .ZN(n12026) );
  XNOR2_X1 U12060 ( .A(n12027), .B(n12028), .ZN(n11786) );
  XNOR2_X1 U12061 ( .A(n12029), .B(n12030), .ZN(n12028) );
  XNOR2_X1 U12062 ( .A(n12031), .B(n12032), .ZN(n11791) );
  XOR2_X1 U12063 ( .A(n12033), .B(n12034), .Z(n12032) );
  NAND2_X1 U12064 ( .A1(b_11_), .A2(a_22_), .ZN(n12034) );
  XNOR2_X1 U12065 ( .A(n12035), .B(n12036), .ZN(n11795) );
  XOR2_X1 U12066 ( .A(n12037), .B(n12038), .Z(n12035) );
  XNOR2_X1 U12067 ( .A(n12039), .B(n12040), .ZN(n11803) );
  NAND2_X1 U12068 ( .A1(n12041), .A2(n12042), .ZN(n12039) );
  XNOR2_X1 U12069 ( .A(n12043), .B(n12044), .ZN(n11807) );
  NAND2_X1 U12070 ( .A1(n12045), .A2(n12046), .ZN(n12043) );
  XOR2_X1 U12071 ( .A(n12047), .B(n12048), .Z(n11811) );
  XOR2_X1 U12072 ( .A(n12049), .B(n12050), .Z(n12048) );
  NAND2_X1 U12073 ( .A1(b_11_), .A2(a_17_), .ZN(n12050) );
  XOR2_X1 U12074 ( .A(n12051), .B(n12052), .Z(n11818) );
  XOR2_X1 U12075 ( .A(n12053), .B(n12054), .Z(n12051) );
  NOR2_X1 U12076 ( .A1(n7782), .A2(n11765), .ZN(n12054) );
  XNOR2_X1 U12077 ( .A(n12055), .B(n12056), .ZN(n11822) );
  XOR2_X1 U12078 ( .A(n12057), .B(n12058), .Z(n12056) );
  NAND2_X1 U12079 ( .A1(b_11_), .A2(a_13_), .ZN(n12058) );
  XNOR2_X1 U12080 ( .A(n12059), .B(n12060), .ZN(n11834) );
  XNOR2_X1 U12081 ( .A(n12061), .B(n12062), .ZN(n12059) );
  NOR2_X1 U12082 ( .A1(n7799), .A2(n11765), .ZN(n12062) );
  XNOR2_X1 U12083 ( .A(n12063), .B(n12064), .ZN(n11839) );
  XNOR2_X1 U12084 ( .A(n12065), .B(n12066), .ZN(n12063) );
  NOR2_X1 U12085 ( .A1(n7870), .A2(n11765), .ZN(n12066) );
  XNOR2_X1 U12086 ( .A(n12067), .B(n12068), .ZN(n11847) );
  XNOR2_X1 U12087 ( .A(n12069), .B(n12070), .ZN(n12067) );
  NOR2_X1 U12088 ( .A1(n7863), .A2(n11765), .ZN(n12070) );
  XNOR2_X1 U12089 ( .A(n12071), .B(n12072), .ZN(n11850) );
  XOR2_X1 U12090 ( .A(n12073), .B(n12074), .Z(n12072) );
  NAND2_X1 U12091 ( .A1(b_11_), .A2(a_6_), .ZN(n12074) );
  XNOR2_X1 U12092 ( .A(n12075), .B(n12076), .ZN(n11855) );
  XOR2_X1 U12093 ( .A(n12077), .B(n12078), .Z(n12075) );
  NOR2_X1 U12094 ( .A1(n7393), .A2(n11765), .ZN(n12078) );
  XNOR2_X1 U12095 ( .A(n12079), .B(n12080), .ZN(n11859) );
  XNOR2_X1 U12096 ( .A(n12081), .B(n12082), .ZN(n12079) );
  NOR2_X1 U12097 ( .A1(n7398), .A2(n11765), .ZN(n12082) );
  XNOR2_X1 U12098 ( .A(n12083), .B(n12084), .ZN(n11862) );
  XOR2_X1 U12099 ( .A(n12085), .B(n12086), .Z(n12084) );
  NAND2_X1 U12100 ( .A1(b_11_), .A2(a_3_), .ZN(n12086) );
  XOR2_X1 U12101 ( .A(n12087), .B(n12088), .Z(n11867) );
  XOR2_X1 U12102 ( .A(n12089), .B(n12090), .Z(n12088) );
  NAND2_X1 U12103 ( .A1(b_11_), .A2(a_2_), .ZN(n12090) );
  XOR2_X1 U12104 ( .A(n12091), .B(n12092), .Z(n11871) );
  XOR2_X1 U12105 ( .A(n12093), .B(n12094), .Z(n12092) );
  NAND2_X1 U12106 ( .A1(b_11_), .A2(a_1_), .ZN(n12094) );
  NAND3_X1 U12107 ( .A1(n12095), .A2(n12096), .A3(n12097), .ZN(n7529) );
  XOR2_X1 U12108 ( .A(n12098), .B(n12099), .Z(n12097) );
  XOR2_X1 U12109 ( .A(n12100), .B(n12101), .Z(n7530) );
  XOR2_X1 U12110 ( .A(n12102), .B(n12103), .Z(n12100) );
  OR2_X1 U12111 ( .A1(n7525), .A2(n7524), .ZN(n7508) );
  XNOR2_X1 U12112 ( .A(n12104), .B(n12105), .ZN(n7524) );
  NAND2_X1 U12113 ( .A1(n12106), .A2(n12107), .ZN(n7525) );
  NAND2_X1 U12114 ( .A1(n12095), .A2(n12096), .ZN(n12107) );
  NAND2_X1 U12115 ( .A1(n12103), .A2(n12108), .ZN(n12096) );
  OR2_X1 U12116 ( .A1(n12102), .A2(n12101), .ZN(n12108) );
  NOR2_X1 U12117 ( .A1(n11765), .A2(n7613), .ZN(n12103) );
  NAND2_X1 U12118 ( .A1(n12101), .A2(n12102), .ZN(n12095) );
  NAND2_X1 U12119 ( .A1(n12109), .A2(n12110), .ZN(n12102) );
  NAND3_X1 U12120 ( .A1(a_1_), .A2(n12111), .A3(b_11_), .ZN(n12110) );
  OR2_X1 U12121 ( .A1(n12093), .A2(n12091), .ZN(n12111) );
  NAND2_X1 U12122 ( .A1(n12091), .A2(n12093), .ZN(n12109) );
  NAND2_X1 U12123 ( .A1(n12112), .A2(n12113), .ZN(n12093) );
  NAND3_X1 U12124 ( .A1(a_2_), .A2(n12114), .A3(b_11_), .ZN(n12113) );
  OR2_X1 U12125 ( .A1(n12089), .A2(n12087), .ZN(n12114) );
  NAND2_X1 U12126 ( .A1(n12087), .A2(n12089), .ZN(n12112) );
  NAND2_X1 U12127 ( .A1(n12115), .A2(n12116), .ZN(n12089) );
  NAND3_X1 U12128 ( .A1(a_3_), .A2(n12117), .A3(b_11_), .ZN(n12116) );
  OR2_X1 U12129 ( .A1(n12085), .A2(n12083), .ZN(n12117) );
  NAND2_X1 U12130 ( .A1(n12083), .A2(n12085), .ZN(n12115) );
  NAND2_X1 U12131 ( .A1(n12118), .A2(n12119), .ZN(n12085) );
  NAND3_X1 U12132 ( .A1(a_4_), .A2(n12120), .A3(b_11_), .ZN(n12119) );
  NAND2_X1 U12133 ( .A1(n12081), .A2(n12080), .ZN(n12120) );
  OR2_X1 U12134 ( .A1(n12080), .A2(n12081), .ZN(n12118) );
  AND2_X1 U12135 ( .A1(n12121), .A2(n12122), .ZN(n12081) );
  NAND3_X1 U12136 ( .A1(a_5_), .A2(n12123), .A3(b_11_), .ZN(n12122) );
  OR2_X1 U12137 ( .A1(n12077), .A2(n12076), .ZN(n12123) );
  NAND2_X1 U12138 ( .A1(n12076), .A2(n12077), .ZN(n12121) );
  NAND2_X1 U12139 ( .A1(n12124), .A2(n12125), .ZN(n12077) );
  NAND3_X1 U12140 ( .A1(a_6_), .A2(n12126), .A3(b_11_), .ZN(n12125) );
  OR2_X1 U12141 ( .A1(n12073), .A2(n12071), .ZN(n12126) );
  NAND2_X1 U12142 ( .A1(n12071), .A2(n12073), .ZN(n12124) );
  NAND2_X1 U12143 ( .A1(n12127), .A2(n12128), .ZN(n12073) );
  NAND3_X1 U12144 ( .A1(a_7_), .A2(n12129), .A3(b_11_), .ZN(n12128) );
  NAND2_X1 U12145 ( .A1(n12069), .A2(n12068), .ZN(n12129) );
  OR2_X1 U12146 ( .A1(n12068), .A2(n12069), .ZN(n12127) );
  AND2_X1 U12147 ( .A1(n12130), .A2(n12131), .ZN(n12069) );
  NAND3_X1 U12148 ( .A1(a_8_), .A2(n12132), .A3(b_11_), .ZN(n12131) );
  OR2_X1 U12149 ( .A1(n11901), .A2(n11899), .ZN(n12132) );
  NAND2_X1 U12150 ( .A1(n11899), .A2(n11901), .ZN(n12130) );
  NAND2_X1 U12151 ( .A1(n12133), .A2(n12134), .ZN(n11901) );
  NAND3_X1 U12152 ( .A1(a_9_), .A2(n12135), .A3(b_11_), .ZN(n12134) );
  NAND2_X1 U12153 ( .A1(n12065), .A2(n12064), .ZN(n12135) );
  OR2_X1 U12154 ( .A1(n12064), .A2(n12065), .ZN(n12133) );
  AND2_X1 U12155 ( .A1(n12136), .A2(n12137), .ZN(n12065) );
  NAND3_X1 U12156 ( .A1(a_10_), .A2(n12138), .A3(b_11_), .ZN(n12137) );
  NAND2_X1 U12157 ( .A1(n12061), .A2(n12060), .ZN(n12138) );
  OR2_X1 U12158 ( .A1(n12060), .A2(n12061), .ZN(n12136) );
  AND2_X1 U12159 ( .A1(n12139), .A2(n12140), .ZN(n12061) );
  NAND2_X1 U12160 ( .A1(n11914), .A2(n12141), .ZN(n12140) );
  OR2_X1 U12161 ( .A1(n11915), .A2(n11916), .ZN(n12141) );
  XNOR2_X1 U12162 ( .A(n12142), .B(n12143), .ZN(n11914) );
  NAND2_X1 U12163 ( .A1(n12144), .A2(n12145), .ZN(n12142) );
  NAND2_X1 U12164 ( .A1(n11916), .A2(n11915), .ZN(n12139) );
  NAND2_X1 U12165 ( .A1(n12146), .A2(n12147), .ZN(n11915) );
  NAND3_X1 U12166 ( .A1(a_12_), .A2(n12148), .A3(b_11_), .ZN(n12147) );
  OR2_X1 U12167 ( .A1(n11923), .A2(n11922), .ZN(n12148) );
  NAND2_X1 U12168 ( .A1(n11922), .A2(n11923), .ZN(n12146) );
  NAND2_X1 U12169 ( .A1(n12149), .A2(n12150), .ZN(n11923) );
  NAND3_X1 U12170 ( .A1(a_13_), .A2(n12151), .A3(b_11_), .ZN(n12150) );
  OR2_X1 U12171 ( .A1(n12057), .A2(n12055), .ZN(n12151) );
  NAND2_X1 U12172 ( .A1(n12055), .A2(n12057), .ZN(n12149) );
  NAND2_X1 U12173 ( .A1(n12152), .A2(n12153), .ZN(n12057) );
  NAND3_X1 U12174 ( .A1(a_14_), .A2(n12154), .A3(b_11_), .ZN(n12153) );
  OR2_X1 U12175 ( .A1(n12053), .A2(n12052), .ZN(n12154) );
  NAND2_X1 U12176 ( .A1(n12052), .A2(n12053), .ZN(n12152) );
  NAND2_X1 U12177 ( .A1(n12155), .A2(n12156), .ZN(n12053) );
  NAND3_X1 U12178 ( .A1(a_15_), .A2(n12157), .A3(b_11_), .ZN(n12156) );
  OR2_X1 U12179 ( .A1(n11937), .A2(n11935), .ZN(n12157) );
  NAND2_X1 U12180 ( .A1(n11935), .A2(n11937), .ZN(n12155) );
  NAND2_X1 U12181 ( .A1(n12158), .A2(n12159), .ZN(n11937) );
  NAND3_X1 U12182 ( .A1(a_16_), .A2(n12160), .A3(b_11_), .ZN(n12159) );
  NAND2_X1 U12183 ( .A1(n11945), .A2(n11944), .ZN(n12160) );
  OR2_X1 U12184 ( .A1(n11944), .A2(n11945), .ZN(n12158) );
  AND2_X1 U12185 ( .A1(n12161), .A2(n12162), .ZN(n11945) );
  NAND3_X1 U12186 ( .A1(a_17_), .A2(n12163), .A3(b_11_), .ZN(n12162) );
  OR2_X1 U12187 ( .A1(n12049), .A2(n12047), .ZN(n12163) );
  NAND2_X1 U12188 ( .A1(n12047), .A2(n12049), .ZN(n12161) );
  NAND2_X1 U12189 ( .A1(n12045), .A2(n12164), .ZN(n12049) );
  NAND2_X1 U12190 ( .A1(n12044), .A2(n12046), .ZN(n12164) );
  NAND2_X1 U12191 ( .A1(n12165), .A2(n12166), .ZN(n12046) );
  NAND2_X1 U12192 ( .A1(b_11_), .A2(a_18_), .ZN(n12166) );
  INV_X1 U12193 ( .A(n12167), .ZN(n12165) );
  XNOR2_X1 U12194 ( .A(n12168), .B(n12169), .ZN(n12044) );
  XNOR2_X1 U12195 ( .A(n12170), .B(n12171), .ZN(n12169) );
  NAND2_X1 U12196 ( .A1(a_18_), .A2(n12167), .ZN(n12045) );
  NAND2_X1 U12197 ( .A1(n12041), .A2(n12172), .ZN(n12167) );
  NAND2_X1 U12198 ( .A1(n12040), .A2(n12042), .ZN(n12172) );
  NAND2_X1 U12199 ( .A1(n12173), .A2(n12174), .ZN(n12042) );
  NAND2_X1 U12200 ( .A1(b_11_), .A2(a_19_), .ZN(n12174) );
  INV_X1 U12201 ( .A(n12175), .ZN(n12173) );
  XNOR2_X1 U12202 ( .A(n12176), .B(n12177), .ZN(n12040) );
  XNOR2_X1 U12203 ( .A(n12178), .B(n12179), .ZN(n12177) );
  NAND2_X1 U12204 ( .A1(a_19_), .A2(n12175), .ZN(n12041) );
  NAND2_X1 U12205 ( .A1(n12180), .A2(n12181), .ZN(n12175) );
  NAND3_X1 U12206 ( .A1(a_20_), .A2(n12182), .A3(b_11_), .ZN(n12181) );
  OR2_X1 U12207 ( .A1(n11962), .A2(n11961), .ZN(n12182) );
  NAND2_X1 U12208 ( .A1(n11961), .A2(n11962), .ZN(n12180) );
  NAND2_X1 U12209 ( .A1(n12183), .A2(n12184), .ZN(n11962) );
  NAND2_X1 U12210 ( .A1(n12038), .A2(n12185), .ZN(n12184) );
  OR2_X1 U12211 ( .A1(n12037), .A2(n12036), .ZN(n12185) );
  NOR2_X1 U12212 ( .A1(n11765), .A2(n7909), .ZN(n12038) );
  NAND2_X1 U12213 ( .A1(n12036), .A2(n12037), .ZN(n12183) );
  NAND2_X1 U12214 ( .A1(n12186), .A2(n12187), .ZN(n12037) );
  NAND3_X1 U12215 ( .A1(a_22_), .A2(n12188), .A3(b_11_), .ZN(n12187) );
  OR2_X1 U12216 ( .A1(n12033), .A2(n12031), .ZN(n12188) );
  NAND2_X1 U12217 ( .A1(n12031), .A2(n12033), .ZN(n12186) );
  NAND2_X1 U12218 ( .A1(n12189), .A2(n12190), .ZN(n12033) );
  NAND2_X1 U12219 ( .A1(n12030), .A2(n12191), .ZN(n12190) );
  OR2_X1 U12220 ( .A1(n12029), .A2(n12027), .ZN(n12191) );
  NOR2_X1 U12221 ( .A1(n11765), .A2(n7916), .ZN(n12030) );
  NAND2_X1 U12222 ( .A1(n12027), .A2(n12029), .ZN(n12189) );
  NAND2_X1 U12223 ( .A1(n12192), .A2(n12193), .ZN(n12029) );
  NAND3_X1 U12224 ( .A1(a_24_), .A2(n12194), .A3(b_11_), .ZN(n12193) );
  NAND2_X1 U12225 ( .A1(n12025), .A2(n12024), .ZN(n12194) );
  OR2_X1 U12226 ( .A1(n12024), .A2(n12025), .ZN(n12192) );
  AND2_X1 U12227 ( .A1(n12195), .A2(n12196), .ZN(n12025) );
  NAND2_X1 U12228 ( .A1(n12022), .A2(n12197), .ZN(n12196) );
  OR2_X1 U12229 ( .A1(n12021), .A2(n12020), .ZN(n12197) );
  NOR2_X1 U12230 ( .A1(n11765), .A2(n7923), .ZN(n12022) );
  NAND2_X1 U12231 ( .A1(n12020), .A2(n12021), .ZN(n12195) );
  NAND2_X1 U12232 ( .A1(n12017), .A2(n12198), .ZN(n12021) );
  NAND2_X1 U12233 ( .A1(n12016), .A2(n12018), .ZN(n12198) );
  NAND2_X1 U12234 ( .A1(n12199), .A2(n12200), .ZN(n12018) );
  NAND2_X1 U12235 ( .A1(b_11_), .A2(a_26_), .ZN(n12200) );
  INV_X1 U12236 ( .A(n12201), .ZN(n12199) );
  XNOR2_X1 U12237 ( .A(n12202), .B(n12203), .ZN(n12016) );
  NAND2_X1 U12238 ( .A1(n12204), .A2(n12205), .ZN(n12202) );
  NAND2_X1 U12239 ( .A1(a_26_), .A2(n12201), .ZN(n12017) );
  NAND2_X1 U12240 ( .A1(n11988), .A2(n12206), .ZN(n12201) );
  NAND2_X1 U12241 ( .A1(n11987), .A2(n11989), .ZN(n12206) );
  NAND2_X1 U12242 ( .A1(n12207), .A2(n12208), .ZN(n11989) );
  NAND2_X1 U12243 ( .A1(b_11_), .A2(a_27_), .ZN(n12208) );
  INV_X1 U12244 ( .A(n12209), .ZN(n12207) );
  XNOR2_X1 U12245 ( .A(n12210), .B(n12211), .ZN(n11987) );
  XOR2_X1 U12246 ( .A(n12212), .B(n12213), .Z(n12210) );
  NAND2_X1 U12247 ( .A1(b_10_), .A2(a_28_), .ZN(n12212) );
  NAND2_X1 U12248 ( .A1(a_27_), .A2(n12209), .ZN(n11988) );
  NAND2_X1 U12249 ( .A1(n12214), .A2(n12215), .ZN(n12209) );
  NAND3_X1 U12250 ( .A1(a_28_), .A2(n12216), .A3(b_11_), .ZN(n12215) );
  NAND2_X1 U12251 ( .A1(n11997), .A2(n11995), .ZN(n12216) );
  OR2_X1 U12252 ( .A1(n11995), .A2(n11997), .ZN(n12214) );
  AND2_X1 U12253 ( .A1(n12217), .A2(n12218), .ZN(n11997) );
  NAND2_X1 U12254 ( .A1(n12012), .A2(n12219), .ZN(n12218) );
  OR2_X1 U12255 ( .A1(n12013), .A2(n12014), .ZN(n12219) );
  NOR2_X1 U12256 ( .A1(n11765), .A2(n7946), .ZN(n12012) );
  NAND2_X1 U12257 ( .A1(n12014), .A2(n12013), .ZN(n12217) );
  NAND2_X1 U12258 ( .A1(n12220), .A2(n12221), .ZN(n12013) );
  NAND2_X1 U12259 ( .A1(b_10_), .A2(n12222), .ZN(n12221) );
  NAND2_X1 U12260 ( .A1(n7272), .A2(n12223), .ZN(n12222) );
  NAND2_X1 U12261 ( .A1(a_30_), .A2(n12224), .ZN(n12223) );
  NAND2_X1 U12262 ( .A1(b_9_), .A2(n12225), .ZN(n12220) );
  NAND2_X1 U12263 ( .A1(n7268), .A2(n12226), .ZN(n12225) );
  NAND2_X1 U12264 ( .A1(a_31_), .A2(n12010), .ZN(n12226) );
  AND3_X1 U12265 ( .A1(b_10_), .A2(n7954), .A3(b_11_), .ZN(n12014) );
  XNOR2_X1 U12266 ( .A(n12227), .B(n12228), .ZN(n11995) );
  XOR2_X1 U12267 ( .A(n12229), .B(n12230), .Z(n12227) );
  XNOR2_X1 U12268 ( .A(n12231), .B(n12232), .ZN(n12020) );
  NAND2_X1 U12269 ( .A1(n12233), .A2(n12234), .ZN(n12231) );
  XNOR2_X1 U12270 ( .A(n12235), .B(n12236), .ZN(n12024) );
  XOR2_X1 U12271 ( .A(n12237), .B(n12238), .Z(n12235) );
  XNOR2_X1 U12272 ( .A(n12239), .B(n12240), .ZN(n12027) );
  XNOR2_X1 U12273 ( .A(n12241), .B(n12242), .ZN(n12239) );
  NOR2_X1 U12274 ( .A1(n7691), .A2(n12010), .ZN(n12242) );
  XNOR2_X1 U12275 ( .A(n12243), .B(n12244), .ZN(n12031) );
  XNOR2_X1 U12276 ( .A(n12245), .B(n12246), .ZN(n12244) );
  XNOR2_X1 U12277 ( .A(n12247), .B(n12248), .ZN(n12036) );
  XOR2_X1 U12278 ( .A(n12249), .B(n12250), .Z(n12248) );
  NAND2_X1 U12279 ( .A1(b_10_), .A2(a_22_), .ZN(n12250) );
  XNOR2_X1 U12280 ( .A(n12251), .B(n12252), .ZN(n11961) );
  XNOR2_X1 U12281 ( .A(n12253), .B(n12254), .ZN(n12251) );
  NOR2_X1 U12282 ( .A1(n7909), .A2(n12010), .ZN(n12254) );
  XNOR2_X1 U12283 ( .A(n12255), .B(n12256), .ZN(n12047) );
  XNOR2_X1 U12284 ( .A(n12257), .B(n12258), .ZN(n12256) );
  XNOR2_X1 U12285 ( .A(n12259), .B(n12260), .ZN(n11944) );
  XOR2_X1 U12286 ( .A(n12261), .B(n12262), .Z(n12259) );
  NOR2_X1 U12287 ( .A1(n7337), .A2(n12010), .ZN(n12262) );
  XNOR2_X1 U12288 ( .A(n12263), .B(n12264), .ZN(n11935) );
  NAND2_X1 U12289 ( .A1(n12265), .A2(n12266), .ZN(n12263) );
  XNOR2_X1 U12290 ( .A(n12267), .B(n12268), .ZN(n12052) );
  NAND2_X1 U12291 ( .A1(n12269), .A2(n12270), .ZN(n12267) );
  XNOR2_X1 U12292 ( .A(n12271), .B(n12272), .ZN(n12055) );
  XNOR2_X1 U12293 ( .A(n12273), .B(n12274), .ZN(n12272) );
  XNOR2_X1 U12294 ( .A(n12275), .B(n12276), .ZN(n11922) );
  XOR2_X1 U12295 ( .A(n12277), .B(n12278), .Z(n12276) );
  NAND2_X1 U12296 ( .A1(b_10_), .A2(a_13_), .ZN(n12278) );
  XOR2_X1 U12297 ( .A(n12279), .B(n12280), .Z(n12060) );
  NAND2_X1 U12298 ( .A1(n12281), .A2(n12282), .ZN(n12279) );
  XOR2_X1 U12299 ( .A(n12283), .B(n12284), .Z(n12064) );
  XNOR2_X1 U12300 ( .A(n12285), .B(n12286), .ZN(n12284) );
  XNOR2_X1 U12301 ( .A(n12287), .B(n12288), .ZN(n11899) );
  NAND2_X1 U12302 ( .A1(n12289), .A2(n12290), .ZN(n12287) );
  XOR2_X1 U12303 ( .A(n12291), .B(n12292), .Z(n12068) );
  NAND2_X1 U12304 ( .A1(n12293), .A2(n12294), .ZN(n12291) );
  XNOR2_X1 U12305 ( .A(n12295), .B(n12296), .ZN(n12071) );
  XNOR2_X1 U12306 ( .A(n12297), .B(n12298), .ZN(n12295) );
  XNOR2_X1 U12307 ( .A(n12299), .B(n12300), .ZN(n12076) );
  XNOR2_X1 U12308 ( .A(n12301), .B(n12302), .ZN(n12300) );
  XNOR2_X1 U12309 ( .A(n12303), .B(n12304), .ZN(n12080) );
  XOR2_X1 U12310 ( .A(n12305), .B(n12306), .Z(n12303) );
  XNOR2_X1 U12311 ( .A(n12307), .B(n12308), .ZN(n12083) );
  XNOR2_X1 U12312 ( .A(n12309), .B(n12310), .ZN(n12308) );
  XNOR2_X1 U12313 ( .A(n12311), .B(n12312), .ZN(n12087) );
  XNOR2_X1 U12314 ( .A(n12313), .B(n12314), .ZN(n12311) );
  XNOR2_X1 U12315 ( .A(n12315), .B(n12316), .ZN(n12091) );
  XNOR2_X1 U12316 ( .A(n12317), .B(n12318), .ZN(n12316) );
  XNOR2_X1 U12317 ( .A(n12319), .B(n12320), .ZN(n12101) );
  XOR2_X1 U12318 ( .A(n12321), .B(n12322), .Z(n12320) );
  NAND2_X1 U12319 ( .A1(b_10_), .A2(a_1_), .ZN(n12322) );
  XOR2_X1 U12320 ( .A(n12099), .B(n12323), .Z(n12106) );
  INV_X1 U12321 ( .A(n12098), .ZN(n12323) );
  XNOR2_X1 U12322 ( .A(n12324), .B(n12325), .ZN(n12099) );
  NOR2_X1 U12323 ( .A1(n7613), .A2(n12010), .ZN(n12325) );
  NAND2_X1 U12324 ( .A1(n12326), .A2(n12327), .ZN(n7251) );
  NAND2_X1 U12325 ( .A1(n12328), .A2(n12329), .ZN(n12327) );
  NAND2_X1 U12326 ( .A1(n12105), .A2(n12104), .ZN(n12326) );
  NAND4_X1 U12327 ( .A1(n12105), .A2(n12328), .A3(n12329), .A4(n12104), .ZN(
        n7252) );
  NAND2_X1 U12328 ( .A1(n12330), .A2(n12331), .ZN(n12104) );
  NAND3_X1 U12329 ( .A1(a_0_), .A2(n12332), .A3(b_10_), .ZN(n12331) );
  OR2_X1 U12330 ( .A1(n12324), .A2(n12098), .ZN(n12332) );
  NAND2_X1 U12331 ( .A1(n12098), .A2(n12324), .ZN(n12330) );
  NAND2_X1 U12332 ( .A1(n12333), .A2(n12334), .ZN(n12324) );
  NAND3_X1 U12333 ( .A1(a_1_), .A2(n12335), .A3(b_10_), .ZN(n12334) );
  OR2_X1 U12334 ( .A1(n12321), .A2(n12319), .ZN(n12335) );
  NAND2_X1 U12335 ( .A1(n12319), .A2(n12321), .ZN(n12333) );
  NAND2_X1 U12336 ( .A1(n12336), .A2(n12337), .ZN(n12321) );
  NAND2_X1 U12337 ( .A1(n12318), .A2(n12338), .ZN(n12337) );
  OR2_X1 U12338 ( .A1(n12317), .A2(n12315), .ZN(n12338) );
  NOR2_X1 U12339 ( .A1(n12010), .A2(n7832), .ZN(n12318) );
  NAND2_X1 U12340 ( .A1(n12315), .A2(n12317), .ZN(n12336) );
  NAND2_X1 U12341 ( .A1(n12339), .A2(n12340), .ZN(n12317) );
  NAND2_X1 U12342 ( .A1(n12314), .A2(n12341), .ZN(n12340) );
  NAND2_X1 U12343 ( .A1(n12313), .A2(n12312), .ZN(n12341) );
  NOR2_X1 U12344 ( .A1(n12010), .A2(n7850), .ZN(n12314) );
  OR2_X1 U12345 ( .A1(n12312), .A2(n12313), .ZN(n12339) );
  AND2_X1 U12346 ( .A1(n12342), .A2(n12343), .ZN(n12313) );
  NAND2_X1 U12347 ( .A1(n12310), .A2(n12344), .ZN(n12343) );
  OR2_X1 U12348 ( .A1(n12309), .A2(n12307), .ZN(n12344) );
  NOR2_X1 U12349 ( .A1(n12010), .A2(n7398), .ZN(n12310) );
  NAND2_X1 U12350 ( .A1(n12307), .A2(n12309), .ZN(n12342) );
  NAND2_X1 U12351 ( .A1(n12345), .A2(n12346), .ZN(n12309) );
  NAND2_X1 U12352 ( .A1(n12306), .A2(n12347), .ZN(n12346) );
  OR2_X1 U12353 ( .A1(n12305), .A2(n12304), .ZN(n12347) );
  NOR2_X1 U12354 ( .A1(n12010), .A2(n7393), .ZN(n12306) );
  NAND2_X1 U12355 ( .A1(n12304), .A2(n12305), .ZN(n12345) );
  NAND2_X1 U12356 ( .A1(n12348), .A2(n12349), .ZN(n12305) );
  NAND2_X1 U12357 ( .A1(n12302), .A2(n12350), .ZN(n12349) );
  OR2_X1 U12358 ( .A1(n12301), .A2(n12299), .ZN(n12350) );
  NOR2_X1 U12359 ( .A1(n12010), .A2(n7388), .ZN(n12302) );
  NAND2_X1 U12360 ( .A1(n12299), .A2(n12301), .ZN(n12348) );
  NAND2_X1 U12361 ( .A1(n12351), .A2(n12352), .ZN(n12301) );
  NAND2_X1 U12362 ( .A1(n12298), .A2(n12353), .ZN(n12352) );
  NAND2_X1 U12363 ( .A1(n12297), .A2(n12296), .ZN(n12353) );
  NOR2_X1 U12364 ( .A1(n12010), .A2(n7863), .ZN(n12298) );
  OR2_X1 U12365 ( .A1(n12296), .A2(n12297), .ZN(n12351) );
  AND2_X1 U12366 ( .A1(n12293), .A2(n12354), .ZN(n12297) );
  NAND2_X1 U12367 ( .A1(n12292), .A2(n12294), .ZN(n12354) );
  NAND2_X1 U12368 ( .A1(n12355), .A2(n12356), .ZN(n12294) );
  NAND2_X1 U12369 ( .A1(b_10_), .A2(a_8_), .ZN(n12356) );
  INV_X1 U12370 ( .A(n12357), .ZN(n12355) );
  XOR2_X1 U12371 ( .A(n12358), .B(n12359), .Z(n12292) );
  XOR2_X1 U12372 ( .A(n12360), .B(n12361), .Z(n12358) );
  NAND2_X1 U12373 ( .A1(a_8_), .A2(n12357), .ZN(n12293) );
  NAND2_X1 U12374 ( .A1(n12289), .A2(n12362), .ZN(n12357) );
  NAND2_X1 U12375 ( .A1(n12288), .A2(n12290), .ZN(n12362) );
  NAND2_X1 U12376 ( .A1(n12363), .A2(n12364), .ZN(n12290) );
  NAND2_X1 U12377 ( .A1(b_10_), .A2(a_9_), .ZN(n12364) );
  INV_X1 U12378 ( .A(n12365), .ZN(n12363) );
  XNOR2_X1 U12379 ( .A(n12366), .B(n12367), .ZN(n12288) );
  XOR2_X1 U12380 ( .A(n12368), .B(n12369), .Z(n12367) );
  NAND2_X1 U12381 ( .A1(a_10_), .A2(b_9_), .ZN(n12369) );
  NAND2_X1 U12382 ( .A1(a_9_), .A2(n12365), .ZN(n12289) );
  NAND2_X1 U12383 ( .A1(n12370), .A2(n12371), .ZN(n12365) );
  NAND2_X1 U12384 ( .A1(n12285), .A2(n12372), .ZN(n12371) );
  OR2_X1 U12385 ( .A1(n12286), .A2(n12283), .ZN(n12372) );
  NAND2_X1 U12386 ( .A1(n12283), .A2(n12286), .ZN(n12370) );
  NAND2_X1 U12387 ( .A1(n12281), .A2(n12373), .ZN(n12286) );
  NAND2_X1 U12388 ( .A1(n12280), .A2(n12282), .ZN(n12373) );
  NAND2_X1 U12389 ( .A1(n12374), .A2(n12375), .ZN(n12282) );
  NAND2_X1 U12390 ( .A1(b_10_), .A2(a_11_), .ZN(n12375) );
  INV_X1 U12391 ( .A(n12376), .ZN(n12374) );
  XNOR2_X1 U12392 ( .A(n12377), .B(n12378), .ZN(n12280) );
  XOR2_X1 U12393 ( .A(n12379), .B(n12380), .Z(n12378) );
  NAND2_X1 U12394 ( .A1(a_12_), .A2(b_9_), .ZN(n12380) );
  NAND2_X1 U12395 ( .A1(a_11_), .A2(n12376), .ZN(n12281) );
  NAND2_X1 U12396 ( .A1(n12144), .A2(n12381), .ZN(n12376) );
  NAND2_X1 U12397 ( .A1(n12143), .A2(n12145), .ZN(n12381) );
  NAND2_X1 U12398 ( .A1(n12382), .A2(n12383), .ZN(n12145) );
  NAND2_X1 U12399 ( .A1(b_10_), .A2(a_12_), .ZN(n12383) );
  INV_X1 U12400 ( .A(n12384), .ZN(n12382) );
  XNOR2_X1 U12401 ( .A(n12385), .B(n12386), .ZN(n12143) );
  XOR2_X1 U12402 ( .A(n12387), .B(n12388), .Z(n12386) );
  NAND2_X1 U12403 ( .A1(a_13_), .A2(b_9_), .ZN(n12388) );
  NAND2_X1 U12404 ( .A1(a_12_), .A2(n12384), .ZN(n12144) );
  NAND2_X1 U12405 ( .A1(n12389), .A2(n12390), .ZN(n12384) );
  NAND3_X1 U12406 ( .A1(a_13_), .A2(n12391), .A3(b_10_), .ZN(n12390) );
  OR2_X1 U12407 ( .A1(n12277), .A2(n12275), .ZN(n12391) );
  NAND2_X1 U12408 ( .A1(n12275), .A2(n12277), .ZN(n12389) );
  NAND2_X1 U12409 ( .A1(n12392), .A2(n12393), .ZN(n12277) );
  NAND2_X1 U12410 ( .A1(n12274), .A2(n12394), .ZN(n12393) );
  OR2_X1 U12411 ( .A1(n12273), .A2(n12271), .ZN(n12394) );
  NOR2_X1 U12412 ( .A1(n12010), .A2(n7782), .ZN(n12274) );
  NAND2_X1 U12413 ( .A1(n12271), .A2(n12273), .ZN(n12392) );
  NAND2_X1 U12414 ( .A1(n12269), .A2(n12395), .ZN(n12273) );
  NAND2_X1 U12415 ( .A1(n12268), .A2(n12270), .ZN(n12395) );
  NAND2_X1 U12416 ( .A1(n12396), .A2(n12397), .ZN(n12270) );
  NAND2_X1 U12417 ( .A1(b_10_), .A2(a_15_), .ZN(n12397) );
  INV_X1 U12418 ( .A(n12398), .ZN(n12396) );
  XNOR2_X1 U12419 ( .A(n12399), .B(n12400), .ZN(n12268) );
  XOR2_X1 U12420 ( .A(n12401), .B(n12402), .Z(n12400) );
  NAND2_X1 U12421 ( .A1(a_16_), .A2(b_9_), .ZN(n12402) );
  NAND2_X1 U12422 ( .A1(a_15_), .A2(n12398), .ZN(n12269) );
  NAND2_X1 U12423 ( .A1(n12265), .A2(n12403), .ZN(n12398) );
  NAND2_X1 U12424 ( .A1(n12264), .A2(n12266), .ZN(n12403) );
  NAND2_X1 U12425 ( .A1(n12404), .A2(n12405), .ZN(n12266) );
  NAND2_X1 U12426 ( .A1(b_10_), .A2(a_16_), .ZN(n12405) );
  INV_X1 U12427 ( .A(n12406), .ZN(n12404) );
  XNOR2_X1 U12428 ( .A(n12407), .B(n12408), .ZN(n12264) );
  XNOR2_X1 U12429 ( .A(n12409), .B(n12410), .ZN(n12407) );
  NOR2_X1 U12430 ( .A1(n12224), .A2(n7337), .ZN(n12410) );
  NAND2_X1 U12431 ( .A1(a_16_), .A2(n12406), .ZN(n12265) );
  NAND2_X1 U12432 ( .A1(n12411), .A2(n12412), .ZN(n12406) );
  NAND3_X1 U12433 ( .A1(a_17_), .A2(n12413), .A3(b_10_), .ZN(n12412) );
  OR2_X1 U12434 ( .A1(n12261), .A2(n12260), .ZN(n12413) );
  NAND2_X1 U12435 ( .A1(n12260), .A2(n12261), .ZN(n12411) );
  NAND2_X1 U12436 ( .A1(n12414), .A2(n12415), .ZN(n12261) );
  NAND2_X1 U12437 ( .A1(n12258), .A2(n12416), .ZN(n12415) );
  OR2_X1 U12438 ( .A1(n12257), .A2(n12255), .ZN(n12416) );
  NOR2_X1 U12439 ( .A1(n12010), .A2(n7764), .ZN(n12258) );
  NAND2_X1 U12440 ( .A1(n12255), .A2(n12257), .ZN(n12414) );
  NAND2_X1 U12441 ( .A1(n12417), .A2(n12418), .ZN(n12257) );
  NAND2_X1 U12442 ( .A1(n12171), .A2(n12419), .ZN(n12418) );
  OR2_X1 U12443 ( .A1(n12170), .A2(n12168), .ZN(n12419) );
  NOR2_X1 U12444 ( .A1(n12010), .A2(n7902), .ZN(n12171) );
  NAND2_X1 U12445 ( .A1(n12168), .A2(n12170), .ZN(n12417) );
  NAND2_X1 U12446 ( .A1(n12420), .A2(n12421), .ZN(n12170) );
  NAND2_X1 U12447 ( .A1(n12179), .A2(n12422), .ZN(n12421) );
  OR2_X1 U12448 ( .A1(n12178), .A2(n12176), .ZN(n12422) );
  NOR2_X1 U12449 ( .A1(n12010), .A2(n7987), .ZN(n12179) );
  NAND2_X1 U12450 ( .A1(n12176), .A2(n12178), .ZN(n12420) );
  NAND2_X1 U12451 ( .A1(n12423), .A2(n12424), .ZN(n12178) );
  NAND3_X1 U12452 ( .A1(a_21_), .A2(n12425), .A3(b_10_), .ZN(n12424) );
  NAND2_X1 U12453 ( .A1(n12253), .A2(n12252), .ZN(n12425) );
  OR2_X1 U12454 ( .A1(n12252), .A2(n12253), .ZN(n12423) );
  AND2_X1 U12455 ( .A1(n12426), .A2(n12427), .ZN(n12253) );
  NAND3_X1 U12456 ( .A1(a_22_), .A2(n12428), .A3(b_10_), .ZN(n12427) );
  OR2_X1 U12457 ( .A1(n12249), .A2(n12247), .ZN(n12428) );
  NAND2_X1 U12458 ( .A1(n12247), .A2(n12249), .ZN(n12426) );
  NAND2_X1 U12459 ( .A1(n12429), .A2(n12430), .ZN(n12249) );
  NAND2_X1 U12460 ( .A1(n12246), .A2(n12431), .ZN(n12430) );
  OR2_X1 U12461 ( .A1(n12245), .A2(n12243), .ZN(n12431) );
  NOR2_X1 U12462 ( .A1(n12010), .A2(n7916), .ZN(n12246) );
  NAND2_X1 U12463 ( .A1(n12243), .A2(n12245), .ZN(n12429) );
  NAND2_X1 U12464 ( .A1(n12432), .A2(n12433), .ZN(n12245) );
  NAND3_X1 U12465 ( .A1(a_24_), .A2(n12434), .A3(b_10_), .ZN(n12433) );
  NAND2_X1 U12466 ( .A1(n12241), .A2(n12240), .ZN(n12434) );
  OR2_X1 U12467 ( .A1(n12240), .A2(n12241), .ZN(n12432) );
  AND2_X1 U12468 ( .A1(n12435), .A2(n12436), .ZN(n12241) );
  NAND2_X1 U12469 ( .A1(n12238), .A2(n12437), .ZN(n12436) );
  OR2_X1 U12470 ( .A1(n12237), .A2(n12236), .ZN(n12437) );
  NOR2_X1 U12471 ( .A1(n12010), .A2(n7923), .ZN(n12238) );
  NAND2_X1 U12472 ( .A1(n12236), .A2(n12237), .ZN(n12435) );
  NAND2_X1 U12473 ( .A1(n12233), .A2(n12438), .ZN(n12237) );
  NAND2_X1 U12474 ( .A1(n12232), .A2(n12234), .ZN(n12438) );
  NAND2_X1 U12475 ( .A1(n12439), .A2(n12440), .ZN(n12234) );
  NAND2_X1 U12476 ( .A1(b_10_), .A2(a_26_), .ZN(n12440) );
  INV_X1 U12477 ( .A(n12441), .ZN(n12439) );
  XNOR2_X1 U12478 ( .A(n12442), .B(n12443), .ZN(n12232) );
  NAND2_X1 U12479 ( .A1(n12444), .A2(n12445), .ZN(n12442) );
  NAND2_X1 U12480 ( .A1(a_26_), .A2(n12441), .ZN(n12233) );
  NAND2_X1 U12481 ( .A1(n12204), .A2(n12446), .ZN(n12441) );
  NAND2_X1 U12482 ( .A1(n12203), .A2(n12205), .ZN(n12446) );
  NAND2_X1 U12483 ( .A1(n12447), .A2(n12448), .ZN(n12205) );
  NAND2_X1 U12484 ( .A1(b_10_), .A2(a_27_), .ZN(n12448) );
  INV_X1 U12485 ( .A(n12449), .ZN(n12447) );
  XNOR2_X1 U12486 ( .A(n12450), .B(n12451), .ZN(n12203) );
  XOR2_X1 U12487 ( .A(n12452), .B(n12453), .Z(n12450) );
  NAND2_X1 U12488 ( .A1(a_28_), .A2(b_9_), .ZN(n12452) );
  NAND2_X1 U12489 ( .A1(a_27_), .A2(n12449), .ZN(n12204) );
  NAND2_X1 U12490 ( .A1(n12454), .A2(n12455), .ZN(n12449) );
  NAND3_X1 U12491 ( .A1(a_28_), .A2(n12456), .A3(b_10_), .ZN(n12455) );
  NAND2_X1 U12492 ( .A1(n12213), .A2(n12211), .ZN(n12456) );
  OR2_X1 U12493 ( .A1(n12211), .A2(n12213), .ZN(n12454) );
  AND2_X1 U12494 ( .A1(n12457), .A2(n12458), .ZN(n12213) );
  NAND2_X1 U12495 ( .A1(n12228), .A2(n12459), .ZN(n12458) );
  OR2_X1 U12496 ( .A1(n12229), .A2(n12230), .ZN(n12459) );
  NOR2_X1 U12497 ( .A1(n12010), .A2(n7946), .ZN(n12228) );
  NAND2_X1 U12498 ( .A1(n12230), .A2(n12229), .ZN(n12457) );
  NAND2_X1 U12499 ( .A1(n12460), .A2(n12461), .ZN(n12229) );
  NAND2_X1 U12500 ( .A1(b_8_), .A2(n12462), .ZN(n12461) );
  NAND2_X1 U12501 ( .A1(n7268), .A2(n12463), .ZN(n12462) );
  NAND2_X1 U12502 ( .A1(a_31_), .A2(n12224), .ZN(n12463) );
  NAND2_X1 U12503 ( .A1(b_9_), .A2(n12464), .ZN(n12460) );
  NAND2_X1 U12504 ( .A1(n7272), .A2(n12465), .ZN(n12464) );
  NAND2_X1 U12505 ( .A1(a_30_), .A2(n12466), .ZN(n12465) );
  AND3_X1 U12506 ( .A1(n7954), .A2(b_9_), .A3(b_10_), .ZN(n12230) );
  XNOR2_X1 U12507 ( .A(n12467), .B(n12468), .ZN(n12211) );
  XOR2_X1 U12508 ( .A(n12469), .B(n12470), .Z(n12467) );
  XNOR2_X1 U12509 ( .A(n12471), .B(n12472), .ZN(n12236) );
  NAND2_X1 U12510 ( .A1(n12473), .A2(n12474), .ZN(n12471) );
  XNOR2_X1 U12511 ( .A(n12475), .B(n12476), .ZN(n12240) );
  XOR2_X1 U12512 ( .A(n12477), .B(n12478), .Z(n12475) );
  XNOR2_X1 U12513 ( .A(n12479), .B(n12480), .ZN(n12243) );
  XNOR2_X1 U12514 ( .A(n12481), .B(n12482), .ZN(n12479) );
  NOR2_X1 U12515 ( .A1(n12224), .A2(n7691), .ZN(n12482) );
  XNOR2_X1 U12516 ( .A(n12483), .B(n12484), .ZN(n12247) );
  XNOR2_X1 U12517 ( .A(n12485), .B(n12486), .ZN(n12484) );
  XOR2_X1 U12518 ( .A(n12487), .B(n12488), .Z(n12252) );
  XNOR2_X1 U12519 ( .A(n12489), .B(n12490), .ZN(n12488) );
  XOR2_X1 U12520 ( .A(n12491), .B(n12492), .Z(n12176) );
  XOR2_X1 U12521 ( .A(n12493), .B(n12494), .Z(n12491) );
  NOR2_X1 U12522 ( .A1(n12224), .A2(n7909), .ZN(n12494) );
  XOR2_X1 U12523 ( .A(n12495), .B(n12496), .Z(n12168) );
  XOR2_X1 U12524 ( .A(n12497), .B(n12498), .Z(n12495) );
  NOR2_X1 U12525 ( .A1(n12224), .A2(n7987), .ZN(n12498) );
  XNOR2_X1 U12526 ( .A(n12499), .B(n12500), .ZN(n12255) );
  XOR2_X1 U12527 ( .A(n12501), .B(n12502), .Z(n12500) );
  NAND2_X1 U12528 ( .A1(a_19_), .A2(b_9_), .ZN(n12502) );
  XNOR2_X1 U12529 ( .A(n12503), .B(n12504), .ZN(n12260) );
  XNOR2_X1 U12530 ( .A(n12505), .B(n12506), .ZN(n12503) );
  NOR2_X1 U12531 ( .A1(n12224), .A2(n7764), .ZN(n12506) );
  XOR2_X1 U12532 ( .A(n12507), .B(n12508), .Z(n12271) );
  XOR2_X1 U12533 ( .A(n12509), .B(n12510), .Z(n12507) );
  NOR2_X1 U12534 ( .A1(n12224), .A2(n7346), .ZN(n12510) );
  XNOR2_X1 U12535 ( .A(n12511), .B(n12512), .ZN(n12275) );
  XOR2_X1 U12536 ( .A(n12513), .B(n12514), .Z(n12512) );
  NAND2_X1 U12537 ( .A1(a_14_), .A2(b_9_), .ZN(n12514) );
  XNOR2_X1 U12538 ( .A(n12515), .B(n12516), .ZN(n12283) );
  XOR2_X1 U12539 ( .A(n12517), .B(n12518), .Z(n12516) );
  NAND2_X1 U12540 ( .A1(a_11_), .A2(b_9_), .ZN(n12518) );
  XNOR2_X1 U12541 ( .A(n12519), .B(n12520), .ZN(n12296) );
  XOR2_X1 U12542 ( .A(n12521), .B(n12522), .Z(n12519) );
  NOR2_X1 U12543 ( .A1(n12224), .A2(n8037), .ZN(n12522) );
  XNOR2_X1 U12544 ( .A(n12523), .B(n12524), .ZN(n12299) );
  XOR2_X1 U12545 ( .A(n12525), .B(n12526), .Z(n12524) );
  NAND2_X1 U12546 ( .A1(a_7_), .A2(b_9_), .ZN(n12526) );
  XNOR2_X1 U12547 ( .A(n12527), .B(n12528), .ZN(n12304) );
  XNOR2_X1 U12548 ( .A(n12529), .B(n12530), .ZN(n12527) );
  NOR2_X1 U12549 ( .A1(n12224), .A2(n7388), .ZN(n12530) );
  XOR2_X1 U12550 ( .A(n12531), .B(n12532), .Z(n12307) );
  XOR2_X1 U12551 ( .A(n12533), .B(n12534), .Z(n12531) );
  NOR2_X1 U12552 ( .A1(n12224), .A2(n7393), .ZN(n12534) );
  XNOR2_X1 U12553 ( .A(n12535), .B(n12536), .ZN(n12312) );
  XOR2_X1 U12554 ( .A(n12537), .B(n12538), .Z(n12535) );
  NOR2_X1 U12555 ( .A1(n12224), .A2(n7398), .ZN(n12538) );
  XOR2_X1 U12556 ( .A(n12539), .B(n12540), .Z(n12315) );
  XOR2_X1 U12557 ( .A(n12541), .B(n12542), .Z(n12539) );
  NOR2_X1 U12558 ( .A1(n12224), .A2(n7850), .ZN(n12542) );
  XOR2_X1 U12559 ( .A(n12543), .B(n12544), .Z(n12319) );
  XOR2_X1 U12560 ( .A(n12545), .B(n12546), .Z(n12543) );
  NOR2_X1 U12561 ( .A1(n12224), .A2(n7832), .ZN(n12546) );
  XOR2_X1 U12562 ( .A(n12547), .B(n12548), .Z(n12098) );
  XOR2_X1 U12563 ( .A(n12549), .B(n12550), .Z(n12547) );
  NOR2_X1 U12564 ( .A1(n12224), .A2(n7411), .ZN(n12550) );
  NAND3_X1 U12565 ( .A1(n12551), .A2(n12552), .A3(n12553), .ZN(n12328) );
  XOR2_X1 U12566 ( .A(n12554), .B(n12555), .Z(n12553) );
  XOR2_X1 U12567 ( .A(n12556), .B(n12557), .Z(n12105) );
  XOR2_X1 U12568 ( .A(n12558), .B(n12559), .Z(n12556) );
  NAND2_X1 U12569 ( .A1(n12560), .A2(n12329), .ZN(n7255) );
  OR2_X1 U12570 ( .A1(n12329), .A2(n12560), .ZN(n7256) );
  XNOR2_X1 U12571 ( .A(n12561), .B(n12562), .ZN(n12560) );
  NAND2_X1 U12572 ( .A1(n12563), .A2(n12564), .ZN(n12329) );
  NAND2_X1 U12573 ( .A1(n12551), .A2(n12552), .ZN(n12564) );
  NAND2_X1 U12574 ( .A1(n12559), .A2(n12565), .ZN(n12552) );
  OR2_X1 U12575 ( .A1(n12558), .A2(n12557), .ZN(n12565) );
  NOR2_X1 U12576 ( .A1(n12224), .A2(n7613), .ZN(n12559) );
  NAND2_X1 U12577 ( .A1(n12557), .A2(n12558), .ZN(n12551) );
  NAND2_X1 U12578 ( .A1(n12566), .A2(n12567), .ZN(n12558) );
  NAND3_X1 U12579 ( .A1(b_9_), .A2(n12568), .A3(a_1_), .ZN(n12567) );
  OR2_X1 U12580 ( .A1(n12549), .A2(n12548), .ZN(n12568) );
  NAND2_X1 U12581 ( .A1(n12548), .A2(n12549), .ZN(n12566) );
  NAND2_X1 U12582 ( .A1(n12569), .A2(n12570), .ZN(n12549) );
  NAND3_X1 U12583 ( .A1(b_9_), .A2(n12571), .A3(a_2_), .ZN(n12570) );
  OR2_X1 U12584 ( .A1(n12545), .A2(n12544), .ZN(n12571) );
  NAND2_X1 U12585 ( .A1(n12544), .A2(n12545), .ZN(n12569) );
  NAND2_X1 U12586 ( .A1(n12572), .A2(n12573), .ZN(n12545) );
  NAND3_X1 U12587 ( .A1(b_9_), .A2(n12574), .A3(a_3_), .ZN(n12573) );
  OR2_X1 U12588 ( .A1(n12541), .A2(n12540), .ZN(n12574) );
  NAND2_X1 U12589 ( .A1(n12540), .A2(n12541), .ZN(n12572) );
  NAND2_X1 U12590 ( .A1(n12575), .A2(n12576), .ZN(n12541) );
  NAND3_X1 U12591 ( .A1(b_9_), .A2(n12577), .A3(a_4_), .ZN(n12576) );
  OR2_X1 U12592 ( .A1(n12537), .A2(n12536), .ZN(n12577) );
  NAND2_X1 U12593 ( .A1(n12536), .A2(n12537), .ZN(n12575) );
  NAND2_X1 U12594 ( .A1(n12578), .A2(n12579), .ZN(n12537) );
  NAND3_X1 U12595 ( .A1(b_9_), .A2(n12580), .A3(a_5_), .ZN(n12579) );
  OR2_X1 U12596 ( .A1(n12533), .A2(n12532), .ZN(n12580) );
  NAND2_X1 U12597 ( .A1(n12532), .A2(n12533), .ZN(n12578) );
  NAND2_X1 U12598 ( .A1(n12581), .A2(n12582), .ZN(n12533) );
  NAND3_X1 U12599 ( .A1(b_9_), .A2(n12583), .A3(a_6_), .ZN(n12582) );
  NAND2_X1 U12600 ( .A1(n12529), .A2(n12528), .ZN(n12583) );
  OR2_X1 U12601 ( .A1(n12528), .A2(n12529), .ZN(n12581) );
  AND2_X1 U12602 ( .A1(n12584), .A2(n12585), .ZN(n12529) );
  NAND3_X1 U12603 ( .A1(b_9_), .A2(n12586), .A3(a_7_), .ZN(n12585) );
  OR2_X1 U12604 ( .A1(n12525), .A2(n12523), .ZN(n12586) );
  NAND2_X1 U12605 ( .A1(n12523), .A2(n12525), .ZN(n12584) );
  NAND2_X1 U12606 ( .A1(n12587), .A2(n12588), .ZN(n12525) );
  NAND3_X1 U12607 ( .A1(b_9_), .A2(n12589), .A3(a_8_), .ZN(n12588) );
  OR2_X1 U12608 ( .A1(n12521), .A2(n12520), .ZN(n12589) );
  NAND2_X1 U12609 ( .A1(n12520), .A2(n12521), .ZN(n12587) );
  NAND2_X1 U12610 ( .A1(n12590), .A2(n12591), .ZN(n12521) );
  NAND2_X1 U12611 ( .A1(n12359), .A2(n12592), .ZN(n12591) );
  OR2_X1 U12612 ( .A1(n12360), .A2(n12361), .ZN(n12592) );
  XNOR2_X1 U12613 ( .A(n12593), .B(n12594), .ZN(n12359) );
  XNOR2_X1 U12614 ( .A(n12595), .B(n12596), .ZN(n12594) );
  NAND2_X1 U12615 ( .A1(n12361), .A2(n12360), .ZN(n12590) );
  NAND2_X1 U12616 ( .A1(n12597), .A2(n12598), .ZN(n12360) );
  NAND3_X1 U12617 ( .A1(b_9_), .A2(n12599), .A3(a_10_), .ZN(n12598) );
  OR2_X1 U12618 ( .A1(n12368), .A2(n12366), .ZN(n12599) );
  NAND2_X1 U12619 ( .A1(n12366), .A2(n12368), .ZN(n12597) );
  NAND2_X1 U12620 ( .A1(n12600), .A2(n12601), .ZN(n12368) );
  NAND3_X1 U12621 ( .A1(b_9_), .A2(n12602), .A3(a_11_), .ZN(n12601) );
  OR2_X1 U12622 ( .A1(n12517), .A2(n12515), .ZN(n12602) );
  NAND2_X1 U12623 ( .A1(n12515), .A2(n12517), .ZN(n12600) );
  NAND2_X1 U12624 ( .A1(n12603), .A2(n12604), .ZN(n12517) );
  NAND3_X1 U12625 ( .A1(b_9_), .A2(n12605), .A3(a_12_), .ZN(n12604) );
  OR2_X1 U12626 ( .A1(n12379), .A2(n12377), .ZN(n12605) );
  NAND2_X1 U12627 ( .A1(n12377), .A2(n12379), .ZN(n12603) );
  NAND2_X1 U12628 ( .A1(n12606), .A2(n12607), .ZN(n12379) );
  NAND3_X1 U12629 ( .A1(b_9_), .A2(n12608), .A3(a_13_), .ZN(n12607) );
  OR2_X1 U12630 ( .A1(n12387), .A2(n12385), .ZN(n12608) );
  NAND2_X1 U12631 ( .A1(n12385), .A2(n12387), .ZN(n12606) );
  NAND2_X1 U12632 ( .A1(n12609), .A2(n12610), .ZN(n12387) );
  NAND3_X1 U12633 ( .A1(b_9_), .A2(n12611), .A3(a_14_), .ZN(n12610) );
  OR2_X1 U12634 ( .A1(n12513), .A2(n12511), .ZN(n12611) );
  NAND2_X1 U12635 ( .A1(n12511), .A2(n12513), .ZN(n12609) );
  NAND2_X1 U12636 ( .A1(n12612), .A2(n12613), .ZN(n12513) );
  NAND3_X1 U12637 ( .A1(b_9_), .A2(n12614), .A3(a_15_), .ZN(n12613) );
  OR2_X1 U12638 ( .A1(n12509), .A2(n12508), .ZN(n12614) );
  NAND2_X1 U12639 ( .A1(n12508), .A2(n12509), .ZN(n12612) );
  NAND2_X1 U12640 ( .A1(n12615), .A2(n12616), .ZN(n12509) );
  NAND3_X1 U12641 ( .A1(b_9_), .A2(n12617), .A3(a_16_), .ZN(n12616) );
  OR2_X1 U12642 ( .A1(n12401), .A2(n12399), .ZN(n12617) );
  NAND2_X1 U12643 ( .A1(n12399), .A2(n12401), .ZN(n12615) );
  NAND2_X1 U12644 ( .A1(n12618), .A2(n12619), .ZN(n12401) );
  NAND3_X1 U12645 ( .A1(b_9_), .A2(n12620), .A3(a_17_), .ZN(n12619) );
  NAND2_X1 U12646 ( .A1(n12409), .A2(n12408), .ZN(n12620) );
  OR2_X1 U12647 ( .A1(n12408), .A2(n12409), .ZN(n12618) );
  AND2_X1 U12648 ( .A1(n12621), .A2(n12622), .ZN(n12409) );
  NAND3_X1 U12649 ( .A1(b_9_), .A2(n12623), .A3(a_18_), .ZN(n12622) );
  NAND2_X1 U12650 ( .A1(n12505), .A2(n12504), .ZN(n12623) );
  OR2_X1 U12651 ( .A1(n12504), .A2(n12505), .ZN(n12621) );
  AND2_X1 U12652 ( .A1(n12624), .A2(n12625), .ZN(n12505) );
  NAND3_X1 U12653 ( .A1(b_9_), .A2(n12626), .A3(a_19_), .ZN(n12625) );
  OR2_X1 U12654 ( .A1(n12501), .A2(n12499), .ZN(n12626) );
  NAND2_X1 U12655 ( .A1(n12499), .A2(n12501), .ZN(n12624) );
  NAND2_X1 U12656 ( .A1(n12627), .A2(n12628), .ZN(n12501) );
  NAND3_X1 U12657 ( .A1(b_9_), .A2(n12629), .A3(a_20_), .ZN(n12628) );
  OR2_X1 U12658 ( .A1(n12497), .A2(n12496), .ZN(n12629) );
  NAND2_X1 U12659 ( .A1(n12496), .A2(n12497), .ZN(n12627) );
  NAND2_X1 U12660 ( .A1(n12630), .A2(n12631), .ZN(n12497) );
  NAND3_X1 U12661 ( .A1(b_9_), .A2(n12632), .A3(a_21_), .ZN(n12631) );
  OR2_X1 U12662 ( .A1(n12493), .A2(n12492), .ZN(n12632) );
  NAND2_X1 U12663 ( .A1(n12492), .A2(n12493), .ZN(n12630) );
  NAND2_X1 U12664 ( .A1(n12633), .A2(n12634), .ZN(n12493) );
  NAND2_X1 U12665 ( .A1(n12490), .A2(n12635), .ZN(n12634) );
  OR2_X1 U12666 ( .A1(n12489), .A2(n12487), .ZN(n12635) );
  NOR2_X1 U12667 ( .A1(n7312), .A2(n12224), .ZN(n12490) );
  NAND2_X1 U12668 ( .A1(n12487), .A2(n12489), .ZN(n12633) );
  NAND2_X1 U12669 ( .A1(n12636), .A2(n12637), .ZN(n12489) );
  NAND2_X1 U12670 ( .A1(n12486), .A2(n12638), .ZN(n12637) );
  OR2_X1 U12671 ( .A1(n12485), .A2(n12483), .ZN(n12638) );
  NOR2_X1 U12672 ( .A1(n7916), .A2(n12224), .ZN(n12486) );
  NAND2_X1 U12673 ( .A1(n12483), .A2(n12485), .ZN(n12636) );
  NAND2_X1 U12674 ( .A1(n12639), .A2(n12640), .ZN(n12485) );
  NAND3_X1 U12675 ( .A1(b_9_), .A2(n12641), .A3(a_24_), .ZN(n12640) );
  NAND2_X1 U12676 ( .A1(n12481), .A2(n12480), .ZN(n12641) );
  OR2_X1 U12677 ( .A1(n12480), .A2(n12481), .ZN(n12639) );
  AND2_X1 U12678 ( .A1(n12642), .A2(n12643), .ZN(n12481) );
  NAND2_X1 U12679 ( .A1(n12478), .A2(n12644), .ZN(n12643) );
  OR2_X1 U12680 ( .A1(n12477), .A2(n12476), .ZN(n12644) );
  NOR2_X1 U12681 ( .A1(n7923), .A2(n12224), .ZN(n12478) );
  NAND2_X1 U12682 ( .A1(n12476), .A2(n12477), .ZN(n12642) );
  NAND2_X1 U12683 ( .A1(n12473), .A2(n12645), .ZN(n12477) );
  NAND2_X1 U12684 ( .A1(n12472), .A2(n12474), .ZN(n12645) );
  NAND2_X1 U12685 ( .A1(n12646), .A2(n12647), .ZN(n12474) );
  NAND2_X1 U12686 ( .A1(a_26_), .A2(b_9_), .ZN(n12647) );
  INV_X1 U12687 ( .A(n12648), .ZN(n12646) );
  XNOR2_X1 U12688 ( .A(n12649), .B(n12650), .ZN(n12472) );
  NAND2_X1 U12689 ( .A1(n12651), .A2(n12652), .ZN(n12649) );
  NAND2_X1 U12690 ( .A1(a_26_), .A2(n12648), .ZN(n12473) );
  NAND2_X1 U12691 ( .A1(n12444), .A2(n12653), .ZN(n12648) );
  NAND2_X1 U12692 ( .A1(n12443), .A2(n12445), .ZN(n12653) );
  NAND2_X1 U12693 ( .A1(n12654), .A2(n12655), .ZN(n12445) );
  NAND2_X1 U12694 ( .A1(a_27_), .A2(b_9_), .ZN(n12655) );
  INV_X1 U12695 ( .A(n12656), .ZN(n12654) );
  XNOR2_X1 U12696 ( .A(n12657), .B(n12658), .ZN(n12443) );
  XOR2_X1 U12697 ( .A(n12659), .B(n12660), .Z(n12657) );
  NAND2_X1 U12698 ( .A1(a_28_), .A2(b_8_), .ZN(n12659) );
  NAND2_X1 U12699 ( .A1(a_27_), .A2(n12656), .ZN(n12444) );
  NAND2_X1 U12700 ( .A1(n12661), .A2(n12662), .ZN(n12656) );
  NAND3_X1 U12701 ( .A1(b_9_), .A2(n12663), .A3(a_28_), .ZN(n12662) );
  NAND2_X1 U12702 ( .A1(n12453), .A2(n12451), .ZN(n12663) );
  OR2_X1 U12703 ( .A1(n12451), .A2(n12453), .ZN(n12661) );
  AND2_X1 U12704 ( .A1(n12664), .A2(n12665), .ZN(n12453) );
  NAND2_X1 U12705 ( .A1(n12468), .A2(n12666), .ZN(n12665) );
  OR2_X1 U12706 ( .A1(n12469), .A2(n12470), .ZN(n12666) );
  NOR2_X1 U12707 ( .A1(n7946), .A2(n12224), .ZN(n12468) );
  NAND2_X1 U12708 ( .A1(n12470), .A2(n12469), .ZN(n12664) );
  NAND2_X1 U12709 ( .A1(n12667), .A2(n12668), .ZN(n12469) );
  NAND2_X1 U12710 ( .A1(b_7_), .A2(n12669), .ZN(n12668) );
  NAND2_X1 U12711 ( .A1(n7268), .A2(n12670), .ZN(n12669) );
  NAND2_X1 U12712 ( .A1(a_31_), .A2(n12466), .ZN(n12670) );
  NAND2_X1 U12713 ( .A1(b_8_), .A2(n12671), .ZN(n12667) );
  NAND2_X1 U12714 ( .A1(n7272), .A2(n12672), .ZN(n12671) );
  NAND2_X1 U12715 ( .A1(a_30_), .A2(n12673), .ZN(n12672) );
  AND3_X1 U12716 ( .A1(n7954), .A2(b_9_), .A3(b_8_), .ZN(n12470) );
  XNOR2_X1 U12717 ( .A(n12674), .B(n12675), .ZN(n12451) );
  XOR2_X1 U12718 ( .A(n12676), .B(n12677), .Z(n12674) );
  XNOR2_X1 U12719 ( .A(n12678), .B(n12679), .ZN(n12476) );
  NAND2_X1 U12720 ( .A1(n12680), .A2(n12681), .ZN(n12678) );
  XNOR2_X1 U12721 ( .A(n12682), .B(n12683), .ZN(n12480) );
  XOR2_X1 U12722 ( .A(n12684), .B(n12685), .Z(n12682) );
  XNOR2_X1 U12723 ( .A(n12686), .B(n12687), .ZN(n12483) );
  XNOR2_X1 U12724 ( .A(n12688), .B(n12689), .ZN(n12686) );
  NOR2_X1 U12725 ( .A1(n12466), .A2(n7691), .ZN(n12689) );
  XNOR2_X1 U12726 ( .A(n12690), .B(n12691), .ZN(n12487) );
  XOR2_X1 U12727 ( .A(n12692), .B(n12693), .Z(n12691) );
  NAND2_X1 U12728 ( .A1(b_8_), .A2(a_23_), .ZN(n12693) );
  XNOR2_X1 U12729 ( .A(n12694), .B(n12695), .ZN(n12492) );
  XNOR2_X1 U12730 ( .A(n12696), .B(n12697), .ZN(n12695) );
  XNOR2_X1 U12731 ( .A(n12698), .B(n12699), .ZN(n12496) );
  XNOR2_X1 U12732 ( .A(n12700), .B(n12701), .ZN(n12698) );
  XNOR2_X1 U12733 ( .A(n12702), .B(n12703), .ZN(n12499) );
  XNOR2_X1 U12734 ( .A(n12704), .B(n12705), .ZN(n12702) );
  XNOR2_X1 U12735 ( .A(n12706), .B(n12707), .ZN(n12504) );
  XOR2_X1 U12736 ( .A(n12708), .B(n12709), .Z(n12706) );
  XOR2_X1 U12737 ( .A(n12710), .B(n12711), .Z(n12408) );
  XOR2_X1 U12738 ( .A(n12712), .B(n12713), .Z(n12711) );
  NAND2_X1 U12739 ( .A1(a_18_), .A2(b_8_), .ZN(n12713) );
  XNOR2_X1 U12740 ( .A(n12714), .B(n12715), .ZN(n12399) );
  NAND2_X1 U12741 ( .A1(n12716), .A2(n12717), .ZN(n12714) );
  XNOR2_X1 U12742 ( .A(n12718), .B(n12719), .ZN(n12508) );
  NAND2_X1 U12743 ( .A1(n12720), .A2(n12721), .ZN(n12718) );
  XNOR2_X1 U12744 ( .A(n12722), .B(n12723), .ZN(n12511) );
  XNOR2_X1 U12745 ( .A(n12724), .B(n12725), .ZN(n12722) );
  XOR2_X1 U12746 ( .A(n12726), .B(n12727), .Z(n12385) );
  XOR2_X1 U12747 ( .A(n12728), .B(n12729), .Z(n12726) );
  NOR2_X1 U12748 ( .A1(n12466), .A2(n7782), .ZN(n12729) );
  XNOR2_X1 U12749 ( .A(n12730), .B(n12731), .ZN(n12377) );
  XNOR2_X1 U12750 ( .A(n12732), .B(n12733), .ZN(n12731) );
  XOR2_X1 U12751 ( .A(n12734), .B(n12735), .Z(n12515) );
  XOR2_X1 U12752 ( .A(n12736), .B(n12737), .Z(n12734) );
  XNOR2_X1 U12753 ( .A(n12738), .B(n12739), .ZN(n12366) );
  XNOR2_X1 U12754 ( .A(n12740), .B(n12741), .ZN(n12738) );
  XNOR2_X1 U12755 ( .A(n12742), .B(n12743), .ZN(n12520) );
  XNOR2_X1 U12756 ( .A(n12744), .B(n12745), .ZN(n12742) );
  XNOR2_X1 U12757 ( .A(n12746), .B(n12747), .ZN(n12523) );
  XOR2_X1 U12758 ( .A(n12748), .B(n12749), .Z(n12747) );
  XOR2_X1 U12759 ( .A(n12750), .B(n12751), .Z(n12528) );
  XNOR2_X1 U12760 ( .A(n12752), .B(n12753), .ZN(n12751) );
  XNOR2_X1 U12761 ( .A(n12754), .B(n12755), .ZN(n12532) );
  XNOR2_X1 U12762 ( .A(n12756), .B(n12757), .ZN(n12755) );
  XNOR2_X1 U12763 ( .A(n12758), .B(n12759), .ZN(n12536) );
  XNOR2_X1 U12764 ( .A(n12760), .B(n12761), .ZN(n12758) );
  NOR2_X1 U12765 ( .A1(n12466), .A2(n7393), .ZN(n12761) );
  XOR2_X1 U12766 ( .A(n12762), .B(n12763), .Z(n12540) );
  XNOR2_X1 U12767 ( .A(n12764), .B(n12765), .ZN(n12763) );
  NAND2_X1 U12768 ( .A1(a_4_), .A2(b_8_), .ZN(n12765) );
  XOR2_X1 U12769 ( .A(n12766), .B(n12767), .Z(n12544) );
  XOR2_X1 U12770 ( .A(n12768), .B(n12769), .Z(n12766) );
  NOR2_X1 U12771 ( .A1(n12466), .A2(n7850), .ZN(n12769) );
  XOR2_X1 U12772 ( .A(n12770), .B(n12771), .Z(n12548) );
  XNOR2_X1 U12773 ( .A(n12772), .B(n12773), .ZN(n12771) );
  NAND2_X1 U12774 ( .A1(a_2_), .A2(b_8_), .ZN(n12773) );
  XOR2_X1 U12775 ( .A(n12774), .B(n12775), .Z(n12557) );
  XNOR2_X1 U12776 ( .A(n12776), .B(n12777), .ZN(n12775) );
  NAND2_X1 U12777 ( .A1(a_1_), .A2(b_8_), .ZN(n12777) );
  XNOR2_X1 U12778 ( .A(n12554), .B(n12555), .ZN(n12563) );
  XNOR2_X1 U12779 ( .A(n12778), .B(n12779), .ZN(n12554) );
  NOR2_X1 U12780 ( .A1(n7613), .A2(n12466), .ZN(n12779) );
  NAND2_X1 U12781 ( .A1(n12780), .A2(n12781), .ZN(n7259) );
  NAND2_X1 U12782 ( .A1(n12782), .A2(n12783), .ZN(n12781) );
  NAND2_X1 U12783 ( .A1(n12562), .A2(n12561), .ZN(n12780) );
  NAND4_X1 U12784 ( .A1(n12562), .A2(n12782), .A3(n12783), .A4(n12561), .ZN(
        n7260) );
  NAND2_X1 U12785 ( .A1(n12784), .A2(n12785), .ZN(n12561) );
  NAND3_X1 U12786 ( .A1(a_0_), .A2(n12786), .A3(b_8_), .ZN(n12785) );
  OR2_X1 U12787 ( .A1(n12778), .A2(n12555), .ZN(n12786) );
  NAND2_X1 U12788 ( .A1(n12555), .A2(n12778), .ZN(n12784) );
  NAND2_X1 U12789 ( .A1(n12787), .A2(n12788), .ZN(n12778) );
  NAND3_X1 U12790 ( .A1(b_8_), .A2(n12789), .A3(a_1_), .ZN(n12788) );
  NAND2_X1 U12791 ( .A1(n12776), .A2(n12774), .ZN(n12789) );
  OR2_X1 U12792 ( .A1(n12774), .A2(n12776), .ZN(n12787) );
  AND2_X1 U12793 ( .A1(n12790), .A2(n12791), .ZN(n12776) );
  NAND3_X1 U12794 ( .A1(b_8_), .A2(n12792), .A3(a_2_), .ZN(n12791) );
  NAND2_X1 U12795 ( .A1(n12772), .A2(n12770), .ZN(n12792) );
  OR2_X1 U12796 ( .A1(n12770), .A2(n12772), .ZN(n12790) );
  AND2_X1 U12797 ( .A1(n12793), .A2(n12794), .ZN(n12772) );
  NAND3_X1 U12798 ( .A1(b_8_), .A2(n12795), .A3(a_3_), .ZN(n12794) );
  OR2_X1 U12799 ( .A1(n12768), .A2(n12767), .ZN(n12795) );
  NAND2_X1 U12800 ( .A1(n12767), .A2(n12768), .ZN(n12793) );
  NAND2_X1 U12801 ( .A1(n12796), .A2(n12797), .ZN(n12768) );
  NAND3_X1 U12802 ( .A1(b_8_), .A2(n12798), .A3(a_4_), .ZN(n12797) );
  NAND2_X1 U12803 ( .A1(n12764), .A2(n12762), .ZN(n12798) );
  OR2_X1 U12804 ( .A1(n12762), .A2(n12764), .ZN(n12796) );
  AND2_X1 U12805 ( .A1(n12799), .A2(n12800), .ZN(n12764) );
  NAND3_X1 U12806 ( .A1(b_8_), .A2(n12801), .A3(a_5_), .ZN(n12800) );
  NAND2_X1 U12807 ( .A1(n12760), .A2(n12759), .ZN(n12801) );
  OR2_X1 U12808 ( .A1(n12759), .A2(n12760), .ZN(n12799) );
  AND2_X1 U12809 ( .A1(n12802), .A2(n12803), .ZN(n12760) );
  NAND2_X1 U12810 ( .A1(n12757), .A2(n12804), .ZN(n12803) );
  OR2_X1 U12811 ( .A1(n12756), .A2(n12754), .ZN(n12804) );
  NOR2_X1 U12812 ( .A1(n7388), .A2(n12466), .ZN(n12757) );
  NAND2_X1 U12813 ( .A1(n12754), .A2(n12756), .ZN(n12802) );
  NAND2_X1 U12814 ( .A1(n12805), .A2(n12806), .ZN(n12756) );
  NAND2_X1 U12815 ( .A1(n12753), .A2(n12807), .ZN(n12806) );
  NAND2_X1 U12816 ( .A1(n12750), .A2(n12752), .ZN(n12807) );
  NOR2_X1 U12817 ( .A1(n7863), .A2(n12466), .ZN(n12753) );
  OR2_X1 U12818 ( .A1(n12750), .A2(n12752), .ZN(n12805) );
  NAND2_X1 U12819 ( .A1(n12808), .A2(n12809), .ZN(n12752) );
  NAND2_X1 U12820 ( .A1(n12810), .A2(n12748), .ZN(n12809) );
  NAND2_X1 U12821 ( .A1(n12746), .A2(n12749), .ZN(n12810) );
  OR2_X1 U12822 ( .A1(n12749), .A2(n12746), .ZN(n12808) );
  XOR2_X1 U12823 ( .A(n12811), .B(n12812), .Z(n12746) );
  XOR2_X1 U12824 ( .A(n12813), .B(n12814), .Z(n12811) );
  NOR2_X1 U12825 ( .A1(n7870), .A2(n12673), .ZN(n12814) );
  NAND2_X1 U12826 ( .A1(n12815), .A2(n12816), .ZN(n12749) );
  NAND2_X1 U12827 ( .A1(n12745), .A2(n12817), .ZN(n12816) );
  NAND2_X1 U12828 ( .A1(n12744), .A2(n12743), .ZN(n12817) );
  NOR2_X1 U12829 ( .A1(n12466), .A2(n7870), .ZN(n12745) );
  OR2_X1 U12830 ( .A1(n12743), .A2(n12744), .ZN(n12815) );
  AND2_X1 U12831 ( .A1(n12818), .A2(n12819), .ZN(n12744) );
  NAND2_X1 U12832 ( .A1(n12596), .A2(n12820), .ZN(n12819) );
  OR2_X1 U12833 ( .A1(n12595), .A2(n12593), .ZN(n12820) );
  NOR2_X1 U12834 ( .A1(n7799), .A2(n12466), .ZN(n12596) );
  NAND2_X1 U12835 ( .A1(n12593), .A2(n12595), .ZN(n12818) );
  NAND2_X1 U12836 ( .A1(n12821), .A2(n12822), .ZN(n12595) );
  NAND2_X1 U12837 ( .A1(n12741), .A2(n12823), .ZN(n12822) );
  NAND2_X1 U12838 ( .A1(n12740), .A2(n12739), .ZN(n12823) );
  NOR2_X1 U12839 ( .A1(n7877), .A2(n12466), .ZN(n12741) );
  OR2_X1 U12840 ( .A1(n12739), .A2(n12740), .ZN(n12821) );
  AND2_X1 U12841 ( .A1(n12824), .A2(n12825), .ZN(n12740) );
  NAND2_X1 U12842 ( .A1(n12737), .A2(n12826), .ZN(n12825) );
  OR2_X1 U12843 ( .A1(n12735), .A2(n12736), .ZN(n12826) );
  NOR2_X1 U12844 ( .A1(n8020), .A2(n12466), .ZN(n12737) );
  NAND2_X1 U12845 ( .A1(n12735), .A2(n12736), .ZN(n12824) );
  NAND2_X1 U12846 ( .A1(n12827), .A2(n12828), .ZN(n12736) );
  NAND2_X1 U12847 ( .A1(n12733), .A2(n12829), .ZN(n12828) );
  OR2_X1 U12848 ( .A1(n12732), .A2(n12730), .ZN(n12829) );
  NOR2_X1 U12849 ( .A1(n7355), .A2(n12466), .ZN(n12733) );
  NAND2_X1 U12850 ( .A1(n12730), .A2(n12732), .ZN(n12827) );
  NAND2_X1 U12851 ( .A1(n12830), .A2(n12831), .ZN(n12732) );
  NAND3_X1 U12852 ( .A1(b_8_), .A2(n12832), .A3(a_14_), .ZN(n12831) );
  OR2_X1 U12853 ( .A1(n12727), .A2(n12728), .ZN(n12832) );
  NAND2_X1 U12854 ( .A1(n12727), .A2(n12728), .ZN(n12830) );
  NAND2_X1 U12855 ( .A1(n12833), .A2(n12834), .ZN(n12728) );
  NAND2_X1 U12856 ( .A1(n12725), .A2(n12835), .ZN(n12834) );
  NAND2_X1 U12857 ( .A1(n12724), .A2(n12723), .ZN(n12835) );
  NOR2_X1 U12858 ( .A1(n7346), .A2(n12466), .ZN(n12725) );
  OR2_X1 U12859 ( .A1(n12723), .A2(n12724), .ZN(n12833) );
  AND2_X1 U12860 ( .A1(n12720), .A2(n12836), .ZN(n12724) );
  NAND2_X1 U12861 ( .A1(n12719), .A2(n12721), .ZN(n12836) );
  NAND2_X1 U12862 ( .A1(n12837), .A2(n12838), .ZN(n12721) );
  NAND2_X1 U12863 ( .A1(a_16_), .A2(b_8_), .ZN(n12838) );
  INV_X1 U12864 ( .A(n12839), .ZN(n12837) );
  XNOR2_X1 U12865 ( .A(n12840), .B(n12841), .ZN(n12719) );
  XNOR2_X1 U12866 ( .A(n12842), .B(n12843), .ZN(n12840) );
  NOR2_X1 U12867 ( .A1(n12673), .A2(n7337), .ZN(n12843) );
  NAND2_X1 U12868 ( .A1(a_16_), .A2(n12839), .ZN(n12720) );
  NAND2_X1 U12869 ( .A1(n12716), .A2(n12844), .ZN(n12839) );
  NAND2_X1 U12870 ( .A1(n12715), .A2(n12717), .ZN(n12844) );
  NAND2_X1 U12871 ( .A1(n12845), .A2(n12846), .ZN(n12717) );
  NAND2_X1 U12872 ( .A1(a_17_), .A2(b_8_), .ZN(n12846) );
  INV_X1 U12873 ( .A(n12847), .ZN(n12845) );
  XNOR2_X1 U12874 ( .A(n12848), .B(n12849), .ZN(n12715) );
  XOR2_X1 U12875 ( .A(n12850), .B(n12851), .Z(n12849) );
  NAND2_X1 U12876 ( .A1(a_18_), .A2(b_7_), .ZN(n12851) );
  NAND2_X1 U12877 ( .A1(a_17_), .A2(n12847), .ZN(n12716) );
  NAND2_X1 U12878 ( .A1(n12852), .A2(n12853), .ZN(n12847) );
  NAND3_X1 U12879 ( .A1(b_8_), .A2(n12854), .A3(a_18_), .ZN(n12853) );
  OR2_X1 U12880 ( .A1(n12710), .A2(n12712), .ZN(n12854) );
  NAND2_X1 U12881 ( .A1(n12710), .A2(n12712), .ZN(n12852) );
  NAND2_X1 U12882 ( .A1(n12855), .A2(n12856), .ZN(n12712) );
  NAND2_X1 U12883 ( .A1(n12709), .A2(n12857), .ZN(n12856) );
  OR2_X1 U12884 ( .A1(n12707), .A2(n12708), .ZN(n12857) );
  NOR2_X1 U12885 ( .A1(n7902), .A2(n12466), .ZN(n12709) );
  NAND2_X1 U12886 ( .A1(n12707), .A2(n12708), .ZN(n12855) );
  NAND2_X1 U12887 ( .A1(n12858), .A2(n12859), .ZN(n12708) );
  NAND2_X1 U12888 ( .A1(n12705), .A2(n12860), .ZN(n12859) );
  NAND2_X1 U12889 ( .A1(n12704), .A2(n12703), .ZN(n12860) );
  NOR2_X1 U12890 ( .A1(n7987), .A2(n12466), .ZN(n12705) );
  OR2_X1 U12891 ( .A1(n12703), .A2(n12704), .ZN(n12858) );
  AND2_X1 U12892 ( .A1(n12861), .A2(n12862), .ZN(n12704) );
  NAND2_X1 U12893 ( .A1(n12701), .A2(n12863), .ZN(n12862) );
  NAND2_X1 U12894 ( .A1(n12700), .A2(n12699), .ZN(n12863) );
  NOR2_X1 U12895 ( .A1(n7909), .A2(n12466), .ZN(n12701) );
  OR2_X1 U12896 ( .A1(n12699), .A2(n12700), .ZN(n12861) );
  AND2_X1 U12897 ( .A1(n12864), .A2(n12865), .ZN(n12700) );
  NAND2_X1 U12898 ( .A1(n12697), .A2(n12866), .ZN(n12865) );
  OR2_X1 U12899 ( .A1(n12696), .A2(n12694), .ZN(n12866) );
  NOR2_X1 U12900 ( .A1(n12466), .A2(n7312), .ZN(n12697) );
  NAND2_X1 U12901 ( .A1(n12694), .A2(n12696), .ZN(n12864) );
  NAND2_X1 U12902 ( .A1(n12867), .A2(n12868), .ZN(n12696) );
  NAND3_X1 U12903 ( .A1(a_23_), .A2(n12869), .A3(b_8_), .ZN(n12868) );
  OR2_X1 U12904 ( .A1(n12692), .A2(n12690), .ZN(n12869) );
  NAND2_X1 U12905 ( .A1(n12690), .A2(n12692), .ZN(n12867) );
  NAND2_X1 U12906 ( .A1(n12870), .A2(n12871), .ZN(n12692) );
  NAND3_X1 U12907 ( .A1(b_8_), .A2(n12872), .A3(a_24_), .ZN(n12871) );
  NAND2_X1 U12908 ( .A1(n12688), .A2(n12687), .ZN(n12872) );
  OR2_X1 U12909 ( .A1(n12687), .A2(n12688), .ZN(n12870) );
  AND2_X1 U12910 ( .A1(n12873), .A2(n12874), .ZN(n12688) );
  NAND2_X1 U12911 ( .A1(n12685), .A2(n12875), .ZN(n12874) );
  OR2_X1 U12912 ( .A1(n12683), .A2(n12684), .ZN(n12875) );
  NOR2_X1 U12913 ( .A1(n12466), .A2(n7923), .ZN(n12685) );
  NAND2_X1 U12914 ( .A1(n12683), .A2(n12684), .ZN(n12873) );
  NAND2_X1 U12915 ( .A1(n12680), .A2(n12876), .ZN(n12684) );
  NAND2_X1 U12916 ( .A1(n12679), .A2(n12681), .ZN(n12876) );
  NAND2_X1 U12917 ( .A1(n12877), .A2(n12878), .ZN(n12681) );
  NAND2_X1 U12918 ( .A1(a_26_), .A2(b_8_), .ZN(n12878) );
  INV_X1 U12919 ( .A(n12879), .ZN(n12877) );
  XNOR2_X1 U12920 ( .A(n12880), .B(n12881), .ZN(n12679) );
  NAND2_X1 U12921 ( .A1(n12882), .A2(n12883), .ZN(n12880) );
  NAND2_X1 U12922 ( .A1(a_26_), .A2(n12879), .ZN(n12680) );
  NAND2_X1 U12923 ( .A1(n12651), .A2(n12884), .ZN(n12879) );
  NAND2_X1 U12924 ( .A1(n12650), .A2(n12652), .ZN(n12884) );
  NAND2_X1 U12925 ( .A1(n12885), .A2(n12886), .ZN(n12652) );
  NAND2_X1 U12926 ( .A1(a_27_), .A2(b_8_), .ZN(n12886) );
  INV_X1 U12927 ( .A(n12887), .ZN(n12885) );
  XNOR2_X1 U12928 ( .A(n12888), .B(n12889), .ZN(n12650) );
  XOR2_X1 U12929 ( .A(n12890), .B(n12891), .Z(n12888) );
  NAND2_X1 U12930 ( .A1(a_28_), .A2(b_7_), .ZN(n12890) );
  NAND2_X1 U12931 ( .A1(a_27_), .A2(n12887), .ZN(n12651) );
  NAND2_X1 U12932 ( .A1(n12892), .A2(n12893), .ZN(n12887) );
  NAND3_X1 U12933 ( .A1(b_8_), .A2(n12894), .A3(a_28_), .ZN(n12893) );
  NAND2_X1 U12934 ( .A1(n12660), .A2(n12658), .ZN(n12894) );
  OR2_X1 U12935 ( .A1(n12658), .A2(n12660), .ZN(n12892) );
  AND2_X1 U12936 ( .A1(n12895), .A2(n12896), .ZN(n12660) );
  NAND2_X1 U12937 ( .A1(n12675), .A2(n12897), .ZN(n12896) );
  OR2_X1 U12938 ( .A1(n12676), .A2(n12677), .ZN(n12897) );
  NOR2_X1 U12939 ( .A1(n12466), .A2(n7946), .ZN(n12675) );
  NAND2_X1 U12940 ( .A1(n12677), .A2(n12676), .ZN(n12895) );
  NAND2_X1 U12941 ( .A1(n12898), .A2(n12899), .ZN(n12676) );
  NAND2_X1 U12942 ( .A1(b_6_), .A2(n12900), .ZN(n12899) );
  NAND2_X1 U12943 ( .A1(n7268), .A2(n12901), .ZN(n12900) );
  NAND2_X1 U12944 ( .A1(a_31_), .A2(n12673), .ZN(n12901) );
  NAND2_X1 U12945 ( .A1(b_7_), .A2(n12902), .ZN(n12898) );
  NAND2_X1 U12946 ( .A1(n7272), .A2(n12903), .ZN(n12902) );
  NAND2_X1 U12947 ( .A1(a_30_), .A2(n12904), .ZN(n12903) );
  AND3_X1 U12948 ( .A1(b_8_), .A2(n7954), .A3(b_7_), .ZN(n12677) );
  XNOR2_X1 U12949 ( .A(n12905), .B(n12906), .ZN(n12658) );
  XOR2_X1 U12950 ( .A(n12907), .B(n12908), .Z(n12905) );
  XNOR2_X1 U12951 ( .A(n12909), .B(n12910), .ZN(n12683) );
  NAND2_X1 U12952 ( .A1(n12911), .A2(n12912), .ZN(n12909) );
  XNOR2_X1 U12953 ( .A(n12913), .B(n12914), .ZN(n12687) );
  XOR2_X1 U12954 ( .A(n12915), .B(n12916), .Z(n12913) );
  XOR2_X1 U12955 ( .A(n12917), .B(n12918), .Z(n12690) );
  XOR2_X1 U12956 ( .A(n12919), .B(n12920), .Z(n12917) );
  XOR2_X1 U12957 ( .A(n12921), .B(n12922), .Z(n12694) );
  XOR2_X1 U12958 ( .A(n12923), .B(n12924), .Z(n12921) );
  NOR2_X1 U12959 ( .A1(n7916), .A2(n12673), .ZN(n12924) );
  XOR2_X1 U12960 ( .A(n12925), .B(n12926), .Z(n12699) );
  NAND2_X1 U12961 ( .A1(n12927), .A2(n12928), .ZN(n12925) );
  XNOR2_X1 U12962 ( .A(n12929), .B(n12930), .ZN(n12703) );
  XOR2_X1 U12963 ( .A(n12931), .B(n12932), .Z(n12929) );
  NOR2_X1 U12964 ( .A1(n12673), .A2(n7909), .ZN(n12932) );
  XNOR2_X1 U12965 ( .A(n12933), .B(n12934), .ZN(n12707) );
  XNOR2_X1 U12966 ( .A(n12935), .B(n12936), .ZN(n12933) );
  NOR2_X1 U12967 ( .A1(n12673), .A2(n7987), .ZN(n12936) );
  XNOR2_X1 U12968 ( .A(n12937), .B(n12938), .ZN(n12710) );
  XOR2_X1 U12969 ( .A(n12939), .B(n12940), .Z(n12938) );
  NAND2_X1 U12970 ( .A1(a_19_), .A2(b_7_), .ZN(n12940) );
  XOR2_X1 U12971 ( .A(n12941), .B(n12942), .Z(n12723) );
  XOR2_X1 U12972 ( .A(n12943), .B(n12944), .Z(n12942) );
  NAND2_X1 U12973 ( .A1(a_16_), .A2(b_7_), .ZN(n12944) );
  XNOR2_X1 U12974 ( .A(n12945), .B(n12946), .ZN(n12727) );
  XNOR2_X1 U12975 ( .A(n12947), .B(n12948), .ZN(n12945) );
  NOR2_X1 U12976 ( .A1(n12673), .A2(n7346), .ZN(n12948) );
  XOR2_X1 U12977 ( .A(n12949), .B(n12950), .Z(n12730) );
  XOR2_X1 U12978 ( .A(n12951), .B(n12952), .Z(n12949) );
  NOR2_X1 U12979 ( .A1(n12673), .A2(n7782), .ZN(n12952) );
  XNOR2_X1 U12980 ( .A(n12953), .B(n12954), .ZN(n12735) );
  XOR2_X1 U12981 ( .A(n12955), .B(n12956), .Z(n12954) );
  NAND2_X1 U12982 ( .A1(a_13_), .A2(b_7_), .ZN(n12956) );
  XNOR2_X1 U12983 ( .A(n12957), .B(n12958), .ZN(n12739) );
  XOR2_X1 U12984 ( .A(n12959), .B(n12960), .Z(n12957) );
  NOR2_X1 U12985 ( .A1(n12673), .A2(n8020), .ZN(n12960) );
  XOR2_X1 U12986 ( .A(n12961), .B(n12962), .Z(n12593) );
  XOR2_X1 U12987 ( .A(n12963), .B(n12964), .Z(n12961) );
  NOR2_X1 U12988 ( .A1(n12673), .A2(n7877), .ZN(n12964) );
  XNOR2_X1 U12989 ( .A(n12965), .B(n12966), .ZN(n12743) );
  XOR2_X1 U12990 ( .A(n12967), .B(n12968), .Z(n12965) );
  NOR2_X1 U12991 ( .A1(n12673), .A2(n7799), .ZN(n12968) );
  XNOR2_X1 U12992 ( .A(n12969), .B(n12970), .ZN(n12750) );
  XOR2_X1 U12993 ( .A(n12971), .B(n12972), .Z(n12969) );
  NOR2_X1 U12994 ( .A1(n12673), .A2(n8037), .ZN(n12972) );
  XOR2_X1 U12995 ( .A(n12973), .B(n12974), .Z(n12754) );
  XOR2_X1 U12996 ( .A(n12975), .B(n12976), .Z(n12973) );
  XNOR2_X1 U12997 ( .A(n12977), .B(n12978), .ZN(n12759) );
  XOR2_X1 U12998 ( .A(n12979), .B(n12980), .Z(n12977) );
  NOR2_X1 U12999 ( .A1(n12673), .A2(n7388), .ZN(n12980) );
  XNOR2_X1 U13000 ( .A(n12981), .B(n12982), .ZN(n12762) );
  XOR2_X1 U13001 ( .A(n12983), .B(n12984), .Z(n12981) );
  NOR2_X1 U13002 ( .A1(n12673), .A2(n7393), .ZN(n12984) );
  XOR2_X1 U13003 ( .A(n12985), .B(n12986), .Z(n12767) );
  XOR2_X1 U13004 ( .A(n12987), .B(n12988), .Z(n12985) );
  NOR2_X1 U13005 ( .A1(n12673), .A2(n7398), .ZN(n12988) );
  XNOR2_X1 U13006 ( .A(n12989), .B(n12990), .ZN(n12770) );
  XOR2_X1 U13007 ( .A(n12991), .B(n12992), .Z(n12989) );
  NOR2_X1 U13008 ( .A1(n12673), .A2(n7850), .ZN(n12992) );
  XNOR2_X1 U13009 ( .A(n12993), .B(n12994), .ZN(n12774) );
  XOR2_X1 U13010 ( .A(n12995), .B(n12996), .Z(n12993) );
  NOR2_X1 U13011 ( .A1(n12673), .A2(n7832), .ZN(n12996) );
  XOR2_X1 U13012 ( .A(n12997), .B(n12998), .Z(n12555) );
  XOR2_X1 U13013 ( .A(n12999), .B(n13000), .Z(n12997) );
  NOR2_X1 U13014 ( .A1(n12673), .A2(n7411), .ZN(n13000) );
  NAND3_X1 U13015 ( .A1(n13001), .A2(n13002), .A3(n13003), .ZN(n12782) );
  XOR2_X1 U13016 ( .A(n13004), .B(n13005), .Z(n13003) );
  INV_X1 U13017 ( .A(n13006), .ZN(n13004) );
  XOR2_X1 U13018 ( .A(n13007), .B(n13008), .Z(n12562) );
  XOR2_X1 U13019 ( .A(n13009), .B(n13010), .Z(n13007) );
  NAND2_X1 U13020 ( .A1(n13011), .A2(n12783), .ZN(n7263) );
  OR2_X1 U13021 ( .A1(n12783), .A2(n13011), .ZN(n7264) );
  XNOR2_X1 U13022 ( .A(n13012), .B(n13013), .ZN(n13011) );
  NAND2_X1 U13023 ( .A1(n13014), .A2(n13015), .ZN(n12783) );
  NAND2_X1 U13024 ( .A1(n13001), .A2(n13002), .ZN(n13015) );
  NAND2_X1 U13025 ( .A1(n13010), .A2(n13016), .ZN(n13002) );
  OR2_X1 U13026 ( .A1(n13008), .A2(n13009), .ZN(n13016) );
  NOR2_X1 U13027 ( .A1(n12673), .A2(n7613), .ZN(n13010) );
  NAND2_X1 U13028 ( .A1(n13008), .A2(n13009), .ZN(n13001) );
  NAND2_X1 U13029 ( .A1(n13017), .A2(n13018), .ZN(n13009) );
  NAND3_X1 U13030 ( .A1(b_7_), .A2(n13019), .A3(a_1_), .ZN(n13018) );
  OR2_X1 U13031 ( .A1(n12998), .A2(n12999), .ZN(n13019) );
  NAND2_X1 U13032 ( .A1(n12998), .A2(n12999), .ZN(n13017) );
  NAND2_X1 U13033 ( .A1(n13020), .A2(n13021), .ZN(n12999) );
  NAND3_X1 U13034 ( .A1(b_7_), .A2(n13022), .A3(a_2_), .ZN(n13021) );
  OR2_X1 U13035 ( .A1(n12994), .A2(n12995), .ZN(n13022) );
  NAND2_X1 U13036 ( .A1(n12994), .A2(n12995), .ZN(n13020) );
  NAND2_X1 U13037 ( .A1(n13023), .A2(n13024), .ZN(n12995) );
  NAND3_X1 U13038 ( .A1(b_7_), .A2(n13025), .A3(a_3_), .ZN(n13024) );
  OR2_X1 U13039 ( .A1(n12990), .A2(n12991), .ZN(n13025) );
  NAND2_X1 U13040 ( .A1(n12990), .A2(n12991), .ZN(n13023) );
  NAND2_X1 U13041 ( .A1(n13026), .A2(n13027), .ZN(n12991) );
  NAND3_X1 U13042 ( .A1(b_7_), .A2(n13028), .A3(a_4_), .ZN(n13027) );
  OR2_X1 U13043 ( .A1(n12986), .A2(n12987), .ZN(n13028) );
  NAND2_X1 U13044 ( .A1(n12986), .A2(n12987), .ZN(n13026) );
  NAND2_X1 U13045 ( .A1(n13029), .A2(n13030), .ZN(n12987) );
  NAND3_X1 U13046 ( .A1(b_7_), .A2(n13031), .A3(a_5_), .ZN(n13030) );
  OR2_X1 U13047 ( .A1(n12982), .A2(n12983), .ZN(n13031) );
  NAND2_X1 U13048 ( .A1(n12982), .A2(n12983), .ZN(n13029) );
  NAND2_X1 U13049 ( .A1(n13032), .A2(n13033), .ZN(n12983) );
  NAND3_X1 U13050 ( .A1(b_7_), .A2(n13034), .A3(a_6_), .ZN(n13033) );
  OR2_X1 U13051 ( .A1(n12978), .A2(n12979), .ZN(n13034) );
  NAND2_X1 U13052 ( .A1(n12978), .A2(n12979), .ZN(n13032) );
  NAND2_X1 U13053 ( .A1(n13035), .A2(n13036), .ZN(n12979) );
  NAND2_X1 U13054 ( .A1(n12974), .A2(n13037), .ZN(n13036) );
  OR2_X1 U13055 ( .A1(n12975), .A2(n12976), .ZN(n13037) );
  XNOR2_X1 U13056 ( .A(n13038), .B(n13039), .ZN(n12974) );
  XOR2_X1 U13057 ( .A(n13040), .B(n13041), .Z(n13039) );
  NAND2_X1 U13058 ( .A1(a_8_), .A2(b_6_), .ZN(n13041) );
  NAND2_X1 U13059 ( .A1(n12976), .A2(n12975), .ZN(n13035) );
  NAND2_X1 U13060 ( .A1(n13042), .A2(n13043), .ZN(n12975) );
  NAND3_X1 U13061 ( .A1(b_7_), .A2(n13044), .A3(a_8_), .ZN(n13043) );
  OR2_X1 U13062 ( .A1(n12970), .A2(n12971), .ZN(n13044) );
  NAND2_X1 U13063 ( .A1(n12970), .A2(n12971), .ZN(n13042) );
  NAND2_X1 U13064 ( .A1(n13045), .A2(n13046), .ZN(n12971) );
  NAND3_X1 U13065 ( .A1(a_9_), .A2(n13047), .A3(b_7_), .ZN(n13046) );
  OR2_X1 U13066 ( .A1(n12812), .A2(n12813), .ZN(n13047) );
  NAND2_X1 U13067 ( .A1(n12812), .A2(n12813), .ZN(n13045) );
  NAND2_X1 U13068 ( .A1(n13048), .A2(n13049), .ZN(n12813) );
  NAND3_X1 U13069 ( .A1(b_7_), .A2(n13050), .A3(a_10_), .ZN(n13049) );
  OR2_X1 U13070 ( .A1(n12966), .A2(n12967), .ZN(n13050) );
  NAND2_X1 U13071 ( .A1(n12966), .A2(n12967), .ZN(n13048) );
  NAND2_X1 U13072 ( .A1(n13051), .A2(n13052), .ZN(n12967) );
  NAND3_X1 U13073 ( .A1(b_7_), .A2(n13053), .A3(a_11_), .ZN(n13052) );
  OR2_X1 U13074 ( .A1(n12962), .A2(n12963), .ZN(n13053) );
  NAND2_X1 U13075 ( .A1(n12962), .A2(n12963), .ZN(n13051) );
  NAND2_X1 U13076 ( .A1(n13054), .A2(n13055), .ZN(n12963) );
  NAND3_X1 U13077 ( .A1(b_7_), .A2(n13056), .A3(a_12_), .ZN(n13055) );
  OR2_X1 U13078 ( .A1(n12958), .A2(n12959), .ZN(n13056) );
  NAND2_X1 U13079 ( .A1(n12958), .A2(n12959), .ZN(n13054) );
  NAND2_X1 U13080 ( .A1(n13057), .A2(n13058), .ZN(n12959) );
  NAND3_X1 U13081 ( .A1(b_7_), .A2(n13059), .A3(a_13_), .ZN(n13058) );
  OR2_X1 U13082 ( .A1(n12955), .A2(n12953), .ZN(n13059) );
  NAND2_X1 U13083 ( .A1(n12953), .A2(n12955), .ZN(n13057) );
  NAND2_X1 U13084 ( .A1(n13060), .A2(n13061), .ZN(n12955) );
  NAND3_X1 U13085 ( .A1(b_7_), .A2(n13062), .A3(a_14_), .ZN(n13061) );
  OR2_X1 U13086 ( .A1(n12950), .A2(n12951), .ZN(n13062) );
  NAND2_X1 U13087 ( .A1(n12950), .A2(n12951), .ZN(n13060) );
  NAND2_X1 U13088 ( .A1(n13063), .A2(n13064), .ZN(n12951) );
  NAND3_X1 U13089 ( .A1(b_7_), .A2(n13065), .A3(a_15_), .ZN(n13064) );
  NAND2_X1 U13090 ( .A1(n12947), .A2(n12946), .ZN(n13065) );
  OR2_X1 U13091 ( .A1(n12946), .A2(n12947), .ZN(n13063) );
  AND2_X1 U13092 ( .A1(n13066), .A2(n13067), .ZN(n12947) );
  NAND3_X1 U13093 ( .A1(b_7_), .A2(n13068), .A3(a_16_), .ZN(n13067) );
  OR2_X1 U13094 ( .A1(n12941), .A2(n12943), .ZN(n13068) );
  NAND2_X1 U13095 ( .A1(n12941), .A2(n12943), .ZN(n13066) );
  NAND2_X1 U13096 ( .A1(n13069), .A2(n13070), .ZN(n12943) );
  NAND3_X1 U13097 ( .A1(b_7_), .A2(n13071), .A3(a_17_), .ZN(n13070) );
  NAND2_X1 U13098 ( .A1(n12842), .A2(n12841), .ZN(n13071) );
  OR2_X1 U13099 ( .A1(n12841), .A2(n12842), .ZN(n13069) );
  AND2_X1 U13100 ( .A1(n13072), .A2(n13073), .ZN(n12842) );
  NAND3_X1 U13101 ( .A1(b_7_), .A2(n13074), .A3(a_18_), .ZN(n13073) );
  OR2_X1 U13102 ( .A1(n12848), .A2(n12850), .ZN(n13074) );
  NAND2_X1 U13103 ( .A1(n12848), .A2(n12850), .ZN(n13072) );
  NAND2_X1 U13104 ( .A1(n13075), .A2(n13076), .ZN(n12850) );
  NAND3_X1 U13105 ( .A1(b_7_), .A2(n13077), .A3(a_19_), .ZN(n13076) );
  OR2_X1 U13106 ( .A1(n12939), .A2(n12937), .ZN(n13077) );
  NAND2_X1 U13107 ( .A1(n12937), .A2(n12939), .ZN(n13075) );
  NAND2_X1 U13108 ( .A1(n13078), .A2(n13079), .ZN(n12939) );
  NAND3_X1 U13109 ( .A1(b_7_), .A2(n13080), .A3(a_20_), .ZN(n13079) );
  NAND2_X1 U13110 ( .A1(n12935), .A2(n12934), .ZN(n13080) );
  OR2_X1 U13111 ( .A1(n12934), .A2(n12935), .ZN(n13078) );
  AND2_X1 U13112 ( .A1(n13081), .A2(n13082), .ZN(n12935) );
  NAND3_X1 U13113 ( .A1(b_7_), .A2(n13083), .A3(a_21_), .ZN(n13082) );
  OR2_X1 U13114 ( .A1(n12930), .A2(n12931), .ZN(n13083) );
  NAND2_X1 U13115 ( .A1(n12930), .A2(n12931), .ZN(n13081) );
  NAND2_X1 U13116 ( .A1(n12927), .A2(n13084), .ZN(n12931) );
  NAND2_X1 U13117 ( .A1(n12926), .A2(n12928), .ZN(n13084) );
  NAND2_X1 U13118 ( .A1(n13085), .A2(n13086), .ZN(n12928) );
  NAND2_X1 U13119 ( .A1(b_7_), .A2(a_22_), .ZN(n13086) );
  INV_X1 U13120 ( .A(n13087), .ZN(n13085) );
  XOR2_X1 U13121 ( .A(n13088), .B(n13089), .Z(n12926) );
  XOR2_X1 U13122 ( .A(n13090), .B(n13091), .Z(n13088) );
  NOR2_X1 U13123 ( .A1(n7916), .A2(n12904), .ZN(n13091) );
  NAND2_X1 U13124 ( .A1(a_22_), .A2(n13087), .ZN(n12927) );
  NAND2_X1 U13125 ( .A1(n13092), .A2(n13093), .ZN(n13087) );
  NAND3_X1 U13126 ( .A1(a_23_), .A2(n13094), .A3(b_7_), .ZN(n13093) );
  OR2_X1 U13127 ( .A1(n12922), .A2(n12923), .ZN(n13094) );
  NAND2_X1 U13128 ( .A1(n12922), .A2(n12923), .ZN(n13092) );
  NAND2_X1 U13129 ( .A1(n13095), .A2(n13096), .ZN(n12923) );
  NAND2_X1 U13130 ( .A1(n12920), .A2(n13097), .ZN(n13096) );
  OR2_X1 U13131 ( .A1(n12918), .A2(n12919), .ZN(n13097) );
  NOR2_X1 U13132 ( .A1(n7691), .A2(n12673), .ZN(n12920) );
  NAND2_X1 U13133 ( .A1(n12918), .A2(n12919), .ZN(n13095) );
  NAND2_X1 U13134 ( .A1(n13098), .A2(n13099), .ZN(n12919) );
  NAND2_X1 U13135 ( .A1(n12916), .A2(n13100), .ZN(n13099) );
  OR2_X1 U13136 ( .A1(n12914), .A2(n12915), .ZN(n13100) );
  NOR2_X1 U13137 ( .A1(n12673), .A2(n7923), .ZN(n12916) );
  NAND2_X1 U13138 ( .A1(n12914), .A2(n12915), .ZN(n13098) );
  NAND2_X1 U13139 ( .A1(n12911), .A2(n13101), .ZN(n12915) );
  NAND2_X1 U13140 ( .A1(n12910), .A2(n12912), .ZN(n13101) );
  NAND2_X1 U13141 ( .A1(n13102), .A2(n13103), .ZN(n12912) );
  NAND2_X1 U13142 ( .A1(a_26_), .A2(b_7_), .ZN(n13103) );
  INV_X1 U13143 ( .A(n13104), .ZN(n13102) );
  XNOR2_X1 U13144 ( .A(n13105), .B(n13106), .ZN(n12910) );
  NAND2_X1 U13145 ( .A1(n13107), .A2(n13108), .ZN(n13105) );
  NAND2_X1 U13146 ( .A1(a_26_), .A2(n13104), .ZN(n12911) );
  NAND2_X1 U13147 ( .A1(n12882), .A2(n13109), .ZN(n13104) );
  NAND2_X1 U13148 ( .A1(n12881), .A2(n12883), .ZN(n13109) );
  NAND2_X1 U13149 ( .A1(n13110), .A2(n13111), .ZN(n12883) );
  NAND2_X1 U13150 ( .A1(a_27_), .A2(b_7_), .ZN(n13111) );
  INV_X1 U13151 ( .A(n13112), .ZN(n13110) );
  XNOR2_X1 U13152 ( .A(n13113), .B(n13114), .ZN(n12881) );
  XOR2_X1 U13153 ( .A(n13115), .B(n13116), .Z(n13113) );
  NAND2_X1 U13154 ( .A1(a_28_), .A2(b_6_), .ZN(n13115) );
  NAND2_X1 U13155 ( .A1(a_27_), .A2(n13112), .ZN(n12882) );
  NAND2_X1 U13156 ( .A1(n13117), .A2(n13118), .ZN(n13112) );
  NAND3_X1 U13157 ( .A1(b_7_), .A2(n13119), .A3(a_28_), .ZN(n13118) );
  NAND2_X1 U13158 ( .A1(n12891), .A2(n12889), .ZN(n13119) );
  OR2_X1 U13159 ( .A1(n12889), .A2(n12891), .ZN(n13117) );
  AND2_X1 U13160 ( .A1(n13120), .A2(n13121), .ZN(n12891) );
  NAND2_X1 U13161 ( .A1(n12906), .A2(n13122), .ZN(n13121) );
  OR2_X1 U13162 ( .A1(n12907), .A2(n12908), .ZN(n13122) );
  NOR2_X1 U13163 ( .A1(n12673), .A2(n7946), .ZN(n12906) );
  NAND2_X1 U13164 ( .A1(n12908), .A2(n12907), .ZN(n13120) );
  NAND2_X1 U13165 ( .A1(n13123), .A2(n13124), .ZN(n12907) );
  NAND2_X1 U13166 ( .A1(b_5_), .A2(n13125), .ZN(n13124) );
  NAND2_X1 U13167 ( .A1(n7268), .A2(n13126), .ZN(n13125) );
  NAND2_X1 U13168 ( .A1(a_31_), .A2(n12904), .ZN(n13126) );
  NAND2_X1 U13169 ( .A1(b_6_), .A2(n13127), .ZN(n13123) );
  NAND2_X1 U13170 ( .A1(n7272), .A2(n13128), .ZN(n13127) );
  NAND2_X1 U13171 ( .A1(a_30_), .A2(n13129), .ZN(n13128) );
  AND3_X1 U13172 ( .A1(b_7_), .A2(n7954), .A3(b_6_), .ZN(n12908) );
  XNOR2_X1 U13173 ( .A(n13130), .B(n13131), .ZN(n12889) );
  XOR2_X1 U13174 ( .A(n13132), .B(n13133), .Z(n13130) );
  XNOR2_X1 U13175 ( .A(n13134), .B(n13135), .ZN(n12914) );
  NAND2_X1 U13176 ( .A1(n13136), .A2(n13137), .ZN(n13134) );
  XNOR2_X1 U13177 ( .A(n13138), .B(n13139), .ZN(n12918) );
  NAND2_X1 U13178 ( .A1(n13140), .A2(n13141), .ZN(n13138) );
  XNOR2_X1 U13179 ( .A(n13142), .B(n13143), .ZN(n12922) );
  XNOR2_X1 U13180 ( .A(n13144), .B(n13145), .ZN(n13143) );
  XNOR2_X1 U13181 ( .A(n13146), .B(n13147), .ZN(n12930) );
  NAND2_X1 U13182 ( .A1(n13148), .A2(n13149), .ZN(n13146) );
  XOR2_X1 U13183 ( .A(n13150), .B(n13151), .Z(n12934) );
  XNOR2_X1 U13184 ( .A(n13152), .B(n13153), .ZN(n13151) );
  XOR2_X1 U13185 ( .A(n13154), .B(n13155), .Z(n12937) );
  XOR2_X1 U13186 ( .A(n13156), .B(n13157), .Z(n13154) );
  NOR2_X1 U13187 ( .A1(n12904), .A2(n7987), .ZN(n13157) );
  XNOR2_X1 U13188 ( .A(n13158), .B(n13159), .ZN(n12848) );
  XNOR2_X1 U13189 ( .A(n13160), .B(n13161), .ZN(n13159) );
  XNOR2_X1 U13190 ( .A(n13162), .B(n13163), .ZN(n12841) );
  XOR2_X1 U13191 ( .A(n13164), .B(n13165), .Z(n13162) );
  XNOR2_X1 U13192 ( .A(n13166), .B(n13167), .ZN(n12941) );
  XNOR2_X1 U13193 ( .A(n13168), .B(n13169), .ZN(n13166) );
  XOR2_X1 U13194 ( .A(n13170), .B(n13171), .Z(n12946) );
  XNOR2_X1 U13195 ( .A(n13172), .B(n13173), .ZN(n13171) );
  XNOR2_X1 U13196 ( .A(n13174), .B(n13175), .ZN(n12950) );
  XNOR2_X1 U13197 ( .A(n13176), .B(n13177), .ZN(n13174) );
  XOR2_X1 U13198 ( .A(n13178), .B(n13179), .Z(n12953) );
  XOR2_X1 U13199 ( .A(n13180), .B(n13181), .Z(n13178) );
  XNOR2_X1 U13200 ( .A(n13182), .B(n13183), .ZN(n12958) );
  XNOR2_X1 U13201 ( .A(n13184), .B(n13185), .ZN(n13182) );
  XNOR2_X1 U13202 ( .A(n13186), .B(n13187), .ZN(n12962) );
  XNOR2_X1 U13203 ( .A(n13188), .B(n13189), .ZN(n13186) );
  XNOR2_X1 U13204 ( .A(n13190), .B(n13191), .ZN(n12966) );
  XNOR2_X1 U13205 ( .A(n13192), .B(n13193), .ZN(n13191) );
  XNOR2_X1 U13206 ( .A(n13194), .B(n13195), .ZN(n12812) );
  XNOR2_X1 U13207 ( .A(n13196), .B(n13197), .ZN(n13194) );
  XNOR2_X1 U13208 ( .A(n13198), .B(n13199), .ZN(n12970) );
  XOR2_X1 U13209 ( .A(n13200), .B(n13201), .Z(n13199) );
  NAND2_X1 U13210 ( .A1(b_6_), .A2(a_9_), .ZN(n13201) );
  XOR2_X1 U13211 ( .A(n13202), .B(n13203), .Z(n12978) );
  XOR2_X1 U13212 ( .A(n13204), .B(n13205), .Z(n13202) );
  NOR2_X1 U13213 ( .A1(n12904), .A2(n7863), .ZN(n13205) );
  XOR2_X1 U13214 ( .A(n13206), .B(n13207), .Z(n12982) );
  XOR2_X1 U13215 ( .A(n13208), .B(n13209), .Z(n13206) );
  XOR2_X1 U13216 ( .A(n13210), .B(n13211), .Z(n12986) );
  XOR2_X1 U13217 ( .A(n13212), .B(n13213), .Z(n13210) );
  NOR2_X1 U13218 ( .A1(n12904), .A2(n7393), .ZN(n13213) );
  XOR2_X1 U13219 ( .A(n13214), .B(n13215), .Z(n12990) );
  XNOR2_X1 U13220 ( .A(n13216), .B(n13217), .ZN(n13215) );
  NAND2_X1 U13221 ( .A1(a_4_), .A2(b_6_), .ZN(n13217) );
  XOR2_X1 U13222 ( .A(n13218), .B(n13219), .Z(n12994) );
  XOR2_X1 U13223 ( .A(n13220), .B(n13221), .Z(n13218) );
  NOR2_X1 U13224 ( .A1(n12904), .A2(n7850), .ZN(n13221) );
  XOR2_X1 U13225 ( .A(n13222), .B(n13223), .Z(n12998) );
  XOR2_X1 U13226 ( .A(n13224), .B(n13225), .Z(n13222) );
  NOR2_X1 U13227 ( .A1(n12904), .A2(n7832), .ZN(n13225) );
  XOR2_X1 U13228 ( .A(n13226), .B(n13227), .Z(n13008) );
  XOR2_X1 U13229 ( .A(n13228), .B(n13229), .Z(n13226) );
  NOR2_X1 U13230 ( .A1(n12904), .A2(n7411), .ZN(n13229) );
  XOR2_X1 U13231 ( .A(n13006), .B(n13005), .Z(n13014) );
  XOR2_X1 U13232 ( .A(n13230), .B(n13231), .Z(n13006) );
  NOR2_X1 U13233 ( .A1(n7613), .A2(n12904), .ZN(n13231) );
  NAND2_X1 U13234 ( .A1(n13232), .A2(n13233), .ZN(n7285) );
  NAND2_X1 U13235 ( .A1(n13234), .A2(n13235), .ZN(n13233) );
  NAND2_X1 U13236 ( .A1(n13013), .A2(n13012), .ZN(n13232) );
  NAND4_X1 U13237 ( .A1(n13013), .A2(n13234), .A3(n13235), .A4(n13012), .ZN(
        n7286) );
  NAND2_X1 U13238 ( .A1(n13236), .A2(n13237), .ZN(n13012) );
  NAND3_X1 U13239 ( .A1(a_0_), .A2(n13238), .A3(b_6_), .ZN(n13237) );
  OR2_X1 U13240 ( .A1(n13005), .A2(n13230), .ZN(n13238) );
  NAND2_X1 U13241 ( .A1(n13005), .A2(n13230), .ZN(n13236) );
  NAND2_X1 U13242 ( .A1(n13239), .A2(n13240), .ZN(n13230) );
  NAND3_X1 U13243 ( .A1(b_6_), .A2(n13241), .A3(a_1_), .ZN(n13240) );
  OR2_X1 U13244 ( .A1(n13228), .A2(n13227), .ZN(n13241) );
  NAND2_X1 U13245 ( .A1(n13227), .A2(n13228), .ZN(n13239) );
  NAND2_X1 U13246 ( .A1(n13242), .A2(n13243), .ZN(n13228) );
  NAND3_X1 U13247 ( .A1(b_6_), .A2(n13244), .A3(a_2_), .ZN(n13243) );
  OR2_X1 U13248 ( .A1(n13224), .A2(n13223), .ZN(n13244) );
  NAND2_X1 U13249 ( .A1(n13223), .A2(n13224), .ZN(n13242) );
  NAND2_X1 U13250 ( .A1(n13245), .A2(n13246), .ZN(n13224) );
  NAND3_X1 U13251 ( .A1(b_6_), .A2(n13247), .A3(a_3_), .ZN(n13246) );
  OR2_X1 U13252 ( .A1(n13220), .A2(n13219), .ZN(n13247) );
  NAND2_X1 U13253 ( .A1(n13219), .A2(n13220), .ZN(n13245) );
  NAND2_X1 U13254 ( .A1(n13248), .A2(n13249), .ZN(n13220) );
  NAND3_X1 U13255 ( .A1(b_6_), .A2(n13250), .A3(a_4_), .ZN(n13249) );
  NAND2_X1 U13256 ( .A1(n13216), .A2(n13214), .ZN(n13250) );
  OR2_X1 U13257 ( .A1(n13214), .A2(n13216), .ZN(n13248) );
  AND2_X1 U13258 ( .A1(n13251), .A2(n13252), .ZN(n13216) );
  NAND3_X1 U13259 ( .A1(b_6_), .A2(n13253), .A3(a_5_), .ZN(n13252) );
  OR2_X1 U13260 ( .A1(n13212), .A2(n13211), .ZN(n13253) );
  NAND2_X1 U13261 ( .A1(n13211), .A2(n13212), .ZN(n13251) );
  NAND2_X1 U13262 ( .A1(n13254), .A2(n13255), .ZN(n13212) );
  NAND2_X1 U13263 ( .A1(n13209), .A2(n13256), .ZN(n13255) );
  OR2_X1 U13264 ( .A1(n13208), .A2(n13207), .ZN(n13256) );
  NAND2_X1 U13265 ( .A1(n13207), .A2(n13208), .ZN(n13254) );
  NAND2_X1 U13266 ( .A1(n13257), .A2(n13258), .ZN(n13208) );
  NAND3_X1 U13267 ( .A1(b_6_), .A2(n13259), .A3(a_7_), .ZN(n13258) );
  OR2_X1 U13268 ( .A1(n13204), .A2(n13203), .ZN(n13259) );
  NAND2_X1 U13269 ( .A1(n13203), .A2(n13204), .ZN(n13257) );
  NAND2_X1 U13270 ( .A1(n13260), .A2(n13261), .ZN(n13204) );
  NAND3_X1 U13271 ( .A1(b_6_), .A2(n13262), .A3(a_8_), .ZN(n13261) );
  OR2_X1 U13272 ( .A1(n13040), .A2(n13038), .ZN(n13262) );
  NAND2_X1 U13273 ( .A1(n13038), .A2(n13040), .ZN(n13260) );
  NAND2_X1 U13274 ( .A1(n13263), .A2(n13264), .ZN(n13040) );
  NAND3_X1 U13275 ( .A1(a_9_), .A2(n13265), .A3(b_6_), .ZN(n13264) );
  OR2_X1 U13276 ( .A1(n13200), .A2(n13198), .ZN(n13265) );
  NAND2_X1 U13277 ( .A1(n13198), .A2(n13200), .ZN(n13263) );
  NAND2_X1 U13278 ( .A1(n13266), .A2(n13267), .ZN(n13200) );
  NAND2_X1 U13279 ( .A1(n13197), .A2(n13268), .ZN(n13267) );
  NAND2_X1 U13280 ( .A1(n13196), .A2(n13195), .ZN(n13268) );
  NOR2_X1 U13281 ( .A1(n7799), .A2(n12904), .ZN(n13197) );
  OR2_X1 U13282 ( .A1(n13195), .A2(n13196), .ZN(n13266) );
  AND2_X1 U13283 ( .A1(n13269), .A2(n13270), .ZN(n13196) );
  NAND2_X1 U13284 ( .A1(n13193), .A2(n13271), .ZN(n13270) );
  OR2_X1 U13285 ( .A1(n13192), .A2(n13190), .ZN(n13271) );
  NOR2_X1 U13286 ( .A1(n7877), .A2(n12904), .ZN(n13193) );
  NAND2_X1 U13287 ( .A1(n13190), .A2(n13192), .ZN(n13269) );
  NAND2_X1 U13288 ( .A1(n13272), .A2(n13273), .ZN(n13192) );
  NAND2_X1 U13289 ( .A1(n13189), .A2(n13274), .ZN(n13273) );
  NAND2_X1 U13290 ( .A1(n13188), .A2(n13187), .ZN(n13274) );
  NOR2_X1 U13291 ( .A1(n8020), .A2(n12904), .ZN(n13189) );
  OR2_X1 U13292 ( .A1(n13187), .A2(n13188), .ZN(n13272) );
  AND2_X1 U13293 ( .A1(n13275), .A2(n13276), .ZN(n13188) );
  NAND2_X1 U13294 ( .A1(n13185), .A2(n13277), .ZN(n13276) );
  NAND2_X1 U13295 ( .A1(n13184), .A2(n13183), .ZN(n13277) );
  NOR2_X1 U13296 ( .A1(n7355), .A2(n12904), .ZN(n13185) );
  OR2_X1 U13297 ( .A1(n13183), .A2(n13184), .ZN(n13275) );
  AND2_X1 U13298 ( .A1(n13278), .A2(n13279), .ZN(n13184) );
  NAND2_X1 U13299 ( .A1(n13181), .A2(n13280), .ZN(n13279) );
  OR2_X1 U13300 ( .A1(n13179), .A2(n13180), .ZN(n13280) );
  NOR2_X1 U13301 ( .A1(n7782), .A2(n12904), .ZN(n13181) );
  NAND2_X1 U13302 ( .A1(n13179), .A2(n13180), .ZN(n13278) );
  NAND2_X1 U13303 ( .A1(n13281), .A2(n13282), .ZN(n13180) );
  NAND2_X1 U13304 ( .A1(n13177), .A2(n13283), .ZN(n13282) );
  NAND2_X1 U13305 ( .A1(n13176), .A2(n13175), .ZN(n13283) );
  NOR2_X1 U13306 ( .A1(n7346), .A2(n12904), .ZN(n13177) );
  OR2_X1 U13307 ( .A1(n13175), .A2(n13176), .ZN(n13281) );
  AND2_X1 U13308 ( .A1(n13284), .A2(n13285), .ZN(n13176) );
  NAND2_X1 U13309 ( .A1(n13173), .A2(n13286), .ZN(n13285) );
  OR2_X1 U13310 ( .A1(n13170), .A2(n13172), .ZN(n13286) );
  NOR2_X1 U13311 ( .A1(n7773), .A2(n12904), .ZN(n13173) );
  NAND2_X1 U13312 ( .A1(n13170), .A2(n13172), .ZN(n13284) );
  NAND2_X1 U13313 ( .A1(n13287), .A2(n13288), .ZN(n13172) );
  NAND2_X1 U13314 ( .A1(n13169), .A2(n13289), .ZN(n13288) );
  NAND2_X1 U13315 ( .A1(n13168), .A2(n13167), .ZN(n13289) );
  NOR2_X1 U13316 ( .A1(n7337), .A2(n12904), .ZN(n13169) );
  OR2_X1 U13317 ( .A1(n13167), .A2(n13168), .ZN(n13287) );
  AND2_X1 U13318 ( .A1(n13290), .A2(n13291), .ZN(n13168) );
  NAND2_X1 U13319 ( .A1(n13165), .A2(n13292), .ZN(n13291) );
  OR2_X1 U13320 ( .A1(n13163), .A2(n13164), .ZN(n13292) );
  NOR2_X1 U13321 ( .A1(n7764), .A2(n12904), .ZN(n13165) );
  NAND2_X1 U13322 ( .A1(n13163), .A2(n13164), .ZN(n13290) );
  NAND2_X1 U13323 ( .A1(n13293), .A2(n13294), .ZN(n13164) );
  NAND2_X1 U13324 ( .A1(n13161), .A2(n13295), .ZN(n13294) );
  OR2_X1 U13325 ( .A1(n13160), .A2(n13158), .ZN(n13295) );
  NOR2_X1 U13326 ( .A1(n7902), .A2(n12904), .ZN(n13161) );
  NAND2_X1 U13327 ( .A1(n13158), .A2(n13160), .ZN(n13293) );
  NAND2_X1 U13328 ( .A1(n13296), .A2(n13297), .ZN(n13160) );
  NAND3_X1 U13329 ( .A1(b_6_), .A2(n13298), .A3(a_20_), .ZN(n13297) );
  OR2_X1 U13330 ( .A1(n13155), .A2(n13156), .ZN(n13298) );
  NAND2_X1 U13331 ( .A1(n13155), .A2(n13156), .ZN(n13296) );
  NAND2_X1 U13332 ( .A1(n13299), .A2(n13300), .ZN(n13156) );
  NAND2_X1 U13333 ( .A1(n13153), .A2(n13301), .ZN(n13300) );
  OR2_X1 U13334 ( .A1(n13150), .A2(n13152), .ZN(n13301) );
  NOR2_X1 U13335 ( .A1(n7909), .A2(n12904), .ZN(n13153) );
  NAND2_X1 U13336 ( .A1(n13150), .A2(n13152), .ZN(n13299) );
  NAND2_X1 U13337 ( .A1(n13148), .A2(n13302), .ZN(n13152) );
  NAND2_X1 U13338 ( .A1(n13147), .A2(n13149), .ZN(n13302) );
  NAND2_X1 U13339 ( .A1(n13303), .A2(n13304), .ZN(n13149) );
  NAND2_X1 U13340 ( .A1(b_6_), .A2(a_22_), .ZN(n13304) );
  INV_X1 U13341 ( .A(n13305), .ZN(n13303) );
  XNOR2_X1 U13342 ( .A(n13306), .B(n13307), .ZN(n13147) );
  XOR2_X1 U13343 ( .A(n13308), .B(n13309), .Z(n13307) );
  NAND2_X1 U13344 ( .A1(b_5_), .A2(a_23_), .ZN(n13309) );
  NAND2_X1 U13345 ( .A1(a_22_), .A2(n13305), .ZN(n13148) );
  NAND2_X1 U13346 ( .A1(n13310), .A2(n13311), .ZN(n13305) );
  NAND3_X1 U13347 ( .A1(a_23_), .A2(n13312), .A3(b_6_), .ZN(n13311) );
  OR2_X1 U13348 ( .A1(n13089), .A2(n13090), .ZN(n13312) );
  NAND2_X1 U13349 ( .A1(n13089), .A2(n13090), .ZN(n13310) );
  NAND2_X1 U13350 ( .A1(n13313), .A2(n13314), .ZN(n13090) );
  NAND2_X1 U13351 ( .A1(n13145), .A2(n13315), .ZN(n13314) );
  OR2_X1 U13352 ( .A1(n13144), .A2(n13142), .ZN(n13315) );
  NOR2_X1 U13353 ( .A1(n7691), .A2(n12904), .ZN(n13145) );
  NAND2_X1 U13354 ( .A1(n13142), .A2(n13144), .ZN(n13313) );
  NAND2_X1 U13355 ( .A1(n13140), .A2(n13316), .ZN(n13144) );
  NAND2_X1 U13356 ( .A1(n13139), .A2(n13141), .ZN(n13316) );
  NAND2_X1 U13357 ( .A1(n13317), .A2(n13318), .ZN(n13141) );
  NAND2_X1 U13358 ( .A1(b_6_), .A2(a_25_), .ZN(n13318) );
  INV_X1 U13359 ( .A(n13319), .ZN(n13317) );
  XNOR2_X1 U13360 ( .A(n13320), .B(n13321), .ZN(n13139) );
  NAND2_X1 U13361 ( .A1(n13322), .A2(n13323), .ZN(n13320) );
  NAND2_X1 U13362 ( .A1(a_25_), .A2(n13319), .ZN(n13140) );
  NAND2_X1 U13363 ( .A1(n13136), .A2(n13324), .ZN(n13319) );
  NAND2_X1 U13364 ( .A1(n13135), .A2(n13137), .ZN(n13324) );
  NAND2_X1 U13365 ( .A1(n13325), .A2(n13326), .ZN(n13137) );
  NAND2_X1 U13366 ( .A1(a_26_), .A2(b_6_), .ZN(n13326) );
  INV_X1 U13367 ( .A(n13327), .ZN(n13325) );
  XNOR2_X1 U13368 ( .A(n13328), .B(n13329), .ZN(n13135) );
  NAND2_X1 U13369 ( .A1(n13330), .A2(n13331), .ZN(n13328) );
  NAND2_X1 U13370 ( .A1(a_26_), .A2(n13327), .ZN(n13136) );
  NAND2_X1 U13371 ( .A1(n13107), .A2(n13332), .ZN(n13327) );
  NAND2_X1 U13372 ( .A1(n13106), .A2(n13108), .ZN(n13332) );
  NAND2_X1 U13373 ( .A1(n13333), .A2(n13334), .ZN(n13108) );
  NAND2_X1 U13374 ( .A1(a_27_), .A2(b_6_), .ZN(n13334) );
  INV_X1 U13375 ( .A(n13335), .ZN(n13333) );
  XNOR2_X1 U13376 ( .A(n13336), .B(n13337), .ZN(n13106) );
  XOR2_X1 U13377 ( .A(n13338), .B(n13339), .Z(n13336) );
  NAND2_X1 U13378 ( .A1(b_5_), .A2(a_28_), .ZN(n13338) );
  NAND2_X1 U13379 ( .A1(a_27_), .A2(n13335), .ZN(n13107) );
  NAND2_X1 U13380 ( .A1(n13340), .A2(n13341), .ZN(n13335) );
  NAND3_X1 U13381 ( .A1(b_6_), .A2(n13342), .A3(a_28_), .ZN(n13341) );
  NAND2_X1 U13382 ( .A1(n13116), .A2(n13114), .ZN(n13342) );
  OR2_X1 U13383 ( .A1(n13114), .A2(n13116), .ZN(n13340) );
  AND2_X1 U13384 ( .A1(n13343), .A2(n13344), .ZN(n13116) );
  NAND2_X1 U13385 ( .A1(n13131), .A2(n13345), .ZN(n13344) );
  OR2_X1 U13386 ( .A1(n13132), .A2(n13133), .ZN(n13345) );
  NOR2_X1 U13387 ( .A1(n12904), .A2(n7946), .ZN(n13131) );
  NAND2_X1 U13388 ( .A1(n13133), .A2(n13132), .ZN(n13343) );
  NAND2_X1 U13389 ( .A1(n13346), .A2(n13347), .ZN(n13132) );
  NAND2_X1 U13390 ( .A1(b_4_), .A2(n13348), .ZN(n13347) );
  NAND2_X1 U13391 ( .A1(n7268), .A2(n13349), .ZN(n13348) );
  NAND2_X1 U13392 ( .A1(a_31_), .A2(n13129), .ZN(n13349) );
  NAND2_X1 U13393 ( .A1(b_5_), .A2(n13350), .ZN(n13346) );
  NAND2_X1 U13394 ( .A1(n7272), .A2(n13351), .ZN(n13350) );
  NAND2_X1 U13395 ( .A1(a_30_), .A2(n13352), .ZN(n13351) );
  AND3_X1 U13396 ( .A1(b_6_), .A2(n7954), .A3(b_5_), .ZN(n13133) );
  XNOR2_X1 U13397 ( .A(n13353), .B(n13354), .ZN(n13114) );
  XOR2_X1 U13398 ( .A(n13355), .B(n13356), .Z(n13353) );
  XNOR2_X1 U13399 ( .A(n13357), .B(n13358), .ZN(n13142) );
  NAND2_X1 U13400 ( .A1(n13359), .A2(n13360), .ZN(n13357) );
  XNOR2_X1 U13401 ( .A(n13361), .B(n13362), .ZN(n13089) );
  XOR2_X1 U13402 ( .A(n13363), .B(n13364), .Z(n13362) );
  NAND2_X1 U13403 ( .A1(a_24_), .A2(b_5_), .ZN(n13364) );
  XNOR2_X1 U13404 ( .A(n13365), .B(n13366), .ZN(n13150) );
  XOR2_X1 U13405 ( .A(n13367), .B(n13368), .Z(n13366) );
  NAND2_X1 U13406 ( .A1(b_5_), .A2(a_22_), .ZN(n13368) );
  XNOR2_X1 U13407 ( .A(n13369), .B(n13370), .ZN(n13155) );
  XOR2_X1 U13408 ( .A(n13371), .B(n13372), .Z(n13370) );
  NAND2_X1 U13409 ( .A1(a_21_), .A2(b_5_), .ZN(n13372) );
  XOR2_X1 U13410 ( .A(n13373), .B(n13374), .Z(n13158) );
  XOR2_X1 U13411 ( .A(n13375), .B(n13376), .Z(n13373) );
  NOR2_X1 U13412 ( .A1(n13129), .A2(n7987), .ZN(n13376) );
  XNOR2_X1 U13413 ( .A(n13377), .B(n13378), .ZN(n13163) );
  XOR2_X1 U13414 ( .A(n13379), .B(n13380), .Z(n13378) );
  NAND2_X1 U13415 ( .A1(a_19_), .A2(b_5_), .ZN(n13380) );
  XNOR2_X1 U13416 ( .A(n13381), .B(n13382), .ZN(n13167) );
  XOR2_X1 U13417 ( .A(n13383), .B(n13384), .Z(n13381) );
  NOR2_X1 U13418 ( .A1(n13129), .A2(n7764), .ZN(n13384) );
  XNOR2_X1 U13419 ( .A(n13385), .B(n13386), .ZN(n13170) );
  XNOR2_X1 U13420 ( .A(n13387), .B(n13388), .ZN(n13385) );
  NOR2_X1 U13421 ( .A1(n13129), .A2(n7337), .ZN(n13388) );
  XNOR2_X1 U13422 ( .A(n13389), .B(n13390), .ZN(n13175) );
  XOR2_X1 U13423 ( .A(n13391), .B(n13392), .Z(n13389) );
  NOR2_X1 U13424 ( .A1(n13129), .A2(n7773), .ZN(n13392) );
  XNOR2_X1 U13425 ( .A(n13393), .B(n13394), .ZN(n13179) );
  XNOR2_X1 U13426 ( .A(n13395), .B(n13396), .ZN(n13393) );
  NOR2_X1 U13427 ( .A1(n13129), .A2(n7346), .ZN(n13396) );
  XNOR2_X1 U13428 ( .A(n13397), .B(n13398), .ZN(n13183) );
  XOR2_X1 U13429 ( .A(n13399), .B(n13400), .Z(n13397) );
  NOR2_X1 U13430 ( .A1(n13129), .A2(n7782), .ZN(n13400) );
  XNOR2_X1 U13431 ( .A(n13401), .B(n13402), .ZN(n13187) );
  XOR2_X1 U13432 ( .A(n13403), .B(n13404), .Z(n13401) );
  NOR2_X1 U13433 ( .A1(n13129), .A2(n7355), .ZN(n13404) );
  XOR2_X1 U13434 ( .A(n13405), .B(n13406), .Z(n13190) );
  XOR2_X1 U13435 ( .A(n13407), .B(n13408), .Z(n13405) );
  NOR2_X1 U13436 ( .A1(n13129), .A2(n8020), .ZN(n13408) );
  XNOR2_X1 U13437 ( .A(n13409), .B(n13410), .ZN(n13195) );
  XOR2_X1 U13438 ( .A(n13411), .B(n13412), .Z(n13409) );
  NOR2_X1 U13439 ( .A1(n13129), .A2(n7877), .ZN(n13412) );
  XOR2_X1 U13440 ( .A(n13413), .B(n13414), .Z(n13198) );
  XOR2_X1 U13441 ( .A(n13415), .B(n13416), .Z(n13413) );
  NOR2_X1 U13442 ( .A1(n13129), .A2(n7799), .ZN(n13416) );
  XNOR2_X1 U13443 ( .A(n13417), .B(n13418), .ZN(n13038) );
  XNOR2_X1 U13444 ( .A(n13419), .B(n13420), .ZN(n13417) );
  NOR2_X1 U13445 ( .A1(n7870), .A2(n13129), .ZN(n13420) );
  XOR2_X1 U13446 ( .A(n13421), .B(n13422), .Z(n13203) );
  XOR2_X1 U13447 ( .A(n13423), .B(n13424), .Z(n13421) );
  NOR2_X1 U13448 ( .A1(n13129), .A2(n8037), .ZN(n13424) );
  XOR2_X1 U13449 ( .A(n13425), .B(n13426), .Z(n13207) );
  XOR2_X1 U13450 ( .A(n13427), .B(n13428), .Z(n13425) );
  NOR2_X1 U13451 ( .A1(n13129), .A2(n7863), .ZN(n13428) );
  XOR2_X1 U13452 ( .A(n13429), .B(n13430), .Z(n13211) );
  XOR2_X1 U13453 ( .A(n13431), .B(n13432), .Z(n13429) );
  NOR2_X1 U13454 ( .A1(n13129), .A2(n7388), .ZN(n13432) );
  XNOR2_X1 U13455 ( .A(n13433), .B(n13434), .ZN(n13214) );
  XOR2_X1 U13456 ( .A(n13435), .B(n13436), .Z(n13433) );
  XOR2_X1 U13457 ( .A(n13437), .B(n13438), .Z(n13219) );
  XOR2_X1 U13458 ( .A(n13439), .B(n13440), .Z(n13437) );
  NOR2_X1 U13459 ( .A1(n13129), .A2(n7398), .ZN(n13440) );
  XOR2_X1 U13460 ( .A(n13441), .B(n13442), .Z(n13223) );
  XOR2_X1 U13461 ( .A(n13443), .B(n13444), .Z(n13441) );
  NOR2_X1 U13462 ( .A1(n13129), .A2(n7850), .ZN(n13444) );
  XOR2_X1 U13463 ( .A(n13445), .B(n13446), .Z(n13227) );
  XOR2_X1 U13464 ( .A(n13447), .B(n13448), .Z(n13445) );
  NOR2_X1 U13465 ( .A1(n13129), .A2(n7832), .ZN(n13448) );
  XOR2_X1 U13466 ( .A(n13449), .B(n13450), .Z(n13005) );
  XOR2_X1 U13467 ( .A(n13451), .B(n13452), .Z(n13449) );
  NOR2_X1 U13468 ( .A1(n13129), .A2(n7411), .ZN(n13452) );
  NAND3_X1 U13469 ( .A1(n13453), .A2(n13454), .A3(n13455), .ZN(n13234) );
  XOR2_X1 U13470 ( .A(n13456), .B(n13457), .Z(n13455) );
  INV_X1 U13471 ( .A(n13458), .ZN(n13456) );
  XOR2_X1 U13472 ( .A(n13459), .B(n13460), .Z(n13013) );
  XOR2_X1 U13473 ( .A(n13461), .B(n13462), .Z(n13459) );
  NAND2_X1 U13474 ( .A1(n13463), .A2(n13235), .ZN(n7331) );
  OR2_X1 U13475 ( .A1(n13235), .A2(n13463), .ZN(n7332) );
  XNOR2_X1 U13476 ( .A(n13464), .B(n13465), .ZN(n13463) );
  NAND2_X1 U13477 ( .A1(n13466), .A2(n13467), .ZN(n13235) );
  NAND2_X1 U13478 ( .A1(n13453), .A2(n13454), .ZN(n13467) );
  NAND2_X1 U13479 ( .A1(n13462), .A2(n13468), .ZN(n13454) );
  OR2_X1 U13480 ( .A1(n13460), .A2(n13461), .ZN(n13468) );
  NOR2_X1 U13481 ( .A1(n13129), .A2(n7613), .ZN(n13462) );
  NAND2_X1 U13482 ( .A1(n13460), .A2(n13461), .ZN(n13453) );
  NAND2_X1 U13483 ( .A1(n13469), .A2(n13470), .ZN(n13461) );
  NAND3_X1 U13484 ( .A1(b_5_), .A2(n13471), .A3(a_1_), .ZN(n13470) );
  OR2_X1 U13485 ( .A1(n13451), .A2(n13450), .ZN(n13471) );
  NAND2_X1 U13486 ( .A1(n13450), .A2(n13451), .ZN(n13469) );
  NAND2_X1 U13487 ( .A1(n13472), .A2(n13473), .ZN(n13451) );
  NAND3_X1 U13488 ( .A1(b_5_), .A2(n13474), .A3(a_2_), .ZN(n13473) );
  OR2_X1 U13489 ( .A1(n13446), .A2(n13447), .ZN(n13474) );
  NAND2_X1 U13490 ( .A1(n13446), .A2(n13447), .ZN(n13472) );
  NAND2_X1 U13491 ( .A1(n13475), .A2(n13476), .ZN(n13447) );
  NAND3_X1 U13492 ( .A1(b_5_), .A2(n13477), .A3(a_3_), .ZN(n13476) );
  OR2_X1 U13493 ( .A1(n13442), .A2(n13443), .ZN(n13477) );
  NAND2_X1 U13494 ( .A1(n13442), .A2(n13443), .ZN(n13475) );
  NAND2_X1 U13495 ( .A1(n13478), .A2(n13479), .ZN(n13443) );
  NAND3_X1 U13496 ( .A1(b_5_), .A2(n13480), .A3(a_4_), .ZN(n13479) );
  OR2_X1 U13497 ( .A1(n13438), .A2(n13439), .ZN(n13480) );
  NAND2_X1 U13498 ( .A1(n13438), .A2(n13439), .ZN(n13478) );
  NAND2_X1 U13499 ( .A1(n13481), .A2(n13482), .ZN(n13439) );
  NAND2_X1 U13500 ( .A1(n13434), .A2(n13483), .ZN(n13482) );
  OR2_X1 U13501 ( .A1(n13435), .A2(n13436), .ZN(n13483) );
  XNOR2_X1 U13502 ( .A(n13484), .B(n13485), .ZN(n13434) );
  XNOR2_X1 U13503 ( .A(n13486), .B(n13487), .ZN(n13484) );
  NOR2_X1 U13504 ( .A1(n13352), .A2(n7388), .ZN(n13487) );
  NAND2_X1 U13505 ( .A1(n13436), .A2(n13435), .ZN(n13481) );
  NAND2_X1 U13506 ( .A1(n13488), .A2(n13489), .ZN(n13435) );
  NAND3_X1 U13507 ( .A1(b_5_), .A2(n13490), .A3(a_6_), .ZN(n13489) );
  OR2_X1 U13508 ( .A1(n13430), .A2(n13431), .ZN(n13490) );
  NAND2_X1 U13509 ( .A1(n13430), .A2(n13431), .ZN(n13488) );
  NAND2_X1 U13510 ( .A1(n13491), .A2(n13492), .ZN(n13431) );
  NAND3_X1 U13511 ( .A1(b_5_), .A2(n13493), .A3(a_7_), .ZN(n13492) );
  OR2_X1 U13512 ( .A1(n13426), .A2(n13427), .ZN(n13493) );
  NAND2_X1 U13513 ( .A1(n13426), .A2(n13427), .ZN(n13491) );
  NAND2_X1 U13514 ( .A1(n13494), .A2(n13495), .ZN(n13427) );
  NAND3_X1 U13515 ( .A1(b_5_), .A2(n13496), .A3(a_8_), .ZN(n13495) );
  OR2_X1 U13516 ( .A1(n13422), .A2(n13423), .ZN(n13496) );
  NAND2_X1 U13517 ( .A1(n13422), .A2(n13423), .ZN(n13494) );
  NAND2_X1 U13518 ( .A1(n13497), .A2(n13498), .ZN(n13423) );
  NAND3_X1 U13519 ( .A1(a_9_), .A2(n13499), .A3(b_5_), .ZN(n13498) );
  NAND2_X1 U13520 ( .A1(n13418), .A2(n13419), .ZN(n13499) );
  OR2_X1 U13521 ( .A1(n13418), .A2(n13419), .ZN(n13497) );
  AND2_X1 U13522 ( .A1(n13500), .A2(n13501), .ZN(n13419) );
  NAND3_X1 U13523 ( .A1(b_5_), .A2(n13502), .A3(a_10_), .ZN(n13501) );
  OR2_X1 U13524 ( .A1(n13414), .A2(n13415), .ZN(n13502) );
  NAND2_X1 U13525 ( .A1(n13414), .A2(n13415), .ZN(n13500) );
  NAND2_X1 U13526 ( .A1(n13503), .A2(n13504), .ZN(n13415) );
  NAND3_X1 U13527 ( .A1(b_5_), .A2(n13505), .A3(a_11_), .ZN(n13504) );
  OR2_X1 U13528 ( .A1(n13410), .A2(n13411), .ZN(n13505) );
  NAND2_X1 U13529 ( .A1(n13410), .A2(n13411), .ZN(n13503) );
  NAND2_X1 U13530 ( .A1(n13506), .A2(n13507), .ZN(n13411) );
  NAND3_X1 U13531 ( .A1(b_5_), .A2(n13508), .A3(a_12_), .ZN(n13507) );
  OR2_X1 U13532 ( .A1(n13406), .A2(n13407), .ZN(n13508) );
  NAND2_X1 U13533 ( .A1(n13406), .A2(n13407), .ZN(n13506) );
  NAND2_X1 U13534 ( .A1(n13509), .A2(n13510), .ZN(n13407) );
  NAND3_X1 U13535 ( .A1(b_5_), .A2(n13511), .A3(a_13_), .ZN(n13510) );
  OR2_X1 U13536 ( .A1(n13402), .A2(n13403), .ZN(n13511) );
  NAND2_X1 U13537 ( .A1(n13402), .A2(n13403), .ZN(n13509) );
  NAND2_X1 U13538 ( .A1(n13512), .A2(n13513), .ZN(n13403) );
  NAND3_X1 U13539 ( .A1(b_5_), .A2(n13514), .A3(a_14_), .ZN(n13513) );
  OR2_X1 U13540 ( .A1(n13398), .A2(n13399), .ZN(n13514) );
  NAND2_X1 U13541 ( .A1(n13398), .A2(n13399), .ZN(n13512) );
  NAND2_X1 U13542 ( .A1(n13515), .A2(n13516), .ZN(n13399) );
  NAND3_X1 U13543 ( .A1(b_5_), .A2(n13517), .A3(a_15_), .ZN(n13516) );
  NAND2_X1 U13544 ( .A1(n13395), .A2(n13394), .ZN(n13517) );
  OR2_X1 U13545 ( .A1(n13394), .A2(n13395), .ZN(n13515) );
  AND2_X1 U13546 ( .A1(n13518), .A2(n13519), .ZN(n13395) );
  NAND3_X1 U13547 ( .A1(b_5_), .A2(n13520), .A3(a_16_), .ZN(n13519) );
  OR2_X1 U13548 ( .A1(n13390), .A2(n13391), .ZN(n13520) );
  NAND2_X1 U13549 ( .A1(n13390), .A2(n13391), .ZN(n13518) );
  NAND2_X1 U13550 ( .A1(n13521), .A2(n13522), .ZN(n13391) );
  NAND3_X1 U13551 ( .A1(b_5_), .A2(n13523), .A3(a_17_), .ZN(n13522) );
  NAND2_X1 U13552 ( .A1(n13387), .A2(n13386), .ZN(n13523) );
  OR2_X1 U13553 ( .A1(n13386), .A2(n13387), .ZN(n13521) );
  AND2_X1 U13554 ( .A1(n13524), .A2(n13525), .ZN(n13387) );
  NAND3_X1 U13555 ( .A1(b_5_), .A2(n13526), .A3(a_18_), .ZN(n13525) );
  OR2_X1 U13556 ( .A1(n13382), .A2(n13383), .ZN(n13526) );
  NAND2_X1 U13557 ( .A1(n13382), .A2(n13383), .ZN(n13524) );
  NAND2_X1 U13558 ( .A1(n13527), .A2(n13528), .ZN(n13383) );
  NAND3_X1 U13559 ( .A1(b_5_), .A2(n13529), .A3(a_19_), .ZN(n13528) );
  OR2_X1 U13560 ( .A1(n13379), .A2(n13377), .ZN(n13529) );
  NAND2_X1 U13561 ( .A1(n13377), .A2(n13379), .ZN(n13527) );
  NAND2_X1 U13562 ( .A1(n13530), .A2(n13531), .ZN(n13379) );
  NAND3_X1 U13563 ( .A1(b_5_), .A2(n13532), .A3(a_20_), .ZN(n13531) );
  OR2_X1 U13564 ( .A1(n13374), .A2(n13375), .ZN(n13532) );
  NAND2_X1 U13565 ( .A1(n13374), .A2(n13375), .ZN(n13530) );
  NAND2_X1 U13566 ( .A1(n13533), .A2(n13534), .ZN(n13375) );
  NAND3_X1 U13567 ( .A1(b_5_), .A2(n13535), .A3(a_21_), .ZN(n13534) );
  OR2_X1 U13568 ( .A1(n13371), .A2(n13369), .ZN(n13535) );
  NAND2_X1 U13569 ( .A1(n13369), .A2(n13371), .ZN(n13533) );
  NAND2_X1 U13570 ( .A1(n13536), .A2(n13537), .ZN(n13371) );
  NAND3_X1 U13571 ( .A1(a_22_), .A2(n13538), .A3(b_5_), .ZN(n13537) );
  OR2_X1 U13572 ( .A1(n13367), .A2(n13365), .ZN(n13538) );
  NAND2_X1 U13573 ( .A1(n13365), .A2(n13367), .ZN(n13536) );
  NAND2_X1 U13574 ( .A1(n13539), .A2(n13540), .ZN(n13367) );
  NAND3_X1 U13575 ( .A1(a_23_), .A2(n13541), .A3(b_5_), .ZN(n13540) );
  OR2_X1 U13576 ( .A1(n13308), .A2(n13306), .ZN(n13541) );
  NAND2_X1 U13577 ( .A1(n13306), .A2(n13308), .ZN(n13539) );
  NAND2_X1 U13578 ( .A1(n13542), .A2(n13543), .ZN(n13308) );
  NAND3_X1 U13579 ( .A1(b_5_), .A2(n13544), .A3(a_24_), .ZN(n13543) );
  OR2_X1 U13580 ( .A1(n13363), .A2(n13361), .ZN(n13544) );
  NAND2_X1 U13581 ( .A1(n13361), .A2(n13363), .ZN(n13542) );
  NAND2_X1 U13582 ( .A1(n13359), .A2(n13545), .ZN(n13363) );
  NAND2_X1 U13583 ( .A1(n13358), .A2(n13360), .ZN(n13545) );
  NAND2_X1 U13584 ( .A1(n13546), .A2(n13547), .ZN(n13360) );
  NAND2_X1 U13585 ( .A1(b_5_), .A2(a_25_), .ZN(n13547) );
  INV_X1 U13586 ( .A(n13548), .ZN(n13546) );
  XNOR2_X1 U13587 ( .A(n13549), .B(n13550), .ZN(n13358) );
  NAND2_X1 U13588 ( .A1(n13551), .A2(n13552), .ZN(n13549) );
  NAND2_X1 U13589 ( .A1(a_25_), .A2(n13548), .ZN(n13359) );
  NAND2_X1 U13590 ( .A1(n13322), .A2(n13553), .ZN(n13548) );
  NAND2_X1 U13591 ( .A1(n13321), .A2(n13323), .ZN(n13553) );
  NAND2_X1 U13592 ( .A1(n13554), .A2(n13555), .ZN(n13323) );
  NAND2_X1 U13593 ( .A1(a_26_), .A2(b_5_), .ZN(n13555) );
  INV_X1 U13594 ( .A(n13556), .ZN(n13554) );
  XNOR2_X1 U13595 ( .A(n13557), .B(n13558), .ZN(n13321) );
  NAND2_X1 U13596 ( .A1(n13559), .A2(n13560), .ZN(n13557) );
  NAND2_X1 U13597 ( .A1(a_26_), .A2(n13556), .ZN(n13322) );
  NAND2_X1 U13598 ( .A1(n13330), .A2(n13561), .ZN(n13556) );
  NAND2_X1 U13599 ( .A1(n13329), .A2(n13331), .ZN(n13561) );
  NAND2_X1 U13600 ( .A1(n13562), .A2(n13563), .ZN(n13331) );
  NAND2_X1 U13601 ( .A1(b_5_), .A2(a_27_), .ZN(n13563) );
  INV_X1 U13602 ( .A(n13564), .ZN(n13562) );
  XNOR2_X1 U13603 ( .A(n13565), .B(n13566), .ZN(n13329) );
  XOR2_X1 U13604 ( .A(n13567), .B(n13568), .Z(n13565) );
  NAND2_X1 U13605 ( .A1(b_4_), .A2(a_28_), .ZN(n13567) );
  NAND2_X1 U13606 ( .A1(a_27_), .A2(n13564), .ZN(n13330) );
  NAND2_X1 U13607 ( .A1(n13569), .A2(n13570), .ZN(n13564) );
  NAND3_X1 U13608 ( .A1(a_28_), .A2(n13571), .A3(b_5_), .ZN(n13570) );
  NAND2_X1 U13609 ( .A1(n13339), .A2(n13337), .ZN(n13571) );
  OR2_X1 U13610 ( .A1(n13337), .A2(n13339), .ZN(n13569) );
  AND2_X1 U13611 ( .A1(n13572), .A2(n13573), .ZN(n13339) );
  NAND2_X1 U13612 ( .A1(n13354), .A2(n13574), .ZN(n13573) );
  OR2_X1 U13613 ( .A1(n13355), .A2(n13356), .ZN(n13574) );
  NOR2_X1 U13614 ( .A1(n13129), .A2(n7946), .ZN(n13354) );
  NAND2_X1 U13615 ( .A1(n13356), .A2(n13355), .ZN(n13572) );
  NAND2_X1 U13616 ( .A1(n13575), .A2(n13576), .ZN(n13355) );
  NAND2_X1 U13617 ( .A1(b_3_), .A2(n13577), .ZN(n13576) );
  NAND2_X1 U13618 ( .A1(n7268), .A2(n13578), .ZN(n13577) );
  NAND2_X1 U13619 ( .A1(a_31_), .A2(n13352), .ZN(n13578) );
  NAND2_X1 U13620 ( .A1(b_4_), .A2(n13579), .ZN(n13575) );
  NAND2_X1 U13621 ( .A1(n7272), .A2(n13580), .ZN(n13579) );
  NAND2_X1 U13622 ( .A1(a_30_), .A2(n13581), .ZN(n13580) );
  AND3_X1 U13623 ( .A1(b_5_), .A2(n7954), .A3(b_4_), .ZN(n13356) );
  XNOR2_X1 U13624 ( .A(n13582), .B(n13583), .ZN(n13337) );
  XOR2_X1 U13625 ( .A(n13584), .B(n13585), .Z(n13582) );
  XOR2_X1 U13626 ( .A(n13586), .B(n13587), .Z(n13361) );
  XOR2_X1 U13627 ( .A(n13588), .B(n13589), .Z(n13586) );
  XOR2_X1 U13628 ( .A(n13590), .B(n13591), .Z(n13306) );
  XOR2_X1 U13629 ( .A(n13592), .B(n13593), .Z(n13590) );
  XOR2_X1 U13630 ( .A(n13594), .B(n13595), .Z(n13365) );
  XOR2_X1 U13631 ( .A(n13596), .B(n13597), .Z(n13594) );
  XNOR2_X1 U13632 ( .A(n13598), .B(n13599), .ZN(n13369) );
  XNOR2_X1 U13633 ( .A(n13600), .B(n13601), .ZN(n13599) );
  XNOR2_X1 U13634 ( .A(n13602), .B(n13603), .ZN(n13374) );
  XNOR2_X1 U13635 ( .A(n13604), .B(n13605), .ZN(n13602) );
  XOR2_X1 U13636 ( .A(n13606), .B(n13607), .Z(n13377) );
  XOR2_X1 U13637 ( .A(n13608), .B(n13609), .Z(n13606) );
  XNOR2_X1 U13638 ( .A(n13610), .B(n13611), .ZN(n13382) );
  XNOR2_X1 U13639 ( .A(n13612), .B(n13613), .ZN(n13610) );
  XNOR2_X1 U13640 ( .A(n13614), .B(n13615), .ZN(n13386) );
  XOR2_X1 U13641 ( .A(n13616), .B(n13617), .Z(n13614) );
  XNOR2_X1 U13642 ( .A(n13618), .B(n13619), .ZN(n13390) );
  XNOR2_X1 U13643 ( .A(n13620), .B(n13621), .ZN(n13618) );
  XNOR2_X1 U13644 ( .A(n13622), .B(n13623), .ZN(n13394) );
  XOR2_X1 U13645 ( .A(n13624), .B(n13625), .Z(n13622) );
  XNOR2_X1 U13646 ( .A(n13626), .B(n13627), .ZN(n13398) );
  XNOR2_X1 U13647 ( .A(n13628), .B(n13629), .ZN(n13626) );
  XNOR2_X1 U13648 ( .A(n13630), .B(n13631), .ZN(n13402) );
  XNOR2_X1 U13649 ( .A(n13632), .B(n13633), .ZN(n13630) );
  XNOR2_X1 U13650 ( .A(n13634), .B(n13635), .ZN(n13406) );
  XNOR2_X1 U13651 ( .A(n13636), .B(n13637), .ZN(n13634) );
  NOR2_X1 U13652 ( .A1(n13352), .A2(n7355), .ZN(n13637) );
  XNOR2_X1 U13653 ( .A(n13638), .B(n13639), .ZN(n13410) );
  XNOR2_X1 U13654 ( .A(n13640), .B(n13641), .ZN(n13638) );
  NOR2_X1 U13655 ( .A1(n13352), .A2(n8020), .ZN(n13641) );
  XOR2_X1 U13656 ( .A(n13642), .B(n13643), .Z(n13414) );
  XNOR2_X1 U13657 ( .A(n13644), .B(n13645), .ZN(n13643) );
  NAND2_X1 U13658 ( .A1(a_11_), .A2(b_4_), .ZN(n13645) );
  XNOR2_X1 U13659 ( .A(n13646), .B(n13647), .ZN(n13418) );
  XNOR2_X1 U13660 ( .A(n13648), .B(n13649), .ZN(n13647) );
  NAND2_X1 U13661 ( .A1(a_10_), .A2(b_4_), .ZN(n13649) );
  XOR2_X1 U13662 ( .A(n13650), .B(n13651), .Z(n13422) );
  XNOR2_X1 U13663 ( .A(n13652), .B(n13653), .ZN(n13651) );
  NAND2_X1 U13664 ( .A1(b_4_), .A2(a_9_), .ZN(n13653) );
  XOR2_X1 U13665 ( .A(n13654), .B(n13655), .Z(n13426) );
  XNOR2_X1 U13666 ( .A(n13656), .B(n13657), .ZN(n13655) );
  NAND2_X1 U13667 ( .A1(a_8_), .A2(b_4_), .ZN(n13657) );
  XOR2_X1 U13668 ( .A(n13658), .B(n13659), .Z(n13430) );
  XOR2_X1 U13669 ( .A(n13660), .B(n13661), .Z(n13658) );
  NOR2_X1 U13670 ( .A1(n13352), .A2(n7863), .ZN(n13661) );
  XOR2_X1 U13671 ( .A(n13662), .B(n13663), .Z(n13438) );
  XOR2_X1 U13672 ( .A(n13664), .B(n13665), .Z(n13662) );
  NOR2_X1 U13673 ( .A1(n13352), .A2(n7393), .ZN(n13665) );
  XOR2_X1 U13674 ( .A(n13666), .B(n13667), .Z(n13442) );
  XOR2_X1 U13675 ( .A(n13668), .B(n13669), .Z(n13666) );
  XOR2_X1 U13676 ( .A(n13670), .B(n13671), .Z(n13446) );
  XOR2_X1 U13677 ( .A(n13672), .B(n13673), .Z(n13670) );
  NOR2_X1 U13678 ( .A1(n13352), .A2(n7850), .ZN(n13673) );
  XOR2_X1 U13679 ( .A(n13674), .B(n13675), .Z(n13450) );
  XOR2_X1 U13680 ( .A(n13676), .B(n13677), .Z(n13674) );
  NOR2_X1 U13681 ( .A1(n13352), .A2(n7832), .ZN(n13677) );
  XOR2_X1 U13682 ( .A(n13678), .B(n13679), .Z(n13460) );
  XOR2_X1 U13683 ( .A(n13680), .B(n13681), .Z(n13678) );
  NOR2_X1 U13684 ( .A1(n13352), .A2(n7411), .ZN(n13681) );
  XOR2_X1 U13685 ( .A(n13458), .B(n13457), .Z(n13466) );
  XOR2_X1 U13686 ( .A(n13682), .B(n13683), .Z(n13458) );
  NOR2_X1 U13687 ( .A1(n7613), .A2(n13352), .ZN(n13683) );
  NAND2_X1 U13688 ( .A1(n13684), .A2(n13685), .ZN(n7378) );
  NAND2_X1 U13689 ( .A1(n13686), .A2(n13687), .ZN(n13685) );
  NAND2_X1 U13690 ( .A1(n13465), .A2(n13464), .ZN(n13684) );
  NAND4_X1 U13691 ( .A1(n13465), .A2(n13686), .A3(n13464), .A4(n13687), .ZN(
        n7379) );
  NAND2_X1 U13692 ( .A1(n13688), .A2(n13689), .ZN(n13464) );
  NAND3_X1 U13693 ( .A1(a_0_), .A2(n13690), .A3(b_4_), .ZN(n13689) );
  OR2_X1 U13694 ( .A1(n13457), .A2(n13682), .ZN(n13690) );
  NAND2_X1 U13695 ( .A1(n13457), .A2(n13682), .ZN(n13688) );
  NAND2_X1 U13696 ( .A1(n13691), .A2(n13692), .ZN(n13682) );
  NAND3_X1 U13697 ( .A1(b_4_), .A2(n13693), .A3(a_1_), .ZN(n13692) );
  OR2_X1 U13698 ( .A1(n13680), .A2(n13679), .ZN(n13693) );
  NAND2_X1 U13699 ( .A1(n13679), .A2(n13680), .ZN(n13691) );
  NAND2_X1 U13700 ( .A1(n13694), .A2(n13695), .ZN(n13680) );
  NAND3_X1 U13701 ( .A1(b_4_), .A2(n13696), .A3(a_2_), .ZN(n13695) );
  OR2_X1 U13702 ( .A1(n13675), .A2(n13676), .ZN(n13696) );
  NAND2_X1 U13703 ( .A1(n13675), .A2(n13676), .ZN(n13694) );
  NAND2_X1 U13704 ( .A1(n13697), .A2(n13698), .ZN(n13676) );
  NAND3_X1 U13705 ( .A1(b_4_), .A2(n13699), .A3(a_3_), .ZN(n13698) );
  OR2_X1 U13706 ( .A1(n13672), .A2(n13671), .ZN(n13699) );
  NAND2_X1 U13707 ( .A1(n13671), .A2(n13672), .ZN(n13697) );
  NAND2_X1 U13708 ( .A1(n13700), .A2(n13701), .ZN(n13672) );
  NAND2_X1 U13709 ( .A1(n13669), .A2(n13702), .ZN(n13701) );
  OR2_X1 U13710 ( .A1(n13668), .A2(n13667), .ZN(n13702) );
  NAND2_X1 U13711 ( .A1(n13667), .A2(n13668), .ZN(n13700) );
  NAND2_X1 U13712 ( .A1(n13703), .A2(n13704), .ZN(n13668) );
  NAND3_X1 U13713 ( .A1(b_4_), .A2(n13705), .A3(a_5_), .ZN(n13704) );
  OR2_X1 U13714 ( .A1(n13664), .A2(n13663), .ZN(n13705) );
  NAND2_X1 U13715 ( .A1(n13663), .A2(n13664), .ZN(n13703) );
  NAND2_X1 U13716 ( .A1(n13706), .A2(n13707), .ZN(n13664) );
  NAND3_X1 U13717 ( .A1(b_4_), .A2(n13708), .A3(a_6_), .ZN(n13707) );
  NAND2_X1 U13718 ( .A1(n13486), .A2(n13485), .ZN(n13708) );
  OR2_X1 U13719 ( .A1(n13485), .A2(n13486), .ZN(n13706) );
  AND2_X1 U13720 ( .A1(n13709), .A2(n13710), .ZN(n13486) );
  NAND3_X1 U13721 ( .A1(b_4_), .A2(n13711), .A3(a_7_), .ZN(n13710) );
  OR2_X1 U13722 ( .A1(n13660), .A2(n13659), .ZN(n13711) );
  NAND2_X1 U13723 ( .A1(n13659), .A2(n13660), .ZN(n13709) );
  NAND2_X1 U13724 ( .A1(n13712), .A2(n13713), .ZN(n13660) );
  NAND3_X1 U13725 ( .A1(b_4_), .A2(n13714), .A3(a_8_), .ZN(n13713) );
  NAND2_X1 U13726 ( .A1(n13656), .A2(n13654), .ZN(n13714) );
  OR2_X1 U13727 ( .A1(n13654), .A2(n13656), .ZN(n13712) );
  AND2_X1 U13728 ( .A1(n13715), .A2(n13716), .ZN(n13656) );
  NAND3_X1 U13729 ( .A1(a_9_), .A2(n13717), .A3(b_4_), .ZN(n13716) );
  NAND2_X1 U13730 ( .A1(n13652), .A2(n13650), .ZN(n13717) );
  OR2_X1 U13731 ( .A1(n13650), .A2(n13652), .ZN(n13715) );
  AND2_X1 U13732 ( .A1(n13718), .A2(n13719), .ZN(n13652) );
  NAND3_X1 U13733 ( .A1(b_4_), .A2(n13720), .A3(a_10_), .ZN(n13719) );
  NAND2_X1 U13734 ( .A1(n13648), .A2(n13646), .ZN(n13720) );
  OR2_X1 U13735 ( .A1(n13646), .A2(n13648), .ZN(n13718) );
  AND2_X1 U13736 ( .A1(n13721), .A2(n13722), .ZN(n13648) );
  NAND3_X1 U13737 ( .A1(b_4_), .A2(n13723), .A3(a_11_), .ZN(n13722) );
  NAND2_X1 U13738 ( .A1(n13644), .A2(n13642), .ZN(n13723) );
  OR2_X1 U13739 ( .A1(n13642), .A2(n13644), .ZN(n13721) );
  AND2_X1 U13740 ( .A1(n13724), .A2(n13725), .ZN(n13644) );
  NAND3_X1 U13741 ( .A1(b_4_), .A2(n13726), .A3(a_12_), .ZN(n13725) );
  NAND2_X1 U13742 ( .A1(n13640), .A2(n13639), .ZN(n13726) );
  OR2_X1 U13743 ( .A1(n13639), .A2(n13640), .ZN(n13724) );
  AND2_X1 U13744 ( .A1(n13727), .A2(n13728), .ZN(n13640) );
  NAND3_X1 U13745 ( .A1(b_4_), .A2(n13729), .A3(a_13_), .ZN(n13728) );
  NAND2_X1 U13746 ( .A1(n13636), .A2(n13635), .ZN(n13729) );
  OR2_X1 U13747 ( .A1(n13635), .A2(n13636), .ZN(n13727) );
  AND2_X1 U13748 ( .A1(n13730), .A2(n13731), .ZN(n13636) );
  NAND2_X1 U13749 ( .A1(n13633), .A2(n13732), .ZN(n13731) );
  NAND2_X1 U13750 ( .A1(n13632), .A2(n13631), .ZN(n13732) );
  NOR2_X1 U13751 ( .A1(n7782), .A2(n13352), .ZN(n13633) );
  OR2_X1 U13752 ( .A1(n13631), .A2(n13632), .ZN(n13730) );
  AND2_X1 U13753 ( .A1(n13733), .A2(n13734), .ZN(n13632) );
  NAND2_X1 U13754 ( .A1(n13628), .A2(n13735), .ZN(n13734) );
  NAND2_X1 U13755 ( .A1(n13629), .A2(n13627), .ZN(n13735) );
  NOR2_X1 U13756 ( .A1(n7346), .A2(n13352), .ZN(n13628) );
  OR2_X1 U13757 ( .A1(n13627), .A2(n13629), .ZN(n13733) );
  AND2_X1 U13758 ( .A1(n13736), .A2(n13737), .ZN(n13629) );
  NAND2_X1 U13759 ( .A1(n13625), .A2(n13738), .ZN(n13737) );
  OR2_X1 U13760 ( .A1(n13623), .A2(n13624), .ZN(n13738) );
  NOR2_X1 U13761 ( .A1(n7773), .A2(n13352), .ZN(n13625) );
  NAND2_X1 U13762 ( .A1(n13623), .A2(n13624), .ZN(n13736) );
  NAND2_X1 U13763 ( .A1(n13739), .A2(n13740), .ZN(n13624) );
  NAND2_X1 U13764 ( .A1(n13620), .A2(n13741), .ZN(n13740) );
  NAND2_X1 U13765 ( .A1(n13621), .A2(n13619), .ZN(n13741) );
  NOR2_X1 U13766 ( .A1(n7337), .A2(n13352), .ZN(n13620) );
  OR2_X1 U13767 ( .A1(n13619), .A2(n13621), .ZN(n13739) );
  AND2_X1 U13768 ( .A1(n13742), .A2(n13743), .ZN(n13621) );
  NAND2_X1 U13769 ( .A1(n13617), .A2(n13744), .ZN(n13743) );
  OR2_X1 U13770 ( .A1(n13615), .A2(n13616), .ZN(n13744) );
  NOR2_X1 U13771 ( .A1(n7764), .A2(n13352), .ZN(n13617) );
  NAND2_X1 U13772 ( .A1(n13615), .A2(n13616), .ZN(n13742) );
  NAND2_X1 U13773 ( .A1(n13745), .A2(n13746), .ZN(n13616) );
  NAND2_X1 U13774 ( .A1(n13613), .A2(n13747), .ZN(n13746) );
  NAND2_X1 U13775 ( .A1(n13612), .A2(n13611), .ZN(n13747) );
  NOR2_X1 U13776 ( .A1(n7902), .A2(n13352), .ZN(n13613) );
  OR2_X1 U13777 ( .A1(n13611), .A2(n13612), .ZN(n13745) );
  AND2_X1 U13778 ( .A1(n13748), .A2(n13749), .ZN(n13612) );
  NAND2_X1 U13779 ( .A1(n13609), .A2(n13750), .ZN(n13749) );
  OR2_X1 U13780 ( .A1(n13607), .A2(n13608), .ZN(n13750) );
  NOR2_X1 U13781 ( .A1(n7987), .A2(n13352), .ZN(n13609) );
  NAND2_X1 U13782 ( .A1(n13607), .A2(n13608), .ZN(n13748) );
  NAND2_X1 U13783 ( .A1(n13751), .A2(n13752), .ZN(n13608) );
  NAND2_X1 U13784 ( .A1(n13604), .A2(n13753), .ZN(n13752) );
  NAND2_X1 U13785 ( .A1(n13605), .A2(n13603), .ZN(n13753) );
  NOR2_X1 U13786 ( .A1(n7909), .A2(n13352), .ZN(n13604) );
  OR2_X1 U13787 ( .A1(n13603), .A2(n13605), .ZN(n13751) );
  AND2_X1 U13788 ( .A1(n13754), .A2(n13755), .ZN(n13605) );
  NAND2_X1 U13789 ( .A1(n13601), .A2(n13756), .ZN(n13755) );
  OR2_X1 U13790 ( .A1(n13598), .A2(n13600), .ZN(n13756) );
  NOR2_X1 U13791 ( .A1(n13352), .A2(n7312), .ZN(n13601) );
  NAND2_X1 U13792 ( .A1(n13598), .A2(n13600), .ZN(n13754) );
  NAND2_X1 U13793 ( .A1(n13757), .A2(n13758), .ZN(n13600) );
  NAND2_X1 U13794 ( .A1(n13597), .A2(n13759), .ZN(n13758) );
  OR2_X1 U13795 ( .A1(n13595), .A2(n13596), .ZN(n13759) );
  NOR2_X1 U13796 ( .A1(n13352), .A2(n7916), .ZN(n13597) );
  NAND2_X1 U13797 ( .A1(n13595), .A2(n13596), .ZN(n13757) );
  NAND2_X1 U13798 ( .A1(n13760), .A2(n13761), .ZN(n13596) );
  NAND2_X1 U13799 ( .A1(n13593), .A2(n13762), .ZN(n13761) );
  OR2_X1 U13800 ( .A1(n13591), .A2(n13592), .ZN(n13762) );
  NOR2_X1 U13801 ( .A1(n7691), .A2(n13352), .ZN(n13593) );
  NAND2_X1 U13802 ( .A1(n13591), .A2(n13592), .ZN(n13760) );
  NAND2_X1 U13803 ( .A1(n13763), .A2(n13764), .ZN(n13592) );
  NAND2_X1 U13804 ( .A1(n13589), .A2(n13765), .ZN(n13764) );
  OR2_X1 U13805 ( .A1(n13587), .A2(n13588), .ZN(n13765) );
  NOR2_X1 U13806 ( .A1(n13352), .A2(n7923), .ZN(n13589) );
  NAND2_X1 U13807 ( .A1(n13587), .A2(n13588), .ZN(n13763) );
  NAND2_X1 U13808 ( .A1(n13551), .A2(n13766), .ZN(n13588) );
  NAND2_X1 U13809 ( .A1(n13550), .A2(n13552), .ZN(n13766) );
  NAND2_X1 U13810 ( .A1(n13767), .A2(n13768), .ZN(n13552) );
  NAND2_X1 U13811 ( .A1(b_4_), .A2(a_26_), .ZN(n13768) );
  INV_X1 U13812 ( .A(n13769), .ZN(n13767) );
  XNOR2_X1 U13813 ( .A(n13770), .B(n13771), .ZN(n13550) );
  NAND2_X1 U13814 ( .A1(n13772), .A2(n13773), .ZN(n13770) );
  NAND2_X1 U13815 ( .A1(a_26_), .A2(n13769), .ZN(n13551) );
  NAND2_X1 U13816 ( .A1(n13559), .A2(n13774), .ZN(n13769) );
  NAND2_X1 U13817 ( .A1(n13558), .A2(n13560), .ZN(n13774) );
  NAND2_X1 U13818 ( .A1(n13775), .A2(n13776), .ZN(n13560) );
  NAND2_X1 U13819 ( .A1(b_4_), .A2(a_27_), .ZN(n13776) );
  INV_X1 U13820 ( .A(n13777), .ZN(n13775) );
  XNOR2_X1 U13821 ( .A(n13778), .B(n13779), .ZN(n13558) );
  XOR2_X1 U13822 ( .A(n13780), .B(n13781), .Z(n13778) );
  NAND2_X1 U13823 ( .A1(b_3_), .A2(a_28_), .ZN(n13780) );
  NAND2_X1 U13824 ( .A1(a_27_), .A2(n13777), .ZN(n13559) );
  NAND2_X1 U13825 ( .A1(n13782), .A2(n13783), .ZN(n13777) );
  NAND3_X1 U13826 ( .A1(a_28_), .A2(n13784), .A3(b_4_), .ZN(n13783) );
  NAND2_X1 U13827 ( .A1(n13568), .A2(n13566), .ZN(n13784) );
  OR2_X1 U13828 ( .A1(n13566), .A2(n13568), .ZN(n13782) );
  AND2_X1 U13829 ( .A1(n13785), .A2(n13786), .ZN(n13568) );
  NAND2_X1 U13830 ( .A1(n13583), .A2(n13787), .ZN(n13786) );
  OR2_X1 U13831 ( .A1(n13584), .A2(n13585), .ZN(n13787) );
  NOR2_X1 U13832 ( .A1(n13352), .A2(n7946), .ZN(n13583) );
  NAND2_X1 U13833 ( .A1(n13585), .A2(n13584), .ZN(n13785) );
  NAND2_X1 U13834 ( .A1(n13788), .A2(n13789), .ZN(n13584) );
  NAND2_X1 U13835 ( .A1(b_2_), .A2(n13790), .ZN(n13789) );
  NAND2_X1 U13836 ( .A1(n7268), .A2(n13791), .ZN(n13790) );
  NAND2_X1 U13837 ( .A1(a_31_), .A2(n13581), .ZN(n13791) );
  NAND2_X1 U13838 ( .A1(b_3_), .A2(n13792), .ZN(n13788) );
  NAND2_X1 U13839 ( .A1(n7272), .A2(n13793), .ZN(n13792) );
  NAND2_X1 U13840 ( .A1(a_30_), .A2(n13794), .ZN(n13793) );
  AND3_X1 U13841 ( .A1(b_4_), .A2(n7954), .A3(b_3_), .ZN(n13585) );
  XNOR2_X1 U13842 ( .A(n13795), .B(n13796), .ZN(n13566) );
  XOR2_X1 U13843 ( .A(n13797), .B(n13798), .Z(n13795) );
  XNOR2_X1 U13844 ( .A(n13799), .B(n13800), .ZN(n13587) );
  NAND2_X1 U13845 ( .A1(n13801), .A2(n13802), .ZN(n13799) );
  XNOR2_X1 U13846 ( .A(n13803), .B(n13804), .ZN(n13591) );
  NAND2_X1 U13847 ( .A1(n13805), .A2(n13806), .ZN(n13803) );
  XNOR2_X1 U13848 ( .A(n13807), .B(n13808), .ZN(n13595) );
  XNOR2_X1 U13849 ( .A(n13809), .B(n13810), .ZN(n13807) );
  NOR2_X1 U13850 ( .A1(n13581), .A2(n7691), .ZN(n13810) );
  XNOR2_X1 U13851 ( .A(n13811), .B(n13812), .ZN(n13598) );
  NAND2_X1 U13852 ( .A1(n13813), .A2(n13814), .ZN(n13811) );
  XNOR2_X1 U13853 ( .A(n13815), .B(n13816), .ZN(n13603) );
  XNOR2_X1 U13854 ( .A(n13817), .B(n13818), .ZN(n13815) );
  NAND2_X1 U13855 ( .A1(b_3_), .A2(a_22_), .ZN(n13817) );
  XNOR2_X1 U13856 ( .A(n13819), .B(n13820), .ZN(n13607) );
  NAND2_X1 U13857 ( .A1(n13821), .A2(n13822), .ZN(n13819) );
  XNOR2_X1 U13858 ( .A(n13823), .B(n13824), .ZN(n13611) );
  XNOR2_X1 U13859 ( .A(n13825), .B(n13826), .ZN(n13823) );
  NAND2_X1 U13860 ( .A1(a_20_), .A2(b_3_), .ZN(n13825) );
  XNOR2_X1 U13861 ( .A(n13827), .B(n13828), .ZN(n13615) );
  NAND2_X1 U13862 ( .A1(n13829), .A2(n13830), .ZN(n13827) );
  XNOR2_X1 U13863 ( .A(n13831), .B(n13832), .ZN(n13619) );
  XNOR2_X1 U13864 ( .A(n13833), .B(n13834), .ZN(n13831) );
  NAND2_X1 U13865 ( .A1(a_18_), .A2(b_3_), .ZN(n13833) );
  XNOR2_X1 U13866 ( .A(n13835), .B(n13836), .ZN(n13623) );
  NAND2_X1 U13867 ( .A1(n13837), .A2(n13838), .ZN(n13835) );
  XNOR2_X1 U13868 ( .A(n13839), .B(n13840), .ZN(n13627) );
  XNOR2_X1 U13869 ( .A(n13841), .B(n13842), .ZN(n13839) );
  NAND2_X1 U13870 ( .A1(a_16_), .A2(b_3_), .ZN(n13841) );
  XOR2_X1 U13871 ( .A(n13843), .B(n13844), .Z(n13631) );
  NAND2_X1 U13872 ( .A1(n13845), .A2(n13846), .ZN(n13843) );
  XNOR2_X1 U13873 ( .A(n13847), .B(n13848), .ZN(n13635) );
  XNOR2_X1 U13874 ( .A(n13849), .B(n13850), .ZN(n13847) );
  NAND2_X1 U13875 ( .A1(a_14_), .A2(b_3_), .ZN(n13849) );
  XOR2_X1 U13876 ( .A(n13851), .B(n13852), .Z(n13639) );
  NAND2_X1 U13877 ( .A1(n13853), .A2(n13854), .ZN(n13851) );
  XNOR2_X1 U13878 ( .A(n13855), .B(n13856), .ZN(n13642) );
  XNOR2_X1 U13879 ( .A(n13857), .B(n13858), .ZN(n13855) );
  NAND2_X1 U13880 ( .A1(a_12_), .A2(b_3_), .ZN(n13857) );
  XOR2_X1 U13881 ( .A(n13859), .B(n13860), .Z(n13646) );
  NAND2_X1 U13882 ( .A1(n13861), .A2(n13862), .ZN(n13859) );
  XNOR2_X1 U13883 ( .A(n13863), .B(n13864), .ZN(n13650) );
  XNOR2_X1 U13884 ( .A(n13865), .B(n13866), .ZN(n13863) );
  NAND2_X1 U13885 ( .A1(a_10_), .A2(b_3_), .ZN(n13865) );
  XOR2_X1 U13886 ( .A(n13867), .B(n13868), .Z(n13654) );
  NAND2_X1 U13887 ( .A1(n13869), .A2(n13870), .ZN(n13867) );
  XOR2_X1 U13888 ( .A(n13871), .B(n13872), .Z(n13659) );
  XNOR2_X1 U13889 ( .A(n13873), .B(n13874), .ZN(n13871) );
  NAND2_X1 U13890 ( .A1(a_8_), .A2(b_3_), .ZN(n13873) );
  XOR2_X1 U13891 ( .A(n13875), .B(n13876), .Z(n13485) );
  NAND2_X1 U13892 ( .A1(n13877), .A2(n13878), .ZN(n13875) );
  XOR2_X1 U13893 ( .A(n13879), .B(n13880), .Z(n13663) );
  XNOR2_X1 U13894 ( .A(n13881), .B(n13882), .ZN(n13879) );
  NAND2_X1 U13895 ( .A1(a_6_), .A2(b_3_), .ZN(n13881) );
  XNOR2_X1 U13896 ( .A(n13883), .B(n13884), .ZN(n13667) );
  NAND2_X1 U13897 ( .A1(n13885), .A2(n13886), .ZN(n13883) );
  XOR2_X1 U13898 ( .A(n13887), .B(n13888), .Z(n13671) );
  XNOR2_X1 U13899 ( .A(n13889), .B(n13890), .ZN(n13887) );
  NAND2_X1 U13900 ( .A1(a_4_), .A2(b_3_), .ZN(n13889) );
  XOR2_X1 U13901 ( .A(n13891), .B(n13892), .Z(n13675) );
  XOR2_X1 U13902 ( .A(n13893), .B(n13894), .Z(n13891) );
  XOR2_X1 U13903 ( .A(n13895), .B(n13896), .Z(n13679) );
  XNOR2_X1 U13904 ( .A(n13897), .B(n13898), .ZN(n13895) );
  NAND2_X1 U13905 ( .A1(a_2_), .A2(b_3_), .ZN(n13897) );
  XNOR2_X1 U13906 ( .A(n13899), .B(n13900), .ZN(n13457) );
  NAND2_X1 U13907 ( .A1(n13901), .A2(n13902), .ZN(n13899) );
  NAND2_X1 U13908 ( .A1(n13903), .A2(n13904), .ZN(n13686) );
  XOR2_X1 U13909 ( .A(n13905), .B(n13906), .Z(n13465) );
  XOR2_X1 U13910 ( .A(n13907), .B(n13908), .Z(n13905) );
  NAND2_X1 U13911 ( .A1(n13909), .A2(n13687), .ZN(n7424) );
  INV_X1 U13912 ( .A(n13910), .ZN(n13687) );
  XOR2_X1 U13913 ( .A(n7513), .B(n13911), .Z(n13909) );
  NAND2_X1 U13914 ( .A1(n13910), .A2(n13912), .ZN(n7425) );
  XOR2_X1 U13915 ( .A(n7514), .B(n7513), .Z(n13912) );
  NOR2_X1 U13916 ( .A1(n13904), .A2(n13903), .ZN(n13910) );
  AND2_X1 U13917 ( .A1(n13913), .A2(n13914), .ZN(n13903) );
  NAND2_X1 U13918 ( .A1(n13907), .A2(n13915), .ZN(n13914) );
  OR2_X1 U13919 ( .A1(n13906), .A2(n13908), .ZN(n13915) );
  NOR2_X1 U13920 ( .A1(n13581), .A2(n7613), .ZN(n13907) );
  NAND2_X1 U13921 ( .A1(n13906), .A2(n13908), .ZN(n13913) );
  NAND2_X1 U13922 ( .A1(n13901), .A2(n13916), .ZN(n13908) );
  NAND2_X1 U13923 ( .A1(n13900), .A2(n13902), .ZN(n13916) );
  NAND2_X1 U13924 ( .A1(n13917), .A2(n13918), .ZN(n13902) );
  NAND2_X1 U13925 ( .A1(a_1_), .A2(b_3_), .ZN(n13918) );
  INV_X1 U13926 ( .A(n13919), .ZN(n13917) );
  XNOR2_X1 U13927 ( .A(n13920), .B(n13921), .ZN(n13900) );
  XNOR2_X1 U13928 ( .A(n13922), .B(n13923), .ZN(n13921) );
  NAND2_X1 U13929 ( .A1(a_1_), .A2(n13919), .ZN(n13901) );
  NAND2_X1 U13930 ( .A1(n13924), .A2(n13925), .ZN(n13919) );
  NAND3_X1 U13931 ( .A1(b_3_), .A2(n13926), .A3(a_2_), .ZN(n13925) );
  OR2_X1 U13932 ( .A1(n13896), .A2(n13898), .ZN(n13926) );
  NAND2_X1 U13933 ( .A1(n13896), .A2(n13898), .ZN(n13924) );
  NAND2_X1 U13934 ( .A1(n13927), .A2(n13928), .ZN(n13898) );
  NAND2_X1 U13935 ( .A1(n13892), .A2(n13929), .ZN(n13928) );
  OR2_X1 U13936 ( .A1(n13893), .A2(n13894), .ZN(n13929) );
  XNOR2_X1 U13937 ( .A(n13930), .B(n13931), .ZN(n13892) );
  NAND2_X1 U13938 ( .A1(n13932), .A2(n13933), .ZN(n13930) );
  NAND2_X1 U13939 ( .A1(n13894), .A2(n13893), .ZN(n13927) );
  NAND2_X1 U13940 ( .A1(n13934), .A2(n13935), .ZN(n13893) );
  NAND3_X1 U13941 ( .A1(b_3_), .A2(n13936), .A3(a_4_), .ZN(n13935) );
  OR2_X1 U13942 ( .A1(n13888), .A2(n13890), .ZN(n13936) );
  NAND2_X1 U13943 ( .A1(n13888), .A2(n13890), .ZN(n13934) );
  NAND2_X1 U13944 ( .A1(n13885), .A2(n13937), .ZN(n13890) );
  NAND2_X1 U13945 ( .A1(n13884), .A2(n13886), .ZN(n13937) );
  NAND2_X1 U13946 ( .A1(n13938), .A2(n13939), .ZN(n13886) );
  NAND2_X1 U13947 ( .A1(a_5_), .A2(b_3_), .ZN(n13939) );
  INV_X1 U13948 ( .A(n13940), .ZN(n13938) );
  XNOR2_X1 U13949 ( .A(n13941), .B(n13942), .ZN(n13884) );
  NAND2_X1 U13950 ( .A1(n13943), .A2(n13944), .ZN(n13941) );
  NAND2_X1 U13951 ( .A1(a_5_), .A2(n13940), .ZN(n13885) );
  NAND2_X1 U13952 ( .A1(n13945), .A2(n13946), .ZN(n13940) );
  NAND3_X1 U13953 ( .A1(b_3_), .A2(n13947), .A3(a_6_), .ZN(n13946) );
  OR2_X1 U13954 ( .A1(n13880), .A2(n13882), .ZN(n13947) );
  NAND2_X1 U13955 ( .A1(n13880), .A2(n13882), .ZN(n13945) );
  NAND2_X1 U13956 ( .A1(n13877), .A2(n13948), .ZN(n13882) );
  NAND2_X1 U13957 ( .A1(n13876), .A2(n13878), .ZN(n13948) );
  NAND2_X1 U13958 ( .A1(n13949), .A2(n13950), .ZN(n13878) );
  NAND2_X1 U13959 ( .A1(a_7_), .A2(b_3_), .ZN(n13950) );
  INV_X1 U13960 ( .A(n13951), .ZN(n13949) );
  XNOR2_X1 U13961 ( .A(n13952), .B(n13953), .ZN(n13876) );
  NAND2_X1 U13962 ( .A1(n13954), .A2(n13955), .ZN(n13952) );
  NAND2_X1 U13963 ( .A1(a_7_), .A2(n13951), .ZN(n13877) );
  NAND2_X1 U13964 ( .A1(n13956), .A2(n13957), .ZN(n13951) );
  NAND3_X1 U13965 ( .A1(b_3_), .A2(n13958), .A3(a_8_), .ZN(n13957) );
  OR2_X1 U13966 ( .A1(n13872), .A2(n13874), .ZN(n13958) );
  NAND2_X1 U13967 ( .A1(n13872), .A2(n13874), .ZN(n13956) );
  NAND2_X1 U13968 ( .A1(n13869), .A2(n13959), .ZN(n13874) );
  NAND2_X1 U13969 ( .A1(n13868), .A2(n13870), .ZN(n13959) );
  NAND2_X1 U13970 ( .A1(n13960), .A2(n13961), .ZN(n13870) );
  NAND2_X1 U13971 ( .A1(b_3_), .A2(a_9_), .ZN(n13961) );
  INV_X1 U13972 ( .A(n13962), .ZN(n13960) );
  XNOR2_X1 U13973 ( .A(n13963), .B(n13964), .ZN(n13868) );
  NAND2_X1 U13974 ( .A1(n13965), .A2(n13966), .ZN(n13963) );
  NAND2_X1 U13975 ( .A1(a_9_), .A2(n13962), .ZN(n13869) );
  NAND2_X1 U13976 ( .A1(n13967), .A2(n13968), .ZN(n13962) );
  NAND3_X1 U13977 ( .A1(b_3_), .A2(n13969), .A3(a_10_), .ZN(n13968) );
  OR2_X1 U13978 ( .A1(n13864), .A2(n13866), .ZN(n13969) );
  NAND2_X1 U13979 ( .A1(n13864), .A2(n13866), .ZN(n13967) );
  NAND2_X1 U13980 ( .A1(n13861), .A2(n13970), .ZN(n13866) );
  NAND2_X1 U13981 ( .A1(n13860), .A2(n13862), .ZN(n13970) );
  NAND2_X1 U13982 ( .A1(n13971), .A2(n13972), .ZN(n13862) );
  NAND2_X1 U13983 ( .A1(a_11_), .A2(b_3_), .ZN(n13972) );
  INV_X1 U13984 ( .A(n13973), .ZN(n13971) );
  XNOR2_X1 U13985 ( .A(n13974), .B(n13975), .ZN(n13860) );
  NAND2_X1 U13986 ( .A1(n13976), .A2(n13977), .ZN(n13974) );
  NAND2_X1 U13987 ( .A1(a_11_), .A2(n13973), .ZN(n13861) );
  NAND2_X1 U13988 ( .A1(n13978), .A2(n13979), .ZN(n13973) );
  NAND3_X1 U13989 ( .A1(b_3_), .A2(n13980), .A3(a_12_), .ZN(n13979) );
  OR2_X1 U13990 ( .A1(n13856), .A2(n13858), .ZN(n13980) );
  NAND2_X1 U13991 ( .A1(n13856), .A2(n13858), .ZN(n13978) );
  NAND2_X1 U13992 ( .A1(n13853), .A2(n13981), .ZN(n13858) );
  NAND2_X1 U13993 ( .A1(n13852), .A2(n13854), .ZN(n13981) );
  NAND2_X1 U13994 ( .A1(n13982), .A2(n13983), .ZN(n13854) );
  NAND2_X1 U13995 ( .A1(a_13_), .A2(b_3_), .ZN(n13983) );
  INV_X1 U13996 ( .A(n13984), .ZN(n13982) );
  XNOR2_X1 U13997 ( .A(n13985), .B(n13986), .ZN(n13852) );
  NAND2_X1 U13998 ( .A1(n13987), .A2(n13988), .ZN(n13985) );
  NAND2_X1 U13999 ( .A1(a_13_), .A2(n13984), .ZN(n13853) );
  NAND2_X1 U14000 ( .A1(n13989), .A2(n13990), .ZN(n13984) );
  NAND3_X1 U14001 ( .A1(b_3_), .A2(n13991), .A3(a_14_), .ZN(n13990) );
  OR2_X1 U14002 ( .A1(n13848), .A2(n13850), .ZN(n13991) );
  NAND2_X1 U14003 ( .A1(n13848), .A2(n13850), .ZN(n13989) );
  NAND2_X1 U14004 ( .A1(n13845), .A2(n13992), .ZN(n13850) );
  NAND2_X1 U14005 ( .A1(n13844), .A2(n13846), .ZN(n13992) );
  NAND2_X1 U14006 ( .A1(n13993), .A2(n13994), .ZN(n13846) );
  NAND2_X1 U14007 ( .A1(a_15_), .A2(b_3_), .ZN(n13994) );
  INV_X1 U14008 ( .A(n13995), .ZN(n13993) );
  XNOR2_X1 U14009 ( .A(n13996), .B(n13997), .ZN(n13844) );
  NAND2_X1 U14010 ( .A1(n13998), .A2(n13999), .ZN(n13996) );
  NAND2_X1 U14011 ( .A1(a_15_), .A2(n13995), .ZN(n13845) );
  NAND2_X1 U14012 ( .A1(n14000), .A2(n14001), .ZN(n13995) );
  NAND3_X1 U14013 ( .A1(b_3_), .A2(n14002), .A3(a_16_), .ZN(n14001) );
  OR2_X1 U14014 ( .A1(n13840), .A2(n13842), .ZN(n14002) );
  NAND2_X1 U14015 ( .A1(n13840), .A2(n13842), .ZN(n14000) );
  NAND2_X1 U14016 ( .A1(n13837), .A2(n14003), .ZN(n13842) );
  NAND2_X1 U14017 ( .A1(n13836), .A2(n13838), .ZN(n14003) );
  NAND2_X1 U14018 ( .A1(n14004), .A2(n14005), .ZN(n13838) );
  NAND2_X1 U14019 ( .A1(a_17_), .A2(b_3_), .ZN(n14005) );
  INV_X1 U14020 ( .A(n14006), .ZN(n14004) );
  XNOR2_X1 U14021 ( .A(n14007), .B(n14008), .ZN(n13836) );
  XNOR2_X1 U14022 ( .A(n14009), .B(n14010), .ZN(n14008) );
  NAND2_X1 U14023 ( .A1(a_17_), .A2(n14006), .ZN(n13837) );
  NAND2_X1 U14024 ( .A1(n14011), .A2(n14012), .ZN(n14006) );
  NAND3_X1 U14025 ( .A1(b_3_), .A2(n14013), .A3(a_18_), .ZN(n14012) );
  OR2_X1 U14026 ( .A1(n13832), .A2(n13834), .ZN(n14013) );
  NAND2_X1 U14027 ( .A1(n13832), .A2(n13834), .ZN(n14011) );
  NAND2_X1 U14028 ( .A1(n13829), .A2(n14014), .ZN(n13834) );
  NAND2_X1 U14029 ( .A1(n13828), .A2(n13830), .ZN(n14014) );
  NAND2_X1 U14030 ( .A1(n14015), .A2(n14016), .ZN(n13830) );
  NAND2_X1 U14031 ( .A1(a_19_), .A2(b_3_), .ZN(n14016) );
  INV_X1 U14032 ( .A(n14017), .ZN(n14015) );
  XNOR2_X1 U14033 ( .A(n14018), .B(n14019), .ZN(n13828) );
  XNOR2_X1 U14034 ( .A(n14020), .B(n14021), .ZN(n14019) );
  NAND2_X1 U14035 ( .A1(a_19_), .A2(n14017), .ZN(n13829) );
  NAND2_X1 U14036 ( .A1(n14022), .A2(n14023), .ZN(n14017) );
  NAND3_X1 U14037 ( .A1(b_3_), .A2(n14024), .A3(a_20_), .ZN(n14023) );
  OR2_X1 U14038 ( .A1(n13824), .A2(n13826), .ZN(n14024) );
  NAND2_X1 U14039 ( .A1(n13824), .A2(n13826), .ZN(n14022) );
  NAND2_X1 U14040 ( .A1(n13821), .A2(n14025), .ZN(n13826) );
  NAND2_X1 U14041 ( .A1(n13820), .A2(n13822), .ZN(n14025) );
  NAND2_X1 U14042 ( .A1(n14026), .A2(n14027), .ZN(n13822) );
  NAND2_X1 U14043 ( .A1(a_21_), .A2(b_3_), .ZN(n14027) );
  INV_X1 U14044 ( .A(n14028), .ZN(n14026) );
  XNOR2_X1 U14045 ( .A(n14029), .B(n14030), .ZN(n13820) );
  XNOR2_X1 U14046 ( .A(n14031), .B(n14032), .ZN(n14030) );
  NAND2_X1 U14047 ( .A1(a_21_), .A2(n14028), .ZN(n13821) );
  NAND2_X1 U14048 ( .A1(n14033), .A2(n14034), .ZN(n14028) );
  NAND3_X1 U14049 ( .A1(a_22_), .A2(n14035), .A3(b_3_), .ZN(n14034) );
  OR2_X1 U14050 ( .A1(n13816), .A2(n13818), .ZN(n14035) );
  NAND2_X1 U14051 ( .A1(n13816), .A2(n13818), .ZN(n14033) );
  NAND2_X1 U14052 ( .A1(n13813), .A2(n14036), .ZN(n13818) );
  NAND2_X1 U14053 ( .A1(n13812), .A2(n13814), .ZN(n14036) );
  NAND2_X1 U14054 ( .A1(n14037), .A2(n14038), .ZN(n13814) );
  NAND2_X1 U14055 ( .A1(b_3_), .A2(a_23_), .ZN(n14038) );
  INV_X1 U14056 ( .A(n14039), .ZN(n14037) );
  XNOR2_X1 U14057 ( .A(n14040), .B(n14041), .ZN(n13812) );
  XNOR2_X1 U14058 ( .A(n14042), .B(n14043), .ZN(n14041) );
  NAND2_X1 U14059 ( .A1(a_23_), .A2(n14039), .ZN(n13813) );
  NAND2_X1 U14060 ( .A1(n14044), .A2(n14045), .ZN(n14039) );
  NAND3_X1 U14061 ( .A1(b_3_), .A2(n14046), .A3(a_24_), .ZN(n14045) );
  NAND2_X1 U14062 ( .A1(n13809), .A2(n13808), .ZN(n14046) );
  OR2_X1 U14063 ( .A1(n13808), .A2(n13809), .ZN(n14044) );
  AND2_X1 U14064 ( .A1(n13805), .A2(n14047), .ZN(n13809) );
  NAND2_X1 U14065 ( .A1(n13804), .A2(n13806), .ZN(n14047) );
  NAND2_X1 U14066 ( .A1(n14048), .A2(n14049), .ZN(n13806) );
  NAND2_X1 U14067 ( .A1(b_3_), .A2(a_25_), .ZN(n14049) );
  INV_X1 U14068 ( .A(n14050), .ZN(n14048) );
  XNOR2_X1 U14069 ( .A(n14051), .B(n14052), .ZN(n13804) );
  XOR2_X1 U14070 ( .A(n14053), .B(n14054), .Z(n14051) );
  NAND2_X1 U14071 ( .A1(b_2_), .A2(a_26_), .ZN(n14053) );
  NAND2_X1 U14072 ( .A1(a_25_), .A2(n14050), .ZN(n13805) );
  NAND2_X1 U14073 ( .A1(n13801), .A2(n14055), .ZN(n14050) );
  NAND2_X1 U14074 ( .A1(n13800), .A2(n13802), .ZN(n14055) );
  NAND2_X1 U14075 ( .A1(n14056), .A2(n14057), .ZN(n13802) );
  NAND2_X1 U14076 ( .A1(b_3_), .A2(a_26_), .ZN(n14057) );
  INV_X1 U14077 ( .A(n14058), .ZN(n14056) );
  XNOR2_X1 U14078 ( .A(n14059), .B(n14060), .ZN(n13800) );
  XNOR2_X1 U14079 ( .A(n14061), .B(n14062), .ZN(n14060) );
  NAND2_X1 U14080 ( .A1(a_26_), .A2(n14058), .ZN(n13801) );
  NAND2_X1 U14081 ( .A1(n13772), .A2(n14063), .ZN(n14058) );
  NAND2_X1 U14082 ( .A1(n13771), .A2(n13773), .ZN(n14063) );
  NAND2_X1 U14083 ( .A1(n14064), .A2(n14065), .ZN(n13773) );
  NAND2_X1 U14084 ( .A1(b_3_), .A2(a_27_), .ZN(n14065) );
  INV_X1 U14085 ( .A(n14066), .ZN(n14064) );
  XOR2_X1 U14086 ( .A(n14067), .B(n14068), .Z(n13771) );
  XNOR2_X1 U14087 ( .A(n14069), .B(n14070), .ZN(n14067) );
  NAND2_X1 U14088 ( .A1(b_2_), .A2(a_28_), .ZN(n14069) );
  NAND2_X1 U14089 ( .A1(a_27_), .A2(n14066), .ZN(n13772) );
  NAND2_X1 U14090 ( .A1(n14071), .A2(n14072), .ZN(n14066) );
  NAND3_X1 U14091 ( .A1(a_28_), .A2(n14073), .A3(b_3_), .ZN(n14072) );
  NAND2_X1 U14092 ( .A1(n13781), .A2(n13779), .ZN(n14073) );
  OR2_X1 U14093 ( .A1(n13779), .A2(n13781), .ZN(n14071) );
  AND2_X1 U14094 ( .A1(n14074), .A2(n14075), .ZN(n13781) );
  NAND2_X1 U14095 ( .A1(n13796), .A2(n14076), .ZN(n14075) );
  OR2_X1 U14096 ( .A1(n13797), .A2(n13798), .ZN(n14076) );
  NOR2_X1 U14097 ( .A1(n13581), .A2(n7946), .ZN(n13796) );
  NAND2_X1 U14098 ( .A1(n13798), .A2(n13797), .ZN(n14074) );
  NAND2_X1 U14099 ( .A1(n14077), .A2(n14078), .ZN(n13797) );
  NAND2_X1 U14100 ( .A1(b_1_), .A2(n14079), .ZN(n14078) );
  NAND2_X1 U14101 ( .A1(n7268), .A2(n14080), .ZN(n14079) );
  NAND2_X1 U14102 ( .A1(a_31_), .A2(n13794), .ZN(n14080) );
  NAND2_X1 U14103 ( .A1(b_2_), .A2(n14081), .ZN(n14077) );
  NAND2_X1 U14104 ( .A1(n7272), .A2(n14082), .ZN(n14081) );
  NAND2_X1 U14105 ( .A1(a_30_), .A2(n14083), .ZN(n14082) );
  AND3_X1 U14106 ( .A1(b_3_), .A2(n7954), .A3(b_2_), .ZN(n13798) );
  XNOR2_X1 U14107 ( .A(n14084), .B(n14085), .ZN(n13779) );
  NOR2_X1 U14108 ( .A1(n7946), .A2(n13794), .ZN(n14085) );
  XOR2_X1 U14109 ( .A(n14086), .B(n14087), .Z(n14084) );
  XOR2_X1 U14110 ( .A(n14088), .B(n14089), .Z(n13808) );
  NAND2_X1 U14111 ( .A1(n14090), .A2(n14091), .ZN(n14088) );
  XNOR2_X1 U14112 ( .A(n14092), .B(n14093), .ZN(n13816) );
  XOR2_X1 U14113 ( .A(n14094), .B(n14095), .Z(n14093) );
  NAND2_X1 U14114 ( .A1(b_2_), .A2(a_23_), .ZN(n14095) );
  XNOR2_X1 U14115 ( .A(n14096), .B(n14097), .ZN(n13824) );
  XOR2_X1 U14116 ( .A(n14098), .B(n14099), .Z(n14096) );
  NAND2_X1 U14117 ( .A1(a_21_), .A2(b_2_), .ZN(n14098) );
  XNOR2_X1 U14118 ( .A(n14100), .B(n14101), .ZN(n13832) );
  XOR2_X1 U14119 ( .A(n14102), .B(n14103), .Z(n14100) );
  NAND2_X1 U14120 ( .A1(a_19_), .A2(b_2_), .ZN(n14102) );
  XNOR2_X1 U14121 ( .A(n14104), .B(n14105), .ZN(n13840) );
  XNOR2_X1 U14122 ( .A(n14106), .B(n14107), .ZN(n14104) );
  XOR2_X1 U14123 ( .A(n14108), .B(n14109), .Z(n13848) );
  XOR2_X1 U14124 ( .A(n14110), .B(n14111), .Z(n14108) );
  XOR2_X1 U14125 ( .A(n14112), .B(n14113), .Z(n13856) );
  XOR2_X1 U14126 ( .A(n14114), .B(n14115), .Z(n14112) );
  XOR2_X1 U14127 ( .A(n14116), .B(n14117), .Z(n13864) );
  XOR2_X1 U14128 ( .A(n14118), .B(n14119), .Z(n14116) );
  XOR2_X1 U14129 ( .A(n14120), .B(n14121), .Z(n13872) );
  XOR2_X1 U14130 ( .A(n14122), .B(n14123), .Z(n14120) );
  XOR2_X1 U14131 ( .A(n14124), .B(n14125), .Z(n13880) );
  XOR2_X1 U14132 ( .A(n14126), .B(n14127), .Z(n14124) );
  XOR2_X1 U14133 ( .A(n14128), .B(n14129), .Z(n13888) );
  XOR2_X1 U14134 ( .A(n14130), .B(n14131), .Z(n14128) );
  XOR2_X1 U14135 ( .A(n14132), .B(n14133), .Z(n13896) );
  XOR2_X1 U14136 ( .A(n14134), .B(n14135), .Z(n14132) );
  XOR2_X1 U14137 ( .A(n14136), .B(n14137), .Z(n13906) );
  XOR2_X1 U14138 ( .A(n14138), .B(n14139), .Z(n14136) );
  XOR2_X1 U14139 ( .A(n14140), .B(n14141), .Z(n13904) );
  NAND2_X1 U14140 ( .A1(n14142), .A2(n14143), .ZN(n14140) );
  NAND2_X1 U14141 ( .A1(n14144), .A2(n14145), .ZN(n7467) );
  OR2_X1 U14142 ( .A1(n7513), .A2(n7514), .ZN(n14145) );
  INV_X1 U14143 ( .A(n13911), .ZN(n7514) );
  NAND2_X1 U14144 ( .A1(n14142), .A2(n14146), .ZN(n13911) );
  NAND2_X1 U14145 ( .A1(n14141), .A2(n14143), .ZN(n14146) );
  NAND2_X1 U14146 ( .A1(n14147), .A2(n14148), .ZN(n14143) );
  NAND2_X1 U14147 ( .A1(b_2_), .A2(a_0_), .ZN(n14148) );
  INV_X1 U14148 ( .A(n14149), .ZN(n14147) );
  XNOR2_X1 U14149 ( .A(n14150), .B(n14151), .ZN(n14141) );
  XNOR2_X1 U14150 ( .A(n14152), .B(n14153), .ZN(n14151) );
  NAND2_X1 U14151 ( .A1(a_0_), .A2(n14149), .ZN(n14142) );
  NAND2_X1 U14152 ( .A1(n14154), .A2(n14155), .ZN(n14149) );
  NAND2_X1 U14153 ( .A1(n14138), .A2(n14156), .ZN(n14155) );
  OR2_X1 U14154 ( .A1(n14139), .A2(n14137), .ZN(n14156) );
  NOR2_X1 U14155 ( .A1(n7411), .A2(n13794), .ZN(n14138) );
  NAND2_X1 U14156 ( .A1(n14137), .A2(n14139), .ZN(n14154) );
  NAND2_X1 U14157 ( .A1(n14157), .A2(n14158), .ZN(n14139) );
  NAND2_X1 U14158 ( .A1(n13922), .A2(n14159), .ZN(n14158) );
  OR2_X1 U14159 ( .A1(n13923), .A2(n13920), .ZN(n14159) );
  NAND2_X1 U14160 ( .A1(n13920), .A2(n13923), .ZN(n14157) );
  NAND2_X1 U14161 ( .A1(n14160), .A2(n14161), .ZN(n13923) );
  NAND2_X1 U14162 ( .A1(n14134), .A2(n14162), .ZN(n14161) );
  OR2_X1 U14163 ( .A1(n14135), .A2(n14133), .ZN(n14162) );
  NOR2_X1 U14164 ( .A1(n7850), .A2(n13794), .ZN(n14134) );
  NAND2_X1 U14165 ( .A1(n14133), .A2(n14135), .ZN(n14160) );
  NAND2_X1 U14166 ( .A1(n13932), .A2(n14163), .ZN(n14135) );
  NAND2_X1 U14167 ( .A1(n13931), .A2(n13933), .ZN(n14163) );
  NAND2_X1 U14168 ( .A1(n14164), .A2(n14165), .ZN(n13933) );
  NAND2_X1 U14169 ( .A1(a_4_), .A2(b_2_), .ZN(n14165) );
  INV_X1 U14170 ( .A(n14166), .ZN(n14164) );
  XOR2_X1 U14171 ( .A(n14167), .B(n14168), .Z(n13931) );
  XNOR2_X1 U14172 ( .A(n14169), .B(n14170), .ZN(n14168) );
  NAND2_X1 U14173 ( .A1(a_5_), .A2(b_1_), .ZN(n14167) );
  NAND2_X1 U14174 ( .A1(a_4_), .A2(n14166), .ZN(n13932) );
  NAND2_X1 U14175 ( .A1(n14171), .A2(n14172), .ZN(n14166) );
  NAND2_X1 U14176 ( .A1(n14130), .A2(n14173), .ZN(n14172) );
  OR2_X1 U14177 ( .A1(n14131), .A2(n14129), .ZN(n14173) );
  NOR2_X1 U14178 ( .A1(n7393), .A2(n13794), .ZN(n14130) );
  NAND2_X1 U14179 ( .A1(n14129), .A2(n14131), .ZN(n14171) );
  NAND2_X1 U14180 ( .A1(n13943), .A2(n14174), .ZN(n14131) );
  NAND2_X1 U14181 ( .A1(n13942), .A2(n13944), .ZN(n14174) );
  NAND2_X1 U14182 ( .A1(n14175), .A2(n14176), .ZN(n13944) );
  NAND2_X1 U14183 ( .A1(a_6_), .A2(b_2_), .ZN(n14176) );
  INV_X1 U14184 ( .A(n14177), .ZN(n14175) );
  XOR2_X1 U14185 ( .A(n14178), .B(n14179), .Z(n13942) );
  XNOR2_X1 U14186 ( .A(n14180), .B(n14181), .ZN(n14179) );
  NAND2_X1 U14187 ( .A1(a_7_), .A2(b_1_), .ZN(n14178) );
  NAND2_X1 U14188 ( .A1(a_6_), .A2(n14177), .ZN(n13943) );
  NAND2_X1 U14189 ( .A1(n14182), .A2(n14183), .ZN(n14177) );
  NAND2_X1 U14190 ( .A1(n14126), .A2(n14184), .ZN(n14183) );
  OR2_X1 U14191 ( .A1(n14127), .A2(n14125), .ZN(n14184) );
  NOR2_X1 U14192 ( .A1(n7863), .A2(n13794), .ZN(n14126) );
  NAND2_X1 U14193 ( .A1(n14125), .A2(n14127), .ZN(n14182) );
  NAND2_X1 U14194 ( .A1(n13954), .A2(n14185), .ZN(n14127) );
  NAND2_X1 U14195 ( .A1(n13953), .A2(n13955), .ZN(n14185) );
  NAND2_X1 U14196 ( .A1(n14186), .A2(n14187), .ZN(n13955) );
  NAND2_X1 U14197 ( .A1(a_8_), .A2(b_2_), .ZN(n14187) );
  INV_X1 U14198 ( .A(n14188), .ZN(n14186) );
  XOR2_X1 U14199 ( .A(n14189), .B(n14190), .Z(n13953) );
  XNOR2_X1 U14200 ( .A(n14191), .B(n14192), .ZN(n14190) );
  NAND2_X1 U14201 ( .A1(b_1_), .A2(a_9_), .ZN(n14189) );
  NAND2_X1 U14202 ( .A1(a_8_), .A2(n14188), .ZN(n13954) );
  NAND2_X1 U14203 ( .A1(n14193), .A2(n14194), .ZN(n14188) );
  NAND2_X1 U14204 ( .A1(n14122), .A2(n14195), .ZN(n14194) );
  OR2_X1 U14205 ( .A1(n14123), .A2(n14121), .ZN(n14195) );
  NOR2_X1 U14206 ( .A1(n13794), .A2(n7870), .ZN(n14122) );
  NAND2_X1 U14207 ( .A1(n14121), .A2(n14123), .ZN(n14193) );
  NAND2_X1 U14208 ( .A1(n13965), .A2(n14196), .ZN(n14123) );
  NAND2_X1 U14209 ( .A1(n13964), .A2(n13966), .ZN(n14196) );
  NAND2_X1 U14210 ( .A1(n14197), .A2(n14198), .ZN(n13966) );
  NAND2_X1 U14211 ( .A1(a_10_), .A2(b_2_), .ZN(n14198) );
  INV_X1 U14212 ( .A(n14199), .ZN(n14197) );
  XOR2_X1 U14213 ( .A(n14200), .B(n14201), .Z(n13964) );
  XNOR2_X1 U14214 ( .A(n14202), .B(n14203), .ZN(n14201) );
  NAND2_X1 U14215 ( .A1(a_11_), .A2(b_1_), .ZN(n14200) );
  NAND2_X1 U14216 ( .A1(a_10_), .A2(n14199), .ZN(n13965) );
  NAND2_X1 U14217 ( .A1(n14204), .A2(n14205), .ZN(n14199) );
  NAND2_X1 U14218 ( .A1(n14118), .A2(n14206), .ZN(n14205) );
  OR2_X1 U14219 ( .A1(n14119), .A2(n14117), .ZN(n14206) );
  NOR2_X1 U14220 ( .A1(n7877), .A2(n13794), .ZN(n14118) );
  NAND2_X1 U14221 ( .A1(n14117), .A2(n14119), .ZN(n14204) );
  NAND2_X1 U14222 ( .A1(n13976), .A2(n14207), .ZN(n14119) );
  NAND2_X1 U14223 ( .A1(n13975), .A2(n13977), .ZN(n14207) );
  NAND2_X1 U14224 ( .A1(n14208), .A2(n14209), .ZN(n13977) );
  NAND2_X1 U14225 ( .A1(a_12_), .A2(b_2_), .ZN(n14209) );
  INV_X1 U14226 ( .A(n14210), .ZN(n14208) );
  XOR2_X1 U14227 ( .A(n14211), .B(n14212), .Z(n13975) );
  XNOR2_X1 U14228 ( .A(n14213), .B(n14214), .ZN(n14212) );
  NAND2_X1 U14229 ( .A1(a_13_), .A2(b_1_), .ZN(n14211) );
  NAND2_X1 U14230 ( .A1(a_12_), .A2(n14210), .ZN(n13976) );
  NAND2_X1 U14231 ( .A1(n14215), .A2(n14216), .ZN(n14210) );
  NAND2_X1 U14232 ( .A1(n14114), .A2(n14217), .ZN(n14216) );
  OR2_X1 U14233 ( .A1(n14115), .A2(n14113), .ZN(n14217) );
  NOR2_X1 U14234 ( .A1(n7355), .A2(n13794), .ZN(n14114) );
  NAND2_X1 U14235 ( .A1(n14113), .A2(n14115), .ZN(n14215) );
  NAND2_X1 U14236 ( .A1(n13987), .A2(n14218), .ZN(n14115) );
  NAND2_X1 U14237 ( .A1(n13986), .A2(n13988), .ZN(n14218) );
  NAND2_X1 U14238 ( .A1(n14219), .A2(n14220), .ZN(n13988) );
  NAND2_X1 U14239 ( .A1(a_14_), .A2(b_2_), .ZN(n14220) );
  INV_X1 U14240 ( .A(n14221), .ZN(n14219) );
  XOR2_X1 U14241 ( .A(n14222), .B(n14223), .Z(n13986) );
  XNOR2_X1 U14242 ( .A(n14224), .B(n14225), .ZN(n14223) );
  NAND2_X1 U14243 ( .A1(a_15_), .A2(b_1_), .ZN(n14222) );
  NAND2_X1 U14244 ( .A1(a_14_), .A2(n14221), .ZN(n13987) );
  NAND2_X1 U14245 ( .A1(n14226), .A2(n14227), .ZN(n14221) );
  NAND2_X1 U14246 ( .A1(n14110), .A2(n14228), .ZN(n14227) );
  OR2_X1 U14247 ( .A1(n14111), .A2(n14109), .ZN(n14228) );
  NOR2_X1 U14248 ( .A1(n7346), .A2(n13794), .ZN(n14110) );
  NAND2_X1 U14249 ( .A1(n14109), .A2(n14111), .ZN(n14226) );
  NAND2_X1 U14250 ( .A1(n13998), .A2(n14229), .ZN(n14111) );
  NAND2_X1 U14251 ( .A1(n13997), .A2(n13999), .ZN(n14229) );
  NAND2_X1 U14252 ( .A1(n14230), .A2(n14231), .ZN(n13999) );
  NAND2_X1 U14253 ( .A1(a_16_), .A2(b_2_), .ZN(n14231) );
  INV_X1 U14254 ( .A(n14232), .ZN(n14230) );
  XOR2_X1 U14255 ( .A(n14233), .B(n14234), .Z(n13997) );
  XNOR2_X1 U14256 ( .A(n14235), .B(n14236), .ZN(n14234) );
  NAND2_X1 U14257 ( .A1(a_17_), .A2(b_1_), .ZN(n14233) );
  NAND2_X1 U14258 ( .A1(a_16_), .A2(n14232), .ZN(n13998) );
  NAND2_X1 U14259 ( .A1(n14237), .A2(n14238), .ZN(n14232) );
  NAND2_X1 U14260 ( .A1(n14106), .A2(n14239), .ZN(n14238) );
  NAND2_X1 U14261 ( .A1(n14107), .A2(n14105), .ZN(n14239) );
  NOR2_X1 U14262 ( .A1(n7337), .A2(n13794), .ZN(n14106) );
  OR2_X1 U14263 ( .A1(n14105), .A2(n14107), .ZN(n14237) );
  AND2_X1 U14264 ( .A1(n14240), .A2(n14241), .ZN(n14107) );
  NAND2_X1 U14265 ( .A1(n14010), .A2(n14242), .ZN(n14241) );
  OR2_X1 U14266 ( .A1(n14009), .A2(n14007), .ZN(n14242) );
  NOR2_X1 U14267 ( .A1(n7764), .A2(n13794), .ZN(n14010) );
  NAND2_X1 U14268 ( .A1(n14007), .A2(n14009), .ZN(n14240) );
  NAND2_X1 U14269 ( .A1(n14243), .A2(n14244), .ZN(n14009) );
  NAND3_X1 U14270 ( .A1(b_2_), .A2(n14245), .A3(a_19_), .ZN(n14244) );
  NAND2_X1 U14271 ( .A1(n14103), .A2(n14101), .ZN(n14245) );
  OR2_X1 U14272 ( .A1(n14101), .A2(n14103), .ZN(n14243) );
  AND2_X1 U14273 ( .A1(n14246), .A2(n14247), .ZN(n14103) );
  NAND2_X1 U14274 ( .A1(n14021), .A2(n14248), .ZN(n14247) );
  OR2_X1 U14275 ( .A1(n14020), .A2(n14018), .ZN(n14248) );
  NOR2_X1 U14276 ( .A1(n7987), .A2(n13794), .ZN(n14021) );
  NAND2_X1 U14277 ( .A1(n14018), .A2(n14020), .ZN(n14246) );
  NAND2_X1 U14278 ( .A1(n14249), .A2(n14250), .ZN(n14020) );
  NAND3_X1 U14279 ( .A1(b_2_), .A2(n14251), .A3(a_21_), .ZN(n14250) );
  NAND2_X1 U14280 ( .A1(n14099), .A2(n14097), .ZN(n14251) );
  OR2_X1 U14281 ( .A1(n14097), .A2(n14099), .ZN(n14249) );
  AND2_X1 U14282 ( .A1(n14252), .A2(n14253), .ZN(n14099) );
  NAND2_X1 U14283 ( .A1(n14032), .A2(n14254), .ZN(n14253) );
  OR2_X1 U14284 ( .A1(n14031), .A2(n14029), .ZN(n14254) );
  NOR2_X1 U14285 ( .A1(n13794), .A2(n7312), .ZN(n14032) );
  NAND2_X1 U14286 ( .A1(n14029), .A2(n14031), .ZN(n14252) );
  NAND2_X1 U14287 ( .A1(n14255), .A2(n14256), .ZN(n14031) );
  NAND3_X1 U14288 ( .A1(a_23_), .A2(n14257), .A3(b_2_), .ZN(n14256) );
  OR2_X1 U14289 ( .A1(n14094), .A2(n14092), .ZN(n14257) );
  NAND2_X1 U14290 ( .A1(n14092), .A2(n14094), .ZN(n14255) );
  NAND2_X1 U14291 ( .A1(n14258), .A2(n14259), .ZN(n14094) );
  NAND2_X1 U14292 ( .A1(n14043), .A2(n14260), .ZN(n14259) );
  OR2_X1 U14293 ( .A1(n14042), .A2(n14040), .ZN(n14260) );
  NOR2_X1 U14294 ( .A1(n7691), .A2(n13794), .ZN(n14043) );
  NAND2_X1 U14295 ( .A1(n14040), .A2(n14042), .ZN(n14258) );
  NAND2_X1 U14296 ( .A1(n14090), .A2(n14261), .ZN(n14042) );
  NAND2_X1 U14297 ( .A1(n14089), .A2(n14091), .ZN(n14261) );
  NAND2_X1 U14298 ( .A1(n14262), .A2(n14263), .ZN(n14091) );
  NAND2_X1 U14299 ( .A1(b_2_), .A2(a_25_), .ZN(n14263) );
  INV_X1 U14300 ( .A(n14264), .ZN(n14262) );
  XOR2_X1 U14301 ( .A(n14265), .B(n14266), .Z(n14089) );
  NOR2_X1 U14302 ( .A1(n14267), .A2(n14268), .ZN(n14266) );
  XOR2_X1 U14303 ( .A(n14269), .B(n14270), .Z(n14265) );
  NAND2_X1 U14304 ( .A1(a_25_), .A2(n14264), .ZN(n14090) );
  NAND2_X1 U14305 ( .A1(n14271), .A2(n14272), .ZN(n14264) );
  NAND3_X1 U14306 ( .A1(a_26_), .A2(n14273), .A3(b_2_), .ZN(n14272) );
  NAND2_X1 U14307 ( .A1(n14054), .A2(n14052), .ZN(n14273) );
  OR2_X1 U14308 ( .A1(n14052), .A2(n14054), .ZN(n14271) );
  AND2_X1 U14309 ( .A1(n14274), .A2(n14275), .ZN(n14054) );
  NAND2_X1 U14310 ( .A1(n14062), .A2(n14276), .ZN(n14275) );
  OR2_X1 U14311 ( .A1(n14061), .A2(n14059), .ZN(n14276) );
  NOR2_X1 U14312 ( .A1(n13794), .A2(n14267), .ZN(n14062) );
  NAND2_X1 U14313 ( .A1(n14059), .A2(n14061), .ZN(n14274) );
  NAND2_X1 U14314 ( .A1(n14277), .A2(n14278), .ZN(n14061) );
  NAND3_X1 U14315 ( .A1(a_28_), .A2(n14279), .A3(b_2_), .ZN(n14278) );
  OR2_X1 U14316 ( .A1(n14068), .A2(n14070), .ZN(n14279) );
  NAND2_X1 U14317 ( .A1(n14068), .A2(n14070), .ZN(n14277) );
  NAND2_X1 U14318 ( .A1(n14280), .A2(n14281), .ZN(n14070) );
  NAND3_X1 U14319 ( .A1(a_29_), .A2(n14282), .A3(b_2_), .ZN(n14281) );
  OR2_X1 U14320 ( .A1(n14086), .A2(n14087), .ZN(n14282) );
  NAND2_X1 U14321 ( .A1(n14087), .A2(n14086), .ZN(n14280) );
  NAND2_X1 U14322 ( .A1(n14283), .A2(n14284), .ZN(n14086) );
  NAND2_X1 U14323 ( .A1(b_0_), .A2(n14285), .ZN(n14284) );
  NAND2_X1 U14324 ( .A1(n7268), .A2(n14286), .ZN(n14285) );
  NAND2_X1 U14325 ( .A1(a_31_), .A2(n14083), .ZN(n14286) );
  NAND2_X1 U14326 ( .A1(b_1_), .A2(n14288), .ZN(n14283) );
  NAND2_X1 U14327 ( .A1(n7272), .A2(n14289), .ZN(n14288) );
  NAND2_X1 U14328 ( .A1(a_30_), .A2(n14268), .ZN(n14289) );
  AND3_X1 U14329 ( .A1(b_2_), .A2(n7954), .A3(b_1_), .ZN(n14087) );
  XNOR2_X1 U14330 ( .A(n14291), .B(n14292), .ZN(n14068) );
  NOR2_X1 U14331 ( .A1(n14287), .A2(n14268), .ZN(n14292) );
  XOR2_X1 U14332 ( .A(n14293), .B(n14294), .Z(n14291) );
  XOR2_X1 U14333 ( .A(n14295), .B(n14296), .Z(n14059) );
  XNOR2_X1 U14334 ( .A(n14297), .B(n14298), .ZN(n14296) );
  NAND2_X1 U14335 ( .A1(b_0_), .A2(a_29_), .ZN(n14295) );
  XNOR2_X1 U14336 ( .A(n14299), .B(n14300), .ZN(n14052) );
  XNOR2_X1 U14337 ( .A(n14301), .B(n14302), .ZN(n14300) );
  NAND2_X1 U14338 ( .A1(b_0_), .A2(a_28_), .ZN(n14299) );
  XOR2_X1 U14339 ( .A(n14303), .B(n14304), .Z(n14040) );
  XNOR2_X1 U14340 ( .A(n14305), .B(n14306), .ZN(n14304) );
  NAND2_X1 U14341 ( .A1(b_0_), .A2(a_26_), .ZN(n14303) );
  XOR2_X1 U14342 ( .A(n14307), .B(n14308), .Z(n14092) );
  NOR2_X1 U14343 ( .A1(n7923), .A2(n14268), .ZN(n14308) );
  XOR2_X1 U14344 ( .A(n14309), .B(n14310), .Z(n14307) );
  XOR2_X1 U14345 ( .A(n14311), .B(n14312), .Z(n14029) );
  XNOR2_X1 U14346 ( .A(n14313), .B(n14314), .ZN(n14312) );
  NAND2_X1 U14347 ( .A1(b_0_), .A2(a_24_), .ZN(n14311) );
  XNOR2_X1 U14348 ( .A(n14315), .B(n14316), .ZN(n14097) );
  NOR2_X1 U14349 ( .A1(n7916), .A2(n14268), .ZN(n14316) );
  XOR2_X1 U14350 ( .A(n14317), .B(n14318), .Z(n14315) );
  XOR2_X1 U14351 ( .A(n14319), .B(n14320), .Z(n14018) );
  XNOR2_X1 U14352 ( .A(n14321), .B(n14322), .ZN(n14320) );
  NAND2_X1 U14353 ( .A1(b_0_), .A2(a_22_), .ZN(n14319) );
  XNOR2_X1 U14354 ( .A(n14323), .B(n14324), .ZN(n14101) );
  NOR2_X1 U14355 ( .A1(n14268), .A2(n7909), .ZN(n14324) );
  XOR2_X1 U14356 ( .A(n14325), .B(n14326), .Z(n14323) );
  XOR2_X1 U14357 ( .A(n14327), .B(n14328), .Z(n14007) );
  XNOR2_X1 U14358 ( .A(n14329), .B(n14330), .ZN(n14328) );
  NAND2_X1 U14359 ( .A1(a_20_), .A2(b_0_), .ZN(n14327) );
  XNOR2_X1 U14360 ( .A(n14331), .B(n14332), .ZN(n14105) );
  NOR2_X1 U14361 ( .A1(n14268), .A2(n7902), .ZN(n14332) );
  XOR2_X1 U14362 ( .A(n14333), .B(n14334), .Z(n14331) );
  XOR2_X1 U14363 ( .A(n14335), .B(n14336), .Z(n14109) );
  NOR2_X1 U14364 ( .A1(n14083), .A2(n7773), .ZN(n14336) );
  XOR2_X1 U14365 ( .A(n14337), .B(n14338), .Z(n14335) );
  XOR2_X1 U14366 ( .A(n14339), .B(n14340), .Z(n14113) );
  NOR2_X1 U14367 ( .A1(n14083), .A2(n7782), .ZN(n14340) );
  XOR2_X1 U14368 ( .A(n14341), .B(n14342), .Z(n14339) );
  XOR2_X1 U14369 ( .A(n14343), .B(n14344), .Z(n14117) );
  NOR2_X1 U14370 ( .A1(n14083), .A2(n8020), .ZN(n14344) );
  XOR2_X1 U14371 ( .A(n14345), .B(n14346), .Z(n14343) );
  XOR2_X1 U14372 ( .A(n14347), .B(n14348), .Z(n14121) );
  NOR2_X1 U14373 ( .A1(n14083), .A2(n7799), .ZN(n14348) );
  XOR2_X1 U14374 ( .A(n14349), .B(n14350), .Z(n14347) );
  XOR2_X1 U14375 ( .A(n14351), .B(n14352), .Z(n14125) );
  NOR2_X1 U14376 ( .A1(n14083), .A2(n8037), .ZN(n14352) );
  XOR2_X1 U14377 ( .A(n14353), .B(n14354), .Z(n14351) );
  XOR2_X1 U14378 ( .A(n14355), .B(n14356), .Z(n14129) );
  NOR2_X1 U14379 ( .A1(n14083), .A2(n7388), .ZN(n14356) );
  XOR2_X1 U14380 ( .A(n14357), .B(n14358), .Z(n14355) );
  XOR2_X1 U14381 ( .A(n14359), .B(n14360), .Z(n14133) );
  NOR2_X1 U14382 ( .A1(n14083), .A2(n7398), .ZN(n14360) );
  XOR2_X1 U14383 ( .A(n14361), .B(n14362), .Z(n14359) );
  XOR2_X1 U14384 ( .A(n14363), .B(n14364), .Z(n13920) );
  XNOR2_X1 U14385 ( .A(n14365), .B(n14366), .ZN(n14364) );
  NAND2_X1 U14386 ( .A1(a_3_), .A2(b_1_), .ZN(n14363) );
  XOR2_X1 U14387 ( .A(n14367), .B(n14368), .Z(n14137) );
  NOR2_X1 U14388 ( .A1(n14083), .A2(n7832), .ZN(n14368) );
  XOR2_X1 U14389 ( .A(n14369), .B(n14370), .Z(n14367) );
  XNOR2_X1 U14390 ( .A(n14371), .B(n14372), .ZN(n7513) );
  NOR2_X1 U14391 ( .A1(n14268), .A2(n7411), .ZN(n14372) );
  XOR2_X1 U14392 ( .A(n14373), .B(n14374), .Z(n14371) );
  XOR2_X1 U14393 ( .A(n7512), .B(n7511), .Z(n14144) );
  NAND2_X1 U14394 ( .A1(n14375), .A2(n14376), .ZN(n7511) );
  NAND3_X1 U14395 ( .A1(b_0_), .A2(n14377), .A3(a_1_), .ZN(n14376) );
  OR2_X1 U14396 ( .A1(n14374), .A2(n14373), .ZN(n14377) );
  NAND2_X1 U14397 ( .A1(n14373), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U14398 ( .A1(n14378), .A2(n14379), .ZN(n14374) );
  NAND2_X1 U14399 ( .A1(n14150), .A2(n14380), .ZN(n14379) );
  OR2_X1 U14400 ( .A1(n14153), .A2(n14152), .ZN(n14380) );
  NOR2_X1 U14401 ( .A1(n7832), .A2(n14268), .ZN(n14150) );
  NAND2_X1 U14402 ( .A1(n14152), .A2(n14153), .ZN(n14378) );
  NAND2_X1 U14403 ( .A1(n14381), .A2(n14382), .ZN(n14153) );
  NAND3_X1 U14404 ( .A1(b_1_), .A2(n14383), .A3(a_2_), .ZN(n14382) );
  OR2_X1 U14405 ( .A1(n14370), .A2(n14369), .ZN(n14383) );
  NAND2_X1 U14406 ( .A1(n14369), .A2(n14370), .ZN(n14381) );
  NAND2_X1 U14407 ( .A1(n14384), .A2(n14385), .ZN(n14370) );
  NAND3_X1 U14408 ( .A1(b_1_), .A2(n14386), .A3(a_3_), .ZN(n14385) );
  OR2_X1 U14409 ( .A1(n14366), .A2(n14365), .ZN(n14386) );
  NAND2_X1 U14410 ( .A1(n14365), .A2(n14366), .ZN(n14384) );
  NAND2_X1 U14411 ( .A1(n14387), .A2(n14388), .ZN(n14366) );
  NAND3_X1 U14412 ( .A1(b_1_), .A2(n14389), .A3(a_4_), .ZN(n14388) );
  OR2_X1 U14413 ( .A1(n14362), .A2(n14361), .ZN(n14389) );
  NAND2_X1 U14414 ( .A1(n14361), .A2(n14362), .ZN(n14387) );
  NAND2_X1 U14415 ( .A1(n14390), .A2(n14391), .ZN(n14362) );
  NAND3_X1 U14416 ( .A1(b_1_), .A2(n14392), .A3(a_5_), .ZN(n14391) );
  OR2_X1 U14417 ( .A1(n14170), .A2(n14169), .ZN(n14392) );
  NAND2_X1 U14418 ( .A1(n14169), .A2(n14170), .ZN(n14390) );
  NAND2_X1 U14419 ( .A1(n14393), .A2(n14394), .ZN(n14170) );
  NAND3_X1 U14420 ( .A1(b_1_), .A2(n14395), .A3(a_6_), .ZN(n14394) );
  OR2_X1 U14421 ( .A1(n14358), .A2(n14357), .ZN(n14395) );
  NAND2_X1 U14422 ( .A1(n14357), .A2(n14358), .ZN(n14393) );
  NAND2_X1 U14423 ( .A1(n14396), .A2(n14397), .ZN(n14358) );
  NAND3_X1 U14424 ( .A1(b_1_), .A2(n14398), .A3(a_7_), .ZN(n14397) );
  OR2_X1 U14425 ( .A1(n14181), .A2(n14180), .ZN(n14398) );
  NAND2_X1 U14426 ( .A1(n14180), .A2(n14181), .ZN(n14396) );
  NAND2_X1 U14427 ( .A1(n14399), .A2(n14400), .ZN(n14181) );
  NAND3_X1 U14428 ( .A1(b_1_), .A2(n14401), .A3(a_8_), .ZN(n14400) );
  OR2_X1 U14429 ( .A1(n14354), .A2(n14353), .ZN(n14401) );
  NAND2_X1 U14430 ( .A1(n14353), .A2(n14354), .ZN(n14399) );
  NAND2_X1 U14431 ( .A1(n14402), .A2(n14403), .ZN(n14354) );
  NAND3_X1 U14432 ( .A1(a_9_), .A2(n14404), .A3(b_1_), .ZN(n14403) );
  OR2_X1 U14433 ( .A1(n14192), .A2(n14191), .ZN(n14404) );
  NAND2_X1 U14434 ( .A1(n14191), .A2(n14192), .ZN(n14402) );
  NAND2_X1 U14435 ( .A1(n14405), .A2(n14406), .ZN(n14192) );
  NAND3_X1 U14436 ( .A1(b_1_), .A2(n14407), .A3(a_10_), .ZN(n14406) );
  OR2_X1 U14437 ( .A1(n14350), .A2(n14349), .ZN(n14407) );
  NAND2_X1 U14438 ( .A1(n14349), .A2(n14350), .ZN(n14405) );
  NAND2_X1 U14439 ( .A1(n14408), .A2(n14409), .ZN(n14350) );
  NAND3_X1 U14440 ( .A1(b_1_), .A2(n14410), .A3(a_11_), .ZN(n14409) );
  OR2_X1 U14441 ( .A1(n14203), .A2(n14202), .ZN(n14410) );
  NAND2_X1 U14442 ( .A1(n14202), .A2(n14203), .ZN(n14408) );
  NAND2_X1 U14443 ( .A1(n14411), .A2(n14412), .ZN(n14203) );
  NAND3_X1 U14444 ( .A1(b_1_), .A2(n14413), .A3(a_12_), .ZN(n14412) );
  OR2_X1 U14445 ( .A1(n14346), .A2(n14345), .ZN(n14413) );
  NAND2_X1 U14446 ( .A1(n14345), .A2(n14346), .ZN(n14411) );
  NAND2_X1 U14447 ( .A1(n14414), .A2(n14415), .ZN(n14346) );
  NAND3_X1 U14448 ( .A1(b_1_), .A2(n14416), .A3(a_13_), .ZN(n14415) );
  OR2_X1 U14449 ( .A1(n14214), .A2(n14213), .ZN(n14416) );
  NAND2_X1 U14450 ( .A1(n14213), .A2(n14214), .ZN(n14414) );
  NAND2_X1 U14451 ( .A1(n14417), .A2(n14418), .ZN(n14214) );
  NAND3_X1 U14452 ( .A1(b_1_), .A2(n14419), .A3(a_14_), .ZN(n14418) );
  OR2_X1 U14453 ( .A1(n14342), .A2(n14341), .ZN(n14419) );
  NAND2_X1 U14454 ( .A1(n14341), .A2(n14342), .ZN(n14417) );
  NAND2_X1 U14455 ( .A1(n14420), .A2(n14421), .ZN(n14342) );
  NAND3_X1 U14456 ( .A1(b_1_), .A2(n14422), .A3(a_15_), .ZN(n14421) );
  OR2_X1 U14457 ( .A1(n14225), .A2(n14224), .ZN(n14422) );
  NAND2_X1 U14458 ( .A1(n14224), .A2(n14225), .ZN(n14420) );
  NAND2_X1 U14459 ( .A1(n14423), .A2(n14424), .ZN(n14225) );
  NAND3_X1 U14460 ( .A1(b_1_), .A2(n14425), .A3(a_16_), .ZN(n14424) );
  OR2_X1 U14461 ( .A1(n14338), .A2(n14337), .ZN(n14425) );
  NAND2_X1 U14462 ( .A1(n14337), .A2(n14338), .ZN(n14423) );
  NAND2_X1 U14463 ( .A1(n14426), .A2(n14427), .ZN(n14338) );
  NAND3_X1 U14464 ( .A1(b_1_), .A2(n14428), .A3(a_17_), .ZN(n14427) );
  OR2_X1 U14465 ( .A1(n14236), .A2(n14235), .ZN(n14428) );
  NAND2_X1 U14466 ( .A1(n14235), .A2(n14236), .ZN(n14426) );
  NAND2_X1 U14467 ( .A1(n14429), .A2(n14430), .ZN(n14236) );
  NAND3_X1 U14468 ( .A1(b_0_), .A2(n14431), .A3(a_19_), .ZN(n14430) );
  OR2_X1 U14469 ( .A1(n14334), .A2(n14333), .ZN(n14431) );
  NAND2_X1 U14470 ( .A1(n14333), .A2(n14334), .ZN(n14429) );
  NAND2_X1 U14471 ( .A1(n14432), .A2(n14433), .ZN(n14334) );
  NAND3_X1 U14472 ( .A1(b_0_), .A2(n14434), .A3(a_20_), .ZN(n14433) );
  OR2_X1 U14473 ( .A1(n14330), .A2(n14329), .ZN(n14434) );
  NAND2_X1 U14474 ( .A1(n14329), .A2(n14330), .ZN(n14432) );
  NAND2_X1 U14475 ( .A1(n14435), .A2(n14436), .ZN(n14330) );
  NAND3_X1 U14476 ( .A1(b_0_), .A2(n14437), .A3(a_21_), .ZN(n14436) );
  NAND2_X1 U14477 ( .A1(n14326), .A2(n14325), .ZN(n14437) );
  INV_X1 U14478 ( .A(n14438), .ZN(n14326) );
  NAND2_X1 U14479 ( .A1(n14439), .A2(n14438), .ZN(n14435) );
  NAND2_X1 U14480 ( .A1(n14440), .A2(n14441), .ZN(n14438) );
  NAND3_X1 U14481 ( .A1(a_22_), .A2(n14442), .A3(b_0_), .ZN(n14441) );
  OR2_X1 U14482 ( .A1(n14322), .A2(n14321), .ZN(n14442) );
  NAND2_X1 U14483 ( .A1(n14321), .A2(n14322), .ZN(n14440) );
  NAND2_X1 U14484 ( .A1(n14443), .A2(n14444), .ZN(n14322) );
  NAND3_X1 U14485 ( .A1(a_23_), .A2(n14445), .A3(b_0_), .ZN(n14444) );
  NAND2_X1 U14486 ( .A1(n14318), .A2(n14317), .ZN(n14445) );
  INV_X1 U14487 ( .A(n14446), .ZN(n14318) );
  NAND2_X1 U14488 ( .A1(n14447), .A2(n14446), .ZN(n14443) );
  NAND2_X1 U14489 ( .A1(n14448), .A2(n14449), .ZN(n14446) );
  NAND3_X1 U14490 ( .A1(a_24_), .A2(n14450), .A3(b_0_), .ZN(n14449) );
  OR2_X1 U14491 ( .A1(n14314), .A2(n14313), .ZN(n14450) );
  NAND2_X1 U14492 ( .A1(n14313), .A2(n14314), .ZN(n14448) );
  NAND2_X1 U14493 ( .A1(n14451), .A2(n14452), .ZN(n14314) );
  NAND3_X1 U14494 ( .A1(a_25_), .A2(n14453), .A3(b_0_), .ZN(n14452) );
  NAND2_X1 U14495 ( .A1(n14310), .A2(n14309), .ZN(n14453) );
  INV_X1 U14496 ( .A(n14454), .ZN(n14310) );
  NAND2_X1 U14497 ( .A1(n14455), .A2(n14454), .ZN(n14451) );
  NAND2_X1 U14498 ( .A1(n14456), .A2(n14457), .ZN(n14454) );
  NAND3_X1 U14499 ( .A1(a_26_), .A2(n14458), .A3(b_0_), .ZN(n14457) );
  OR2_X1 U14500 ( .A1(n14306), .A2(n14305), .ZN(n14458) );
  NAND2_X1 U14501 ( .A1(n14305), .A2(n14306), .ZN(n14456) );
  NAND2_X1 U14502 ( .A1(n14459), .A2(n14460), .ZN(n14306) );
  NAND3_X1 U14503 ( .A1(a_27_), .A2(n14461), .A3(b_0_), .ZN(n14460) );
  NAND2_X1 U14504 ( .A1(n14270), .A2(n14269), .ZN(n14461) );
  INV_X1 U14505 ( .A(n14462), .ZN(n14270) );
  NAND2_X1 U14506 ( .A1(n14463), .A2(n14462), .ZN(n14459) );
  NAND2_X1 U14507 ( .A1(n14464), .A2(n14465), .ZN(n14462) );
  NAND3_X1 U14508 ( .A1(a_28_), .A2(n14466), .A3(b_0_), .ZN(n14465) );
  OR2_X1 U14509 ( .A1(n14302), .A2(n14301), .ZN(n14466) );
  NAND2_X1 U14510 ( .A1(n14301), .A2(n14302), .ZN(n14464) );
  NAND2_X1 U14511 ( .A1(n14467), .A2(n14468), .ZN(n14302) );
  NAND3_X1 U14512 ( .A1(a_29_), .A2(n14469), .A3(b_0_), .ZN(n14468) );
  OR2_X1 U14513 ( .A1(n14298), .A2(n14297), .ZN(n14469) );
  NAND2_X1 U14514 ( .A1(n14297), .A2(n14298), .ZN(n14467) );
  NAND2_X1 U14515 ( .A1(n14294), .A2(n14470), .ZN(n14298) );
  NAND3_X1 U14516 ( .A1(b_0_), .A2(a_30_), .A3(n14293), .ZN(n14470) );
  NOR2_X1 U14517 ( .A1(n14083), .A2(n7946), .ZN(n14293) );
  NAND3_X1 U14518 ( .A1(b_1_), .A2(n7954), .A3(b_0_), .ZN(n14294) );
  INV_X1 U14519 ( .A(a_31_), .ZN(n14290) );
  NOR2_X1 U14520 ( .A1(n14083), .A2(n14471), .ZN(n14297) );
  NOR2_X1 U14521 ( .A1(n14083), .A2(n14267), .ZN(n14301) );
  INV_X1 U14522 ( .A(n14269), .ZN(n14463) );
  NAND2_X1 U14523 ( .A1(b_1_), .A2(a_26_), .ZN(n14269) );
  NOR2_X1 U14524 ( .A1(n14083), .A2(n7923), .ZN(n14305) );
  INV_X1 U14525 ( .A(n14309), .ZN(n14455) );
  NAND2_X1 U14526 ( .A1(b_1_), .A2(a_24_), .ZN(n14309) );
  NOR2_X1 U14527 ( .A1(n14083), .A2(n7916), .ZN(n14313) );
  INV_X1 U14528 ( .A(n14317), .ZN(n14447) );
  NAND2_X1 U14529 ( .A1(b_1_), .A2(a_22_), .ZN(n14317) );
  NOR2_X1 U14530 ( .A1(n7909), .A2(n14083), .ZN(n14321) );
  INV_X1 U14531 ( .A(n14325), .ZN(n14439) );
  NAND2_X1 U14532 ( .A1(a_20_), .A2(b_1_), .ZN(n14325) );
  NOR2_X1 U14533 ( .A1(n7902), .A2(n14083), .ZN(n14329) );
  NOR2_X1 U14534 ( .A1(n7764), .A2(n14083), .ZN(n14333) );
  NOR2_X1 U14535 ( .A1(n7764), .A2(n14268), .ZN(n14235) );
  NOR2_X1 U14536 ( .A1(n7337), .A2(n14268), .ZN(n14337) );
  NOR2_X1 U14537 ( .A1(n7773), .A2(n14268), .ZN(n14224) );
  NOR2_X1 U14538 ( .A1(n7346), .A2(n14268), .ZN(n14341) );
  NOR2_X1 U14539 ( .A1(n7782), .A2(n14268), .ZN(n14213) );
  NOR2_X1 U14540 ( .A1(n7355), .A2(n14268), .ZN(n14345) );
  NOR2_X1 U14541 ( .A1(n8020), .A2(n14268), .ZN(n14202) );
  NOR2_X1 U14542 ( .A1(n7877), .A2(n14268), .ZN(n14349) );
  NOR2_X1 U14543 ( .A1(n7799), .A2(n14268), .ZN(n14191) );
  NOR2_X1 U14544 ( .A1(n14268), .A2(n7870), .ZN(n14353) );
  NOR2_X1 U14545 ( .A1(n8037), .A2(n14268), .ZN(n14180) );
  NOR2_X1 U14546 ( .A1(n7863), .A2(n14268), .ZN(n14357) );
  NOR2_X1 U14547 ( .A1(n7388), .A2(n14268), .ZN(n14169) );
  NOR2_X1 U14548 ( .A1(n7393), .A2(n14268), .ZN(n14361) );
  NOR2_X1 U14549 ( .A1(n7398), .A2(n14268), .ZN(n14365) );
  NOR2_X1 U14550 ( .A1(n7850), .A2(n14268), .ZN(n14369) );
  INV_X1 U14551 ( .A(b_0_), .ZN(n14268) );
  NOR2_X1 U14552 ( .A1(n14083), .A2(n7613), .ZN(n14373) );
  INV_X1 U14553 ( .A(a_0_), .ZN(n7613) );
  NAND3_X1 U14554 ( .A1(n14472), .A2(n14473), .A3(n14474), .ZN(Result_add_9_)
         );
  NAND2_X1 U14555 ( .A1(n12361), .A2(n14475), .ZN(n14474) );
  INV_X1 U14556 ( .A(n14476), .ZN(n12361) );
  NAND3_X1 U14557 ( .A1(n14477), .A2(n7870), .A3(b_9_), .ZN(n14473) );
  NAND2_X1 U14558 ( .A1(n14478), .A2(n12224), .ZN(n14472) );
  XOR2_X1 U14559 ( .A(n14475), .B(a_9_), .Z(n14478) );
  XOR2_X1 U14560 ( .A(n14479), .B(n14480), .Z(Result_add_8_) );
  AND2_X1 U14561 ( .A1(n14481), .A2(n12748), .ZN(n14480) );
  NAND3_X1 U14562 ( .A1(n14482), .A2(n14483), .A3(n14484), .ZN(Result_add_7_)
         );
  NAND2_X1 U14563 ( .A1(n12976), .A2(n14485), .ZN(n14484) );
  INV_X1 U14564 ( .A(n14486), .ZN(n12976) );
  OR3_X1 U14565 ( .A1(n14485), .A2(a_7_), .A3(n12673), .ZN(n14483) );
  NAND2_X1 U14566 ( .A1(n14487), .A2(n12673), .ZN(n14482) );
  XOR2_X1 U14567 ( .A(n14485), .B(a_7_), .Z(n14487) );
  XNOR2_X1 U14568 ( .A(n14488), .B(n14489), .ZN(Result_add_6_) );
  NOR2_X1 U14569 ( .A1(n14490), .A2(n13209), .ZN(n14489) );
  NAND3_X1 U14570 ( .A1(n14491), .A2(n14492), .A3(n14493), .ZN(Result_add_5_)
         );
  NAND2_X1 U14571 ( .A1(n13436), .A2(n14494), .ZN(n14493) );
  INV_X1 U14572 ( .A(n14495), .ZN(n13436) );
  NAND3_X1 U14573 ( .A1(n14496), .A2(n7393), .A3(b_5_), .ZN(n14492) );
  NAND2_X1 U14574 ( .A1(n14497), .A2(n13129), .ZN(n14491) );
  XOR2_X1 U14575 ( .A(n14494), .B(a_5_), .Z(n14497) );
  XNOR2_X1 U14576 ( .A(n14498), .B(n14499), .ZN(Result_add_4_) );
  NOR2_X1 U14577 ( .A1(n14500), .A2(n13669), .ZN(n14499) );
  NAND3_X1 U14578 ( .A1(n14501), .A2(n14502), .A3(n14503), .ZN(Result_add_3_)
         );
  NAND2_X1 U14579 ( .A1(n13894), .A2(n14504), .ZN(n14503) );
  INV_X1 U14580 ( .A(n14505), .ZN(n13894) );
  NAND3_X1 U14581 ( .A1(n14506), .A2(n7850), .A3(b_3_), .ZN(n14502) );
  NAND2_X1 U14582 ( .A1(n14507), .A2(n13581), .ZN(n14501) );
  XOR2_X1 U14583 ( .A(n14504), .B(a_3_), .Z(n14507) );
  XOR2_X1 U14584 ( .A(b_31_), .B(a_31_), .Z(Result_add_31_) );
  NAND3_X1 U14585 ( .A1(n14508), .A2(n14509), .A3(n7277), .ZN(Result_add_30_)
         );
  NAND2_X1 U14586 ( .A1(Result_mul_63_), .A2(n7724), .ZN(n7277) );
  INV_X1 U14587 ( .A(n14510), .ZN(n7724) );
  NAND2_X1 U14588 ( .A1(n14511), .A2(n7274), .ZN(n14509) );
  XOR2_X1 U14589 ( .A(n14287), .B(n14512), .Z(n14511) );
  NAND3_X1 U14590 ( .A1(n14512), .A2(n14287), .A3(b_30_), .ZN(n14508) );
  XNOR2_X1 U14591 ( .A(n14513), .B(n14514), .ZN(Result_add_2_) );
  NOR2_X1 U14592 ( .A1(n14515), .A2(n13922), .ZN(n14514) );
  NAND3_X1 U14593 ( .A1(n14516), .A2(n14517), .A3(n14518), .ZN(Result_add_29_)
         );
  NAND2_X1 U14594 ( .A1(n7956), .A2(n14519), .ZN(n14518) );
  INV_X1 U14595 ( .A(n14520), .ZN(n7956) );
  NAND3_X1 U14596 ( .A1(n14521), .A2(n7946), .A3(b_29_), .ZN(n14517) );
  NAND2_X1 U14597 ( .A1(n14522), .A2(n7725), .ZN(n14516) );
  XOR2_X1 U14598 ( .A(n7946), .B(n14521), .Z(n14522) );
  INV_X1 U14599 ( .A(n14519), .ZN(n14521) );
  XNOR2_X1 U14600 ( .A(n14523), .B(n14524), .ZN(Result_add_28_) );
  NAND2_X1 U14601 ( .A1(n8169), .A2(n14525), .ZN(n14523) );
  NAND3_X1 U14602 ( .A1(n14526), .A2(n14527), .A3(n14528), .ZN(Result_add_27_)
         );
  NAND2_X1 U14603 ( .A1(n8381), .A2(n14529), .ZN(n14528) );
  INV_X1 U14604 ( .A(n14530), .ZN(n8381) );
  OR3_X1 U14605 ( .A1(n14529), .A2(a_27_), .A3(n8183), .ZN(n14527) );
  NAND2_X1 U14606 ( .A1(n14531), .A2(n8183), .ZN(n14526) );
  XOR2_X1 U14607 ( .A(n14529), .B(a_27_), .Z(n14531) );
  XOR2_X1 U14608 ( .A(n14532), .B(n14533), .Z(Result_add_26_) );
  AND2_X1 U14609 ( .A1(n14534), .A2(n8827), .ZN(n14533) );
  NAND3_X1 U14610 ( .A1(n14535), .A2(n14536), .A3(n14537), .ZN(Result_add_25_)
         );
  NAND2_X1 U14611 ( .A1(n8864), .A2(n14538), .ZN(n14537) );
  INV_X1 U14612 ( .A(n14539), .ZN(n8864) );
  OR3_X1 U14613 ( .A1(n14538), .A2(a_25_), .A3(n8639), .ZN(n14536) );
  NAND2_X1 U14614 ( .A1(n14540), .A2(n8639), .ZN(n14535) );
  XOR2_X1 U14615 ( .A(n14538), .B(a_25_), .Z(n14540) );
  XNOR2_X1 U14616 ( .A(n14541), .B(n14542), .ZN(Result_add_24_) );
  NOR2_X1 U14617 ( .A1(n14543), .A2(n9087), .ZN(n14542) );
  NAND3_X1 U14618 ( .A1(n14544), .A2(n14545), .A3(n14546), .ZN(Result_add_23_)
         );
  NAND2_X1 U14619 ( .A1(n9332), .A2(n14547), .ZN(n14546) );
  NAND3_X1 U14620 ( .A1(n14548), .A2(n7916), .A3(b_23_), .ZN(n14545) );
  NAND2_X1 U14621 ( .A1(n14549), .A2(n9071), .ZN(n14544) );
  XOR2_X1 U14622 ( .A(n14547), .B(a_23_), .Z(n14549) );
  XNOR2_X1 U14623 ( .A(n14550), .B(n14551), .ZN(Result_add_22_) );
  NOR2_X1 U14624 ( .A1(n14552), .A2(n9561), .ZN(n14551) );
  NAND3_X1 U14625 ( .A1(n14553), .A2(n14554), .A3(n14555), .ZN(Result_add_21_)
         );
  NAND2_X1 U14626 ( .A1(n9774), .A2(n14556), .ZN(n14555) );
  INV_X1 U14627 ( .A(n14557), .ZN(n9774) );
  NAND3_X1 U14628 ( .A1(n14558), .A2(n7909), .A3(b_21_), .ZN(n14554) );
  NAND2_X1 U14629 ( .A1(n14559), .A2(n9537), .ZN(n14553) );
  XOR2_X1 U14630 ( .A(n14556), .B(a_21_), .Z(n14559) );
  XOR2_X1 U14631 ( .A(n14560), .B(n14561), .Z(Result_add_20_) );
  AND2_X1 U14632 ( .A1(n14562), .A2(n10163), .ZN(n14561) );
  NAND2_X1 U14633 ( .A1(n14563), .A2(n14564), .ZN(Result_add_1_) );
  NAND2_X1 U14634 ( .A1(n14565), .A2(n14566), .ZN(n14564) );
  OR2_X1 U14635 ( .A1(n14152), .A2(n14567), .ZN(n14565) );
  NAND2_X1 U14636 ( .A1(n14568), .A2(n14569), .ZN(n14563) );
  XOR2_X1 U14637 ( .A(b_1_), .B(a_1_), .Z(n14568) );
  NAND3_X1 U14638 ( .A1(n14570), .A2(n14571), .A3(n14572), .ZN(Result_add_19_)
         );
  NAND2_X1 U14639 ( .A1(n10243), .A2(n14573), .ZN(n14572) );
  INV_X1 U14640 ( .A(n14574), .ZN(n10243) );
  OR3_X1 U14641 ( .A1(n14573), .A2(a_19_), .A3(n9964), .ZN(n14571) );
  NAND2_X1 U14642 ( .A1(n14575), .A2(n9964), .ZN(n14570) );
  XOR2_X1 U14643 ( .A(n14573), .B(a_19_), .Z(n14575) );
  XNOR2_X1 U14644 ( .A(n14576), .B(n14577), .ZN(Result_add_18_) );
  NOR2_X1 U14645 ( .A1(n14578), .A2(n10460), .ZN(n14577) );
  NAND3_X1 U14646 ( .A1(n14579), .A2(n14580), .A3(n14581), .ZN(Result_add_17_)
         );
  NAND2_X1 U14647 ( .A1(n10723), .A2(n14582), .ZN(n14581) );
  INV_X1 U14648 ( .A(n14583), .ZN(n10723) );
  NAND3_X1 U14649 ( .A1(n14584), .A2(n7337), .A3(b_17_), .ZN(n14580) );
  NAND2_X1 U14650 ( .A1(n14585), .A2(n10420), .ZN(n14579) );
  XOR2_X1 U14651 ( .A(n14582), .B(a_17_), .Z(n14585) );
  XNOR2_X1 U14652 ( .A(n14586), .B(n14587), .ZN(Result_add_16_) );
  NOR2_X1 U14653 ( .A1(n14588), .A2(n10910), .ZN(n14587) );
  NAND3_X1 U14654 ( .A1(n14589), .A2(n14590), .A3(n14591), .ZN(Result_add_15_)
         );
  NAND2_X1 U14655 ( .A1(n11150), .A2(n14592), .ZN(n14591) );
  NAND3_X1 U14656 ( .A1(n14593), .A2(n7346), .A3(b_15_), .ZN(n14590) );
  NAND2_X1 U14657 ( .A1(n14594), .A2(n10863), .ZN(n14589) );
  XOR2_X1 U14658 ( .A(n14592), .B(a_15_), .Z(n14594) );
  XNOR2_X1 U14659 ( .A(n14595), .B(n14596), .ZN(Result_add_14_) );
  NOR2_X1 U14660 ( .A1(n14597), .A2(n11370), .ZN(n14596) );
  NAND3_X1 U14661 ( .A1(n14598), .A2(n14599), .A3(n14600), .ZN(Result_add_13_)
         );
  NAND2_X1 U14662 ( .A1(n11615), .A2(n14601), .ZN(n14600) );
  INV_X1 U14663 ( .A(n14602), .ZN(n11615) );
  NAND3_X1 U14664 ( .A1(n14603), .A2(n7355), .A3(b_13_), .ZN(n14599) );
  NAND2_X1 U14665 ( .A1(n14604), .A2(n11322), .ZN(n14598) );
  XOR2_X1 U14666 ( .A(n14601), .B(a_13_), .Z(n14604) );
  XNOR2_X1 U14667 ( .A(n14605), .B(n14606), .ZN(Result_add_12_) );
  NOR2_X1 U14668 ( .A1(n14607), .A2(n11824), .ZN(n14606) );
  NAND3_X1 U14669 ( .A1(n14608), .A2(n14609), .A3(n14610), .ZN(Result_add_11_)
         );
  NAND2_X1 U14670 ( .A1(n11916), .A2(n14611), .ZN(n14610) );
  INV_X1 U14671 ( .A(n14612), .ZN(n11916) );
  NAND3_X1 U14672 ( .A1(n14613), .A2(n7877), .A3(b_11_), .ZN(n14609) );
  NAND2_X1 U14673 ( .A1(n14614), .A2(n11765), .ZN(n14608) );
  XOR2_X1 U14674 ( .A(n14611), .B(a_11_), .Z(n14614) );
  XNOR2_X1 U14675 ( .A(n14615), .B(n14616), .ZN(Result_add_10_) );
  NOR2_X1 U14676 ( .A1(n14617), .A2(n12285), .ZN(n14616) );
  XOR2_X1 U14677 ( .A(n14618), .B(n14619), .Z(Result_add_0_) );
  NOR2_X1 U14678 ( .A1(n14620), .A2(n14621), .ZN(n14619) );
  INV_X1 U14679 ( .A(n7512), .ZN(n14621) );
  NAND2_X1 U14680 ( .A1(b_0_), .A2(a_0_), .ZN(n7512) );
  NOR2_X1 U14681 ( .A1(b_0_), .A2(a_0_), .ZN(n14620) );
  NOR2_X1 U14682 ( .A1(n14567), .A2(n14622), .ZN(n14618) );
  NOR2_X1 U14683 ( .A1(n14152), .A2(n14566), .ZN(n14622) );
  INV_X1 U14684 ( .A(n14569), .ZN(n14566) );
  NOR2_X1 U14685 ( .A1(n13922), .A2(n14623), .ZN(n14569) );
  NOR2_X1 U14686 ( .A1(n14515), .A2(n14513), .ZN(n14623) );
  AND2_X1 U14687 ( .A1(n14505), .A2(n14624), .ZN(n14513) );
  NAND2_X1 U14688 ( .A1(n14625), .A2(n14504), .ZN(n14624) );
  INV_X1 U14689 ( .A(n14506), .ZN(n14504) );
  NOR2_X1 U14690 ( .A1(n13669), .A2(n14626), .ZN(n14506) );
  NOR2_X1 U14691 ( .A1(n14500), .A2(n14498), .ZN(n14626) );
  AND2_X1 U14692 ( .A1(n14495), .A2(n14627), .ZN(n14498) );
  NAND2_X1 U14693 ( .A1(n14628), .A2(n14494), .ZN(n14627) );
  INV_X1 U14694 ( .A(n14496), .ZN(n14494) );
  NOR2_X1 U14695 ( .A1(n13209), .A2(n14629), .ZN(n14496) );
  NOR2_X1 U14696 ( .A1(n14490), .A2(n14488), .ZN(n14629) );
  AND2_X1 U14697 ( .A1(n14486), .A2(n14630), .ZN(n14488) );
  NAND2_X1 U14698 ( .A1(n14631), .A2(n14485), .ZN(n14630) );
  NAND2_X1 U14699 ( .A1(n12748), .A2(n14632), .ZN(n14485) );
  NAND2_X1 U14700 ( .A1(n14481), .A2(n14479), .ZN(n14632) );
  NAND2_X1 U14701 ( .A1(n14476), .A2(n14633), .ZN(n14479) );
  NAND2_X1 U14702 ( .A1(n14634), .A2(n14475), .ZN(n14633) );
  INV_X1 U14703 ( .A(n14477), .ZN(n14475) );
  NOR2_X1 U14704 ( .A1(n12285), .A2(n14635), .ZN(n14477) );
  NOR2_X1 U14705 ( .A1(n14617), .A2(n14615), .ZN(n14635) );
  AND2_X1 U14706 ( .A1(n14612), .A2(n14636), .ZN(n14615) );
  NAND2_X1 U14707 ( .A1(n14637), .A2(n14611), .ZN(n14636) );
  INV_X1 U14708 ( .A(n14613), .ZN(n14611) );
  NOR2_X1 U14709 ( .A1(n11824), .A2(n14638), .ZN(n14613) );
  NOR2_X1 U14710 ( .A1(n14607), .A2(n14605), .ZN(n14638) );
  AND2_X1 U14711 ( .A1(n14602), .A2(n14639), .ZN(n14605) );
  NAND2_X1 U14712 ( .A1(n14640), .A2(n14601), .ZN(n14639) );
  INV_X1 U14713 ( .A(n14603), .ZN(n14601) );
  NOR2_X1 U14714 ( .A1(n11370), .A2(n14641), .ZN(n14603) );
  NOR2_X1 U14715 ( .A1(n14597), .A2(n14595), .ZN(n14641) );
  NOR2_X1 U14716 ( .A1(n11150), .A2(n14642), .ZN(n14595) );
  AND2_X1 U14717 ( .A1(n14643), .A2(n14592), .ZN(n14642) );
  INV_X1 U14718 ( .A(n14593), .ZN(n14592) );
  NOR2_X1 U14719 ( .A1(n10910), .A2(n14644), .ZN(n14593) );
  NOR2_X1 U14720 ( .A1(n14588), .A2(n14586), .ZN(n14644) );
  AND2_X1 U14721 ( .A1(n14583), .A2(n14645), .ZN(n14586) );
  NAND2_X1 U14722 ( .A1(n14646), .A2(n14582), .ZN(n14645) );
  INV_X1 U14723 ( .A(n14584), .ZN(n14582) );
  NOR2_X1 U14724 ( .A1(n10460), .A2(n14647), .ZN(n14584) );
  NOR2_X1 U14725 ( .A1(n14578), .A2(n14576), .ZN(n14647) );
  AND2_X1 U14726 ( .A1(n14574), .A2(n14648), .ZN(n14576) );
  NAND2_X1 U14727 ( .A1(n14649), .A2(n14573), .ZN(n14648) );
  NAND2_X1 U14728 ( .A1(n10163), .A2(n14650), .ZN(n14573) );
  NAND2_X1 U14729 ( .A1(n14562), .A2(n14560), .ZN(n14650) );
  NAND2_X1 U14730 ( .A1(n14557), .A2(n14651), .ZN(n14560) );
  NAND2_X1 U14731 ( .A1(n14652), .A2(n14556), .ZN(n14651) );
  INV_X1 U14732 ( .A(n14558), .ZN(n14556) );
  NOR2_X1 U14733 ( .A1(n9561), .A2(n14653), .ZN(n14558) );
  NOR2_X1 U14734 ( .A1(n14552), .A2(n14550), .ZN(n14653) );
  NOR2_X1 U14735 ( .A1(n9332), .A2(n14654), .ZN(n14550) );
  AND2_X1 U14736 ( .A1(n14655), .A2(n14547), .ZN(n14654) );
  INV_X1 U14737 ( .A(n14548), .ZN(n14547) );
  NOR2_X1 U14738 ( .A1(n9087), .A2(n14656), .ZN(n14548) );
  NOR2_X1 U14739 ( .A1(n14543), .A2(n14541), .ZN(n14656) );
  AND2_X1 U14740 ( .A1(n14539), .A2(n14657), .ZN(n14541) );
  NAND2_X1 U14741 ( .A1(n14658), .A2(n14538), .ZN(n14657) );
  NAND2_X1 U14742 ( .A1(n8827), .A2(n14659), .ZN(n14538) );
  NAND2_X1 U14743 ( .A1(n14534), .A2(n14532), .ZN(n14659) );
  NAND2_X1 U14744 ( .A1(n14530), .A2(n14660), .ZN(n14532) );
  NAND2_X1 U14745 ( .A1(n14661), .A2(n14529), .ZN(n14660) );
  NAND2_X1 U14746 ( .A1(n8169), .A2(n14662), .ZN(n14529) );
  NAND2_X1 U14747 ( .A1(n14525), .A2(n14524), .ZN(n14662) );
  NAND2_X1 U14748 ( .A1(n14520), .A2(n14663), .ZN(n14524) );
  NAND2_X1 U14749 ( .A1(n14664), .A2(n14519), .ZN(n14663) );
  NAND2_X1 U14750 ( .A1(n14510), .A2(n14665), .ZN(n14519) );
  NAND2_X1 U14751 ( .A1(Result_mul_63_), .A2(n14666), .ZN(n14665) );
  NAND2_X1 U14752 ( .A1(n7274), .A2(n14287), .ZN(n14666) );
  INV_X1 U14753 ( .A(a_30_), .ZN(n14287) );
  INV_X1 U14754 ( .A(n14512), .ZN(Result_mul_63_) );
  NAND2_X1 U14755 ( .A1(b_31_), .A2(a_31_), .ZN(n14512) );
  NAND2_X1 U14756 ( .A1(b_30_), .A2(a_30_), .ZN(n14510) );
  NAND2_X1 U14757 ( .A1(n7725), .A2(n7946), .ZN(n14664) );
  INV_X1 U14758 ( .A(b_29_), .ZN(n7725) );
  NAND2_X1 U14759 ( .A1(b_29_), .A2(a_29_), .ZN(n14520) );
  NAND2_X1 U14760 ( .A1(n7953), .A2(n14471), .ZN(n14525) );
  INV_X1 U14761 ( .A(a_28_), .ZN(n14471) );
  INV_X1 U14762 ( .A(b_28_), .ZN(n7953) );
  NAND2_X1 U14763 ( .A1(b_28_), .A2(a_28_), .ZN(n8169) );
  NAND2_X1 U14764 ( .A1(n8183), .A2(n14267), .ZN(n14661) );
  INV_X1 U14765 ( .A(a_27_), .ZN(n14267) );
  NAND2_X1 U14766 ( .A1(b_27_), .A2(a_27_), .ZN(n14530) );
  NAND2_X1 U14767 ( .A1(n8403), .A2(n7295), .ZN(n14534) );
  INV_X1 U14768 ( .A(a_26_), .ZN(n7295) );
  INV_X1 U14769 ( .A(b_26_), .ZN(n8403) );
  NAND2_X1 U14770 ( .A1(b_26_), .A2(a_26_), .ZN(n8827) );
  NAND2_X1 U14771 ( .A1(n8639), .A2(n7923), .ZN(n14658) );
  INV_X1 U14772 ( .A(b_25_), .ZN(n8639) );
  NAND2_X1 U14773 ( .A1(b_25_), .A2(a_25_), .ZN(n14539) );
  NOR2_X1 U14774 ( .A1(b_24_), .A2(a_24_), .ZN(n14543) );
  NOR2_X1 U14775 ( .A1(n8848), .A2(n7691), .ZN(n9087) );
  INV_X1 U14776 ( .A(b_24_), .ZN(n8848) );
  NAND2_X1 U14777 ( .A1(n9071), .A2(n7916), .ZN(n14655) );
  NOR2_X1 U14778 ( .A1(n9071), .A2(n7916), .ZN(n9332) );
  INV_X1 U14779 ( .A(b_23_), .ZN(n9071) );
  NOR2_X1 U14780 ( .A1(b_22_), .A2(a_22_), .ZN(n14552) );
  NOR2_X1 U14781 ( .A1(n9312), .A2(n7312), .ZN(n9561) );
  INV_X1 U14782 ( .A(a_22_), .ZN(n7312) );
  NAND2_X1 U14783 ( .A1(n9537), .A2(n7909), .ZN(n14652) );
  INV_X1 U14784 ( .A(b_21_), .ZN(n9537) );
  NAND2_X1 U14785 ( .A1(b_21_), .A2(a_21_), .ZN(n14557) );
  NAND2_X1 U14786 ( .A1(n9746), .A2(n7987), .ZN(n14562) );
  INV_X1 U14787 ( .A(b_20_), .ZN(n9746) );
  NAND2_X1 U14788 ( .A1(b_20_), .A2(a_20_), .ZN(n10163) );
  NAND2_X1 U14789 ( .A1(n9964), .A2(n7902), .ZN(n14649) );
  INV_X1 U14790 ( .A(a_19_), .ZN(n7902) );
  INV_X1 U14791 ( .A(b_19_), .ZN(n9964) );
  NAND2_X1 U14792 ( .A1(b_19_), .A2(a_19_), .ZN(n14574) );
  NOR2_X1 U14793 ( .A1(b_18_), .A2(a_18_), .ZN(n14578) );
  NOR2_X1 U14794 ( .A1(n10207), .A2(n7764), .ZN(n10460) );
  INV_X1 U14795 ( .A(b_18_), .ZN(n10207) );
  NAND2_X1 U14796 ( .A1(n10420), .A2(n7337), .ZN(n14646) );
  INV_X1 U14797 ( .A(b_17_), .ZN(n10420) );
  NAND2_X1 U14798 ( .A1(b_17_), .A2(a_17_), .ZN(n14583) );
  NOR2_X1 U14799 ( .A1(b_16_), .A2(a_16_), .ZN(n14588) );
  NOR2_X1 U14800 ( .A1(n10683), .A2(n7773), .ZN(n10910) );
  INV_X1 U14801 ( .A(a_16_), .ZN(n7773) );
  NAND2_X1 U14802 ( .A1(n10863), .A2(n7346), .ZN(n14643) );
  NOR2_X1 U14803 ( .A1(n10863), .A2(n7346), .ZN(n11150) );
  INV_X1 U14804 ( .A(b_15_), .ZN(n10863) );
  NOR2_X1 U14805 ( .A1(b_14_), .A2(a_14_), .ZN(n14597) );
  NOR2_X1 U14806 ( .A1(n11103), .A2(n7782), .ZN(n11370) );
  INV_X1 U14807 ( .A(a_14_), .ZN(n7782) );
  INV_X1 U14808 ( .A(b_14_), .ZN(n11103) );
  NAND2_X1 U14809 ( .A1(n11322), .A2(n7355), .ZN(n14640) );
  INV_X1 U14810 ( .A(a_13_), .ZN(n7355) );
  INV_X1 U14811 ( .A(b_13_), .ZN(n11322) );
  NAND2_X1 U14812 ( .A1(b_13_), .A2(a_13_), .ZN(n14602) );
  NOR2_X1 U14813 ( .A1(b_12_), .A2(a_12_), .ZN(n14607) );
  NOR2_X1 U14814 ( .A1(n11559), .A2(n8020), .ZN(n11824) );
  INV_X1 U14815 ( .A(a_12_), .ZN(n8020) );
  INV_X1 U14816 ( .A(b_12_), .ZN(n11559) );
  NAND2_X1 U14817 ( .A1(n11765), .A2(n7877), .ZN(n14637) );
  INV_X1 U14818 ( .A(a_11_), .ZN(n7877) );
  INV_X1 U14819 ( .A(b_11_), .ZN(n11765) );
  NAND2_X1 U14820 ( .A1(b_11_), .A2(a_11_), .ZN(n14612) );
  NOR2_X1 U14821 ( .A1(b_10_), .A2(a_10_), .ZN(n14617) );
  NOR2_X1 U14822 ( .A1(n12010), .A2(n7799), .ZN(n12285) );
  INV_X1 U14823 ( .A(a_10_), .ZN(n7799) );
  INV_X1 U14824 ( .A(b_10_), .ZN(n12010) );
  NAND2_X1 U14825 ( .A1(n12224), .A2(n7870), .ZN(n14634) );
  INV_X1 U14826 ( .A(b_9_), .ZN(n12224) );
  NAND2_X1 U14827 ( .A1(a_9_), .A2(b_9_), .ZN(n14476) );
  NAND2_X1 U14828 ( .A1(n12466), .A2(n8037), .ZN(n14481) );
  INV_X1 U14829 ( .A(a_8_), .ZN(n8037) );
  INV_X1 U14830 ( .A(b_8_), .ZN(n12466) );
  NAND2_X1 U14831 ( .A1(a_8_), .A2(b_8_), .ZN(n12748) );
  NAND2_X1 U14832 ( .A1(n12673), .A2(n7863), .ZN(n14631) );
  INV_X1 U14833 ( .A(a_7_), .ZN(n7863) );
  NAND2_X1 U14834 ( .A1(a_7_), .A2(b_7_), .ZN(n14486) );
  NOR2_X1 U14835 ( .A1(b_6_), .A2(a_6_), .ZN(n14490) );
  NOR2_X1 U14836 ( .A1(n7388), .A2(n12904), .ZN(n13209) );
  INV_X1 U14837 ( .A(b_6_), .ZN(n12904) );
  INV_X1 U14838 ( .A(a_6_), .ZN(n7388) );
  NAND2_X1 U14839 ( .A1(n13129), .A2(n7393), .ZN(n14628) );
  INV_X1 U14840 ( .A(a_5_), .ZN(n7393) );
  INV_X1 U14841 ( .A(b_5_), .ZN(n13129) );
  NAND2_X1 U14842 ( .A1(a_5_), .A2(b_5_), .ZN(n14495) );
  NOR2_X1 U14843 ( .A1(b_4_), .A2(a_4_), .ZN(n14500) );
  NOR2_X1 U14844 ( .A1(n7398), .A2(n13352), .ZN(n13669) );
  INV_X1 U14845 ( .A(b_4_), .ZN(n13352) );
  INV_X1 U14846 ( .A(a_4_), .ZN(n7398) );
  NAND2_X1 U14847 ( .A1(n13581), .A2(n7850), .ZN(n14625) );
  INV_X1 U14848 ( .A(a_3_), .ZN(n7850) );
  INV_X1 U14849 ( .A(b_3_), .ZN(n13581) );
  NAND2_X1 U14850 ( .A1(a_3_), .A2(b_3_), .ZN(n14505) );
  NOR2_X1 U14851 ( .A1(b_2_), .A2(a_2_), .ZN(n14515) );
  NOR2_X1 U14852 ( .A1(n7832), .A2(n13794), .ZN(n13922) );
  INV_X1 U14853 ( .A(b_2_), .ZN(n13794) );
  INV_X1 U14854 ( .A(a_2_), .ZN(n7832) );
  NOR2_X1 U14855 ( .A1(n7411), .A2(n14083), .ZN(n14152) );
  INV_X1 U14856 ( .A(b_1_), .ZN(n14083) );
  INV_X1 U14857 ( .A(a_1_), .ZN(n7411) );
  NOR2_X1 U14858 ( .A1(b_1_), .A2(a_1_), .ZN(n14567) );
endmodule

