module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, N421, N430, N431, N432 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92, N95, N99, N102, N105, N108, N112, N115;
output N223, N329, N370, N421, N430, N431, N432;
wire new_n595_, new_n614_, new_n445_, new_n699_, new_n236_, new_n238_, new_n479_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n738_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n670_, new_n456_, new_n691_, new_n170_, new_n246_, new_n682_, new_n812_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n853_, new_n602_, new_n114_, new_n188_, new_n240_, new_n660_, new_n413_, new_n695_, new_n526_, new_n442_, new_n677_, new_n642_, new_n211_, new_n123_, new_n127_, new_n342_, new_n552_, new_n649_, new_n678_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n500_, new_n786_, new_n799_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n580_, new_n484_, new_n832_, new_n766_, new_n272_, new_n282_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n110_, new_n315_, new_n685_, new_n124_, new_n326_, new_n554_, new_n648_, new_n164_, new_n230_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n849_, new_n855_, new_n606_, new_n589_, new_n796_, new_n248_, new_n350_, new_n117_, new_n655_, new_n630_, new_n759_, new_n167_, new_n385_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n297_, new_n361_, new_n565_, new_n764_, new_n150_, new_n683_, new_n108_, new_n137_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n530_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n158_, new_n763_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n271_, new_n674_, new_n274_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n650_, new_n708_, new_n750_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n506_, new_n680_, new_n256_, new_n778_, new_n452_, new_n381_, new_n656_, new_n820_, new_n771_, new_n388_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n657_, new_n652_, new_n314_, new_n582_, new_n118_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n346_, new_n396_, new_n198_, new_n438_, new_n696_, new_n208_, new_n632_, new_n671_, new_n528_, new_n179_, new_n572_, new_n850_, new_n436_, new_n397_, new_n729_, new_n399_, new_n596_, new_n870_, new_n805_, new_n559_, new_n762_, new_n838_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n295_, new_n359_, new_n132_, new_n794_, new_n628_, new_n166_, new_n162_, new_n745_, new_n457_, new_n161_, new_n553_, new_n668_, new_n333_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n276_, new_n688_, new_n155_, new_n384_, new_n410_, new_n851_, new_n543_, new_n113_, new_n775_, new_n371_, new_n509_, new_n454_, new_n202_, new_n296_, new_n661_, new_n308_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n259_, new_n362_, new_n654_, new_n713_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n130_, new_n505_, new_n619_, new_n471_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n352_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n126_, new_n810_, new_n808_, new_n177_, new_n493_, new_n547_, new_n264_, new_n665_, new_n800_, new_n379_, new_n719_, new_n869_, new_n273_, new_n586_, new_n270_, new_n570_, new_n598_, new_n824_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n302_, new_n191_, new_n755_, new_n225_, new_n387_, new_n544_, new_n476_, new_n615_, new_n722_, new_n112_, new_n856_, new_n121_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n737_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n631_, new_n453_, new_n516_, new_n163_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n440_, new_n733_, new_n122_, new_n531_, new_n593_, new_n111_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n115_, new_n307_, new_n852_, new_n190_, new_n597_, new_n408_, new_n470_, new_n213_, new_n134_, new_n769_, new_n651_, new_n433_, new_n871_, new_n435_, new_n109_, new_n776_, new_n265_, new_n732_, new_n687_, new_n370_, new_n689_, new_n584_, new_n815_, new_n278_, new_n304_, new_n523_, new_n638_, new_n712_, new_n550_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n129_, new_n711_, new_n644_, new_n731_, new_n599_, new_n412_, new_n607_, new_n645_, new_n327_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n818_, new_n574_, new_n319_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n754_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n803_, new_n330_, new_n727_, new_n375_, new_n294_, new_n760_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n357_, new_n320_, new_n780_, new_n245_, new_n643_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n560_, new_n865_, new_n128_, new_n358_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n425_, new_n175_, new_n226_, new_n802_, new_n697_, new_n185_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n434_, new_n200_, new_n422_, new_n581_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n686_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n120_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n356_, new_n647_, new_n229_, new_n536_, new_n464_, new_n204_, new_n181_, new_n135_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n108_, N56 );
and g001 ( new_n109_, keyIn_0_4, N50 );
not g002 ( new_n110_, new_n109_ );
or g003 ( new_n111_, keyIn_0_4, N50 );
and g004 ( new_n112_, new_n110_, new_n111_ );
or g005 ( new_n113_, new_n112_, new_n108_ );
and g006 ( new_n114_, new_n113_, keyIn_0_10 );
not g007 ( new_n115_, new_n114_ );
or g008 ( new_n116_, new_n113_, keyIn_0_10 );
and g009 ( new_n117_, new_n115_, new_n116_ );
not g010 ( new_n118_, new_n117_ );
or g011 ( new_n119_, keyIn_0_1, N24 );
not g012 ( new_n120_, new_n119_ );
not g013 ( new_n121_, N30 );
and g014 ( new_n122_, keyIn_0_1, N24 );
or g015 ( new_n123_, new_n122_, new_n121_ );
or g016 ( new_n124_, new_n123_, new_n120_ );
or g017 ( new_n125_, new_n124_, keyIn_0_8 );
and g018 ( new_n126_, new_n124_, keyIn_0_8 );
not g019 ( new_n127_, new_n126_ );
and g020 ( new_n128_, new_n127_, new_n125_ );
or g021 ( new_n129_, keyIn_0_2, N37 );
not g022 ( new_n130_, new_n129_ );
not g023 ( new_n131_, N43 );
and g024 ( new_n132_, keyIn_0_2, N37 );
or g025 ( new_n133_, new_n132_, new_n131_ );
or g026 ( new_n134_, new_n133_, new_n130_ );
or g027 ( new_n135_, new_n134_, keyIn_0_9 );
not g028 ( new_n136_, keyIn_0_9 );
not g029 ( new_n137_, new_n132_ );
and g030 ( new_n138_, new_n137_, N43 );
and g031 ( new_n139_, new_n138_, new_n129_ );
or g032 ( new_n140_, new_n139_, new_n136_ );
and g033 ( new_n141_, new_n140_, new_n135_ );
or g034 ( new_n142_, new_n128_, new_n141_ );
or g035 ( new_n143_, new_n142_, new_n118_ );
not g036 ( new_n144_, keyIn_0_13 );
not g037 ( new_n145_, keyIn_0_7 );
and g038 ( new_n146_, new_n145_, N102 );
not g039 ( new_n147_, new_n146_ );
or g040 ( new_n148_, new_n145_, N102 );
and g041 ( new_n149_, new_n148_, N108 );
and g042 ( new_n150_, new_n149_, new_n147_ );
or g043 ( new_n151_, new_n150_, new_n144_ );
not g044 ( new_n152_, N108 );
not g045 ( new_n153_, N102 );
and g046 ( new_n154_, new_n153_, keyIn_0_7 );
or g047 ( new_n155_, new_n154_, new_n152_ );
or g048 ( new_n156_, new_n155_, new_n146_ );
or g049 ( new_n157_, new_n156_, keyIn_0_13 );
and g050 ( new_n158_, new_n157_, new_n151_ );
not g051 ( new_n159_, keyIn_0_0 );
and g052 ( new_n160_, new_n159_, N1 );
not g053 ( new_n161_, new_n160_ );
or g054 ( new_n162_, new_n159_, N1 );
and g055 ( new_n163_, new_n162_, N4 );
and g056 ( new_n164_, new_n163_, new_n161_ );
not g057 ( new_n165_, N11 );
and g058 ( new_n166_, new_n165_, N17 );
not g059 ( new_n167_, N63 );
and g060 ( new_n168_, new_n167_, N69 );
or g061 ( new_n169_, new_n166_, new_n168_ );
or g062 ( new_n170_, new_n164_, new_n169_ );
or g063 ( new_n171_, new_n158_, new_n170_ );
not g064 ( new_n172_, N76 );
and g065 ( new_n173_, new_n172_, keyIn_0_5 );
not g066 ( new_n174_, keyIn_0_5 );
and g067 ( new_n175_, new_n174_, N76 );
or g068 ( new_n176_, new_n173_, new_n175_ );
and g069 ( new_n177_, new_n176_, N82 );
or g070 ( new_n178_, new_n177_, keyIn_0_11 );
not g071 ( new_n179_, keyIn_0_11 );
not g072 ( new_n180_, N82 );
or g073 ( new_n181_, new_n174_, N76 );
or g074 ( new_n182_, new_n172_, keyIn_0_5 );
and g075 ( new_n183_, new_n181_, new_n182_ );
or g076 ( new_n184_, new_n183_, new_n180_ );
or g077 ( new_n185_, new_n184_, new_n179_ );
and g078 ( new_n186_, new_n185_, new_n178_ );
not g079 ( new_n187_, keyIn_0_12 );
or g080 ( new_n188_, keyIn_0_6, N89 );
not g081 ( new_n189_, new_n188_ );
not g082 ( new_n190_, N95 );
and g083 ( new_n191_, keyIn_0_6, N89 );
or g084 ( new_n192_, new_n191_, new_n190_ );
or g085 ( new_n193_, new_n192_, new_n189_ );
or g086 ( new_n194_, new_n193_, new_n187_ );
and g087 ( new_n195_, new_n193_, new_n187_ );
not g088 ( new_n196_, new_n195_ );
and g089 ( new_n197_, new_n196_, new_n194_ );
or g090 ( new_n198_, new_n186_, new_n197_ );
or g091 ( new_n199_, new_n198_, new_n171_ );
or g092 ( new_n200_, new_n199_, new_n143_ );
or g093 ( new_n201_, new_n200_, keyIn_0_14 );
not g094 ( new_n202_, keyIn_0_14 );
not g095 ( new_n203_, new_n125_ );
or g096 ( new_n204_, new_n203_, new_n126_ );
not g097 ( new_n205_, new_n135_ );
and g098 ( new_n206_, new_n134_, keyIn_0_9 );
or g099 ( new_n207_, new_n205_, new_n206_ );
and g100 ( new_n208_, new_n204_, new_n207_ );
and g101 ( new_n209_, new_n208_, new_n117_ );
and g102 ( new_n210_, new_n156_, keyIn_0_13 );
and g103 ( new_n211_, new_n150_, new_n144_ );
or g104 ( new_n212_, new_n210_, new_n211_ );
not g105 ( new_n213_, new_n170_ );
and g106 ( new_n214_, new_n212_, new_n213_ );
and g107 ( new_n215_, new_n184_, new_n179_ );
and g108 ( new_n216_, new_n177_, keyIn_0_11 );
or g109 ( new_n217_, new_n215_, new_n216_ );
not g110 ( new_n218_, new_n194_ );
or g111 ( new_n219_, new_n218_, new_n195_ );
and g112 ( new_n220_, new_n219_, new_n217_ );
and g113 ( new_n221_, new_n220_, new_n214_ );
and g114 ( new_n222_, new_n209_, new_n221_ );
or g115 ( new_n223_, new_n222_, new_n202_ );
and g116 ( N223, new_n201_, new_n223_ );
not g117 ( new_n225_, keyIn_0_28 );
not g118 ( new_n226_, keyIn_0_24 );
not g119 ( new_n227_, keyIn_0_18 );
or g120 ( new_n228_, N223, keyIn_0_15 );
not g121 ( new_n229_, keyIn_0_15 );
and g122 ( new_n230_, new_n222_, new_n202_ );
and g123 ( new_n231_, new_n200_, keyIn_0_14 );
or g124 ( new_n232_, new_n231_, new_n230_ );
or g125 ( new_n233_, new_n232_, new_n229_ );
and g126 ( new_n234_, new_n228_, new_n233_ );
and g127 ( new_n235_, new_n234_, new_n207_ );
and g128 ( new_n236_, new_n232_, new_n229_ );
and g129 ( new_n237_, N223, keyIn_0_15 );
or g130 ( new_n238_, new_n236_, new_n237_ );
and g131 ( new_n239_, new_n238_, new_n141_ );
or g132 ( new_n240_, new_n239_, new_n235_ );
and g133 ( new_n241_, new_n240_, new_n227_ );
not g134 ( new_n242_, new_n241_ );
or g135 ( new_n243_, new_n240_, new_n227_ );
and g136 ( new_n244_, new_n242_, new_n243_ );
not g137 ( new_n245_, N47 );
and g138 ( new_n246_, new_n131_, keyIn_0_3 );
not g139 ( new_n247_, new_n246_ );
or g140 ( new_n248_, new_n131_, keyIn_0_3 );
and g141 ( new_n249_, new_n247_, new_n248_ );
and g142 ( new_n250_, new_n249_, new_n245_ );
not g143 ( new_n251_, new_n250_ );
or g144 ( new_n252_, new_n244_, new_n251_ );
and g145 ( new_n253_, new_n252_, new_n226_ );
not g146 ( new_n254_, new_n253_ );
or g147 ( new_n255_, new_n252_, new_n226_ );
and g148 ( new_n256_, new_n254_, new_n255_ );
or g149 ( new_n257_, new_n234_, new_n164_ );
not g150 ( new_n258_, new_n164_ );
or g151 ( new_n259_, new_n238_, new_n258_ );
and g152 ( new_n260_, new_n259_, new_n257_ );
or g153 ( new_n261_, new_n260_, keyIn_0_16 );
not g154 ( new_n262_, keyIn_0_16 );
and g155 ( new_n263_, new_n238_, new_n258_ );
and g156 ( new_n264_, new_n234_, new_n164_ );
or g157 ( new_n265_, new_n263_, new_n264_ );
or g158 ( new_n266_, new_n265_, new_n262_ );
and g159 ( new_n267_, new_n266_, new_n261_ );
not g160 ( new_n268_, N8 );
and g161 ( new_n269_, new_n268_, N4 );
not g162 ( new_n270_, new_n269_ );
or g163 ( new_n271_, new_n267_, new_n270_ );
and g164 ( new_n272_, new_n271_, keyIn_0_22 );
not g165 ( new_n273_, keyIn_0_22 );
and g166 ( new_n274_, new_n265_, new_n262_ );
and g167 ( new_n275_, new_n260_, keyIn_0_16 );
or g168 ( new_n276_, new_n274_, new_n275_ );
and g169 ( new_n277_, new_n276_, new_n269_ );
and g170 ( new_n278_, new_n277_, new_n273_ );
or g171 ( new_n279_, new_n272_, new_n278_ );
not g172 ( new_n280_, new_n166_ );
and g173 ( new_n281_, new_n238_, new_n280_ );
not g174 ( new_n282_, keyIn_0_17 );
and g175 ( new_n283_, new_n234_, new_n166_ );
or g176 ( new_n284_, new_n283_, new_n282_ );
or g177 ( new_n285_, new_n284_, new_n281_ );
or g178 ( new_n286_, new_n234_, new_n166_ );
or g179 ( new_n287_, new_n238_, new_n280_ );
and g180 ( new_n288_, new_n287_, new_n286_ );
or g181 ( new_n289_, new_n288_, keyIn_0_17 );
and g182 ( new_n290_, new_n289_, new_n285_ );
not g183 ( new_n291_, N21 );
and g184 ( new_n292_, new_n291_, N17 );
not g185 ( new_n293_, new_n292_ );
or g186 ( new_n294_, new_n290_, new_n293_ );
and g187 ( new_n295_, new_n294_, keyIn_0_23 );
not g188 ( new_n296_, keyIn_0_23 );
and g189 ( new_n297_, new_n287_, keyIn_0_17 );
and g190 ( new_n298_, new_n297_, new_n286_ );
or g191 ( new_n299_, new_n281_, new_n283_ );
and g192 ( new_n300_, new_n299_, new_n282_ );
or g193 ( new_n301_, new_n300_, new_n298_ );
and g194 ( new_n302_, new_n301_, new_n292_ );
and g195 ( new_n303_, new_n302_, new_n296_ );
or g196 ( new_n304_, new_n303_, new_n295_ );
and g197 ( new_n305_, new_n279_, new_n304_ );
and g198 ( new_n306_, new_n305_, new_n256_ );
not g199 ( new_n307_, keyIn_0_21 );
or g200 ( new_n308_, new_n234_, new_n212_ );
or g201 ( new_n309_, new_n238_, new_n158_ );
and g202 ( new_n310_, new_n309_, new_n308_ );
or g203 ( new_n311_, new_n310_, new_n307_ );
and g204 ( new_n312_, new_n238_, new_n158_ );
and g205 ( new_n313_, new_n234_, new_n212_ );
or g206 ( new_n314_, new_n312_, new_n313_ );
or g207 ( new_n315_, new_n314_, keyIn_0_21 );
and g208 ( new_n316_, new_n315_, new_n311_ );
not g209 ( new_n317_, N112 );
and g210 ( new_n318_, new_n317_, N108 );
not g211 ( new_n319_, new_n318_ );
or g212 ( new_n320_, new_n316_, new_n319_ );
and g213 ( new_n321_, new_n320_, keyIn_0_27 );
not g214 ( new_n322_, keyIn_0_27 );
and g215 ( new_n323_, new_n314_, keyIn_0_21 );
and g216 ( new_n324_, new_n310_, new_n307_ );
or g217 ( new_n325_, new_n323_, new_n324_ );
and g218 ( new_n326_, new_n325_, new_n318_ );
and g219 ( new_n327_, new_n326_, new_n322_ );
or g220 ( new_n328_, new_n321_, new_n327_ );
and g221 ( new_n329_, new_n234_, new_n219_ );
and g222 ( new_n330_, new_n238_, new_n197_ );
or g223 ( new_n331_, new_n330_, new_n329_ );
not g224 ( new_n332_, new_n331_ );
not g225 ( new_n333_, N99 );
and g226 ( new_n334_, new_n333_, N95 );
and g227 ( new_n335_, new_n332_, new_n334_ );
not g228 ( new_n336_, new_n335_ );
and g229 ( new_n337_, new_n234_, new_n204_ );
and g230 ( new_n338_, new_n238_, new_n128_ );
or g231 ( new_n339_, new_n338_, new_n337_ );
not g232 ( new_n340_, new_n339_ );
not g233 ( new_n341_, N34 );
and g234 ( new_n342_, new_n341_, N30 );
and g235 ( new_n343_, new_n340_, new_n342_ );
not g236 ( new_n344_, new_n343_ );
and g237 ( new_n345_, new_n234_, new_n217_ );
and g238 ( new_n346_, new_n238_, new_n186_ );
or g239 ( new_n347_, new_n346_, new_n345_ );
not g240 ( new_n348_, new_n347_ );
not g241 ( new_n349_, N86 );
and g242 ( new_n350_, new_n349_, N82 );
and g243 ( new_n351_, new_n348_, new_n350_ );
not g244 ( new_n352_, new_n351_ );
and g245 ( new_n353_, new_n344_, new_n352_ );
and g246 ( new_n354_, new_n353_, new_n336_ );
and g247 ( new_n355_, new_n328_, new_n354_ );
not g248 ( new_n356_, keyIn_0_25 );
not g249 ( new_n357_, keyIn_0_19 );
or g250 ( new_n358_, new_n234_, new_n117_ );
or g251 ( new_n359_, new_n238_, new_n118_ );
and g252 ( new_n360_, new_n359_, new_n358_ );
or g253 ( new_n361_, new_n360_, new_n357_ );
and g254 ( new_n362_, new_n238_, new_n118_ );
and g255 ( new_n363_, new_n234_, new_n117_ );
or g256 ( new_n364_, new_n362_, new_n363_ );
or g257 ( new_n365_, new_n364_, keyIn_0_19 );
and g258 ( new_n366_, new_n365_, new_n361_ );
not g259 ( new_n367_, N60 );
and g260 ( new_n368_, new_n367_, N56 );
not g261 ( new_n369_, new_n368_ );
or g262 ( new_n370_, new_n366_, new_n369_ );
and g263 ( new_n371_, new_n370_, new_n356_ );
and g264 ( new_n372_, new_n364_, keyIn_0_19 );
and g265 ( new_n373_, new_n360_, new_n357_ );
or g266 ( new_n374_, new_n372_, new_n373_ );
and g267 ( new_n375_, new_n374_, new_n368_ );
and g268 ( new_n376_, new_n375_, keyIn_0_25 );
or g269 ( new_n377_, new_n371_, new_n376_ );
or g270 ( new_n378_, new_n234_, new_n168_ );
not g271 ( new_n379_, new_n168_ );
or g272 ( new_n380_, new_n238_, new_n379_ );
and g273 ( new_n381_, new_n380_, keyIn_0_20 );
and g274 ( new_n382_, new_n381_, new_n378_ );
not g275 ( new_n383_, keyIn_0_20 );
and g276 ( new_n384_, new_n238_, new_n379_ );
and g277 ( new_n385_, new_n234_, new_n168_ );
or g278 ( new_n386_, new_n384_, new_n385_ );
and g279 ( new_n387_, new_n386_, new_n383_ );
or g280 ( new_n388_, new_n387_, new_n382_ );
not g281 ( new_n389_, N73 );
and g282 ( new_n390_, new_n389_, N69 );
and g283 ( new_n391_, new_n388_, new_n390_ );
or g284 ( new_n392_, new_n391_, keyIn_0_26 );
not g285 ( new_n393_, keyIn_0_26 );
or g286 ( new_n394_, new_n385_, new_n383_ );
or g287 ( new_n395_, new_n394_, new_n384_ );
and g288 ( new_n396_, new_n380_, new_n378_ );
or g289 ( new_n397_, new_n396_, keyIn_0_20 );
and g290 ( new_n398_, new_n397_, new_n395_ );
not g291 ( new_n399_, new_n390_ );
or g292 ( new_n400_, new_n398_, new_n399_ );
or g293 ( new_n401_, new_n400_, new_n393_ );
and g294 ( new_n402_, new_n392_, new_n401_ );
and g295 ( new_n403_, new_n377_, new_n402_ );
and g296 ( new_n404_, new_n355_, new_n403_ );
and g297 ( new_n405_, new_n404_, new_n306_ );
and g298 ( new_n406_, new_n405_, new_n225_ );
not g299 ( new_n407_, new_n406_ );
or g300 ( new_n408_, new_n405_, new_n225_ );
and g301 ( N329, new_n407_, new_n408_ );
not g302 ( new_n410_, keyIn_0_44 );
not g303 ( new_n411_, keyIn_0_41 );
not g304 ( new_n412_, keyIn_0_35 );
and g305 ( new_n413_, new_n400_, new_n393_ );
and g306 ( new_n414_, new_n391_, keyIn_0_26 );
or g307 ( new_n415_, new_n414_, new_n413_ );
or g308 ( new_n416_, N329, keyIn_0_31 );
not g309 ( new_n417_, keyIn_0_31 );
not g310 ( new_n418_, new_n255_ );
or g311 ( new_n419_, new_n418_, new_n253_ );
or g312 ( new_n420_, new_n277_, new_n273_ );
or g313 ( new_n421_, new_n271_, keyIn_0_22 );
and g314 ( new_n422_, new_n421_, new_n420_ );
or g315 ( new_n423_, new_n302_, new_n296_ );
or g316 ( new_n424_, new_n294_, keyIn_0_23 );
and g317 ( new_n425_, new_n423_, new_n424_ );
or g318 ( new_n426_, new_n422_, new_n425_ );
or g319 ( new_n427_, new_n426_, new_n419_ );
or g320 ( new_n428_, new_n326_, new_n322_ );
or g321 ( new_n429_, new_n320_, keyIn_0_27 );
and g322 ( new_n430_, new_n429_, new_n428_ );
not g323 ( new_n431_, new_n354_ );
or g324 ( new_n432_, new_n430_, new_n431_ );
or g325 ( new_n433_, new_n375_, keyIn_0_25 );
or g326 ( new_n434_, new_n370_, new_n356_ );
and g327 ( new_n435_, new_n434_, new_n433_ );
or g328 ( new_n436_, new_n415_, new_n435_ );
or g329 ( new_n437_, new_n436_, new_n432_ );
or g330 ( new_n438_, new_n437_, new_n427_ );
and g331 ( new_n439_, new_n438_, keyIn_0_28 );
or g332 ( new_n440_, new_n439_, new_n406_ );
or g333 ( new_n441_, new_n440_, new_n417_ );
and g334 ( new_n442_, new_n441_, new_n416_ );
and g335 ( new_n443_, new_n442_, new_n415_ );
and g336 ( new_n444_, new_n440_, new_n417_ );
and g337 ( new_n445_, N329, keyIn_0_31 );
or g338 ( new_n446_, new_n444_, new_n445_ );
and g339 ( new_n447_, new_n446_, new_n402_ );
or g340 ( new_n448_, new_n447_, new_n443_ );
and g341 ( new_n449_, new_n448_, new_n412_ );
not g342 ( new_n450_, new_n449_ );
or g343 ( new_n451_, new_n448_, new_n412_ );
not g344 ( new_n452_, N79 );
and g345 ( new_n453_, new_n452_, N69 );
and g346 ( new_n454_, new_n388_, new_n453_ );
not g347 ( new_n455_, new_n454_ );
and g348 ( new_n456_, new_n455_, keyIn_0_29 );
not g349 ( new_n457_, new_n456_ );
or g350 ( new_n458_, new_n455_, keyIn_0_29 );
and g351 ( new_n459_, new_n457_, new_n458_ );
and g352 ( new_n460_, new_n451_, new_n459_ );
and g353 ( new_n461_, new_n460_, new_n450_ );
not g354 ( new_n462_, new_n461_ );
and g355 ( new_n463_, new_n462_, new_n411_ );
and g356 ( new_n464_, new_n461_, keyIn_0_41 );
or g357 ( new_n465_, new_n463_, new_n464_ );
not g358 ( new_n466_, keyIn_0_32 );
and g359 ( new_n467_, new_n446_, new_n304_ );
and g360 ( new_n468_, new_n442_, new_n425_ );
or g361 ( new_n469_, new_n467_, new_n468_ );
and g362 ( new_n470_, new_n469_, new_n466_ );
or g363 ( new_n471_, new_n442_, new_n425_ );
or g364 ( new_n472_, new_n446_, new_n304_ );
and g365 ( new_n473_, new_n472_, new_n471_ );
and g366 ( new_n474_, new_n473_, keyIn_0_32 );
not g367 ( new_n475_, N27 );
and g368 ( new_n476_, new_n475_, N17 );
and g369 ( new_n477_, new_n301_, new_n476_ );
not g370 ( new_n478_, new_n477_ );
or g371 ( new_n479_, new_n474_, new_n478_ );
or g372 ( new_n480_, new_n479_, new_n470_ );
and g373 ( new_n481_, new_n480_, keyIn_0_38 );
not g374 ( new_n482_, keyIn_0_38 );
not g375 ( new_n483_, new_n470_ );
or g376 ( new_n484_, new_n469_, new_n466_ );
and g377 ( new_n485_, new_n484_, new_n477_ );
and g378 ( new_n486_, new_n485_, new_n483_ );
and g379 ( new_n487_, new_n486_, new_n482_ );
or g380 ( new_n488_, new_n481_, new_n487_ );
or g381 ( new_n489_, new_n446_, new_n377_ );
or g382 ( new_n490_, new_n442_, new_n435_ );
and g383 ( new_n491_, new_n489_, new_n490_ );
and g384 ( new_n492_, new_n491_, keyIn_0_34 );
not g385 ( new_n493_, new_n492_ );
or g386 ( new_n494_, new_n491_, keyIn_0_34 );
not g387 ( new_n495_, N66 );
and g388 ( new_n496_, new_n495_, N56 );
and g389 ( new_n497_, new_n374_, new_n496_ );
and g390 ( new_n498_, new_n494_, new_n497_ );
and g391 ( new_n499_, new_n498_, new_n493_ );
or g392 ( new_n500_, new_n499_, keyIn_0_40 );
and g393 ( new_n501_, new_n497_, keyIn_0_40 );
and g394 ( new_n502_, new_n493_, new_n501_ );
and g395 ( new_n503_, new_n502_, new_n494_ );
not g396 ( new_n504_, new_n503_ );
and g397 ( new_n505_, new_n500_, new_n504_ );
not g398 ( new_n506_, new_n505_ );
and g399 ( new_n507_, new_n506_, new_n488_ );
and g400 ( new_n508_, new_n507_, new_n465_ );
not g401 ( new_n509_, keyIn_0_43 );
not g402 ( new_n510_, keyIn_0_37 );
or g403 ( new_n511_, new_n442_, new_n430_ );
or g404 ( new_n512_, new_n446_, new_n328_ );
and g405 ( new_n513_, new_n512_, new_n511_ );
and g406 ( new_n514_, new_n513_, new_n510_ );
and g407 ( new_n515_, new_n446_, new_n328_ );
and g408 ( new_n516_, new_n442_, new_n430_ );
or g409 ( new_n517_, new_n515_, new_n516_ );
and g410 ( new_n518_, new_n517_, keyIn_0_37 );
not g411 ( new_n519_, N115 );
and g412 ( new_n520_, new_n519_, N108 );
and g413 ( new_n521_, new_n325_, new_n520_ );
not g414 ( new_n522_, new_n521_ );
and g415 ( new_n523_, new_n522_, keyIn_0_30 );
not g416 ( new_n524_, new_n523_ );
or g417 ( new_n525_, new_n522_, keyIn_0_30 );
and g418 ( new_n526_, new_n524_, new_n525_ );
or g419 ( new_n527_, new_n518_, new_n526_ );
or g420 ( new_n528_, new_n527_, new_n514_ );
and g421 ( new_n529_, new_n528_, new_n509_ );
not g422 ( new_n530_, new_n529_ );
or g423 ( new_n531_, new_n446_, new_n344_ );
or g424 ( new_n532_, new_n442_, new_n343_ );
and g425 ( new_n533_, new_n531_, new_n532_ );
and g426 ( new_n534_, new_n533_, keyIn_0_33 );
not g427 ( new_n535_, new_n534_ );
or g428 ( new_n536_, new_n533_, keyIn_0_33 );
not g429 ( new_n537_, N40 );
and g430 ( new_n538_, new_n537_, N30 );
and g431 ( new_n539_, new_n340_, new_n538_ );
and g432 ( new_n540_, new_n536_, new_n539_ );
and g433 ( new_n541_, new_n540_, new_n535_ );
and g434 ( new_n542_, new_n541_, keyIn_0_39 );
not g435 ( new_n543_, new_n542_ );
not g436 ( new_n544_, new_n514_ );
or g437 ( new_n545_, new_n513_, new_n510_ );
not g438 ( new_n546_, new_n526_ );
and g439 ( new_n547_, new_n545_, new_n546_ );
and g440 ( new_n548_, new_n547_, new_n544_ );
and g441 ( new_n549_, new_n548_, keyIn_0_43 );
not g442 ( new_n550_, new_n549_ );
and g443 ( new_n551_, new_n543_, new_n550_ );
and g444 ( new_n552_, new_n551_, new_n530_ );
not g445 ( new_n553_, keyIn_0_42 );
not g446 ( new_n554_, keyIn_0_36 );
or g447 ( new_n555_, new_n446_, new_n336_ );
or g448 ( new_n556_, new_n442_, new_n335_ );
and g449 ( new_n557_, new_n555_, new_n556_ );
and g450 ( new_n558_, new_n557_, new_n554_ );
not g451 ( new_n559_, new_n558_ );
or g452 ( new_n560_, new_n557_, new_n554_ );
not g453 ( new_n561_, N105 );
and g454 ( new_n562_, new_n561_, N95 );
and g455 ( new_n563_, new_n332_, new_n562_ );
and g456 ( new_n564_, new_n560_, new_n563_ );
and g457 ( new_n565_, new_n564_, new_n559_ );
or g458 ( new_n566_, new_n565_, new_n553_ );
and g459 ( new_n567_, new_n442_, new_n351_ );
not g460 ( new_n568_, new_n567_ );
and g461 ( new_n569_, new_n446_, new_n352_ );
not g462 ( new_n570_, new_n569_ );
not g463 ( new_n571_, N92 );
and g464 ( new_n572_, new_n571_, N82 );
and g465 ( new_n573_, new_n348_, new_n572_ );
and g466 ( new_n574_, new_n570_, new_n573_ );
and g467 ( new_n575_, new_n574_, new_n568_ );
and g468 ( new_n576_, new_n442_, new_n422_ );
not g469 ( new_n577_, new_n576_ );
and g470 ( new_n578_, new_n446_, new_n279_ );
not g471 ( new_n579_, new_n578_ );
not g472 ( new_n580_, N14 );
and g473 ( new_n581_, new_n580_, N4 );
and g474 ( new_n582_, new_n276_, new_n581_ );
and g475 ( new_n583_, new_n579_, new_n582_ );
and g476 ( new_n584_, new_n583_, new_n577_ );
and g477 ( new_n585_, new_n442_, new_n419_ );
not g478 ( new_n586_, new_n585_ );
and g479 ( new_n587_, new_n446_, new_n256_ );
not g480 ( new_n588_, new_n587_ );
not g481 ( new_n589_, new_n244_ );
not g482 ( new_n590_, N53 );
and g483 ( new_n591_, new_n249_, new_n590_ );
and g484 ( new_n592_, new_n589_, new_n591_ );
and g485 ( new_n593_, new_n588_, new_n592_ );
and g486 ( new_n594_, new_n593_, new_n586_ );
or g487 ( new_n595_, new_n584_, new_n594_ );
or g488 ( new_n596_, new_n595_, new_n575_ );
not g489 ( new_n597_, new_n596_ );
and g490 ( new_n598_, new_n566_, new_n597_ );
or g491 ( new_n599_, new_n541_, keyIn_0_39 );
and g492 ( new_n600_, new_n565_, new_n553_ );
not g493 ( new_n601_, new_n600_ );
and g494 ( new_n602_, new_n601_, new_n599_ );
and g495 ( new_n603_, new_n602_, new_n598_ );
and g496 ( new_n604_, new_n552_, new_n603_ );
and g497 ( new_n605_, new_n508_, new_n604_ );
and g498 ( new_n606_, new_n605_, new_n410_ );
not g499 ( new_n607_, new_n465_ );
or g500 ( new_n608_, new_n486_, new_n482_ );
or g501 ( new_n609_, new_n480_, keyIn_0_38 );
and g502 ( new_n610_, new_n609_, new_n608_ );
or g503 ( new_n611_, new_n610_, new_n505_ );
or g504 ( new_n612_, new_n611_, new_n607_ );
or g505 ( new_n613_, new_n542_, new_n549_ );
or g506 ( new_n614_, new_n613_, new_n529_ );
and g507 ( new_n615_, new_n442_, new_n335_ );
and g508 ( new_n616_, new_n446_, new_n336_ );
or g509 ( new_n617_, new_n616_, new_n615_ );
and g510 ( new_n618_, new_n617_, keyIn_0_36 );
not g511 ( new_n619_, new_n563_ );
or g512 ( new_n620_, new_n618_, new_n619_ );
or g513 ( new_n621_, new_n620_, new_n558_ );
and g514 ( new_n622_, new_n621_, keyIn_0_42 );
or g515 ( new_n623_, new_n622_, new_n596_ );
not g516 ( new_n624_, keyIn_0_39 );
not g517 ( new_n625_, keyIn_0_33 );
and g518 ( new_n626_, new_n442_, new_n343_ );
and g519 ( new_n627_, new_n446_, new_n344_ );
or g520 ( new_n628_, new_n627_, new_n626_ );
and g521 ( new_n629_, new_n628_, new_n625_ );
not g522 ( new_n630_, new_n539_ );
or g523 ( new_n631_, new_n629_, new_n630_ );
or g524 ( new_n632_, new_n631_, new_n534_ );
and g525 ( new_n633_, new_n632_, new_n624_ );
or g526 ( new_n634_, new_n633_, new_n600_ );
or g527 ( new_n635_, new_n623_, new_n634_ );
or g528 ( new_n636_, new_n635_, new_n614_ );
or g529 ( new_n637_, new_n636_, new_n612_ );
and g530 ( new_n638_, new_n637_, keyIn_0_44 );
or g531 ( N370, new_n638_, new_n606_ );
not g532 ( new_n640_, keyIn_0_58 );
or g533 ( new_n641_, new_n637_, keyIn_0_44 );
or g534 ( new_n642_, new_n605_, new_n410_ );
and g535 ( new_n643_, new_n641_, new_n642_ );
or g536 ( new_n644_, new_n643_, keyIn_0_45 );
not g537 ( new_n645_, keyIn_0_45 );
or g538 ( new_n646_, N370, new_n645_ );
and g539 ( new_n647_, new_n644_, new_n646_ );
and g540 ( new_n648_, new_n647_, N14 );
and g541 ( new_n649_, N329, N8 );
not g542 ( new_n650_, N4 );
and g543 ( new_n651_, N223, N1 );
or g544 ( new_n652_, new_n651_, new_n650_ );
or g545 ( new_n653_, new_n649_, new_n652_ );
or g546 ( new_n654_, new_n648_, new_n653_ );
and g547 ( new_n655_, N370, new_n645_ );
and g548 ( new_n656_, new_n643_, keyIn_0_45 );
or g549 ( new_n657_, new_n655_, new_n656_ );
or g550 ( new_n658_, new_n657_, new_n590_ );
or g551 ( new_n659_, new_n658_, keyIn_0_48 );
not g552 ( new_n660_, keyIn_0_48 );
and g553 ( new_n661_, new_n647_, N53 );
or g554 ( new_n662_, new_n661_, new_n660_ );
and g555 ( new_n663_, new_n659_, new_n662_ );
and g556 ( new_n664_, N329, N47 );
and g557 ( new_n665_, N223, N37 );
or g558 ( new_n666_, new_n665_, new_n131_ );
or g559 ( new_n667_, new_n664_, new_n666_ );
or g560 ( new_n668_, new_n663_, new_n667_ );
and g561 ( new_n669_, new_n668_, keyIn_0_53 );
not g562 ( new_n670_, keyIn_0_53 );
and g563 ( new_n671_, new_n661_, new_n660_ );
and g564 ( new_n672_, new_n658_, keyIn_0_48 );
or g565 ( new_n673_, new_n672_, new_n671_ );
not g566 ( new_n674_, new_n667_ );
and g567 ( new_n675_, new_n673_, new_n674_ );
and g568 ( new_n676_, new_n675_, new_n670_ );
or g569 ( new_n677_, new_n669_, new_n676_ );
and g570 ( new_n678_, new_n647_, N66 );
and g571 ( new_n679_, new_n678_, keyIn_0_49 );
not g572 ( new_n680_, new_n679_ );
or g573 ( new_n681_, new_n678_, keyIn_0_49 );
and g574 ( new_n682_, N329, N60 );
and g575 ( new_n683_, N223, N50 );
or g576 ( new_n684_, new_n683_, new_n108_ );
or g577 ( new_n685_, new_n682_, new_n684_ );
not g578 ( new_n686_, new_n685_ );
and g579 ( new_n687_, new_n681_, new_n686_ );
and g580 ( new_n688_, new_n687_, new_n680_ );
or g581 ( new_n689_, new_n688_, keyIn_0_54 );
not g582 ( new_n690_, new_n689_ );
and g583 ( new_n691_, new_n688_, keyIn_0_54 );
or g584 ( new_n692_, new_n690_, new_n691_ );
and g585 ( new_n693_, new_n692_, new_n677_ );
not g586 ( new_n694_, new_n693_ );
not g587 ( new_n695_, keyIn_0_46 );
or g588 ( new_n696_, new_n657_, new_n475_ );
and g589 ( new_n697_, new_n696_, new_n695_ );
and g590 ( new_n698_, new_n647_, N27 );
and g591 ( new_n699_, new_n698_, keyIn_0_46 );
and g592 ( new_n700_, N329, N21 );
not g593 ( new_n701_, new_n700_ );
and g594 ( new_n702_, N223, N11 );
not g595 ( new_n703_, new_n702_ );
and g596 ( new_n704_, new_n703_, N17 );
and g597 ( new_n705_, new_n701_, new_n704_ );
not g598 ( new_n706_, new_n705_ );
or g599 ( new_n707_, new_n699_, new_n706_ );
or g600 ( new_n708_, new_n707_, new_n697_ );
or g601 ( new_n709_, new_n708_, keyIn_0_51 );
not g602 ( new_n710_, keyIn_0_51 );
not g603 ( new_n711_, new_n697_ );
not g604 ( new_n712_, new_n699_ );
and g605 ( new_n713_, new_n712_, new_n705_ );
and g606 ( new_n714_, new_n713_, new_n711_ );
or g607 ( new_n715_, new_n714_, new_n710_ );
and g608 ( new_n716_, new_n715_, new_n709_ );
not g609 ( new_n717_, keyIn_0_52 );
not g610 ( new_n718_, keyIn_0_47 );
or g611 ( new_n719_, new_n657_, new_n537_ );
or g612 ( new_n720_, new_n719_, new_n718_ );
and g613 ( new_n721_, new_n647_, N40 );
or g614 ( new_n722_, new_n721_, keyIn_0_47 );
and g615 ( new_n723_, new_n720_, new_n722_ );
and g616 ( new_n724_, N329, N34 );
and g617 ( new_n725_, N223, N24 );
or g618 ( new_n726_, new_n725_, new_n121_ );
or g619 ( new_n727_, new_n724_, new_n726_ );
or g620 ( new_n728_, new_n723_, new_n727_ );
and g621 ( new_n729_, new_n728_, new_n717_ );
and g622 ( new_n730_, new_n721_, keyIn_0_47 );
and g623 ( new_n731_, new_n719_, new_n718_ );
or g624 ( new_n732_, new_n731_, new_n730_ );
not g625 ( new_n733_, new_n727_ );
and g626 ( new_n734_, new_n732_, new_n733_ );
and g627 ( new_n735_, new_n734_, keyIn_0_52 );
or g628 ( new_n736_, new_n729_, new_n735_ );
or g629 ( new_n737_, new_n716_, new_n736_ );
and g630 ( new_n738_, new_n647_, N115 );
and g631 ( new_n739_, N329, N112 );
and g632 ( new_n740_, N223, N102 );
or g633 ( new_n741_, new_n740_, new_n152_ );
or g634 ( new_n742_, new_n739_, new_n741_ );
or g635 ( new_n743_, new_n738_, new_n742_ );
and g636 ( new_n744_, new_n647_, N92 );
and g637 ( new_n745_, N329, N86 );
and g638 ( new_n746_, N223, N76 );
or g639 ( new_n747_, new_n746_, new_n180_ );
or g640 ( new_n748_, new_n745_, new_n747_ );
or g641 ( new_n749_, new_n744_, new_n748_ );
and g642 ( new_n750_, new_n647_, N105 );
and g643 ( new_n751_, N329, N99 );
and g644 ( new_n752_, N223, N89 );
or g645 ( new_n753_, new_n752_, new_n190_ );
or g646 ( new_n754_, new_n751_, new_n753_ );
or g647 ( new_n755_, new_n750_, new_n754_ );
and g648 ( new_n756_, new_n749_, new_n755_ );
and g649 ( new_n757_, new_n756_, new_n743_ );
not g650 ( new_n758_, new_n757_ );
and g651 ( new_n759_, new_n647_, N79 );
and g652 ( new_n760_, new_n759_, keyIn_0_50 );
not g653 ( new_n761_, new_n760_ );
or g654 ( new_n762_, new_n759_, keyIn_0_50 );
and g655 ( new_n763_, N329, N73 );
not g656 ( new_n764_, new_n763_ );
and g657 ( new_n765_, N223, N63 );
not g658 ( new_n766_, new_n765_ );
and g659 ( new_n767_, new_n766_, N69 );
and g660 ( new_n768_, new_n764_, new_n767_ );
and g661 ( new_n769_, new_n762_, new_n768_ );
and g662 ( new_n770_, new_n769_, new_n761_ );
and g663 ( new_n771_, new_n770_, keyIn_0_55 );
not g664 ( new_n772_, keyIn_0_55 );
not g665 ( new_n773_, keyIn_0_50 );
or g666 ( new_n774_, new_n657_, new_n452_ );
and g667 ( new_n775_, new_n774_, new_n773_ );
not g668 ( new_n776_, new_n768_ );
or g669 ( new_n777_, new_n775_, new_n776_ );
or g670 ( new_n778_, new_n777_, new_n760_ );
and g671 ( new_n779_, new_n778_, new_n772_ );
or g672 ( new_n780_, new_n779_, new_n771_ );
or g673 ( new_n781_, new_n780_, new_n758_ );
or g674 ( new_n782_, new_n737_, new_n781_ );
or g675 ( new_n783_, new_n782_, new_n694_ );
and g676 ( new_n784_, new_n783_, keyIn_0_56 );
not g677 ( new_n785_, keyIn_0_56 );
and g678 ( new_n786_, new_n714_, new_n710_ );
and g679 ( new_n787_, new_n708_, keyIn_0_51 );
or g680 ( new_n788_, new_n786_, new_n787_ );
or g681 ( new_n789_, new_n734_, keyIn_0_52 );
or g682 ( new_n790_, new_n728_, new_n717_ );
and g683 ( new_n791_, new_n790_, new_n789_ );
and g684 ( new_n792_, new_n788_, new_n791_ );
or g685 ( new_n793_, new_n778_, new_n772_ );
or g686 ( new_n794_, new_n770_, keyIn_0_55 );
and g687 ( new_n795_, new_n793_, new_n794_ );
and g688 ( new_n796_, new_n795_, new_n757_ );
and g689 ( new_n797_, new_n792_, new_n796_ );
and g690 ( new_n798_, new_n797_, new_n693_ );
and g691 ( new_n799_, new_n798_, new_n785_ );
or g692 ( new_n800_, new_n784_, new_n799_ );
and g693 ( new_n801_, new_n800_, new_n654_ );
and g694 ( new_n802_, new_n801_, new_n640_ );
not g695 ( new_n803_, new_n654_ );
or g696 ( new_n804_, new_n798_, new_n785_ );
not g697 ( new_n805_, new_n799_ );
and g698 ( new_n806_, new_n805_, new_n804_ );
or g699 ( new_n807_, new_n806_, new_n803_ );
and g700 ( new_n808_, new_n807_, keyIn_0_58 );
or g701 ( N421, new_n808_, new_n802_ );
not g702 ( new_n810_, keyIn_0_61 );
not g703 ( new_n811_, keyIn_0_57 );
or g704 ( new_n812_, new_n675_, new_n670_ );
or g705 ( new_n813_, new_n668_, keyIn_0_53 );
and g706 ( new_n814_, new_n813_, new_n812_ );
and g707 ( new_n815_, new_n814_, new_n811_ );
not g708 ( new_n816_, new_n815_ );
or g709 ( new_n817_, new_n814_, new_n811_ );
and g710 ( new_n818_, new_n817_, new_n791_ );
and g711 ( new_n819_, new_n818_, new_n816_ );
or g712 ( new_n820_, new_n819_, keyIn_0_59 );
not g713 ( new_n821_, keyIn_0_59 );
and g714 ( new_n822_, new_n677_, keyIn_0_57 );
or g715 ( new_n823_, new_n822_, new_n736_ );
or g716 ( new_n824_, new_n823_, new_n815_ );
or g717 ( new_n825_, new_n824_, new_n821_ );
and g718 ( new_n826_, new_n825_, new_n820_ );
and g719 ( new_n827_, new_n792_, new_n692_ );
not g720 ( new_n828_, new_n827_ );
or g721 ( new_n829_, new_n826_, new_n828_ );
and g722 ( new_n830_, new_n829_, new_n810_ );
and g723 ( new_n831_, new_n824_, new_n821_ );
and g724 ( new_n832_, new_n819_, keyIn_0_59 );
or g725 ( new_n833_, new_n831_, new_n832_ );
and g726 ( new_n834_, new_n833_, new_n827_ );
and g727 ( new_n835_, new_n834_, keyIn_0_61 );
or g728 ( N430, new_n830_, new_n835_ );
not g729 ( new_n837_, keyIn_0_62 );
not g730 ( new_n838_, keyIn_0_60 );
and g731 ( new_n839_, new_n677_, new_n791_ );
and g732 ( new_n840_, new_n692_, new_n780_ );
and g733 ( new_n841_, new_n840_, new_n839_ );
or g734 ( new_n842_, new_n841_, new_n838_ );
or g735 ( new_n843_, new_n736_, new_n814_ );
not g736 ( new_n844_, new_n691_ );
and g737 ( new_n845_, new_n844_, new_n689_ );
or g738 ( new_n846_, new_n845_, new_n795_ );
or g739 ( new_n847_, new_n843_, new_n846_ );
or g740 ( new_n848_, new_n847_, keyIn_0_60 );
and g741 ( new_n849_, new_n848_, new_n842_ );
not g742 ( new_n850_, new_n749_ );
and g743 ( new_n851_, new_n693_, new_n850_ );
or g744 ( new_n852_, new_n851_, new_n737_ );
or g745 ( new_n853_, new_n849_, new_n852_ );
and g746 ( new_n854_, new_n853_, new_n837_ );
not g747 ( new_n855_, new_n853_ );
and g748 ( new_n856_, new_n855_, keyIn_0_62 );
or g749 ( N431, new_n856_, new_n854_ );
and g750 ( new_n858_, new_n847_, keyIn_0_60 );
and g751 ( new_n859_, new_n841_, new_n838_ );
or g752 ( new_n860_, new_n858_, new_n859_ );
or g753 ( new_n861_, new_n850_, new_n755_ );
or g754 ( new_n862_, new_n843_, new_n861_ );
and g755 ( new_n863_, new_n862_, new_n788_ );
and g756 ( new_n864_, new_n860_, new_n863_ );
and g757 ( new_n865_, new_n864_, new_n833_ );
and g758 ( new_n866_, new_n865_, keyIn_0_63 );
not g759 ( new_n867_, keyIn_0_63 );
not g760 ( new_n868_, new_n863_ );
or g761 ( new_n869_, new_n849_, new_n868_ );
or g762 ( new_n870_, new_n869_, new_n826_ );
and g763 ( new_n871_, new_n870_, new_n867_ );
or g764 ( N432, new_n871_, new_n866_ );
endmodule