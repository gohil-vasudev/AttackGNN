module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063;

  NAND2_X1 U534 ( .A1(n518), .A2(n519), .ZN(Result_9_) );
  NAND2_X1 U535 ( .A1(n520), .A2(n521), .ZN(n519) );
  XNOR2_X1 U536 ( .A(n522), .B(n523), .ZN(n520) );
  XOR2_X1 U537 ( .A(n524), .B(n525), .Z(n523) );
  NAND2_X1 U538 ( .A1(b_7_), .A2(a_1_), .ZN(n525) );
  NAND2_X1 U539 ( .A1(n526), .A2(n527), .ZN(n518) );
  NAND2_X1 U540 ( .A1(n528), .A2(n529), .ZN(n527) );
  INV_X1 U541 ( .A(n530), .ZN(n529) );
  NOR2_X1 U542 ( .A1(n531), .A2(n532), .ZN(n530) );
  NOR2_X1 U543 ( .A1(n533), .A2(n534), .ZN(n531) );
  NAND2_X1 U544 ( .A1(n535), .A2(n532), .ZN(n528) );
  INV_X1 U545 ( .A(n536), .ZN(n532) );
  XNOR2_X1 U546 ( .A(n537), .B(a_1_), .ZN(n535) );
  NAND2_X1 U547 ( .A1(n538), .A2(n539), .ZN(Result_8_) );
  NAND2_X1 U548 ( .A1(n540), .A2(n521), .ZN(n539) );
  XOR2_X1 U549 ( .A(n541), .B(n542), .Z(n540) );
  XNOR2_X1 U550 ( .A(n543), .B(n544), .ZN(n542) );
  NAND2_X1 U551 ( .A1(n545), .A2(n526), .ZN(n538) );
  XNOR2_X1 U552 ( .A(n546), .B(n547), .ZN(n545) );
  NOR2_X1 U553 ( .A1(n534), .A2(n548), .ZN(n546) );
  NOR2_X1 U554 ( .A1(n533), .A2(n536), .ZN(n548) );
  NAND2_X1 U555 ( .A1(n549), .A2(n550), .ZN(n536) );
  NAND2_X1 U556 ( .A1(n551), .A2(n552), .ZN(n550) );
  NOR2_X1 U557 ( .A1(b_1_), .A2(a_1_), .ZN(n534) );
  NOR2_X1 U558 ( .A1(n526), .A2(n553), .ZN(Result_7_) );
  XNOR2_X1 U559 ( .A(n554), .B(n555), .ZN(n553) );
  NOR2_X1 U560 ( .A1(n556), .A2(n557), .ZN(Result_6_) );
  NAND2_X1 U561 ( .A1(n521), .A2(n558), .ZN(n557) );
  INV_X1 U562 ( .A(n559), .ZN(n558) );
  NOR2_X1 U563 ( .A1(n560), .A2(n561), .ZN(n556) );
  NOR2_X1 U564 ( .A1(n555), .A2(n554), .ZN(n560) );
  INV_X1 U565 ( .A(n562), .ZN(n555) );
  NOR2_X1 U566 ( .A1(n526), .A2(n563), .ZN(Result_5_) );
  XNOR2_X1 U567 ( .A(n559), .B(n564), .ZN(n563) );
  NOR2_X1 U568 ( .A1(n565), .A2(n566), .ZN(n564) );
  NOR2_X1 U569 ( .A1(n567), .A2(n568), .ZN(n566) );
  NOR2_X1 U570 ( .A1(n526), .A2(n569), .ZN(Result_4_) );
  XNOR2_X1 U571 ( .A(n570), .B(n571), .ZN(n569) );
  NOR2_X1 U572 ( .A1(n526), .A2(n572), .ZN(Result_3_) );
  XNOR2_X1 U573 ( .A(n573), .B(n574), .ZN(n572) );
  NOR2_X1 U574 ( .A1(n575), .A2(n576), .ZN(n573) );
  INV_X1 U575 ( .A(n577), .ZN(n576) );
  NOR2_X1 U576 ( .A1(n578), .A2(n579), .ZN(n575) );
  NOR2_X1 U577 ( .A1(n526), .A2(n580), .ZN(Result_2_) );
  XNOR2_X1 U578 ( .A(n581), .B(n582), .ZN(n580) );
  NOR2_X1 U579 ( .A1(n526), .A2(n583), .ZN(Result_1_) );
  XOR2_X1 U580 ( .A(n584), .B(n585), .Z(n583) );
  NOR2_X1 U581 ( .A1(n581), .A2(n582), .ZN(n585) );
  NAND2_X1 U582 ( .A1(n586), .A2(n587), .ZN(n584) );
  NAND2_X1 U583 ( .A1(n588), .A2(n589), .ZN(Result_15_) );
  NAND2_X1 U584 ( .A1(n590), .A2(n521), .ZN(n589) );
  NAND2_X1 U585 ( .A1(n526), .A2(n591), .ZN(n588) );
  NAND2_X1 U586 ( .A1(n592), .A2(n593), .ZN(n591) );
  NAND2_X1 U587 ( .A1(b_7_), .A2(n594), .ZN(n593) );
  NAND2_X1 U588 ( .A1(n595), .A2(n596), .ZN(Result_14_) );
  NAND2_X1 U589 ( .A1(n526), .A2(n597), .ZN(n596) );
  NAND2_X1 U590 ( .A1(n598), .A2(n599), .ZN(n597) );
  NOR2_X1 U591 ( .A1(n600), .A2(n601), .ZN(n598) );
  NOR2_X1 U592 ( .A1(n602), .A2(n603), .ZN(n601) );
  NAND2_X1 U593 ( .A1(n604), .A2(n605), .ZN(n603) );
  INV_X1 U594 ( .A(n590), .ZN(n604) );
  NOR2_X1 U595 ( .A1(b_6_), .A2(n606), .ZN(n600) );
  XNOR2_X1 U596 ( .A(n590), .B(a_6_), .ZN(n606) );
  NAND2_X1 U597 ( .A1(n607), .A2(n521), .ZN(n595) );
  XOR2_X1 U598 ( .A(n608), .B(n609), .Z(n607) );
  NAND2_X1 U599 ( .A1(b_7_), .A2(a_6_), .ZN(n609) );
  NAND2_X1 U600 ( .A1(n610), .A2(n611), .ZN(Result_13_) );
  NAND2_X1 U601 ( .A1(n526), .A2(n612), .ZN(n611) );
  NAND2_X1 U602 ( .A1(n613), .A2(n614), .ZN(n612) );
  NAND2_X1 U603 ( .A1(n615), .A2(n616), .ZN(n614) );
  NOR2_X1 U604 ( .A1(n617), .A2(n618), .ZN(n613) );
  NOR2_X1 U605 ( .A1(b_5_), .A2(n619), .ZN(n618) );
  XNOR2_X1 U606 ( .A(n620), .B(n621), .ZN(n619) );
  NOR2_X1 U607 ( .A1(n622), .A2(n623), .ZN(n617) );
  NAND2_X1 U608 ( .A1(n621), .A2(n620), .ZN(n623) );
  INV_X1 U609 ( .A(n616), .ZN(n621) );
  NAND2_X1 U610 ( .A1(n624), .A2(n521), .ZN(n610) );
  XNOR2_X1 U611 ( .A(n625), .B(n626), .ZN(n624) );
  XNOR2_X1 U612 ( .A(n627), .B(n599), .ZN(n626) );
  NAND2_X1 U613 ( .A1(n628), .A2(n629), .ZN(Result_12_) );
  NAND2_X1 U614 ( .A1(n630), .A2(n521), .ZN(n629) );
  XNOR2_X1 U615 ( .A(n631), .B(n632), .ZN(n630) );
  NAND2_X1 U616 ( .A1(n633), .A2(n634), .ZN(n631) );
  NAND2_X1 U617 ( .A1(n526), .A2(n635), .ZN(n628) );
  XNOR2_X1 U618 ( .A(n636), .B(n637), .ZN(n635) );
  NAND2_X1 U619 ( .A1(n638), .A2(n639), .ZN(n636) );
  NAND2_X1 U620 ( .A1(n640), .A2(n641), .ZN(Result_11_) );
  NAND2_X1 U621 ( .A1(n526), .A2(n642), .ZN(n641) );
  NAND2_X1 U622 ( .A1(n643), .A2(n644), .ZN(n642) );
  NAND2_X1 U623 ( .A1(n645), .A2(n646), .ZN(n644) );
  NOR2_X1 U624 ( .A1(n647), .A2(n648), .ZN(n643) );
  NOR2_X1 U625 ( .A1(b_3_), .A2(n649), .ZN(n648) );
  XNOR2_X1 U626 ( .A(a_3_), .B(n646), .ZN(n649) );
  INV_X1 U627 ( .A(n650), .ZN(n647) );
  NAND2_X1 U628 ( .A1(b_3_), .A2(n651), .ZN(n650) );
  NOR2_X1 U629 ( .A1(n646), .A2(a_3_), .ZN(n651) );
  NAND2_X1 U630 ( .A1(n652), .A2(n521), .ZN(n640) );
  XOR2_X1 U631 ( .A(n653), .B(n654), .Z(n652) );
  XOR2_X1 U632 ( .A(n655), .B(n656), .Z(n653) );
  NOR2_X1 U633 ( .A1(n657), .A2(n658), .ZN(n656) );
  NAND2_X1 U634 ( .A1(n659), .A2(n660), .ZN(Result_10_) );
  NAND2_X1 U635 ( .A1(n661), .A2(n521), .ZN(n660) );
  XNOR2_X1 U636 ( .A(n662), .B(n663), .ZN(n661) );
  XOR2_X1 U637 ( .A(n664), .B(n665), .Z(n663) );
  NAND2_X1 U638 ( .A1(b_7_), .A2(a_2_), .ZN(n665) );
  NAND2_X1 U639 ( .A1(n526), .A2(n666), .ZN(n659) );
  XNOR2_X1 U640 ( .A(n552), .B(n667), .ZN(n666) );
  NAND2_X1 U641 ( .A1(n551), .A2(n549), .ZN(n667) );
  NAND2_X1 U642 ( .A1(n668), .A2(n669), .ZN(n551) );
  NAND2_X1 U643 ( .A1(n670), .A2(n671), .ZN(n552) );
  NAND2_X1 U644 ( .A1(n672), .A2(n646), .ZN(n671) );
  NAND2_X1 U645 ( .A1(n638), .A2(n673), .ZN(n646) );
  NAND2_X1 U646 ( .A1(n639), .A2(n637), .ZN(n673) );
  NAND2_X1 U647 ( .A1(n674), .A2(n675), .ZN(n637) );
  NAND2_X1 U648 ( .A1(n676), .A2(n616), .ZN(n675) );
  NAND2_X1 U649 ( .A1(n677), .A2(n678), .ZN(n616) );
  NAND2_X1 U650 ( .A1(n590), .A2(n679), .ZN(n678) );
  NAND2_X1 U651 ( .A1(n602), .A2(n605), .ZN(n679) );
  INV_X1 U652 ( .A(n680), .ZN(n677) );
  NAND2_X1 U653 ( .A1(n622), .A2(n620), .ZN(n676) );
  NAND2_X1 U654 ( .A1(n681), .A2(n682), .ZN(n639) );
  NAND2_X1 U655 ( .A1(n683), .A2(n657), .ZN(n672) );
  INV_X1 U656 ( .A(n645), .ZN(n670) );
  NOR2_X1 U657 ( .A1(n526), .A2(n684), .ZN(Result_0_) );
  NOR2_X1 U658 ( .A1(n685), .A2(n686), .ZN(n684) );
  NAND2_X1 U659 ( .A1(n586), .A2(n687), .ZN(n686) );
  NAND2_X1 U660 ( .A1(n688), .A2(n689), .ZN(n586) );
  INV_X1 U661 ( .A(n690), .ZN(n689) );
  NAND2_X1 U662 ( .A1(n687), .A2(n691), .ZN(n690) );
  NAND2_X1 U663 ( .A1(n692), .A2(b_0_), .ZN(n687) );
  NOR2_X1 U664 ( .A1(n693), .A2(n694), .ZN(n688) );
  NOR2_X1 U665 ( .A1(n582), .A2(n695), .ZN(n685) );
  NAND2_X1 U666 ( .A1(n587), .A2(n696), .ZN(n695) );
  INV_X1 U667 ( .A(n581), .ZN(n696) );
  NOR2_X1 U668 ( .A1(n697), .A2(n698), .ZN(n581) );
  INV_X1 U669 ( .A(n699), .ZN(n698) );
  NAND2_X1 U670 ( .A1(n700), .A2(n701), .ZN(n699) );
  NAND2_X1 U671 ( .A1(n577), .A2(n702), .ZN(n697) );
  NAND2_X1 U672 ( .A1(n578), .A2(n574), .ZN(n702) );
  NOR2_X1 U673 ( .A1(n570), .A2(n571), .ZN(n574) );
  INV_X1 U674 ( .A(n703), .ZN(n571) );
  NAND2_X1 U675 ( .A1(n704), .A2(n705), .ZN(n703) );
  NAND2_X1 U676 ( .A1(n559), .A2(n568), .ZN(n705) );
  NOR2_X1 U677 ( .A1(n706), .A2(n554), .ZN(n559) );
  NAND2_X1 U678 ( .A1(n707), .A2(n708), .ZN(n554) );
  NAND2_X1 U679 ( .A1(n541), .A2(n709), .ZN(n708) );
  NAND2_X1 U680 ( .A1(n544), .A2(n543), .ZN(n709) );
  XNOR2_X1 U681 ( .A(n710), .B(n711), .ZN(n541) );
  XOR2_X1 U682 ( .A(n712), .B(n713), .Z(n710) );
  NOR2_X1 U683 ( .A1(n714), .A2(n602), .ZN(n713) );
  INV_X1 U684 ( .A(n715), .ZN(n707) );
  NOR2_X1 U685 ( .A1(n543), .A2(n544), .ZN(n715) );
  NOR2_X1 U686 ( .A1(n658), .A2(n716), .ZN(n544) );
  NAND2_X1 U687 ( .A1(n717), .A2(n718), .ZN(n543) );
  NAND2_X1 U688 ( .A1(n719), .A2(b_7_), .ZN(n718) );
  NOR2_X1 U689 ( .A1(n720), .A2(n714), .ZN(n719) );
  NOR2_X1 U690 ( .A1(n522), .A2(n524), .ZN(n720) );
  NAND2_X1 U691 ( .A1(n522), .A2(n524), .ZN(n717) );
  NAND2_X1 U692 ( .A1(n721), .A2(n722), .ZN(n524) );
  NAND2_X1 U693 ( .A1(n723), .A2(b_7_), .ZN(n722) );
  NOR2_X1 U694 ( .A1(n724), .A2(n669), .ZN(n723) );
  NOR2_X1 U695 ( .A1(n662), .A2(n664), .ZN(n724) );
  NAND2_X1 U696 ( .A1(n662), .A2(n664), .ZN(n721) );
  NAND2_X1 U697 ( .A1(n725), .A2(n726), .ZN(n664) );
  NAND2_X1 U698 ( .A1(n727), .A2(b_7_), .ZN(n726) );
  NOR2_X1 U699 ( .A1(n728), .A2(n657), .ZN(n727) );
  NOR2_X1 U700 ( .A1(n654), .A2(n655), .ZN(n728) );
  NAND2_X1 U701 ( .A1(n654), .A2(n655), .ZN(n725) );
  NAND2_X1 U702 ( .A1(n633), .A2(n729), .ZN(n655) );
  NAND2_X1 U703 ( .A1(n632), .A2(n634), .ZN(n729) );
  NAND2_X1 U704 ( .A1(n730), .A2(n731), .ZN(n634) );
  NAND2_X1 U705 ( .A1(b_7_), .A2(a_4_), .ZN(n731) );
  XNOR2_X1 U706 ( .A(n732), .B(n733), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n734), .B(n735), .ZN(n732) );
  INV_X1 U708 ( .A(n736), .ZN(n633) );
  NOR2_X1 U709 ( .A1(n682), .A2(n730), .ZN(n736) );
  NOR2_X1 U710 ( .A1(n737), .A2(n738), .ZN(n730) );
  INV_X1 U711 ( .A(n739), .ZN(n738) );
  NAND2_X1 U712 ( .A1(n627), .A2(n740), .ZN(n739) );
  NAND2_X1 U713 ( .A1(n625), .A2(n599), .ZN(n740) );
  NOR2_X1 U714 ( .A1(n658), .A2(n620), .ZN(n627) );
  NOR2_X1 U715 ( .A1(n599), .A2(n625), .ZN(n737) );
  XNOR2_X1 U716 ( .A(n680), .B(n741), .ZN(n625) );
  NOR2_X1 U717 ( .A1(n594), .A2(n622), .ZN(n741) );
  NAND2_X1 U718 ( .A1(n680), .A2(n590), .ZN(n599) );
  NOR2_X1 U719 ( .A1(n658), .A2(n594), .ZN(n590) );
  INV_X1 U720 ( .A(b_7_), .ZN(n658) );
  NOR2_X1 U721 ( .A1(n602), .A2(n605), .ZN(n680) );
  XOR2_X1 U722 ( .A(n742), .B(n743), .Z(n654) );
  XOR2_X1 U723 ( .A(n744), .B(n745), .Z(n743) );
  XNOR2_X1 U724 ( .A(n746), .B(n747), .ZN(n662) );
  XOR2_X1 U725 ( .A(n748), .B(n749), .Z(n747) );
  XNOR2_X1 U726 ( .A(n750), .B(n751), .ZN(n522) );
  XNOR2_X1 U727 ( .A(n752), .B(n753), .ZN(n751) );
  NAND2_X1 U728 ( .A1(n562), .A2(n561), .ZN(n706) );
  XOR2_X1 U729 ( .A(n754), .B(n755), .Z(n561) );
  XOR2_X1 U730 ( .A(n756), .B(n757), .Z(n562) );
  XNOR2_X1 U731 ( .A(n758), .B(n759), .ZN(n757) );
  NOR2_X1 U732 ( .A1(n565), .A2(n760), .ZN(n704) );
  NOR2_X1 U733 ( .A1(n761), .A2(n762), .ZN(n760) );
  INV_X1 U734 ( .A(n763), .ZN(n565) );
  NAND2_X1 U735 ( .A1(n567), .A2(n568), .ZN(n763) );
  XOR2_X1 U736 ( .A(n762), .B(n761), .Z(n568) );
  XOR2_X1 U737 ( .A(n764), .B(n765), .Z(n761) );
  XNOR2_X1 U738 ( .A(n766), .B(n767), .ZN(n764) );
  NAND2_X1 U739 ( .A1(n768), .A2(n769), .ZN(n762) );
  NAND2_X1 U740 ( .A1(n770), .A2(n771), .ZN(n769) );
  NAND2_X1 U741 ( .A1(n772), .A2(n773), .ZN(n771) );
  INV_X1 U742 ( .A(n774), .ZN(n768) );
  NOR2_X1 U743 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U744 ( .A1(n755), .A2(n754), .ZN(n567) );
  NAND2_X1 U745 ( .A1(n775), .A2(n776), .ZN(n754) );
  NAND2_X1 U746 ( .A1(n756), .A2(n777), .ZN(n776) );
  NAND2_X1 U747 ( .A1(n759), .A2(n758), .ZN(n777) );
  XOR2_X1 U748 ( .A(n778), .B(n779), .Z(n756) );
  XOR2_X1 U749 ( .A(n780), .B(n781), .Z(n779) );
  NAND2_X1 U750 ( .A1(b_5_), .A2(a_1_), .ZN(n781) );
  INV_X1 U751 ( .A(n782), .ZN(n775) );
  NOR2_X1 U752 ( .A1(n758), .A2(n759), .ZN(n782) );
  NOR2_X1 U753 ( .A1(n716), .A2(n602), .ZN(n759) );
  NAND2_X1 U754 ( .A1(n783), .A2(n784), .ZN(n758) );
  NAND2_X1 U755 ( .A1(n785), .A2(b_6_), .ZN(n784) );
  NOR2_X1 U756 ( .A1(n786), .A2(n714), .ZN(n785) );
  NOR2_X1 U757 ( .A1(n712), .A2(n711), .ZN(n786) );
  NAND2_X1 U758 ( .A1(n711), .A2(n712), .ZN(n783) );
  NAND2_X1 U759 ( .A1(n787), .A2(n788), .ZN(n712) );
  NAND2_X1 U760 ( .A1(n753), .A2(n789), .ZN(n788) );
  INV_X1 U761 ( .A(n790), .ZN(n789) );
  NOR2_X1 U762 ( .A1(n750), .A2(n752), .ZN(n790) );
  NOR2_X1 U763 ( .A1(n669), .A2(n602), .ZN(n753) );
  NAND2_X1 U764 ( .A1(n750), .A2(n752), .ZN(n787) );
  NAND2_X1 U765 ( .A1(n791), .A2(n792), .ZN(n752) );
  INV_X1 U766 ( .A(n793), .ZN(n792) );
  NOR2_X1 U767 ( .A1(n749), .A2(n794), .ZN(n793) );
  NOR2_X1 U768 ( .A1(n748), .A2(n746), .ZN(n794) );
  NAND2_X1 U769 ( .A1(a_3_), .A2(b_6_), .ZN(n749) );
  NAND2_X1 U770 ( .A1(n746), .A2(n748), .ZN(n791) );
  NAND2_X1 U771 ( .A1(n795), .A2(n796), .ZN(n748) );
  NAND2_X1 U772 ( .A1(n745), .A2(n797), .ZN(n796) );
  NAND2_X1 U773 ( .A1(n798), .A2(n799), .ZN(n797) );
  INV_X1 U774 ( .A(n744), .ZN(n799) );
  NOR2_X1 U775 ( .A1(n682), .A2(n602), .ZN(n745) );
  NAND2_X1 U776 ( .A1(n744), .A2(n742), .ZN(n795) );
  INV_X1 U777 ( .A(n798), .ZN(n742) );
  XOR2_X1 U778 ( .A(n800), .B(n801), .Z(n798) );
  XOR2_X1 U779 ( .A(n674), .B(n802), .Z(n800) );
  NOR2_X1 U780 ( .A1(n803), .A2(n804), .ZN(n744) );
  NOR2_X1 U781 ( .A1(n805), .A2(n735), .ZN(n804) );
  NOR2_X1 U782 ( .A1(n608), .A2(n806), .ZN(n735) );
  NAND2_X1 U783 ( .A1(b_6_), .A2(a_7_), .ZN(n608) );
  INV_X1 U784 ( .A(n807), .ZN(n805) );
  NAND2_X1 U785 ( .A1(n734), .A2(n733), .ZN(n807) );
  NOR2_X1 U786 ( .A1(n733), .A2(n734), .ZN(n803) );
  NOR2_X1 U787 ( .A1(n620), .A2(n602), .ZN(n734) );
  XNOR2_X1 U788 ( .A(n806), .B(n808), .ZN(n733) );
  NOR2_X1 U789 ( .A1(n594), .A2(n681), .ZN(n808) );
  XNOR2_X1 U790 ( .A(n809), .B(n810), .ZN(n746) );
  NAND2_X1 U791 ( .A1(n811), .A2(n812), .ZN(n809) );
  XNOR2_X1 U792 ( .A(n813), .B(n814), .ZN(n750) );
  XOR2_X1 U793 ( .A(n815), .B(n816), .Z(n814) );
  NAND2_X1 U794 ( .A1(a_3_), .A2(b_5_), .ZN(n816) );
  XNOR2_X1 U795 ( .A(n817), .B(n818), .ZN(n711) );
  XOR2_X1 U796 ( .A(n819), .B(n820), .Z(n818) );
  NAND2_X1 U797 ( .A1(a_2_), .A2(b_5_), .ZN(n820) );
  XNOR2_X1 U798 ( .A(n770), .B(n821), .ZN(n755) );
  XNOR2_X1 U799 ( .A(n773), .B(n772), .ZN(n821) );
  NOR2_X1 U800 ( .A1(n716), .A2(n622), .ZN(n772) );
  NAND2_X1 U801 ( .A1(n822), .A2(n823), .ZN(n773) );
  NAND2_X1 U802 ( .A1(n824), .A2(b_5_), .ZN(n823) );
  NOR2_X1 U803 ( .A1(n825), .A2(n714), .ZN(n824) );
  NOR2_X1 U804 ( .A1(n780), .A2(n778), .ZN(n825) );
  NAND2_X1 U805 ( .A1(n778), .A2(n780), .ZN(n822) );
  NAND2_X1 U806 ( .A1(n826), .A2(n827), .ZN(n780) );
  NAND2_X1 U807 ( .A1(n828), .A2(a_2_), .ZN(n827) );
  NOR2_X1 U808 ( .A1(n829), .A2(n622), .ZN(n828) );
  NOR2_X1 U809 ( .A1(n817), .A2(n819), .ZN(n829) );
  NAND2_X1 U810 ( .A1(n817), .A2(n819), .ZN(n826) );
  NAND2_X1 U811 ( .A1(n830), .A2(n831), .ZN(n819) );
  NAND2_X1 U812 ( .A1(n832), .A2(a_3_), .ZN(n831) );
  NOR2_X1 U813 ( .A1(n833), .A2(n622), .ZN(n832) );
  INV_X1 U814 ( .A(b_5_), .ZN(n622) );
  NOR2_X1 U815 ( .A1(n813), .A2(n815), .ZN(n833) );
  NAND2_X1 U816 ( .A1(n813), .A2(n815), .ZN(n830) );
  NAND2_X1 U817 ( .A1(n811), .A2(n834), .ZN(n815) );
  NAND2_X1 U818 ( .A1(n810), .A2(n812), .ZN(n834) );
  NAND2_X1 U819 ( .A1(n835), .A2(n836), .ZN(n812) );
  NAND2_X1 U820 ( .A1(a_4_), .A2(b_5_), .ZN(n836) );
  INV_X1 U821 ( .A(n837), .ZN(n835) );
  XOR2_X1 U822 ( .A(n838), .B(n839), .Z(n810) );
  XOR2_X1 U823 ( .A(n840), .B(n841), .Z(n839) );
  NAND2_X1 U824 ( .A1(a_4_), .A2(n837), .ZN(n811) );
  NAND2_X1 U825 ( .A1(n842), .A2(n843), .ZN(n837) );
  NAND2_X1 U826 ( .A1(n802), .A2(n844), .ZN(n843) );
  INV_X1 U827 ( .A(n845), .ZN(n844) );
  NOR2_X1 U828 ( .A1(n801), .A2(n615), .ZN(n845) );
  NOR2_X1 U829 ( .A1(n846), .A2(n806), .ZN(n802) );
  NAND2_X1 U830 ( .A1(b_5_), .A2(a_6_), .ZN(n806) );
  NAND2_X1 U831 ( .A1(a_7_), .A2(b_4_), .ZN(n846) );
  NAND2_X1 U832 ( .A1(n615), .A2(n801), .ZN(n842) );
  XOR2_X1 U833 ( .A(n847), .B(n848), .Z(n801) );
  INV_X1 U834 ( .A(n674), .ZN(n615) );
  NAND2_X1 U835 ( .A1(a_5_), .A2(b_5_), .ZN(n674) );
  XOR2_X1 U836 ( .A(n849), .B(n850), .Z(n813) );
  XOR2_X1 U837 ( .A(n851), .B(n638), .Z(n849) );
  XNOR2_X1 U838 ( .A(n852), .B(n853), .ZN(n817) );
  XNOR2_X1 U839 ( .A(n854), .B(n855), .ZN(n853) );
  XOR2_X1 U840 ( .A(n856), .B(n857), .Z(n778) );
  XOR2_X1 U841 ( .A(n858), .B(n859), .Z(n857) );
  XOR2_X1 U842 ( .A(n860), .B(n861), .Z(n770) );
  XNOR2_X1 U843 ( .A(n862), .B(n863), .ZN(n860) );
  XNOR2_X1 U844 ( .A(n864), .B(n865), .ZN(n570) );
  NAND2_X1 U845 ( .A1(n579), .A2(n578), .ZN(n577) );
  XOR2_X1 U846 ( .A(n701), .B(n700), .Z(n578) );
  XOR2_X1 U847 ( .A(n866), .B(n867), .Z(n700) );
  XOR2_X1 U848 ( .A(n868), .B(n869), .Z(n867) );
  NAND2_X1 U849 ( .A1(a_0_), .A2(b_2_), .ZN(n869) );
  NAND2_X1 U850 ( .A1(n870), .A2(n871), .ZN(n701) );
  NAND2_X1 U851 ( .A1(n872), .A2(n873), .ZN(n871) );
  INV_X1 U852 ( .A(n874), .ZN(n873) );
  NOR2_X1 U853 ( .A1(n875), .A2(n876), .ZN(n874) );
  NAND2_X1 U854 ( .A1(n876), .A2(n875), .ZN(n870) );
  NOR2_X1 U855 ( .A1(n864), .A2(n865), .ZN(n579) );
  XNOR2_X1 U856 ( .A(n877), .B(n872), .ZN(n865) );
  XNOR2_X1 U857 ( .A(n878), .B(n879), .ZN(n872) );
  XNOR2_X1 U858 ( .A(n880), .B(n881), .ZN(n878) );
  XOR2_X1 U859 ( .A(n876), .B(n875), .Z(n877) );
  NAND2_X1 U860 ( .A1(n882), .A2(n883), .ZN(n875) );
  NAND2_X1 U861 ( .A1(n884), .A2(n885), .ZN(n883) );
  INV_X1 U862 ( .A(n886), .ZN(n885) );
  NOR2_X1 U863 ( .A1(n887), .A2(n888), .ZN(n886) );
  NAND2_X1 U864 ( .A1(n888), .A2(n887), .ZN(n882) );
  NOR2_X1 U865 ( .A1(n716), .A2(n683), .ZN(n876) );
  NOR2_X1 U866 ( .A1(n889), .A2(n890), .ZN(n864) );
  INV_X1 U867 ( .A(n891), .ZN(n890) );
  NAND2_X1 U868 ( .A1(n767), .A2(n892), .ZN(n891) );
  NAND2_X1 U869 ( .A1(n765), .A2(n766), .ZN(n892) );
  NOR2_X1 U870 ( .A1(n716), .A2(n681), .ZN(n767) );
  NOR2_X1 U871 ( .A1(n765), .A2(n766), .ZN(n889) );
  NOR2_X1 U872 ( .A1(n893), .A2(n894), .ZN(n766) );
  INV_X1 U873 ( .A(n895), .ZN(n894) );
  NAND2_X1 U874 ( .A1(n863), .A2(n896), .ZN(n895) );
  NAND2_X1 U875 ( .A1(n861), .A2(n862), .ZN(n896) );
  NOR2_X1 U876 ( .A1(n681), .A2(n714), .ZN(n863) );
  NOR2_X1 U877 ( .A1(n861), .A2(n862), .ZN(n893) );
  NOR2_X1 U878 ( .A1(n897), .A2(n898), .ZN(n862) );
  INV_X1 U879 ( .A(n899), .ZN(n898) );
  NAND2_X1 U880 ( .A1(n859), .A2(n900), .ZN(n899) );
  NAND2_X1 U881 ( .A1(n858), .A2(n856), .ZN(n900) );
  NOR2_X1 U882 ( .A1(n669), .A2(n681), .ZN(n859) );
  NOR2_X1 U883 ( .A1(n856), .A2(n858), .ZN(n897) );
  NOR2_X1 U884 ( .A1(n901), .A2(n902), .ZN(n858) );
  INV_X1 U885 ( .A(n903), .ZN(n902) );
  NAND2_X1 U886 ( .A1(n855), .A2(n904), .ZN(n903) );
  NAND2_X1 U887 ( .A1(n852), .A2(n854), .ZN(n904) );
  NOR2_X1 U888 ( .A1(n657), .A2(n681), .ZN(n855) );
  NOR2_X1 U889 ( .A1(n852), .A2(n854), .ZN(n901) );
  NAND2_X1 U890 ( .A1(n905), .A2(n906), .ZN(n854) );
  INV_X1 U891 ( .A(n907), .ZN(n906) );
  NOR2_X1 U892 ( .A1(n850), .A2(n908), .ZN(n907) );
  NOR2_X1 U893 ( .A1(n638), .A2(n851), .ZN(n908) );
  XNOR2_X1 U894 ( .A(n909), .B(n910), .ZN(n850) );
  XNOR2_X1 U895 ( .A(n911), .B(n912), .ZN(n910) );
  NAND2_X1 U896 ( .A1(n851), .A2(n638), .ZN(n905) );
  NAND2_X1 U897 ( .A1(b_4_), .A2(a_4_), .ZN(n638) );
  NOR2_X1 U898 ( .A1(n913), .A2(n914), .ZN(n851) );
  INV_X1 U899 ( .A(n915), .ZN(n914) );
  NAND2_X1 U900 ( .A1(n838), .A2(n916), .ZN(n915) );
  NAND2_X1 U901 ( .A1(n841), .A2(n840), .ZN(n916) );
  NOR2_X1 U902 ( .A1(n681), .A2(n620), .ZN(n838) );
  NOR2_X1 U903 ( .A1(n840), .A2(n841), .ZN(n913) );
  NAND2_X1 U904 ( .A1(n917), .A2(n918), .ZN(n841) );
  NAND2_X1 U905 ( .A1(n919), .A2(n920), .ZN(n918) );
  INV_X1 U906 ( .A(n912), .ZN(n917) );
  NAND2_X1 U907 ( .A1(n848), .A2(n847), .ZN(n840) );
  NOR2_X1 U908 ( .A1(n681), .A2(n605), .ZN(n847) );
  NOR2_X1 U909 ( .A1(n683), .A2(n594), .ZN(n848) );
  XNOR2_X1 U910 ( .A(n921), .B(n922), .ZN(n852) );
  XOR2_X1 U911 ( .A(n923), .B(n924), .Z(n921) );
  XOR2_X1 U912 ( .A(n925), .B(n926), .Z(n856) );
  XNOR2_X1 U913 ( .A(n927), .B(n645), .ZN(n925) );
  XOR2_X1 U914 ( .A(n928), .B(n929), .Z(n861) );
  XNOR2_X1 U915 ( .A(n930), .B(n931), .ZN(n928) );
  XOR2_X1 U916 ( .A(n884), .B(n932), .Z(n765) );
  XNOR2_X1 U917 ( .A(n887), .B(n888), .ZN(n932) );
  NOR2_X1 U918 ( .A1(n683), .A2(n714), .ZN(n888) );
  NAND2_X1 U919 ( .A1(n933), .A2(n934), .ZN(n887) );
  NAND2_X1 U920 ( .A1(n929), .A2(n935), .ZN(n934) );
  INV_X1 U921 ( .A(n936), .ZN(n935) );
  NOR2_X1 U922 ( .A1(n931), .A2(n930), .ZN(n936) );
  XOR2_X1 U923 ( .A(n937), .B(n938), .Z(n929) );
  XOR2_X1 U924 ( .A(n939), .B(n940), .Z(n937) );
  NAND2_X1 U925 ( .A1(n931), .A2(n930), .ZN(n933) );
  NOR2_X1 U926 ( .A1(n941), .A2(n942), .ZN(n930) );
  NOR2_X1 U927 ( .A1(n943), .A2(n645), .ZN(n942) );
  NOR2_X1 U928 ( .A1(n657), .A2(n683), .ZN(n645) );
  NOR2_X1 U929 ( .A1(n926), .A2(n927), .ZN(n943) );
  INV_X1 U930 ( .A(n944), .ZN(n941) );
  NAND2_X1 U931 ( .A1(n926), .A2(n927), .ZN(n944) );
  NOR2_X1 U932 ( .A1(n945), .A2(n946), .ZN(n927) );
  INV_X1 U933 ( .A(n947), .ZN(n946) );
  NAND2_X1 U934 ( .A1(n922), .A2(n948), .ZN(n947) );
  NAND2_X1 U935 ( .A1(n923), .A2(n924), .ZN(n948) );
  XNOR2_X1 U936 ( .A(n949), .B(n950), .ZN(n922) );
  NAND2_X1 U937 ( .A1(n951), .A2(n952), .ZN(n949) );
  NOR2_X1 U938 ( .A1(n924), .A2(n923), .ZN(n945) );
  NOR2_X1 U939 ( .A1(n953), .A2(n954), .ZN(n923) );
  INV_X1 U940 ( .A(n955), .ZN(n954) );
  NAND2_X1 U941 ( .A1(n912), .A2(n956), .ZN(n955) );
  NAND2_X1 U942 ( .A1(n911), .A2(n909), .ZN(n956) );
  NOR2_X1 U943 ( .A1(n919), .A2(n920), .ZN(n912) );
  NAND2_X1 U944 ( .A1(b_3_), .A2(a_6_), .ZN(n919) );
  NOR2_X1 U945 ( .A1(n909), .A2(n911), .ZN(n953) );
  NAND2_X1 U946 ( .A1(n957), .A2(n958), .ZN(n911) );
  NAND2_X1 U947 ( .A1(n959), .A2(n960), .ZN(n958) );
  NAND2_X1 U948 ( .A1(b_1_), .A2(a_7_), .ZN(n960) );
  NAND2_X1 U949 ( .A1(b_2_), .A2(a_6_), .ZN(n959) );
  NAND2_X1 U950 ( .A1(b_3_), .A2(a_5_), .ZN(n909) );
  NAND2_X1 U951 ( .A1(b_3_), .A2(a_4_), .ZN(n924) );
  XOR2_X1 U952 ( .A(n961), .B(n962), .Z(n926) );
  NAND2_X1 U953 ( .A1(n963), .A2(n964), .ZN(n961) );
  NOR2_X1 U954 ( .A1(n669), .A2(n683), .ZN(n931) );
  XOR2_X1 U955 ( .A(n965), .B(n966), .Z(n884) );
  XNOR2_X1 U956 ( .A(n549), .B(n967), .ZN(n966) );
  NAND2_X1 U957 ( .A1(n968), .A2(n969), .ZN(n587) );
  NAND2_X1 U958 ( .A1(b_0_), .A2(n970), .ZN(n969) );
  NAND2_X1 U959 ( .A1(n971), .A2(n691), .ZN(n968) );
  INV_X1 U960 ( .A(n693), .ZN(n971) );
  XOR2_X1 U961 ( .A(n693), .B(n691), .Z(n582) );
  NAND2_X1 U962 ( .A1(n972), .A2(n973), .ZN(n691) );
  NOR2_X1 U963 ( .A1(n974), .A2(n975), .ZN(n972) );
  NOR2_X1 U964 ( .A1(b_0_), .A2(n970), .ZN(n975) );
  INV_X1 U965 ( .A(n692), .ZN(n970) );
  NOR2_X1 U966 ( .A1(n976), .A2(n694), .ZN(n974) );
  NOR2_X1 U967 ( .A1(n977), .A2(n978), .ZN(n976) );
  NOR2_X1 U968 ( .A1(n692), .A2(n714), .ZN(n978) );
  NOR2_X1 U969 ( .A1(n716), .A2(n537), .ZN(n692) );
  NOR2_X1 U970 ( .A1(n669), .A2(n979), .ZN(n977) );
  INV_X1 U971 ( .A(n533), .ZN(n979) );
  NOR2_X1 U972 ( .A1(n868), .A2(n980), .ZN(n693) );
  NOR2_X1 U973 ( .A1(n866), .A2(n668), .ZN(n980) );
  XOR2_X1 U974 ( .A(n981), .B(n982), .Z(n866) );
  NOR2_X1 U975 ( .A1(n694), .A2(n669), .ZN(n982) );
  NAND2_X1 U976 ( .A1(n533), .A2(n973), .ZN(n981) );
  INV_X1 U977 ( .A(n983), .ZN(n973) );
  NAND2_X1 U978 ( .A1(n984), .A2(n985), .ZN(n983) );
  NAND2_X1 U979 ( .A1(n986), .A2(b_1_), .ZN(n985) );
  NOR2_X1 U980 ( .A1(n987), .A2(n669), .ZN(n986) );
  NOR2_X1 U981 ( .A1(n988), .A2(n989), .ZN(n987) );
  NAND2_X1 U982 ( .A1(n988), .A2(n989), .ZN(n984) );
  NOR2_X1 U983 ( .A1(n537), .A2(n714), .ZN(n533) );
  NAND2_X1 U984 ( .A1(n990), .A2(n991), .ZN(n868) );
  NAND2_X1 U985 ( .A1(n880), .A2(n992), .ZN(n991) );
  INV_X1 U986 ( .A(n993), .ZN(n992) );
  NOR2_X1 U987 ( .A1(n879), .A2(n881), .ZN(n993) );
  NOR2_X1 U988 ( .A1(n668), .A2(n714), .ZN(n880) );
  INV_X1 U989 ( .A(a_1_), .ZN(n714) );
  NAND2_X1 U990 ( .A1(n879), .A2(n881), .ZN(n990) );
  NOR2_X1 U991 ( .A1(n994), .A2(n995), .ZN(n881) );
  INV_X1 U992 ( .A(n996), .ZN(n995) );
  NAND2_X1 U993 ( .A1(n997), .A2(n549), .ZN(n996) );
  NAND2_X1 U994 ( .A1(b_2_), .A2(a_2_), .ZN(n549) );
  NAND2_X1 U995 ( .A1(n965), .A2(n967), .ZN(n997) );
  NOR2_X1 U996 ( .A1(n965), .A2(n967), .ZN(n994) );
  NOR2_X1 U997 ( .A1(n998), .A2(n999), .ZN(n967) );
  NOR2_X1 U998 ( .A1(n1000), .A2(n940), .ZN(n999) );
  NOR2_X1 U999 ( .A1(n668), .A2(n657), .ZN(n940) );
  INV_X1 U1000 ( .A(n1001), .ZN(n1000) );
  NAND2_X1 U1001 ( .A1(n938), .A2(n939), .ZN(n1001) );
  NOR2_X1 U1002 ( .A1(n939), .A2(n938), .ZN(n998) );
  XOR2_X1 U1003 ( .A(n1002), .B(n1003), .Z(n938) );
  NOR2_X1 U1004 ( .A1(n694), .A2(n620), .ZN(n1003) );
  XOR2_X1 U1005 ( .A(n1004), .B(n1005), .Z(n1002) );
  NAND2_X1 U1006 ( .A1(n963), .A2(n1006), .ZN(n939) );
  NAND2_X1 U1007 ( .A1(n962), .A2(n964), .ZN(n1006) );
  NAND2_X1 U1008 ( .A1(n1007), .A2(n1008), .ZN(n964) );
  NAND2_X1 U1009 ( .A1(b_2_), .A2(a_4_), .ZN(n1008) );
  INV_X1 U1010 ( .A(n1009), .ZN(n1007) );
  XNOR2_X1 U1011 ( .A(n1010), .B(n1011), .ZN(n962) );
  XOR2_X1 U1012 ( .A(n1012), .B(n1013), .Z(n1010) );
  NAND2_X1 U1013 ( .A1(a_4_), .A2(n1009), .ZN(n963) );
  NAND2_X1 U1014 ( .A1(n951), .A2(n1014), .ZN(n1009) );
  NAND2_X1 U1015 ( .A1(n950), .A2(n952), .ZN(n1014) );
  NAND2_X1 U1016 ( .A1(n957), .A2(n1015), .ZN(n952) );
  NAND2_X1 U1017 ( .A1(b_2_), .A2(a_5_), .ZN(n1015) );
  INV_X1 U1018 ( .A(n1016), .ZN(n957) );
  INV_X1 U1019 ( .A(n1017), .ZN(n950) );
  NAND2_X1 U1020 ( .A1(n1013), .A2(n1018), .ZN(n1017) );
  NAND2_X1 U1021 ( .A1(n1019), .A2(n1020), .ZN(n1018) );
  NAND2_X1 U1022 ( .A1(n1016), .A2(a_5_), .ZN(n951) );
  NOR2_X1 U1023 ( .A1(n920), .A2(n1020), .ZN(n1016) );
  NAND2_X1 U1024 ( .A1(b_2_), .A2(a_7_), .ZN(n920) );
  XOR2_X1 U1025 ( .A(n1021), .B(n1022), .Z(n965) );
  XNOR2_X1 U1026 ( .A(n1023), .B(n1024), .ZN(n1022) );
  NAND2_X1 U1027 ( .A1(a_4_), .A2(b_0_), .ZN(n1021) );
  XOR2_X1 U1028 ( .A(n1025), .B(n1026), .Z(n879) );
  XNOR2_X1 U1029 ( .A(n988), .B(n989), .ZN(n1026) );
  NAND2_X1 U1030 ( .A1(n1027), .A2(n1028), .ZN(n989) );
  NAND2_X1 U1031 ( .A1(n1029), .A2(a_4_), .ZN(n1028) );
  NOR2_X1 U1032 ( .A1(n1030), .A2(n694), .ZN(n1029) );
  NOR2_X1 U1033 ( .A1(n1023), .A2(n1024), .ZN(n1030) );
  NAND2_X1 U1034 ( .A1(n1023), .A2(n1024), .ZN(n1027) );
  NAND2_X1 U1035 ( .A1(n1031), .A2(n1032), .ZN(n1024) );
  NAND2_X1 U1036 ( .A1(n1033), .A2(a_5_), .ZN(n1032) );
  NOR2_X1 U1037 ( .A1(n1034), .A2(n694), .ZN(n1033) );
  NOR2_X1 U1038 ( .A1(n1004), .A2(n1005), .ZN(n1034) );
  NAND2_X1 U1039 ( .A1(n1004), .A2(n1005), .ZN(n1031) );
  NAND2_X1 U1040 ( .A1(n1013), .A2(n1035), .ZN(n1005) );
  NAND2_X1 U1041 ( .A1(n1011), .A2(n1012), .ZN(n1035) );
  NOR2_X1 U1042 ( .A1(n537), .A2(n620), .ZN(n1012) );
  NOR2_X1 U1043 ( .A1(n694), .A2(n605), .ZN(n1011) );
  INV_X1 U1044 ( .A(n1036), .ZN(n1013) );
  NOR2_X1 U1045 ( .A1(n1019), .A2(n1020), .ZN(n1036) );
  NAND2_X1 U1046 ( .A1(b_1_), .A2(a_6_), .ZN(n1020) );
  NAND2_X1 U1047 ( .A1(a_7_), .A2(b_0_), .ZN(n1019) );
  NOR2_X1 U1048 ( .A1(n537), .A2(n682), .ZN(n1004) );
  NOR2_X1 U1049 ( .A1(n537), .A2(n657), .ZN(n1023) );
  NOR2_X1 U1050 ( .A1(n657), .A2(n694), .ZN(n988) );
  NAND2_X1 U1051 ( .A1(b_1_), .A2(a_2_), .ZN(n1025) );
  INV_X1 U1052 ( .A(n521), .ZN(n526) );
  NAND2_X1 U1053 ( .A1(n1037), .A2(n1038), .ZN(n521) );
  NAND2_X1 U1054 ( .A1(n1039), .A2(n547), .ZN(n1038) );
  NAND2_X1 U1055 ( .A1(b_0_), .A2(n716), .ZN(n547) );
  INV_X1 U1056 ( .A(a_0_), .ZN(n716) );
  NAND2_X1 U1057 ( .A1(n1040), .A2(n1041), .ZN(n1039) );
  NAND2_X1 U1058 ( .A1(a_1_), .A2(n537), .ZN(n1041) );
  NAND2_X1 U1059 ( .A1(n1042), .A2(n1043), .ZN(n1040) );
  NAND2_X1 U1060 ( .A1(b_2_), .A2(n669), .ZN(n1043) );
  INV_X1 U1061 ( .A(a_2_), .ZN(n669) );
  NOR2_X1 U1062 ( .A1(n1044), .A2(n1045), .ZN(n1042) );
  NOR2_X1 U1063 ( .A1(a_1_), .A2(n537), .ZN(n1045) );
  INV_X1 U1064 ( .A(b_1_), .ZN(n537) );
  NOR2_X1 U1065 ( .A1(n1046), .A2(n1047), .ZN(n1044) );
  NAND2_X1 U1066 ( .A1(n1048), .A2(n1049), .ZN(n1047) );
  NAND2_X1 U1067 ( .A1(n1050), .A2(n1051), .ZN(n1049) );
  NAND2_X1 U1068 ( .A1(b_4_), .A2(n682), .ZN(n1051) );
  INV_X1 U1069 ( .A(a_4_), .ZN(n682) );
  NOR2_X1 U1070 ( .A1(n1052), .A2(n1053), .ZN(n1050) );
  NOR2_X1 U1071 ( .A1(a_3_), .A2(n683), .ZN(n1053) );
  INV_X1 U1072 ( .A(b_3_), .ZN(n683) );
  NOR2_X1 U1073 ( .A1(n1054), .A2(n1055), .ZN(n1052) );
  NAND2_X1 U1074 ( .A1(n1056), .A2(n1057), .ZN(n1055) );
  NAND2_X1 U1075 ( .A1(n1058), .A2(n1059), .ZN(n1057) );
  NAND2_X1 U1076 ( .A1(b_5_), .A2(n620), .ZN(n1059) );
  NOR2_X1 U1077 ( .A1(n1060), .A2(n1061), .ZN(n1058) );
  NOR2_X1 U1078 ( .A1(a_6_), .A2(n1062), .ZN(n1061) );
  NOR2_X1 U1079 ( .A1(n1063), .A2(n602), .ZN(n1060) );
  INV_X1 U1080 ( .A(b_6_), .ZN(n602) );
  NOR2_X1 U1081 ( .A1(n592), .A2(n605), .ZN(n1063) );
  INV_X1 U1082 ( .A(a_6_), .ZN(n605) );
  INV_X1 U1083 ( .A(n1062), .ZN(n592) );
  NOR2_X1 U1084 ( .A1(n594), .A2(b_7_), .ZN(n1062) );
  INV_X1 U1085 ( .A(a_7_), .ZN(n594) );
  NAND2_X1 U1086 ( .A1(a_4_), .A2(n681), .ZN(n1056) );
  INV_X1 U1087 ( .A(b_4_), .ZN(n681) );
  NOR2_X1 U1088 ( .A1(b_5_), .A2(n620), .ZN(n1054) );
  INV_X1 U1089 ( .A(a_5_), .ZN(n620) );
  NAND2_X1 U1090 ( .A1(a_2_), .A2(n668), .ZN(n1048) );
  INV_X1 U1091 ( .A(b_2_), .ZN(n668) );
  NOR2_X1 U1092 ( .A1(b_3_), .A2(n657), .ZN(n1046) );
  INV_X1 U1093 ( .A(a_3_), .ZN(n657) );
  NAND2_X1 U1094 ( .A1(a_0_), .A2(n694), .ZN(n1037) );
  INV_X1 U1095 ( .A(b_0_), .ZN(n694) );
endmodule

