module add_mul_comp_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, 
        a_18_, a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, 
        a_28_, a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, 
        b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, 
        b_17_, b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, 
        b_27_, b_28_, b_29_, b_30_, b_31_, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151;

  OR2_X1 U7557 ( .A1(n8036), .A2(n7535), .ZN(n7493) );
  INV_X1 U7558 ( .A(n7493), .ZN(n7494) );
  INV_X2 U7559 ( .A(b_25_), .ZN(n7609) );
  INV_X2 U7560 ( .A(b_7_), .ZN(n7874) );
  INV_X2 U7561 ( .A(b_27_), .ZN(n7582) );
  INV_X2 U7562 ( .A(b_16_), .ZN(n11315) );
  INV_X2 U7563 ( .A(b_5_), .ZN(n7901) );
  INV_X2 U7564 ( .A(b_22_), .ZN(n9968) );
  INV_X2 U7565 ( .A(b_4_), .ZN(n8054) );
  INV_X2 U7566 ( .A(a_1_), .ZN(n7957) );
  INV_X2 U7567 ( .A(a_24_), .ZN(n8041) );
  INV_X2 U7568 ( .A(a_18_), .ZN(n8047) );
  INV_X2 U7569 ( .A(a_20_), .ZN(n8044) );
  INV_X2 U7570 ( .A(a_25_), .ZN(n8039) );
  INV_X2 U7571 ( .A(a_23_), .ZN(n8042) );
  INV_X2 U7572 ( .A(a_17_), .ZN(n7732) );
  NAND2_X2 U7573 ( .A1(a_30_), .A2(n8036), .ZN(n7531) );
  NAND2_X2 U7574 ( .A1(a_31_), .A2(n7535), .ZN(n7527) );
  INV_X2 U7575 ( .A(a_21_), .ZN(n7665) );
  INV_X4 U7576 ( .A(n7519), .ZN(n7495) );
  NAND2_X2 U7577 ( .A1(n15059), .A2(n15060), .ZN(n7519) );
  INV_X2 U7578 ( .A(a_29_), .ZN(n7545) );
  NOR2_X1 U7579 ( .A1(n7495), .A2(n7496), .ZN(Result_9_) );
  XOR2_X1 U7580 ( .A(n7497), .B(n7498), .Z(n7496) );
  NAND2_X1 U7581 ( .A1(n7499), .A2(n7500), .ZN(n7498) );
  NOR2_X1 U7582 ( .A1(n7495), .A2(n7501), .ZN(Result_8_) );
  XOR2_X1 U7583 ( .A(n7502), .B(n7503), .Z(n7501) );
  NAND2_X1 U7584 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
  NOR2_X1 U7585 ( .A1(n7495), .A2(n7506), .ZN(Result_7_) );
  XOR2_X1 U7586 ( .A(n7507), .B(n7508), .Z(n7506) );
  NAND2_X1 U7587 ( .A1(n7509), .A2(n7510), .ZN(n7508) );
  NOR2_X1 U7588 ( .A1(n7495), .A2(n7511), .ZN(Result_6_) );
  XOR2_X1 U7589 ( .A(n7512), .B(n7513), .Z(n7511) );
  NAND2_X1 U7590 ( .A1(n7514), .A2(n7515), .ZN(n7513) );
  NAND2_X1 U7591 ( .A1(n7516), .A2(n7517), .ZN(Result_63_) );
  NAND2_X1 U7592 ( .A1(n7518), .A2(n7519), .ZN(n7517) );
  NAND2_X1 U7593 ( .A1(n7520), .A2(n7495), .ZN(n7516) );
  XOR2_X1 U7594 ( .A(b_31_), .B(a_31_), .Z(n7520) );
  NAND2_X1 U7595 ( .A1(n7521), .A2(n7522), .ZN(Result_62_) );
  NAND2_X1 U7596 ( .A1(n7523), .A2(n7519), .ZN(n7522) );
  NAND2_X1 U7597 ( .A1(n7524), .A2(n7525), .ZN(n7523) );
  NAND2_X1 U7598 ( .A1(b_30_), .A2(n7526), .ZN(n7525) );
  NAND2_X1 U7599 ( .A1(n7527), .A2(n7528), .ZN(n7526) );
  NAND2_X1 U7600 ( .A1(a_31_), .A2(n7529), .ZN(n7528) );
  NAND2_X1 U7601 ( .A1(b_31_), .A2(n7530), .ZN(n7524) );
  NAND2_X1 U7602 ( .A1(n7531), .A2(n7532), .ZN(n7530) );
  NAND2_X1 U7603 ( .A1(n7533), .A2(n7495), .ZN(n7521) );
  XNOR2_X1 U7604 ( .A(n7518), .B(n7534), .ZN(n7533) );
  XOR2_X1 U7605 ( .A(n7535), .B(b_30_), .Z(n7534) );
  NAND2_X1 U7606 ( .A1(n7536), .A2(n7537), .ZN(Result_61_) );
  NAND2_X1 U7607 ( .A1(n7495), .A2(n7538), .ZN(n7537) );
  NAND3_X1 U7608 ( .A1(n7539), .A2(n7540), .A3(n7541), .ZN(n7538) );
  NAND2_X1 U7609 ( .A1(n7542), .A2(n7543), .ZN(n7541) );
  NAND3_X1 U7610 ( .A1(n7544), .A2(n7545), .A3(b_29_), .ZN(n7540) );
  NAND2_X1 U7611 ( .A1(n7546), .A2(n7547), .ZN(n7539) );
  XOR2_X1 U7612 ( .A(n7545), .B(n7544), .Z(n7546) );
  INV_X1 U7613 ( .A(n7543), .ZN(n7544) );
  NAND2_X1 U7614 ( .A1(n7548), .A2(n7519), .ZN(n7536) );
  XOR2_X1 U7615 ( .A(n7549), .B(n7550), .Z(n7548) );
  NOR2_X1 U7616 ( .A1(n7529), .A2(n7545), .ZN(n7550) );
  XOR2_X1 U7617 ( .A(n7551), .B(n7552), .Z(n7549) );
  NAND2_X1 U7618 ( .A1(n7553), .A2(n7554), .ZN(Result_60_) );
  NAND2_X1 U7619 ( .A1(n7555), .A2(n7519), .ZN(n7554) );
  XOR2_X1 U7620 ( .A(n7556), .B(n7557), .Z(n7555) );
  XOR2_X1 U7621 ( .A(n7558), .B(n7559), .Z(n7557) );
  NOR2_X1 U7622 ( .A1(n7529), .A2(n7560), .ZN(n7559) );
  NAND2_X1 U7623 ( .A1(n7495), .A2(n7561), .ZN(n7553) );
  XNOR2_X1 U7624 ( .A(n7562), .B(n7563), .ZN(n7561) );
  NAND2_X1 U7625 ( .A1(n7564), .A2(n7565), .ZN(n7562) );
  NOR2_X1 U7626 ( .A1(n7495), .A2(n7566), .ZN(Result_5_) );
  XOR2_X1 U7627 ( .A(n7567), .B(n7568), .Z(n7566) );
  NAND2_X1 U7628 ( .A1(n7569), .A2(n7570), .ZN(n7568) );
  NAND2_X1 U7629 ( .A1(n7571), .A2(n7572), .ZN(Result_59_) );
  NAND2_X1 U7630 ( .A1(n7495), .A2(n7573), .ZN(n7572) );
  NAND3_X1 U7631 ( .A1(n7574), .A2(n7575), .A3(n7576), .ZN(n7573) );
  NAND2_X1 U7632 ( .A1(n7577), .A2(n7578), .ZN(n7576) );
  NAND3_X1 U7633 ( .A1(n7579), .A2(n7580), .A3(b_27_), .ZN(n7575) );
  NAND2_X1 U7634 ( .A1(n7581), .A2(n7582), .ZN(n7574) );
  XOR2_X1 U7635 ( .A(n7580), .B(n7579), .Z(n7581) );
  INV_X1 U7636 ( .A(n7578), .ZN(n7579) );
  NAND2_X1 U7637 ( .A1(n7583), .A2(n7519), .ZN(n7571) );
  XNOR2_X1 U7638 ( .A(n7584), .B(n7585), .ZN(n7583) );
  NAND2_X1 U7639 ( .A1(n7586), .A2(n7587), .ZN(n7584) );
  NAND2_X1 U7640 ( .A1(n7588), .A2(n7589), .ZN(Result_58_) );
  NAND2_X1 U7641 ( .A1(n7590), .A2(n7519), .ZN(n7589) );
  XOR2_X1 U7642 ( .A(n7591), .B(n7592), .Z(n7590) );
  XOR2_X1 U7643 ( .A(n7593), .B(n7594), .Z(n7591) );
  NOR2_X1 U7644 ( .A1(n7529), .A2(n7595), .ZN(n7594) );
  NAND2_X1 U7645 ( .A1(n7495), .A2(n7596), .ZN(n7588) );
  XOR2_X1 U7646 ( .A(n7597), .B(n7598), .Z(n7596) );
  AND2_X1 U7647 ( .A1(n7599), .A2(n7600), .ZN(n7598) );
  NAND2_X1 U7648 ( .A1(n7601), .A2(n7602), .ZN(Result_57_) );
  NAND2_X1 U7649 ( .A1(n7495), .A2(n7603), .ZN(n7602) );
  NAND3_X1 U7650 ( .A1(n7604), .A2(n7605), .A3(n7606), .ZN(n7603) );
  NAND2_X1 U7651 ( .A1(n7607), .A2(n7608), .ZN(n7606) );
  OR3_X1 U7652 ( .A1(n7608), .A2(a_25_), .A3(n7609), .ZN(n7605) );
  NAND2_X1 U7653 ( .A1(n7610), .A2(n7609), .ZN(n7604) );
  XOR2_X1 U7654 ( .A(n7608), .B(a_25_), .Z(n7610) );
  NAND2_X1 U7655 ( .A1(n7611), .A2(n7519), .ZN(n7601) );
  XNOR2_X1 U7656 ( .A(n7612), .B(n7613), .ZN(n7611) );
  NAND2_X1 U7657 ( .A1(n7614), .A2(n7615), .ZN(n7612) );
  NAND2_X1 U7658 ( .A1(n7616), .A2(n7617), .ZN(Result_56_) );
  NAND2_X1 U7659 ( .A1(n7618), .A2(n7519), .ZN(n7617) );
  XOR2_X1 U7660 ( .A(n7619), .B(n7620), .Z(n7618) );
  XNOR2_X1 U7661 ( .A(n7621), .B(n7622), .ZN(n7620) );
  NAND2_X1 U7662 ( .A1(a_24_), .A2(b_31_), .ZN(n7621) );
  NAND2_X1 U7663 ( .A1(n7495), .A2(n7623), .ZN(n7616) );
  XOR2_X1 U7664 ( .A(n7624), .B(n7625), .Z(n7623) );
  AND2_X1 U7665 ( .A1(n7626), .A2(n7627), .ZN(n7625) );
  NAND2_X1 U7666 ( .A1(n7628), .A2(n7629), .ZN(Result_55_) );
  NAND2_X1 U7667 ( .A1(n7495), .A2(n7630), .ZN(n7629) );
  NAND3_X1 U7668 ( .A1(n7631), .A2(n7632), .A3(n7633), .ZN(n7630) );
  NAND2_X1 U7669 ( .A1(n7634), .A2(n7635), .ZN(n7633) );
  OR3_X1 U7670 ( .A1(n7635), .A2(a_23_), .A3(n7636), .ZN(n7632) );
  NAND2_X1 U7671 ( .A1(n7637), .A2(n7636), .ZN(n7631) );
  XOR2_X1 U7672 ( .A(n7635), .B(a_23_), .Z(n7637) );
  NAND2_X1 U7673 ( .A1(n7638), .A2(n7519), .ZN(n7628) );
  XNOR2_X1 U7674 ( .A(n7639), .B(n7640), .ZN(n7638) );
  NAND2_X1 U7675 ( .A1(n7641), .A2(n7642), .ZN(n7639) );
  NAND2_X1 U7676 ( .A1(n7643), .A2(n7644), .ZN(Result_54_) );
  NAND2_X1 U7677 ( .A1(n7645), .A2(n7519), .ZN(n7644) );
  XOR2_X1 U7678 ( .A(n7646), .B(n7647), .Z(n7645) );
  XOR2_X1 U7679 ( .A(n7648), .B(n7649), .Z(n7647) );
  NOR2_X1 U7680 ( .A1(n7529), .A2(n7650), .ZN(n7649) );
  NAND2_X1 U7681 ( .A1(n7495), .A2(n7651), .ZN(n7643) );
  XNOR2_X1 U7682 ( .A(n7652), .B(n7653), .ZN(n7651) );
  NOR2_X1 U7683 ( .A1(n7654), .A2(n7655), .ZN(n7653) );
  NAND2_X1 U7684 ( .A1(n7656), .A2(n7657), .ZN(Result_53_) );
  NAND2_X1 U7685 ( .A1(n7495), .A2(n7658), .ZN(n7657) );
  NAND3_X1 U7686 ( .A1(n7659), .A2(n7660), .A3(n7661), .ZN(n7658) );
  NAND2_X1 U7687 ( .A1(n7662), .A2(n7663), .ZN(n7661) );
  NAND3_X1 U7688 ( .A1(n7664), .A2(n7665), .A3(b_21_), .ZN(n7660) );
  NAND2_X1 U7689 ( .A1(n7666), .A2(n7667), .ZN(n7659) );
  XOR2_X1 U7690 ( .A(n7663), .B(a_21_), .Z(n7666) );
  NAND2_X1 U7691 ( .A1(n7668), .A2(n7519), .ZN(n7656) );
  XOR2_X1 U7692 ( .A(n7669), .B(n7670), .Z(n7668) );
  XNOR2_X1 U7693 ( .A(n7671), .B(n7672), .ZN(n7670) );
  NAND2_X1 U7694 ( .A1(a_21_), .A2(b_31_), .ZN(n7672) );
  NAND2_X1 U7695 ( .A1(n7673), .A2(n7674), .ZN(Result_52_) );
  NAND2_X1 U7696 ( .A1(n7675), .A2(n7519), .ZN(n7674) );
  XOR2_X1 U7697 ( .A(n7676), .B(n7677), .Z(n7675) );
  XNOR2_X1 U7698 ( .A(n7678), .B(n7679), .ZN(n7677) );
  NAND2_X1 U7699 ( .A1(a_20_), .A2(b_31_), .ZN(n7679) );
  NAND2_X1 U7700 ( .A1(n7495), .A2(n7680), .ZN(n7673) );
  XOR2_X1 U7701 ( .A(n7681), .B(n7682), .Z(n7680) );
  AND2_X1 U7702 ( .A1(n7683), .A2(n7684), .ZN(n7682) );
  NAND2_X1 U7703 ( .A1(n7685), .A2(n7686), .ZN(Result_51_) );
  NAND2_X1 U7704 ( .A1(n7495), .A2(n7687), .ZN(n7686) );
  NAND3_X1 U7705 ( .A1(n7688), .A2(n7689), .A3(n7690), .ZN(n7687) );
  NAND2_X1 U7706 ( .A1(n7691), .A2(n7692), .ZN(n7690) );
  OR3_X1 U7707 ( .A1(n7692), .A2(a_19_), .A3(n7693), .ZN(n7689) );
  NAND2_X1 U7708 ( .A1(n7694), .A2(n7693), .ZN(n7688) );
  XOR2_X1 U7709 ( .A(n7692), .B(a_19_), .Z(n7694) );
  NAND2_X1 U7710 ( .A1(n7695), .A2(n7519), .ZN(n7685) );
  XNOR2_X1 U7711 ( .A(n7696), .B(n7697), .ZN(n7695) );
  XOR2_X1 U7712 ( .A(n7698), .B(n7699), .Z(n7697) );
  NAND2_X1 U7713 ( .A1(a_19_), .A2(b_31_), .ZN(n7699) );
  NAND2_X1 U7714 ( .A1(n7700), .A2(n7701), .ZN(Result_50_) );
  NAND2_X1 U7715 ( .A1(n7702), .A2(n7519), .ZN(n7701) );
  XOR2_X1 U7716 ( .A(n7703), .B(n7704), .Z(n7702) );
  XNOR2_X1 U7717 ( .A(n7705), .B(n7706), .ZN(n7704) );
  NAND2_X1 U7718 ( .A1(a_18_), .A2(b_31_), .ZN(n7706) );
  NAND2_X1 U7719 ( .A1(n7495), .A2(n7707), .ZN(n7700) );
  XOR2_X1 U7720 ( .A(n7708), .B(n7709), .Z(n7707) );
  AND2_X1 U7721 ( .A1(n7710), .A2(n7711), .ZN(n7709) );
  NOR2_X1 U7722 ( .A1(n7495), .A2(n7712), .ZN(Result_4_) );
  XOR2_X1 U7723 ( .A(n7713), .B(n7714), .Z(n7712) );
  NAND2_X1 U7724 ( .A1(n7715), .A2(n7716), .ZN(n7714) );
  NAND2_X1 U7725 ( .A1(n7717), .A2(n7718), .ZN(Result_49_) );
  NAND2_X1 U7726 ( .A1(n7495), .A2(n7719), .ZN(n7718) );
  NAND3_X1 U7727 ( .A1(n7720), .A2(n7721), .A3(n7722), .ZN(n7719) );
  NAND2_X1 U7728 ( .A1(n7723), .A2(n7724), .ZN(n7722) );
  OR3_X1 U7729 ( .A1(n7724), .A2(a_17_), .A3(n7725), .ZN(n7721) );
  NAND2_X1 U7730 ( .A1(n7726), .A2(n7725), .ZN(n7720) );
  XOR2_X1 U7731 ( .A(n7724), .B(a_17_), .Z(n7726) );
  NAND2_X1 U7732 ( .A1(n7727), .A2(n7519), .ZN(n7717) );
  XOR2_X1 U7733 ( .A(n7728), .B(n7729), .Z(n7727) );
  XOR2_X1 U7734 ( .A(n7730), .B(n7731), .Z(n7728) );
  NOR2_X1 U7735 ( .A1(n7529), .A2(n7732), .ZN(n7731) );
  NAND2_X1 U7736 ( .A1(n7733), .A2(n7734), .ZN(Result_48_) );
  NAND2_X1 U7737 ( .A1(n7735), .A2(n7519), .ZN(n7734) );
  XOR2_X1 U7738 ( .A(n7736), .B(n7737), .Z(n7735) );
  XNOR2_X1 U7739 ( .A(n7738), .B(n7739), .ZN(n7737) );
  NAND2_X1 U7740 ( .A1(a_16_), .A2(b_31_), .ZN(n7739) );
  NAND2_X1 U7741 ( .A1(n7495), .A2(n7740), .ZN(n7733) );
  XNOR2_X1 U7742 ( .A(n7741), .B(n7742), .ZN(n7740) );
  NOR2_X1 U7743 ( .A1(n7743), .A2(n7744), .ZN(n7742) );
  NAND2_X1 U7744 ( .A1(n7745), .A2(n7746), .ZN(Result_47_) );
  NAND2_X1 U7745 ( .A1(n7495), .A2(n7747), .ZN(n7746) );
  NAND3_X1 U7746 ( .A1(n7748), .A2(n7749), .A3(n7750), .ZN(n7747) );
  NAND2_X1 U7747 ( .A1(n7751), .A2(n7752), .ZN(n7750) );
  NAND3_X1 U7748 ( .A1(n7753), .A2(n7754), .A3(b_15_), .ZN(n7749) );
  NAND2_X1 U7749 ( .A1(n7755), .A2(n7756), .ZN(n7748) );
  XOR2_X1 U7750 ( .A(n7752), .B(a_15_), .Z(n7755) );
  NAND2_X1 U7751 ( .A1(n7757), .A2(n7519), .ZN(n7745) );
  XNOR2_X1 U7752 ( .A(n7758), .B(n7759), .ZN(n7757) );
  XOR2_X1 U7753 ( .A(n7760), .B(n7761), .Z(n7759) );
  NAND2_X1 U7754 ( .A1(a_15_), .A2(b_31_), .ZN(n7761) );
  NAND2_X1 U7755 ( .A1(n7762), .A2(n7763), .ZN(Result_46_) );
  NAND2_X1 U7756 ( .A1(n7764), .A2(n7519), .ZN(n7763) );
  XOR2_X1 U7757 ( .A(n7765), .B(n7766), .Z(n7764) );
  XNOR2_X1 U7758 ( .A(n7767), .B(n7768), .ZN(n7766) );
  NAND2_X1 U7759 ( .A1(a_14_), .A2(b_31_), .ZN(n7768) );
  NAND2_X1 U7760 ( .A1(n7495), .A2(n7769), .ZN(n7762) );
  XOR2_X1 U7761 ( .A(n7770), .B(n7771), .Z(n7769) );
  AND2_X1 U7762 ( .A1(n7772), .A2(n7773), .ZN(n7771) );
  NAND2_X1 U7763 ( .A1(n7774), .A2(n7775), .ZN(Result_45_) );
  NAND2_X1 U7764 ( .A1(n7495), .A2(n7776), .ZN(n7775) );
  NAND3_X1 U7765 ( .A1(n7777), .A2(n7778), .A3(n7779), .ZN(n7776) );
  NAND2_X1 U7766 ( .A1(n7780), .A2(n7781), .ZN(n7779) );
  OR3_X1 U7767 ( .A1(n7781), .A2(a_13_), .A3(n7782), .ZN(n7778) );
  NAND2_X1 U7768 ( .A1(n7783), .A2(n7782), .ZN(n7777) );
  XOR2_X1 U7769 ( .A(n7781), .B(a_13_), .Z(n7783) );
  NAND2_X1 U7770 ( .A1(n7784), .A2(n7519), .ZN(n7774) );
  XOR2_X1 U7771 ( .A(n7785), .B(n7786), .Z(n7784) );
  XOR2_X1 U7772 ( .A(n7787), .B(n7788), .Z(n7785) );
  NOR2_X1 U7773 ( .A1(n7529), .A2(n7789), .ZN(n7788) );
  NAND2_X1 U7774 ( .A1(n7790), .A2(n7791), .ZN(Result_44_) );
  NAND2_X1 U7775 ( .A1(n7792), .A2(n7519), .ZN(n7791) );
  XOR2_X1 U7776 ( .A(n7793), .B(n7794), .Z(n7792) );
  XNOR2_X1 U7777 ( .A(n7795), .B(n7796), .ZN(n7794) );
  NAND2_X1 U7778 ( .A1(a_12_), .A2(b_31_), .ZN(n7796) );
  NAND2_X1 U7779 ( .A1(n7495), .A2(n7797), .ZN(n7790) );
  XNOR2_X1 U7780 ( .A(n7798), .B(n7799), .ZN(n7797) );
  NOR2_X1 U7781 ( .A1(n7800), .A2(n7801), .ZN(n7799) );
  NAND2_X1 U7782 ( .A1(n7802), .A2(n7803), .ZN(Result_43_) );
  NAND2_X1 U7783 ( .A1(n7495), .A2(n7804), .ZN(n7803) );
  NAND3_X1 U7784 ( .A1(n7805), .A2(n7806), .A3(n7807), .ZN(n7804) );
  NAND2_X1 U7785 ( .A1(n7808), .A2(n7809), .ZN(n7807) );
  NAND3_X1 U7786 ( .A1(n7810), .A2(n7811), .A3(b_11_), .ZN(n7806) );
  NAND2_X1 U7787 ( .A1(n7812), .A2(n7813), .ZN(n7805) );
  XOR2_X1 U7788 ( .A(n7809), .B(a_11_), .Z(n7812) );
  NAND2_X1 U7789 ( .A1(n7814), .A2(n7519), .ZN(n7802) );
  XNOR2_X1 U7790 ( .A(n7815), .B(n7816), .ZN(n7814) );
  XOR2_X1 U7791 ( .A(n7817), .B(n7818), .Z(n7816) );
  NAND2_X1 U7792 ( .A1(a_11_), .A2(b_31_), .ZN(n7818) );
  NAND2_X1 U7793 ( .A1(n7819), .A2(n7820), .ZN(Result_42_) );
  NAND2_X1 U7794 ( .A1(n7821), .A2(n7519), .ZN(n7820) );
  XOR2_X1 U7795 ( .A(n7822), .B(n7823), .Z(n7821) );
  XNOR2_X1 U7796 ( .A(n7824), .B(n7825), .ZN(n7823) );
  NAND2_X1 U7797 ( .A1(a_10_), .A2(b_31_), .ZN(n7825) );
  NAND2_X1 U7798 ( .A1(n7495), .A2(n7826), .ZN(n7819) );
  XOR2_X1 U7799 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND2_X1 U7800 ( .A1(n7829), .A2(n7830), .ZN(n7828) );
  NAND2_X1 U7801 ( .A1(n7831), .A2(n7832), .ZN(Result_41_) );
  NAND2_X1 U7802 ( .A1(n7495), .A2(n7833), .ZN(n7832) );
  NAND3_X1 U7803 ( .A1(n7834), .A2(n7835), .A3(n7836), .ZN(n7833) );
  NAND2_X1 U7804 ( .A1(n7837), .A2(n7838), .ZN(n7836) );
  OR3_X1 U7805 ( .A1(n7838), .A2(a_9_), .A3(n7839), .ZN(n7835) );
  NAND2_X1 U7806 ( .A1(n7840), .A2(n7839), .ZN(n7834) );
  XOR2_X1 U7807 ( .A(n7838), .B(a_9_), .Z(n7840) );
  NAND2_X1 U7808 ( .A1(n7841), .A2(n7519), .ZN(n7831) );
  XOR2_X1 U7809 ( .A(n7842), .B(n7843), .Z(n7841) );
  XNOR2_X1 U7810 ( .A(n7844), .B(n7845), .ZN(n7843) );
  NAND2_X1 U7811 ( .A1(a_9_), .A2(b_31_), .ZN(n7845) );
  NAND2_X1 U7812 ( .A1(n7846), .A2(n7847), .ZN(Result_40_) );
  NAND2_X1 U7813 ( .A1(n7848), .A2(n7519), .ZN(n7847) );
  XOR2_X1 U7814 ( .A(n7849), .B(n7850), .Z(n7848) );
  XNOR2_X1 U7815 ( .A(n7851), .B(n7852), .ZN(n7850) );
  NAND2_X1 U7816 ( .A1(a_8_), .A2(b_31_), .ZN(n7852) );
  NAND2_X1 U7817 ( .A1(n7495), .A2(n7853), .ZN(n7846) );
  XNOR2_X1 U7818 ( .A(n7854), .B(n7855), .ZN(n7853) );
  NOR2_X1 U7819 ( .A1(n7856), .A2(n7857), .ZN(n7855) );
  NOR2_X1 U7820 ( .A1(n7495), .A2(n7858), .ZN(Result_3_) );
  XOR2_X1 U7821 ( .A(n7859), .B(n7860), .Z(n7858) );
  NAND2_X1 U7822 ( .A1(n7861), .A2(n7862), .ZN(n7860) );
  NAND2_X1 U7823 ( .A1(n7863), .A2(n7864), .ZN(Result_39_) );
  NAND2_X1 U7824 ( .A1(n7495), .A2(n7865), .ZN(n7864) );
  NAND3_X1 U7825 ( .A1(n7866), .A2(n7867), .A3(n7868), .ZN(n7865) );
  NAND2_X1 U7826 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
  NAND3_X1 U7827 ( .A1(n7871), .A2(n7872), .A3(b_7_), .ZN(n7867) );
  NAND2_X1 U7828 ( .A1(n7873), .A2(n7874), .ZN(n7866) );
  XOR2_X1 U7829 ( .A(n7870), .B(a_7_), .Z(n7873) );
  NAND2_X1 U7830 ( .A1(n7875), .A2(n7519), .ZN(n7863) );
  XNOR2_X1 U7831 ( .A(n7876), .B(n7877), .ZN(n7875) );
  XOR2_X1 U7832 ( .A(n7878), .B(n7879), .Z(n7877) );
  NAND2_X1 U7833 ( .A1(a_7_), .A2(b_31_), .ZN(n7879) );
  NAND2_X1 U7834 ( .A1(n7880), .A2(n7881), .ZN(Result_38_) );
  NAND2_X1 U7835 ( .A1(n7882), .A2(n7519), .ZN(n7881) );
  XOR2_X1 U7836 ( .A(n7883), .B(n7884), .Z(n7882) );
  XOR2_X1 U7837 ( .A(n7885), .B(n7886), .Z(n7883) );
  NOR2_X1 U7838 ( .A1(n7529), .A2(n7887), .ZN(n7886) );
  NAND2_X1 U7839 ( .A1(n7495), .A2(n7888), .ZN(n7880) );
  XOR2_X1 U7840 ( .A(n7889), .B(n7890), .Z(n7888) );
  AND2_X1 U7841 ( .A1(n7891), .A2(n7892), .ZN(n7890) );
  NAND2_X1 U7842 ( .A1(n7893), .A2(n7894), .ZN(Result_37_) );
  NAND2_X1 U7843 ( .A1(n7495), .A2(n7895), .ZN(n7894) );
  NAND3_X1 U7844 ( .A1(n7896), .A2(n7897), .A3(n7898), .ZN(n7895) );
  NAND2_X1 U7845 ( .A1(n7899), .A2(n7900), .ZN(n7898) );
  OR3_X1 U7846 ( .A1(n7900), .A2(a_5_), .A3(n7901), .ZN(n7897) );
  NAND2_X1 U7847 ( .A1(n7902), .A2(n7901), .ZN(n7896) );
  XOR2_X1 U7848 ( .A(n7900), .B(a_5_), .Z(n7902) );
  NAND2_X1 U7849 ( .A1(n7903), .A2(n7519), .ZN(n7893) );
  XOR2_X1 U7850 ( .A(n7904), .B(n7905), .Z(n7903) );
  XOR2_X1 U7851 ( .A(n7906), .B(n7907), .Z(n7904) );
  NOR2_X1 U7852 ( .A1(n7529), .A2(n7908), .ZN(n7907) );
  NAND2_X1 U7853 ( .A1(n7909), .A2(n7910), .ZN(Result_36_) );
  NAND2_X1 U7854 ( .A1(n7911), .A2(n7519), .ZN(n7910) );
  XOR2_X1 U7855 ( .A(n7912), .B(n7913), .Z(n7911) );
  XOR2_X1 U7856 ( .A(n7914), .B(n7915), .Z(n7912) );
  NOR2_X1 U7857 ( .A1(n7529), .A2(n7916), .ZN(n7915) );
  NAND2_X1 U7858 ( .A1(n7495), .A2(n7917), .ZN(n7909) );
  XOR2_X1 U7859 ( .A(n7918), .B(n7919), .Z(n7917) );
  AND2_X1 U7860 ( .A1(n7920), .A2(n7921), .ZN(n7919) );
  NAND2_X1 U7861 ( .A1(n7922), .A2(n7923), .ZN(Result_35_) );
  NAND2_X1 U7862 ( .A1(n7495), .A2(n7924), .ZN(n7923) );
  NAND3_X1 U7863 ( .A1(n7925), .A2(n7926), .A3(n7927), .ZN(n7924) );
  NAND2_X1 U7864 ( .A1(n7928), .A2(n7929), .ZN(n7927) );
  OR3_X1 U7865 ( .A1(n7929), .A2(a_3_), .A3(n7930), .ZN(n7926) );
  NAND2_X1 U7866 ( .A1(n7931), .A2(n7930), .ZN(n7925) );
  XOR2_X1 U7867 ( .A(n7929), .B(a_3_), .Z(n7931) );
  NAND2_X1 U7868 ( .A1(n7932), .A2(n7519), .ZN(n7922) );
  XOR2_X1 U7869 ( .A(n7933), .B(n7934), .Z(n7932) );
  XOR2_X1 U7870 ( .A(n7935), .B(n7936), .Z(n7933) );
  NOR2_X1 U7871 ( .A1(n7529), .A2(n7937), .ZN(n7936) );
  NAND2_X1 U7872 ( .A1(n7938), .A2(n7939), .ZN(Result_34_) );
  NAND2_X1 U7873 ( .A1(n7940), .A2(n7519), .ZN(n7939) );
  XOR2_X1 U7874 ( .A(n7941), .B(n7942), .Z(n7940) );
  XNOR2_X1 U7875 ( .A(n7943), .B(n7944), .ZN(n7942) );
  NAND2_X1 U7876 ( .A1(a_2_), .A2(b_31_), .ZN(n7944) );
  NAND2_X1 U7877 ( .A1(n7495), .A2(n7945), .ZN(n7938) );
  XOR2_X1 U7878 ( .A(n7946), .B(n7947), .Z(n7945) );
  AND2_X1 U7879 ( .A1(n7948), .A2(n7949), .ZN(n7947) );
  NAND2_X1 U7880 ( .A1(n7950), .A2(n7951), .ZN(Result_33_) );
  NAND2_X1 U7881 ( .A1(n7952), .A2(n7519), .ZN(n7951) );
  XOR2_X1 U7882 ( .A(n7953), .B(n7954), .Z(n7952) );
  XOR2_X1 U7883 ( .A(n7955), .B(n7956), .Z(n7953) );
  NOR2_X1 U7884 ( .A1(n7957), .A2(n7529), .ZN(n7956) );
  NAND2_X1 U7885 ( .A1(n7958), .A2(n7495), .ZN(n7950) );
  NAND2_X1 U7886 ( .A1(n7959), .A2(n7960), .ZN(n7958) );
  NAND2_X1 U7887 ( .A1(n7961), .A2(n7962), .ZN(n7960) );
  OR2_X1 U7888 ( .A1(n7963), .A2(n7964), .ZN(n7961) );
  NAND2_X1 U7889 ( .A1(n7965), .A2(n7966), .ZN(n7959) );
  INV_X1 U7890 ( .A(n7962), .ZN(n7966) );
  XOR2_X1 U7891 ( .A(b_1_), .B(a_1_), .Z(n7965) );
  NAND2_X1 U7892 ( .A1(n7967), .A2(n7968), .ZN(Result_32_) );
  NAND2_X1 U7893 ( .A1(n7969), .A2(n7519), .ZN(n7968) );
  XOR2_X1 U7894 ( .A(n7970), .B(n7971), .Z(n7969) );
  XNOR2_X1 U7895 ( .A(n7972), .B(n7973), .ZN(n7971) );
  NAND2_X1 U7896 ( .A1(a_0_), .A2(b_31_), .ZN(n7973) );
  NAND2_X1 U7897 ( .A1(n7974), .A2(n7495), .ZN(n7967) );
  XNOR2_X1 U7898 ( .A(n7975), .B(n7976), .ZN(n7974) );
  NOR2_X1 U7899 ( .A1(n7964), .A2(n7977), .ZN(n7975) );
  NOR2_X1 U7900 ( .A1(n7963), .A2(n7962), .ZN(n7977) );
  NAND2_X1 U7901 ( .A1(n7949), .A2(n7978), .ZN(n7962) );
  NAND2_X1 U7902 ( .A1(n7948), .A2(n7946), .ZN(n7978) );
  NAND2_X1 U7903 ( .A1(n7979), .A2(n7980), .ZN(n7946) );
  NAND2_X1 U7904 ( .A1(n7981), .A2(n7929), .ZN(n7980) );
  NAND2_X1 U7905 ( .A1(n7921), .A2(n7982), .ZN(n7929) );
  NAND2_X1 U7906 ( .A1(n7920), .A2(n7918), .ZN(n7982) );
  NAND2_X1 U7907 ( .A1(n7983), .A2(n7984), .ZN(n7918) );
  NAND2_X1 U7908 ( .A1(n7985), .A2(n7900), .ZN(n7984) );
  NAND2_X1 U7909 ( .A1(n7892), .A2(n7986), .ZN(n7900) );
  NAND2_X1 U7910 ( .A1(n7891), .A2(n7889), .ZN(n7986) );
  NAND2_X1 U7911 ( .A1(n7987), .A2(n7988), .ZN(n7889) );
  NAND2_X1 U7912 ( .A1(n7989), .A2(n7870), .ZN(n7988) );
  INV_X1 U7913 ( .A(n7871), .ZN(n7870) );
  NOR2_X1 U7914 ( .A1(n7857), .A2(n7990), .ZN(n7871) );
  NOR2_X1 U7915 ( .A1(n7856), .A2(n7854), .ZN(n7990) );
  AND2_X1 U7916 ( .A1(n7991), .A2(n7992), .ZN(n7854) );
  NAND2_X1 U7917 ( .A1(n7993), .A2(n7838), .ZN(n7992) );
  NAND2_X1 U7918 ( .A1(n7830), .A2(n7994), .ZN(n7838) );
  NAND2_X1 U7919 ( .A1(n7829), .A2(n7827), .ZN(n7994) );
  NAND2_X1 U7920 ( .A1(n7995), .A2(n7996), .ZN(n7827) );
  NAND2_X1 U7921 ( .A1(n7997), .A2(n7809), .ZN(n7996) );
  INV_X1 U7922 ( .A(n7810), .ZN(n7809) );
  NOR2_X1 U7923 ( .A1(n7801), .A2(n7998), .ZN(n7810) );
  NOR2_X1 U7924 ( .A1(n7800), .A2(n7798), .ZN(n7998) );
  AND2_X1 U7925 ( .A1(n7999), .A2(n8000), .ZN(n7798) );
  NAND2_X1 U7926 ( .A1(n8001), .A2(n7781), .ZN(n8000) );
  NAND2_X1 U7927 ( .A1(n7773), .A2(n8002), .ZN(n7781) );
  NAND2_X1 U7928 ( .A1(n7772), .A2(n7770), .ZN(n8002) );
  NAND2_X1 U7929 ( .A1(n8003), .A2(n8004), .ZN(n7770) );
  NAND2_X1 U7930 ( .A1(n8005), .A2(n7752), .ZN(n8004) );
  INV_X1 U7931 ( .A(n7753), .ZN(n7752) );
  NOR2_X1 U7932 ( .A1(n7744), .A2(n8006), .ZN(n7753) );
  NOR2_X1 U7933 ( .A1(n7743), .A2(n7741), .ZN(n8006) );
  AND2_X1 U7934 ( .A1(n8007), .A2(n8008), .ZN(n7741) );
  NAND2_X1 U7935 ( .A1(n8009), .A2(n7724), .ZN(n8008) );
  NAND2_X1 U7936 ( .A1(n7711), .A2(n8010), .ZN(n7724) );
  NAND2_X1 U7937 ( .A1(n7710), .A2(n7708), .ZN(n8010) );
  NAND2_X1 U7938 ( .A1(n8011), .A2(n8012), .ZN(n7708) );
  NAND2_X1 U7939 ( .A1(n8013), .A2(n7692), .ZN(n8012) );
  NAND2_X1 U7940 ( .A1(n7684), .A2(n8014), .ZN(n7692) );
  NAND2_X1 U7941 ( .A1(n7683), .A2(n7681), .ZN(n8014) );
  NAND2_X1 U7942 ( .A1(n8015), .A2(n8016), .ZN(n7681) );
  NAND2_X1 U7943 ( .A1(n8017), .A2(n7663), .ZN(n8016) );
  INV_X1 U7944 ( .A(n7664), .ZN(n7663) );
  NOR2_X1 U7945 ( .A1(n7655), .A2(n8018), .ZN(n7664) );
  NOR2_X1 U7946 ( .A1(n7654), .A2(n7652), .ZN(n8018) );
  NOR2_X1 U7947 ( .A1(n7634), .A2(n8019), .ZN(n7652) );
  AND2_X1 U7948 ( .A1(n8020), .A2(n7635), .ZN(n8019) );
  NAND2_X1 U7949 ( .A1(n7627), .A2(n8021), .ZN(n7635) );
  NAND2_X1 U7950 ( .A1(n7626), .A2(n7624), .ZN(n8021) );
  NAND2_X1 U7951 ( .A1(n8022), .A2(n8023), .ZN(n7624) );
  NAND2_X1 U7952 ( .A1(n8024), .A2(n7608), .ZN(n8023) );
  NAND2_X1 U7953 ( .A1(n7600), .A2(n8025), .ZN(n7608) );
  NAND2_X1 U7954 ( .A1(n7599), .A2(n7597), .ZN(n8025) );
  NAND2_X1 U7955 ( .A1(n8026), .A2(n8027), .ZN(n7597) );
  NAND2_X1 U7956 ( .A1(n8028), .A2(n7578), .ZN(n8027) );
  NAND2_X1 U7957 ( .A1(n7564), .A2(n8029), .ZN(n7578) );
  NAND2_X1 U7958 ( .A1(n7565), .A2(n7563), .ZN(n8029) );
  NAND2_X1 U7959 ( .A1(n8030), .A2(n8031), .ZN(n7563) );
  NAND2_X1 U7960 ( .A1(n8032), .A2(n7543), .ZN(n8031) );
  NAND2_X1 U7961 ( .A1(n8033), .A2(n8034), .ZN(n7543) );
  NAND2_X1 U7962 ( .A1(b_30_), .A2(n8035), .ZN(n8034) );
  OR2_X1 U7963 ( .A1(a_30_), .A2(n7518), .ZN(n8035) );
  NOR2_X1 U7964 ( .A1(n8036), .A2(n7529), .ZN(n7518) );
  INV_X1 U7965 ( .A(b_31_), .ZN(n7529) );
  NAND2_X1 U7966 ( .A1(n7494), .A2(b_31_), .ZN(n8033) );
  NAND2_X1 U7967 ( .A1(n7547), .A2(n7545), .ZN(n8032) );
  NAND2_X1 U7968 ( .A1(n8037), .A2(n7560), .ZN(n7565) );
  NAND2_X1 U7969 ( .A1(n7582), .A2(n7580), .ZN(n8028) );
  NAND2_X1 U7970 ( .A1(n8038), .A2(n7595), .ZN(n7599) );
  NAND2_X1 U7971 ( .A1(n7609), .A2(n8039), .ZN(n8024) );
  NAND2_X1 U7972 ( .A1(n8040), .A2(n8041), .ZN(n7626) );
  NAND2_X1 U7973 ( .A1(n7636), .A2(n8042), .ZN(n8020) );
  NOR2_X1 U7974 ( .A1(b_22_), .A2(a_22_), .ZN(n7654) );
  NAND2_X1 U7975 ( .A1(n7667), .A2(n7665), .ZN(n8017) );
  NAND2_X1 U7976 ( .A1(n8043), .A2(n8044), .ZN(n7683) );
  NAND2_X1 U7977 ( .A1(n7693), .A2(n8045), .ZN(n8013) );
  NAND2_X1 U7978 ( .A1(n8046), .A2(n8047), .ZN(n7710) );
  NAND2_X1 U7979 ( .A1(n7725), .A2(n7732), .ZN(n8009) );
  NOR2_X1 U7980 ( .A1(b_16_), .A2(a_16_), .ZN(n7743) );
  NAND2_X1 U7981 ( .A1(n7756), .A2(n7754), .ZN(n8005) );
  NAND2_X1 U7982 ( .A1(n8048), .A2(n8049), .ZN(n7772) );
  NAND2_X1 U7983 ( .A1(n7782), .A2(n7789), .ZN(n8001) );
  NOR2_X1 U7984 ( .A1(b_12_), .A2(a_12_), .ZN(n7800) );
  NAND2_X1 U7985 ( .A1(n7813), .A2(n7811), .ZN(n7997) );
  NAND2_X1 U7986 ( .A1(n8050), .A2(n8051), .ZN(n7829) );
  NAND2_X1 U7987 ( .A1(n7839), .A2(n8052), .ZN(n7993) );
  NOR2_X1 U7988 ( .A1(b_8_), .A2(a_8_), .ZN(n7856) );
  NAND2_X1 U7989 ( .A1(n7874), .A2(n7872), .ZN(n7989) );
  NAND2_X1 U7990 ( .A1(n8053), .A2(n7887), .ZN(n7891) );
  NAND2_X1 U7991 ( .A1(n7901), .A2(n7908), .ZN(n7985) );
  NAND2_X1 U7992 ( .A1(n8054), .A2(n7916), .ZN(n7920) );
  NAND2_X1 U7993 ( .A1(n7930), .A2(n7937), .ZN(n7981) );
  NAND2_X1 U7994 ( .A1(n8055), .A2(n8056), .ZN(n7948) );
  NOR2_X1 U7995 ( .A1(b_1_), .A2(a_1_), .ZN(n7964) );
  NOR2_X1 U7996 ( .A1(n7495), .A2(n8057), .ZN(Result_31_) );
  XNOR2_X1 U7997 ( .A(n8058), .B(n8059), .ZN(n8057) );
  NOR3_X1 U7998 ( .A1(n8060), .A2(n8061), .A3(n7495), .ZN(Result_30_) );
  NOR2_X1 U7999 ( .A1(n8062), .A2(n8063), .ZN(n8060) );
  AND2_X1 U8000 ( .A1(n8059), .A2(n8058), .ZN(n8062) );
  NOR2_X1 U8001 ( .A1(n7495), .A2(n8064), .ZN(Result_2_) );
  XOR2_X1 U8002 ( .A(n8065), .B(n8066), .Z(n8064) );
  NAND2_X1 U8003 ( .A1(n8067), .A2(n8068), .ZN(n8066) );
  NOR2_X1 U8004 ( .A1(n7495), .A2(n8069), .ZN(Result_29_) );
  XNOR2_X1 U8005 ( .A(n8061), .B(n8070), .ZN(n8069) );
  AND2_X1 U8006 ( .A1(n8071), .A2(n8072), .ZN(n8070) );
  NOR2_X1 U8007 ( .A1(n7495), .A2(n8073), .ZN(Result_28_) );
  XOR2_X1 U8008 ( .A(n8074), .B(n8075), .Z(n8073) );
  NOR2_X1 U8009 ( .A1(n8076), .A2(n8077), .ZN(n8075) );
  NOR2_X1 U8010 ( .A1(n7495), .A2(n8078), .ZN(Result_27_) );
  XOR2_X1 U8011 ( .A(n8079), .B(n8080), .Z(n8078) );
  NOR2_X1 U8012 ( .A1(n8081), .A2(n8082), .ZN(n8080) );
  NOR2_X1 U8013 ( .A1(n7495), .A2(n8083), .ZN(Result_26_) );
  XOR2_X1 U8014 ( .A(n8084), .B(n8085), .Z(n8083) );
  NAND2_X1 U8015 ( .A1(n8086), .A2(n8087), .ZN(n8084) );
  NOR2_X1 U8016 ( .A1(n7495), .A2(n8088), .ZN(Result_25_) );
  XOR2_X1 U8017 ( .A(n8089), .B(n8090), .Z(n8088) );
  NAND2_X1 U8018 ( .A1(n8091), .A2(n8092), .ZN(n8090) );
  NOR2_X1 U8019 ( .A1(n7495), .A2(n8093), .ZN(Result_24_) );
  XOR2_X1 U8020 ( .A(n8094), .B(n8095), .Z(n8093) );
  NAND2_X1 U8021 ( .A1(n8096), .A2(n8097), .ZN(n8095) );
  NOR2_X1 U8022 ( .A1(n7495), .A2(n8098), .ZN(Result_23_) );
  XOR2_X1 U8023 ( .A(n8099), .B(n8100), .Z(n8098) );
  NAND2_X1 U8024 ( .A1(n8101), .A2(n8102), .ZN(n8100) );
  NOR2_X1 U8025 ( .A1(n7495), .A2(n8103), .ZN(Result_22_) );
  XOR2_X1 U8026 ( .A(n8104), .B(n8105), .Z(n8103) );
  NAND2_X1 U8027 ( .A1(n8106), .A2(n8107), .ZN(n8105) );
  NOR2_X1 U8028 ( .A1(n7495), .A2(n8108), .ZN(Result_21_) );
  XOR2_X1 U8029 ( .A(n8109), .B(n8110), .Z(n8108) );
  NAND2_X1 U8030 ( .A1(n8111), .A2(n8112), .ZN(n8110) );
  NOR2_X1 U8031 ( .A1(n7495), .A2(n8113), .ZN(Result_20_) );
  XOR2_X1 U8032 ( .A(n8114), .B(n8115), .Z(n8113) );
  NAND2_X1 U8033 ( .A1(n8116), .A2(n8117), .ZN(n8115) );
  NOR2_X1 U8034 ( .A1(n7495), .A2(n8118), .ZN(Result_1_) );
  XOR2_X1 U8035 ( .A(n8119), .B(n8120), .Z(n8118) );
  NAND2_X1 U8036 ( .A1(n8121), .A2(n8122), .ZN(n8120) );
  NOR2_X1 U8037 ( .A1(n7495), .A2(n8123), .ZN(Result_19_) );
  XOR2_X1 U8038 ( .A(n8124), .B(n8125), .Z(n8123) );
  NAND2_X1 U8039 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  NOR2_X1 U8040 ( .A1(n7495), .A2(n8128), .ZN(Result_18_) );
  XOR2_X1 U8041 ( .A(n8129), .B(n8130), .Z(n8128) );
  NAND2_X1 U8042 ( .A1(n8131), .A2(n8132), .ZN(n8130) );
  NOR2_X1 U8043 ( .A1(n7495), .A2(n8133), .ZN(Result_17_) );
  XOR2_X1 U8044 ( .A(n8134), .B(n8135), .Z(n8133) );
  NAND2_X1 U8045 ( .A1(n8136), .A2(n8137), .ZN(n8135) );
  NOR2_X1 U8046 ( .A1(n7495), .A2(n8138), .ZN(Result_16_) );
  XOR2_X1 U8047 ( .A(n8139), .B(n8140), .Z(n8138) );
  NAND2_X1 U8048 ( .A1(n8141), .A2(n8142), .ZN(n8140) );
  NOR2_X1 U8049 ( .A1(n7495), .A2(n8143), .ZN(Result_15_) );
  XOR2_X1 U8050 ( .A(n8144), .B(n8145), .Z(n8143) );
  NAND2_X1 U8051 ( .A1(n8146), .A2(n8147), .ZN(n8145) );
  NOR2_X1 U8052 ( .A1(n7495), .A2(n8148), .ZN(Result_14_) );
  XOR2_X1 U8053 ( .A(n8149), .B(n8150), .Z(n8148) );
  NAND2_X1 U8054 ( .A1(n8151), .A2(n8152), .ZN(n8150) );
  NOR2_X1 U8055 ( .A1(n7495), .A2(n8153), .ZN(Result_13_) );
  XOR2_X1 U8056 ( .A(n8154), .B(n8155), .Z(n8153) );
  NAND2_X1 U8057 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  NOR2_X1 U8058 ( .A1(n7495), .A2(n8158), .ZN(Result_12_) );
  XOR2_X1 U8059 ( .A(n8159), .B(n8160), .Z(n8158) );
  NAND2_X1 U8060 ( .A1(n8161), .A2(n8162), .ZN(n8160) );
  NOR2_X1 U8061 ( .A1(n7495), .A2(n8163), .ZN(Result_11_) );
  XOR2_X1 U8062 ( .A(n8164), .B(n8165), .Z(n8163) );
  NAND2_X1 U8063 ( .A1(n8166), .A2(n8167), .ZN(n8165) );
  NOR2_X1 U8064 ( .A1(n7495), .A2(n8168), .ZN(Result_10_) );
  XOR2_X1 U8065 ( .A(n8169), .B(n8170), .Z(n8168) );
  NAND2_X1 U8066 ( .A1(n8171), .A2(n8172), .ZN(n8170) );
  NOR2_X1 U8067 ( .A1(n7495), .A2(n8173), .ZN(Result_0_) );
  AND3_X1 U8068 ( .A1(n8174), .A2(n8175), .A3(n8122), .ZN(n8173) );
  NAND4_X1 U8069 ( .A1(b_0_), .A2(n8175), .A3(n8176), .A4(n8177), .ZN(n8122)
         );
  NAND2_X1 U8070 ( .A1(n8119), .A2(n8121), .ZN(n8174) );
  NAND2_X1 U8071 ( .A1(n8178), .A2(n8179), .ZN(n8121) );
  NAND2_X1 U8072 ( .A1(b_0_), .A2(n8175), .ZN(n8179) );
  NAND2_X1 U8073 ( .A1(n8180), .A2(n8181), .ZN(n8175) );
  NAND2_X1 U8074 ( .A1(n8176), .A2(n8177), .ZN(n8178) );
  NAND2_X1 U8075 ( .A1(n8067), .A2(n8182), .ZN(n8119) );
  NAND2_X1 U8076 ( .A1(n8068), .A2(n8065), .ZN(n8182) );
  NAND2_X1 U8077 ( .A1(n7861), .A2(n8183), .ZN(n8065) );
  NAND2_X1 U8078 ( .A1(n7862), .A2(n7859), .ZN(n8183) );
  NAND2_X1 U8079 ( .A1(n7715), .A2(n8184), .ZN(n7859) );
  NAND2_X1 U8080 ( .A1(n7716), .A2(n7713), .ZN(n8184) );
  NAND2_X1 U8081 ( .A1(n7569), .A2(n8185), .ZN(n7713) );
  NAND2_X1 U8082 ( .A1(n7570), .A2(n7567), .ZN(n8185) );
  NAND2_X1 U8083 ( .A1(n7514), .A2(n8186), .ZN(n7567) );
  NAND2_X1 U8084 ( .A1(n7515), .A2(n7512), .ZN(n8186) );
  NAND2_X1 U8085 ( .A1(n7509), .A2(n8187), .ZN(n7512) );
  NAND2_X1 U8086 ( .A1(n7510), .A2(n7507), .ZN(n8187) );
  NAND2_X1 U8087 ( .A1(n7504), .A2(n8188), .ZN(n7507) );
  NAND2_X1 U8088 ( .A1(n7505), .A2(n7502), .ZN(n8188) );
  NAND2_X1 U8089 ( .A1(n7499), .A2(n8189), .ZN(n7502) );
  NAND2_X1 U8090 ( .A1(n7500), .A2(n7497), .ZN(n8189) );
  NAND2_X1 U8091 ( .A1(n8171), .A2(n8190), .ZN(n7497) );
  NAND2_X1 U8092 ( .A1(n8169), .A2(n8172), .ZN(n8190) );
  NAND2_X1 U8093 ( .A1(n8191), .A2(n8192), .ZN(n8172) );
  XNOR2_X1 U8094 ( .A(n8193), .B(n8194), .ZN(n8191) );
  NAND2_X1 U8095 ( .A1(n8166), .A2(n8195), .ZN(n8169) );
  NAND2_X1 U8096 ( .A1(n8164), .A2(n8167), .ZN(n8195) );
  NAND2_X1 U8097 ( .A1(n8196), .A2(n8197), .ZN(n8167) );
  NAND2_X1 U8098 ( .A1(n8198), .A2(n8192), .ZN(n8197) );
  NAND2_X1 U8099 ( .A1(n8199), .A2(n8200), .ZN(n8196) );
  NAND2_X1 U8100 ( .A1(n8161), .A2(n8201), .ZN(n8164) );
  NAND2_X1 U8101 ( .A1(n8159), .A2(n8162), .ZN(n8201) );
  NAND2_X1 U8102 ( .A1(n8202), .A2(n8203), .ZN(n8162) );
  XNOR2_X1 U8103 ( .A(n8200), .B(n8199), .ZN(n8202) );
  NAND2_X1 U8104 ( .A1(n8156), .A2(n8204), .ZN(n8159) );
  NAND2_X1 U8105 ( .A1(n8154), .A2(n8157), .ZN(n8204) );
  NAND2_X1 U8106 ( .A1(n8205), .A2(n8206), .ZN(n8157) );
  NAND2_X1 U8107 ( .A1(n8207), .A2(n8203), .ZN(n8206) );
  NAND2_X1 U8108 ( .A1(n8208), .A2(n8209), .ZN(n8205) );
  NAND2_X1 U8109 ( .A1(n8151), .A2(n8210), .ZN(n8154) );
  NAND2_X1 U8110 ( .A1(n8152), .A2(n8149), .ZN(n8210) );
  NAND2_X1 U8111 ( .A1(n8146), .A2(n8211), .ZN(n8149) );
  NAND2_X1 U8112 ( .A1(n8147), .A2(n8144), .ZN(n8211) );
  NAND2_X1 U8113 ( .A1(n8141), .A2(n8212), .ZN(n8144) );
  NAND2_X1 U8114 ( .A1(n8139), .A2(n8142), .ZN(n8212) );
  NAND2_X1 U8115 ( .A1(n8213), .A2(n8214), .ZN(n8142) );
  NAND2_X1 U8116 ( .A1(n8215), .A2(n8216), .ZN(n8214) );
  XNOR2_X1 U8117 ( .A(n8217), .B(n8218), .ZN(n8213) );
  NAND2_X1 U8118 ( .A1(n8136), .A2(n8219), .ZN(n8139) );
  NAND2_X1 U8119 ( .A1(n8137), .A2(n8134), .ZN(n8219) );
  NAND2_X1 U8120 ( .A1(n8131), .A2(n8220), .ZN(n8134) );
  NAND2_X1 U8121 ( .A1(n8129), .A2(n8132), .ZN(n8220) );
  NAND2_X1 U8122 ( .A1(n8221), .A2(n8222), .ZN(n8132) );
  NAND2_X1 U8123 ( .A1(n8223), .A2(n8224), .ZN(n8222) );
  XNOR2_X1 U8124 ( .A(n8225), .B(n8226), .ZN(n8221) );
  NAND2_X1 U8125 ( .A1(n8126), .A2(n8227), .ZN(n8129) );
  NAND2_X1 U8126 ( .A1(n8124), .A2(n8127), .ZN(n8227) );
  NAND2_X1 U8127 ( .A1(n8228), .A2(n8229), .ZN(n8127) );
  NAND2_X1 U8128 ( .A1(n8230), .A2(n8231), .ZN(n8229) );
  XNOR2_X1 U8129 ( .A(n8223), .B(n8224), .ZN(n8228) );
  NAND2_X1 U8130 ( .A1(n8117), .A2(n8232), .ZN(n8124) );
  NAND2_X1 U8131 ( .A1(n8114), .A2(n8116), .ZN(n8232) );
  NAND2_X1 U8132 ( .A1(n8233), .A2(n8234), .ZN(n8116) );
  XNOR2_X1 U8133 ( .A(n8231), .B(n8230), .ZN(n8233) );
  NAND2_X1 U8134 ( .A1(n8112), .A2(n8235), .ZN(n8114) );
  NAND2_X1 U8135 ( .A1(n8109), .A2(n8111), .ZN(n8235) );
  NAND2_X1 U8136 ( .A1(n8236), .A2(n8237), .ZN(n8111) );
  NAND2_X1 U8137 ( .A1(n8238), .A2(n8234), .ZN(n8237) );
  NAND2_X1 U8138 ( .A1(n8239), .A2(n8240), .ZN(n8236) );
  NAND2_X1 U8139 ( .A1(n8106), .A2(n8241), .ZN(n8109) );
  NAND2_X1 U8140 ( .A1(n8104), .A2(n8107), .ZN(n8241) );
  NAND2_X1 U8141 ( .A1(n8242), .A2(n8243), .ZN(n8107) );
  NAND2_X1 U8142 ( .A1(n8244), .A2(n8245), .ZN(n8243) );
  XNOR2_X1 U8143 ( .A(n8240), .B(n8239), .ZN(n8242) );
  NAND2_X1 U8144 ( .A1(n8101), .A2(n8246), .ZN(n8104) );
  NAND2_X1 U8145 ( .A1(n8099), .A2(n8102), .ZN(n8246) );
  NAND2_X1 U8146 ( .A1(n8247), .A2(n8248), .ZN(n8102) );
  NAND2_X1 U8147 ( .A1(n8249), .A2(n8250), .ZN(n8248) );
  XNOR2_X1 U8148 ( .A(n8245), .B(n8244), .ZN(n8247) );
  NAND2_X1 U8149 ( .A1(n8097), .A2(n8251), .ZN(n8099) );
  NAND2_X1 U8150 ( .A1(n8094), .A2(n8096), .ZN(n8251) );
  NAND2_X1 U8151 ( .A1(n8252), .A2(n8253), .ZN(n8096) );
  XOR2_X1 U8152 ( .A(n8250), .B(n8254), .Z(n8252) );
  NAND2_X1 U8153 ( .A1(n8092), .A2(n8255), .ZN(n8094) );
  NAND2_X1 U8154 ( .A1(n8089), .A2(n8091), .ZN(n8255) );
  NAND2_X1 U8155 ( .A1(n8256), .A2(n8257), .ZN(n8091) );
  NAND2_X1 U8156 ( .A1(n8258), .A2(n8253), .ZN(n8257) );
  NAND2_X1 U8157 ( .A1(n8259), .A2(n8260), .ZN(n8256) );
  NAND2_X1 U8158 ( .A1(n8087), .A2(n8261), .ZN(n8089) );
  NAND2_X1 U8159 ( .A1(n8085), .A2(n8086), .ZN(n8261) );
  NAND2_X1 U8160 ( .A1(n8262), .A2(n8263), .ZN(n8086) );
  XNOR2_X1 U8161 ( .A(n8259), .B(n8260), .ZN(n8262) );
  NAND2_X1 U8162 ( .A1(n8264), .A2(n8265), .ZN(n8085) );
  OR2_X1 U8163 ( .A1(n8079), .A2(n8081), .ZN(n8265) );
  AND2_X1 U8164 ( .A1(n8266), .A2(n8267), .ZN(n8081) );
  NOR2_X1 U8165 ( .A1(n8268), .A2(n8076), .ZN(n8079) );
  NOR2_X1 U8166 ( .A1(n8269), .A2(n8270), .ZN(n8076) );
  NOR2_X1 U8167 ( .A1(n8077), .A2(n8074), .ZN(n8268) );
  AND2_X1 U8168 ( .A1(n8071), .A2(n8271), .ZN(n8074) );
  NAND2_X1 U8169 ( .A1(n8061), .A2(n8072), .ZN(n8271) );
  NAND2_X1 U8170 ( .A1(n8272), .A2(n8273), .ZN(n8072) );
  NAND2_X1 U8171 ( .A1(n8274), .A2(n8275), .ZN(n8273) );
  XNOR2_X1 U8172 ( .A(n8276), .B(n8277), .ZN(n8272) );
  AND3_X1 U8173 ( .A1(n8063), .A2(n8059), .A3(n8058), .ZN(n8061) );
  XNOR2_X1 U8174 ( .A(n8278), .B(n8279), .ZN(n8058) );
  XOR2_X1 U8175 ( .A(n8280), .B(n8281), .Z(n8279) );
  NAND2_X1 U8176 ( .A1(a_0_), .A2(b_30_), .ZN(n8281) );
  NAND2_X1 U8177 ( .A1(n8282), .A2(n8283), .ZN(n8059) );
  NAND3_X1 U8178 ( .A1(b_31_), .A2(n8284), .A3(a_0_), .ZN(n8283) );
  NAND2_X1 U8179 ( .A1(n7972), .A2(n7970), .ZN(n8284) );
  OR2_X1 U8180 ( .A1(n7970), .A2(n7972), .ZN(n8282) );
  AND2_X1 U8181 ( .A1(n8285), .A2(n8286), .ZN(n7972) );
  NAND3_X1 U8182 ( .A1(a_1_), .A2(n8287), .A3(b_31_), .ZN(n8286) );
  OR2_X1 U8183 ( .A1(n7955), .A2(n7954), .ZN(n8287) );
  NAND2_X1 U8184 ( .A1(n7954), .A2(n7955), .ZN(n8285) );
  NAND2_X1 U8185 ( .A1(n8288), .A2(n8289), .ZN(n7955) );
  NAND3_X1 U8186 ( .A1(b_31_), .A2(n8290), .A3(a_2_), .ZN(n8289) );
  NAND2_X1 U8187 ( .A1(n7943), .A2(n7941), .ZN(n8290) );
  OR2_X1 U8188 ( .A1(n7941), .A2(n7943), .ZN(n8288) );
  AND2_X1 U8189 ( .A1(n8291), .A2(n8292), .ZN(n7943) );
  NAND3_X1 U8190 ( .A1(b_31_), .A2(n8293), .A3(a_3_), .ZN(n8292) );
  OR2_X1 U8191 ( .A1(n7935), .A2(n7934), .ZN(n8293) );
  NAND2_X1 U8192 ( .A1(n7934), .A2(n7935), .ZN(n8291) );
  NAND2_X1 U8193 ( .A1(n8294), .A2(n8295), .ZN(n7935) );
  NAND3_X1 U8194 ( .A1(b_31_), .A2(n8296), .A3(a_4_), .ZN(n8295) );
  OR2_X1 U8195 ( .A1(n7914), .A2(n7913), .ZN(n8296) );
  NAND2_X1 U8196 ( .A1(n7913), .A2(n7914), .ZN(n8294) );
  NAND2_X1 U8197 ( .A1(n8297), .A2(n8298), .ZN(n7914) );
  NAND3_X1 U8198 ( .A1(b_31_), .A2(n8299), .A3(a_5_), .ZN(n8298) );
  OR2_X1 U8199 ( .A1(n7906), .A2(n7905), .ZN(n8299) );
  NAND2_X1 U8200 ( .A1(n7905), .A2(n7906), .ZN(n8297) );
  NAND2_X1 U8201 ( .A1(n8300), .A2(n8301), .ZN(n7906) );
  NAND3_X1 U8202 ( .A1(b_31_), .A2(n8302), .A3(a_6_), .ZN(n8301) );
  OR2_X1 U8203 ( .A1(n7885), .A2(n7884), .ZN(n8302) );
  NAND2_X1 U8204 ( .A1(n7884), .A2(n7885), .ZN(n8300) );
  NAND2_X1 U8205 ( .A1(n8303), .A2(n8304), .ZN(n7885) );
  NAND3_X1 U8206 ( .A1(b_31_), .A2(n8305), .A3(a_7_), .ZN(n8304) );
  OR2_X1 U8207 ( .A1(n7878), .A2(n7876), .ZN(n8305) );
  NAND2_X1 U8208 ( .A1(n7876), .A2(n7878), .ZN(n8303) );
  NAND2_X1 U8209 ( .A1(n8306), .A2(n8307), .ZN(n7878) );
  NAND3_X1 U8210 ( .A1(b_31_), .A2(n8308), .A3(a_8_), .ZN(n8307) );
  NAND2_X1 U8211 ( .A1(n7851), .A2(n7849), .ZN(n8308) );
  OR2_X1 U8212 ( .A1(n7849), .A2(n7851), .ZN(n8306) );
  AND2_X1 U8213 ( .A1(n8309), .A2(n8310), .ZN(n7851) );
  NAND3_X1 U8214 ( .A1(b_31_), .A2(n8311), .A3(a_9_), .ZN(n8310) );
  NAND2_X1 U8215 ( .A1(n7844), .A2(n7842), .ZN(n8311) );
  OR2_X1 U8216 ( .A1(n7842), .A2(n7844), .ZN(n8309) );
  AND2_X1 U8217 ( .A1(n8312), .A2(n8313), .ZN(n7844) );
  NAND3_X1 U8218 ( .A1(b_31_), .A2(n8314), .A3(a_10_), .ZN(n8313) );
  NAND2_X1 U8219 ( .A1(n7824), .A2(n7822), .ZN(n8314) );
  OR2_X1 U8220 ( .A1(n7822), .A2(n7824), .ZN(n8312) );
  AND2_X1 U8221 ( .A1(n8315), .A2(n8316), .ZN(n7824) );
  NAND3_X1 U8222 ( .A1(b_31_), .A2(n8317), .A3(a_11_), .ZN(n8316) );
  OR2_X1 U8223 ( .A1(n7817), .A2(n7815), .ZN(n8317) );
  NAND2_X1 U8224 ( .A1(n7815), .A2(n7817), .ZN(n8315) );
  NAND2_X1 U8225 ( .A1(n8318), .A2(n8319), .ZN(n7817) );
  NAND3_X1 U8226 ( .A1(b_31_), .A2(n8320), .A3(a_12_), .ZN(n8319) );
  NAND2_X1 U8227 ( .A1(n7795), .A2(n7793), .ZN(n8320) );
  OR2_X1 U8228 ( .A1(n7793), .A2(n7795), .ZN(n8318) );
  AND2_X1 U8229 ( .A1(n8321), .A2(n8322), .ZN(n7795) );
  NAND3_X1 U8230 ( .A1(b_31_), .A2(n8323), .A3(a_13_), .ZN(n8322) );
  OR2_X1 U8231 ( .A1(n7787), .A2(n7786), .ZN(n8323) );
  NAND2_X1 U8232 ( .A1(n7786), .A2(n7787), .ZN(n8321) );
  NAND2_X1 U8233 ( .A1(n8324), .A2(n8325), .ZN(n7787) );
  NAND3_X1 U8234 ( .A1(b_31_), .A2(n8326), .A3(a_14_), .ZN(n8325) );
  NAND2_X1 U8235 ( .A1(n7767), .A2(n7765), .ZN(n8326) );
  OR2_X1 U8236 ( .A1(n7765), .A2(n7767), .ZN(n8324) );
  AND2_X1 U8237 ( .A1(n8327), .A2(n8328), .ZN(n7767) );
  NAND3_X1 U8238 ( .A1(b_31_), .A2(n8329), .A3(a_15_), .ZN(n8328) );
  OR2_X1 U8239 ( .A1(n7760), .A2(n7758), .ZN(n8329) );
  NAND2_X1 U8240 ( .A1(n7758), .A2(n7760), .ZN(n8327) );
  NAND2_X1 U8241 ( .A1(n8330), .A2(n8331), .ZN(n7760) );
  NAND3_X1 U8242 ( .A1(b_31_), .A2(n8332), .A3(a_16_), .ZN(n8331) );
  NAND2_X1 U8243 ( .A1(n7738), .A2(n7736), .ZN(n8332) );
  OR2_X1 U8244 ( .A1(n7736), .A2(n7738), .ZN(n8330) );
  AND2_X1 U8245 ( .A1(n8333), .A2(n8334), .ZN(n7738) );
  NAND3_X1 U8246 ( .A1(b_31_), .A2(n8335), .A3(a_17_), .ZN(n8334) );
  OR2_X1 U8247 ( .A1(n7730), .A2(n7729), .ZN(n8335) );
  NAND2_X1 U8248 ( .A1(n7729), .A2(n7730), .ZN(n8333) );
  NAND2_X1 U8249 ( .A1(n8336), .A2(n8337), .ZN(n7730) );
  NAND3_X1 U8250 ( .A1(b_31_), .A2(n8338), .A3(a_18_), .ZN(n8337) );
  NAND2_X1 U8251 ( .A1(n7705), .A2(n7703), .ZN(n8338) );
  OR2_X1 U8252 ( .A1(n7703), .A2(n7705), .ZN(n8336) );
  AND2_X1 U8253 ( .A1(n8339), .A2(n8340), .ZN(n7705) );
  NAND3_X1 U8254 ( .A1(b_31_), .A2(n8341), .A3(a_19_), .ZN(n8340) );
  OR2_X1 U8255 ( .A1(n7698), .A2(n7696), .ZN(n8341) );
  NAND2_X1 U8256 ( .A1(n7696), .A2(n7698), .ZN(n8339) );
  NAND2_X1 U8257 ( .A1(n8342), .A2(n8343), .ZN(n7698) );
  NAND3_X1 U8258 ( .A1(b_31_), .A2(n8344), .A3(a_20_), .ZN(n8343) );
  NAND2_X1 U8259 ( .A1(n7678), .A2(n7676), .ZN(n8344) );
  OR2_X1 U8260 ( .A1(n7676), .A2(n7678), .ZN(n8342) );
  AND2_X1 U8261 ( .A1(n8345), .A2(n8346), .ZN(n7678) );
  NAND3_X1 U8262 ( .A1(b_31_), .A2(n8347), .A3(a_21_), .ZN(n8346) );
  NAND2_X1 U8263 ( .A1(n7671), .A2(n7669), .ZN(n8347) );
  OR2_X1 U8264 ( .A1(n7669), .A2(n7671), .ZN(n8345) );
  AND2_X1 U8265 ( .A1(n8348), .A2(n8349), .ZN(n7671) );
  NAND3_X1 U8266 ( .A1(b_31_), .A2(n8350), .A3(a_22_), .ZN(n8349) );
  NAND2_X1 U8267 ( .A1(n7648), .A2(n7646), .ZN(n8350) );
  OR2_X1 U8268 ( .A1(n7646), .A2(n7648), .ZN(n8348) );
  AND2_X1 U8269 ( .A1(n7641), .A2(n8351), .ZN(n7648) );
  NAND2_X1 U8270 ( .A1(n7640), .A2(n7642), .ZN(n8351) );
  NAND2_X1 U8271 ( .A1(n8352), .A2(n8353), .ZN(n7642) );
  NAND2_X1 U8272 ( .A1(a_23_), .A2(b_31_), .ZN(n8353) );
  INV_X1 U8273 ( .A(n8354), .ZN(n8352) );
  XOR2_X1 U8274 ( .A(n8355), .B(n8356), .Z(n7640) );
  XOR2_X1 U8275 ( .A(n8357), .B(n8358), .Z(n8355) );
  NOR2_X1 U8276 ( .A1(n8359), .A2(n8041), .ZN(n8358) );
  NAND2_X1 U8277 ( .A1(a_23_), .A2(n8354), .ZN(n7641) );
  NAND2_X1 U8278 ( .A1(n8360), .A2(n8361), .ZN(n8354) );
  NAND3_X1 U8279 ( .A1(b_31_), .A2(n8362), .A3(a_24_), .ZN(n8361) );
  OR2_X1 U8280 ( .A1(n7622), .A2(n7619), .ZN(n8362) );
  NAND2_X1 U8281 ( .A1(n7619), .A2(n7622), .ZN(n8360) );
  NAND2_X1 U8282 ( .A1(n7614), .A2(n8363), .ZN(n7622) );
  NAND2_X1 U8283 ( .A1(n7613), .A2(n7615), .ZN(n8363) );
  NAND2_X1 U8284 ( .A1(n8364), .A2(n8365), .ZN(n7615) );
  NAND2_X1 U8285 ( .A1(a_25_), .A2(b_31_), .ZN(n8365) );
  INV_X1 U8286 ( .A(n8366), .ZN(n8364) );
  XNOR2_X1 U8287 ( .A(n8367), .B(n8368), .ZN(n7613) );
  NAND2_X1 U8288 ( .A1(n8369), .A2(n8370), .ZN(n8367) );
  NAND2_X1 U8289 ( .A1(a_25_), .A2(n8366), .ZN(n7614) );
  NAND2_X1 U8290 ( .A1(n8371), .A2(n8372), .ZN(n8366) );
  NAND3_X1 U8291 ( .A1(b_31_), .A2(n8373), .A3(a_26_), .ZN(n8372) );
  OR2_X1 U8292 ( .A1(n7593), .A2(n7592), .ZN(n8373) );
  NAND2_X1 U8293 ( .A1(n7592), .A2(n7593), .ZN(n8371) );
  NAND2_X1 U8294 ( .A1(n7586), .A2(n8374), .ZN(n7593) );
  NAND2_X1 U8295 ( .A1(n7585), .A2(n7587), .ZN(n8374) );
  NAND2_X1 U8296 ( .A1(n8375), .A2(n8376), .ZN(n7587) );
  NAND2_X1 U8297 ( .A1(a_27_), .A2(b_31_), .ZN(n8376) );
  INV_X1 U8298 ( .A(n8377), .ZN(n8375) );
  XNOR2_X1 U8299 ( .A(n8378), .B(n8379), .ZN(n7585) );
  XOR2_X1 U8300 ( .A(n8380), .B(n8381), .Z(n8378) );
  NAND2_X1 U8301 ( .A1(a_28_), .A2(b_30_), .ZN(n8380) );
  NAND2_X1 U8302 ( .A1(a_27_), .A2(n8377), .ZN(n7586) );
  NAND2_X1 U8303 ( .A1(n8382), .A2(n8383), .ZN(n8377) );
  NAND3_X1 U8304 ( .A1(b_31_), .A2(n8384), .A3(a_28_), .ZN(n8383) );
  NAND2_X1 U8305 ( .A1(n7558), .A2(n7556), .ZN(n8384) );
  OR2_X1 U8306 ( .A1(n7556), .A2(n7558), .ZN(n8382) );
  AND2_X1 U8307 ( .A1(n8385), .A2(n8386), .ZN(n7558) );
  NAND3_X1 U8308 ( .A1(b_31_), .A2(n8387), .A3(a_29_), .ZN(n8386) );
  OR2_X1 U8309 ( .A1(n7551), .A2(n7552), .ZN(n8387) );
  NAND2_X1 U8310 ( .A1(n7552), .A2(n7551), .ZN(n8385) );
  NAND2_X1 U8311 ( .A1(n8388), .A2(n8389), .ZN(n7551) );
  NAND2_X1 U8312 ( .A1(b_29_), .A2(n8390), .ZN(n8389) );
  NAND2_X1 U8313 ( .A1(n7527), .A2(n8391), .ZN(n8390) );
  NAND2_X1 U8314 ( .A1(a_31_), .A2(n8359), .ZN(n8391) );
  NAND2_X1 U8315 ( .A1(b_30_), .A2(n8392), .ZN(n8388) );
  NAND2_X1 U8316 ( .A1(n7531), .A2(n8393), .ZN(n8392) );
  NAND2_X1 U8317 ( .A1(a_30_), .A2(n7547), .ZN(n8393) );
  AND3_X1 U8318 ( .A1(b_30_), .A2(b_31_), .A3(n7494), .ZN(n7552) );
  XNOR2_X1 U8319 ( .A(n8394), .B(n8395), .ZN(n7556) );
  XOR2_X1 U8320 ( .A(n8396), .B(n8397), .Z(n8394) );
  XNOR2_X1 U8321 ( .A(n8398), .B(n8399), .ZN(n7592) );
  NAND2_X1 U8322 ( .A1(n8400), .A2(n8401), .ZN(n8398) );
  XOR2_X1 U8323 ( .A(n8402), .B(n8403), .Z(n7619) );
  XOR2_X1 U8324 ( .A(n8404), .B(n8405), .Z(n8402) );
  XOR2_X1 U8325 ( .A(n8406), .B(n8407), .Z(n7646) );
  XNOR2_X1 U8326 ( .A(n8408), .B(n8409), .ZN(n8407) );
  XNOR2_X1 U8327 ( .A(n8410), .B(n8411), .ZN(n7669) );
  XOR2_X1 U8328 ( .A(n8412), .B(n8413), .Z(n8410) );
  NOR2_X1 U8329 ( .A1(n8359), .A2(n7650), .ZN(n8413) );
  XNOR2_X1 U8330 ( .A(n8414), .B(n8415), .ZN(n7676) );
  XOR2_X1 U8331 ( .A(n8416), .B(n8417), .Z(n8414) );
  XNOR2_X1 U8332 ( .A(n8418), .B(n8419), .ZN(n7696) );
  XOR2_X1 U8333 ( .A(n8420), .B(n8421), .Z(n8419) );
  NAND2_X1 U8334 ( .A1(a_20_), .A2(b_30_), .ZN(n8421) );
  XOR2_X1 U8335 ( .A(n8422), .B(n8423), .Z(n7703) );
  XNOR2_X1 U8336 ( .A(n8424), .B(n8425), .ZN(n8423) );
  XNOR2_X1 U8337 ( .A(n8426), .B(n8427), .ZN(n7729) );
  XNOR2_X1 U8338 ( .A(n8428), .B(n8429), .ZN(n8426) );
  NOR2_X1 U8339 ( .A1(n8359), .A2(n8047), .ZN(n8429) );
  XOR2_X1 U8340 ( .A(n8430), .B(n8431), .Z(n7736) );
  XNOR2_X1 U8341 ( .A(n8432), .B(n8433), .ZN(n8431) );
  XNOR2_X1 U8342 ( .A(n8434), .B(n8435), .ZN(n7758) );
  XNOR2_X1 U8343 ( .A(n8436), .B(n8437), .ZN(n8434) );
  NOR2_X1 U8344 ( .A1(n8359), .A2(n8438), .ZN(n8437) );
  XOR2_X1 U8345 ( .A(n8439), .B(n8440), .Z(n7765) );
  XNOR2_X1 U8346 ( .A(n8441), .B(n8442), .ZN(n8440) );
  XNOR2_X1 U8347 ( .A(n8443), .B(n8444), .ZN(n7786) );
  XNOR2_X1 U8348 ( .A(n8445), .B(n8446), .ZN(n8443) );
  NOR2_X1 U8349 ( .A1(n8359), .A2(n8049), .ZN(n8446) );
  XNOR2_X1 U8350 ( .A(n8447), .B(n8448), .ZN(n7793) );
  XOR2_X1 U8351 ( .A(n8449), .B(n8450), .Z(n8447) );
  XNOR2_X1 U8352 ( .A(n8451), .B(n8452), .ZN(n7815) );
  XOR2_X1 U8353 ( .A(n8453), .B(n8454), .Z(n8452) );
  NAND2_X1 U8354 ( .A1(a_12_), .A2(b_30_), .ZN(n8454) );
  XOR2_X1 U8355 ( .A(n8455), .B(n8456), .Z(n7822) );
  XNOR2_X1 U8356 ( .A(n8457), .B(n8458), .ZN(n8456) );
  XNOR2_X1 U8357 ( .A(n8459), .B(n8460), .ZN(n7842) );
  XOR2_X1 U8358 ( .A(n8461), .B(n8462), .Z(n8459) );
  NOR2_X1 U8359 ( .A1(n8359), .A2(n8051), .ZN(n8462) );
  XNOR2_X1 U8360 ( .A(n8463), .B(n8464), .ZN(n7849) );
  XOR2_X1 U8361 ( .A(n8465), .B(n8466), .Z(n8463) );
  XNOR2_X1 U8362 ( .A(n8467), .B(n8468), .ZN(n7876) );
  XOR2_X1 U8363 ( .A(n8469), .B(n8470), .Z(n8468) );
  NAND2_X1 U8364 ( .A1(a_8_), .A2(b_30_), .ZN(n8470) );
  XNOR2_X1 U8365 ( .A(n8471), .B(n8472), .ZN(n7884) );
  XNOR2_X1 U8366 ( .A(n8473), .B(n8474), .ZN(n8472) );
  XNOR2_X1 U8367 ( .A(n8475), .B(n8476), .ZN(n7905) );
  XNOR2_X1 U8368 ( .A(n8477), .B(n8478), .ZN(n8475) );
  NOR2_X1 U8369 ( .A1(n8359), .A2(n7887), .ZN(n8478) );
  XNOR2_X1 U8370 ( .A(n8479), .B(n8480), .ZN(n7913) );
  XNOR2_X1 U8371 ( .A(n8481), .B(n8482), .ZN(n8479) );
  XNOR2_X1 U8372 ( .A(n8483), .B(n8484), .ZN(n7934) );
  XOR2_X1 U8373 ( .A(n8485), .B(n8486), .Z(n8484) );
  NAND2_X1 U8374 ( .A1(a_4_), .A2(b_30_), .ZN(n8486) );
  XOR2_X1 U8375 ( .A(n8487), .B(n8488), .Z(n7941) );
  XNOR2_X1 U8376 ( .A(n8489), .B(n8490), .ZN(n8488) );
  XNOR2_X1 U8377 ( .A(n8491), .B(n8492), .ZN(n7954) );
  XNOR2_X1 U8378 ( .A(n8493), .B(n8494), .ZN(n8491) );
  NOR2_X1 U8379 ( .A1(n8359), .A2(n8056), .ZN(n8494) );
  XNOR2_X1 U8380 ( .A(n8495), .B(n8496), .ZN(n7970) );
  XOR2_X1 U8381 ( .A(n8497), .B(n8498), .Z(n8495) );
  NOR2_X1 U8382 ( .A1(n7957), .A2(n8359), .ZN(n8498) );
  XOR2_X1 U8383 ( .A(n8275), .B(n8274), .Z(n8063) );
  NAND4_X1 U8384 ( .A1(n8274), .A2(n8499), .A3(n8275), .A4(n8270), .ZN(n8071)
         );
  NAND2_X1 U8385 ( .A1(n8500), .A2(n8501), .ZN(n8275) );
  NAND3_X1 U8386 ( .A1(b_30_), .A2(n8502), .A3(a_0_), .ZN(n8501) );
  OR2_X1 U8387 ( .A1(n8280), .A2(n8278), .ZN(n8502) );
  NAND2_X1 U8388 ( .A1(n8278), .A2(n8280), .ZN(n8500) );
  NAND2_X1 U8389 ( .A1(n8503), .A2(n8504), .ZN(n8280) );
  NAND3_X1 U8390 ( .A1(a_1_), .A2(n8505), .A3(b_30_), .ZN(n8504) );
  OR2_X1 U8391 ( .A1(n8496), .A2(n8497), .ZN(n8505) );
  NAND2_X1 U8392 ( .A1(n8496), .A2(n8497), .ZN(n8503) );
  NAND2_X1 U8393 ( .A1(n8506), .A2(n8507), .ZN(n8497) );
  NAND3_X1 U8394 ( .A1(b_30_), .A2(n8508), .A3(a_2_), .ZN(n8507) );
  NAND2_X1 U8395 ( .A1(n8493), .A2(n8492), .ZN(n8508) );
  OR2_X1 U8396 ( .A1(n8492), .A2(n8493), .ZN(n8506) );
  AND2_X1 U8397 ( .A1(n8509), .A2(n8510), .ZN(n8493) );
  NAND2_X1 U8398 ( .A1(n8490), .A2(n8511), .ZN(n8510) );
  OR2_X1 U8399 ( .A1(n8487), .A2(n8489), .ZN(n8511) );
  NOR2_X1 U8400 ( .A1(n7937), .A2(n8359), .ZN(n8490) );
  NAND2_X1 U8401 ( .A1(n8487), .A2(n8489), .ZN(n8509) );
  NAND2_X1 U8402 ( .A1(n8512), .A2(n8513), .ZN(n8489) );
  NAND3_X1 U8403 ( .A1(b_30_), .A2(n8514), .A3(a_4_), .ZN(n8513) );
  OR2_X1 U8404 ( .A1(n8485), .A2(n8483), .ZN(n8514) );
  NAND2_X1 U8405 ( .A1(n8483), .A2(n8485), .ZN(n8512) );
  NAND2_X1 U8406 ( .A1(n8515), .A2(n8516), .ZN(n8485) );
  NAND2_X1 U8407 ( .A1(n8482), .A2(n8517), .ZN(n8516) );
  NAND2_X1 U8408 ( .A1(n8481), .A2(n8480), .ZN(n8517) );
  NOR2_X1 U8409 ( .A1(n7908), .A2(n8359), .ZN(n8482) );
  OR2_X1 U8410 ( .A1(n8480), .A2(n8481), .ZN(n8515) );
  AND2_X1 U8411 ( .A1(n8518), .A2(n8519), .ZN(n8481) );
  NAND3_X1 U8412 ( .A1(b_30_), .A2(n8520), .A3(a_6_), .ZN(n8519) );
  NAND2_X1 U8413 ( .A1(n8477), .A2(n8476), .ZN(n8520) );
  OR2_X1 U8414 ( .A1(n8476), .A2(n8477), .ZN(n8518) );
  AND2_X1 U8415 ( .A1(n8521), .A2(n8522), .ZN(n8477) );
  NAND2_X1 U8416 ( .A1(n8474), .A2(n8523), .ZN(n8522) );
  OR2_X1 U8417 ( .A1(n8473), .A2(n8471), .ZN(n8523) );
  NOR2_X1 U8418 ( .A1(n7872), .A2(n8359), .ZN(n8474) );
  NAND2_X1 U8419 ( .A1(n8471), .A2(n8473), .ZN(n8521) );
  NAND2_X1 U8420 ( .A1(n8524), .A2(n8525), .ZN(n8473) );
  NAND3_X1 U8421 ( .A1(b_30_), .A2(n8526), .A3(a_8_), .ZN(n8525) );
  OR2_X1 U8422 ( .A1(n8469), .A2(n8467), .ZN(n8526) );
  NAND2_X1 U8423 ( .A1(n8467), .A2(n8469), .ZN(n8524) );
  NAND2_X1 U8424 ( .A1(n8527), .A2(n8528), .ZN(n8469) );
  NAND2_X1 U8425 ( .A1(n8466), .A2(n8529), .ZN(n8528) );
  OR2_X1 U8426 ( .A1(n8464), .A2(n8465), .ZN(n8529) );
  NOR2_X1 U8427 ( .A1(n8052), .A2(n8359), .ZN(n8466) );
  NAND2_X1 U8428 ( .A1(n8464), .A2(n8465), .ZN(n8527) );
  NAND2_X1 U8429 ( .A1(n8530), .A2(n8531), .ZN(n8465) );
  NAND3_X1 U8430 ( .A1(b_30_), .A2(n8532), .A3(a_10_), .ZN(n8531) );
  OR2_X1 U8431 ( .A1(n8460), .A2(n8461), .ZN(n8532) );
  NAND2_X1 U8432 ( .A1(n8460), .A2(n8461), .ZN(n8530) );
  NAND2_X1 U8433 ( .A1(n8533), .A2(n8534), .ZN(n8461) );
  NAND2_X1 U8434 ( .A1(n8458), .A2(n8535), .ZN(n8534) );
  OR2_X1 U8435 ( .A1(n8455), .A2(n8457), .ZN(n8535) );
  NOR2_X1 U8436 ( .A1(n7811), .A2(n8359), .ZN(n8458) );
  NAND2_X1 U8437 ( .A1(n8455), .A2(n8457), .ZN(n8533) );
  NAND2_X1 U8438 ( .A1(n8536), .A2(n8537), .ZN(n8457) );
  NAND3_X1 U8439 ( .A1(b_30_), .A2(n8538), .A3(a_12_), .ZN(n8537) );
  OR2_X1 U8440 ( .A1(n8453), .A2(n8451), .ZN(n8538) );
  NAND2_X1 U8441 ( .A1(n8451), .A2(n8453), .ZN(n8536) );
  NAND2_X1 U8442 ( .A1(n8539), .A2(n8540), .ZN(n8453) );
  NAND2_X1 U8443 ( .A1(n8450), .A2(n8541), .ZN(n8540) );
  OR2_X1 U8444 ( .A1(n8448), .A2(n8449), .ZN(n8541) );
  NOR2_X1 U8445 ( .A1(n7789), .A2(n8359), .ZN(n8450) );
  NAND2_X1 U8446 ( .A1(n8448), .A2(n8449), .ZN(n8539) );
  NAND2_X1 U8447 ( .A1(n8542), .A2(n8543), .ZN(n8449) );
  NAND3_X1 U8448 ( .A1(b_30_), .A2(n8544), .A3(a_14_), .ZN(n8543) );
  NAND2_X1 U8449 ( .A1(n8445), .A2(n8444), .ZN(n8544) );
  OR2_X1 U8450 ( .A1(n8444), .A2(n8445), .ZN(n8542) );
  AND2_X1 U8451 ( .A1(n8545), .A2(n8546), .ZN(n8445) );
  NAND2_X1 U8452 ( .A1(n8442), .A2(n8547), .ZN(n8546) );
  OR2_X1 U8453 ( .A1(n8439), .A2(n8441), .ZN(n8547) );
  NOR2_X1 U8454 ( .A1(n7754), .A2(n8359), .ZN(n8442) );
  NAND2_X1 U8455 ( .A1(n8439), .A2(n8441), .ZN(n8545) );
  NAND2_X1 U8456 ( .A1(n8548), .A2(n8549), .ZN(n8441) );
  NAND3_X1 U8457 ( .A1(b_30_), .A2(n8550), .A3(a_16_), .ZN(n8549) );
  NAND2_X1 U8458 ( .A1(n8436), .A2(n8435), .ZN(n8550) );
  OR2_X1 U8459 ( .A1(n8435), .A2(n8436), .ZN(n8548) );
  AND2_X1 U8460 ( .A1(n8551), .A2(n8552), .ZN(n8436) );
  NAND2_X1 U8461 ( .A1(n8433), .A2(n8553), .ZN(n8552) );
  OR2_X1 U8462 ( .A1(n8430), .A2(n8432), .ZN(n8553) );
  NOR2_X1 U8463 ( .A1(n7732), .A2(n8359), .ZN(n8433) );
  NAND2_X1 U8464 ( .A1(n8430), .A2(n8432), .ZN(n8551) );
  NAND2_X1 U8465 ( .A1(n8554), .A2(n8555), .ZN(n8432) );
  NAND3_X1 U8466 ( .A1(b_30_), .A2(n8556), .A3(a_18_), .ZN(n8555) );
  NAND2_X1 U8467 ( .A1(n8428), .A2(n8427), .ZN(n8556) );
  OR2_X1 U8468 ( .A1(n8427), .A2(n8428), .ZN(n8554) );
  AND2_X1 U8469 ( .A1(n8557), .A2(n8558), .ZN(n8428) );
  NAND2_X1 U8470 ( .A1(n8425), .A2(n8559), .ZN(n8558) );
  OR2_X1 U8471 ( .A1(n8422), .A2(n8424), .ZN(n8559) );
  NOR2_X1 U8472 ( .A1(n8045), .A2(n8359), .ZN(n8425) );
  NAND2_X1 U8473 ( .A1(n8422), .A2(n8424), .ZN(n8557) );
  NAND2_X1 U8474 ( .A1(n8560), .A2(n8561), .ZN(n8424) );
  NAND3_X1 U8475 ( .A1(b_30_), .A2(n8562), .A3(a_20_), .ZN(n8561) );
  OR2_X1 U8476 ( .A1(n8420), .A2(n8418), .ZN(n8562) );
  NAND2_X1 U8477 ( .A1(n8418), .A2(n8420), .ZN(n8560) );
  NAND2_X1 U8478 ( .A1(n8563), .A2(n8564), .ZN(n8420) );
  NAND2_X1 U8479 ( .A1(n8417), .A2(n8565), .ZN(n8564) );
  OR2_X1 U8480 ( .A1(n8415), .A2(n8416), .ZN(n8565) );
  NOR2_X1 U8481 ( .A1(n7665), .A2(n8359), .ZN(n8417) );
  NAND2_X1 U8482 ( .A1(n8415), .A2(n8416), .ZN(n8563) );
  NAND2_X1 U8483 ( .A1(n8566), .A2(n8567), .ZN(n8416) );
  NAND3_X1 U8484 ( .A1(b_30_), .A2(n8568), .A3(a_22_), .ZN(n8567) );
  OR2_X1 U8485 ( .A1(n8411), .A2(n8412), .ZN(n8568) );
  NAND2_X1 U8486 ( .A1(n8411), .A2(n8412), .ZN(n8566) );
  NAND2_X1 U8487 ( .A1(n8569), .A2(n8570), .ZN(n8412) );
  NAND2_X1 U8488 ( .A1(n8409), .A2(n8571), .ZN(n8570) );
  OR2_X1 U8489 ( .A1(n8406), .A2(n8408), .ZN(n8571) );
  NOR2_X1 U8490 ( .A1(n8042), .A2(n8359), .ZN(n8409) );
  NAND2_X1 U8491 ( .A1(n8406), .A2(n8408), .ZN(n8569) );
  NAND2_X1 U8492 ( .A1(n8572), .A2(n8573), .ZN(n8408) );
  NAND3_X1 U8493 ( .A1(b_30_), .A2(n8574), .A3(a_24_), .ZN(n8573) );
  OR2_X1 U8494 ( .A1(n8356), .A2(n8357), .ZN(n8574) );
  NAND2_X1 U8495 ( .A1(n8356), .A2(n8357), .ZN(n8572) );
  NAND2_X1 U8496 ( .A1(n8575), .A2(n8576), .ZN(n8357) );
  NAND2_X1 U8497 ( .A1(n8405), .A2(n8577), .ZN(n8576) );
  OR2_X1 U8498 ( .A1(n8403), .A2(n8404), .ZN(n8577) );
  NOR2_X1 U8499 ( .A1(n8039), .A2(n8359), .ZN(n8405) );
  NAND2_X1 U8500 ( .A1(n8403), .A2(n8404), .ZN(n8575) );
  NAND2_X1 U8501 ( .A1(n8369), .A2(n8578), .ZN(n8404) );
  NAND2_X1 U8502 ( .A1(n8368), .A2(n8370), .ZN(n8578) );
  NAND2_X1 U8503 ( .A1(n8579), .A2(n8580), .ZN(n8370) );
  NAND2_X1 U8504 ( .A1(a_26_), .A2(b_30_), .ZN(n8580) );
  INV_X1 U8505 ( .A(n8581), .ZN(n8579) );
  XNOR2_X1 U8506 ( .A(n8582), .B(n8583), .ZN(n8368) );
  NAND2_X1 U8507 ( .A1(n8584), .A2(n8585), .ZN(n8582) );
  NAND2_X1 U8508 ( .A1(a_26_), .A2(n8581), .ZN(n8369) );
  NAND2_X1 U8509 ( .A1(n8400), .A2(n8586), .ZN(n8581) );
  NAND2_X1 U8510 ( .A1(n8399), .A2(n8401), .ZN(n8586) );
  NAND2_X1 U8511 ( .A1(n8587), .A2(n8588), .ZN(n8401) );
  NAND2_X1 U8512 ( .A1(a_27_), .A2(b_30_), .ZN(n8588) );
  INV_X1 U8513 ( .A(n8589), .ZN(n8587) );
  XNOR2_X1 U8514 ( .A(n8590), .B(n8591), .ZN(n8399) );
  XOR2_X1 U8515 ( .A(n8592), .B(n8593), .Z(n8590) );
  NAND2_X1 U8516 ( .A1(a_28_), .A2(b_29_), .ZN(n8592) );
  NAND2_X1 U8517 ( .A1(a_27_), .A2(n8589), .ZN(n8400) );
  NAND2_X1 U8518 ( .A1(n8594), .A2(n8595), .ZN(n8589) );
  NAND3_X1 U8519 ( .A1(b_30_), .A2(n8596), .A3(a_28_), .ZN(n8595) );
  NAND2_X1 U8520 ( .A1(n8381), .A2(n8379), .ZN(n8596) );
  OR2_X1 U8521 ( .A1(n8379), .A2(n8381), .ZN(n8594) );
  AND2_X1 U8522 ( .A1(n8597), .A2(n8598), .ZN(n8381) );
  NAND2_X1 U8523 ( .A1(n8395), .A2(n8599), .ZN(n8598) );
  OR2_X1 U8524 ( .A1(n8396), .A2(n8397), .ZN(n8599) );
  NOR2_X1 U8525 ( .A1(n7545), .A2(n8359), .ZN(n8395) );
  NAND2_X1 U8526 ( .A1(n8397), .A2(n8396), .ZN(n8597) );
  NAND2_X1 U8527 ( .A1(n8600), .A2(n8601), .ZN(n8396) );
  NAND2_X1 U8528 ( .A1(b_28_), .A2(n8602), .ZN(n8601) );
  NAND2_X1 U8529 ( .A1(n7527), .A2(n8603), .ZN(n8602) );
  NAND2_X1 U8530 ( .A1(a_31_), .A2(n7547), .ZN(n8603) );
  NAND2_X1 U8531 ( .A1(b_29_), .A2(n8604), .ZN(n8600) );
  NAND2_X1 U8532 ( .A1(n7531), .A2(n8605), .ZN(n8604) );
  NAND2_X1 U8533 ( .A1(a_30_), .A2(n8037), .ZN(n8605) );
  AND3_X1 U8534 ( .A1(b_29_), .A2(b_30_), .A3(n7494), .ZN(n8397) );
  XNOR2_X1 U8535 ( .A(n8606), .B(n7542), .ZN(n8379) );
  XOR2_X1 U8536 ( .A(n8607), .B(n8608), .Z(n8606) );
  XNOR2_X1 U8537 ( .A(n8609), .B(n8610), .ZN(n8403) );
  NAND2_X1 U8538 ( .A1(n8611), .A2(n8612), .ZN(n8609) );
  XNOR2_X1 U8539 ( .A(n8613), .B(n8614), .ZN(n8356) );
  XNOR2_X1 U8540 ( .A(n8615), .B(n8616), .ZN(n8613) );
  XNOR2_X1 U8541 ( .A(n8617), .B(n8618), .ZN(n8406) );
  XOR2_X1 U8542 ( .A(n8619), .B(n8620), .Z(n8618) );
  NAND2_X1 U8543 ( .A1(a_24_), .A2(b_29_), .ZN(n8620) );
  XNOR2_X1 U8544 ( .A(n8621), .B(n8622), .ZN(n8411) );
  XNOR2_X1 U8545 ( .A(n8623), .B(n8624), .ZN(n8622) );
  XNOR2_X1 U8546 ( .A(n8625), .B(n8626), .ZN(n8415) );
  XOR2_X1 U8547 ( .A(n8627), .B(n8628), .Z(n8626) );
  NAND2_X1 U8548 ( .A1(a_22_), .A2(b_29_), .ZN(n8628) );
  XOR2_X1 U8549 ( .A(n8629), .B(n8630), .Z(n8418) );
  XOR2_X1 U8550 ( .A(n8631), .B(n8632), .Z(n8629) );
  XNOR2_X1 U8551 ( .A(n8633), .B(n8634), .ZN(n8422) );
  XNOR2_X1 U8552 ( .A(n8635), .B(n8636), .ZN(n8633) );
  NOR2_X1 U8553 ( .A1(n7547), .A2(n8044), .ZN(n8636) );
  XOR2_X1 U8554 ( .A(n8637), .B(n8638), .Z(n8427) );
  XNOR2_X1 U8555 ( .A(n8639), .B(n8640), .ZN(n8638) );
  XNOR2_X1 U8556 ( .A(n8641), .B(n8642), .ZN(n8430) );
  XNOR2_X1 U8557 ( .A(n8643), .B(n8644), .ZN(n8641) );
  NOR2_X1 U8558 ( .A1(n7547), .A2(n8047), .ZN(n8644) );
  XNOR2_X1 U8559 ( .A(n8645), .B(n8646), .ZN(n8435) );
  XOR2_X1 U8560 ( .A(n8647), .B(n8648), .Z(n8645) );
  XNOR2_X1 U8561 ( .A(n8649), .B(n8650), .ZN(n8439) );
  XOR2_X1 U8562 ( .A(n8651), .B(n8652), .Z(n8650) );
  NAND2_X1 U8563 ( .A1(a_16_), .A2(b_29_), .ZN(n8652) );
  XOR2_X1 U8564 ( .A(n8653), .B(n8654), .Z(n8444) );
  XNOR2_X1 U8565 ( .A(n8655), .B(n8656), .ZN(n8654) );
  XNOR2_X1 U8566 ( .A(n8657), .B(n8658), .ZN(n8448) );
  XNOR2_X1 U8567 ( .A(n8659), .B(n8660), .ZN(n8657) );
  NOR2_X1 U8568 ( .A1(n7547), .A2(n8049), .ZN(n8660) );
  XOR2_X1 U8569 ( .A(n8661), .B(n8662), .Z(n8451) );
  XOR2_X1 U8570 ( .A(n8663), .B(n8664), .Z(n8661) );
  XNOR2_X1 U8571 ( .A(n8665), .B(n8666), .ZN(n8455) );
  XNOR2_X1 U8572 ( .A(n8667), .B(n8668), .ZN(n8665) );
  NOR2_X1 U8573 ( .A1(n7547), .A2(n8669), .ZN(n8668) );
  XNOR2_X1 U8574 ( .A(n8670), .B(n8671), .ZN(n8460) );
  XNOR2_X1 U8575 ( .A(n8672), .B(n8673), .ZN(n8671) );
  XNOR2_X1 U8576 ( .A(n8674), .B(n8675), .ZN(n8464) );
  XNOR2_X1 U8577 ( .A(n8676), .B(n8677), .ZN(n8674) );
  NOR2_X1 U8578 ( .A1(n7547), .A2(n8051), .ZN(n8677) );
  XOR2_X1 U8579 ( .A(n8678), .B(n8679), .Z(n8467) );
  XOR2_X1 U8580 ( .A(n8680), .B(n8681), .Z(n8678) );
  XOR2_X1 U8581 ( .A(n8682), .B(n8683), .Z(n8471) );
  XOR2_X1 U8582 ( .A(n8684), .B(n8685), .Z(n8682) );
  NOR2_X1 U8583 ( .A1(n7547), .A2(n8686), .ZN(n8685) );
  XOR2_X1 U8584 ( .A(n8687), .B(n8688), .Z(n8476) );
  XNOR2_X1 U8585 ( .A(n8689), .B(n8690), .ZN(n8688) );
  XNOR2_X1 U8586 ( .A(n8691), .B(n8692), .ZN(n8480) );
  XOR2_X1 U8587 ( .A(n8693), .B(n8694), .Z(n8691) );
  NOR2_X1 U8588 ( .A1(n7547), .A2(n7887), .ZN(n8694) );
  XOR2_X1 U8589 ( .A(n8695), .B(n8696), .Z(n8483) );
  XOR2_X1 U8590 ( .A(n8697), .B(n8698), .Z(n8695) );
  XNOR2_X1 U8591 ( .A(n8699), .B(n8700), .ZN(n8487) );
  XNOR2_X1 U8592 ( .A(n8701), .B(n8702), .ZN(n8699) );
  NOR2_X1 U8593 ( .A1(n7547), .A2(n7916), .ZN(n8702) );
  XOR2_X1 U8594 ( .A(n8703), .B(n8704), .Z(n8492) );
  XOR2_X1 U8595 ( .A(n8705), .B(n8706), .Z(n8704) );
  NAND2_X1 U8596 ( .A1(a_3_), .A2(b_29_), .ZN(n8706) );
  XNOR2_X1 U8597 ( .A(n8707), .B(n8708), .ZN(n8496) );
  XOR2_X1 U8598 ( .A(n8709), .B(n8710), .Z(n8708) );
  XNOR2_X1 U8599 ( .A(n8711), .B(n8712), .ZN(n8278) );
  XNOR2_X1 U8600 ( .A(n8713), .B(n8714), .ZN(n8711) );
  NOR2_X1 U8601 ( .A1(n7957), .A2(n7547), .ZN(n8714) );
  NAND2_X1 U8602 ( .A1(n8276), .A2(n8277), .ZN(n8499) );
  XNOR2_X1 U8603 ( .A(n8715), .B(n8716), .ZN(n8274) );
  NAND2_X1 U8604 ( .A1(n8717), .A2(n8718), .ZN(n8715) );
  AND2_X1 U8605 ( .A1(n8270), .A2(n8269), .ZN(n8077) );
  NAND2_X1 U8606 ( .A1(n8266), .A2(n8719), .ZN(n8269) );
  NAND2_X1 U8607 ( .A1(n8720), .A2(n8721), .ZN(n8719) );
  OR2_X1 U8608 ( .A1(n8277), .A2(n8276), .ZN(n8270) );
  AND2_X1 U8609 ( .A1(n8717), .A2(n8722), .ZN(n8276) );
  NAND2_X1 U8610 ( .A1(n8716), .A2(n8718), .ZN(n8722) );
  NAND2_X1 U8611 ( .A1(n8723), .A2(n8724), .ZN(n8718) );
  NAND2_X1 U8612 ( .A1(a_0_), .A2(b_29_), .ZN(n8724) );
  INV_X1 U8613 ( .A(n8725), .ZN(n8723) );
  XOR2_X1 U8614 ( .A(n8726), .B(n8727), .Z(n8716) );
  XOR2_X1 U8615 ( .A(n8728), .B(n8729), .Z(n8726) );
  NAND2_X1 U8616 ( .A1(a_0_), .A2(n8725), .ZN(n8717) );
  NAND2_X1 U8617 ( .A1(n8730), .A2(n8731), .ZN(n8725) );
  NAND3_X1 U8618 ( .A1(a_1_), .A2(n8732), .A3(b_29_), .ZN(n8731) );
  NAND2_X1 U8619 ( .A1(n8713), .A2(n8712), .ZN(n8732) );
  OR2_X1 U8620 ( .A1(n8712), .A2(n8713), .ZN(n8730) );
  AND2_X1 U8621 ( .A1(n8733), .A2(n8734), .ZN(n8713) );
  NAND2_X1 U8622 ( .A1(n8709), .A2(n8735), .ZN(n8734) );
  NAND2_X1 U8623 ( .A1(n8736), .A2(n8710), .ZN(n8735) );
  INV_X1 U8624 ( .A(n8707), .ZN(n8736) );
  NAND2_X1 U8625 ( .A1(n8737), .A2(n8738), .ZN(n8709) );
  NAND3_X1 U8626 ( .A1(b_29_), .A2(n8739), .A3(a_3_), .ZN(n8738) );
  OR2_X1 U8627 ( .A1(n8705), .A2(n8703), .ZN(n8739) );
  NAND2_X1 U8628 ( .A1(n8703), .A2(n8705), .ZN(n8737) );
  NAND2_X1 U8629 ( .A1(n8740), .A2(n8741), .ZN(n8705) );
  NAND3_X1 U8630 ( .A1(b_29_), .A2(n8742), .A3(a_4_), .ZN(n8741) );
  NAND2_X1 U8631 ( .A1(n8701), .A2(n8700), .ZN(n8742) );
  OR2_X1 U8632 ( .A1(n8700), .A2(n8701), .ZN(n8740) );
  AND2_X1 U8633 ( .A1(n8743), .A2(n8744), .ZN(n8701) );
  NAND2_X1 U8634 ( .A1(n8698), .A2(n8745), .ZN(n8744) );
  OR2_X1 U8635 ( .A1(n8697), .A2(n8696), .ZN(n8745) );
  NOR2_X1 U8636 ( .A1(n7908), .A2(n7547), .ZN(n8698) );
  NAND2_X1 U8637 ( .A1(n8696), .A2(n8697), .ZN(n8743) );
  NAND2_X1 U8638 ( .A1(n8746), .A2(n8747), .ZN(n8697) );
  NAND3_X1 U8639 ( .A1(b_29_), .A2(n8748), .A3(a_6_), .ZN(n8747) );
  OR2_X1 U8640 ( .A1(n8693), .A2(n8692), .ZN(n8748) );
  NAND2_X1 U8641 ( .A1(n8692), .A2(n8693), .ZN(n8746) );
  NAND2_X1 U8642 ( .A1(n8749), .A2(n8750), .ZN(n8693) );
  NAND2_X1 U8643 ( .A1(n8690), .A2(n8751), .ZN(n8750) );
  OR2_X1 U8644 ( .A1(n8689), .A2(n8687), .ZN(n8751) );
  NOR2_X1 U8645 ( .A1(n7872), .A2(n7547), .ZN(n8690) );
  NAND2_X1 U8646 ( .A1(n8687), .A2(n8689), .ZN(n8749) );
  NAND2_X1 U8647 ( .A1(n8752), .A2(n8753), .ZN(n8689) );
  NAND3_X1 U8648 ( .A1(b_29_), .A2(n8754), .A3(a_8_), .ZN(n8753) );
  OR2_X1 U8649 ( .A1(n8684), .A2(n8683), .ZN(n8754) );
  NAND2_X1 U8650 ( .A1(n8683), .A2(n8684), .ZN(n8752) );
  NAND2_X1 U8651 ( .A1(n8755), .A2(n8756), .ZN(n8684) );
  NAND2_X1 U8652 ( .A1(n8681), .A2(n8757), .ZN(n8756) );
  OR2_X1 U8653 ( .A1(n8680), .A2(n8679), .ZN(n8757) );
  NOR2_X1 U8654 ( .A1(n8052), .A2(n7547), .ZN(n8681) );
  NAND2_X1 U8655 ( .A1(n8679), .A2(n8680), .ZN(n8755) );
  NAND2_X1 U8656 ( .A1(n8758), .A2(n8759), .ZN(n8680) );
  NAND3_X1 U8657 ( .A1(b_29_), .A2(n8760), .A3(a_10_), .ZN(n8759) );
  NAND2_X1 U8658 ( .A1(n8676), .A2(n8675), .ZN(n8760) );
  OR2_X1 U8659 ( .A1(n8675), .A2(n8676), .ZN(n8758) );
  AND2_X1 U8660 ( .A1(n8761), .A2(n8762), .ZN(n8676) );
  NAND2_X1 U8661 ( .A1(n8673), .A2(n8763), .ZN(n8762) );
  OR2_X1 U8662 ( .A1(n8672), .A2(n8670), .ZN(n8763) );
  NOR2_X1 U8663 ( .A1(n7811), .A2(n7547), .ZN(n8673) );
  NAND2_X1 U8664 ( .A1(n8670), .A2(n8672), .ZN(n8761) );
  NAND2_X1 U8665 ( .A1(n8764), .A2(n8765), .ZN(n8672) );
  NAND3_X1 U8666 ( .A1(b_29_), .A2(n8766), .A3(a_12_), .ZN(n8765) );
  NAND2_X1 U8667 ( .A1(n8667), .A2(n8666), .ZN(n8766) );
  OR2_X1 U8668 ( .A1(n8666), .A2(n8667), .ZN(n8764) );
  AND2_X1 U8669 ( .A1(n8767), .A2(n8768), .ZN(n8667) );
  NAND2_X1 U8670 ( .A1(n8664), .A2(n8769), .ZN(n8768) );
  OR2_X1 U8671 ( .A1(n8663), .A2(n8662), .ZN(n8769) );
  NOR2_X1 U8672 ( .A1(n7789), .A2(n7547), .ZN(n8664) );
  NAND2_X1 U8673 ( .A1(n8662), .A2(n8663), .ZN(n8767) );
  NAND2_X1 U8674 ( .A1(n8770), .A2(n8771), .ZN(n8663) );
  NAND3_X1 U8675 ( .A1(b_29_), .A2(n8772), .A3(a_14_), .ZN(n8771) );
  NAND2_X1 U8676 ( .A1(n8659), .A2(n8658), .ZN(n8772) );
  OR2_X1 U8677 ( .A1(n8658), .A2(n8659), .ZN(n8770) );
  AND2_X1 U8678 ( .A1(n8773), .A2(n8774), .ZN(n8659) );
  NAND2_X1 U8679 ( .A1(n8656), .A2(n8775), .ZN(n8774) );
  OR2_X1 U8680 ( .A1(n8655), .A2(n8653), .ZN(n8775) );
  NOR2_X1 U8681 ( .A1(n7754), .A2(n7547), .ZN(n8656) );
  NAND2_X1 U8682 ( .A1(n8653), .A2(n8655), .ZN(n8773) );
  NAND2_X1 U8683 ( .A1(n8776), .A2(n8777), .ZN(n8655) );
  NAND3_X1 U8684 ( .A1(b_29_), .A2(n8778), .A3(a_16_), .ZN(n8777) );
  OR2_X1 U8685 ( .A1(n8651), .A2(n8649), .ZN(n8778) );
  NAND2_X1 U8686 ( .A1(n8649), .A2(n8651), .ZN(n8776) );
  NAND2_X1 U8687 ( .A1(n8779), .A2(n8780), .ZN(n8651) );
  NAND2_X1 U8688 ( .A1(n8648), .A2(n8781), .ZN(n8780) );
  OR2_X1 U8689 ( .A1(n8647), .A2(n8646), .ZN(n8781) );
  NOR2_X1 U8690 ( .A1(n7732), .A2(n7547), .ZN(n8648) );
  NAND2_X1 U8691 ( .A1(n8646), .A2(n8647), .ZN(n8779) );
  NAND2_X1 U8692 ( .A1(n8782), .A2(n8783), .ZN(n8647) );
  NAND3_X1 U8693 ( .A1(b_29_), .A2(n8784), .A3(a_18_), .ZN(n8783) );
  NAND2_X1 U8694 ( .A1(n8643), .A2(n8642), .ZN(n8784) );
  OR2_X1 U8695 ( .A1(n8642), .A2(n8643), .ZN(n8782) );
  AND2_X1 U8696 ( .A1(n8785), .A2(n8786), .ZN(n8643) );
  NAND2_X1 U8697 ( .A1(n8640), .A2(n8787), .ZN(n8786) );
  OR2_X1 U8698 ( .A1(n8639), .A2(n8637), .ZN(n8787) );
  NOR2_X1 U8699 ( .A1(n8045), .A2(n7547), .ZN(n8640) );
  NAND2_X1 U8700 ( .A1(n8637), .A2(n8639), .ZN(n8785) );
  NAND2_X1 U8701 ( .A1(n8788), .A2(n8789), .ZN(n8639) );
  NAND3_X1 U8702 ( .A1(b_29_), .A2(n8790), .A3(a_20_), .ZN(n8789) );
  NAND2_X1 U8703 ( .A1(n8635), .A2(n8634), .ZN(n8790) );
  OR2_X1 U8704 ( .A1(n8634), .A2(n8635), .ZN(n8788) );
  AND2_X1 U8705 ( .A1(n8791), .A2(n8792), .ZN(n8635) );
  NAND2_X1 U8706 ( .A1(n8632), .A2(n8793), .ZN(n8792) );
  OR2_X1 U8707 ( .A1(n8631), .A2(n8630), .ZN(n8793) );
  NOR2_X1 U8708 ( .A1(n7665), .A2(n7547), .ZN(n8632) );
  NAND2_X1 U8709 ( .A1(n8630), .A2(n8631), .ZN(n8791) );
  NAND2_X1 U8710 ( .A1(n8794), .A2(n8795), .ZN(n8631) );
  NAND3_X1 U8711 ( .A1(b_29_), .A2(n8796), .A3(a_22_), .ZN(n8795) );
  OR2_X1 U8712 ( .A1(n8627), .A2(n8625), .ZN(n8796) );
  NAND2_X1 U8713 ( .A1(n8625), .A2(n8627), .ZN(n8794) );
  NAND2_X1 U8714 ( .A1(n8797), .A2(n8798), .ZN(n8627) );
  NAND2_X1 U8715 ( .A1(n8624), .A2(n8799), .ZN(n8798) );
  OR2_X1 U8716 ( .A1(n8623), .A2(n8621), .ZN(n8799) );
  NOR2_X1 U8717 ( .A1(n8042), .A2(n7547), .ZN(n8624) );
  NAND2_X1 U8718 ( .A1(n8621), .A2(n8623), .ZN(n8797) );
  NAND2_X1 U8719 ( .A1(n8800), .A2(n8801), .ZN(n8623) );
  NAND3_X1 U8720 ( .A1(b_29_), .A2(n8802), .A3(a_24_), .ZN(n8801) );
  OR2_X1 U8721 ( .A1(n8619), .A2(n8617), .ZN(n8802) );
  NAND2_X1 U8722 ( .A1(n8617), .A2(n8619), .ZN(n8800) );
  NAND2_X1 U8723 ( .A1(n8803), .A2(n8804), .ZN(n8619) );
  NAND2_X1 U8724 ( .A1(n8616), .A2(n8805), .ZN(n8804) );
  NAND2_X1 U8725 ( .A1(n8615), .A2(n8614), .ZN(n8805) );
  NOR2_X1 U8726 ( .A1(n8039), .A2(n7547), .ZN(n8616) );
  OR2_X1 U8727 ( .A1(n8614), .A2(n8615), .ZN(n8803) );
  AND2_X1 U8728 ( .A1(n8611), .A2(n8806), .ZN(n8615) );
  NAND2_X1 U8729 ( .A1(n8610), .A2(n8612), .ZN(n8806) );
  NAND2_X1 U8730 ( .A1(n8807), .A2(n8808), .ZN(n8612) );
  NAND2_X1 U8731 ( .A1(a_26_), .A2(b_29_), .ZN(n8808) );
  INV_X1 U8732 ( .A(n8809), .ZN(n8807) );
  XNOR2_X1 U8733 ( .A(n8810), .B(n8811), .ZN(n8610) );
  NAND2_X1 U8734 ( .A1(n8812), .A2(n8813), .ZN(n8810) );
  NAND2_X1 U8735 ( .A1(a_26_), .A2(n8809), .ZN(n8611) );
  NAND2_X1 U8736 ( .A1(n8584), .A2(n8814), .ZN(n8809) );
  NAND2_X1 U8737 ( .A1(n8583), .A2(n8585), .ZN(n8814) );
  NAND2_X1 U8738 ( .A1(n8815), .A2(n8816), .ZN(n8585) );
  NAND2_X1 U8739 ( .A1(a_27_), .A2(b_29_), .ZN(n8816) );
  INV_X1 U8740 ( .A(n8817), .ZN(n8815) );
  XOR2_X1 U8741 ( .A(n8818), .B(n8819), .Z(n8583) );
  XOR2_X1 U8742 ( .A(n7564), .B(n8820), .Z(n8818) );
  NAND2_X1 U8743 ( .A1(a_27_), .A2(n8817), .ZN(n8584) );
  NAND2_X1 U8744 ( .A1(n8821), .A2(n8822), .ZN(n8817) );
  NAND3_X1 U8745 ( .A1(b_29_), .A2(n8823), .A3(a_28_), .ZN(n8822) );
  NAND2_X1 U8746 ( .A1(n8593), .A2(n8591), .ZN(n8823) );
  OR2_X1 U8747 ( .A1(n8591), .A2(n8593), .ZN(n8821) );
  AND2_X1 U8748 ( .A1(n8824), .A2(n8825), .ZN(n8593) );
  NAND2_X1 U8749 ( .A1(n7542), .A2(n8826), .ZN(n8825) );
  OR2_X1 U8750 ( .A1(n8607), .A2(n8608), .ZN(n8826) );
  INV_X1 U8751 ( .A(n8030), .ZN(n7542) );
  NAND2_X1 U8752 ( .A1(a_29_), .A2(b_29_), .ZN(n8030) );
  NAND2_X1 U8753 ( .A1(n8608), .A2(n8607), .ZN(n8824) );
  NAND2_X1 U8754 ( .A1(n8827), .A2(n8828), .ZN(n8607) );
  NAND2_X1 U8755 ( .A1(b_27_), .A2(n8829), .ZN(n8828) );
  NAND2_X1 U8756 ( .A1(n7527), .A2(n8830), .ZN(n8829) );
  NAND2_X1 U8757 ( .A1(a_31_), .A2(n8037), .ZN(n8830) );
  NAND2_X1 U8758 ( .A1(b_28_), .A2(n8831), .ZN(n8827) );
  NAND2_X1 U8759 ( .A1(n7531), .A2(n8832), .ZN(n8831) );
  NAND2_X1 U8760 ( .A1(a_30_), .A2(n7582), .ZN(n8832) );
  AND3_X1 U8761 ( .A1(b_28_), .A2(b_29_), .A3(n7494), .ZN(n8608) );
  XNOR2_X1 U8762 ( .A(n8833), .B(n8834), .ZN(n8591) );
  XOR2_X1 U8763 ( .A(n8835), .B(n8836), .Z(n8833) );
  XOR2_X1 U8764 ( .A(n8837), .B(n8838), .Z(n8614) );
  NAND2_X1 U8765 ( .A1(n8839), .A2(n8840), .ZN(n8837) );
  XOR2_X1 U8766 ( .A(n8841), .B(n8842), .Z(n8617) );
  XOR2_X1 U8767 ( .A(n8843), .B(n8844), .Z(n8841) );
  XOR2_X1 U8768 ( .A(n8845), .B(n8846), .Z(n8621) );
  XOR2_X1 U8769 ( .A(n8847), .B(n8848), .Z(n8845) );
  NOR2_X1 U8770 ( .A1(n8037), .A2(n8041), .ZN(n8848) );
  XNOR2_X1 U8771 ( .A(n8849), .B(n8850), .ZN(n8625) );
  XNOR2_X1 U8772 ( .A(n8851), .B(n8852), .ZN(n8850) );
  XNOR2_X1 U8773 ( .A(n8853), .B(n8854), .ZN(n8630) );
  XNOR2_X1 U8774 ( .A(n8855), .B(n8856), .ZN(n8853) );
  NOR2_X1 U8775 ( .A1(n8037), .A2(n7650), .ZN(n8856) );
  XOR2_X1 U8776 ( .A(n8857), .B(n8858), .Z(n8634) );
  XNOR2_X1 U8777 ( .A(n8859), .B(n8860), .ZN(n8858) );
  XNOR2_X1 U8778 ( .A(n8861), .B(n8862), .ZN(n8637) );
  XNOR2_X1 U8779 ( .A(n8863), .B(n8864), .ZN(n8861) );
  NOR2_X1 U8780 ( .A1(n8037), .A2(n8044), .ZN(n8864) );
  XOR2_X1 U8781 ( .A(n8865), .B(n8866), .Z(n8642) );
  XNOR2_X1 U8782 ( .A(n8867), .B(n8868), .ZN(n8866) );
  XNOR2_X1 U8783 ( .A(n8869), .B(n8870), .ZN(n8646) );
  XNOR2_X1 U8784 ( .A(n8871), .B(n8872), .ZN(n8869) );
  NOR2_X1 U8785 ( .A1(n8037), .A2(n8047), .ZN(n8872) );
  XOR2_X1 U8786 ( .A(n8873), .B(n8874), .Z(n8649) );
  XOR2_X1 U8787 ( .A(n8875), .B(n8876), .Z(n8873) );
  XNOR2_X1 U8788 ( .A(n8877), .B(n8878), .ZN(n8653) );
  XOR2_X1 U8789 ( .A(n8879), .B(n8880), .Z(n8878) );
  NAND2_X1 U8790 ( .A1(a_16_), .A2(b_28_), .ZN(n8880) );
  XOR2_X1 U8791 ( .A(n8881), .B(n8882), .Z(n8658) );
  XNOR2_X1 U8792 ( .A(n8883), .B(n8884), .ZN(n8882) );
  XNOR2_X1 U8793 ( .A(n8885), .B(n8886), .ZN(n8662) );
  XNOR2_X1 U8794 ( .A(n8887), .B(n8888), .ZN(n8885) );
  NOR2_X1 U8795 ( .A1(n8037), .A2(n8049), .ZN(n8888) );
  XNOR2_X1 U8796 ( .A(n8889), .B(n8890), .ZN(n8666) );
  XOR2_X1 U8797 ( .A(n8891), .B(n8892), .Z(n8889) );
  XNOR2_X1 U8798 ( .A(n8893), .B(n8894), .ZN(n8670) );
  XOR2_X1 U8799 ( .A(n8895), .B(n8896), .Z(n8894) );
  NAND2_X1 U8800 ( .A1(a_12_), .A2(b_28_), .ZN(n8896) );
  XOR2_X1 U8801 ( .A(n8897), .B(n8898), .Z(n8675) );
  XNOR2_X1 U8802 ( .A(n8899), .B(n8900), .ZN(n8898) );
  XNOR2_X1 U8803 ( .A(n8901), .B(n8902), .ZN(n8679) );
  XOR2_X1 U8804 ( .A(n8903), .B(n8904), .Z(n8901) );
  NAND2_X1 U8805 ( .A1(a_10_), .A2(b_28_), .ZN(n8903) );
  XNOR2_X1 U8806 ( .A(n8905), .B(n8906), .ZN(n8683) );
  XNOR2_X1 U8807 ( .A(n8907), .B(n8908), .ZN(n8905) );
  XNOR2_X1 U8808 ( .A(n8909), .B(n8910), .ZN(n8687) );
  XOR2_X1 U8809 ( .A(n8911), .B(n8912), .Z(n8910) );
  NAND2_X1 U8810 ( .A1(a_8_), .A2(b_28_), .ZN(n8912) );
  XNOR2_X1 U8811 ( .A(n8913), .B(n8914), .ZN(n8692) );
  XNOR2_X1 U8812 ( .A(n8915), .B(n8916), .ZN(n8914) );
  XNOR2_X1 U8813 ( .A(n8917), .B(n8918), .ZN(n8696) );
  XNOR2_X1 U8814 ( .A(n8919), .B(n8920), .ZN(n8917) );
  NOR2_X1 U8815 ( .A1(n8037), .A2(n7887), .ZN(n8920) );
  XNOR2_X1 U8816 ( .A(n8921), .B(n8922), .ZN(n8700) );
  XOR2_X1 U8817 ( .A(n8923), .B(n8924), .Z(n8921) );
  XNOR2_X1 U8818 ( .A(n8925), .B(n8926), .ZN(n8703) );
  XOR2_X1 U8819 ( .A(n8927), .B(n8928), .Z(n8926) );
  NAND2_X1 U8820 ( .A1(a_4_), .A2(b_28_), .ZN(n8928) );
  NAND2_X1 U8821 ( .A1(n8929), .A2(n8707), .ZN(n8733) );
  XNOR2_X1 U8822 ( .A(n8930), .B(n8931), .ZN(n8707) );
  XOR2_X1 U8823 ( .A(n8932), .B(n8933), .Z(n8931) );
  NAND2_X1 U8824 ( .A1(a_3_), .A2(b_28_), .ZN(n8933) );
  INV_X1 U8825 ( .A(n8710), .ZN(n8929) );
  NAND2_X1 U8826 ( .A1(a_2_), .A2(b_29_), .ZN(n8710) );
  XNOR2_X1 U8827 ( .A(n8934), .B(n8935), .ZN(n8712) );
  XOR2_X1 U8828 ( .A(n8936), .B(n8937), .Z(n8934) );
  XOR2_X1 U8829 ( .A(n8938), .B(n8939), .Z(n8277) );
  XNOR2_X1 U8830 ( .A(n8940), .B(n8941), .ZN(n8938) );
  NOR2_X1 U8831 ( .A1(n8037), .A2(n8942), .ZN(n8941) );
  INV_X1 U8832 ( .A(n8082), .ZN(n8264) );
  NOR2_X1 U8833 ( .A1(n8267), .A2(n8266), .ZN(n8082) );
  OR2_X1 U8834 ( .A1(n8721), .A2(n8720), .ZN(n8266) );
  AND2_X1 U8835 ( .A1(n8943), .A2(n8944), .ZN(n8720) );
  NAND3_X1 U8836 ( .A1(b_28_), .A2(n8945), .A3(a_0_), .ZN(n8944) );
  NAND2_X1 U8837 ( .A1(n8940), .A2(n8939), .ZN(n8945) );
  OR2_X1 U8838 ( .A1(n8939), .A2(n8940), .ZN(n8943) );
  AND2_X1 U8839 ( .A1(n8946), .A2(n8947), .ZN(n8940) );
  NAND2_X1 U8840 ( .A1(n8729), .A2(n8948), .ZN(n8947) );
  OR2_X1 U8841 ( .A1(n8728), .A2(n8727), .ZN(n8948) );
  NOR2_X1 U8842 ( .A1(n8037), .A2(n7957), .ZN(n8729) );
  NAND2_X1 U8843 ( .A1(n8727), .A2(n8728), .ZN(n8946) );
  NAND2_X1 U8844 ( .A1(n8949), .A2(n8950), .ZN(n8728) );
  NAND2_X1 U8845 ( .A1(n8936), .A2(n8951), .ZN(n8950) );
  OR2_X1 U8846 ( .A1(n8935), .A2(n8937), .ZN(n8951) );
  NAND2_X1 U8847 ( .A1(n8952), .A2(n8953), .ZN(n8936) );
  NAND3_X1 U8848 ( .A1(b_28_), .A2(n8954), .A3(a_3_), .ZN(n8953) );
  OR2_X1 U8849 ( .A1(n8932), .A2(n8930), .ZN(n8954) );
  NAND2_X1 U8850 ( .A1(n8930), .A2(n8932), .ZN(n8952) );
  NAND2_X1 U8851 ( .A1(n8955), .A2(n8956), .ZN(n8932) );
  NAND3_X1 U8852 ( .A1(b_28_), .A2(n8957), .A3(a_4_), .ZN(n8956) );
  OR2_X1 U8853 ( .A1(n8927), .A2(n8925), .ZN(n8957) );
  NAND2_X1 U8854 ( .A1(n8925), .A2(n8927), .ZN(n8955) );
  NAND2_X1 U8855 ( .A1(n8958), .A2(n8959), .ZN(n8927) );
  NAND2_X1 U8856 ( .A1(n8924), .A2(n8960), .ZN(n8959) );
  OR2_X1 U8857 ( .A1(n8923), .A2(n8922), .ZN(n8960) );
  NOR2_X1 U8858 ( .A1(n7908), .A2(n8037), .ZN(n8924) );
  NAND2_X1 U8859 ( .A1(n8922), .A2(n8923), .ZN(n8958) );
  NAND2_X1 U8860 ( .A1(n8961), .A2(n8962), .ZN(n8923) );
  NAND3_X1 U8861 ( .A1(b_28_), .A2(n8963), .A3(a_6_), .ZN(n8962) );
  NAND2_X1 U8862 ( .A1(n8919), .A2(n8918), .ZN(n8963) );
  OR2_X1 U8863 ( .A1(n8918), .A2(n8919), .ZN(n8961) );
  AND2_X1 U8864 ( .A1(n8964), .A2(n8965), .ZN(n8919) );
  NAND2_X1 U8865 ( .A1(n8916), .A2(n8966), .ZN(n8965) );
  OR2_X1 U8866 ( .A1(n8915), .A2(n8913), .ZN(n8966) );
  NOR2_X1 U8867 ( .A1(n7872), .A2(n8037), .ZN(n8916) );
  NAND2_X1 U8868 ( .A1(n8913), .A2(n8915), .ZN(n8964) );
  NAND2_X1 U8869 ( .A1(n8967), .A2(n8968), .ZN(n8915) );
  NAND3_X1 U8870 ( .A1(b_28_), .A2(n8969), .A3(a_8_), .ZN(n8968) );
  OR2_X1 U8871 ( .A1(n8911), .A2(n8909), .ZN(n8969) );
  NAND2_X1 U8872 ( .A1(n8909), .A2(n8911), .ZN(n8967) );
  NAND2_X1 U8873 ( .A1(n8970), .A2(n8971), .ZN(n8911) );
  NAND2_X1 U8874 ( .A1(n8908), .A2(n8972), .ZN(n8971) );
  NAND2_X1 U8875 ( .A1(n8907), .A2(n8906), .ZN(n8972) );
  NOR2_X1 U8876 ( .A1(n8052), .A2(n8037), .ZN(n8908) );
  OR2_X1 U8877 ( .A1(n8906), .A2(n8907), .ZN(n8970) );
  AND2_X1 U8878 ( .A1(n8973), .A2(n8974), .ZN(n8907) );
  NAND3_X1 U8879 ( .A1(b_28_), .A2(n8975), .A3(a_10_), .ZN(n8974) );
  NAND2_X1 U8880 ( .A1(n8904), .A2(n8902), .ZN(n8975) );
  OR2_X1 U8881 ( .A1(n8902), .A2(n8904), .ZN(n8973) );
  AND2_X1 U8882 ( .A1(n8976), .A2(n8977), .ZN(n8904) );
  NAND2_X1 U8883 ( .A1(n8900), .A2(n8978), .ZN(n8977) );
  OR2_X1 U8884 ( .A1(n8899), .A2(n8897), .ZN(n8978) );
  NOR2_X1 U8885 ( .A1(n7811), .A2(n8037), .ZN(n8900) );
  NAND2_X1 U8886 ( .A1(n8897), .A2(n8899), .ZN(n8976) );
  NAND2_X1 U8887 ( .A1(n8979), .A2(n8980), .ZN(n8899) );
  NAND3_X1 U8888 ( .A1(b_28_), .A2(n8981), .A3(a_12_), .ZN(n8980) );
  OR2_X1 U8889 ( .A1(n8895), .A2(n8893), .ZN(n8981) );
  NAND2_X1 U8890 ( .A1(n8893), .A2(n8895), .ZN(n8979) );
  NAND2_X1 U8891 ( .A1(n8982), .A2(n8983), .ZN(n8895) );
  NAND2_X1 U8892 ( .A1(n8892), .A2(n8984), .ZN(n8983) );
  OR2_X1 U8893 ( .A1(n8891), .A2(n8890), .ZN(n8984) );
  NOR2_X1 U8894 ( .A1(n7789), .A2(n8037), .ZN(n8892) );
  NAND2_X1 U8895 ( .A1(n8890), .A2(n8891), .ZN(n8982) );
  NAND2_X1 U8896 ( .A1(n8985), .A2(n8986), .ZN(n8891) );
  NAND3_X1 U8897 ( .A1(b_28_), .A2(n8987), .A3(a_14_), .ZN(n8986) );
  NAND2_X1 U8898 ( .A1(n8887), .A2(n8886), .ZN(n8987) );
  OR2_X1 U8899 ( .A1(n8886), .A2(n8887), .ZN(n8985) );
  AND2_X1 U8900 ( .A1(n8988), .A2(n8989), .ZN(n8887) );
  NAND2_X1 U8901 ( .A1(n8884), .A2(n8990), .ZN(n8989) );
  OR2_X1 U8902 ( .A1(n8883), .A2(n8881), .ZN(n8990) );
  NOR2_X1 U8903 ( .A1(n7754), .A2(n8037), .ZN(n8884) );
  NAND2_X1 U8904 ( .A1(n8881), .A2(n8883), .ZN(n8988) );
  NAND2_X1 U8905 ( .A1(n8991), .A2(n8992), .ZN(n8883) );
  NAND3_X1 U8906 ( .A1(b_28_), .A2(n8993), .A3(a_16_), .ZN(n8992) );
  OR2_X1 U8907 ( .A1(n8879), .A2(n8877), .ZN(n8993) );
  NAND2_X1 U8908 ( .A1(n8877), .A2(n8879), .ZN(n8991) );
  NAND2_X1 U8909 ( .A1(n8994), .A2(n8995), .ZN(n8879) );
  NAND2_X1 U8910 ( .A1(n8876), .A2(n8996), .ZN(n8995) );
  OR2_X1 U8911 ( .A1(n8875), .A2(n8874), .ZN(n8996) );
  NOR2_X1 U8912 ( .A1(n7732), .A2(n8037), .ZN(n8876) );
  NAND2_X1 U8913 ( .A1(n8874), .A2(n8875), .ZN(n8994) );
  NAND2_X1 U8914 ( .A1(n8997), .A2(n8998), .ZN(n8875) );
  NAND3_X1 U8915 ( .A1(b_28_), .A2(n8999), .A3(a_18_), .ZN(n8998) );
  NAND2_X1 U8916 ( .A1(n8871), .A2(n8870), .ZN(n8999) );
  OR2_X1 U8917 ( .A1(n8870), .A2(n8871), .ZN(n8997) );
  AND2_X1 U8918 ( .A1(n9000), .A2(n9001), .ZN(n8871) );
  NAND2_X1 U8919 ( .A1(n8868), .A2(n9002), .ZN(n9001) );
  OR2_X1 U8920 ( .A1(n8867), .A2(n8865), .ZN(n9002) );
  NOR2_X1 U8921 ( .A1(n8045), .A2(n8037), .ZN(n8868) );
  NAND2_X1 U8922 ( .A1(n8865), .A2(n8867), .ZN(n9000) );
  NAND2_X1 U8923 ( .A1(n9003), .A2(n9004), .ZN(n8867) );
  NAND3_X1 U8924 ( .A1(b_28_), .A2(n9005), .A3(a_20_), .ZN(n9004) );
  NAND2_X1 U8925 ( .A1(n8863), .A2(n8862), .ZN(n9005) );
  OR2_X1 U8926 ( .A1(n8862), .A2(n8863), .ZN(n9003) );
  AND2_X1 U8927 ( .A1(n9006), .A2(n9007), .ZN(n8863) );
  NAND2_X1 U8928 ( .A1(n8860), .A2(n9008), .ZN(n9007) );
  OR2_X1 U8929 ( .A1(n8859), .A2(n8857), .ZN(n9008) );
  NOR2_X1 U8930 ( .A1(n7665), .A2(n8037), .ZN(n8860) );
  NAND2_X1 U8931 ( .A1(n8857), .A2(n8859), .ZN(n9006) );
  NAND2_X1 U8932 ( .A1(n9009), .A2(n9010), .ZN(n8859) );
  NAND3_X1 U8933 ( .A1(b_28_), .A2(n9011), .A3(a_22_), .ZN(n9010) );
  NAND2_X1 U8934 ( .A1(n8855), .A2(n8854), .ZN(n9011) );
  OR2_X1 U8935 ( .A1(n8854), .A2(n8855), .ZN(n9009) );
  AND2_X1 U8936 ( .A1(n9012), .A2(n9013), .ZN(n8855) );
  NAND2_X1 U8937 ( .A1(n8852), .A2(n9014), .ZN(n9013) );
  OR2_X1 U8938 ( .A1(n8851), .A2(n8849), .ZN(n9014) );
  NOR2_X1 U8939 ( .A1(n8042), .A2(n8037), .ZN(n8852) );
  NAND2_X1 U8940 ( .A1(n8849), .A2(n8851), .ZN(n9012) );
  NAND2_X1 U8941 ( .A1(n9015), .A2(n9016), .ZN(n8851) );
  NAND3_X1 U8942 ( .A1(b_28_), .A2(n9017), .A3(a_24_), .ZN(n9016) );
  OR2_X1 U8943 ( .A1(n8847), .A2(n8846), .ZN(n9017) );
  NAND2_X1 U8944 ( .A1(n8846), .A2(n8847), .ZN(n9015) );
  NAND2_X1 U8945 ( .A1(n9018), .A2(n9019), .ZN(n8847) );
  NAND2_X1 U8946 ( .A1(n8844), .A2(n9020), .ZN(n9019) );
  OR2_X1 U8947 ( .A1(n8843), .A2(n8842), .ZN(n9020) );
  NOR2_X1 U8948 ( .A1(n8039), .A2(n8037), .ZN(n8844) );
  NAND2_X1 U8949 ( .A1(n8842), .A2(n8843), .ZN(n9018) );
  NAND2_X1 U8950 ( .A1(n8839), .A2(n9021), .ZN(n8843) );
  NAND2_X1 U8951 ( .A1(n8838), .A2(n8840), .ZN(n9021) );
  NAND2_X1 U8952 ( .A1(n9022), .A2(n9023), .ZN(n8840) );
  NAND2_X1 U8953 ( .A1(a_26_), .A2(b_28_), .ZN(n9023) );
  INV_X1 U8954 ( .A(n9024), .ZN(n9022) );
  XOR2_X1 U8955 ( .A(n9025), .B(n9026), .Z(n8838) );
  XOR2_X1 U8956 ( .A(n9027), .B(n7577), .Z(n9025) );
  NAND2_X1 U8957 ( .A1(a_26_), .A2(n9024), .ZN(n8839) );
  NAND2_X1 U8958 ( .A1(n8812), .A2(n9028), .ZN(n9024) );
  NAND2_X1 U8959 ( .A1(n8811), .A2(n8813), .ZN(n9028) );
  NAND2_X1 U8960 ( .A1(n9029), .A2(n9030), .ZN(n8813) );
  NAND2_X1 U8961 ( .A1(a_27_), .A2(b_28_), .ZN(n9030) );
  INV_X1 U8962 ( .A(n9031), .ZN(n9029) );
  XNOR2_X1 U8963 ( .A(n9032), .B(n9033), .ZN(n8811) );
  XOR2_X1 U8964 ( .A(n9034), .B(n9035), .Z(n9032) );
  NAND2_X1 U8965 ( .A1(b_27_), .A2(a_28_), .ZN(n9034) );
  NAND2_X1 U8966 ( .A1(a_27_), .A2(n9031), .ZN(n8812) );
  NAND2_X1 U8967 ( .A1(n9036), .A2(n9037), .ZN(n9031) );
  NAND2_X1 U8968 ( .A1(n8819), .A2(n9038), .ZN(n9037) );
  NAND2_X1 U8969 ( .A1(n8820), .A2(n7564), .ZN(n9038) );
  INV_X1 U8970 ( .A(n9039), .ZN(n8820) );
  XOR2_X1 U8971 ( .A(n9040), .B(n9041), .Z(n8819) );
  XOR2_X1 U8972 ( .A(n9042), .B(n9043), .Z(n9040) );
  NAND2_X1 U8973 ( .A1(n9044), .A2(n9039), .ZN(n9036) );
  NAND2_X1 U8974 ( .A1(n9045), .A2(n9046), .ZN(n9039) );
  NAND2_X1 U8975 ( .A1(n8834), .A2(n9047), .ZN(n9046) );
  OR2_X1 U8976 ( .A1(n8835), .A2(n8836), .ZN(n9047) );
  NOR2_X1 U8977 ( .A1(n8037), .A2(n7545), .ZN(n8834) );
  NAND2_X1 U8978 ( .A1(n8836), .A2(n8835), .ZN(n9045) );
  NAND2_X1 U8979 ( .A1(n9048), .A2(n9049), .ZN(n8835) );
  NAND2_X1 U8980 ( .A1(b_26_), .A2(n9050), .ZN(n9049) );
  NAND2_X1 U8981 ( .A1(n7527), .A2(n9051), .ZN(n9050) );
  NAND2_X1 U8982 ( .A1(a_31_), .A2(n7582), .ZN(n9051) );
  NAND2_X1 U8983 ( .A1(b_27_), .A2(n9052), .ZN(n9048) );
  NAND2_X1 U8984 ( .A1(n7531), .A2(n9053), .ZN(n9052) );
  NAND2_X1 U8985 ( .A1(a_30_), .A2(n8038), .ZN(n9053) );
  AND3_X1 U8986 ( .A1(b_28_), .A2(b_27_), .A3(n7494), .ZN(n8836) );
  INV_X1 U8987 ( .A(n7564), .ZN(n9044) );
  NAND2_X1 U8988 ( .A1(b_28_), .A2(a_28_), .ZN(n7564) );
  XNOR2_X1 U8989 ( .A(n9054), .B(n9055), .ZN(n8842) );
  NAND2_X1 U8990 ( .A1(n9056), .A2(n9057), .ZN(n9054) );
  XNOR2_X1 U8991 ( .A(n9058), .B(n9059), .ZN(n8846) );
  XNOR2_X1 U8992 ( .A(n9060), .B(n9061), .ZN(n9058) );
  XNOR2_X1 U8993 ( .A(n9062), .B(n9063), .ZN(n8849) );
  XOR2_X1 U8994 ( .A(n9064), .B(n9065), .Z(n9063) );
  NAND2_X1 U8995 ( .A1(a_24_), .A2(b_27_), .ZN(n9065) );
  XOR2_X1 U8996 ( .A(n9066), .B(n9067), .Z(n8854) );
  XNOR2_X1 U8997 ( .A(n9068), .B(n9069), .ZN(n9067) );
  XNOR2_X1 U8998 ( .A(n9070), .B(n9071), .ZN(n8857) );
  XOR2_X1 U8999 ( .A(n9072), .B(n9073), .Z(n9071) );
  NAND2_X1 U9000 ( .A1(a_22_), .A2(b_27_), .ZN(n9073) );
  XNOR2_X1 U9001 ( .A(n9074), .B(n9075), .ZN(n8862) );
  XOR2_X1 U9002 ( .A(n9076), .B(n9077), .Z(n9074) );
  XNOR2_X1 U9003 ( .A(n9078), .B(n9079), .ZN(n8865) );
  XNOR2_X1 U9004 ( .A(n9080), .B(n9081), .ZN(n9078) );
  NOR2_X1 U9005 ( .A1(n7582), .A2(n8044), .ZN(n9081) );
  XOR2_X1 U9006 ( .A(n9082), .B(n9083), .Z(n8870) );
  XNOR2_X1 U9007 ( .A(n9084), .B(n9085), .ZN(n9083) );
  XNOR2_X1 U9008 ( .A(n9086), .B(n9087), .ZN(n8874) );
  XNOR2_X1 U9009 ( .A(n9088), .B(n9089), .ZN(n9086) );
  NOR2_X1 U9010 ( .A1(n7582), .A2(n8047), .ZN(n9089) );
  XOR2_X1 U9011 ( .A(n9090), .B(n9091), .Z(n8877) );
  XOR2_X1 U9012 ( .A(n9092), .B(n9093), .Z(n9090) );
  XNOR2_X1 U9013 ( .A(n9094), .B(n9095), .ZN(n8881) );
  XNOR2_X1 U9014 ( .A(n9096), .B(n9097), .ZN(n9094) );
  NOR2_X1 U9015 ( .A1(n7582), .A2(n8438), .ZN(n9097) );
  XOR2_X1 U9016 ( .A(n9098), .B(n9099), .Z(n8886) );
  XNOR2_X1 U9017 ( .A(n9100), .B(n9101), .ZN(n9099) );
  XNOR2_X1 U9018 ( .A(n9102), .B(n9103), .ZN(n8890) );
  XNOR2_X1 U9019 ( .A(n9104), .B(n9105), .ZN(n9102) );
  NOR2_X1 U9020 ( .A1(n7582), .A2(n8049), .ZN(n9105) );
  XNOR2_X1 U9021 ( .A(n9106), .B(n9107), .ZN(n8893) );
  XNOR2_X1 U9022 ( .A(n9108), .B(n9109), .ZN(n9106) );
  XNOR2_X1 U9023 ( .A(n9110), .B(n9111), .ZN(n8897) );
  XOR2_X1 U9024 ( .A(n9112), .B(n9113), .Z(n9111) );
  NAND2_X1 U9025 ( .A1(a_12_), .A2(b_27_), .ZN(n9113) );
  XOR2_X1 U9026 ( .A(n9114), .B(n9115), .Z(n8902) );
  XNOR2_X1 U9027 ( .A(n9116), .B(n9117), .ZN(n9115) );
  XNOR2_X1 U9028 ( .A(n9118), .B(n9119), .ZN(n8906) );
  XOR2_X1 U9029 ( .A(n9120), .B(n9121), .Z(n9118) );
  NOR2_X1 U9030 ( .A1(n7582), .A2(n8051), .ZN(n9121) );
  XOR2_X1 U9031 ( .A(n9122), .B(n9123), .Z(n8909) );
  XOR2_X1 U9032 ( .A(n9124), .B(n9125), .Z(n9122) );
  XOR2_X1 U9033 ( .A(n9126), .B(n9127), .Z(n8913) );
  XOR2_X1 U9034 ( .A(n9128), .B(n9129), .Z(n9126) );
  NOR2_X1 U9035 ( .A1(n7582), .A2(n8686), .ZN(n9129) );
  XOR2_X1 U9036 ( .A(n9130), .B(n9131), .Z(n8918) );
  XOR2_X1 U9037 ( .A(n9132), .B(n9133), .Z(n9131) );
  NAND2_X1 U9038 ( .A1(a_7_), .A2(b_27_), .ZN(n9133) );
  XNOR2_X1 U9039 ( .A(n9134), .B(n9135), .ZN(n8922) );
  XNOR2_X1 U9040 ( .A(n9136), .B(n9137), .ZN(n9134) );
  NOR2_X1 U9041 ( .A1(n7582), .A2(n7887), .ZN(n9137) );
  XNOR2_X1 U9042 ( .A(n9138), .B(n9139), .ZN(n8925) );
  XNOR2_X1 U9043 ( .A(n9140), .B(n9141), .ZN(n9139) );
  XNOR2_X1 U9044 ( .A(n9142), .B(n9143), .ZN(n8930) );
  XNOR2_X1 U9045 ( .A(n9144), .B(n9145), .ZN(n9142) );
  NOR2_X1 U9046 ( .A1(n7582), .A2(n7916), .ZN(n9145) );
  NAND2_X1 U9047 ( .A1(n8937), .A2(n8935), .ZN(n8949) );
  XNOR2_X1 U9048 ( .A(n9146), .B(n9147), .ZN(n8935) );
  NAND2_X1 U9049 ( .A1(n9148), .A2(n9149), .ZN(n9146) );
  NOR2_X1 U9050 ( .A1(n8056), .A2(n8037), .ZN(n8937) );
  XNOR2_X1 U9051 ( .A(n9150), .B(n9151), .ZN(n8727) );
  NAND2_X1 U9052 ( .A1(n9152), .A2(n9153), .ZN(n9150) );
  XNOR2_X1 U9053 ( .A(n9154), .B(n9155), .ZN(n8939) );
  XOR2_X1 U9054 ( .A(n9156), .B(n9157), .Z(n9154) );
  NOR2_X1 U9055 ( .A1(n7957), .A2(n7582), .ZN(n9157) );
  XNOR2_X1 U9056 ( .A(n9158), .B(n9159), .ZN(n8721) );
  XNOR2_X1 U9057 ( .A(n9160), .B(n9161), .ZN(n9158) );
  NAND2_X1 U9058 ( .A1(n9162), .A2(n8263), .ZN(n8267) );
  INV_X1 U9059 ( .A(n9163), .ZN(n8263) );
  NAND2_X1 U9060 ( .A1(n9164), .A2(n9165), .ZN(n9162) );
  NAND2_X1 U9061 ( .A1(n9163), .A2(n9166), .ZN(n8087) );
  XOR2_X1 U9062 ( .A(n8260), .B(n8259), .Z(n9166) );
  NOR2_X1 U9063 ( .A1(n9165), .A2(n9164), .ZN(n9163) );
  XOR2_X1 U9064 ( .A(n9167), .B(n9168), .Z(n9164) );
  XNOR2_X1 U9065 ( .A(n9169), .B(n9170), .ZN(n9167) );
  NOR2_X1 U9066 ( .A1(n8038), .A2(n8942), .ZN(n9170) );
  NAND2_X1 U9067 ( .A1(n9171), .A2(n9172), .ZN(n9165) );
  NAND2_X1 U9068 ( .A1(n9160), .A2(n9173), .ZN(n9172) );
  NAND2_X1 U9069 ( .A1(n9161), .A2(n9159), .ZN(n9173) );
  AND2_X1 U9070 ( .A1(n9174), .A2(n9175), .ZN(n9160) );
  NAND3_X1 U9071 ( .A1(a_1_), .A2(n9176), .A3(b_27_), .ZN(n9175) );
  OR2_X1 U9072 ( .A1(n9156), .A2(n9155), .ZN(n9176) );
  NAND2_X1 U9073 ( .A1(n9155), .A2(n9156), .ZN(n9174) );
  NAND2_X1 U9074 ( .A1(n9152), .A2(n9177), .ZN(n9156) );
  NAND2_X1 U9075 ( .A1(n9151), .A2(n9153), .ZN(n9177) );
  NAND2_X1 U9076 ( .A1(n9178), .A2(n9179), .ZN(n9153) );
  NAND2_X1 U9077 ( .A1(a_2_), .A2(b_27_), .ZN(n9179) );
  INV_X1 U9078 ( .A(n9180), .ZN(n9178) );
  XNOR2_X1 U9079 ( .A(n9181), .B(n9182), .ZN(n9151) );
  XNOR2_X1 U9080 ( .A(n9183), .B(n9184), .ZN(n9181) );
  NOR2_X1 U9081 ( .A1(n8038), .A2(n7937), .ZN(n9184) );
  NAND2_X1 U9082 ( .A1(a_2_), .A2(n9180), .ZN(n9152) );
  NAND2_X1 U9083 ( .A1(n9148), .A2(n9185), .ZN(n9180) );
  NAND2_X1 U9084 ( .A1(n9147), .A2(n9149), .ZN(n9185) );
  NAND2_X1 U9085 ( .A1(n9186), .A2(n9187), .ZN(n9149) );
  NAND2_X1 U9086 ( .A1(a_3_), .A2(b_27_), .ZN(n9187) );
  INV_X1 U9087 ( .A(n9188), .ZN(n9186) );
  XNOR2_X1 U9088 ( .A(n9189), .B(n9190), .ZN(n9147) );
  XNOR2_X1 U9089 ( .A(n9191), .B(n9192), .ZN(n9190) );
  NAND2_X1 U9090 ( .A1(a_3_), .A2(n9188), .ZN(n9148) );
  NAND2_X1 U9091 ( .A1(n9193), .A2(n9194), .ZN(n9188) );
  NAND3_X1 U9092 ( .A1(b_27_), .A2(n9195), .A3(a_4_), .ZN(n9194) );
  NAND2_X1 U9093 ( .A1(n9144), .A2(n9143), .ZN(n9195) );
  OR2_X1 U9094 ( .A1(n9143), .A2(n9144), .ZN(n9193) );
  AND2_X1 U9095 ( .A1(n9196), .A2(n9197), .ZN(n9144) );
  NAND2_X1 U9096 ( .A1(n9141), .A2(n9198), .ZN(n9197) );
  OR2_X1 U9097 ( .A1(n9140), .A2(n9138), .ZN(n9198) );
  NOR2_X1 U9098 ( .A1(n7908), .A2(n7582), .ZN(n9141) );
  NAND2_X1 U9099 ( .A1(n9138), .A2(n9140), .ZN(n9196) );
  NAND2_X1 U9100 ( .A1(n9199), .A2(n9200), .ZN(n9140) );
  NAND3_X1 U9101 ( .A1(b_27_), .A2(n9201), .A3(a_6_), .ZN(n9200) );
  NAND2_X1 U9102 ( .A1(n9136), .A2(n9135), .ZN(n9201) );
  OR2_X1 U9103 ( .A1(n9135), .A2(n9136), .ZN(n9199) );
  AND2_X1 U9104 ( .A1(n9202), .A2(n9203), .ZN(n9136) );
  NAND3_X1 U9105 ( .A1(b_27_), .A2(n9204), .A3(a_7_), .ZN(n9203) );
  OR2_X1 U9106 ( .A1(n9132), .A2(n9130), .ZN(n9204) );
  NAND2_X1 U9107 ( .A1(n9130), .A2(n9132), .ZN(n9202) );
  NAND2_X1 U9108 ( .A1(n9205), .A2(n9206), .ZN(n9132) );
  NAND3_X1 U9109 ( .A1(b_27_), .A2(n9207), .A3(a_8_), .ZN(n9206) );
  OR2_X1 U9110 ( .A1(n9128), .A2(n9127), .ZN(n9207) );
  NAND2_X1 U9111 ( .A1(n9127), .A2(n9128), .ZN(n9205) );
  NAND2_X1 U9112 ( .A1(n9208), .A2(n9209), .ZN(n9128) );
  NAND2_X1 U9113 ( .A1(n9125), .A2(n9210), .ZN(n9209) );
  OR2_X1 U9114 ( .A1(n9124), .A2(n9123), .ZN(n9210) );
  NOR2_X1 U9115 ( .A1(n8052), .A2(n7582), .ZN(n9125) );
  NAND2_X1 U9116 ( .A1(n9123), .A2(n9124), .ZN(n9208) );
  NAND2_X1 U9117 ( .A1(n9211), .A2(n9212), .ZN(n9124) );
  NAND3_X1 U9118 ( .A1(b_27_), .A2(n9213), .A3(a_10_), .ZN(n9212) );
  OR2_X1 U9119 ( .A1(n9120), .A2(n9119), .ZN(n9213) );
  NAND2_X1 U9120 ( .A1(n9119), .A2(n9120), .ZN(n9211) );
  NAND2_X1 U9121 ( .A1(n9214), .A2(n9215), .ZN(n9120) );
  NAND2_X1 U9122 ( .A1(n9117), .A2(n9216), .ZN(n9215) );
  OR2_X1 U9123 ( .A1(n9116), .A2(n9114), .ZN(n9216) );
  NOR2_X1 U9124 ( .A1(n7811), .A2(n7582), .ZN(n9117) );
  NAND2_X1 U9125 ( .A1(n9114), .A2(n9116), .ZN(n9214) );
  NAND2_X1 U9126 ( .A1(n9217), .A2(n9218), .ZN(n9116) );
  NAND3_X1 U9127 ( .A1(b_27_), .A2(n9219), .A3(a_12_), .ZN(n9218) );
  OR2_X1 U9128 ( .A1(n9112), .A2(n9110), .ZN(n9219) );
  NAND2_X1 U9129 ( .A1(n9110), .A2(n9112), .ZN(n9217) );
  NAND2_X1 U9130 ( .A1(n9220), .A2(n9221), .ZN(n9112) );
  NAND2_X1 U9131 ( .A1(n9109), .A2(n9222), .ZN(n9221) );
  NAND2_X1 U9132 ( .A1(n9108), .A2(n9107), .ZN(n9222) );
  NOR2_X1 U9133 ( .A1(n7789), .A2(n7582), .ZN(n9109) );
  OR2_X1 U9134 ( .A1(n9107), .A2(n9108), .ZN(n9220) );
  AND2_X1 U9135 ( .A1(n9223), .A2(n9224), .ZN(n9108) );
  NAND3_X1 U9136 ( .A1(b_27_), .A2(n9225), .A3(a_14_), .ZN(n9224) );
  NAND2_X1 U9137 ( .A1(n9104), .A2(n9103), .ZN(n9225) );
  OR2_X1 U9138 ( .A1(n9103), .A2(n9104), .ZN(n9223) );
  AND2_X1 U9139 ( .A1(n9226), .A2(n9227), .ZN(n9104) );
  NAND2_X1 U9140 ( .A1(n9101), .A2(n9228), .ZN(n9227) );
  OR2_X1 U9141 ( .A1(n9100), .A2(n9098), .ZN(n9228) );
  NOR2_X1 U9142 ( .A1(n7754), .A2(n7582), .ZN(n9101) );
  NAND2_X1 U9143 ( .A1(n9098), .A2(n9100), .ZN(n9226) );
  NAND2_X1 U9144 ( .A1(n9229), .A2(n9230), .ZN(n9100) );
  NAND3_X1 U9145 ( .A1(b_27_), .A2(n9231), .A3(a_16_), .ZN(n9230) );
  NAND2_X1 U9146 ( .A1(n9096), .A2(n9095), .ZN(n9231) );
  OR2_X1 U9147 ( .A1(n9095), .A2(n9096), .ZN(n9229) );
  AND2_X1 U9148 ( .A1(n9232), .A2(n9233), .ZN(n9096) );
  NAND2_X1 U9149 ( .A1(n9093), .A2(n9234), .ZN(n9233) );
  OR2_X1 U9150 ( .A1(n9092), .A2(n9091), .ZN(n9234) );
  NOR2_X1 U9151 ( .A1(n7732), .A2(n7582), .ZN(n9093) );
  NAND2_X1 U9152 ( .A1(n9091), .A2(n9092), .ZN(n9232) );
  NAND2_X1 U9153 ( .A1(n9235), .A2(n9236), .ZN(n9092) );
  NAND3_X1 U9154 ( .A1(b_27_), .A2(n9237), .A3(a_18_), .ZN(n9236) );
  NAND2_X1 U9155 ( .A1(n9088), .A2(n9087), .ZN(n9237) );
  OR2_X1 U9156 ( .A1(n9087), .A2(n9088), .ZN(n9235) );
  AND2_X1 U9157 ( .A1(n9238), .A2(n9239), .ZN(n9088) );
  NAND2_X1 U9158 ( .A1(n9085), .A2(n9240), .ZN(n9239) );
  OR2_X1 U9159 ( .A1(n9084), .A2(n9082), .ZN(n9240) );
  NOR2_X1 U9160 ( .A1(n8045), .A2(n7582), .ZN(n9085) );
  NAND2_X1 U9161 ( .A1(n9082), .A2(n9084), .ZN(n9238) );
  NAND2_X1 U9162 ( .A1(n9241), .A2(n9242), .ZN(n9084) );
  NAND3_X1 U9163 ( .A1(b_27_), .A2(n9243), .A3(a_20_), .ZN(n9242) );
  NAND2_X1 U9164 ( .A1(n9080), .A2(n9079), .ZN(n9243) );
  OR2_X1 U9165 ( .A1(n9079), .A2(n9080), .ZN(n9241) );
  AND2_X1 U9166 ( .A1(n9244), .A2(n9245), .ZN(n9080) );
  NAND2_X1 U9167 ( .A1(n9077), .A2(n9246), .ZN(n9245) );
  OR2_X1 U9168 ( .A1(n9076), .A2(n9075), .ZN(n9246) );
  NOR2_X1 U9169 ( .A1(n7665), .A2(n7582), .ZN(n9077) );
  NAND2_X1 U9170 ( .A1(n9075), .A2(n9076), .ZN(n9244) );
  NAND2_X1 U9171 ( .A1(n9247), .A2(n9248), .ZN(n9076) );
  NAND3_X1 U9172 ( .A1(b_27_), .A2(n9249), .A3(a_22_), .ZN(n9248) );
  OR2_X1 U9173 ( .A1(n9072), .A2(n9070), .ZN(n9249) );
  NAND2_X1 U9174 ( .A1(n9070), .A2(n9072), .ZN(n9247) );
  NAND2_X1 U9175 ( .A1(n9250), .A2(n9251), .ZN(n9072) );
  NAND2_X1 U9176 ( .A1(n9069), .A2(n9252), .ZN(n9251) );
  OR2_X1 U9177 ( .A1(n9068), .A2(n9066), .ZN(n9252) );
  NOR2_X1 U9178 ( .A1(n8042), .A2(n7582), .ZN(n9069) );
  NAND2_X1 U9179 ( .A1(n9066), .A2(n9068), .ZN(n9250) );
  NAND2_X1 U9180 ( .A1(n9253), .A2(n9254), .ZN(n9068) );
  NAND3_X1 U9181 ( .A1(b_27_), .A2(n9255), .A3(a_24_), .ZN(n9254) );
  OR2_X1 U9182 ( .A1(n9064), .A2(n9062), .ZN(n9255) );
  NAND2_X1 U9183 ( .A1(n9062), .A2(n9064), .ZN(n9253) );
  NAND2_X1 U9184 ( .A1(n9256), .A2(n9257), .ZN(n9064) );
  NAND2_X1 U9185 ( .A1(n9061), .A2(n9258), .ZN(n9257) );
  NAND2_X1 U9186 ( .A1(n9060), .A2(n9059), .ZN(n9258) );
  NOR2_X1 U9187 ( .A1(n8039), .A2(n7582), .ZN(n9061) );
  OR2_X1 U9188 ( .A1(n9059), .A2(n9060), .ZN(n9256) );
  AND2_X1 U9189 ( .A1(n9056), .A2(n9259), .ZN(n9060) );
  NAND2_X1 U9190 ( .A1(n9055), .A2(n9057), .ZN(n9259) );
  NAND2_X1 U9191 ( .A1(n9260), .A2(n9261), .ZN(n9057) );
  NAND2_X1 U9192 ( .A1(a_26_), .A2(b_27_), .ZN(n9261) );
  INV_X1 U9193 ( .A(n9262), .ZN(n9260) );
  XNOR2_X1 U9194 ( .A(n9263), .B(n9264), .ZN(n9055) );
  NAND2_X1 U9195 ( .A1(n9265), .A2(n9266), .ZN(n9263) );
  NAND2_X1 U9196 ( .A1(a_26_), .A2(n9262), .ZN(n9056) );
  NAND2_X1 U9197 ( .A1(n9267), .A2(n9268), .ZN(n9262) );
  NAND2_X1 U9198 ( .A1(n9026), .A2(n9269), .ZN(n9268) );
  OR2_X1 U9199 ( .A1(n9027), .A2(n7577), .ZN(n9269) );
  XNOR2_X1 U9200 ( .A(n9270), .B(n9271), .ZN(n9026) );
  XOR2_X1 U9201 ( .A(n9272), .B(n9273), .Z(n9270) );
  NAND2_X1 U9202 ( .A1(b_26_), .A2(a_28_), .ZN(n9272) );
  NAND2_X1 U9203 ( .A1(n7577), .A2(n9027), .ZN(n9267) );
  NAND2_X1 U9204 ( .A1(n9274), .A2(n9275), .ZN(n9027) );
  NAND3_X1 U9205 ( .A1(a_28_), .A2(n9276), .A3(b_27_), .ZN(n9275) );
  NAND2_X1 U9206 ( .A1(n9035), .A2(n9033), .ZN(n9276) );
  OR2_X1 U9207 ( .A1(n9033), .A2(n9035), .ZN(n9274) );
  AND2_X1 U9208 ( .A1(n9277), .A2(n9278), .ZN(n9035) );
  NAND2_X1 U9209 ( .A1(n9041), .A2(n9279), .ZN(n9278) );
  OR2_X1 U9210 ( .A1(n9042), .A2(n9043), .ZN(n9279) );
  NOR2_X1 U9211 ( .A1(n7582), .A2(n7545), .ZN(n9041) );
  NAND2_X1 U9212 ( .A1(n9043), .A2(n9042), .ZN(n9277) );
  NAND2_X1 U9213 ( .A1(n9280), .A2(n9281), .ZN(n9042) );
  NAND2_X1 U9214 ( .A1(b_25_), .A2(n9282), .ZN(n9281) );
  NAND2_X1 U9215 ( .A1(n7527), .A2(n9283), .ZN(n9282) );
  NAND2_X1 U9216 ( .A1(a_31_), .A2(n8038), .ZN(n9283) );
  NAND2_X1 U9217 ( .A1(b_26_), .A2(n9284), .ZN(n9280) );
  NAND2_X1 U9218 ( .A1(n7531), .A2(n9285), .ZN(n9284) );
  NAND2_X1 U9219 ( .A1(a_30_), .A2(n7609), .ZN(n9285) );
  AND3_X1 U9220 ( .A1(b_26_), .A2(b_27_), .A3(n7494), .ZN(n9043) );
  XNOR2_X1 U9221 ( .A(n9286), .B(n9287), .ZN(n9033) );
  XOR2_X1 U9222 ( .A(n9288), .B(n9289), .Z(n9286) );
  INV_X1 U9223 ( .A(n8026), .ZN(n7577) );
  NAND2_X1 U9224 ( .A1(a_27_), .A2(b_27_), .ZN(n8026) );
  XNOR2_X1 U9225 ( .A(n9290), .B(n9291), .ZN(n9059) );
  XOR2_X1 U9226 ( .A(n9292), .B(n9293), .Z(n9290) );
  XOR2_X1 U9227 ( .A(n9294), .B(n9295), .Z(n9062) );
  XOR2_X1 U9228 ( .A(n9296), .B(n9297), .Z(n9294) );
  XNOR2_X1 U9229 ( .A(n9298), .B(n9299), .ZN(n9066) );
  XNOR2_X1 U9230 ( .A(n9300), .B(n9301), .ZN(n9298) );
  NOR2_X1 U9231 ( .A1(n8038), .A2(n8041), .ZN(n9301) );
  XNOR2_X1 U9232 ( .A(n9302), .B(n9303), .ZN(n9070) );
  XNOR2_X1 U9233 ( .A(n9304), .B(n9305), .ZN(n9303) );
  XNOR2_X1 U9234 ( .A(n9306), .B(n9307), .ZN(n9075) );
  XOR2_X1 U9235 ( .A(n9308), .B(n9309), .Z(n9307) );
  NAND2_X1 U9236 ( .A1(a_22_), .A2(b_26_), .ZN(n9309) );
  XNOR2_X1 U9237 ( .A(n9310), .B(n9311), .ZN(n9079) );
  XOR2_X1 U9238 ( .A(n9312), .B(n9313), .Z(n9310) );
  XNOR2_X1 U9239 ( .A(n9314), .B(n9315), .ZN(n9082) );
  XNOR2_X1 U9240 ( .A(n9316), .B(n9317), .ZN(n9314) );
  NOR2_X1 U9241 ( .A1(n8038), .A2(n8044), .ZN(n9317) );
  XOR2_X1 U9242 ( .A(n9318), .B(n9319), .Z(n9087) );
  XNOR2_X1 U9243 ( .A(n9320), .B(n9321), .ZN(n9319) );
  XNOR2_X1 U9244 ( .A(n9322), .B(n9323), .ZN(n9091) );
  XNOR2_X1 U9245 ( .A(n9324), .B(n9325), .ZN(n9322) );
  NOR2_X1 U9246 ( .A1(n8038), .A2(n8047), .ZN(n9325) );
  XNOR2_X1 U9247 ( .A(n9326), .B(n9327), .ZN(n9095) );
  XOR2_X1 U9248 ( .A(n9328), .B(n9329), .Z(n9326) );
  XNOR2_X1 U9249 ( .A(n9330), .B(n9331), .ZN(n9098) );
  XOR2_X1 U9250 ( .A(n9332), .B(n9333), .Z(n9331) );
  NAND2_X1 U9251 ( .A1(a_16_), .A2(b_26_), .ZN(n9333) );
  XOR2_X1 U9252 ( .A(n9334), .B(n9335), .Z(n9103) );
  XNOR2_X1 U9253 ( .A(n9336), .B(n9337), .ZN(n9335) );
  XNOR2_X1 U9254 ( .A(n9338), .B(n9339), .ZN(n9107) );
  XOR2_X1 U9255 ( .A(n9340), .B(n9341), .Z(n9338) );
  NOR2_X1 U9256 ( .A1(n8038), .A2(n8049), .ZN(n9341) );
  XOR2_X1 U9257 ( .A(n9342), .B(n9343), .Z(n9110) );
  XOR2_X1 U9258 ( .A(n9344), .B(n9345), .Z(n9342) );
  XNOR2_X1 U9259 ( .A(n9346), .B(n9347), .ZN(n9114) );
  XOR2_X1 U9260 ( .A(n9348), .B(n9349), .Z(n9347) );
  NAND2_X1 U9261 ( .A1(a_12_), .A2(b_26_), .ZN(n9349) );
  XNOR2_X1 U9262 ( .A(n9350), .B(n9351), .ZN(n9119) );
  XNOR2_X1 U9263 ( .A(n9352), .B(n9353), .ZN(n9351) );
  XNOR2_X1 U9264 ( .A(n9354), .B(n9355), .ZN(n9123) );
  XNOR2_X1 U9265 ( .A(n9356), .B(n9357), .ZN(n9354) );
  NOR2_X1 U9266 ( .A1(n8038), .A2(n8051), .ZN(n9357) );
  XNOR2_X1 U9267 ( .A(n9358), .B(n9359), .ZN(n9127) );
  XNOR2_X1 U9268 ( .A(n9360), .B(n9361), .ZN(n9358) );
  XNOR2_X1 U9269 ( .A(n9362), .B(n9363), .ZN(n9130) );
  XOR2_X1 U9270 ( .A(n9364), .B(n9365), .Z(n9363) );
  NAND2_X1 U9271 ( .A1(a_8_), .A2(b_26_), .ZN(n9365) );
  XOR2_X1 U9272 ( .A(n9366), .B(n9367), .Z(n9135) );
  NAND2_X1 U9273 ( .A1(n9368), .A2(n9369), .ZN(n9366) );
  XNOR2_X1 U9274 ( .A(n9370), .B(n9371), .ZN(n9138) );
  XOR2_X1 U9275 ( .A(n9372), .B(n9373), .Z(n9370) );
  NAND2_X1 U9276 ( .A1(a_6_), .A2(b_26_), .ZN(n9372) );
  XOR2_X1 U9277 ( .A(n9374), .B(n9375), .Z(n9143) );
  XOR2_X1 U9278 ( .A(n9376), .B(n9377), .Z(n9375) );
  NAND2_X1 U9279 ( .A1(a_5_), .A2(b_26_), .ZN(n9377) );
  XNOR2_X1 U9280 ( .A(n9378), .B(n9379), .ZN(n9155) );
  XNOR2_X1 U9281 ( .A(n9380), .B(n9381), .ZN(n9379) );
  OR2_X1 U9282 ( .A1(n9159), .A2(n9161), .ZN(n9171) );
  NOR2_X1 U9283 ( .A1(n8942), .A2(n7582), .ZN(n9161) );
  XNOR2_X1 U9284 ( .A(n9382), .B(n9383), .ZN(n9159) );
  XNOR2_X1 U9285 ( .A(n9384), .B(n9385), .ZN(n9382) );
  NAND4_X1 U9286 ( .A1(n8259), .A2(n8258), .A3(n8260), .A4(n8253), .ZN(n8092)
         );
  INV_X1 U9287 ( .A(n9386), .ZN(n8253) );
  NAND2_X1 U9288 ( .A1(n9387), .A2(n9388), .ZN(n8260) );
  NAND3_X1 U9289 ( .A1(b_26_), .A2(n9389), .A3(a_0_), .ZN(n9388) );
  NAND2_X1 U9290 ( .A1(n9169), .A2(n9168), .ZN(n9389) );
  OR2_X1 U9291 ( .A1(n9168), .A2(n9169), .ZN(n9387) );
  AND2_X1 U9292 ( .A1(n9390), .A2(n9391), .ZN(n9169) );
  NAND2_X1 U9293 ( .A1(n9385), .A2(n9392), .ZN(n9391) );
  NAND2_X1 U9294 ( .A1(n9384), .A2(n9383), .ZN(n9392) );
  NOR2_X1 U9295 ( .A1(n8038), .A2(n7957), .ZN(n9385) );
  OR2_X1 U9296 ( .A1(n9383), .A2(n9384), .ZN(n9390) );
  AND2_X1 U9297 ( .A1(n9393), .A2(n9394), .ZN(n9384) );
  NAND2_X1 U9298 ( .A1(n9381), .A2(n9395), .ZN(n9394) );
  OR2_X1 U9299 ( .A1(n9380), .A2(n9378), .ZN(n9395) );
  NOR2_X1 U9300 ( .A1(n8056), .A2(n8038), .ZN(n9381) );
  NAND2_X1 U9301 ( .A1(n9378), .A2(n9380), .ZN(n9393) );
  NAND2_X1 U9302 ( .A1(n9396), .A2(n9397), .ZN(n9380) );
  NAND3_X1 U9303 ( .A1(b_26_), .A2(n9398), .A3(a_3_), .ZN(n9397) );
  NAND2_X1 U9304 ( .A1(n9183), .A2(n9182), .ZN(n9398) );
  OR2_X1 U9305 ( .A1(n9182), .A2(n9183), .ZN(n9396) );
  AND2_X1 U9306 ( .A1(n9399), .A2(n9400), .ZN(n9183) );
  NAND2_X1 U9307 ( .A1(n9192), .A2(n9401), .ZN(n9400) );
  OR2_X1 U9308 ( .A1(n9191), .A2(n9189), .ZN(n9401) );
  NOR2_X1 U9309 ( .A1(n7916), .A2(n8038), .ZN(n9192) );
  NAND2_X1 U9310 ( .A1(n9189), .A2(n9191), .ZN(n9399) );
  NAND2_X1 U9311 ( .A1(n9402), .A2(n9403), .ZN(n9191) );
  NAND3_X1 U9312 ( .A1(b_26_), .A2(n9404), .A3(a_5_), .ZN(n9403) );
  OR2_X1 U9313 ( .A1(n9376), .A2(n9374), .ZN(n9404) );
  NAND2_X1 U9314 ( .A1(n9374), .A2(n9376), .ZN(n9402) );
  NAND2_X1 U9315 ( .A1(n9405), .A2(n9406), .ZN(n9376) );
  NAND3_X1 U9316 ( .A1(b_26_), .A2(n9407), .A3(a_6_), .ZN(n9406) );
  NAND2_X1 U9317 ( .A1(n9373), .A2(n9371), .ZN(n9407) );
  OR2_X1 U9318 ( .A1(n9371), .A2(n9373), .ZN(n9405) );
  AND2_X1 U9319 ( .A1(n9368), .A2(n9408), .ZN(n9373) );
  NAND2_X1 U9320 ( .A1(n9367), .A2(n9369), .ZN(n9408) );
  NAND2_X1 U9321 ( .A1(n9409), .A2(n9410), .ZN(n9369) );
  NAND2_X1 U9322 ( .A1(a_7_), .A2(b_26_), .ZN(n9410) );
  INV_X1 U9323 ( .A(n9411), .ZN(n9409) );
  XOR2_X1 U9324 ( .A(n9412), .B(n9413), .Z(n9367) );
  XOR2_X1 U9325 ( .A(n9414), .B(n9415), .Z(n9412) );
  NOR2_X1 U9326 ( .A1(n7609), .A2(n8686), .ZN(n9415) );
  NAND2_X1 U9327 ( .A1(a_7_), .A2(n9411), .ZN(n9368) );
  NAND2_X1 U9328 ( .A1(n9416), .A2(n9417), .ZN(n9411) );
  NAND3_X1 U9329 ( .A1(b_26_), .A2(n9418), .A3(a_8_), .ZN(n9417) );
  OR2_X1 U9330 ( .A1(n9364), .A2(n9362), .ZN(n9418) );
  NAND2_X1 U9331 ( .A1(n9362), .A2(n9364), .ZN(n9416) );
  NAND2_X1 U9332 ( .A1(n9419), .A2(n9420), .ZN(n9364) );
  NAND2_X1 U9333 ( .A1(n9361), .A2(n9421), .ZN(n9420) );
  NAND2_X1 U9334 ( .A1(n9360), .A2(n9359), .ZN(n9421) );
  NOR2_X1 U9335 ( .A1(n8052), .A2(n8038), .ZN(n9361) );
  OR2_X1 U9336 ( .A1(n9359), .A2(n9360), .ZN(n9419) );
  AND2_X1 U9337 ( .A1(n9422), .A2(n9423), .ZN(n9360) );
  NAND3_X1 U9338 ( .A1(b_26_), .A2(n9424), .A3(a_10_), .ZN(n9423) );
  NAND2_X1 U9339 ( .A1(n9356), .A2(n9355), .ZN(n9424) );
  OR2_X1 U9340 ( .A1(n9355), .A2(n9356), .ZN(n9422) );
  AND2_X1 U9341 ( .A1(n9425), .A2(n9426), .ZN(n9356) );
  NAND2_X1 U9342 ( .A1(n9353), .A2(n9427), .ZN(n9426) );
  OR2_X1 U9343 ( .A1(n9352), .A2(n9350), .ZN(n9427) );
  NOR2_X1 U9344 ( .A1(n7811), .A2(n8038), .ZN(n9353) );
  NAND2_X1 U9345 ( .A1(n9350), .A2(n9352), .ZN(n9425) );
  NAND2_X1 U9346 ( .A1(n9428), .A2(n9429), .ZN(n9352) );
  NAND3_X1 U9347 ( .A1(b_26_), .A2(n9430), .A3(a_12_), .ZN(n9429) );
  OR2_X1 U9348 ( .A1(n9348), .A2(n9346), .ZN(n9430) );
  NAND2_X1 U9349 ( .A1(n9346), .A2(n9348), .ZN(n9428) );
  NAND2_X1 U9350 ( .A1(n9431), .A2(n9432), .ZN(n9348) );
  NAND2_X1 U9351 ( .A1(n9345), .A2(n9433), .ZN(n9432) );
  OR2_X1 U9352 ( .A1(n9344), .A2(n9343), .ZN(n9433) );
  NOR2_X1 U9353 ( .A1(n7789), .A2(n8038), .ZN(n9345) );
  NAND2_X1 U9354 ( .A1(n9343), .A2(n9344), .ZN(n9431) );
  NAND2_X1 U9355 ( .A1(n9434), .A2(n9435), .ZN(n9344) );
  NAND3_X1 U9356 ( .A1(b_26_), .A2(n9436), .A3(a_14_), .ZN(n9435) );
  OR2_X1 U9357 ( .A1(n9340), .A2(n9339), .ZN(n9436) );
  NAND2_X1 U9358 ( .A1(n9339), .A2(n9340), .ZN(n9434) );
  NAND2_X1 U9359 ( .A1(n9437), .A2(n9438), .ZN(n9340) );
  NAND2_X1 U9360 ( .A1(n9337), .A2(n9439), .ZN(n9438) );
  OR2_X1 U9361 ( .A1(n9336), .A2(n9334), .ZN(n9439) );
  NOR2_X1 U9362 ( .A1(n7754), .A2(n8038), .ZN(n9337) );
  NAND2_X1 U9363 ( .A1(n9334), .A2(n9336), .ZN(n9437) );
  NAND2_X1 U9364 ( .A1(n9440), .A2(n9441), .ZN(n9336) );
  NAND3_X1 U9365 ( .A1(b_26_), .A2(n9442), .A3(a_16_), .ZN(n9441) );
  OR2_X1 U9366 ( .A1(n9332), .A2(n9330), .ZN(n9442) );
  NAND2_X1 U9367 ( .A1(n9330), .A2(n9332), .ZN(n9440) );
  NAND2_X1 U9368 ( .A1(n9443), .A2(n9444), .ZN(n9332) );
  NAND2_X1 U9369 ( .A1(n9329), .A2(n9445), .ZN(n9444) );
  OR2_X1 U9370 ( .A1(n9328), .A2(n9327), .ZN(n9445) );
  NOR2_X1 U9371 ( .A1(n7732), .A2(n8038), .ZN(n9329) );
  NAND2_X1 U9372 ( .A1(n9327), .A2(n9328), .ZN(n9443) );
  NAND2_X1 U9373 ( .A1(n9446), .A2(n9447), .ZN(n9328) );
  NAND3_X1 U9374 ( .A1(b_26_), .A2(n9448), .A3(a_18_), .ZN(n9447) );
  NAND2_X1 U9375 ( .A1(n9324), .A2(n9323), .ZN(n9448) );
  OR2_X1 U9376 ( .A1(n9323), .A2(n9324), .ZN(n9446) );
  AND2_X1 U9377 ( .A1(n9449), .A2(n9450), .ZN(n9324) );
  NAND2_X1 U9378 ( .A1(n9321), .A2(n9451), .ZN(n9450) );
  OR2_X1 U9379 ( .A1(n9320), .A2(n9318), .ZN(n9451) );
  NOR2_X1 U9380 ( .A1(n8045), .A2(n8038), .ZN(n9321) );
  NAND2_X1 U9381 ( .A1(n9318), .A2(n9320), .ZN(n9449) );
  NAND2_X1 U9382 ( .A1(n9452), .A2(n9453), .ZN(n9320) );
  NAND3_X1 U9383 ( .A1(b_26_), .A2(n9454), .A3(a_20_), .ZN(n9453) );
  NAND2_X1 U9384 ( .A1(n9316), .A2(n9315), .ZN(n9454) );
  OR2_X1 U9385 ( .A1(n9315), .A2(n9316), .ZN(n9452) );
  AND2_X1 U9386 ( .A1(n9455), .A2(n9456), .ZN(n9316) );
  NAND2_X1 U9387 ( .A1(n9313), .A2(n9457), .ZN(n9456) );
  OR2_X1 U9388 ( .A1(n9312), .A2(n9311), .ZN(n9457) );
  NOR2_X1 U9389 ( .A1(n7665), .A2(n8038), .ZN(n9313) );
  NAND2_X1 U9390 ( .A1(n9311), .A2(n9312), .ZN(n9455) );
  NAND2_X1 U9391 ( .A1(n9458), .A2(n9459), .ZN(n9312) );
  NAND3_X1 U9392 ( .A1(b_26_), .A2(n9460), .A3(a_22_), .ZN(n9459) );
  OR2_X1 U9393 ( .A1(n9308), .A2(n9306), .ZN(n9460) );
  NAND2_X1 U9394 ( .A1(n9306), .A2(n9308), .ZN(n9458) );
  NAND2_X1 U9395 ( .A1(n9461), .A2(n9462), .ZN(n9308) );
  NAND2_X1 U9396 ( .A1(n9305), .A2(n9463), .ZN(n9462) );
  OR2_X1 U9397 ( .A1(n9304), .A2(n9302), .ZN(n9463) );
  NOR2_X1 U9398 ( .A1(n8042), .A2(n8038), .ZN(n9305) );
  NAND2_X1 U9399 ( .A1(n9302), .A2(n9304), .ZN(n9461) );
  NAND2_X1 U9400 ( .A1(n9464), .A2(n9465), .ZN(n9304) );
  NAND3_X1 U9401 ( .A1(b_26_), .A2(n9466), .A3(a_24_), .ZN(n9465) );
  NAND2_X1 U9402 ( .A1(n9300), .A2(n9299), .ZN(n9466) );
  OR2_X1 U9403 ( .A1(n9299), .A2(n9300), .ZN(n9464) );
  AND2_X1 U9404 ( .A1(n9467), .A2(n9468), .ZN(n9300) );
  NAND2_X1 U9405 ( .A1(n9297), .A2(n9469), .ZN(n9468) );
  OR2_X1 U9406 ( .A1(n9296), .A2(n9295), .ZN(n9469) );
  NOR2_X1 U9407 ( .A1(n8039), .A2(n8038), .ZN(n9297) );
  NAND2_X1 U9408 ( .A1(n9295), .A2(n9296), .ZN(n9467) );
  NAND2_X1 U9409 ( .A1(n9470), .A2(n9471), .ZN(n9296) );
  NAND2_X1 U9410 ( .A1(n9291), .A2(n9472), .ZN(n9471) );
  OR2_X1 U9411 ( .A1(n9292), .A2(n9293), .ZN(n9472) );
  XNOR2_X1 U9412 ( .A(n9473), .B(n9474), .ZN(n9291) );
  NAND2_X1 U9413 ( .A1(n9475), .A2(n9476), .ZN(n9473) );
  NAND2_X1 U9414 ( .A1(n9293), .A2(n9292), .ZN(n9470) );
  NAND2_X1 U9415 ( .A1(n9265), .A2(n9477), .ZN(n9292) );
  NAND2_X1 U9416 ( .A1(n9264), .A2(n9266), .ZN(n9477) );
  NAND2_X1 U9417 ( .A1(n9478), .A2(n9479), .ZN(n9266) );
  NAND2_X1 U9418 ( .A1(b_26_), .A2(a_27_), .ZN(n9479) );
  INV_X1 U9419 ( .A(n9480), .ZN(n9478) );
  XNOR2_X1 U9420 ( .A(n9481), .B(n9482), .ZN(n9264) );
  XOR2_X1 U9421 ( .A(n9483), .B(n9484), .Z(n9481) );
  NAND2_X1 U9422 ( .A1(b_25_), .A2(a_28_), .ZN(n9483) );
  NAND2_X1 U9423 ( .A1(a_27_), .A2(n9480), .ZN(n9265) );
  NAND2_X1 U9424 ( .A1(n9485), .A2(n9486), .ZN(n9480) );
  NAND3_X1 U9425 ( .A1(a_28_), .A2(n9487), .A3(b_26_), .ZN(n9486) );
  NAND2_X1 U9426 ( .A1(n9273), .A2(n9271), .ZN(n9487) );
  OR2_X1 U9427 ( .A1(n9271), .A2(n9273), .ZN(n9485) );
  AND2_X1 U9428 ( .A1(n9488), .A2(n9489), .ZN(n9273) );
  NAND2_X1 U9429 ( .A1(n9287), .A2(n9490), .ZN(n9489) );
  OR2_X1 U9430 ( .A1(n9288), .A2(n9289), .ZN(n9490) );
  NOR2_X1 U9431 ( .A1(n8038), .A2(n7545), .ZN(n9287) );
  NAND2_X1 U9432 ( .A1(n9289), .A2(n9288), .ZN(n9488) );
  NAND2_X1 U9433 ( .A1(n9491), .A2(n9492), .ZN(n9288) );
  NAND2_X1 U9434 ( .A1(b_24_), .A2(n9493), .ZN(n9492) );
  NAND2_X1 U9435 ( .A1(n7527), .A2(n9494), .ZN(n9493) );
  NAND2_X1 U9436 ( .A1(a_31_), .A2(n7609), .ZN(n9494) );
  NAND2_X1 U9437 ( .A1(b_25_), .A2(n9495), .ZN(n9491) );
  NAND2_X1 U9438 ( .A1(n7531), .A2(n9496), .ZN(n9495) );
  NAND2_X1 U9439 ( .A1(a_30_), .A2(n8040), .ZN(n9496) );
  AND3_X1 U9440 ( .A1(b_26_), .A2(b_25_), .A3(n7494), .ZN(n9289) );
  XNOR2_X1 U9441 ( .A(n9497), .B(n9498), .ZN(n9271) );
  XOR2_X1 U9442 ( .A(n9499), .B(n9500), .Z(n9497) );
  INV_X1 U9443 ( .A(n7600), .ZN(n9293) );
  NAND2_X1 U9444 ( .A1(b_26_), .A2(a_26_), .ZN(n7600) );
  XNOR2_X1 U9445 ( .A(n9501), .B(n9502), .ZN(n9295) );
  NAND2_X1 U9446 ( .A1(n9503), .A2(n9504), .ZN(n9501) );
  XNOR2_X1 U9447 ( .A(n9505), .B(n9506), .ZN(n9299) );
  XOR2_X1 U9448 ( .A(n9507), .B(n7607), .Z(n9505) );
  XNOR2_X1 U9449 ( .A(n9508), .B(n9509), .ZN(n9302) );
  XNOR2_X1 U9450 ( .A(n9510), .B(n9511), .ZN(n9508) );
  NOR2_X1 U9451 ( .A1(n7609), .A2(n8041), .ZN(n9511) );
  XNOR2_X1 U9452 ( .A(n9512), .B(n9513), .ZN(n9306) );
  XNOR2_X1 U9453 ( .A(n9514), .B(n9515), .ZN(n9513) );
  XNOR2_X1 U9454 ( .A(n9516), .B(n9517), .ZN(n9311) );
  XOR2_X1 U9455 ( .A(n9518), .B(n9519), .Z(n9517) );
  NAND2_X1 U9456 ( .A1(a_22_), .A2(b_25_), .ZN(n9519) );
  XNOR2_X1 U9457 ( .A(n9520), .B(n9521), .ZN(n9315) );
  XOR2_X1 U9458 ( .A(n9522), .B(n9523), .Z(n9520) );
  XNOR2_X1 U9459 ( .A(n9524), .B(n9525), .ZN(n9318) );
  XNOR2_X1 U9460 ( .A(n9526), .B(n9527), .ZN(n9524) );
  NOR2_X1 U9461 ( .A1(n7609), .A2(n8044), .ZN(n9527) );
  XOR2_X1 U9462 ( .A(n9528), .B(n9529), .Z(n9323) );
  XNOR2_X1 U9463 ( .A(n9530), .B(n9531), .ZN(n9529) );
  XNOR2_X1 U9464 ( .A(n9532), .B(n9533), .ZN(n9327) );
  XNOR2_X1 U9465 ( .A(n9534), .B(n9535), .ZN(n9532) );
  NOR2_X1 U9466 ( .A1(n7609), .A2(n8047), .ZN(n9535) );
  XOR2_X1 U9467 ( .A(n9536), .B(n9537), .Z(n9330) );
  XOR2_X1 U9468 ( .A(n9538), .B(n9539), .Z(n9536) );
  XNOR2_X1 U9469 ( .A(n9540), .B(n9541), .ZN(n9334) );
  XOR2_X1 U9470 ( .A(n9542), .B(n9543), .Z(n9541) );
  NAND2_X1 U9471 ( .A1(a_16_), .A2(b_25_), .ZN(n9543) );
  XNOR2_X1 U9472 ( .A(n9544), .B(n9545), .ZN(n9339) );
  XNOR2_X1 U9473 ( .A(n9546), .B(n9547), .ZN(n9545) );
  XNOR2_X1 U9474 ( .A(n9548), .B(n9549), .ZN(n9343) );
  XNOR2_X1 U9475 ( .A(n9550), .B(n9551), .ZN(n9548) );
  NOR2_X1 U9476 ( .A1(n7609), .A2(n8049), .ZN(n9551) );
  XOR2_X1 U9477 ( .A(n9552), .B(n9553), .Z(n9346) );
  XOR2_X1 U9478 ( .A(n9554), .B(n9555), .Z(n9552) );
  XOR2_X1 U9479 ( .A(n9556), .B(n9557), .Z(n9350) );
  XOR2_X1 U9480 ( .A(n9558), .B(n9559), .Z(n9556) );
  NOR2_X1 U9481 ( .A1(n7609), .A2(n8669), .ZN(n9559) );
  XOR2_X1 U9482 ( .A(n9560), .B(n9561), .Z(n9355) );
  XOR2_X1 U9483 ( .A(n9562), .B(n9563), .Z(n9561) );
  NAND2_X1 U9484 ( .A1(a_11_), .A2(b_25_), .ZN(n9563) );
  XNOR2_X1 U9485 ( .A(n9564), .B(n9565), .ZN(n9359) );
  XOR2_X1 U9486 ( .A(n9566), .B(n9567), .Z(n9564) );
  NOR2_X1 U9487 ( .A1(n7609), .A2(n8051), .ZN(n9567) );
  XOR2_X1 U9488 ( .A(n9568), .B(n9569), .Z(n9362) );
  XOR2_X1 U9489 ( .A(n9570), .B(n9571), .Z(n9568) );
  XNOR2_X1 U9490 ( .A(n9572), .B(n9573), .ZN(n9371) );
  XOR2_X1 U9491 ( .A(n9574), .B(n9575), .Z(n9572) );
  NOR2_X1 U9492 ( .A1(n7609), .A2(n7872), .ZN(n9575) );
  XNOR2_X1 U9493 ( .A(n9576), .B(n9577), .ZN(n9374) );
  XOR2_X1 U9494 ( .A(n9578), .B(n9579), .Z(n9577) );
  XOR2_X1 U9495 ( .A(n9580), .B(n9581), .Z(n9189) );
  XOR2_X1 U9496 ( .A(n9582), .B(n9583), .Z(n9580) );
  NOR2_X1 U9497 ( .A1(n7609), .A2(n7908), .ZN(n9583) );
  XNOR2_X1 U9498 ( .A(n9584), .B(n9585), .ZN(n9182) );
  XOR2_X1 U9499 ( .A(n9586), .B(n9587), .Z(n9584) );
  NOR2_X1 U9500 ( .A1(n7609), .A2(n7916), .ZN(n9587) );
  XNOR2_X1 U9501 ( .A(n9588), .B(n9589), .ZN(n9378) );
  XOR2_X1 U9502 ( .A(n9590), .B(n9591), .Z(n9589) );
  NAND2_X1 U9503 ( .A1(a_3_), .A2(b_25_), .ZN(n9591) );
  XOR2_X1 U9504 ( .A(n9592), .B(n9593), .Z(n9383) );
  XOR2_X1 U9505 ( .A(n9594), .B(n9595), .Z(n9593) );
  NAND2_X1 U9506 ( .A1(a_2_), .A2(b_25_), .ZN(n9595) );
  XNOR2_X1 U9507 ( .A(n9596), .B(n9597), .ZN(n9168) );
  XOR2_X1 U9508 ( .A(n9598), .B(n9599), .Z(n9596) );
  NOR2_X1 U9509 ( .A1(n7957), .A2(n7609), .ZN(n9599) );
  NAND2_X1 U9510 ( .A1(n9600), .A2(n9601), .ZN(n8258) );
  XNOR2_X1 U9511 ( .A(n9602), .B(n9603), .ZN(n8259) );
  XNOR2_X1 U9512 ( .A(n9604), .B(n9605), .ZN(n9603) );
  NAND2_X1 U9513 ( .A1(n9606), .A2(n9386), .ZN(n8097) );
  NOR2_X1 U9514 ( .A1(n9601), .A2(n9600), .ZN(n9386) );
  AND2_X1 U9515 ( .A1(n9607), .A2(n9608), .ZN(n9600) );
  NAND2_X1 U9516 ( .A1(n9605), .A2(n9609), .ZN(n9608) );
  OR2_X1 U9517 ( .A1(n9604), .A2(n9602), .ZN(n9609) );
  NOR2_X1 U9518 ( .A1(n8942), .A2(n7609), .ZN(n9605) );
  NAND2_X1 U9519 ( .A1(n9602), .A2(n9604), .ZN(n9607) );
  NAND2_X1 U9520 ( .A1(n9610), .A2(n9611), .ZN(n9604) );
  NAND3_X1 U9521 ( .A1(a_1_), .A2(n9612), .A3(b_25_), .ZN(n9611) );
  OR2_X1 U9522 ( .A1(n9598), .A2(n9597), .ZN(n9612) );
  NAND2_X1 U9523 ( .A1(n9597), .A2(n9598), .ZN(n9610) );
  NAND2_X1 U9524 ( .A1(n9613), .A2(n9614), .ZN(n9598) );
  NAND3_X1 U9525 ( .A1(b_25_), .A2(n9615), .A3(a_2_), .ZN(n9614) );
  OR2_X1 U9526 ( .A1(n9594), .A2(n9592), .ZN(n9615) );
  NAND2_X1 U9527 ( .A1(n9592), .A2(n9594), .ZN(n9613) );
  NAND2_X1 U9528 ( .A1(n9616), .A2(n9617), .ZN(n9594) );
  NAND3_X1 U9529 ( .A1(b_25_), .A2(n9618), .A3(a_3_), .ZN(n9617) );
  OR2_X1 U9530 ( .A1(n9590), .A2(n9588), .ZN(n9618) );
  NAND2_X1 U9531 ( .A1(n9588), .A2(n9590), .ZN(n9616) );
  NAND2_X1 U9532 ( .A1(n9619), .A2(n9620), .ZN(n9590) );
  NAND3_X1 U9533 ( .A1(b_25_), .A2(n9621), .A3(a_4_), .ZN(n9620) );
  OR2_X1 U9534 ( .A1(n9586), .A2(n9585), .ZN(n9621) );
  NAND2_X1 U9535 ( .A1(n9585), .A2(n9586), .ZN(n9619) );
  NAND2_X1 U9536 ( .A1(n9622), .A2(n9623), .ZN(n9586) );
  NAND3_X1 U9537 ( .A1(b_25_), .A2(n9624), .A3(a_5_), .ZN(n9623) );
  OR2_X1 U9538 ( .A1(n9582), .A2(n9581), .ZN(n9624) );
  NAND2_X1 U9539 ( .A1(n9581), .A2(n9582), .ZN(n9622) );
  NAND2_X1 U9540 ( .A1(n9625), .A2(n9626), .ZN(n9582) );
  NAND2_X1 U9541 ( .A1(n9578), .A2(n9627), .ZN(n9626) );
  NAND2_X1 U9542 ( .A1(n9628), .A2(n9579), .ZN(n9627) );
  INV_X1 U9543 ( .A(n9576), .ZN(n9628) );
  NAND2_X1 U9544 ( .A1(n9629), .A2(n9630), .ZN(n9578) );
  NAND3_X1 U9545 ( .A1(b_25_), .A2(n9631), .A3(a_7_), .ZN(n9630) );
  OR2_X1 U9546 ( .A1(n9574), .A2(n9573), .ZN(n9631) );
  NAND2_X1 U9547 ( .A1(n9573), .A2(n9574), .ZN(n9629) );
  NAND2_X1 U9548 ( .A1(n9632), .A2(n9633), .ZN(n9574) );
  NAND3_X1 U9549 ( .A1(b_25_), .A2(n9634), .A3(a_8_), .ZN(n9633) );
  OR2_X1 U9550 ( .A1(n9414), .A2(n9413), .ZN(n9634) );
  NAND2_X1 U9551 ( .A1(n9413), .A2(n9414), .ZN(n9632) );
  NAND2_X1 U9552 ( .A1(n9635), .A2(n9636), .ZN(n9414) );
  NAND2_X1 U9553 ( .A1(n9571), .A2(n9637), .ZN(n9636) );
  OR2_X1 U9554 ( .A1(n9570), .A2(n9569), .ZN(n9637) );
  NOR2_X1 U9555 ( .A1(n8052), .A2(n7609), .ZN(n9571) );
  NAND2_X1 U9556 ( .A1(n9569), .A2(n9570), .ZN(n9635) );
  NAND2_X1 U9557 ( .A1(n9638), .A2(n9639), .ZN(n9570) );
  NAND3_X1 U9558 ( .A1(b_25_), .A2(n9640), .A3(a_10_), .ZN(n9639) );
  OR2_X1 U9559 ( .A1(n9566), .A2(n9565), .ZN(n9640) );
  NAND2_X1 U9560 ( .A1(n9565), .A2(n9566), .ZN(n9638) );
  NAND2_X1 U9561 ( .A1(n9641), .A2(n9642), .ZN(n9566) );
  NAND3_X1 U9562 ( .A1(b_25_), .A2(n9643), .A3(a_11_), .ZN(n9642) );
  OR2_X1 U9563 ( .A1(n9562), .A2(n9560), .ZN(n9643) );
  NAND2_X1 U9564 ( .A1(n9560), .A2(n9562), .ZN(n9641) );
  NAND2_X1 U9565 ( .A1(n9644), .A2(n9645), .ZN(n9562) );
  NAND3_X1 U9566 ( .A1(b_25_), .A2(n9646), .A3(a_12_), .ZN(n9645) );
  OR2_X1 U9567 ( .A1(n9558), .A2(n9557), .ZN(n9646) );
  NAND2_X1 U9568 ( .A1(n9557), .A2(n9558), .ZN(n9644) );
  NAND2_X1 U9569 ( .A1(n9647), .A2(n9648), .ZN(n9558) );
  NAND2_X1 U9570 ( .A1(n9555), .A2(n9649), .ZN(n9648) );
  OR2_X1 U9571 ( .A1(n9554), .A2(n9553), .ZN(n9649) );
  NOR2_X1 U9572 ( .A1(n7789), .A2(n7609), .ZN(n9555) );
  NAND2_X1 U9573 ( .A1(n9553), .A2(n9554), .ZN(n9647) );
  NAND2_X1 U9574 ( .A1(n9650), .A2(n9651), .ZN(n9554) );
  NAND3_X1 U9575 ( .A1(b_25_), .A2(n9652), .A3(a_14_), .ZN(n9651) );
  NAND2_X1 U9576 ( .A1(n9550), .A2(n9549), .ZN(n9652) );
  OR2_X1 U9577 ( .A1(n9549), .A2(n9550), .ZN(n9650) );
  AND2_X1 U9578 ( .A1(n9653), .A2(n9654), .ZN(n9550) );
  NAND2_X1 U9579 ( .A1(n9547), .A2(n9655), .ZN(n9654) );
  OR2_X1 U9580 ( .A1(n9546), .A2(n9544), .ZN(n9655) );
  NOR2_X1 U9581 ( .A1(n7754), .A2(n7609), .ZN(n9547) );
  NAND2_X1 U9582 ( .A1(n9544), .A2(n9546), .ZN(n9653) );
  NAND2_X1 U9583 ( .A1(n9656), .A2(n9657), .ZN(n9546) );
  NAND3_X1 U9584 ( .A1(b_25_), .A2(n9658), .A3(a_16_), .ZN(n9657) );
  OR2_X1 U9585 ( .A1(n9542), .A2(n9540), .ZN(n9658) );
  NAND2_X1 U9586 ( .A1(n9540), .A2(n9542), .ZN(n9656) );
  NAND2_X1 U9587 ( .A1(n9659), .A2(n9660), .ZN(n9542) );
  NAND2_X1 U9588 ( .A1(n9539), .A2(n9661), .ZN(n9660) );
  OR2_X1 U9589 ( .A1(n9538), .A2(n9537), .ZN(n9661) );
  NOR2_X1 U9590 ( .A1(n7732), .A2(n7609), .ZN(n9539) );
  NAND2_X1 U9591 ( .A1(n9537), .A2(n9538), .ZN(n9659) );
  NAND2_X1 U9592 ( .A1(n9662), .A2(n9663), .ZN(n9538) );
  NAND3_X1 U9593 ( .A1(b_25_), .A2(n9664), .A3(a_18_), .ZN(n9663) );
  NAND2_X1 U9594 ( .A1(n9534), .A2(n9533), .ZN(n9664) );
  OR2_X1 U9595 ( .A1(n9533), .A2(n9534), .ZN(n9662) );
  AND2_X1 U9596 ( .A1(n9665), .A2(n9666), .ZN(n9534) );
  NAND2_X1 U9597 ( .A1(n9531), .A2(n9667), .ZN(n9666) );
  OR2_X1 U9598 ( .A1(n9530), .A2(n9528), .ZN(n9667) );
  NOR2_X1 U9599 ( .A1(n8045), .A2(n7609), .ZN(n9531) );
  NAND2_X1 U9600 ( .A1(n9528), .A2(n9530), .ZN(n9665) );
  NAND2_X1 U9601 ( .A1(n9668), .A2(n9669), .ZN(n9530) );
  NAND3_X1 U9602 ( .A1(b_25_), .A2(n9670), .A3(a_20_), .ZN(n9669) );
  NAND2_X1 U9603 ( .A1(n9526), .A2(n9525), .ZN(n9670) );
  OR2_X1 U9604 ( .A1(n9525), .A2(n9526), .ZN(n9668) );
  AND2_X1 U9605 ( .A1(n9671), .A2(n9672), .ZN(n9526) );
  NAND2_X1 U9606 ( .A1(n9523), .A2(n9673), .ZN(n9672) );
  OR2_X1 U9607 ( .A1(n9522), .A2(n9521), .ZN(n9673) );
  NOR2_X1 U9608 ( .A1(n7665), .A2(n7609), .ZN(n9523) );
  NAND2_X1 U9609 ( .A1(n9521), .A2(n9522), .ZN(n9671) );
  NAND2_X1 U9610 ( .A1(n9674), .A2(n9675), .ZN(n9522) );
  NAND3_X1 U9611 ( .A1(b_25_), .A2(n9676), .A3(a_22_), .ZN(n9675) );
  OR2_X1 U9612 ( .A1(n9518), .A2(n9516), .ZN(n9676) );
  NAND2_X1 U9613 ( .A1(n9516), .A2(n9518), .ZN(n9674) );
  NAND2_X1 U9614 ( .A1(n9677), .A2(n9678), .ZN(n9518) );
  NAND2_X1 U9615 ( .A1(n9515), .A2(n9679), .ZN(n9678) );
  OR2_X1 U9616 ( .A1(n9514), .A2(n9512), .ZN(n9679) );
  NOR2_X1 U9617 ( .A1(n8042), .A2(n7609), .ZN(n9515) );
  NAND2_X1 U9618 ( .A1(n9512), .A2(n9514), .ZN(n9677) );
  NAND2_X1 U9619 ( .A1(n9680), .A2(n9681), .ZN(n9514) );
  NAND3_X1 U9620 ( .A1(b_25_), .A2(n9682), .A3(a_24_), .ZN(n9681) );
  NAND2_X1 U9621 ( .A1(n9510), .A2(n9509), .ZN(n9682) );
  OR2_X1 U9622 ( .A1(n9509), .A2(n9510), .ZN(n9680) );
  AND2_X1 U9623 ( .A1(n9683), .A2(n9684), .ZN(n9510) );
  NAND2_X1 U9624 ( .A1(n7607), .A2(n9685), .ZN(n9684) );
  OR2_X1 U9625 ( .A1(n9507), .A2(n9506), .ZN(n9685) );
  INV_X1 U9626 ( .A(n8022), .ZN(n7607) );
  NAND2_X1 U9627 ( .A1(a_25_), .A2(b_25_), .ZN(n8022) );
  NAND2_X1 U9628 ( .A1(n9506), .A2(n9507), .ZN(n9683) );
  NAND2_X1 U9629 ( .A1(n9503), .A2(n9686), .ZN(n9507) );
  NAND2_X1 U9630 ( .A1(n9502), .A2(n9504), .ZN(n9686) );
  NAND2_X1 U9631 ( .A1(n9687), .A2(n9688), .ZN(n9504) );
  NAND2_X1 U9632 ( .A1(b_25_), .A2(a_26_), .ZN(n9688) );
  INV_X1 U9633 ( .A(n9689), .ZN(n9687) );
  XNOR2_X1 U9634 ( .A(n9690), .B(n9691), .ZN(n9502) );
  NAND2_X1 U9635 ( .A1(n9692), .A2(n9693), .ZN(n9690) );
  NAND2_X1 U9636 ( .A1(a_26_), .A2(n9689), .ZN(n9503) );
  NAND2_X1 U9637 ( .A1(n9475), .A2(n9694), .ZN(n9689) );
  NAND2_X1 U9638 ( .A1(n9474), .A2(n9476), .ZN(n9694) );
  NAND2_X1 U9639 ( .A1(n9695), .A2(n9696), .ZN(n9476) );
  NAND2_X1 U9640 ( .A1(b_25_), .A2(a_27_), .ZN(n9696) );
  INV_X1 U9641 ( .A(n9697), .ZN(n9695) );
  XNOR2_X1 U9642 ( .A(n9698), .B(n9699), .ZN(n9474) );
  XOR2_X1 U9643 ( .A(n9700), .B(n9701), .Z(n9698) );
  NAND2_X1 U9644 ( .A1(b_24_), .A2(a_28_), .ZN(n9700) );
  NAND2_X1 U9645 ( .A1(a_27_), .A2(n9697), .ZN(n9475) );
  NAND2_X1 U9646 ( .A1(n9702), .A2(n9703), .ZN(n9697) );
  NAND3_X1 U9647 ( .A1(a_28_), .A2(n9704), .A3(b_25_), .ZN(n9703) );
  NAND2_X1 U9648 ( .A1(n9484), .A2(n9482), .ZN(n9704) );
  OR2_X1 U9649 ( .A1(n9482), .A2(n9484), .ZN(n9702) );
  AND2_X1 U9650 ( .A1(n9705), .A2(n9706), .ZN(n9484) );
  NAND2_X1 U9651 ( .A1(n9498), .A2(n9707), .ZN(n9706) );
  OR2_X1 U9652 ( .A1(n9499), .A2(n9500), .ZN(n9707) );
  NOR2_X1 U9653 ( .A1(n7609), .A2(n7545), .ZN(n9498) );
  NAND2_X1 U9654 ( .A1(n9500), .A2(n9499), .ZN(n9705) );
  NAND2_X1 U9655 ( .A1(n9708), .A2(n9709), .ZN(n9499) );
  NAND2_X1 U9656 ( .A1(b_23_), .A2(n9710), .ZN(n9709) );
  NAND2_X1 U9657 ( .A1(n7527), .A2(n9711), .ZN(n9710) );
  NAND2_X1 U9658 ( .A1(a_31_), .A2(n8040), .ZN(n9711) );
  NAND2_X1 U9659 ( .A1(b_24_), .A2(n9712), .ZN(n9708) );
  NAND2_X1 U9660 ( .A1(n7531), .A2(n9713), .ZN(n9712) );
  NAND2_X1 U9661 ( .A1(a_30_), .A2(n7636), .ZN(n9713) );
  AND3_X1 U9662 ( .A1(b_24_), .A2(b_25_), .A3(n7494), .ZN(n9500) );
  XNOR2_X1 U9663 ( .A(n9714), .B(n9715), .ZN(n9482) );
  XOR2_X1 U9664 ( .A(n9716), .B(n9717), .Z(n9714) );
  XNOR2_X1 U9665 ( .A(n9718), .B(n9719), .ZN(n9506) );
  NAND2_X1 U9666 ( .A1(n9720), .A2(n9721), .ZN(n9718) );
  XNOR2_X1 U9667 ( .A(n9722), .B(n9723), .ZN(n9509) );
  XOR2_X1 U9668 ( .A(n9724), .B(n9725), .Z(n9722) );
  XOR2_X1 U9669 ( .A(n9726), .B(n9727), .Z(n9512) );
  XOR2_X1 U9670 ( .A(n9728), .B(n9729), .Z(n9726) );
  XOR2_X1 U9671 ( .A(n9730), .B(n9731), .Z(n9516) );
  XOR2_X1 U9672 ( .A(n9732), .B(n9733), .Z(n9730) );
  XNOR2_X1 U9673 ( .A(n9734), .B(n9735), .ZN(n9521) );
  XOR2_X1 U9674 ( .A(n9736), .B(n9737), .Z(n9735) );
  NAND2_X1 U9675 ( .A1(a_22_), .A2(b_24_), .ZN(n9737) );
  XNOR2_X1 U9676 ( .A(n9738), .B(n9739), .ZN(n9525) );
  XOR2_X1 U9677 ( .A(n9740), .B(n9741), .Z(n9738) );
  XNOR2_X1 U9678 ( .A(n9742), .B(n9743), .ZN(n9528) );
  XNOR2_X1 U9679 ( .A(n9744), .B(n9745), .ZN(n9742) );
  NOR2_X1 U9680 ( .A1(n8040), .A2(n8044), .ZN(n9745) );
  XOR2_X1 U9681 ( .A(n9746), .B(n9747), .Z(n9533) );
  XNOR2_X1 U9682 ( .A(n9748), .B(n9749), .ZN(n9747) );
  XNOR2_X1 U9683 ( .A(n9750), .B(n9751), .ZN(n9537) );
  XNOR2_X1 U9684 ( .A(n9752), .B(n9753), .ZN(n9750) );
  NOR2_X1 U9685 ( .A1(n8040), .A2(n8047), .ZN(n9753) );
  XOR2_X1 U9686 ( .A(n9754), .B(n9755), .Z(n9540) );
  XOR2_X1 U9687 ( .A(n9756), .B(n9757), .Z(n9754) );
  XOR2_X1 U9688 ( .A(n9758), .B(n9759), .Z(n9544) );
  XOR2_X1 U9689 ( .A(n9760), .B(n9761), .Z(n9758) );
  NOR2_X1 U9690 ( .A1(n8040), .A2(n8438), .ZN(n9761) );
  XOR2_X1 U9691 ( .A(n9762), .B(n9763), .Z(n9549) );
  XNOR2_X1 U9692 ( .A(n9764), .B(n9765), .ZN(n9763) );
  XNOR2_X1 U9693 ( .A(n9766), .B(n9767), .ZN(n9553) );
  XOR2_X1 U9694 ( .A(n9768), .B(n9769), .Z(n9766) );
  NAND2_X1 U9695 ( .A1(a_14_), .A2(b_24_), .ZN(n9768) );
  XNOR2_X1 U9696 ( .A(n9770), .B(n9771), .ZN(n9557) );
  XNOR2_X1 U9697 ( .A(n9772), .B(n9773), .ZN(n9770) );
  XNOR2_X1 U9698 ( .A(n9774), .B(n9775), .ZN(n9560) );
  XOR2_X1 U9699 ( .A(n9776), .B(n9777), .Z(n9775) );
  NAND2_X1 U9700 ( .A1(a_12_), .A2(b_24_), .ZN(n9777) );
  XNOR2_X1 U9701 ( .A(n9778), .B(n9779), .ZN(n9565) );
  NAND2_X1 U9702 ( .A1(n9780), .A2(n9781), .ZN(n9778) );
  XNOR2_X1 U9703 ( .A(n9782), .B(n9783), .ZN(n9569) );
  XNOR2_X1 U9704 ( .A(n9784), .B(n9785), .ZN(n9783) );
  NOR2_X1 U9705 ( .A1(n8040), .A2(n8051), .ZN(n9785) );
  XNOR2_X1 U9706 ( .A(n9786), .B(n9787), .ZN(n9413) );
  XNOR2_X1 U9707 ( .A(n9788), .B(n9789), .ZN(n9787) );
  XNOR2_X1 U9708 ( .A(n9790), .B(n9791), .ZN(n9573) );
  XOR2_X1 U9709 ( .A(n9792), .B(n9793), .Z(n9790) );
  NAND2_X1 U9710 ( .A1(a_8_), .A2(b_24_), .ZN(n9792) );
  NAND2_X1 U9711 ( .A1(n9794), .A2(n9576), .ZN(n9625) );
  XNOR2_X1 U9712 ( .A(n9795), .B(n9796), .ZN(n9576) );
  NAND2_X1 U9713 ( .A1(n9797), .A2(n9798), .ZN(n9795) );
  INV_X1 U9714 ( .A(n9579), .ZN(n9794) );
  NAND2_X1 U9715 ( .A1(a_6_), .A2(b_25_), .ZN(n9579) );
  XNOR2_X1 U9716 ( .A(n9799), .B(n9800), .ZN(n9581) );
  XNOR2_X1 U9717 ( .A(n9801), .B(n9802), .ZN(n9799) );
  XNOR2_X1 U9718 ( .A(n9803), .B(n9804), .ZN(n9585) );
  XNOR2_X1 U9719 ( .A(n9805), .B(n9806), .ZN(n9804) );
  XNOR2_X1 U9720 ( .A(n9807), .B(n9808), .ZN(n9588) );
  XOR2_X1 U9721 ( .A(n9809), .B(n9810), .Z(n9807) );
  NAND2_X1 U9722 ( .A1(a_4_), .A2(b_24_), .ZN(n9809) );
  XNOR2_X1 U9723 ( .A(n9811), .B(n9812), .ZN(n9592) );
  NAND2_X1 U9724 ( .A1(n9813), .A2(n9814), .ZN(n9811) );
  XNOR2_X1 U9725 ( .A(n9815), .B(n9816), .ZN(n9597) );
  NAND2_X1 U9726 ( .A1(n9817), .A2(n9818), .ZN(n9815) );
  XNOR2_X1 U9727 ( .A(n9819), .B(n9820), .ZN(n9602) );
  NAND2_X1 U9728 ( .A1(n9821), .A2(n9822), .ZN(n9819) );
  XOR2_X1 U9729 ( .A(n9823), .B(n9824), .Z(n9601) );
  NAND2_X1 U9730 ( .A1(n9825), .A2(n9826), .ZN(n9823) );
  XOR2_X1 U9731 ( .A(n8249), .B(n8250), .Z(n9606) );
  NAND3_X1 U9732 ( .A1(n8249), .A2(n8250), .A3(n9827), .ZN(n8101) );
  XOR2_X1 U9733 ( .A(n8245), .B(n8244), .Z(n9827) );
  NAND2_X1 U9734 ( .A1(n9825), .A2(n9828), .ZN(n8250) );
  NAND2_X1 U9735 ( .A1(n9824), .A2(n9826), .ZN(n9828) );
  NAND2_X1 U9736 ( .A1(n9829), .A2(n9830), .ZN(n9826) );
  NAND2_X1 U9737 ( .A1(a_0_), .A2(b_24_), .ZN(n9830) );
  INV_X1 U9738 ( .A(n9831), .ZN(n9829) );
  XNOR2_X1 U9739 ( .A(n9832), .B(n9833), .ZN(n9824) );
  XOR2_X1 U9740 ( .A(n9834), .B(n9835), .Z(n9833) );
  NAND2_X1 U9741 ( .A1(b_23_), .A2(a_1_), .ZN(n9835) );
  NAND2_X1 U9742 ( .A1(a_0_), .A2(n9831), .ZN(n9825) );
  NAND2_X1 U9743 ( .A1(n9821), .A2(n9836), .ZN(n9831) );
  NAND2_X1 U9744 ( .A1(n9820), .A2(n9822), .ZN(n9836) );
  NAND2_X1 U9745 ( .A1(n9837), .A2(n9838), .ZN(n9822) );
  NAND2_X1 U9746 ( .A1(b_24_), .A2(a_1_), .ZN(n9838) );
  INV_X1 U9747 ( .A(n9839), .ZN(n9837) );
  XNOR2_X1 U9748 ( .A(n9840), .B(n9841), .ZN(n9820) );
  XNOR2_X1 U9749 ( .A(n9842), .B(n9843), .ZN(n9840) );
  NOR2_X1 U9750 ( .A1(n7636), .A2(n8056), .ZN(n9843) );
  NAND2_X1 U9751 ( .A1(a_1_), .A2(n9839), .ZN(n9821) );
  NAND2_X1 U9752 ( .A1(n9817), .A2(n9844), .ZN(n9839) );
  NAND2_X1 U9753 ( .A1(n9816), .A2(n9818), .ZN(n9844) );
  NAND2_X1 U9754 ( .A1(n9845), .A2(n9846), .ZN(n9818) );
  NAND2_X1 U9755 ( .A1(a_2_), .A2(b_24_), .ZN(n9846) );
  INV_X1 U9756 ( .A(n9847), .ZN(n9845) );
  XNOR2_X1 U9757 ( .A(n9848), .B(n9849), .ZN(n9816) );
  XOR2_X1 U9758 ( .A(n9850), .B(n9851), .Z(n9849) );
  NAND2_X1 U9759 ( .A1(a_3_), .A2(b_23_), .ZN(n9851) );
  NAND2_X1 U9760 ( .A1(a_2_), .A2(n9847), .ZN(n9817) );
  NAND2_X1 U9761 ( .A1(n9813), .A2(n9852), .ZN(n9847) );
  NAND2_X1 U9762 ( .A1(n9812), .A2(n9814), .ZN(n9852) );
  NAND2_X1 U9763 ( .A1(n9853), .A2(n9854), .ZN(n9814) );
  NAND2_X1 U9764 ( .A1(a_3_), .A2(b_24_), .ZN(n9854) );
  INV_X1 U9765 ( .A(n9855), .ZN(n9853) );
  XNOR2_X1 U9766 ( .A(n9856), .B(n9857), .ZN(n9812) );
  XOR2_X1 U9767 ( .A(n9858), .B(n9859), .Z(n9857) );
  NAND2_X1 U9768 ( .A1(a_4_), .A2(b_23_), .ZN(n9859) );
  NAND2_X1 U9769 ( .A1(a_3_), .A2(n9855), .ZN(n9813) );
  NAND2_X1 U9770 ( .A1(n9860), .A2(n9861), .ZN(n9855) );
  NAND3_X1 U9771 ( .A1(b_24_), .A2(n9862), .A3(a_4_), .ZN(n9861) );
  NAND2_X1 U9772 ( .A1(n9810), .A2(n9808), .ZN(n9862) );
  OR2_X1 U9773 ( .A1(n9808), .A2(n9810), .ZN(n9860) );
  AND2_X1 U9774 ( .A1(n9863), .A2(n9864), .ZN(n9810) );
  NAND2_X1 U9775 ( .A1(n9806), .A2(n9865), .ZN(n9864) );
  OR2_X1 U9776 ( .A1(n9805), .A2(n9803), .ZN(n9865) );
  NOR2_X1 U9777 ( .A1(n7908), .A2(n8040), .ZN(n9806) );
  NAND2_X1 U9778 ( .A1(n9803), .A2(n9805), .ZN(n9863) );
  NAND2_X1 U9779 ( .A1(n9866), .A2(n9867), .ZN(n9805) );
  NAND2_X1 U9780 ( .A1(n9802), .A2(n9868), .ZN(n9867) );
  NAND2_X1 U9781 ( .A1(n9800), .A2(n9801), .ZN(n9868) );
  NAND2_X1 U9782 ( .A1(n9797), .A2(n9869), .ZN(n9802) );
  NAND2_X1 U9783 ( .A1(n9796), .A2(n9798), .ZN(n9869) );
  NAND2_X1 U9784 ( .A1(n9870), .A2(n9871), .ZN(n9798) );
  NAND2_X1 U9785 ( .A1(a_7_), .A2(b_24_), .ZN(n9871) );
  INV_X1 U9786 ( .A(n9872), .ZN(n9870) );
  XNOR2_X1 U9787 ( .A(n9873), .B(n9874), .ZN(n9796) );
  XNOR2_X1 U9788 ( .A(n9875), .B(n9876), .ZN(n9874) );
  NAND2_X1 U9789 ( .A1(a_7_), .A2(n9872), .ZN(n9797) );
  NAND2_X1 U9790 ( .A1(n9877), .A2(n9878), .ZN(n9872) );
  NAND3_X1 U9791 ( .A1(b_24_), .A2(n9879), .A3(a_8_), .ZN(n9878) );
  NAND2_X1 U9792 ( .A1(n9793), .A2(n9791), .ZN(n9879) );
  OR2_X1 U9793 ( .A1(n9791), .A2(n9793), .ZN(n9877) );
  AND2_X1 U9794 ( .A1(n9880), .A2(n9881), .ZN(n9793) );
  NAND2_X1 U9795 ( .A1(n9789), .A2(n9882), .ZN(n9881) );
  OR2_X1 U9796 ( .A1(n9788), .A2(n9786), .ZN(n9882) );
  NOR2_X1 U9797 ( .A1(n8052), .A2(n8040), .ZN(n9789) );
  NAND2_X1 U9798 ( .A1(n9786), .A2(n9788), .ZN(n9880) );
  NAND2_X1 U9799 ( .A1(n9883), .A2(n9884), .ZN(n9788) );
  NAND3_X1 U9800 ( .A1(b_24_), .A2(n9885), .A3(a_10_), .ZN(n9884) );
  OR2_X1 U9801 ( .A1(n9784), .A2(n9782), .ZN(n9885) );
  NAND2_X1 U9802 ( .A1(n9782), .A2(n9784), .ZN(n9883) );
  NAND2_X1 U9803 ( .A1(n9780), .A2(n9886), .ZN(n9784) );
  NAND2_X1 U9804 ( .A1(n9779), .A2(n9781), .ZN(n9886) );
  NAND2_X1 U9805 ( .A1(n9887), .A2(n9888), .ZN(n9781) );
  NAND2_X1 U9806 ( .A1(a_11_), .A2(b_24_), .ZN(n9888) );
  INV_X1 U9807 ( .A(n9889), .ZN(n9887) );
  XNOR2_X1 U9808 ( .A(n9890), .B(n9891), .ZN(n9779) );
  XNOR2_X1 U9809 ( .A(n9892), .B(n9893), .ZN(n9890) );
  NOR2_X1 U9810 ( .A1(n7636), .A2(n8669), .ZN(n9893) );
  NAND2_X1 U9811 ( .A1(a_11_), .A2(n9889), .ZN(n9780) );
  NAND2_X1 U9812 ( .A1(n9894), .A2(n9895), .ZN(n9889) );
  NAND3_X1 U9813 ( .A1(b_24_), .A2(n9896), .A3(a_12_), .ZN(n9895) );
  OR2_X1 U9814 ( .A1(n9776), .A2(n9774), .ZN(n9896) );
  NAND2_X1 U9815 ( .A1(n9774), .A2(n9776), .ZN(n9894) );
  NAND2_X1 U9816 ( .A1(n9897), .A2(n9898), .ZN(n9776) );
  NAND2_X1 U9817 ( .A1(n9773), .A2(n9899), .ZN(n9898) );
  NAND2_X1 U9818 ( .A1(n9772), .A2(n9771), .ZN(n9899) );
  NOR2_X1 U9819 ( .A1(n7789), .A2(n8040), .ZN(n9773) );
  OR2_X1 U9820 ( .A1(n9771), .A2(n9772), .ZN(n9897) );
  AND2_X1 U9821 ( .A1(n9900), .A2(n9901), .ZN(n9772) );
  NAND3_X1 U9822 ( .A1(b_24_), .A2(n9902), .A3(a_14_), .ZN(n9901) );
  NAND2_X1 U9823 ( .A1(n9769), .A2(n9767), .ZN(n9902) );
  OR2_X1 U9824 ( .A1(n9767), .A2(n9769), .ZN(n9900) );
  AND2_X1 U9825 ( .A1(n9903), .A2(n9904), .ZN(n9769) );
  NAND2_X1 U9826 ( .A1(n9765), .A2(n9905), .ZN(n9904) );
  OR2_X1 U9827 ( .A1(n9764), .A2(n9762), .ZN(n9905) );
  NOR2_X1 U9828 ( .A1(n7754), .A2(n8040), .ZN(n9765) );
  NAND2_X1 U9829 ( .A1(n9762), .A2(n9764), .ZN(n9903) );
  NAND2_X1 U9830 ( .A1(n9906), .A2(n9907), .ZN(n9764) );
  NAND3_X1 U9831 ( .A1(b_24_), .A2(n9908), .A3(a_16_), .ZN(n9907) );
  OR2_X1 U9832 ( .A1(n9760), .A2(n9759), .ZN(n9908) );
  NAND2_X1 U9833 ( .A1(n9759), .A2(n9760), .ZN(n9906) );
  NAND2_X1 U9834 ( .A1(n9909), .A2(n9910), .ZN(n9760) );
  NAND2_X1 U9835 ( .A1(n9757), .A2(n9911), .ZN(n9910) );
  OR2_X1 U9836 ( .A1(n9756), .A2(n9755), .ZN(n9911) );
  NOR2_X1 U9837 ( .A1(n7732), .A2(n8040), .ZN(n9757) );
  NAND2_X1 U9838 ( .A1(n9755), .A2(n9756), .ZN(n9909) );
  NAND2_X1 U9839 ( .A1(n9912), .A2(n9913), .ZN(n9756) );
  NAND3_X1 U9840 ( .A1(b_24_), .A2(n9914), .A3(a_18_), .ZN(n9913) );
  NAND2_X1 U9841 ( .A1(n9752), .A2(n9751), .ZN(n9914) );
  OR2_X1 U9842 ( .A1(n9751), .A2(n9752), .ZN(n9912) );
  AND2_X1 U9843 ( .A1(n9915), .A2(n9916), .ZN(n9752) );
  NAND2_X1 U9844 ( .A1(n9749), .A2(n9917), .ZN(n9916) );
  OR2_X1 U9845 ( .A1(n9748), .A2(n9746), .ZN(n9917) );
  NOR2_X1 U9846 ( .A1(n8045), .A2(n8040), .ZN(n9749) );
  NAND2_X1 U9847 ( .A1(n9746), .A2(n9748), .ZN(n9915) );
  NAND2_X1 U9848 ( .A1(n9918), .A2(n9919), .ZN(n9748) );
  NAND3_X1 U9849 ( .A1(b_24_), .A2(n9920), .A3(a_20_), .ZN(n9919) );
  NAND2_X1 U9850 ( .A1(n9744), .A2(n9743), .ZN(n9920) );
  OR2_X1 U9851 ( .A1(n9743), .A2(n9744), .ZN(n9918) );
  AND2_X1 U9852 ( .A1(n9921), .A2(n9922), .ZN(n9744) );
  NAND2_X1 U9853 ( .A1(n9741), .A2(n9923), .ZN(n9922) );
  OR2_X1 U9854 ( .A1(n9740), .A2(n9739), .ZN(n9923) );
  NOR2_X1 U9855 ( .A1(n7665), .A2(n8040), .ZN(n9741) );
  NAND2_X1 U9856 ( .A1(n9739), .A2(n9740), .ZN(n9921) );
  NAND2_X1 U9857 ( .A1(n9924), .A2(n9925), .ZN(n9740) );
  NAND3_X1 U9858 ( .A1(b_24_), .A2(n9926), .A3(a_22_), .ZN(n9925) );
  OR2_X1 U9859 ( .A1(n9736), .A2(n9734), .ZN(n9926) );
  NAND2_X1 U9860 ( .A1(n9734), .A2(n9736), .ZN(n9924) );
  NAND2_X1 U9861 ( .A1(n9927), .A2(n9928), .ZN(n9736) );
  NAND2_X1 U9862 ( .A1(n9733), .A2(n9929), .ZN(n9928) );
  OR2_X1 U9863 ( .A1(n9732), .A2(n9731), .ZN(n9929) );
  NOR2_X1 U9864 ( .A1(n8042), .A2(n8040), .ZN(n9733) );
  NAND2_X1 U9865 ( .A1(n9731), .A2(n9732), .ZN(n9927) );
  NAND2_X1 U9866 ( .A1(n9930), .A2(n9931), .ZN(n9732) );
  NAND2_X1 U9867 ( .A1(n9727), .A2(n9932), .ZN(n9931) );
  OR2_X1 U9868 ( .A1(n9728), .A2(n9729), .ZN(n9932) );
  XOR2_X1 U9869 ( .A(n9933), .B(n9934), .Z(n9727) );
  XOR2_X1 U9870 ( .A(n9935), .B(n9936), .Z(n9933) );
  NAND2_X1 U9871 ( .A1(n9729), .A2(n9728), .ZN(n9930) );
  NAND2_X1 U9872 ( .A1(n9937), .A2(n9938), .ZN(n9728) );
  NAND2_X1 U9873 ( .A1(n9725), .A2(n9939), .ZN(n9938) );
  OR2_X1 U9874 ( .A1(n9724), .A2(n9723), .ZN(n9939) );
  NOR2_X1 U9875 ( .A1(n8040), .A2(n8039), .ZN(n9725) );
  NAND2_X1 U9876 ( .A1(n9723), .A2(n9724), .ZN(n9937) );
  NAND2_X1 U9877 ( .A1(n9720), .A2(n9940), .ZN(n9724) );
  NAND2_X1 U9878 ( .A1(n9719), .A2(n9721), .ZN(n9940) );
  NAND2_X1 U9879 ( .A1(n9941), .A2(n9942), .ZN(n9721) );
  NAND2_X1 U9880 ( .A1(b_24_), .A2(a_26_), .ZN(n9942) );
  INV_X1 U9881 ( .A(n9943), .ZN(n9941) );
  XNOR2_X1 U9882 ( .A(n9944), .B(n9945), .ZN(n9719) );
  NAND2_X1 U9883 ( .A1(n9946), .A2(n9947), .ZN(n9944) );
  NAND2_X1 U9884 ( .A1(a_26_), .A2(n9943), .ZN(n9720) );
  NAND2_X1 U9885 ( .A1(n9692), .A2(n9948), .ZN(n9943) );
  NAND2_X1 U9886 ( .A1(n9691), .A2(n9693), .ZN(n9948) );
  NAND2_X1 U9887 ( .A1(n9949), .A2(n9950), .ZN(n9693) );
  NAND2_X1 U9888 ( .A1(b_24_), .A2(a_27_), .ZN(n9950) );
  INV_X1 U9889 ( .A(n9951), .ZN(n9949) );
  XNOR2_X1 U9890 ( .A(n9952), .B(n9953), .ZN(n9691) );
  XOR2_X1 U9891 ( .A(n9954), .B(n9955), .Z(n9952) );
  NAND2_X1 U9892 ( .A1(b_23_), .A2(a_28_), .ZN(n9954) );
  NAND2_X1 U9893 ( .A1(a_27_), .A2(n9951), .ZN(n9692) );
  NAND2_X1 U9894 ( .A1(n9956), .A2(n9957), .ZN(n9951) );
  NAND3_X1 U9895 ( .A1(a_28_), .A2(n9958), .A3(b_24_), .ZN(n9957) );
  NAND2_X1 U9896 ( .A1(n9701), .A2(n9699), .ZN(n9958) );
  OR2_X1 U9897 ( .A1(n9699), .A2(n9701), .ZN(n9956) );
  AND2_X1 U9898 ( .A1(n9959), .A2(n9960), .ZN(n9701) );
  NAND2_X1 U9899 ( .A1(n9715), .A2(n9961), .ZN(n9960) );
  OR2_X1 U9900 ( .A1(n9716), .A2(n9717), .ZN(n9961) );
  NOR2_X1 U9901 ( .A1(n8040), .A2(n7545), .ZN(n9715) );
  NAND2_X1 U9902 ( .A1(n9717), .A2(n9716), .ZN(n9959) );
  NAND2_X1 U9903 ( .A1(n9962), .A2(n9963), .ZN(n9716) );
  NAND2_X1 U9904 ( .A1(b_22_), .A2(n9964), .ZN(n9963) );
  NAND2_X1 U9905 ( .A1(n7527), .A2(n9965), .ZN(n9964) );
  NAND2_X1 U9906 ( .A1(a_31_), .A2(n7636), .ZN(n9965) );
  NAND2_X1 U9907 ( .A1(b_23_), .A2(n9966), .ZN(n9962) );
  NAND2_X1 U9908 ( .A1(n7531), .A2(n9967), .ZN(n9966) );
  NAND2_X1 U9909 ( .A1(a_30_), .A2(n9968), .ZN(n9967) );
  AND3_X1 U9910 ( .A1(b_24_), .A2(b_23_), .A3(n7494), .ZN(n9717) );
  XNOR2_X1 U9911 ( .A(n9969), .B(n9970), .ZN(n9699) );
  XOR2_X1 U9912 ( .A(n9971), .B(n9972), .Z(n9969) );
  XNOR2_X1 U9913 ( .A(n9973), .B(n9974), .ZN(n9723) );
  NAND2_X1 U9914 ( .A1(n9975), .A2(n9976), .ZN(n9973) );
  INV_X1 U9915 ( .A(n7627), .ZN(n9729) );
  NAND2_X1 U9916 ( .A1(b_24_), .A2(a_24_), .ZN(n7627) );
  XNOR2_X1 U9917 ( .A(n9977), .B(n9978), .ZN(n9731) );
  XNOR2_X1 U9918 ( .A(n9979), .B(n9980), .ZN(n9977) );
  NOR2_X1 U9919 ( .A1(n8041), .A2(n7636), .ZN(n9980) );
  XNOR2_X1 U9920 ( .A(n9981), .B(n9982), .ZN(n9734) );
  XNOR2_X1 U9921 ( .A(n9983), .B(n7634), .ZN(n9982) );
  XNOR2_X1 U9922 ( .A(n9984), .B(n9985), .ZN(n9739) );
  XOR2_X1 U9923 ( .A(n9986), .B(n9987), .Z(n9985) );
  NAND2_X1 U9924 ( .A1(a_22_), .A2(b_23_), .ZN(n9987) );
  XNOR2_X1 U9925 ( .A(n9988), .B(n9989), .ZN(n9743) );
  XOR2_X1 U9926 ( .A(n9990), .B(n9991), .Z(n9988) );
  XNOR2_X1 U9927 ( .A(n9992), .B(n9993), .ZN(n9746) );
  XNOR2_X1 U9928 ( .A(n9994), .B(n9995), .ZN(n9992) );
  NOR2_X1 U9929 ( .A1(n7636), .A2(n8044), .ZN(n9995) );
  XOR2_X1 U9930 ( .A(n9996), .B(n9997), .Z(n9751) );
  XNOR2_X1 U9931 ( .A(n9998), .B(n9999), .ZN(n9997) );
  XNOR2_X1 U9932 ( .A(n10000), .B(n10001), .ZN(n9755) );
  XNOR2_X1 U9933 ( .A(n10002), .B(n10003), .ZN(n10000) );
  NOR2_X1 U9934 ( .A1(n7636), .A2(n8047), .ZN(n10003) );
  XNOR2_X1 U9935 ( .A(n10004), .B(n10005), .ZN(n9759) );
  XNOR2_X1 U9936 ( .A(n10006), .B(n10007), .ZN(n10004) );
  XNOR2_X1 U9937 ( .A(n10008), .B(n10009), .ZN(n9762) );
  XOR2_X1 U9938 ( .A(n10010), .B(n10011), .Z(n10009) );
  NAND2_X1 U9939 ( .A1(a_16_), .A2(b_23_), .ZN(n10011) );
  XOR2_X1 U9940 ( .A(n10012), .B(n10013), .Z(n9767) );
  XOR2_X1 U9941 ( .A(n10014), .B(n10015), .Z(n10013) );
  NAND2_X1 U9942 ( .A1(a_15_), .A2(b_23_), .ZN(n10015) );
  XOR2_X1 U9943 ( .A(n10016), .B(n10017), .Z(n9771) );
  NAND2_X1 U9944 ( .A1(n10018), .A2(n10019), .ZN(n10016) );
  XOR2_X1 U9945 ( .A(n10020), .B(n10021), .Z(n9774) );
  XOR2_X1 U9946 ( .A(n10022), .B(n10023), .Z(n10020) );
  XOR2_X1 U9947 ( .A(n10024), .B(n10025), .Z(n9782) );
  XOR2_X1 U9948 ( .A(n10026), .B(n10027), .Z(n10024) );
  NOR2_X1 U9949 ( .A1(n7636), .A2(n7811), .ZN(n10027) );
  XNOR2_X1 U9950 ( .A(n10028), .B(n10029), .ZN(n9786) );
  NAND2_X1 U9951 ( .A1(n10030), .A2(n10031), .ZN(n10028) );
  XOR2_X1 U9952 ( .A(n10032), .B(n10033), .Z(n9791) );
  XNOR2_X1 U9953 ( .A(n10034), .B(n10035), .ZN(n10033) );
  OR2_X1 U9954 ( .A1(n9801), .A2(n9800), .ZN(n9866) );
  XNOR2_X1 U9955 ( .A(n10036), .B(n10037), .ZN(n9800) );
  XOR2_X1 U9956 ( .A(n10038), .B(n10039), .Z(n10036) );
  NOR2_X1 U9957 ( .A1(n7636), .A2(n7872), .ZN(n10039) );
  NAND2_X1 U9958 ( .A1(a_6_), .A2(b_24_), .ZN(n9801) );
  XNOR2_X1 U9959 ( .A(n10040), .B(n10041), .ZN(n9803) );
  NAND2_X1 U9960 ( .A1(n10042), .A2(n10043), .ZN(n10040) );
  XOR2_X1 U9961 ( .A(n10044), .B(n10045), .Z(n9808) );
  XOR2_X1 U9962 ( .A(n10046), .B(n10047), .Z(n10045) );
  NAND2_X1 U9963 ( .A1(a_5_), .A2(b_23_), .ZN(n10047) );
  INV_X1 U9964 ( .A(n8254), .ZN(n8249) );
  XOR2_X1 U9965 ( .A(n10048), .B(n10049), .Z(n8254) );
  XNOR2_X1 U9966 ( .A(n10050), .B(n10051), .ZN(n10048) );
  NOR2_X1 U9967 ( .A1(n7636), .A2(n8942), .ZN(n10051) );
  NAND3_X1 U9968 ( .A1(n10052), .A2(n8245), .A3(n8244), .ZN(n8106) );
  XNOR2_X1 U9969 ( .A(n10053), .B(n10054), .ZN(n8244) );
  NAND2_X1 U9970 ( .A1(n10055), .A2(n10056), .ZN(n10053) );
  NAND2_X1 U9971 ( .A1(n10057), .A2(n10058), .ZN(n8245) );
  NAND3_X1 U9972 ( .A1(b_23_), .A2(n10059), .A3(a_0_), .ZN(n10058) );
  NAND2_X1 U9973 ( .A1(n10050), .A2(n10049), .ZN(n10059) );
  OR2_X1 U9974 ( .A1(n10049), .A2(n10050), .ZN(n10057) );
  AND2_X1 U9975 ( .A1(n10060), .A2(n10061), .ZN(n10050) );
  NAND3_X1 U9976 ( .A1(a_1_), .A2(n10062), .A3(b_23_), .ZN(n10061) );
  OR2_X1 U9977 ( .A1(n9834), .A2(n9832), .ZN(n10062) );
  NAND2_X1 U9978 ( .A1(n9832), .A2(n9834), .ZN(n10060) );
  NAND2_X1 U9979 ( .A1(n10063), .A2(n10064), .ZN(n9834) );
  NAND3_X1 U9980 ( .A1(b_23_), .A2(n10065), .A3(a_2_), .ZN(n10064) );
  NAND2_X1 U9981 ( .A1(n9842), .A2(n9841), .ZN(n10065) );
  OR2_X1 U9982 ( .A1(n9841), .A2(n9842), .ZN(n10063) );
  AND2_X1 U9983 ( .A1(n10066), .A2(n10067), .ZN(n9842) );
  NAND3_X1 U9984 ( .A1(b_23_), .A2(n10068), .A3(a_3_), .ZN(n10067) );
  OR2_X1 U9985 ( .A1(n9850), .A2(n9848), .ZN(n10068) );
  NAND2_X1 U9986 ( .A1(n9848), .A2(n9850), .ZN(n10066) );
  NAND2_X1 U9987 ( .A1(n10069), .A2(n10070), .ZN(n9850) );
  NAND3_X1 U9988 ( .A1(b_23_), .A2(n10071), .A3(a_4_), .ZN(n10070) );
  OR2_X1 U9989 ( .A1(n9858), .A2(n9856), .ZN(n10071) );
  NAND2_X1 U9990 ( .A1(n9856), .A2(n9858), .ZN(n10069) );
  NAND2_X1 U9991 ( .A1(n10072), .A2(n10073), .ZN(n9858) );
  NAND3_X1 U9992 ( .A1(b_23_), .A2(n10074), .A3(a_5_), .ZN(n10073) );
  OR2_X1 U9993 ( .A1(n10046), .A2(n10044), .ZN(n10074) );
  NAND2_X1 U9994 ( .A1(n10044), .A2(n10046), .ZN(n10072) );
  NAND2_X1 U9995 ( .A1(n10042), .A2(n10075), .ZN(n10046) );
  NAND2_X1 U9996 ( .A1(n10041), .A2(n10043), .ZN(n10075) );
  NAND2_X1 U9997 ( .A1(n10076), .A2(n10077), .ZN(n10043) );
  NAND2_X1 U9998 ( .A1(a_6_), .A2(b_23_), .ZN(n10077) );
  INV_X1 U9999 ( .A(n10078), .ZN(n10076) );
  XNOR2_X1 U10000 ( .A(n10079), .B(n10080), .ZN(n10041) );
  XNOR2_X1 U10001 ( .A(n10081), .B(n10082), .ZN(n10080) );
  NAND2_X1 U10002 ( .A1(a_6_), .A2(n10078), .ZN(n10042) );
  NAND2_X1 U10003 ( .A1(n10083), .A2(n10084), .ZN(n10078) );
  NAND3_X1 U10004 ( .A1(b_23_), .A2(n10085), .A3(a_7_), .ZN(n10084) );
  OR2_X1 U10005 ( .A1(n10038), .A2(n10037), .ZN(n10085) );
  NAND2_X1 U10006 ( .A1(n10037), .A2(n10038), .ZN(n10083) );
  NAND2_X1 U10007 ( .A1(n10086), .A2(n10087), .ZN(n10038) );
  NAND2_X1 U10008 ( .A1(n9876), .A2(n10088), .ZN(n10087) );
  OR2_X1 U10009 ( .A1(n9875), .A2(n9873), .ZN(n10088) );
  NOR2_X1 U10010 ( .A1(n8686), .A2(n7636), .ZN(n9876) );
  NAND2_X1 U10011 ( .A1(n9873), .A2(n9875), .ZN(n10086) );
  NAND2_X1 U10012 ( .A1(n10089), .A2(n10090), .ZN(n9875) );
  NAND2_X1 U10013 ( .A1(n10035), .A2(n10091), .ZN(n10090) );
  OR2_X1 U10014 ( .A1(n10034), .A2(n10032), .ZN(n10091) );
  NOR2_X1 U10015 ( .A1(n8052), .A2(n7636), .ZN(n10035) );
  NAND2_X1 U10016 ( .A1(n10032), .A2(n10034), .ZN(n10089) );
  NAND2_X1 U10017 ( .A1(n10030), .A2(n10092), .ZN(n10034) );
  NAND2_X1 U10018 ( .A1(n10029), .A2(n10031), .ZN(n10092) );
  NAND2_X1 U10019 ( .A1(n10093), .A2(n10094), .ZN(n10031) );
  NAND2_X1 U10020 ( .A1(a_10_), .A2(b_23_), .ZN(n10094) );
  INV_X1 U10021 ( .A(n10095), .ZN(n10093) );
  XNOR2_X1 U10022 ( .A(n10096), .B(n10097), .ZN(n10029) );
  XNOR2_X1 U10023 ( .A(n10098), .B(n10099), .ZN(n10097) );
  NAND2_X1 U10024 ( .A1(a_10_), .A2(n10095), .ZN(n10030) );
  NAND2_X1 U10025 ( .A1(n10100), .A2(n10101), .ZN(n10095) );
  NAND3_X1 U10026 ( .A1(b_23_), .A2(n10102), .A3(a_11_), .ZN(n10101) );
  OR2_X1 U10027 ( .A1(n10026), .A2(n10025), .ZN(n10102) );
  NAND2_X1 U10028 ( .A1(n10025), .A2(n10026), .ZN(n10100) );
  NAND2_X1 U10029 ( .A1(n10103), .A2(n10104), .ZN(n10026) );
  NAND3_X1 U10030 ( .A1(b_23_), .A2(n10105), .A3(a_12_), .ZN(n10104) );
  NAND2_X1 U10031 ( .A1(n9892), .A2(n9891), .ZN(n10105) );
  OR2_X1 U10032 ( .A1(n9891), .A2(n9892), .ZN(n10103) );
  AND2_X1 U10033 ( .A1(n10106), .A2(n10107), .ZN(n9892) );
  NAND2_X1 U10034 ( .A1(n10023), .A2(n10108), .ZN(n10107) );
  OR2_X1 U10035 ( .A1(n10022), .A2(n10021), .ZN(n10108) );
  NOR2_X1 U10036 ( .A1(n7789), .A2(n7636), .ZN(n10023) );
  NAND2_X1 U10037 ( .A1(n10021), .A2(n10022), .ZN(n10106) );
  NAND2_X1 U10038 ( .A1(n10018), .A2(n10109), .ZN(n10022) );
  NAND2_X1 U10039 ( .A1(n10017), .A2(n10019), .ZN(n10109) );
  NAND2_X1 U10040 ( .A1(n10110), .A2(n10111), .ZN(n10019) );
  NAND2_X1 U10041 ( .A1(a_14_), .A2(b_23_), .ZN(n10111) );
  INV_X1 U10042 ( .A(n10112), .ZN(n10110) );
  XOR2_X1 U10043 ( .A(n10113), .B(n10114), .Z(n10017) );
  XOR2_X1 U10044 ( .A(n10115), .B(n10116), .Z(n10113) );
  NAND2_X1 U10045 ( .A1(a_14_), .A2(n10112), .ZN(n10018) );
  NAND2_X1 U10046 ( .A1(n10117), .A2(n10118), .ZN(n10112) );
  NAND3_X1 U10047 ( .A1(b_23_), .A2(n10119), .A3(a_15_), .ZN(n10118) );
  OR2_X1 U10048 ( .A1(n10014), .A2(n10012), .ZN(n10119) );
  NAND2_X1 U10049 ( .A1(n10012), .A2(n10014), .ZN(n10117) );
  NAND2_X1 U10050 ( .A1(n10120), .A2(n10121), .ZN(n10014) );
  NAND3_X1 U10051 ( .A1(b_23_), .A2(n10122), .A3(a_16_), .ZN(n10121) );
  OR2_X1 U10052 ( .A1(n10010), .A2(n10008), .ZN(n10122) );
  NAND2_X1 U10053 ( .A1(n10008), .A2(n10010), .ZN(n10120) );
  NAND2_X1 U10054 ( .A1(n10123), .A2(n10124), .ZN(n10010) );
  NAND2_X1 U10055 ( .A1(n10007), .A2(n10125), .ZN(n10124) );
  NAND2_X1 U10056 ( .A1(n10006), .A2(n10005), .ZN(n10125) );
  NOR2_X1 U10057 ( .A1(n7732), .A2(n7636), .ZN(n10007) );
  OR2_X1 U10058 ( .A1(n10005), .A2(n10006), .ZN(n10123) );
  AND2_X1 U10059 ( .A1(n10126), .A2(n10127), .ZN(n10006) );
  NAND3_X1 U10060 ( .A1(b_23_), .A2(n10128), .A3(a_18_), .ZN(n10127) );
  NAND2_X1 U10061 ( .A1(n10002), .A2(n10001), .ZN(n10128) );
  OR2_X1 U10062 ( .A1(n10001), .A2(n10002), .ZN(n10126) );
  AND2_X1 U10063 ( .A1(n10129), .A2(n10130), .ZN(n10002) );
  NAND2_X1 U10064 ( .A1(n9999), .A2(n10131), .ZN(n10130) );
  OR2_X1 U10065 ( .A1(n9998), .A2(n9996), .ZN(n10131) );
  NOR2_X1 U10066 ( .A1(n8045), .A2(n7636), .ZN(n9999) );
  NAND2_X1 U10067 ( .A1(n9996), .A2(n9998), .ZN(n10129) );
  NAND2_X1 U10068 ( .A1(n10132), .A2(n10133), .ZN(n9998) );
  NAND3_X1 U10069 ( .A1(b_23_), .A2(n10134), .A3(a_20_), .ZN(n10133) );
  NAND2_X1 U10070 ( .A1(n9994), .A2(n9993), .ZN(n10134) );
  OR2_X1 U10071 ( .A1(n9993), .A2(n9994), .ZN(n10132) );
  AND2_X1 U10072 ( .A1(n10135), .A2(n10136), .ZN(n9994) );
  NAND2_X1 U10073 ( .A1(n9991), .A2(n10137), .ZN(n10136) );
  OR2_X1 U10074 ( .A1(n9990), .A2(n9989), .ZN(n10137) );
  NOR2_X1 U10075 ( .A1(n7665), .A2(n7636), .ZN(n9991) );
  NAND2_X1 U10076 ( .A1(n9989), .A2(n9990), .ZN(n10135) );
  NAND2_X1 U10077 ( .A1(n10138), .A2(n10139), .ZN(n9990) );
  NAND3_X1 U10078 ( .A1(b_23_), .A2(n10140), .A3(a_22_), .ZN(n10139) );
  OR2_X1 U10079 ( .A1(n9986), .A2(n9984), .ZN(n10140) );
  NAND2_X1 U10080 ( .A1(n9984), .A2(n9986), .ZN(n10138) );
  NAND2_X1 U10081 ( .A1(n10141), .A2(n10142), .ZN(n9986) );
  NAND2_X1 U10082 ( .A1(n7634), .A2(n10143), .ZN(n10142) );
  OR2_X1 U10083 ( .A1(n9983), .A2(n9981), .ZN(n10143) );
  NOR2_X1 U10084 ( .A1(n8042), .A2(n7636), .ZN(n7634) );
  NAND2_X1 U10085 ( .A1(n9981), .A2(n9983), .ZN(n10141) );
  NAND2_X1 U10086 ( .A1(n10144), .A2(n10145), .ZN(n9983) );
  NAND3_X1 U10087 ( .A1(a_24_), .A2(n10146), .A3(b_23_), .ZN(n10145) );
  NAND2_X1 U10088 ( .A1(n9979), .A2(n9978), .ZN(n10146) );
  OR2_X1 U10089 ( .A1(n9978), .A2(n9979), .ZN(n10144) );
  AND2_X1 U10090 ( .A1(n10147), .A2(n10148), .ZN(n9979) );
  NAND2_X1 U10091 ( .A1(n9936), .A2(n10149), .ZN(n10148) );
  OR2_X1 U10092 ( .A1(n9935), .A2(n9934), .ZN(n10149) );
  NOR2_X1 U10093 ( .A1(n7636), .A2(n8039), .ZN(n9936) );
  NAND2_X1 U10094 ( .A1(n9934), .A2(n9935), .ZN(n10147) );
  NAND2_X1 U10095 ( .A1(n9975), .A2(n10150), .ZN(n9935) );
  NAND2_X1 U10096 ( .A1(n9974), .A2(n9976), .ZN(n10150) );
  NAND2_X1 U10097 ( .A1(n10151), .A2(n10152), .ZN(n9976) );
  NAND2_X1 U10098 ( .A1(b_23_), .A2(a_26_), .ZN(n10152) );
  INV_X1 U10099 ( .A(n10153), .ZN(n10151) );
  XNOR2_X1 U10100 ( .A(n10154), .B(n10155), .ZN(n9974) );
  NAND2_X1 U10101 ( .A1(n10156), .A2(n10157), .ZN(n10154) );
  NAND2_X1 U10102 ( .A1(a_26_), .A2(n10153), .ZN(n9975) );
  NAND2_X1 U10103 ( .A1(n9946), .A2(n10158), .ZN(n10153) );
  NAND2_X1 U10104 ( .A1(n9945), .A2(n9947), .ZN(n10158) );
  NAND2_X1 U10105 ( .A1(n10159), .A2(n10160), .ZN(n9947) );
  NAND2_X1 U10106 ( .A1(b_23_), .A2(a_27_), .ZN(n10160) );
  INV_X1 U10107 ( .A(n10161), .ZN(n10159) );
  XNOR2_X1 U10108 ( .A(n10162), .B(n10163), .ZN(n9945) );
  XOR2_X1 U10109 ( .A(n10164), .B(n10165), .Z(n10162) );
  NAND2_X1 U10110 ( .A1(b_22_), .A2(a_28_), .ZN(n10164) );
  NAND2_X1 U10111 ( .A1(a_27_), .A2(n10161), .ZN(n9946) );
  NAND2_X1 U10112 ( .A1(n10166), .A2(n10167), .ZN(n10161) );
  NAND3_X1 U10113 ( .A1(a_28_), .A2(n10168), .A3(b_23_), .ZN(n10167) );
  NAND2_X1 U10114 ( .A1(n9955), .A2(n9953), .ZN(n10168) );
  OR2_X1 U10115 ( .A1(n9953), .A2(n9955), .ZN(n10166) );
  AND2_X1 U10116 ( .A1(n10169), .A2(n10170), .ZN(n9955) );
  NAND2_X1 U10117 ( .A1(n9970), .A2(n10171), .ZN(n10170) );
  OR2_X1 U10118 ( .A1(n9971), .A2(n9972), .ZN(n10171) );
  NOR2_X1 U10119 ( .A1(n7636), .A2(n7545), .ZN(n9970) );
  NAND2_X1 U10120 ( .A1(n9972), .A2(n9971), .ZN(n10169) );
  NAND2_X1 U10121 ( .A1(n10172), .A2(n10173), .ZN(n9971) );
  NAND2_X1 U10122 ( .A1(b_21_), .A2(n10174), .ZN(n10173) );
  NAND2_X1 U10123 ( .A1(n7527), .A2(n10175), .ZN(n10174) );
  NAND2_X1 U10124 ( .A1(a_31_), .A2(n9968), .ZN(n10175) );
  NAND2_X1 U10125 ( .A1(b_22_), .A2(n10176), .ZN(n10172) );
  NAND2_X1 U10126 ( .A1(n7531), .A2(n10177), .ZN(n10176) );
  NAND2_X1 U10127 ( .A1(a_30_), .A2(n7667), .ZN(n10177) );
  AND3_X1 U10128 ( .A1(b_22_), .A2(b_23_), .A3(n7494), .ZN(n9972) );
  XNOR2_X1 U10129 ( .A(n10178), .B(n10179), .ZN(n9953) );
  XOR2_X1 U10130 ( .A(n10180), .B(n10181), .Z(n10178) );
  XNOR2_X1 U10131 ( .A(n10182), .B(n10183), .ZN(n9934) );
  NAND2_X1 U10132 ( .A1(n10184), .A2(n10185), .ZN(n10182) );
  XNOR2_X1 U10133 ( .A(n10186), .B(n10187), .ZN(n9978) );
  XOR2_X1 U10134 ( .A(n10188), .B(n10189), .Z(n10186) );
  XNOR2_X1 U10135 ( .A(n10190), .B(n10191), .ZN(n9981) );
  XNOR2_X1 U10136 ( .A(n10192), .B(n10193), .ZN(n10190) );
  NOR2_X1 U10137 ( .A1(n8041), .A2(n9968), .ZN(n10193) );
  XNOR2_X1 U10138 ( .A(n10194), .B(n10195), .ZN(n9984) );
  XNOR2_X1 U10139 ( .A(n10196), .B(n10197), .ZN(n10195) );
  XNOR2_X1 U10140 ( .A(n10198), .B(n10199), .ZN(n9989) );
  XNOR2_X1 U10141 ( .A(n10200), .B(n7655), .ZN(n10199) );
  XNOR2_X1 U10142 ( .A(n10201), .B(n10202), .ZN(n9993) );
  XOR2_X1 U10143 ( .A(n10203), .B(n10204), .Z(n10201) );
  XNOR2_X1 U10144 ( .A(n10205), .B(n10206), .ZN(n9996) );
  XNOR2_X1 U10145 ( .A(n10207), .B(n10208), .ZN(n10205) );
  NOR2_X1 U10146 ( .A1(n9968), .A2(n8044), .ZN(n10208) );
  XOR2_X1 U10147 ( .A(n10209), .B(n10210), .Z(n10001) );
  XNOR2_X1 U10148 ( .A(n10211), .B(n10212), .ZN(n10210) );
  XNOR2_X1 U10149 ( .A(n10213), .B(n10214), .ZN(n10005) );
  XOR2_X1 U10150 ( .A(n10215), .B(n10216), .Z(n10213) );
  NOR2_X1 U10151 ( .A1(n9968), .A2(n8047), .ZN(n10216) );
  XOR2_X1 U10152 ( .A(n10217), .B(n10218), .Z(n10008) );
  XOR2_X1 U10153 ( .A(n10219), .B(n10220), .Z(n10217) );
  XNOR2_X1 U10154 ( .A(n10221), .B(n10222), .ZN(n10012) );
  XOR2_X1 U10155 ( .A(n10223), .B(n10224), .Z(n10222) );
  NAND2_X1 U10156 ( .A1(a_16_), .A2(b_22_), .ZN(n10224) );
  XNOR2_X1 U10157 ( .A(n10225), .B(n10226), .ZN(n10021) );
  XNOR2_X1 U10158 ( .A(n10227), .B(n10228), .ZN(n10225) );
  NOR2_X1 U10159 ( .A1(n9968), .A2(n8049), .ZN(n10228) );
  XOR2_X1 U10160 ( .A(n10229), .B(n10230), .Z(n9891) );
  XNOR2_X1 U10161 ( .A(n10231), .B(n10232), .ZN(n10230) );
  XNOR2_X1 U10162 ( .A(n10233), .B(n10234), .ZN(n10025) );
  XNOR2_X1 U10163 ( .A(n10235), .B(n10236), .ZN(n10233) );
  NOR2_X1 U10164 ( .A1(n9968), .A2(n8669), .ZN(n10236) );
  XNOR2_X1 U10165 ( .A(n10237), .B(n10238), .ZN(n10032) );
  XNOR2_X1 U10166 ( .A(n10239), .B(n10240), .ZN(n10237) );
  NOR2_X1 U10167 ( .A1(n9968), .A2(n8051), .ZN(n10240) );
  XNOR2_X1 U10168 ( .A(n10241), .B(n10242), .ZN(n9873) );
  XOR2_X1 U10169 ( .A(n10243), .B(n10244), .Z(n10242) );
  NAND2_X1 U10170 ( .A1(a_9_), .A2(b_22_), .ZN(n10244) );
  XNOR2_X1 U10171 ( .A(n10245), .B(n10246), .ZN(n10037) );
  XNOR2_X1 U10172 ( .A(n10247), .B(n10248), .ZN(n10245) );
  XNOR2_X1 U10173 ( .A(n10249), .B(n10250), .ZN(n10044) );
  XNOR2_X1 U10174 ( .A(n10251), .B(n10252), .ZN(n10249) );
  NOR2_X1 U10175 ( .A1(n9968), .A2(n7887), .ZN(n10252) );
  XNOR2_X1 U10176 ( .A(n10253), .B(n10254), .ZN(n9856) );
  XNOR2_X1 U10177 ( .A(n10255), .B(n10256), .ZN(n10254) );
  XOR2_X1 U10178 ( .A(n10257), .B(n10258), .Z(n9848) );
  XOR2_X1 U10179 ( .A(n10259), .B(n10260), .Z(n10257) );
  XNOR2_X1 U10180 ( .A(n10261), .B(n10262), .ZN(n9841) );
  XOR2_X1 U10181 ( .A(n10263), .B(n10264), .Z(n10261) );
  XOR2_X1 U10182 ( .A(n10265), .B(n10266), .Z(n9832) );
  XOR2_X1 U10183 ( .A(n10267), .B(n10268), .Z(n10265) );
  XNOR2_X1 U10184 ( .A(n10269), .B(n10270), .ZN(n10049) );
  XOR2_X1 U10185 ( .A(n10271), .B(n10272), .Z(n10269) );
  NOR2_X1 U10186 ( .A1(n7957), .A2(n9968), .ZN(n10272) );
  XOR2_X1 U10187 ( .A(n8240), .B(n8239), .Z(n10052) );
  NAND4_X1 U10188 ( .A1(n8239), .A2(n8238), .A3(n8240), .A4(n8234), .ZN(n8112)
         );
  INV_X1 U10189 ( .A(n10273), .ZN(n8234) );
  NAND2_X1 U10190 ( .A1(n10055), .A2(n10274), .ZN(n8240) );
  NAND2_X1 U10191 ( .A1(n10054), .A2(n10056), .ZN(n10274) );
  NAND2_X1 U10192 ( .A1(n10275), .A2(n10276), .ZN(n10056) );
  NAND2_X1 U10193 ( .A1(a_0_), .A2(b_22_), .ZN(n10276) );
  INV_X1 U10194 ( .A(n10277), .ZN(n10275) );
  XOR2_X1 U10195 ( .A(n10278), .B(n10279), .Z(n10054) );
  XOR2_X1 U10196 ( .A(n10280), .B(n10281), .Z(n10278) );
  NOR2_X1 U10197 ( .A1(n7957), .A2(n7667), .ZN(n10281) );
  NAND2_X1 U10198 ( .A1(a_0_), .A2(n10277), .ZN(n10055) );
  NAND2_X1 U10199 ( .A1(n10282), .A2(n10283), .ZN(n10277) );
  NAND3_X1 U10200 ( .A1(a_1_), .A2(n10284), .A3(b_22_), .ZN(n10283) );
  OR2_X1 U10201 ( .A1(n10271), .A2(n10270), .ZN(n10284) );
  NAND2_X1 U10202 ( .A1(n10270), .A2(n10271), .ZN(n10282) );
  NAND2_X1 U10203 ( .A1(n10285), .A2(n10286), .ZN(n10271) );
  NAND2_X1 U10204 ( .A1(n10268), .A2(n10287), .ZN(n10286) );
  OR2_X1 U10205 ( .A1(n10267), .A2(n10266), .ZN(n10287) );
  NOR2_X1 U10206 ( .A1(n8056), .A2(n9968), .ZN(n10268) );
  NAND2_X1 U10207 ( .A1(n10266), .A2(n10267), .ZN(n10285) );
  NAND2_X1 U10208 ( .A1(n10288), .A2(n10289), .ZN(n10267) );
  NAND2_X1 U10209 ( .A1(n10264), .A2(n10290), .ZN(n10289) );
  OR2_X1 U10210 ( .A1(n10263), .A2(n10262), .ZN(n10290) );
  NOR2_X1 U10211 ( .A1(n7937), .A2(n9968), .ZN(n10264) );
  NAND2_X1 U10212 ( .A1(n10262), .A2(n10263), .ZN(n10288) );
  NAND2_X1 U10213 ( .A1(n10291), .A2(n10292), .ZN(n10263) );
  NAND2_X1 U10214 ( .A1(n10260), .A2(n10293), .ZN(n10292) );
  OR2_X1 U10215 ( .A1(n10259), .A2(n10258), .ZN(n10293) );
  NOR2_X1 U10216 ( .A1(n7916), .A2(n9968), .ZN(n10260) );
  NAND2_X1 U10217 ( .A1(n10258), .A2(n10259), .ZN(n10291) );
  NAND2_X1 U10218 ( .A1(n10294), .A2(n10295), .ZN(n10259) );
  NAND2_X1 U10219 ( .A1(n10256), .A2(n10296), .ZN(n10295) );
  OR2_X1 U10220 ( .A1(n10255), .A2(n10253), .ZN(n10296) );
  NOR2_X1 U10221 ( .A1(n7908), .A2(n9968), .ZN(n10256) );
  NAND2_X1 U10222 ( .A1(n10253), .A2(n10255), .ZN(n10294) );
  NAND2_X1 U10223 ( .A1(n10297), .A2(n10298), .ZN(n10255) );
  NAND3_X1 U10224 ( .A1(b_22_), .A2(n10299), .A3(a_6_), .ZN(n10298) );
  NAND2_X1 U10225 ( .A1(n10251), .A2(n10250), .ZN(n10299) );
  OR2_X1 U10226 ( .A1(n10250), .A2(n10251), .ZN(n10297) );
  AND2_X1 U10227 ( .A1(n10300), .A2(n10301), .ZN(n10251) );
  NAND2_X1 U10228 ( .A1(n10082), .A2(n10302), .ZN(n10301) );
  OR2_X1 U10229 ( .A1(n10081), .A2(n10079), .ZN(n10302) );
  NOR2_X1 U10230 ( .A1(n7872), .A2(n9968), .ZN(n10082) );
  NAND2_X1 U10231 ( .A1(n10079), .A2(n10081), .ZN(n10300) );
  NAND2_X1 U10232 ( .A1(n10303), .A2(n10304), .ZN(n10081) );
  NAND2_X1 U10233 ( .A1(n10248), .A2(n10305), .ZN(n10304) );
  NAND2_X1 U10234 ( .A1(n10247), .A2(n10246), .ZN(n10305) );
  NOR2_X1 U10235 ( .A1(n8686), .A2(n9968), .ZN(n10248) );
  OR2_X1 U10236 ( .A1(n10246), .A2(n10247), .ZN(n10303) );
  AND2_X1 U10237 ( .A1(n10306), .A2(n10307), .ZN(n10247) );
  NAND3_X1 U10238 ( .A1(b_22_), .A2(n10308), .A3(a_9_), .ZN(n10307) );
  OR2_X1 U10239 ( .A1(n10243), .A2(n10241), .ZN(n10308) );
  NAND2_X1 U10240 ( .A1(n10241), .A2(n10243), .ZN(n10306) );
  NAND2_X1 U10241 ( .A1(n10309), .A2(n10310), .ZN(n10243) );
  NAND3_X1 U10242 ( .A1(b_22_), .A2(n10311), .A3(a_10_), .ZN(n10310) );
  NAND2_X1 U10243 ( .A1(n10239), .A2(n10238), .ZN(n10311) );
  OR2_X1 U10244 ( .A1(n10238), .A2(n10239), .ZN(n10309) );
  AND2_X1 U10245 ( .A1(n10312), .A2(n10313), .ZN(n10239) );
  NAND2_X1 U10246 ( .A1(n10099), .A2(n10314), .ZN(n10313) );
  OR2_X1 U10247 ( .A1(n10098), .A2(n10096), .ZN(n10314) );
  NOR2_X1 U10248 ( .A1(n7811), .A2(n9968), .ZN(n10099) );
  NAND2_X1 U10249 ( .A1(n10096), .A2(n10098), .ZN(n10312) );
  NAND2_X1 U10250 ( .A1(n10315), .A2(n10316), .ZN(n10098) );
  NAND3_X1 U10251 ( .A1(b_22_), .A2(n10317), .A3(a_12_), .ZN(n10316) );
  NAND2_X1 U10252 ( .A1(n10235), .A2(n10234), .ZN(n10317) );
  OR2_X1 U10253 ( .A1(n10234), .A2(n10235), .ZN(n10315) );
  AND2_X1 U10254 ( .A1(n10318), .A2(n10319), .ZN(n10235) );
  NAND2_X1 U10255 ( .A1(n10232), .A2(n10320), .ZN(n10319) );
  OR2_X1 U10256 ( .A1(n10231), .A2(n10229), .ZN(n10320) );
  NOR2_X1 U10257 ( .A1(n7789), .A2(n9968), .ZN(n10232) );
  NAND2_X1 U10258 ( .A1(n10229), .A2(n10231), .ZN(n10318) );
  NAND2_X1 U10259 ( .A1(n10321), .A2(n10322), .ZN(n10231) );
  NAND3_X1 U10260 ( .A1(b_22_), .A2(n10323), .A3(a_14_), .ZN(n10322) );
  NAND2_X1 U10261 ( .A1(n10227), .A2(n10226), .ZN(n10323) );
  OR2_X1 U10262 ( .A1(n10226), .A2(n10227), .ZN(n10321) );
  AND2_X1 U10263 ( .A1(n10324), .A2(n10325), .ZN(n10227) );
  NAND2_X1 U10264 ( .A1(n10116), .A2(n10326), .ZN(n10325) );
  OR2_X1 U10265 ( .A1(n10115), .A2(n10114), .ZN(n10326) );
  NOR2_X1 U10266 ( .A1(n7754), .A2(n9968), .ZN(n10116) );
  NAND2_X1 U10267 ( .A1(n10114), .A2(n10115), .ZN(n10324) );
  NAND2_X1 U10268 ( .A1(n10327), .A2(n10328), .ZN(n10115) );
  NAND3_X1 U10269 ( .A1(b_22_), .A2(n10329), .A3(a_16_), .ZN(n10328) );
  OR2_X1 U10270 ( .A1(n10223), .A2(n10221), .ZN(n10329) );
  NAND2_X1 U10271 ( .A1(n10221), .A2(n10223), .ZN(n10327) );
  NAND2_X1 U10272 ( .A1(n10330), .A2(n10331), .ZN(n10223) );
  NAND2_X1 U10273 ( .A1(n10220), .A2(n10332), .ZN(n10331) );
  OR2_X1 U10274 ( .A1(n10219), .A2(n10218), .ZN(n10332) );
  NOR2_X1 U10275 ( .A1(n7732), .A2(n9968), .ZN(n10220) );
  NAND2_X1 U10276 ( .A1(n10218), .A2(n10219), .ZN(n10330) );
  NAND2_X1 U10277 ( .A1(n10333), .A2(n10334), .ZN(n10219) );
  NAND3_X1 U10278 ( .A1(b_22_), .A2(n10335), .A3(a_18_), .ZN(n10334) );
  OR2_X1 U10279 ( .A1(n10215), .A2(n10214), .ZN(n10335) );
  NAND2_X1 U10280 ( .A1(n10214), .A2(n10215), .ZN(n10333) );
  NAND2_X1 U10281 ( .A1(n10336), .A2(n10337), .ZN(n10215) );
  NAND2_X1 U10282 ( .A1(n10212), .A2(n10338), .ZN(n10337) );
  OR2_X1 U10283 ( .A1(n10211), .A2(n10209), .ZN(n10338) );
  NOR2_X1 U10284 ( .A1(n8045), .A2(n9968), .ZN(n10212) );
  NAND2_X1 U10285 ( .A1(n10209), .A2(n10211), .ZN(n10336) );
  NAND2_X1 U10286 ( .A1(n10339), .A2(n10340), .ZN(n10211) );
  NAND3_X1 U10287 ( .A1(b_22_), .A2(n10341), .A3(a_20_), .ZN(n10340) );
  NAND2_X1 U10288 ( .A1(n10207), .A2(n10206), .ZN(n10341) );
  OR2_X1 U10289 ( .A1(n10206), .A2(n10207), .ZN(n10339) );
  AND2_X1 U10290 ( .A1(n10342), .A2(n10343), .ZN(n10207) );
  NAND2_X1 U10291 ( .A1(n10204), .A2(n10344), .ZN(n10343) );
  OR2_X1 U10292 ( .A1(n10203), .A2(n10202), .ZN(n10344) );
  NOR2_X1 U10293 ( .A1(n7665), .A2(n9968), .ZN(n10204) );
  NAND2_X1 U10294 ( .A1(n10202), .A2(n10203), .ZN(n10342) );
  NAND2_X1 U10295 ( .A1(n10345), .A2(n10346), .ZN(n10203) );
  NAND2_X1 U10296 ( .A1(n10198), .A2(n10347), .ZN(n10346) );
  OR2_X1 U10297 ( .A1(n10200), .A2(n7655), .ZN(n10347) );
  XNOR2_X1 U10298 ( .A(n10348), .B(n10349), .ZN(n10198) );
  XNOR2_X1 U10299 ( .A(n10350), .B(n10351), .ZN(n10349) );
  NAND2_X1 U10300 ( .A1(n7655), .A2(n10200), .ZN(n10345) );
  NAND2_X1 U10301 ( .A1(n10352), .A2(n10353), .ZN(n10200) );
  NAND2_X1 U10302 ( .A1(n10197), .A2(n10354), .ZN(n10353) );
  OR2_X1 U10303 ( .A1(n10196), .A2(n10194), .ZN(n10354) );
  NOR2_X1 U10304 ( .A1(n9968), .A2(n8042), .ZN(n10197) );
  NAND2_X1 U10305 ( .A1(n10194), .A2(n10196), .ZN(n10352) );
  NAND2_X1 U10306 ( .A1(n10355), .A2(n10356), .ZN(n10196) );
  NAND3_X1 U10307 ( .A1(a_24_), .A2(n10357), .A3(b_22_), .ZN(n10356) );
  NAND2_X1 U10308 ( .A1(n10192), .A2(n10191), .ZN(n10357) );
  OR2_X1 U10309 ( .A1(n10191), .A2(n10192), .ZN(n10355) );
  AND2_X1 U10310 ( .A1(n10358), .A2(n10359), .ZN(n10192) );
  NAND2_X1 U10311 ( .A1(n10189), .A2(n10360), .ZN(n10359) );
  OR2_X1 U10312 ( .A1(n10188), .A2(n10187), .ZN(n10360) );
  NOR2_X1 U10313 ( .A1(n9968), .A2(n8039), .ZN(n10189) );
  NAND2_X1 U10314 ( .A1(n10187), .A2(n10188), .ZN(n10358) );
  NAND2_X1 U10315 ( .A1(n10184), .A2(n10361), .ZN(n10188) );
  NAND2_X1 U10316 ( .A1(n10183), .A2(n10185), .ZN(n10361) );
  NAND2_X1 U10317 ( .A1(n10362), .A2(n10363), .ZN(n10185) );
  NAND2_X1 U10318 ( .A1(b_22_), .A2(a_26_), .ZN(n10363) );
  INV_X1 U10319 ( .A(n10364), .ZN(n10362) );
  XNOR2_X1 U10320 ( .A(n10365), .B(n10366), .ZN(n10183) );
  NAND2_X1 U10321 ( .A1(n10367), .A2(n10368), .ZN(n10365) );
  NAND2_X1 U10322 ( .A1(a_26_), .A2(n10364), .ZN(n10184) );
  NAND2_X1 U10323 ( .A1(n10156), .A2(n10369), .ZN(n10364) );
  NAND2_X1 U10324 ( .A1(n10155), .A2(n10157), .ZN(n10369) );
  NAND2_X1 U10325 ( .A1(n10370), .A2(n10371), .ZN(n10157) );
  NAND2_X1 U10326 ( .A1(b_22_), .A2(a_27_), .ZN(n10371) );
  INV_X1 U10327 ( .A(n10372), .ZN(n10370) );
  XNOR2_X1 U10328 ( .A(n10373), .B(n10374), .ZN(n10155) );
  XOR2_X1 U10329 ( .A(n10375), .B(n10376), .Z(n10373) );
  NAND2_X1 U10330 ( .A1(b_21_), .A2(a_28_), .ZN(n10375) );
  NAND2_X1 U10331 ( .A1(a_27_), .A2(n10372), .ZN(n10156) );
  NAND2_X1 U10332 ( .A1(n10377), .A2(n10378), .ZN(n10372) );
  NAND3_X1 U10333 ( .A1(a_28_), .A2(n10379), .A3(b_22_), .ZN(n10378) );
  NAND2_X1 U10334 ( .A1(n10165), .A2(n10163), .ZN(n10379) );
  OR2_X1 U10335 ( .A1(n10163), .A2(n10165), .ZN(n10377) );
  AND2_X1 U10336 ( .A1(n10380), .A2(n10381), .ZN(n10165) );
  NAND2_X1 U10337 ( .A1(n10179), .A2(n10382), .ZN(n10381) );
  OR2_X1 U10338 ( .A1(n10180), .A2(n10181), .ZN(n10382) );
  NOR2_X1 U10339 ( .A1(n9968), .A2(n7545), .ZN(n10179) );
  NAND2_X1 U10340 ( .A1(n10181), .A2(n10180), .ZN(n10380) );
  NAND2_X1 U10341 ( .A1(n10383), .A2(n10384), .ZN(n10180) );
  NAND2_X1 U10342 ( .A1(b_20_), .A2(n10385), .ZN(n10384) );
  NAND2_X1 U10343 ( .A1(n7527), .A2(n10386), .ZN(n10385) );
  NAND2_X1 U10344 ( .A1(a_31_), .A2(n7667), .ZN(n10386) );
  NAND2_X1 U10345 ( .A1(b_21_), .A2(n10387), .ZN(n10383) );
  NAND2_X1 U10346 ( .A1(n7531), .A2(n10388), .ZN(n10387) );
  NAND2_X1 U10347 ( .A1(a_30_), .A2(n8043), .ZN(n10388) );
  AND3_X1 U10348 ( .A1(b_22_), .A2(b_21_), .A3(n7494), .ZN(n10181) );
  XNOR2_X1 U10349 ( .A(n10389), .B(n10390), .ZN(n10163) );
  XOR2_X1 U10350 ( .A(n10391), .B(n10392), .Z(n10389) );
  XNOR2_X1 U10351 ( .A(n10393), .B(n10394), .ZN(n10187) );
  NAND2_X1 U10352 ( .A1(n10395), .A2(n10396), .ZN(n10393) );
  XNOR2_X1 U10353 ( .A(n10397), .B(n10398), .ZN(n10191) );
  XOR2_X1 U10354 ( .A(n10399), .B(n10400), .Z(n10397) );
  XNOR2_X1 U10355 ( .A(n10401), .B(n10402), .ZN(n10194) );
  XNOR2_X1 U10356 ( .A(n10403), .B(n10404), .ZN(n10401) );
  NOR2_X1 U10357 ( .A1(n8041), .A2(n7667), .ZN(n10404) );
  NOR2_X1 U10358 ( .A1(n9968), .A2(n7650), .ZN(n7655) );
  XNOR2_X1 U10359 ( .A(n10405), .B(n10406), .ZN(n10202) );
  XOR2_X1 U10360 ( .A(n10407), .B(n10408), .Z(n10406) );
  NAND2_X1 U10361 ( .A1(b_21_), .A2(a_22_), .ZN(n10408) );
  XNOR2_X1 U10362 ( .A(n10409), .B(n10410), .ZN(n10206) );
  XOR2_X1 U10363 ( .A(n10411), .B(n7662), .Z(n10409) );
  XNOR2_X1 U10364 ( .A(n10412), .B(n10413), .ZN(n10209) );
  XNOR2_X1 U10365 ( .A(n10414), .B(n10415), .ZN(n10412) );
  NOR2_X1 U10366 ( .A1(n7667), .A2(n8044), .ZN(n10415) );
  XNOR2_X1 U10367 ( .A(n10416), .B(n10417), .ZN(n10214) );
  XNOR2_X1 U10368 ( .A(n10418), .B(n10419), .ZN(n10417) );
  XNOR2_X1 U10369 ( .A(n10420), .B(n10421), .ZN(n10218) );
  XNOR2_X1 U10370 ( .A(n10422), .B(n10423), .ZN(n10420) );
  NOR2_X1 U10371 ( .A1(n7667), .A2(n8047), .ZN(n10423) );
  XNOR2_X1 U10372 ( .A(n10424), .B(n10425), .ZN(n10221) );
  XNOR2_X1 U10373 ( .A(n10426), .B(n10427), .ZN(n10425) );
  XNOR2_X1 U10374 ( .A(n10428), .B(n10429), .ZN(n10114) );
  XNOR2_X1 U10375 ( .A(n10430), .B(n10431), .ZN(n10428) );
  NOR2_X1 U10376 ( .A1(n7667), .A2(n8438), .ZN(n10431) );
  XNOR2_X1 U10377 ( .A(n10432), .B(n10433), .ZN(n10226) );
  XOR2_X1 U10378 ( .A(n10434), .B(n10435), .Z(n10432) );
  XNOR2_X1 U10379 ( .A(n10436), .B(n10437), .ZN(n10229) );
  XNOR2_X1 U10380 ( .A(n10438), .B(n10439), .ZN(n10436) );
  NOR2_X1 U10381 ( .A1(n7667), .A2(n8049), .ZN(n10439) );
  XNOR2_X1 U10382 ( .A(n10440), .B(n10441), .ZN(n10234) );
  XOR2_X1 U10383 ( .A(n10442), .B(n10443), .Z(n10440) );
  XNOR2_X1 U10384 ( .A(n10444), .B(n10445), .ZN(n10096) );
  XOR2_X1 U10385 ( .A(n10446), .B(n10447), .Z(n10445) );
  NAND2_X1 U10386 ( .A1(a_12_), .A2(b_21_), .ZN(n10447) );
  XOR2_X1 U10387 ( .A(n10448), .B(n10449), .Z(n10238) );
  XNOR2_X1 U10388 ( .A(n10450), .B(n10451), .ZN(n10449) );
  XOR2_X1 U10389 ( .A(n10452), .B(n10453), .Z(n10241) );
  XOR2_X1 U10390 ( .A(n10454), .B(n10455), .Z(n10452) );
  XNOR2_X1 U10391 ( .A(n10456), .B(n10457), .ZN(n10246) );
  XOR2_X1 U10392 ( .A(n10458), .B(n10459), .Z(n10456) );
  NOR2_X1 U10393 ( .A1(n7667), .A2(n8052), .ZN(n10459) );
  XNOR2_X1 U10394 ( .A(n10460), .B(n10461), .ZN(n10079) );
  XOR2_X1 U10395 ( .A(n10462), .B(n10463), .Z(n10461) );
  NAND2_X1 U10396 ( .A1(a_8_), .A2(b_21_), .ZN(n10463) );
  XOR2_X1 U10397 ( .A(n10464), .B(n10465), .Z(n10250) );
  XOR2_X1 U10398 ( .A(n10466), .B(n10467), .Z(n10465) );
  NAND2_X1 U10399 ( .A1(a_7_), .A2(b_21_), .ZN(n10467) );
  XNOR2_X1 U10400 ( .A(n10468), .B(n10469), .ZN(n10253) );
  XNOR2_X1 U10401 ( .A(n10470), .B(n10471), .ZN(n10468) );
  NOR2_X1 U10402 ( .A1(n7667), .A2(n7887), .ZN(n10471) );
  XNOR2_X1 U10403 ( .A(n10472), .B(n10473), .ZN(n10258) );
  XNOR2_X1 U10404 ( .A(n10474), .B(n10475), .ZN(n10472) );
  NOR2_X1 U10405 ( .A1(n7667), .A2(n7908), .ZN(n10475) );
  XNOR2_X1 U10406 ( .A(n10476), .B(n10477), .ZN(n10262) );
  XNOR2_X1 U10407 ( .A(n10478), .B(n10479), .ZN(n10476) );
  NOR2_X1 U10408 ( .A1(n7667), .A2(n7916), .ZN(n10479) );
  XNOR2_X1 U10409 ( .A(n10480), .B(n10481), .ZN(n10266) );
  XOR2_X1 U10410 ( .A(n10482), .B(n10483), .Z(n10481) );
  NAND2_X1 U10411 ( .A1(a_3_), .A2(b_21_), .ZN(n10483) );
  XNOR2_X1 U10412 ( .A(n10484), .B(n10485), .ZN(n10270) );
  XOR2_X1 U10413 ( .A(n10486), .B(n10487), .Z(n10485) );
  NAND2_X1 U10414 ( .A1(a_2_), .A2(b_21_), .ZN(n10487) );
  NAND2_X1 U10415 ( .A1(n10488), .A2(n10489), .ZN(n8238) );
  XNOR2_X1 U10416 ( .A(n10490), .B(n10491), .ZN(n8239) );
  XNOR2_X1 U10417 ( .A(n10492), .B(n10493), .ZN(n10491) );
  NAND2_X1 U10418 ( .A1(n10494), .A2(n10273), .ZN(n8117) );
  NOR2_X1 U10419 ( .A1(n10489), .A2(n10488), .ZN(n10273) );
  AND2_X1 U10420 ( .A1(n10495), .A2(n10496), .ZN(n10488) );
  NAND2_X1 U10421 ( .A1(n10493), .A2(n10497), .ZN(n10496) );
  OR2_X1 U10422 ( .A1(n10492), .A2(n10490), .ZN(n10497) );
  NOR2_X1 U10423 ( .A1(n8942), .A2(n7667), .ZN(n10493) );
  NAND2_X1 U10424 ( .A1(n10490), .A2(n10492), .ZN(n10495) );
  NAND2_X1 U10425 ( .A1(n10498), .A2(n10499), .ZN(n10492) );
  NAND3_X1 U10426 ( .A1(a_1_), .A2(n10500), .A3(b_21_), .ZN(n10499) );
  OR2_X1 U10427 ( .A1(n10280), .A2(n10279), .ZN(n10500) );
  NAND2_X1 U10428 ( .A1(n10279), .A2(n10280), .ZN(n10498) );
  NAND2_X1 U10429 ( .A1(n10501), .A2(n10502), .ZN(n10280) );
  NAND3_X1 U10430 ( .A1(b_21_), .A2(n10503), .A3(a_2_), .ZN(n10502) );
  OR2_X1 U10431 ( .A1(n10486), .A2(n10484), .ZN(n10503) );
  NAND2_X1 U10432 ( .A1(n10484), .A2(n10486), .ZN(n10501) );
  NAND2_X1 U10433 ( .A1(n10504), .A2(n10505), .ZN(n10486) );
  NAND3_X1 U10434 ( .A1(b_21_), .A2(n10506), .A3(a_3_), .ZN(n10505) );
  OR2_X1 U10435 ( .A1(n10482), .A2(n10480), .ZN(n10506) );
  NAND2_X1 U10436 ( .A1(n10480), .A2(n10482), .ZN(n10504) );
  NAND2_X1 U10437 ( .A1(n10507), .A2(n10508), .ZN(n10482) );
  NAND3_X1 U10438 ( .A1(b_21_), .A2(n10509), .A3(a_4_), .ZN(n10508) );
  NAND2_X1 U10439 ( .A1(n10478), .A2(n10477), .ZN(n10509) );
  OR2_X1 U10440 ( .A1(n10477), .A2(n10478), .ZN(n10507) );
  AND2_X1 U10441 ( .A1(n10510), .A2(n10511), .ZN(n10478) );
  NAND3_X1 U10442 ( .A1(b_21_), .A2(n10512), .A3(a_5_), .ZN(n10511) );
  NAND2_X1 U10443 ( .A1(n10474), .A2(n10473), .ZN(n10512) );
  OR2_X1 U10444 ( .A1(n10473), .A2(n10474), .ZN(n10510) );
  AND2_X1 U10445 ( .A1(n10513), .A2(n10514), .ZN(n10474) );
  NAND3_X1 U10446 ( .A1(b_21_), .A2(n10515), .A3(a_6_), .ZN(n10514) );
  NAND2_X1 U10447 ( .A1(n10470), .A2(n10469), .ZN(n10515) );
  OR2_X1 U10448 ( .A1(n10469), .A2(n10470), .ZN(n10513) );
  AND2_X1 U10449 ( .A1(n10516), .A2(n10517), .ZN(n10470) );
  NAND3_X1 U10450 ( .A1(b_21_), .A2(n10518), .A3(a_7_), .ZN(n10517) );
  OR2_X1 U10451 ( .A1(n10466), .A2(n10464), .ZN(n10518) );
  NAND2_X1 U10452 ( .A1(n10464), .A2(n10466), .ZN(n10516) );
  NAND2_X1 U10453 ( .A1(n10519), .A2(n10520), .ZN(n10466) );
  NAND3_X1 U10454 ( .A1(b_21_), .A2(n10521), .A3(a_8_), .ZN(n10520) );
  OR2_X1 U10455 ( .A1(n10462), .A2(n10460), .ZN(n10521) );
  NAND2_X1 U10456 ( .A1(n10460), .A2(n10462), .ZN(n10519) );
  NAND2_X1 U10457 ( .A1(n10522), .A2(n10523), .ZN(n10462) );
  NAND3_X1 U10458 ( .A1(b_21_), .A2(n10524), .A3(a_9_), .ZN(n10523) );
  OR2_X1 U10459 ( .A1(n10458), .A2(n10457), .ZN(n10524) );
  NAND2_X1 U10460 ( .A1(n10457), .A2(n10458), .ZN(n10522) );
  NAND2_X1 U10461 ( .A1(n10525), .A2(n10526), .ZN(n10458) );
  NAND2_X1 U10462 ( .A1(n10455), .A2(n10527), .ZN(n10526) );
  OR2_X1 U10463 ( .A1(n10454), .A2(n10453), .ZN(n10527) );
  NOR2_X1 U10464 ( .A1(n8051), .A2(n7667), .ZN(n10455) );
  NAND2_X1 U10465 ( .A1(n10453), .A2(n10454), .ZN(n10525) );
  NAND2_X1 U10466 ( .A1(n10528), .A2(n10529), .ZN(n10454) );
  NAND2_X1 U10467 ( .A1(n10451), .A2(n10530), .ZN(n10529) );
  OR2_X1 U10468 ( .A1(n10450), .A2(n10448), .ZN(n10530) );
  NOR2_X1 U10469 ( .A1(n7811), .A2(n7667), .ZN(n10451) );
  NAND2_X1 U10470 ( .A1(n10448), .A2(n10450), .ZN(n10528) );
  NAND2_X1 U10471 ( .A1(n10531), .A2(n10532), .ZN(n10450) );
  NAND3_X1 U10472 ( .A1(b_21_), .A2(n10533), .A3(a_12_), .ZN(n10532) );
  OR2_X1 U10473 ( .A1(n10446), .A2(n10444), .ZN(n10533) );
  NAND2_X1 U10474 ( .A1(n10444), .A2(n10446), .ZN(n10531) );
  NAND2_X1 U10475 ( .A1(n10534), .A2(n10535), .ZN(n10446) );
  NAND2_X1 U10476 ( .A1(n10443), .A2(n10536), .ZN(n10535) );
  OR2_X1 U10477 ( .A1(n10442), .A2(n10441), .ZN(n10536) );
  NOR2_X1 U10478 ( .A1(n7789), .A2(n7667), .ZN(n10443) );
  NAND2_X1 U10479 ( .A1(n10441), .A2(n10442), .ZN(n10534) );
  NAND2_X1 U10480 ( .A1(n10537), .A2(n10538), .ZN(n10442) );
  NAND3_X1 U10481 ( .A1(b_21_), .A2(n10539), .A3(a_14_), .ZN(n10538) );
  NAND2_X1 U10482 ( .A1(n10438), .A2(n10437), .ZN(n10539) );
  OR2_X1 U10483 ( .A1(n10437), .A2(n10438), .ZN(n10537) );
  AND2_X1 U10484 ( .A1(n10540), .A2(n10541), .ZN(n10438) );
  NAND2_X1 U10485 ( .A1(n10435), .A2(n10542), .ZN(n10541) );
  OR2_X1 U10486 ( .A1(n10434), .A2(n10433), .ZN(n10542) );
  NOR2_X1 U10487 ( .A1(n7754), .A2(n7667), .ZN(n10435) );
  NAND2_X1 U10488 ( .A1(n10433), .A2(n10434), .ZN(n10540) );
  NAND2_X1 U10489 ( .A1(n10543), .A2(n10544), .ZN(n10434) );
  NAND3_X1 U10490 ( .A1(b_21_), .A2(n10545), .A3(a_16_), .ZN(n10544) );
  NAND2_X1 U10491 ( .A1(n10430), .A2(n10429), .ZN(n10545) );
  OR2_X1 U10492 ( .A1(n10429), .A2(n10430), .ZN(n10543) );
  AND2_X1 U10493 ( .A1(n10546), .A2(n10547), .ZN(n10430) );
  NAND2_X1 U10494 ( .A1(n10427), .A2(n10548), .ZN(n10547) );
  OR2_X1 U10495 ( .A1(n10426), .A2(n10424), .ZN(n10548) );
  NOR2_X1 U10496 ( .A1(n7732), .A2(n7667), .ZN(n10427) );
  NAND2_X1 U10497 ( .A1(n10424), .A2(n10426), .ZN(n10546) );
  NAND2_X1 U10498 ( .A1(n10549), .A2(n10550), .ZN(n10426) );
  NAND3_X1 U10499 ( .A1(b_21_), .A2(n10551), .A3(a_18_), .ZN(n10550) );
  NAND2_X1 U10500 ( .A1(n10422), .A2(n10421), .ZN(n10551) );
  OR2_X1 U10501 ( .A1(n10421), .A2(n10422), .ZN(n10549) );
  AND2_X1 U10502 ( .A1(n10552), .A2(n10553), .ZN(n10422) );
  NAND2_X1 U10503 ( .A1(n10419), .A2(n10554), .ZN(n10553) );
  OR2_X1 U10504 ( .A1(n10418), .A2(n10416), .ZN(n10554) );
  NOR2_X1 U10505 ( .A1(n8045), .A2(n7667), .ZN(n10419) );
  NAND2_X1 U10506 ( .A1(n10416), .A2(n10418), .ZN(n10552) );
  NAND2_X1 U10507 ( .A1(n10555), .A2(n10556), .ZN(n10418) );
  NAND3_X1 U10508 ( .A1(b_21_), .A2(n10557), .A3(a_20_), .ZN(n10556) );
  NAND2_X1 U10509 ( .A1(n10414), .A2(n10413), .ZN(n10557) );
  OR2_X1 U10510 ( .A1(n10413), .A2(n10414), .ZN(n10555) );
  AND2_X1 U10511 ( .A1(n10558), .A2(n10559), .ZN(n10414) );
  NAND2_X1 U10512 ( .A1(n7662), .A2(n10560), .ZN(n10559) );
  OR2_X1 U10513 ( .A1(n10411), .A2(n10410), .ZN(n10560) );
  INV_X1 U10514 ( .A(n8015), .ZN(n7662) );
  NAND2_X1 U10515 ( .A1(a_21_), .A2(b_21_), .ZN(n8015) );
  NAND2_X1 U10516 ( .A1(n10410), .A2(n10411), .ZN(n10558) );
  NAND2_X1 U10517 ( .A1(n10561), .A2(n10562), .ZN(n10411) );
  NAND3_X1 U10518 ( .A1(a_22_), .A2(n10563), .A3(b_21_), .ZN(n10562) );
  OR2_X1 U10519 ( .A1(n10407), .A2(n10405), .ZN(n10563) );
  NAND2_X1 U10520 ( .A1(n10405), .A2(n10407), .ZN(n10561) );
  NAND2_X1 U10521 ( .A1(n10564), .A2(n10565), .ZN(n10407) );
  NAND2_X1 U10522 ( .A1(n10351), .A2(n10566), .ZN(n10565) );
  OR2_X1 U10523 ( .A1(n10350), .A2(n10348), .ZN(n10566) );
  NOR2_X1 U10524 ( .A1(n7667), .A2(n8042), .ZN(n10351) );
  NAND2_X1 U10525 ( .A1(n10348), .A2(n10350), .ZN(n10564) );
  NAND2_X1 U10526 ( .A1(n10567), .A2(n10568), .ZN(n10350) );
  NAND3_X1 U10527 ( .A1(a_24_), .A2(n10569), .A3(b_21_), .ZN(n10568) );
  NAND2_X1 U10528 ( .A1(n10403), .A2(n10402), .ZN(n10569) );
  OR2_X1 U10529 ( .A1(n10402), .A2(n10403), .ZN(n10567) );
  AND2_X1 U10530 ( .A1(n10570), .A2(n10571), .ZN(n10403) );
  NAND2_X1 U10531 ( .A1(n10400), .A2(n10572), .ZN(n10571) );
  OR2_X1 U10532 ( .A1(n10399), .A2(n10398), .ZN(n10572) );
  NOR2_X1 U10533 ( .A1(n7667), .A2(n8039), .ZN(n10400) );
  NAND2_X1 U10534 ( .A1(n10398), .A2(n10399), .ZN(n10570) );
  NAND2_X1 U10535 ( .A1(n10395), .A2(n10573), .ZN(n10399) );
  NAND2_X1 U10536 ( .A1(n10394), .A2(n10396), .ZN(n10573) );
  NAND2_X1 U10537 ( .A1(n10574), .A2(n10575), .ZN(n10396) );
  NAND2_X1 U10538 ( .A1(b_21_), .A2(a_26_), .ZN(n10575) );
  INV_X1 U10539 ( .A(n10576), .ZN(n10574) );
  XNOR2_X1 U10540 ( .A(n10577), .B(n10578), .ZN(n10394) );
  NAND2_X1 U10541 ( .A1(n10579), .A2(n10580), .ZN(n10577) );
  NAND2_X1 U10542 ( .A1(a_26_), .A2(n10576), .ZN(n10395) );
  NAND2_X1 U10543 ( .A1(n10367), .A2(n10581), .ZN(n10576) );
  NAND2_X1 U10544 ( .A1(n10366), .A2(n10368), .ZN(n10581) );
  NAND2_X1 U10545 ( .A1(n10582), .A2(n10583), .ZN(n10368) );
  NAND2_X1 U10546 ( .A1(b_21_), .A2(a_27_), .ZN(n10583) );
  INV_X1 U10547 ( .A(n10584), .ZN(n10582) );
  XNOR2_X1 U10548 ( .A(n10585), .B(n10586), .ZN(n10366) );
  XOR2_X1 U10549 ( .A(n10587), .B(n10588), .Z(n10585) );
  NAND2_X1 U10550 ( .A1(b_20_), .A2(a_28_), .ZN(n10587) );
  NAND2_X1 U10551 ( .A1(a_27_), .A2(n10584), .ZN(n10367) );
  NAND2_X1 U10552 ( .A1(n10589), .A2(n10590), .ZN(n10584) );
  NAND3_X1 U10553 ( .A1(a_28_), .A2(n10591), .A3(b_21_), .ZN(n10590) );
  NAND2_X1 U10554 ( .A1(n10376), .A2(n10374), .ZN(n10591) );
  OR2_X1 U10555 ( .A1(n10374), .A2(n10376), .ZN(n10589) );
  AND2_X1 U10556 ( .A1(n10592), .A2(n10593), .ZN(n10376) );
  NAND2_X1 U10557 ( .A1(n10390), .A2(n10594), .ZN(n10593) );
  OR2_X1 U10558 ( .A1(n10391), .A2(n10392), .ZN(n10594) );
  NOR2_X1 U10559 ( .A1(n7667), .A2(n7545), .ZN(n10390) );
  NAND2_X1 U10560 ( .A1(n10392), .A2(n10391), .ZN(n10592) );
  NAND2_X1 U10561 ( .A1(n10595), .A2(n10596), .ZN(n10391) );
  NAND2_X1 U10562 ( .A1(b_19_), .A2(n10597), .ZN(n10596) );
  NAND2_X1 U10563 ( .A1(n7527), .A2(n10598), .ZN(n10597) );
  NAND2_X1 U10564 ( .A1(a_31_), .A2(n8043), .ZN(n10598) );
  NAND2_X1 U10565 ( .A1(b_20_), .A2(n10599), .ZN(n10595) );
  NAND2_X1 U10566 ( .A1(n7531), .A2(n10600), .ZN(n10599) );
  NAND2_X1 U10567 ( .A1(a_30_), .A2(n7693), .ZN(n10600) );
  AND3_X1 U10568 ( .A1(b_20_), .A2(b_21_), .A3(n7494), .ZN(n10392) );
  XNOR2_X1 U10569 ( .A(n10601), .B(n10602), .ZN(n10374) );
  XOR2_X1 U10570 ( .A(n10603), .B(n10604), .Z(n10601) );
  XNOR2_X1 U10571 ( .A(n10605), .B(n10606), .ZN(n10398) );
  NAND2_X1 U10572 ( .A1(n10607), .A2(n10608), .ZN(n10605) );
  XNOR2_X1 U10573 ( .A(n10609), .B(n10610), .ZN(n10402) );
  XOR2_X1 U10574 ( .A(n10611), .B(n10612), .Z(n10609) );
  XNOR2_X1 U10575 ( .A(n10613), .B(n10614), .ZN(n10348) );
  XNOR2_X1 U10576 ( .A(n10615), .B(n10616), .ZN(n10613) );
  NOR2_X1 U10577 ( .A1(n8041), .A2(n8043), .ZN(n10616) );
  XNOR2_X1 U10578 ( .A(n10617), .B(n10618), .ZN(n10405) );
  XNOR2_X1 U10579 ( .A(n10619), .B(n10620), .ZN(n10618) );
  XNOR2_X1 U10580 ( .A(n10621), .B(n10622), .ZN(n10410) );
  XOR2_X1 U10581 ( .A(n10623), .B(n10624), .Z(n10622) );
  NAND2_X1 U10582 ( .A1(b_20_), .A2(a_22_), .ZN(n10624) );
  XNOR2_X1 U10583 ( .A(n10625), .B(n10626), .ZN(n10413) );
  XOR2_X1 U10584 ( .A(n10627), .B(n10628), .Z(n10625) );
  XOR2_X1 U10585 ( .A(n10629), .B(n10630), .Z(n10416) );
  XOR2_X1 U10586 ( .A(n10631), .B(n10632), .Z(n10629) );
  XNOR2_X1 U10587 ( .A(n10633), .B(n10634), .ZN(n10421) );
  XOR2_X1 U10588 ( .A(n10635), .B(n10636), .Z(n10633) );
  XNOR2_X1 U10589 ( .A(n10637), .B(n10638), .ZN(n10424) );
  XNOR2_X1 U10590 ( .A(n10639), .B(n10640), .ZN(n10637) );
  NOR2_X1 U10591 ( .A1(n8043), .A2(n8047), .ZN(n10640) );
  XOR2_X1 U10592 ( .A(n10641), .B(n10642), .Z(n10429) );
  XNOR2_X1 U10593 ( .A(n10643), .B(n10644), .ZN(n10642) );
  XNOR2_X1 U10594 ( .A(n10645), .B(n10646), .ZN(n10433) );
  XNOR2_X1 U10595 ( .A(n10647), .B(n10648), .ZN(n10645) );
  NOR2_X1 U10596 ( .A1(n8043), .A2(n8438), .ZN(n10648) );
  XOR2_X1 U10597 ( .A(n10649), .B(n10650), .Z(n10437) );
  XNOR2_X1 U10598 ( .A(n10651), .B(n10652), .ZN(n10650) );
  XNOR2_X1 U10599 ( .A(n10653), .B(n10654), .ZN(n10441) );
  XNOR2_X1 U10600 ( .A(n10655), .B(n10656), .ZN(n10653) );
  NOR2_X1 U10601 ( .A1(n8043), .A2(n8049), .ZN(n10656) );
  XNOR2_X1 U10602 ( .A(n10657), .B(n10658), .ZN(n10444) );
  XNOR2_X1 U10603 ( .A(n10659), .B(n10660), .ZN(n10658) );
  XNOR2_X1 U10604 ( .A(n10661), .B(n10662), .ZN(n10448) );
  XOR2_X1 U10605 ( .A(n10663), .B(n10664), .Z(n10662) );
  NAND2_X1 U10606 ( .A1(a_12_), .A2(b_20_), .ZN(n10664) );
  XNOR2_X1 U10607 ( .A(n10665), .B(n10666), .ZN(n10453) );
  XOR2_X1 U10608 ( .A(n10667), .B(n10668), .Z(n10666) );
  NAND2_X1 U10609 ( .A1(a_11_), .A2(b_20_), .ZN(n10668) );
  XNOR2_X1 U10610 ( .A(n10669), .B(n10670), .ZN(n10457) );
  XNOR2_X1 U10611 ( .A(n10671), .B(n10672), .ZN(n10669) );
  XOR2_X1 U10612 ( .A(n10673), .B(n10674), .Z(n10460) );
  XOR2_X1 U10613 ( .A(n10675), .B(n10676), .Z(n10673) );
  XNOR2_X1 U10614 ( .A(n10677), .B(n10678), .ZN(n10464) );
  XNOR2_X1 U10615 ( .A(n10679), .B(n10680), .ZN(n10677) );
  NOR2_X1 U10616 ( .A1(n8043), .A2(n8686), .ZN(n10680) );
  XOR2_X1 U10617 ( .A(n10681), .B(n10682), .Z(n10469) );
  NAND2_X1 U10618 ( .A1(n10683), .A2(n10684), .ZN(n10681) );
  XOR2_X1 U10619 ( .A(n10685), .B(n10686), .Z(n10473) );
  NAND2_X1 U10620 ( .A1(n10687), .A2(n10688), .ZN(n10685) );
  XOR2_X1 U10621 ( .A(n10689), .B(n10690), .Z(n10477) );
  XNOR2_X1 U10622 ( .A(n10691), .B(n10692), .ZN(n10690) );
  XNOR2_X1 U10623 ( .A(n10693), .B(n10694), .ZN(n10480) );
  XOR2_X1 U10624 ( .A(n10695), .B(n10696), .Z(n10694) );
  NAND2_X1 U10625 ( .A1(a_4_), .A2(b_20_), .ZN(n10696) );
  XNOR2_X1 U10626 ( .A(n10697), .B(n10698), .ZN(n10484) );
  NAND2_X1 U10627 ( .A1(n10699), .A2(n10700), .ZN(n10697) );
  XNOR2_X1 U10628 ( .A(n10701), .B(n10702), .ZN(n10279) );
  NAND2_X1 U10629 ( .A1(n10703), .A2(n10704), .ZN(n10701) );
  XNOR2_X1 U10630 ( .A(n10705), .B(n10706), .ZN(n10490) );
  XNOR2_X1 U10631 ( .A(n10707), .B(n10708), .ZN(n10705) );
  XNOR2_X1 U10632 ( .A(n10709), .B(n10710), .ZN(n10489) );
  XOR2_X1 U10633 ( .A(n10711), .B(n10712), .Z(n10709) );
  NOR2_X1 U10634 ( .A1(n8043), .A2(n8942), .ZN(n10712) );
  XOR2_X1 U10635 ( .A(n8231), .B(n8230), .Z(n10494) );
  NAND3_X1 U10636 ( .A1(n8230), .A2(n8231), .A3(n10713), .ZN(n8126) );
  XOR2_X1 U10637 ( .A(n8224), .B(n8223), .Z(n10713) );
  NAND2_X1 U10638 ( .A1(n10714), .A2(n10715), .ZN(n8231) );
  NAND3_X1 U10639 ( .A1(b_20_), .A2(n10716), .A3(a_0_), .ZN(n10715) );
  OR2_X1 U10640 ( .A1(n10711), .A2(n10710), .ZN(n10716) );
  NAND2_X1 U10641 ( .A1(n10710), .A2(n10711), .ZN(n10714) );
  NAND2_X1 U10642 ( .A1(n10717), .A2(n10718), .ZN(n10711) );
  NAND2_X1 U10643 ( .A1(n10708), .A2(n10719), .ZN(n10718) );
  NAND2_X1 U10644 ( .A1(n10707), .A2(n10706), .ZN(n10719) );
  NOR2_X1 U10645 ( .A1(n8043), .A2(n7957), .ZN(n10708) );
  OR2_X1 U10646 ( .A1(n10706), .A2(n10707), .ZN(n10717) );
  AND2_X1 U10647 ( .A1(n10703), .A2(n10720), .ZN(n10707) );
  NAND2_X1 U10648 ( .A1(n10702), .A2(n10704), .ZN(n10720) );
  NAND2_X1 U10649 ( .A1(n10721), .A2(n10722), .ZN(n10704) );
  NAND2_X1 U10650 ( .A1(a_2_), .A2(b_20_), .ZN(n10722) );
  INV_X1 U10651 ( .A(n10723), .ZN(n10721) );
  XNOR2_X1 U10652 ( .A(n10724), .B(n10725), .ZN(n10702) );
  XOR2_X1 U10653 ( .A(n10726), .B(n10727), .Z(n10725) );
  NAND2_X1 U10654 ( .A1(a_3_), .A2(b_19_), .ZN(n10727) );
  NAND2_X1 U10655 ( .A1(a_2_), .A2(n10723), .ZN(n10703) );
  NAND2_X1 U10656 ( .A1(n10699), .A2(n10728), .ZN(n10723) );
  NAND2_X1 U10657 ( .A1(n10698), .A2(n10700), .ZN(n10728) );
  NAND2_X1 U10658 ( .A1(n10729), .A2(n10730), .ZN(n10700) );
  NAND2_X1 U10659 ( .A1(a_3_), .A2(b_20_), .ZN(n10730) );
  INV_X1 U10660 ( .A(n10731), .ZN(n10729) );
  XOR2_X1 U10661 ( .A(n10732), .B(n10733), .Z(n10698) );
  XOR2_X1 U10662 ( .A(n10734), .B(n10735), .Z(n10732) );
  NOR2_X1 U10663 ( .A1(n7693), .A2(n7916), .ZN(n10735) );
  NAND2_X1 U10664 ( .A1(a_3_), .A2(n10731), .ZN(n10699) );
  NAND2_X1 U10665 ( .A1(n10736), .A2(n10737), .ZN(n10731) );
  NAND3_X1 U10666 ( .A1(b_20_), .A2(n10738), .A3(a_4_), .ZN(n10737) );
  OR2_X1 U10667 ( .A1(n10695), .A2(n10693), .ZN(n10738) );
  NAND2_X1 U10668 ( .A1(n10693), .A2(n10695), .ZN(n10736) );
  NAND2_X1 U10669 ( .A1(n10739), .A2(n10740), .ZN(n10695) );
  NAND2_X1 U10670 ( .A1(n10692), .A2(n10741), .ZN(n10740) );
  OR2_X1 U10671 ( .A1(n10691), .A2(n10689), .ZN(n10741) );
  NOR2_X1 U10672 ( .A1(n7908), .A2(n8043), .ZN(n10692) );
  NAND2_X1 U10673 ( .A1(n10689), .A2(n10691), .ZN(n10739) );
  NAND2_X1 U10674 ( .A1(n10687), .A2(n10742), .ZN(n10691) );
  NAND2_X1 U10675 ( .A1(n10686), .A2(n10688), .ZN(n10742) );
  NAND2_X1 U10676 ( .A1(n10743), .A2(n10744), .ZN(n10688) );
  NAND2_X1 U10677 ( .A1(a_6_), .A2(b_20_), .ZN(n10744) );
  INV_X1 U10678 ( .A(n10745), .ZN(n10743) );
  XNOR2_X1 U10679 ( .A(n10746), .B(n10747), .ZN(n10686) );
  XOR2_X1 U10680 ( .A(n10748), .B(n10749), .Z(n10747) );
  NAND2_X1 U10681 ( .A1(a_7_), .A2(b_19_), .ZN(n10749) );
  NAND2_X1 U10682 ( .A1(a_6_), .A2(n10745), .ZN(n10687) );
  NAND2_X1 U10683 ( .A1(n10683), .A2(n10750), .ZN(n10745) );
  NAND2_X1 U10684 ( .A1(n10682), .A2(n10684), .ZN(n10750) );
  NAND2_X1 U10685 ( .A1(n10751), .A2(n10752), .ZN(n10684) );
  NAND2_X1 U10686 ( .A1(a_7_), .A2(b_20_), .ZN(n10752) );
  INV_X1 U10687 ( .A(n10753), .ZN(n10751) );
  XOR2_X1 U10688 ( .A(n10754), .B(n10755), .Z(n10682) );
  XOR2_X1 U10689 ( .A(n10756), .B(n10757), .Z(n10754) );
  NOR2_X1 U10690 ( .A1(n7693), .A2(n8686), .ZN(n10757) );
  NAND2_X1 U10691 ( .A1(a_7_), .A2(n10753), .ZN(n10683) );
  NAND2_X1 U10692 ( .A1(n10758), .A2(n10759), .ZN(n10753) );
  NAND3_X1 U10693 ( .A1(b_20_), .A2(n10760), .A3(a_8_), .ZN(n10759) );
  NAND2_X1 U10694 ( .A1(n10679), .A2(n10678), .ZN(n10760) );
  OR2_X1 U10695 ( .A1(n10678), .A2(n10679), .ZN(n10758) );
  AND2_X1 U10696 ( .A1(n10761), .A2(n10762), .ZN(n10679) );
  NAND2_X1 U10697 ( .A1(n10675), .A2(n10763), .ZN(n10762) );
  OR2_X1 U10698 ( .A1(n10676), .A2(n10674), .ZN(n10763) );
  NOR2_X1 U10699 ( .A1(n8052), .A2(n8043), .ZN(n10675) );
  NAND2_X1 U10700 ( .A1(n10674), .A2(n10676), .ZN(n10761) );
  NAND2_X1 U10701 ( .A1(n10764), .A2(n10765), .ZN(n10676) );
  NAND2_X1 U10702 ( .A1(n10672), .A2(n10766), .ZN(n10765) );
  NAND2_X1 U10703 ( .A1(n10671), .A2(n10670), .ZN(n10766) );
  NOR2_X1 U10704 ( .A1(n8051), .A2(n8043), .ZN(n10672) );
  OR2_X1 U10705 ( .A1(n10670), .A2(n10671), .ZN(n10764) );
  AND2_X1 U10706 ( .A1(n10767), .A2(n10768), .ZN(n10671) );
  NAND3_X1 U10707 ( .A1(b_20_), .A2(n10769), .A3(a_11_), .ZN(n10768) );
  OR2_X1 U10708 ( .A1(n10667), .A2(n10665), .ZN(n10769) );
  NAND2_X1 U10709 ( .A1(n10665), .A2(n10667), .ZN(n10767) );
  NAND2_X1 U10710 ( .A1(n10770), .A2(n10771), .ZN(n10667) );
  NAND3_X1 U10711 ( .A1(b_20_), .A2(n10772), .A3(a_12_), .ZN(n10771) );
  OR2_X1 U10712 ( .A1(n10663), .A2(n10661), .ZN(n10772) );
  NAND2_X1 U10713 ( .A1(n10661), .A2(n10663), .ZN(n10770) );
  NAND2_X1 U10714 ( .A1(n10773), .A2(n10774), .ZN(n10663) );
  NAND2_X1 U10715 ( .A1(n10660), .A2(n10775), .ZN(n10774) );
  OR2_X1 U10716 ( .A1(n10659), .A2(n10657), .ZN(n10775) );
  NOR2_X1 U10717 ( .A1(n7789), .A2(n8043), .ZN(n10660) );
  NAND2_X1 U10718 ( .A1(n10657), .A2(n10659), .ZN(n10773) );
  NAND2_X1 U10719 ( .A1(n10776), .A2(n10777), .ZN(n10659) );
  NAND3_X1 U10720 ( .A1(b_20_), .A2(n10778), .A3(a_14_), .ZN(n10777) );
  NAND2_X1 U10721 ( .A1(n10655), .A2(n10654), .ZN(n10778) );
  OR2_X1 U10722 ( .A1(n10654), .A2(n10655), .ZN(n10776) );
  AND2_X1 U10723 ( .A1(n10779), .A2(n10780), .ZN(n10655) );
  NAND2_X1 U10724 ( .A1(n10652), .A2(n10781), .ZN(n10780) );
  OR2_X1 U10725 ( .A1(n10651), .A2(n10649), .ZN(n10781) );
  NOR2_X1 U10726 ( .A1(n7754), .A2(n8043), .ZN(n10652) );
  NAND2_X1 U10727 ( .A1(n10649), .A2(n10651), .ZN(n10779) );
  NAND2_X1 U10728 ( .A1(n10782), .A2(n10783), .ZN(n10651) );
  NAND3_X1 U10729 ( .A1(b_20_), .A2(n10784), .A3(a_16_), .ZN(n10783) );
  NAND2_X1 U10730 ( .A1(n10647), .A2(n10646), .ZN(n10784) );
  OR2_X1 U10731 ( .A1(n10646), .A2(n10647), .ZN(n10782) );
  AND2_X1 U10732 ( .A1(n10785), .A2(n10786), .ZN(n10647) );
  NAND2_X1 U10733 ( .A1(n10644), .A2(n10787), .ZN(n10786) );
  OR2_X1 U10734 ( .A1(n10643), .A2(n10641), .ZN(n10787) );
  NOR2_X1 U10735 ( .A1(n7732), .A2(n8043), .ZN(n10644) );
  NAND2_X1 U10736 ( .A1(n10641), .A2(n10643), .ZN(n10785) );
  NAND2_X1 U10737 ( .A1(n10788), .A2(n10789), .ZN(n10643) );
  NAND3_X1 U10738 ( .A1(b_20_), .A2(n10790), .A3(a_18_), .ZN(n10789) );
  NAND2_X1 U10739 ( .A1(n10639), .A2(n10638), .ZN(n10790) );
  OR2_X1 U10740 ( .A1(n10638), .A2(n10639), .ZN(n10788) );
  AND2_X1 U10741 ( .A1(n10791), .A2(n10792), .ZN(n10639) );
  NAND2_X1 U10742 ( .A1(n10636), .A2(n10793), .ZN(n10792) );
  OR2_X1 U10743 ( .A1(n10635), .A2(n10634), .ZN(n10793) );
  NOR2_X1 U10744 ( .A1(n8045), .A2(n8043), .ZN(n10636) );
  NAND2_X1 U10745 ( .A1(n10634), .A2(n10635), .ZN(n10791) );
  NAND2_X1 U10746 ( .A1(n10794), .A2(n10795), .ZN(n10635) );
  NAND2_X1 U10747 ( .A1(n10630), .A2(n10796), .ZN(n10795) );
  OR2_X1 U10748 ( .A1(n10631), .A2(n10632), .ZN(n10796) );
  XNOR2_X1 U10749 ( .A(n10797), .B(n10798), .ZN(n10630) );
  XNOR2_X1 U10750 ( .A(n10799), .B(n10800), .ZN(n10797) );
  NAND2_X1 U10751 ( .A1(n10632), .A2(n10631), .ZN(n10794) );
  NAND2_X1 U10752 ( .A1(n10801), .A2(n10802), .ZN(n10631) );
  NAND2_X1 U10753 ( .A1(n10628), .A2(n10803), .ZN(n10802) );
  OR2_X1 U10754 ( .A1(n10627), .A2(n10626), .ZN(n10803) );
  NOR2_X1 U10755 ( .A1(n8043), .A2(n7665), .ZN(n10628) );
  NAND2_X1 U10756 ( .A1(n10626), .A2(n10627), .ZN(n10801) );
  NAND2_X1 U10757 ( .A1(n10804), .A2(n10805), .ZN(n10627) );
  NAND3_X1 U10758 ( .A1(a_22_), .A2(n10806), .A3(b_20_), .ZN(n10805) );
  OR2_X1 U10759 ( .A1(n10623), .A2(n10621), .ZN(n10806) );
  NAND2_X1 U10760 ( .A1(n10621), .A2(n10623), .ZN(n10804) );
  NAND2_X1 U10761 ( .A1(n10807), .A2(n10808), .ZN(n10623) );
  NAND2_X1 U10762 ( .A1(n10620), .A2(n10809), .ZN(n10808) );
  OR2_X1 U10763 ( .A1(n10619), .A2(n10617), .ZN(n10809) );
  NOR2_X1 U10764 ( .A1(n8043), .A2(n8042), .ZN(n10620) );
  NAND2_X1 U10765 ( .A1(n10617), .A2(n10619), .ZN(n10807) );
  NAND2_X1 U10766 ( .A1(n10810), .A2(n10811), .ZN(n10619) );
  NAND3_X1 U10767 ( .A1(a_24_), .A2(n10812), .A3(b_20_), .ZN(n10811) );
  NAND2_X1 U10768 ( .A1(n10615), .A2(n10614), .ZN(n10812) );
  OR2_X1 U10769 ( .A1(n10614), .A2(n10615), .ZN(n10810) );
  AND2_X1 U10770 ( .A1(n10813), .A2(n10814), .ZN(n10615) );
  NAND2_X1 U10771 ( .A1(n10612), .A2(n10815), .ZN(n10814) );
  OR2_X1 U10772 ( .A1(n10611), .A2(n10610), .ZN(n10815) );
  NOR2_X1 U10773 ( .A1(n8043), .A2(n8039), .ZN(n10612) );
  NAND2_X1 U10774 ( .A1(n10610), .A2(n10611), .ZN(n10813) );
  NAND2_X1 U10775 ( .A1(n10607), .A2(n10816), .ZN(n10611) );
  NAND2_X1 U10776 ( .A1(n10606), .A2(n10608), .ZN(n10816) );
  NAND2_X1 U10777 ( .A1(n10817), .A2(n10818), .ZN(n10608) );
  NAND2_X1 U10778 ( .A1(b_20_), .A2(a_26_), .ZN(n10818) );
  INV_X1 U10779 ( .A(n10819), .ZN(n10817) );
  XNOR2_X1 U10780 ( .A(n10820), .B(n10821), .ZN(n10606) );
  NAND2_X1 U10781 ( .A1(n10822), .A2(n10823), .ZN(n10820) );
  NAND2_X1 U10782 ( .A1(a_26_), .A2(n10819), .ZN(n10607) );
  NAND2_X1 U10783 ( .A1(n10579), .A2(n10824), .ZN(n10819) );
  NAND2_X1 U10784 ( .A1(n10578), .A2(n10580), .ZN(n10824) );
  NAND2_X1 U10785 ( .A1(n10825), .A2(n10826), .ZN(n10580) );
  NAND2_X1 U10786 ( .A1(b_20_), .A2(a_27_), .ZN(n10826) );
  INV_X1 U10787 ( .A(n10827), .ZN(n10825) );
  XNOR2_X1 U10788 ( .A(n10828), .B(n10829), .ZN(n10578) );
  XOR2_X1 U10789 ( .A(n10830), .B(n10831), .Z(n10828) );
  NAND2_X1 U10790 ( .A1(b_19_), .A2(a_28_), .ZN(n10830) );
  NAND2_X1 U10791 ( .A1(a_27_), .A2(n10827), .ZN(n10579) );
  NAND2_X1 U10792 ( .A1(n10832), .A2(n10833), .ZN(n10827) );
  NAND3_X1 U10793 ( .A1(a_28_), .A2(n10834), .A3(b_20_), .ZN(n10833) );
  NAND2_X1 U10794 ( .A1(n10588), .A2(n10586), .ZN(n10834) );
  OR2_X1 U10795 ( .A1(n10586), .A2(n10588), .ZN(n10832) );
  AND2_X1 U10796 ( .A1(n10835), .A2(n10836), .ZN(n10588) );
  NAND2_X1 U10797 ( .A1(n10602), .A2(n10837), .ZN(n10836) );
  OR2_X1 U10798 ( .A1(n10603), .A2(n10604), .ZN(n10837) );
  NOR2_X1 U10799 ( .A1(n8043), .A2(n7545), .ZN(n10602) );
  NAND2_X1 U10800 ( .A1(n10604), .A2(n10603), .ZN(n10835) );
  NAND2_X1 U10801 ( .A1(n10838), .A2(n10839), .ZN(n10603) );
  NAND2_X1 U10802 ( .A1(b_18_), .A2(n10840), .ZN(n10839) );
  NAND2_X1 U10803 ( .A1(n7527), .A2(n10841), .ZN(n10840) );
  NAND2_X1 U10804 ( .A1(a_31_), .A2(n7693), .ZN(n10841) );
  NAND2_X1 U10805 ( .A1(b_19_), .A2(n10842), .ZN(n10838) );
  NAND2_X1 U10806 ( .A1(n7531), .A2(n10843), .ZN(n10842) );
  NAND2_X1 U10807 ( .A1(a_30_), .A2(n8046), .ZN(n10843) );
  AND3_X1 U10808 ( .A1(b_20_), .A2(b_19_), .A3(n7494), .ZN(n10604) );
  XNOR2_X1 U10809 ( .A(n10844), .B(n10845), .ZN(n10586) );
  XOR2_X1 U10810 ( .A(n10846), .B(n10847), .Z(n10844) );
  XNOR2_X1 U10811 ( .A(n10848), .B(n10849), .ZN(n10610) );
  NAND2_X1 U10812 ( .A1(n10850), .A2(n10851), .ZN(n10848) );
  XNOR2_X1 U10813 ( .A(n10852), .B(n10853), .ZN(n10614) );
  XOR2_X1 U10814 ( .A(n10854), .B(n10855), .Z(n10852) );
  XNOR2_X1 U10815 ( .A(n10856), .B(n10857), .ZN(n10617) );
  XNOR2_X1 U10816 ( .A(n10858), .B(n10859), .ZN(n10856) );
  NOR2_X1 U10817 ( .A1(n8041), .A2(n7693), .ZN(n10859) );
  XNOR2_X1 U10818 ( .A(n10860), .B(n10861), .ZN(n10621) );
  XNOR2_X1 U10819 ( .A(n10862), .B(n10863), .ZN(n10861) );
  XNOR2_X1 U10820 ( .A(n10864), .B(n10865), .ZN(n10626) );
  XOR2_X1 U10821 ( .A(n10866), .B(n10867), .Z(n10865) );
  NAND2_X1 U10822 ( .A1(b_19_), .A2(a_22_), .ZN(n10867) );
  INV_X1 U10823 ( .A(n7684), .ZN(n10632) );
  NAND2_X1 U10824 ( .A1(b_20_), .A2(a_20_), .ZN(n7684) );
  XNOR2_X1 U10825 ( .A(n10868), .B(n10869), .ZN(n10634) );
  XOR2_X1 U10826 ( .A(n10870), .B(n10871), .Z(n10868) );
  NAND2_X1 U10827 ( .A1(b_19_), .A2(a_20_), .ZN(n10870) );
  XNOR2_X1 U10828 ( .A(n10872), .B(n10873), .ZN(n10638) );
  XOR2_X1 U10829 ( .A(n10874), .B(n7691), .Z(n10872) );
  XNOR2_X1 U10830 ( .A(n10875), .B(n10876), .ZN(n10641) );
  XNOR2_X1 U10831 ( .A(n10877), .B(n10878), .ZN(n10875) );
  NOR2_X1 U10832 ( .A1(n7693), .A2(n8047), .ZN(n10878) );
  XNOR2_X1 U10833 ( .A(n10879), .B(n10880), .ZN(n10646) );
  XOR2_X1 U10834 ( .A(n10881), .B(n10882), .Z(n10879) );
  XNOR2_X1 U10835 ( .A(n10883), .B(n10884), .ZN(n10649) );
  XOR2_X1 U10836 ( .A(n10885), .B(n10886), .Z(n10884) );
  NAND2_X1 U10837 ( .A1(a_16_), .A2(b_19_), .ZN(n10886) );
  XOR2_X1 U10838 ( .A(n10887), .B(n10888), .Z(n10654) );
  XNOR2_X1 U10839 ( .A(n10889), .B(n10890), .ZN(n10888) );
  XNOR2_X1 U10840 ( .A(n10891), .B(n10892), .ZN(n10657) );
  XNOR2_X1 U10841 ( .A(n10893), .B(n10894), .ZN(n10891) );
  NOR2_X1 U10842 ( .A1(n7693), .A2(n8049), .ZN(n10894) );
  XOR2_X1 U10843 ( .A(n10895), .B(n10896), .Z(n10661) );
  XOR2_X1 U10844 ( .A(n10897), .B(n10898), .Z(n10895) );
  XNOR2_X1 U10845 ( .A(n10899), .B(n10900), .ZN(n10665) );
  XOR2_X1 U10846 ( .A(n10901), .B(n10902), .Z(n10900) );
  NAND2_X1 U10847 ( .A1(a_12_), .A2(b_19_), .ZN(n10902) );
  XOR2_X1 U10848 ( .A(n10903), .B(n10904), .Z(n10670) );
  NAND2_X1 U10849 ( .A1(n10905), .A2(n10906), .ZN(n10903) );
  XNOR2_X1 U10850 ( .A(n10907), .B(n10908), .ZN(n10674) );
  NAND2_X1 U10851 ( .A1(n10909), .A2(n10910), .ZN(n10907) );
  XNOR2_X1 U10852 ( .A(n10911), .B(n10912), .ZN(n10678) );
  XOR2_X1 U10853 ( .A(n10913), .B(n10914), .Z(n10911) );
  NOR2_X1 U10854 ( .A1(n7693), .A2(n8052), .ZN(n10914) );
  XNOR2_X1 U10855 ( .A(n10915), .B(n10916), .ZN(n10689) );
  XNOR2_X1 U10856 ( .A(n10917), .B(n10918), .ZN(n10915) );
  NOR2_X1 U10857 ( .A1(n7693), .A2(n7887), .ZN(n10918) );
  XNOR2_X1 U10858 ( .A(n10919), .B(n10920), .ZN(n10693) );
  XOR2_X1 U10859 ( .A(n10921), .B(n10922), .Z(n10920) );
  NAND2_X1 U10860 ( .A1(a_5_), .A2(b_19_), .ZN(n10922) );
  XOR2_X1 U10861 ( .A(n10923), .B(n10924), .Z(n10706) );
  XOR2_X1 U10862 ( .A(n10925), .B(n10926), .Z(n10924) );
  NAND2_X1 U10863 ( .A1(a_2_), .A2(b_19_), .ZN(n10926) );
  XNOR2_X1 U10864 ( .A(n10927), .B(n10928), .ZN(n10710) );
  XOR2_X1 U10865 ( .A(n10929), .B(n10930), .Z(n10928) );
  NAND2_X1 U10866 ( .A1(b_19_), .A2(a_1_), .ZN(n10930) );
  XNOR2_X1 U10867 ( .A(n10931), .B(n10932), .ZN(n8230) );
  XOR2_X1 U10868 ( .A(n10933), .B(n10934), .Z(n10932) );
  NAND2_X1 U10869 ( .A1(a_0_), .A2(b_19_), .ZN(n10934) );
  NAND3_X1 U10870 ( .A1(n10935), .A2(n8224), .A3(n8223), .ZN(n8131) );
  XOR2_X1 U10871 ( .A(n10936), .B(n10937), .Z(n8223) );
  XOR2_X1 U10872 ( .A(n10938), .B(n10939), .Z(n10936) );
  NOR2_X1 U10873 ( .A1(n8046), .A2(n8942), .ZN(n10939) );
  NAND2_X1 U10874 ( .A1(n10940), .A2(n10941), .ZN(n8224) );
  NAND3_X1 U10875 ( .A1(b_19_), .A2(n10942), .A3(a_0_), .ZN(n10941) );
  OR2_X1 U10876 ( .A1(n10933), .A2(n10931), .ZN(n10942) );
  NAND2_X1 U10877 ( .A1(n10931), .A2(n10933), .ZN(n10940) );
  NAND2_X1 U10878 ( .A1(n10943), .A2(n10944), .ZN(n10933) );
  NAND3_X1 U10879 ( .A1(a_1_), .A2(n10945), .A3(b_19_), .ZN(n10944) );
  OR2_X1 U10880 ( .A1(n10929), .A2(n10927), .ZN(n10945) );
  NAND2_X1 U10881 ( .A1(n10927), .A2(n10929), .ZN(n10943) );
  NAND2_X1 U10882 ( .A1(n10946), .A2(n10947), .ZN(n10929) );
  NAND3_X1 U10883 ( .A1(b_19_), .A2(n10948), .A3(a_2_), .ZN(n10947) );
  OR2_X1 U10884 ( .A1(n10925), .A2(n10923), .ZN(n10948) );
  NAND2_X1 U10885 ( .A1(n10923), .A2(n10925), .ZN(n10946) );
  NAND2_X1 U10886 ( .A1(n10949), .A2(n10950), .ZN(n10925) );
  NAND3_X1 U10887 ( .A1(b_19_), .A2(n10951), .A3(a_3_), .ZN(n10950) );
  OR2_X1 U10888 ( .A1(n10726), .A2(n10724), .ZN(n10951) );
  NAND2_X1 U10889 ( .A1(n10724), .A2(n10726), .ZN(n10949) );
  NAND2_X1 U10890 ( .A1(n10952), .A2(n10953), .ZN(n10726) );
  NAND3_X1 U10891 ( .A1(b_19_), .A2(n10954), .A3(a_4_), .ZN(n10953) );
  OR2_X1 U10892 ( .A1(n10734), .A2(n10733), .ZN(n10954) );
  NAND2_X1 U10893 ( .A1(n10733), .A2(n10734), .ZN(n10952) );
  NAND2_X1 U10894 ( .A1(n10955), .A2(n10956), .ZN(n10734) );
  NAND3_X1 U10895 ( .A1(b_19_), .A2(n10957), .A3(a_5_), .ZN(n10956) );
  OR2_X1 U10896 ( .A1(n10921), .A2(n10919), .ZN(n10957) );
  NAND2_X1 U10897 ( .A1(n10919), .A2(n10921), .ZN(n10955) );
  NAND2_X1 U10898 ( .A1(n10958), .A2(n10959), .ZN(n10921) );
  NAND3_X1 U10899 ( .A1(b_19_), .A2(n10960), .A3(a_6_), .ZN(n10959) );
  NAND2_X1 U10900 ( .A1(n10917), .A2(n10916), .ZN(n10960) );
  OR2_X1 U10901 ( .A1(n10916), .A2(n10917), .ZN(n10958) );
  AND2_X1 U10902 ( .A1(n10961), .A2(n10962), .ZN(n10917) );
  NAND3_X1 U10903 ( .A1(b_19_), .A2(n10963), .A3(a_7_), .ZN(n10962) );
  OR2_X1 U10904 ( .A1(n10748), .A2(n10746), .ZN(n10963) );
  NAND2_X1 U10905 ( .A1(n10746), .A2(n10748), .ZN(n10961) );
  NAND2_X1 U10906 ( .A1(n10964), .A2(n10965), .ZN(n10748) );
  NAND3_X1 U10907 ( .A1(b_19_), .A2(n10966), .A3(a_8_), .ZN(n10965) );
  OR2_X1 U10908 ( .A1(n10756), .A2(n10755), .ZN(n10966) );
  NAND2_X1 U10909 ( .A1(n10755), .A2(n10756), .ZN(n10964) );
  NAND2_X1 U10910 ( .A1(n10967), .A2(n10968), .ZN(n10756) );
  NAND3_X1 U10911 ( .A1(b_19_), .A2(n10969), .A3(a_9_), .ZN(n10968) );
  OR2_X1 U10912 ( .A1(n10913), .A2(n10912), .ZN(n10969) );
  NAND2_X1 U10913 ( .A1(n10912), .A2(n10913), .ZN(n10967) );
  NAND2_X1 U10914 ( .A1(n10909), .A2(n10970), .ZN(n10913) );
  NAND2_X1 U10915 ( .A1(n10908), .A2(n10910), .ZN(n10970) );
  NAND2_X1 U10916 ( .A1(n10971), .A2(n10972), .ZN(n10910) );
  NAND2_X1 U10917 ( .A1(a_10_), .A2(b_19_), .ZN(n10972) );
  INV_X1 U10918 ( .A(n10973), .ZN(n10971) );
  XNOR2_X1 U10919 ( .A(n10974), .B(n10975), .ZN(n10908) );
  XNOR2_X1 U10920 ( .A(n10976), .B(n10977), .ZN(n10974) );
  NAND2_X1 U10921 ( .A1(a_10_), .A2(n10973), .ZN(n10909) );
  NAND2_X1 U10922 ( .A1(n10905), .A2(n10978), .ZN(n10973) );
  NAND2_X1 U10923 ( .A1(n10904), .A2(n10906), .ZN(n10978) );
  NAND2_X1 U10924 ( .A1(n10979), .A2(n10980), .ZN(n10906) );
  NAND2_X1 U10925 ( .A1(a_11_), .A2(b_19_), .ZN(n10980) );
  INV_X1 U10926 ( .A(n10981), .ZN(n10979) );
  XNOR2_X1 U10927 ( .A(n10982), .B(n10983), .ZN(n10904) );
  XNOR2_X1 U10928 ( .A(n10984), .B(n10985), .ZN(n10983) );
  NAND2_X1 U10929 ( .A1(a_11_), .A2(n10981), .ZN(n10905) );
  NAND2_X1 U10930 ( .A1(n10986), .A2(n10987), .ZN(n10981) );
  NAND3_X1 U10931 ( .A1(b_19_), .A2(n10988), .A3(a_12_), .ZN(n10987) );
  OR2_X1 U10932 ( .A1(n10901), .A2(n10899), .ZN(n10988) );
  NAND2_X1 U10933 ( .A1(n10899), .A2(n10901), .ZN(n10986) );
  NAND2_X1 U10934 ( .A1(n10989), .A2(n10990), .ZN(n10901) );
  NAND2_X1 U10935 ( .A1(n10898), .A2(n10991), .ZN(n10990) );
  OR2_X1 U10936 ( .A1(n10897), .A2(n10896), .ZN(n10991) );
  NOR2_X1 U10937 ( .A1(n7789), .A2(n7693), .ZN(n10898) );
  NAND2_X1 U10938 ( .A1(n10896), .A2(n10897), .ZN(n10989) );
  NAND2_X1 U10939 ( .A1(n10992), .A2(n10993), .ZN(n10897) );
  NAND3_X1 U10940 ( .A1(b_19_), .A2(n10994), .A3(a_14_), .ZN(n10993) );
  NAND2_X1 U10941 ( .A1(n10893), .A2(n10892), .ZN(n10994) );
  OR2_X1 U10942 ( .A1(n10892), .A2(n10893), .ZN(n10992) );
  AND2_X1 U10943 ( .A1(n10995), .A2(n10996), .ZN(n10893) );
  NAND2_X1 U10944 ( .A1(n10890), .A2(n10997), .ZN(n10996) );
  OR2_X1 U10945 ( .A1(n10889), .A2(n10887), .ZN(n10997) );
  NOR2_X1 U10946 ( .A1(n7754), .A2(n7693), .ZN(n10890) );
  NAND2_X1 U10947 ( .A1(n10887), .A2(n10889), .ZN(n10995) );
  NAND2_X1 U10948 ( .A1(n10998), .A2(n10999), .ZN(n10889) );
  NAND3_X1 U10949 ( .A1(b_19_), .A2(n11000), .A3(a_16_), .ZN(n10999) );
  OR2_X1 U10950 ( .A1(n10885), .A2(n10883), .ZN(n11000) );
  NAND2_X1 U10951 ( .A1(n10883), .A2(n10885), .ZN(n10998) );
  NAND2_X1 U10952 ( .A1(n11001), .A2(n11002), .ZN(n10885) );
  NAND2_X1 U10953 ( .A1(n10882), .A2(n11003), .ZN(n11002) );
  OR2_X1 U10954 ( .A1(n10881), .A2(n10880), .ZN(n11003) );
  NOR2_X1 U10955 ( .A1(n7732), .A2(n7693), .ZN(n10882) );
  NAND2_X1 U10956 ( .A1(n10880), .A2(n10881), .ZN(n11001) );
  NAND2_X1 U10957 ( .A1(n11004), .A2(n11005), .ZN(n10881) );
  NAND3_X1 U10958 ( .A1(b_19_), .A2(n11006), .A3(a_18_), .ZN(n11005) );
  NAND2_X1 U10959 ( .A1(n10877), .A2(n10876), .ZN(n11006) );
  OR2_X1 U10960 ( .A1(n10876), .A2(n10877), .ZN(n11004) );
  AND2_X1 U10961 ( .A1(n11007), .A2(n11008), .ZN(n10877) );
  NAND2_X1 U10962 ( .A1(n7691), .A2(n11009), .ZN(n11008) );
  OR2_X1 U10963 ( .A1(n10874), .A2(n10873), .ZN(n11009) );
  INV_X1 U10964 ( .A(n8011), .ZN(n7691) );
  NAND2_X1 U10965 ( .A1(a_19_), .A2(b_19_), .ZN(n8011) );
  NAND2_X1 U10966 ( .A1(n10873), .A2(n10874), .ZN(n11007) );
  NAND2_X1 U10967 ( .A1(n11010), .A2(n11011), .ZN(n10874) );
  NAND3_X1 U10968 ( .A1(a_20_), .A2(n11012), .A3(b_19_), .ZN(n11011) );
  NAND2_X1 U10969 ( .A1(n10871), .A2(n10869), .ZN(n11012) );
  OR2_X1 U10970 ( .A1(n10869), .A2(n10871), .ZN(n11010) );
  AND2_X1 U10971 ( .A1(n11013), .A2(n11014), .ZN(n10871) );
  NAND2_X1 U10972 ( .A1(n10800), .A2(n11015), .ZN(n11014) );
  NAND2_X1 U10973 ( .A1(n10799), .A2(n10798), .ZN(n11015) );
  NOR2_X1 U10974 ( .A1(n7693), .A2(n7665), .ZN(n10800) );
  OR2_X1 U10975 ( .A1(n10798), .A2(n10799), .ZN(n11013) );
  AND2_X1 U10976 ( .A1(n11016), .A2(n11017), .ZN(n10799) );
  NAND3_X1 U10977 ( .A1(a_22_), .A2(n11018), .A3(b_19_), .ZN(n11017) );
  OR2_X1 U10978 ( .A1(n10866), .A2(n10864), .ZN(n11018) );
  NAND2_X1 U10979 ( .A1(n10864), .A2(n10866), .ZN(n11016) );
  NAND2_X1 U10980 ( .A1(n11019), .A2(n11020), .ZN(n10866) );
  NAND2_X1 U10981 ( .A1(n10863), .A2(n11021), .ZN(n11020) );
  OR2_X1 U10982 ( .A1(n10862), .A2(n10860), .ZN(n11021) );
  NOR2_X1 U10983 ( .A1(n7693), .A2(n8042), .ZN(n10863) );
  NAND2_X1 U10984 ( .A1(n10860), .A2(n10862), .ZN(n11019) );
  NAND2_X1 U10985 ( .A1(n11022), .A2(n11023), .ZN(n10862) );
  NAND3_X1 U10986 ( .A1(a_24_), .A2(n11024), .A3(b_19_), .ZN(n11023) );
  NAND2_X1 U10987 ( .A1(n10858), .A2(n10857), .ZN(n11024) );
  OR2_X1 U10988 ( .A1(n10857), .A2(n10858), .ZN(n11022) );
  AND2_X1 U10989 ( .A1(n11025), .A2(n11026), .ZN(n10858) );
  NAND2_X1 U10990 ( .A1(n10855), .A2(n11027), .ZN(n11026) );
  OR2_X1 U10991 ( .A1(n10854), .A2(n10853), .ZN(n11027) );
  NOR2_X1 U10992 ( .A1(n7693), .A2(n8039), .ZN(n10855) );
  NAND2_X1 U10993 ( .A1(n10853), .A2(n10854), .ZN(n11025) );
  NAND2_X1 U10994 ( .A1(n10850), .A2(n11028), .ZN(n10854) );
  NAND2_X1 U10995 ( .A1(n10849), .A2(n10851), .ZN(n11028) );
  NAND2_X1 U10996 ( .A1(n11029), .A2(n11030), .ZN(n10851) );
  NAND2_X1 U10997 ( .A1(b_19_), .A2(a_26_), .ZN(n11030) );
  INV_X1 U10998 ( .A(n11031), .ZN(n11029) );
  XNOR2_X1 U10999 ( .A(n11032), .B(n11033), .ZN(n10849) );
  NAND2_X1 U11000 ( .A1(n11034), .A2(n11035), .ZN(n11032) );
  NAND2_X1 U11001 ( .A1(a_26_), .A2(n11031), .ZN(n10850) );
  NAND2_X1 U11002 ( .A1(n10822), .A2(n11036), .ZN(n11031) );
  NAND2_X1 U11003 ( .A1(n10821), .A2(n10823), .ZN(n11036) );
  NAND2_X1 U11004 ( .A1(n11037), .A2(n11038), .ZN(n10823) );
  NAND2_X1 U11005 ( .A1(b_19_), .A2(a_27_), .ZN(n11038) );
  INV_X1 U11006 ( .A(n11039), .ZN(n11037) );
  XNOR2_X1 U11007 ( .A(n11040), .B(n11041), .ZN(n10821) );
  XOR2_X1 U11008 ( .A(n11042), .B(n11043), .Z(n11040) );
  NAND2_X1 U11009 ( .A1(b_18_), .A2(a_28_), .ZN(n11042) );
  NAND2_X1 U11010 ( .A1(a_27_), .A2(n11039), .ZN(n10822) );
  NAND2_X1 U11011 ( .A1(n11044), .A2(n11045), .ZN(n11039) );
  NAND3_X1 U11012 ( .A1(a_28_), .A2(n11046), .A3(b_19_), .ZN(n11045) );
  NAND2_X1 U11013 ( .A1(n10831), .A2(n10829), .ZN(n11046) );
  OR2_X1 U11014 ( .A1(n10829), .A2(n10831), .ZN(n11044) );
  AND2_X1 U11015 ( .A1(n11047), .A2(n11048), .ZN(n10831) );
  NAND2_X1 U11016 ( .A1(n10845), .A2(n11049), .ZN(n11048) );
  OR2_X1 U11017 ( .A1(n10846), .A2(n10847), .ZN(n11049) );
  NOR2_X1 U11018 ( .A1(n7693), .A2(n7545), .ZN(n10845) );
  NAND2_X1 U11019 ( .A1(n10847), .A2(n10846), .ZN(n11047) );
  NAND2_X1 U11020 ( .A1(n11050), .A2(n11051), .ZN(n10846) );
  NAND2_X1 U11021 ( .A1(b_17_), .A2(n11052), .ZN(n11051) );
  NAND2_X1 U11022 ( .A1(n7527), .A2(n11053), .ZN(n11052) );
  NAND2_X1 U11023 ( .A1(a_31_), .A2(n8046), .ZN(n11053) );
  NAND2_X1 U11024 ( .A1(b_18_), .A2(n11054), .ZN(n11050) );
  NAND2_X1 U11025 ( .A1(n7531), .A2(n11055), .ZN(n11054) );
  NAND2_X1 U11026 ( .A1(a_30_), .A2(n7725), .ZN(n11055) );
  AND3_X1 U11027 ( .A1(b_18_), .A2(b_19_), .A3(n7494), .ZN(n10847) );
  XNOR2_X1 U11028 ( .A(n11056), .B(n11057), .ZN(n10829) );
  XOR2_X1 U11029 ( .A(n11058), .B(n11059), .Z(n11056) );
  XNOR2_X1 U11030 ( .A(n11060), .B(n11061), .ZN(n10853) );
  NAND2_X1 U11031 ( .A1(n11062), .A2(n11063), .ZN(n11060) );
  XNOR2_X1 U11032 ( .A(n11064), .B(n11065), .ZN(n10857) );
  XOR2_X1 U11033 ( .A(n11066), .B(n11067), .Z(n11064) );
  XNOR2_X1 U11034 ( .A(n11068), .B(n11069), .ZN(n10860) );
  XNOR2_X1 U11035 ( .A(n11070), .B(n11071), .ZN(n11068) );
  NOR2_X1 U11036 ( .A1(n8041), .A2(n8046), .ZN(n11071) );
  XNOR2_X1 U11037 ( .A(n11072), .B(n11073), .ZN(n10864) );
  XOR2_X1 U11038 ( .A(n11074), .B(n11075), .Z(n11073) );
  NAND2_X1 U11039 ( .A1(b_18_), .A2(a_23_), .ZN(n11075) );
  XOR2_X1 U11040 ( .A(n11076), .B(n11077), .Z(n10798) );
  NAND2_X1 U11041 ( .A1(n11078), .A2(n11079), .ZN(n11076) );
  XNOR2_X1 U11042 ( .A(n11080), .B(n11081), .ZN(n10869) );
  XOR2_X1 U11043 ( .A(n11082), .B(n11083), .Z(n11080) );
  XNOR2_X1 U11044 ( .A(n11084), .B(n11085), .ZN(n10873) );
  XNOR2_X1 U11045 ( .A(n11086), .B(n11087), .ZN(n11084) );
  NOR2_X1 U11046 ( .A1(n8044), .A2(n8046), .ZN(n11087) );
  XOR2_X1 U11047 ( .A(n11088), .B(n11089), .Z(n10876) );
  XNOR2_X1 U11048 ( .A(n11090), .B(n11091), .ZN(n11089) );
  XOR2_X1 U11049 ( .A(n11092), .B(n11093), .Z(n10880) );
  XOR2_X1 U11050 ( .A(n11094), .B(n11095), .Z(n11092) );
  XNOR2_X1 U11051 ( .A(n11096), .B(n11097), .ZN(n10883) );
  XNOR2_X1 U11052 ( .A(n11098), .B(n11099), .ZN(n11097) );
  XNOR2_X1 U11053 ( .A(n11100), .B(n11101), .ZN(n10887) );
  XOR2_X1 U11054 ( .A(n11102), .B(n11103), .Z(n11101) );
  NAND2_X1 U11055 ( .A1(a_16_), .A2(b_18_), .ZN(n11103) );
  XOR2_X1 U11056 ( .A(n11104), .B(n11105), .Z(n10892) );
  XNOR2_X1 U11057 ( .A(n11106), .B(n11107), .ZN(n11105) );
  XNOR2_X1 U11058 ( .A(n11108), .B(n11109), .ZN(n10896) );
  XNOR2_X1 U11059 ( .A(n11110), .B(n11111), .ZN(n11108) );
  NOR2_X1 U11060 ( .A1(n8046), .A2(n8049), .ZN(n11111) );
  XNOR2_X1 U11061 ( .A(n11112), .B(n11113), .ZN(n10899) );
  XNOR2_X1 U11062 ( .A(n11114), .B(n11115), .ZN(n11112) );
  NOR2_X1 U11063 ( .A1(n8046), .A2(n7789), .ZN(n11115) );
  XNOR2_X1 U11064 ( .A(n11116), .B(n11117), .ZN(n10912) );
  XNOR2_X1 U11065 ( .A(n11118), .B(n11119), .ZN(n11116) );
  NOR2_X1 U11066 ( .A1(n8046), .A2(n8051), .ZN(n11119) );
  XNOR2_X1 U11067 ( .A(n11120), .B(n11121), .ZN(n10755) );
  NAND2_X1 U11068 ( .A1(n11122), .A2(n11123), .ZN(n11120) );
  XNOR2_X1 U11069 ( .A(n11124), .B(n11125), .ZN(n10746) );
  NAND2_X1 U11070 ( .A1(n11126), .A2(n11127), .ZN(n11124) );
  XOR2_X1 U11071 ( .A(n11128), .B(n11129), .Z(n10916) );
  NAND2_X1 U11072 ( .A1(n11130), .A2(n11131), .ZN(n11128) );
  XNOR2_X1 U11073 ( .A(n11132), .B(n11133), .ZN(n10919) );
  NAND2_X1 U11074 ( .A1(n11134), .A2(n11135), .ZN(n11132) );
  XNOR2_X1 U11075 ( .A(n11136), .B(n11137), .ZN(n10733) );
  NAND2_X1 U11076 ( .A1(n11138), .A2(n11139), .ZN(n11136) );
  XNOR2_X1 U11077 ( .A(n11140), .B(n11141), .ZN(n10724) );
  NAND2_X1 U11078 ( .A1(n11142), .A2(n11143), .ZN(n11140) );
  XNOR2_X1 U11079 ( .A(n11144), .B(n11145), .ZN(n10923) );
  NAND2_X1 U11080 ( .A1(n11146), .A2(n11147), .ZN(n11144) );
  XNOR2_X1 U11081 ( .A(n11148), .B(n11149), .ZN(n10927) );
  NAND2_X1 U11082 ( .A1(n11150), .A2(n11151), .ZN(n11148) );
  XNOR2_X1 U11083 ( .A(n11152), .B(n11153), .ZN(n10931) );
  XNOR2_X1 U11084 ( .A(n11154), .B(n11155), .ZN(n11153) );
  XOR2_X1 U11085 ( .A(n8225), .B(n8226), .Z(n10935) );
  NAND2_X1 U11086 ( .A1(n11156), .A2(n11157), .ZN(n8137) );
  NAND2_X1 U11087 ( .A1(n8226), .A2(n8225), .ZN(n11157) );
  XOR2_X1 U11088 ( .A(n8216), .B(n11158), .Z(n11156) );
  NAND3_X1 U11089 ( .A1(n8226), .A2(n8225), .A3(n11159), .ZN(n8136) );
  XOR2_X1 U11090 ( .A(n8216), .B(n8215), .Z(n11159) );
  NAND2_X1 U11091 ( .A1(n11160), .A2(n11161), .ZN(n8225) );
  NAND3_X1 U11092 ( .A1(b_18_), .A2(n11162), .A3(a_0_), .ZN(n11161) );
  OR2_X1 U11093 ( .A1(n10937), .A2(n10938), .ZN(n11162) );
  NAND2_X1 U11094 ( .A1(n10937), .A2(n10938), .ZN(n11160) );
  NAND2_X1 U11095 ( .A1(n11163), .A2(n11164), .ZN(n10938) );
  NAND2_X1 U11096 ( .A1(n11155), .A2(n11165), .ZN(n11164) );
  OR2_X1 U11097 ( .A1(n11152), .A2(n11154), .ZN(n11165) );
  NOR2_X1 U11098 ( .A1(n8046), .A2(n7957), .ZN(n11155) );
  NAND2_X1 U11099 ( .A1(n11152), .A2(n11154), .ZN(n11163) );
  NAND2_X1 U11100 ( .A1(n11150), .A2(n11166), .ZN(n11154) );
  NAND2_X1 U11101 ( .A1(n11149), .A2(n11151), .ZN(n11166) );
  NAND2_X1 U11102 ( .A1(n11167), .A2(n11168), .ZN(n11151) );
  NAND2_X1 U11103 ( .A1(a_2_), .A2(b_18_), .ZN(n11168) );
  INV_X1 U11104 ( .A(n11169), .ZN(n11167) );
  XNOR2_X1 U11105 ( .A(n11170), .B(n11171), .ZN(n11149) );
  XOR2_X1 U11106 ( .A(n11172), .B(n11173), .Z(n11171) );
  NAND2_X1 U11107 ( .A1(a_3_), .A2(b_17_), .ZN(n11173) );
  NAND2_X1 U11108 ( .A1(a_2_), .A2(n11169), .ZN(n11150) );
  NAND2_X1 U11109 ( .A1(n11146), .A2(n11174), .ZN(n11169) );
  NAND2_X1 U11110 ( .A1(n11145), .A2(n11147), .ZN(n11174) );
  NAND2_X1 U11111 ( .A1(n11175), .A2(n11176), .ZN(n11147) );
  NAND2_X1 U11112 ( .A1(a_3_), .A2(b_18_), .ZN(n11176) );
  INV_X1 U11113 ( .A(n11177), .ZN(n11175) );
  XNOR2_X1 U11114 ( .A(n11178), .B(n11179), .ZN(n11145) );
  XNOR2_X1 U11115 ( .A(n11180), .B(n11181), .ZN(n11178) );
  NOR2_X1 U11116 ( .A1(n7725), .A2(n7916), .ZN(n11181) );
  NAND2_X1 U11117 ( .A1(a_3_), .A2(n11177), .ZN(n11146) );
  NAND2_X1 U11118 ( .A1(n11142), .A2(n11182), .ZN(n11177) );
  NAND2_X1 U11119 ( .A1(n11141), .A2(n11143), .ZN(n11182) );
  NAND2_X1 U11120 ( .A1(n11183), .A2(n11184), .ZN(n11143) );
  NAND2_X1 U11121 ( .A1(a_4_), .A2(b_18_), .ZN(n11184) );
  INV_X1 U11122 ( .A(n11185), .ZN(n11183) );
  XNOR2_X1 U11123 ( .A(n11186), .B(n11187), .ZN(n11141) );
  XOR2_X1 U11124 ( .A(n11188), .B(n11189), .Z(n11187) );
  NAND2_X1 U11125 ( .A1(a_5_), .A2(b_17_), .ZN(n11189) );
  NAND2_X1 U11126 ( .A1(a_4_), .A2(n11185), .ZN(n11142) );
  NAND2_X1 U11127 ( .A1(n11138), .A2(n11190), .ZN(n11185) );
  NAND2_X1 U11128 ( .A1(n11137), .A2(n11139), .ZN(n11190) );
  NAND2_X1 U11129 ( .A1(n11191), .A2(n11192), .ZN(n11139) );
  NAND2_X1 U11130 ( .A1(a_5_), .A2(b_18_), .ZN(n11192) );
  INV_X1 U11131 ( .A(n11193), .ZN(n11191) );
  XNOR2_X1 U11132 ( .A(n11194), .B(n11195), .ZN(n11137) );
  XOR2_X1 U11133 ( .A(n11196), .B(n11197), .Z(n11195) );
  NAND2_X1 U11134 ( .A1(a_6_), .A2(b_17_), .ZN(n11197) );
  NAND2_X1 U11135 ( .A1(a_5_), .A2(n11193), .ZN(n11138) );
  NAND2_X1 U11136 ( .A1(n11134), .A2(n11198), .ZN(n11193) );
  NAND2_X1 U11137 ( .A1(n11133), .A2(n11135), .ZN(n11198) );
  NAND2_X1 U11138 ( .A1(n11199), .A2(n11200), .ZN(n11135) );
  NAND2_X1 U11139 ( .A1(a_6_), .A2(b_18_), .ZN(n11200) );
  INV_X1 U11140 ( .A(n11201), .ZN(n11199) );
  XNOR2_X1 U11141 ( .A(n11202), .B(n11203), .ZN(n11133) );
  XOR2_X1 U11142 ( .A(n11204), .B(n11205), .Z(n11203) );
  NAND2_X1 U11143 ( .A1(a_7_), .A2(b_17_), .ZN(n11205) );
  NAND2_X1 U11144 ( .A1(a_6_), .A2(n11201), .ZN(n11134) );
  NAND2_X1 U11145 ( .A1(n11130), .A2(n11206), .ZN(n11201) );
  NAND2_X1 U11146 ( .A1(n11129), .A2(n11131), .ZN(n11206) );
  NAND2_X1 U11147 ( .A1(n11207), .A2(n11208), .ZN(n11131) );
  NAND2_X1 U11148 ( .A1(a_7_), .A2(b_18_), .ZN(n11208) );
  INV_X1 U11149 ( .A(n11209), .ZN(n11207) );
  XNOR2_X1 U11150 ( .A(n11210), .B(n11211), .ZN(n11129) );
  XOR2_X1 U11151 ( .A(n11212), .B(n11213), .Z(n11211) );
  NAND2_X1 U11152 ( .A1(a_8_), .A2(b_17_), .ZN(n11213) );
  NAND2_X1 U11153 ( .A1(a_7_), .A2(n11209), .ZN(n11130) );
  NAND2_X1 U11154 ( .A1(n11126), .A2(n11214), .ZN(n11209) );
  NAND2_X1 U11155 ( .A1(n11125), .A2(n11127), .ZN(n11214) );
  NAND2_X1 U11156 ( .A1(n11215), .A2(n11216), .ZN(n11127) );
  NAND2_X1 U11157 ( .A1(a_8_), .A2(b_18_), .ZN(n11216) );
  INV_X1 U11158 ( .A(n11217), .ZN(n11215) );
  XNOR2_X1 U11159 ( .A(n11218), .B(n11219), .ZN(n11125) );
  XNOR2_X1 U11160 ( .A(n11220), .B(n11221), .ZN(n11218) );
  NOR2_X1 U11161 ( .A1(n7725), .A2(n8052), .ZN(n11221) );
  NAND2_X1 U11162 ( .A1(a_8_), .A2(n11217), .ZN(n11126) );
  NAND2_X1 U11163 ( .A1(n11122), .A2(n11222), .ZN(n11217) );
  NAND2_X1 U11164 ( .A1(n11121), .A2(n11123), .ZN(n11222) );
  NAND2_X1 U11165 ( .A1(n11223), .A2(n11224), .ZN(n11123) );
  NAND2_X1 U11166 ( .A1(a_9_), .A2(b_18_), .ZN(n11224) );
  INV_X1 U11167 ( .A(n11225), .ZN(n11223) );
  XNOR2_X1 U11168 ( .A(n11226), .B(n11227), .ZN(n11121) );
  XNOR2_X1 U11169 ( .A(n11228), .B(n11229), .ZN(n11226) );
  NOR2_X1 U11170 ( .A1(n7725), .A2(n8051), .ZN(n11229) );
  NAND2_X1 U11171 ( .A1(a_9_), .A2(n11225), .ZN(n11122) );
  NAND2_X1 U11172 ( .A1(n11230), .A2(n11231), .ZN(n11225) );
  NAND3_X1 U11173 ( .A1(b_18_), .A2(n11232), .A3(a_10_), .ZN(n11231) );
  NAND2_X1 U11174 ( .A1(n11118), .A2(n11117), .ZN(n11232) );
  OR2_X1 U11175 ( .A1(n11117), .A2(n11118), .ZN(n11230) );
  AND2_X1 U11176 ( .A1(n11233), .A2(n11234), .ZN(n11118) );
  NAND2_X1 U11177 ( .A1(n10976), .A2(n11235), .ZN(n11234) );
  NAND2_X1 U11178 ( .A1(n10977), .A2(n10975), .ZN(n11235) );
  NOR2_X1 U11179 ( .A1(n7811), .A2(n8046), .ZN(n10976) );
  OR2_X1 U11180 ( .A1(n10975), .A2(n10977), .ZN(n11233) );
  AND2_X1 U11181 ( .A1(n11236), .A2(n11237), .ZN(n10977) );
  NAND2_X1 U11182 ( .A1(n10985), .A2(n11238), .ZN(n11237) );
  OR2_X1 U11183 ( .A1(n10982), .A2(n10984), .ZN(n11238) );
  NOR2_X1 U11184 ( .A1(n8669), .A2(n8046), .ZN(n10985) );
  NAND2_X1 U11185 ( .A1(n10982), .A2(n10984), .ZN(n11236) );
  NAND2_X1 U11186 ( .A1(n11239), .A2(n11240), .ZN(n10984) );
  NAND3_X1 U11187 ( .A1(b_18_), .A2(n11241), .A3(a_13_), .ZN(n11240) );
  NAND2_X1 U11188 ( .A1(n11114), .A2(n11113), .ZN(n11241) );
  OR2_X1 U11189 ( .A1(n11113), .A2(n11114), .ZN(n11239) );
  AND2_X1 U11190 ( .A1(n11242), .A2(n11243), .ZN(n11114) );
  NAND3_X1 U11191 ( .A1(b_18_), .A2(n11244), .A3(a_14_), .ZN(n11243) );
  NAND2_X1 U11192 ( .A1(n11110), .A2(n11109), .ZN(n11244) );
  OR2_X1 U11193 ( .A1(n11109), .A2(n11110), .ZN(n11242) );
  AND2_X1 U11194 ( .A1(n11245), .A2(n11246), .ZN(n11110) );
  NAND2_X1 U11195 ( .A1(n11107), .A2(n11247), .ZN(n11246) );
  OR2_X1 U11196 ( .A1(n11104), .A2(n11106), .ZN(n11247) );
  NOR2_X1 U11197 ( .A1(n7754), .A2(n8046), .ZN(n11107) );
  NAND2_X1 U11198 ( .A1(n11104), .A2(n11106), .ZN(n11245) );
  NAND2_X1 U11199 ( .A1(n11248), .A2(n11249), .ZN(n11106) );
  NAND3_X1 U11200 ( .A1(b_18_), .A2(n11250), .A3(a_16_), .ZN(n11249) );
  OR2_X1 U11201 ( .A1(n11102), .A2(n11100), .ZN(n11250) );
  NAND2_X1 U11202 ( .A1(n11100), .A2(n11102), .ZN(n11248) );
  NAND2_X1 U11203 ( .A1(n11251), .A2(n11252), .ZN(n11102) );
  NAND2_X1 U11204 ( .A1(n11099), .A2(n11253), .ZN(n11252) );
  OR2_X1 U11205 ( .A1(n11096), .A2(n11098), .ZN(n11253) );
  NOR2_X1 U11206 ( .A1(n7732), .A2(n8046), .ZN(n11099) );
  NAND2_X1 U11207 ( .A1(n11096), .A2(n11098), .ZN(n11251) );
  NAND2_X1 U11208 ( .A1(n11254), .A2(n11255), .ZN(n11098) );
  NAND2_X1 U11209 ( .A1(n11093), .A2(n11256), .ZN(n11255) );
  OR2_X1 U11210 ( .A1(n11094), .A2(n11095), .ZN(n11256) );
  XNOR2_X1 U11211 ( .A(n11257), .B(n11258), .ZN(n11093) );
  XNOR2_X1 U11212 ( .A(n11259), .B(n11260), .ZN(n11258) );
  NAND2_X1 U11213 ( .A1(n11095), .A2(n11094), .ZN(n11254) );
  NAND2_X1 U11214 ( .A1(n11261), .A2(n11262), .ZN(n11094) );
  NAND2_X1 U11215 ( .A1(n11091), .A2(n11263), .ZN(n11262) );
  OR2_X1 U11216 ( .A1(n11088), .A2(n11090), .ZN(n11263) );
  NOR2_X1 U11217 ( .A1(n8046), .A2(n8045), .ZN(n11091) );
  NAND2_X1 U11218 ( .A1(n11088), .A2(n11090), .ZN(n11261) );
  NAND2_X1 U11219 ( .A1(n11264), .A2(n11265), .ZN(n11090) );
  NAND3_X1 U11220 ( .A1(a_20_), .A2(n11266), .A3(b_18_), .ZN(n11265) );
  NAND2_X1 U11221 ( .A1(n11086), .A2(n11085), .ZN(n11266) );
  OR2_X1 U11222 ( .A1(n11085), .A2(n11086), .ZN(n11264) );
  AND2_X1 U11223 ( .A1(n11267), .A2(n11268), .ZN(n11086) );
  NAND2_X1 U11224 ( .A1(n11082), .A2(n11269), .ZN(n11268) );
  OR2_X1 U11225 ( .A1(n11081), .A2(n11083), .ZN(n11269) );
  NOR2_X1 U11226 ( .A1(n8046), .A2(n7665), .ZN(n11082) );
  NAND2_X1 U11227 ( .A1(n11081), .A2(n11083), .ZN(n11267) );
  NAND2_X1 U11228 ( .A1(n11078), .A2(n11270), .ZN(n11083) );
  NAND2_X1 U11229 ( .A1(n11077), .A2(n11079), .ZN(n11270) );
  NAND2_X1 U11230 ( .A1(n11271), .A2(n11272), .ZN(n11079) );
  NAND2_X1 U11231 ( .A1(b_18_), .A2(a_22_), .ZN(n11272) );
  INV_X1 U11232 ( .A(n11273), .ZN(n11271) );
  XNOR2_X1 U11233 ( .A(n11274), .B(n11275), .ZN(n11077) );
  XNOR2_X1 U11234 ( .A(n11276), .B(n11277), .ZN(n11275) );
  NAND2_X1 U11235 ( .A1(a_22_), .A2(n11273), .ZN(n11078) );
  NAND2_X1 U11236 ( .A1(n11278), .A2(n11279), .ZN(n11273) );
  NAND3_X1 U11237 ( .A1(a_23_), .A2(n11280), .A3(b_18_), .ZN(n11279) );
  OR2_X1 U11238 ( .A1(n11072), .A2(n11074), .ZN(n11280) );
  NAND2_X1 U11239 ( .A1(n11072), .A2(n11074), .ZN(n11278) );
  NAND2_X1 U11240 ( .A1(n11281), .A2(n11282), .ZN(n11074) );
  NAND3_X1 U11241 ( .A1(a_24_), .A2(n11283), .A3(b_18_), .ZN(n11282) );
  NAND2_X1 U11242 ( .A1(n11070), .A2(n11069), .ZN(n11283) );
  OR2_X1 U11243 ( .A1(n11069), .A2(n11070), .ZN(n11281) );
  AND2_X1 U11244 ( .A1(n11284), .A2(n11285), .ZN(n11070) );
  NAND2_X1 U11245 ( .A1(n11067), .A2(n11286), .ZN(n11285) );
  OR2_X1 U11246 ( .A1(n11065), .A2(n11066), .ZN(n11286) );
  NOR2_X1 U11247 ( .A1(n8046), .A2(n8039), .ZN(n11067) );
  NAND2_X1 U11248 ( .A1(n11065), .A2(n11066), .ZN(n11284) );
  NAND2_X1 U11249 ( .A1(n11062), .A2(n11287), .ZN(n11066) );
  NAND2_X1 U11250 ( .A1(n11061), .A2(n11063), .ZN(n11287) );
  NAND2_X1 U11251 ( .A1(n11288), .A2(n11289), .ZN(n11063) );
  NAND2_X1 U11252 ( .A1(b_18_), .A2(a_26_), .ZN(n11289) );
  INV_X1 U11253 ( .A(n11290), .ZN(n11288) );
  XNOR2_X1 U11254 ( .A(n11291), .B(n11292), .ZN(n11061) );
  NAND2_X1 U11255 ( .A1(n11293), .A2(n11294), .ZN(n11291) );
  NAND2_X1 U11256 ( .A1(a_26_), .A2(n11290), .ZN(n11062) );
  NAND2_X1 U11257 ( .A1(n11034), .A2(n11295), .ZN(n11290) );
  NAND2_X1 U11258 ( .A1(n11033), .A2(n11035), .ZN(n11295) );
  NAND2_X1 U11259 ( .A1(n11296), .A2(n11297), .ZN(n11035) );
  NAND2_X1 U11260 ( .A1(b_18_), .A2(a_27_), .ZN(n11297) );
  INV_X1 U11261 ( .A(n11298), .ZN(n11296) );
  XNOR2_X1 U11262 ( .A(n11299), .B(n11300), .ZN(n11033) );
  XOR2_X1 U11263 ( .A(n11301), .B(n11302), .Z(n11299) );
  NAND2_X1 U11264 ( .A1(b_17_), .A2(a_28_), .ZN(n11301) );
  NAND2_X1 U11265 ( .A1(a_27_), .A2(n11298), .ZN(n11034) );
  NAND2_X1 U11266 ( .A1(n11303), .A2(n11304), .ZN(n11298) );
  NAND3_X1 U11267 ( .A1(a_28_), .A2(n11305), .A3(b_18_), .ZN(n11304) );
  NAND2_X1 U11268 ( .A1(n11043), .A2(n11041), .ZN(n11305) );
  OR2_X1 U11269 ( .A1(n11041), .A2(n11043), .ZN(n11303) );
  AND2_X1 U11270 ( .A1(n11306), .A2(n11307), .ZN(n11043) );
  NAND2_X1 U11271 ( .A1(n11057), .A2(n11308), .ZN(n11307) );
  OR2_X1 U11272 ( .A1(n11058), .A2(n11059), .ZN(n11308) );
  NOR2_X1 U11273 ( .A1(n8046), .A2(n7545), .ZN(n11057) );
  NAND2_X1 U11274 ( .A1(n11059), .A2(n11058), .ZN(n11306) );
  NAND2_X1 U11275 ( .A1(n11309), .A2(n11310), .ZN(n11058) );
  NAND2_X1 U11276 ( .A1(b_16_), .A2(n11311), .ZN(n11310) );
  NAND2_X1 U11277 ( .A1(n7527), .A2(n11312), .ZN(n11311) );
  NAND2_X1 U11278 ( .A1(a_31_), .A2(n7725), .ZN(n11312) );
  NAND2_X1 U11279 ( .A1(b_17_), .A2(n11313), .ZN(n11309) );
  NAND2_X1 U11280 ( .A1(n7531), .A2(n11314), .ZN(n11313) );
  NAND2_X1 U11281 ( .A1(a_30_), .A2(n11315), .ZN(n11314) );
  AND3_X1 U11282 ( .A1(b_18_), .A2(b_17_), .A3(n7494), .ZN(n11059) );
  XNOR2_X1 U11283 ( .A(n11316), .B(n11317), .ZN(n11041) );
  XOR2_X1 U11284 ( .A(n11318), .B(n11319), .Z(n11316) );
  XNOR2_X1 U11285 ( .A(n11320), .B(n11321), .ZN(n11065) );
  NAND2_X1 U11286 ( .A1(n11322), .A2(n11323), .ZN(n11320) );
  XNOR2_X1 U11287 ( .A(n11324), .B(n11325), .ZN(n11069) );
  XOR2_X1 U11288 ( .A(n11326), .B(n11327), .Z(n11324) );
  XNOR2_X1 U11289 ( .A(n11328), .B(n11329), .ZN(n11072) );
  XNOR2_X1 U11290 ( .A(n11330), .B(n11331), .ZN(n11328) );
  NOR2_X1 U11291 ( .A1(n8041), .A2(n7725), .ZN(n11331) );
  XNOR2_X1 U11292 ( .A(n11332), .B(n11333), .ZN(n11081) );
  XOR2_X1 U11293 ( .A(n11334), .B(n11335), .Z(n11333) );
  NAND2_X1 U11294 ( .A1(b_17_), .A2(a_22_), .ZN(n11335) );
  XNOR2_X1 U11295 ( .A(n11336), .B(n11337), .ZN(n11085) );
  XOR2_X1 U11296 ( .A(n11338), .B(n11339), .Z(n11336) );
  XNOR2_X1 U11297 ( .A(n11340), .B(n11341), .ZN(n11088) );
  XNOR2_X1 U11298 ( .A(n11342), .B(n11343), .ZN(n11340) );
  NOR2_X1 U11299 ( .A1(n8044), .A2(n7725), .ZN(n11343) );
  INV_X1 U11300 ( .A(n7711), .ZN(n11095) );
  NAND2_X1 U11301 ( .A1(b_18_), .A2(a_18_), .ZN(n7711) );
  XNOR2_X1 U11302 ( .A(n11344), .B(n11345), .ZN(n11096) );
  XNOR2_X1 U11303 ( .A(n11346), .B(n11347), .ZN(n11344) );
  NOR2_X1 U11304 ( .A1(n8047), .A2(n7725), .ZN(n11347) );
  XOR2_X1 U11305 ( .A(n11348), .B(n11349), .Z(n11100) );
  XOR2_X1 U11306 ( .A(n11350), .B(n7723), .Z(n11348) );
  XNOR2_X1 U11307 ( .A(n11351), .B(n11352), .ZN(n11104) );
  XOR2_X1 U11308 ( .A(n11353), .B(n11354), .Z(n11352) );
  NAND2_X1 U11309 ( .A1(a_16_), .A2(b_17_), .ZN(n11354) );
  XOR2_X1 U11310 ( .A(n11355), .B(n11356), .Z(n11109) );
  XNOR2_X1 U11311 ( .A(n11357), .B(n11358), .ZN(n11356) );
  XNOR2_X1 U11312 ( .A(n11359), .B(n11360), .ZN(n11113) );
  XOR2_X1 U11313 ( .A(n11361), .B(n11362), .Z(n11359) );
  XNOR2_X1 U11314 ( .A(n11363), .B(n11364), .ZN(n10982) );
  XNOR2_X1 U11315 ( .A(n11365), .B(n11366), .ZN(n11363) );
  NOR2_X1 U11316 ( .A1(n7725), .A2(n7789), .ZN(n11366) );
  XOR2_X1 U11317 ( .A(n11367), .B(n11368), .Z(n10975) );
  XOR2_X1 U11318 ( .A(n11369), .B(n11370), .Z(n11368) );
  NAND2_X1 U11319 ( .A1(a_12_), .A2(b_17_), .ZN(n11370) );
  XOR2_X1 U11320 ( .A(n11371), .B(n11372), .Z(n11117) );
  XOR2_X1 U11321 ( .A(n11373), .B(n11374), .Z(n11372) );
  NAND2_X1 U11322 ( .A1(a_11_), .A2(b_17_), .ZN(n11374) );
  XNOR2_X1 U11323 ( .A(n11375), .B(n11376), .ZN(n11152) );
  XOR2_X1 U11324 ( .A(n11377), .B(n11378), .Z(n11376) );
  NAND2_X1 U11325 ( .A1(a_2_), .A2(b_17_), .ZN(n11378) );
  XNOR2_X1 U11326 ( .A(n11379), .B(n11380), .ZN(n10937) );
  XOR2_X1 U11327 ( .A(n11381), .B(n11382), .Z(n11380) );
  NAND2_X1 U11328 ( .A1(b_17_), .A2(a_1_), .ZN(n11382) );
  XNOR2_X1 U11329 ( .A(n11383), .B(n11384), .ZN(n8226) );
  XOR2_X1 U11330 ( .A(n11385), .B(n11386), .Z(n11384) );
  NAND2_X1 U11331 ( .A1(a_0_), .A2(b_17_), .ZN(n11386) );
  NAND3_X1 U11332 ( .A1(n8215), .A2(n8216), .A3(n11387), .ZN(n8141) );
  XOR2_X1 U11333 ( .A(n8218), .B(n8217), .Z(n11387) );
  NAND2_X1 U11334 ( .A1(n11388), .A2(n11389), .ZN(n8216) );
  NAND3_X1 U11335 ( .A1(b_17_), .A2(n11390), .A3(a_0_), .ZN(n11389) );
  OR2_X1 U11336 ( .A1(n11385), .A2(n11383), .ZN(n11390) );
  NAND2_X1 U11337 ( .A1(n11383), .A2(n11385), .ZN(n11388) );
  NAND2_X1 U11338 ( .A1(n11391), .A2(n11392), .ZN(n11385) );
  NAND3_X1 U11339 ( .A1(a_1_), .A2(n11393), .A3(b_17_), .ZN(n11392) );
  OR2_X1 U11340 ( .A1(n11381), .A2(n11379), .ZN(n11393) );
  NAND2_X1 U11341 ( .A1(n11379), .A2(n11381), .ZN(n11391) );
  NAND2_X1 U11342 ( .A1(n11394), .A2(n11395), .ZN(n11381) );
  NAND3_X1 U11343 ( .A1(b_17_), .A2(n11396), .A3(a_2_), .ZN(n11395) );
  OR2_X1 U11344 ( .A1(n11377), .A2(n11375), .ZN(n11396) );
  NAND2_X1 U11345 ( .A1(n11375), .A2(n11377), .ZN(n11394) );
  NAND2_X1 U11346 ( .A1(n11397), .A2(n11398), .ZN(n11377) );
  NAND3_X1 U11347 ( .A1(b_17_), .A2(n11399), .A3(a_3_), .ZN(n11398) );
  OR2_X1 U11348 ( .A1(n11172), .A2(n11170), .ZN(n11399) );
  NAND2_X1 U11349 ( .A1(n11170), .A2(n11172), .ZN(n11397) );
  NAND2_X1 U11350 ( .A1(n11400), .A2(n11401), .ZN(n11172) );
  NAND3_X1 U11351 ( .A1(b_17_), .A2(n11402), .A3(a_4_), .ZN(n11401) );
  NAND2_X1 U11352 ( .A1(n11180), .A2(n11179), .ZN(n11402) );
  OR2_X1 U11353 ( .A1(n11179), .A2(n11180), .ZN(n11400) );
  AND2_X1 U11354 ( .A1(n11403), .A2(n11404), .ZN(n11180) );
  NAND3_X1 U11355 ( .A1(b_17_), .A2(n11405), .A3(a_5_), .ZN(n11404) );
  OR2_X1 U11356 ( .A1(n11188), .A2(n11186), .ZN(n11405) );
  NAND2_X1 U11357 ( .A1(n11186), .A2(n11188), .ZN(n11403) );
  NAND2_X1 U11358 ( .A1(n11406), .A2(n11407), .ZN(n11188) );
  NAND3_X1 U11359 ( .A1(b_17_), .A2(n11408), .A3(a_6_), .ZN(n11407) );
  OR2_X1 U11360 ( .A1(n11196), .A2(n11194), .ZN(n11408) );
  NAND2_X1 U11361 ( .A1(n11194), .A2(n11196), .ZN(n11406) );
  NAND2_X1 U11362 ( .A1(n11409), .A2(n11410), .ZN(n11196) );
  NAND3_X1 U11363 ( .A1(b_17_), .A2(n11411), .A3(a_7_), .ZN(n11410) );
  OR2_X1 U11364 ( .A1(n11204), .A2(n11202), .ZN(n11411) );
  NAND2_X1 U11365 ( .A1(n11202), .A2(n11204), .ZN(n11409) );
  NAND2_X1 U11366 ( .A1(n11412), .A2(n11413), .ZN(n11204) );
  NAND3_X1 U11367 ( .A1(b_17_), .A2(n11414), .A3(a_8_), .ZN(n11413) );
  OR2_X1 U11368 ( .A1(n11212), .A2(n11210), .ZN(n11414) );
  NAND2_X1 U11369 ( .A1(n11210), .A2(n11212), .ZN(n11412) );
  NAND2_X1 U11370 ( .A1(n11415), .A2(n11416), .ZN(n11212) );
  NAND3_X1 U11371 ( .A1(b_17_), .A2(n11417), .A3(a_9_), .ZN(n11416) );
  NAND2_X1 U11372 ( .A1(n11220), .A2(n11219), .ZN(n11417) );
  OR2_X1 U11373 ( .A1(n11219), .A2(n11220), .ZN(n11415) );
  AND2_X1 U11374 ( .A1(n11418), .A2(n11419), .ZN(n11220) );
  NAND3_X1 U11375 ( .A1(b_17_), .A2(n11420), .A3(a_10_), .ZN(n11419) );
  NAND2_X1 U11376 ( .A1(n11228), .A2(n11227), .ZN(n11420) );
  OR2_X1 U11377 ( .A1(n11227), .A2(n11228), .ZN(n11418) );
  AND2_X1 U11378 ( .A1(n11421), .A2(n11422), .ZN(n11228) );
  NAND3_X1 U11379 ( .A1(b_17_), .A2(n11423), .A3(a_11_), .ZN(n11422) );
  OR2_X1 U11380 ( .A1(n11373), .A2(n11371), .ZN(n11423) );
  NAND2_X1 U11381 ( .A1(n11371), .A2(n11373), .ZN(n11421) );
  NAND2_X1 U11382 ( .A1(n11424), .A2(n11425), .ZN(n11373) );
  NAND3_X1 U11383 ( .A1(b_17_), .A2(n11426), .A3(a_12_), .ZN(n11425) );
  OR2_X1 U11384 ( .A1(n11369), .A2(n11367), .ZN(n11426) );
  NAND2_X1 U11385 ( .A1(n11367), .A2(n11369), .ZN(n11424) );
  NAND2_X1 U11386 ( .A1(n11427), .A2(n11428), .ZN(n11369) );
  NAND3_X1 U11387 ( .A1(b_17_), .A2(n11429), .A3(a_13_), .ZN(n11428) );
  NAND2_X1 U11388 ( .A1(n11365), .A2(n11364), .ZN(n11429) );
  OR2_X1 U11389 ( .A1(n11364), .A2(n11365), .ZN(n11427) );
  AND2_X1 U11390 ( .A1(n11430), .A2(n11431), .ZN(n11365) );
  NAND2_X1 U11391 ( .A1(n11362), .A2(n11432), .ZN(n11431) );
  OR2_X1 U11392 ( .A1(n11361), .A2(n11360), .ZN(n11432) );
  NOR2_X1 U11393 ( .A1(n8049), .A2(n7725), .ZN(n11362) );
  NAND2_X1 U11394 ( .A1(n11360), .A2(n11361), .ZN(n11430) );
  NAND2_X1 U11395 ( .A1(n11433), .A2(n11434), .ZN(n11361) );
  NAND2_X1 U11396 ( .A1(n11358), .A2(n11435), .ZN(n11434) );
  OR2_X1 U11397 ( .A1(n11357), .A2(n11355), .ZN(n11435) );
  NOR2_X1 U11398 ( .A1(n7754), .A2(n7725), .ZN(n11358) );
  NAND2_X1 U11399 ( .A1(n11355), .A2(n11357), .ZN(n11433) );
  NAND2_X1 U11400 ( .A1(n11436), .A2(n11437), .ZN(n11357) );
  NAND3_X1 U11401 ( .A1(b_17_), .A2(n11438), .A3(a_16_), .ZN(n11437) );
  OR2_X1 U11402 ( .A1(n11353), .A2(n11351), .ZN(n11438) );
  NAND2_X1 U11403 ( .A1(n11351), .A2(n11353), .ZN(n11436) );
  NAND2_X1 U11404 ( .A1(n11439), .A2(n11440), .ZN(n11353) );
  NAND2_X1 U11405 ( .A1(n7723), .A2(n11441), .ZN(n11440) );
  OR2_X1 U11406 ( .A1(n11350), .A2(n11349), .ZN(n11441) );
  INV_X1 U11407 ( .A(n8007), .ZN(n7723) );
  NAND2_X1 U11408 ( .A1(a_17_), .A2(b_17_), .ZN(n8007) );
  NAND2_X1 U11409 ( .A1(n11349), .A2(n11350), .ZN(n11439) );
  NAND2_X1 U11410 ( .A1(n11442), .A2(n11443), .ZN(n11350) );
  NAND3_X1 U11411 ( .A1(a_18_), .A2(n11444), .A3(b_17_), .ZN(n11443) );
  NAND2_X1 U11412 ( .A1(n11346), .A2(n11345), .ZN(n11444) );
  OR2_X1 U11413 ( .A1(n11345), .A2(n11346), .ZN(n11442) );
  AND2_X1 U11414 ( .A1(n11445), .A2(n11446), .ZN(n11346) );
  NAND2_X1 U11415 ( .A1(n11260), .A2(n11447), .ZN(n11446) );
  OR2_X1 U11416 ( .A1(n11259), .A2(n11257), .ZN(n11447) );
  NOR2_X1 U11417 ( .A1(n7725), .A2(n8045), .ZN(n11260) );
  NAND2_X1 U11418 ( .A1(n11257), .A2(n11259), .ZN(n11445) );
  NAND2_X1 U11419 ( .A1(n11448), .A2(n11449), .ZN(n11259) );
  NAND3_X1 U11420 ( .A1(a_20_), .A2(n11450), .A3(b_17_), .ZN(n11449) );
  NAND2_X1 U11421 ( .A1(n11342), .A2(n11341), .ZN(n11450) );
  OR2_X1 U11422 ( .A1(n11341), .A2(n11342), .ZN(n11448) );
  AND2_X1 U11423 ( .A1(n11451), .A2(n11452), .ZN(n11342) );
  NAND2_X1 U11424 ( .A1(n11339), .A2(n11453), .ZN(n11452) );
  OR2_X1 U11425 ( .A1(n11338), .A2(n11337), .ZN(n11453) );
  NOR2_X1 U11426 ( .A1(n7725), .A2(n7665), .ZN(n11339) );
  NAND2_X1 U11427 ( .A1(n11337), .A2(n11338), .ZN(n11451) );
  NAND2_X1 U11428 ( .A1(n11454), .A2(n11455), .ZN(n11338) );
  NAND3_X1 U11429 ( .A1(a_22_), .A2(n11456), .A3(b_17_), .ZN(n11455) );
  OR2_X1 U11430 ( .A1(n11334), .A2(n11332), .ZN(n11456) );
  NAND2_X1 U11431 ( .A1(n11332), .A2(n11334), .ZN(n11454) );
  NAND2_X1 U11432 ( .A1(n11457), .A2(n11458), .ZN(n11334) );
  NAND2_X1 U11433 ( .A1(n11277), .A2(n11459), .ZN(n11458) );
  OR2_X1 U11434 ( .A1(n11276), .A2(n11274), .ZN(n11459) );
  NOR2_X1 U11435 ( .A1(n7725), .A2(n8042), .ZN(n11277) );
  NAND2_X1 U11436 ( .A1(n11274), .A2(n11276), .ZN(n11457) );
  NAND2_X1 U11437 ( .A1(n11460), .A2(n11461), .ZN(n11276) );
  NAND3_X1 U11438 ( .A1(a_24_), .A2(n11462), .A3(b_17_), .ZN(n11461) );
  NAND2_X1 U11439 ( .A1(n11330), .A2(n11329), .ZN(n11462) );
  OR2_X1 U11440 ( .A1(n11329), .A2(n11330), .ZN(n11460) );
  AND2_X1 U11441 ( .A1(n11463), .A2(n11464), .ZN(n11330) );
  NAND2_X1 U11442 ( .A1(n11327), .A2(n11465), .ZN(n11464) );
  OR2_X1 U11443 ( .A1(n11326), .A2(n11325), .ZN(n11465) );
  NOR2_X1 U11444 ( .A1(n7725), .A2(n8039), .ZN(n11327) );
  NAND2_X1 U11445 ( .A1(n11325), .A2(n11326), .ZN(n11463) );
  NAND2_X1 U11446 ( .A1(n11322), .A2(n11466), .ZN(n11326) );
  NAND2_X1 U11447 ( .A1(n11321), .A2(n11323), .ZN(n11466) );
  NAND2_X1 U11448 ( .A1(n11467), .A2(n11468), .ZN(n11323) );
  NAND2_X1 U11449 ( .A1(b_17_), .A2(a_26_), .ZN(n11468) );
  INV_X1 U11450 ( .A(n11469), .ZN(n11467) );
  XNOR2_X1 U11451 ( .A(n11470), .B(n11471), .ZN(n11321) );
  NAND2_X1 U11452 ( .A1(n11472), .A2(n11473), .ZN(n11470) );
  NAND2_X1 U11453 ( .A1(a_26_), .A2(n11469), .ZN(n11322) );
  NAND2_X1 U11454 ( .A1(n11293), .A2(n11474), .ZN(n11469) );
  NAND2_X1 U11455 ( .A1(n11292), .A2(n11294), .ZN(n11474) );
  NAND2_X1 U11456 ( .A1(n11475), .A2(n11476), .ZN(n11294) );
  NAND2_X1 U11457 ( .A1(b_17_), .A2(a_27_), .ZN(n11476) );
  INV_X1 U11458 ( .A(n11477), .ZN(n11475) );
  XNOR2_X1 U11459 ( .A(n11478), .B(n11479), .ZN(n11292) );
  XOR2_X1 U11460 ( .A(n11480), .B(n11481), .Z(n11478) );
  NAND2_X1 U11461 ( .A1(b_16_), .A2(a_28_), .ZN(n11480) );
  NAND2_X1 U11462 ( .A1(a_27_), .A2(n11477), .ZN(n11293) );
  NAND2_X1 U11463 ( .A1(n11482), .A2(n11483), .ZN(n11477) );
  NAND3_X1 U11464 ( .A1(a_28_), .A2(n11484), .A3(b_17_), .ZN(n11483) );
  NAND2_X1 U11465 ( .A1(n11302), .A2(n11300), .ZN(n11484) );
  OR2_X1 U11466 ( .A1(n11300), .A2(n11302), .ZN(n11482) );
  AND2_X1 U11467 ( .A1(n11485), .A2(n11486), .ZN(n11302) );
  NAND2_X1 U11468 ( .A1(n11317), .A2(n11487), .ZN(n11486) );
  OR2_X1 U11469 ( .A1(n11318), .A2(n11319), .ZN(n11487) );
  NOR2_X1 U11470 ( .A1(n7725), .A2(n7545), .ZN(n11317) );
  NAND2_X1 U11471 ( .A1(n11319), .A2(n11318), .ZN(n11485) );
  NAND2_X1 U11472 ( .A1(n11488), .A2(n11489), .ZN(n11318) );
  NAND2_X1 U11473 ( .A1(b_15_), .A2(n11490), .ZN(n11489) );
  NAND2_X1 U11474 ( .A1(n7527), .A2(n11491), .ZN(n11490) );
  NAND2_X1 U11475 ( .A1(a_31_), .A2(n11315), .ZN(n11491) );
  NAND2_X1 U11476 ( .A1(b_16_), .A2(n11492), .ZN(n11488) );
  NAND2_X1 U11477 ( .A1(n7531), .A2(n11493), .ZN(n11492) );
  NAND2_X1 U11478 ( .A1(a_30_), .A2(n7756), .ZN(n11493) );
  AND3_X1 U11479 ( .A1(b_16_), .A2(b_17_), .A3(n7494), .ZN(n11319) );
  XNOR2_X1 U11480 ( .A(n11494), .B(n11495), .ZN(n11300) );
  XOR2_X1 U11481 ( .A(n11496), .B(n11497), .Z(n11494) );
  XNOR2_X1 U11482 ( .A(n11498), .B(n11499), .ZN(n11325) );
  NAND2_X1 U11483 ( .A1(n11500), .A2(n11501), .ZN(n11498) );
  XNOR2_X1 U11484 ( .A(n11502), .B(n11503), .ZN(n11329) );
  XOR2_X1 U11485 ( .A(n11504), .B(n11505), .Z(n11502) );
  XNOR2_X1 U11486 ( .A(n11506), .B(n11507), .ZN(n11274) );
  XNOR2_X1 U11487 ( .A(n11508), .B(n11509), .ZN(n11506) );
  NOR2_X1 U11488 ( .A1(n8041), .A2(n11315), .ZN(n11509) );
  XNOR2_X1 U11489 ( .A(n11510), .B(n11511), .ZN(n11332) );
  XNOR2_X1 U11490 ( .A(n11512), .B(n11513), .ZN(n11511) );
  XNOR2_X1 U11491 ( .A(n11514), .B(n11515), .ZN(n11337) );
  XNOR2_X1 U11492 ( .A(n11516), .B(n11517), .ZN(n11514) );
  NOR2_X1 U11493 ( .A1(n7650), .A2(n11315), .ZN(n11517) );
  XNOR2_X1 U11494 ( .A(n11518), .B(n11519), .ZN(n11341) );
  XOR2_X1 U11495 ( .A(n11520), .B(n11521), .Z(n11518) );
  XNOR2_X1 U11496 ( .A(n11522), .B(n11523), .ZN(n11257) );
  XNOR2_X1 U11497 ( .A(n11524), .B(n11525), .ZN(n11522) );
  NOR2_X1 U11498 ( .A1(n8044), .A2(n11315), .ZN(n11525) );
  XOR2_X1 U11499 ( .A(n11526), .B(n11527), .Z(n11345) );
  XNOR2_X1 U11500 ( .A(n11528), .B(n11529), .ZN(n11527) );
  XNOR2_X1 U11501 ( .A(n11530), .B(n11531), .ZN(n11349) );
  XNOR2_X1 U11502 ( .A(n11532), .B(n11533), .ZN(n11530) );
  NOR2_X1 U11503 ( .A1(n8047), .A2(n11315), .ZN(n11533) );
  XOR2_X1 U11504 ( .A(n11534), .B(n11535), .Z(n11351) );
  XOR2_X1 U11505 ( .A(n11536), .B(n11537), .Z(n11534) );
  XNOR2_X1 U11506 ( .A(n11538), .B(n11539), .ZN(n11355) );
  XNOR2_X1 U11507 ( .A(n11540), .B(n7744), .ZN(n11539) );
  XNOR2_X1 U11508 ( .A(n11541), .B(n11542), .ZN(n11360) );
  NAND2_X1 U11509 ( .A1(n11543), .A2(n11544), .ZN(n11541) );
  XNOR2_X1 U11510 ( .A(n11545), .B(n11546), .ZN(n11364) );
  XOR2_X1 U11511 ( .A(n11547), .B(n11548), .Z(n11545) );
  XNOR2_X1 U11512 ( .A(n11549), .B(n11550), .ZN(n11367) );
  XNOR2_X1 U11513 ( .A(n11551), .B(n11552), .ZN(n11549) );
  XNOR2_X1 U11514 ( .A(n11553), .B(n11554), .ZN(n11371) );
  XNOR2_X1 U11515 ( .A(n11555), .B(n11556), .ZN(n11553) );
  XNOR2_X1 U11516 ( .A(n11557), .B(n11558), .ZN(n11227) );
  XOR2_X1 U11517 ( .A(n11559), .B(n11560), .Z(n11557) );
  XNOR2_X1 U11518 ( .A(n11561), .B(n11562), .ZN(n11219) );
  XOR2_X1 U11519 ( .A(n11563), .B(n11564), .Z(n11561) );
  XNOR2_X1 U11520 ( .A(n11565), .B(n11566), .ZN(n11210) );
  XNOR2_X1 U11521 ( .A(n11567), .B(n11568), .ZN(n11566) );
  XNOR2_X1 U11522 ( .A(n11569), .B(n11570), .ZN(n11202) );
  XNOR2_X1 U11523 ( .A(n11571), .B(n11572), .ZN(n11569) );
  NOR2_X1 U11524 ( .A1(n11315), .A2(n8686), .ZN(n11572) );
  XNOR2_X1 U11525 ( .A(n11573), .B(n11574), .ZN(n11194) );
  XNOR2_X1 U11526 ( .A(n11575), .B(n11576), .ZN(n11574) );
  XNOR2_X1 U11527 ( .A(n11577), .B(n11578), .ZN(n11186) );
  XOR2_X1 U11528 ( .A(n11579), .B(n11580), .Z(n11578) );
  NAND2_X1 U11529 ( .A1(a_6_), .A2(b_16_), .ZN(n11580) );
  XOR2_X1 U11530 ( .A(n11581), .B(n11582), .Z(n11179) );
  NAND2_X1 U11531 ( .A1(n11583), .A2(n11584), .ZN(n11581) );
  XNOR2_X1 U11532 ( .A(n11585), .B(n11586), .ZN(n11170) );
  XNOR2_X1 U11533 ( .A(n11587), .B(n11588), .ZN(n11585) );
  XOR2_X1 U11534 ( .A(n11589), .B(n11590), .Z(n11375) );
  XOR2_X1 U11535 ( .A(n11591), .B(n11592), .Z(n11589) );
  XOR2_X1 U11536 ( .A(n11593), .B(n11594), .Z(n11379) );
  XOR2_X1 U11537 ( .A(n11595), .B(n11596), .Z(n11593) );
  XNOR2_X1 U11538 ( .A(n11597), .B(n11598), .ZN(n11383) );
  XNOR2_X1 U11539 ( .A(n11599), .B(n11600), .ZN(n11597) );
  INV_X1 U11540 ( .A(n11158), .ZN(n8215) );
  XOR2_X1 U11541 ( .A(n11601), .B(n11602), .Z(n11158) );
  XOR2_X1 U11542 ( .A(n11603), .B(n11604), .Z(n11602) );
  NAND2_X1 U11543 ( .A1(a_0_), .A2(b_16_), .ZN(n11604) );
  NAND2_X1 U11544 ( .A1(n11605), .A2(n11606), .ZN(n8147) );
  NAND2_X1 U11545 ( .A1(n8218), .A2(n8217), .ZN(n11606) );
  XOR2_X1 U11546 ( .A(n11607), .B(n11608), .Z(n11605) );
  NAND3_X1 U11547 ( .A1(n8218), .A2(n8217), .A3(n11609), .ZN(n8146) );
  XOR2_X1 U11548 ( .A(n11610), .B(n11607), .Z(n11609) );
  NAND2_X1 U11549 ( .A1(n11611), .A2(n11612), .ZN(n8217) );
  NAND3_X1 U11550 ( .A1(b_16_), .A2(n11613), .A3(a_0_), .ZN(n11612) );
  OR2_X1 U11551 ( .A1(n11603), .A2(n11601), .ZN(n11613) );
  NAND2_X1 U11552 ( .A1(n11601), .A2(n11603), .ZN(n11611) );
  NAND2_X1 U11553 ( .A1(n11614), .A2(n11615), .ZN(n11603) );
  NAND2_X1 U11554 ( .A1(n11600), .A2(n11616), .ZN(n11615) );
  NAND2_X1 U11555 ( .A1(n11599), .A2(n11598), .ZN(n11616) );
  NOR2_X1 U11556 ( .A1(n11315), .A2(n7957), .ZN(n11600) );
  OR2_X1 U11557 ( .A1(n11598), .A2(n11599), .ZN(n11614) );
  AND2_X1 U11558 ( .A1(n11617), .A2(n11618), .ZN(n11599) );
  NAND2_X1 U11559 ( .A1(n11596), .A2(n11619), .ZN(n11618) );
  OR2_X1 U11560 ( .A1(n11594), .A2(n11595), .ZN(n11619) );
  NOR2_X1 U11561 ( .A1(n8056), .A2(n11315), .ZN(n11596) );
  NAND2_X1 U11562 ( .A1(n11594), .A2(n11595), .ZN(n11617) );
  NAND2_X1 U11563 ( .A1(n11620), .A2(n11621), .ZN(n11595) );
  NAND2_X1 U11564 ( .A1(n11592), .A2(n11622), .ZN(n11621) );
  OR2_X1 U11565 ( .A1(n11590), .A2(n11591), .ZN(n11622) );
  NOR2_X1 U11566 ( .A1(n7937), .A2(n11315), .ZN(n11592) );
  NAND2_X1 U11567 ( .A1(n11590), .A2(n11591), .ZN(n11620) );
  NAND2_X1 U11568 ( .A1(n11623), .A2(n11624), .ZN(n11591) );
  NAND2_X1 U11569 ( .A1(n11588), .A2(n11625), .ZN(n11624) );
  NAND2_X1 U11570 ( .A1(n11587), .A2(n11586), .ZN(n11625) );
  NOR2_X1 U11571 ( .A1(n7916), .A2(n11315), .ZN(n11588) );
  OR2_X1 U11572 ( .A1(n11586), .A2(n11587), .ZN(n11623) );
  AND2_X1 U11573 ( .A1(n11583), .A2(n11626), .ZN(n11587) );
  NAND2_X1 U11574 ( .A1(n11582), .A2(n11584), .ZN(n11626) );
  NAND2_X1 U11575 ( .A1(n11627), .A2(n11628), .ZN(n11584) );
  NAND2_X1 U11576 ( .A1(a_5_), .A2(b_16_), .ZN(n11628) );
  INV_X1 U11577 ( .A(n11629), .ZN(n11627) );
  XOR2_X1 U11578 ( .A(n11630), .B(n11631), .Z(n11582) );
  XOR2_X1 U11579 ( .A(n11632), .B(n11633), .Z(n11630) );
  NOR2_X1 U11580 ( .A1(n7756), .A2(n7887), .ZN(n11633) );
  NAND2_X1 U11581 ( .A1(a_5_), .A2(n11629), .ZN(n11583) );
  NAND2_X1 U11582 ( .A1(n11634), .A2(n11635), .ZN(n11629) );
  NAND3_X1 U11583 ( .A1(b_16_), .A2(n11636), .A3(a_6_), .ZN(n11635) );
  OR2_X1 U11584 ( .A1(n11579), .A2(n11577), .ZN(n11636) );
  NAND2_X1 U11585 ( .A1(n11577), .A2(n11579), .ZN(n11634) );
  NAND2_X1 U11586 ( .A1(n11637), .A2(n11638), .ZN(n11579) );
  NAND2_X1 U11587 ( .A1(n11576), .A2(n11639), .ZN(n11638) );
  OR2_X1 U11588 ( .A1(n11573), .A2(n11575), .ZN(n11639) );
  NOR2_X1 U11589 ( .A1(n7872), .A2(n11315), .ZN(n11576) );
  NAND2_X1 U11590 ( .A1(n11573), .A2(n11575), .ZN(n11637) );
  NAND2_X1 U11591 ( .A1(n11640), .A2(n11641), .ZN(n11575) );
  NAND3_X1 U11592 ( .A1(b_16_), .A2(n11642), .A3(a_8_), .ZN(n11641) );
  NAND2_X1 U11593 ( .A1(n11571), .A2(n11570), .ZN(n11642) );
  OR2_X1 U11594 ( .A1(n11570), .A2(n11571), .ZN(n11640) );
  AND2_X1 U11595 ( .A1(n11643), .A2(n11644), .ZN(n11571) );
  NAND2_X1 U11596 ( .A1(n11568), .A2(n11645), .ZN(n11644) );
  OR2_X1 U11597 ( .A1(n11567), .A2(n11565), .ZN(n11645) );
  NOR2_X1 U11598 ( .A1(n8052), .A2(n11315), .ZN(n11568) );
  NAND2_X1 U11599 ( .A1(n11565), .A2(n11567), .ZN(n11643) );
  NAND2_X1 U11600 ( .A1(n11646), .A2(n11647), .ZN(n11567) );
  NAND2_X1 U11601 ( .A1(n11564), .A2(n11648), .ZN(n11647) );
  OR2_X1 U11602 ( .A1(n11562), .A2(n11563), .ZN(n11648) );
  NOR2_X1 U11603 ( .A1(n8051), .A2(n11315), .ZN(n11564) );
  NAND2_X1 U11604 ( .A1(n11562), .A2(n11563), .ZN(n11646) );
  NAND2_X1 U11605 ( .A1(n11649), .A2(n11650), .ZN(n11563) );
  NAND2_X1 U11606 ( .A1(n11560), .A2(n11651), .ZN(n11650) );
  OR2_X1 U11607 ( .A1(n11558), .A2(n11559), .ZN(n11651) );
  NOR2_X1 U11608 ( .A1(n7811), .A2(n11315), .ZN(n11560) );
  NAND2_X1 U11609 ( .A1(n11558), .A2(n11559), .ZN(n11649) );
  NAND2_X1 U11610 ( .A1(n11652), .A2(n11653), .ZN(n11559) );
  NAND2_X1 U11611 ( .A1(n11556), .A2(n11654), .ZN(n11653) );
  NAND2_X1 U11612 ( .A1(n11555), .A2(n11554), .ZN(n11654) );
  NOR2_X1 U11613 ( .A1(n8669), .A2(n11315), .ZN(n11556) );
  OR2_X1 U11614 ( .A1(n11554), .A2(n11555), .ZN(n11652) );
  AND2_X1 U11615 ( .A1(n11655), .A2(n11656), .ZN(n11555) );
  NAND2_X1 U11616 ( .A1(n11552), .A2(n11657), .ZN(n11656) );
  NAND2_X1 U11617 ( .A1(n11551), .A2(n11550), .ZN(n11657) );
  NOR2_X1 U11618 ( .A1(n7789), .A2(n11315), .ZN(n11552) );
  OR2_X1 U11619 ( .A1(n11550), .A2(n11551), .ZN(n11655) );
  AND2_X1 U11620 ( .A1(n11658), .A2(n11659), .ZN(n11551) );
  NAND2_X1 U11621 ( .A1(n11548), .A2(n11660), .ZN(n11659) );
  OR2_X1 U11622 ( .A1(n11546), .A2(n11547), .ZN(n11660) );
  NOR2_X1 U11623 ( .A1(n8049), .A2(n11315), .ZN(n11548) );
  NAND2_X1 U11624 ( .A1(n11546), .A2(n11547), .ZN(n11658) );
  NAND2_X1 U11625 ( .A1(n11543), .A2(n11661), .ZN(n11547) );
  NAND2_X1 U11626 ( .A1(n11542), .A2(n11544), .ZN(n11661) );
  NAND2_X1 U11627 ( .A1(n11662), .A2(n11663), .ZN(n11544) );
  NAND2_X1 U11628 ( .A1(a_15_), .A2(b_16_), .ZN(n11663) );
  INV_X1 U11629 ( .A(n11664), .ZN(n11662) );
  XNOR2_X1 U11630 ( .A(n11665), .B(n11666), .ZN(n11542) );
  XOR2_X1 U11631 ( .A(n11667), .B(n11668), .Z(n11666) );
  NAND2_X1 U11632 ( .A1(b_15_), .A2(a_16_), .ZN(n11668) );
  NAND2_X1 U11633 ( .A1(a_15_), .A2(n11664), .ZN(n11543) );
  NAND2_X1 U11634 ( .A1(n11669), .A2(n11670), .ZN(n11664) );
  NAND2_X1 U11635 ( .A1(n11538), .A2(n11671), .ZN(n11670) );
  OR2_X1 U11636 ( .A1(n11540), .A2(n7744), .ZN(n11671) );
  XOR2_X1 U11637 ( .A(n11672), .B(n11673), .Z(n11538) );
  XOR2_X1 U11638 ( .A(n11674), .B(n11675), .Z(n11672) );
  NAND2_X1 U11639 ( .A1(n7744), .A2(n11540), .ZN(n11669) );
  NAND2_X1 U11640 ( .A1(n11676), .A2(n11677), .ZN(n11540) );
  NAND2_X1 U11641 ( .A1(n11537), .A2(n11678), .ZN(n11677) );
  OR2_X1 U11642 ( .A1(n11535), .A2(n11536), .ZN(n11678) );
  NOR2_X1 U11643 ( .A1(n11315), .A2(n7732), .ZN(n11537) );
  NAND2_X1 U11644 ( .A1(n11535), .A2(n11536), .ZN(n11676) );
  NAND2_X1 U11645 ( .A1(n11679), .A2(n11680), .ZN(n11536) );
  NAND3_X1 U11646 ( .A1(a_18_), .A2(n11681), .A3(b_16_), .ZN(n11680) );
  NAND2_X1 U11647 ( .A1(n11532), .A2(n11531), .ZN(n11681) );
  OR2_X1 U11648 ( .A1(n11531), .A2(n11532), .ZN(n11679) );
  AND2_X1 U11649 ( .A1(n11682), .A2(n11683), .ZN(n11532) );
  NAND2_X1 U11650 ( .A1(n11529), .A2(n11684), .ZN(n11683) );
  OR2_X1 U11651 ( .A1(n11526), .A2(n11528), .ZN(n11684) );
  NOR2_X1 U11652 ( .A1(n11315), .A2(n8045), .ZN(n11529) );
  NAND2_X1 U11653 ( .A1(n11526), .A2(n11528), .ZN(n11682) );
  NAND2_X1 U11654 ( .A1(n11685), .A2(n11686), .ZN(n11528) );
  NAND3_X1 U11655 ( .A1(a_20_), .A2(n11687), .A3(b_16_), .ZN(n11686) );
  NAND2_X1 U11656 ( .A1(n11524), .A2(n11523), .ZN(n11687) );
  OR2_X1 U11657 ( .A1(n11523), .A2(n11524), .ZN(n11685) );
  AND2_X1 U11658 ( .A1(n11688), .A2(n11689), .ZN(n11524) );
  NAND2_X1 U11659 ( .A1(n11521), .A2(n11690), .ZN(n11689) );
  OR2_X1 U11660 ( .A1(n11519), .A2(n11520), .ZN(n11690) );
  NOR2_X1 U11661 ( .A1(n11315), .A2(n7665), .ZN(n11521) );
  NAND2_X1 U11662 ( .A1(n11519), .A2(n11520), .ZN(n11688) );
  NAND2_X1 U11663 ( .A1(n11691), .A2(n11692), .ZN(n11520) );
  NAND3_X1 U11664 ( .A1(a_22_), .A2(n11693), .A3(b_16_), .ZN(n11692) );
  NAND2_X1 U11665 ( .A1(n11516), .A2(n11515), .ZN(n11693) );
  OR2_X1 U11666 ( .A1(n11515), .A2(n11516), .ZN(n11691) );
  AND2_X1 U11667 ( .A1(n11694), .A2(n11695), .ZN(n11516) );
  NAND2_X1 U11668 ( .A1(n11513), .A2(n11696), .ZN(n11695) );
  OR2_X1 U11669 ( .A1(n11510), .A2(n11512), .ZN(n11696) );
  NOR2_X1 U11670 ( .A1(n11315), .A2(n8042), .ZN(n11513) );
  NAND2_X1 U11671 ( .A1(n11510), .A2(n11512), .ZN(n11694) );
  NAND2_X1 U11672 ( .A1(n11697), .A2(n11698), .ZN(n11512) );
  NAND3_X1 U11673 ( .A1(a_24_), .A2(n11699), .A3(b_16_), .ZN(n11698) );
  NAND2_X1 U11674 ( .A1(n11508), .A2(n11507), .ZN(n11699) );
  OR2_X1 U11675 ( .A1(n11507), .A2(n11508), .ZN(n11697) );
  AND2_X1 U11676 ( .A1(n11700), .A2(n11701), .ZN(n11508) );
  NAND2_X1 U11677 ( .A1(n11505), .A2(n11702), .ZN(n11701) );
  OR2_X1 U11678 ( .A1(n11503), .A2(n11504), .ZN(n11702) );
  NOR2_X1 U11679 ( .A1(n11315), .A2(n8039), .ZN(n11505) );
  NAND2_X1 U11680 ( .A1(n11503), .A2(n11504), .ZN(n11700) );
  NAND2_X1 U11681 ( .A1(n11500), .A2(n11703), .ZN(n11504) );
  NAND2_X1 U11682 ( .A1(n11499), .A2(n11501), .ZN(n11703) );
  NAND2_X1 U11683 ( .A1(n11704), .A2(n11705), .ZN(n11501) );
  NAND2_X1 U11684 ( .A1(b_16_), .A2(a_26_), .ZN(n11705) );
  INV_X1 U11685 ( .A(n11706), .ZN(n11704) );
  XNOR2_X1 U11686 ( .A(n11707), .B(n11708), .ZN(n11499) );
  NAND2_X1 U11687 ( .A1(n11709), .A2(n11710), .ZN(n11707) );
  NAND2_X1 U11688 ( .A1(a_26_), .A2(n11706), .ZN(n11500) );
  NAND2_X1 U11689 ( .A1(n11472), .A2(n11711), .ZN(n11706) );
  NAND2_X1 U11690 ( .A1(n11471), .A2(n11473), .ZN(n11711) );
  NAND2_X1 U11691 ( .A1(n11712), .A2(n11713), .ZN(n11473) );
  NAND2_X1 U11692 ( .A1(b_16_), .A2(a_27_), .ZN(n11713) );
  INV_X1 U11693 ( .A(n11714), .ZN(n11712) );
  XNOR2_X1 U11694 ( .A(n11715), .B(n11716), .ZN(n11471) );
  XOR2_X1 U11695 ( .A(n11717), .B(n11718), .Z(n11715) );
  NAND2_X1 U11696 ( .A1(b_15_), .A2(a_28_), .ZN(n11717) );
  NAND2_X1 U11697 ( .A1(a_27_), .A2(n11714), .ZN(n11472) );
  NAND2_X1 U11698 ( .A1(n11719), .A2(n11720), .ZN(n11714) );
  NAND3_X1 U11699 ( .A1(a_28_), .A2(n11721), .A3(b_16_), .ZN(n11720) );
  NAND2_X1 U11700 ( .A1(n11481), .A2(n11479), .ZN(n11721) );
  OR2_X1 U11701 ( .A1(n11479), .A2(n11481), .ZN(n11719) );
  AND2_X1 U11702 ( .A1(n11722), .A2(n11723), .ZN(n11481) );
  NAND2_X1 U11703 ( .A1(n11495), .A2(n11724), .ZN(n11723) );
  OR2_X1 U11704 ( .A1(n11496), .A2(n11497), .ZN(n11724) );
  NOR2_X1 U11705 ( .A1(n11315), .A2(n7545), .ZN(n11495) );
  NAND2_X1 U11706 ( .A1(n11497), .A2(n11496), .ZN(n11722) );
  NAND2_X1 U11707 ( .A1(n11725), .A2(n11726), .ZN(n11496) );
  NAND2_X1 U11708 ( .A1(b_14_), .A2(n11727), .ZN(n11726) );
  NAND2_X1 U11709 ( .A1(n7527), .A2(n11728), .ZN(n11727) );
  NAND2_X1 U11710 ( .A1(a_31_), .A2(n7756), .ZN(n11728) );
  NAND2_X1 U11711 ( .A1(b_15_), .A2(n11729), .ZN(n11725) );
  NAND2_X1 U11712 ( .A1(n7531), .A2(n11730), .ZN(n11729) );
  NAND2_X1 U11713 ( .A1(a_30_), .A2(n8048), .ZN(n11730) );
  AND3_X1 U11714 ( .A1(b_16_), .A2(b_15_), .A3(n7494), .ZN(n11497) );
  XNOR2_X1 U11715 ( .A(n11731), .B(n11732), .ZN(n11479) );
  XOR2_X1 U11716 ( .A(n11733), .B(n11734), .Z(n11731) );
  XNOR2_X1 U11717 ( .A(n11735), .B(n11736), .ZN(n11503) );
  NAND2_X1 U11718 ( .A1(n11737), .A2(n11738), .ZN(n11735) );
  XNOR2_X1 U11719 ( .A(n11739), .B(n11740), .ZN(n11507) );
  XOR2_X1 U11720 ( .A(n11741), .B(n11742), .Z(n11739) );
  XNOR2_X1 U11721 ( .A(n11743), .B(n11744), .ZN(n11510) );
  XNOR2_X1 U11722 ( .A(n11745), .B(n11746), .ZN(n11743) );
  NOR2_X1 U11723 ( .A1(n8041), .A2(n7756), .ZN(n11746) );
  XOR2_X1 U11724 ( .A(n11747), .B(n11748), .Z(n11515) );
  XNOR2_X1 U11725 ( .A(n11749), .B(n11750), .ZN(n11748) );
  XNOR2_X1 U11726 ( .A(n11751), .B(n11752), .ZN(n11519) );
  XNOR2_X1 U11727 ( .A(n11753), .B(n11754), .ZN(n11751) );
  NOR2_X1 U11728 ( .A1(n7650), .A2(n7756), .ZN(n11754) );
  XNOR2_X1 U11729 ( .A(n11755), .B(n11756), .ZN(n11523) );
  XOR2_X1 U11730 ( .A(n11757), .B(n11758), .Z(n11755) );
  XNOR2_X1 U11731 ( .A(n11759), .B(n11760), .ZN(n11526) );
  XNOR2_X1 U11732 ( .A(n11761), .B(n11762), .ZN(n11759) );
  NOR2_X1 U11733 ( .A1(n8044), .A2(n7756), .ZN(n11762) );
  XOR2_X1 U11734 ( .A(n11763), .B(n11764), .Z(n11531) );
  XNOR2_X1 U11735 ( .A(n11765), .B(n11766), .ZN(n11764) );
  XNOR2_X1 U11736 ( .A(n11767), .B(n11768), .ZN(n11535) );
  XNOR2_X1 U11737 ( .A(n11769), .B(n11770), .ZN(n11767) );
  NOR2_X1 U11738 ( .A1(n8047), .A2(n7756), .ZN(n11770) );
  NOR2_X1 U11739 ( .A1(n11315), .A2(n8438), .ZN(n7744) );
  XNOR2_X1 U11740 ( .A(n11771), .B(n11772), .ZN(n11546) );
  XOR2_X1 U11741 ( .A(n8003), .B(n11773), .Z(n11772) );
  XOR2_X1 U11742 ( .A(n11774), .B(n11775), .Z(n11550) );
  NAND2_X1 U11743 ( .A1(n11776), .A2(n11777), .ZN(n11774) );
  XOR2_X1 U11744 ( .A(n11778), .B(n11779), .Z(n11554) );
  XOR2_X1 U11745 ( .A(n11780), .B(n11781), .Z(n11779) );
  NAND2_X1 U11746 ( .A1(a_13_), .A2(b_15_), .ZN(n11781) );
  XNOR2_X1 U11747 ( .A(n11782), .B(n11783), .ZN(n11558) );
  XOR2_X1 U11748 ( .A(n11784), .B(n11785), .Z(n11783) );
  NAND2_X1 U11749 ( .A1(a_12_), .A2(b_15_), .ZN(n11785) );
  XNOR2_X1 U11750 ( .A(n11786), .B(n11787), .ZN(n11562) );
  XNOR2_X1 U11751 ( .A(n11788), .B(n11789), .ZN(n11786) );
  NOR2_X1 U11752 ( .A1(n7756), .A2(n7811), .ZN(n11789) );
  XNOR2_X1 U11753 ( .A(n11790), .B(n11791), .ZN(n11565) );
  XOR2_X1 U11754 ( .A(n11792), .B(n11793), .Z(n11791) );
  NAND2_X1 U11755 ( .A1(a_10_), .A2(b_15_), .ZN(n11793) );
  XOR2_X1 U11756 ( .A(n11794), .B(n11795), .Z(n11570) );
  XOR2_X1 U11757 ( .A(n11796), .B(n11797), .Z(n11795) );
  NAND2_X1 U11758 ( .A1(a_9_), .A2(b_15_), .ZN(n11797) );
  XNOR2_X1 U11759 ( .A(n11798), .B(n11799), .ZN(n11573) );
  XNOR2_X1 U11760 ( .A(n11800), .B(n11801), .ZN(n11798) );
  NOR2_X1 U11761 ( .A1(n7756), .A2(n8686), .ZN(n11801) );
  XOR2_X1 U11762 ( .A(n11802), .B(n11803), .Z(n11577) );
  XOR2_X1 U11763 ( .A(n11804), .B(n11805), .Z(n11802) );
  NOR2_X1 U11764 ( .A1(n7756), .A2(n7872), .ZN(n11805) );
  XNOR2_X1 U11765 ( .A(n11806), .B(n11807), .ZN(n11586) );
  XNOR2_X1 U11766 ( .A(n11808), .B(n11809), .ZN(n11806) );
  NAND2_X1 U11767 ( .A1(a_5_), .A2(b_15_), .ZN(n11808) );
  XNOR2_X1 U11768 ( .A(n11810), .B(n11811), .ZN(n11590) );
  XNOR2_X1 U11769 ( .A(n11812), .B(n11813), .ZN(n11810) );
  NOR2_X1 U11770 ( .A1(n7756), .A2(n7916), .ZN(n11813) );
  XNOR2_X1 U11771 ( .A(n11814), .B(n11815), .ZN(n11594) );
  XOR2_X1 U11772 ( .A(n11816), .B(n11817), .Z(n11815) );
  NAND2_X1 U11773 ( .A1(a_3_), .A2(b_15_), .ZN(n11817) );
  XNOR2_X1 U11774 ( .A(n11818), .B(n11819), .ZN(n11598) );
  XOR2_X1 U11775 ( .A(n11820), .B(n11821), .Z(n11818) );
  NOR2_X1 U11776 ( .A1(n7756), .A2(n8056), .ZN(n11821) );
  XNOR2_X1 U11777 ( .A(n11822), .B(n11823), .ZN(n11601) );
  XOR2_X1 U11778 ( .A(n11824), .B(n11825), .Z(n11823) );
  NAND2_X1 U11779 ( .A1(b_15_), .A2(a_1_), .ZN(n11825) );
  XNOR2_X1 U11780 ( .A(n11826), .B(n11827), .ZN(n8218) );
  XOR2_X1 U11781 ( .A(n11828), .B(n11829), .Z(n11827) );
  NAND2_X1 U11782 ( .A1(a_0_), .A2(b_15_), .ZN(n11829) );
  NAND2_X1 U11783 ( .A1(n11830), .A2(n11831), .ZN(n8152) );
  NAND2_X1 U11784 ( .A1(n11610), .A2(n11607), .ZN(n11831) );
  XNOR2_X1 U11785 ( .A(n8209), .B(n8208), .ZN(n11830) );
  NAND3_X1 U11786 ( .A1(n11610), .A2(n11607), .A3(n11832), .ZN(n8151) );
  XOR2_X1 U11787 ( .A(n8209), .B(n8208), .Z(n11832) );
  NAND2_X1 U11788 ( .A1(n11833), .A2(n11834), .ZN(n11607) );
  NAND3_X1 U11789 ( .A1(b_15_), .A2(n11835), .A3(a_0_), .ZN(n11834) );
  OR2_X1 U11790 ( .A1(n11828), .A2(n11826), .ZN(n11835) );
  NAND2_X1 U11791 ( .A1(n11826), .A2(n11828), .ZN(n11833) );
  NAND2_X1 U11792 ( .A1(n11836), .A2(n11837), .ZN(n11828) );
  NAND3_X1 U11793 ( .A1(a_1_), .A2(n11838), .A3(b_15_), .ZN(n11837) );
  OR2_X1 U11794 ( .A1(n11822), .A2(n11824), .ZN(n11838) );
  NAND2_X1 U11795 ( .A1(n11822), .A2(n11824), .ZN(n11836) );
  NAND2_X1 U11796 ( .A1(n11839), .A2(n11840), .ZN(n11824) );
  NAND3_X1 U11797 ( .A1(b_15_), .A2(n11841), .A3(a_2_), .ZN(n11840) );
  OR2_X1 U11798 ( .A1(n11819), .A2(n11820), .ZN(n11841) );
  NAND2_X1 U11799 ( .A1(n11819), .A2(n11820), .ZN(n11839) );
  NAND2_X1 U11800 ( .A1(n11842), .A2(n11843), .ZN(n11820) );
  NAND3_X1 U11801 ( .A1(b_15_), .A2(n11844), .A3(a_3_), .ZN(n11843) );
  OR2_X1 U11802 ( .A1(n11816), .A2(n11814), .ZN(n11844) );
  NAND2_X1 U11803 ( .A1(n11814), .A2(n11816), .ZN(n11842) );
  NAND2_X1 U11804 ( .A1(n11845), .A2(n11846), .ZN(n11816) );
  NAND3_X1 U11805 ( .A1(b_15_), .A2(n11847), .A3(a_4_), .ZN(n11846) );
  NAND2_X1 U11806 ( .A1(n11812), .A2(n11811), .ZN(n11847) );
  OR2_X1 U11807 ( .A1(n11811), .A2(n11812), .ZN(n11845) );
  AND2_X1 U11808 ( .A1(n11848), .A2(n11849), .ZN(n11812) );
  NAND3_X1 U11809 ( .A1(b_15_), .A2(n11850), .A3(a_5_), .ZN(n11849) );
  OR2_X1 U11810 ( .A1(n11807), .A2(n11809), .ZN(n11850) );
  NAND2_X1 U11811 ( .A1(n11807), .A2(n11809), .ZN(n11848) );
  NAND2_X1 U11812 ( .A1(n11851), .A2(n11852), .ZN(n11809) );
  NAND3_X1 U11813 ( .A1(b_15_), .A2(n11853), .A3(a_6_), .ZN(n11852) );
  OR2_X1 U11814 ( .A1(n11631), .A2(n11632), .ZN(n11853) );
  NAND2_X1 U11815 ( .A1(n11631), .A2(n11632), .ZN(n11851) );
  NAND2_X1 U11816 ( .A1(n11854), .A2(n11855), .ZN(n11632) );
  NAND3_X1 U11817 ( .A1(b_15_), .A2(n11856), .A3(a_7_), .ZN(n11855) );
  OR2_X1 U11818 ( .A1(n11803), .A2(n11804), .ZN(n11856) );
  NAND2_X1 U11819 ( .A1(n11803), .A2(n11804), .ZN(n11854) );
  NAND2_X1 U11820 ( .A1(n11857), .A2(n11858), .ZN(n11804) );
  NAND3_X1 U11821 ( .A1(b_15_), .A2(n11859), .A3(a_8_), .ZN(n11858) );
  NAND2_X1 U11822 ( .A1(n11800), .A2(n11799), .ZN(n11859) );
  OR2_X1 U11823 ( .A1(n11799), .A2(n11800), .ZN(n11857) );
  AND2_X1 U11824 ( .A1(n11860), .A2(n11861), .ZN(n11800) );
  NAND3_X1 U11825 ( .A1(b_15_), .A2(n11862), .A3(a_9_), .ZN(n11861) );
  OR2_X1 U11826 ( .A1(n11794), .A2(n11796), .ZN(n11862) );
  NAND2_X1 U11827 ( .A1(n11794), .A2(n11796), .ZN(n11860) );
  NAND2_X1 U11828 ( .A1(n11863), .A2(n11864), .ZN(n11796) );
  NAND3_X1 U11829 ( .A1(b_15_), .A2(n11865), .A3(a_10_), .ZN(n11864) );
  OR2_X1 U11830 ( .A1(n11790), .A2(n11792), .ZN(n11865) );
  NAND2_X1 U11831 ( .A1(n11790), .A2(n11792), .ZN(n11863) );
  NAND2_X1 U11832 ( .A1(n11866), .A2(n11867), .ZN(n11792) );
  NAND3_X1 U11833 ( .A1(b_15_), .A2(n11868), .A3(a_11_), .ZN(n11867) );
  NAND2_X1 U11834 ( .A1(n11788), .A2(n11787), .ZN(n11868) );
  OR2_X1 U11835 ( .A1(n11787), .A2(n11788), .ZN(n11866) );
  AND2_X1 U11836 ( .A1(n11869), .A2(n11870), .ZN(n11788) );
  NAND3_X1 U11837 ( .A1(b_15_), .A2(n11871), .A3(a_12_), .ZN(n11870) );
  OR2_X1 U11838 ( .A1(n11784), .A2(n11782), .ZN(n11871) );
  NAND2_X1 U11839 ( .A1(n11782), .A2(n11784), .ZN(n11869) );
  NAND2_X1 U11840 ( .A1(n11872), .A2(n11873), .ZN(n11784) );
  NAND3_X1 U11841 ( .A1(b_15_), .A2(n11874), .A3(a_13_), .ZN(n11873) );
  OR2_X1 U11842 ( .A1(n11778), .A2(n11780), .ZN(n11874) );
  NAND2_X1 U11843 ( .A1(n11778), .A2(n11780), .ZN(n11872) );
  NAND2_X1 U11844 ( .A1(n11776), .A2(n11875), .ZN(n11780) );
  NAND2_X1 U11845 ( .A1(n11775), .A2(n11777), .ZN(n11875) );
  NAND2_X1 U11846 ( .A1(n11876), .A2(n11877), .ZN(n11777) );
  NAND2_X1 U11847 ( .A1(a_14_), .A2(b_15_), .ZN(n11877) );
  INV_X1 U11848 ( .A(n11878), .ZN(n11876) );
  XOR2_X1 U11849 ( .A(n11879), .B(n11880), .Z(n11775) );
  XOR2_X1 U11850 ( .A(n11881), .B(n11882), .Z(n11879) );
  NAND2_X1 U11851 ( .A1(a_14_), .A2(n11878), .ZN(n11776) );
  NAND2_X1 U11852 ( .A1(n11883), .A2(n11884), .ZN(n11878) );
  NAND2_X1 U11853 ( .A1(n11771), .A2(n11885), .ZN(n11884) );
  OR2_X1 U11854 ( .A1(n11773), .A2(n7751), .ZN(n11885) );
  XNOR2_X1 U11855 ( .A(n11886), .B(n11887), .ZN(n11771) );
  XNOR2_X1 U11856 ( .A(n11888), .B(n11889), .ZN(n11887) );
  NAND2_X1 U11857 ( .A1(n7751), .A2(n11773), .ZN(n11883) );
  NAND2_X1 U11858 ( .A1(n11890), .A2(n11891), .ZN(n11773) );
  NAND3_X1 U11859 ( .A1(a_16_), .A2(n11892), .A3(b_15_), .ZN(n11891) );
  OR2_X1 U11860 ( .A1(n11667), .A2(n11665), .ZN(n11892) );
  NAND2_X1 U11861 ( .A1(n11665), .A2(n11667), .ZN(n11890) );
  NAND2_X1 U11862 ( .A1(n11893), .A2(n11894), .ZN(n11667) );
  NAND2_X1 U11863 ( .A1(n11675), .A2(n11895), .ZN(n11894) );
  OR2_X1 U11864 ( .A1(n11673), .A2(n11674), .ZN(n11895) );
  NOR2_X1 U11865 ( .A1(n7756), .A2(n7732), .ZN(n11675) );
  NAND2_X1 U11866 ( .A1(n11673), .A2(n11674), .ZN(n11893) );
  NAND2_X1 U11867 ( .A1(n11896), .A2(n11897), .ZN(n11674) );
  NAND3_X1 U11868 ( .A1(a_18_), .A2(n11898), .A3(b_15_), .ZN(n11897) );
  NAND2_X1 U11869 ( .A1(n11769), .A2(n11768), .ZN(n11898) );
  OR2_X1 U11870 ( .A1(n11768), .A2(n11769), .ZN(n11896) );
  AND2_X1 U11871 ( .A1(n11899), .A2(n11900), .ZN(n11769) );
  NAND2_X1 U11872 ( .A1(n11766), .A2(n11901), .ZN(n11900) );
  OR2_X1 U11873 ( .A1(n11763), .A2(n11765), .ZN(n11901) );
  NOR2_X1 U11874 ( .A1(n7756), .A2(n8045), .ZN(n11766) );
  NAND2_X1 U11875 ( .A1(n11763), .A2(n11765), .ZN(n11899) );
  NAND2_X1 U11876 ( .A1(n11902), .A2(n11903), .ZN(n11765) );
  NAND3_X1 U11877 ( .A1(a_20_), .A2(n11904), .A3(b_15_), .ZN(n11903) );
  NAND2_X1 U11878 ( .A1(n11761), .A2(n11760), .ZN(n11904) );
  OR2_X1 U11879 ( .A1(n11760), .A2(n11761), .ZN(n11902) );
  AND2_X1 U11880 ( .A1(n11905), .A2(n11906), .ZN(n11761) );
  NAND2_X1 U11881 ( .A1(n11758), .A2(n11907), .ZN(n11906) );
  OR2_X1 U11882 ( .A1(n11756), .A2(n11757), .ZN(n11907) );
  NOR2_X1 U11883 ( .A1(n7756), .A2(n7665), .ZN(n11758) );
  NAND2_X1 U11884 ( .A1(n11756), .A2(n11757), .ZN(n11905) );
  NAND2_X1 U11885 ( .A1(n11908), .A2(n11909), .ZN(n11757) );
  NAND3_X1 U11886 ( .A1(a_22_), .A2(n11910), .A3(b_15_), .ZN(n11909) );
  NAND2_X1 U11887 ( .A1(n11753), .A2(n11752), .ZN(n11910) );
  OR2_X1 U11888 ( .A1(n11752), .A2(n11753), .ZN(n11908) );
  AND2_X1 U11889 ( .A1(n11911), .A2(n11912), .ZN(n11753) );
  NAND2_X1 U11890 ( .A1(n11750), .A2(n11913), .ZN(n11912) );
  OR2_X1 U11891 ( .A1(n11747), .A2(n11749), .ZN(n11913) );
  NOR2_X1 U11892 ( .A1(n7756), .A2(n8042), .ZN(n11750) );
  NAND2_X1 U11893 ( .A1(n11747), .A2(n11749), .ZN(n11911) );
  NAND2_X1 U11894 ( .A1(n11914), .A2(n11915), .ZN(n11749) );
  NAND3_X1 U11895 ( .A1(a_24_), .A2(n11916), .A3(b_15_), .ZN(n11915) );
  NAND2_X1 U11896 ( .A1(n11745), .A2(n11744), .ZN(n11916) );
  OR2_X1 U11897 ( .A1(n11744), .A2(n11745), .ZN(n11914) );
  AND2_X1 U11898 ( .A1(n11917), .A2(n11918), .ZN(n11745) );
  NAND2_X1 U11899 ( .A1(n11742), .A2(n11919), .ZN(n11918) );
  OR2_X1 U11900 ( .A1(n11740), .A2(n11741), .ZN(n11919) );
  NOR2_X1 U11901 ( .A1(n7756), .A2(n8039), .ZN(n11742) );
  NAND2_X1 U11902 ( .A1(n11740), .A2(n11741), .ZN(n11917) );
  NAND2_X1 U11903 ( .A1(n11737), .A2(n11920), .ZN(n11741) );
  NAND2_X1 U11904 ( .A1(n11736), .A2(n11738), .ZN(n11920) );
  NAND2_X1 U11905 ( .A1(n11921), .A2(n11922), .ZN(n11738) );
  NAND2_X1 U11906 ( .A1(b_15_), .A2(a_26_), .ZN(n11922) );
  INV_X1 U11907 ( .A(n11923), .ZN(n11921) );
  XNOR2_X1 U11908 ( .A(n11924), .B(n11925), .ZN(n11736) );
  NAND2_X1 U11909 ( .A1(n11926), .A2(n11927), .ZN(n11924) );
  NAND2_X1 U11910 ( .A1(a_26_), .A2(n11923), .ZN(n11737) );
  NAND2_X1 U11911 ( .A1(n11709), .A2(n11928), .ZN(n11923) );
  NAND2_X1 U11912 ( .A1(n11708), .A2(n11710), .ZN(n11928) );
  NAND2_X1 U11913 ( .A1(n11929), .A2(n11930), .ZN(n11710) );
  NAND2_X1 U11914 ( .A1(b_15_), .A2(a_27_), .ZN(n11930) );
  INV_X1 U11915 ( .A(n11931), .ZN(n11929) );
  XNOR2_X1 U11916 ( .A(n11932), .B(n11933), .ZN(n11708) );
  XOR2_X1 U11917 ( .A(n11934), .B(n11935), .Z(n11932) );
  NAND2_X1 U11918 ( .A1(b_14_), .A2(a_28_), .ZN(n11934) );
  NAND2_X1 U11919 ( .A1(a_27_), .A2(n11931), .ZN(n11709) );
  NAND2_X1 U11920 ( .A1(n11936), .A2(n11937), .ZN(n11931) );
  NAND3_X1 U11921 ( .A1(a_28_), .A2(n11938), .A3(b_15_), .ZN(n11937) );
  NAND2_X1 U11922 ( .A1(n11718), .A2(n11716), .ZN(n11938) );
  OR2_X1 U11923 ( .A1(n11716), .A2(n11718), .ZN(n11936) );
  AND2_X1 U11924 ( .A1(n11939), .A2(n11940), .ZN(n11718) );
  NAND2_X1 U11925 ( .A1(n11732), .A2(n11941), .ZN(n11940) );
  OR2_X1 U11926 ( .A1(n11733), .A2(n11734), .ZN(n11941) );
  NOR2_X1 U11927 ( .A1(n7756), .A2(n7545), .ZN(n11732) );
  NAND2_X1 U11928 ( .A1(n11734), .A2(n11733), .ZN(n11939) );
  NAND2_X1 U11929 ( .A1(n11942), .A2(n11943), .ZN(n11733) );
  NAND2_X1 U11930 ( .A1(b_13_), .A2(n11944), .ZN(n11943) );
  NAND2_X1 U11931 ( .A1(n7527), .A2(n11945), .ZN(n11944) );
  NAND2_X1 U11932 ( .A1(a_31_), .A2(n8048), .ZN(n11945) );
  NAND2_X1 U11933 ( .A1(b_14_), .A2(n11946), .ZN(n11942) );
  NAND2_X1 U11934 ( .A1(n7531), .A2(n11947), .ZN(n11946) );
  NAND2_X1 U11935 ( .A1(a_30_), .A2(n7782), .ZN(n11947) );
  AND3_X1 U11936 ( .A1(b_14_), .A2(b_15_), .A3(n7494), .ZN(n11734) );
  XNOR2_X1 U11937 ( .A(n11948), .B(n11949), .ZN(n11716) );
  XOR2_X1 U11938 ( .A(n11950), .B(n11951), .Z(n11948) );
  XNOR2_X1 U11939 ( .A(n11952), .B(n11953), .ZN(n11740) );
  NAND2_X1 U11940 ( .A1(n11954), .A2(n11955), .ZN(n11952) );
  XNOR2_X1 U11941 ( .A(n11956), .B(n11957), .ZN(n11744) );
  XOR2_X1 U11942 ( .A(n11958), .B(n11959), .Z(n11956) );
  XNOR2_X1 U11943 ( .A(n11960), .B(n11961), .ZN(n11747) );
  XNOR2_X1 U11944 ( .A(n11962), .B(n11963), .ZN(n11960) );
  NOR2_X1 U11945 ( .A1(n8041), .A2(n8048), .ZN(n11963) );
  XOR2_X1 U11946 ( .A(n11964), .B(n11965), .Z(n11752) );
  XNOR2_X1 U11947 ( .A(n11966), .B(n11967), .ZN(n11965) );
  XNOR2_X1 U11948 ( .A(n11968), .B(n11969), .ZN(n11756) );
  XOR2_X1 U11949 ( .A(n11970), .B(n11971), .Z(n11969) );
  NAND2_X1 U11950 ( .A1(b_14_), .A2(a_22_), .ZN(n11971) );
  XNOR2_X1 U11951 ( .A(n11972), .B(n11973), .ZN(n11760) );
  XOR2_X1 U11952 ( .A(n11974), .B(n11975), .Z(n11972) );
  XNOR2_X1 U11953 ( .A(n11976), .B(n11977), .ZN(n11763) );
  XNOR2_X1 U11954 ( .A(n11978), .B(n11979), .ZN(n11976) );
  NOR2_X1 U11955 ( .A1(n8044), .A2(n8048), .ZN(n11979) );
  XOR2_X1 U11956 ( .A(n11980), .B(n11981), .Z(n11768) );
  XNOR2_X1 U11957 ( .A(n11982), .B(n11983), .ZN(n11981) );
  XNOR2_X1 U11958 ( .A(n11984), .B(n11985), .ZN(n11673) );
  XNOR2_X1 U11959 ( .A(n11986), .B(n11987), .ZN(n11984) );
  NOR2_X1 U11960 ( .A1(n8047), .A2(n8048), .ZN(n11987) );
  XOR2_X1 U11961 ( .A(n11988), .B(n11989), .Z(n11665) );
  XOR2_X1 U11962 ( .A(n11990), .B(n11991), .Z(n11988) );
  NOR2_X1 U11963 ( .A1(n7732), .A2(n8048), .ZN(n11991) );
  INV_X1 U11964 ( .A(n8003), .ZN(n7751) );
  NAND2_X1 U11965 ( .A1(a_15_), .A2(b_15_), .ZN(n8003) );
  XOR2_X1 U11966 ( .A(n11992), .B(n11993), .Z(n11778) );
  XOR2_X1 U11967 ( .A(n11994), .B(n11995), .Z(n11992) );
  XNOR2_X1 U11968 ( .A(n11996), .B(n11997), .ZN(n11782) );
  NAND2_X1 U11969 ( .A1(n11998), .A2(n11999), .ZN(n11996) );
  XNOR2_X1 U11970 ( .A(n12000), .B(n12001), .ZN(n11787) );
  XOR2_X1 U11971 ( .A(n12002), .B(n12003), .Z(n12000) );
  XNOR2_X1 U11972 ( .A(n12004), .B(n12005), .ZN(n11790) );
  XNOR2_X1 U11973 ( .A(n12006), .B(n12007), .ZN(n12004) );
  NOR2_X1 U11974 ( .A1(n8048), .A2(n7811), .ZN(n12007) );
  XNOR2_X1 U11975 ( .A(n12008), .B(n12009), .ZN(n11794) );
  XNOR2_X1 U11976 ( .A(n12010), .B(n12011), .ZN(n12008) );
  XOR2_X1 U11977 ( .A(n12012), .B(n12013), .Z(n11799) );
  XOR2_X1 U11978 ( .A(n12014), .B(n12015), .Z(n12013) );
  NAND2_X1 U11979 ( .A1(a_9_), .A2(b_14_), .ZN(n12015) );
  XNOR2_X1 U11980 ( .A(n12016), .B(n12017), .ZN(n11803) );
  NAND2_X1 U11981 ( .A1(n12018), .A2(n12019), .ZN(n12016) );
  XNOR2_X1 U11982 ( .A(n12020), .B(n12021), .ZN(n11631) );
  NAND2_X1 U11983 ( .A1(n12022), .A2(n12023), .ZN(n12020) );
  XNOR2_X1 U11984 ( .A(n12024), .B(n12025), .ZN(n11807) );
  NAND2_X1 U11985 ( .A1(n12026), .A2(n12027), .ZN(n12024) );
  XOR2_X1 U11986 ( .A(n12028), .B(n12029), .Z(n11811) );
  NAND2_X1 U11987 ( .A1(n12030), .A2(n12031), .ZN(n12028) );
  XNOR2_X1 U11988 ( .A(n12032), .B(n12033), .ZN(n11814) );
  XNOR2_X1 U11989 ( .A(n12034), .B(n12035), .ZN(n12033) );
  XNOR2_X1 U11990 ( .A(n12036), .B(n12037), .ZN(n11819) );
  XNOR2_X1 U11991 ( .A(n12038), .B(n12039), .ZN(n12037) );
  XNOR2_X1 U11992 ( .A(n12040), .B(n12041), .ZN(n11822) );
  XNOR2_X1 U11993 ( .A(n12042), .B(n12043), .ZN(n12040) );
  NOR2_X1 U11994 ( .A1(n8048), .A2(n8056), .ZN(n12043) );
  XNOR2_X1 U11995 ( .A(n12044), .B(n12045), .ZN(n11826) );
  XNOR2_X1 U11996 ( .A(n12046), .B(n12047), .ZN(n12045) );
  INV_X1 U11997 ( .A(n11608), .ZN(n11610) );
  XOR2_X1 U11998 ( .A(n12048), .B(n12049), .Z(n11608) );
  XOR2_X1 U11999 ( .A(n12050), .B(n12051), .Z(n12049) );
  NAND2_X1 U12000 ( .A1(a_0_), .A2(b_14_), .ZN(n12051) );
  NAND4_X1 U12001 ( .A1(n8208), .A2(n8207), .A3(n8209), .A4(n8203), .ZN(n8156)
         );
  INV_X1 U12002 ( .A(n12052), .ZN(n8203) );
  NAND2_X1 U12003 ( .A1(n12053), .A2(n12054), .ZN(n8209) );
  NAND3_X1 U12004 ( .A1(b_14_), .A2(n12055), .A3(a_0_), .ZN(n12054) );
  OR2_X1 U12005 ( .A1(n12050), .A2(n12048), .ZN(n12055) );
  NAND2_X1 U12006 ( .A1(n12048), .A2(n12050), .ZN(n12053) );
  NAND2_X1 U12007 ( .A1(n12056), .A2(n12057), .ZN(n12050) );
  NAND2_X1 U12008 ( .A1(n12047), .A2(n12058), .ZN(n12057) );
  OR2_X1 U12009 ( .A1(n12046), .A2(n12044), .ZN(n12058) );
  NOR2_X1 U12010 ( .A1(n8048), .A2(n7957), .ZN(n12047) );
  NAND2_X1 U12011 ( .A1(n12044), .A2(n12046), .ZN(n12056) );
  NAND2_X1 U12012 ( .A1(n12059), .A2(n12060), .ZN(n12046) );
  NAND3_X1 U12013 ( .A1(b_14_), .A2(n12061), .A3(a_2_), .ZN(n12060) );
  NAND2_X1 U12014 ( .A1(n12042), .A2(n12041), .ZN(n12061) );
  OR2_X1 U12015 ( .A1(n12041), .A2(n12042), .ZN(n12059) );
  AND2_X1 U12016 ( .A1(n12062), .A2(n12063), .ZN(n12042) );
  NAND2_X1 U12017 ( .A1(n12039), .A2(n12064), .ZN(n12063) );
  OR2_X1 U12018 ( .A1(n12038), .A2(n12036), .ZN(n12064) );
  NOR2_X1 U12019 ( .A1(n7937), .A2(n8048), .ZN(n12039) );
  NAND2_X1 U12020 ( .A1(n12036), .A2(n12038), .ZN(n12062) );
  NAND2_X1 U12021 ( .A1(n12065), .A2(n12066), .ZN(n12038) );
  NAND2_X1 U12022 ( .A1(n12035), .A2(n12067), .ZN(n12066) );
  OR2_X1 U12023 ( .A1(n12034), .A2(n12032), .ZN(n12067) );
  NOR2_X1 U12024 ( .A1(n7916), .A2(n8048), .ZN(n12035) );
  NAND2_X1 U12025 ( .A1(n12032), .A2(n12034), .ZN(n12065) );
  NAND2_X1 U12026 ( .A1(n12030), .A2(n12068), .ZN(n12034) );
  NAND2_X1 U12027 ( .A1(n12029), .A2(n12031), .ZN(n12068) );
  NAND2_X1 U12028 ( .A1(n12069), .A2(n12070), .ZN(n12031) );
  NAND2_X1 U12029 ( .A1(a_5_), .A2(b_14_), .ZN(n12070) );
  INV_X1 U12030 ( .A(n12071), .ZN(n12069) );
  XNOR2_X1 U12031 ( .A(n12072), .B(n12073), .ZN(n12029) );
  XOR2_X1 U12032 ( .A(n12074), .B(n12075), .Z(n12073) );
  NAND2_X1 U12033 ( .A1(a_6_), .A2(b_13_), .ZN(n12075) );
  NAND2_X1 U12034 ( .A1(a_5_), .A2(n12071), .ZN(n12030) );
  NAND2_X1 U12035 ( .A1(n12026), .A2(n12076), .ZN(n12071) );
  NAND2_X1 U12036 ( .A1(n12025), .A2(n12027), .ZN(n12076) );
  NAND2_X1 U12037 ( .A1(n12077), .A2(n12078), .ZN(n12027) );
  NAND2_X1 U12038 ( .A1(a_6_), .A2(b_14_), .ZN(n12078) );
  INV_X1 U12039 ( .A(n12079), .ZN(n12077) );
  XNOR2_X1 U12040 ( .A(n12080), .B(n12081), .ZN(n12025) );
  XOR2_X1 U12041 ( .A(n12082), .B(n12083), .Z(n12081) );
  NAND2_X1 U12042 ( .A1(a_7_), .A2(b_13_), .ZN(n12083) );
  NAND2_X1 U12043 ( .A1(a_6_), .A2(n12079), .ZN(n12026) );
  NAND2_X1 U12044 ( .A1(n12022), .A2(n12084), .ZN(n12079) );
  NAND2_X1 U12045 ( .A1(n12021), .A2(n12023), .ZN(n12084) );
  NAND2_X1 U12046 ( .A1(n12085), .A2(n12086), .ZN(n12023) );
  NAND2_X1 U12047 ( .A1(a_7_), .A2(b_14_), .ZN(n12086) );
  INV_X1 U12048 ( .A(n12087), .ZN(n12085) );
  XNOR2_X1 U12049 ( .A(n12088), .B(n12089), .ZN(n12021) );
  XNOR2_X1 U12050 ( .A(n12090), .B(n12091), .ZN(n12088) );
  NOR2_X1 U12051 ( .A1(n7782), .A2(n8686), .ZN(n12091) );
  NAND2_X1 U12052 ( .A1(a_7_), .A2(n12087), .ZN(n12022) );
  NAND2_X1 U12053 ( .A1(n12018), .A2(n12092), .ZN(n12087) );
  NAND2_X1 U12054 ( .A1(n12017), .A2(n12019), .ZN(n12092) );
  NAND2_X1 U12055 ( .A1(n12093), .A2(n12094), .ZN(n12019) );
  NAND2_X1 U12056 ( .A1(a_8_), .A2(b_14_), .ZN(n12094) );
  INV_X1 U12057 ( .A(n12095), .ZN(n12093) );
  XNOR2_X1 U12058 ( .A(n12096), .B(n12097), .ZN(n12017) );
  XOR2_X1 U12059 ( .A(n12098), .B(n12099), .Z(n12097) );
  NAND2_X1 U12060 ( .A1(a_9_), .A2(b_13_), .ZN(n12099) );
  NAND2_X1 U12061 ( .A1(a_8_), .A2(n12095), .ZN(n12018) );
  NAND2_X1 U12062 ( .A1(n12100), .A2(n12101), .ZN(n12095) );
  NAND3_X1 U12063 ( .A1(b_14_), .A2(n12102), .A3(a_9_), .ZN(n12101) );
  OR2_X1 U12064 ( .A1(n12014), .A2(n12012), .ZN(n12102) );
  NAND2_X1 U12065 ( .A1(n12012), .A2(n12014), .ZN(n12100) );
  NAND2_X1 U12066 ( .A1(n12103), .A2(n12104), .ZN(n12014) );
  NAND2_X1 U12067 ( .A1(n12011), .A2(n12105), .ZN(n12104) );
  NAND2_X1 U12068 ( .A1(n12010), .A2(n12009), .ZN(n12105) );
  NOR2_X1 U12069 ( .A1(n8051), .A2(n8048), .ZN(n12011) );
  OR2_X1 U12070 ( .A1(n12009), .A2(n12010), .ZN(n12103) );
  AND2_X1 U12071 ( .A1(n12106), .A2(n12107), .ZN(n12010) );
  NAND3_X1 U12072 ( .A1(b_14_), .A2(n12108), .A3(a_11_), .ZN(n12107) );
  NAND2_X1 U12073 ( .A1(n12006), .A2(n12005), .ZN(n12108) );
  OR2_X1 U12074 ( .A1(n12005), .A2(n12006), .ZN(n12106) );
  AND2_X1 U12075 ( .A1(n12109), .A2(n12110), .ZN(n12006) );
  NAND2_X1 U12076 ( .A1(n12003), .A2(n12111), .ZN(n12110) );
  OR2_X1 U12077 ( .A1(n12002), .A2(n12001), .ZN(n12111) );
  NOR2_X1 U12078 ( .A1(n8669), .A2(n8048), .ZN(n12003) );
  NAND2_X1 U12079 ( .A1(n12001), .A2(n12002), .ZN(n12109) );
  NAND2_X1 U12080 ( .A1(n11998), .A2(n12112), .ZN(n12002) );
  NAND2_X1 U12081 ( .A1(n11997), .A2(n11999), .ZN(n12112) );
  NAND2_X1 U12082 ( .A1(n12113), .A2(n12114), .ZN(n11999) );
  NAND2_X1 U12083 ( .A1(a_13_), .A2(b_14_), .ZN(n12114) );
  INV_X1 U12084 ( .A(n12115), .ZN(n12113) );
  XOR2_X1 U12085 ( .A(n12116), .B(n12117), .Z(n11997) );
  XOR2_X1 U12086 ( .A(n12118), .B(n12119), .Z(n12116) );
  NOR2_X1 U12087 ( .A1(n8049), .A2(n7782), .ZN(n12119) );
  NAND2_X1 U12088 ( .A1(a_13_), .A2(n12115), .ZN(n11998) );
  NAND2_X1 U12089 ( .A1(n12120), .A2(n12121), .ZN(n12115) );
  NAND2_X1 U12090 ( .A1(n11993), .A2(n12122), .ZN(n12121) );
  OR2_X1 U12091 ( .A1(n11994), .A2(n11995), .ZN(n12122) );
  XNOR2_X1 U12092 ( .A(n12123), .B(n12124), .ZN(n11993) );
  XOR2_X1 U12093 ( .A(n12125), .B(n12126), .Z(n12124) );
  NAND2_X1 U12094 ( .A1(b_13_), .A2(a_15_), .ZN(n12126) );
  NAND2_X1 U12095 ( .A1(n11995), .A2(n11994), .ZN(n12120) );
  NAND2_X1 U12096 ( .A1(n12127), .A2(n12128), .ZN(n11994) );
  NAND2_X1 U12097 ( .A1(n11882), .A2(n12129), .ZN(n12128) );
  OR2_X1 U12098 ( .A1(n11881), .A2(n11880), .ZN(n12129) );
  NOR2_X1 U12099 ( .A1(n8048), .A2(n7754), .ZN(n11882) );
  NAND2_X1 U12100 ( .A1(n11880), .A2(n11881), .ZN(n12127) );
  NAND2_X1 U12101 ( .A1(n12130), .A2(n12131), .ZN(n11881) );
  NAND2_X1 U12102 ( .A1(n11889), .A2(n12132), .ZN(n12131) );
  OR2_X1 U12103 ( .A1(n11888), .A2(n11886), .ZN(n12132) );
  NOR2_X1 U12104 ( .A1(n8048), .A2(n8438), .ZN(n11889) );
  NAND2_X1 U12105 ( .A1(n11886), .A2(n11888), .ZN(n12130) );
  NAND2_X1 U12106 ( .A1(n12133), .A2(n12134), .ZN(n11888) );
  NAND3_X1 U12107 ( .A1(a_17_), .A2(n12135), .A3(b_14_), .ZN(n12134) );
  OR2_X1 U12108 ( .A1(n11990), .A2(n11989), .ZN(n12135) );
  NAND2_X1 U12109 ( .A1(n11989), .A2(n11990), .ZN(n12133) );
  NAND2_X1 U12110 ( .A1(n12136), .A2(n12137), .ZN(n11990) );
  NAND3_X1 U12111 ( .A1(a_18_), .A2(n12138), .A3(b_14_), .ZN(n12137) );
  NAND2_X1 U12112 ( .A1(n11986), .A2(n11985), .ZN(n12138) );
  OR2_X1 U12113 ( .A1(n11985), .A2(n11986), .ZN(n12136) );
  AND2_X1 U12114 ( .A1(n12139), .A2(n12140), .ZN(n11986) );
  NAND2_X1 U12115 ( .A1(n11983), .A2(n12141), .ZN(n12140) );
  OR2_X1 U12116 ( .A1(n11982), .A2(n11980), .ZN(n12141) );
  NOR2_X1 U12117 ( .A1(n8048), .A2(n8045), .ZN(n11983) );
  NAND2_X1 U12118 ( .A1(n11980), .A2(n11982), .ZN(n12139) );
  NAND2_X1 U12119 ( .A1(n12142), .A2(n12143), .ZN(n11982) );
  NAND3_X1 U12120 ( .A1(a_20_), .A2(n12144), .A3(b_14_), .ZN(n12143) );
  NAND2_X1 U12121 ( .A1(n11978), .A2(n11977), .ZN(n12144) );
  OR2_X1 U12122 ( .A1(n11977), .A2(n11978), .ZN(n12142) );
  AND2_X1 U12123 ( .A1(n12145), .A2(n12146), .ZN(n11978) );
  NAND2_X1 U12124 ( .A1(n11975), .A2(n12147), .ZN(n12146) );
  OR2_X1 U12125 ( .A1(n11974), .A2(n11973), .ZN(n12147) );
  NOR2_X1 U12126 ( .A1(n8048), .A2(n7665), .ZN(n11975) );
  NAND2_X1 U12127 ( .A1(n11973), .A2(n11974), .ZN(n12145) );
  NAND2_X1 U12128 ( .A1(n12148), .A2(n12149), .ZN(n11974) );
  NAND3_X1 U12129 ( .A1(a_22_), .A2(n12150), .A3(b_14_), .ZN(n12149) );
  OR2_X1 U12130 ( .A1(n11970), .A2(n11968), .ZN(n12150) );
  NAND2_X1 U12131 ( .A1(n11968), .A2(n11970), .ZN(n12148) );
  NAND2_X1 U12132 ( .A1(n12151), .A2(n12152), .ZN(n11970) );
  NAND2_X1 U12133 ( .A1(n11967), .A2(n12153), .ZN(n12152) );
  OR2_X1 U12134 ( .A1(n11966), .A2(n11964), .ZN(n12153) );
  NOR2_X1 U12135 ( .A1(n8048), .A2(n8042), .ZN(n11967) );
  NAND2_X1 U12136 ( .A1(n11964), .A2(n11966), .ZN(n12151) );
  NAND2_X1 U12137 ( .A1(n12154), .A2(n12155), .ZN(n11966) );
  NAND3_X1 U12138 ( .A1(a_24_), .A2(n12156), .A3(b_14_), .ZN(n12155) );
  NAND2_X1 U12139 ( .A1(n11962), .A2(n11961), .ZN(n12156) );
  OR2_X1 U12140 ( .A1(n11961), .A2(n11962), .ZN(n12154) );
  AND2_X1 U12141 ( .A1(n12157), .A2(n12158), .ZN(n11962) );
  NAND2_X1 U12142 ( .A1(n11959), .A2(n12159), .ZN(n12158) );
  OR2_X1 U12143 ( .A1(n11958), .A2(n11957), .ZN(n12159) );
  NOR2_X1 U12144 ( .A1(n8048), .A2(n8039), .ZN(n11959) );
  NAND2_X1 U12145 ( .A1(n11957), .A2(n11958), .ZN(n12157) );
  NAND2_X1 U12146 ( .A1(n11954), .A2(n12160), .ZN(n11958) );
  NAND2_X1 U12147 ( .A1(n11953), .A2(n11955), .ZN(n12160) );
  NAND2_X1 U12148 ( .A1(n12161), .A2(n12162), .ZN(n11955) );
  NAND2_X1 U12149 ( .A1(b_14_), .A2(a_26_), .ZN(n12162) );
  INV_X1 U12150 ( .A(n12163), .ZN(n12161) );
  XNOR2_X1 U12151 ( .A(n12164), .B(n12165), .ZN(n11953) );
  NAND2_X1 U12152 ( .A1(n12166), .A2(n12167), .ZN(n12164) );
  NAND2_X1 U12153 ( .A1(a_26_), .A2(n12163), .ZN(n11954) );
  NAND2_X1 U12154 ( .A1(n11926), .A2(n12168), .ZN(n12163) );
  NAND2_X1 U12155 ( .A1(n11925), .A2(n11927), .ZN(n12168) );
  NAND2_X1 U12156 ( .A1(n12169), .A2(n12170), .ZN(n11927) );
  NAND2_X1 U12157 ( .A1(b_14_), .A2(a_27_), .ZN(n12170) );
  INV_X1 U12158 ( .A(n12171), .ZN(n12169) );
  XNOR2_X1 U12159 ( .A(n12172), .B(n12173), .ZN(n11925) );
  XOR2_X1 U12160 ( .A(n12174), .B(n12175), .Z(n12172) );
  NAND2_X1 U12161 ( .A1(b_13_), .A2(a_28_), .ZN(n12174) );
  NAND2_X1 U12162 ( .A1(a_27_), .A2(n12171), .ZN(n11926) );
  NAND2_X1 U12163 ( .A1(n12176), .A2(n12177), .ZN(n12171) );
  NAND3_X1 U12164 ( .A1(a_28_), .A2(n12178), .A3(b_14_), .ZN(n12177) );
  NAND2_X1 U12165 ( .A1(n11935), .A2(n11933), .ZN(n12178) );
  OR2_X1 U12166 ( .A1(n11933), .A2(n11935), .ZN(n12176) );
  AND2_X1 U12167 ( .A1(n12179), .A2(n12180), .ZN(n11935) );
  NAND2_X1 U12168 ( .A1(n11949), .A2(n12181), .ZN(n12180) );
  OR2_X1 U12169 ( .A1(n11950), .A2(n11951), .ZN(n12181) );
  NOR2_X1 U12170 ( .A1(n8048), .A2(n7545), .ZN(n11949) );
  NAND2_X1 U12171 ( .A1(n11951), .A2(n11950), .ZN(n12179) );
  NAND2_X1 U12172 ( .A1(n12182), .A2(n12183), .ZN(n11950) );
  NAND2_X1 U12173 ( .A1(b_12_), .A2(n12184), .ZN(n12183) );
  NAND2_X1 U12174 ( .A1(n7527), .A2(n12185), .ZN(n12184) );
  NAND2_X1 U12175 ( .A1(a_31_), .A2(n7782), .ZN(n12185) );
  NAND2_X1 U12176 ( .A1(b_13_), .A2(n12186), .ZN(n12182) );
  NAND2_X1 U12177 ( .A1(n7531), .A2(n12187), .ZN(n12186) );
  NAND2_X1 U12178 ( .A1(a_30_), .A2(n12188), .ZN(n12187) );
  AND3_X1 U12179 ( .A1(b_14_), .A2(b_13_), .A3(n7494), .ZN(n11951) );
  XNOR2_X1 U12180 ( .A(n12189), .B(n12190), .ZN(n11933) );
  XOR2_X1 U12181 ( .A(n12191), .B(n12192), .Z(n12189) );
  XNOR2_X1 U12182 ( .A(n12193), .B(n12194), .ZN(n11957) );
  NAND2_X1 U12183 ( .A1(n12195), .A2(n12196), .ZN(n12193) );
  XNOR2_X1 U12184 ( .A(n12197), .B(n12198), .ZN(n11961) );
  XOR2_X1 U12185 ( .A(n12199), .B(n12200), .Z(n12197) );
  XNOR2_X1 U12186 ( .A(n12201), .B(n12202), .ZN(n11964) );
  XNOR2_X1 U12187 ( .A(n12203), .B(n12204), .ZN(n12201) );
  NOR2_X1 U12188 ( .A1(n8041), .A2(n7782), .ZN(n12204) );
  XNOR2_X1 U12189 ( .A(n12205), .B(n12206), .ZN(n11968) );
  XNOR2_X1 U12190 ( .A(n12207), .B(n12208), .ZN(n12206) );
  XNOR2_X1 U12191 ( .A(n12209), .B(n12210), .ZN(n11973) );
  XOR2_X1 U12192 ( .A(n12211), .B(n12212), .Z(n12210) );
  NAND2_X1 U12193 ( .A1(b_13_), .A2(a_22_), .ZN(n12212) );
  XNOR2_X1 U12194 ( .A(n12213), .B(n12214), .ZN(n11977) );
  XOR2_X1 U12195 ( .A(n12215), .B(n12216), .Z(n12213) );
  XNOR2_X1 U12196 ( .A(n12217), .B(n12218), .ZN(n11980) );
  XNOR2_X1 U12197 ( .A(n12219), .B(n12220), .ZN(n12217) );
  NOR2_X1 U12198 ( .A1(n8044), .A2(n7782), .ZN(n12220) );
  XOR2_X1 U12199 ( .A(n12221), .B(n12222), .Z(n11985) );
  XNOR2_X1 U12200 ( .A(n12223), .B(n12224), .ZN(n12222) );
  XNOR2_X1 U12201 ( .A(n12225), .B(n12226), .ZN(n11989) );
  XNOR2_X1 U12202 ( .A(n12227), .B(n12228), .ZN(n12225) );
  XNOR2_X1 U12203 ( .A(n12229), .B(n12230), .ZN(n11886) );
  XOR2_X1 U12204 ( .A(n12231), .B(n12232), .Z(n12229) );
  NAND2_X1 U12205 ( .A1(b_13_), .A2(a_17_), .ZN(n12231) );
  XNOR2_X1 U12206 ( .A(n12233), .B(n12234), .ZN(n11880) );
  XNOR2_X1 U12207 ( .A(n12235), .B(n12236), .ZN(n12233) );
  NOR2_X1 U12208 ( .A1(n8438), .A2(n7782), .ZN(n12236) );
  INV_X1 U12209 ( .A(n7773), .ZN(n11995) );
  NAND2_X1 U12210 ( .A1(b_14_), .A2(a_14_), .ZN(n7773) );
  XOR2_X1 U12211 ( .A(n12237), .B(n12238), .Z(n12001) );
  XOR2_X1 U12212 ( .A(n12239), .B(n7780), .Z(n12237) );
  XNOR2_X1 U12213 ( .A(n12240), .B(n12241), .ZN(n12005) );
  XNOR2_X1 U12214 ( .A(n12242), .B(n12243), .ZN(n12240) );
  NAND2_X1 U12215 ( .A1(a_12_), .A2(b_13_), .ZN(n12242) );
  XNOR2_X1 U12216 ( .A(n12244), .B(n12245), .ZN(n12009) );
  XOR2_X1 U12217 ( .A(n12246), .B(n12247), .Z(n12244) );
  NOR2_X1 U12218 ( .A1(n7782), .A2(n7811), .ZN(n12247) );
  XNOR2_X1 U12219 ( .A(n12248), .B(n12249), .ZN(n12012) );
  XNOR2_X1 U12220 ( .A(n12250), .B(n12251), .ZN(n12248) );
  NOR2_X1 U12221 ( .A1(n7782), .A2(n8051), .ZN(n12251) );
  XNOR2_X1 U12222 ( .A(n12252), .B(n12253), .ZN(n12032) );
  XNOR2_X1 U12223 ( .A(n12254), .B(n12255), .ZN(n12252) );
  NOR2_X1 U12224 ( .A1(n7782), .A2(n7908), .ZN(n12255) );
  XNOR2_X1 U12225 ( .A(n12256), .B(n12257), .ZN(n12036) );
  XOR2_X1 U12226 ( .A(n12258), .B(n12259), .Z(n12257) );
  NAND2_X1 U12227 ( .A1(a_4_), .A2(b_13_), .ZN(n12259) );
  XOR2_X1 U12228 ( .A(n12260), .B(n12261), .Z(n12041) );
  XOR2_X1 U12229 ( .A(n12262), .B(n12263), .Z(n12261) );
  NAND2_X1 U12230 ( .A1(a_3_), .A2(b_13_), .ZN(n12263) );
  XNOR2_X1 U12231 ( .A(n12264), .B(n12265), .ZN(n12044) );
  XNOR2_X1 U12232 ( .A(n12266), .B(n12267), .ZN(n12264) );
  NOR2_X1 U12233 ( .A1(n7782), .A2(n8056), .ZN(n12267) );
  XNOR2_X1 U12234 ( .A(n12268), .B(n12269), .ZN(n12048) );
  XOR2_X1 U12235 ( .A(n12270), .B(n12271), .Z(n12269) );
  NAND2_X1 U12236 ( .A1(b_13_), .A2(a_1_), .ZN(n12271) );
  NAND2_X1 U12237 ( .A1(n12272), .A2(n12273), .ZN(n8207) );
  XNOR2_X1 U12238 ( .A(n12274), .B(n12275), .ZN(n8208) );
  XNOR2_X1 U12239 ( .A(n12276), .B(n12277), .ZN(n12275) );
  NAND2_X1 U12240 ( .A1(n12052), .A2(n12278), .ZN(n8161) );
  XOR2_X1 U12241 ( .A(n8200), .B(n8199), .Z(n12278) );
  NOR2_X1 U12242 ( .A1(n12273), .A2(n12272), .ZN(n12052) );
  AND2_X1 U12243 ( .A1(n12279), .A2(n12280), .ZN(n12272) );
  NAND2_X1 U12244 ( .A1(n12277), .A2(n12281), .ZN(n12280) );
  OR2_X1 U12245 ( .A1(n12276), .A2(n12274), .ZN(n12281) );
  NOR2_X1 U12246 ( .A1(n8942), .A2(n7782), .ZN(n12277) );
  NAND2_X1 U12247 ( .A1(n12274), .A2(n12276), .ZN(n12279) );
  NAND2_X1 U12248 ( .A1(n12282), .A2(n12283), .ZN(n12276) );
  NAND3_X1 U12249 ( .A1(a_1_), .A2(n12284), .A3(b_13_), .ZN(n12283) );
  OR2_X1 U12250 ( .A1(n12270), .A2(n12268), .ZN(n12284) );
  NAND2_X1 U12251 ( .A1(n12268), .A2(n12270), .ZN(n12282) );
  NAND2_X1 U12252 ( .A1(n12285), .A2(n12286), .ZN(n12270) );
  NAND3_X1 U12253 ( .A1(b_13_), .A2(n12287), .A3(a_2_), .ZN(n12286) );
  NAND2_X1 U12254 ( .A1(n12266), .A2(n12265), .ZN(n12287) );
  OR2_X1 U12255 ( .A1(n12265), .A2(n12266), .ZN(n12285) );
  AND2_X1 U12256 ( .A1(n12288), .A2(n12289), .ZN(n12266) );
  NAND3_X1 U12257 ( .A1(b_13_), .A2(n12290), .A3(a_3_), .ZN(n12289) );
  OR2_X1 U12258 ( .A1(n12262), .A2(n12260), .ZN(n12290) );
  NAND2_X1 U12259 ( .A1(n12260), .A2(n12262), .ZN(n12288) );
  NAND2_X1 U12260 ( .A1(n12291), .A2(n12292), .ZN(n12262) );
  NAND3_X1 U12261 ( .A1(b_13_), .A2(n12293), .A3(a_4_), .ZN(n12292) );
  OR2_X1 U12262 ( .A1(n12258), .A2(n12256), .ZN(n12293) );
  NAND2_X1 U12263 ( .A1(n12256), .A2(n12258), .ZN(n12291) );
  NAND2_X1 U12264 ( .A1(n12294), .A2(n12295), .ZN(n12258) );
  NAND3_X1 U12265 ( .A1(b_13_), .A2(n12296), .A3(a_5_), .ZN(n12295) );
  NAND2_X1 U12266 ( .A1(n12254), .A2(n12253), .ZN(n12296) );
  OR2_X1 U12267 ( .A1(n12253), .A2(n12254), .ZN(n12294) );
  AND2_X1 U12268 ( .A1(n12297), .A2(n12298), .ZN(n12254) );
  NAND3_X1 U12269 ( .A1(b_13_), .A2(n12299), .A3(a_6_), .ZN(n12298) );
  OR2_X1 U12270 ( .A1(n12074), .A2(n12072), .ZN(n12299) );
  NAND2_X1 U12271 ( .A1(n12072), .A2(n12074), .ZN(n12297) );
  NAND2_X1 U12272 ( .A1(n12300), .A2(n12301), .ZN(n12074) );
  NAND3_X1 U12273 ( .A1(b_13_), .A2(n12302), .A3(a_7_), .ZN(n12301) );
  OR2_X1 U12274 ( .A1(n12082), .A2(n12080), .ZN(n12302) );
  NAND2_X1 U12275 ( .A1(n12080), .A2(n12082), .ZN(n12300) );
  NAND2_X1 U12276 ( .A1(n12303), .A2(n12304), .ZN(n12082) );
  NAND3_X1 U12277 ( .A1(b_13_), .A2(n12305), .A3(a_8_), .ZN(n12304) );
  NAND2_X1 U12278 ( .A1(n12090), .A2(n12089), .ZN(n12305) );
  OR2_X1 U12279 ( .A1(n12089), .A2(n12090), .ZN(n12303) );
  AND2_X1 U12280 ( .A1(n12306), .A2(n12307), .ZN(n12090) );
  NAND3_X1 U12281 ( .A1(b_13_), .A2(n12308), .A3(a_9_), .ZN(n12307) );
  OR2_X1 U12282 ( .A1(n12098), .A2(n12096), .ZN(n12308) );
  NAND2_X1 U12283 ( .A1(n12096), .A2(n12098), .ZN(n12306) );
  NAND2_X1 U12284 ( .A1(n12309), .A2(n12310), .ZN(n12098) );
  NAND3_X1 U12285 ( .A1(b_13_), .A2(n12311), .A3(a_10_), .ZN(n12310) );
  NAND2_X1 U12286 ( .A1(n12250), .A2(n12249), .ZN(n12311) );
  OR2_X1 U12287 ( .A1(n12249), .A2(n12250), .ZN(n12309) );
  AND2_X1 U12288 ( .A1(n12312), .A2(n12313), .ZN(n12250) );
  NAND3_X1 U12289 ( .A1(b_13_), .A2(n12314), .A3(a_11_), .ZN(n12313) );
  OR2_X1 U12290 ( .A1(n12246), .A2(n12245), .ZN(n12314) );
  NAND2_X1 U12291 ( .A1(n12245), .A2(n12246), .ZN(n12312) );
  NAND2_X1 U12292 ( .A1(n12315), .A2(n12316), .ZN(n12246) );
  NAND3_X1 U12293 ( .A1(b_13_), .A2(n12317), .A3(a_12_), .ZN(n12316) );
  OR2_X1 U12294 ( .A1(n12243), .A2(n12241), .ZN(n12317) );
  NAND2_X1 U12295 ( .A1(n12241), .A2(n12243), .ZN(n12315) );
  NAND2_X1 U12296 ( .A1(n12318), .A2(n12319), .ZN(n12243) );
  NAND2_X1 U12297 ( .A1(n12238), .A2(n12320), .ZN(n12319) );
  OR2_X1 U12298 ( .A1(n12239), .A2(n7780), .ZN(n12320) );
  XNOR2_X1 U12299 ( .A(n12321), .B(n12322), .ZN(n12238) );
  NAND2_X1 U12300 ( .A1(n12323), .A2(n12324), .ZN(n12321) );
  NAND2_X1 U12301 ( .A1(n7780), .A2(n12239), .ZN(n12318) );
  NAND2_X1 U12302 ( .A1(n12325), .A2(n12326), .ZN(n12239) );
  NAND3_X1 U12303 ( .A1(a_14_), .A2(n12327), .A3(b_13_), .ZN(n12326) );
  OR2_X1 U12304 ( .A1(n12118), .A2(n12117), .ZN(n12327) );
  NAND2_X1 U12305 ( .A1(n12117), .A2(n12118), .ZN(n12325) );
  NAND2_X1 U12306 ( .A1(n12328), .A2(n12329), .ZN(n12118) );
  NAND3_X1 U12307 ( .A1(a_15_), .A2(n12330), .A3(b_13_), .ZN(n12329) );
  OR2_X1 U12308 ( .A1(n12125), .A2(n12123), .ZN(n12330) );
  NAND2_X1 U12309 ( .A1(n12123), .A2(n12125), .ZN(n12328) );
  NAND2_X1 U12310 ( .A1(n12331), .A2(n12332), .ZN(n12125) );
  NAND3_X1 U12311 ( .A1(a_16_), .A2(n12333), .A3(b_13_), .ZN(n12332) );
  NAND2_X1 U12312 ( .A1(n12235), .A2(n12234), .ZN(n12333) );
  OR2_X1 U12313 ( .A1(n12234), .A2(n12235), .ZN(n12331) );
  AND2_X1 U12314 ( .A1(n12334), .A2(n12335), .ZN(n12235) );
  NAND3_X1 U12315 ( .A1(a_17_), .A2(n12336), .A3(b_13_), .ZN(n12335) );
  NAND2_X1 U12316 ( .A1(n12232), .A2(n12230), .ZN(n12336) );
  OR2_X1 U12317 ( .A1(n12230), .A2(n12232), .ZN(n12334) );
  AND2_X1 U12318 ( .A1(n12337), .A2(n12338), .ZN(n12232) );
  NAND2_X1 U12319 ( .A1(n12228), .A2(n12339), .ZN(n12338) );
  NAND2_X1 U12320 ( .A1(n12227), .A2(n12226), .ZN(n12339) );
  NOR2_X1 U12321 ( .A1(n7782), .A2(n8047), .ZN(n12228) );
  OR2_X1 U12322 ( .A1(n12226), .A2(n12227), .ZN(n12337) );
  AND2_X1 U12323 ( .A1(n12340), .A2(n12341), .ZN(n12227) );
  NAND2_X1 U12324 ( .A1(n12224), .A2(n12342), .ZN(n12341) );
  OR2_X1 U12325 ( .A1(n12223), .A2(n12221), .ZN(n12342) );
  NOR2_X1 U12326 ( .A1(n7782), .A2(n8045), .ZN(n12224) );
  NAND2_X1 U12327 ( .A1(n12221), .A2(n12223), .ZN(n12340) );
  NAND2_X1 U12328 ( .A1(n12343), .A2(n12344), .ZN(n12223) );
  NAND3_X1 U12329 ( .A1(a_20_), .A2(n12345), .A3(b_13_), .ZN(n12344) );
  NAND2_X1 U12330 ( .A1(n12219), .A2(n12218), .ZN(n12345) );
  OR2_X1 U12331 ( .A1(n12218), .A2(n12219), .ZN(n12343) );
  AND2_X1 U12332 ( .A1(n12346), .A2(n12347), .ZN(n12219) );
  NAND2_X1 U12333 ( .A1(n12216), .A2(n12348), .ZN(n12347) );
  OR2_X1 U12334 ( .A1(n12215), .A2(n12214), .ZN(n12348) );
  NOR2_X1 U12335 ( .A1(n7782), .A2(n7665), .ZN(n12216) );
  NAND2_X1 U12336 ( .A1(n12214), .A2(n12215), .ZN(n12346) );
  NAND2_X1 U12337 ( .A1(n12349), .A2(n12350), .ZN(n12215) );
  NAND3_X1 U12338 ( .A1(a_22_), .A2(n12351), .A3(b_13_), .ZN(n12350) );
  OR2_X1 U12339 ( .A1(n12211), .A2(n12209), .ZN(n12351) );
  NAND2_X1 U12340 ( .A1(n12209), .A2(n12211), .ZN(n12349) );
  NAND2_X1 U12341 ( .A1(n12352), .A2(n12353), .ZN(n12211) );
  NAND2_X1 U12342 ( .A1(n12208), .A2(n12354), .ZN(n12353) );
  OR2_X1 U12343 ( .A1(n12207), .A2(n12205), .ZN(n12354) );
  NOR2_X1 U12344 ( .A1(n7782), .A2(n8042), .ZN(n12208) );
  NAND2_X1 U12345 ( .A1(n12205), .A2(n12207), .ZN(n12352) );
  NAND2_X1 U12346 ( .A1(n12355), .A2(n12356), .ZN(n12207) );
  NAND3_X1 U12347 ( .A1(a_24_), .A2(n12357), .A3(b_13_), .ZN(n12356) );
  NAND2_X1 U12348 ( .A1(n12203), .A2(n12202), .ZN(n12357) );
  OR2_X1 U12349 ( .A1(n12202), .A2(n12203), .ZN(n12355) );
  AND2_X1 U12350 ( .A1(n12358), .A2(n12359), .ZN(n12203) );
  NAND2_X1 U12351 ( .A1(n12200), .A2(n12360), .ZN(n12359) );
  OR2_X1 U12352 ( .A1(n12199), .A2(n12198), .ZN(n12360) );
  NOR2_X1 U12353 ( .A1(n7782), .A2(n8039), .ZN(n12200) );
  NAND2_X1 U12354 ( .A1(n12198), .A2(n12199), .ZN(n12358) );
  NAND2_X1 U12355 ( .A1(n12195), .A2(n12361), .ZN(n12199) );
  NAND2_X1 U12356 ( .A1(n12194), .A2(n12196), .ZN(n12361) );
  NAND2_X1 U12357 ( .A1(n12362), .A2(n12363), .ZN(n12196) );
  NAND2_X1 U12358 ( .A1(b_13_), .A2(a_26_), .ZN(n12363) );
  INV_X1 U12359 ( .A(n12364), .ZN(n12362) );
  XNOR2_X1 U12360 ( .A(n12365), .B(n12366), .ZN(n12194) );
  NAND2_X1 U12361 ( .A1(n12367), .A2(n12368), .ZN(n12365) );
  NAND2_X1 U12362 ( .A1(a_26_), .A2(n12364), .ZN(n12195) );
  NAND2_X1 U12363 ( .A1(n12166), .A2(n12369), .ZN(n12364) );
  NAND2_X1 U12364 ( .A1(n12165), .A2(n12167), .ZN(n12369) );
  NAND2_X1 U12365 ( .A1(n12370), .A2(n12371), .ZN(n12167) );
  NAND2_X1 U12366 ( .A1(b_13_), .A2(a_27_), .ZN(n12371) );
  INV_X1 U12367 ( .A(n12372), .ZN(n12370) );
  XNOR2_X1 U12368 ( .A(n12373), .B(n12374), .ZN(n12165) );
  XOR2_X1 U12369 ( .A(n12375), .B(n12376), .Z(n12373) );
  NAND2_X1 U12370 ( .A1(b_12_), .A2(a_28_), .ZN(n12375) );
  NAND2_X1 U12371 ( .A1(a_27_), .A2(n12372), .ZN(n12166) );
  NAND2_X1 U12372 ( .A1(n12377), .A2(n12378), .ZN(n12372) );
  NAND3_X1 U12373 ( .A1(a_28_), .A2(n12379), .A3(b_13_), .ZN(n12378) );
  NAND2_X1 U12374 ( .A1(n12175), .A2(n12173), .ZN(n12379) );
  OR2_X1 U12375 ( .A1(n12173), .A2(n12175), .ZN(n12377) );
  AND2_X1 U12376 ( .A1(n12380), .A2(n12381), .ZN(n12175) );
  NAND2_X1 U12377 ( .A1(n12190), .A2(n12382), .ZN(n12381) );
  OR2_X1 U12378 ( .A1(n12191), .A2(n12192), .ZN(n12382) );
  NOR2_X1 U12379 ( .A1(n7782), .A2(n7545), .ZN(n12190) );
  NAND2_X1 U12380 ( .A1(n12192), .A2(n12191), .ZN(n12380) );
  NAND2_X1 U12381 ( .A1(n12383), .A2(n12384), .ZN(n12191) );
  NAND2_X1 U12382 ( .A1(b_11_), .A2(n12385), .ZN(n12384) );
  NAND2_X1 U12383 ( .A1(n7527), .A2(n12386), .ZN(n12385) );
  NAND2_X1 U12384 ( .A1(a_31_), .A2(n12188), .ZN(n12386) );
  NAND2_X1 U12385 ( .A1(b_12_), .A2(n12387), .ZN(n12383) );
  NAND2_X1 U12386 ( .A1(n7531), .A2(n12388), .ZN(n12387) );
  NAND2_X1 U12387 ( .A1(a_30_), .A2(n7813), .ZN(n12388) );
  AND3_X1 U12388 ( .A1(b_12_), .A2(b_13_), .A3(n7494), .ZN(n12192) );
  XNOR2_X1 U12389 ( .A(n12389), .B(n12390), .ZN(n12173) );
  XOR2_X1 U12390 ( .A(n12391), .B(n12392), .Z(n12389) );
  XNOR2_X1 U12391 ( .A(n12393), .B(n12394), .ZN(n12198) );
  NAND2_X1 U12392 ( .A1(n12395), .A2(n12396), .ZN(n12393) );
  XNOR2_X1 U12393 ( .A(n12397), .B(n12398), .ZN(n12202) );
  XOR2_X1 U12394 ( .A(n12399), .B(n12400), .Z(n12397) );
  XNOR2_X1 U12395 ( .A(n12401), .B(n12402), .ZN(n12205) );
  XNOR2_X1 U12396 ( .A(n12403), .B(n12404), .ZN(n12401) );
  NOR2_X1 U12397 ( .A1(n8041), .A2(n12188), .ZN(n12404) );
  XNOR2_X1 U12398 ( .A(n12405), .B(n12406), .ZN(n12209) );
  XNOR2_X1 U12399 ( .A(n12407), .B(n12408), .ZN(n12406) );
  XNOR2_X1 U12400 ( .A(n12409), .B(n12410), .ZN(n12214) );
  XOR2_X1 U12401 ( .A(n12411), .B(n12412), .Z(n12410) );
  NAND2_X1 U12402 ( .A1(b_12_), .A2(a_22_), .ZN(n12412) );
  XNOR2_X1 U12403 ( .A(n12413), .B(n12414), .ZN(n12218) );
  XOR2_X1 U12404 ( .A(n12415), .B(n12416), .Z(n12413) );
  XNOR2_X1 U12405 ( .A(n12417), .B(n12418), .ZN(n12221) );
  XNOR2_X1 U12406 ( .A(n12419), .B(n12420), .ZN(n12417) );
  NOR2_X1 U12407 ( .A1(n8044), .A2(n12188), .ZN(n12420) );
  XOR2_X1 U12408 ( .A(n12421), .B(n12422), .Z(n12226) );
  NAND2_X1 U12409 ( .A1(n12423), .A2(n12424), .ZN(n12421) );
  XNOR2_X1 U12410 ( .A(n12425), .B(n12426), .ZN(n12230) );
  XOR2_X1 U12411 ( .A(n12427), .B(n12428), .Z(n12425) );
  XNOR2_X1 U12412 ( .A(n12429), .B(n12430), .ZN(n12234) );
  XOR2_X1 U12413 ( .A(n12431), .B(n12432), .Z(n12429) );
  XNOR2_X1 U12414 ( .A(n12433), .B(n12434), .ZN(n12123) );
  XNOR2_X1 U12415 ( .A(n12435), .B(n12436), .ZN(n12433) );
  NOR2_X1 U12416 ( .A1(n8438), .A2(n12188), .ZN(n12436) );
  XNOR2_X1 U12417 ( .A(n12437), .B(n12438), .ZN(n12117) );
  NAND2_X1 U12418 ( .A1(n12439), .A2(n12440), .ZN(n12437) );
  INV_X1 U12419 ( .A(n7999), .ZN(n7780) );
  NAND2_X1 U12420 ( .A1(a_13_), .A2(b_13_), .ZN(n7999) );
  XNOR2_X1 U12421 ( .A(n12441), .B(n12442), .ZN(n12241) );
  XNOR2_X1 U12422 ( .A(n12443), .B(n12444), .ZN(n12442) );
  XNOR2_X1 U12423 ( .A(n12445), .B(n12446), .ZN(n12245) );
  XNOR2_X1 U12424 ( .A(n12447), .B(n7801), .ZN(n12446) );
  XOR2_X1 U12425 ( .A(n12448), .B(n12449), .Z(n12249) );
  NAND2_X1 U12426 ( .A1(n12450), .A2(n12451), .ZN(n12448) );
  XNOR2_X1 U12427 ( .A(n12452), .B(n12453), .ZN(n12096) );
  NAND2_X1 U12428 ( .A1(n12454), .A2(n12455), .ZN(n12452) );
  XNOR2_X1 U12429 ( .A(n12456), .B(n12457), .ZN(n12089) );
  XOR2_X1 U12430 ( .A(n12458), .B(n12459), .Z(n12456) );
  XOR2_X1 U12431 ( .A(n12460), .B(n12461), .Z(n12080) );
  XOR2_X1 U12432 ( .A(n12462), .B(n12463), .Z(n12460) );
  NOR2_X1 U12433 ( .A1(n12188), .A2(n8686), .ZN(n12463) );
  XNOR2_X1 U12434 ( .A(n12464), .B(n12465), .ZN(n12072) );
  NAND2_X1 U12435 ( .A1(n12466), .A2(n12467), .ZN(n12464) );
  XNOR2_X1 U12436 ( .A(n12468), .B(n12469), .ZN(n12253) );
  XOR2_X1 U12437 ( .A(n12470), .B(n12471), .Z(n12468) );
  XNOR2_X1 U12438 ( .A(n12472), .B(n12473), .ZN(n12256) );
  XNOR2_X1 U12439 ( .A(n12474), .B(n12475), .ZN(n12472) );
  NOR2_X1 U12440 ( .A1(n12188), .A2(n7908), .ZN(n12475) );
  XNOR2_X1 U12441 ( .A(n12476), .B(n12477), .ZN(n12260) );
  XNOR2_X1 U12442 ( .A(n12478), .B(n12479), .ZN(n12477) );
  XNOR2_X1 U12443 ( .A(n12480), .B(n12481), .ZN(n12265) );
  XOR2_X1 U12444 ( .A(n12482), .B(n12483), .Z(n12480) );
  NOR2_X1 U12445 ( .A1(n12188), .A2(n7937), .ZN(n12483) );
  XNOR2_X1 U12446 ( .A(n12484), .B(n12485), .ZN(n12268) );
  XNOR2_X1 U12447 ( .A(n12486), .B(n12487), .ZN(n12484) );
  XNOR2_X1 U12448 ( .A(n12488), .B(n12489), .ZN(n12274) );
  XNOR2_X1 U12449 ( .A(n12490), .B(n12491), .ZN(n12489) );
  XOR2_X1 U12450 ( .A(n12492), .B(n12493), .Z(n12273) );
  XNOR2_X1 U12451 ( .A(n12494), .B(n12495), .ZN(n12492) );
  NOR2_X1 U12452 ( .A1(n12188), .A2(n8942), .ZN(n12495) );
  NAND4_X1 U12453 ( .A1(n8199), .A2(n8198), .A3(n8200), .A4(n8192), .ZN(n8166)
         );
  INV_X1 U12454 ( .A(n12496), .ZN(n8192) );
  NAND2_X1 U12455 ( .A1(n12497), .A2(n12498), .ZN(n8200) );
  NAND3_X1 U12456 ( .A1(b_12_), .A2(n12499), .A3(a_0_), .ZN(n12498) );
  NAND2_X1 U12457 ( .A1(n12494), .A2(n12493), .ZN(n12499) );
  OR2_X1 U12458 ( .A1(n12493), .A2(n12494), .ZN(n12497) );
  AND2_X1 U12459 ( .A1(n12500), .A2(n12501), .ZN(n12494) );
  NAND2_X1 U12460 ( .A1(n12491), .A2(n12502), .ZN(n12501) );
  OR2_X1 U12461 ( .A1(n12490), .A2(n12488), .ZN(n12502) );
  NOR2_X1 U12462 ( .A1(n12188), .A2(n7957), .ZN(n12491) );
  NAND2_X1 U12463 ( .A1(n12488), .A2(n12490), .ZN(n12500) );
  NAND2_X1 U12464 ( .A1(n12503), .A2(n12504), .ZN(n12490) );
  NAND2_X1 U12465 ( .A1(n12487), .A2(n12505), .ZN(n12504) );
  NAND2_X1 U12466 ( .A1(n12486), .A2(n12485), .ZN(n12505) );
  NOR2_X1 U12467 ( .A1(n8056), .A2(n12188), .ZN(n12487) );
  OR2_X1 U12468 ( .A1(n12485), .A2(n12486), .ZN(n12503) );
  AND2_X1 U12469 ( .A1(n12506), .A2(n12507), .ZN(n12486) );
  NAND3_X1 U12470 ( .A1(b_12_), .A2(n12508), .A3(a_3_), .ZN(n12507) );
  OR2_X1 U12471 ( .A1(n12482), .A2(n12481), .ZN(n12508) );
  NAND2_X1 U12472 ( .A1(n12481), .A2(n12482), .ZN(n12506) );
  NAND2_X1 U12473 ( .A1(n12509), .A2(n12510), .ZN(n12482) );
  NAND2_X1 U12474 ( .A1(n12479), .A2(n12511), .ZN(n12510) );
  OR2_X1 U12475 ( .A1(n12478), .A2(n12476), .ZN(n12511) );
  NOR2_X1 U12476 ( .A1(n7916), .A2(n12188), .ZN(n12479) );
  NAND2_X1 U12477 ( .A1(n12476), .A2(n12478), .ZN(n12509) );
  NAND2_X1 U12478 ( .A1(n12512), .A2(n12513), .ZN(n12478) );
  NAND3_X1 U12479 ( .A1(b_12_), .A2(n12514), .A3(a_5_), .ZN(n12513) );
  NAND2_X1 U12480 ( .A1(n12474), .A2(n12473), .ZN(n12514) );
  OR2_X1 U12481 ( .A1(n12473), .A2(n12474), .ZN(n12512) );
  AND2_X1 U12482 ( .A1(n12515), .A2(n12516), .ZN(n12474) );
  NAND2_X1 U12483 ( .A1(n12471), .A2(n12517), .ZN(n12516) );
  OR2_X1 U12484 ( .A1(n12470), .A2(n12469), .ZN(n12517) );
  NOR2_X1 U12485 ( .A1(n7887), .A2(n12188), .ZN(n12471) );
  NAND2_X1 U12486 ( .A1(n12469), .A2(n12470), .ZN(n12515) );
  NAND2_X1 U12487 ( .A1(n12466), .A2(n12518), .ZN(n12470) );
  NAND2_X1 U12488 ( .A1(n12465), .A2(n12467), .ZN(n12518) );
  NAND2_X1 U12489 ( .A1(n12519), .A2(n12520), .ZN(n12467) );
  NAND2_X1 U12490 ( .A1(a_7_), .A2(b_12_), .ZN(n12520) );
  INV_X1 U12491 ( .A(n12521), .ZN(n12519) );
  XNOR2_X1 U12492 ( .A(n12522), .B(n12523), .ZN(n12465) );
  XOR2_X1 U12493 ( .A(n12524), .B(n12525), .Z(n12523) );
  NAND2_X1 U12494 ( .A1(a_8_), .A2(b_11_), .ZN(n12525) );
  NAND2_X1 U12495 ( .A1(a_7_), .A2(n12521), .ZN(n12466) );
  NAND2_X1 U12496 ( .A1(n12526), .A2(n12527), .ZN(n12521) );
  NAND3_X1 U12497 ( .A1(b_12_), .A2(n12528), .A3(a_8_), .ZN(n12527) );
  OR2_X1 U12498 ( .A1(n12462), .A2(n12461), .ZN(n12528) );
  NAND2_X1 U12499 ( .A1(n12461), .A2(n12462), .ZN(n12526) );
  NAND2_X1 U12500 ( .A1(n12529), .A2(n12530), .ZN(n12462) );
  NAND2_X1 U12501 ( .A1(n12459), .A2(n12531), .ZN(n12530) );
  OR2_X1 U12502 ( .A1(n12458), .A2(n12457), .ZN(n12531) );
  NOR2_X1 U12503 ( .A1(n8052), .A2(n12188), .ZN(n12459) );
  NAND2_X1 U12504 ( .A1(n12457), .A2(n12458), .ZN(n12529) );
  NAND2_X1 U12505 ( .A1(n12454), .A2(n12532), .ZN(n12458) );
  NAND2_X1 U12506 ( .A1(n12453), .A2(n12455), .ZN(n12532) );
  NAND2_X1 U12507 ( .A1(n12533), .A2(n12534), .ZN(n12455) );
  NAND2_X1 U12508 ( .A1(a_10_), .A2(b_12_), .ZN(n12534) );
  INV_X1 U12509 ( .A(n12535), .ZN(n12533) );
  XOR2_X1 U12510 ( .A(n12536), .B(n12537), .Z(n12453) );
  XOR2_X1 U12511 ( .A(n12538), .B(n7808), .Z(n12536) );
  NAND2_X1 U12512 ( .A1(a_10_), .A2(n12535), .ZN(n12454) );
  NAND2_X1 U12513 ( .A1(n12450), .A2(n12539), .ZN(n12535) );
  NAND2_X1 U12514 ( .A1(n12449), .A2(n12451), .ZN(n12539) );
  NAND2_X1 U12515 ( .A1(n12540), .A2(n12541), .ZN(n12451) );
  NAND2_X1 U12516 ( .A1(a_11_), .A2(b_12_), .ZN(n12541) );
  INV_X1 U12517 ( .A(n12542), .ZN(n12540) );
  XOR2_X1 U12518 ( .A(n12543), .B(n12544), .Z(n12449) );
  XOR2_X1 U12519 ( .A(n12545), .B(n12546), .Z(n12543) );
  NOR2_X1 U12520 ( .A1(n8669), .A2(n7813), .ZN(n12546) );
  NAND2_X1 U12521 ( .A1(a_11_), .A2(n12542), .ZN(n12450) );
  NAND2_X1 U12522 ( .A1(n12547), .A2(n12548), .ZN(n12542) );
  NAND2_X1 U12523 ( .A1(n12445), .A2(n12549), .ZN(n12548) );
  OR2_X1 U12524 ( .A1(n12447), .A2(n7801), .ZN(n12549) );
  XNOR2_X1 U12525 ( .A(n12550), .B(n12551), .ZN(n12445) );
  XOR2_X1 U12526 ( .A(n12552), .B(n12553), .Z(n12551) );
  NAND2_X1 U12527 ( .A1(b_11_), .A2(a_13_), .ZN(n12553) );
  NAND2_X1 U12528 ( .A1(n7801), .A2(n12447), .ZN(n12547) );
  NAND2_X1 U12529 ( .A1(n12554), .A2(n12555), .ZN(n12447) );
  NAND2_X1 U12530 ( .A1(n12444), .A2(n12556), .ZN(n12555) );
  OR2_X1 U12531 ( .A1(n12443), .A2(n12441), .ZN(n12556) );
  NOR2_X1 U12532 ( .A1(n12188), .A2(n7789), .ZN(n12444) );
  NAND2_X1 U12533 ( .A1(n12441), .A2(n12443), .ZN(n12554) );
  NAND2_X1 U12534 ( .A1(n12323), .A2(n12557), .ZN(n12443) );
  NAND2_X1 U12535 ( .A1(n12322), .A2(n12324), .ZN(n12557) );
  NAND2_X1 U12536 ( .A1(n12558), .A2(n12559), .ZN(n12324) );
  NAND2_X1 U12537 ( .A1(b_12_), .A2(a_14_), .ZN(n12559) );
  INV_X1 U12538 ( .A(n12560), .ZN(n12558) );
  XNOR2_X1 U12539 ( .A(n12561), .B(n12562), .ZN(n12322) );
  XOR2_X1 U12540 ( .A(n12563), .B(n12564), .Z(n12562) );
  NAND2_X1 U12541 ( .A1(b_11_), .A2(a_15_), .ZN(n12564) );
  NAND2_X1 U12542 ( .A1(a_14_), .A2(n12560), .ZN(n12323) );
  NAND2_X1 U12543 ( .A1(n12439), .A2(n12565), .ZN(n12560) );
  NAND2_X1 U12544 ( .A1(n12438), .A2(n12440), .ZN(n12565) );
  NAND2_X1 U12545 ( .A1(n12566), .A2(n12567), .ZN(n12440) );
  NAND2_X1 U12546 ( .A1(b_12_), .A2(a_15_), .ZN(n12567) );
  INV_X1 U12547 ( .A(n12568), .ZN(n12566) );
  XNOR2_X1 U12548 ( .A(n12569), .B(n12570), .ZN(n12438) );
  XNOR2_X1 U12549 ( .A(n12571), .B(n12572), .ZN(n12569) );
  NOR2_X1 U12550 ( .A1(n8438), .A2(n7813), .ZN(n12572) );
  NAND2_X1 U12551 ( .A1(a_15_), .A2(n12568), .ZN(n12439) );
  NAND2_X1 U12552 ( .A1(n12573), .A2(n12574), .ZN(n12568) );
  NAND3_X1 U12553 ( .A1(a_16_), .A2(n12575), .A3(b_12_), .ZN(n12574) );
  NAND2_X1 U12554 ( .A1(n12435), .A2(n12434), .ZN(n12575) );
  OR2_X1 U12555 ( .A1(n12434), .A2(n12435), .ZN(n12573) );
  AND2_X1 U12556 ( .A1(n12576), .A2(n12577), .ZN(n12435) );
  NAND2_X1 U12557 ( .A1(n12431), .A2(n12578), .ZN(n12577) );
  OR2_X1 U12558 ( .A1(n12432), .A2(n12430), .ZN(n12578) );
  NOR2_X1 U12559 ( .A1(n12188), .A2(n7732), .ZN(n12431) );
  NAND2_X1 U12560 ( .A1(n12430), .A2(n12432), .ZN(n12576) );
  NAND2_X1 U12561 ( .A1(n12579), .A2(n12580), .ZN(n12432) );
  NAND2_X1 U12562 ( .A1(n12427), .A2(n12581), .ZN(n12580) );
  OR2_X1 U12563 ( .A1(n12428), .A2(n12426), .ZN(n12581) );
  NOR2_X1 U12564 ( .A1(n12188), .A2(n8047), .ZN(n12427) );
  NAND2_X1 U12565 ( .A1(n12426), .A2(n12428), .ZN(n12579) );
  NAND2_X1 U12566 ( .A1(n12423), .A2(n12582), .ZN(n12428) );
  NAND2_X1 U12567 ( .A1(n12422), .A2(n12424), .ZN(n12582) );
  NAND2_X1 U12568 ( .A1(n12583), .A2(n12584), .ZN(n12424) );
  NAND2_X1 U12569 ( .A1(b_12_), .A2(a_19_), .ZN(n12584) );
  INV_X1 U12570 ( .A(n12585), .ZN(n12583) );
  XOR2_X1 U12571 ( .A(n12586), .B(n12587), .Z(n12422) );
  XOR2_X1 U12572 ( .A(n12588), .B(n12589), .Z(n12586) );
  NOR2_X1 U12573 ( .A1(n8044), .A2(n7813), .ZN(n12589) );
  NAND2_X1 U12574 ( .A1(a_19_), .A2(n12585), .ZN(n12423) );
  NAND2_X1 U12575 ( .A1(n12590), .A2(n12591), .ZN(n12585) );
  NAND3_X1 U12576 ( .A1(a_20_), .A2(n12592), .A3(b_12_), .ZN(n12591) );
  NAND2_X1 U12577 ( .A1(n12419), .A2(n12418), .ZN(n12592) );
  OR2_X1 U12578 ( .A1(n12418), .A2(n12419), .ZN(n12590) );
  AND2_X1 U12579 ( .A1(n12593), .A2(n12594), .ZN(n12419) );
  NAND2_X1 U12580 ( .A1(n12416), .A2(n12595), .ZN(n12594) );
  OR2_X1 U12581 ( .A1(n12415), .A2(n12414), .ZN(n12595) );
  NOR2_X1 U12582 ( .A1(n12188), .A2(n7665), .ZN(n12416) );
  NAND2_X1 U12583 ( .A1(n12414), .A2(n12415), .ZN(n12593) );
  NAND2_X1 U12584 ( .A1(n12596), .A2(n12597), .ZN(n12415) );
  NAND3_X1 U12585 ( .A1(a_22_), .A2(n12598), .A3(b_12_), .ZN(n12597) );
  OR2_X1 U12586 ( .A1(n12411), .A2(n12409), .ZN(n12598) );
  NAND2_X1 U12587 ( .A1(n12409), .A2(n12411), .ZN(n12596) );
  NAND2_X1 U12588 ( .A1(n12599), .A2(n12600), .ZN(n12411) );
  NAND2_X1 U12589 ( .A1(n12408), .A2(n12601), .ZN(n12600) );
  OR2_X1 U12590 ( .A1(n12407), .A2(n12405), .ZN(n12601) );
  NOR2_X1 U12591 ( .A1(n12188), .A2(n8042), .ZN(n12408) );
  NAND2_X1 U12592 ( .A1(n12405), .A2(n12407), .ZN(n12599) );
  NAND2_X1 U12593 ( .A1(n12602), .A2(n12603), .ZN(n12407) );
  NAND3_X1 U12594 ( .A1(a_24_), .A2(n12604), .A3(b_12_), .ZN(n12603) );
  NAND2_X1 U12595 ( .A1(n12403), .A2(n12402), .ZN(n12604) );
  OR2_X1 U12596 ( .A1(n12402), .A2(n12403), .ZN(n12602) );
  AND2_X1 U12597 ( .A1(n12605), .A2(n12606), .ZN(n12403) );
  NAND2_X1 U12598 ( .A1(n12400), .A2(n12607), .ZN(n12606) );
  OR2_X1 U12599 ( .A1(n12399), .A2(n12398), .ZN(n12607) );
  NOR2_X1 U12600 ( .A1(n12188), .A2(n8039), .ZN(n12400) );
  NAND2_X1 U12601 ( .A1(n12398), .A2(n12399), .ZN(n12605) );
  NAND2_X1 U12602 ( .A1(n12395), .A2(n12608), .ZN(n12399) );
  NAND2_X1 U12603 ( .A1(n12394), .A2(n12396), .ZN(n12608) );
  NAND2_X1 U12604 ( .A1(n12609), .A2(n12610), .ZN(n12396) );
  NAND2_X1 U12605 ( .A1(b_12_), .A2(a_26_), .ZN(n12610) );
  INV_X1 U12606 ( .A(n12611), .ZN(n12609) );
  XNOR2_X1 U12607 ( .A(n12612), .B(n12613), .ZN(n12394) );
  NAND2_X1 U12608 ( .A1(n12614), .A2(n12615), .ZN(n12612) );
  NAND2_X1 U12609 ( .A1(a_26_), .A2(n12611), .ZN(n12395) );
  NAND2_X1 U12610 ( .A1(n12367), .A2(n12616), .ZN(n12611) );
  NAND2_X1 U12611 ( .A1(n12366), .A2(n12368), .ZN(n12616) );
  NAND2_X1 U12612 ( .A1(n12617), .A2(n12618), .ZN(n12368) );
  NAND2_X1 U12613 ( .A1(b_12_), .A2(a_27_), .ZN(n12618) );
  INV_X1 U12614 ( .A(n12619), .ZN(n12617) );
  XNOR2_X1 U12615 ( .A(n12620), .B(n12621), .ZN(n12366) );
  XOR2_X1 U12616 ( .A(n12622), .B(n12623), .Z(n12620) );
  NAND2_X1 U12617 ( .A1(b_11_), .A2(a_28_), .ZN(n12622) );
  NAND2_X1 U12618 ( .A1(a_27_), .A2(n12619), .ZN(n12367) );
  NAND2_X1 U12619 ( .A1(n12624), .A2(n12625), .ZN(n12619) );
  NAND3_X1 U12620 ( .A1(a_28_), .A2(n12626), .A3(b_12_), .ZN(n12625) );
  NAND2_X1 U12621 ( .A1(n12376), .A2(n12374), .ZN(n12626) );
  OR2_X1 U12622 ( .A1(n12374), .A2(n12376), .ZN(n12624) );
  AND2_X1 U12623 ( .A1(n12627), .A2(n12628), .ZN(n12376) );
  NAND2_X1 U12624 ( .A1(n12390), .A2(n12629), .ZN(n12628) );
  OR2_X1 U12625 ( .A1(n12391), .A2(n12392), .ZN(n12629) );
  NOR2_X1 U12626 ( .A1(n12188), .A2(n7545), .ZN(n12390) );
  NAND2_X1 U12627 ( .A1(n12392), .A2(n12391), .ZN(n12627) );
  NAND2_X1 U12628 ( .A1(n12630), .A2(n12631), .ZN(n12391) );
  NAND2_X1 U12629 ( .A1(b_10_), .A2(n12632), .ZN(n12631) );
  NAND2_X1 U12630 ( .A1(n7527), .A2(n12633), .ZN(n12632) );
  NAND2_X1 U12631 ( .A1(a_31_), .A2(n7813), .ZN(n12633) );
  NAND2_X1 U12632 ( .A1(b_11_), .A2(n12634), .ZN(n12630) );
  NAND2_X1 U12633 ( .A1(n7531), .A2(n12635), .ZN(n12634) );
  NAND2_X1 U12634 ( .A1(a_30_), .A2(n8050), .ZN(n12635) );
  AND3_X1 U12635 ( .A1(b_12_), .A2(b_11_), .A3(n7494), .ZN(n12392) );
  XNOR2_X1 U12636 ( .A(n12636), .B(n12637), .ZN(n12374) );
  XOR2_X1 U12637 ( .A(n12638), .B(n12639), .Z(n12636) );
  XNOR2_X1 U12638 ( .A(n12640), .B(n12641), .ZN(n12398) );
  NAND2_X1 U12639 ( .A1(n12642), .A2(n12643), .ZN(n12640) );
  XNOR2_X1 U12640 ( .A(n12644), .B(n12645), .ZN(n12402) );
  XOR2_X1 U12641 ( .A(n12646), .B(n12647), .Z(n12644) );
  XNOR2_X1 U12642 ( .A(n12648), .B(n12649), .ZN(n12405) );
  XNOR2_X1 U12643 ( .A(n12650), .B(n12651), .ZN(n12648) );
  NOR2_X1 U12644 ( .A1(n8041), .A2(n7813), .ZN(n12651) );
  XNOR2_X1 U12645 ( .A(n12652), .B(n12653), .ZN(n12409) );
  XNOR2_X1 U12646 ( .A(n12654), .B(n12655), .ZN(n12653) );
  XNOR2_X1 U12647 ( .A(n12656), .B(n12657), .ZN(n12414) );
  XOR2_X1 U12648 ( .A(n12658), .B(n12659), .Z(n12657) );
  NAND2_X1 U12649 ( .A1(b_11_), .A2(a_22_), .ZN(n12659) );
  XNOR2_X1 U12650 ( .A(n12660), .B(n12661), .ZN(n12418) );
  XOR2_X1 U12651 ( .A(n12662), .B(n12663), .Z(n12660) );
  XNOR2_X1 U12652 ( .A(n12664), .B(n12665), .ZN(n12426) );
  NAND2_X1 U12653 ( .A1(n12666), .A2(n12667), .ZN(n12664) );
  XNOR2_X1 U12654 ( .A(n12668), .B(n12669), .ZN(n12430) );
  NAND2_X1 U12655 ( .A1(n12670), .A2(n12671), .ZN(n12668) );
  XOR2_X1 U12656 ( .A(n12672), .B(n12673), .Z(n12434) );
  XOR2_X1 U12657 ( .A(n12674), .B(n12675), .Z(n12673) );
  NAND2_X1 U12658 ( .A1(b_11_), .A2(a_17_), .ZN(n12675) );
  XOR2_X1 U12659 ( .A(n12676), .B(n12677), .Z(n12441) );
  XOR2_X1 U12660 ( .A(n12678), .B(n12679), .Z(n12676) );
  NOR2_X1 U12661 ( .A1(n8049), .A2(n7813), .ZN(n12679) );
  NOR2_X1 U12662 ( .A1(n12188), .A2(n8669), .ZN(n7801) );
  XNOR2_X1 U12663 ( .A(n12680), .B(n12681), .ZN(n12457) );
  XNOR2_X1 U12664 ( .A(n12682), .B(n12683), .ZN(n12680) );
  NOR2_X1 U12665 ( .A1(n7813), .A2(n8051), .ZN(n12683) );
  XNOR2_X1 U12666 ( .A(n12684), .B(n12685), .ZN(n12461) );
  XOR2_X1 U12667 ( .A(n12686), .B(n12687), .Z(n12685) );
  NAND2_X1 U12668 ( .A1(a_9_), .A2(b_11_), .ZN(n12687) );
  XNOR2_X1 U12669 ( .A(n12688), .B(n12689), .ZN(n12469) );
  XOR2_X1 U12670 ( .A(n12690), .B(n12691), .Z(n12689) );
  NAND2_X1 U12671 ( .A1(a_7_), .A2(b_11_), .ZN(n12691) );
  XNOR2_X1 U12672 ( .A(n12692), .B(n12693), .ZN(n12473) );
  XOR2_X1 U12673 ( .A(n12694), .B(n12695), .Z(n12692) );
  NOR2_X1 U12674 ( .A1(n7813), .A2(n7887), .ZN(n12695) );
  XNOR2_X1 U12675 ( .A(n12696), .B(n12697), .ZN(n12476) );
  XOR2_X1 U12676 ( .A(n12698), .B(n12699), .Z(n12697) );
  NAND2_X1 U12677 ( .A1(a_5_), .A2(b_11_), .ZN(n12699) );
  XNOR2_X1 U12678 ( .A(n12700), .B(n12701), .ZN(n12481) );
  XOR2_X1 U12679 ( .A(n12702), .B(n12703), .Z(n12701) );
  NAND2_X1 U12680 ( .A1(a_4_), .A2(b_11_), .ZN(n12703) );
  XNOR2_X1 U12681 ( .A(n12704), .B(n12705), .ZN(n12485) );
  XOR2_X1 U12682 ( .A(n12706), .B(n12707), .Z(n12704) );
  NOR2_X1 U12683 ( .A1(n7813), .A2(n7937), .ZN(n12707) );
  XNOR2_X1 U12684 ( .A(n12708), .B(n12709), .ZN(n12488) );
  XOR2_X1 U12685 ( .A(n12710), .B(n12711), .Z(n12709) );
  NAND2_X1 U12686 ( .A1(a_2_), .A2(b_11_), .ZN(n12711) );
  XNOR2_X1 U12687 ( .A(n12712), .B(n12713), .ZN(n12493) );
  XOR2_X1 U12688 ( .A(n12714), .B(n12715), .Z(n12712) );
  NOR2_X1 U12689 ( .A1(n7957), .A2(n7813), .ZN(n12715) );
  NAND2_X1 U12690 ( .A1(n12716), .A2(n12717), .ZN(n8198) );
  XNOR2_X1 U12691 ( .A(n12718), .B(n12719), .ZN(n8199) );
  XNOR2_X1 U12692 ( .A(n12720), .B(n12721), .ZN(n12719) );
  NAND2_X1 U12693 ( .A1(n12496), .A2(n12722), .ZN(n8171) );
  XOR2_X1 U12694 ( .A(n8193), .B(n8194), .Z(n12722) );
  NOR2_X1 U12695 ( .A1(n12717), .A2(n12716), .ZN(n12496) );
  AND2_X1 U12696 ( .A1(n12723), .A2(n12724), .ZN(n12716) );
  NAND2_X1 U12697 ( .A1(n12721), .A2(n12725), .ZN(n12724) );
  OR2_X1 U12698 ( .A1(n12720), .A2(n12718), .ZN(n12725) );
  NOR2_X1 U12699 ( .A1(n8942), .A2(n7813), .ZN(n12721) );
  NAND2_X1 U12700 ( .A1(n12718), .A2(n12720), .ZN(n12723) );
  NAND2_X1 U12701 ( .A1(n12726), .A2(n12727), .ZN(n12720) );
  NAND3_X1 U12702 ( .A1(a_1_), .A2(n12728), .A3(b_11_), .ZN(n12727) );
  OR2_X1 U12703 ( .A1(n12714), .A2(n12713), .ZN(n12728) );
  NAND2_X1 U12704 ( .A1(n12713), .A2(n12714), .ZN(n12726) );
  NAND2_X1 U12705 ( .A1(n12729), .A2(n12730), .ZN(n12714) );
  NAND3_X1 U12706 ( .A1(b_11_), .A2(n12731), .A3(a_2_), .ZN(n12730) );
  OR2_X1 U12707 ( .A1(n12710), .A2(n12708), .ZN(n12731) );
  NAND2_X1 U12708 ( .A1(n12708), .A2(n12710), .ZN(n12729) );
  NAND2_X1 U12709 ( .A1(n12732), .A2(n12733), .ZN(n12710) );
  NAND3_X1 U12710 ( .A1(b_11_), .A2(n12734), .A3(a_3_), .ZN(n12733) );
  OR2_X1 U12711 ( .A1(n12706), .A2(n12705), .ZN(n12734) );
  NAND2_X1 U12712 ( .A1(n12705), .A2(n12706), .ZN(n12732) );
  NAND2_X1 U12713 ( .A1(n12735), .A2(n12736), .ZN(n12706) );
  NAND3_X1 U12714 ( .A1(b_11_), .A2(n12737), .A3(a_4_), .ZN(n12736) );
  OR2_X1 U12715 ( .A1(n12702), .A2(n12700), .ZN(n12737) );
  NAND2_X1 U12716 ( .A1(n12700), .A2(n12702), .ZN(n12735) );
  NAND2_X1 U12717 ( .A1(n12738), .A2(n12739), .ZN(n12702) );
  NAND3_X1 U12718 ( .A1(b_11_), .A2(n12740), .A3(a_5_), .ZN(n12739) );
  OR2_X1 U12719 ( .A1(n12698), .A2(n12696), .ZN(n12740) );
  NAND2_X1 U12720 ( .A1(n12696), .A2(n12698), .ZN(n12738) );
  NAND2_X1 U12721 ( .A1(n12741), .A2(n12742), .ZN(n12698) );
  NAND3_X1 U12722 ( .A1(b_11_), .A2(n12743), .A3(a_6_), .ZN(n12742) );
  OR2_X1 U12723 ( .A1(n12694), .A2(n12693), .ZN(n12743) );
  NAND2_X1 U12724 ( .A1(n12693), .A2(n12694), .ZN(n12741) );
  NAND2_X1 U12725 ( .A1(n12744), .A2(n12745), .ZN(n12694) );
  NAND3_X1 U12726 ( .A1(b_11_), .A2(n12746), .A3(a_7_), .ZN(n12745) );
  OR2_X1 U12727 ( .A1(n12690), .A2(n12688), .ZN(n12746) );
  NAND2_X1 U12728 ( .A1(n12688), .A2(n12690), .ZN(n12744) );
  NAND2_X1 U12729 ( .A1(n12747), .A2(n12748), .ZN(n12690) );
  NAND3_X1 U12730 ( .A1(b_11_), .A2(n12749), .A3(a_8_), .ZN(n12748) );
  OR2_X1 U12731 ( .A1(n12524), .A2(n12522), .ZN(n12749) );
  NAND2_X1 U12732 ( .A1(n12522), .A2(n12524), .ZN(n12747) );
  NAND2_X1 U12733 ( .A1(n12750), .A2(n12751), .ZN(n12524) );
  NAND3_X1 U12734 ( .A1(b_11_), .A2(n12752), .A3(a_9_), .ZN(n12751) );
  OR2_X1 U12735 ( .A1(n12686), .A2(n12684), .ZN(n12752) );
  NAND2_X1 U12736 ( .A1(n12684), .A2(n12686), .ZN(n12750) );
  NAND2_X1 U12737 ( .A1(n12753), .A2(n12754), .ZN(n12686) );
  NAND3_X1 U12738 ( .A1(b_11_), .A2(n12755), .A3(a_10_), .ZN(n12754) );
  NAND2_X1 U12739 ( .A1(n12682), .A2(n12681), .ZN(n12755) );
  OR2_X1 U12740 ( .A1(n12681), .A2(n12682), .ZN(n12753) );
  AND2_X1 U12741 ( .A1(n12756), .A2(n12757), .ZN(n12682) );
  NAND2_X1 U12742 ( .A1(n12537), .A2(n12758), .ZN(n12757) );
  OR2_X1 U12743 ( .A1(n12538), .A2(n7808), .ZN(n12758) );
  XNOR2_X1 U12744 ( .A(n12759), .B(n12760), .ZN(n12537) );
  NAND2_X1 U12745 ( .A1(n12761), .A2(n12762), .ZN(n12759) );
  NAND2_X1 U12746 ( .A1(n7808), .A2(n12538), .ZN(n12756) );
  NAND2_X1 U12747 ( .A1(n12763), .A2(n12764), .ZN(n12538) );
  NAND3_X1 U12748 ( .A1(a_12_), .A2(n12765), .A3(b_11_), .ZN(n12764) );
  OR2_X1 U12749 ( .A1(n12545), .A2(n12544), .ZN(n12765) );
  NAND2_X1 U12750 ( .A1(n12544), .A2(n12545), .ZN(n12763) );
  NAND2_X1 U12751 ( .A1(n12766), .A2(n12767), .ZN(n12545) );
  NAND3_X1 U12752 ( .A1(a_13_), .A2(n12768), .A3(b_11_), .ZN(n12767) );
  OR2_X1 U12753 ( .A1(n12552), .A2(n12550), .ZN(n12768) );
  NAND2_X1 U12754 ( .A1(n12550), .A2(n12552), .ZN(n12766) );
  NAND2_X1 U12755 ( .A1(n12769), .A2(n12770), .ZN(n12552) );
  NAND3_X1 U12756 ( .A1(a_14_), .A2(n12771), .A3(b_11_), .ZN(n12770) );
  OR2_X1 U12757 ( .A1(n12678), .A2(n12677), .ZN(n12771) );
  NAND2_X1 U12758 ( .A1(n12677), .A2(n12678), .ZN(n12769) );
  NAND2_X1 U12759 ( .A1(n12772), .A2(n12773), .ZN(n12678) );
  NAND3_X1 U12760 ( .A1(a_15_), .A2(n12774), .A3(b_11_), .ZN(n12773) );
  OR2_X1 U12761 ( .A1(n12563), .A2(n12561), .ZN(n12774) );
  NAND2_X1 U12762 ( .A1(n12561), .A2(n12563), .ZN(n12772) );
  NAND2_X1 U12763 ( .A1(n12775), .A2(n12776), .ZN(n12563) );
  NAND3_X1 U12764 ( .A1(a_16_), .A2(n12777), .A3(b_11_), .ZN(n12776) );
  NAND2_X1 U12765 ( .A1(n12571), .A2(n12570), .ZN(n12777) );
  OR2_X1 U12766 ( .A1(n12570), .A2(n12571), .ZN(n12775) );
  AND2_X1 U12767 ( .A1(n12778), .A2(n12779), .ZN(n12571) );
  NAND3_X1 U12768 ( .A1(a_17_), .A2(n12780), .A3(b_11_), .ZN(n12779) );
  OR2_X1 U12769 ( .A1(n12674), .A2(n12672), .ZN(n12780) );
  NAND2_X1 U12770 ( .A1(n12672), .A2(n12674), .ZN(n12778) );
  NAND2_X1 U12771 ( .A1(n12670), .A2(n12781), .ZN(n12674) );
  NAND2_X1 U12772 ( .A1(n12669), .A2(n12671), .ZN(n12781) );
  NAND2_X1 U12773 ( .A1(n12782), .A2(n12783), .ZN(n12671) );
  NAND2_X1 U12774 ( .A1(b_11_), .A2(a_18_), .ZN(n12783) );
  INV_X1 U12775 ( .A(n12784), .ZN(n12782) );
  XNOR2_X1 U12776 ( .A(n12785), .B(n12786), .ZN(n12669) );
  XNOR2_X1 U12777 ( .A(n12787), .B(n12788), .ZN(n12786) );
  NAND2_X1 U12778 ( .A1(a_18_), .A2(n12784), .ZN(n12670) );
  NAND2_X1 U12779 ( .A1(n12666), .A2(n12789), .ZN(n12784) );
  NAND2_X1 U12780 ( .A1(n12665), .A2(n12667), .ZN(n12789) );
  NAND2_X1 U12781 ( .A1(n12790), .A2(n12791), .ZN(n12667) );
  NAND2_X1 U12782 ( .A1(b_11_), .A2(a_19_), .ZN(n12791) );
  INV_X1 U12783 ( .A(n12792), .ZN(n12790) );
  XNOR2_X1 U12784 ( .A(n12793), .B(n12794), .ZN(n12665) );
  XNOR2_X1 U12785 ( .A(n12795), .B(n12796), .ZN(n12794) );
  NAND2_X1 U12786 ( .A1(a_19_), .A2(n12792), .ZN(n12666) );
  NAND2_X1 U12787 ( .A1(n12797), .A2(n12798), .ZN(n12792) );
  NAND3_X1 U12788 ( .A1(a_20_), .A2(n12799), .A3(b_11_), .ZN(n12798) );
  OR2_X1 U12789 ( .A1(n12588), .A2(n12587), .ZN(n12799) );
  NAND2_X1 U12790 ( .A1(n12587), .A2(n12588), .ZN(n12797) );
  NAND2_X1 U12791 ( .A1(n12800), .A2(n12801), .ZN(n12588) );
  NAND2_X1 U12792 ( .A1(n12663), .A2(n12802), .ZN(n12801) );
  OR2_X1 U12793 ( .A1(n12662), .A2(n12661), .ZN(n12802) );
  NOR2_X1 U12794 ( .A1(n7813), .A2(n7665), .ZN(n12663) );
  NAND2_X1 U12795 ( .A1(n12661), .A2(n12662), .ZN(n12800) );
  NAND2_X1 U12796 ( .A1(n12803), .A2(n12804), .ZN(n12662) );
  NAND3_X1 U12797 ( .A1(a_22_), .A2(n12805), .A3(b_11_), .ZN(n12804) );
  OR2_X1 U12798 ( .A1(n12658), .A2(n12656), .ZN(n12805) );
  NAND2_X1 U12799 ( .A1(n12656), .A2(n12658), .ZN(n12803) );
  NAND2_X1 U12800 ( .A1(n12806), .A2(n12807), .ZN(n12658) );
  NAND2_X1 U12801 ( .A1(n12655), .A2(n12808), .ZN(n12807) );
  OR2_X1 U12802 ( .A1(n12654), .A2(n12652), .ZN(n12808) );
  NOR2_X1 U12803 ( .A1(n7813), .A2(n8042), .ZN(n12655) );
  NAND2_X1 U12804 ( .A1(n12652), .A2(n12654), .ZN(n12806) );
  NAND2_X1 U12805 ( .A1(n12809), .A2(n12810), .ZN(n12654) );
  NAND3_X1 U12806 ( .A1(a_24_), .A2(n12811), .A3(b_11_), .ZN(n12810) );
  NAND2_X1 U12807 ( .A1(n12650), .A2(n12649), .ZN(n12811) );
  OR2_X1 U12808 ( .A1(n12649), .A2(n12650), .ZN(n12809) );
  AND2_X1 U12809 ( .A1(n12812), .A2(n12813), .ZN(n12650) );
  NAND2_X1 U12810 ( .A1(n12647), .A2(n12814), .ZN(n12813) );
  OR2_X1 U12811 ( .A1(n12646), .A2(n12645), .ZN(n12814) );
  NOR2_X1 U12812 ( .A1(n7813), .A2(n8039), .ZN(n12647) );
  NAND2_X1 U12813 ( .A1(n12645), .A2(n12646), .ZN(n12812) );
  NAND2_X1 U12814 ( .A1(n12642), .A2(n12815), .ZN(n12646) );
  NAND2_X1 U12815 ( .A1(n12641), .A2(n12643), .ZN(n12815) );
  NAND2_X1 U12816 ( .A1(n12816), .A2(n12817), .ZN(n12643) );
  NAND2_X1 U12817 ( .A1(b_11_), .A2(a_26_), .ZN(n12817) );
  INV_X1 U12818 ( .A(n12818), .ZN(n12816) );
  XNOR2_X1 U12819 ( .A(n12819), .B(n12820), .ZN(n12641) );
  NAND2_X1 U12820 ( .A1(n12821), .A2(n12822), .ZN(n12819) );
  NAND2_X1 U12821 ( .A1(a_26_), .A2(n12818), .ZN(n12642) );
  NAND2_X1 U12822 ( .A1(n12614), .A2(n12823), .ZN(n12818) );
  NAND2_X1 U12823 ( .A1(n12613), .A2(n12615), .ZN(n12823) );
  NAND2_X1 U12824 ( .A1(n12824), .A2(n12825), .ZN(n12615) );
  NAND2_X1 U12825 ( .A1(b_11_), .A2(a_27_), .ZN(n12825) );
  INV_X1 U12826 ( .A(n12826), .ZN(n12824) );
  XNOR2_X1 U12827 ( .A(n12827), .B(n12828), .ZN(n12613) );
  XOR2_X1 U12828 ( .A(n12829), .B(n12830), .Z(n12827) );
  NAND2_X1 U12829 ( .A1(b_10_), .A2(a_28_), .ZN(n12829) );
  NAND2_X1 U12830 ( .A1(a_27_), .A2(n12826), .ZN(n12614) );
  NAND2_X1 U12831 ( .A1(n12831), .A2(n12832), .ZN(n12826) );
  NAND3_X1 U12832 ( .A1(a_28_), .A2(n12833), .A3(b_11_), .ZN(n12832) );
  NAND2_X1 U12833 ( .A1(n12623), .A2(n12621), .ZN(n12833) );
  OR2_X1 U12834 ( .A1(n12621), .A2(n12623), .ZN(n12831) );
  AND2_X1 U12835 ( .A1(n12834), .A2(n12835), .ZN(n12623) );
  NAND2_X1 U12836 ( .A1(n12637), .A2(n12836), .ZN(n12835) );
  OR2_X1 U12837 ( .A1(n12638), .A2(n12639), .ZN(n12836) );
  NOR2_X1 U12838 ( .A1(n7813), .A2(n7545), .ZN(n12637) );
  NAND2_X1 U12839 ( .A1(n12639), .A2(n12638), .ZN(n12834) );
  NAND2_X1 U12840 ( .A1(n12837), .A2(n12838), .ZN(n12638) );
  NAND2_X1 U12841 ( .A1(b_10_), .A2(n12839), .ZN(n12838) );
  NAND2_X1 U12842 ( .A1(n7531), .A2(n12840), .ZN(n12839) );
  NAND2_X1 U12843 ( .A1(a_30_), .A2(n7839), .ZN(n12840) );
  NAND2_X1 U12844 ( .A1(b_9_), .A2(n12841), .ZN(n12837) );
  NAND2_X1 U12845 ( .A1(n7527), .A2(n12842), .ZN(n12841) );
  NAND2_X1 U12846 ( .A1(a_31_), .A2(n8050), .ZN(n12842) );
  AND3_X1 U12847 ( .A1(b_10_), .A2(b_11_), .A3(n7494), .ZN(n12639) );
  XNOR2_X1 U12848 ( .A(n12843), .B(n12844), .ZN(n12621) );
  XOR2_X1 U12849 ( .A(n12845), .B(n12846), .Z(n12843) );
  XNOR2_X1 U12850 ( .A(n12847), .B(n12848), .ZN(n12645) );
  NAND2_X1 U12851 ( .A1(n12849), .A2(n12850), .ZN(n12847) );
  XNOR2_X1 U12852 ( .A(n12851), .B(n12852), .ZN(n12649) );
  XOR2_X1 U12853 ( .A(n12853), .B(n12854), .Z(n12851) );
  XNOR2_X1 U12854 ( .A(n12855), .B(n12856), .ZN(n12652) );
  XNOR2_X1 U12855 ( .A(n12857), .B(n12858), .ZN(n12855) );
  NOR2_X1 U12856 ( .A1(n8041), .A2(n8050), .ZN(n12858) );
  XNOR2_X1 U12857 ( .A(n12859), .B(n12860), .ZN(n12656) );
  XNOR2_X1 U12858 ( .A(n12861), .B(n12862), .ZN(n12860) );
  XNOR2_X1 U12859 ( .A(n12863), .B(n12864), .ZN(n12661) );
  XNOR2_X1 U12860 ( .A(n12865), .B(n12866), .ZN(n12863) );
  NOR2_X1 U12861 ( .A1(n7650), .A2(n8050), .ZN(n12866) );
  XNOR2_X1 U12862 ( .A(n12867), .B(n12868), .ZN(n12587) );
  XNOR2_X1 U12863 ( .A(n12869), .B(n12870), .ZN(n12867) );
  NOR2_X1 U12864 ( .A1(n7665), .A2(n8050), .ZN(n12870) );
  XNOR2_X1 U12865 ( .A(n12871), .B(n12872), .ZN(n12672) );
  XNOR2_X1 U12866 ( .A(n12873), .B(n12874), .ZN(n12872) );
  XNOR2_X1 U12867 ( .A(n12875), .B(n12876), .ZN(n12570) );
  XOR2_X1 U12868 ( .A(n12877), .B(n12878), .Z(n12875) );
  NOR2_X1 U12869 ( .A1(n7732), .A2(n8050), .ZN(n12878) );
  XNOR2_X1 U12870 ( .A(n12879), .B(n12880), .ZN(n12561) );
  NAND2_X1 U12871 ( .A1(n12881), .A2(n12882), .ZN(n12879) );
  XNOR2_X1 U12872 ( .A(n12883), .B(n12884), .ZN(n12677) );
  NAND2_X1 U12873 ( .A1(n12885), .A2(n12886), .ZN(n12883) );
  XNOR2_X1 U12874 ( .A(n12887), .B(n12888), .ZN(n12550) );
  XNOR2_X1 U12875 ( .A(n12889), .B(n12890), .ZN(n12888) );
  XNOR2_X1 U12876 ( .A(n12891), .B(n12892), .ZN(n12544) );
  XOR2_X1 U12877 ( .A(n12893), .B(n12894), .Z(n12892) );
  NAND2_X1 U12878 ( .A1(b_10_), .A2(a_13_), .ZN(n12894) );
  INV_X1 U12879 ( .A(n7995), .ZN(n7808) );
  NAND2_X1 U12880 ( .A1(a_11_), .A2(b_11_), .ZN(n7995) );
  XOR2_X1 U12881 ( .A(n12895), .B(n12896), .Z(n12681) );
  NAND2_X1 U12882 ( .A1(n12897), .A2(n12898), .ZN(n12895) );
  XOR2_X1 U12883 ( .A(n12899), .B(n12900), .Z(n12684) );
  XOR2_X1 U12884 ( .A(n12901), .B(n12902), .Z(n12899) );
  XNOR2_X1 U12885 ( .A(n12903), .B(n12904), .ZN(n12522) );
  NAND2_X1 U12886 ( .A1(n12905), .A2(n12906), .ZN(n12903) );
  XNOR2_X1 U12887 ( .A(n12907), .B(n12908), .ZN(n12688) );
  NAND2_X1 U12888 ( .A1(n12909), .A2(n12910), .ZN(n12907) );
  XNOR2_X1 U12889 ( .A(n12911), .B(n12912), .ZN(n12693) );
  XNOR2_X1 U12890 ( .A(n12913), .B(n12914), .ZN(n12912) );
  XNOR2_X1 U12891 ( .A(n12915), .B(n12916), .ZN(n12696) );
  XNOR2_X1 U12892 ( .A(n12917), .B(n12918), .ZN(n12915) );
  XOR2_X1 U12893 ( .A(n12919), .B(n12920), .Z(n12700) );
  XOR2_X1 U12894 ( .A(n12921), .B(n12922), .Z(n12919) );
  XNOR2_X1 U12895 ( .A(n12923), .B(n12924), .ZN(n12705) );
  XNOR2_X1 U12896 ( .A(n12925), .B(n12926), .ZN(n12924) );
  XNOR2_X1 U12897 ( .A(n12927), .B(n12928), .ZN(n12708) );
  XNOR2_X1 U12898 ( .A(n12929), .B(n12930), .ZN(n12927) );
  XNOR2_X1 U12899 ( .A(n12931), .B(n12932), .ZN(n12713) );
  XNOR2_X1 U12900 ( .A(n12933), .B(n12934), .ZN(n12932) );
  XNOR2_X1 U12901 ( .A(n12935), .B(n12936), .ZN(n12718) );
  XNOR2_X1 U12902 ( .A(n12937), .B(n12938), .ZN(n12935) );
  NOR2_X1 U12903 ( .A1(n7957), .A2(n8050), .ZN(n12938) );
  XNOR2_X1 U12904 ( .A(n12939), .B(n12940), .ZN(n12717) );
  XNOR2_X1 U12905 ( .A(n12941), .B(n12942), .ZN(n12940) );
  NAND2_X1 U12906 ( .A1(a_0_), .A2(b_10_), .ZN(n12942) );
  NAND2_X1 U12907 ( .A1(n12943), .A2(n12944), .ZN(n7500) );
  NAND2_X1 U12908 ( .A1(n12945), .A2(n12946), .ZN(n12944) );
  NAND2_X1 U12909 ( .A1(n8194), .A2(n8193), .ZN(n12943) );
  NAND4_X1 U12910 ( .A1(n8194), .A2(n12945), .A3(n8193), .A4(n12946), .ZN(
        n7499) );
  NAND2_X1 U12911 ( .A1(n12947), .A2(n12948), .ZN(n8193) );
  NAND3_X1 U12912 ( .A1(b_10_), .A2(n12949), .A3(a_0_), .ZN(n12948) );
  NAND2_X1 U12913 ( .A1(n12941), .A2(n12939), .ZN(n12949) );
  OR2_X1 U12914 ( .A1(n12939), .A2(n12941), .ZN(n12947) );
  AND2_X1 U12915 ( .A1(n12950), .A2(n12951), .ZN(n12941) );
  NAND3_X1 U12916 ( .A1(a_1_), .A2(n12952), .A3(b_10_), .ZN(n12951) );
  NAND2_X1 U12917 ( .A1(n12937), .A2(n12936), .ZN(n12952) );
  OR2_X1 U12918 ( .A1(n12936), .A2(n12937), .ZN(n12950) );
  AND2_X1 U12919 ( .A1(n12953), .A2(n12954), .ZN(n12937) );
  NAND2_X1 U12920 ( .A1(n12934), .A2(n12955), .ZN(n12954) );
  OR2_X1 U12921 ( .A1(n12933), .A2(n12931), .ZN(n12955) );
  NOR2_X1 U12922 ( .A1(n8056), .A2(n8050), .ZN(n12934) );
  NAND2_X1 U12923 ( .A1(n12931), .A2(n12933), .ZN(n12953) );
  NAND2_X1 U12924 ( .A1(n12956), .A2(n12957), .ZN(n12933) );
  NAND2_X1 U12925 ( .A1(n12929), .A2(n12958), .ZN(n12957) );
  NAND2_X1 U12926 ( .A1(n12930), .A2(n12928), .ZN(n12958) );
  NOR2_X1 U12927 ( .A1(n7937), .A2(n8050), .ZN(n12929) );
  OR2_X1 U12928 ( .A1(n12928), .A2(n12930), .ZN(n12956) );
  AND2_X1 U12929 ( .A1(n12959), .A2(n12960), .ZN(n12930) );
  NAND2_X1 U12930 ( .A1(n12926), .A2(n12961), .ZN(n12960) );
  OR2_X1 U12931 ( .A1(n12925), .A2(n12923), .ZN(n12961) );
  NOR2_X1 U12932 ( .A1(n7916), .A2(n8050), .ZN(n12926) );
  NAND2_X1 U12933 ( .A1(n12923), .A2(n12925), .ZN(n12959) );
  NAND2_X1 U12934 ( .A1(n12962), .A2(n12963), .ZN(n12925) );
  NAND2_X1 U12935 ( .A1(n12922), .A2(n12964), .ZN(n12963) );
  OR2_X1 U12936 ( .A1(n12920), .A2(n12921), .ZN(n12964) );
  NOR2_X1 U12937 ( .A1(n7908), .A2(n8050), .ZN(n12922) );
  NAND2_X1 U12938 ( .A1(n12920), .A2(n12921), .ZN(n12962) );
  NAND2_X1 U12939 ( .A1(n12965), .A2(n12966), .ZN(n12921) );
  NAND2_X1 U12940 ( .A1(n12918), .A2(n12967), .ZN(n12966) );
  NAND2_X1 U12941 ( .A1(n12917), .A2(n12916), .ZN(n12967) );
  NOR2_X1 U12942 ( .A1(n7887), .A2(n8050), .ZN(n12918) );
  OR2_X1 U12943 ( .A1(n12916), .A2(n12917), .ZN(n12965) );
  AND2_X1 U12944 ( .A1(n12968), .A2(n12969), .ZN(n12917) );
  NAND2_X1 U12945 ( .A1(n12914), .A2(n12970), .ZN(n12969) );
  OR2_X1 U12946 ( .A1(n12913), .A2(n12911), .ZN(n12970) );
  NOR2_X1 U12947 ( .A1(n7872), .A2(n8050), .ZN(n12914) );
  NAND2_X1 U12948 ( .A1(n12911), .A2(n12913), .ZN(n12968) );
  NAND2_X1 U12949 ( .A1(n12909), .A2(n12971), .ZN(n12913) );
  NAND2_X1 U12950 ( .A1(n12908), .A2(n12910), .ZN(n12971) );
  NAND2_X1 U12951 ( .A1(n12972), .A2(n12973), .ZN(n12910) );
  NAND2_X1 U12952 ( .A1(a_8_), .A2(b_10_), .ZN(n12973) );
  INV_X1 U12953 ( .A(n12974), .ZN(n12972) );
  XOR2_X1 U12954 ( .A(n12975), .B(n12976), .Z(n12908) );
  XOR2_X1 U12955 ( .A(n12977), .B(n7837), .Z(n12975) );
  NAND2_X1 U12956 ( .A1(a_8_), .A2(n12974), .ZN(n12909) );
  NAND2_X1 U12957 ( .A1(n12905), .A2(n12978), .ZN(n12974) );
  NAND2_X1 U12958 ( .A1(n12904), .A2(n12906), .ZN(n12978) );
  NAND2_X1 U12959 ( .A1(n12979), .A2(n12980), .ZN(n12906) );
  NAND2_X1 U12960 ( .A1(a_9_), .A2(b_10_), .ZN(n12980) );
  INV_X1 U12961 ( .A(n12981), .ZN(n12979) );
  XOR2_X1 U12962 ( .A(n12982), .B(n12983), .Z(n12904) );
  XOR2_X1 U12963 ( .A(n12984), .B(n12985), .Z(n12982) );
  NOR2_X1 U12964 ( .A1(n8051), .A2(n7839), .ZN(n12985) );
  NAND2_X1 U12965 ( .A1(a_9_), .A2(n12981), .ZN(n12905) );
  NAND2_X1 U12966 ( .A1(n12986), .A2(n12987), .ZN(n12981) );
  NAND2_X1 U12967 ( .A1(n12900), .A2(n12988), .ZN(n12987) );
  OR2_X1 U12968 ( .A1(n12901), .A2(n12902), .ZN(n12988) );
  XNOR2_X1 U12969 ( .A(n12989), .B(n12990), .ZN(n12900) );
  XOR2_X1 U12970 ( .A(n12991), .B(n12992), .Z(n12990) );
  NAND2_X1 U12971 ( .A1(b_9_), .A2(a_11_), .ZN(n12992) );
  NAND2_X1 U12972 ( .A1(n12902), .A2(n12901), .ZN(n12986) );
  NAND2_X1 U12973 ( .A1(n12897), .A2(n12993), .ZN(n12901) );
  NAND2_X1 U12974 ( .A1(n12896), .A2(n12898), .ZN(n12993) );
  NAND2_X1 U12975 ( .A1(n12994), .A2(n12995), .ZN(n12898) );
  NAND2_X1 U12976 ( .A1(b_10_), .A2(a_11_), .ZN(n12995) );
  INV_X1 U12977 ( .A(n12996), .ZN(n12994) );
  XOR2_X1 U12978 ( .A(n12997), .B(n12998), .Z(n12896) );
  XOR2_X1 U12979 ( .A(n12999), .B(n13000), .Z(n12997) );
  NOR2_X1 U12980 ( .A1(n8669), .A2(n7839), .ZN(n13000) );
  NAND2_X1 U12981 ( .A1(a_11_), .A2(n12996), .ZN(n12897) );
  NAND2_X1 U12982 ( .A1(n12761), .A2(n13001), .ZN(n12996) );
  NAND2_X1 U12983 ( .A1(n12760), .A2(n12762), .ZN(n13001) );
  NAND2_X1 U12984 ( .A1(n13002), .A2(n13003), .ZN(n12762) );
  NAND2_X1 U12985 ( .A1(b_10_), .A2(a_12_), .ZN(n13003) );
  INV_X1 U12986 ( .A(n13004), .ZN(n13002) );
  XNOR2_X1 U12987 ( .A(n13005), .B(n13006), .ZN(n12760) );
  XOR2_X1 U12988 ( .A(n13007), .B(n13008), .Z(n13006) );
  NAND2_X1 U12989 ( .A1(b_9_), .A2(a_13_), .ZN(n13008) );
  NAND2_X1 U12990 ( .A1(a_12_), .A2(n13004), .ZN(n12761) );
  NAND2_X1 U12991 ( .A1(n13009), .A2(n13010), .ZN(n13004) );
  NAND3_X1 U12992 ( .A1(a_13_), .A2(n13011), .A3(b_10_), .ZN(n13010) );
  OR2_X1 U12993 ( .A1(n12893), .A2(n12891), .ZN(n13011) );
  NAND2_X1 U12994 ( .A1(n12891), .A2(n12893), .ZN(n13009) );
  NAND2_X1 U12995 ( .A1(n13012), .A2(n13013), .ZN(n12893) );
  NAND2_X1 U12996 ( .A1(n12890), .A2(n13014), .ZN(n13013) );
  OR2_X1 U12997 ( .A1(n12889), .A2(n12887), .ZN(n13014) );
  NOR2_X1 U12998 ( .A1(n8050), .A2(n8049), .ZN(n12890) );
  NAND2_X1 U12999 ( .A1(n12887), .A2(n12889), .ZN(n13012) );
  NAND2_X1 U13000 ( .A1(n12885), .A2(n13015), .ZN(n12889) );
  NAND2_X1 U13001 ( .A1(n12884), .A2(n12886), .ZN(n13015) );
  NAND2_X1 U13002 ( .A1(n13016), .A2(n13017), .ZN(n12886) );
  NAND2_X1 U13003 ( .A1(b_10_), .A2(a_15_), .ZN(n13017) );
  INV_X1 U13004 ( .A(n13018), .ZN(n13016) );
  XNOR2_X1 U13005 ( .A(n13019), .B(n13020), .ZN(n12884) );
  XOR2_X1 U13006 ( .A(n13021), .B(n13022), .Z(n13020) );
  NAND2_X1 U13007 ( .A1(b_9_), .A2(a_16_), .ZN(n13022) );
  NAND2_X1 U13008 ( .A1(a_15_), .A2(n13018), .ZN(n12885) );
  NAND2_X1 U13009 ( .A1(n12881), .A2(n13023), .ZN(n13018) );
  NAND2_X1 U13010 ( .A1(n12880), .A2(n12882), .ZN(n13023) );
  NAND2_X1 U13011 ( .A1(n13024), .A2(n13025), .ZN(n12882) );
  NAND2_X1 U13012 ( .A1(b_10_), .A2(a_16_), .ZN(n13025) );
  INV_X1 U13013 ( .A(n13026), .ZN(n13024) );
  XNOR2_X1 U13014 ( .A(n13027), .B(n13028), .ZN(n12880) );
  XNOR2_X1 U13015 ( .A(n13029), .B(n13030), .ZN(n13027) );
  NOR2_X1 U13016 ( .A1(n7732), .A2(n7839), .ZN(n13030) );
  NAND2_X1 U13017 ( .A1(a_16_), .A2(n13026), .ZN(n12881) );
  NAND2_X1 U13018 ( .A1(n13031), .A2(n13032), .ZN(n13026) );
  NAND3_X1 U13019 ( .A1(a_17_), .A2(n13033), .A3(b_10_), .ZN(n13032) );
  OR2_X1 U13020 ( .A1(n12876), .A2(n12877), .ZN(n13033) );
  NAND2_X1 U13021 ( .A1(n12876), .A2(n12877), .ZN(n13031) );
  NAND2_X1 U13022 ( .A1(n13034), .A2(n13035), .ZN(n12877) );
  NAND2_X1 U13023 ( .A1(n12874), .A2(n13036), .ZN(n13035) );
  OR2_X1 U13024 ( .A1(n12873), .A2(n12871), .ZN(n13036) );
  NOR2_X1 U13025 ( .A1(n8050), .A2(n8047), .ZN(n12874) );
  NAND2_X1 U13026 ( .A1(n12871), .A2(n12873), .ZN(n13034) );
  NAND2_X1 U13027 ( .A1(n13037), .A2(n13038), .ZN(n12873) );
  NAND2_X1 U13028 ( .A1(n12788), .A2(n13039), .ZN(n13038) );
  OR2_X1 U13029 ( .A1(n12787), .A2(n12785), .ZN(n13039) );
  NOR2_X1 U13030 ( .A1(n8050), .A2(n8045), .ZN(n12788) );
  NAND2_X1 U13031 ( .A1(n12785), .A2(n12787), .ZN(n13037) );
  NAND2_X1 U13032 ( .A1(n13040), .A2(n13041), .ZN(n12787) );
  NAND2_X1 U13033 ( .A1(n12796), .A2(n13042), .ZN(n13041) );
  OR2_X1 U13034 ( .A1(n12795), .A2(n12793), .ZN(n13042) );
  NOR2_X1 U13035 ( .A1(n8050), .A2(n8044), .ZN(n12796) );
  NAND2_X1 U13036 ( .A1(n12793), .A2(n12795), .ZN(n13040) );
  NAND2_X1 U13037 ( .A1(n13043), .A2(n13044), .ZN(n12795) );
  NAND3_X1 U13038 ( .A1(a_21_), .A2(n13045), .A3(b_10_), .ZN(n13044) );
  NAND2_X1 U13039 ( .A1(n12869), .A2(n12868), .ZN(n13045) );
  OR2_X1 U13040 ( .A1(n12868), .A2(n12869), .ZN(n13043) );
  AND2_X1 U13041 ( .A1(n13046), .A2(n13047), .ZN(n12869) );
  NAND3_X1 U13042 ( .A1(a_22_), .A2(n13048), .A3(b_10_), .ZN(n13047) );
  NAND2_X1 U13043 ( .A1(n12865), .A2(n12864), .ZN(n13048) );
  OR2_X1 U13044 ( .A1(n12864), .A2(n12865), .ZN(n13046) );
  AND2_X1 U13045 ( .A1(n13049), .A2(n13050), .ZN(n12865) );
  NAND2_X1 U13046 ( .A1(n12862), .A2(n13051), .ZN(n13050) );
  OR2_X1 U13047 ( .A1(n12859), .A2(n12861), .ZN(n13051) );
  NOR2_X1 U13048 ( .A1(n8050), .A2(n8042), .ZN(n12862) );
  NAND2_X1 U13049 ( .A1(n12859), .A2(n12861), .ZN(n13049) );
  NAND2_X1 U13050 ( .A1(n13052), .A2(n13053), .ZN(n12861) );
  NAND3_X1 U13051 ( .A1(a_24_), .A2(n13054), .A3(b_10_), .ZN(n13053) );
  NAND2_X1 U13052 ( .A1(n12857), .A2(n12856), .ZN(n13054) );
  OR2_X1 U13053 ( .A1(n12856), .A2(n12857), .ZN(n13052) );
  AND2_X1 U13054 ( .A1(n13055), .A2(n13056), .ZN(n12857) );
  NAND2_X1 U13055 ( .A1(n12854), .A2(n13057), .ZN(n13056) );
  OR2_X1 U13056 ( .A1(n12852), .A2(n12853), .ZN(n13057) );
  NOR2_X1 U13057 ( .A1(n8050), .A2(n8039), .ZN(n12854) );
  NAND2_X1 U13058 ( .A1(n12852), .A2(n12853), .ZN(n13055) );
  NAND2_X1 U13059 ( .A1(n12849), .A2(n13058), .ZN(n12853) );
  NAND2_X1 U13060 ( .A1(n12848), .A2(n12850), .ZN(n13058) );
  NAND2_X1 U13061 ( .A1(n13059), .A2(n13060), .ZN(n12850) );
  NAND2_X1 U13062 ( .A1(b_10_), .A2(a_26_), .ZN(n13060) );
  INV_X1 U13063 ( .A(n13061), .ZN(n13059) );
  XNOR2_X1 U13064 ( .A(n13062), .B(n13063), .ZN(n12848) );
  NAND2_X1 U13065 ( .A1(n13064), .A2(n13065), .ZN(n13062) );
  NAND2_X1 U13066 ( .A1(a_26_), .A2(n13061), .ZN(n12849) );
  NAND2_X1 U13067 ( .A1(n12821), .A2(n13066), .ZN(n13061) );
  NAND2_X1 U13068 ( .A1(n12820), .A2(n12822), .ZN(n13066) );
  NAND2_X1 U13069 ( .A1(n13067), .A2(n13068), .ZN(n12822) );
  NAND2_X1 U13070 ( .A1(b_10_), .A2(a_27_), .ZN(n13068) );
  INV_X1 U13071 ( .A(n13069), .ZN(n13067) );
  XNOR2_X1 U13072 ( .A(n13070), .B(n13071), .ZN(n12820) );
  XOR2_X1 U13073 ( .A(n13072), .B(n13073), .Z(n13070) );
  NAND2_X1 U13074 ( .A1(b_9_), .A2(a_28_), .ZN(n13072) );
  NAND2_X1 U13075 ( .A1(a_27_), .A2(n13069), .ZN(n12821) );
  NAND2_X1 U13076 ( .A1(n13074), .A2(n13075), .ZN(n13069) );
  NAND3_X1 U13077 ( .A1(a_28_), .A2(n13076), .A3(b_10_), .ZN(n13075) );
  NAND2_X1 U13078 ( .A1(n12830), .A2(n12828), .ZN(n13076) );
  OR2_X1 U13079 ( .A1(n12828), .A2(n12830), .ZN(n13074) );
  AND2_X1 U13080 ( .A1(n13077), .A2(n13078), .ZN(n12830) );
  NAND2_X1 U13081 ( .A1(n12844), .A2(n13079), .ZN(n13078) );
  OR2_X1 U13082 ( .A1(n12845), .A2(n12846), .ZN(n13079) );
  NOR2_X1 U13083 ( .A1(n8050), .A2(n7545), .ZN(n12844) );
  NAND2_X1 U13084 ( .A1(n12846), .A2(n12845), .ZN(n13077) );
  NAND2_X1 U13085 ( .A1(n13080), .A2(n13081), .ZN(n12845) );
  NAND2_X1 U13086 ( .A1(b_8_), .A2(n13082), .ZN(n13081) );
  NAND2_X1 U13087 ( .A1(n7527), .A2(n13083), .ZN(n13082) );
  NAND2_X1 U13088 ( .A1(a_31_), .A2(n7839), .ZN(n13083) );
  NAND2_X1 U13089 ( .A1(b_9_), .A2(n13084), .ZN(n13080) );
  NAND2_X1 U13090 ( .A1(n7531), .A2(n13085), .ZN(n13084) );
  NAND2_X1 U13091 ( .A1(a_30_), .A2(n13086), .ZN(n13085) );
  AND3_X1 U13092 ( .A1(b_9_), .A2(b_10_), .A3(n7494), .ZN(n12846) );
  XNOR2_X1 U13093 ( .A(n13087), .B(n13088), .ZN(n12828) );
  XOR2_X1 U13094 ( .A(n13089), .B(n13090), .Z(n13087) );
  XNOR2_X1 U13095 ( .A(n13091), .B(n13092), .ZN(n12852) );
  NAND2_X1 U13096 ( .A1(n13093), .A2(n13094), .ZN(n13091) );
  XNOR2_X1 U13097 ( .A(n13095), .B(n13096), .ZN(n12856) );
  XOR2_X1 U13098 ( .A(n13097), .B(n13098), .Z(n13095) );
  XNOR2_X1 U13099 ( .A(n13099), .B(n13100), .ZN(n12859) );
  XNOR2_X1 U13100 ( .A(n13101), .B(n13102), .ZN(n13099) );
  NOR2_X1 U13101 ( .A1(n8041), .A2(n7839), .ZN(n13102) );
  XOR2_X1 U13102 ( .A(n13103), .B(n13104), .Z(n12864) );
  XNOR2_X1 U13103 ( .A(n13105), .B(n13106), .ZN(n13104) );
  XNOR2_X1 U13104 ( .A(n13107), .B(n13108), .ZN(n12868) );
  XOR2_X1 U13105 ( .A(n13109), .B(n13110), .Z(n13107) );
  XOR2_X1 U13106 ( .A(n13111), .B(n13112), .Z(n12793) );
  XOR2_X1 U13107 ( .A(n13113), .B(n13114), .Z(n13111) );
  NOR2_X1 U13108 ( .A1(n7665), .A2(n7839), .ZN(n13114) );
  XOR2_X1 U13109 ( .A(n13115), .B(n13116), .Z(n12785) );
  XOR2_X1 U13110 ( .A(n13117), .B(n13118), .Z(n13115) );
  NOR2_X1 U13111 ( .A1(n8044), .A2(n7839), .ZN(n13118) );
  XNOR2_X1 U13112 ( .A(n13119), .B(n13120), .ZN(n12871) );
  XOR2_X1 U13113 ( .A(n13121), .B(n13122), .Z(n13120) );
  NAND2_X1 U13114 ( .A1(b_9_), .A2(a_19_), .ZN(n13122) );
  XNOR2_X1 U13115 ( .A(n13123), .B(n13124), .ZN(n12876) );
  XNOR2_X1 U13116 ( .A(n13125), .B(n13126), .ZN(n13123) );
  NOR2_X1 U13117 ( .A1(n8047), .A2(n7839), .ZN(n13126) );
  XOR2_X1 U13118 ( .A(n13127), .B(n13128), .Z(n12887) );
  XOR2_X1 U13119 ( .A(n13129), .B(n13130), .Z(n13127) );
  NOR2_X1 U13120 ( .A1(n7754), .A2(n7839), .ZN(n13130) );
  XNOR2_X1 U13121 ( .A(n13131), .B(n13132), .ZN(n12891) );
  XOR2_X1 U13122 ( .A(n13133), .B(n13134), .Z(n13132) );
  NAND2_X1 U13123 ( .A1(b_9_), .A2(a_14_), .ZN(n13134) );
  INV_X1 U13124 ( .A(n7830), .ZN(n12902) );
  NAND2_X1 U13125 ( .A1(b_10_), .A2(a_10_), .ZN(n7830) );
  XOR2_X1 U13126 ( .A(n13135), .B(n13136), .Z(n12911) );
  XNOR2_X1 U13127 ( .A(n13137), .B(n13138), .ZN(n13135) );
  NAND2_X1 U13128 ( .A1(a_8_), .A2(b_9_), .ZN(n13137) );
  XOR2_X1 U13129 ( .A(n13139), .B(n13140), .Z(n12916) );
  XOR2_X1 U13130 ( .A(n13141), .B(n13142), .Z(n13140) );
  NAND2_X1 U13131 ( .A1(a_7_), .A2(b_9_), .ZN(n13142) );
  XNOR2_X1 U13132 ( .A(n13143), .B(n13144), .ZN(n12920) );
  XNOR2_X1 U13133 ( .A(n13145), .B(n13146), .ZN(n13143) );
  NOR2_X1 U13134 ( .A1(n7839), .A2(n7887), .ZN(n13146) );
  XOR2_X1 U13135 ( .A(n13147), .B(n13148), .Z(n12923) );
  XOR2_X1 U13136 ( .A(n13149), .B(n13150), .Z(n13147) );
  NOR2_X1 U13137 ( .A1(n7839), .A2(n7908), .ZN(n13150) );
  XNOR2_X1 U13138 ( .A(n13151), .B(n13152), .ZN(n12928) );
  XOR2_X1 U13139 ( .A(n13153), .B(n13154), .Z(n13151) );
  NOR2_X1 U13140 ( .A1(n7839), .A2(n7916), .ZN(n13154) );
  XOR2_X1 U13141 ( .A(n13155), .B(n13156), .Z(n12931) );
  XOR2_X1 U13142 ( .A(n13157), .B(n13158), .Z(n13155) );
  NOR2_X1 U13143 ( .A1(n7839), .A2(n7937), .ZN(n13158) );
  XNOR2_X1 U13144 ( .A(n13159), .B(n13160), .ZN(n12936) );
  XOR2_X1 U13145 ( .A(n13161), .B(n13162), .Z(n13159) );
  NOR2_X1 U13146 ( .A1(n7839), .A2(n8056), .ZN(n13162) );
  XNOR2_X1 U13147 ( .A(n13163), .B(n13164), .ZN(n12939) );
  XOR2_X1 U13148 ( .A(n13165), .B(n13166), .Z(n13163) );
  NAND2_X1 U13149 ( .A1(n13167), .A2(n13168), .ZN(n12945) );
  XOR2_X1 U13150 ( .A(n13169), .B(n13170), .Z(n8194) );
  XOR2_X1 U13151 ( .A(n13171), .B(n13172), .Z(n13169) );
  NAND2_X1 U13152 ( .A1(n13173), .A2(n12946), .ZN(n7505) );
  INV_X1 U13153 ( .A(n13174), .ZN(n12946) );
  XNOR2_X1 U13154 ( .A(n13175), .B(n13176), .ZN(n13173) );
  NAND2_X1 U13155 ( .A1(n13174), .A2(n13177), .ZN(n7504) );
  XOR2_X1 U13156 ( .A(n13175), .B(n13176), .Z(n13177) );
  NOR2_X1 U13157 ( .A1(n13168), .A2(n13167), .ZN(n13174) );
  AND2_X1 U13158 ( .A1(n13178), .A2(n13179), .ZN(n13167) );
  NAND2_X1 U13159 ( .A1(n13172), .A2(n13180), .ZN(n13179) );
  OR2_X1 U13160 ( .A1(n13170), .A2(n13171), .ZN(n13180) );
  NOR2_X1 U13161 ( .A1(n8942), .A2(n7839), .ZN(n13172) );
  NAND2_X1 U13162 ( .A1(n13170), .A2(n13171), .ZN(n13178) );
  NAND2_X1 U13163 ( .A1(n13181), .A2(n13182), .ZN(n13171) );
  NAND2_X1 U13164 ( .A1(n13166), .A2(n13183), .ZN(n13182) );
  OR2_X1 U13165 ( .A1(n13164), .A2(n13165), .ZN(n13183) );
  NOR2_X1 U13166 ( .A1(n7839), .A2(n7957), .ZN(n13166) );
  NAND2_X1 U13167 ( .A1(n13164), .A2(n13165), .ZN(n13181) );
  NAND2_X1 U13168 ( .A1(n13184), .A2(n13185), .ZN(n13165) );
  NAND3_X1 U13169 ( .A1(b_9_), .A2(n13186), .A3(a_2_), .ZN(n13185) );
  OR2_X1 U13170 ( .A1(n13160), .A2(n13161), .ZN(n13186) );
  NAND2_X1 U13171 ( .A1(n13160), .A2(n13161), .ZN(n13184) );
  NAND2_X1 U13172 ( .A1(n13187), .A2(n13188), .ZN(n13161) );
  NAND3_X1 U13173 ( .A1(b_9_), .A2(n13189), .A3(a_3_), .ZN(n13188) );
  OR2_X1 U13174 ( .A1(n13156), .A2(n13157), .ZN(n13189) );
  NAND2_X1 U13175 ( .A1(n13156), .A2(n13157), .ZN(n13187) );
  NAND2_X1 U13176 ( .A1(n13190), .A2(n13191), .ZN(n13157) );
  NAND3_X1 U13177 ( .A1(b_9_), .A2(n13192), .A3(a_4_), .ZN(n13191) );
  OR2_X1 U13178 ( .A1(n13152), .A2(n13153), .ZN(n13192) );
  NAND2_X1 U13179 ( .A1(n13152), .A2(n13153), .ZN(n13190) );
  NAND2_X1 U13180 ( .A1(n13193), .A2(n13194), .ZN(n13153) );
  NAND3_X1 U13181 ( .A1(b_9_), .A2(n13195), .A3(a_5_), .ZN(n13194) );
  OR2_X1 U13182 ( .A1(n13148), .A2(n13149), .ZN(n13195) );
  NAND2_X1 U13183 ( .A1(n13148), .A2(n13149), .ZN(n13193) );
  NAND2_X1 U13184 ( .A1(n13196), .A2(n13197), .ZN(n13149) );
  NAND3_X1 U13185 ( .A1(b_9_), .A2(n13198), .A3(a_6_), .ZN(n13197) );
  NAND2_X1 U13186 ( .A1(n13145), .A2(n13144), .ZN(n13198) );
  OR2_X1 U13187 ( .A1(n13144), .A2(n13145), .ZN(n13196) );
  AND2_X1 U13188 ( .A1(n13199), .A2(n13200), .ZN(n13145) );
  NAND3_X1 U13189 ( .A1(b_9_), .A2(n13201), .A3(a_7_), .ZN(n13200) );
  OR2_X1 U13190 ( .A1(n13139), .A2(n13141), .ZN(n13201) );
  NAND2_X1 U13191 ( .A1(n13139), .A2(n13141), .ZN(n13199) );
  NAND2_X1 U13192 ( .A1(n13202), .A2(n13203), .ZN(n13141) );
  NAND3_X1 U13193 ( .A1(b_9_), .A2(n13204), .A3(a_8_), .ZN(n13203) );
  OR2_X1 U13194 ( .A1(n13136), .A2(n13138), .ZN(n13204) );
  NAND2_X1 U13195 ( .A1(n13136), .A2(n13138), .ZN(n13202) );
  NAND2_X1 U13196 ( .A1(n13205), .A2(n13206), .ZN(n13138) );
  NAND2_X1 U13197 ( .A1(n12976), .A2(n13207), .ZN(n13206) );
  OR2_X1 U13198 ( .A1(n12977), .A2(n7837), .ZN(n13207) );
  XNOR2_X1 U13199 ( .A(n13208), .B(n13209), .ZN(n12976) );
  XNOR2_X1 U13200 ( .A(n13210), .B(n13211), .ZN(n13209) );
  NAND2_X1 U13201 ( .A1(n7837), .A2(n12977), .ZN(n13205) );
  NAND2_X1 U13202 ( .A1(n13212), .A2(n13213), .ZN(n12977) );
  NAND3_X1 U13203 ( .A1(a_10_), .A2(n13214), .A3(b_9_), .ZN(n13213) );
  OR2_X1 U13204 ( .A1(n12983), .A2(n12984), .ZN(n13214) );
  NAND2_X1 U13205 ( .A1(n12983), .A2(n12984), .ZN(n13212) );
  NAND2_X1 U13206 ( .A1(n13215), .A2(n13216), .ZN(n12984) );
  NAND3_X1 U13207 ( .A1(a_11_), .A2(n13217), .A3(b_9_), .ZN(n13216) );
  OR2_X1 U13208 ( .A1(n12991), .A2(n12989), .ZN(n13217) );
  NAND2_X1 U13209 ( .A1(n12989), .A2(n12991), .ZN(n13215) );
  NAND2_X1 U13210 ( .A1(n13218), .A2(n13219), .ZN(n12991) );
  NAND3_X1 U13211 ( .A1(a_12_), .A2(n13220), .A3(b_9_), .ZN(n13219) );
  OR2_X1 U13212 ( .A1(n12998), .A2(n12999), .ZN(n13220) );
  NAND2_X1 U13213 ( .A1(n12998), .A2(n12999), .ZN(n13218) );
  NAND2_X1 U13214 ( .A1(n13221), .A2(n13222), .ZN(n12999) );
  NAND3_X1 U13215 ( .A1(a_13_), .A2(n13223), .A3(b_9_), .ZN(n13222) );
  OR2_X1 U13216 ( .A1(n13007), .A2(n13005), .ZN(n13223) );
  NAND2_X1 U13217 ( .A1(n13005), .A2(n13007), .ZN(n13221) );
  NAND2_X1 U13218 ( .A1(n13224), .A2(n13225), .ZN(n13007) );
  NAND3_X1 U13219 ( .A1(a_14_), .A2(n13226), .A3(b_9_), .ZN(n13225) );
  OR2_X1 U13220 ( .A1(n13131), .A2(n13133), .ZN(n13226) );
  NAND2_X1 U13221 ( .A1(n13131), .A2(n13133), .ZN(n13224) );
  NAND2_X1 U13222 ( .A1(n13227), .A2(n13228), .ZN(n13133) );
  NAND3_X1 U13223 ( .A1(a_15_), .A2(n13229), .A3(b_9_), .ZN(n13228) );
  OR2_X1 U13224 ( .A1(n13128), .A2(n13129), .ZN(n13229) );
  NAND2_X1 U13225 ( .A1(n13128), .A2(n13129), .ZN(n13227) );
  NAND2_X1 U13226 ( .A1(n13230), .A2(n13231), .ZN(n13129) );
  NAND3_X1 U13227 ( .A1(a_16_), .A2(n13232), .A3(b_9_), .ZN(n13231) );
  OR2_X1 U13228 ( .A1(n13021), .A2(n13019), .ZN(n13232) );
  NAND2_X1 U13229 ( .A1(n13019), .A2(n13021), .ZN(n13230) );
  NAND2_X1 U13230 ( .A1(n13233), .A2(n13234), .ZN(n13021) );
  NAND3_X1 U13231 ( .A1(a_17_), .A2(n13235), .A3(b_9_), .ZN(n13234) );
  NAND2_X1 U13232 ( .A1(n13029), .A2(n13028), .ZN(n13235) );
  OR2_X1 U13233 ( .A1(n13028), .A2(n13029), .ZN(n13233) );
  AND2_X1 U13234 ( .A1(n13236), .A2(n13237), .ZN(n13029) );
  NAND3_X1 U13235 ( .A1(a_18_), .A2(n13238), .A3(b_9_), .ZN(n13237) );
  NAND2_X1 U13236 ( .A1(n13125), .A2(n13124), .ZN(n13238) );
  OR2_X1 U13237 ( .A1(n13124), .A2(n13125), .ZN(n13236) );
  AND2_X1 U13238 ( .A1(n13239), .A2(n13240), .ZN(n13125) );
  NAND3_X1 U13239 ( .A1(a_19_), .A2(n13241), .A3(b_9_), .ZN(n13240) );
  OR2_X1 U13240 ( .A1(n13119), .A2(n13121), .ZN(n13241) );
  NAND2_X1 U13241 ( .A1(n13119), .A2(n13121), .ZN(n13239) );
  NAND2_X1 U13242 ( .A1(n13242), .A2(n13243), .ZN(n13121) );
  NAND3_X1 U13243 ( .A1(a_20_), .A2(n13244), .A3(b_9_), .ZN(n13243) );
  OR2_X1 U13244 ( .A1(n13116), .A2(n13117), .ZN(n13244) );
  NAND2_X1 U13245 ( .A1(n13116), .A2(n13117), .ZN(n13242) );
  NAND2_X1 U13246 ( .A1(n13245), .A2(n13246), .ZN(n13117) );
  NAND3_X1 U13247 ( .A1(a_21_), .A2(n13247), .A3(b_9_), .ZN(n13246) );
  OR2_X1 U13248 ( .A1(n13112), .A2(n13113), .ZN(n13247) );
  NAND2_X1 U13249 ( .A1(n13112), .A2(n13113), .ZN(n13245) );
  NAND2_X1 U13250 ( .A1(n13248), .A2(n13249), .ZN(n13113) );
  NAND2_X1 U13251 ( .A1(n13110), .A2(n13250), .ZN(n13249) );
  OR2_X1 U13252 ( .A1(n13108), .A2(n13109), .ZN(n13250) );
  NOR2_X1 U13253 ( .A1(n7839), .A2(n7650), .ZN(n13110) );
  NAND2_X1 U13254 ( .A1(n13108), .A2(n13109), .ZN(n13248) );
  NAND2_X1 U13255 ( .A1(n13251), .A2(n13252), .ZN(n13109) );
  NAND2_X1 U13256 ( .A1(n13106), .A2(n13253), .ZN(n13252) );
  OR2_X1 U13257 ( .A1(n13103), .A2(n13105), .ZN(n13253) );
  NOR2_X1 U13258 ( .A1(n7839), .A2(n8042), .ZN(n13106) );
  NAND2_X1 U13259 ( .A1(n13103), .A2(n13105), .ZN(n13251) );
  NAND2_X1 U13260 ( .A1(n13254), .A2(n13255), .ZN(n13105) );
  NAND3_X1 U13261 ( .A1(a_24_), .A2(n13256), .A3(b_9_), .ZN(n13255) );
  NAND2_X1 U13262 ( .A1(n13101), .A2(n13100), .ZN(n13256) );
  OR2_X1 U13263 ( .A1(n13100), .A2(n13101), .ZN(n13254) );
  AND2_X1 U13264 ( .A1(n13257), .A2(n13258), .ZN(n13101) );
  NAND2_X1 U13265 ( .A1(n13098), .A2(n13259), .ZN(n13258) );
  OR2_X1 U13266 ( .A1(n13096), .A2(n13097), .ZN(n13259) );
  NOR2_X1 U13267 ( .A1(n7839), .A2(n8039), .ZN(n13098) );
  NAND2_X1 U13268 ( .A1(n13096), .A2(n13097), .ZN(n13257) );
  NAND2_X1 U13269 ( .A1(n13093), .A2(n13260), .ZN(n13097) );
  NAND2_X1 U13270 ( .A1(n13092), .A2(n13094), .ZN(n13260) );
  NAND2_X1 U13271 ( .A1(n13261), .A2(n13262), .ZN(n13094) );
  NAND2_X1 U13272 ( .A1(b_9_), .A2(a_26_), .ZN(n13262) );
  INV_X1 U13273 ( .A(n13263), .ZN(n13261) );
  XNOR2_X1 U13274 ( .A(n13264), .B(n13265), .ZN(n13092) );
  NAND2_X1 U13275 ( .A1(n13266), .A2(n13267), .ZN(n13264) );
  NAND2_X1 U13276 ( .A1(a_26_), .A2(n13263), .ZN(n13093) );
  NAND2_X1 U13277 ( .A1(n13064), .A2(n13268), .ZN(n13263) );
  NAND2_X1 U13278 ( .A1(n13063), .A2(n13065), .ZN(n13268) );
  NAND2_X1 U13279 ( .A1(n13269), .A2(n13270), .ZN(n13065) );
  NAND2_X1 U13280 ( .A1(b_9_), .A2(a_27_), .ZN(n13270) );
  INV_X1 U13281 ( .A(n13271), .ZN(n13269) );
  XNOR2_X1 U13282 ( .A(n13272), .B(n13273), .ZN(n13063) );
  XOR2_X1 U13283 ( .A(n13274), .B(n13275), .Z(n13272) );
  NAND2_X1 U13284 ( .A1(b_8_), .A2(a_28_), .ZN(n13274) );
  NAND2_X1 U13285 ( .A1(a_27_), .A2(n13271), .ZN(n13064) );
  NAND2_X1 U13286 ( .A1(n13276), .A2(n13277), .ZN(n13271) );
  NAND3_X1 U13287 ( .A1(a_28_), .A2(n13278), .A3(b_9_), .ZN(n13277) );
  NAND2_X1 U13288 ( .A1(n13073), .A2(n13071), .ZN(n13278) );
  OR2_X1 U13289 ( .A1(n13071), .A2(n13073), .ZN(n13276) );
  AND2_X1 U13290 ( .A1(n13279), .A2(n13280), .ZN(n13073) );
  NAND2_X1 U13291 ( .A1(n13088), .A2(n13281), .ZN(n13280) );
  OR2_X1 U13292 ( .A1(n13089), .A2(n13090), .ZN(n13281) );
  NOR2_X1 U13293 ( .A1(n7839), .A2(n7545), .ZN(n13088) );
  NAND2_X1 U13294 ( .A1(n13090), .A2(n13089), .ZN(n13279) );
  NAND2_X1 U13295 ( .A1(n13282), .A2(n13283), .ZN(n13089) );
  NAND2_X1 U13296 ( .A1(b_7_), .A2(n13284), .ZN(n13283) );
  NAND2_X1 U13297 ( .A1(n7527), .A2(n13285), .ZN(n13284) );
  NAND2_X1 U13298 ( .A1(a_31_), .A2(n13086), .ZN(n13285) );
  NAND2_X1 U13299 ( .A1(b_8_), .A2(n13286), .ZN(n13282) );
  NAND2_X1 U13300 ( .A1(n7531), .A2(n13287), .ZN(n13286) );
  NAND2_X1 U13301 ( .A1(a_30_), .A2(n7874), .ZN(n13287) );
  AND3_X1 U13302 ( .A1(b_8_), .A2(b_9_), .A3(n7494), .ZN(n13090) );
  XNOR2_X1 U13303 ( .A(n13288), .B(n13289), .ZN(n13071) );
  XOR2_X1 U13304 ( .A(n13290), .B(n13291), .Z(n13288) );
  XNOR2_X1 U13305 ( .A(n13292), .B(n13293), .ZN(n13096) );
  NAND2_X1 U13306 ( .A1(n13294), .A2(n13295), .ZN(n13292) );
  XNOR2_X1 U13307 ( .A(n13296), .B(n13297), .ZN(n13100) );
  XOR2_X1 U13308 ( .A(n13298), .B(n13299), .Z(n13296) );
  XNOR2_X1 U13309 ( .A(n13300), .B(n13301), .ZN(n13103) );
  XNOR2_X1 U13310 ( .A(n13302), .B(n13303), .ZN(n13300) );
  NOR2_X1 U13311 ( .A1(n8041), .A2(n13086), .ZN(n13303) );
  XNOR2_X1 U13312 ( .A(n13304), .B(n13305), .ZN(n13108) );
  XOR2_X1 U13313 ( .A(n13306), .B(n13307), .Z(n13305) );
  NAND2_X1 U13314 ( .A1(b_8_), .A2(a_23_), .ZN(n13307) );
  XNOR2_X1 U13315 ( .A(n13308), .B(n13309), .ZN(n13112) );
  XNOR2_X1 U13316 ( .A(n13310), .B(n13311), .ZN(n13309) );
  XNOR2_X1 U13317 ( .A(n13312), .B(n13313), .ZN(n13116) );
  XNOR2_X1 U13318 ( .A(n13314), .B(n13315), .ZN(n13312) );
  XNOR2_X1 U13319 ( .A(n13316), .B(n13317), .ZN(n13119) );
  XNOR2_X1 U13320 ( .A(n13318), .B(n13319), .ZN(n13316) );
  XNOR2_X1 U13321 ( .A(n13320), .B(n13321), .ZN(n13124) );
  XOR2_X1 U13322 ( .A(n13322), .B(n13323), .Z(n13320) );
  XOR2_X1 U13323 ( .A(n13324), .B(n13325), .Z(n13028) );
  XOR2_X1 U13324 ( .A(n13326), .B(n13327), .Z(n13325) );
  NAND2_X1 U13325 ( .A1(b_8_), .A2(a_18_), .ZN(n13327) );
  XNOR2_X1 U13326 ( .A(n13328), .B(n13329), .ZN(n13019) );
  NAND2_X1 U13327 ( .A1(n13330), .A2(n13331), .ZN(n13328) );
  XNOR2_X1 U13328 ( .A(n13332), .B(n13333), .ZN(n13128) );
  NAND2_X1 U13329 ( .A1(n13334), .A2(n13335), .ZN(n13332) );
  XNOR2_X1 U13330 ( .A(n13336), .B(n13337), .ZN(n13131) );
  XNOR2_X1 U13331 ( .A(n13338), .B(n13339), .ZN(n13336) );
  XNOR2_X1 U13332 ( .A(n13340), .B(n13341), .ZN(n13005) );
  XOR2_X1 U13333 ( .A(n13342), .B(n13343), .Z(n13341) );
  NAND2_X1 U13334 ( .A1(b_8_), .A2(a_14_), .ZN(n13343) );
  XNOR2_X1 U13335 ( .A(n13344), .B(n13345), .ZN(n12998) );
  XNOR2_X1 U13336 ( .A(n13346), .B(n13347), .ZN(n13344) );
  XNOR2_X1 U13337 ( .A(n13348), .B(n13349), .ZN(n12989) );
  XNOR2_X1 U13338 ( .A(n13350), .B(n13351), .ZN(n13349) );
  XNOR2_X1 U13339 ( .A(n13352), .B(n13353), .ZN(n12983) );
  XNOR2_X1 U13340 ( .A(n13354), .B(n13355), .ZN(n13352) );
  INV_X1 U13341 ( .A(n7991), .ZN(n7837) );
  NAND2_X1 U13342 ( .A1(a_9_), .A2(b_9_), .ZN(n7991) );
  XNOR2_X1 U13343 ( .A(n13356), .B(n13357), .ZN(n13136) );
  XNOR2_X1 U13344 ( .A(n13358), .B(n13359), .ZN(n13356) );
  XOR2_X1 U13345 ( .A(n13360), .B(n13361), .Z(n13139) );
  XNOR2_X1 U13346 ( .A(n13362), .B(n7857), .ZN(n13361) );
  XNOR2_X1 U13347 ( .A(n13363), .B(n13364), .ZN(n13144) );
  XOR2_X1 U13348 ( .A(n13365), .B(n13366), .Z(n13363) );
  XNOR2_X1 U13349 ( .A(n13367), .B(n13368), .ZN(n13148) );
  XNOR2_X1 U13350 ( .A(n13369), .B(n13370), .ZN(n13368) );
  XNOR2_X1 U13351 ( .A(n13371), .B(n13372), .ZN(n13152) );
  XNOR2_X1 U13352 ( .A(n13373), .B(n13374), .ZN(n13371) );
  NOR2_X1 U13353 ( .A1(n13086), .A2(n7908), .ZN(n13374) );
  XNOR2_X1 U13354 ( .A(n13375), .B(n13376), .ZN(n13156) );
  XOR2_X1 U13355 ( .A(n13377), .B(n13378), .Z(n13376) );
  NAND2_X1 U13356 ( .A1(a_4_), .A2(b_8_), .ZN(n13378) );
  XOR2_X1 U13357 ( .A(n13379), .B(n13380), .Z(n13160) );
  XOR2_X1 U13358 ( .A(n13381), .B(n13382), .Z(n13379) );
  NOR2_X1 U13359 ( .A1(n13086), .A2(n7937), .ZN(n13382) );
  XOR2_X1 U13360 ( .A(n13383), .B(n13384), .Z(n13164) );
  XNOR2_X1 U13361 ( .A(n13385), .B(n13386), .ZN(n13384) );
  NAND2_X1 U13362 ( .A1(a_2_), .A2(b_8_), .ZN(n13386) );
  XOR2_X1 U13363 ( .A(n13387), .B(n13388), .Z(n13170) );
  XOR2_X1 U13364 ( .A(n13389), .B(n13390), .Z(n13387) );
  NOR2_X1 U13365 ( .A1(n7957), .A2(n13086), .ZN(n13390) );
  XNOR2_X1 U13366 ( .A(n13391), .B(n13392), .ZN(n13168) );
  XOR2_X1 U13367 ( .A(n13393), .B(n13394), .Z(n13391) );
  NOR2_X1 U13368 ( .A1(n13086), .A2(n8942), .ZN(n13394) );
  NAND2_X1 U13369 ( .A1(n13395), .A2(n13396), .ZN(n7510) );
  NAND2_X1 U13370 ( .A1(n13397), .A2(n13398), .ZN(n13396) );
  NAND2_X1 U13371 ( .A1(n13176), .A2(n13175), .ZN(n13395) );
  NAND4_X1 U13372 ( .A1(n13176), .A2(n13397), .A3(n13175), .A4(n13398), .ZN(
        n7509) );
  NAND2_X1 U13373 ( .A1(n13399), .A2(n13400), .ZN(n13175) );
  NAND3_X1 U13374 ( .A1(b_8_), .A2(n13401), .A3(a_0_), .ZN(n13400) );
  OR2_X1 U13375 ( .A1(n13393), .A2(n13392), .ZN(n13401) );
  NAND2_X1 U13376 ( .A1(n13392), .A2(n13393), .ZN(n13399) );
  NAND2_X1 U13377 ( .A1(n13402), .A2(n13403), .ZN(n13393) );
  NAND3_X1 U13378 ( .A1(a_1_), .A2(n13404), .A3(b_8_), .ZN(n13403) );
  OR2_X1 U13379 ( .A1(n13389), .A2(n13388), .ZN(n13404) );
  NAND2_X1 U13380 ( .A1(n13388), .A2(n13389), .ZN(n13402) );
  NAND2_X1 U13381 ( .A1(n13405), .A2(n13406), .ZN(n13389) );
  NAND3_X1 U13382 ( .A1(b_8_), .A2(n13407), .A3(a_2_), .ZN(n13406) );
  NAND2_X1 U13383 ( .A1(n13385), .A2(n13383), .ZN(n13407) );
  OR2_X1 U13384 ( .A1(n13383), .A2(n13385), .ZN(n13405) );
  AND2_X1 U13385 ( .A1(n13408), .A2(n13409), .ZN(n13385) );
  NAND3_X1 U13386 ( .A1(b_8_), .A2(n13410), .A3(a_3_), .ZN(n13409) );
  OR2_X1 U13387 ( .A1(n13381), .A2(n13380), .ZN(n13410) );
  NAND2_X1 U13388 ( .A1(n13380), .A2(n13381), .ZN(n13408) );
  NAND2_X1 U13389 ( .A1(n13411), .A2(n13412), .ZN(n13381) );
  NAND3_X1 U13390 ( .A1(b_8_), .A2(n13413), .A3(a_4_), .ZN(n13412) );
  OR2_X1 U13391 ( .A1(n13377), .A2(n13375), .ZN(n13413) );
  NAND2_X1 U13392 ( .A1(n13375), .A2(n13377), .ZN(n13411) );
  NAND2_X1 U13393 ( .A1(n13414), .A2(n13415), .ZN(n13377) );
  NAND3_X1 U13394 ( .A1(b_8_), .A2(n13416), .A3(a_5_), .ZN(n13415) );
  NAND2_X1 U13395 ( .A1(n13373), .A2(n13372), .ZN(n13416) );
  OR2_X1 U13396 ( .A1(n13372), .A2(n13373), .ZN(n13414) );
  AND2_X1 U13397 ( .A1(n13417), .A2(n13418), .ZN(n13373) );
  NAND2_X1 U13398 ( .A1(n13370), .A2(n13419), .ZN(n13418) );
  OR2_X1 U13399 ( .A1(n13369), .A2(n13367), .ZN(n13419) );
  NOR2_X1 U13400 ( .A1(n7887), .A2(n13086), .ZN(n13370) );
  NAND2_X1 U13401 ( .A1(n13367), .A2(n13369), .ZN(n13417) );
  NAND2_X1 U13402 ( .A1(n13420), .A2(n13421), .ZN(n13369) );
  NAND2_X1 U13403 ( .A1(n13366), .A2(n13422), .ZN(n13421) );
  NAND2_X1 U13404 ( .A1(n13364), .A2(n13365), .ZN(n13422) );
  NOR2_X1 U13405 ( .A1(n7872), .A2(n13086), .ZN(n13366) );
  OR2_X1 U13406 ( .A1(n13364), .A2(n13365), .ZN(n13420) );
  NAND2_X1 U13407 ( .A1(n13423), .A2(n13424), .ZN(n13365) );
  NAND2_X1 U13408 ( .A1(n13360), .A2(n13425), .ZN(n13424) );
  NAND2_X1 U13409 ( .A1(n7857), .A2(n13362), .ZN(n13425) );
  XNOR2_X1 U13410 ( .A(n13426), .B(n13427), .ZN(n13360) );
  XOR2_X1 U13411 ( .A(n13428), .B(n13429), .Z(n13426) );
  NOR2_X1 U13412 ( .A1(n8052), .A2(n7874), .ZN(n13429) );
  OR2_X1 U13413 ( .A1(n13362), .A2(n7857), .ZN(n13423) );
  NOR2_X1 U13414 ( .A1(n13086), .A2(n8686), .ZN(n7857) );
  NAND2_X1 U13415 ( .A1(n13430), .A2(n13431), .ZN(n13362) );
  NAND2_X1 U13416 ( .A1(n13359), .A2(n13432), .ZN(n13431) );
  NAND2_X1 U13417 ( .A1(n13358), .A2(n13357), .ZN(n13432) );
  NOR2_X1 U13418 ( .A1(n13086), .A2(n8052), .ZN(n13359) );
  OR2_X1 U13419 ( .A1(n13357), .A2(n13358), .ZN(n13430) );
  AND2_X1 U13420 ( .A1(n13433), .A2(n13434), .ZN(n13358) );
  NAND2_X1 U13421 ( .A1(n13211), .A2(n13435), .ZN(n13434) );
  OR2_X1 U13422 ( .A1(n13210), .A2(n13208), .ZN(n13435) );
  NOR2_X1 U13423 ( .A1(n13086), .A2(n8051), .ZN(n13211) );
  NAND2_X1 U13424 ( .A1(n13208), .A2(n13210), .ZN(n13433) );
  NAND2_X1 U13425 ( .A1(n13436), .A2(n13437), .ZN(n13210) );
  NAND2_X1 U13426 ( .A1(n13355), .A2(n13438), .ZN(n13437) );
  NAND2_X1 U13427 ( .A1(n13354), .A2(n13353), .ZN(n13438) );
  NOR2_X1 U13428 ( .A1(n13086), .A2(n7811), .ZN(n13355) );
  OR2_X1 U13429 ( .A1(n13353), .A2(n13354), .ZN(n13436) );
  AND2_X1 U13430 ( .A1(n13439), .A2(n13440), .ZN(n13354) );
  NAND2_X1 U13431 ( .A1(n13351), .A2(n13441), .ZN(n13440) );
  OR2_X1 U13432 ( .A1(n13348), .A2(n13350), .ZN(n13441) );
  NOR2_X1 U13433 ( .A1(n13086), .A2(n8669), .ZN(n13351) );
  NAND2_X1 U13434 ( .A1(n13348), .A2(n13350), .ZN(n13439) );
  NAND2_X1 U13435 ( .A1(n13442), .A2(n13443), .ZN(n13350) );
  NAND2_X1 U13436 ( .A1(n13347), .A2(n13444), .ZN(n13443) );
  NAND2_X1 U13437 ( .A1(n13346), .A2(n13345), .ZN(n13444) );
  NOR2_X1 U13438 ( .A1(n13086), .A2(n7789), .ZN(n13347) );
  OR2_X1 U13439 ( .A1(n13345), .A2(n13346), .ZN(n13442) );
  AND2_X1 U13440 ( .A1(n13445), .A2(n13446), .ZN(n13346) );
  NAND3_X1 U13441 ( .A1(a_14_), .A2(n13447), .A3(b_8_), .ZN(n13446) );
  OR2_X1 U13442 ( .A1(n13340), .A2(n13342), .ZN(n13447) );
  NAND2_X1 U13443 ( .A1(n13340), .A2(n13342), .ZN(n13445) );
  NAND2_X1 U13444 ( .A1(n13448), .A2(n13449), .ZN(n13342) );
  NAND2_X1 U13445 ( .A1(n13339), .A2(n13450), .ZN(n13449) );
  NAND2_X1 U13446 ( .A1(n13338), .A2(n13337), .ZN(n13450) );
  NOR2_X1 U13447 ( .A1(n13086), .A2(n7754), .ZN(n13339) );
  OR2_X1 U13448 ( .A1(n13337), .A2(n13338), .ZN(n13448) );
  AND2_X1 U13449 ( .A1(n13334), .A2(n13451), .ZN(n13338) );
  NAND2_X1 U13450 ( .A1(n13333), .A2(n13335), .ZN(n13451) );
  NAND2_X1 U13451 ( .A1(n13452), .A2(n13453), .ZN(n13335) );
  NAND2_X1 U13452 ( .A1(b_8_), .A2(a_16_), .ZN(n13453) );
  INV_X1 U13453 ( .A(n13454), .ZN(n13452) );
  XNOR2_X1 U13454 ( .A(n13455), .B(n13456), .ZN(n13333) );
  XNOR2_X1 U13455 ( .A(n13457), .B(n13458), .ZN(n13455) );
  NOR2_X1 U13456 ( .A1(n7732), .A2(n7874), .ZN(n13458) );
  NAND2_X1 U13457 ( .A1(a_16_), .A2(n13454), .ZN(n13334) );
  NAND2_X1 U13458 ( .A1(n13330), .A2(n13459), .ZN(n13454) );
  NAND2_X1 U13459 ( .A1(n13329), .A2(n13331), .ZN(n13459) );
  NAND2_X1 U13460 ( .A1(n13460), .A2(n13461), .ZN(n13331) );
  NAND2_X1 U13461 ( .A1(b_8_), .A2(a_17_), .ZN(n13461) );
  INV_X1 U13462 ( .A(n13462), .ZN(n13460) );
  XNOR2_X1 U13463 ( .A(n13463), .B(n13464), .ZN(n13329) );
  XOR2_X1 U13464 ( .A(n13465), .B(n13466), .Z(n13464) );
  NAND2_X1 U13465 ( .A1(b_7_), .A2(a_18_), .ZN(n13466) );
  NAND2_X1 U13466 ( .A1(a_17_), .A2(n13462), .ZN(n13330) );
  NAND2_X1 U13467 ( .A1(n13467), .A2(n13468), .ZN(n13462) );
  NAND3_X1 U13468 ( .A1(a_18_), .A2(n13469), .A3(b_8_), .ZN(n13468) );
  OR2_X1 U13469 ( .A1(n13324), .A2(n13326), .ZN(n13469) );
  NAND2_X1 U13470 ( .A1(n13324), .A2(n13326), .ZN(n13467) );
  NAND2_X1 U13471 ( .A1(n13470), .A2(n13471), .ZN(n13326) );
  NAND2_X1 U13472 ( .A1(n13323), .A2(n13472), .ZN(n13471) );
  OR2_X1 U13473 ( .A1(n13321), .A2(n13322), .ZN(n13472) );
  NOR2_X1 U13474 ( .A1(n13086), .A2(n8045), .ZN(n13323) );
  NAND2_X1 U13475 ( .A1(n13321), .A2(n13322), .ZN(n13470) );
  NAND2_X1 U13476 ( .A1(n13473), .A2(n13474), .ZN(n13322) );
  NAND2_X1 U13477 ( .A1(n13319), .A2(n13475), .ZN(n13474) );
  NAND2_X1 U13478 ( .A1(n13318), .A2(n13317), .ZN(n13475) );
  NOR2_X1 U13479 ( .A1(n13086), .A2(n8044), .ZN(n13319) );
  OR2_X1 U13480 ( .A1(n13317), .A2(n13318), .ZN(n13473) );
  AND2_X1 U13481 ( .A1(n13476), .A2(n13477), .ZN(n13318) );
  NAND2_X1 U13482 ( .A1(n13315), .A2(n13478), .ZN(n13477) );
  NAND2_X1 U13483 ( .A1(n13314), .A2(n13313), .ZN(n13478) );
  NOR2_X1 U13484 ( .A1(n13086), .A2(n7665), .ZN(n13315) );
  OR2_X1 U13485 ( .A1(n13313), .A2(n13314), .ZN(n13476) );
  AND2_X1 U13486 ( .A1(n13479), .A2(n13480), .ZN(n13314) );
  NAND2_X1 U13487 ( .A1(n13311), .A2(n13481), .ZN(n13480) );
  OR2_X1 U13488 ( .A1(n13310), .A2(n13308), .ZN(n13481) );
  NOR2_X1 U13489 ( .A1(n13086), .A2(n7650), .ZN(n13311) );
  NAND2_X1 U13490 ( .A1(n13308), .A2(n13310), .ZN(n13479) );
  NAND2_X1 U13491 ( .A1(n13482), .A2(n13483), .ZN(n13310) );
  NAND3_X1 U13492 ( .A1(a_23_), .A2(n13484), .A3(b_8_), .ZN(n13483) );
  OR2_X1 U13493 ( .A1(n13306), .A2(n13304), .ZN(n13484) );
  NAND2_X1 U13494 ( .A1(n13304), .A2(n13306), .ZN(n13482) );
  NAND2_X1 U13495 ( .A1(n13485), .A2(n13486), .ZN(n13306) );
  NAND3_X1 U13496 ( .A1(a_24_), .A2(n13487), .A3(b_8_), .ZN(n13486) );
  NAND2_X1 U13497 ( .A1(n13302), .A2(n13301), .ZN(n13487) );
  OR2_X1 U13498 ( .A1(n13301), .A2(n13302), .ZN(n13485) );
  AND2_X1 U13499 ( .A1(n13488), .A2(n13489), .ZN(n13302) );
  NAND2_X1 U13500 ( .A1(n13299), .A2(n13490), .ZN(n13489) );
  OR2_X1 U13501 ( .A1(n13297), .A2(n13298), .ZN(n13490) );
  NOR2_X1 U13502 ( .A1(n13086), .A2(n8039), .ZN(n13299) );
  NAND2_X1 U13503 ( .A1(n13297), .A2(n13298), .ZN(n13488) );
  NAND2_X1 U13504 ( .A1(n13294), .A2(n13491), .ZN(n13298) );
  NAND2_X1 U13505 ( .A1(n13293), .A2(n13295), .ZN(n13491) );
  NAND2_X1 U13506 ( .A1(n13492), .A2(n13493), .ZN(n13295) );
  NAND2_X1 U13507 ( .A1(b_8_), .A2(a_26_), .ZN(n13493) );
  INV_X1 U13508 ( .A(n13494), .ZN(n13492) );
  XNOR2_X1 U13509 ( .A(n13495), .B(n13496), .ZN(n13293) );
  NAND2_X1 U13510 ( .A1(n13497), .A2(n13498), .ZN(n13495) );
  NAND2_X1 U13511 ( .A1(a_26_), .A2(n13494), .ZN(n13294) );
  NAND2_X1 U13512 ( .A1(n13266), .A2(n13499), .ZN(n13494) );
  NAND2_X1 U13513 ( .A1(n13265), .A2(n13267), .ZN(n13499) );
  NAND2_X1 U13514 ( .A1(n13500), .A2(n13501), .ZN(n13267) );
  NAND2_X1 U13515 ( .A1(b_8_), .A2(a_27_), .ZN(n13501) );
  INV_X1 U13516 ( .A(n13502), .ZN(n13500) );
  XNOR2_X1 U13517 ( .A(n13503), .B(n13504), .ZN(n13265) );
  XOR2_X1 U13518 ( .A(n13505), .B(n13506), .Z(n13503) );
  NAND2_X1 U13519 ( .A1(b_7_), .A2(a_28_), .ZN(n13505) );
  NAND2_X1 U13520 ( .A1(a_27_), .A2(n13502), .ZN(n13266) );
  NAND2_X1 U13521 ( .A1(n13507), .A2(n13508), .ZN(n13502) );
  NAND3_X1 U13522 ( .A1(a_28_), .A2(n13509), .A3(b_8_), .ZN(n13508) );
  NAND2_X1 U13523 ( .A1(n13275), .A2(n13273), .ZN(n13509) );
  OR2_X1 U13524 ( .A1(n13273), .A2(n13275), .ZN(n13507) );
  AND2_X1 U13525 ( .A1(n13510), .A2(n13511), .ZN(n13275) );
  NAND2_X1 U13526 ( .A1(n13289), .A2(n13512), .ZN(n13511) );
  OR2_X1 U13527 ( .A1(n13290), .A2(n13291), .ZN(n13512) );
  NOR2_X1 U13528 ( .A1(n13086), .A2(n7545), .ZN(n13289) );
  NAND2_X1 U13529 ( .A1(n13291), .A2(n13290), .ZN(n13510) );
  NAND2_X1 U13530 ( .A1(n13513), .A2(n13514), .ZN(n13290) );
  NAND2_X1 U13531 ( .A1(b_6_), .A2(n13515), .ZN(n13514) );
  NAND2_X1 U13532 ( .A1(n7527), .A2(n13516), .ZN(n13515) );
  NAND2_X1 U13533 ( .A1(a_31_), .A2(n7874), .ZN(n13516) );
  NAND2_X1 U13534 ( .A1(b_7_), .A2(n13517), .ZN(n13513) );
  NAND2_X1 U13535 ( .A1(n7531), .A2(n13518), .ZN(n13517) );
  NAND2_X1 U13536 ( .A1(a_30_), .A2(n8053), .ZN(n13518) );
  AND3_X1 U13537 ( .A1(b_8_), .A2(b_7_), .A3(n7494), .ZN(n13291) );
  XNOR2_X1 U13538 ( .A(n13519), .B(n13520), .ZN(n13273) );
  XOR2_X1 U13539 ( .A(n13521), .B(n13522), .Z(n13519) );
  XNOR2_X1 U13540 ( .A(n13523), .B(n13524), .ZN(n13297) );
  NAND2_X1 U13541 ( .A1(n13525), .A2(n13526), .ZN(n13523) );
  XNOR2_X1 U13542 ( .A(n13527), .B(n13528), .ZN(n13301) );
  XOR2_X1 U13543 ( .A(n13529), .B(n13530), .Z(n13527) );
  XOR2_X1 U13544 ( .A(n13531), .B(n13532), .Z(n13304) );
  XOR2_X1 U13545 ( .A(n13533), .B(n13534), .Z(n13531) );
  XOR2_X1 U13546 ( .A(n13535), .B(n13536), .Z(n13308) );
  XOR2_X1 U13547 ( .A(n13537), .B(n13538), .Z(n13535) );
  NOR2_X1 U13548 ( .A1(n8042), .A2(n7874), .ZN(n13538) );
  XOR2_X1 U13549 ( .A(n13539), .B(n13540), .Z(n13313) );
  NAND2_X1 U13550 ( .A1(n13541), .A2(n13542), .ZN(n13539) );
  XNOR2_X1 U13551 ( .A(n13543), .B(n13544), .ZN(n13317) );
  XOR2_X1 U13552 ( .A(n13545), .B(n13546), .Z(n13543) );
  NOR2_X1 U13553 ( .A1(n7665), .A2(n7874), .ZN(n13546) );
  XNOR2_X1 U13554 ( .A(n13547), .B(n13548), .ZN(n13321) );
  XNOR2_X1 U13555 ( .A(n13549), .B(n13550), .ZN(n13547) );
  NOR2_X1 U13556 ( .A1(n8044), .A2(n7874), .ZN(n13550) );
  XNOR2_X1 U13557 ( .A(n13551), .B(n13552), .ZN(n13324) );
  XOR2_X1 U13558 ( .A(n13553), .B(n13554), .Z(n13552) );
  NAND2_X1 U13559 ( .A1(b_7_), .A2(a_19_), .ZN(n13554) );
  XNOR2_X1 U13560 ( .A(n13555), .B(n13556), .ZN(n13337) );
  XOR2_X1 U13561 ( .A(n13557), .B(n13558), .Z(n13555) );
  NOR2_X1 U13562 ( .A1(n8438), .A2(n7874), .ZN(n13558) );
  XNOR2_X1 U13563 ( .A(n13559), .B(n13560), .ZN(n13340) );
  XOR2_X1 U13564 ( .A(n13561), .B(n13562), .Z(n13560) );
  NAND2_X1 U13565 ( .A1(b_7_), .A2(a_15_), .ZN(n13562) );
  XNOR2_X1 U13566 ( .A(n13563), .B(n13564), .ZN(n13345) );
  XOR2_X1 U13567 ( .A(n13565), .B(n13566), .Z(n13563) );
  NOR2_X1 U13568 ( .A1(n8049), .A2(n7874), .ZN(n13566) );
  XNOR2_X1 U13569 ( .A(n13567), .B(n13568), .ZN(n13348) );
  XOR2_X1 U13570 ( .A(n13569), .B(n13570), .Z(n13568) );
  NAND2_X1 U13571 ( .A1(b_7_), .A2(a_13_), .ZN(n13570) );
  XNOR2_X1 U13572 ( .A(n13571), .B(n13572), .ZN(n13353) );
  XOR2_X1 U13573 ( .A(n13573), .B(n13574), .Z(n13571) );
  NOR2_X1 U13574 ( .A1(n8669), .A2(n7874), .ZN(n13574) );
  XOR2_X1 U13575 ( .A(n13575), .B(n13576), .Z(n13208) );
  XOR2_X1 U13576 ( .A(n13577), .B(n13578), .Z(n13575) );
  NOR2_X1 U13577 ( .A1(n7811), .A2(n7874), .ZN(n13578) );
  XNOR2_X1 U13578 ( .A(n13579), .B(n13580), .ZN(n13357) );
  XOR2_X1 U13579 ( .A(n13581), .B(n13582), .Z(n13579) );
  NOR2_X1 U13580 ( .A1(n8051), .A2(n7874), .ZN(n13582) );
  XNOR2_X1 U13581 ( .A(n13583), .B(n13584), .ZN(n13364) );
  XOR2_X1 U13582 ( .A(n13585), .B(n13586), .Z(n13583) );
  NOR2_X1 U13583 ( .A1(n8686), .A2(n7874), .ZN(n13586) );
  XOR2_X1 U13584 ( .A(n13587), .B(n13588), .Z(n13367) );
  XOR2_X1 U13585 ( .A(n13589), .B(n7869), .Z(n13587) );
  XNOR2_X1 U13586 ( .A(n13590), .B(n13591), .ZN(n13372) );
  XOR2_X1 U13587 ( .A(n13592), .B(n13593), .Z(n13590) );
  NOR2_X1 U13588 ( .A1(n7874), .A2(n7887), .ZN(n13593) );
  XOR2_X1 U13589 ( .A(n13594), .B(n13595), .Z(n13375) );
  XOR2_X1 U13590 ( .A(n13596), .B(n13597), .Z(n13594) );
  NOR2_X1 U13591 ( .A1(n7874), .A2(n7908), .ZN(n13597) );
  XOR2_X1 U13592 ( .A(n13598), .B(n13599), .Z(n13380) );
  XOR2_X1 U13593 ( .A(n13600), .B(n13601), .Z(n13598) );
  NOR2_X1 U13594 ( .A1(n7874), .A2(n7916), .ZN(n13601) );
  XNOR2_X1 U13595 ( .A(n13602), .B(n13603), .ZN(n13383) );
  XOR2_X1 U13596 ( .A(n13604), .B(n13605), .Z(n13602) );
  NOR2_X1 U13597 ( .A1(n7874), .A2(n7937), .ZN(n13605) );
  XOR2_X1 U13598 ( .A(n13606), .B(n13607), .Z(n13388) );
  XOR2_X1 U13599 ( .A(n13608), .B(n13609), .Z(n13606) );
  NOR2_X1 U13600 ( .A1(n7874), .A2(n8056), .ZN(n13609) );
  XOR2_X1 U13601 ( .A(n13610), .B(n13611), .Z(n13392) );
  XOR2_X1 U13602 ( .A(n13612), .B(n13613), .Z(n13610) );
  NAND2_X1 U13603 ( .A1(n13614), .A2(n13615), .ZN(n13397) );
  XOR2_X1 U13604 ( .A(n13616), .B(n13617), .Z(n13176) );
  XOR2_X1 U13605 ( .A(n13618), .B(n13619), .Z(n13616) );
  NAND2_X1 U13606 ( .A1(n13620), .A2(n13398), .ZN(n7515) );
  INV_X1 U13607 ( .A(n13621), .ZN(n13398) );
  XNOR2_X1 U13608 ( .A(n13622), .B(n13623), .ZN(n13620) );
  NAND2_X1 U13609 ( .A1(n13621), .A2(n13624), .ZN(n7514) );
  XOR2_X1 U13610 ( .A(n13622), .B(n13623), .Z(n13624) );
  NOR2_X1 U13611 ( .A1(n13615), .A2(n13614), .ZN(n13621) );
  AND2_X1 U13612 ( .A1(n13625), .A2(n13626), .ZN(n13614) );
  NAND2_X1 U13613 ( .A1(n13619), .A2(n13627), .ZN(n13626) );
  OR2_X1 U13614 ( .A1(n13617), .A2(n13618), .ZN(n13627) );
  NOR2_X1 U13615 ( .A1(n8942), .A2(n7874), .ZN(n13619) );
  NAND2_X1 U13616 ( .A1(n13617), .A2(n13618), .ZN(n13625) );
  NAND2_X1 U13617 ( .A1(n13628), .A2(n13629), .ZN(n13618) );
  NAND2_X1 U13618 ( .A1(n13613), .A2(n13630), .ZN(n13629) );
  OR2_X1 U13619 ( .A1(n13611), .A2(n13612), .ZN(n13630) );
  NOR2_X1 U13620 ( .A1(n7874), .A2(n7957), .ZN(n13613) );
  NAND2_X1 U13621 ( .A1(n13611), .A2(n13612), .ZN(n13628) );
  NAND2_X1 U13622 ( .A1(n13631), .A2(n13632), .ZN(n13612) );
  NAND3_X1 U13623 ( .A1(b_7_), .A2(n13633), .A3(a_2_), .ZN(n13632) );
  OR2_X1 U13624 ( .A1(n13607), .A2(n13608), .ZN(n13633) );
  NAND2_X1 U13625 ( .A1(n13607), .A2(n13608), .ZN(n13631) );
  NAND2_X1 U13626 ( .A1(n13634), .A2(n13635), .ZN(n13608) );
  NAND3_X1 U13627 ( .A1(b_7_), .A2(n13636), .A3(a_3_), .ZN(n13635) );
  OR2_X1 U13628 ( .A1(n13603), .A2(n13604), .ZN(n13636) );
  NAND2_X1 U13629 ( .A1(n13603), .A2(n13604), .ZN(n13634) );
  NAND2_X1 U13630 ( .A1(n13637), .A2(n13638), .ZN(n13604) );
  NAND3_X1 U13631 ( .A1(b_7_), .A2(n13639), .A3(a_4_), .ZN(n13638) );
  OR2_X1 U13632 ( .A1(n13599), .A2(n13600), .ZN(n13639) );
  NAND2_X1 U13633 ( .A1(n13599), .A2(n13600), .ZN(n13637) );
  NAND2_X1 U13634 ( .A1(n13640), .A2(n13641), .ZN(n13600) );
  NAND3_X1 U13635 ( .A1(b_7_), .A2(n13642), .A3(a_5_), .ZN(n13641) );
  OR2_X1 U13636 ( .A1(n13595), .A2(n13596), .ZN(n13642) );
  NAND2_X1 U13637 ( .A1(n13595), .A2(n13596), .ZN(n13640) );
  NAND2_X1 U13638 ( .A1(n13643), .A2(n13644), .ZN(n13596) );
  NAND3_X1 U13639 ( .A1(b_7_), .A2(n13645), .A3(a_6_), .ZN(n13644) );
  OR2_X1 U13640 ( .A1(n13591), .A2(n13592), .ZN(n13645) );
  NAND2_X1 U13641 ( .A1(n13591), .A2(n13592), .ZN(n13643) );
  NAND2_X1 U13642 ( .A1(n13646), .A2(n13647), .ZN(n13592) );
  NAND2_X1 U13643 ( .A1(n13588), .A2(n13648), .ZN(n13647) );
  OR2_X1 U13644 ( .A1(n13589), .A2(n7869), .ZN(n13648) );
  XNOR2_X1 U13645 ( .A(n13649), .B(n13650), .ZN(n13588) );
  XOR2_X1 U13646 ( .A(n13651), .B(n13652), .Z(n13650) );
  NAND2_X1 U13647 ( .A1(b_6_), .A2(a_8_), .ZN(n13652) );
  NAND2_X1 U13648 ( .A1(n7869), .A2(n13589), .ZN(n13646) );
  NAND2_X1 U13649 ( .A1(n13653), .A2(n13654), .ZN(n13589) );
  NAND3_X1 U13650 ( .A1(a_8_), .A2(n13655), .A3(b_7_), .ZN(n13654) );
  OR2_X1 U13651 ( .A1(n13584), .A2(n13585), .ZN(n13655) );
  NAND2_X1 U13652 ( .A1(n13584), .A2(n13585), .ZN(n13653) );
  NAND2_X1 U13653 ( .A1(n13656), .A2(n13657), .ZN(n13585) );
  NAND3_X1 U13654 ( .A1(a_9_), .A2(n13658), .A3(b_7_), .ZN(n13657) );
  OR2_X1 U13655 ( .A1(n13427), .A2(n13428), .ZN(n13658) );
  NAND2_X1 U13656 ( .A1(n13427), .A2(n13428), .ZN(n13656) );
  NAND2_X1 U13657 ( .A1(n13659), .A2(n13660), .ZN(n13428) );
  NAND3_X1 U13658 ( .A1(a_10_), .A2(n13661), .A3(b_7_), .ZN(n13660) );
  OR2_X1 U13659 ( .A1(n13580), .A2(n13581), .ZN(n13661) );
  NAND2_X1 U13660 ( .A1(n13580), .A2(n13581), .ZN(n13659) );
  NAND2_X1 U13661 ( .A1(n13662), .A2(n13663), .ZN(n13581) );
  NAND3_X1 U13662 ( .A1(a_11_), .A2(n13664), .A3(b_7_), .ZN(n13663) );
  OR2_X1 U13663 ( .A1(n13576), .A2(n13577), .ZN(n13664) );
  NAND2_X1 U13664 ( .A1(n13576), .A2(n13577), .ZN(n13662) );
  NAND2_X1 U13665 ( .A1(n13665), .A2(n13666), .ZN(n13577) );
  NAND3_X1 U13666 ( .A1(a_12_), .A2(n13667), .A3(b_7_), .ZN(n13666) );
  OR2_X1 U13667 ( .A1(n13572), .A2(n13573), .ZN(n13667) );
  NAND2_X1 U13668 ( .A1(n13572), .A2(n13573), .ZN(n13665) );
  NAND2_X1 U13669 ( .A1(n13668), .A2(n13669), .ZN(n13573) );
  NAND3_X1 U13670 ( .A1(a_13_), .A2(n13670), .A3(b_7_), .ZN(n13669) );
  OR2_X1 U13671 ( .A1(n13569), .A2(n13567), .ZN(n13670) );
  NAND2_X1 U13672 ( .A1(n13567), .A2(n13569), .ZN(n13668) );
  NAND2_X1 U13673 ( .A1(n13671), .A2(n13672), .ZN(n13569) );
  NAND3_X1 U13674 ( .A1(a_14_), .A2(n13673), .A3(b_7_), .ZN(n13672) );
  OR2_X1 U13675 ( .A1(n13564), .A2(n13565), .ZN(n13673) );
  NAND2_X1 U13676 ( .A1(n13564), .A2(n13565), .ZN(n13671) );
  NAND2_X1 U13677 ( .A1(n13674), .A2(n13675), .ZN(n13565) );
  NAND3_X1 U13678 ( .A1(a_15_), .A2(n13676), .A3(b_7_), .ZN(n13675) );
  OR2_X1 U13679 ( .A1(n13561), .A2(n13559), .ZN(n13676) );
  NAND2_X1 U13680 ( .A1(n13559), .A2(n13561), .ZN(n13674) );
  NAND2_X1 U13681 ( .A1(n13677), .A2(n13678), .ZN(n13561) );
  NAND3_X1 U13682 ( .A1(a_16_), .A2(n13679), .A3(b_7_), .ZN(n13678) );
  OR2_X1 U13683 ( .A1(n13556), .A2(n13557), .ZN(n13679) );
  NAND2_X1 U13684 ( .A1(n13556), .A2(n13557), .ZN(n13677) );
  NAND2_X1 U13685 ( .A1(n13680), .A2(n13681), .ZN(n13557) );
  NAND3_X1 U13686 ( .A1(a_17_), .A2(n13682), .A3(b_7_), .ZN(n13681) );
  NAND2_X1 U13687 ( .A1(n13457), .A2(n13456), .ZN(n13682) );
  OR2_X1 U13688 ( .A1(n13456), .A2(n13457), .ZN(n13680) );
  AND2_X1 U13689 ( .A1(n13683), .A2(n13684), .ZN(n13457) );
  NAND3_X1 U13690 ( .A1(a_18_), .A2(n13685), .A3(b_7_), .ZN(n13684) );
  OR2_X1 U13691 ( .A1(n13463), .A2(n13465), .ZN(n13685) );
  NAND2_X1 U13692 ( .A1(n13463), .A2(n13465), .ZN(n13683) );
  NAND2_X1 U13693 ( .A1(n13686), .A2(n13687), .ZN(n13465) );
  NAND3_X1 U13694 ( .A1(a_19_), .A2(n13688), .A3(b_7_), .ZN(n13687) );
  OR2_X1 U13695 ( .A1(n13553), .A2(n13551), .ZN(n13688) );
  NAND2_X1 U13696 ( .A1(n13551), .A2(n13553), .ZN(n13686) );
  NAND2_X1 U13697 ( .A1(n13689), .A2(n13690), .ZN(n13553) );
  NAND3_X1 U13698 ( .A1(a_20_), .A2(n13691), .A3(b_7_), .ZN(n13690) );
  NAND2_X1 U13699 ( .A1(n13549), .A2(n13548), .ZN(n13691) );
  OR2_X1 U13700 ( .A1(n13548), .A2(n13549), .ZN(n13689) );
  AND2_X1 U13701 ( .A1(n13692), .A2(n13693), .ZN(n13549) );
  NAND3_X1 U13702 ( .A1(a_21_), .A2(n13694), .A3(b_7_), .ZN(n13693) );
  OR2_X1 U13703 ( .A1(n13544), .A2(n13545), .ZN(n13694) );
  NAND2_X1 U13704 ( .A1(n13544), .A2(n13545), .ZN(n13692) );
  NAND2_X1 U13705 ( .A1(n13541), .A2(n13695), .ZN(n13545) );
  NAND2_X1 U13706 ( .A1(n13540), .A2(n13542), .ZN(n13695) );
  NAND2_X1 U13707 ( .A1(n13696), .A2(n13697), .ZN(n13542) );
  NAND2_X1 U13708 ( .A1(b_7_), .A2(a_22_), .ZN(n13697) );
  INV_X1 U13709 ( .A(n13698), .ZN(n13696) );
  XOR2_X1 U13710 ( .A(n13699), .B(n13700), .Z(n13540) );
  XOR2_X1 U13711 ( .A(n13701), .B(n13702), .Z(n13699) );
  NOR2_X1 U13712 ( .A1(n8042), .A2(n8053), .ZN(n13702) );
  NAND2_X1 U13713 ( .A1(a_22_), .A2(n13698), .ZN(n13541) );
  NAND2_X1 U13714 ( .A1(n13703), .A2(n13704), .ZN(n13698) );
  NAND3_X1 U13715 ( .A1(a_23_), .A2(n13705), .A3(b_7_), .ZN(n13704) );
  OR2_X1 U13716 ( .A1(n13536), .A2(n13537), .ZN(n13705) );
  NAND2_X1 U13717 ( .A1(n13536), .A2(n13537), .ZN(n13703) );
  NAND2_X1 U13718 ( .A1(n13706), .A2(n13707), .ZN(n13537) );
  NAND2_X1 U13719 ( .A1(n13534), .A2(n13708), .ZN(n13707) );
  OR2_X1 U13720 ( .A1(n13532), .A2(n13533), .ZN(n13708) );
  NOR2_X1 U13721 ( .A1(n7874), .A2(n8041), .ZN(n13534) );
  NAND2_X1 U13722 ( .A1(n13532), .A2(n13533), .ZN(n13706) );
  NAND2_X1 U13723 ( .A1(n13709), .A2(n13710), .ZN(n13533) );
  NAND2_X1 U13724 ( .A1(n13530), .A2(n13711), .ZN(n13710) );
  OR2_X1 U13725 ( .A1(n13528), .A2(n13529), .ZN(n13711) );
  NOR2_X1 U13726 ( .A1(n7874), .A2(n8039), .ZN(n13530) );
  NAND2_X1 U13727 ( .A1(n13528), .A2(n13529), .ZN(n13709) );
  NAND2_X1 U13728 ( .A1(n13525), .A2(n13712), .ZN(n13529) );
  NAND2_X1 U13729 ( .A1(n13524), .A2(n13526), .ZN(n13712) );
  NAND2_X1 U13730 ( .A1(n13713), .A2(n13714), .ZN(n13526) );
  NAND2_X1 U13731 ( .A1(b_7_), .A2(a_26_), .ZN(n13714) );
  INV_X1 U13732 ( .A(n13715), .ZN(n13713) );
  XNOR2_X1 U13733 ( .A(n13716), .B(n13717), .ZN(n13524) );
  NAND2_X1 U13734 ( .A1(n13718), .A2(n13719), .ZN(n13716) );
  NAND2_X1 U13735 ( .A1(a_26_), .A2(n13715), .ZN(n13525) );
  NAND2_X1 U13736 ( .A1(n13497), .A2(n13720), .ZN(n13715) );
  NAND2_X1 U13737 ( .A1(n13496), .A2(n13498), .ZN(n13720) );
  NAND2_X1 U13738 ( .A1(n13721), .A2(n13722), .ZN(n13498) );
  NAND2_X1 U13739 ( .A1(b_7_), .A2(a_27_), .ZN(n13722) );
  INV_X1 U13740 ( .A(n13723), .ZN(n13721) );
  XNOR2_X1 U13741 ( .A(n13724), .B(n13725), .ZN(n13496) );
  XOR2_X1 U13742 ( .A(n13726), .B(n13727), .Z(n13724) );
  NAND2_X1 U13743 ( .A1(b_6_), .A2(a_28_), .ZN(n13726) );
  NAND2_X1 U13744 ( .A1(a_27_), .A2(n13723), .ZN(n13497) );
  NAND2_X1 U13745 ( .A1(n13728), .A2(n13729), .ZN(n13723) );
  NAND3_X1 U13746 ( .A1(a_28_), .A2(n13730), .A3(b_7_), .ZN(n13729) );
  NAND2_X1 U13747 ( .A1(n13506), .A2(n13504), .ZN(n13730) );
  OR2_X1 U13748 ( .A1(n13504), .A2(n13506), .ZN(n13728) );
  AND2_X1 U13749 ( .A1(n13731), .A2(n13732), .ZN(n13506) );
  NAND2_X1 U13750 ( .A1(n13520), .A2(n13733), .ZN(n13732) );
  OR2_X1 U13751 ( .A1(n13521), .A2(n13522), .ZN(n13733) );
  NOR2_X1 U13752 ( .A1(n7874), .A2(n7545), .ZN(n13520) );
  NAND2_X1 U13753 ( .A1(n13522), .A2(n13521), .ZN(n13731) );
  NAND2_X1 U13754 ( .A1(n13734), .A2(n13735), .ZN(n13521) );
  NAND2_X1 U13755 ( .A1(b_5_), .A2(n13736), .ZN(n13735) );
  NAND2_X1 U13756 ( .A1(n7527), .A2(n13737), .ZN(n13736) );
  NAND2_X1 U13757 ( .A1(a_31_), .A2(n8053), .ZN(n13737) );
  NAND2_X1 U13758 ( .A1(b_6_), .A2(n13738), .ZN(n13734) );
  NAND2_X1 U13759 ( .A1(n7531), .A2(n13739), .ZN(n13738) );
  NAND2_X1 U13760 ( .A1(a_30_), .A2(n7901), .ZN(n13739) );
  AND3_X1 U13761 ( .A1(b_6_), .A2(b_7_), .A3(n7494), .ZN(n13522) );
  XNOR2_X1 U13762 ( .A(n13740), .B(n13741), .ZN(n13504) );
  XOR2_X1 U13763 ( .A(n13742), .B(n13743), .Z(n13740) );
  XNOR2_X1 U13764 ( .A(n13744), .B(n13745), .ZN(n13528) );
  NAND2_X1 U13765 ( .A1(n13746), .A2(n13747), .ZN(n13744) );
  XNOR2_X1 U13766 ( .A(n13748), .B(n13749), .ZN(n13532) );
  NAND2_X1 U13767 ( .A1(n13750), .A2(n13751), .ZN(n13748) );
  XNOR2_X1 U13768 ( .A(n13752), .B(n13753), .ZN(n13536) );
  XNOR2_X1 U13769 ( .A(n13754), .B(n13755), .ZN(n13753) );
  XNOR2_X1 U13770 ( .A(n13756), .B(n13757), .ZN(n13544) );
  NAND2_X1 U13771 ( .A1(n13758), .A2(n13759), .ZN(n13756) );
  XOR2_X1 U13772 ( .A(n13760), .B(n13761), .Z(n13548) );
  XNOR2_X1 U13773 ( .A(n13762), .B(n13763), .ZN(n13761) );
  XOR2_X1 U13774 ( .A(n13764), .B(n13765), .Z(n13551) );
  XOR2_X1 U13775 ( .A(n13766), .B(n13767), .Z(n13764) );
  NOR2_X1 U13776 ( .A1(n8044), .A2(n8053), .ZN(n13767) );
  XNOR2_X1 U13777 ( .A(n13768), .B(n13769), .ZN(n13463) );
  XNOR2_X1 U13778 ( .A(n13770), .B(n13771), .ZN(n13768) );
  XNOR2_X1 U13779 ( .A(n13772), .B(n13773), .ZN(n13456) );
  XOR2_X1 U13780 ( .A(n13774), .B(n13775), .Z(n13772) );
  XNOR2_X1 U13781 ( .A(n13776), .B(n13777), .ZN(n13556) );
  XNOR2_X1 U13782 ( .A(n13778), .B(n13779), .ZN(n13776) );
  XNOR2_X1 U13783 ( .A(n13780), .B(n13781), .ZN(n13559) );
  XNOR2_X1 U13784 ( .A(n13782), .B(n13783), .ZN(n13781) );
  XNOR2_X1 U13785 ( .A(n13784), .B(n13785), .ZN(n13564) );
  XNOR2_X1 U13786 ( .A(n13786), .B(n13787), .ZN(n13784) );
  XOR2_X1 U13787 ( .A(n13788), .B(n13789), .Z(n13567) );
  XOR2_X1 U13788 ( .A(n13790), .B(n13791), .Z(n13788) );
  XNOR2_X1 U13789 ( .A(n13792), .B(n13793), .ZN(n13572) );
  XNOR2_X1 U13790 ( .A(n13794), .B(n13795), .ZN(n13792) );
  XNOR2_X1 U13791 ( .A(n13796), .B(n13797), .ZN(n13576) );
  XNOR2_X1 U13792 ( .A(n13798), .B(n13799), .ZN(n13796) );
  XNOR2_X1 U13793 ( .A(n13800), .B(n13801), .ZN(n13580) );
  XNOR2_X1 U13794 ( .A(n13802), .B(n13803), .ZN(n13801) );
  XNOR2_X1 U13795 ( .A(n13804), .B(n13805), .ZN(n13427) );
  XNOR2_X1 U13796 ( .A(n13806), .B(n13807), .ZN(n13804) );
  XNOR2_X1 U13797 ( .A(n13808), .B(n13809), .ZN(n13584) );
  XOR2_X1 U13798 ( .A(n13810), .B(n13811), .Z(n13809) );
  NAND2_X1 U13799 ( .A1(b_6_), .A2(a_9_), .ZN(n13811) );
  INV_X1 U13800 ( .A(n7987), .ZN(n7869) );
  NAND2_X1 U13801 ( .A1(a_7_), .A2(b_7_), .ZN(n7987) );
  XOR2_X1 U13802 ( .A(n13812), .B(n13813), .Z(n13591) );
  XOR2_X1 U13803 ( .A(n13814), .B(n13815), .Z(n13812) );
  NOR2_X1 U13804 ( .A1(n7872), .A2(n8053), .ZN(n13815) );
  XOR2_X1 U13805 ( .A(n13816), .B(n13817), .Z(n13595) );
  XOR2_X1 U13806 ( .A(n13818), .B(n13819), .Z(n13816) );
  XOR2_X1 U13807 ( .A(n13820), .B(n13821), .Z(n13599) );
  XOR2_X1 U13808 ( .A(n13822), .B(n13823), .Z(n13820) );
  NOR2_X1 U13809 ( .A1(n8053), .A2(n7908), .ZN(n13823) );
  XOR2_X1 U13810 ( .A(n13824), .B(n13825), .Z(n13603) );
  XNOR2_X1 U13811 ( .A(n13826), .B(n13827), .ZN(n13825) );
  NAND2_X1 U13812 ( .A1(a_4_), .A2(b_6_), .ZN(n13827) );
  XOR2_X1 U13813 ( .A(n13828), .B(n13829), .Z(n13607) );
  XOR2_X1 U13814 ( .A(n13830), .B(n13831), .Z(n13828) );
  NOR2_X1 U13815 ( .A1(n8053), .A2(n7937), .ZN(n13831) );
  XOR2_X1 U13816 ( .A(n13832), .B(n13833), .Z(n13611) );
  XOR2_X1 U13817 ( .A(n13834), .B(n13835), .Z(n13832) );
  NOR2_X1 U13818 ( .A1(n8053), .A2(n8056), .ZN(n13835) );
  XOR2_X1 U13819 ( .A(n13836), .B(n13837), .Z(n13617) );
  XOR2_X1 U13820 ( .A(n13838), .B(n13839), .Z(n13836) );
  NOR2_X1 U13821 ( .A1(n7957), .A2(n8053), .ZN(n13839) );
  XNOR2_X1 U13822 ( .A(n13840), .B(n13841), .ZN(n13615) );
  XOR2_X1 U13823 ( .A(n13842), .B(n13843), .Z(n13840) );
  NOR2_X1 U13824 ( .A1(n8053), .A2(n8942), .ZN(n13843) );
  NAND2_X1 U13825 ( .A1(n13844), .A2(n13845), .ZN(n7570) );
  NAND2_X1 U13826 ( .A1(n13846), .A2(n13847), .ZN(n13845) );
  NAND2_X1 U13827 ( .A1(n13623), .A2(n13622), .ZN(n13844) );
  NAND4_X1 U13828 ( .A1(n13623), .A2(n13846), .A3(n13622), .A4(n13847), .ZN(
        n7569) );
  NAND2_X1 U13829 ( .A1(n13848), .A2(n13849), .ZN(n13622) );
  NAND3_X1 U13830 ( .A1(b_6_), .A2(n13850), .A3(a_0_), .ZN(n13849) );
  OR2_X1 U13831 ( .A1(n13841), .A2(n13842), .ZN(n13850) );
  NAND2_X1 U13832 ( .A1(n13841), .A2(n13842), .ZN(n13848) );
  NAND2_X1 U13833 ( .A1(n13851), .A2(n13852), .ZN(n13842) );
  NAND3_X1 U13834 ( .A1(a_1_), .A2(n13853), .A3(b_6_), .ZN(n13852) );
  OR2_X1 U13835 ( .A1(n13838), .A2(n13837), .ZN(n13853) );
  NAND2_X1 U13836 ( .A1(n13837), .A2(n13838), .ZN(n13851) );
  NAND2_X1 U13837 ( .A1(n13854), .A2(n13855), .ZN(n13838) );
  NAND3_X1 U13838 ( .A1(b_6_), .A2(n13856), .A3(a_2_), .ZN(n13855) );
  OR2_X1 U13839 ( .A1(n13834), .A2(n13833), .ZN(n13856) );
  NAND2_X1 U13840 ( .A1(n13833), .A2(n13834), .ZN(n13854) );
  NAND2_X1 U13841 ( .A1(n13857), .A2(n13858), .ZN(n13834) );
  NAND3_X1 U13842 ( .A1(b_6_), .A2(n13859), .A3(a_3_), .ZN(n13858) );
  OR2_X1 U13843 ( .A1(n13830), .A2(n13829), .ZN(n13859) );
  NAND2_X1 U13844 ( .A1(n13829), .A2(n13830), .ZN(n13857) );
  NAND2_X1 U13845 ( .A1(n13860), .A2(n13861), .ZN(n13830) );
  NAND3_X1 U13846 ( .A1(b_6_), .A2(n13862), .A3(a_4_), .ZN(n13861) );
  NAND2_X1 U13847 ( .A1(n13826), .A2(n13824), .ZN(n13862) );
  OR2_X1 U13848 ( .A1(n13824), .A2(n13826), .ZN(n13860) );
  AND2_X1 U13849 ( .A1(n13863), .A2(n13864), .ZN(n13826) );
  NAND3_X1 U13850 ( .A1(b_6_), .A2(n13865), .A3(a_5_), .ZN(n13864) );
  OR2_X1 U13851 ( .A1(n13822), .A2(n13821), .ZN(n13865) );
  NAND2_X1 U13852 ( .A1(n13821), .A2(n13822), .ZN(n13863) );
  NAND2_X1 U13853 ( .A1(n13866), .A2(n13867), .ZN(n13822) );
  NAND2_X1 U13854 ( .A1(n13817), .A2(n13868), .ZN(n13867) );
  OR2_X1 U13855 ( .A1(n13818), .A2(n13819), .ZN(n13868) );
  XNOR2_X1 U13856 ( .A(n13869), .B(n13870), .ZN(n13817) );
  XNOR2_X1 U13857 ( .A(n13871), .B(n13872), .ZN(n13869) );
  NOR2_X1 U13858 ( .A1(n7872), .A2(n7901), .ZN(n13872) );
  NAND2_X1 U13859 ( .A1(n13819), .A2(n13818), .ZN(n13866) );
  NAND2_X1 U13860 ( .A1(n13873), .A2(n13874), .ZN(n13818) );
  NAND3_X1 U13861 ( .A1(a_7_), .A2(n13875), .A3(b_6_), .ZN(n13874) );
  OR2_X1 U13862 ( .A1(n13814), .A2(n13813), .ZN(n13875) );
  NAND2_X1 U13863 ( .A1(n13813), .A2(n13814), .ZN(n13873) );
  NAND2_X1 U13864 ( .A1(n13876), .A2(n13877), .ZN(n13814) );
  NAND3_X1 U13865 ( .A1(a_8_), .A2(n13878), .A3(b_6_), .ZN(n13877) );
  OR2_X1 U13866 ( .A1(n13651), .A2(n13649), .ZN(n13878) );
  NAND2_X1 U13867 ( .A1(n13649), .A2(n13651), .ZN(n13876) );
  NAND2_X1 U13868 ( .A1(n13879), .A2(n13880), .ZN(n13651) );
  NAND3_X1 U13869 ( .A1(a_9_), .A2(n13881), .A3(b_6_), .ZN(n13880) );
  OR2_X1 U13870 ( .A1(n13810), .A2(n13808), .ZN(n13881) );
  NAND2_X1 U13871 ( .A1(n13808), .A2(n13810), .ZN(n13879) );
  NAND2_X1 U13872 ( .A1(n13882), .A2(n13883), .ZN(n13810) );
  NAND2_X1 U13873 ( .A1(n13807), .A2(n13884), .ZN(n13883) );
  NAND2_X1 U13874 ( .A1(n13806), .A2(n13805), .ZN(n13884) );
  NOR2_X1 U13875 ( .A1(n8053), .A2(n8051), .ZN(n13807) );
  OR2_X1 U13876 ( .A1(n13805), .A2(n13806), .ZN(n13882) );
  AND2_X1 U13877 ( .A1(n13885), .A2(n13886), .ZN(n13806) );
  NAND2_X1 U13878 ( .A1(n13803), .A2(n13887), .ZN(n13886) );
  OR2_X1 U13879 ( .A1(n13802), .A2(n13800), .ZN(n13887) );
  NOR2_X1 U13880 ( .A1(n8053), .A2(n7811), .ZN(n13803) );
  NAND2_X1 U13881 ( .A1(n13800), .A2(n13802), .ZN(n13885) );
  NAND2_X1 U13882 ( .A1(n13888), .A2(n13889), .ZN(n13802) );
  NAND2_X1 U13883 ( .A1(n13799), .A2(n13890), .ZN(n13889) );
  NAND2_X1 U13884 ( .A1(n13798), .A2(n13797), .ZN(n13890) );
  NOR2_X1 U13885 ( .A1(n8053), .A2(n8669), .ZN(n13799) );
  OR2_X1 U13886 ( .A1(n13797), .A2(n13798), .ZN(n13888) );
  AND2_X1 U13887 ( .A1(n13891), .A2(n13892), .ZN(n13798) );
  NAND2_X1 U13888 ( .A1(n13795), .A2(n13893), .ZN(n13892) );
  NAND2_X1 U13889 ( .A1(n13794), .A2(n13793), .ZN(n13893) );
  NOR2_X1 U13890 ( .A1(n8053), .A2(n7789), .ZN(n13795) );
  OR2_X1 U13891 ( .A1(n13793), .A2(n13794), .ZN(n13891) );
  AND2_X1 U13892 ( .A1(n13894), .A2(n13895), .ZN(n13794) );
  NAND2_X1 U13893 ( .A1(n13791), .A2(n13896), .ZN(n13895) );
  OR2_X1 U13894 ( .A1(n13789), .A2(n13790), .ZN(n13896) );
  NOR2_X1 U13895 ( .A1(n8053), .A2(n8049), .ZN(n13791) );
  NAND2_X1 U13896 ( .A1(n13789), .A2(n13790), .ZN(n13894) );
  NAND2_X1 U13897 ( .A1(n13897), .A2(n13898), .ZN(n13790) );
  NAND2_X1 U13898 ( .A1(n13787), .A2(n13899), .ZN(n13898) );
  NAND2_X1 U13899 ( .A1(n13786), .A2(n13785), .ZN(n13899) );
  NOR2_X1 U13900 ( .A1(n8053), .A2(n7754), .ZN(n13787) );
  OR2_X1 U13901 ( .A1(n13785), .A2(n13786), .ZN(n13897) );
  AND2_X1 U13902 ( .A1(n13900), .A2(n13901), .ZN(n13786) );
  NAND2_X1 U13903 ( .A1(n13783), .A2(n13902), .ZN(n13901) );
  OR2_X1 U13904 ( .A1(n13780), .A2(n13782), .ZN(n13902) );
  NOR2_X1 U13905 ( .A1(n8053), .A2(n8438), .ZN(n13783) );
  NAND2_X1 U13906 ( .A1(n13780), .A2(n13782), .ZN(n13900) );
  NAND2_X1 U13907 ( .A1(n13903), .A2(n13904), .ZN(n13782) );
  NAND2_X1 U13908 ( .A1(n13779), .A2(n13905), .ZN(n13904) );
  NAND2_X1 U13909 ( .A1(n13778), .A2(n13777), .ZN(n13905) );
  NOR2_X1 U13910 ( .A1(n8053), .A2(n7732), .ZN(n13779) );
  OR2_X1 U13911 ( .A1(n13777), .A2(n13778), .ZN(n13903) );
  AND2_X1 U13912 ( .A1(n13906), .A2(n13907), .ZN(n13778) );
  NAND2_X1 U13913 ( .A1(n13774), .A2(n13908), .ZN(n13907) );
  OR2_X1 U13914 ( .A1(n13773), .A2(n13775), .ZN(n13908) );
  NOR2_X1 U13915 ( .A1(n8053), .A2(n8047), .ZN(n13774) );
  NAND2_X1 U13916 ( .A1(n13773), .A2(n13775), .ZN(n13906) );
  NAND2_X1 U13917 ( .A1(n13909), .A2(n13910), .ZN(n13775) );
  NAND2_X1 U13918 ( .A1(n13771), .A2(n13911), .ZN(n13910) );
  NAND2_X1 U13919 ( .A1(n13770), .A2(n13769), .ZN(n13911) );
  NOR2_X1 U13920 ( .A1(n8053), .A2(n8045), .ZN(n13771) );
  OR2_X1 U13921 ( .A1(n13769), .A2(n13770), .ZN(n13909) );
  AND2_X1 U13922 ( .A1(n13912), .A2(n13913), .ZN(n13770) );
  NAND3_X1 U13923 ( .A1(a_20_), .A2(n13914), .A3(b_6_), .ZN(n13913) );
  OR2_X1 U13924 ( .A1(n13765), .A2(n13766), .ZN(n13914) );
  NAND2_X1 U13925 ( .A1(n13765), .A2(n13766), .ZN(n13912) );
  NAND2_X1 U13926 ( .A1(n13915), .A2(n13916), .ZN(n13766) );
  NAND2_X1 U13927 ( .A1(n13763), .A2(n13917), .ZN(n13916) );
  OR2_X1 U13928 ( .A1(n13760), .A2(n13762), .ZN(n13917) );
  NOR2_X1 U13929 ( .A1(n8053), .A2(n7665), .ZN(n13763) );
  NAND2_X1 U13930 ( .A1(n13760), .A2(n13762), .ZN(n13915) );
  NAND2_X1 U13931 ( .A1(n13758), .A2(n13918), .ZN(n13762) );
  NAND2_X1 U13932 ( .A1(n13757), .A2(n13759), .ZN(n13918) );
  NAND2_X1 U13933 ( .A1(n13919), .A2(n13920), .ZN(n13759) );
  NAND2_X1 U13934 ( .A1(b_6_), .A2(a_22_), .ZN(n13920) );
  INV_X1 U13935 ( .A(n13921), .ZN(n13919) );
  XNOR2_X1 U13936 ( .A(n13922), .B(n13923), .ZN(n13757) );
  XOR2_X1 U13937 ( .A(n13924), .B(n13925), .Z(n13923) );
  NAND2_X1 U13938 ( .A1(b_5_), .A2(a_23_), .ZN(n13925) );
  NAND2_X1 U13939 ( .A1(a_22_), .A2(n13921), .ZN(n13758) );
  NAND2_X1 U13940 ( .A1(n13926), .A2(n13927), .ZN(n13921) );
  NAND3_X1 U13941 ( .A1(a_23_), .A2(n13928), .A3(b_6_), .ZN(n13927) );
  OR2_X1 U13942 ( .A1(n13700), .A2(n13701), .ZN(n13928) );
  NAND2_X1 U13943 ( .A1(n13700), .A2(n13701), .ZN(n13926) );
  NAND2_X1 U13944 ( .A1(n13929), .A2(n13930), .ZN(n13701) );
  NAND2_X1 U13945 ( .A1(n13755), .A2(n13931), .ZN(n13930) );
  OR2_X1 U13946 ( .A1(n13754), .A2(n13752), .ZN(n13931) );
  NOR2_X1 U13947 ( .A1(n8053), .A2(n8041), .ZN(n13755) );
  NAND2_X1 U13948 ( .A1(n13752), .A2(n13754), .ZN(n13929) );
  NAND2_X1 U13949 ( .A1(n13750), .A2(n13932), .ZN(n13754) );
  NAND2_X1 U13950 ( .A1(n13749), .A2(n13751), .ZN(n13932) );
  NAND2_X1 U13951 ( .A1(n13933), .A2(n13934), .ZN(n13751) );
  NAND2_X1 U13952 ( .A1(b_6_), .A2(a_25_), .ZN(n13934) );
  INV_X1 U13953 ( .A(n13935), .ZN(n13933) );
  XNOR2_X1 U13954 ( .A(n13936), .B(n13937), .ZN(n13749) );
  NAND2_X1 U13955 ( .A1(n13938), .A2(n13939), .ZN(n13936) );
  NAND2_X1 U13956 ( .A1(a_25_), .A2(n13935), .ZN(n13750) );
  NAND2_X1 U13957 ( .A1(n13746), .A2(n13940), .ZN(n13935) );
  NAND2_X1 U13958 ( .A1(n13745), .A2(n13747), .ZN(n13940) );
  NAND2_X1 U13959 ( .A1(n13941), .A2(n13942), .ZN(n13747) );
  NAND2_X1 U13960 ( .A1(b_6_), .A2(a_26_), .ZN(n13942) );
  INV_X1 U13961 ( .A(n13943), .ZN(n13941) );
  XNOR2_X1 U13962 ( .A(n13944), .B(n13945), .ZN(n13745) );
  NAND2_X1 U13963 ( .A1(n13946), .A2(n13947), .ZN(n13944) );
  NAND2_X1 U13964 ( .A1(a_26_), .A2(n13943), .ZN(n13746) );
  NAND2_X1 U13965 ( .A1(n13718), .A2(n13948), .ZN(n13943) );
  NAND2_X1 U13966 ( .A1(n13717), .A2(n13719), .ZN(n13948) );
  NAND2_X1 U13967 ( .A1(n13949), .A2(n13950), .ZN(n13719) );
  NAND2_X1 U13968 ( .A1(b_6_), .A2(a_27_), .ZN(n13950) );
  INV_X1 U13969 ( .A(n13951), .ZN(n13949) );
  XNOR2_X1 U13970 ( .A(n13952), .B(n13953), .ZN(n13717) );
  XOR2_X1 U13971 ( .A(n13954), .B(n13955), .Z(n13952) );
  NAND2_X1 U13972 ( .A1(b_5_), .A2(a_28_), .ZN(n13954) );
  NAND2_X1 U13973 ( .A1(a_27_), .A2(n13951), .ZN(n13718) );
  NAND2_X1 U13974 ( .A1(n13956), .A2(n13957), .ZN(n13951) );
  NAND3_X1 U13975 ( .A1(a_28_), .A2(n13958), .A3(b_6_), .ZN(n13957) );
  NAND2_X1 U13976 ( .A1(n13727), .A2(n13725), .ZN(n13958) );
  OR2_X1 U13977 ( .A1(n13725), .A2(n13727), .ZN(n13956) );
  AND2_X1 U13978 ( .A1(n13959), .A2(n13960), .ZN(n13727) );
  NAND2_X1 U13979 ( .A1(n13741), .A2(n13961), .ZN(n13960) );
  OR2_X1 U13980 ( .A1(n13742), .A2(n13743), .ZN(n13961) );
  NOR2_X1 U13981 ( .A1(n8053), .A2(n7545), .ZN(n13741) );
  NAND2_X1 U13982 ( .A1(n13743), .A2(n13742), .ZN(n13959) );
  NAND2_X1 U13983 ( .A1(n13962), .A2(n13963), .ZN(n13742) );
  NAND2_X1 U13984 ( .A1(b_4_), .A2(n13964), .ZN(n13963) );
  NAND2_X1 U13985 ( .A1(n7527), .A2(n13965), .ZN(n13964) );
  NAND2_X1 U13986 ( .A1(a_31_), .A2(n7901), .ZN(n13965) );
  NAND2_X1 U13987 ( .A1(b_5_), .A2(n13966), .ZN(n13962) );
  NAND2_X1 U13988 ( .A1(n7531), .A2(n13967), .ZN(n13966) );
  NAND2_X1 U13989 ( .A1(a_30_), .A2(n8054), .ZN(n13967) );
  AND3_X1 U13990 ( .A1(b_6_), .A2(b_5_), .A3(n7494), .ZN(n13743) );
  XNOR2_X1 U13991 ( .A(n13968), .B(n13969), .ZN(n13725) );
  XOR2_X1 U13992 ( .A(n13970), .B(n13971), .Z(n13968) );
  XNOR2_X1 U13993 ( .A(n13972), .B(n13973), .ZN(n13752) );
  NAND2_X1 U13994 ( .A1(n13974), .A2(n13975), .ZN(n13972) );
  XNOR2_X1 U13995 ( .A(n13976), .B(n13977), .ZN(n13700) );
  XOR2_X1 U13996 ( .A(n13978), .B(n13979), .Z(n13977) );
  NAND2_X1 U13997 ( .A1(b_5_), .A2(a_24_), .ZN(n13979) );
  XNOR2_X1 U13998 ( .A(n13980), .B(n13981), .ZN(n13760) );
  XOR2_X1 U13999 ( .A(n13982), .B(n13983), .Z(n13981) );
  NAND2_X1 U14000 ( .A1(b_5_), .A2(a_22_), .ZN(n13983) );
  XNOR2_X1 U14001 ( .A(n13984), .B(n13985), .ZN(n13765) );
  XNOR2_X1 U14002 ( .A(n13986), .B(n13987), .ZN(n13984) );
  NOR2_X1 U14003 ( .A1(n7665), .A2(n7901), .ZN(n13987) );
  XNOR2_X1 U14004 ( .A(n13988), .B(n13989), .ZN(n13769) );
  XOR2_X1 U14005 ( .A(n13990), .B(n13991), .Z(n13988) );
  NOR2_X1 U14006 ( .A1(n8044), .A2(n7901), .ZN(n13991) );
  XNOR2_X1 U14007 ( .A(n13992), .B(n13993), .ZN(n13773) );
  XOR2_X1 U14008 ( .A(n13994), .B(n13995), .Z(n13993) );
  NAND2_X1 U14009 ( .A1(b_5_), .A2(a_19_), .ZN(n13995) );
  XNOR2_X1 U14010 ( .A(n13996), .B(n13997), .ZN(n13777) );
  XOR2_X1 U14011 ( .A(n13998), .B(n13999), .Z(n13996) );
  NOR2_X1 U14012 ( .A1(n8047), .A2(n7901), .ZN(n13999) );
  XNOR2_X1 U14013 ( .A(n14000), .B(n14001), .ZN(n13780) );
  XNOR2_X1 U14014 ( .A(n14002), .B(n14003), .ZN(n14000) );
  NOR2_X1 U14015 ( .A1(n7732), .A2(n7901), .ZN(n14003) );
  XNOR2_X1 U14016 ( .A(n14004), .B(n14005), .ZN(n13785) );
  XOR2_X1 U14017 ( .A(n14006), .B(n14007), .Z(n14004) );
  NOR2_X1 U14018 ( .A1(n8438), .A2(n7901), .ZN(n14007) );
  XNOR2_X1 U14019 ( .A(n14008), .B(n14009), .ZN(n13789) );
  XNOR2_X1 U14020 ( .A(n14010), .B(n14011), .ZN(n14008) );
  NOR2_X1 U14021 ( .A1(n7754), .A2(n7901), .ZN(n14011) );
  XNOR2_X1 U14022 ( .A(n14012), .B(n14013), .ZN(n13793) );
  XOR2_X1 U14023 ( .A(n14014), .B(n14015), .Z(n14012) );
  NOR2_X1 U14024 ( .A1(n8049), .A2(n7901), .ZN(n14015) );
  XNOR2_X1 U14025 ( .A(n14016), .B(n14017), .ZN(n13797) );
  XOR2_X1 U14026 ( .A(n14018), .B(n14019), .Z(n14016) );
  NOR2_X1 U14027 ( .A1(n7789), .A2(n7901), .ZN(n14019) );
  XOR2_X1 U14028 ( .A(n14020), .B(n14021), .Z(n13800) );
  XOR2_X1 U14029 ( .A(n14022), .B(n14023), .Z(n14020) );
  NOR2_X1 U14030 ( .A1(n8669), .A2(n7901), .ZN(n14023) );
  XNOR2_X1 U14031 ( .A(n14024), .B(n14025), .ZN(n13805) );
  XOR2_X1 U14032 ( .A(n14026), .B(n14027), .Z(n14024) );
  NOR2_X1 U14033 ( .A1(n7811), .A2(n7901), .ZN(n14027) );
  XOR2_X1 U14034 ( .A(n14028), .B(n14029), .Z(n13808) );
  XOR2_X1 U14035 ( .A(n14030), .B(n14031), .Z(n14028) );
  NOR2_X1 U14036 ( .A1(n8051), .A2(n7901), .ZN(n14031) );
  XNOR2_X1 U14037 ( .A(n14032), .B(n14033), .ZN(n13649) );
  XNOR2_X1 U14038 ( .A(n14034), .B(n14035), .ZN(n14032) );
  NOR2_X1 U14039 ( .A1(n8052), .A2(n7901), .ZN(n14035) );
  XOR2_X1 U14040 ( .A(n14036), .B(n14037), .Z(n13813) );
  XOR2_X1 U14041 ( .A(n14038), .B(n14039), .Z(n14036) );
  NOR2_X1 U14042 ( .A1(n8686), .A2(n7901), .ZN(n14039) );
  INV_X1 U14043 ( .A(n7892), .ZN(n13819) );
  NAND2_X1 U14044 ( .A1(b_6_), .A2(a_6_), .ZN(n7892) );
  XOR2_X1 U14045 ( .A(n14040), .B(n14041), .Z(n13821) );
  XOR2_X1 U14046 ( .A(n14042), .B(n14043), .Z(n14040) );
  NOR2_X1 U14047 ( .A1(n7887), .A2(n7901), .ZN(n14043) );
  XNOR2_X1 U14048 ( .A(n14044), .B(n14045), .ZN(n13824) );
  XOR2_X1 U14049 ( .A(n14046), .B(n7899), .Z(n14044) );
  XOR2_X1 U14050 ( .A(n14047), .B(n14048), .Z(n13829) );
  XOR2_X1 U14051 ( .A(n14049), .B(n14050), .Z(n14047) );
  NOR2_X1 U14052 ( .A1(n7901), .A2(n7916), .ZN(n14050) );
  XOR2_X1 U14053 ( .A(n14051), .B(n14052), .Z(n13833) );
  XOR2_X1 U14054 ( .A(n14053), .B(n14054), .Z(n14051) );
  NOR2_X1 U14055 ( .A1(n7901), .A2(n7937), .ZN(n14054) );
  XOR2_X1 U14056 ( .A(n14055), .B(n14056), .Z(n13837) );
  XOR2_X1 U14057 ( .A(n14057), .B(n14058), .Z(n14055) );
  NOR2_X1 U14058 ( .A1(n7901), .A2(n8056), .ZN(n14058) );
  XOR2_X1 U14059 ( .A(n14059), .B(n14060), .Z(n13841) );
  XOR2_X1 U14060 ( .A(n14061), .B(n14062), .Z(n14059) );
  NAND2_X1 U14061 ( .A1(n14063), .A2(n14064), .ZN(n13846) );
  XOR2_X1 U14062 ( .A(n14065), .B(n14066), .Z(n13623) );
  XOR2_X1 U14063 ( .A(n14067), .B(n14068), .Z(n14065) );
  NAND2_X1 U14064 ( .A1(n14069), .A2(n13847), .ZN(n7716) );
  INV_X1 U14065 ( .A(n14070), .ZN(n13847) );
  XNOR2_X1 U14066 ( .A(n14071), .B(n14072), .ZN(n14069) );
  NAND2_X1 U14067 ( .A1(n14070), .A2(n14073), .ZN(n7715) );
  XOR2_X1 U14068 ( .A(n14071), .B(n14072), .Z(n14073) );
  NOR2_X1 U14069 ( .A1(n14064), .A2(n14063), .ZN(n14070) );
  AND2_X1 U14070 ( .A1(n14074), .A2(n14075), .ZN(n14063) );
  NAND2_X1 U14071 ( .A1(n14068), .A2(n14076), .ZN(n14075) );
  OR2_X1 U14072 ( .A1(n14066), .A2(n14067), .ZN(n14076) );
  NOR2_X1 U14073 ( .A1(n8942), .A2(n7901), .ZN(n14068) );
  NAND2_X1 U14074 ( .A1(n14066), .A2(n14067), .ZN(n14074) );
  NAND2_X1 U14075 ( .A1(n14077), .A2(n14078), .ZN(n14067) );
  NAND2_X1 U14076 ( .A1(n14062), .A2(n14079), .ZN(n14078) );
  OR2_X1 U14077 ( .A1(n14061), .A2(n14060), .ZN(n14079) );
  NOR2_X1 U14078 ( .A1(n7901), .A2(n7957), .ZN(n14062) );
  NAND2_X1 U14079 ( .A1(n14060), .A2(n14061), .ZN(n14077) );
  NAND2_X1 U14080 ( .A1(n14080), .A2(n14081), .ZN(n14061) );
  NAND3_X1 U14081 ( .A1(b_5_), .A2(n14082), .A3(a_2_), .ZN(n14081) );
  OR2_X1 U14082 ( .A1(n14056), .A2(n14057), .ZN(n14082) );
  NAND2_X1 U14083 ( .A1(n14056), .A2(n14057), .ZN(n14080) );
  NAND2_X1 U14084 ( .A1(n14083), .A2(n14084), .ZN(n14057) );
  NAND3_X1 U14085 ( .A1(b_5_), .A2(n14085), .A3(a_3_), .ZN(n14084) );
  OR2_X1 U14086 ( .A1(n14052), .A2(n14053), .ZN(n14085) );
  NAND2_X1 U14087 ( .A1(n14052), .A2(n14053), .ZN(n14083) );
  NAND2_X1 U14088 ( .A1(n14086), .A2(n14087), .ZN(n14053) );
  NAND3_X1 U14089 ( .A1(b_5_), .A2(n14088), .A3(a_4_), .ZN(n14087) );
  OR2_X1 U14090 ( .A1(n14048), .A2(n14049), .ZN(n14088) );
  NAND2_X1 U14091 ( .A1(n14048), .A2(n14049), .ZN(n14086) );
  NAND2_X1 U14092 ( .A1(n14089), .A2(n14090), .ZN(n14049) );
  NAND2_X1 U14093 ( .A1(n14045), .A2(n14091), .ZN(n14090) );
  OR2_X1 U14094 ( .A1(n14046), .A2(n7899), .ZN(n14091) );
  XNOR2_X1 U14095 ( .A(n14092), .B(n14093), .ZN(n14045) );
  XNOR2_X1 U14096 ( .A(n14094), .B(n14095), .ZN(n14092) );
  NOR2_X1 U14097 ( .A1(n7887), .A2(n8054), .ZN(n14095) );
  NAND2_X1 U14098 ( .A1(n7899), .A2(n14046), .ZN(n14089) );
  NAND2_X1 U14099 ( .A1(n14096), .A2(n14097), .ZN(n14046) );
  NAND3_X1 U14100 ( .A1(a_6_), .A2(n14098), .A3(b_5_), .ZN(n14097) );
  OR2_X1 U14101 ( .A1(n14041), .A2(n14042), .ZN(n14098) );
  NAND2_X1 U14102 ( .A1(n14041), .A2(n14042), .ZN(n14096) );
  NAND2_X1 U14103 ( .A1(n14099), .A2(n14100), .ZN(n14042) );
  NAND3_X1 U14104 ( .A1(a_7_), .A2(n14101), .A3(b_5_), .ZN(n14100) );
  NAND2_X1 U14105 ( .A1(n13870), .A2(n13871), .ZN(n14101) );
  OR2_X1 U14106 ( .A1(n13870), .A2(n13871), .ZN(n14099) );
  AND2_X1 U14107 ( .A1(n14102), .A2(n14103), .ZN(n13871) );
  NAND3_X1 U14108 ( .A1(a_8_), .A2(n14104), .A3(b_5_), .ZN(n14103) );
  OR2_X1 U14109 ( .A1(n14037), .A2(n14038), .ZN(n14104) );
  NAND2_X1 U14110 ( .A1(n14037), .A2(n14038), .ZN(n14102) );
  NAND2_X1 U14111 ( .A1(n14105), .A2(n14106), .ZN(n14038) );
  NAND3_X1 U14112 ( .A1(a_9_), .A2(n14107), .A3(b_5_), .ZN(n14106) );
  NAND2_X1 U14113 ( .A1(n14033), .A2(n14034), .ZN(n14107) );
  OR2_X1 U14114 ( .A1(n14033), .A2(n14034), .ZN(n14105) );
  AND2_X1 U14115 ( .A1(n14108), .A2(n14109), .ZN(n14034) );
  NAND3_X1 U14116 ( .A1(a_10_), .A2(n14110), .A3(b_5_), .ZN(n14109) );
  OR2_X1 U14117 ( .A1(n14029), .A2(n14030), .ZN(n14110) );
  NAND2_X1 U14118 ( .A1(n14029), .A2(n14030), .ZN(n14108) );
  NAND2_X1 U14119 ( .A1(n14111), .A2(n14112), .ZN(n14030) );
  NAND3_X1 U14120 ( .A1(a_11_), .A2(n14113), .A3(b_5_), .ZN(n14112) );
  OR2_X1 U14121 ( .A1(n14025), .A2(n14026), .ZN(n14113) );
  NAND2_X1 U14122 ( .A1(n14025), .A2(n14026), .ZN(n14111) );
  NAND2_X1 U14123 ( .A1(n14114), .A2(n14115), .ZN(n14026) );
  NAND3_X1 U14124 ( .A1(a_12_), .A2(n14116), .A3(b_5_), .ZN(n14115) );
  OR2_X1 U14125 ( .A1(n14021), .A2(n14022), .ZN(n14116) );
  NAND2_X1 U14126 ( .A1(n14021), .A2(n14022), .ZN(n14114) );
  NAND2_X1 U14127 ( .A1(n14117), .A2(n14118), .ZN(n14022) );
  NAND3_X1 U14128 ( .A1(a_13_), .A2(n14119), .A3(b_5_), .ZN(n14118) );
  OR2_X1 U14129 ( .A1(n14017), .A2(n14018), .ZN(n14119) );
  NAND2_X1 U14130 ( .A1(n14017), .A2(n14018), .ZN(n14117) );
  NAND2_X1 U14131 ( .A1(n14120), .A2(n14121), .ZN(n14018) );
  NAND3_X1 U14132 ( .A1(a_14_), .A2(n14122), .A3(b_5_), .ZN(n14121) );
  OR2_X1 U14133 ( .A1(n14013), .A2(n14014), .ZN(n14122) );
  NAND2_X1 U14134 ( .A1(n14013), .A2(n14014), .ZN(n14120) );
  NAND2_X1 U14135 ( .A1(n14123), .A2(n14124), .ZN(n14014) );
  NAND3_X1 U14136 ( .A1(a_15_), .A2(n14125), .A3(b_5_), .ZN(n14124) );
  NAND2_X1 U14137 ( .A1(n14010), .A2(n14009), .ZN(n14125) );
  OR2_X1 U14138 ( .A1(n14009), .A2(n14010), .ZN(n14123) );
  AND2_X1 U14139 ( .A1(n14126), .A2(n14127), .ZN(n14010) );
  NAND3_X1 U14140 ( .A1(a_16_), .A2(n14128), .A3(b_5_), .ZN(n14127) );
  OR2_X1 U14141 ( .A1(n14005), .A2(n14006), .ZN(n14128) );
  NAND2_X1 U14142 ( .A1(n14005), .A2(n14006), .ZN(n14126) );
  NAND2_X1 U14143 ( .A1(n14129), .A2(n14130), .ZN(n14006) );
  NAND3_X1 U14144 ( .A1(a_17_), .A2(n14131), .A3(b_5_), .ZN(n14130) );
  NAND2_X1 U14145 ( .A1(n14002), .A2(n14001), .ZN(n14131) );
  OR2_X1 U14146 ( .A1(n14001), .A2(n14002), .ZN(n14129) );
  AND2_X1 U14147 ( .A1(n14132), .A2(n14133), .ZN(n14002) );
  NAND3_X1 U14148 ( .A1(a_18_), .A2(n14134), .A3(b_5_), .ZN(n14133) );
  OR2_X1 U14149 ( .A1(n13997), .A2(n13998), .ZN(n14134) );
  NAND2_X1 U14150 ( .A1(n13997), .A2(n13998), .ZN(n14132) );
  NAND2_X1 U14151 ( .A1(n14135), .A2(n14136), .ZN(n13998) );
  NAND3_X1 U14152 ( .A1(a_19_), .A2(n14137), .A3(b_5_), .ZN(n14136) );
  OR2_X1 U14153 ( .A1(n13994), .A2(n13992), .ZN(n14137) );
  NAND2_X1 U14154 ( .A1(n13992), .A2(n13994), .ZN(n14135) );
  NAND2_X1 U14155 ( .A1(n14138), .A2(n14139), .ZN(n13994) );
  NAND3_X1 U14156 ( .A1(a_20_), .A2(n14140), .A3(b_5_), .ZN(n14139) );
  OR2_X1 U14157 ( .A1(n13989), .A2(n13990), .ZN(n14140) );
  NAND2_X1 U14158 ( .A1(n13989), .A2(n13990), .ZN(n14138) );
  NAND2_X1 U14159 ( .A1(n14141), .A2(n14142), .ZN(n13990) );
  NAND3_X1 U14160 ( .A1(a_21_), .A2(n14143), .A3(b_5_), .ZN(n14142) );
  NAND2_X1 U14161 ( .A1(n13986), .A2(n13985), .ZN(n14143) );
  OR2_X1 U14162 ( .A1(n13985), .A2(n13986), .ZN(n14141) );
  AND2_X1 U14163 ( .A1(n14144), .A2(n14145), .ZN(n13986) );
  NAND3_X1 U14164 ( .A1(a_22_), .A2(n14146), .A3(b_5_), .ZN(n14145) );
  OR2_X1 U14165 ( .A1(n13982), .A2(n13980), .ZN(n14146) );
  NAND2_X1 U14166 ( .A1(n13980), .A2(n13982), .ZN(n14144) );
  NAND2_X1 U14167 ( .A1(n14147), .A2(n14148), .ZN(n13982) );
  NAND3_X1 U14168 ( .A1(a_23_), .A2(n14149), .A3(b_5_), .ZN(n14148) );
  OR2_X1 U14169 ( .A1(n13924), .A2(n13922), .ZN(n14149) );
  NAND2_X1 U14170 ( .A1(n13922), .A2(n13924), .ZN(n14147) );
  NAND2_X1 U14171 ( .A1(n14150), .A2(n14151), .ZN(n13924) );
  NAND3_X1 U14172 ( .A1(a_24_), .A2(n14152), .A3(b_5_), .ZN(n14151) );
  OR2_X1 U14173 ( .A1(n13978), .A2(n13976), .ZN(n14152) );
  NAND2_X1 U14174 ( .A1(n13976), .A2(n13978), .ZN(n14150) );
  NAND2_X1 U14175 ( .A1(n13974), .A2(n14153), .ZN(n13978) );
  NAND2_X1 U14176 ( .A1(n13973), .A2(n13975), .ZN(n14153) );
  NAND2_X1 U14177 ( .A1(n14154), .A2(n14155), .ZN(n13975) );
  NAND2_X1 U14178 ( .A1(b_5_), .A2(a_25_), .ZN(n14155) );
  INV_X1 U14179 ( .A(n14156), .ZN(n14154) );
  XNOR2_X1 U14180 ( .A(n14157), .B(n14158), .ZN(n13973) );
  NAND2_X1 U14181 ( .A1(n14159), .A2(n14160), .ZN(n14157) );
  NAND2_X1 U14182 ( .A1(a_25_), .A2(n14156), .ZN(n13974) );
  NAND2_X1 U14183 ( .A1(n13938), .A2(n14161), .ZN(n14156) );
  NAND2_X1 U14184 ( .A1(n13937), .A2(n13939), .ZN(n14161) );
  NAND2_X1 U14185 ( .A1(n14162), .A2(n14163), .ZN(n13939) );
  NAND2_X1 U14186 ( .A1(b_5_), .A2(a_26_), .ZN(n14163) );
  INV_X1 U14187 ( .A(n14164), .ZN(n14162) );
  XNOR2_X1 U14188 ( .A(n14165), .B(n14166), .ZN(n13937) );
  NAND2_X1 U14189 ( .A1(n14167), .A2(n14168), .ZN(n14165) );
  NAND2_X1 U14190 ( .A1(a_26_), .A2(n14164), .ZN(n13938) );
  NAND2_X1 U14191 ( .A1(n13946), .A2(n14169), .ZN(n14164) );
  NAND2_X1 U14192 ( .A1(n13945), .A2(n13947), .ZN(n14169) );
  NAND2_X1 U14193 ( .A1(n14170), .A2(n14171), .ZN(n13947) );
  NAND2_X1 U14194 ( .A1(b_5_), .A2(a_27_), .ZN(n14171) );
  INV_X1 U14195 ( .A(n14172), .ZN(n14170) );
  XNOR2_X1 U14196 ( .A(n14173), .B(n14174), .ZN(n13945) );
  XOR2_X1 U14197 ( .A(n14175), .B(n14176), .Z(n14173) );
  NAND2_X1 U14198 ( .A1(b_4_), .A2(a_28_), .ZN(n14175) );
  NAND2_X1 U14199 ( .A1(a_27_), .A2(n14172), .ZN(n13946) );
  NAND2_X1 U14200 ( .A1(n14177), .A2(n14178), .ZN(n14172) );
  NAND3_X1 U14201 ( .A1(a_28_), .A2(n14179), .A3(b_5_), .ZN(n14178) );
  NAND2_X1 U14202 ( .A1(n13955), .A2(n13953), .ZN(n14179) );
  OR2_X1 U14203 ( .A1(n13953), .A2(n13955), .ZN(n14177) );
  AND2_X1 U14204 ( .A1(n14180), .A2(n14181), .ZN(n13955) );
  NAND2_X1 U14205 ( .A1(n13969), .A2(n14182), .ZN(n14181) );
  OR2_X1 U14206 ( .A1(n13970), .A2(n13971), .ZN(n14182) );
  NOR2_X1 U14207 ( .A1(n7901), .A2(n7545), .ZN(n13969) );
  NAND2_X1 U14208 ( .A1(n13971), .A2(n13970), .ZN(n14180) );
  NAND2_X1 U14209 ( .A1(n14183), .A2(n14184), .ZN(n13970) );
  NAND2_X1 U14210 ( .A1(b_3_), .A2(n14185), .ZN(n14184) );
  NAND2_X1 U14211 ( .A1(n7527), .A2(n14186), .ZN(n14185) );
  NAND2_X1 U14212 ( .A1(a_31_), .A2(n8054), .ZN(n14186) );
  NAND2_X1 U14213 ( .A1(b_4_), .A2(n14187), .ZN(n14183) );
  NAND2_X1 U14214 ( .A1(n7531), .A2(n14188), .ZN(n14187) );
  NAND2_X1 U14215 ( .A1(a_30_), .A2(n7930), .ZN(n14188) );
  AND3_X1 U14216 ( .A1(b_4_), .A2(b_5_), .A3(n7494), .ZN(n13971) );
  XNOR2_X1 U14217 ( .A(n14189), .B(n14190), .ZN(n13953) );
  XOR2_X1 U14218 ( .A(n14191), .B(n14192), .Z(n14189) );
  XOR2_X1 U14219 ( .A(n14193), .B(n14194), .Z(n13976) );
  XOR2_X1 U14220 ( .A(n14195), .B(n14196), .Z(n14193) );
  XOR2_X1 U14221 ( .A(n14197), .B(n14198), .Z(n13922) );
  XOR2_X1 U14222 ( .A(n14199), .B(n14200), .Z(n14197) );
  XOR2_X1 U14223 ( .A(n14201), .B(n14202), .Z(n13980) );
  XOR2_X1 U14224 ( .A(n14203), .B(n14204), .Z(n14201) );
  XOR2_X1 U14225 ( .A(n14205), .B(n14206), .Z(n13985) );
  XNOR2_X1 U14226 ( .A(n14207), .B(n14208), .ZN(n14206) );
  XNOR2_X1 U14227 ( .A(n14209), .B(n14210), .ZN(n13989) );
  XNOR2_X1 U14228 ( .A(n14211), .B(n14212), .ZN(n14209) );
  XOR2_X1 U14229 ( .A(n14213), .B(n14214), .Z(n13992) );
  XOR2_X1 U14230 ( .A(n14215), .B(n14216), .Z(n14213) );
  XNOR2_X1 U14231 ( .A(n14217), .B(n14218), .ZN(n13997) );
  XNOR2_X1 U14232 ( .A(n14219), .B(n14220), .ZN(n14217) );
  XNOR2_X1 U14233 ( .A(n14221), .B(n14222), .ZN(n14001) );
  XOR2_X1 U14234 ( .A(n14223), .B(n14224), .Z(n14221) );
  XNOR2_X1 U14235 ( .A(n14225), .B(n14226), .ZN(n14005) );
  XNOR2_X1 U14236 ( .A(n14227), .B(n14228), .ZN(n14225) );
  XNOR2_X1 U14237 ( .A(n14229), .B(n14230), .ZN(n14009) );
  XOR2_X1 U14238 ( .A(n14231), .B(n14232), .Z(n14229) );
  XNOR2_X1 U14239 ( .A(n14233), .B(n14234), .ZN(n14013) );
  XNOR2_X1 U14240 ( .A(n14235), .B(n14236), .ZN(n14233) );
  XNOR2_X1 U14241 ( .A(n14237), .B(n14238), .ZN(n14017) );
  XNOR2_X1 U14242 ( .A(n14239), .B(n14240), .ZN(n14237) );
  XNOR2_X1 U14243 ( .A(n14241), .B(n14242), .ZN(n14021) );
  XNOR2_X1 U14244 ( .A(n14243), .B(n14244), .ZN(n14241) );
  NOR2_X1 U14245 ( .A1(n7789), .A2(n8054), .ZN(n14244) );
  XNOR2_X1 U14246 ( .A(n14245), .B(n14246), .ZN(n14025) );
  XNOR2_X1 U14247 ( .A(n14247), .B(n14248), .ZN(n14245) );
  NOR2_X1 U14248 ( .A1(n8669), .A2(n8054), .ZN(n14248) );
  XOR2_X1 U14249 ( .A(n14249), .B(n14250), .Z(n14029) );
  XNOR2_X1 U14250 ( .A(n14251), .B(n14252), .ZN(n14250) );
  NAND2_X1 U14251 ( .A1(b_4_), .A2(a_11_), .ZN(n14252) );
  XNOR2_X1 U14252 ( .A(n14253), .B(n14254), .ZN(n14033) );
  XNOR2_X1 U14253 ( .A(n14255), .B(n14256), .ZN(n14254) );
  NAND2_X1 U14254 ( .A1(b_4_), .A2(a_10_), .ZN(n14256) );
  XOR2_X1 U14255 ( .A(n14257), .B(n14258), .Z(n14037) );
  XNOR2_X1 U14256 ( .A(n14259), .B(n14260), .ZN(n14258) );
  NAND2_X1 U14257 ( .A1(b_4_), .A2(a_9_), .ZN(n14260) );
  XNOR2_X1 U14258 ( .A(n14261), .B(n14262), .ZN(n13870) );
  XOR2_X1 U14259 ( .A(n14263), .B(n14264), .Z(n14261) );
  NOR2_X1 U14260 ( .A1(n8686), .A2(n8054), .ZN(n14264) );
  XOR2_X1 U14261 ( .A(n14265), .B(n14266), .Z(n14041) );
  XOR2_X1 U14262 ( .A(n14267), .B(n14268), .Z(n14265) );
  NOR2_X1 U14263 ( .A1(n7872), .A2(n8054), .ZN(n14268) );
  INV_X1 U14264 ( .A(n7983), .ZN(n7899) );
  NAND2_X1 U14265 ( .A1(a_5_), .A2(b_5_), .ZN(n7983) );
  XOR2_X1 U14266 ( .A(n14269), .B(n14270), .Z(n14048) );
  XOR2_X1 U14267 ( .A(n14271), .B(n14272), .Z(n14269) );
  NOR2_X1 U14268 ( .A1(n7908), .A2(n8054), .ZN(n14272) );
  XOR2_X1 U14269 ( .A(n14273), .B(n14274), .Z(n14052) );
  XOR2_X1 U14270 ( .A(n14275), .B(n14276), .Z(n14273) );
  XOR2_X1 U14271 ( .A(n14277), .B(n14278), .Z(n14056) );
  XOR2_X1 U14272 ( .A(n14279), .B(n14280), .Z(n14277) );
  NOR2_X1 U14273 ( .A1(n8054), .A2(n7937), .ZN(n14280) );
  XOR2_X1 U14274 ( .A(n14281), .B(n14282), .Z(n14060) );
  XOR2_X1 U14275 ( .A(n14283), .B(n14284), .Z(n14281) );
  NOR2_X1 U14276 ( .A1(n8054), .A2(n8056), .ZN(n14284) );
  XOR2_X1 U14277 ( .A(n14285), .B(n14286), .Z(n14066) );
  XOR2_X1 U14278 ( .A(n14287), .B(n14288), .Z(n14285) );
  NOR2_X1 U14279 ( .A1(n7957), .A2(n8054), .ZN(n14288) );
  XNOR2_X1 U14280 ( .A(n14289), .B(n14290), .ZN(n14064) );
  XOR2_X1 U14281 ( .A(n14291), .B(n14292), .Z(n14289) );
  NOR2_X1 U14282 ( .A1(n8054), .A2(n8942), .ZN(n14292) );
  NAND2_X1 U14283 ( .A1(n14293), .A2(n14294), .ZN(n7862) );
  NAND2_X1 U14284 ( .A1(n14295), .A2(n14296), .ZN(n14294) );
  NAND2_X1 U14285 ( .A1(n14072), .A2(n14071), .ZN(n14293) );
  NAND4_X1 U14286 ( .A1(n14072), .A2(n14295), .A3(n14071), .A4(n14296), .ZN(
        n7861) );
  NAND2_X1 U14287 ( .A1(n14297), .A2(n14298), .ZN(n14071) );
  NAND3_X1 U14288 ( .A1(b_4_), .A2(n14299), .A3(a_0_), .ZN(n14298) );
  OR2_X1 U14289 ( .A1(n14291), .A2(n14290), .ZN(n14299) );
  NAND2_X1 U14290 ( .A1(n14290), .A2(n14291), .ZN(n14297) );
  NAND2_X1 U14291 ( .A1(n14300), .A2(n14301), .ZN(n14291) );
  NAND3_X1 U14292 ( .A1(a_1_), .A2(n14302), .A3(b_4_), .ZN(n14301) );
  OR2_X1 U14293 ( .A1(n14287), .A2(n14286), .ZN(n14302) );
  NAND2_X1 U14294 ( .A1(n14286), .A2(n14287), .ZN(n14300) );
  NAND2_X1 U14295 ( .A1(n14303), .A2(n14304), .ZN(n14287) );
  NAND3_X1 U14296 ( .A1(b_4_), .A2(n14305), .A3(a_2_), .ZN(n14304) );
  OR2_X1 U14297 ( .A1(n14282), .A2(n14283), .ZN(n14305) );
  NAND2_X1 U14298 ( .A1(n14282), .A2(n14283), .ZN(n14303) );
  NAND2_X1 U14299 ( .A1(n14306), .A2(n14307), .ZN(n14283) );
  NAND3_X1 U14300 ( .A1(b_4_), .A2(n14308), .A3(a_3_), .ZN(n14307) );
  OR2_X1 U14301 ( .A1(n14279), .A2(n14278), .ZN(n14308) );
  NAND2_X1 U14302 ( .A1(n14278), .A2(n14279), .ZN(n14306) );
  NAND2_X1 U14303 ( .A1(n14309), .A2(n14310), .ZN(n14279) );
  NAND2_X1 U14304 ( .A1(n14274), .A2(n14311), .ZN(n14310) );
  OR2_X1 U14305 ( .A1(n14275), .A2(n14276), .ZN(n14311) );
  XNOR2_X1 U14306 ( .A(n14312), .B(n14313), .ZN(n14274) );
  NAND2_X1 U14307 ( .A1(n14314), .A2(n14315), .ZN(n14312) );
  NAND2_X1 U14308 ( .A1(n14276), .A2(n14275), .ZN(n14309) );
  NAND2_X1 U14309 ( .A1(n14316), .A2(n14317), .ZN(n14275) );
  NAND3_X1 U14310 ( .A1(a_5_), .A2(n14318), .A3(b_4_), .ZN(n14317) );
  OR2_X1 U14311 ( .A1(n14271), .A2(n14270), .ZN(n14318) );
  NAND2_X1 U14312 ( .A1(n14270), .A2(n14271), .ZN(n14316) );
  NAND2_X1 U14313 ( .A1(n14319), .A2(n14320), .ZN(n14271) );
  NAND3_X1 U14314 ( .A1(a_6_), .A2(n14321), .A3(b_4_), .ZN(n14320) );
  NAND2_X1 U14315 ( .A1(n14094), .A2(n14093), .ZN(n14321) );
  OR2_X1 U14316 ( .A1(n14093), .A2(n14094), .ZN(n14319) );
  AND2_X1 U14317 ( .A1(n14322), .A2(n14323), .ZN(n14094) );
  NAND3_X1 U14318 ( .A1(a_7_), .A2(n14324), .A3(b_4_), .ZN(n14323) );
  OR2_X1 U14319 ( .A1(n14267), .A2(n14266), .ZN(n14324) );
  NAND2_X1 U14320 ( .A1(n14266), .A2(n14267), .ZN(n14322) );
  NAND2_X1 U14321 ( .A1(n14325), .A2(n14326), .ZN(n14267) );
  NAND3_X1 U14322 ( .A1(a_8_), .A2(n14327), .A3(b_4_), .ZN(n14326) );
  OR2_X1 U14323 ( .A1(n14263), .A2(n14262), .ZN(n14327) );
  NAND2_X1 U14324 ( .A1(n14262), .A2(n14263), .ZN(n14325) );
  NAND2_X1 U14325 ( .A1(n14328), .A2(n14329), .ZN(n14263) );
  NAND3_X1 U14326 ( .A1(a_9_), .A2(n14330), .A3(b_4_), .ZN(n14329) );
  NAND2_X1 U14327 ( .A1(n14259), .A2(n14257), .ZN(n14330) );
  OR2_X1 U14328 ( .A1(n14257), .A2(n14259), .ZN(n14328) );
  AND2_X1 U14329 ( .A1(n14331), .A2(n14332), .ZN(n14259) );
  NAND3_X1 U14330 ( .A1(a_10_), .A2(n14333), .A3(b_4_), .ZN(n14332) );
  NAND2_X1 U14331 ( .A1(n14255), .A2(n14253), .ZN(n14333) );
  OR2_X1 U14332 ( .A1(n14253), .A2(n14255), .ZN(n14331) );
  AND2_X1 U14333 ( .A1(n14334), .A2(n14335), .ZN(n14255) );
  NAND3_X1 U14334 ( .A1(a_11_), .A2(n14336), .A3(b_4_), .ZN(n14335) );
  NAND2_X1 U14335 ( .A1(n14251), .A2(n14249), .ZN(n14336) );
  OR2_X1 U14336 ( .A1(n14249), .A2(n14251), .ZN(n14334) );
  AND2_X1 U14337 ( .A1(n14337), .A2(n14338), .ZN(n14251) );
  NAND3_X1 U14338 ( .A1(a_12_), .A2(n14339), .A3(b_4_), .ZN(n14338) );
  NAND2_X1 U14339 ( .A1(n14247), .A2(n14246), .ZN(n14339) );
  OR2_X1 U14340 ( .A1(n14246), .A2(n14247), .ZN(n14337) );
  AND2_X1 U14341 ( .A1(n14340), .A2(n14341), .ZN(n14247) );
  NAND3_X1 U14342 ( .A1(a_13_), .A2(n14342), .A3(b_4_), .ZN(n14341) );
  NAND2_X1 U14343 ( .A1(n14243), .A2(n14242), .ZN(n14342) );
  OR2_X1 U14344 ( .A1(n14242), .A2(n14243), .ZN(n14340) );
  AND2_X1 U14345 ( .A1(n14343), .A2(n14344), .ZN(n14243) );
  NAND2_X1 U14346 ( .A1(n14240), .A2(n14345), .ZN(n14344) );
  NAND2_X1 U14347 ( .A1(n14239), .A2(n14238), .ZN(n14345) );
  NOR2_X1 U14348 ( .A1(n8054), .A2(n8049), .ZN(n14240) );
  OR2_X1 U14349 ( .A1(n14238), .A2(n14239), .ZN(n14343) );
  AND2_X1 U14350 ( .A1(n14346), .A2(n14347), .ZN(n14239) );
  NAND2_X1 U14351 ( .A1(n14236), .A2(n14348), .ZN(n14347) );
  NAND2_X1 U14352 ( .A1(n14235), .A2(n14234), .ZN(n14348) );
  NOR2_X1 U14353 ( .A1(n8054), .A2(n7754), .ZN(n14236) );
  OR2_X1 U14354 ( .A1(n14234), .A2(n14235), .ZN(n14346) );
  AND2_X1 U14355 ( .A1(n14349), .A2(n14350), .ZN(n14235) );
  NAND2_X1 U14356 ( .A1(n14232), .A2(n14351), .ZN(n14350) );
  OR2_X1 U14357 ( .A1(n14230), .A2(n14231), .ZN(n14351) );
  NOR2_X1 U14358 ( .A1(n8054), .A2(n8438), .ZN(n14232) );
  NAND2_X1 U14359 ( .A1(n14230), .A2(n14231), .ZN(n14349) );
  NAND2_X1 U14360 ( .A1(n14352), .A2(n14353), .ZN(n14231) );
  NAND2_X1 U14361 ( .A1(n14228), .A2(n14354), .ZN(n14353) );
  NAND2_X1 U14362 ( .A1(n14227), .A2(n14226), .ZN(n14354) );
  NOR2_X1 U14363 ( .A1(n8054), .A2(n7732), .ZN(n14228) );
  OR2_X1 U14364 ( .A1(n14226), .A2(n14227), .ZN(n14352) );
  AND2_X1 U14365 ( .A1(n14355), .A2(n14356), .ZN(n14227) );
  NAND2_X1 U14366 ( .A1(n14224), .A2(n14357), .ZN(n14356) );
  OR2_X1 U14367 ( .A1(n14222), .A2(n14223), .ZN(n14357) );
  NOR2_X1 U14368 ( .A1(n8054), .A2(n8047), .ZN(n14224) );
  NAND2_X1 U14369 ( .A1(n14222), .A2(n14223), .ZN(n14355) );
  NAND2_X1 U14370 ( .A1(n14358), .A2(n14359), .ZN(n14223) );
  NAND2_X1 U14371 ( .A1(n14220), .A2(n14360), .ZN(n14359) );
  NAND2_X1 U14372 ( .A1(n14219), .A2(n14218), .ZN(n14360) );
  NOR2_X1 U14373 ( .A1(n8054), .A2(n8045), .ZN(n14220) );
  OR2_X1 U14374 ( .A1(n14218), .A2(n14219), .ZN(n14358) );
  AND2_X1 U14375 ( .A1(n14361), .A2(n14362), .ZN(n14219) );
  NAND2_X1 U14376 ( .A1(n14216), .A2(n14363), .ZN(n14362) );
  OR2_X1 U14377 ( .A1(n14214), .A2(n14215), .ZN(n14363) );
  NOR2_X1 U14378 ( .A1(n8054), .A2(n8044), .ZN(n14216) );
  NAND2_X1 U14379 ( .A1(n14214), .A2(n14215), .ZN(n14361) );
  NAND2_X1 U14380 ( .A1(n14364), .A2(n14365), .ZN(n14215) );
  NAND2_X1 U14381 ( .A1(n14211), .A2(n14366), .ZN(n14365) );
  NAND2_X1 U14382 ( .A1(n14212), .A2(n14210), .ZN(n14366) );
  NOR2_X1 U14383 ( .A1(n8054), .A2(n7665), .ZN(n14211) );
  OR2_X1 U14384 ( .A1(n14210), .A2(n14212), .ZN(n14364) );
  AND2_X1 U14385 ( .A1(n14367), .A2(n14368), .ZN(n14212) );
  NAND2_X1 U14386 ( .A1(n14208), .A2(n14369), .ZN(n14368) );
  OR2_X1 U14387 ( .A1(n14205), .A2(n14207), .ZN(n14369) );
  NOR2_X1 U14388 ( .A1(n8054), .A2(n7650), .ZN(n14208) );
  NAND2_X1 U14389 ( .A1(n14205), .A2(n14207), .ZN(n14367) );
  NAND2_X1 U14390 ( .A1(n14370), .A2(n14371), .ZN(n14207) );
  NAND2_X1 U14391 ( .A1(n14204), .A2(n14372), .ZN(n14371) );
  OR2_X1 U14392 ( .A1(n14202), .A2(n14203), .ZN(n14372) );
  NOR2_X1 U14393 ( .A1(n8054), .A2(n8042), .ZN(n14204) );
  NAND2_X1 U14394 ( .A1(n14202), .A2(n14203), .ZN(n14370) );
  NAND2_X1 U14395 ( .A1(n14373), .A2(n14374), .ZN(n14203) );
  NAND2_X1 U14396 ( .A1(n14200), .A2(n14375), .ZN(n14374) );
  OR2_X1 U14397 ( .A1(n14198), .A2(n14199), .ZN(n14375) );
  NOR2_X1 U14398 ( .A1(n8054), .A2(n8041), .ZN(n14200) );
  NAND2_X1 U14399 ( .A1(n14198), .A2(n14199), .ZN(n14373) );
  NAND2_X1 U14400 ( .A1(n14376), .A2(n14377), .ZN(n14199) );
  NAND2_X1 U14401 ( .A1(n14196), .A2(n14378), .ZN(n14377) );
  OR2_X1 U14402 ( .A1(n14194), .A2(n14195), .ZN(n14378) );
  NOR2_X1 U14403 ( .A1(n8054), .A2(n8039), .ZN(n14196) );
  NAND2_X1 U14404 ( .A1(n14194), .A2(n14195), .ZN(n14376) );
  NAND2_X1 U14405 ( .A1(n14159), .A2(n14379), .ZN(n14195) );
  NAND2_X1 U14406 ( .A1(n14158), .A2(n14160), .ZN(n14379) );
  NAND2_X1 U14407 ( .A1(n14380), .A2(n14381), .ZN(n14160) );
  NAND2_X1 U14408 ( .A1(b_4_), .A2(a_26_), .ZN(n14381) );
  INV_X1 U14409 ( .A(n14382), .ZN(n14380) );
  XNOR2_X1 U14410 ( .A(n14383), .B(n14384), .ZN(n14158) );
  NAND2_X1 U14411 ( .A1(n14385), .A2(n14386), .ZN(n14383) );
  NAND2_X1 U14412 ( .A1(a_26_), .A2(n14382), .ZN(n14159) );
  NAND2_X1 U14413 ( .A1(n14167), .A2(n14387), .ZN(n14382) );
  NAND2_X1 U14414 ( .A1(n14166), .A2(n14168), .ZN(n14387) );
  NAND2_X1 U14415 ( .A1(n14388), .A2(n14389), .ZN(n14168) );
  NAND2_X1 U14416 ( .A1(b_4_), .A2(a_27_), .ZN(n14389) );
  INV_X1 U14417 ( .A(n14390), .ZN(n14388) );
  XNOR2_X1 U14418 ( .A(n14391), .B(n14392), .ZN(n14166) );
  XOR2_X1 U14419 ( .A(n14393), .B(n14394), .Z(n14391) );
  NAND2_X1 U14420 ( .A1(b_3_), .A2(a_28_), .ZN(n14393) );
  NAND2_X1 U14421 ( .A1(a_27_), .A2(n14390), .ZN(n14167) );
  NAND2_X1 U14422 ( .A1(n14395), .A2(n14396), .ZN(n14390) );
  NAND3_X1 U14423 ( .A1(a_28_), .A2(n14397), .A3(b_4_), .ZN(n14396) );
  NAND2_X1 U14424 ( .A1(n14176), .A2(n14174), .ZN(n14397) );
  OR2_X1 U14425 ( .A1(n14174), .A2(n14176), .ZN(n14395) );
  AND2_X1 U14426 ( .A1(n14398), .A2(n14399), .ZN(n14176) );
  NAND2_X1 U14427 ( .A1(n14190), .A2(n14400), .ZN(n14399) );
  OR2_X1 U14428 ( .A1(n14191), .A2(n14192), .ZN(n14400) );
  NOR2_X1 U14429 ( .A1(n8054), .A2(n7545), .ZN(n14190) );
  NAND2_X1 U14430 ( .A1(n14192), .A2(n14191), .ZN(n14398) );
  NAND2_X1 U14431 ( .A1(n14401), .A2(n14402), .ZN(n14191) );
  NAND2_X1 U14432 ( .A1(b_2_), .A2(n14403), .ZN(n14402) );
  NAND2_X1 U14433 ( .A1(n7527), .A2(n14404), .ZN(n14403) );
  NAND2_X1 U14434 ( .A1(a_31_), .A2(n7930), .ZN(n14404) );
  NAND2_X1 U14435 ( .A1(b_3_), .A2(n14405), .ZN(n14401) );
  NAND2_X1 U14436 ( .A1(n7531), .A2(n14406), .ZN(n14405) );
  NAND2_X1 U14437 ( .A1(a_30_), .A2(n8055), .ZN(n14406) );
  AND3_X1 U14438 ( .A1(b_4_), .A2(b_3_), .A3(n7494), .ZN(n14192) );
  XNOR2_X1 U14439 ( .A(n14407), .B(n14408), .ZN(n14174) );
  XOR2_X1 U14440 ( .A(n14409), .B(n14410), .Z(n14407) );
  XNOR2_X1 U14441 ( .A(n14411), .B(n14412), .ZN(n14194) );
  NAND2_X1 U14442 ( .A1(n14413), .A2(n14414), .ZN(n14411) );
  XNOR2_X1 U14443 ( .A(n14415), .B(n14416), .ZN(n14198) );
  NAND2_X1 U14444 ( .A1(n14417), .A2(n14418), .ZN(n14415) );
  XNOR2_X1 U14445 ( .A(n14419), .B(n14420), .ZN(n14202) );
  XNOR2_X1 U14446 ( .A(n14421), .B(n14422), .ZN(n14419) );
  NOR2_X1 U14447 ( .A1(n8041), .A2(n7930), .ZN(n14422) );
  XNOR2_X1 U14448 ( .A(n14423), .B(n14424), .ZN(n14205) );
  NAND2_X1 U14449 ( .A1(n14425), .A2(n14426), .ZN(n14423) );
  XNOR2_X1 U14450 ( .A(n14427), .B(n14428), .ZN(n14210) );
  XNOR2_X1 U14451 ( .A(n14429), .B(n14430), .ZN(n14427) );
  NAND2_X1 U14452 ( .A1(b_3_), .A2(a_22_), .ZN(n14429) );
  XNOR2_X1 U14453 ( .A(n14431), .B(n14432), .ZN(n14214) );
  NAND2_X1 U14454 ( .A1(n14433), .A2(n14434), .ZN(n14431) );
  XNOR2_X1 U14455 ( .A(n14435), .B(n14436), .ZN(n14218) );
  XNOR2_X1 U14456 ( .A(n14437), .B(n14438), .ZN(n14435) );
  NAND2_X1 U14457 ( .A1(b_3_), .A2(a_20_), .ZN(n14437) );
  XNOR2_X1 U14458 ( .A(n14439), .B(n14440), .ZN(n14222) );
  NAND2_X1 U14459 ( .A1(n14441), .A2(n14442), .ZN(n14439) );
  XNOR2_X1 U14460 ( .A(n14443), .B(n14444), .ZN(n14226) );
  XNOR2_X1 U14461 ( .A(n14445), .B(n14446), .ZN(n14443) );
  NAND2_X1 U14462 ( .A1(b_3_), .A2(a_18_), .ZN(n14445) );
  XNOR2_X1 U14463 ( .A(n14447), .B(n14448), .ZN(n14230) );
  NAND2_X1 U14464 ( .A1(n14449), .A2(n14450), .ZN(n14447) );
  XNOR2_X1 U14465 ( .A(n14451), .B(n14452), .ZN(n14234) );
  XNOR2_X1 U14466 ( .A(n14453), .B(n14454), .ZN(n14451) );
  NAND2_X1 U14467 ( .A1(b_3_), .A2(a_16_), .ZN(n14453) );
  XOR2_X1 U14468 ( .A(n14455), .B(n14456), .Z(n14238) );
  NAND2_X1 U14469 ( .A1(n14457), .A2(n14458), .ZN(n14455) );
  XNOR2_X1 U14470 ( .A(n14459), .B(n14460), .ZN(n14242) );
  XNOR2_X1 U14471 ( .A(n14461), .B(n14462), .ZN(n14459) );
  NAND2_X1 U14472 ( .A1(b_3_), .A2(a_14_), .ZN(n14461) );
  XOR2_X1 U14473 ( .A(n14463), .B(n14464), .Z(n14246) );
  NAND2_X1 U14474 ( .A1(n14465), .A2(n14466), .ZN(n14463) );
  XNOR2_X1 U14475 ( .A(n14467), .B(n14468), .ZN(n14249) );
  XNOR2_X1 U14476 ( .A(n14469), .B(n14470), .ZN(n14467) );
  NAND2_X1 U14477 ( .A1(b_3_), .A2(a_12_), .ZN(n14469) );
  XOR2_X1 U14478 ( .A(n14471), .B(n14472), .Z(n14253) );
  NAND2_X1 U14479 ( .A1(n14473), .A2(n14474), .ZN(n14471) );
  XNOR2_X1 U14480 ( .A(n14475), .B(n14476), .ZN(n14257) );
  XNOR2_X1 U14481 ( .A(n14477), .B(n14478), .ZN(n14475) );
  NAND2_X1 U14482 ( .A1(b_3_), .A2(a_10_), .ZN(n14477) );
  XNOR2_X1 U14483 ( .A(n14479), .B(n14480), .ZN(n14262) );
  NAND2_X1 U14484 ( .A1(n14481), .A2(n14482), .ZN(n14479) );
  XOR2_X1 U14485 ( .A(n14483), .B(n14484), .Z(n14266) );
  XNOR2_X1 U14486 ( .A(n14485), .B(n14486), .ZN(n14483) );
  NAND2_X1 U14487 ( .A1(b_3_), .A2(a_8_), .ZN(n14485) );
  XOR2_X1 U14488 ( .A(n14487), .B(n14488), .Z(n14093) );
  NAND2_X1 U14489 ( .A1(n14489), .A2(n14490), .ZN(n14487) );
  XOR2_X1 U14490 ( .A(n14491), .B(n14492), .Z(n14270) );
  XNOR2_X1 U14491 ( .A(n14493), .B(n14494), .ZN(n14491) );
  NAND2_X1 U14492 ( .A1(b_3_), .A2(a_6_), .ZN(n14493) );
  INV_X1 U14493 ( .A(n7921), .ZN(n14276) );
  NAND2_X1 U14494 ( .A1(b_4_), .A2(a_4_), .ZN(n7921) );
  XOR2_X1 U14495 ( .A(n14495), .B(n14496), .Z(n14278) );
  XNOR2_X1 U14496 ( .A(n14497), .B(n14498), .ZN(n14495) );
  NAND2_X1 U14497 ( .A1(b_3_), .A2(a_4_), .ZN(n14497) );
  XOR2_X1 U14498 ( .A(n14499), .B(n14500), .Z(n14282) );
  XOR2_X1 U14499 ( .A(n14501), .B(n7928), .Z(n14499) );
  XOR2_X1 U14500 ( .A(n14502), .B(n14503), .Z(n14286) );
  XNOR2_X1 U14501 ( .A(n14504), .B(n14505), .ZN(n14502) );
  NAND2_X1 U14502 ( .A1(a_2_), .A2(b_3_), .ZN(n14504) );
  XOR2_X1 U14503 ( .A(n14506), .B(n14507), .Z(n14290) );
  XOR2_X1 U14504 ( .A(n14508), .B(n14509), .Z(n14506) );
  NAND2_X1 U14505 ( .A1(n14510), .A2(n14511), .ZN(n14295) );
  XOR2_X1 U14506 ( .A(n14512), .B(n14513), .Z(n14072) );
  XOR2_X1 U14507 ( .A(n14514), .B(n14515), .Z(n14512) );
  NAND2_X1 U14508 ( .A1(n14516), .A2(n14296), .ZN(n8068) );
  INV_X1 U14509 ( .A(n14517), .ZN(n14296) );
  XNOR2_X1 U14510 ( .A(n8176), .B(n8177), .ZN(n14516) );
  NAND2_X1 U14511 ( .A1(n14517), .A2(n14518), .ZN(n8067) );
  XOR2_X1 U14512 ( .A(n8177), .B(n8176), .Z(n14518) );
  NAND3_X1 U14513 ( .A1(n14519), .A2(n14520), .A3(n14521), .ZN(n8176) );
  XNOR2_X1 U14514 ( .A(n8180), .B(n8181), .ZN(n14521) );
  NOR2_X1 U14515 ( .A1(n7957), .A2(n14522), .ZN(n8181) );
  NOR2_X1 U14516 ( .A1(n8942), .A2(n14523), .ZN(n8180) );
  NAND3_X1 U14517 ( .A1(a_2_), .A2(b_0_), .A3(n7963), .ZN(n14520) );
  NAND2_X1 U14518 ( .A1(n14524), .A2(n14525), .ZN(n8177) );
  NAND2_X1 U14519 ( .A1(n14526), .A2(b_2_), .ZN(n14525) );
  NOR2_X1 U14520 ( .A1(n14511), .A2(n14510), .ZN(n14517) );
  AND2_X1 U14521 ( .A1(n14527), .A2(n14528), .ZN(n14510) );
  NAND2_X1 U14522 ( .A1(n14514), .A2(n14529), .ZN(n14528) );
  OR2_X1 U14523 ( .A1(n14513), .A2(n14515), .ZN(n14529) );
  NOR2_X1 U14524 ( .A1(n8942), .A2(n7930), .ZN(n14514) );
  NAND2_X1 U14525 ( .A1(n14513), .A2(n14515), .ZN(n14527) );
  NAND2_X1 U14526 ( .A1(n14530), .A2(n14531), .ZN(n14515) );
  NAND2_X1 U14527 ( .A1(n14509), .A2(n14532), .ZN(n14531) );
  OR2_X1 U14528 ( .A1(n14507), .A2(n14508), .ZN(n14532) );
  NOR2_X1 U14529 ( .A1(n7930), .A2(n7957), .ZN(n14509) );
  NAND2_X1 U14530 ( .A1(n14507), .A2(n14508), .ZN(n14530) );
  NAND2_X1 U14531 ( .A1(n14533), .A2(n14534), .ZN(n14508) );
  NAND3_X1 U14532 ( .A1(b_3_), .A2(n14535), .A3(a_2_), .ZN(n14534) );
  OR2_X1 U14533 ( .A1(n14503), .A2(n14505), .ZN(n14535) );
  NAND2_X1 U14534 ( .A1(n14503), .A2(n14505), .ZN(n14533) );
  NAND2_X1 U14535 ( .A1(n14536), .A2(n14537), .ZN(n14505) );
  NAND2_X1 U14536 ( .A1(n14500), .A2(n14538), .ZN(n14537) );
  OR2_X1 U14537 ( .A1(n14501), .A2(n7928), .ZN(n14538) );
  XNOR2_X1 U14538 ( .A(n14539), .B(n14540), .ZN(n14500) );
  NAND2_X1 U14539 ( .A1(n14541), .A2(n14542), .ZN(n14539) );
  NAND2_X1 U14540 ( .A1(n7928), .A2(n14501), .ZN(n14536) );
  NAND2_X1 U14541 ( .A1(n14543), .A2(n14544), .ZN(n14501) );
  NAND3_X1 U14542 ( .A1(a_4_), .A2(n14545), .A3(b_3_), .ZN(n14544) );
  OR2_X1 U14543 ( .A1(n14496), .A2(n14498), .ZN(n14545) );
  NAND2_X1 U14544 ( .A1(n14496), .A2(n14498), .ZN(n14543) );
  NAND2_X1 U14545 ( .A1(n14314), .A2(n14546), .ZN(n14498) );
  NAND2_X1 U14546 ( .A1(n14313), .A2(n14315), .ZN(n14546) );
  NAND2_X1 U14547 ( .A1(n14547), .A2(n14548), .ZN(n14315) );
  NAND2_X1 U14548 ( .A1(b_3_), .A2(a_5_), .ZN(n14548) );
  INV_X1 U14549 ( .A(n14549), .ZN(n14547) );
  XNOR2_X1 U14550 ( .A(n14550), .B(n14551), .ZN(n14313) );
  NAND2_X1 U14551 ( .A1(n14552), .A2(n14553), .ZN(n14550) );
  NAND2_X1 U14552 ( .A1(a_5_), .A2(n14549), .ZN(n14314) );
  NAND2_X1 U14553 ( .A1(n14554), .A2(n14555), .ZN(n14549) );
  NAND3_X1 U14554 ( .A1(a_6_), .A2(n14556), .A3(b_3_), .ZN(n14555) );
  OR2_X1 U14555 ( .A1(n14492), .A2(n14494), .ZN(n14556) );
  NAND2_X1 U14556 ( .A1(n14492), .A2(n14494), .ZN(n14554) );
  NAND2_X1 U14557 ( .A1(n14489), .A2(n14557), .ZN(n14494) );
  NAND2_X1 U14558 ( .A1(n14488), .A2(n14490), .ZN(n14557) );
  NAND2_X1 U14559 ( .A1(n14558), .A2(n14559), .ZN(n14490) );
  NAND2_X1 U14560 ( .A1(b_3_), .A2(a_7_), .ZN(n14559) );
  INV_X1 U14561 ( .A(n14560), .ZN(n14558) );
  XNOR2_X1 U14562 ( .A(n14561), .B(n14562), .ZN(n14488) );
  NAND2_X1 U14563 ( .A1(n14563), .A2(n14564), .ZN(n14561) );
  NAND2_X1 U14564 ( .A1(a_7_), .A2(n14560), .ZN(n14489) );
  NAND2_X1 U14565 ( .A1(n14565), .A2(n14566), .ZN(n14560) );
  NAND3_X1 U14566 ( .A1(a_8_), .A2(n14567), .A3(b_3_), .ZN(n14566) );
  OR2_X1 U14567 ( .A1(n14484), .A2(n14486), .ZN(n14567) );
  NAND2_X1 U14568 ( .A1(n14484), .A2(n14486), .ZN(n14565) );
  NAND2_X1 U14569 ( .A1(n14481), .A2(n14568), .ZN(n14486) );
  NAND2_X1 U14570 ( .A1(n14480), .A2(n14482), .ZN(n14568) );
  NAND2_X1 U14571 ( .A1(n14569), .A2(n14570), .ZN(n14482) );
  NAND2_X1 U14572 ( .A1(b_3_), .A2(a_9_), .ZN(n14570) );
  INV_X1 U14573 ( .A(n14571), .ZN(n14569) );
  XNOR2_X1 U14574 ( .A(n14572), .B(n14573), .ZN(n14480) );
  NAND2_X1 U14575 ( .A1(n14574), .A2(n14575), .ZN(n14572) );
  NAND2_X1 U14576 ( .A1(a_9_), .A2(n14571), .ZN(n14481) );
  NAND2_X1 U14577 ( .A1(n14576), .A2(n14577), .ZN(n14571) );
  NAND3_X1 U14578 ( .A1(a_10_), .A2(n14578), .A3(b_3_), .ZN(n14577) );
  OR2_X1 U14579 ( .A1(n14476), .A2(n14478), .ZN(n14578) );
  NAND2_X1 U14580 ( .A1(n14476), .A2(n14478), .ZN(n14576) );
  NAND2_X1 U14581 ( .A1(n14473), .A2(n14579), .ZN(n14478) );
  NAND2_X1 U14582 ( .A1(n14472), .A2(n14474), .ZN(n14579) );
  NAND2_X1 U14583 ( .A1(n14580), .A2(n14581), .ZN(n14474) );
  NAND2_X1 U14584 ( .A1(b_3_), .A2(a_11_), .ZN(n14581) );
  INV_X1 U14585 ( .A(n14582), .ZN(n14580) );
  XNOR2_X1 U14586 ( .A(n14583), .B(n14584), .ZN(n14472) );
  NAND2_X1 U14587 ( .A1(n14585), .A2(n14586), .ZN(n14583) );
  NAND2_X1 U14588 ( .A1(a_11_), .A2(n14582), .ZN(n14473) );
  NAND2_X1 U14589 ( .A1(n14587), .A2(n14588), .ZN(n14582) );
  NAND3_X1 U14590 ( .A1(a_12_), .A2(n14589), .A3(b_3_), .ZN(n14588) );
  OR2_X1 U14591 ( .A1(n14468), .A2(n14470), .ZN(n14589) );
  NAND2_X1 U14592 ( .A1(n14468), .A2(n14470), .ZN(n14587) );
  NAND2_X1 U14593 ( .A1(n14465), .A2(n14590), .ZN(n14470) );
  NAND2_X1 U14594 ( .A1(n14464), .A2(n14466), .ZN(n14590) );
  NAND2_X1 U14595 ( .A1(n14591), .A2(n14592), .ZN(n14466) );
  NAND2_X1 U14596 ( .A1(b_3_), .A2(a_13_), .ZN(n14592) );
  INV_X1 U14597 ( .A(n14593), .ZN(n14591) );
  XNOR2_X1 U14598 ( .A(n14594), .B(n14595), .ZN(n14464) );
  NAND2_X1 U14599 ( .A1(n14596), .A2(n14597), .ZN(n14594) );
  NAND2_X1 U14600 ( .A1(a_13_), .A2(n14593), .ZN(n14465) );
  NAND2_X1 U14601 ( .A1(n14598), .A2(n14599), .ZN(n14593) );
  NAND3_X1 U14602 ( .A1(a_14_), .A2(n14600), .A3(b_3_), .ZN(n14599) );
  OR2_X1 U14603 ( .A1(n14460), .A2(n14462), .ZN(n14600) );
  NAND2_X1 U14604 ( .A1(n14460), .A2(n14462), .ZN(n14598) );
  NAND2_X1 U14605 ( .A1(n14457), .A2(n14601), .ZN(n14462) );
  NAND2_X1 U14606 ( .A1(n14456), .A2(n14458), .ZN(n14601) );
  NAND2_X1 U14607 ( .A1(n14602), .A2(n14603), .ZN(n14458) );
  NAND2_X1 U14608 ( .A1(b_3_), .A2(a_15_), .ZN(n14603) );
  INV_X1 U14609 ( .A(n14604), .ZN(n14602) );
  XNOR2_X1 U14610 ( .A(n14605), .B(n14606), .ZN(n14456) );
  NAND2_X1 U14611 ( .A1(n14607), .A2(n14608), .ZN(n14605) );
  NAND2_X1 U14612 ( .A1(a_15_), .A2(n14604), .ZN(n14457) );
  NAND2_X1 U14613 ( .A1(n14609), .A2(n14610), .ZN(n14604) );
  NAND3_X1 U14614 ( .A1(a_16_), .A2(n14611), .A3(b_3_), .ZN(n14610) );
  OR2_X1 U14615 ( .A1(n14452), .A2(n14454), .ZN(n14611) );
  NAND2_X1 U14616 ( .A1(n14452), .A2(n14454), .ZN(n14609) );
  NAND2_X1 U14617 ( .A1(n14449), .A2(n14612), .ZN(n14454) );
  NAND2_X1 U14618 ( .A1(n14448), .A2(n14450), .ZN(n14612) );
  NAND2_X1 U14619 ( .A1(n14613), .A2(n14614), .ZN(n14450) );
  NAND2_X1 U14620 ( .A1(b_3_), .A2(a_17_), .ZN(n14614) );
  INV_X1 U14621 ( .A(n14615), .ZN(n14613) );
  XNOR2_X1 U14622 ( .A(n14616), .B(n14617), .ZN(n14448) );
  XNOR2_X1 U14623 ( .A(n14618), .B(n14619), .ZN(n14617) );
  NAND2_X1 U14624 ( .A1(a_17_), .A2(n14615), .ZN(n14449) );
  NAND2_X1 U14625 ( .A1(n14620), .A2(n14621), .ZN(n14615) );
  NAND3_X1 U14626 ( .A1(a_18_), .A2(n14622), .A3(b_3_), .ZN(n14621) );
  OR2_X1 U14627 ( .A1(n14444), .A2(n14446), .ZN(n14622) );
  NAND2_X1 U14628 ( .A1(n14444), .A2(n14446), .ZN(n14620) );
  NAND2_X1 U14629 ( .A1(n14441), .A2(n14623), .ZN(n14446) );
  NAND2_X1 U14630 ( .A1(n14440), .A2(n14442), .ZN(n14623) );
  NAND2_X1 U14631 ( .A1(n14624), .A2(n14625), .ZN(n14442) );
  NAND2_X1 U14632 ( .A1(b_3_), .A2(a_19_), .ZN(n14625) );
  INV_X1 U14633 ( .A(n14626), .ZN(n14624) );
  XNOR2_X1 U14634 ( .A(n14627), .B(n14628), .ZN(n14440) );
  XNOR2_X1 U14635 ( .A(n14629), .B(n14630), .ZN(n14628) );
  NAND2_X1 U14636 ( .A1(a_19_), .A2(n14626), .ZN(n14441) );
  NAND2_X1 U14637 ( .A1(n14631), .A2(n14632), .ZN(n14626) );
  NAND3_X1 U14638 ( .A1(a_20_), .A2(n14633), .A3(b_3_), .ZN(n14632) );
  OR2_X1 U14639 ( .A1(n14436), .A2(n14438), .ZN(n14633) );
  NAND2_X1 U14640 ( .A1(n14436), .A2(n14438), .ZN(n14631) );
  NAND2_X1 U14641 ( .A1(n14433), .A2(n14634), .ZN(n14438) );
  NAND2_X1 U14642 ( .A1(n14432), .A2(n14434), .ZN(n14634) );
  NAND2_X1 U14643 ( .A1(n14635), .A2(n14636), .ZN(n14434) );
  NAND2_X1 U14644 ( .A1(b_3_), .A2(a_21_), .ZN(n14636) );
  INV_X1 U14645 ( .A(n14637), .ZN(n14635) );
  XNOR2_X1 U14646 ( .A(n14638), .B(n14639), .ZN(n14432) );
  XNOR2_X1 U14647 ( .A(n14640), .B(n14641), .ZN(n14639) );
  NAND2_X1 U14648 ( .A1(a_21_), .A2(n14637), .ZN(n14433) );
  NAND2_X1 U14649 ( .A1(n14642), .A2(n14643), .ZN(n14637) );
  NAND3_X1 U14650 ( .A1(a_22_), .A2(n14644), .A3(b_3_), .ZN(n14643) );
  OR2_X1 U14651 ( .A1(n14428), .A2(n14430), .ZN(n14644) );
  NAND2_X1 U14652 ( .A1(n14428), .A2(n14430), .ZN(n14642) );
  NAND2_X1 U14653 ( .A1(n14425), .A2(n14645), .ZN(n14430) );
  NAND2_X1 U14654 ( .A1(n14424), .A2(n14426), .ZN(n14645) );
  NAND2_X1 U14655 ( .A1(n14646), .A2(n14647), .ZN(n14426) );
  NAND2_X1 U14656 ( .A1(b_3_), .A2(a_23_), .ZN(n14647) );
  INV_X1 U14657 ( .A(n14648), .ZN(n14646) );
  XNOR2_X1 U14658 ( .A(n14649), .B(n14650), .ZN(n14424) );
  XNOR2_X1 U14659 ( .A(n14651), .B(n14652), .ZN(n14650) );
  NAND2_X1 U14660 ( .A1(a_23_), .A2(n14648), .ZN(n14425) );
  NAND2_X1 U14661 ( .A1(n14653), .A2(n14654), .ZN(n14648) );
  NAND3_X1 U14662 ( .A1(a_24_), .A2(n14655), .A3(b_3_), .ZN(n14654) );
  NAND2_X1 U14663 ( .A1(n14421), .A2(n14420), .ZN(n14655) );
  OR2_X1 U14664 ( .A1(n14420), .A2(n14421), .ZN(n14653) );
  AND2_X1 U14665 ( .A1(n14417), .A2(n14656), .ZN(n14421) );
  NAND2_X1 U14666 ( .A1(n14416), .A2(n14418), .ZN(n14656) );
  NAND2_X1 U14667 ( .A1(n14657), .A2(n14658), .ZN(n14418) );
  NAND2_X1 U14668 ( .A1(b_3_), .A2(a_25_), .ZN(n14658) );
  INV_X1 U14669 ( .A(n14659), .ZN(n14657) );
  XNOR2_X1 U14670 ( .A(n14660), .B(n14661), .ZN(n14416) );
  XOR2_X1 U14671 ( .A(n14662), .B(n14663), .Z(n14660) );
  NAND2_X1 U14672 ( .A1(b_2_), .A2(a_26_), .ZN(n14662) );
  NAND2_X1 U14673 ( .A1(a_25_), .A2(n14659), .ZN(n14417) );
  NAND2_X1 U14674 ( .A1(n14413), .A2(n14664), .ZN(n14659) );
  NAND2_X1 U14675 ( .A1(n14412), .A2(n14414), .ZN(n14664) );
  NAND2_X1 U14676 ( .A1(n14665), .A2(n14666), .ZN(n14414) );
  NAND2_X1 U14677 ( .A1(b_3_), .A2(a_26_), .ZN(n14666) );
  INV_X1 U14678 ( .A(n14667), .ZN(n14665) );
  XNOR2_X1 U14679 ( .A(n14668), .B(n14669), .ZN(n14412) );
  XNOR2_X1 U14680 ( .A(n14670), .B(n14671), .ZN(n14669) );
  NAND2_X1 U14681 ( .A1(a_26_), .A2(n14667), .ZN(n14413) );
  NAND2_X1 U14682 ( .A1(n14385), .A2(n14672), .ZN(n14667) );
  NAND2_X1 U14683 ( .A1(n14384), .A2(n14386), .ZN(n14672) );
  NAND2_X1 U14684 ( .A1(n14673), .A2(n14674), .ZN(n14386) );
  NAND2_X1 U14685 ( .A1(b_3_), .A2(a_27_), .ZN(n14674) );
  INV_X1 U14686 ( .A(n14675), .ZN(n14673) );
  XOR2_X1 U14687 ( .A(n14676), .B(n14677), .Z(n14384) );
  XNOR2_X1 U14688 ( .A(n14678), .B(n14679), .ZN(n14676) );
  NAND2_X1 U14689 ( .A1(b_2_), .A2(a_28_), .ZN(n14678) );
  NAND2_X1 U14690 ( .A1(a_27_), .A2(n14675), .ZN(n14385) );
  NAND2_X1 U14691 ( .A1(n14680), .A2(n14681), .ZN(n14675) );
  NAND3_X1 U14692 ( .A1(a_28_), .A2(n14682), .A3(b_3_), .ZN(n14681) );
  NAND2_X1 U14693 ( .A1(n14394), .A2(n14392), .ZN(n14682) );
  OR2_X1 U14694 ( .A1(n14392), .A2(n14394), .ZN(n14680) );
  AND2_X1 U14695 ( .A1(n14683), .A2(n14684), .ZN(n14394) );
  NAND2_X1 U14696 ( .A1(n14408), .A2(n14685), .ZN(n14684) );
  OR2_X1 U14697 ( .A1(n14409), .A2(n14410), .ZN(n14685) );
  NOR2_X1 U14698 ( .A1(n7930), .A2(n7545), .ZN(n14408) );
  NAND2_X1 U14699 ( .A1(n14410), .A2(n14409), .ZN(n14683) );
  NAND2_X1 U14700 ( .A1(n14686), .A2(n14687), .ZN(n14409) );
  NAND2_X1 U14701 ( .A1(b_1_), .A2(n14688), .ZN(n14687) );
  NAND2_X1 U14702 ( .A1(n7527), .A2(n14689), .ZN(n14688) );
  NAND2_X1 U14703 ( .A1(a_31_), .A2(n8055), .ZN(n14689) );
  NAND2_X1 U14704 ( .A1(b_2_), .A2(n14690), .ZN(n14686) );
  NAND2_X1 U14705 ( .A1(n7531), .A2(n14691), .ZN(n14690) );
  NAND2_X1 U14706 ( .A1(a_30_), .A2(n14523), .ZN(n14691) );
  AND3_X1 U14707 ( .A1(b_2_), .A2(b_3_), .A3(n7494), .ZN(n14410) );
  XNOR2_X1 U14708 ( .A(n14692), .B(n14693), .ZN(n14392) );
  NOR2_X1 U14709 ( .A1(n7545), .A2(n8055), .ZN(n14693) );
  XOR2_X1 U14710 ( .A(n14694), .B(n14695), .Z(n14692) );
  XOR2_X1 U14711 ( .A(n14696), .B(n14697), .Z(n14420) );
  NAND2_X1 U14712 ( .A1(n14698), .A2(n14699), .ZN(n14696) );
  XNOR2_X1 U14713 ( .A(n14700), .B(n14701), .ZN(n14428) );
  XOR2_X1 U14714 ( .A(n14702), .B(n14703), .Z(n14701) );
  NAND2_X1 U14715 ( .A1(b_2_), .A2(a_23_), .ZN(n14703) );
  XNOR2_X1 U14716 ( .A(n14704), .B(n14705), .ZN(n14436) );
  XNOR2_X1 U14717 ( .A(n14706), .B(n14707), .ZN(n14704) );
  NOR2_X1 U14718 ( .A1(n7665), .A2(n8055), .ZN(n14707) );
  XNOR2_X1 U14719 ( .A(n14708), .B(n14709), .ZN(n14444) );
  XOR2_X1 U14720 ( .A(n14710), .B(n14711), .Z(n14708) );
  NAND2_X1 U14721 ( .A1(b_2_), .A2(a_19_), .ZN(n14710) );
  XNOR2_X1 U14722 ( .A(n14712), .B(n14713), .ZN(n14452) );
  XNOR2_X1 U14723 ( .A(n14714), .B(n14715), .ZN(n14712) );
  XOR2_X1 U14724 ( .A(n14716), .B(n14717), .Z(n14460) );
  XOR2_X1 U14725 ( .A(n14718), .B(n14719), .Z(n14716) );
  XOR2_X1 U14726 ( .A(n14720), .B(n14721), .Z(n14468) );
  XOR2_X1 U14727 ( .A(n14722), .B(n14723), .Z(n14720) );
  XOR2_X1 U14728 ( .A(n14724), .B(n14725), .Z(n14476) );
  XOR2_X1 U14729 ( .A(n14726), .B(n14727), .Z(n14724) );
  XOR2_X1 U14730 ( .A(n14728), .B(n14729), .Z(n14484) );
  XOR2_X1 U14731 ( .A(n14730), .B(n14731), .Z(n14728) );
  XOR2_X1 U14732 ( .A(n14732), .B(n14733), .Z(n14492) );
  XOR2_X1 U14733 ( .A(n14734), .B(n14735), .Z(n14732) );
  XOR2_X1 U14734 ( .A(n14736), .B(n14737), .Z(n14496) );
  XOR2_X1 U14735 ( .A(n14738), .B(n14739), .Z(n14736) );
  INV_X1 U14736 ( .A(n7979), .ZN(n7928) );
  NAND2_X1 U14737 ( .A1(a_3_), .A2(b_3_), .ZN(n7979) );
  XOR2_X1 U14738 ( .A(n14740), .B(n14741), .Z(n14503) );
  XOR2_X1 U14739 ( .A(n14742), .B(n14743), .Z(n14740) );
  XNOR2_X1 U14740 ( .A(n14744), .B(n14745), .ZN(n14507) );
  XOR2_X1 U14741 ( .A(n14746), .B(n7949), .Z(n14745) );
  XOR2_X1 U14742 ( .A(n14747), .B(n14748), .Z(n14513) );
  XOR2_X1 U14743 ( .A(n14749), .B(n14750), .Z(n14747) );
  XOR2_X1 U14744 ( .A(n14526), .B(n14751), .Z(n14511) );
  XNOR2_X1 U14745 ( .A(n14524), .B(n14752), .ZN(n14751) );
  NAND2_X1 U14746 ( .A1(a_0_), .A2(b_2_), .ZN(n14752) );
  AND2_X1 U14747 ( .A1(n14753), .A2(n14754), .ZN(n14524) );
  NAND2_X1 U14748 ( .A1(n14749), .A2(n14755), .ZN(n14754) );
  OR2_X1 U14749 ( .A1(n14750), .A2(n14748), .ZN(n14755) );
  NOR2_X1 U14750 ( .A1(n8055), .A2(n7957), .ZN(n14749) );
  NAND2_X1 U14751 ( .A1(n14748), .A2(n14750), .ZN(n14753) );
  NAND2_X1 U14752 ( .A1(n14756), .A2(n14757), .ZN(n14750) );
  NAND2_X1 U14753 ( .A1(n14744), .A2(n14758), .ZN(n14757) );
  OR2_X1 U14754 ( .A1(n14746), .A2(n14759), .ZN(n14758) );
  XOR2_X1 U14755 ( .A(n14760), .B(n14761), .Z(n14744) );
  XNOR2_X1 U14756 ( .A(n14762), .B(n14763), .ZN(n14761) );
  NAND2_X1 U14757 ( .A1(b_1_), .A2(a_3_), .ZN(n14760) );
  NAND2_X1 U14758 ( .A1(n14759), .A2(n14746), .ZN(n14756) );
  NAND2_X1 U14759 ( .A1(n14764), .A2(n14765), .ZN(n14746) );
  NAND2_X1 U14760 ( .A1(n14742), .A2(n14766), .ZN(n14765) );
  OR2_X1 U14761 ( .A1(n14743), .A2(n14741), .ZN(n14766) );
  NOR2_X1 U14762 ( .A1(n8055), .A2(n7937), .ZN(n14742) );
  NAND2_X1 U14763 ( .A1(n14741), .A2(n14743), .ZN(n14764) );
  NAND2_X1 U14764 ( .A1(n14541), .A2(n14767), .ZN(n14743) );
  NAND2_X1 U14765 ( .A1(n14540), .A2(n14542), .ZN(n14767) );
  NAND2_X1 U14766 ( .A1(n14768), .A2(n14769), .ZN(n14542) );
  NAND2_X1 U14767 ( .A1(b_2_), .A2(a_4_), .ZN(n14769) );
  INV_X1 U14768 ( .A(n14770), .ZN(n14768) );
  XOR2_X1 U14769 ( .A(n14771), .B(n14772), .Z(n14540) );
  XNOR2_X1 U14770 ( .A(n14773), .B(n14774), .ZN(n14772) );
  NAND2_X1 U14771 ( .A1(b_1_), .A2(a_5_), .ZN(n14771) );
  NAND2_X1 U14772 ( .A1(a_4_), .A2(n14770), .ZN(n14541) );
  NAND2_X1 U14773 ( .A1(n14775), .A2(n14776), .ZN(n14770) );
  NAND2_X1 U14774 ( .A1(n14738), .A2(n14777), .ZN(n14776) );
  OR2_X1 U14775 ( .A1(n14739), .A2(n14737), .ZN(n14777) );
  NOR2_X1 U14776 ( .A1(n8055), .A2(n7908), .ZN(n14738) );
  NAND2_X1 U14777 ( .A1(n14737), .A2(n14739), .ZN(n14775) );
  NAND2_X1 U14778 ( .A1(n14552), .A2(n14778), .ZN(n14739) );
  NAND2_X1 U14779 ( .A1(n14551), .A2(n14553), .ZN(n14778) );
  NAND2_X1 U14780 ( .A1(n14779), .A2(n14780), .ZN(n14553) );
  NAND2_X1 U14781 ( .A1(b_2_), .A2(a_6_), .ZN(n14780) );
  INV_X1 U14782 ( .A(n14781), .ZN(n14779) );
  XOR2_X1 U14783 ( .A(n14782), .B(n14783), .Z(n14551) );
  XNOR2_X1 U14784 ( .A(n14784), .B(n14785), .ZN(n14783) );
  NAND2_X1 U14785 ( .A1(b_1_), .A2(a_7_), .ZN(n14782) );
  NAND2_X1 U14786 ( .A1(a_6_), .A2(n14781), .ZN(n14552) );
  NAND2_X1 U14787 ( .A1(n14786), .A2(n14787), .ZN(n14781) );
  NAND2_X1 U14788 ( .A1(n14734), .A2(n14788), .ZN(n14787) );
  OR2_X1 U14789 ( .A1(n14735), .A2(n14733), .ZN(n14788) );
  NOR2_X1 U14790 ( .A1(n8055), .A2(n7872), .ZN(n14734) );
  NAND2_X1 U14791 ( .A1(n14733), .A2(n14735), .ZN(n14786) );
  NAND2_X1 U14792 ( .A1(n14563), .A2(n14789), .ZN(n14735) );
  NAND2_X1 U14793 ( .A1(n14562), .A2(n14564), .ZN(n14789) );
  NAND2_X1 U14794 ( .A1(n14790), .A2(n14791), .ZN(n14564) );
  NAND2_X1 U14795 ( .A1(b_2_), .A2(a_8_), .ZN(n14791) );
  INV_X1 U14796 ( .A(n14792), .ZN(n14790) );
  XOR2_X1 U14797 ( .A(n14793), .B(n14794), .Z(n14562) );
  XNOR2_X1 U14798 ( .A(n14795), .B(n14796), .ZN(n14794) );
  NAND2_X1 U14799 ( .A1(b_1_), .A2(a_9_), .ZN(n14793) );
  NAND2_X1 U14800 ( .A1(a_8_), .A2(n14792), .ZN(n14563) );
  NAND2_X1 U14801 ( .A1(n14797), .A2(n14798), .ZN(n14792) );
  NAND2_X1 U14802 ( .A1(n14730), .A2(n14799), .ZN(n14798) );
  OR2_X1 U14803 ( .A1(n14731), .A2(n14729), .ZN(n14799) );
  NOR2_X1 U14804 ( .A1(n8055), .A2(n8052), .ZN(n14730) );
  NAND2_X1 U14805 ( .A1(n14729), .A2(n14731), .ZN(n14797) );
  NAND2_X1 U14806 ( .A1(n14574), .A2(n14800), .ZN(n14731) );
  NAND2_X1 U14807 ( .A1(n14573), .A2(n14575), .ZN(n14800) );
  NAND2_X1 U14808 ( .A1(n14801), .A2(n14802), .ZN(n14575) );
  NAND2_X1 U14809 ( .A1(b_2_), .A2(a_10_), .ZN(n14802) );
  INV_X1 U14810 ( .A(n14803), .ZN(n14801) );
  XOR2_X1 U14811 ( .A(n14804), .B(n14805), .Z(n14573) );
  XNOR2_X1 U14812 ( .A(n14806), .B(n14807), .ZN(n14805) );
  NAND2_X1 U14813 ( .A1(b_1_), .A2(a_11_), .ZN(n14804) );
  NAND2_X1 U14814 ( .A1(a_10_), .A2(n14803), .ZN(n14574) );
  NAND2_X1 U14815 ( .A1(n14808), .A2(n14809), .ZN(n14803) );
  NAND2_X1 U14816 ( .A1(n14726), .A2(n14810), .ZN(n14809) );
  OR2_X1 U14817 ( .A1(n14727), .A2(n14725), .ZN(n14810) );
  NOR2_X1 U14818 ( .A1(n8055), .A2(n7811), .ZN(n14726) );
  NAND2_X1 U14819 ( .A1(n14725), .A2(n14727), .ZN(n14808) );
  NAND2_X1 U14820 ( .A1(n14585), .A2(n14811), .ZN(n14727) );
  NAND2_X1 U14821 ( .A1(n14584), .A2(n14586), .ZN(n14811) );
  NAND2_X1 U14822 ( .A1(n14812), .A2(n14813), .ZN(n14586) );
  NAND2_X1 U14823 ( .A1(b_2_), .A2(a_12_), .ZN(n14813) );
  INV_X1 U14824 ( .A(n14814), .ZN(n14812) );
  XOR2_X1 U14825 ( .A(n14815), .B(n14816), .Z(n14584) );
  XNOR2_X1 U14826 ( .A(n14817), .B(n14818), .ZN(n14816) );
  NAND2_X1 U14827 ( .A1(b_1_), .A2(a_13_), .ZN(n14815) );
  NAND2_X1 U14828 ( .A1(a_12_), .A2(n14814), .ZN(n14585) );
  NAND2_X1 U14829 ( .A1(n14819), .A2(n14820), .ZN(n14814) );
  NAND2_X1 U14830 ( .A1(n14722), .A2(n14821), .ZN(n14820) );
  OR2_X1 U14831 ( .A1(n14723), .A2(n14721), .ZN(n14821) );
  NOR2_X1 U14832 ( .A1(n8055), .A2(n7789), .ZN(n14722) );
  NAND2_X1 U14833 ( .A1(n14721), .A2(n14723), .ZN(n14819) );
  NAND2_X1 U14834 ( .A1(n14596), .A2(n14822), .ZN(n14723) );
  NAND2_X1 U14835 ( .A1(n14595), .A2(n14597), .ZN(n14822) );
  NAND2_X1 U14836 ( .A1(n14823), .A2(n14824), .ZN(n14597) );
  NAND2_X1 U14837 ( .A1(b_2_), .A2(a_14_), .ZN(n14824) );
  INV_X1 U14838 ( .A(n14825), .ZN(n14823) );
  XOR2_X1 U14839 ( .A(n14826), .B(n14827), .Z(n14595) );
  XNOR2_X1 U14840 ( .A(n14828), .B(n14829), .ZN(n14827) );
  NAND2_X1 U14841 ( .A1(b_1_), .A2(a_15_), .ZN(n14826) );
  NAND2_X1 U14842 ( .A1(a_14_), .A2(n14825), .ZN(n14596) );
  NAND2_X1 U14843 ( .A1(n14830), .A2(n14831), .ZN(n14825) );
  NAND2_X1 U14844 ( .A1(n14718), .A2(n14832), .ZN(n14831) );
  OR2_X1 U14845 ( .A1(n14719), .A2(n14717), .ZN(n14832) );
  NOR2_X1 U14846 ( .A1(n8055), .A2(n7754), .ZN(n14718) );
  NAND2_X1 U14847 ( .A1(n14717), .A2(n14719), .ZN(n14830) );
  NAND2_X1 U14848 ( .A1(n14607), .A2(n14833), .ZN(n14719) );
  NAND2_X1 U14849 ( .A1(n14606), .A2(n14608), .ZN(n14833) );
  NAND2_X1 U14850 ( .A1(n14834), .A2(n14835), .ZN(n14608) );
  NAND2_X1 U14851 ( .A1(b_2_), .A2(a_16_), .ZN(n14835) );
  INV_X1 U14852 ( .A(n14836), .ZN(n14834) );
  XOR2_X1 U14853 ( .A(n14837), .B(n14838), .Z(n14606) );
  XNOR2_X1 U14854 ( .A(n14839), .B(n14840), .ZN(n14838) );
  NAND2_X1 U14855 ( .A1(b_1_), .A2(a_17_), .ZN(n14837) );
  NAND2_X1 U14856 ( .A1(a_16_), .A2(n14836), .ZN(n14607) );
  NAND2_X1 U14857 ( .A1(n14841), .A2(n14842), .ZN(n14836) );
  NAND2_X1 U14858 ( .A1(n14714), .A2(n14843), .ZN(n14842) );
  NAND2_X1 U14859 ( .A1(n14715), .A2(n14713), .ZN(n14843) );
  NOR2_X1 U14860 ( .A1(n8055), .A2(n7732), .ZN(n14714) );
  OR2_X1 U14861 ( .A1(n14713), .A2(n14715), .ZN(n14841) );
  AND2_X1 U14862 ( .A1(n14844), .A2(n14845), .ZN(n14715) );
  NAND2_X1 U14863 ( .A1(n14619), .A2(n14846), .ZN(n14845) );
  OR2_X1 U14864 ( .A1(n14618), .A2(n14616), .ZN(n14846) );
  NOR2_X1 U14865 ( .A1(n8055), .A2(n8047), .ZN(n14619) );
  NAND2_X1 U14866 ( .A1(n14616), .A2(n14618), .ZN(n14844) );
  NAND2_X1 U14867 ( .A1(n14847), .A2(n14848), .ZN(n14618) );
  NAND3_X1 U14868 ( .A1(a_19_), .A2(n14849), .A3(b_2_), .ZN(n14848) );
  NAND2_X1 U14869 ( .A1(n14711), .A2(n14709), .ZN(n14849) );
  OR2_X1 U14870 ( .A1(n14709), .A2(n14711), .ZN(n14847) );
  AND2_X1 U14871 ( .A1(n14850), .A2(n14851), .ZN(n14711) );
  NAND2_X1 U14872 ( .A1(n14630), .A2(n14852), .ZN(n14851) );
  OR2_X1 U14873 ( .A1(n14629), .A2(n14627), .ZN(n14852) );
  NOR2_X1 U14874 ( .A1(n8055), .A2(n8044), .ZN(n14630) );
  NAND2_X1 U14875 ( .A1(n14627), .A2(n14629), .ZN(n14850) );
  NAND2_X1 U14876 ( .A1(n14853), .A2(n14854), .ZN(n14629) );
  NAND3_X1 U14877 ( .A1(a_21_), .A2(n14855), .A3(b_2_), .ZN(n14854) );
  NAND2_X1 U14878 ( .A1(n14706), .A2(n14705), .ZN(n14855) );
  OR2_X1 U14879 ( .A1(n14705), .A2(n14706), .ZN(n14853) );
  AND2_X1 U14880 ( .A1(n14856), .A2(n14857), .ZN(n14706) );
  NAND2_X1 U14881 ( .A1(n14641), .A2(n14858), .ZN(n14857) );
  OR2_X1 U14882 ( .A1(n14640), .A2(n14638), .ZN(n14858) );
  NOR2_X1 U14883 ( .A1(n8055), .A2(n7650), .ZN(n14641) );
  NAND2_X1 U14884 ( .A1(n14638), .A2(n14640), .ZN(n14856) );
  NAND2_X1 U14885 ( .A1(n14859), .A2(n14860), .ZN(n14640) );
  NAND3_X1 U14886 ( .A1(a_23_), .A2(n14861), .A3(b_2_), .ZN(n14860) );
  OR2_X1 U14887 ( .A1(n14702), .A2(n14700), .ZN(n14861) );
  NAND2_X1 U14888 ( .A1(n14700), .A2(n14702), .ZN(n14859) );
  NAND2_X1 U14889 ( .A1(n14862), .A2(n14863), .ZN(n14702) );
  NAND2_X1 U14890 ( .A1(n14652), .A2(n14864), .ZN(n14863) );
  OR2_X1 U14891 ( .A1(n14651), .A2(n14649), .ZN(n14864) );
  NOR2_X1 U14892 ( .A1(n8055), .A2(n8041), .ZN(n14652) );
  NAND2_X1 U14893 ( .A1(n14649), .A2(n14651), .ZN(n14862) );
  NAND2_X1 U14894 ( .A1(n14698), .A2(n14865), .ZN(n14651) );
  NAND2_X1 U14895 ( .A1(n14697), .A2(n14699), .ZN(n14865) );
  NAND2_X1 U14896 ( .A1(n14866), .A2(n14867), .ZN(n14699) );
  NAND2_X1 U14897 ( .A1(b_2_), .A2(a_25_), .ZN(n14867) );
  INV_X1 U14898 ( .A(n14868), .ZN(n14866) );
  XOR2_X1 U14899 ( .A(n14869), .B(n14870), .Z(n14697) );
  NOR2_X1 U14900 ( .A1(n14522), .A2(n7580), .ZN(n14870) );
  XOR2_X1 U14901 ( .A(n14871), .B(n14872), .Z(n14869) );
  NAND2_X1 U14902 ( .A1(a_25_), .A2(n14868), .ZN(n14698) );
  NAND2_X1 U14903 ( .A1(n14873), .A2(n14874), .ZN(n14868) );
  NAND3_X1 U14904 ( .A1(a_26_), .A2(n14875), .A3(b_2_), .ZN(n14874) );
  NAND2_X1 U14905 ( .A1(n14663), .A2(n14661), .ZN(n14875) );
  OR2_X1 U14906 ( .A1(n14661), .A2(n14663), .ZN(n14873) );
  AND2_X1 U14907 ( .A1(n14876), .A2(n14877), .ZN(n14663) );
  NAND2_X1 U14908 ( .A1(n14671), .A2(n14878), .ZN(n14877) );
  OR2_X1 U14909 ( .A1(n14670), .A2(n14668), .ZN(n14878) );
  NOR2_X1 U14910 ( .A1(n8055), .A2(n7580), .ZN(n14671) );
  NAND2_X1 U14911 ( .A1(n14668), .A2(n14670), .ZN(n14876) );
  NAND2_X1 U14912 ( .A1(n14879), .A2(n14880), .ZN(n14670) );
  NAND3_X1 U14913 ( .A1(a_28_), .A2(n14881), .A3(b_2_), .ZN(n14880) );
  OR2_X1 U14914 ( .A1(n14677), .A2(n14679), .ZN(n14881) );
  NAND2_X1 U14915 ( .A1(n14677), .A2(n14679), .ZN(n14879) );
  NAND2_X1 U14916 ( .A1(n14882), .A2(n14883), .ZN(n14679) );
  NAND3_X1 U14917 ( .A1(a_29_), .A2(n14884), .A3(b_2_), .ZN(n14883) );
  OR2_X1 U14918 ( .A1(n14694), .A2(n14695), .ZN(n14884) );
  NAND2_X1 U14919 ( .A1(n14695), .A2(n14694), .ZN(n14882) );
  NAND2_X1 U14920 ( .A1(n14885), .A2(n14886), .ZN(n14694) );
  NAND2_X1 U14921 ( .A1(b_0_), .A2(n14887), .ZN(n14886) );
  NAND2_X1 U14922 ( .A1(n7527), .A2(n14888), .ZN(n14887) );
  NAND2_X1 U14923 ( .A1(a_31_), .A2(n14523), .ZN(n14888) );
  NAND2_X1 U14924 ( .A1(b_1_), .A2(n14889), .ZN(n14885) );
  NAND2_X1 U14925 ( .A1(n7531), .A2(n14890), .ZN(n14889) );
  NAND2_X1 U14926 ( .A1(a_30_), .A2(n14522), .ZN(n14890) );
  AND3_X1 U14927 ( .A1(b_2_), .A2(b_1_), .A3(n7494), .ZN(n14695) );
  XNOR2_X1 U14928 ( .A(n14891), .B(n14892), .ZN(n14677) );
  NOR2_X1 U14929 ( .A1(n14522), .A2(n7535), .ZN(n14892) );
  XOR2_X1 U14930 ( .A(n14893), .B(n14894), .Z(n14891) );
  XOR2_X1 U14931 ( .A(n14895), .B(n14896), .Z(n14668) );
  XNOR2_X1 U14932 ( .A(n14897), .B(n14898), .ZN(n14896) );
  NAND2_X1 U14933 ( .A1(a_29_), .A2(b_0_), .ZN(n14895) );
  XNOR2_X1 U14934 ( .A(n14899), .B(n14900), .ZN(n14661) );
  XNOR2_X1 U14935 ( .A(n14901), .B(n14902), .ZN(n14900) );
  NAND2_X1 U14936 ( .A1(a_28_), .A2(b_0_), .ZN(n14899) );
  XOR2_X1 U14937 ( .A(n14903), .B(n14904), .Z(n14649) );
  XNOR2_X1 U14938 ( .A(n14905), .B(n14906), .ZN(n14904) );
  NAND2_X1 U14939 ( .A1(a_26_), .A2(b_0_), .ZN(n14903) );
  XOR2_X1 U14940 ( .A(n14907), .B(n14908), .Z(n14700) );
  NOR2_X1 U14941 ( .A1(n14522), .A2(n8039), .ZN(n14908) );
  XOR2_X1 U14942 ( .A(n14909), .B(n14910), .Z(n14907) );
  XOR2_X1 U14943 ( .A(n14911), .B(n14912), .Z(n14638) );
  XNOR2_X1 U14944 ( .A(n14913), .B(n14914), .ZN(n14912) );
  NAND2_X1 U14945 ( .A1(a_24_), .A2(b_0_), .ZN(n14911) );
  XNOR2_X1 U14946 ( .A(n14915), .B(n14916), .ZN(n14705) );
  NOR2_X1 U14947 ( .A1(n14522), .A2(n8042), .ZN(n14916) );
  XOR2_X1 U14948 ( .A(n14917), .B(n14918), .Z(n14915) );
  XOR2_X1 U14949 ( .A(n14919), .B(n14920), .Z(n14627) );
  XNOR2_X1 U14950 ( .A(n14921), .B(n14922), .ZN(n14920) );
  NAND2_X1 U14951 ( .A1(a_22_), .A2(b_0_), .ZN(n14919) );
  XNOR2_X1 U14952 ( .A(n14923), .B(n14924), .ZN(n14709) );
  NOR2_X1 U14953 ( .A1(n14522), .A2(n7665), .ZN(n14924) );
  XOR2_X1 U14954 ( .A(n14925), .B(n14926), .Z(n14923) );
  XOR2_X1 U14955 ( .A(n14927), .B(n14928), .Z(n14616) );
  XNOR2_X1 U14956 ( .A(n14929), .B(n14930), .ZN(n14928) );
  NAND2_X1 U14957 ( .A1(a_20_), .A2(b_0_), .ZN(n14927) );
  XNOR2_X1 U14958 ( .A(n14931), .B(n14932), .ZN(n14713) );
  NOR2_X1 U14959 ( .A1(n14522), .A2(n8045), .ZN(n14932) );
  XOR2_X1 U14960 ( .A(n14933), .B(n14934), .Z(n14931) );
  XOR2_X1 U14961 ( .A(n14935), .B(n14936), .Z(n14717) );
  NOR2_X1 U14962 ( .A1(n8438), .A2(n14523), .ZN(n14936) );
  XOR2_X1 U14963 ( .A(n14937), .B(n14938), .Z(n14935) );
  XOR2_X1 U14964 ( .A(n14939), .B(n14940), .Z(n14721) );
  NOR2_X1 U14965 ( .A1(n8049), .A2(n14523), .ZN(n14940) );
  XOR2_X1 U14966 ( .A(n14941), .B(n14942), .Z(n14939) );
  XOR2_X1 U14967 ( .A(n14943), .B(n14944), .Z(n14725) );
  NOR2_X1 U14968 ( .A1(n8669), .A2(n14523), .ZN(n14944) );
  XOR2_X1 U14969 ( .A(n14945), .B(n14946), .Z(n14943) );
  XOR2_X1 U14970 ( .A(n14947), .B(n14948), .Z(n14729) );
  NOR2_X1 U14971 ( .A1(n8051), .A2(n14523), .ZN(n14948) );
  XOR2_X1 U14972 ( .A(n14949), .B(n14950), .Z(n14947) );
  XOR2_X1 U14973 ( .A(n14951), .B(n14952), .Z(n14733) );
  NOR2_X1 U14974 ( .A1(n8686), .A2(n14523), .ZN(n14952) );
  XOR2_X1 U14975 ( .A(n14953), .B(n14954), .Z(n14951) );
  XOR2_X1 U14976 ( .A(n14955), .B(n14956), .Z(n14737) );
  NOR2_X1 U14977 ( .A1(n7887), .A2(n14523), .ZN(n14956) );
  XOR2_X1 U14978 ( .A(n14957), .B(n14958), .Z(n14955) );
  XOR2_X1 U14979 ( .A(n14959), .B(n14960), .Z(n14741) );
  NOR2_X1 U14980 ( .A1(n7916), .A2(n14523), .ZN(n14960) );
  XOR2_X1 U14981 ( .A(n14961), .B(n14962), .Z(n14959) );
  INV_X1 U14982 ( .A(n7949), .ZN(n14759) );
  NAND2_X1 U14983 ( .A1(b_2_), .A2(a_2_), .ZN(n7949) );
  XOR2_X1 U14984 ( .A(n14963), .B(n14964), .Z(n14748) );
  XOR2_X1 U14985 ( .A(n14965), .B(n14966), .Z(n14963) );
  XNOR2_X1 U14986 ( .A(n14967), .B(n14968), .ZN(n14526) );
  AND2_X1 U14987 ( .A1(n7963), .A2(n14519), .ZN(n14968) );
  AND2_X1 U14988 ( .A1(n14969), .A2(n14970), .ZN(n14519) );
  NAND2_X1 U14989 ( .A1(n14964), .A2(n14971), .ZN(n14970) );
  OR2_X1 U14990 ( .A1(n14966), .A2(n14965), .ZN(n14971) );
  NOR2_X1 U14991 ( .A1(n14523), .A2(n8056), .ZN(n14964) );
  NAND2_X1 U14992 ( .A1(n14965), .A2(n14966), .ZN(n14969) );
  NAND2_X1 U14993 ( .A1(n14972), .A2(n14973), .ZN(n14966) );
  NAND3_X1 U14994 ( .A1(a_3_), .A2(n14974), .A3(b_1_), .ZN(n14973) );
  OR2_X1 U14995 ( .A1(n14763), .A2(n14762), .ZN(n14974) );
  NAND2_X1 U14996 ( .A1(n14762), .A2(n14763), .ZN(n14972) );
  NAND2_X1 U14997 ( .A1(n14975), .A2(n14976), .ZN(n14763) );
  NAND3_X1 U14998 ( .A1(a_4_), .A2(n14977), .A3(b_1_), .ZN(n14976) );
  OR2_X1 U14999 ( .A1(n14962), .A2(n14961), .ZN(n14977) );
  NAND2_X1 U15000 ( .A1(n14961), .A2(n14962), .ZN(n14975) );
  NAND2_X1 U15001 ( .A1(n14978), .A2(n14979), .ZN(n14962) );
  NAND3_X1 U15002 ( .A1(a_5_), .A2(n14980), .A3(b_1_), .ZN(n14979) );
  OR2_X1 U15003 ( .A1(n14774), .A2(n14773), .ZN(n14980) );
  NAND2_X1 U15004 ( .A1(n14773), .A2(n14774), .ZN(n14978) );
  NAND2_X1 U15005 ( .A1(n14981), .A2(n14982), .ZN(n14774) );
  NAND3_X1 U15006 ( .A1(a_6_), .A2(n14983), .A3(b_1_), .ZN(n14982) );
  OR2_X1 U15007 ( .A1(n14958), .A2(n14957), .ZN(n14983) );
  NAND2_X1 U15008 ( .A1(n14957), .A2(n14958), .ZN(n14981) );
  NAND2_X1 U15009 ( .A1(n14984), .A2(n14985), .ZN(n14958) );
  NAND3_X1 U15010 ( .A1(a_7_), .A2(n14986), .A3(b_1_), .ZN(n14985) );
  OR2_X1 U15011 ( .A1(n14785), .A2(n14784), .ZN(n14986) );
  NAND2_X1 U15012 ( .A1(n14784), .A2(n14785), .ZN(n14984) );
  NAND2_X1 U15013 ( .A1(n14987), .A2(n14988), .ZN(n14785) );
  NAND3_X1 U15014 ( .A1(a_8_), .A2(n14989), .A3(b_1_), .ZN(n14988) );
  OR2_X1 U15015 ( .A1(n14954), .A2(n14953), .ZN(n14989) );
  NAND2_X1 U15016 ( .A1(n14953), .A2(n14954), .ZN(n14987) );
  NAND2_X1 U15017 ( .A1(n14990), .A2(n14991), .ZN(n14954) );
  NAND3_X1 U15018 ( .A1(a_9_), .A2(n14992), .A3(b_1_), .ZN(n14991) );
  OR2_X1 U15019 ( .A1(n14796), .A2(n14795), .ZN(n14992) );
  NAND2_X1 U15020 ( .A1(n14795), .A2(n14796), .ZN(n14990) );
  NAND2_X1 U15021 ( .A1(n14993), .A2(n14994), .ZN(n14796) );
  NAND3_X1 U15022 ( .A1(a_10_), .A2(n14995), .A3(b_1_), .ZN(n14994) );
  OR2_X1 U15023 ( .A1(n14950), .A2(n14949), .ZN(n14995) );
  NAND2_X1 U15024 ( .A1(n14949), .A2(n14950), .ZN(n14993) );
  NAND2_X1 U15025 ( .A1(n14996), .A2(n14997), .ZN(n14950) );
  NAND3_X1 U15026 ( .A1(a_11_), .A2(n14998), .A3(b_1_), .ZN(n14997) );
  OR2_X1 U15027 ( .A1(n14807), .A2(n14806), .ZN(n14998) );
  NAND2_X1 U15028 ( .A1(n14806), .A2(n14807), .ZN(n14996) );
  NAND2_X1 U15029 ( .A1(n14999), .A2(n15000), .ZN(n14807) );
  NAND3_X1 U15030 ( .A1(a_12_), .A2(n15001), .A3(b_1_), .ZN(n15000) );
  OR2_X1 U15031 ( .A1(n14946), .A2(n14945), .ZN(n15001) );
  NAND2_X1 U15032 ( .A1(n14945), .A2(n14946), .ZN(n14999) );
  NAND2_X1 U15033 ( .A1(n15002), .A2(n15003), .ZN(n14946) );
  NAND3_X1 U15034 ( .A1(a_13_), .A2(n15004), .A3(b_1_), .ZN(n15003) );
  OR2_X1 U15035 ( .A1(n14818), .A2(n14817), .ZN(n15004) );
  NAND2_X1 U15036 ( .A1(n14817), .A2(n14818), .ZN(n15002) );
  NAND2_X1 U15037 ( .A1(n15005), .A2(n15006), .ZN(n14818) );
  NAND3_X1 U15038 ( .A1(a_14_), .A2(n15007), .A3(b_1_), .ZN(n15006) );
  OR2_X1 U15039 ( .A1(n14942), .A2(n14941), .ZN(n15007) );
  NAND2_X1 U15040 ( .A1(n14941), .A2(n14942), .ZN(n15005) );
  NAND2_X1 U15041 ( .A1(n15008), .A2(n15009), .ZN(n14942) );
  NAND3_X1 U15042 ( .A1(a_15_), .A2(n15010), .A3(b_1_), .ZN(n15009) );
  OR2_X1 U15043 ( .A1(n14829), .A2(n14828), .ZN(n15010) );
  NAND2_X1 U15044 ( .A1(n14828), .A2(n14829), .ZN(n15008) );
  NAND2_X1 U15045 ( .A1(n15011), .A2(n15012), .ZN(n14829) );
  NAND3_X1 U15046 ( .A1(a_16_), .A2(n15013), .A3(b_1_), .ZN(n15012) );
  OR2_X1 U15047 ( .A1(n14938), .A2(n14937), .ZN(n15013) );
  NAND2_X1 U15048 ( .A1(n14937), .A2(n14938), .ZN(n15011) );
  NAND2_X1 U15049 ( .A1(n15014), .A2(n15015), .ZN(n14938) );
  NAND3_X1 U15050 ( .A1(a_17_), .A2(n15016), .A3(b_1_), .ZN(n15015) );
  OR2_X1 U15051 ( .A1(n14840), .A2(n14839), .ZN(n15016) );
  NAND2_X1 U15052 ( .A1(n14839), .A2(n14840), .ZN(n15014) );
  NAND2_X1 U15053 ( .A1(n15017), .A2(n15018), .ZN(n14840) );
  NAND3_X1 U15054 ( .A1(b_0_), .A2(n15019), .A3(a_19_), .ZN(n15018) );
  OR2_X1 U15055 ( .A1(n14934), .A2(n14933), .ZN(n15019) );
  NAND2_X1 U15056 ( .A1(n14933), .A2(n14934), .ZN(n15017) );
  NAND2_X1 U15057 ( .A1(n15020), .A2(n15021), .ZN(n14934) );
  NAND3_X1 U15058 ( .A1(b_0_), .A2(n15022), .A3(a_20_), .ZN(n15021) );
  OR2_X1 U15059 ( .A1(n14930), .A2(n14929), .ZN(n15022) );
  NAND2_X1 U15060 ( .A1(n14929), .A2(n14930), .ZN(n15020) );
  NAND2_X1 U15061 ( .A1(n15023), .A2(n15024), .ZN(n14930) );
  NAND3_X1 U15062 ( .A1(b_0_), .A2(n15025), .A3(a_21_), .ZN(n15024) );
  NAND2_X1 U15063 ( .A1(n14926), .A2(n14925), .ZN(n15025) );
  INV_X1 U15064 ( .A(n15026), .ZN(n14926) );
  NAND2_X1 U15065 ( .A1(n15027), .A2(n15026), .ZN(n15023) );
  NAND2_X1 U15066 ( .A1(n15028), .A2(n15029), .ZN(n15026) );
  NAND3_X1 U15067 ( .A1(b_0_), .A2(n15030), .A3(a_22_), .ZN(n15029) );
  OR2_X1 U15068 ( .A1(n14922), .A2(n14921), .ZN(n15030) );
  NAND2_X1 U15069 ( .A1(n14921), .A2(n14922), .ZN(n15028) );
  NAND2_X1 U15070 ( .A1(n15031), .A2(n15032), .ZN(n14922) );
  NAND3_X1 U15071 ( .A1(b_0_), .A2(n15033), .A3(a_23_), .ZN(n15032) );
  NAND2_X1 U15072 ( .A1(n14918), .A2(n14917), .ZN(n15033) );
  INV_X1 U15073 ( .A(n15034), .ZN(n14918) );
  NAND2_X1 U15074 ( .A1(n15035), .A2(n15034), .ZN(n15031) );
  NAND2_X1 U15075 ( .A1(n15036), .A2(n15037), .ZN(n15034) );
  NAND3_X1 U15076 ( .A1(b_0_), .A2(n15038), .A3(a_24_), .ZN(n15037) );
  OR2_X1 U15077 ( .A1(n14914), .A2(n14913), .ZN(n15038) );
  NAND2_X1 U15078 ( .A1(n14913), .A2(n14914), .ZN(n15036) );
  NAND2_X1 U15079 ( .A1(n15039), .A2(n15040), .ZN(n14914) );
  NAND3_X1 U15080 ( .A1(b_0_), .A2(n15041), .A3(a_25_), .ZN(n15040) );
  NAND2_X1 U15081 ( .A1(n14910), .A2(n14909), .ZN(n15041) );
  INV_X1 U15082 ( .A(n15042), .ZN(n14910) );
  NAND2_X1 U15083 ( .A1(n15043), .A2(n15042), .ZN(n15039) );
  NAND2_X1 U15084 ( .A1(n15044), .A2(n15045), .ZN(n15042) );
  NAND3_X1 U15085 ( .A1(b_0_), .A2(n15046), .A3(a_26_), .ZN(n15045) );
  OR2_X1 U15086 ( .A1(n14906), .A2(n14905), .ZN(n15046) );
  NAND2_X1 U15087 ( .A1(n14905), .A2(n14906), .ZN(n15044) );
  NAND2_X1 U15088 ( .A1(n15047), .A2(n15048), .ZN(n14906) );
  NAND3_X1 U15089 ( .A1(b_0_), .A2(n15049), .A3(a_27_), .ZN(n15048) );
  NAND2_X1 U15090 ( .A1(n14872), .A2(n14871), .ZN(n15049) );
  INV_X1 U15091 ( .A(n15050), .ZN(n14872) );
  NAND2_X1 U15092 ( .A1(n15051), .A2(n15050), .ZN(n15047) );
  NAND2_X1 U15093 ( .A1(n15052), .A2(n15053), .ZN(n15050) );
  NAND3_X1 U15094 ( .A1(b_0_), .A2(n15054), .A3(a_28_), .ZN(n15053) );
  OR2_X1 U15095 ( .A1(n14902), .A2(n14901), .ZN(n15054) );
  NAND2_X1 U15096 ( .A1(n14901), .A2(n14902), .ZN(n15052) );
  NAND2_X1 U15097 ( .A1(n15055), .A2(n15056), .ZN(n14902) );
  NAND3_X1 U15098 ( .A1(b_0_), .A2(n15057), .A3(a_29_), .ZN(n15056) );
  OR2_X1 U15099 ( .A1(n14898), .A2(n14897), .ZN(n15057) );
  NAND2_X1 U15100 ( .A1(n14897), .A2(n14898), .ZN(n15055) );
  NAND2_X1 U15101 ( .A1(n14894), .A2(n15058), .ZN(n14898) );
  NAND3_X1 U15102 ( .A1(a_30_), .A2(b_0_), .A3(n14893), .ZN(n15058) );
  NOR2_X1 U15103 ( .A1(n14523), .A2(n7545), .ZN(n14893) );
  NAND3_X1 U15104 ( .A1(b_1_), .A2(b_0_), .A3(n7494), .ZN(n14894) );
  NOR2_X1 U15105 ( .A1(n14523), .A2(n7560), .ZN(n14897) );
  NOR2_X1 U15106 ( .A1(n14523), .A2(n7580), .ZN(n14901) );
  INV_X1 U15107 ( .A(n14871), .ZN(n15051) );
  NAND2_X1 U15108 ( .A1(b_1_), .A2(a_26_), .ZN(n14871) );
  NOR2_X1 U15109 ( .A1(n14523), .A2(n8039), .ZN(n14905) );
  INV_X1 U15110 ( .A(n14909), .ZN(n15043) );
  NAND2_X1 U15111 ( .A1(b_1_), .A2(a_24_), .ZN(n14909) );
  NOR2_X1 U15112 ( .A1(n14523), .A2(n8042), .ZN(n14913) );
  INV_X1 U15113 ( .A(n14917), .ZN(n15035) );
  NAND2_X1 U15114 ( .A1(b_1_), .A2(a_22_), .ZN(n14917) );
  NOR2_X1 U15115 ( .A1(n14523), .A2(n7665), .ZN(n14921) );
  INV_X1 U15116 ( .A(n14925), .ZN(n15027) );
  NAND2_X1 U15117 ( .A1(b_1_), .A2(a_20_), .ZN(n14925) );
  NOR2_X1 U15118 ( .A1(n14523), .A2(n8045), .ZN(n14929) );
  NOR2_X1 U15119 ( .A1(n14523), .A2(n8047), .ZN(n14933) );
  NOR2_X1 U15120 ( .A1(n8047), .A2(n14522), .ZN(n14839) );
  NOR2_X1 U15121 ( .A1(n7732), .A2(n14522), .ZN(n14937) );
  NOR2_X1 U15122 ( .A1(n8438), .A2(n14522), .ZN(n14828) );
  NOR2_X1 U15123 ( .A1(n7754), .A2(n14522), .ZN(n14941) );
  NOR2_X1 U15124 ( .A1(n8049), .A2(n14522), .ZN(n14817) );
  NOR2_X1 U15125 ( .A1(n7789), .A2(n14522), .ZN(n14945) );
  NOR2_X1 U15126 ( .A1(n8669), .A2(n14522), .ZN(n14806) );
  NOR2_X1 U15127 ( .A1(n7811), .A2(n14522), .ZN(n14949) );
  NOR2_X1 U15128 ( .A1(n8051), .A2(n14522), .ZN(n14795) );
  NOR2_X1 U15129 ( .A1(n8052), .A2(n14522), .ZN(n14953) );
  NOR2_X1 U15130 ( .A1(n8686), .A2(n14522), .ZN(n14784) );
  NOR2_X1 U15131 ( .A1(n7872), .A2(n14522), .ZN(n14957) );
  NOR2_X1 U15132 ( .A1(n7887), .A2(n14522), .ZN(n14773) );
  NOR2_X1 U15133 ( .A1(n7908), .A2(n14522), .ZN(n14961) );
  NOR2_X1 U15134 ( .A1(n7916), .A2(n14522), .ZN(n14762) );
  NOR2_X1 U15135 ( .A1(n7937), .A2(n14522), .ZN(n14965) );
  NOR2_X1 U15136 ( .A1(n14523), .A2(n7957), .ZN(n7963) );
  NAND2_X1 U15137 ( .A1(a_2_), .A2(b_0_), .ZN(n14967) );
  NAND2_X1 U15138 ( .A1(n15061), .A2(n7976), .ZN(n15060) );
  NAND2_X1 U15139 ( .A1(b_0_), .A2(n8942), .ZN(n7976) );
  INV_X1 U15140 ( .A(a_0_), .ZN(n8942) );
  NAND2_X1 U15141 ( .A1(n15062), .A2(n15063), .ZN(n15061) );
  NAND2_X1 U15142 ( .A1(a_1_), .A2(n14523), .ZN(n15063) );
  INV_X1 U15143 ( .A(b_1_), .ZN(n14523) );
  NAND3_X1 U15144 ( .A1(n15064), .A2(n15065), .A3(n15066), .ZN(n15062) );
  NAND2_X1 U15145 ( .A1(b_2_), .A2(n8056), .ZN(n15066) );
  INV_X1 U15146 ( .A(a_2_), .ZN(n8056) );
  NAND3_X1 U15147 ( .A1(n15067), .A2(n15068), .A3(n15069), .ZN(n15065) );
  NAND2_X1 U15148 ( .A1(a_3_), .A2(n7930), .ZN(n15069) );
  INV_X1 U15149 ( .A(b_3_), .ZN(n7930) );
  NAND3_X1 U15150 ( .A1(n15070), .A2(n15071), .A3(n15072), .ZN(n15068) );
  NAND2_X1 U15151 ( .A1(b_4_), .A2(n7916), .ZN(n15072) );
  INV_X1 U15152 ( .A(a_4_), .ZN(n7916) );
  NAND3_X1 U15153 ( .A1(n15073), .A2(n15074), .A3(n15075), .ZN(n15071) );
  NAND2_X1 U15154 ( .A1(a_5_), .A2(n7901), .ZN(n15075) );
  NAND3_X1 U15155 ( .A1(n15076), .A2(n15077), .A3(n15078), .ZN(n15074) );
  NAND2_X1 U15156 ( .A1(b_6_), .A2(n7887), .ZN(n15078) );
  INV_X1 U15157 ( .A(a_6_), .ZN(n7887) );
  NAND3_X1 U15158 ( .A1(n15079), .A2(n15080), .A3(n15081), .ZN(n15077) );
  NAND2_X1 U15159 ( .A1(a_7_), .A2(n7874), .ZN(n15081) );
  NAND3_X1 U15160 ( .A1(n15082), .A2(n15083), .A3(n15084), .ZN(n15080) );
  NAND2_X1 U15161 ( .A1(b_8_), .A2(n8686), .ZN(n15084) );
  INV_X1 U15162 ( .A(a_8_), .ZN(n8686) );
  NAND3_X1 U15163 ( .A1(n15085), .A2(n15086), .A3(n15087), .ZN(n15083) );
  NAND2_X1 U15164 ( .A1(a_9_), .A2(n7839), .ZN(n15087) );
  INV_X1 U15165 ( .A(b_9_), .ZN(n7839) );
  NAND3_X1 U15166 ( .A1(n15088), .A2(n15089), .A3(n15090), .ZN(n15086) );
  NAND2_X1 U15167 ( .A1(b_9_), .A2(n8052), .ZN(n15090) );
  INV_X1 U15168 ( .A(a_9_), .ZN(n8052) );
  NAND3_X1 U15169 ( .A1(n15091), .A2(n15092), .A3(n15093), .ZN(n15089) );
  NAND2_X1 U15170 ( .A1(a_11_), .A2(n7813), .ZN(n15093) );
  INV_X1 U15171 ( .A(b_11_), .ZN(n7813) );
  NAND3_X1 U15172 ( .A1(n15094), .A2(n15095), .A3(n15096), .ZN(n15092) );
  NAND2_X1 U15173 ( .A1(b_12_), .A2(n8669), .ZN(n15096) );
  INV_X1 U15174 ( .A(a_12_), .ZN(n8669) );
  NAND3_X1 U15175 ( .A1(n15097), .A2(n15098), .A3(n15099), .ZN(n15095) );
  NAND2_X1 U15176 ( .A1(a_13_), .A2(n7782), .ZN(n15099) );
  INV_X1 U15177 ( .A(b_13_), .ZN(n7782) );
  NAND3_X1 U15178 ( .A1(n15100), .A2(n15101), .A3(n15102), .ZN(n15098) );
  NAND2_X1 U15179 ( .A1(b_14_), .A2(n8049), .ZN(n15102) );
  INV_X1 U15180 ( .A(a_14_), .ZN(n8049) );
  NAND3_X1 U15181 ( .A1(n15103), .A2(n15104), .A3(n15105), .ZN(n15101) );
  NAND2_X1 U15182 ( .A1(a_15_), .A2(n7756), .ZN(n15105) );
  INV_X1 U15183 ( .A(b_15_), .ZN(n7756) );
  NAND3_X1 U15184 ( .A1(n15106), .A2(n15107), .A3(n15108), .ZN(n15104) );
  NAND2_X1 U15185 ( .A1(b_16_), .A2(n8438), .ZN(n15108) );
  INV_X1 U15186 ( .A(a_16_), .ZN(n8438) );
  NAND3_X1 U15187 ( .A1(n15109), .A2(n15110), .A3(n15111), .ZN(n15107) );
  NAND2_X1 U15188 ( .A1(a_17_), .A2(n7725), .ZN(n15111) );
  INV_X1 U15189 ( .A(b_17_), .ZN(n7725) );
  NAND3_X1 U15190 ( .A1(n15112), .A2(n15113), .A3(n15114), .ZN(n15110) );
  NAND2_X1 U15191 ( .A1(b_18_), .A2(n8047), .ZN(n15114) );
  NAND3_X1 U15192 ( .A1(n15115), .A2(n15116), .A3(n15117), .ZN(n15113) );
  NAND2_X1 U15193 ( .A1(a_19_), .A2(n7693), .ZN(n15117) );
  INV_X1 U15194 ( .A(b_19_), .ZN(n7693) );
  NAND3_X1 U15195 ( .A1(n15118), .A2(n15119), .A3(n15120), .ZN(n15116) );
  NAND2_X1 U15196 ( .A1(b_20_), .A2(n8044), .ZN(n15120) );
  NAND3_X1 U15197 ( .A1(n15121), .A2(n15122), .A3(n15123), .ZN(n15119) );
  NAND2_X1 U15198 ( .A1(a_21_), .A2(n7667), .ZN(n15123) );
  INV_X1 U15199 ( .A(b_21_), .ZN(n7667) );
  NAND3_X1 U15200 ( .A1(n15124), .A2(n15125), .A3(n15126), .ZN(n15122) );
  NAND2_X1 U15201 ( .A1(b_22_), .A2(n7650), .ZN(n15126) );
  INV_X1 U15202 ( .A(a_22_), .ZN(n7650) );
  NAND3_X1 U15203 ( .A1(n15127), .A2(n15128), .A3(n15129), .ZN(n15125) );
  NAND2_X1 U15204 ( .A1(a_23_), .A2(n7636), .ZN(n15129) );
  INV_X1 U15205 ( .A(b_23_), .ZN(n7636) );
  NAND3_X1 U15206 ( .A1(n15130), .A2(n15131), .A3(n15132), .ZN(n15128) );
  NAND2_X1 U15207 ( .A1(b_24_), .A2(n8041), .ZN(n15132) );
  NAND3_X1 U15208 ( .A1(n15133), .A2(n15134), .A3(n15135), .ZN(n15131) );
  NAND2_X1 U15209 ( .A1(a_25_), .A2(n7609), .ZN(n15135) );
  NAND3_X1 U15210 ( .A1(n15136), .A2(n15137), .A3(n15138), .ZN(n15134) );
  NAND2_X1 U15211 ( .A1(b_26_), .A2(n7595), .ZN(n15138) );
  INV_X1 U15212 ( .A(a_26_), .ZN(n7595) );
  NAND3_X1 U15213 ( .A1(n15139), .A2(n15140), .A3(n15141), .ZN(n15137) );
  NAND2_X1 U15214 ( .A1(a_27_), .A2(n7582), .ZN(n15141) );
  NAND3_X1 U15215 ( .A1(n15142), .A2(n15143), .A3(n15144), .ZN(n15140) );
  NAND2_X1 U15216 ( .A1(b_28_), .A2(n7560), .ZN(n15144) );
  INV_X1 U15217 ( .A(a_28_), .ZN(n7560) );
  NAND3_X1 U15218 ( .A1(n15145), .A2(n15146), .A3(n15147), .ZN(n15143) );
  NAND2_X1 U15219 ( .A1(a_29_), .A2(n7547), .ZN(n15147) );
  INV_X1 U15220 ( .A(b_29_), .ZN(n7547) );
  NAND4_X1 U15221 ( .A1(n15148), .A2(n15149), .A3(n15150), .A4(n15151), .ZN(
        n15146) );
  NAND2_X1 U15222 ( .A1(b_31_), .A2(n7532), .ZN(n15151) );
  NAND2_X1 U15223 ( .A1(a_30_), .A2(n8359), .ZN(n7532) );
  OR2_X1 U15224 ( .A1(n8359), .A2(n7494), .ZN(n15150) );
  INV_X1 U15225 ( .A(b_30_), .ZN(n8359) );
  NAND2_X1 U15226 ( .A1(b_29_), .A2(n7545), .ZN(n15149) );
  NAND2_X1 U15227 ( .A1(n7535), .A2(n8036), .ZN(n15148) );
  INV_X1 U15228 ( .A(a_31_), .ZN(n8036) );
  INV_X1 U15229 ( .A(a_30_), .ZN(n7535) );
  NAND2_X1 U15230 ( .A1(a_28_), .A2(n8037), .ZN(n15145) );
  INV_X1 U15231 ( .A(b_28_), .ZN(n8037) );
  NAND2_X1 U15232 ( .A1(b_27_), .A2(n7580), .ZN(n15142) );
  INV_X1 U15233 ( .A(a_27_), .ZN(n7580) );
  NAND2_X1 U15234 ( .A1(a_26_), .A2(n8038), .ZN(n15139) );
  INV_X1 U15235 ( .A(b_26_), .ZN(n8038) );
  NAND2_X1 U15236 ( .A1(b_25_), .A2(n8039), .ZN(n15136) );
  NAND2_X1 U15237 ( .A1(a_24_), .A2(n8040), .ZN(n15133) );
  INV_X1 U15238 ( .A(b_24_), .ZN(n8040) );
  NAND2_X1 U15239 ( .A1(b_23_), .A2(n8042), .ZN(n15130) );
  NAND2_X1 U15240 ( .A1(a_22_), .A2(n9968), .ZN(n15127) );
  NAND2_X1 U15241 ( .A1(b_21_), .A2(n7665), .ZN(n15124) );
  NAND2_X1 U15242 ( .A1(a_20_), .A2(n8043), .ZN(n15121) );
  INV_X1 U15243 ( .A(b_20_), .ZN(n8043) );
  NAND2_X1 U15244 ( .A1(b_19_), .A2(n8045), .ZN(n15118) );
  INV_X1 U15245 ( .A(a_19_), .ZN(n8045) );
  NAND2_X1 U15246 ( .A1(a_18_), .A2(n8046), .ZN(n15115) );
  INV_X1 U15247 ( .A(b_18_), .ZN(n8046) );
  NAND2_X1 U15248 ( .A1(b_17_), .A2(n7732), .ZN(n15112) );
  NAND2_X1 U15249 ( .A1(a_16_), .A2(n11315), .ZN(n15109) );
  NAND2_X1 U15250 ( .A1(b_15_), .A2(n7754), .ZN(n15106) );
  INV_X1 U15251 ( .A(a_15_), .ZN(n7754) );
  NAND2_X1 U15252 ( .A1(a_14_), .A2(n8048), .ZN(n15103) );
  INV_X1 U15253 ( .A(b_14_), .ZN(n8048) );
  NAND2_X1 U15254 ( .A1(b_13_), .A2(n7789), .ZN(n15100) );
  INV_X1 U15255 ( .A(a_13_), .ZN(n7789) );
  NAND2_X1 U15256 ( .A1(a_12_), .A2(n12188), .ZN(n15097) );
  INV_X1 U15257 ( .A(b_12_), .ZN(n12188) );
  NAND2_X1 U15258 ( .A1(b_11_), .A2(n7811), .ZN(n15094) );
  INV_X1 U15259 ( .A(a_11_), .ZN(n7811) );
  NAND2_X1 U15260 ( .A1(a_10_), .A2(n8050), .ZN(n15091) );
  INV_X1 U15261 ( .A(b_10_), .ZN(n8050) );
  NAND2_X1 U15262 ( .A1(b_10_), .A2(n8051), .ZN(n15088) );
  INV_X1 U15263 ( .A(a_10_), .ZN(n8051) );
  NAND2_X1 U15264 ( .A1(a_8_), .A2(n13086), .ZN(n15085) );
  INV_X1 U15265 ( .A(b_8_), .ZN(n13086) );
  NAND2_X1 U15266 ( .A1(b_7_), .A2(n7872), .ZN(n15082) );
  INV_X1 U15267 ( .A(a_7_), .ZN(n7872) );
  NAND2_X1 U15268 ( .A1(a_6_), .A2(n8053), .ZN(n15079) );
  INV_X1 U15269 ( .A(b_6_), .ZN(n8053) );
  NAND2_X1 U15270 ( .A1(b_5_), .A2(n7908), .ZN(n15076) );
  INV_X1 U15271 ( .A(a_5_), .ZN(n7908) );
  NAND2_X1 U15272 ( .A1(a_4_), .A2(n8054), .ZN(n15073) );
  NAND2_X1 U15273 ( .A1(b_3_), .A2(n7937), .ZN(n15070) );
  INV_X1 U15274 ( .A(a_3_), .ZN(n7937) );
  NAND2_X1 U15275 ( .A1(a_2_), .A2(n8055), .ZN(n15067) );
  INV_X1 U15276 ( .A(b_2_), .ZN(n8055) );
  NAND2_X1 U15277 ( .A1(b_1_), .A2(n7957), .ZN(n15064) );
  NAND2_X1 U15278 ( .A1(a_0_), .A2(n14522), .ZN(n15059) );
  INV_X1 U15279 ( .A(b_0_), .ZN(n14522) );
endmodule

