module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n798_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n481_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n796_, new_n350_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n429_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1020_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n917_, new_n426_, new_n1036_, new_n398_, new_n646_, new_n395_, new_n538_, new_n383_, new_n854_, new_n541_, new_n458_, new_n1026_, new_n447_, new_n473_, new_n790_, new_n1081_, new_n587_, new_n783_, new_n739_, new_n969_, new_n835_, new_n996_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n628_, new_n409_, new_n745_, new_n457_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n1002_, new_n834_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n998_, new_n1056_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n499_, new_n533_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n597_, new_n978_, new_n408_, new_n470_, new_n1072_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n681_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n377_, new_n539_, new_n905_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n780_, new_n984_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n877_, new_n348_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1023_, new_n951_, new_n709_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n647_, new_n889_, new_n536_, new_n464_, new_n573_, new_n765_, new_n405_;

and g000 ( N388, N29, N42, N75 );
and g001 ( N389, N29, N36, N80 );
nand g002 ( new_n345_, N29, N36, N42 );
not g003 ( N390, new_n345_ );
and g004 ( N391, N85, N86 );
not g005 ( new_n348_, N1 );
not g006 ( new_n349_, N8 );
not g007 ( new_n350_, N13 );
not g008 ( new_n351_, N17 );
nor g009 ( N418, new_n348_, new_n349_, new_n350_, new_n351_ );
nand g010 ( new_n353_, N1, N13, N17, N26 );
nor g011 ( new_n354_, N390, new_n353_ );
xor g012 ( N419, new_n354_, keyIn_0_8 );
nand g013 ( N420, N59, N75, N80 );
nand g014 ( N421, N36, N59, N80 );
nand g015 ( N422, N36, N42, N59 );
not g016 ( new_n359_, N90 );
nor g017 ( new_n360_, N87, N88 );
nor g018 ( N423, new_n360_, new_n359_ );
nor g019 ( new_n362_, new_n353_, new_n345_ );
xor g020 ( N446, new_n362_, keyIn_0_25 );
not g021 ( new_n364_, keyIn_0_0 );
nand g022 ( new_n365_, new_n364_, N1, N26, N51 );
nand g023 ( new_n366_, N1, N26, N51 );
nand g024 ( new_n367_, new_n366_, keyIn_0_0 );
nand g025 ( new_n368_, new_n367_, new_n365_ );
not g026 ( N447, new_n368_ );
not g027 ( new_n370_, N55 );
nor g028 ( new_n371_, new_n348_, new_n349_, new_n350_, new_n370_ );
nand g029 ( new_n372_, new_n371_, N29, N68 );
xnor g030 ( N448, new_n372_, keyIn_0_12 );
and g031 ( new_n374_, N59, N68 );
nand g032 ( new_n375_, new_n371_, N74, new_n374_ );
xnor g033 ( N449, new_n375_, keyIn_0_13 );
not g034 ( new_n377_, N89 );
nor g035 ( N450, new_n360_, new_n377_ );
xor g036 ( new_n379_, N101, N106 );
xnor g037 ( new_n380_, new_n379_, keyIn_0_16 );
xor g038 ( new_n381_, new_n380_, keyIn_0_29 );
xnor g039 ( new_n382_, N91, N96 );
xnor g040 ( new_n383_, new_n382_, keyIn_0_15 );
xor g041 ( new_n384_, new_n383_, keyIn_0_28 );
nand g042 ( new_n385_, new_n381_, new_n384_ );
or g043 ( new_n386_, new_n385_, keyIn_0_42 );
nand g044 ( new_n387_, new_n385_, keyIn_0_42 );
nand g045 ( new_n388_, new_n380_, new_n383_ );
xnor g046 ( new_n389_, new_n388_, keyIn_0_30 );
nand g047 ( new_n390_, new_n386_, new_n387_, new_n389_ );
xnor g048 ( new_n391_, new_n390_, keyIn_0_52 );
nor g049 ( new_n392_, new_n391_, N130 );
xor g050 ( new_n393_, new_n392_, keyIn_0_71 );
nand g051 ( new_n394_, new_n391_, N130 );
xor g052 ( new_n395_, new_n394_, keyIn_0_70 );
nand g053 ( new_n396_, new_n393_, new_n395_ );
xnor g054 ( new_n397_, new_n396_, keyIn_0_94 );
xor g055 ( new_n398_, N111, N116 );
xnor g056 ( new_n399_, new_n398_, keyIn_0_17 );
xor g057 ( new_n400_, new_n399_, keyIn_0_31 );
xnor g058 ( new_n401_, N121, N126 );
xnor g059 ( new_n402_, new_n401_, keyIn_0_18 );
xor g060 ( new_n403_, new_n402_, keyIn_0_32 );
nand g061 ( new_n404_, new_n400_, new_n403_ );
xor g062 ( new_n405_, new_n404_, keyIn_0_43 );
nand g063 ( new_n406_, new_n399_, new_n402_ );
xor g064 ( new_n407_, new_n406_, keyIn_0_33 );
nand g065 ( new_n408_, new_n405_, new_n407_ );
xor g066 ( new_n409_, new_n408_, keyIn_0_53 );
nor g067 ( new_n410_, new_n409_, N135 );
xor g068 ( new_n411_, new_n410_, keyIn_0_73 );
nand g069 ( new_n412_, new_n409_, N135 );
xnor g070 ( new_n413_, new_n412_, keyIn_0_72 );
nand g071 ( new_n414_, new_n411_, new_n413_ );
xor g072 ( new_n415_, new_n414_, keyIn_0_95 );
nand g073 ( new_n416_, new_n415_, new_n397_ );
xor g074 ( new_n417_, new_n416_, keyIn_0_106 );
nor g075 ( new_n418_, new_n415_, new_n397_ );
xor g076 ( new_n419_, new_n418_, keyIn_0_116 );
nand g077 ( new_n420_, new_n419_, new_n417_ );
xnor g078 ( N767, new_n420_, keyIn_0_139 );
xnor g079 ( new_n422_, N171, N177 );
xnor g080 ( new_n423_, new_n422_, keyIn_0_22 );
xor g081 ( new_n424_, new_n423_, keyIn_0_36 );
xor g082 ( new_n425_, N159, N165 );
xnor g083 ( new_n426_, new_n425_, keyIn_0_21 );
xor g084 ( new_n427_, new_n426_, keyIn_0_35 );
nand g085 ( new_n428_, new_n427_, new_n424_ );
xnor g086 ( new_n429_, new_n428_, keyIn_0_49 );
nand g087 ( new_n430_, new_n426_, new_n423_ );
xor g088 ( new_n431_, new_n430_, keyIn_0_37 );
nand g089 ( new_n432_, new_n429_, new_n431_ );
xnor g090 ( new_n433_, new_n432_, keyIn_0_68 );
nor g091 ( new_n434_, new_n433_, N130 );
xor g092 ( new_n435_, new_n434_, keyIn_0_91 );
nand g093 ( new_n436_, new_n433_, N130 );
xnor g094 ( new_n437_, new_n436_, keyIn_0_90 );
nand g095 ( new_n438_, new_n435_, new_n437_ );
xor g096 ( new_n439_, new_n438_, keyIn_0_104 );
not g097 ( new_n440_, N207 );
xor g098 ( new_n441_, N195, N201 );
xnor g099 ( new_n442_, new_n441_, keyIn_0_24 );
xnor g100 ( new_n443_, new_n442_, keyIn_0_39 );
xor g101 ( new_n444_, N183, N189 );
xnor g102 ( new_n445_, new_n444_, keyIn_0_23 );
xnor g103 ( new_n446_, new_n445_, keyIn_0_38 );
nand g104 ( new_n447_, new_n443_, new_n446_ );
or g105 ( new_n448_, new_n447_, keyIn_0_50 );
nand g106 ( new_n449_, new_n447_, keyIn_0_50 );
nand g107 ( new_n450_, new_n442_, new_n445_ );
xnor g108 ( new_n451_, new_n450_, keyIn_0_40 );
nand g109 ( new_n452_, new_n448_, new_n449_, new_n451_ );
xor g110 ( new_n453_, new_n452_, keyIn_0_69 );
nor g111 ( new_n454_, new_n453_, new_n440_ );
xor g112 ( new_n455_, new_n454_, keyIn_0_92 );
nand g113 ( new_n456_, new_n453_, new_n440_ );
xor g114 ( new_n457_, new_n456_, keyIn_0_93 );
nand g115 ( new_n458_, new_n455_, new_n457_ );
xnor g116 ( new_n459_, new_n458_, keyIn_0_105 );
nor g117 ( new_n460_, new_n439_, new_n459_ );
xor g118 ( new_n461_, new_n460_, keyIn_0_115 );
nand g119 ( new_n462_, new_n439_, new_n459_ );
xnor g120 ( new_n463_, new_n462_, keyIn_0_117 );
nand g121 ( new_n464_, new_n461_, new_n463_ );
xnor g122 ( N768, new_n464_, keyIn_0_140 );
not g123 ( new_n466_, keyIn_0_137 );
not g124 ( new_n467_, keyIn_0_103 );
not g125 ( new_n468_, keyIn_0_63 );
not g126 ( new_n469_, keyIn_0_26 );
nand g127 ( new_n470_, new_n368_, keyIn_0_9 );
not g128 ( new_n471_, keyIn_0_9 );
nand g129 ( new_n472_, new_n367_, new_n471_, new_n365_ );
nand g130 ( new_n473_, new_n470_, new_n472_ );
nand g131 ( new_n474_, new_n473_, new_n469_ );
nand g132 ( new_n475_, new_n470_, keyIn_0_26, new_n472_ );
nand g133 ( new_n476_, new_n474_, new_n475_ );
nand g134 ( new_n477_, N59, N156 );
xnor g135 ( new_n478_, new_n477_, keyIn_0_5 );
nand g136 ( new_n479_, new_n476_, N17, new_n478_ );
nand g137 ( new_n480_, new_n479_, keyIn_0_48 );
not g138 ( new_n481_, keyIn_0_48 );
nand g139 ( new_n482_, new_n476_, new_n481_, N17, new_n478_ );
nand g140 ( new_n483_, new_n480_, new_n482_ );
nand g141 ( new_n484_, new_n483_, N1 );
nand g142 ( new_n485_, new_n484_, new_n468_ );
nand g143 ( new_n486_, new_n483_, keyIn_0_63, N1 );
nand g144 ( new_n487_, new_n485_, new_n486_ );
nand g145 ( new_n488_, new_n487_, N153 );
nand g146 ( new_n489_, new_n488_, keyIn_0_88 );
not g147 ( new_n490_, keyIn_0_88 );
nand g148 ( new_n491_, new_n487_, new_n490_, N153 );
nand g149 ( new_n492_, new_n489_, new_n491_ );
not g150 ( new_n493_, keyIn_0_47 );
not g151 ( new_n494_, keyIn_0_20 );
nor g152 ( new_n495_, N17, N42 );
xor g153 ( new_n496_, new_n495_, keyIn_0_6 );
nand g154 ( new_n497_, N17, N42 );
xor g155 ( new_n498_, new_n497_, keyIn_0_7 );
nand g156 ( new_n499_, new_n496_, new_n498_ );
nor g157 ( new_n500_, new_n499_, new_n494_ );
and g158 ( new_n501_, new_n499_, new_n494_ );
nor g159 ( new_n502_, new_n501_, new_n500_, new_n477_ );
nand g160 ( new_n503_, new_n502_, new_n493_, new_n476_ );
not g161 ( new_n504_, keyIn_0_1 );
nand g162 ( new_n505_, N1, N8, N17, N51 );
xnor g163 ( new_n506_, new_n505_, new_n504_ );
xnor g164 ( new_n507_, new_n506_, keyIn_0_10 );
nand g165 ( new_n508_, N42, N59, N75 );
xor g166 ( new_n509_, new_n508_, keyIn_0_3 );
xnor g167 ( new_n510_, new_n509_, keyIn_0_14 );
nand g168 ( new_n511_, new_n510_, new_n507_ );
xnor g169 ( new_n512_, new_n511_, keyIn_0_34 );
nand g170 ( new_n513_, new_n502_, new_n476_ );
nand g171 ( new_n514_, new_n513_, keyIn_0_47 );
nand g172 ( new_n515_, new_n514_, new_n512_, new_n503_ );
nand g173 ( new_n516_, new_n515_, keyIn_0_54 );
not g174 ( new_n517_, keyIn_0_54 );
nand g175 ( new_n518_, new_n514_, new_n512_, new_n517_, new_n503_ );
nand g176 ( new_n519_, new_n516_, keyIn_0_89, N126, new_n518_ );
not g177 ( new_n520_, keyIn_0_89 );
nand g178 ( new_n521_, new_n516_, N126, new_n518_ );
nand g179 ( new_n522_, new_n521_, new_n520_ );
nand g180 ( new_n523_, new_n522_, new_n519_ );
nand g181 ( new_n524_, new_n492_, new_n523_ );
nand g182 ( new_n525_, new_n524_, new_n467_ );
nand g183 ( new_n526_, new_n492_, keyIn_0_103, new_n523_ );
nand g184 ( new_n527_, N29, N75, N80 );
xor g185 ( new_n528_, new_n527_, keyIn_0_2 );
nand g186 ( new_n529_, new_n476_, new_n528_ );
nor g187 ( new_n530_, new_n529_, new_n370_ );
not g188 ( new_n531_, new_n530_ );
or g189 ( new_n532_, new_n531_, keyIn_0_46 );
nand g190 ( new_n533_, new_n531_, keyIn_0_46 );
xor g191 ( new_n534_, keyIn_0_4, N268 );
xor g192 ( new_n535_, new_n534_, keyIn_0_19 );
nand g193 ( new_n536_, new_n532_, new_n533_, new_n535_ );
xnor g194 ( new_n537_, new_n536_, keyIn_0_67 );
nand g195 ( new_n538_, new_n525_, new_n526_, new_n537_ );
nand g196 ( new_n539_, new_n538_, keyIn_0_114 );
not g197 ( new_n540_, keyIn_0_114 );
nand g198 ( new_n541_, new_n525_, new_n540_, new_n526_, new_n537_ );
nand g199 ( new_n542_, new_n539_, new_n466_, N201, new_n541_ );
nand g200 ( new_n543_, new_n539_, N201, new_n541_ );
nand g201 ( new_n544_, new_n543_, keyIn_0_137 );
nand g202 ( new_n545_, new_n544_, new_n542_ );
not g203 ( new_n546_, keyIn_0_138 );
not g204 ( new_n547_, N201 );
nand g205 ( new_n548_, new_n539_, new_n541_ );
nand g206 ( new_n549_, new_n548_, new_n546_, new_n547_ );
nand g207 ( new_n550_, new_n548_, new_n547_ );
nand g208 ( new_n551_, new_n550_, keyIn_0_138 );
nand g209 ( new_n552_, new_n545_, new_n549_, new_n551_ );
xor g210 ( new_n553_, new_n552_, keyIn_0_163 );
nor g211 ( new_n554_, new_n553_, N261 );
xor g212 ( new_n555_, new_n554_, keyIn_0_184 );
nand g213 ( new_n556_, new_n553_, N261 );
xor g214 ( new_n557_, new_n556_, keyIn_0_185 );
and g215 ( new_n558_, new_n555_, new_n557_ );
or g216 ( new_n559_, new_n558_, keyIn_0_202 );
nand g217 ( new_n560_, new_n558_, keyIn_0_202 );
nand g218 ( new_n561_, new_n559_, N219, new_n560_ );
xnor g219 ( new_n562_, new_n561_, keyIn_0_210 );
nand g220 ( new_n563_, N121, N210 );
nand g221 ( new_n564_, new_n562_, new_n563_ );
or g222 ( new_n565_, new_n564_, keyIn_0_216 );
nand g223 ( new_n566_, new_n564_, keyIn_0_216 );
nand g224 ( new_n567_, new_n553_, N228 );
nand g225 ( new_n568_, new_n544_, keyIn_0_162, new_n542_ );
not g226 ( new_n569_, keyIn_0_162 );
nand g227 ( new_n570_, new_n545_, new_n569_ );
nand g228 ( new_n571_, new_n570_, new_n568_ );
nand g229 ( new_n572_, new_n571_, N237 );
and g230 ( new_n573_, new_n567_, new_n572_ );
and g231 ( new_n574_, new_n573_, keyIn_0_203 );
nor g232 ( new_n575_, new_n573_, keyIn_0_203 );
nand g233 ( new_n576_, new_n539_, N246, new_n541_ );
nand g234 ( new_n577_, N255, N267 );
nand g235 ( new_n578_, new_n576_, new_n577_ );
xor g236 ( new_n579_, new_n578_, keyIn_0_164 );
nand g237 ( new_n580_, new_n371_, N42, N72, new_n374_ );
xor g238 ( new_n581_, new_n580_, keyIn_0_11 );
nand g239 ( new_n582_, new_n581_, N73 );
xnor g240 ( new_n583_, new_n582_, keyIn_0_27 );
xnor g241 ( new_n584_, new_n583_, keyIn_0_41 );
xnor g242 ( new_n585_, new_n584_, keyIn_0_51 );
and g243 ( new_n586_, new_n585_, N201 );
nor g244 ( new_n587_, new_n574_, new_n575_, new_n579_, new_n586_ );
nand g245 ( new_n588_, new_n565_, new_n566_, new_n587_ );
xnor g246 ( N850, new_n588_, keyIn_0_222 );
not g247 ( new_n590_, keyIn_0_196 );
not g248 ( new_n591_, keyIn_0_187 );
not g249 ( new_n592_, N189 );
not g250 ( new_n593_, keyIn_0_101 );
not g251 ( new_n594_, keyIn_0_84 );
nand g252 ( new_n595_, new_n487_, new_n594_, N146 );
nand g253 ( new_n596_, new_n487_, N146 );
nand g254 ( new_n597_, new_n596_, keyIn_0_84 );
nand g255 ( new_n598_, new_n597_, new_n595_ );
not g256 ( new_n599_, keyIn_0_85 );
nand g257 ( new_n600_, new_n516_, N116, new_n518_ );
nand g258 ( new_n601_, new_n600_, new_n599_ );
nand g259 ( new_n602_, new_n516_, keyIn_0_85, N116, new_n518_ );
nand g260 ( new_n603_, new_n601_, new_n602_ );
nand g261 ( new_n604_, new_n598_, new_n593_, new_n603_ );
nand g262 ( new_n605_, new_n598_, new_n603_ );
nand g263 ( new_n606_, new_n605_, keyIn_0_101 );
xnor g264 ( new_n607_, new_n536_, keyIn_0_65 );
nand g265 ( new_n608_, new_n606_, keyIn_0_112, new_n604_, new_n607_ );
not g266 ( new_n609_, keyIn_0_112 );
nand g267 ( new_n610_, new_n606_, new_n604_, new_n607_ );
nand g268 ( new_n611_, new_n610_, new_n609_ );
nand g269 ( new_n612_, new_n611_, keyIn_0_134, new_n592_, new_n608_ );
not g270 ( new_n613_, keyIn_0_134 );
nand g271 ( new_n614_, new_n611_, new_n592_, new_n608_ );
nand g272 ( new_n615_, new_n614_, new_n613_ );
and g273 ( new_n616_, new_n615_, new_n612_ );
not g274 ( new_n617_, keyIn_0_159 );
not g275 ( new_n618_, keyIn_0_113 );
not g276 ( new_n619_, keyIn_0_102 );
not g277 ( new_n620_, keyIn_0_86 );
nand g278 ( new_n621_, new_n487_, N149 );
nand g279 ( new_n622_, new_n621_, new_n620_ );
nand g280 ( new_n623_, new_n487_, keyIn_0_86, N149 );
nand g281 ( new_n624_, new_n622_, new_n623_ );
nand g282 ( new_n625_, new_n516_, keyIn_0_87, N121, new_n518_ );
not g283 ( new_n626_, keyIn_0_87 );
nand g284 ( new_n627_, new_n516_, N121, new_n518_ );
nand g285 ( new_n628_, new_n627_, new_n626_ );
nand g286 ( new_n629_, new_n628_, new_n625_ );
nand g287 ( new_n630_, new_n624_, new_n629_ );
nand g288 ( new_n631_, new_n630_, new_n619_ );
nand g289 ( new_n632_, new_n624_, keyIn_0_102, new_n629_ );
xnor g290 ( new_n633_, new_n536_, keyIn_0_66 );
nand g291 ( new_n634_, new_n631_, new_n632_, new_n633_ );
nand g292 ( new_n635_, new_n634_, new_n618_ );
nand g293 ( new_n636_, new_n631_, keyIn_0_113, new_n632_, new_n633_ );
nand g294 ( new_n637_, new_n635_, new_n636_ );
nand g295 ( new_n638_, new_n637_, N195 );
nand g296 ( new_n639_, new_n638_, keyIn_0_135 );
not g297 ( new_n640_, keyIn_0_135 );
nand g298 ( new_n641_, new_n637_, new_n640_, N195 );
nand g299 ( new_n642_, new_n639_, new_n641_ );
nand g300 ( new_n643_, new_n642_, new_n617_ );
nand g301 ( new_n644_, new_n639_, keyIn_0_159, new_n641_ );
nand g302 ( new_n645_, new_n643_, new_n644_ );
nand g303 ( new_n646_, new_n645_, new_n616_ );
nand g304 ( new_n647_, new_n646_, new_n591_ );
nand g305 ( new_n648_, new_n645_, keyIn_0_187, new_n616_ );
nand g306 ( new_n649_, new_n647_, new_n648_ );
nand g307 ( new_n650_, new_n551_, N261, new_n549_ );
not g308 ( new_n651_, N195 );
nand g309 ( new_n652_, new_n635_, keyIn_0_136, new_n651_, new_n636_ );
not g310 ( new_n653_, keyIn_0_136 );
nand g311 ( new_n654_, new_n635_, new_n651_, new_n636_ );
nand g312 ( new_n655_, new_n654_, new_n653_ );
nand g313 ( new_n656_, new_n615_, new_n655_, new_n612_, new_n652_ );
nor g314 ( new_n657_, new_n650_, new_n656_ );
nor g315 ( new_n658_, new_n657_, keyIn_0_167 );
not g316 ( new_n659_, keyIn_0_167 );
nor g317 ( new_n660_, new_n650_, new_n656_, new_n659_ );
nor g318 ( new_n661_, new_n658_, new_n660_ );
not g319 ( new_n662_, new_n656_ );
nand g320 ( new_n663_, new_n571_, new_n662_ );
and g321 ( new_n664_, new_n663_, keyIn_0_188 );
nor g322 ( new_n665_, new_n661_, new_n664_ );
not g323 ( new_n666_, keyIn_0_156 );
not g324 ( new_n667_, keyIn_0_133 );
nand g325 ( new_n668_, new_n611_, new_n608_ );
nand g326 ( new_n669_, new_n668_, N189 );
nand g327 ( new_n670_, new_n669_, new_n667_ );
nand g328 ( new_n671_, new_n668_, keyIn_0_133, N189 );
nand g329 ( new_n672_, new_n670_, new_n671_ );
nand g330 ( new_n673_, new_n672_, new_n666_ );
nand g331 ( new_n674_, new_n670_, keyIn_0_156, new_n671_ );
nand g332 ( new_n675_, new_n673_, new_n674_ );
nand g333 ( new_n676_, new_n675_, keyIn_0_177 );
not g334 ( new_n677_, keyIn_0_177 );
nand g335 ( new_n678_, new_n673_, new_n677_, new_n674_ );
nand g336 ( new_n679_, new_n676_, new_n678_ );
or g337 ( new_n680_, new_n663_, keyIn_0_188 );
nand g338 ( new_n681_, new_n665_, new_n649_, new_n679_, new_n680_ );
nand g339 ( new_n682_, new_n681_, new_n590_ );
and g340 ( new_n683_, new_n680_, new_n679_ );
nand g341 ( new_n684_, new_n683_, keyIn_0_196, new_n665_, new_n649_ );
nand g342 ( new_n685_, new_n682_, new_n684_ );
nand g343 ( new_n686_, new_n487_, N143 );
xor g344 ( new_n687_, new_n686_, keyIn_0_82 );
and g345 ( new_n688_, new_n516_, new_n518_ );
nand g346 ( new_n689_, new_n688_, N111 );
xor g347 ( new_n690_, new_n689_, keyIn_0_83 );
nand g348 ( new_n691_, new_n690_, new_n687_ );
xor g349 ( new_n692_, new_n691_, keyIn_0_100 );
xnor g350 ( new_n693_, new_n536_, keyIn_0_64 );
nand g351 ( new_n694_, new_n692_, new_n693_ );
xnor g352 ( new_n695_, new_n694_, keyIn_0_111 );
nor g353 ( new_n696_, new_n695_, N183 );
xnor g354 ( new_n697_, new_n696_, keyIn_0_131 );
nand g355 ( new_n698_, new_n695_, N183 );
xnor g356 ( new_n699_, new_n698_, keyIn_0_130 );
nand g357 ( new_n700_, new_n697_, new_n699_ );
xnor g358 ( new_n701_, new_n700_, keyIn_0_154 );
nand g359 ( new_n702_, new_n701_, new_n685_ );
xnor g360 ( new_n703_, new_n702_, keyIn_0_204 );
nor g361 ( new_n704_, new_n701_, new_n685_ );
xnor g362 ( new_n705_, new_n704_, keyIn_0_205 );
nand g363 ( new_n706_, new_n705_, new_n703_ );
xnor g364 ( new_n707_, new_n706_, keyIn_0_213 );
nand g365 ( new_n708_, new_n707_, N219 );
xnor g366 ( new_n709_, new_n708_, keyIn_0_219 );
nand g367 ( new_n710_, N106, N210 );
nand g368 ( new_n711_, new_n709_, new_n710_ );
or g369 ( new_n712_, new_n711_, keyIn_0_230 );
nand g370 ( new_n713_, new_n711_, keyIn_0_230 );
not g371 ( new_n714_, new_n701_ );
nand g372 ( new_n715_, new_n714_, N228 );
xnor g373 ( new_n716_, new_n715_, keyIn_0_175 );
not g374 ( new_n717_, keyIn_0_153 );
xnor g375 ( new_n718_, new_n699_, new_n717_ );
nand g376 ( new_n719_, new_n718_, N237 );
xnor g377 ( new_n720_, new_n719_, keyIn_0_176 );
and g378 ( new_n721_, new_n716_, new_n720_ );
nor g379 ( new_n722_, new_n721_, keyIn_0_197 );
and g380 ( new_n723_, new_n721_, keyIn_0_197 );
and g381 ( new_n724_, new_n695_, N246 );
or g382 ( new_n725_, new_n724_, keyIn_0_132 );
nand g383 ( new_n726_, new_n724_, keyIn_0_132 );
nand g384 ( new_n727_, new_n585_, N183 );
nand g385 ( new_n728_, new_n725_, new_n726_, new_n727_ );
xnor g386 ( new_n729_, new_n728_, keyIn_0_155 );
nor g387 ( new_n730_, new_n723_, new_n722_, new_n729_ );
nand g388 ( new_n731_, new_n712_, new_n713_, new_n730_ );
xor g389 ( N863, new_n731_, keyIn_0_240 );
nand g390 ( new_n733_, new_n655_, new_n652_ );
not g391 ( new_n734_, new_n733_ );
nand g392 ( new_n735_, new_n571_, new_n734_ );
xor g393 ( new_n736_, new_n735_, keyIn_0_186 );
xor g394 ( new_n737_, new_n645_, keyIn_0_180 );
nor g395 ( new_n738_, new_n650_, new_n733_ );
xnor g396 ( new_n739_, new_n738_, keyIn_0_166 );
nand g397 ( new_n740_, new_n736_, new_n737_, new_n739_ );
xor g398 ( new_n741_, new_n740_, keyIn_0_198 );
nand g399 ( new_n742_, new_n672_, new_n616_ );
xnor g400 ( new_n743_, new_n742_, keyIn_0_157 );
nor g401 ( new_n744_, new_n741_, new_n743_ );
xnor g402 ( new_n745_, new_n744_, keyIn_0_206 );
nand g403 ( new_n746_, new_n741_, new_n743_ );
xnor g404 ( new_n747_, new_n746_, keyIn_0_207 );
nand g405 ( new_n748_, new_n745_, new_n747_ );
xor g406 ( new_n749_, new_n748_, keyIn_0_214 );
nand g407 ( new_n750_, new_n749_, N219 );
xnor g408 ( new_n751_, new_n750_, keyIn_0_220 );
nand g409 ( new_n752_, N111, N210 );
nand g410 ( new_n753_, new_n751_, new_n752_ );
or g411 ( new_n754_, new_n753_, keyIn_0_231 );
nand g412 ( new_n755_, new_n753_, keyIn_0_231 );
nand g413 ( new_n756_, new_n743_, N228 );
xor g414 ( new_n757_, new_n756_, keyIn_0_178 );
not g415 ( new_n758_, N237 );
nor g416 ( new_n759_, new_n675_, new_n758_ );
xnor g417 ( new_n760_, new_n759_, keyIn_0_179 );
nand g418 ( new_n761_, new_n757_, new_n760_ );
xor g419 ( new_n762_, new_n761_, keyIn_0_199 );
nand g420 ( new_n763_, new_n668_, N246 );
nand g421 ( new_n764_, N255, N259 );
nand g422 ( new_n765_, new_n763_, new_n764_ );
nor g423 ( new_n766_, new_n765_, keyIn_0_158 );
and g424 ( new_n767_, new_n765_, keyIn_0_158 );
and g425 ( new_n768_, new_n585_, N189 );
nor g426 ( new_n769_, new_n762_, new_n766_, new_n767_, new_n768_ );
nand g427 ( new_n770_, new_n754_, new_n755_, new_n769_ );
xor g428 ( N864, new_n770_, keyIn_0_241 );
xnor g429 ( new_n772_, new_n571_, keyIn_0_183 );
xnor g430 ( new_n773_, new_n650_, keyIn_0_165 );
nand g431 ( new_n774_, new_n772_, new_n773_ );
xnor g432 ( new_n775_, new_n774_, keyIn_0_200 );
nand g433 ( new_n776_, new_n734_, new_n642_ );
xor g434 ( new_n777_, new_n776_, keyIn_0_160 );
not g435 ( new_n778_, new_n777_ );
nand g436 ( new_n779_, new_n775_, new_n778_ );
xor g437 ( new_n780_, new_n779_, keyIn_0_208 );
nor g438 ( new_n781_, new_n775_, new_n778_ );
xnor g439 ( new_n782_, new_n781_, keyIn_0_209 );
and g440 ( new_n783_, new_n780_, new_n782_ );
or g441 ( new_n784_, new_n783_, keyIn_0_215 );
nand g442 ( new_n785_, new_n783_, keyIn_0_215 );
nand g443 ( new_n786_, new_n784_, N219, new_n785_ );
xor g444 ( new_n787_, new_n786_, keyIn_0_221 );
nand g445 ( new_n788_, N116, N210 );
nand g446 ( new_n789_, new_n787_, new_n788_ );
xnor g447 ( new_n790_, new_n789_, keyIn_0_232 );
nand g448 ( new_n791_, new_n777_, N228 );
xor g449 ( new_n792_, new_n791_, keyIn_0_181 );
nand g450 ( new_n793_, new_n645_, N237 );
xor g451 ( new_n794_, new_n793_, keyIn_0_182 );
nand g452 ( new_n795_, new_n792_, new_n794_ );
xnor g453 ( new_n796_, new_n795_, keyIn_0_201 );
nand g454 ( new_n797_, new_n637_, N246 );
nand g455 ( new_n798_, N255, N260 );
nand g456 ( new_n799_, new_n797_, new_n798_ );
nor g457 ( new_n800_, new_n799_, keyIn_0_161 );
and g458 ( new_n801_, new_n799_, keyIn_0_161 );
and g459 ( new_n802_, new_n585_, N195 );
nor g460 ( new_n803_, new_n801_, new_n800_, new_n802_ );
nand g461 ( new_n804_, new_n790_, new_n796_, new_n803_ );
xor g462 ( N865, new_n804_, keyIn_0_242 );
not g463 ( new_n806_, keyIn_0_225 );
not g464 ( new_n807_, keyIn_0_211 );
nand g465 ( new_n808_, new_n682_, new_n807_, new_n684_, new_n697_ );
nand g466 ( new_n809_, new_n682_, new_n684_, new_n697_ );
nand g467 ( new_n810_, new_n809_, keyIn_0_211 );
nand g468 ( new_n811_, new_n810_, new_n808_ );
not g469 ( new_n812_, keyIn_0_174 );
xnor g470 ( new_n813_, new_n718_, new_n812_ );
nand g471 ( new_n814_, new_n811_, keyIn_0_212, new_n813_ );
not g472 ( new_n815_, keyIn_0_212 );
nand g473 ( new_n816_, new_n811_, new_n813_ );
nand g474 ( new_n817_, new_n816_, new_n815_ );
nand g475 ( new_n818_, new_n688_, N96 );
xor g476 ( new_n819_, new_n818_, keyIn_0_76 );
nand g477 ( new_n820_, N51, N138 );
nand g478 ( new_n821_, new_n819_, new_n820_ );
xor g479 ( new_n822_, new_n821_, keyIn_0_97 );
nor g480 ( new_n823_, new_n529_, new_n351_ );
not g481 ( new_n824_, new_n823_ );
or g482 ( new_n825_, new_n824_, keyIn_0_45 );
nand g483 ( new_n826_, new_n824_, keyIn_0_45 );
nand g484 ( new_n827_, new_n825_, new_n534_, new_n826_ );
xor g485 ( new_n828_, new_n827_, keyIn_0_58 );
nand g486 ( new_n829_, new_n476_, N55, new_n478_ );
xor g487 ( new_n830_, new_n829_, keyIn_0_44 );
nand g488 ( new_n831_, new_n830_, N146 );
xor g489 ( new_n832_, new_n831_, keyIn_0_57 );
nand g490 ( new_n833_, new_n828_, new_n832_ );
xor g491 ( new_n834_, new_n833_, keyIn_0_77 );
nand g492 ( new_n835_, new_n822_, new_n834_ );
xnor g493 ( new_n836_, new_n835_, keyIn_0_108 );
nor g494 ( new_n837_, new_n836_, N165 );
xor g495 ( new_n838_, new_n837_, keyIn_0_122 );
not g496 ( new_n839_, N171 );
nand g497 ( new_n840_, new_n688_, N101 );
xor g498 ( new_n841_, new_n840_, keyIn_0_78 );
nand g499 ( new_n842_, N17, N138 );
nand g500 ( new_n843_, new_n841_, new_n842_ );
xnor g501 ( new_n844_, new_n843_, keyIn_0_98 );
xor g502 ( new_n845_, new_n827_, keyIn_0_60 );
nand g503 ( new_n846_, new_n830_, N149 );
xnor g504 ( new_n847_, new_n846_, keyIn_0_59 );
nand g505 ( new_n848_, new_n845_, new_n847_ );
xor g506 ( new_n849_, new_n848_, keyIn_0_79 );
nand g507 ( new_n850_, new_n844_, new_n849_ );
xnor g508 ( new_n851_, new_n850_, keyIn_0_109 );
nand g509 ( new_n852_, new_n851_, new_n839_ );
xor g510 ( new_n853_, new_n852_, keyIn_0_125 );
not g511 ( new_n854_, keyIn_0_99 );
nand g512 ( new_n855_, new_n688_, N106 );
or g513 ( new_n856_, new_n855_, keyIn_0_80 );
nand g514 ( new_n857_, new_n855_, keyIn_0_80 );
nand g515 ( new_n858_, N138, N152 );
nand g516 ( new_n859_, new_n856_, new_n857_, new_n858_ );
nand g517 ( new_n860_, new_n859_, new_n854_ );
xor g518 ( new_n861_, new_n827_, keyIn_0_62 );
nand g519 ( new_n862_, new_n830_, N153 );
xnor g520 ( new_n863_, new_n862_, keyIn_0_61 );
nand g521 ( new_n864_, new_n861_, new_n863_ );
xnor g522 ( new_n865_, new_n864_, keyIn_0_81 );
or g523 ( new_n866_, new_n859_, new_n854_ );
nand g524 ( new_n867_, new_n866_, new_n865_, new_n860_ );
xnor g525 ( new_n868_, new_n867_, keyIn_0_110 );
or g526 ( new_n869_, new_n868_, N177 );
xor g527 ( new_n870_, new_n869_, keyIn_0_128 );
and g528 ( new_n871_, new_n838_, new_n853_, new_n870_ );
nand g529 ( new_n872_, new_n817_, new_n806_, new_n814_, new_n871_ );
nand g530 ( new_n873_, new_n817_, new_n814_, new_n871_ );
nand g531 ( new_n874_, new_n873_, keyIn_0_225 );
nand g532 ( new_n875_, new_n868_, N177 );
xor g533 ( new_n876_, new_n875_, keyIn_0_127 );
xor g534 ( new_n877_, new_n876_, keyIn_0_150 );
nand g535 ( new_n878_, new_n877_, new_n838_, new_n853_ );
xor g536 ( new_n879_, new_n878_, keyIn_0_191 );
nor g537 ( new_n880_, new_n851_, new_n839_ );
xnor g538 ( new_n881_, new_n880_, keyIn_0_124 );
xnor g539 ( new_n882_, new_n881_, keyIn_0_147 );
and g540 ( new_n883_, new_n882_, new_n838_ );
and g541 ( new_n884_, new_n883_, keyIn_0_190 );
nor g542 ( new_n885_, new_n883_, keyIn_0_190 );
nand g543 ( new_n886_, new_n836_, N165 );
xnor g544 ( new_n887_, new_n886_, keyIn_0_121 );
xor g545 ( new_n888_, new_n887_, keyIn_0_144 );
xnor g546 ( new_n889_, new_n888_, keyIn_0_168 );
nor g547 ( new_n890_, new_n879_, new_n889_, new_n884_, new_n885_ );
nand g548 ( new_n891_, new_n874_, keyIn_0_226, new_n872_, new_n890_ );
not g549 ( new_n892_, keyIn_0_226 );
nand g550 ( new_n893_, new_n874_, new_n872_, new_n890_ );
nand g551 ( new_n894_, new_n893_, new_n892_ );
nand g552 ( new_n895_, new_n894_, new_n891_ );
nand g553 ( new_n896_, new_n688_, N91 );
xor g554 ( new_n897_, new_n896_, keyIn_0_74 );
nand g555 ( new_n898_, N8, N138 );
nand g556 ( new_n899_, new_n897_, new_n898_ );
or g557 ( new_n900_, new_n899_, keyIn_0_96 );
nand g558 ( new_n901_, new_n899_, keyIn_0_96 );
xor g559 ( new_n902_, new_n827_, keyIn_0_56 );
nand g560 ( new_n903_, new_n830_, N143 );
xor g561 ( new_n904_, new_n903_, keyIn_0_55 );
nand g562 ( new_n905_, new_n902_, new_n904_ );
xor g563 ( new_n906_, new_n905_, keyIn_0_75 );
nand g564 ( new_n907_, new_n900_, new_n901_, new_n906_ );
xnor g565 ( new_n908_, new_n907_, keyIn_0_107 );
nor g566 ( new_n909_, new_n908_, N159 );
xnor g567 ( new_n910_, new_n909_, keyIn_0_119 );
nand g568 ( new_n911_, new_n895_, new_n910_ );
or g569 ( new_n912_, new_n911_, keyIn_0_243 );
nand g570 ( new_n913_, new_n911_, keyIn_0_243 );
nand g571 ( new_n914_, new_n908_, N159 );
xnor g572 ( new_n915_, new_n914_, keyIn_0_118 );
xor g573 ( new_n916_, new_n915_, keyIn_0_141 );
nand g574 ( new_n917_, new_n912_, new_n913_, new_n916_ );
xor g575 ( N866, new_n917_, keyIn_0_248 );
nand g576 ( new_n919_, new_n817_, new_n814_ );
nand g577 ( new_n920_, new_n870_, new_n876_ );
xnor g578 ( new_n921_, new_n920_, keyIn_0_151 );
not g579 ( new_n922_, new_n921_ );
nand g580 ( new_n923_, new_n919_, new_n922_ );
xnor g581 ( new_n924_, new_n923_, keyIn_0_217 );
nand g582 ( new_n925_, new_n817_, new_n814_, new_n921_ );
xnor g583 ( new_n926_, new_n925_, keyIn_0_218 );
nand g584 ( new_n927_, new_n924_, new_n926_ );
or g585 ( new_n928_, new_n927_, keyIn_0_229 );
nand g586 ( new_n929_, new_n927_, keyIn_0_229 );
nand g587 ( new_n930_, new_n928_, N219, new_n929_ );
xnor g588 ( new_n931_, new_n930_, keyIn_0_239 );
nand g589 ( new_n932_, N101, N210 );
nand g590 ( new_n933_, new_n931_, new_n932_ );
xor g591 ( new_n934_, new_n933_, keyIn_0_247 );
nand g592 ( new_n935_, new_n921_, N228 );
xnor g593 ( new_n936_, new_n935_, keyIn_0_172 );
nand g594 ( new_n937_, new_n877_, N237 );
xor g595 ( new_n938_, new_n937_, keyIn_0_173 );
nand g596 ( new_n939_, new_n936_, new_n938_ );
nor g597 ( new_n940_, new_n939_, keyIn_0_195 );
and g598 ( new_n941_, new_n939_, keyIn_0_195 );
nand g599 ( new_n942_, new_n868_, N246 );
or g600 ( new_n943_, new_n942_, keyIn_0_129 );
nand g601 ( new_n944_, new_n942_, keyIn_0_129 );
nand g602 ( new_n945_, new_n585_, N177 );
nand g603 ( new_n946_, new_n943_, new_n944_, new_n945_ );
xor g604 ( new_n947_, new_n946_, keyIn_0_152 );
nor g605 ( new_n948_, new_n941_, new_n940_, new_n947_ );
nand g606 ( new_n949_, new_n934_, new_n948_ );
nand g607 ( new_n950_, new_n949_, keyIn_0_249 );
not g608 ( new_n951_, keyIn_0_249 );
nand g609 ( new_n952_, new_n934_, new_n951_, new_n948_ );
nand g610 ( N874, new_n950_, new_n952_ );
not g611 ( new_n954_, keyIn_0_253 );
not g612 ( new_n955_, keyIn_0_250 );
nand g613 ( new_n956_, new_n910_, new_n915_ );
xor g614 ( new_n957_, new_n956_, keyIn_0_142 );
nand g615 ( new_n958_, new_n895_, new_n957_ );
xnor g616 ( new_n959_, new_n958_, keyIn_0_234 );
not g617 ( new_n960_, new_n957_ );
nand g618 ( new_n961_, new_n894_, new_n891_, new_n960_ );
xnor g619 ( new_n962_, new_n961_, keyIn_0_233 );
nand g620 ( new_n963_, new_n959_, new_n962_, keyIn_0_244 );
not g621 ( new_n964_, keyIn_0_244 );
nand g622 ( new_n965_, new_n959_, new_n962_ );
nand g623 ( new_n966_, new_n965_, new_n964_ );
nand g624 ( new_n967_, new_n966_, N219, new_n963_ );
not g625 ( new_n968_, N210 );
or g626 ( new_n969_, new_n535_, new_n968_ );
nand g627 ( new_n970_, new_n967_, new_n955_, new_n969_ );
nand g628 ( new_n971_, new_n967_, new_n969_ );
nand g629 ( new_n972_, new_n971_, keyIn_0_250 );
nand g630 ( new_n973_, new_n972_, new_n970_ );
nand g631 ( new_n974_, new_n957_, N228 );
or g632 ( new_n975_, new_n916_, new_n758_ );
nand g633 ( new_n976_, new_n974_, new_n975_ );
nor g634 ( new_n977_, new_n976_, keyIn_0_192 );
and g635 ( new_n978_, new_n976_, keyIn_0_192 );
nand g636 ( new_n979_, new_n908_, N246 );
xor g637 ( new_n980_, new_n979_, keyIn_0_120 );
nand g638 ( new_n981_, new_n585_, N159 );
nand g639 ( new_n982_, new_n980_, new_n981_ );
xnor g640 ( new_n983_, new_n982_, keyIn_0_143 );
nor g641 ( new_n984_, new_n978_, new_n977_, new_n983_ );
nand g642 ( new_n985_, new_n973_, new_n954_, new_n984_ );
nand g643 ( new_n986_, new_n973_, new_n984_ );
nand g644 ( new_n987_, new_n986_, keyIn_0_253 );
nand g645 ( N878, new_n987_, new_n985_ );
not g646 ( new_n989_, keyIn_0_245 );
not g647 ( new_n990_, keyIn_0_224 );
and g648 ( new_n991_, new_n853_, new_n870_ );
nand g649 ( new_n992_, new_n817_, new_n814_, new_n991_ );
nand g650 ( new_n993_, new_n992_, new_n990_ );
nand g651 ( new_n994_, new_n817_, keyIn_0_224, new_n814_, new_n991_ );
nand g652 ( new_n995_, new_n993_, new_n994_ );
and g653 ( new_n996_, new_n877_, new_n853_ );
and g654 ( new_n997_, new_n996_, keyIn_0_189 );
nor g655 ( new_n998_, new_n996_, keyIn_0_189 );
xor g656 ( new_n999_, new_n882_, keyIn_0_169 );
nor g657 ( new_n1000_, new_n999_, new_n997_, new_n998_ );
nand g658 ( new_n1001_, new_n995_, new_n1000_ );
nand g659 ( new_n1002_, new_n1001_, keyIn_0_227 );
not g660 ( new_n1003_, keyIn_0_227 );
nand g661 ( new_n1004_, new_n995_, new_n1003_, new_n1000_ );
nand g662 ( new_n1005_, new_n1002_, new_n1004_ );
nand g663 ( new_n1006_, new_n838_, new_n887_ );
xor g664 ( new_n1007_, new_n1006_, keyIn_0_145 );
nand g665 ( new_n1008_, new_n1005_, keyIn_0_236, new_n1007_ );
not g666 ( new_n1009_, keyIn_0_236 );
nand g667 ( new_n1010_, new_n1005_, new_n1007_ );
nand g668 ( new_n1011_, new_n1010_, new_n1009_ );
nand g669 ( new_n1012_, new_n1011_, new_n1008_ );
not g670 ( new_n1013_, new_n1007_ );
nand g671 ( new_n1014_, new_n1002_, new_n1004_, new_n1013_ );
xnor g672 ( new_n1015_, new_n1014_, keyIn_0_235 );
nand g673 ( new_n1016_, new_n1012_, new_n1015_, new_n989_ );
nand g674 ( new_n1017_, new_n1012_, new_n1015_ );
nand g675 ( new_n1018_, new_n1017_, keyIn_0_245 );
nand g676 ( new_n1019_, new_n1018_, N219, new_n1016_ );
nand g677 ( new_n1020_, N91, N210 );
nand g678 ( new_n1021_, new_n1019_, keyIn_0_251, new_n1020_ );
not g679 ( new_n1022_, keyIn_0_251 );
nand g680 ( new_n1023_, new_n1019_, new_n1020_ );
nand g681 ( new_n1024_, new_n1023_, new_n1022_ );
nand g682 ( new_n1025_, new_n1024_, new_n1021_ );
nand g683 ( new_n1026_, new_n1007_, N228 );
nand g684 ( new_n1027_, new_n888_, N237 );
nand g685 ( new_n1028_, new_n1026_, new_n1027_ );
nor g686 ( new_n1029_, new_n1028_, keyIn_0_193 );
and g687 ( new_n1030_, new_n1028_, keyIn_0_193 );
nand g688 ( new_n1031_, new_n836_, N246 );
xnor g689 ( new_n1032_, new_n1031_, keyIn_0_123 );
nand g690 ( new_n1033_, new_n585_, N165 );
nand g691 ( new_n1034_, new_n1032_, new_n1033_ );
xor g692 ( new_n1035_, new_n1034_, keyIn_0_146 );
nor g693 ( new_n1036_, new_n1030_, new_n1029_, new_n1035_ );
nand g694 ( new_n1037_, new_n1025_, keyIn_0_254, new_n1036_ );
not g695 ( new_n1038_, keyIn_0_254 );
nand g696 ( new_n1039_, new_n1025_, new_n1036_ );
nand g697 ( new_n1040_, new_n1039_, new_n1038_ );
nand g698 ( N879, new_n1040_, new_n1037_ );
not g699 ( new_n1042_, keyIn_0_252 );
not g700 ( new_n1043_, keyIn_0_246 );
not g701 ( new_n1044_, keyIn_0_228 );
nand g702 ( new_n1045_, new_n817_, new_n814_, new_n870_ );
or g703 ( new_n1046_, new_n1045_, keyIn_0_223 );
nand g704 ( new_n1047_, new_n1045_, keyIn_0_223 );
xor g705 ( new_n1048_, new_n877_, keyIn_0_171 );
nand g706 ( new_n1049_, new_n1046_, new_n1047_, new_n1048_ );
nand g707 ( new_n1050_, new_n1049_, new_n1044_ );
nand g708 ( new_n1051_, new_n1046_, keyIn_0_228, new_n1047_, new_n1048_ );
nand g709 ( new_n1052_, new_n1050_, new_n1051_ );
nand g710 ( new_n1053_, new_n853_, new_n881_ );
xnor g711 ( new_n1054_, new_n1053_, keyIn_0_148 );
not g712 ( new_n1055_, new_n1054_ );
nand g713 ( new_n1056_, new_n1052_, new_n1055_ );
xnor g714 ( new_n1057_, new_n1056_, keyIn_0_237 );
nand g715 ( new_n1058_, new_n1050_, new_n1051_, new_n1054_ );
xor g716 ( new_n1059_, new_n1058_, keyIn_0_238 );
nand g717 ( new_n1060_, new_n1057_, new_n1059_, new_n1043_ );
nand g718 ( new_n1061_, new_n1057_, new_n1059_ );
nand g719 ( new_n1062_, new_n1061_, keyIn_0_246 );
nand g720 ( new_n1063_, new_n1062_, N219, new_n1060_ );
nand g721 ( new_n1064_, N96, N210 );
nand g722 ( new_n1065_, new_n1063_, new_n1064_ );
nand g723 ( new_n1066_, new_n1065_, new_n1042_ );
nand g724 ( new_n1067_, new_n1063_, keyIn_0_252, new_n1064_ );
nand g725 ( new_n1068_, new_n882_, N237 );
xnor g726 ( new_n1069_, new_n1068_, keyIn_0_170 );
nand g727 ( new_n1070_, new_n1054_, N228 );
nand g728 ( new_n1071_, new_n1069_, new_n1070_ );
nor g729 ( new_n1072_, new_n1071_, keyIn_0_194 );
and g730 ( new_n1073_, new_n1071_, keyIn_0_194 );
not g731 ( new_n1074_, N246 );
nor g732 ( new_n1075_, new_n851_, new_n1074_ );
or g733 ( new_n1076_, new_n1075_, keyIn_0_126 );
nand g734 ( new_n1077_, new_n1075_, keyIn_0_126 );
nand g735 ( new_n1078_, new_n585_, N171 );
nand g736 ( new_n1079_, new_n1076_, new_n1077_, new_n1078_ );
xnor g737 ( new_n1080_, new_n1079_, keyIn_0_149 );
nor g738 ( new_n1081_, new_n1073_, new_n1072_, new_n1080_ );
nand g739 ( new_n1082_, new_n1066_, new_n1067_, new_n1081_ );
nand g740 ( new_n1083_, new_n1082_, keyIn_0_255 );
not g741 ( new_n1084_, keyIn_0_255 );
nand g742 ( new_n1085_, new_n1066_, new_n1084_, new_n1067_, new_n1081_ );
nand g743 ( N880, new_n1083_, new_n1085_ );
endmodule