module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n1105_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n1145_, new_n657_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1020_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n398_, new_n646_, new_n1132_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n1106_, new_n473_, new_n1147_, new_n790_, new_n1081_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n943_, new_n874_, new_n402_, new_n663_, new_n579_, new_n347_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n745_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1136_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n1056_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n905_, new_n539_, new_n803_, new_n727_, new_n375_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n780_, new_n984_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n877_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n866_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

nand g000 ( new_n343_, N29, N42, N75 );
not g001 ( N388, new_n343_ );
nand g002 ( new_n345_, N29, N36, N80 );
not g003 ( N389, new_n345_ );
nand g004 ( new_n347_, N29, N36, N42 );
not g005 ( N390, new_n347_ );
nand g006 ( new_n349_, N85, N86 );
not g007 ( N391, new_n349_ );
nand g008 ( new_n351_, N1, N8, N13, N17 );
not g009 ( N418, new_n351_ );
nand g010 ( new_n353_, N1, N13, N17, N26 );
nor g011 ( new_n354_, N390, new_n353_ );
xor g012 ( N419, new_n354_, keyIn_0_8 );
nand g013 ( N420, N59, N75, N80 );
nand g014 ( N421, N36, N59, N80 );
nand g015 ( N422, N36, N42, N59 );
not g016 ( new_n359_, N90 );
nor g017 ( new_n360_, N87, N88 );
nor g018 ( N423, new_n360_, new_n359_ );
nor g019 ( new_n362_, new_n353_, new_n347_ );
xor g020 ( N446, new_n362_, keyIn_0_25 );
not g021 ( new_n364_, keyIn_0_0 );
nand g022 ( new_n365_, new_n364_, N1, N26, N51 );
nand g023 ( new_n366_, N1, N26, N51 );
nand g024 ( new_n367_, new_n366_, keyIn_0_0 );
nand g025 ( new_n368_, new_n367_, new_n365_ );
not g026 ( N447, new_n368_ );
nand g027 ( new_n370_, N1, N8, N13, N55 );
not g028 ( new_n371_, new_n370_ );
nand g029 ( new_n372_, new_n371_, N29, N68 );
xnor g030 ( N448, new_n372_, keyIn_0_12 );
nand g031 ( new_n374_, N59, N68 );
not g032 ( new_n375_, new_n374_ );
nand g033 ( new_n376_, new_n371_, N74, new_n375_ );
xnor g034 ( N449, new_n376_, keyIn_0_13 );
not g035 ( new_n378_, N89 );
nor g036 ( N450, new_n360_, new_n378_ );
not g037 ( new_n380_, N135 );
xnor g038 ( new_n381_, N121, N126 );
xnor g039 ( new_n382_, new_n381_, keyIn_0_18 );
xor g040 ( new_n383_, new_n382_, keyIn_0_32 );
xor g041 ( new_n384_, N111, N116 );
xnor g042 ( new_n385_, new_n384_, keyIn_0_17 );
xor g043 ( new_n386_, new_n385_, keyIn_0_31 );
nand g044 ( new_n387_, new_n386_, new_n383_ );
xor g045 ( new_n388_, new_n387_, keyIn_0_43 );
nand g046 ( new_n389_, new_n385_, new_n382_ );
xor g047 ( new_n390_, new_n389_, keyIn_0_33 );
nand g048 ( new_n391_, new_n388_, new_n390_ );
xnor g049 ( new_n392_, new_n391_, keyIn_0_53 );
nand g050 ( new_n393_, new_n392_, new_n380_ );
xnor g051 ( new_n394_, new_n393_, keyIn_0_73 );
not g052 ( new_n395_, new_n392_ );
nand g053 ( new_n396_, new_n395_, N135 );
xnor g054 ( new_n397_, new_n396_, keyIn_0_72 );
nand g055 ( new_n398_, new_n397_, new_n394_ );
xnor g056 ( new_n399_, new_n398_, keyIn_0_95 );
not g057 ( new_n400_, new_n399_ );
not g058 ( new_n401_, N130 );
not g059 ( new_n402_, keyIn_0_42 );
xnor g060 ( new_n403_, N91, N96 );
xnor g061 ( new_n404_, new_n403_, keyIn_0_15 );
xor g062 ( new_n405_, new_n404_, keyIn_0_28 );
xor g063 ( new_n406_, N101, N106 );
xnor g064 ( new_n407_, new_n406_, keyIn_0_16 );
xor g065 ( new_n408_, new_n407_, keyIn_0_29 );
nand g066 ( new_n409_, new_n408_, new_n402_, new_n405_ );
nand g067 ( new_n410_, new_n408_, new_n405_ );
nand g068 ( new_n411_, new_n410_, keyIn_0_42 );
nand g069 ( new_n412_, new_n407_, new_n404_ );
xnor g070 ( new_n413_, new_n412_, keyIn_0_30 );
nand g071 ( new_n414_, new_n411_, new_n409_, new_n413_ );
xor g072 ( new_n415_, new_n414_, keyIn_0_52 );
nand g073 ( new_n416_, new_n415_, new_n401_ );
xnor g074 ( new_n417_, new_n416_, keyIn_0_71 );
not g075 ( new_n418_, new_n415_ );
nand g076 ( new_n419_, new_n418_, N130 );
xor g077 ( new_n420_, new_n419_, keyIn_0_70 );
nand g078 ( new_n421_, new_n420_, new_n417_ );
xnor g079 ( new_n422_, new_n421_, keyIn_0_94 );
nand g080 ( new_n423_, new_n400_, new_n422_ );
xor g081 ( new_n424_, new_n423_, keyIn_0_106 );
not g082 ( new_n425_, new_n422_ );
nand g083 ( new_n426_, new_n425_, new_n399_ );
xnor g084 ( new_n427_, new_n426_, keyIn_0_116 );
nand g085 ( new_n428_, new_n424_, new_n427_ );
xnor g086 ( N767, new_n428_, keyIn_0_139 );
xnor g087 ( new_n430_, N171, N177 );
xnor g088 ( new_n431_, new_n430_, keyIn_0_22 );
xor g089 ( new_n432_, new_n431_, keyIn_0_36 );
xor g090 ( new_n433_, N159, N165 );
xnor g091 ( new_n434_, new_n433_, keyIn_0_21 );
xor g092 ( new_n435_, new_n434_, keyIn_0_35 );
nand g093 ( new_n436_, new_n435_, new_n432_ );
xnor g094 ( new_n437_, new_n436_, keyIn_0_49 );
nand g095 ( new_n438_, new_n434_, new_n431_ );
xor g096 ( new_n439_, new_n438_, keyIn_0_37 );
nand g097 ( new_n440_, new_n437_, new_n439_ );
xor g098 ( new_n441_, new_n440_, keyIn_0_68 );
nand g099 ( new_n442_, new_n441_, new_n401_ );
xnor g100 ( new_n443_, new_n442_, keyIn_0_91 );
not g101 ( new_n444_, new_n441_ );
nand g102 ( new_n445_, new_n444_, N130 );
xnor g103 ( new_n446_, new_n445_, keyIn_0_90 );
nand g104 ( new_n447_, new_n446_, new_n443_ );
xor g105 ( new_n448_, new_n447_, keyIn_0_104 );
not g106 ( new_n449_, keyIn_0_50 );
xor g107 ( new_n450_, N195, N201 );
xnor g108 ( new_n451_, new_n450_, keyIn_0_24 );
xnor g109 ( new_n452_, new_n451_, keyIn_0_39 );
xor g110 ( new_n453_, N183, N189 );
xnor g111 ( new_n454_, new_n453_, keyIn_0_23 );
xnor g112 ( new_n455_, new_n454_, keyIn_0_38 );
nand g113 ( new_n456_, new_n452_, new_n455_, new_n449_ );
nand g114 ( new_n457_, new_n452_, new_n455_ );
nand g115 ( new_n458_, new_n457_, keyIn_0_50 );
nand g116 ( new_n459_, new_n451_, new_n454_ );
xnor g117 ( new_n460_, new_n459_, keyIn_0_40 );
nand g118 ( new_n461_, new_n458_, new_n456_, new_n460_ );
xnor g119 ( new_n462_, new_n461_, keyIn_0_69 );
nand g120 ( new_n463_, new_n462_, N207 );
xnor g121 ( new_n464_, new_n463_, keyIn_0_92 );
not g122 ( new_n465_, N207 );
not g123 ( new_n466_, new_n462_ );
nand g124 ( new_n467_, new_n466_, new_n465_ );
xor g125 ( new_n468_, new_n467_, keyIn_0_93 );
nand g126 ( new_n469_, new_n468_, new_n464_ );
xnor g127 ( new_n470_, new_n469_, keyIn_0_105 );
nor g128 ( new_n471_, new_n448_, new_n470_ );
xor g129 ( new_n472_, new_n471_, keyIn_0_115 );
nand g130 ( new_n473_, new_n448_, new_n470_ );
xnor g131 ( new_n474_, new_n473_, keyIn_0_117 );
nand g132 ( new_n475_, new_n472_, new_n474_ );
xnor g133 ( N768, new_n475_, keyIn_0_140 );
not g134 ( new_n477_, keyIn_0_216 );
not g135 ( new_n478_, keyIn_0_202 );
not g136 ( new_n479_, N261 );
not g137 ( new_n480_, keyIn_0_103 );
not g138 ( new_n481_, keyIn_0_48 );
nand g139 ( new_n482_, new_n368_, keyIn_0_9 );
not g140 ( new_n483_, keyIn_0_9 );
nand g141 ( new_n484_, new_n367_, new_n483_, new_n365_ );
nand g142 ( new_n485_, new_n482_, keyIn_0_26, new_n484_ );
not g143 ( new_n486_, keyIn_0_26 );
nand g144 ( new_n487_, new_n482_, new_n484_ );
nand g145 ( new_n488_, new_n487_, new_n486_ );
nand g146 ( new_n489_, new_n488_, new_n485_ );
nand g147 ( new_n490_, N59, N156 );
xnor g148 ( new_n491_, new_n490_, keyIn_0_5 );
nand g149 ( new_n492_, new_n489_, new_n481_, N17, new_n491_ );
nand g150 ( new_n493_, new_n489_, N17, new_n491_ );
nand g151 ( new_n494_, new_n493_, keyIn_0_48 );
nand g152 ( new_n495_, new_n494_, new_n492_ );
nand g153 ( new_n496_, new_n495_, keyIn_0_63, N1 );
not g154 ( new_n497_, keyIn_0_63 );
nand g155 ( new_n498_, new_n495_, N1 );
nand g156 ( new_n499_, new_n498_, new_n497_ );
nand g157 ( new_n500_, new_n499_, new_n496_ );
nand g158 ( new_n501_, new_n500_, N153 );
nand g159 ( new_n502_, new_n501_, keyIn_0_88 );
not g160 ( new_n503_, keyIn_0_88 );
nand g161 ( new_n504_, new_n500_, new_n503_, N153 );
nand g162 ( new_n505_, new_n502_, new_n504_ );
not g163 ( new_n506_, keyIn_0_89 );
not g164 ( new_n507_, keyIn_0_54 );
not g165 ( new_n508_, keyIn_0_47 );
nor g166 ( new_n509_, N17, N42 );
xnor g167 ( new_n510_, new_n509_, keyIn_0_6 );
nand g168 ( new_n511_, N17, N42 );
xnor g169 ( new_n512_, new_n511_, keyIn_0_7 );
nor g170 ( new_n513_, new_n510_, new_n512_ );
nand g171 ( new_n514_, new_n513_, keyIn_0_20 );
nor g172 ( new_n515_, new_n513_, keyIn_0_20 );
nor g173 ( new_n516_, new_n515_, new_n490_ );
nand g174 ( new_n517_, new_n516_, new_n489_, new_n508_, new_n514_ );
nand g175 ( new_n518_, new_n516_, new_n489_, new_n514_ );
nand g176 ( new_n519_, new_n518_, keyIn_0_47 );
not g177 ( new_n520_, keyIn_0_1 );
nand g178 ( new_n521_, N1, N8, N17, N51 );
xnor g179 ( new_n522_, new_n521_, new_n520_ );
xnor g180 ( new_n523_, new_n522_, keyIn_0_10 );
not g181 ( new_n524_, keyIn_0_3 );
nand g182 ( new_n525_, N42, N59, N75 );
xnor g183 ( new_n526_, new_n525_, new_n524_ );
xnor g184 ( new_n527_, new_n526_, keyIn_0_14 );
nand g185 ( new_n528_, new_n523_, new_n527_ );
xnor g186 ( new_n529_, new_n528_, keyIn_0_34 );
nand g187 ( new_n530_, new_n529_, new_n519_, new_n507_, new_n517_ );
nand g188 ( new_n531_, new_n529_, new_n519_, new_n517_ );
nand g189 ( new_n532_, new_n531_, keyIn_0_54 );
nand g190 ( new_n533_, new_n532_, N126, new_n530_ );
nand g191 ( new_n534_, new_n533_, new_n506_ );
nand g192 ( new_n535_, new_n532_, keyIn_0_89, N126, new_n530_ );
nand g193 ( new_n536_, new_n534_, new_n535_ );
nand g194 ( new_n537_, new_n505_, new_n536_ );
nand g195 ( new_n538_, new_n537_, new_n480_ );
nand g196 ( new_n539_, new_n505_, keyIn_0_103, new_n536_ );
not g197 ( new_n540_, keyIn_0_46 );
nand g198 ( new_n541_, N29, N75, N80 );
xor g199 ( new_n542_, new_n541_, keyIn_0_2 );
nand g200 ( new_n543_, new_n489_, new_n542_ );
not g201 ( new_n544_, new_n543_ );
nand g202 ( new_n545_, new_n544_, new_n540_, N55 );
nand g203 ( new_n546_, new_n544_, N55 );
nand g204 ( new_n547_, new_n546_, keyIn_0_46 );
xor g205 ( new_n548_, keyIn_0_4, N268 );
xor g206 ( new_n549_, new_n548_, keyIn_0_19 );
nand g207 ( new_n550_, new_n547_, new_n545_, new_n549_ );
xnor g208 ( new_n551_, new_n550_, keyIn_0_67 );
nand g209 ( new_n552_, new_n538_, new_n539_, new_n551_ );
nand g210 ( new_n553_, new_n552_, keyIn_0_114 );
not g211 ( new_n554_, keyIn_0_114 );
nand g212 ( new_n555_, new_n538_, new_n554_, new_n539_, new_n551_ );
nand g213 ( new_n556_, new_n553_, N201, new_n555_ );
nand g214 ( new_n557_, new_n556_, keyIn_0_137 );
not g215 ( new_n558_, keyIn_0_137 );
nand g216 ( new_n559_, new_n553_, new_n558_, N201, new_n555_ );
nand g217 ( new_n560_, new_n557_, new_n559_ );
not g218 ( new_n561_, keyIn_0_138 );
not g219 ( new_n562_, N201 );
nand g220 ( new_n563_, new_n553_, new_n555_ );
nand g221 ( new_n564_, new_n563_, new_n561_, new_n562_ );
nand g222 ( new_n565_, new_n563_, new_n562_ );
nand g223 ( new_n566_, new_n565_, keyIn_0_138 );
nand g224 ( new_n567_, new_n560_, new_n564_, new_n566_ );
xnor g225 ( new_n568_, new_n567_, keyIn_0_163 );
nand g226 ( new_n569_, new_n568_, new_n479_ );
xnor g227 ( new_n570_, new_n569_, keyIn_0_184 );
not g228 ( new_n571_, new_n568_ );
nand g229 ( new_n572_, new_n571_, N261 );
xor g230 ( new_n573_, new_n572_, keyIn_0_185 );
nand g231 ( new_n574_, new_n573_, new_n570_ );
nand g232 ( new_n575_, new_n574_, new_n478_ );
nand g233 ( new_n576_, new_n573_, keyIn_0_202, new_n570_ );
nand g234 ( new_n577_, new_n575_, N219, new_n576_ );
xnor g235 ( new_n578_, new_n577_, keyIn_0_210 );
nand g236 ( new_n579_, N121, N210 );
nand g237 ( new_n580_, new_n578_, new_n477_, new_n579_ );
nand g238 ( new_n581_, new_n578_, new_n579_ );
nand g239 ( new_n582_, new_n581_, keyIn_0_216 );
nand g240 ( new_n583_, new_n571_, N228 );
nand g241 ( new_n584_, new_n557_, keyIn_0_162, new_n559_ );
not g242 ( new_n585_, keyIn_0_162 );
nand g243 ( new_n586_, new_n560_, new_n585_ );
nand g244 ( new_n587_, new_n586_, new_n584_ );
nand g245 ( new_n588_, new_n587_, N237 );
nand g246 ( new_n589_, new_n583_, keyIn_0_203, new_n588_ );
not g247 ( new_n590_, keyIn_0_203 );
nand g248 ( new_n591_, new_n583_, new_n588_ );
nand g249 ( new_n592_, new_n591_, new_n590_ );
nand g250 ( new_n593_, new_n553_, N246, new_n555_ );
nand g251 ( new_n594_, N255, N267 );
nand g252 ( new_n595_, new_n593_, new_n594_ );
xnor g253 ( new_n596_, new_n595_, keyIn_0_164 );
nand g254 ( new_n597_, new_n371_, N42, N72, new_n375_ );
xor g255 ( new_n598_, new_n597_, keyIn_0_11 );
nand g256 ( new_n599_, new_n598_, N73 );
xnor g257 ( new_n600_, new_n599_, keyIn_0_27 );
xnor g258 ( new_n601_, new_n600_, keyIn_0_41 );
xnor g259 ( new_n602_, new_n601_, keyIn_0_51 );
nand g260 ( new_n603_, new_n602_, N201 );
nand g261 ( new_n604_, new_n592_, new_n589_, new_n596_, new_n603_ );
not g262 ( new_n605_, new_n604_ );
nand g263 ( new_n606_, new_n582_, new_n580_, new_n605_ );
xnor g264 ( N850, new_n606_, keyIn_0_222 );
not g265 ( new_n608_, keyIn_0_230 );
not g266 ( new_n609_, keyIn_0_196 );
not g267 ( new_n610_, N189 );
not g268 ( new_n611_, keyIn_0_112 );
not g269 ( new_n612_, keyIn_0_101 );
not g270 ( new_n613_, keyIn_0_84 );
nand g271 ( new_n614_, new_n500_, new_n613_, N146 );
nand g272 ( new_n615_, new_n500_, N146 );
nand g273 ( new_n616_, new_n615_, keyIn_0_84 );
nand g274 ( new_n617_, new_n616_, new_n614_ );
not g275 ( new_n618_, keyIn_0_85 );
nand g276 ( new_n619_, new_n532_, N116, new_n530_ );
xnor g277 ( new_n620_, new_n619_, new_n618_ );
nand g278 ( new_n621_, new_n617_, new_n620_, new_n612_ );
nand g279 ( new_n622_, new_n617_, new_n620_ );
nand g280 ( new_n623_, new_n622_, keyIn_0_101 );
xnor g281 ( new_n624_, new_n550_, keyIn_0_65 );
nand g282 ( new_n625_, new_n623_, new_n621_, new_n624_ );
nand g283 ( new_n626_, new_n625_, new_n611_ );
nand g284 ( new_n627_, new_n623_, keyIn_0_112, new_n621_, new_n624_ );
nand g285 ( new_n628_, new_n626_, new_n610_, new_n627_ );
xnor g286 ( new_n629_, new_n628_, keyIn_0_134 );
not g287 ( new_n630_, keyIn_0_113 );
not g288 ( new_n631_, keyIn_0_102 );
not g289 ( new_n632_, keyIn_0_86 );
nand g290 ( new_n633_, new_n500_, N149 );
nand g291 ( new_n634_, new_n633_, new_n632_ );
nand g292 ( new_n635_, new_n500_, keyIn_0_86, N149 );
nand g293 ( new_n636_, new_n634_, new_n635_ );
not g294 ( new_n637_, keyIn_0_87 );
nand g295 ( new_n638_, new_n532_, N121, new_n530_ );
xnor g296 ( new_n639_, new_n638_, new_n637_ );
nand g297 ( new_n640_, new_n636_, new_n639_ );
nand g298 ( new_n641_, new_n640_, new_n631_ );
nand g299 ( new_n642_, new_n636_, new_n639_, keyIn_0_102 );
xnor g300 ( new_n643_, new_n550_, keyIn_0_66 );
nand g301 ( new_n644_, new_n641_, new_n642_, new_n643_ );
nand g302 ( new_n645_, new_n644_, new_n630_ );
nand g303 ( new_n646_, new_n641_, keyIn_0_113, new_n642_, new_n643_ );
nand g304 ( new_n647_, new_n645_, new_n646_ );
nand g305 ( new_n648_, new_n647_, N195 );
nand g306 ( new_n649_, new_n648_, keyIn_0_135 );
not g307 ( new_n650_, keyIn_0_135 );
nand g308 ( new_n651_, new_n647_, new_n650_, N195 );
nand g309 ( new_n652_, new_n649_, keyIn_0_159, new_n651_ );
not g310 ( new_n653_, keyIn_0_159 );
nand g311 ( new_n654_, new_n649_, new_n651_ );
nand g312 ( new_n655_, new_n654_, new_n653_ );
nand g313 ( new_n656_, new_n655_, new_n652_ );
nand g314 ( new_n657_, new_n656_, keyIn_0_187, new_n629_ );
not g315 ( new_n658_, keyIn_0_187 );
nand g316 ( new_n659_, new_n656_, new_n629_ );
nand g317 ( new_n660_, new_n659_, new_n658_ );
nand g318 ( new_n661_, new_n660_, new_n657_ );
not g319 ( new_n662_, keyIn_0_167 );
not g320 ( new_n663_, keyIn_0_134 );
nand g321 ( new_n664_, new_n628_, new_n663_ );
nand g322 ( new_n665_, new_n626_, keyIn_0_134, new_n610_, new_n627_ );
not g323 ( new_n666_, keyIn_0_136 );
not g324 ( new_n667_, N195 );
nand g325 ( new_n668_, new_n645_, new_n667_, new_n646_ );
nand g326 ( new_n669_, new_n668_, new_n666_ );
nand g327 ( new_n670_, new_n645_, keyIn_0_136, new_n667_, new_n646_ );
nand g328 ( new_n671_, new_n664_, new_n669_, new_n665_, new_n670_ );
nand g329 ( new_n672_, new_n566_, N261, new_n564_ );
nor g330 ( new_n673_, new_n672_, new_n671_, new_n662_ );
nor g331 ( new_n674_, new_n672_, new_n671_ );
nor g332 ( new_n675_, new_n674_, keyIn_0_167 );
nor g333 ( new_n676_, new_n675_, new_n673_ );
not g334 ( new_n677_, new_n671_ );
nand g335 ( new_n678_, new_n587_, new_n677_ );
nand g336 ( new_n679_, new_n678_, keyIn_0_188 );
not g337 ( new_n680_, new_n679_ );
nor g338 ( new_n681_, new_n680_, new_n676_ );
not g339 ( new_n682_, keyIn_0_177 );
not g340 ( new_n683_, keyIn_0_156 );
not g341 ( new_n684_, keyIn_0_133 );
nand g342 ( new_n685_, new_n626_, new_n627_ );
nand g343 ( new_n686_, new_n685_, N189 );
nand g344 ( new_n687_, new_n686_, new_n684_ );
nand g345 ( new_n688_, new_n685_, keyIn_0_133, N189 );
nand g346 ( new_n689_, new_n687_, new_n688_ );
nand g347 ( new_n690_, new_n689_, new_n683_ );
nand g348 ( new_n691_, new_n687_, keyIn_0_156, new_n688_ );
nand g349 ( new_n692_, new_n690_, new_n682_, new_n691_ );
nand g350 ( new_n693_, new_n690_, new_n691_ );
nand g351 ( new_n694_, new_n693_, keyIn_0_177 );
nand g352 ( new_n695_, new_n694_, new_n692_ );
not g353 ( new_n696_, keyIn_0_188 );
nand g354 ( new_n697_, new_n587_, new_n696_, new_n677_ );
nand g355 ( new_n698_, new_n681_, new_n661_, new_n695_, new_n697_ );
nand g356 ( new_n699_, new_n698_, new_n609_ );
nand g357 ( new_n700_, new_n695_, new_n697_ );
not g358 ( new_n701_, new_n700_ );
nand g359 ( new_n702_, new_n701_, keyIn_0_196, new_n661_, new_n681_ );
nand g360 ( new_n703_, new_n699_, new_n702_ );
nand g361 ( new_n704_, new_n500_, N143 );
xor g362 ( new_n705_, new_n704_, keyIn_0_82 );
xnor g363 ( new_n706_, new_n531_, new_n507_ );
nand g364 ( new_n707_, new_n706_, N111 );
xor g365 ( new_n708_, new_n707_, keyIn_0_83 );
nand g366 ( new_n709_, new_n708_, new_n705_ );
xor g367 ( new_n710_, new_n709_, keyIn_0_100 );
xnor g368 ( new_n711_, new_n550_, keyIn_0_64 );
nand g369 ( new_n712_, new_n710_, new_n711_ );
xnor g370 ( new_n713_, new_n712_, keyIn_0_111 );
nand g371 ( new_n714_, new_n713_, N183 );
xnor g372 ( new_n715_, new_n714_, keyIn_0_130 );
not g373 ( new_n716_, N183 );
not g374 ( new_n717_, new_n713_ );
nand g375 ( new_n718_, new_n717_, new_n716_ );
xor g376 ( new_n719_, new_n718_, keyIn_0_131 );
nand g377 ( new_n720_, new_n719_, new_n715_ );
xnor g378 ( new_n721_, new_n720_, keyIn_0_154 );
nand g379 ( new_n722_, new_n721_, new_n703_ );
xnor g380 ( new_n723_, new_n722_, keyIn_0_204 );
not g381 ( new_n724_, new_n721_ );
nand g382 ( new_n725_, new_n724_, new_n699_, new_n702_ );
xor g383 ( new_n726_, new_n725_, keyIn_0_205 );
nand g384 ( new_n727_, new_n726_, new_n723_ );
xnor g385 ( new_n728_, new_n727_, keyIn_0_213 );
nand g386 ( new_n729_, new_n728_, N219 );
xnor g387 ( new_n730_, new_n729_, keyIn_0_219 );
nand g388 ( new_n731_, N106, N210 );
nand g389 ( new_n732_, new_n730_, new_n608_, new_n731_ );
nand g390 ( new_n733_, new_n730_, new_n731_ );
nand g391 ( new_n734_, new_n733_, keyIn_0_230 );
not g392 ( new_n735_, keyIn_0_197 );
nand g393 ( new_n736_, new_n724_, N228 );
xnor g394 ( new_n737_, new_n736_, keyIn_0_175 );
xor g395 ( new_n738_, new_n715_, keyIn_0_153 );
nand g396 ( new_n739_, new_n738_, N237 );
xnor g397 ( new_n740_, new_n739_, keyIn_0_176 );
nand g398 ( new_n741_, new_n737_, new_n740_ );
nand g399 ( new_n742_, new_n741_, new_n735_ );
nand g400 ( new_n743_, new_n737_, keyIn_0_197, new_n740_ );
not g401 ( new_n744_, keyIn_0_132 );
nand g402 ( new_n745_, new_n713_, N246 );
nand g403 ( new_n746_, new_n745_, new_n744_ );
nand g404 ( new_n747_, new_n713_, keyIn_0_132, N246 );
nand g405 ( new_n748_, new_n602_, N183 );
nand g406 ( new_n749_, new_n746_, new_n747_, new_n748_ );
xor g407 ( new_n750_, new_n749_, keyIn_0_155 );
nand g408 ( new_n751_, new_n743_, new_n750_ );
not g409 ( new_n752_, new_n751_ );
nand g410 ( new_n753_, new_n734_, new_n732_, new_n742_, new_n752_ );
xor g411 ( N863, new_n753_, keyIn_0_240 );
not g412 ( new_n755_, keyIn_0_231 );
xnor g413 ( new_n756_, new_n668_, keyIn_0_136 );
nand g414 ( new_n757_, new_n587_, new_n756_ );
xor g415 ( new_n758_, new_n757_, keyIn_0_186 );
xor g416 ( new_n759_, new_n656_, keyIn_0_180 );
nand g417 ( new_n760_, new_n756_, N261, new_n564_, new_n566_ );
xor g418 ( new_n761_, new_n760_, keyIn_0_166 );
nand g419 ( new_n762_, new_n758_, new_n759_, new_n761_ );
xnor g420 ( new_n763_, new_n762_, keyIn_0_198 );
nand g421 ( new_n764_, new_n689_, new_n629_ );
xor g422 ( new_n765_, new_n764_, keyIn_0_157 );
nand g423 ( new_n766_, new_n763_, new_n765_ );
xor g424 ( new_n767_, new_n766_, keyIn_0_206 );
not g425 ( new_n768_, new_n763_ );
not g426 ( new_n769_, new_n765_ );
nand g427 ( new_n770_, new_n768_, new_n769_ );
xnor g428 ( new_n771_, new_n770_, keyIn_0_207 );
nand g429 ( new_n772_, new_n771_, new_n767_ );
xor g430 ( new_n773_, new_n772_, keyIn_0_214 );
nand g431 ( new_n774_, new_n773_, N219 );
xnor g432 ( new_n775_, new_n774_, keyIn_0_220 );
nand g433 ( new_n776_, N111, N210 );
nand g434 ( new_n777_, new_n775_, new_n755_, new_n776_ );
nand g435 ( new_n778_, new_n775_, new_n776_ );
nand g436 ( new_n779_, new_n778_, keyIn_0_231 );
nand g437 ( new_n780_, new_n769_, N228 );
xor g438 ( new_n781_, new_n780_, keyIn_0_178 );
nand g439 ( new_n782_, new_n690_, N237, new_n691_ );
xor g440 ( new_n783_, new_n782_, keyIn_0_179 );
nand g441 ( new_n784_, new_n781_, new_n783_ );
xnor g442 ( new_n785_, new_n784_, keyIn_0_199 );
not g443 ( new_n786_, keyIn_0_158 );
nand g444 ( new_n787_, new_n685_, N246 );
nand g445 ( new_n788_, N255, N259 );
nand g446 ( new_n789_, new_n787_, new_n786_, new_n788_ );
nand g447 ( new_n790_, new_n787_, new_n788_ );
nand g448 ( new_n791_, new_n790_, keyIn_0_158 );
nand g449 ( new_n792_, new_n602_, N189 );
nand g450 ( new_n793_, new_n785_, new_n789_, new_n791_, new_n792_ );
not g451 ( new_n794_, new_n793_ );
nand g452 ( new_n795_, new_n779_, new_n777_, new_n794_ );
xor g453 ( N864, new_n795_, keyIn_0_241 );
not g454 ( new_n797_, keyIn_0_215 );
xnor g455 ( new_n798_, new_n587_, keyIn_0_183 );
xnor g456 ( new_n799_, new_n672_, keyIn_0_165 );
nand g457 ( new_n800_, new_n798_, new_n799_ );
xor g458 ( new_n801_, new_n800_, keyIn_0_200 );
not g459 ( new_n802_, new_n801_ );
nand g460 ( new_n803_, new_n654_, new_n756_ );
xor g461 ( new_n804_, new_n803_, keyIn_0_160 );
not g462 ( new_n805_, new_n804_ );
nand g463 ( new_n806_, new_n802_, new_n805_ );
xor g464 ( new_n807_, new_n806_, keyIn_0_208 );
nand g465 ( new_n808_, new_n801_, new_n804_ );
xor g466 ( new_n809_, new_n808_, keyIn_0_209 );
nand g467 ( new_n810_, new_n807_, new_n809_ );
nand g468 ( new_n811_, new_n810_, new_n797_ );
nand g469 ( new_n812_, new_n807_, keyIn_0_215, new_n809_ );
nand g470 ( new_n813_, new_n811_, N219, new_n812_ );
xor g471 ( new_n814_, new_n813_, keyIn_0_221 );
nand g472 ( new_n815_, N116, N210 );
nand g473 ( new_n816_, new_n814_, new_n815_ );
xnor g474 ( new_n817_, new_n816_, keyIn_0_232 );
nand g475 ( new_n818_, new_n804_, N228 );
xor g476 ( new_n819_, new_n818_, keyIn_0_181 );
nand g477 ( new_n820_, new_n656_, N237 );
xor g478 ( new_n821_, new_n820_, keyIn_0_182 );
nand g479 ( new_n822_, new_n819_, new_n821_ );
xnor g480 ( new_n823_, new_n822_, keyIn_0_201 );
not g481 ( new_n824_, keyIn_0_161 );
nand g482 ( new_n825_, new_n647_, N246 );
nand g483 ( new_n826_, N255, N260 );
nand g484 ( new_n827_, new_n825_, new_n824_, new_n826_ );
nand g485 ( new_n828_, new_n825_, new_n826_ );
nand g486 ( new_n829_, new_n828_, keyIn_0_161 );
nand g487 ( new_n830_, new_n602_, N195 );
nand g488 ( new_n831_, new_n829_, new_n827_, new_n830_ );
not g489 ( new_n832_, new_n831_ );
nand g490 ( new_n833_, new_n817_, new_n823_, new_n832_ );
xor g491 ( N865, new_n833_, keyIn_0_242 );
not g492 ( new_n835_, keyIn_0_243 );
not g493 ( new_n836_, keyIn_0_226 );
not g494 ( new_n837_, keyIn_0_225 );
not g495 ( new_n838_, keyIn_0_212 );
not g496 ( new_n839_, keyIn_0_211 );
nand g497 ( new_n840_, new_n699_, new_n839_, new_n702_, new_n719_ );
nand g498 ( new_n841_, new_n699_, new_n702_, new_n719_ );
nand g499 ( new_n842_, new_n841_, keyIn_0_211 );
nand g500 ( new_n843_, new_n842_, new_n840_ );
not g501 ( new_n844_, keyIn_0_174 );
xnor g502 ( new_n845_, new_n738_, new_n844_ );
nand g503 ( new_n846_, new_n843_, new_n845_ );
nand g504 ( new_n847_, new_n846_, new_n838_ );
nand g505 ( new_n848_, new_n843_, keyIn_0_212, new_n845_ );
not g506 ( new_n849_, N171 );
nand g507 ( new_n850_, new_n706_, N101 );
xor g508 ( new_n851_, new_n850_, keyIn_0_78 );
nand g509 ( new_n852_, N17, N138 );
nand g510 ( new_n853_, new_n851_, new_n852_ );
xnor g511 ( new_n854_, new_n853_, keyIn_0_98 );
nand g512 ( new_n855_, new_n489_, N55, new_n491_ );
xor g513 ( new_n856_, new_n855_, keyIn_0_44 );
nand g514 ( new_n857_, new_n856_, N149 );
xnor g515 ( new_n858_, new_n857_, keyIn_0_59 );
not g516 ( new_n859_, keyIn_0_45 );
nand g517 ( new_n860_, new_n544_, new_n859_, N17 );
nand g518 ( new_n861_, new_n544_, N17 );
nand g519 ( new_n862_, new_n861_, keyIn_0_45 );
nand g520 ( new_n863_, new_n862_, new_n548_, new_n860_ );
xor g521 ( new_n864_, new_n863_, keyIn_0_60 );
nand g522 ( new_n865_, new_n864_, new_n858_ );
xor g523 ( new_n866_, new_n865_, keyIn_0_79 );
nand g524 ( new_n867_, new_n854_, new_n866_ );
xnor g525 ( new_n868_, new_n867_, keyIn_0_109 );
nand g526 ( new_n869_, new_n868_, new_n849_ );
xor g527 ( new_n870_, new_n869_, keyIn_0_125 );
not g528 ( new_n871_, N165 );
nand g529 ( new_n872_, new_n706_, N96 );
xor g530 ( new_n873_, new_n872_, keyIn_0_76 );
nand g531 ( new_n874_, N51, N138 );
nand g532 ( new_n875_, new_n873_, new_n874_ );
xor g533 ( new_n876_, new_n875_, keyIn_0_97 );
xor g534 ( new_n877_, new_n863_, keyIn_0_58 );
nand g535 ( new_n878_, new_n856_, N146 );
xor g536 ( new_n879_, new_n878_, keyIn_0_57 );
nand g537 ( new_n880_, new_n879_, new_n877_ );
xor g538 ( new_n881_, new_n880_, keyIn_0_77 );
nand g539 ( new_n882_, new_n876_, new_n881_ );
xor g540 ( new_n883_, new_n882_, keyIn_0_108 );
nand g541 ( new_n884_, new_n883_, new_n871_ );
xnor g542 ( new_n885_, new_n884_, keyIn_0_122 );
nand g543 ( new_n886_, new_n885_, new_n870_ );
not g544 ( new_n887_, new_n886_ );
not g545 ( new_n888_, N177 );
not g546 ( new_n889_, keyIn_0_99 );
not g547 ( new_n890_, keyIn_0_80 );
nand g548 ( new_n891_, new_n706_, new_n890_, N106 );
nand g549 ( new_n892_, new_n706_, N106 );
nand g550 ( new_n893_, new_n892_, keyIn_0_80 );
nand g551 ( new_n894_, N138, N152 );
nand g552 ( new_n895_, new_n893_, new_n891_, new_n894_ );
nand g553 ( new_n896_, new_n895_, new_n889_ );
nand g554 ( new_n897_, new_n856_, N153 );
xnor g555 ( new_n898_, new_n897_, keyIn_0_61 );
xor g556 ( new_n899_, new_n863_, keyIn_0_62 );
nand g557 ( new_n900_, new_n899_, new_n898_ );
xnor g558 ( new_n901_, new_n900_, keyIn_0_81 );
nand g559 ( new_n902_, new_n893_, keyIn_0_99, new_n891_, new_n894_ );
nand g560 ( new_n903_, new_n901_, new_n896_, new_n902_ );
xor g561 ( new_n904_, new_n903_, keyIn_0_110 );
nand g562 ( new_n905_, new_n904_, new_n888_ );
xor g563 ( new_n906_, new_n905_, keyIn_0_128 );
nand g564 ( new_n907_, new_n887_, new_n906_ );
not g565 ( new_n908_, new_n907_ );
nand g566 ( new_n909_, new_n847_, new_n837_, new_n848_, new_n908_ );
nand g567 ( new_n910_, new_n847_, new_n848_, new_n908_ );
nand g568 ( new_n911_, new_n910_, keyIn_0_225 );
not g569 ( new_n912_, new_n904_ );
nand g570 ( new_n913_, new_n912_, N177 );
xor g571 ( new_n914_, new_n913_, keyIn_0_127 );
xor g572 ( new_n915_, new_n914_, keyIn_0_150 );
nand g573 ( new_n916_, new_n887_, new_n915_ );
xnor g574 ( new_n917_, new_n916_, keyIn_0_191 );
not g575 ( new_n918_, new_n868_ );
nand g576 ( new_n919_, new_n918_, N171 );
xor g577 ( new_n920_, new_n919_, keyIn_0_124 );
xnor g578 ( new_n921_, new_n920_, keyIn_0_147 );
nand g579 ( new_n922_, new_n921_, keyIn_0_190, new_n885_ );
not g580 ( new_n923_, new_n883_ );
nand g581 ( new_n924_, new_n923_, N165 );
xor g582 ( new_n925_, new_n924_, keyIn_0_121 );
xnor g583 ( new_n926_, new_n925_, keyIn_0_144 );
xor g584 ( new_n927_, new_n926_, keyIn_0_168 );
not g585 ( new_n928_, keyIn_0_190 );
nand g586 ( new_n929_, new_n921_, new_n885_ );
nand g587 ( new_n930_, new_n929_, new_n928_ );
nand g588 ( new_n931_, new_n927_, new_n917_, new_n922_, new_n930_ );
not g589 ( new_n932_, new_n931_ );
nand g590 ( new_n933_, new_n911_, new_n909_, new_n932_ );
xnor g591 ( new_n934_, new_n933_, new_n836_ );
not g592 ( new_n935_, N159 );
not g593 ( new_n936_, keyIn_0_96 );
nand g594 ( new_n937_, new_n706_, N91 );
xor g595 ( new_n938_, new_n937_, keyIn_0_74 );
nand g596 ( new_n939_, N8, N138 );
nand g597 ( new_n940_, new_n938_, new_n936_, new_n939_ );
nand g598 ( new_n941_, new_n938_, new_n939_ );
nand g599 ( new_n942_, new_n941_, keyIn_0_96 );
xor g600 ( new_n943_, new_n863_, keyIn_0_56 );
nand g601 ( new_n944_, new_n856_, N143 );
xor g602 ( new_n945_, new_n944_, keyIn_0_55 );
nand g603 ( new_n946_, new_n945_, new_n943_ );
xor g604 ( new_n947_, new_n946_, keyIn_0_75 );
nand g605 ( new_n948_, new_n942_, new_n940_, new_n947_ );
xor g606 ( new_n949_, new_n948_, keyIn_0_107 );
nand g607 ( new_n950_, new_n949_, new_n935_ );
xor g608 ( new_n951_, new_n950_, keyIn_0_119 );
nand g609 ( new_n952_, new_n934_, new_n835_, new_n951_ );
nand g610 ( new_n953_, new_n934_, new_n951_ );
nand g611 ( new_n954_, new_n953_, keyIn_0_243 );
not g612 ( new_n955_, new_n949_ );
nand g613 ( new_n956_, new_n955_, N159 );
xnor g614 ( new_n957_, new_n956_, keyIn_0_118 );
xor g615 ( new_n958_, new_n957_, keyIn_0_141 );
nand g616 ( new_n959_, new_n954_, new_n952_, new_n958_ );
xor g617 ( N866, new_n959_, keyIn_0_248 );
not g618 ( new_n961_, keyIn_0_247 );
not g619 ( new_n962_, keyIn_0_229 );
nand g620 ( new_n963_, new_n847_, new_n848_ );
nand g621 ( new_n964_, new_n914_, new_n906_ );
xnor g622 ( new_n965_, new_n964_, keyIn_0_151 );
not g623 ( new_n966_, new_n965_ );
nand g624 ( new_n967_, new_n963_, new_n966_ );
xnor g625 ( new_n968_, new_n967_, keyIn_0_217 );
not g626 ( new_n969_, new_n963_ );
nand g627 ( new_n970_, new_n969_, new_n965_ );
xnor g628 ( new_n971_, new_n970_, keyIn_0_218 );
nand g629 ( new_n972_, new_n971_, new_n962_, new_n968_ );
nand g630 ( new_n973_, new_n971_, new_n968_ );
nand g631 ( new_n974_, new_n973_, keyIn_0_229 );
nand g632 ( new_n975_, new_n974_, N219, new_n972_ );
xnor g633 ( new_n976_, new_n975_, keyIn_0_239 );
nand g634 ( new_n977_, N101, N210 );
nand g635 ( new_n978_, new_n976_, new_n977_ );
xnor g636 ( new_n979_, new_n978_, new_n961_ );
not g637 ( new_n980_, keyIn_0_195 );
nand g638 ( new_n981_, new_n965_, N228 );
xnor g639 ( new_n982_, new_n981_, keyIn_0_172 );
nand g640 ( new_n983_, new_n915_, N237 );
xor g641 ( new_n984_, new_n983_, keyIn_0_173 );
nand g642 ( new_n985_, new_n984_, new_n982_, new_n980_ );
nand g643 ( new_n986_, new_n984_, new_n982_ );
nand g644 ( new_n987_, new_n986_, keyIn_0_195 );
not g645 ( new_n988_, keyIn_0_129 );
nand g646 ( new_n989_, new_n912_, new_n988_, N246 );
nand g647 ( new_n990_, new_n912_, N246 );
nand g648 ( new_n991_, new_n990_, keyIn_0_129 );
nand g649 ( new_n992_, new_n602_, N177 );
nand g650 ( new_n993_, new_n991_, new_n989_, new_n992_ );
xnor g651 ( new_n994_, new_n993_, keyIn_0_152 );
nand g652 ( new_n995_, new_n987_, new_n985_, new_n994_ );
not g653 ( new_n996_, new_n995_ );
nand g654 ( new_n997_, new_n979_, new_n996_ );
xnor g655 ( N874, new_n997_, keyIn_0_249 );
not g656 ( new_n999_, keyIn_0_234 );
nand g657 ( new_n1000_, new_n957_, new_n951_ );
xor g658 ( new_n1001_, new_n1000_, keyIn_0_142 );
nand g659 ( new_n1002_, new_n934_, new_n999_, new_n1001_ );
nand g660 ( new_n1003_, new_n934_, new_n1001_ );
nand g661 ( new_n1004_, new_n1003_, keyIn_0_234 );
nand g662 ( new_n1005_, new_n1004_, new_n1002_ );
not g663 ( new_n1006_, keyIn_0_233 );
xnor g664 ( new_n1007_, new_n933_, keyIn_0_226 );
not g665 ( new_n1008_, new_n1001_ );
nand g666 ( new_n1009_, new_n1007_, new_n1006_, new_n1008_ );
nand g667 ( new_n1010_, new_n1007_, new_n1008_ );
nand g668 ( new_n1011_, new_n1010_, keyIn_0_233 );
nand g669 ( new_n1012_, new_n1011_, new_n1009_ );
nand g670 ( new_n1013_, new_n1005_, new_n1012_, keyIn_0_244 );
not g671 ( new_n1014_, keyIn_0_244 );
nand g672 ( new_n1015_, new_n1005_, new_n1012_ );
nand g673 ( new_n1016_, new_n1015_, new_n1014_ );
nand g674 ( new_n1017_, new_n1016_, N219, new_n1013_ );
not g675 ( new_n1018_, new_n549_ );
nand g676 ( new_n1019_, new_n1018_, N210 );
nand g677 ( new_n1020_, new_n1017_, new_n1019_ );
nand g678 ( new_n1021_, new_n1020_, keyIn_0_250 );
not g679 ( new_n1022_, keyIn_0_250 );
nand g680 ( new_n1023_, new_n1017_, new_n1022_, new_n1019_ );
nand g681 ( new_n1024_, new_n1021_, new_n1023_ );
not g682 ( new_n1025_, keyIn_0_192 );
nand g683 ( new_n1026_, new_n1001_, N228 );
not g684 ( new_n1027_, new_n958_ );
nand g685 ( new_n1028_, new_n1027_, N237 );
nand g686 ( new_n1029_, new_n1026_, new_n1025_, new_n1028_ );
nand g687 ( new_n1030_, new_n1026_, new_n1028_ );
nand g688 ( new_n1031_, new_n1030_, keyIn_0_192 );
nand g689 ( new_n1032_, new_n955_, N246 );
xor g690 ( new_n1033_, new_n1032_, keyIn_0_120 );
nand g691 ( new_n1034_, new_n602_, N159 );
nand g692 ( new_n1035_, new_n1033_, new_n1034_ );
xor g693 ( new_n1036_, new_n1035_, keyIn_0_143 );
nand g694 ( new_n1037_, new_n1031_, new_n1029_, new_n1036_ );
not g695 ( new_n1038_, new_n1037_ );
nand g696 ( new_n1039_, new_n1024_, new_n1038_ );
nand g697 ( new_n1040_, new_n1039_, keyIn_0_253 );
not g698 ( new_n1041_, keyIn_0_253 );
nand g699 ( new_n1042_, new_n1024_, new_n1041_, new_n1038_ );
nand g700 ( N878, new_n1040_, new_n1042_ );
not g701 ( new_n1044_, keyIn_0_254 );
not g702 ( new_n1045_, keyIn_0_251 );
not g703 ( new_n1046_, keyIn_0_245 );
nand g704 ( new_n1047_, new_n870_, new_n906_ );
not g705 ( new_n1048_, new_n1047_ );
nand g706 ( new_n1049_, new_n847_, keyIn_0_224, new_n848_, new_n1048_ );
not g707 ( new_n1050_, keyIn_0_224 );
nand g708 ( new_n1051_, new_n847_, new_n848_, new_n1048_ );
nand g709 ( new_n1052_, new_n1051_, new_n1050_ );
nand g710 ( new_n1053_, new_n1052_, new_n1049_ );
nand g711 ( new_n1054_, new_n915_, keyIn_0_189, new_n870_ );
not g712 ( new_n1055_, keyIn_0_189 );
nand g713 ( new_n1056_, new_n915_, new_n870_ );
nand g714 ( new_n1057_, new_n1056_, new_n1055_ );
xnor g715 ( new_n1058_, new_n921_, keyIn_0_169 );
nand g716 ( new_n1059_, new_n1058_, new_n1054_, new_n1057_ );
not g717 ( new_n1060_, new_n1059_ );
nand g718 ( new_n1061_, new_n1053_, new_n1060_ );
nand g719 ( new_n1062_, new_n1061_, keyIn_0_227 );
not g720 ( new_n1063_, keyIn_0_227 );
nand g721 ( new_n1064_, new_n1053_, new_n1063_, new_n1060_ );
not g722 ( new_n1065_, new_n925_ );
nand g723 ( new_n1066_, new_n1065_, new_n885_ );
xor g724 ( new_n1067_, new_n1066_, keyIn_0_145 );
not g725 ( new_n1068_, new_n1067_ );
nand g726 ( new_n1069_, new_n1062_, new_n1064_, new_n1068_ );
xnor g727 ( new_n1070_, new_n1069_, keyIn_0_235 );
nand g728 ( new_n1071_, new_n1062_, new_n1064_ );
nand g729 ( new_n1072_, new_n1071_, keyIn_0_236, new_n1067_ );
not g730 ( new_n1073_, keyIn_0_236 );
nand g731 ( new_n1074_, new_n1071_, new_n1067_ );
nand g732 ( new_n1075_, new_n1074_, new_n1073_ );
nand g733 ( new_n1076_, new_n1075_, new_n1072_ );
nand g734 ( new_n1077_, new_n1076_, new_n1070_, new_n1046_ );
nand g735 ( new_n1078_, new_n1076_, new_n1070_ );
nand g736 ( new_n1079_, new_n1078_, keyIn_0_245 );
nand g737 ( new_n1080_, new_n1079_, N219, new_n1077_ );
nand g738 ( new_n1081_, N91, N210 );
nand g739 ( new_n1082_, new_n1080_, new_n1081_ );
nand g740 ( new_n1083_, new_n1082_, new_n1045_ );
nand g741 ( new_n1084_, new_n1080_, keyIn_0_251, new_n1081_ );
nand g742 ( new_n1085_, new_n1083_, new_n1084_ );
not g743 ( new_n1086_, keyIn_0_193 );
nand g744 ( new_n1087_, new_n1067_, N228 );
nand g745 ( new_n1088_, new_n926_, N237 );
nand g746 ( new_n1089_, new_n1087_, new_n1086_, new_n1088_ );
nand g747 ( new_n1090_, new_n1087_, new_n1088_ );
nand g748 ( new_n1091_, new_n1090_, keyIn_0_193 );
nand g749 ( new_n1092_, new_n923_, N246 );
xnor g750 ( new_n1093_, new_n1092_, keyIn_0_123 );
nand g751 ( new_n1094_, new_n602_, N165 );
nand g752 ( new_n1095_, new_n1093_, new_n1094_ );
xnor g753 ( new_n1096_, new_n1095_, keyIn_0_146 );
nand g754 ( new_n1097_, new_n1091_, new_n1089_, new_n1096_ );
not g755 ( new_n1098_, new_n1097_ );
nand g756 ( new_n1099_, new_n1085_, new_n1098_ );
nand g757 ( new_n1100_, new_n1099_, new_n1044_ );
nand g758 ( new_n1101_, new_n1085_, keyIn_0_254, new_n1098_ );
nand g759 ( N879, new_n1100_, new_n1101_ );
not g760 ( new_n1103_, keyIn_0_252 );
not g761 ( new_n1104_, keyIn_0_246 );
not g762 ( new_n1105_, keyIn_0_223 );
nand g763 ( new_n1106_, new_n969_, new_n1105_, new_n906_ );
nand g764 ( new_n1107_, new_n847_, new_n848_, new_n906_ );
nand g765 ( new_n1108_, new_n1107_, keyIn_0_223 );
xor g766 ( new_n1109_, new_n915_, keyIn_0_171 );
nand g767 ( new_n1110_, new_n1106_, keyIn_0_228, new_n1108_, new_n1109_ );
not g768 ( new_n1111_, keyIn_0_228 );
nand g769 ( new_n1112_, new_n1106_, new_n1108_, new_n1109_ );
nand g770 ( new_n1113_, new_n1112_, new_n1111_ );
nand g771 ( new_n1114_, new_n1113_, new_n1110_ );
nand g772 ( new_n1115_, new_n920_, new_n870_ );
xnor g773 ( new_n1116_, new_n1115_, keyIn_0_148 );
not g774 ( new_n1117_, new_n1116_ );
nand g775 ( new_n1118_, new_n1114_, new_n1117_ );
xnor g776 ( new_n1119_, new_n1118_, keyIn_0_237 );
nand g777 ( new_n1120_, new_n1113_, new_n1110_, new_n1116_ );
xor g778 ( new_n1121_, new_n1120_, keyIn_0_238 );
nand g779 ( new_n1122_, new_n1119_, new_n1121_, new_n1104_ );
nand g780 ( new_n1123_, new_n1119_, new_n1121_ );
nand g781 ( new_n1124_, new_n1123_, keyIn_0_246 );
nand g782 ( new_n1125_, new_n1124_, N219, new_n1122_ );
nand g783 ( new_n1126_, N96, N210 );
nand g784 ( new_n1127_, new_n1125_, new_n1126_ );
nand g785 ( new_n1128_, new_n1127_, new_n1103_ );
nand g786 ( new_n1129_, new_n1125_, keyIn_0_252, new_n1126_ );
not g787 ( new_n1130_, keyIn_0_194 );
nand g788 ( new_n1131_, new_n921_, N237 );
xnor g789 ( new_n1132_, new_n1131_, keyIn_0_170 );
nand g790 ( new_n1133_, new_n1116_, N228 );
nand g791 ( new_n1134_, new_n1132_, new_n1130_, new_n1133_ );
nand g792 ( new_n1135_, new_n1132_, new_n1133_ );
nand g793 ( new_n1136_, new_n1135_, keyIn_0_194 );
not g794 ( new_n1137_, keyIn_0_126 );
nand g795 ( new_n1138_, new_n918_, N246 );
nand g796 ( new_n1139_, new_n1138_, new_n1137_ );
nand g797 ( new_n1140_, new_n918_, keyIn_0_126, N246 );
nand g798 ( new_n1141_, new_n602_, N171 );
nand g799 ( new_n1142_, new_n1139_, new_n1140_, new_n1141_ );
xor g800 ( new_n1143_, new_n1142_, keyIn_0_149 );
nand g801 ( new_n1144_, new_n1136_, new_n1134_, new_n1143_ );
not g802 ( new_n1145_, new_n1144_ );
nand g803 ( new_n1146_, new_n1128_, new_n1129_, new_n1145_ );
nand g804 ( new_n1147_, new_n1146_, keyIn_0_255 );
not g805 ( new_n1148_, keyIn_0_255 );
nand g806 ( new_n1149_, new_n1128_, new_n1148_, new_n1129_, new_n1145_ );
nand g807 ( N880, new_n1147_, new_n1149_ );
endmodule