module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999;

  AND2_X1 U2020 ( .A1(n1988), .A2(n1989), .ZN(Result_9_) );
  XOR2_X1 U2021 ( .A(n1990), .B(n1991), .Z(n1988) );
  AND2_X1 U2022 ( .A1(n1992), .A2(n1993), .ZN(n1991) );
  OR2_X1 U2023 ( .A1(n1994), .A2(n1995), .ZN(n1993) );
  INV_X1 U2024 ( .A(n1996), .ZN(n1992) );
  AND2_X1 U2025 ( .A1(n1997), .A2(n1989), .ZN(Result_8_) );
  XOR2_X1 U2026 ( .A(n1998), .B(n1999), .Z(n1997) );
  AND2_X1 U2027 ( .A1(n1989), .A2(n2000), .ZN(Result_7_) );
  XOR2_X1 U2028 ( .A(n2001), .B(n2002), .Z(n2000) );
  AND2_X1 U2029 ( .A1(n2003), .A2(n2004), .ZN(n2002) );
  OR2_X1 U2030 ( .A1(n2005), .A2(n2006), .ZN(n2004) );
  INV_X1 U2031 ( .A(n2007), .ZN(n2003) );
  AND2_X1 U2032 ( .A1(n2008), .A2(n1989), .ZN(Result_6_) );
  XOR2_X1 U2033 ( .A(n2009), .B(n2010), .Z(n2008) );
  AND2_X1 U2034 ( .A1(n1989), .A2(n2011), .ZN(Result_5_) );
  XOR2_X1 U2035 ( .A(n2012), .B(n2013), .Z(n2011) );
  AND2_X1 U2036 ( .A1(n2014), .A2(n2015), .ZN(n2013) );
  OR2_X1 U2037 ( .A1(n2016), .A2(n2017), .ZN(n2015) );
  INV_X1 U2038 ( .A(n2018), .ZN(n2014) );
  AND2_X1 U2039 ( .A1(n2019), .A2(n1989), .ZN(Result_4_) );
  XOR2_X1 U2040 ( .A(n2020), .B(n2021), .Z(n2019) );
  AND2_X1 U2041 ( .A1(n1989), .A2(n2022), .ZN(Result_3_) );
  XOR2_X1 U2042 ( .A(n2023), .B(n2024), .Z(n2022) );
  AND2_X1 U2043 ( .A1(n2025), .A2(n2026), .ZN(n2024) );
  OR2_X1 U2044 ( .A1(n2027), .A2(n2028), .ZN(n2026) );
  INV_X1 U2045 ( .A(n2029), .ZN(n2025) );
  OR2_X1 U2046 ( .A1(n2030), .A2(n2031), .ZN(Result_31_) );
  AND2_X1 U2047 ( .A1(n2032), .A2(n1989), .ZN(n2031) );
  AND2_X1 U2048 ( .A1(n2033), .A2(n2034), .ZN(n2030) );
  XNOR2_X1 U2049 ( .A(n2035), .B(a_15_), .ZN(n2033) );
  OR2_X1 U2050 ( .A1(n2036), .A2(n2037), .ZN(Result_30_) );
  OR2_X1 U2051 ( .A1(n2038), .A2(n2039), .ZN(n2037) );
  AND2_X1 U2052 ( .A1(n2040), .A2(n1989), .ZN(n2039) );
  AND2_X1 U2053 ( .A1(b_15_), .A2(n2041), .ZN(n2040) );
  OR2_X1 U2054 ( .A1(n2042), .A2(n2043), .ZN(n2041) );
  AND2_X1 U2055 ( .A1(n2044), .A2(n2034), .ZN(n2038) );
  OR2_X1 U2056 ( .A1(n2045), .A2(n2046), .ZN(n2044) );
  AND2_X1 U2057 ( .A1(n2047), .A2(n2032), .ZN(n2046) );
  AND2_X1 U2058 ( .A1(n2048), .A2(n2049), .ZN(n2047) );
  AND2_X1 U2059 ( .A1(n2042), .A2(n2050), .ZN(n2045) );
  AND2_X1 U2060 ( .A1(n2051), .A2(b_14_), .ZN(n2036) );
  AND2_X1 U2061 ( .A1(n2052), .A2(n2053), .ZN(n2051) );
  OR2_X1 U2062 ( .A1(n1989), .A2(n2054), .ZN(n2053) );
  XNOR2_X1 U2063 ( .A(a_14_), .B(n2032), .ZN(n2054) );
  INV_X1 U2064 ( .A(n2050), .ZN(n2032) );
  OR2_X1 U2065 ( .A1(n2034), .A2(n2055), .ZN(n2052) );
  OR2_X1 U2066 ( .A1(n2056), .A2(n2057), .ZN(n2055) );
  AND2_X1 U2067 ( .A1(a_15_), .A2(n2035), .ZN(n2057) );
  AND2_X1 U2068 ( .A1(n2058), .A2(n1989), .ZN(Result_2_) );
  XOR2_X1 U2069 ( .A(n2059), .B(n2060), .Z(n2058) );
  OR2_X1 U2070 ( .A1(n2061), .A2(n2062), .ZN(Result_29_) );
  AND2_X1 U2071 ( .A1(n2063), .A2(n1989), .ZN(n2062) );
  XOR2_X1 U2072 ( .A(n2064), .B(n2065), .Z(n2063) );
  XNOR2_X1 U2073 ( .A(n2066), .B(n2067), .ZN(n2065) );
  AND2_X1 U2074 ( .A1(n2068), .A2(n2034), .ZN(n2061) );
  OR2_X1 U2075 ( .A1(n2069), .A2(n2070), .ZN(n2068) );
  OR2_X1 U2076 ( .A1(n2071), .A2(n2072), .ZN(n2070) );
  AND2_X1 U2077 ( .A1(n2073), .A2(n2074), .ZN(n2072) );
  INV_X1 U2078 ( .A(n2075), .ZN(n2071) );
  OR2_X1 U2079 ( .A1(n2076), .A2(n2074), .ZN(n2075) );
  AND2_X1 U2080 ( .A1(n2077), .A2(n2078), .ZN(n2069) );
  XNOR2_X1 U2081 ( .A(n2074), .B(a_13_), .ZN(n2077) );
  OR2_X1 U2082 ( .A1(n2079), .A2(n2080), .ZN(Result_28_) );
  AND2_X1 U2083 ( .A1(n2081), .A2(n1989), .ZN(n2080) );
  XNOR2_X1 U2084 ( .A(n2082), .B(n2083), .ZN(n2081) );
  XOR2_X1 U2085 ( .A(n2084), .B(n2085), .Z(n2083) );
  AND2_X1 U2086 ( .A1(n2086), .A2(n2034), .ZN(n2079) );
  XOR2_X1 U2087 ( .A(n2087), .B(n2088), .Z(n2086) );
  OR2_X1 U2088 ( .A1(n2089), .A2(n2090), .ZN(n2088) );
  OR2_X1 U2089 ( .A1(n2091), .A2(n2092), .ZN(Result_27_) );
  AND2_X1 U2090 ( .A1(n2093), .A2(n1989), .ZN(n2092) );
  XNOR2_X1 U2091 ( .A(n2094), .B(n2095), .ZN(n2093) );
  XOR2_X1 U2092 ( .A(n2096), .B(n2097), .Z(n2095) );
  AND2_X1 U2093 ( .A1(n2098), .A2(n2034), .ZN(n2091) );
  OR2_X1 U2094 ( .A1(n2099), .A2(n2100), .ZN(n2098) );
  OR2_X1 U2095 ( .A1(n2101), .A2(n2102), .ZN(n2100) );
  INV_X1 U2096 ( .A(n2103), .ZN(n2102) );
  OR2_X1 U2097 ( .A1(n2104), .A2(n2105), .ZN(n2103) );
  AND2_X1 U2098 ( .A1(n2106), .A2(n2104), .ZN(n2101) );
  AND2_X1 U2099 ( .A1(n2107), .A2(n2108), .ZN(n2099) );
  XNOR2_X1 U2100 ( .A(a_11_), .B(n2104), .ZN(n2107) );
  OR2_X1 U2101 ( .A1(n2109), .A2(n2110), .ZN(Result_26_) );
  AND2_X1 U2102 ( .A1(n2111), .A2(n1989), .ZN(n2110) );
  XNOR2_X1 U2103 ( .A(n2112), .B(n2113), .ZN(n2111) );
  XOR2_X1 U2104 ( .A(n2114), .B(n2115), .Z(n2113) );
  AND2_X1 U2105 ( .A1(n2116), .A2(n2034), .ZN(n2109) );
  XOR2_X1 U2106 ( .A(n2117), .B(n2118), .Z(n2116) );
  OR2_X1 U2107 ( .A1(n2119), .A2(n2120), .ZN(n2118) );
  OR2_X1 U2108 ( .A1(n2121), .A2(n2122), .ZN(Result_25_) );
  AND2_X1 U2109 ( .A1(n2123), .A2(n1989), .ZN(n2122) );
  XNOR2_X1 U2110 ( .A(n2124), .B(n2125), .ZN(n2123) );
  XOR2_X1 U2111 ( .A(n2126), .B(n2127), .Z(n2125) );
  AND2_X1 U2112 ( .A1(n2128), .A2(n2034), .ZN(n2121) );
  OR2_X1 U2113 ( .A1(n2129), .A2(n2130), .ZN(n2128) );
  OR2_X1 U2114 ( .A1(n2131), .A2(n2132), .ZN(n2130) );
  INV_X1 U2115 ( .A(n2133), .ZN(n2132) );
  OR2_X1 U2116 ( .A1(n2134), .A2(n2135), .ZN(n2133) );
  AND2_X1 U2117 ( .A1(n2136), .A2(n2134), .ZN(n2131) );
  AND2_X1 U2118 ( .A1(n2137), .A2(n2138), .ZN(n2129) );
  XNOR2_X1 U2119 ( .A(a_9_), .B(n2134), .ZN(n2137) );
  OR2_X1 U2120 ( .A1(n2139), .A2(n2140), .ZN(Result_24_) );
  AND2_X1 U2121 ( .A1(n2141), .A2(n1989), .ZN(n2140) );
  XNOR2_X1 U2122 ( .A(n2142), .B(n2143), .ZN(n2141) );
  XOR2_X1 U2123 ( .A(n2144), .B(n2145), .Z(n2143) );
  AND2_X1 U2124 ( .A1(n2146), .A2(n2034), .ZN(n2139) );
  XOR2_X1 U2125 ( .A(n2147), .B(n2148), .Z(n2146) );
  OR2_X1 U2126 ( .A1(n2149), .A2(n2150), .ZN(n2148) );
  OR2_X1 U2127 ( .A1(n2151), .A2(n2152), .ZN(Result_23_) );
  AND2_X1 U2128 ( .A1(n2153), .A2(n1989), .ZN(n2152) );
  XNOR2_X1 U2129 ( .A(n2154), .B(n2155), .ZN(n2153) );
  XOR2_X1 U2130 ( .A(n2156), .B(n2157), .Z(n2155) );
  AND2_X1 U2131 ( .A1(n2158), .A2(n2034), .ZN(n2151) );
  OR2_X1 U2132 ( .A1(n2159), .A2(n2160), .ZN(n2158) );
  OR2_X1 U2133 ( .A1(n2161), .A2(n2162), .ZN(n2160) );
  INV_X1 U2134 ( .A(n2163), .ZN(n2162) );
  OR2_X1 U2135 ( .A1(n2164), .A2(n2165), .ZN(n2163) );
  AND2_X1 U2136 ( .A1(n2166), .A2(n2164), .ZN(n2161) );
  AND2_X1 U2137 ( .A1(n2167), .A2(n2168), .ZN(n2159) );
  XNOR2_X1 U2138 ( .A(a_7_), .B(n2164), .ZN(n2167) );
  OR2_X1 U2139 ( .A1(n2169), .A2(n2170), .ZN(Result_22_) );
  AND2_X1 U2140 ( .A1(n2171), .A2(n1989), .ZN(n2170) );
  XNOR2_X1 U2141 ( .A(n2172), .B(n2173), .ZN(n2171) );
  XOR2_X1 U2142 ( .A(n2174), .B(n2175), .Z(n2173) );
  AND2_X1 U2143 ( .A1(n2176), .A2(n2034), .ZN(n2169) );
  XOR2_X1 U2144 ( .A(n2177), .B(n2178), .Z(n2176) );
  OR2_X1 U2145 ( .A1(n2179), .A2(n2180), .ZN(n2178) );
  OR2_X1 U2146 ( .A1(n2181), .A2(n2182), .ZN(Result_21_) );
  AND2_X1 U2147 ( .A1(n2183), .A2(n1989), .ZN(n2182) );
  XNOR2_X1 U2148 ( .A(n2184), .B(n2185), .ZN(n2183) );
  XOR2_X1 U2149 ( .A(n2186), .B(n2187), .Z(n2185) );
  AND2_X1 U2150 ( .A1(n2188), .A2(n2034), .ZN(n2181) );
  OR2_X1 U2151 ( .A1(n2189), .A2(n2190), .ZN(n2188) );
  OR2_X1 U2152 ( .A1(n2191), .A2(n2192), .ZN(n2190) );
  INV_X1 U2153 ( .A(n2193), .ZN(n2192) );
  OR2_X1 U2154 ( .A1(n2194), .A2(n2195), .ZN(n2193) );
  AND2_X1 U2155 ( .A1(n2196), .A2(n2194), .ZN(n2191) );
  AND2_X1 U2156 ( .A1(n2197), .A2(n2198), .ZN(n2189) );
  XNOR2_X1 U2157 ( .A(a_5_), .B(n2194), .ZN(n2197) );
  OR2_X1 U2158 ( .A1(n2199), .A2(n2200), .ZN(Result_20_) );
  AND2_X1 U2159 ( .A1(n2201), .A2(n1989), .ZN(n2200) );
  XNOR2_X1 U2160 ( .A(n2202), .B(n2203), .ZN(n2201) );
  XOR2_X1 U2161 ( .A(n2204), .B(n2205), .Z(n2203) );
  AND2_X1 U2162 ( .A1(n2206), .A2(n2034), .ZN(n2199) );
  XOR2_X1 U2163 ( .A(n2207), .B(n2208), .Z(n2206) );
  OR2_X1 U2164 ( .A1(n2209), .A2(n2210), .ZN(n2208) );
  AND2_X1 U2165 ( .A1(n1989), .A2(n2211), .ZN(Result_1_) );
  XNOR2_X1 U2166 ( .A(n2212), .B(n2213), .ZN(n2211) );
  OR2_X1 U2167 ( .A1(n2214), .A2(n2215), .ZN(n2213) );
  AND2_X1 U2168 ( .A1(n2216), .A2(n2217), .ZN(n2215) );
  OR2_X1 U2169 ( .A1(n2218), .A2(n2219), .ZN(Result_19_) );
  AND2_X1 U2170 ( .A1(n2220), .A2(n1989), .ZN(n2219) );
  XNOR2_X1 U2171 ( .A(n2221), .B(n2222), .ZN(n2220) );
  XOR2_X1 U2172 ( .A(n2223), .B(n2224), .Z(n2222) );
  AND2_X1 U2173 ( .A1(n2225), .A2(n2034), .ZN(n2218) );
  OR2_X1 U2174 ( .A1(n2226), .A2(n2227), .ZN(n2225) );
  OR2_X1 U2175 ( .A1(n2228), .A2(n2229), .ZN(n2227) );
  INV_X1 U2176 ( .A(n2230), .ZN(n2229) );
  OR2_X1 U2177 ( .A1(n2231), .A2(n2232), .ZN(n2230) );
  AND2_X1 U2178 ( .A1(n2233), .A2(n2231), .ZN(n2228) );
  AND2_X1 U2179 ( .A1(n2234), .A2(n2235), .ZN(n2226) );
  XNOR2_X1 U2180 ( .A(a_3_), .B(n2231), .ZN(n2234) );
  OR2_X1 U2181 ( .A1(n2236), .A2(n2237), .ZN(Result_18_) );
  AND2_X1 U2182 ( .A1(n2238), .A2(n1989), .ZN(n2237) );
  XNOR2_X1 U2183 ( .A(n2239), .B(n2240), .ZN(n2238) );
  XOR2_X1 U2184 ( .A(n2241), .B(n2242), .Z(n2240) );
  AND2_X1 U2185 ( .A1(n2243), .A2(n2034), .ZN(n2236) );
  XOR2_X1 U2186 ( .A(n2244), .B(n2245), .Z(n2243) );
  OR2_X1 U2187 ( .A1(n2246), .A2(n2247), .ZN(n2245) );
  OR2_X1 U2188 ( .A1(n2248), .A2(n2249), .ZN(Result_17_) );
  AND2_X1 U2189 ( .A1(n2250), .A2(n1989), .ZN(n2249) );
  XNOR2_X1 U2190 ( .A(n2251), .B(n2252), .ZN(n2250) );
  XOR2_X1 U2191 ( .A(n2253), .B(n2254), .Z(n2252) );
  AND2_X1 U2192 ( .A1(n2255), .A2(n2034), .ZN(n2248) );
  XOR2_X1 U2193 ( .A(n2256), .B(n2257), .Z(n2255) );
  AND2_X1 U2194 ( .A1(n2258), .A2(n2259), .ZN(n2257) );
  INV_X1 U2195 ( .A(n2260), .ZN(n2258) );
  OR2_X1 U2196 ( .A1(n2261), .A2(n2262), .ZN(Result_16_) );
  AND2_X1 U2197 ( .A1(n2263), .A2(n1989), .ZN(n2262) );
  XNOR2_X1 U2198 ( .A(n2264), .B(n2265), .ZN(n2263) );
  XOR2_X1 U2199 ( .A(n2266), .B(n2267), .Z(n2265) );
  AND2_X1 U2200 ( .A1(n2268), .A2(n2034), .ZN(n2261) );
  XOR2_X1 U2201 ( .A(n2269), .B(n2270), .Z(n2268) );
  OR2_X1 U2202 ( .A1(a_0_), .A2(n2271), .ZN(n2270) );
  OR2_X1 U2203 ( .A1(n2272), .A2(n2273), .ZN(n2269) );
  AND2_X1 U2204 ( .A1(n2274), .A2(n2275), .ZN(n2273) );
  AND2_X1 U2205 ( .A1(n2256), .A2(n2276), .ZN(n2272) );
  OR2_X1 U2206 ( .A1(n2277), .A2(n2246), .ZN(n2256) );
  AND2_X1 U2207 ( .A1(n2278), .A2(n2279), .ZN(n2246) );
  AND2_X1 U2208 ( .A1(n2244), .A2(n2280), .ZN(n2277) );
  OR2_X1 U2209 ( .A1(n2281), .A2(n2282), .ZN(n2244) );
  AND2_X1 U2210 ( .A1(n2283), .A2(n2235), .ZN(n2282) );
  AND2_X1 U2211 ( .A1(n2231), .A2(n2232), .ZN(n2281) );
  OR2_X1 U2212 ( .A1(n2284), .A2(n2209), .ZN(n2231) );
  AND2_X1 U2213 ( .A1(n2285), .A2(n2286), .ZN(n2209) );
  AND2_X1 U2214 ( .A1(n2207), .A2(n2287), .ZN(n2284) );
  OR2_X1 U2215 ( .A1(n2288), .A2(n2289), .ZN(n2207) );
  AND2_X1 U2216 ( .A1(n2290), .A2(n2198), .ZN(n2289) );
  AND2_X1 U2217 ( .A1(n2194), .A2(n2195), .ZN(n2288) );
  OR2_X1 U2218 ( .A1(n2291), .A2(n2179), .ZN(n2194) );
  AND2_X1 U2219 ( .A1(n2292), .A2(n2293), .ZN(n2179) );
  AND2_X1 U2220 ( .A1(n2177), .A2(n2294), .ZN(n2291) );
  OR2_X1 U2221 ( .A1(n2295), .A2(n2296), .ZN(n2177) );
  AND2_X1 U2222 ( .A1(n2297), .A2(n2168), .ZN(n2296) );
  AND2_X1 U2223 ( .A1(n2164), .A2(n2165), .ZN(n2295) );
  OR2_X1 U2224 ( .A1(n2298), .A2(n2149), .ZN(n2164) );
  AND2_X1 U2225 ( .A1(n2299), .A2(n2300), .ZN(n2149) );
  AND2_X1 U2226 ( .A1(n2147), .A2(n2301), .ZN(n2298) );
  OR2_X1 U2227 ( .A1(n2302), .A2(n2303), .ZN(n2147) );
  AND2_X1 U2228 ( .A1(n2304), .A2(n2138), .ZN(n2303) );
  AND2_X1 U2229 ( .A1(n2134), .A2(n2135), .ZN(n2302) );
  OR2_X1 U2230 ( .A1(n2305), .A2(n2120), .ZN(n2134) );
  AND2_X1 U2231 ( .A1(n2306), .A2(n2307), .ZN(n2120) );
  AND2_X1 U2232 ( .A1(n2117), .A2(n2308), .ZN(n2305) );
  OR2_X1 U2233 ( .A1(n2309), .A2(n2310), .ZN(n2117) );
  AND2_X1 U2234 ( .A1(n2311), .A2(n2108), .ZN(n2310) );
  AND2_X1 U2235 ( .A1(n2104), .A2(n2105), .ZN(n2309) );
  OR2_X1 U2236 ( .A1(n2312), .A2(n2090), .ZN(n2104) );
  AND2_X1 U2237 ( .A1(n2313), .A2(n2314), .ZN(n2090) );
  AND2_X1 U2238 ( .A1(n2087), .A2(n2315), .ZN(n2312) );
  OR2_X1 U2239 ( .A1(n2316), .A2(n2317), .ZN(n2087) );
  AND2_X1 U2240 ( .A1(n2318), .A2(n2078), .ZN(n2317) );
  AND2_X1 U2241 ( .A1(n2074), .A2(n2076), .ZN(n2316) );
  AND2_X1 U2242 ( .A1(n2319), .A2(n2320), .ZN(n2074) );
  OR2_X1 U2243 ( .A1(n2049), .A2(n2321), .ZN(n2320) );
  AND2_X1 U2244 ( .A1(n2048), .A2(n2050), .ZN(n2321) );
  OR2_X1 U2245 ( .A1(n2322), .A2(n2035), .ZN(n2050) );
  AND2_X1 U2246 ( .A1(n1989), .A2(n2323), .ZN(Result_15_) );
  XNOR2_X1 U2247 ( .A(n2324), .B(n2325), .ZN(n2323) );
  AND2_X1 U2248 ( .A1(n2326), .A2(n1989), .ZN(Result_14_) );
  AND2_X1 U2249 ( .A1(n2327), .A2(n2328), .ZN(n2326) );
  OR2_X1 U2250 ( .A1(n2329), .A2(n2330), .ZN(n2327) );
  AND2_X1 U2251 ( .A1(n2331), .A2(n2325), .ZN(n2329) );
  AND2_X1 U2252 ( .A1(n1989), .A2(n2332), .ZN(Result_13_) );
  XOR2_X1 U2253 ( .A(n2328), .B(n2333), .Z(n2332) );
  OR2_X1 U2254 ( .A1(n2334), .A2(n2335), .ZN(n2333) );
  AND2_X1 U2255 ( .A1(n2336), .A2(n2337), .ZN(n2335) );
  INV_X1 U2256 ( .A(n2338), .ZN(n2328) );
  AND2_X1 U2257 ( .A1(n2339), .A2(n1989), .ZN(Result_12_) );
  XOR2_X1 U2258 ( .A(n2340), .B(n2341), .Z(n2339) );
  AND2_X1 U2259 ( .A1(n2342), .A2(n2343), .ZN(n2341) );
  OR2_X1 U2260 ( .A1(n2344), .A2(n2345), .ZN(n2343) );
  INV_X1 U2261 ( .A(n2346), .ZN(n2342) );
  AND2_X1 U2262 ( .A1(n2347), .A2(n1989), .ZN(Result_11_) );
  XOR2_X1 U2263 ( .A(n2348), .B(n2349), .Z(n2347) );
  AND2_X1 U2264 ( .A1(n2350), .A2(n2351), .ZN(n2349) );
  OR2_X1 U2265 ( .A1(n2352), .A2(n2353), .ZN(n2351) );
  AND2_X1 U2266 ( .A1(n2354), .A2(n2355), .ZN(n2352) );
  INV_X1 U2267 ( .A(n2356), .ZN(n2350) );
  AND2_X1 U2268 ( .A1(n2357), .A2(n1989), .ZN(Result_10_) );
  XOR2_X1 U2269 ( .A(n2358), .B(n2359), .Z(n2357) );
  AND2_X1 U2270 ( .A1(n2360), .A2(n2361), .ZN(n2359) );
  OR2_X1 U2271 ( .A1(n2362), .A2(n2363), .ZN(n2361) );
  AND2_X1 U2272 ( .A1(n2364), .A2(n2365), .ZN(n2362) );
  INV_X1 U2273 ( .A(n2366), .ZN(n2360) );
  AND2_X1 U2274 ( .A1(n1989), .A2(n2367), .ZN(Result_0_) );
  OR2_X1 U2275 ( .A1(n2368), .A2(n2369), .ZN(n2367) );
  OR2_X1 U2276 ( .A1(n2214), .A2(n2370), .ZN(n2369) );
  AND2_X1 U2277 ( .A1(n2371), .A2(b_0_), .ZN(n2370) );
  INV_X1 U2278 ( .A(n2372), .ZN(n2214) );
  OR2_X1 U2279 ( .A1(n2216), .A2(n2217), .ZN(n2372) );
  OR2_X1 U2280 ( .A1(n2373), .A2(n2374), .ZN(n2217) );
  AND2_X1 U2281 ( .A1(n2212), .A2(n2375), .ZN(n2368) );
  INV_X1 U2282 ( .A(n2216), .ZN(n2375) );
  OR2_X1 U2283 ( .A1(n2371), .A2(n2271), .ZN(n2216) );
  AND2_X1 U2284 ( .A1(n2059), .A2(n2060), .ZN(n2212) );
  XOR2_X1 U2285 ( .A(n2374), .B(n2373), .Z(n2060) );
  AND2_X1 U2286 ( .A1(n2376), .A2(n2377), .ZN(n2373) );
  AND2_X1 U2287 ( .A1(n2378), .A2(n2379), .ZN(n2377) );
  XNOR2_X1 U2288 ( .A(n2371), .B(n2380), .ZN(n2376) );
  AND2_X1 U2289 ( .A1(b_0_), .A2(a_1_), .ZN(n2380) );
  AND2_X1 U2290 ( .A1(b_1_), .A2(a_0_), .ZN(n2371) );
  AND2_X1 U2291 ( .A1(n2381), .A2(n2382), .ZN(n2374) );
  INV_X1 U2292 ( .A(n2383), .ZN(n2382) );
  AND2_X1 U2293 ( .A1(n2384), .A2(n2385), .ZN(n2383) );
  OR2_X1 U2294 ( .A1(n2386), .A2(n2387), .ZN(n2059) );
  OR2_X1 U2295 ( .A1(n2388), .A2(n2029), .ZN(n2386) );
  AND2_X1 U2296 ( .A1(n2027), .A2(n2028), .ZN(n2029) );
  AND2_X1 U2297 ( .A1(n2389), .A2(n2390), .ZN(n2028) );
  INV_X1 U2298 ( .A(n2391), .ZN(n2389) );
  AND2_X1 U2299 ( .A1(n2023), .A2(n2027), .ZN(n2388) );
  INV_X1 U2300 ( .A(n2392), .ZN(n2027) );
  OR2_X1 U2301 ( .A1(n2393), .A2(n2387), .ZN(n2392) );
  INV_X1 U2302 ( .A(n2394), .ZN(n2387) );
  OR2_X1 U2303 ( .A1(n2395), .A2(n2396), .ZN(n2394) );
  AND2_X1 U2304 ( .A1(n2395), .A2(n2396), .ZN(n2393) );
  OR2_X1 U2305 ( .A1(n2397), .A2(n2398), .ZN(n2396) );
  AND2_X1 U2306 ( .A1(n2399), .A2(n2400), .ZN(n2398) );
  AND2_X1 U2307 ( .A1(n2401), .A2(n2402), .ZN(n2397) );
  OR2_X1 U2308 ( .A1(n2400), .A2(n2399), .ZN(n2402) );
  XNOR2_X1 U2309 ( .A(n2385), .B(n2403), .ZN(n2395) );
  XNOR2_X1 U2310 ( .A(n2381), .B(n2384), .ZN(n2403) );
  AND2_X1 U2311 ( .A1(b_2_), .A2(a_0_), .ZN(n2384) );
  OR2_X1 U2312 ( .A1(n2404), .A2(n2405), .ZN(n2381) );
  AND2_X1 U2313 ( .A1(n2406), .A2(n2407), .ZN(n2405) );
  AND2_X1 U2314 ( .A1(n2408), .A2(n2409), .ZN(n2404) );
  OR2_X1 U2315 ( .A1(n2407), .A2(n2406), .ZN(n2409) );
  XOR2_X1 U2316 ( .A(n2410), .B(n2379), .Z(n2385) );
  OR2_X1 U2317 ( .A1(n2411), .A2(n2412), .ZN(n2379) );
  AND2_X1 U2318 ( .A1(n2413), .A2(n2414), .ZN(n2412) );
  AND2_X1 U2319 ( .A1(n2415), .A2(n2416), .ZN(n2411) );
  OR2_X1 U2320 ( .A1(n2414), .A2(n2413), .ZN(n2415) );
  OR2_X1 U2321 ( .A1(n2417), .A2(n2418), .ZN(n2410) );
  INV_X1 U2322 ( .A(n2378), .ZN(n2418) );
  OR2_X1 U2323 ( .A1(n2276), .A2(n2419), .ZN(n2378) );
  AND2_X1 U2324 ( .A1(n2419), .A2(n2276), .ZN(n2417) );
  OR2_X1 U2325 ( .A1(n2275), .A2(n2274), .ZN(n2276) );
  OR2_X1 U2326 ( .A1(n2278), .A2(n2271), .ZN(n2419) );
  AND2_X1 U2327 ( .A1(n2020), .A2(n2021), .ZN(n2023) );
  XNOR2_X1 U2328 ( .A(n2390), .B(n2391), .ZN(n2021) );
  OR2_X1 U2329 ( .A1(n2420), .A2(n2421), .ZN(n2391) );
  AND2_X1 U2330 ( .A1(n2422), .A2(n2423), .ZN(n2421) );
  AND2_X1 U2331 ( .A1(n2424), .A2(n2425), .ZN(n2420) );
  OR2_X1 U2332 ( .A1(n2423), .A2(n2422), .ZN(n2425) );
  XNOR2_X1 U2333 ( .A(n2401), .B(n2426), .ZN(n2390) );
  XOR2_X1 U2334 ( .A(n2400), .B(n2399), .Z(n2426) );
  OR2_X1 U2335 ( .A1(n2235), .A2(n2427), .ZN(n2399) );
  OR2_X1 U2336 ( .A1(n2428), .A2(n2429), .ZN(n2400) );
  AND2_X1 U2337 ( .A1(n2430), .A2(n2431), .ZN(n2429) );
  AND2_X1 U2338 ( .A1(n2432), .A2(n2433), .ZN(n2428) );
  OR2_X1 U2339 ( .A1(n2431), .A2(n2430), .ZN(n2433) );
  XOR2_X1 U2340 ( .A(n2408), .B(n2434), .Z(n2401) );
  XOR2_X1 U2341 ( .A(n2407), .B(n2406), .Z(n2434) );
  OR2_X1 U2342 ( .A1(n2279), .A2(n2274), .ZN(n2406) );
  OR2_X1 U2343 ( .A1(n2435), .A2(n2436), .ZN(n2407) );
  AND2_X1 U2344 ( .A1(n2437), .A2(n2280), .ZN(n2436) );
  AND2_X1 U2345 ( .A1(n2438), .A2(n2439), .ZN(n2435) );
  OR2_X1 U2346 ( .A1(n2280), .A2(n2437), .ZN(n2439) );
  XOR2_X1 U2347 ( .A(n2413), .B(n2440), .Z(n2408) );
  XOR2_X1 U2348 ( .A(n2414), .B(n2416), .Z(n2440) );
  OR2_X1 U2349 ( .A1(n2283), .A2(n2271), .ZN(n2416) );
  OR2_X1 U2350 ( .A1(n2441), .A2(n2442), .ZN(n2414) );
  AND2_X1 U2351 ( .A1(n2443), .A2(n2444), .ZN(n2442) );
  AND2_X1 U2352 ( .A1(n2445), .A2(n2446), .ZN(n2441) );
  OR2_X1 U2353 ( .A1(n2444), .A2(n2443), .ZN(n2445) );
  OR2_X1 U2354 ( .A1(n2275), .A2(n2278), .ZN(n2413) );
  OR2_X1 U2355 ( .A1(n2447), .A2(n2448), .ZN(n2020) );
  OR2_X1 U2356 ( .A1(n2449), .A2(n2018), .ZN(n2447) );
  AND2_X1 U2357 ( .A1(n2016), .A2(n2017), .ZN(n2018) );
  AND2_X1 U2358 ( .A1(n2450), .A2(n2451), .ZN(n2017) );
  INV_X1 U2359 ( .A(n2452), .ZN(n2450) );
  AND2_X1 U2360 ( .A1(n2012), .A2(n2016), .ZN(n2449) );
  INV_X1 U2361 ( .A(n2453), .ZN(n2016) );
  OR2_X1 U2362 ( .A1(n2454), .A2(n2448), .ZN(n2453) );
  INV_X1 U2363 ( .A(n2455), .ZN(n2448) );
  OR2_X1 U2364 ( .A1(n2456), .A2(n2457), .ZN(n2455) );
  AND2_X1 U2365 ( .A1(n2456), .A2(n2457), .ZN(n2454) );
  OR2_X1 U2366 ( .A1(n2458), .A2(n2459), .ZN(n2457) );
  AND2_X1 U2367 ( .A1(n2460), .A2(n2461), .ZN(n2459) );
  AND2_X1 U2368 ( .A1(n2462), .A2(n2463), .ZN(n2458) );
  OR2_X1 U2369 ( .A1(n2461), .A2(n2460), .ZN(n2463) );
  XOR2_X1 U2370 ( .A(n2424), .B(n2464), .Z(n2456) );
  XOR2_X1 U2371 ( .A(n2423), .B(n2422), .Z(n2464) );
  OR2_X1 U2372 ( .A1(n2286), .A2(n2427), .ZN(n2422) );
  OR2_X1 U2373 ( .A1(n2465), .A2(n2466), .ZN(n2423) );
  AND2_X1 U2374 ( .A1(n2467), .A2(n2468), .ZN(n2466) );
  AND2_X1 U2375 ( .A1(n2469), .A2(n2470), .ZN(n2465) );
  OR2_X1 U2376 ( .A1(n2468), .A2(n2467), .ZN(n2470) );
  XOR2_X1 U2377 ( .A(n2432), .B(n2471), .Z(n2424) );
  XOR2_X1 U2378 ( .A(n2431), .B(n2430), .Z(n2471) );
  OR2_X1 U2379 ( .A1(n2235), .A2(n2274), .ZN(n2430) );
  OR2_X1 U2380 ( .A1(n2472), .A2(n2473), .ZN(n2431) );
  AND2_X1 U2381 ( .A1(n2474), .A2(n2475), .ZN(n2473) );
  AND2_X1 U2382 ( .A1(n2476), .A2(n2477), .ZN(n2472) );
  OR2_X1 U2383 ( .A1(n2475), .A2(n2474), .ZN(n2477) );
  XNOR2_X1 U2384 ( .A(n2478), .B(n2438), .ZN(n2432) );
  XOR2_X1 U2385 ( .A(n2443), .B(n2479), .Z(n2438) );
  XOR2_X1 U2386 ( .A(n2444), .B(n2446), .Z(n2479) );
  OR2_X1 U2387 ( .A1(n2285), .A2(n2271), .ZN(n2446) );
  OR2_X1 U2388 ( .A1(n2480), .A2(n2481), .ZN(n2444) );
  AND2_X1 U2389 ( .A1(n2482), .A2(n2483), .ZN(n2481) );
  AND2_X1 U2390 ( .A1(n2484), .A2(n2485), .ZN(n2480) );
  OR2_X1 U2391 ( .A1(n2483), .A2(n2482), .ZN(n2484) );
  OR2_X1 U2392 ( .A1(n2275), .A2(n2283), .ZN(n2443) );
  XNOR2_X1 U2393 ( .A(n2280), .B(n2437), .ZN(n2478) );
  OR2_X1 U2394 ( .A1(n2486), .A2(n2487), .ZN(n2437) );
  AND2_X1 U2395 ( .A1(n2488), .A2(n2489), .ZN(n2487) );
  AND2_X1 U2396 ( .A1(n2490), .A2(n2491), .ZN(n2486) );
  OR2_X1 U2397 ( .A1(n2489), .A2(n2488), .ZN(n2491) );
  INV_X1 U2398 ( .A(n2247), .ZN(n2280) );
  AND2_X1 U2399 ( .A1(b_2_), .A2(a_2_), .ZN(n2247) );
  AND2_X1 U2400 ( .A1(n2009), .A2(n2010), .ZN(n2012) );
  XNOR2_X1 U2401 ( .A(n2451), .B(n2452), .ZN(n2010) );
  OR2_X1 U2402 ( .A1(n2492), .A2(n2493), .ZN(n2452) );
  AND2_X1 U2403 ( .A1(n2494), .A2(n2495), .ZN(n2493) );
  AND2_X1 U2404 ( .A1(n2496), .A2(n2497), .ZN(n2492) );
  OR2_X1 U2405 ( .A1(n2495), .A2(n2494), .ZN(n2497) );
  XNOR2_X1 U2406 ( .A(n2462), .B(n2498), .ZN(n2451) );
  XOR2_X1 U2407 ( .A(n2461), .B(n2460), .Z(n2498) );
  OR2_X1 U2408 ( .A1(n2198), .A2(n2427), .ZN(n2460) );
  OR2_X1 U2409 ( .A1(n2499), .A2(n2500), .ZN(n2461) );
  AND2_X1 U2410 ( .A1(n2501), .A2(n2502), .ZN(n2500) );
  AND2_X1 U2411 ( .A1(n2503), .A2(n2504), .ZN(n2499) );
  OR2_X1 U2412 ( .A1(n2502), .A2(n2501), .ZN(n2504) );
  XOR2_X1 U2413 ( .A(n2469), .B(n2505), .Z(n2462) );
  XOR2_X1 U2414 ( .A(n2468), .B(n2467), .Z(n2505) );
  OR2_X1 U2415 ( .A1(n2286), .A2(n2274), .ZN(n2467) );
  OR2_X1 U2416 ( .A1(n2506), .A2(n2507), .ZN(n2468) );
  AND2_X1 U2417 ( .A1(n2508), .A2(n2509), .ZN(n2507) );
  AND2_X1 U2418 ( .A1(n2510), .A2(n2511), .ZN(n2506) );
  OR2_X1 U2419 ( .A1(n2509), .A2(n2508), .ZN(n2511) );
  XOR2_X1 U2420 ( .A(n2476), .B(n2512), .Z(n2469) );
  XOR2_X1 U2421 ( .A(n2475), .B(n2474), .Z(n2512) );
  OR2_X1 U2422 ( .A1(n2235), .A2(n2278), .ZN(n2474) );
  OR2_X1 U2423 ( .A1(n2513), .A2(n2514), .ZN(n2475) );
  AND2_X1 U2424 ( .A1(n2232), .A2(n2515), .ZN(n2514) );
  AND2_X1 U2425 ( .A1(n2516), .A2(n2517), .ZN(n2513) );
  OR2_X1 U2426 ( .A1(n2515), .A2(n2232), .ZN(n2517) );
  XOR2_X1 U2427 ( .A(n2490), .B(n2518), .Z(n2476) );
  XOR2_X1 U2428 ( .A(n2489), .B(n2488), .Z(n2518) );
  OR2_X1 U2429 ( .A1(n2279), .A2(n2283), .ZN(n2488) );
  OR2_X1 U2430 ( .A1(n2519), .A2(n2520), .ZN(n2489) );
  AND2_X1 U2431 ( .A1(n2521), .A2(n2522), .ZN(n2520) );
  AND2_X1 U2432 ( .A1(n2523), .A2(n2524), .ZN(n2519) );
  OR2_X1 U2433 ( .A1(n2522), .A2(n2521), .ZN(n2524) );
  XOR2_X1 U2434 ( .A(n2482), .B(n2525), .Z(n2490) );
  XOR2_X1 U2435 ( .A(n2483), .B(n2485), .Z(n2525) );
  OR2_X1 U2436 ( .A1(n2290), .A2(n2271), .ZN(n2485) );
  OR2_X1 U2437 ( .A1(n2526), .A2(n2527), .ZN(n2483) );
  AND2_X1 U2438 ( .A1(n2528), .A2(n2529), .ZN(n2527) );
  AND2_X1 U2439 ( .A1(n2530), .A2(n2531), .ZN(n2526) );
  OR2_X1 U2440 ( .A1(n2529), .A2(n2528), .ZN(n2530) );
  OR2_X1 U2441 ( .A1(n2275), .A2(n2285), .ZN(n2482) );
  OR2_X1 U2442 ( .A1(n2532), .A2(n2533), .ZN(n2009) );
  OR2_X1 U2443 ( .A1(n2534), .A2(n2007), .ZN(n2532) );
  AND2_X1 U2444 ( .A1(n2005), .A2(n2006), .ZN(n2007) );
  AND2_X1 U2445 ( .A1(n2535), .A2(n2536), .ZN(n2006) );
  INV_X1 U2446 ( .A(n2537), .ZN(n2535) );
  AND2_X1 U2447 ( .A1(n2001), .A2(n2005), .ZN(n2534) );
  INV_X1 U2448 ( .A(n2538), .ZN(n2005) );
  OR2_X1 U2449 ( .A1(n2539), .A2(n2533), .ZN(n2538) );
  INV_X1 U2450 ( .A(n2540), .ZN(n2533) );
  OR2_X1 U2451 ( .A1(n2541), .A2(n2542), .ZN(n2540) );
  AND2_X1 U2452 ( .A1(n2541), .A2(n2542), .ZN(n2539) );
  OR2_X1 U2453 ( .A1(n2543), .A2(n2544), .ZN(n2542) );
  AND2_X1 U2454 ( .A1(n2545), .A2(n2546), .ZN(n2544) );
  AND2_X1 U2455 ( .A1(n2547), .A2(n2548), .ZN(n2543) );
  OR2_X1 U2456 ( .A1(n2546), .A2(n2545), .ZN(n2548) );
  XOR2_X1 U2457 ( .A(n2496), .B(n2549), .Z(n2541) );
  XOR2_X1 U2458 ( .A(n2495), .B(n2494), .Z(n2549) );
  OR2_X1 U2459 ( .A1(n2293), .A2(n2427), .ZN(n2494) );
  OR2_X1 U2460 ( .A1(n2550), .A2(n2551), .ZN(n2495) );
  AND2_X1 U2461 ( .A1(n2552), .A2(n2553), .ZN(n2551) );
  AND2_X1 U2462 ( .A1(n2554), .A2(n2555), .ZN(n2550) );
  OR2_X1 U2463 ( .A1(n2553), .A2(n2552), .ZN(n2555) );
  XOR2_X1 U2464 ( .A(n2503), .B(n2556), .Z(n2496) );
  XOR2_X1 U2465 ( .A(n2502), .B(n2501), .Z(n2556) );
  OR2_X1 U2466 ( .A1(n2198), .A2(n2274), .ZN(n2501) );
  OR2_X1 U2467 ( .A1(n2557), .A2(n2558), .ZN(n2502) );
  AND2_X1 U2468 ( .A1(n2559), .A2(n2560), .ZN(n2558) );
  AND2_X1 U2469 ( .A1(n2561), .A2(n2562), .ZN(n2557) );
  OR2_X1 U2470 ( .A1(n2560), .A2(n2559), .ZN(n2562) );
  XOR2_X1 U2471 ( .A(n2510), .B(n2563), .Z(n2503) );
  XOR2_X1 U2472 ( .A(n2509), .B(n2508), .Z(n2563) );
  OR2_X1 U2473 ( .A1(n2286), .A2(n2278), .ZN(n2508) );
  OR2_X1 U2474 ( .A1(n2564), .A2(n2565), .ZN(n2509) );
  AND2_X1 U2475 ( .A1(n2566), .A2(n2567), .ZN(n2565) );
  AND2_X1 U2476 ( .A1(n2568), .A2(n2569), .ZN(n2564) );
  OR2_X1 U2477 ( .A1(n2567), .A2(n2566), .ZN(n2569) );
  XOR2_X1 U2478 ( .A(n2516), .B(n2570), .Z(n2510) );
  XOR2_X1 U2479 ( .A(n2515), .B(n2232), .Z(n2570) );
  OR2_X1 U2480 ( .A1(n2235), .A2(n2283), .ZN(n2232) );
  OR2_X1 U2481 ( .A1(n2571), .A2(n2572), .ZN(n2515) );
  AND2_X1 U2482 ( .A1(n2573), .A2(n2574), .ZN(n2572) );
  AND2_X1 U2483 ( .A1(n2575), .A2(n2576), .ZN(n2571) );
  OR2_X1 U2484 ( .A1(n2574), .A2(n2573), .ZN(n2576) );
  XOR2_X1 U2485 ( .A(n2523), .B(n2577), .Z(n2516) );
  XOR2_X1 U2486 ( .A(n2522), .B(n2521), .Z(n2577) );
  OR2_X1 U2487 ( .A1(n2279), .A2(n2285), .ZN(n2521) );
  OR2_X1 U2488 ( .A1(n2578), .A2(n2579), .ZN(n2522) );
  AND2_X1 U2489 ( .A1(n2580), .A2(n2581), .ZN(n2579) );
  AND2_X1 U2490 ( .A1(n2582), .A2(n2583), .ZN(n2578) );
  OR2_X1 U2491 ( .A1(n2581), .A2(n2580), .ZN(n2583) );
  XOR2_X1 U2492 ( .A(n2528), .B(n2584), .Z(n2523) );
  XOR2_X1 U2493 ( .A(n2529), .B(n2531), .Z(n2584) );
  OR2_X1 U2494 ( .A1(n2292), .A2(n2271), .ZN(n2531) );
  OR2_X1 U2495 ( .A1(n2585), .A2(n2586), .ZN(n2529) );
  AND2_X1 U2496 ( .A1(n2587), .A2(n2588), .ZN(n2586) );
  AND2_X1 U2497 ( .A1(n2589), .A2(n2590), .ZN(n2585) );
  OR2_X1 U2498 ( .A1(n2588), .A2(n2587), .ZN(n2589) );
  OR2_X1 U2499 ( .A1(n2275), .A2(n2290), .ZN(n2528) );
  AND2_X1 U2500 ( .A1(n1998), .A2(n1999), .ZN(n2001) );
  XNOR2_X1 U2501 ( .A(n2536), .B(n2537), .ZN(n1999) );
  OR2_X1 U2502 ( .A1(n2591), .A2(n2592), .ZN(n2537) );
  AND2_X1 U2503 ( .A1(n2593), .A2(n2594), .ZN(n2592) );
  AND2_X1 U2504 ( .A1(n2595), .A2(n2596), .ZN(n2591) );
  OR2_X1 U2505 ( .A1(n2594), .A2(n2593), .ZN(n2596) );
  XNOR2_X1 U2506 ( .A(n2547), .B(n2597), .ZN(n2536) );
  XOR2_X1 U2507 ( .A(n2546), .B(n2545), .Z(n2597) );
  OR2_X1 U2508 ( .A1(n2168), .A2(n2427), .ZN(n2545) );
  OR2_X1 U2509 ( .A1(n2598), .A2(n2599), .ZN(n2546) );
  AND2_X1 U2510 ( .A1(n2600), .A2(n2601), .ZN(n2599) );
  AND2_X1 U2511 ( .A1(n2602), .A2(n2603), .ZN(n2598) );
  OR2_X1 U2512 ( .A1(n2601), .A2(n2600), .ZN(n2603) );
  XOR2_X1 U2513 ( .A(n2554), .B(n2604), .Z(n2547) );
  XOR2_X1 U2514 ( .A(n2553), .B(n2552), .Z(n2604) );
  OR2_X1 U2515 ( .A1(n2293), .A2(n2274), .ZN(n2552) );
  OR2_X1 U2516 ( .A1(n2605), .A2(n2606), .ZN(n2553) );
  AND2_X1 U2517 ( .A1(n2607), .A2(n2608), .ZN(n2606) );
  AND2_X1 U2518 ( .A1(n2609), .A2(n2610), .ZN(n2605) );
  OR2_X1 U2519 ( .A1(n2608), .A2(n2607), .ZN(n2610) );
  XOR2_X1 U2520 ( .A(n2561), .B(n2611), .Z(n2554) );
  XOR2_X1 U2521 ( .A(n2560), .B(n2559), .Z(n2611) );
  OR2_X1 U2522 ( .A1(n2198), .A2(n2278), .ZN(n2559) );
  OR2_X1 U2523 ( .A1(n2612), .A2(n2613), .ZN(n2560) );
  AND2_X1 U2524 ( .A1(n2614), .A2(n2615), .ZN(n2613) );
  AND2_X1 U2525 ( .A1(n2616), .A2(n2617), .ZN(n2612) );
  OR2_X1 U2526 ( .A1(n2615), .A2(n2614), .ZN(n2617) );
  XOR2_X1 U2527 ( .A(n2568), .B(n2618), .Z(n2561) );
  XOR2_X1 U2528 ( .A(n2567), .B(n2566), .Z(n2618) );
  OR2_X1 U2529 ( .A1(n2286), .A2(n2283), .ZN(n2566) );
  OR2_X1 U2530 ( .A1(n2619), .A2(n2620), .ZN(n2567) );
  AND2_X1 U2531 ( .A1(n2621), .A2(n2287), .ZN(n2620) );
  AND2_X1 U2532 ( .A1(n2622), .A2(n2623), .ZN(n2619) );
  OR2_X1 U2533 ( .A1(n2287), .A2(n2621), .ZN(n2623) );
  XOR2_X1 U2534 ( .A(n2575), .B(n2624), .Z(n2568) );
  XOR2_X1 U2535 ( .A(n2574), .B(n2573), .Z(n2624) );
  OR2_X1 U2536 ( .A1(n2285), .A2(n2235), .ZN(n2573) );
  OR2_X1 U2537 ( .A1(n2625), .A2(n2626), .ZN(n2574) );
  AND2_X1 U2538 ( .A1(n2627), .A2(n2628), .ZN(n2626) );
  AND2_X1 U2539 ( .A1(n2629), .A2(n2630), .ZN(n2625) );
  OR2_X1 U2540 ( .A1(n2628), .A2(n2627), .ZN(n2630) );
  XOR2_X1 U2541 ( .A(n2582), .B(n2631), .Z(n2575) );
  XOR2_X1 U2542 ( .A(n2581), .B(n2580), .Z(n2631) );
  OR2_X1 U2543 ( .A1(n2279), .A2(n2290), .ZN(n2580) );
  OR2_X1 U2544 ( .A1(n2632), .A2(n2633), .ZN(n2581) );
  AND2_X1 U2545 ( .A1(n2634), .A2(n2635), .ZN(n2633) );
  AND2_X1 U2546 ( .A1(n2636), .A2(n2637), .ZN(n2632) );
  OR2_X1 U2547 ( .A1(n2635), .A2(n2634), .ZN(n2637) );
  XOR2_X1 U2548 ( .A(n2587), .B(n2638), .Z(n2582) );
  XOR2_X1 U2549 ( .A(n2588), .B(n2590), .Z(n2638) );
  OR2_X1 U2550 ( .A1(n2297), .A2(n2271), .ZN(n2590) );
  OR2_X1 U2551 ( .A1(n2639), .A2(n2640), .ZN(n2588) );
  AND2_X1 U2552 ( .A1(n2641), .A2(n2642), .ZN(n2640) );
  AND2_X1 U2553 ( .A1(n2643), .A2(n2644), .ZN(n2639) );
  OR2_X1 U2554 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  OR2_X1 U2555 ( .A1(n2275), .A2(n2292), .ZN(n2587) );
  OR2_X1 U2556 ( .A1(n2645), .A2(n2646), .ZN(n1998) );
  OR2_X1 U2557 ( .A1(n2647), .A2(n1996), .ZN(n2645) );
  AND2_X1 U2558 ( .A1(n1994), .A2(n1995), .ZN(n1996) );
  AND2_X1 U2559 ( .A1(n2648), .A2(n2649), .ZN(n1995) );
  INV_X1 U2560 ( .A(n2650), .ZN(n2648) );
  AND2_X1 U2561 ( .A1(n1994), .A2(n1990), .ZN(n2647) );
  OR2_X1 U2562 ( .A1(n2651), .A2(n2366), .ZN(n1990) );
  AND2_X1 U2563 ( .A1(n2364), .A2(n2652), .ZN(n2366) );
  AND2_X1 U2564 ( .A1(n2365), .A2(n2363), .ZN(n2652) );
  INV_X1 U2565 ( .A(n2653), .ZN(n2364) );
  AND2_X1 U2566 ( .A1(n2363), .A2(n2358), .ZN(n2651) );
  OR2_X1 U2567 ( .A1(n2654), .A2(n2356), .ZN(n2358) );
  AND2_X1 U2568 ( .A1(n2354), .A2(n2655), .ZN(n2356) );
  AND2_X1 U2569 ( .A1(n2355), .A2(n2353), .ZN(n2655) );
  INV_X1 U2570 ( .A(n2656), .ZN(n2354) );
  AND2_X1 U2571 ( .A1(n2353), .A2(n2348), .ZN(n2654) );
  OR2_X1 U2572 ( .A1(n2657), .A2(n2346), .ZN(n2348) );
  AND2_X1 U2573 ( .A1(n2345), .A2(n2344), .ZN(n2346) );
  AND2_X1 U2574 ( .A1(n2345), .A2(n2340), .ZN(n2657) );
  OR2_X1 U2575 ( .A1(n2658), .A2(n2334), .ZN(n2340) );
  AND2_X1 U2576 ( .A1(n2659), .A2(n2660), .ZN(n2334) );
  INV_X1 U2577 ( .A(n2337), .ZN(n2660) );
  OR2_X1 U2578 ( .A1(n2661), .A2(n2662), .ZN(n2337) );
  AND2_X1 U2579 ( .A1(n2338), .A2(n2659), .ZN(n2658) );
  INV_X1 U2580 ( .A(n2336), .ZN(n2659) );
  OR2_X1 U2581 ( .A1(n2663), .A2(n2344), .ZN(n2336) );
  INV_X1 U2582 ( .A(n2664), .ZN(n2344) );
  OR2_X1 U2583 ( .A1(n2665), .A2(n2666), .ZN(n2664) );
  AND2_X1 U2584 ( .A1(n2665), .A2(n2666), .ZN(n2663) );
  OR2_X1 U2585 ( .A1(n2667), .A2(n2668), .ZN(n2666) );
  AND2_X1 U2586 ( .A1(n2669), .A2(n2670), .ZN(n2668) );
  AND2_X1 U2587 ( .A1(n2671), .A2(n2672), .ZN(n2667) );
  OR2_X1 U2588 ( .A1(n2670), .A2(n2669), .ZN(n2672) );
  XOR2_X1 U2589 ( .A(n2673), .B(n2674), .Z(n2665) );
  XOR2_X1 U2590 ( .A(n2675), .B(n2676), .Z(n2674) );
  AND2_X1 U2591 ( .A1(n2331), .A2(n2677), .ZN(n2338) );
  AND2_X1 U2592 ( .A1(n2325), .A2(n2330), .ZN(n2677) );
  XOR2_X1 U2593 ( .A(n2662), .B(n2661), .Z(n2330) );
  OR2_X1 U2594 ( .A1(n2678), .A2(n2679), .ZN(n2661) );
  AND2_X1 U2595 ( .A1(n2680), .A2(n2681), .ZN(n2679) );
  AND2_X1 U2596 ( .A1(n2682), .A2(n2683), .ZN(n2678) );
  OR2_X1 U2597 ( .A1(n2680), .A2(n2681), .ZN(n2683) );
  XOR2_X1 U2598 ( .A(n2671), .B(n2684), .Z(n2662) );
  XOR2_X1 U2599 ( .A(n2670), .B(n2669), .Z(n2684) );
  OR2_X1 U2600 ( .A1(n2078), .A2(n2427), .ZN(n2669) );
  OR2_X1 U2601 ( .A1(n2685), .A2(n2686), .ZN(n2670) );
  AND2_X1 U2602 ( .A1(n2687), .A2(n2688), .ZN(n2686) );
  AND2_X1 U2603 ( .A1(n2689), .A2(n2690), .ZN(n2685) );
  OR2_X1 U2604 ( .A1(n2688), .A2(n2687), .ZN(n2690) );
  XOR2_X1 U2605 ( .A(n2691), .B(n2692), .Z(n2671) );
  XOR2_X1 U2606 ( .A(n2693), .B(n2694), .Z(n2692) );
  XNOR2_X1 U2607 ( .A(n2682), .B(n2695), .ZN(n2325) );
  XOR2_X1 U2608 ( .A(n2681), .B(n2680), .Z(n2695) );
  OR2_X1 U2609 ( .A1(n2049), .A2(n2427), .ZN(n2680) );
  OR2_X1 U2610 ( .A1(n2696), .A2(n2697), .ZN(n2681) );
  AND2_X1 U2611 ( .A1(n2698), .A2(n2699), .ZN(n2697) );
  AND2_X1 U2612 ( .A1(n2700), .A2(n2701), .ZN(n2696) );
  OR2_X1 U2613 ( .A1(n2699), .A2(n2698), .ZN(n2701) );
  XOR2_X1 U2614 ( .A(n2689), .B(n2702), .Z(n2682) );
  XOR2_X1 U2615 ( .A(n2688), .B(n2687), .Z(n2702) );
  OR2_X1 U2616 ( .A1(n2078), .A2(n2274), .ZN(n2687) );
  OR2_X1 U2617 ( .A1(n2703), .A2(n2704), .ZN(n2688) );
  AND2_X1 U2618 ( .A1(n2705), .A2(n2706), .ZN(n2704) );
  AND2_X1 U2619 ( .A1(n2707), .A2(n2708), .ZN(n2703) );
  OR2_X1 U2620 ( .A1(n2706), .A2(n2705), .ZN(n2708) );
  XOR2_X1 U2621 ( .A(n2709), .B(n2710), .Z(n2689) );
  XOR2_X1 U2622 ( .A(n2711), .B(n2712), .Z(n2710) );
  INV_X1 U2623 ( .A(n2324), .ZN(n2331) );
  OR2_X1 U2624 ( .A1(n2713), .A2(n2714), .ZN(n2324) );
  AND2_X1 U2625 ( .A1(n2267), .A2(n2266), .ZN(n2714) );
  AND2_X1 U2626 ( .A1(n2264), .A2(n2715), .ZN(n2713) );
  OR2_X1 U2627 ( .A1(n2267), .A2(n2266), .ZN(n2715) );
  OR2_X1 U2628 ( .A1(n2716), .A2(n2717), .ZN(n2266) );
  AND2_X1 U2629 ( .A1(n2254), .A2(n2253), .ZN(n2717) );
  AND2_X1 U2630 ( .A1(n2251), .A2(n2718), .ZN(n2716) );
  OR2_X1 U2631 ( .A1(n2254), .A2(n2253), .ZN(n2718) );
  OR2_X1 U2632 ( .A1(n2719), .A2(n2720), .ZN(n2253) );
  AND2_X1 U2633 ( .A1(n2242), .A2(n2241), .ZN(n2720) );
  AND2_X1 U2634 ( .A1(n2239), .A2(n2721), .ZN(n2719) );
  OR2_X1 U2635 ( .A1(n2242), .A2(n2241), .ZN(n2721) );
  OR2_X1 U2636 ( .A1(n2722), .A2(n2723), .ZN(n2241) );
  AND2_X1 U2637 ( .A1(n2224), .A2(n2223), .ZN(n2723) );
  AND2_X1 U2638 ( .A1(n2221), .A2(n2724), .ZN(n2722) );
  OR2_X1 U2639 ( .A1(n2224), .A2(n2223), .ZN(n2724) );
  OR2_X1 U2640 ( .A1(n2725), .A2(n2726), .ZN(n2223) );
  AND2_X1 U2641 ( .A1(n2205), .A2(n2204), .ZN(n2726) );
  AND2_X1 U2642 ( .A1(n2202), .A2(n2727), .ZN(n2725) );
  OR2_X1 U2643 ( .A1(n2205), .A2(n2204), .ZN(n2727) );
  OR2_X1 U2644 ( .A1(n2728), .A2(n2729), .ZN(n2204) );
  AND2_X1 U2645 ( .A1(n2187), .A2(n2186), .ZN(n2729) );
  AND2_X1 U2646 ( .A1(n2184), .A2(n2730), .ZN(n2728) );
  OR2_X1 U2647 ( .A1(n2187), .A2(n2186), .ZN(n2730) );
  OR2_X1 U2648 ( .A1(n2731), .A2(n2732), .ZN(n2186) );
  AND2_X1 U2649 ( .A1(n2175), .A2(n2174), .ZN(n2732) );
  AND2_X1 U2650 ( .A1(n2172), .A2(n2733), .ZN(n2731) );
  OR2_X1 U2651 ( .A1(n2175), .A2(n2174), .ZN(n2733) );
  OR2_X1 U2652 ( .A1(n2734), .A2(n2735), .ZN(n2174) );
  AND2_X1 U2653 ( .A1(n2157), .A2(n2156), .ZN(n2735) );
  AND2_X1 U2654 ( .A1(n2154), .A2(n2736), .ZN(n2734) );
  OR2_X1 U2655 ( .A1(n2157), .A2(n2156), .ZN(n2736) );
  OR2_X1 U2656 ( .A1(n2737), .A2(n2738), .ZN(n2156) );
  AND2_X1 U2657 ( .A1(n2145), .A2(n2144), .ZN(n2738) );
  AND2_X1 U2658 ( .A1(n2142), .A2(n2739), .ZN(n2737) );
  OR2_X1 U2659 ( .A1(n2145), .A2(n2144), .ZN(n2739) );
  OR2_X1 U2660 ( .A1(n2740), .A2(n2741), .ZN(n2144) );
  AND2_X1 U2661 ( .A1(n2127), .A2(n2126), .ZN(n2741) );
  AND2_X1 U2662 ( .A1(n2124), .A2(n2742), .ZN(n2740) );
  OR2_X1 U2663 ( .A1(n2127), .A2(n2126), .ZN(n2742) );
  OR2_X1 U2664 ( .A1(n2743), .A2(n2744), .ZN(n2126) );
  AND2_X1 U2665 ( .A1(n2115), .A2(n2114), .ZN(n2744) );
  AND2_X1 U2666 ( .A1(n2112), .A2(n2745), .ZN(n2743) );
  OR2_X1 U2667 ( .A1(n2115), .A2(n2114), .ZN(n2745) );
  OR2_X1 U2668 ( .A1(n2746), .A2(n2747), .ZN(n2114) );
  AND2_X1 U2669 ( .A1(n2097), .A2(n2096), .ZN(n2747) );
  AND2_X1 U2670 ( .A1(n2094), .A2(n2748), .ZN(n2746) );
  OR2_X1 U2671 ( .A1(n2097), .A2(n2096), .ZN(n2748) );
  OR2_X1 U2672 ( .A1(n2749), .A2(n2750), .ZN(n2096) );
  AND2_X1 U2673 ( .A1(n2085), .A2(n2084), .ZN(n2750) );
  AND2_X1 U2674 ( .A1(n2082), .A2(n2751), .ZN(n2749) );
  OR2_X1 U2675 ( .A1(n2085), .A2(n2084), .ZN(n2751) );
  OR2_X1 U2676 ( .A1(n2752), .A2(n2753), .ZN(n2084) );
  AND2_X1 U2677 ( .A1(n2064), .A2(n2067), .ZN(n2753) );
  AND2_X1 U2678 ( .A1(n2066), .A2(n2754), .ZN(n2752) );
  OR2_X1 U2679 ( .A1(n2064), .A2(n2067), .ZN(n2754) );
  OR2_X1 U2680 ( .A1(n2318), .A2(n2035), .ZN(n2067) );
  OR2_X1 U2681 ( .A1(n2049), .A2(n2319), .ZN(n2064) );
  OR2_X1 U2682 ( .A1(n2035), .A2(n2755), .ZN(n2319) );
  INV_X1 U2683 ( .A(n2756), .ZN(n2066) );
  OR2_X1 U2684 ( .A1(n2757), .A2(n2758), .ZN(n2756) );
  AND2_X1 U2685 ( .A1(b_14_), .A2(n2759), .ZN(n2758) );
  OR2_X1 U2686 ( .A1(n2760), .A2(n2043), .ZN(n2759) );
  AND2_X1 U2687 ( .A1(a_14_), .A2(n2078), .ZN(n2760) );
  AND2_X1 U2688 ( .A1(b_13_), .A2(n2761), .ZN(n2757) );
  OR2_X1 U2689 ( .A1(n2762), .A2(n2056), .ZN(n2761) );
  AND2_X1 U2690 ( .A1(a_15_), .A2(n2049), .ZN(n2762) );
  OR2_X1 U2691 ( .A1(n2313), .A2(n2035), .ZN(n2085) );
  XNOR2_X1 U2692 ( .A(n2763), .B(n2764), .ZN(n2082) );
  XNOR2_X1 U2693 ( .A(n2765), .B(n2766), .ZN(n2764) );
  OR2_X1 U2694 ( .A1(n2311), .A2(n2035), .ZN(n2097) );
  XNOR2_X1 U2695 ( .A(n2767), .B(n2768), .ZN(n2094) );
  XNOR2_X1 U2696 ( .A(n2769), .B(n2770), .ZN(n2767) );
  OR2_X1 U2697 ( .A1(n2306), .A2(n2035), .ZN(n2115) );
  XOR2_X1 U2698 ( .A(n2771), .B(n2772), .Z(n2112) );
  XOR2_X1 U2699 ( .A(n2773), .B(n2774), .Z(n2772) );
  OR2_X1 U2700 ( .A1(n2304), .A2(n2035), .ZN(n2127) );
  XOR2_X1 U2701 ( .A(n2775), .B(n2776), .Z(n2124) );
  XOR2_X1 U2702 ( .A(n2777), .B(n2778), .Z(n2776) );
  OR2_X1 U2703 ( .A1(n2299), .A2(n2035), .ZN(n2145) );
  XOR2_X1 U2704 ( .A(n2779), .B(n2780), .Z(n2142) );
  XOR2_X1 U2705 ( .A(n2781), .B(n2782), .Z(n2780) );
  OR2_X1 U2706 ( .A1(n2297), .A2(n2035), .ZN(n2157) );
  XOR2_X1 U2707 ( .A(n2783), .B(n2784), .Z(n2154) );
  XOR2_X1 U2708 ( .A(n2785), .B(n2786), .Z(n2784) );
  OR2_X1 U2709 ( .A1(n2292), .A2(n2035), .ZN(n2175) );
  XOR2_X1 U2710 ( .A(n2787), .B(n2788), .Z(n2172) );
  XOR2_X1 U2711 ( .A(n2789), .B(n2790), .Z(n2788) );
  OR2_X1 U2712 ( .A1(n2290), .A2(n2035), .ZN(n2187) );
  XOR2_X1 U2713 ( .A(n2791), .B(n2792), .Z(n2184) );
  XOR2_X1 U2714 ( .A(n2793), .B(n2794), .Z(n2792) );
  OR2_X1 U2715 ( .A1(n2285), .A2(n2035), .ZN(n2205) );
  XOR2_X1 U2716 ( .A(n2795), .B(n2796), .Z(n2202) );
  XOR2_X1 U2717 ( .A(n2797), .B(n2798), .Z(n2796) );
  OR2_X1 U2718 ( .A1(n2283), .A2(n2035), .ZN(n2224) );
  XOR2_X1 U2719 ( .A(n2799), .B(n2800), .Z(n2221) );
  XOR2_X1 U2720 ( .A(n2801), .B(n2802), .Z(n2800) );
  OR2_X1 U2721 ( .A1(n2278), .A2(n2035), .ZN(n2242) );
  XOR2_X1 U2722 ( .A(n2803), .B(n2804), .Z(n2239) );
  XOR2_X1 U2723 ( .A(n2805), .B(n2806), .Z(n2804) );
  OR2_X1 U2724 ( .A1(n2274), .A2(n2035), .ZN(n2254) );
  XOR2_X1 U2725 ( .A(n2807), .B(n2808), .Z(n2251) );
  XOR2_X1 U2726 ( .A(n2809), .B(n2810), .Z(n2808) );
  OR2_X1 U2727 ( .A1(n2427), .A2(n2035), .ZN(n2267) );
  INV_X1 U2728 ( .A(b_15_), .ZN(n2035) );
  XOR2_X1 U2729 ( .A(n2700), .B(n2811), .Z(n2264) );
  XOR2_X1 U2730 ( .A(n2699), .B(n2698), .Z(n2811) );
  OR2_X1 U2731 ( .A1(n2049), .A2(n2274), .ZN(n2698) );
  OR2_X1 U2732 ( .A1(n2812), .A2(n2813), .ZN(n2699) );
  AND2_X1 U2733 ( .A1(n2810), .A2(n2809), .ZN(n2813) );
  AND2_X1 U2734 ( .A1(n2807), .A2(n2814), .ZN(n2812) );
  OR2_X1 U2735 ( .A1(n2809), .A2(n2810), .ZN(n2814) );
  OR2_X1 U2736 ( .A1(n2049), .A2(n2278), .ZN(n2810) );
  OR2_X1 U2737 ( .A1(n2815), .A2(n2816), .ZN(n2809) );
  AND2_X1 U2738 ( .A1(n2806), .A2(n2805), .ZN(n2816) );
  AND2_X1 U2739 ( .A1(n2803), .A2(n2817), .ZN(n2815) );
  OR2_X1 U2740 ( .A1(n2805), .A2(n2806), .ZN(n2817) );
  OR2_X1 U2741 ( .A1(n2049), .A2(n2283), .ZN(n2806) );
  OR2_X1 U2742 ( .A1(n2818), .A2(n2819), .ZN(n2805) );
  AND2_X1 U2743 ( .A1(n2802), .A2(n2801), .ZN(n2819) );
  AND2_X1 U2744 ( .A1(n2799), .A2(n2820), .ZN(n2818) );
  OR2_X1 U2745 ( .A1(n2801), .A2(n2802), .ZN(n2820) );
  OR2_X1 U2746 ( .A1(n2049), .A2(n2285), .ZN(n2802) );
  OR2_X1 U2747 ( .A1(n2821), .A2(n2822), .ZN(n2801) );
  AND2_X1 U2748 ( .A1(n2798), .A2(n2797), .ZN(n2822) );
  AND2_X1 U2749 ( .A1(n2795), .A2(n2823), .ZN(n2821) );
  OR2_X1 U2750 ( .A1(n2797), .A2(n2798), .ZN(n2823) );
  OR2_X1 U2751 ( .A1(n2049), .A2(n2290), .ZN(n2798) );
  OR2_X1 U2752 ( .A1(n2824), .A2(n2825), .ZN(n2797) );
  AND2_X1 U2753 ( .A1(n2794), .A2(n2793), .ZN(n2825) );
  AND2_X1 U2754 ( .A1(n2791), .A2(n2826), .ZN(n2824) );
  OR2_X1 U2755 ( .A1(n2793), .A2(n2794), .ZN(n2826) );
  OR2_X1 U2756 ( .A1(n2049), .A2(n2292), .ZN(n2794) );
  OR2_X1 U2757 ( .A1(n2827), .A2(n2828), .ZN(n2793) );
  AND2_X1 U2758 ( .A1(n2790), .A2(n2789), .ZN(n2828) );
  AND2_X1 U2759 ( .A1(n2787), .A2(n2829), .ZN(n2827) );
  OR2_X1 U2760 ( .A1(n2789), .A2(n2790), .ZN(n2829) );
  OR2_X1 U2761 ( .A1(n2049), .A2(n2297), .ZN(n2790) );
  OR2_X1 U2762 ( .A1(n2830), .A2(n2831), .ZN(n2789) );
  AND2_X1 U2763 ( .A1(n2786), .A2(n2785), .ZN(n2831) );
  AND2_X1 U2764 ( .A1(n2783), .A2(n2832), .ZN(n2830) );
  OR2_X1 U2765 ( .A1(n2785), .A2(n2786), .ZN(n2832) );
  OR2_X1 U2766 ( .A1(n2049), .A2(n2299), .ZN(n2786) );
  OR2_X1 U2767 ( .A1(n2833), .A2(n2834), .ZN(n2785) );
  AND2_X1 U2768 ( .A1(n2782), .A2(n2781), .ZN(n2834) );
  AND2_X1 U2769 ( .A1(n2779), .A2(n2835), .ZN(n2833) );
  OR2_X1 U2770 ( .A1(n2781), .A2(n2782), .ZN(n2835) );
  OR2_X1 U2771 ( .A1(n2049), .A2(n2304), .ZN(n2782) );
  OR2_X1 U2772 ( .A1(n2836), .A2(n2837), .ZN(n2781) );
  AND2_X1 U2773 ( .A1(n2778), .A2(n2777), .ZN(n2837) );
  AND2_X1 U2774 ( .A1(n2775), .A2(n2838), .ZN(n2836) );
  OR2_X1 U2775 ( .A1(n2777), .A2(n2778), .ZN(n2838) );
  OR2_X1 U2776 ( .A1(n2049), .A2(n2306), .ZN(n2778) );
  OR2_X1 U2777 ( .A1(n2839), .A2(n2840), .ZN(n2777) );
  AND2_X1 U2778 ( .A1(n2774), .A2(n2773), .ZN(n2840) );
  AND2_X1 U2779 ( .A1(n2771), .A2(n2841), .ZN(n2839) );
  OR2_X1 U2780 ( .A1(n2773), .A2(n2774), .ZN(n2841) );
  OR2_X1 U2781 ( .A1(n2049), .A2(n2311), .ZN(n2774) );
  OR2_X1 U2782 ( .A1(n2842), .A2(n2843), .ZN(n2773) );
  AND2_X1 U2783 ( .A1(n2770), .A2(n2769), .ZN(n2843) );
  AND2_X1 U2784 ( .A1(n2768), .A2(n2844), .ZN(n2842) );
  OR2_X1 U2785 ( .A1(n2769), .A2(n2770), .ZN(n2844) );
  OR2_X1 U2786 ( .A1(n2049), .A2(n2313), .ZN(n2770) );
  OR2_X1 U2787 ( .A1(n2845), .A2(n2846), .ZN(n2769) );
  AND2_X1 U2788 ( .A1(n2763), .A2(n2766), .ZN(n2846) );
  AND2_X1 U2789 ( .A1(n2765), .A2(n2847), .ZN(n2845) );
  OR2_X1 U2790 ( .A1(n2766), .A2(n2763), .ZN(n2847) );
  OR2_X1 U2791 ( .A1(n2049), .A2(n2318), .ZN(n2763) );
  OR2_X1 U2792 ( .A1(n2755), .A2(n2848), .ZN(n2766) );
  OR2_X1 U2793 ( .A1(n2049), .A2(n2078), .ZN(n2848) );
  INV_X1 U2794 ( .A(n2849), .ZN(n2765) );
  OR2_X1 U2795 ( .A1(n2850), .A2(n2851), .ZN(n2849) );
  AND2_X1 U2796 ( .A1(b_13_), .A2(n2852), .ZN(n2851) );
  OR2_X1 U2797 ( .A1(n2853), .A2(n2043), .ZN(n2852) );
  AND2_X1 U2798 ( .A1(a_14_), .A2(n2314), .ZN(n2853) );
  AND2_X1 U2799 ( .A1(b_12_), .A2(n2854), .ZN(n2850) );
  OR2_X1 U2800 ( .A1(n2855), .A2(n2056), .ZN(n2854) );
  AND2_X1 U2801 ( .A1(a_15_), .A2(n2078), .ZN(n2855) );
  XNOR2_X1 U2802 ( .A(n2076), .B(n2856), .ZN(n2768) );
  XNOR2_X1 U2803 ( .A(n2857), .B(n2858), .ZN(n2856) );
  XNOR2_X1 U2804 ( .A(n2859), .B(n2860), .ZN(n2771) );
  XNOR2_X1 U2805 ( .A(n2861), .B(n2862), .ZN(n2859) );
  XOR2_X1 U2806 ( .A(n2863), .B(n2864), .Z(n2775) );
  XOR2_X1 U2807 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR2_X1 U2808 ( .A(n2867), .B(n2868), .Z(n2779) );
  XOR2_X1 U2809 ( .A(n2869), .B(n2870), .Z(n2868) );
  XOR2_X1 U2810 ( .A(n2871), .B(n2872), .Z(n2783) );
  XOR2_X1 U2811 ( .A(n2873), .B(n2874), .Z(n2872) );
  XOR2_X1 U2812 ( .A(n2875), .B(n2876), .Z(n2787) );
  XOR2_X1 U2813 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR2_X1 U2814 ( .A(n2879), .B(n2880), .Z(n2791) );
  XOR2_X1 U2815 ( .A(n2881), .B(n2882), .Z(n2880) );
  XOR2_X1 U2816 ( .A(n2883), .B(n2884), .Z(n2795) );
  XOR2_X1 U2817 ( .A(n2885), .B(n2886), .Z(n2884) );
  XOR2_X1 U2818 ( .A(n2887), .B(n2888), .Z(n2799) );
  XOR2_X1 U2819 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR2_X1 U2820 ( .A(n2891), .B(n2892), .Z(n2803) );
  XOR2_X1 U2821 ( .A(n2893), .B(n2894), .Z(n2892) );
  XOR2_X1 U2822 ( .A(n2895), .B(n2896), .Z(n2807) );
  XOR2_X1 U2823 ( .A(n2897), .B(n2898), .Z(n2896) );
  XOR2_X1 U2824 ( .A(n2707), .B(n2899), .Z(n2700) );
  XOR2_X1 U2825 ( .A(n2706), .B(n2705), .Z(n2899) );
  OR2_X1 U2826 ( .A1(n2078), .A2(n2278), .ZN(n2705) );
  OR2_X1 U2827 ( .A1(n2900), .A2(n2901), .ZN(n2706) );
  AND2_X1 U2828 ( .A1(n2898), .A2(n2897), .ZN(n2901) );
  AND2_X1 U2829 ( .A1(n2895), .A2(n2902), .ZN(n2900) );
  OR2_X1 U2830 ( .A1(n2897), .A2(n2898), .ZN(n2902) );
  OR2_X1 U2831 ( .A1(n2078), .A2(n2283), .ZN(n2898) );
  OR2_X1 U2832 ( .A1(n2903), .A2(n2904), .ZN(n2897) );
  AND2_X1 U2833 ( .A1(n2894), .A2(n2893), .ZN(n2904) );
  AND2_X1 U2834 ( .A1(n2891), .A2(n2905), .ZN(n2903) );
  OR2_X1 U2835 ( .A1(n2893), .A2(n2894), .ZN(n2905) );
  OR2_X1 U2836 ( .A1(n2078), .A2(n2285), .ZN(n2894) );
  OR2_X1 U2837 ( .A1(n2906), .A2(n2907), .ZN(n2893) );
  AND2_X1 U2838 ( .A1(n2890), .A2(n2889), .ZN(n2907) );
  AND2_X1 U2839 ( .A1(n2887), .A2(n2908), .ZN(n2906) );
  OR2_X1 U2840 ( .A1(n2889), .A2(n2890), .ZN(n2908) );
  OR2_X1 U2841 ( .A1(n2078), .A2(n2290), .ZN(n2890) );
  OR2_X1 U2842 ( .A1(n2909), .A2(n2910), .ZN(n2889) );
  AND2_X1 U2843 ( .A1(n2886), .A2(n2885), .ZN(n2910) );
  AND2_X1 U2844 ( .A1(n2883), .A2(n2911), .ZN(n2909) );
  OR2_X1 U2845 ( .A1(n2885), .A2(n2886), .ZN(n2911) );
  OR2_X1 U2846 ( .A1(n2078), .A2(n2292), .ZN(n2886) );
  OR2_X1 U2847 ( .A1(n2912), .A2(n2913), .ZN(n2885) );
  AND2_X1 U2848 ( .A1(n2882), .A2(n2881), .ZN(n2913) );
  AND2_X1 U2849 ( .A1(n2879), .A2(n2914), .ZN(n2912) );
  OR2_X1 U2850 ( .A1(n2881), .A2(n2882), .ZN(n2914) );
  OR2_X1 U2851 ( .A1(n2078), .A2(n2297), .ZN(n2882) );
  OR2_X1 U2852 ( .A1(n2915), .A2(n2916), .ZN(n2881) );
  AND2_X1 U2853 ( .A1(n2878), .A2(n2877), .ZN(n2916) );
  AND2_X1 U2854 ( .A1(n2875), .A2(n2917), .ZN(n2915) );
  OR2_X1 U2855 ( .A1(n2877), .A2(n2878), .ZN(n2917) );
  OR2_X1 U2856 ( .A1(n2078), .A2(n2299), .ZN(n2878) );
  OR2_X1 U2857 ( .A1(n2918), .A2(n2919), .ZN(n2877) );
  AND2_X1 U2858 ( .A1(n2874), .A2(n2873), .ZN(n2919) );
  AND2_X1 U2859 ( .A1(n2871), .A2(n2920), .ZN(n2918) );
  OR2_X1 U2860 ( .A1(n2873), .A2(n2874), .ZN(n2920) );
  OR2_X1 U2861 ( .A1(n2078), .A2(n2304), .ZN(n2874) );
  OR2_X1 U2862 ( .A1(n2921), .A2(n2922), .ZN(n2873) );
  AND2_X1 U2863 ( .A1(n2870), .A2(n2869), .ZN(n2922) );
  AND2_X1 U2864 ( .A1(n2867), .A2(n2923), .ZN(n2921) );
  OR2_X1 U2865 ( .A1(n2869), .A2(n2870), .ZN(n2923) );
  OR2_X1 U2866 ( .A1(n2078), .A2(n2306), .ZN(n2870) );
  OR2_X1 U2867 ( .A1(n2924), .A2(n2925), .ZN(n2869) );
  AND2_X1 U2868 ( .A1(n2866), .A2(n2865), .ZN(n2925) );
  AND2_X1 U2869 ( .A1(n2863), .A2(n2926), .ZN(n2924) );
  OR2_X1 U2870 ( .A1(n2865), .A2(n2866), .ZN(n2926) );
  OR2_X1 U2871 ( .A1(n2078), .A2(n2311), .ZN(n2866) );
  OR2_X1 U2872 ( .A1(n2927), .A2(n2928), .ZN(n2865) );
  AND2_X1 U2873 ( .A1(n2862), .A2(n2861), .ZN(n2928) );
  AND2_X1 U2874 ( .A1(n2860), .A2(n2929), .ZN(n2927) );
  OR2_X1 U2875 ( .A1(n2861), .A2(n2862), .ZN(n2929) );
  OR2_X1 U2876 ( .A1(n2078), .A2(n2313), .ZN(n2862) );
  OR2_X1 U2877 ( .A1(n2930), .A2(n2931), .ZN(n2861) );
  AND2_X1 U2878 ( .A1(n2076), .A2(n2858), .ZN(n2931) );
  AND2_X1 U2879 ( .A1(n2857), .A2(n2932), .ZN(n2930) );
  OR2_X1 U2880 ( .A1(n2858), .A2(n2076), .ZN(n2932) );
  OR2_X1 U2881 ( .A1(n2078), .A2(n2318), .ZN(n2076) );
  OR2_X1 U2882 ( .A1(n2755), .A2(n2933), .ZN(n2858) );
  OR2_X1 U2883 ( .A1(n2078), .A2(n2314), .ZN(n2933) );
  INV_X1 U2884 ( .A(b_13_), .ZN(n2078) );
  INV_X1 U2885 ( .A(n2934), .ZN(n2857) );
  OR2_X1 U2886 ( .A1(n2935), .A2(n2936), .ZN(n2934) );
  AND2_X1 U2887 ( .A1(b_12_), .A2(n2937), .ZN(n2936) );
  OR2_X1 U2888 ( .A1(n2938), .A2(n2043), .ZN(n2937) );
  AND2_X1 U2889 ( .A1(a_14_), .A2(n2108), .ZN(n2938) );
  AND2_X1 U2890 ( .A1(b_11_), .A2(n2939), .ZN(n2935) );
  OR2_X1 U2891 ( .A1(n2940), .A2(n2056), .ZN(n2939) );
  AND2_X1 U2892 ( .A1(a_15_), .A2(n2314), .ZN(n2940) );
  XNOR2_X1 U2893 ( .A(n2941), .B(n2942), .ZN(n2860) );
  XNOR2_X1 U2894 ( .A(n2943), .B(n2944), .ZN(n2942) );
  XNOR2_X1 U2895 ( .A(n2945), .B(n2946), .ZN(n2863) );
  XNOR2_X1 U2896 ( .A(n2947), .B(n2315), .ZN(n2945) );
  XOR2_X1 U2897 ( .A(n2948), .B(n2949), .Z(n2867) );
  XOR2_X1 U2898 ( .A(n2950), .B(n2951), .Z(n2949) );
  XOR2_X1 U2899 ( .A(n2952), .B(n2953), .Z(n2871) );
  XOR2_X1 U2900 ( .A(n2954), .B(n2955), .Z(n2953) );
  XOR2_X1 U2901 ( .A(n2956), .B(n2957), .Z(n2875) );
  XOR2_X1 U2902 ( .A(n2958), .B(n2959), .Z(n2957) );
  XOR2_X1 U2903 ( .A(n2960), .B(n2961), .Z(n2879) );
  XOR2_X1 U2904 ( .A(n2962), .B(n2963), .Z(n2961) );
  XOR2_X1 U2905 ( .A(n2964), .B(n2965), .Z(n2883) );
  XOR2_X1 U2906 ( .A(n2966), .B(n2967), .Z(n2965) );
  XOR2_X1 U2907 ( .A(n2968), .B(n2969), .Z(n2887) );
  XOR2_X1 U2908 ( .A(n2970), .B(n2971), .Z(n2969) );
  XOR2_X1 U2909 ( .A(n2972), .B(n2973), .Z(n2891) );
  XOR2_X1 U2910 ( .A(n2974), .B(n2975), .Z(n2973) );
  XOR2_X1 U2911 ( .A(n2976), .B(n2977), .Z(n2895) );
  XOR2_X1 U2912 ( .A(n2978), .B(n2979), .Z(n2977) );
  XOR2_X1 U2913 ( .A(n2980), .B(n2981), .Z(n2707) );
  XOR2_X1 U2914 ( .A(n2982), .B(n2983), .Z(n2981) );
  XNOR2_X1 U2915 ( .A(n2355), .B(n2656), .ZN(n2345) );
  OR2_X1 U2916 ( .A1(n2984), .A2(n2985), .ZN(n2656) );
  AND2_X1 U2917 ( .A1(n2676), .A2(n2675), .ZN(n2985) );
  AND2_X1 U2918 ( .A1(n2673), .A2(n2986), .ZN(n2984) );
  OR2_X1 U2919 ( .A1(n2675), .A2(n2676), .ZN(n2986) );
  OR2_X1 U2920 ( .A1(n2314), .A2(n2427), .ZN(n2676) );
  OR2_X1 U2921 ( .A1(n2987), .A2(n2988), .ZN(n2675) );
  AND2_X1 U2922 ( .A1(n2694), .A2(n2693), .ZN(n2988) );
  AND2_X1 U2923 ( .A1(n2691), .A2(n2989), .ZN(n2987) );
  OR2_X1 U2924 ( .A1(n2693), .A2(n2694), .ZN(n2989) );
  OR2_X1 U2925 ( .A1(n2314), .A2(n2274), .ZN(n2694) );
  OR2_X1 U2926 ( .A1(n2990), .A2(n2991), .ZN(n2693) );
  AND2_X1 U2927 ( .A1(n2712), .A2(n2711), .ZN(n2991) );
  AND2_X1 U2928 ( .A1(n2709), .A2(n2992), .ZN(n2990) );
  OR2_X1 U2929 ( .A1(n2711), .A2(n2712), .ZN(n2992) );
  OR2_X1 U2930 ( .A1(n2314), .A2(n2278), .ZN(n2712) );
  OR2_X1 U2931 ( .A1(n2993), .A2(n2994), .ZN(n2711) );
  AND2_X1 U2932 ( .A1(n2983), .A2(n2982), .ZN(n2994) );
  AND2_X1 U2933 ( .A1(n2980), .A2(n2995), .ZN(n2993) );
  OR2_X1 U2934 ( .A1(n2982), .A2(n2983), .ZN(n2995) );
  OR2_X1 U2935 ( .A1(n2314), .A2(n2283), .ZN(n2983) );
  OR2_X1 U2936 ( .A1(n2996), .A2(n2997), .ZN(n2982) );
  AND2_X1 U2937 ( .A1(n2979), .A2(n2978), .ZN(n2997) );
  AND2_X1 U2938 ( .A1(n2976), .A2(n2998), .ZN(n2996) );
  OR2_X1 U2939 ( .A1(n2978), .A2(n2979), .ZN(n2998) );
  OR2_X1 U2940 ( .A1(n2314), .A2(n2285), .ZN(n2979) );
  OR2_X1 U2941 ( .A1(n2999), .A2(n3000), .ZN(n2978) );
  AND2_X1 U2942 ( .A1(n2975), .A2(n2974), .ZN(n3000) );
  AND2_X1 U2943 ( .A1(n2972), .A2(n3001), .ZN(n2999) );
  OR2_X1 U2944 ( .A1(n2974), .A2(n2975), .ZN(n3001) );
  OR2_X1 U2945 ( .A1(n2314), .A2(n2290), .ZN(n2975) );
  OR2_X1 U2946 ( .A1(n3002), .A2(n3003), .ZN(n2974) );
  AND2_X1 U2947 ( .A1(n2971), .A2(n2970), .ZN(n3003) );
  AND2_X1 U2948 ( .A1(n2968), .A2(n3004), .ZN(n3002) );
  OR2_X1 U2949 ( .A1(n2970), .A2(n2971), .ZN(n3004) );
  OR2_X1 U2950 ( .A1(n2314), .A2(n2292), .ZN(n2971) );
  OR2_X1 U2951 ( .A1(n3005), .A2(n3006), .ZN(n2970) );
  AND2_X1 U2952 ( .A1(n2967), .A2(n2966), .ZN(n3006) );
  AND2_X1 U2953 ( .A1(n2964), .A2(n3007), .ZN(n3005) );
  OR2_X1 U2954 ( .A1(n2966), .A2(n2967), .ZN(n3007) );
  OR2_X1 U2955 ( .A1(n2314), .A2(n2297), .ZN(n2967) );
  OR2_X1 U2956 ( .A1(n3008), .A2(n3009), .ZN(n2966) );
  AND2_X1 U2957 ( .A1(n2963), .A2(n2962), .ZN(n3009) );
  AND2_X1 U2958 ( .A1(n2960), .A2(n3010), .ZN(n3008) );
  OR2_X1 U2959 ( .A1(n2962), .A2(n2963), .ZN(n3010) );
  OR2_X1 U2960 ( .A1(n2314), .A2(n2299), .ZN(n2963) );
  OR2_X1 U2961 ( .A1(n3011), .A2(n3012), .ZN(n2962) );
  AND2_X1 U2962 ( .A1(n2959), .A2(n2958), .ZN(n3012) );
  AND2_X1 U2963 ( .A1(n2956), .A2(n3013), .ZN(n3011) );
  OR2_X1 U2964 ( .A1(n2958), .A2(n2959), .ZN(n3013) );
  OR2_X1 U2965 ( .A1(n2314), .A2(n2304), .ZN(n2959) );
  OR2_X1 U2966 ( .A1(n3014), .A2(n3015), .ZN(n2958) );
  AND2_X1 U2967 ( .A1(n2955), .A2(n2954), .ZN(n3015) );
  AND2_X1 U2968 ( .A1(n2952), .A2(n3016), .ZN(n3014) );
  OR2_X1 U2969 ( .A1(n2954), .A2(n2955), .ZN(n3016) );
  OR2_X1 U2970 ( .A1(n2314), .A2(n2306), .ZN(n2955) );
  OR2_X1 U2971 ( .A1(n3017), .A2(n3018), .ZN(n2954) );
  AND2_X1 U2972 ( .A1(n2951), .A2(n2950), .ZN(n3018) );
  AND2_X1 U2973 ( .A1(n2948), .A2(n3019), .ZN(n3017) );
  OR2_X1 U2974 ( .A1(n2950), .A2(n2951), .ZN(n3019) );
  OR2_X1 U2975 ( .A1(n2314), .A2(n2311), .ZN(n2951) );
  OR2_X1 U2976 ( .A1(n3020), .A2(n3021), .ZN(n2950) );
  AND2_X1 U2977 ( .A1(n2315), .A2(n2947), .ZN(n3021) );
  AND2_X1 U2978 ( .A1(n2946), .A2(n3022), .ZN(n3020) );
  OR2_X1 U2979 ( .A1(n2947), .A2(n2315), .ZN(n3022) );
  INV_X1 U2980 ( .A(n2089), .ZN(n2315) );
  AND2_X1 U2981 ( .A1(a_12_), .A2(b_12_), .ZN(n2089) );
  OR2_X1 U2982 ( .A1(n3023), .A2(n3024), .ZN(n2947) );
  AND2_X1 U2983 ( .A1(n2941), .A2(n2944), .ZN(n3024) );
  AND2_X1 U2984 ( .A1(n2943), .A2(n3025), .ZN(n3023) );
  OR2_X1 U2985 ( .A1(n2944), .A2(n2941), .ZN(n3025) );
  OR2_X1 U2986 ( .A1(n2318), .A2(n2314), .ZN(n2941) );
  OR2_X1 U2987 ( .A1(n2755), .A2(n3026), .ZN(n2944) );
  OR2_X1 U2988 ( .A1(n2314), .A2(n2108), .ZN(n3026) );
  INV_X1 U2989 ( .A(b_12_), .ZN(n2314) );
  INV_X1 U2990 ( .A(n3027), .ZN(n2943) );
  OR2_X1 U2991 ( .A1(n3028), .A2(n3029), .ZN(n3027) );
  AND2_X1 U2992 ( .A1(b_11_), .A2(n3030), .ZN(n3029) );
  OR2_X1 U2993 ( .A1(n3031), .A2(n2043), .ZN(n3030) );
  AND2_X1 U2994 ( .A1(a_14_), .A2(n2307), .ZN(n3031) );
  AND2_X1 U2995 ( .A1(b_10_), .A2(n3032), .ZN(n3028) );
  OR2_X1 U2996 ( .A1(n3033), .A2(n2056), .ZN(n3032) );
  AND2_X1 U2997 ( .A1(a_15_), .A2(n2108), .ZN(n3033) );
  XNOR2_X1 U2998 ( .A(n3034), .B(n3035), .ZN(n2946) );
  XNOR2_X1 U2999 ( .A(n3036), .B(n3037), .ZN(n3035) );
  XNOR2_X1 U3000 ( .A(n3038), .B(n3039), .ZN(n2948) );
  XNOR2_X1 U3001 ( .A(n3040), .B(n3041), .ZN(n3038) );
  XOR2_X1 U3002 ( .A(n3042), .B(n3043), .Z(n2952) );
  XOR2_X1 U3003 ( .A(n3044), .B(n2105), .Z(n3043) );
  XOR2_X1 U3004 ( .A(n3045), .B(n3046), .Z(n2956) );
  XOR2_X1 U3005 ( .A(n3047), .B(n3048), .Z(n3046) );
  XOR2_X1 U3006 ( .A(n3049), .B(n3050), .Z(n2960) );
  XOR2_X1 U3007 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR2_X1 U3008 ( .A(n3053), .B(n3054), .Z(n2964) );
  XOR2_X1 U3009 ( .A(n3055), .B(n3056), .Z(n3054) );
  XOR2_X1 U3010 ( .A(n3057), .B(n3058), .Z(n2968) );
  XOR2_X1 U3011 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR2_X1 U3012 ( .A(n3061), .B(n3062), .Z(n2972) );
  XOR2_X1 U3013 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR2_X1 U3014 ( .A(n3065), .B(n3066), .Z(n2976) );
  XOR2_X1 U3015 ( .A(n3067), .B(n3068), .Z(n3066) );
  XOR2_X1 U3016 ( .A(n3069), .B(n3070), .Z(n2980) );
  XOR2_X1 U3017 ( .A(n3071), .B(n3072), .Z(n3070) );
  XOR2_X1 U3018 ( .A(n3073), .B(n3074), .Z(n2709) );
  XOR2_X1 U3019 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR2_X1 U3020 ( .A(n3077), .B(n3078), .Z(n2691) );
  XOR2_X1 U3021 ( .A(n3079), .B(n3080), .Z(n3078) );
  XOR2_X1 U3022 ( .A(n3081), .B(n3082), .Z(n2673) );
  XOR2_X1 U3023 ( .A(n3083), .B(n3084), .Z(n3082) );
  XNOR2_X1 U3024 ( .A(n3085), .B(n3086), .ZN(n2355) );
  XOR2_X1 U3025 ( .A(n3087), .B(n3088), .Z(n3086) );
  XNOR2_X1 U3026 ( .A(n2365), .B(n2653), .ZN(n2353) );
  OR2_X1 U3027 ( .A1(n3089), .A2(n3090), .ZN(n2653) );
  AND2_X1 U3028 ( .A1(n3088), .A2(n3087), .ZN(n3090) );
  AND2_X1 U3029 ( .A1(n3085), .A2(n3091), .ZN(n3089) );
  OR2_X1 U3030 ( .A1(n3087), .A2(n3088), .ZN(n3091) );
  OR2_X1 U3031 ( .A1(n2108), .A2(n2427), .ZN(n3088) );
  OR2_X1 U3032 ( .A1(n3092), .A2(n3093), .ZN(n3087) );
  AND2_X1 U3033 ( .A1(n3084), .A2(n3083), .ZN(n3093) );
  AND2_X1 U3034 ( .A1(n3081), .A2(n3094), .ZN(n3092) );
  OR2_X1 U3035 ( .A1(n3083), .A2(n3084), .ZN(n3094) );
  OR2_X1 U3036 ( .A1(n2108), .A2(n2274), .ZN(n3084) );
  OR2_X1 U3037 ( .A1(n3095), .A2(n3096), .ZN(n3083) );
  AND2_X1 U3038 ( .A1(n3080), .A2(n3079), .ZN(n3096) );
  AND2_X1 U3039 ( .A1(n3077), .A2(n3097), .ZN(n3095) );
  OR2_X1 U3040 ( .A1(n3079), .A2(n3080), .ZN(n3097) );
  OR2_X1 U3041 ( .A1(n2108), .A2(n2278), .ZN(n3080) );
  OR2_X1 U3042 ( .A1(n3098), .A2(n3099), .ZN(n3079) );
  AND2_X1 U3043 ( .A1(n3076), .A2(n3075), .ZN(n3099) );
  AND2_X1 U3044 ( .A1(n3073), .A2(n3100), .ZN(n3098) );
  OR2_X1 U3045 ( .A1(n3075), .A2(n3076), .ZN(n3100) );
  OR2_X1 U3046 ( .A1(n2108), .A2(n2283), .ZN(n3076) );
  OR2_X1 U3047 ( .A1(n3101), .A2(n3102), .ZN(n3075) );
  AND2_X1 U3048 ( .A1(n3072), .A2(n3071), .ZN(n3102) );
  AND2_X1 U3049 ( .A1(n3069), .A2(n3103), .ZN(n3101) );
  OR2_X1 U3050 ( .A1(n3071), .A2(n3072), .ZN(n3103) );
  OR2_X1 U3051 ( .A1(n2108), .A2(n2285), .ZN(n3072) );
  OR2_X1 U3052 ( .A1(n3104), .A2(n3105), .ZN(n3071) );
  AND2_X1 U3053 ( .A1(n3068), .A2(n3067), .ZN(n3105) );
  AND2_X1 U3054 ( .A1(n3065), .A2(n3106), .ZN(n3104) );
  OR2_X1 U3055 ( .A1(n3067), .A2(n3068), .ZN(n3106) );
  OR2_X1 U3056 ( .A1(n2108), .A2(n2290), .ZN(n3068) );
  OR2_X1 U3057 ( .A1(n3107), .A2(n3108), .ZN(n3067) );
  AND2_X1 U3058 ( .A1(n3064), .A2(n3063), .ZN(n3108) );
  AND2_X1 U3059 ( .A1(n3061), .A2(n3109), .ZN(n3107) );
  OR2_X1 U3060 ( .A1(n3063), .A2(n3064), .ZN(n3109) );
  OR2_X1 U3061 ( .A1(n2108), .A2(n2292), .ZN(n3064) );
  OR2_X1 U3062 ( .A1(n3110), .A2(n3111), .ZN(n3063) );
  AND2_X1 U3063 ( .A1(n3060), .A2(n3059), .ZN(n3111) );
  AND2_X1 U3064 ( .A1(n3057), .A2(n3112), .ZN(n3110) );
  OR2_X1 U3065 ( .A1(n3059), .A2(n3060), .ZN(n3112) );
  OR2_X1 U3066 ( .A1(n2108), .A2(n2297), .ZN(n3060) );
  OR2_X1 U3067 ( .A1(n3113), .A2(n3114), .ZN(n3059) );
  AND2_X1 U3068 ( .A1(n3056), .A2(n3055), .ZN(n3114) );
  AND2_X1 U3069 ( .A1(n3053), .A2(n3115), .ZN(n3113) );
  OR2_X1 U3070 ( .A1(n3055), .A2(n3056), .ZN(n3115) );
  OR2_X1 U3071 ( .A1(n2108), .A2(n2299), .ZN(n3056) );
  OR2_X1 U3072 ( .A1(n3116), .A2(n3117), .ZN(n3055) );
  AND2_X1 U3073 ( .A1(n3052), .A2(n3051), .ZN(n3117) );
  AND2_X1 U3074 ( .A1(n3049), .A2(n3118), .ZN(n3116) );
  OR2_X1 U3075 ( .A1(n3051), .A2(n3052), .ZN(n3118) );
  OR2_X1 U3076 ( .A1(n2108), .A2(n2304), .ZN(n3052) );
  OR2_X1 U3077 ( .A1(n3119), .A2(n3120), .ZN(n3051) );
  AND2_X1 U3078 ( .A1(n3048), .A2(n3047), .ZN(n3120) );
  AND2_X1 U3079 ( .A1(n3045), .A2(n3121), .ZN(n3119) );
  OR2_X1 U3080 ( .A1(n3047), .A2(n3048), .ZN(n3121) );
  OR2_X1 U3081 ( .A1(n2108), .A2(n2306), .ZN(n3048) );
  OR2_X1 U3082 ( .A1(n3122), .A2(n3123), .ZN(n3047) );
  AND2_X1 U3083 ( .A1(n2105), .A2(n3044), .ZN(n3123) );
  AND2_X1 U3084 ( .A1(n3042), .A2(n3124), .ZN(n3122) );
  OR2_X1 U3085 ( .A1(n3044), .A2(n2105), .ZN(n3124) );
  OR2_X1 U3086 ( .A1(n2108), .A2(n2311), .ZN(n2105) );
  OR2_X1 U3087 ( .A1(n3125), .A2(n3126), .ZN(n3044) );
  AND2_X1 U3088 ( .A1(n3041), .A2(n3040), .ZN(n3126) );
  AND2_X1 U3089 ( .A1(n3039), .A2(n3127), .ZN(n3125) );
  OR2_X1 U3090 ( .A1(n3040), .A2(n3041), .ZN(n3127) );
  OR2_X1 U3091 ( .A1(n2313), .A2(n2108), .ZN(n3041) );
  OR2_X1 U3092 ( .A1(n3128), .A2(n3129), .ZN(n3040) );
  AND2_X1 U3093 ( .A1(n3034), .A2(n3037), .ZN(n3129) );
  AND2_X1 U3094 ( .A1(n3036), .A2(n3130), .ZN(n3128) );
  OR2_X1 U3095 ( .A1(n3037), .A2(n3034), .ZN(n3130) );
  OR2_X1 U3096 ( .A1(n2318), .A2(n2108), .ZN(n3034) );
  OR2_X1 U3097 ( .A1(n2755), .A2(n3131), .ZN(n3037) );
  OR2_X1 U3098 ( .A1(n2108), .A2(n2307), .ZN(n3131) );
  INV_X1 U3099 ( .A(b_11_), .ZN(n2108) );
  INV_X1 U3100 ( .A(n3132), .ZN(n3036) );
  OR2_X1 U3101 ( .A1(n3133), .A2(n3134), .ZN(n3132) );
  AND2_X1 U3102 ( .A1(b_9_), .A2(n3135), .ZN(n3134) );
  OR2_X1 U3103 ( .A1(n3136), .A2(n2056), .ZN(n3135) );
  AND2_X1 U3104 ( .A1(a_15_), .A2(n2307), .ZN(n3136) );
  AND2_X1 U3105 ( .A1(b_10_), .A2(n3137), .ZN(n3133) );
  OR2_X1 U3106 ( .A1(n3138), .A2(n2043), .ZN(n3137) );
  AND2_X1 U3107 ( .A1(a_14_), .A2(n2138), .ZN(n3138) );
  XNOR2_X1 U3108 ( .A(n3139), .B(n3140), .ZN(n3039) );
  XNOR2_X1 U3109 ( .A(n3141), .B(n3142), .ZN(n3140) );
  XNOR2_X1 U3110 ( .A(n3143), .B(n3144), .ZN(n3042) );
  XNOR2_X1 U3111 ( .A(n3145), .B(n3146), .ZN(n3143) );
  XOR2_X1 U3112 ( .A(n3147), .B(n3148), .Z(n3045) );
  XOR2_X1 U3113 ( .A(n3149), .B(n3150), .Z(n3148) );
  XOR2_X1 U3114 ( .A(n3151), .B(n3152), .Z(n3049) );
  XNOR2_X1 U3115 ( .A(n3153), .B(n2119), .ZN(n3152) );
  XOR2_X1 U3116 ( .A(n3154), .B(n3155), .Z(n3053) );
  XOR2_X1 U3117 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR2_X1 U3118 ( .A(n3158), .B(n3159), .Z(n3057) );
  XOR2_X1 U3119 ( .A(n3160), .B(n3161), .Z(n3159) );
  XOR2_X1 U3120 ( .A(n3162), .B(n3163), .Z(n3061) );
  XOR2_X1 U3121 ( .A(n3164), .B(n3165), .Z(n3163) );
  XOR2_X1 U3122 ( .A(n3166), .B(n3167), .Z(n3065) );
  XOR2_X1 U3123 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR2_X1 U3124 ( .A(n3170), .B(n3171), .Z(n3069) );
  XOR2_X1 U3125 ( .A(n3172), .B(n3173), .Z(n3171) );
  XOR2_X1 U3126 ( .A(n3174), .B(n3175), .Z(n3073) );
  XOR2_X1 U3127 ( .A(n3176), .B(n3177), .Z(n3175) );
  XOR2_X1 U3128 ( .A(n3178), .B(n3179), .Z(n3077) );
  XOR2_X1 U3129 ( .A(n3180), .B(n3181), .Z(n3179) );
  XOR2_X1 U3130 ( .A(n3182), .B(n3183), .Z(n3081) );
  XOR2_X1 U3131 ( .A(n3184), .B(n3185), .Z(n3183) );
  XOR2_X1 U3132 ( .A(n3186), .B(n3187), .Z(n3085) );
  XOR2_X1 U3133 ( .A(n3188), .B(n3189), .Z(n3187) );
  XNOR2_X1 U3134 ( .A(n3190), .B(n3191), .ZN(n2365) );
  XOR2_X1 U3135 ( .A(n3192), .B(n3193), .Z(n3191) );
  XNOR2_X1 U3136 ( .A(n2649), .B(n2650), .ZN(n2363) );
  OR2_X1 U3137 ( .A1(n3194), .A2(n3195), .ZN(n2650) );
  AND2_X1 U3138 ( .A1(n3193), .A2(n3192), .ZN(n3195) );
  AND2_X1 U3139 ( .A1(n3190), .A2(n3196), .ZN(n3194) );
  OR2_X1 U3140 ( .A1(n3192), .A2(n3193), .ZN(n3196) );
  OR2_X1 U3141 ( .A1(n2307), .A2(n2427), .ZN(n3193) );
  OR2_X1 U3142 ( .A1(n3197), .A2(n3198), .ZN(n3192) );
  AND2_X1 U3143 ( .A1(n3189), .A2(n3188), .ZN(n3198) );
  AND2_X1 U3144 ( .A1(n3186), .A2(n3199), .ZN(n3197) );
  OR2_X1 U3145 ( .A1(n3188), .A2(n3189), .ZN(n3199) );
  OR2_X1 U3146 ( .A1(n2307), .A2(n2274), .ZN(n3189) );
  OR2_X1 U3147 ( .A1(n3200), .A2(n3201), .ZN(n3188) );
  AND2_X1 U3148 ( .A1(n3185), .A2(n3184), .ZN(n3201) );
  AND2_X1 U3149 ( .A1(n3182), .A2(n3202), .ZN(n3200) );
  OR2_X1 U3150 ( .A1(n3184), .A2(n3185), .ZN(n3202) );
  OR2_X1 U3151 ( .A1(n2307), .A2(n2278), .ZN(n3185) );
  OR2_X1 U3152 ( .A1(n3203), .A2(n3204), .ZN(n3184) );
  AND2_X1 U3153 ( .A1(n3178), .A2(n3181), .ZN(n3204) );
  AND2_X1 U3154 ( .A1(n3205), .A2(n3180), .ZN(n3203) );
  OR2_X1 U3155 ( .A1(n3206), .A2(n3207), .ZN(n3180) );
  AND2_X1 U3156 ( .A1(n3177), .A2(n3176), .ZN(n3207) );
  AND2_X1 U3157 ( .A1(n3174), .A2(n3208), .ZN(n3206) );
  OR2_X1 U3158 ( .A1(n3176), .A2(n3177), .ZN(n3208) );
  OR2_X1 U3159 ( .A1(n2307), .A2(n2285), .ZN(n3177) );
  OR2_X1 U3160 ( .A1(n3209), .A2(n3210), .ZN(n3176) );
  AND2_X1 U3161 ( .A1(n3170), .A2(n3173), .ZN(n3210) );
  AND2_X1 U3162 ( .A1(n3211), .A2(n3172), .ZN(n3209) );
  OR2_X1 U3163 ( .A1(n3212), .A2(n3213), .ZN(n3172) );
  AND2_X1 U3164 ( .A1(n3166), .A2(n3169), .ZN(n3213) );
  AND2_X1 U3165 ( .A1(n3214), .A2(n3168), .ZN(n3212) );
  OR2_X1 U3166 ( .A1(n3215), .A2(n3216), .ZN(n3168) );
  AND2_X1 U3167 ( .A1(n3162), .A2(n3165), .ZN(n3216) );
  AND2_X1 U3168 ( .A1(n3217), .A2(n3164), .ZN(n3215) );
  OR2_X1 U3169 ( .A1(n3218), .A2(n3219), .ZN(n3164) );
  AND2_X1 U3170 ( .A1(n3158), .A2(n3161), .ZN(n3219) );
  AND2_X1 U3171 ( .A1(n3220), .A2(n3160), .ZN(n3218) );
  OR2_X1 U3172 ( .A1(n3221), .A2(n3222), .ZN(n3160) );
  AND2_X1 U3173 ( .A1(n3154), .A2(n3157), .ZN(n3222) );
  AND2_X1 U3174 ( .A1(n3223), .A2(n3156), .ZN(n3221) );
  OR2_X1 U3175 ( .A1(n3224), .A2(n3225), .ZN(n3156) );
  AND2_X1 U3176 ( .A1(n3151), .A2(n2308), .ZN(n3225) );
  AND2_X1 U3177 ( .A1(n3226), .A2(n3153), .ZN(n3224) );
  OR2_X1 U3178 ( .A1(n3227), .A2(n3228), .ZN(n3153) );
  AND2_X1 U3179 ( .A1(n3147), .A2(n3150), .ZN(n3228) );
  AND2_X1 U3180 ( .A1(n3229), .A2(n3149), .ZN(n3227) );
  OR2_X1 U3181 ( .A1(n3230), .A2(n3231), .ZN(n3149) );
  AND2_X1 U3182 ( .A1(n3144), .A2(n3146), .ZN(n3231) );
  AND2_X1 U3183 ( .A1(n3232), .A2(n3145), .ZN(n3230) );
  OR2_X1 U3184 ( .A1(n3233), .A2(n3234), .ZN(n3145) );
  AND2_X1 U3185 ( .A1(n3139), .A2(n3142), .ZN(n3234) );
  AND2_X1 U3186 ( .A1(n3141), .A2(n3235), .ZN(n3233) );
  OR2_X1 U3187 ( .A1(n3142), .A2(n3139), .ZN(n3235) );
  OR2_X1 U3188 ( .A1(n2318), .A2(n2307), .ZN(n3139) );
  OR2_X1 U3189 ( .A1(n2755), .A2(n3236), .ZN(n3142) );
  OR2_X1 U3190 ( .A1(n2307), .A2(n2138), .ZN(n3236) );
  INV_X1 U3191 ( .A(n3237), .ZN(n3141) );
  OR2_X1 U3192 ( .A1(n3238), .A2(n3239), .ZN(n3237) );
  AND2_X1 U3193 ( .A1(b_9_), .A2(n3240), .ZN(n3239) );
  OR2_X1 U3194 ( .A1(n3241), .A2(n2043), .ZN(n3240) );
  AND2_X1 U3195 ( .A1(a_14_), .A2(n2300), .ZN(n3241) );
  AND2_X1 U3196 ( .A1(b_8_), .A2(n3242), .ZN(n3238) );
  OR2_X1 U3197 ( .A1(n3243), .A2(n2056), .ZN(n3242) );
  AND2_X1 U3198 ( .A1(a_15_), .A2(n2138), .ZN(n3243) );
  OR2_X1 U3199 ( .A1(n3146), .A2(n3144), .ZN(n3232) );
  XNOR2_X1 U3200 ( .A(n3244), .B(n3245), .ZN(n3144) );
  XNOR2_X1 U3201 ( .A(n3246), .B(n3247), .ZN(n3245) );
  OR2_X1 U3202 ( .A1(n2313), .A2(n2307), .ZN(n3146) );
  OR2_X1 U3203 ( .A1(n3150), .A2(n3147), .ZN(n3229) );
  XNOR2_X1 U3204 ( .A(n3248), .B(n3249), .ZN(n3147) );
  XNOR2_X1 U3205 ( .A(n3250), .B(n3251), .ZN(n3248) );
  OR2_X1 U3206 ( .A1(n2311), .A2(n2307), .ZN(n3150) );
  OR2_X1 U3207 ( .A1(n2308), .A2(n3151), .ZN(n3226) );
  XOR2_X1 U3208 ( .A(n3252), .B(n3253), .Z(n3151) );
  XOR2_X1 U3209 ( .A(n3254), .B(n3255), .Z(n3253) );
  INV_X1 U3210 ( .A(n2119), .ZN(n2308) );
  AND2_X1 U3211 ( .A1(a_10_), .A2(b_10_), .ZN(n2119) );
  OR2_X1 U3212 ( .A1(n3157), .A2(n3154), .ZN(n3223) );
  XOR2_X1 U3213 ( .A(n3256), .B(n3257), .Z(n3154) );
  XOR2_X1 U3214 ( .A(n3258), .B(n3259), .Z(n3257) );
  OR2_X1 U3215 ( .A1(n2307), .A2(n2304), .ZN(n3157) );
  OR2_X1 U3216 ( .A1(n3161), .A2(n3158), .ZN(n3220) );
  XOR2_X1 U3217 ( .A(n3260), .B(n3261), .Z(n3158) );
  XOR2_X1 U3218 ( .A(n3262), .B(n2135), .Z(n3261) );
  OR2_X1 U3219 ( .A1(n2307), .A2(n2299), .ZN(n3161) );
  OR2_X1 U3220 ( .A1(n3165), .A2(n3162), .ZN(n3217) );
  XOR2_X1 U3221 ( .A(n3263), .B(n3264), .Z(n3162) );
  XOR2_X1 U3222 ( .A(n3265), .B(n3266), .Z(n3264) );
  OR2_X1 U3223 ( .A1(n2307), .A2(n2297), .ZN(n3165) );
  OR2_X1 U3224 ( .A1(n3169), .A2(n3166), .ZN(n3214) );
  XOR2_X1 U3225 ( .A(n3267), .B(n3268), .Z(n3166) );
  XOR2_X1 U3226 ( .A(n3269), .B(n3270), .Z(n3268) );
  OR2_X1 U3227 ( .A1(n2307), .A2(n2292), .ZN(n3169) );
  OR2_X1 U3228 ( .A1(n3173), .A2(n3170), .ZN(n3211) );
  XOR2_X1 U3229 ( .A(n3271), .B(n3272), .Z(n3170) );
  XOR2_X1 U3230 ( .A(n3273), .B(n3274), .Z(n3272) );
  OR2_X1 U3231 ( .A1(n2307), .A2(n2290), .ZN(n3173) );
  XOR2_X1 U3232 ( .A(n3275), .B(n3276), .Z(n3174) );
  XOR2_X1 U3233 ( .A(n3277), .B(n3278), .Z(n3276) );
  OR2_X1 U3234 ( .A1(n3181), .A2(n3178), .ZN(n3205) );
  XOR2_X1 U3235 ( .A(n3279), .B(n3280), .Z(n3178) );
  XOR2_X1 U3236 ( .A(n3281), .B(n3282), .Z(n3280) );
  OR2_X1 U3237 ( .A1(n2307), .A2(n2283), .ZN(n3181) );
  INV_X1 U3238 ( .A(b_10_), .ZN(n2307) );
  XOR2_X1 U3239 ( .A(n3283), .B(n3284), .Z(n3182) );
  XOR2_X1 U3240 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR2_X1 U3241 ( .A(n3287), .B(n3288), .Z(n3186) );
  XOR2_X1 U3242 ( .A(n3289), .B(n3290), .Z(n3288) );
  XOR2_X1 U3243 ( .A(n3291), .B(n3292), .Z(n3190) );
  XOR2_X1 U3244 ( .A(n3293), .B(n3294), .Z(n3292) );
  XNOR2_X1 U3245 ( .A(n3295), .B(n3296), .ZN(n2649) );
  XOR2_X1 U3246 ( .A(n3297), .B(n3298), .Z(n3296) );
  INV_X1 U3247 ( .A(n3299), .ZN(n1994) );
  OR2_X1 U3248 ( .A1(n3300), .A2(n2646), .ZN(n3299) );
  INV_X1 U3249 ( .A(n3301), .ZN(n2646) );
  OR2_X1 U3250 ( .A1(n3302), .A2(n3303), .ZN(n3301) );
  AND2_X1 U3251 ( .A1(n3302), .A2(n3303), .ZN(n3300) );
  OR2_X1 U3252 ( .A1(n3304), .A2(n3305), .ZN(n3303) );
  AND2_X1 U3253 ( .A1(n3298), .A2(n3297), .ZN(n3305) );
  AND2_X1 U3254 ( .A1(n3295), .A2(n3306), .ZN(n3304) );
  OR2_X1 U3255 ( .A1(n3297), .A2(n3298), .ZN(n3306) );
  OR2_X1 U3256 ( .A1(n2138), .A2(n2427), .ZN(n3298) );
  OR2_X1 U3257 ( .A1(n3307), .A2(n3308), .ZN(n3297) );
  AND2_X1 U3258 ( .A1(n3294), .A2(n3293), .ZN(n3308) );
  AND2_X1 U3259 ( .A1(n3291), .A2(n3309), .ZN(n3307) );
  OR2_X1 U3260 ( .A1(n3293), .A2(n3294), .ZN(n3309) );
  OR2_X1 U3261 ( .A1(n2138), .A2(n2274), .ZN(n3294) );
  OR2_X1 U3262 ( .A1(n3310), .A2(n3311), .ZN(n3293) );
  AND2_X1 U3263 ( .A1(n3290), .A2(n3289), .ZN(n3311) );
  AND2_X1 U3264 ( .A1(n3287), .A2(n3312), .ZN(n3310) );
  OR2_X1 U3265 ( .A1(n3289), .A2(n3290), .ZN(n3312) );
  OR2_X1 U3266 ( .A1(n2138), .A2(n2278), .ZN(n3290) );
  OR2_X1 U3267 ( .A1(n3313), .A2(n3314), .ZN(n3289) );
  AND2_X1 U3268 ( .A1(n3286), .A2(n3285), .ZN(n3314) );
  AND2_X1 U3269 ( .A1(n3283), .A2(n3315), .ZN(n3313) );
  OR2_X1 U3270 ( .A1(n3285), .A2(n3286), .ZN(n3315) );
  OR2_X1 U3271 ( .A1(n2138), .A2(n2283), .ZN(n3286) );
  OR2_X1 U3272 ( .A1(n3316), .A2(n3317), .ZN(n3285) );
  AND2_X1 U3273 ( .A1(n3279), .A2(n3282), .ZN(n3317) );
  AND2_X1 U3274 ( .A1(n3318), .A2(n3281), .ZN(n3316) );
  OR2_X1 U3275 ( .A1(n3319), .A2(n3320), .ZN(n3281) );
  AND2_X1 U3276 ( .A1(n3278), .A2(n3277), .ZN(n3320) );
  AND2_X1 U3277 ( .A1(n3275), .A2(n3321), .ZN(n3319) );
  OR2_X1 U3278 ( .A1(n3277), .A2(n3278), .ZN(n3321) );
  OR2_X1 U3279 ( .A1(n2138), .A2(n2290), .ZN(n3278) );
  OR2_X1 U3280 ( .A1(n3322), .A2(n3323), .ZN(n3277) );
  AND2_X1 U3281 ( .A1(n3271), .A2(n3274), .ZN(n3323) );
  AND2_X1 U3282 ( .A1(n3324), .A2(n3273), .ZN(n3322) );
  OR2_X1 U3283 ( .A1(n3325), .A2(n3326), .ZN(n3273) );
  AND2_X1 U3284 ( .A1(n3267), .A2(n3270), .ZN(n3326) );
  AND2_X1 U3285 ( .A1(n3327), .A2(n3269), .ZN(n3325) );
  OR2_X1 U3286 ( .A1(n3328), .A2(n3329), .ZN(n3269) );
  AND2_X1 U3287 ( .A1(n3263), .A2(n3266), .ZN(n3329) );
  AND2_X1 U3288 ( .A1(n3330), .A2(n3265), .ZN(n3328) );
  OR2_X1 U3289 ( .A1(n3331), .A2(n3332), .ZN(n3265) );
  AND2_X1 U3290 ( .A1(n3260), .A2(n2135), .ZN(n3332) );
  AND2_X1 U3291 ( .A1(n3333), .A2(n3262), .ZN(n3331) );
  OR2_X1 U3292 ( .A1(n3334), .A2(n3335), .ZN(n3262) );
  AND2_X1 U3293 ( .A1(n3256), .A2(n3259), .ZN(n3335) );
  AND2_X1 U3294 ( .A1(n3336), .A2(n3258), .ZN(n3334) );
  OR2_X1 U3295 ( .A1(n3337), .A2(n3338), .ZN(n3258) );
  AND2_X1 U3296 ( .A1(n3252), .A2(n3255), .ZN(n3338) );
  AND2_X1 U3297 ( .A1(n3339), .A2(n3254), .ZN(n3337) );
  OR2_X1 U3298 ( .A1(n3340), .A2(n3341), .ZN(n3254) );
  AND2_X1 U3299 ( .A1(n3249), .A2(n3251), .ZN(n3341) );
  AND2_X1 U3300 ( .A1(n3342), .A2(n3250), .ZN(n3340) );
  OR2_X1 U3301 ( .A1(n3343), .A2(n3344), .ZN(n3250) );
  AND2_X1 U3302 ( .A1(n3244), .A2(n3247), .ZN(n3344) );
  AND2_X1 U3303 ( .A1(n3246), .A2(n3345), .ZN(n3343) );
  OR2_X1 U3304 ( .A1(n3247), .A2(n3244), .ZN(n3345) );
  OR2_X1 U3305 ( .A1(n2318), .A2(n2138), .ZN(n3244) );
  OR2_X1 U3306 ( .A1(n2755), .A2(n3346), .ZN(n3247) );
  OR2_X1 U3307 ( .A1(n2138), .A2(n2300), .ZN(n3346) );
  INV_X1 U3308 ( .A(n3347), .ZN(n3246) );
  OR2_X1 U3309 ( .A1(n3348), .A2(n3349), .ZN(n3347) );
  AND2_X1 U3310 ( .A1(b_8_), .A2(n3350), .ZN(n3349) );
  OR2_X1 U3311 ( .A1(n3351), .A2(n2043), .ZN(n3350) );
  AND2_X1 U3312 ( .A1(a_14_), .A2(n2168), .ZN(n3351) );
  AND2_X1 U3313 ( .A1(b_7_), .A2(n3352), .ZN(n3348) );
  OR2_X1 U3314 ( .A1(n3353), .A2(n2056), .ZN(n3352) );
  AND2_X1 U3315 ( .A1(a_15_), .A2(n2300), .ZN(n3353) );
  OR2_X1 U3316 ( .A1(n3251), .A2(n3249), .ZN(n3342) );
  XNOR2_X1 U3317 ( .A(n3354), .B(n3355), .ZN(n3249) );
  XNOR2_X1 U3318 ( .A(n3356), .B(n3357), .ZN(n3355) );
  OR2_X1 U3319 ( .A1(n2313), .A2(n2138), .ZN(n3251) );
  OR2_X1 U3320 ( .A1(n3255), .A2(n3252), .ZN(n3339) );
  XNOR2_X1 U3321 ( .A(n3358), .B(n3359), .ZN(n3252) );
  XNOR2_X1 U3322 ( .A(n3360), .B(n3361), .ZN(n3358) );
  OR2_X1 U3323 ( .A1(n2311), .A2(n2138), .ZN(n3255) );
  OR2_X1 U3324 ( .A1(n3259), .A2(n3256), .ZN(n3336) );
  XOR2_X1 U3325 ( .A(n3362), .B(n3363), .Z(n3256) );
  XOR2_X1 U3326 ( .A(n3364), .B(n3365), .Z(n3363) );
  OR2_X1 U3327 ( .A1(n2306), .A2(n2138), .ZN(n3259) );
  OR2_X1 U3328 ( .A1(n2135), .A2(n3260), .ZN(n3333) );
  XOR2_X1 U3329 ( .A(n3366), .B(n3367), .Z(n3260) );
  XOR2_X1 U3330 ( .A(n3368), .B(n3369), .Z(n3367) );
  OR2_X1 U3331 ( .A1(n2138), .A2(n2304), .ZN(n2135) );
  OR2_X1 U3332 ( .A1(n3266), .A2(n3263), .ZN(n3330) );
  XOR2_X1 U3333 ( .A(n3370), .B(n3371), .Z(n3263) );
  XOR2_X1 U3334 ( .A(n3372), .B(n3373), .Z(n3371) );
  OR2_X1 U3335 ( .A1(n2138), .A2(n2299), .ZN(n3266) );
  OR2_X1 U3336 ( .A1(n3270), .A2(n3267), .ZN(n3327) );
  XNOR2_X1 U3337 ( .A(n3374), .B(n3375), .ZN(n3267) );
  XNOR2_X1 U3338 ( .A(n2301), .B(n3376), .ZN(n3374) );
  OR2_X1 U3339 ( .A1(n2138), .A2(n2297), .ZN(n3270) );
  OR2_X1 U3340 ( .A1(n3274), .A2(n3271), .ZN(n3324) );
  XOR2_X1 U3341 ( .A(n3377), .B(n3378), .Z(n3271) );
  XOR2_X1 U3342 ( .A(n3379), .B(n3380), .Z(n3378) );
  OR2_X1 U3343 ( .A1(n2138), .A2(n2292), .ZN(n3274) );
  XOR2_X1 U3344 ( .A(n3381), .B(n3382), .Z(n3275) );
  XOR2_X1 U3345 ( .A(n3383), .B(n3384), .Z(n3382) );
  OR2_X1 U3346 ( .A1(n3282), .A2(n3279), .ZN(n3318) );
  XOR2_X1 U3347 ( .A(n3385), .B(n3386), .Z(n3279) );
  XOR2_X1 U3348 ( .A(n3387), .B(n3388), .Z(n3386) );
  OR2_X1 U3349 ( .A1(n2138), .A2(n2285), .ZN(n3282) );
  INV_X1 U3350 ( .A(b_9_), .ZN(n2138) );
  XOR2_X1 U3351 ( .A(n3389), .B(n3390), .Z(n3283) );
  XOR2_X1 U3352 ( .A(n3391), .B(n3392), .Z(n3390) );
  XOR2_X1 U3353 ( .A(n3393), .B(n3394), .Z(n3287) );
  XOR2_X1 U3354 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR2_X1 U3355 ( .A(n3397), .B(n3398), .Z(n3291) );
  XOR2_X1 U3356 ( .A(n3399), .B(n3400), .Z(n3398) );
  XOR2_X1 U3357 ( .A(n3401), .B(n3402), .Z(n3295) );
  XOR2_X1 U3358 ( .A(n3403), .B(n3404), .Z(n3402) );
  XOR2_X1 U3359 ( .A(n2595), .B(n3405), .Z(n3302) );
  XOR2_X1 U3360 ( .A(n2594), .B(n2593), .Z(n3405) );
  OR2_X1 U3361 ( .A1(n2300), .A2(n2427), .ZN(n2593) );
  OR2_X1 U3362 ( .A1(n3406), .A2(n3407), .ZN(n2594) );
  AND2_X1 U3363 ( .A1(n3404), .A2(n3403), .ZN(n3407) );
  AND2_X1 U3364 ( .A1(n3401), .A2(n3408), .ZN(n3406) );
  OR2_X1 U3365 ( .A1(n3403), .A2(n3404), .ZN(n3408) );
  OR2_X1 U3366 ( .A1(n2300), .A2(n2274), .ZN(n3404) );
  OR2_X1 U3367 ( .A1(n3409), .A2(n3410), .ZN(n3403) );
  AND2_X1 U3368 ( .A1(n3400), .A2(n3399), .ZN(n3410) );
  AND2_X1 U3369 ( .A1(n3397), .A2(n3411), .ZN(n3409) );
  OR2_X1 U3370 ( .A1(n3399), .A2(n3400), .ZN(n3411) );
  OR2_X1 U3371 ( .A1(n2300), .A2(n2278), .ZN(n3400) );
  OR2_X1 U3372 ( .A1(n3412), .A2(n3413), .ZN(n3399) );
  AND2_X1 U3373 ( .A1(n3396), .A2(n3395), .ZN(n3413) );
  AND2_X1 U3374 ( .A1(n3393), .A2(n3414), .ZN(n3412) );
  OR2_X1 U3375 ( .A1(n3395), .A2(n3396), .ZN(n3414) );
  OR2_X1 U3376 ( .A1(n2300), .A2(n2283), .ZN(n3396) );
  OR2_X1 U3377 ( .A1(n3415), .A2(n3416), .ZN(n3395) );
  AND2_X1 U3378 ( .A1(n3392), .A2(n3391), .ZN(n3416) );
  AND2_X1 U3379 ( .A1(n3389), .A2(n3417), .ZN(n3415) );
  OR2_X1 U3380 ( .A1(n3391), .A2(n3392), .ZN(n3417) );
  OR2_X1 U3381 ( .A1(n2300), .A2(n2285), .ZN(n3392) );
  OR2_X1 U3382 ( .A1(n3418), .A2(n3419), .ZN(n3391) );
  AND2_X1 U3383 ( .A1(n3385), .A2(n3388), .ZN(n3419) );
  AND2_X1 U3384 ( .A1(n3420), .A2(n3387), .ZN(n3418) );
  OR2_X1 U3385 ( .A1(n3421), .A2(n3422), .ZN(n3387) );
  AND2_X1 U3386 ( .A1(n3384), .A2(n3383), .ZN(n3422) );
  AND2_X1 U3387 ( .A1(n3381), .A2(n3423), .ZN(n3421) );
  OR2_X1 U3388 ( .A1(n3383), .A2(n3384), .ZN(n3423) );
  OR2_X1 U3389 ( .A1(n2300), .A2(n2292), .ZN(n3384) );
  OR2_X1 U3390 ( .A1(n3424), .A2(n3425), .ZN(n3383) );
  AND2_X1 U3391 ( .A1(n3377), .A2(n3380), .ZN(n3425) );
  AND2_X1 U3392 ( .A1(n3426), .A2(n3379), .ZN(n3424) );
  OR2_X1 U3393 ( .A1(n3427), .A2(n3428), .ZN(n3379) );
  AND2_X1 U3394 ( .A1(n3375), .A2(n2301), .ZN(n3428) );
  AND2_X1 U3395 ( .A1(n3429), .A2(n3376), .ZN(n3427) );
  OR2_X1 U3396 ( .A1(n3430), .A2(n3431), .ZN(n3376) );
  AND2_X1 U3397 ( .A1(n3370), .A2(n3373), .ZN(n3431) );
  AND2_X1 U3398 ( .A1(n3432), .A2(n3372), .ZN(n3430) );
  OR2_X1 U3399 ( .A1(n3433), .A2(n3434), .ZN(n3372) );
  AND2_X1 U3400 ( .A1(n3366), .A2(n3369), .ZN(n3434) );
  AND2_X1 U3401 ( .A1(n3435), .A2(n3368), .ZN(n3433) );
  OR2_X1 U3402 ( .A1(n3436), .A2(n3437), .ZN(n3368) );
  AND2_X1 U3403 ( .A1(n3362), .A2(n3365), .ZN(n3437) );
  AND2_X1 U3404 ( .A1(n3438), .A2(n3364), .ZN(n3436) );
  OR2_X1 U3405 ( .A1(n3439), .A2(n3440), .ZN(n3364) );
  AND2_X1 U3406 ( .A1(n3359), .A2(n3361), .ZN(n3440) );
  AND2_X1 U3407 ( .A1(n3441), .A2(n3360), .ZN(n3439) );
  OR2_X1 U3408 ( .A1(n3442), .A2(n3443), .ZN(n3360) );
  AND2_X1 U3409 ( .A1(n3354), .A2(n3357), .ZN(n3443) );
  AND2_X1 U3410 ( .A1(n3356), .A2(n3444), .ZN(n3442) );
  OR2_X1 U3411 ( .A1(n3357), .A2(n3354), .ZN(n3444) );
  OR2_X1 U3412 ( .A1(n2318), .A2(n2300), .ZN(n3354) );
  OR2_X1 U3413 ( .A1(n2755), .A2(n3445), .ZN(n3357) );
  OR2_X1 U3414 ( .A1(n2300), .A2(n2168), .ZN(n3445) );
  INV_X1 U3415 ( .A(n3446), .ZN(n3356) );
  OR2_X1 U3416 ( .A1(n3447), .A2(n3448), .ZN(n3446) );
  AND2_X1 U3417 ( .A1(b_7_), .A2(n3449), .ZN(n3448) );
  OR2_X1 U3418 ( .A1(n3450), .A2(n2043), .ZN(n3449) );
  AND2_X1 U3419 ( .A1(a_14_), .A2(n2293), .ZN(n3450) );
  AND2_X1 U3420 ( .A1(b_6_), .A2(n3451), .ZN(n3447) );
  OR2_X1 U3421 ( .A1(n3452), .A2(n2056), .ZN(n3451) );
  AND2_X1 U3422 ( .A1(a_15_), .A2(n2168), .ZN(n3452) );
  OR2_X1 U3423 ( .A1(n3361), .A2(n3359), .ZN(n3441) );
  XNOR2_X1 U3424 ( .A(n3453), .B(n3454), .ZN(n3359) );
  XNOR2_X1 U3425 ( .A(n3455), .B(n3456), .ZN(n3454) );
  OR2_X1 U3426 ( .A1(n2313), .A2(n2300), .ZN(n3361) );
  OR2_X1 U3427 ( .A1(n3365), .A2(n3362), .ZN(n3438) );
  XNOR2_X1 U3428 ( .A(n3457), .B(n3458), .ZN(n3362) );
  XNOR2_X1 U3429 ( .A(n3459), .B(n3460), .ZN(n3457) );
  OR2_X1 U3430 ( .A1(n2311), .A2(n2300), .ZN(n3365) );
  OR2_X1 U3431 ( .A1(n3369), .A2(n3366), .ZN(n3435) );
  XOR2_X1 U3432 ( .A(n3461), .B(n3462), .Z(n3366) );
  XOR2_X1 U3433 ( .A(n3463), .B(n3464), .Z(n3462) );
  OR2_X1 U3434 ( .A1(n2306), .A2(n2300), .ZN(n3369) );
  OR2_X1 U3435 ( .A1(n3373), .A2(n3370), .ZN(n3432) );
  XOR2_X1 U3436 ( .A(n3465), .B(n3466), .Z(n3370) );
  XOR2_X1 U3437 ( .A(n3467), .B(n3468), .Z(n3466) );
  OR2_X1 U3438 ( .A1(n2304), .A2(n2300), .ZN(n3373) );
  OR2_X1 U3439 ( .A1(n2301), .A2(n3375), .ZN(n3429) );
  XOR2_X1 U3440 ( .A(n3469), .B(n3470), .Z(n3375) );
  XOR2_X1 U3441 ( .A(n3471), .B(n3472), .Z(n3470) );
  INV_X1 U3442 ( .A(n2150), .ZN(n2301) );
  AND2_X1 U3443 ( .A1(a_8_), .A2(b_8_), .ZN(n2150) );
  OR2_X1 U3444 ( .A1(n3380), .A2(n3377), .ZN(n3426) );
  XOR2_X1 U3445 ( .A(n3473), .B(n3474), .Z(n3377) );
  XOR2_X1 U3446 ( .A(n3475), .B(n3476), .Z(n3474) );
  OR2_X1 U3447 ( .A1(n2300), .A2(n2297), .ZN(n3380) );
  XOR2_X1 U3448 ( .A(n3477), .B(n3478), .Z(n3381) );
  XOR2_X1 U3449 ( .A(n3479), .B(n2165), .Z(n3478) );
  OR2_X1 U3450 ( .A1(n3388), .A2(n3385), .ZN(n3420) );
  XOR2_X1 U3451 ( .A(n3480), .B(n3481), .Z(n3385) );
  XOR2_X1 U3452 ( .A(n3482), .B(n3483), .Z(n3481) );
  OR2_X1 U3453 ( .A1(n2300), .A2(n2290), .ZN(n3388) );
  INV_X1 U3454 ( .A(b_8_), .ZN(n2300) );
  XOR2_X1 U3455 ( .A(n3484), .B(n3485), .Z(n3389) );
  XOR2_X1 U3456 ( .A(n3486), .B(n3487), .Z(n3485) );
  XOR2_X1 U3457 ( .A(n3488), .B(n3489), .Z(n3393) );
  XOR2_X1 U3458 ( .A(n3490), .B(n3491), .Z(n3489) );
  XOR2_X1 U3459 ( .A(n3492), .B(n3493), .Z(n3397) );
  XOR2_X1 U3460 ( .A(n3494), .B(n3495), .Z(n3493) );
  XOR2_X1 U3461 ( .A(n3496), .B(n3497), .Z(n3401) );
  XOR2_X1 U3462 ( .A(n3498), .B(n3499), .Z(n3497) );
  XOR2_X1 U3463 ( .A(n2602), .B(n3500), .Z(n2595) );
  XOR2_X1 U3464 ( .A(n2601), .B(n2600), .Z(n3500) );
  OR2_X1 U3465 ( .A1(n2168), .A2(n2274), .ZN(n2600) );
  OR2_X1 U3466 ( .A1(n3501), .A2(n3502), .ZN(n2601) );
  AND2_X1 U3467 ( .A1(n3499), .A2(n3498), .ZN(n3502) );
  AND2_X1 U3468 ( .A1(n3496), .A2(n3503), .ZN(n3501) );
  OR2_X1 U3469 ( .A1(n3498), .A2(n3499), .ZN(n3503) );
  OR2_X1 U3470 ( .A1(n2168), .A2(n2278), .ZN(n3499) );
  OR2_X1 U3471 ( .A1(n3504), .A2(n3505), .ZN(n3498) );
  AND2_X1 U3472 ( .A1(n3495), .A2(n3494), .ZN(n3505) );
  AND2_X1 U3473 ( .A1(n3492), .A2(n3506), .ZN(n3504) );
  OR2_X1 U3474 ( .A1(n3494), .A2(n3495), .ZN(n3506) );
  OR2_X1 U3475 ( .A1(n2168), .A2(n2283), .ZN(n3495) );
  OR2_X1 U3476 ( .A1(n3507), .A2(n3508), .ZN(n3494) );
  AND2_X1 U3477 ( .A1(n3491), .A2(n3490), .ZN(n3508) );
  AND2_X1 U3478 ( .A1(n3488), .A2(n3509), .ZN(n3507) );
  OR2_X1 U3479 ( .A1(n3490), .A2(n3491), .ZN(n3509) );
  OR2_X1 U3480 ( .A1(n2168), .A2(n2285), .ZN(n3491) );
  OR2_X1 U3481 ( .A1(n3510), .A2(n3511), .ZN(n3490) );
  AND2_X1 U3482 ( .A1(n3487), .A2(n3486), .ZN(n3511) );
  AND2_X1 U3483 ( .A1(n3484), .A2(n3512), .ZN(n3510) );
  OR2_X1 U3484 ( .A1(n3486), .A2(n3487), .ZN(n3512) );
  OR2_X1 U3485 ( .A1(n2168), .A2(n2290), .ZN(n3487) );
  OR2_X1 U3486 ( .A1(n3513), .A2(n3514), .ZN(n3486) );
  AND2_X1 U3487 ( .A1(n3480), .A2(n3483), .ZN(n3514) );
  AND2_X1 U3488 ( .A1(n3515), .A2(n3482), .ZN(n3513) );
  OR2_X1 U3489 ( .A1(n3516), .A2(n3517), .ZN(n3482) );
  AND2_X1 U3490 ( .A1(n2165), .A2(n3479), .ZN(n3517) );
  AND2_X1 U3491 ( .A1(n3477), .A2(n3518), .ZN(n3516) );
  OR2_X1 U3492 ( .A1(n3479), .A2(n2165), .ZN(n3518) );
  OR2_X1 U3493 ( .A1(n2168), .A2(n2297), .ZN(n2165) );
  OR2_X1 U3494 ( .A1(n3519), .A2(n3520), .ZN(n3479) );
  AND2_X1 U3495 ( .A1(n3473), .A2(n3476), .ZN(n3520) );
  AND2_X1 U3496 ( .A1(n3521), .A2(n3475), .ZN(n3519) );
  OR2_X1 U3497 ( .A1(n3522), .A2(n3523), .ZN(n3475) );
  AND2_X1 U3498 ( .A1(n3469), .A2(n3472), .ZN(n3523) );
  AND2_X1 U3499 ( .A1(n3524), .A2(n3471), .ZN(n3522) );
  OR2_X1 U3500 ( .A1(n3525), .A2(n3526), .ZN(n3471) );
  AND2_X1 U3501 ( .A1(n3465), .A2(n3468), .ZN(n3526) );
  AND2_X1 U3502 ( .A1(n3527), .A2(n3467), .ZN(n3525) );
  OR2_X1 U3503 ( .A1(n3528), .A2(n3529), .ZN(n3467) );
  AND2_X1 U3504 ( .A1(n3461), .A2(n3464), .ZN(n3529) );
  AND2_X1 U3505 ( .A1(n3530), .A2(n3463), .ZN(n3528) );
  OR2_X1 U3506 ( .A1(n3531), .A2(n3532), .ZN(n3463) );
  AND2_X1 U3507 ( .A1(n3458), .A2(n3460), .ZN(n3532) );
  AND2_X1 U3508 ( .A1(n3533), .A2(n3459), .ZN(n3531) );
  OR2_X1 U3509 ( .A1(n3534), .A2(n3535), .ZN(n3459) );
  AND2_X1 U3510 ( .A1(n3453), .A2(n3456), .ZN(n3535) );
  AND2_X1 U3511 ( .A1(n3455), .A2(n3536), .ZN(n3534) );
  OR2_X1 U3512 ( .A1(n3456), .A2(n3453), .ZN(n3536) );
  OR2_X1 U3513 ( .A1(n2318), .A2(n2168), .ZN(n3453) );
  OR2_X1 U3514 ( .A1(n2755), .A2(n3537), .ZN(n3456) );
  OR2_X1 U3515 ( .A1(n2168), .A2(n2293), .ZN(n3537) );
  INV_X1 U3516 ( .A(n3538), .ZN(n3455) );
  OR2_X1 U3517 ( .A1(n3539), .A2(n3540), .ZN(n3538) );
  AND2_X1 U3518 ( .A1(b_6_), .A2(n3541), .ZN(n3540) );
  OR2_X1 U3519 ( .A1(n3542), .A2(n2043), .ZN(n3541) );
  AND2_X1 U3520 ( .A1(a_14_), .A2(n2198), .ZN(n3542) );
  AND2_X1 U3521 ( .A1(b_5_), .A2(n3543), .ZN(n3539) );
  OR2_X1 U3522 ( .A1(n3544), .A2(n2056), .ZN(n3543) );
  AND2_X1 U3523 ( .A1(a_15_), .A2(n2293), .ZN(n3544) );
  OR2_X1 U3524 ( .A1(n3460), .A2(n3458), .ZN(n3533) );
  XNOR2_X1 U3525 ( .A(n3545), .B(n3546), .ZN(n3458) );
  XNOR2_X1 U3526 ( .A(n3547), .B(n3548), .ZN(n3546) );
  OR2_X1 U3527 ( .A1(n2313), .A2(n2168), .ZN(n3460) );
  OR2_X1 U3528 ( .A1(n3464), .A2(n3461), .ZN(n3530) );
  XNOR2_X1 U3529 ( .A(n3549), .B(n3550), .ZN(n3461) );
  XNOR2_X1 U3530 ( .A(n3551), .B(n3552), .ZN(n3549) );
  OR2_X1 U3531 ( .A1(n2311), .A2(n2168), .ZN(n3464) );
  OR2_X1 U3532 ( .A1(n3468), .A2(n3465), .ZN(n3527) );
  XOR2_X1 U3533 ( .A(n3553), .B(n3554), .Z(n3465) );
  XOR2_X1 U3534 ( .A(n3555), .B(n3556), .Z(n3554) );
  OR2_X1 U3535 ( .A1(n2306), .A2(n2168), .ZN(n3468) );
  OR2_X1 U3536 ( .A1(n3472), .A2(n3469), .ZN(n3524) );
  XOR2_X1 U3537 ( .A(n3557), .B(n3558), .Z(n3469) );
  XOR2_X1 U3538 ( .A(n3559), .B(n3560), .Z(n3558) );
  OR2_X1 U3539 ( .A1(n2304), .A2(n2168), .ZN(n3472) );
  OR2_X1 U3540 ( .A1(n3476), .A2(n3473), .ZN(n3521) );
  XOR2_X1 U3541 ( .A(n3561), .B(n3562), .Z(n3473) );
  XOR2_X1 U3542 ( .A(n3563), .B(n3564), .Z(n3562) );
  OR2_X1 U3543 ( .A1(n2299), .A2(n2168), .ZN(n3476) );
  XOR2_X1 U3544 ( .A(n3565), .B(n3566), .Z(n3477) );
  XOR2_X1 U3545 ( .A(n3567), .B(n3568), .Z(n3566) );
  OR2_X1 U3546 ( .A1(n3483), .A2(n3480), .ZN(n3515) );
  XOR2_X1 U3547 ( .A(n3569), .B(n3570), .Z(n3480) );
  XOR2_X1 U3548 ( .A(n3571), .B(n3572), .Z(n3570) );
  OR2_X1 U3549 ( .A1(n2168), .A2(n2292), .ZN(n3483) );
  INV_X1 U3550 ( .A(b_7_), .ZN(n2168) );
  XNOR2_X1 U3551 ( .A(n3573), .B(n3574), .ZN(n3484) );
  XNOR2_X1 U3552 ( .A(n2294), .B(n3575), .ZN(n3573) );
  XOR2_X1 U3553 ( .A(n3576), .B(n3577), .Z(n3488) );
  XOR2_X1 U3554 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR2_X1 U3555 ( .A(n3580), .B(n3581), .Z(n3492) );
  XOR2_X1 U3556 ( .A(n3582), .B(n3583), .Z(n3581) );
  XOR2_X1 U3557 ( .A(n3584), .B(n3585), .Z(n3496) );
  XOR2_X1 U3558 ( .A(n3586), .B(n3587), .Z(n3585) );
  XOR2_X1 U3559 ( .A(n2609), .B(n3588), .Z(n2602) );
  XOR2_X1 U3560 ( .A(n2608), .B(n2607), .Z(n3588) );
  OR2_X1 U3561 ( .A1(n2293), .A2(n2278), .ZN(n2607) );
  OR2_X1 U3562 ( .A1(n3589), .A2(n3590), .ZN(n2608) );
  AND2_X1 U3563 ( .A1(n3587), .A2(n3586), .ZN(n3590) );
  AND2_X1 U3564 ( .A1(n3584), .A2(n3591), .ZN(n3589) );
  OR2_X1 U3565 ( .A1(n3586), .A2(n3587), .ZN(n3591) );
  OR2_X1 U3566 ( .A1(n2293), .A2(n2283), .ZN(n3587) );
  OR2_X1 U3567 ( .A1(n3592), .A2(n3593), .ZN(n3586) );
  AND2_X1 U3568 ( .A1(n3583), .A2(n3582), .ZN(n3593) );
  AND2_X1 U3569 ( .A1(n3580), .A2(n3594), .ZN(n3592) );
  OR2_X1 U3570 ( .A1(n3582), .A2(n3583), .ZN(n3594) );
  OR2_X1 U3571 ( .A1(n2293), .A2(n2285), .ZN(n3583) );
  OR2_X1 U3572 ( .A1(n3595), .A2(n3596), .ZN(n3582) );
  AND2_X1 U3573 ( .A1(n3579), .A2(n3578), .ZN(n3596) );
  AND2_X1 U3574 ( .A1(n3576), .A2(n3597), .ZN(n3595) );
  OR2_X1 U3575 ( .A1(n3578), .A2(n3579), .ZN(n3597) );
  OR2_X1 U3576 ( .A1(n2293), .A2(n2290), .ZN(n3579) );
  OR2_X1 U3577 ( .A1(n3598), .A2(n3599), .ZN(n3578) );
  AND2_X1 U3578 ( .A1(n3575), .A2(n2294), .ZN(n3599) );
  AND2_X1 U3579 ( .A1(n3574), .A2(n3600), .ZN(n3598) );
  OR2_X1 U3580 ( .A1(n2294), .A2(n3575), .ZN(n3600) );
  OR2_X1 U3581 ( .A1(n3601), .A2(n3602), .ZN(n3575) );
  AND2_X1 U3582 ( .A1(n3569), .A2(n3572), .ZN(n3602) );
  AND2_X1 U3583 ( .A1(n3603), .A2(n3571), .ZN(n3601) );
  OR2_X1 U3584 ( .A1(n3604), .A2(n3605), .ZN(n3571) );
  AND2_X1 U3585 ( .A1(n3568), .A2(n3567), .ZN(n3605) );
  AND2_X1 U3586 ( .A1(n3565), .A2(n3606), .ZN(n3604) );
  OR2_X1 U3587 ( .A1(n3567), .A2(n3568), .ZN(n3606) );
  OR2_X1 U3588 ( .A1(n2299), .A2(n2293), .ZN(n3568) );
  OR2_X1 U3589 ( .A1(n3607), .A2(n3608), .ZN(n3567) );
  AND2_X1 U3590 ( .A1(n3561), .A2(n3564), .ZN(n3608) );
  AND2_X1 U3591 ( .A1(n3609), .A2(n3563), .ZN(n3607) );
  OR2_X1 U3592 ( .A1(n3610), .A2(n3611), .ZN(n3563) );
  AND2_X1 U3593 ( .A1(n3557), .A2(n3560), .ZN(n3611) );
  AND2_X1 U3594 ( .A1(n3612), .A2(n3559), .ZN(n3610) );
  OR2_X1 U3595 ( .A1(n3613), .A2(n3614), .ZN(n3559) );
  AND2_X1 U3596 ( .A1(n3553), .A2(n3556), .ZN(n3614) );
  AND2_X1 U3597 ( .A1(n3615), .A2(n3555), .ZN(n3613) );
  OR2_X1 U3598 ( .A1(n3616), .A2(n3617), .ZN(n3555) );
  AND2_X1 U3599 ( .A1(n3550), .A2(n3552), .ZN(n3617) );
  AND2_X1 U3600 ( .A1(n3618), .A2(n3551), .ZN(n3616) );
  OR2_X1 U3601 ( .A1(n3619), .A2(n3620), .ZN(n3551) );
  AND2_X1 U3602 ( .A1(n3545), .A2(n3548), .ZN(n3620) );
  AND2_X1 U3603 ( .A1(n3547), .A2(n3621), .ZN(n3619) );
  OR2_X1 U3604 ( .A1(n3548), .A2(n3545), .ZN(n3621) );
  OR2_X1 U3605 ( .A1(n2318), .A2(n2293), .ZN(n3545) );
  OR2_X1 U3606 ( .A1(n2755), .A2(n3622), .ZN(n3548) );
  OR2_X1 U3607 ( .A1(n2293), .A2(n2198), .ZN(n3622) );
  INV_X1 U3608 ( .A(n3623), .ZN(n3547) );
  OR2_X1 U3609 ( .A1(n3624), .A2(n3625), .ZN(n3623) );
  AND2_X1 U3610 ( .A1(b_5_), .A2(n3626), .ZN(n3625) );
  OR2_X1 U3611 ( .A1(n3627), .A2(n2043), .ZN(n3626) );
  AND2_X1 U3612 ( .A1(a_14_), .A2(n2286), .ZN(n3627) );
  AND2_X1 U3613 ( .A1(b_4_), .A2(n3628), .ZN(n3624) );
  OR2_X1 U3614 ( .A1(n3629), .A2(n2056), .ZN(n3628) );
  AND2_X1 U3615 ( .A1(a_15_), .A2(n2198), .ZN(n3629) );
  OR2_X1 U3616 ( .A1(n3552), .A2(n3550), .ZN(n3618) );
  XNOR2_X1 U3617 ( .A(n3630), .B(n3631), .ZN(n3550) );
  XNOR2_X1 U3618 ( .A(n3632), .B(n3633), .ZN(n3631) );
  OR2_X1 U3619 ( .A1(n2313), .A2(n2293), .ZN(n3552) );
  OR2_X1 U3620 ( .A1(n3556), .A2(n3553), .ZN(n3615) );
  XNOR2_X1 U3621 ( .A(n3634), .B(n3635), .ZN(n3553) );
  XNOR2_X1 U3622 ( .A(n3636), .B(n3637), .ZN(n3634) );
  OR2_X1 U3623 ( .A1(n2311), .A2(n2293), .ZN(n3556) );
  OR2_X1 U3624 ( .A1(n3560), .A2(n3557), .ZN(n3612) );
  XOR2_X1 U3625 ( .A(n3638), .B(n3639), .Z(n3557) );
  XOR2_X1 U3626 ( .A(n3640), .B(n3641), .Z(n3639) );
  OR2_X1 U3627 ( .A1(n2306), .A2(n2293), .ZN(n3560) );
  OR2_X1 U3628 ( .A1(n3564), .A2(n3561), .ZN(n3609) );
  XOR2_X1 U3629 ( .A(n3642), .B(n3643), .Z(n3561) );
  XOR2_X1 U3630 ( .A(n3644), .B(n3645), .Z(n3643) );
  OR2_X1 U3631 ( .A1(n2304), .A2(n2293), .ZN(n3564) );
  XOR2_X1 U3632 ( .A(n3646), .B(n3647), .Z(n3565) );
  XOR2_X1 U3633 ( .A(n3648), .B(n3649), .Z(n3647) );
  OR2_X1 U3634 ( .A1(n3572), .A2(n3569), .ZN(n3603) );
  XOR2_X1 U3635 ( .A(n3650), .B(n3651), .Z(n3569) );
  XOR2_X1 U3636 ( .A(n3652), .B(n3653), .Z(n3651) );
  OR2_X1 U3637 ( .A1(n2297), .A2(n2293), .ZN(n3572) );
  INV_X1 U3638 ( .A(b_6_), .ZN(n2293) );
  INV_X1 U3639 ( .A(n2180), .ZN(n2294) );
  AND2_X1 U3640 ( .A1(a_6_), .A2(b_6_), .ZN(n2180) );
  XOR2_X1 U3641 ( .A(n3654), .B(n3655), .Z(n3574) );
  XOR2_X1 U3642 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR2_X1 U3643 ( .A(n3658), .B(n3659), .Z(n3576) );
  XOR2_X1 U3644 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR2_X1 U3645 ( .A(n3662), .B(n3663), .Z(n3580) );
  XOR2_X1 U3646 ( .A(n3664), .B(n2195), .Z(n3663) );
  XOR2_X1 U3647 ( .A(n3665), .B(n3666), .Z(n3584) );
  XOR2_X1 U3648 ( .A(n3667), .B(n3668), .Z(n3666) );
  XOR2_X1 U3649 ( .A(n2616), .B(n3669), .Z(n2609) );
  XOR2_X1 U3650 ( .A(n2615), .B(n2614), .Z(n3669) );
  OR2_X1 U3651 ( .A1(n2198), .A2(n2283), .ZN(n2614) );
  OR2_X1 U3652 ( .A1(n3670), .A2(n3671), .ZN(n2615) );
  AND2_X1 U3653 ( .A1(n3668), .A2(n3667), .ZN(n3671) );
  AND2_X1 U3654 ( .A1(n3665), .A2(n3672), .ZN(n3670) );
  OR2_X1 U3655 ( .A1(n3667), .A2(n3668), .ZN(n3672) );
  OR2_X1 U3656 ( .A1(n2198), .A2(n2285), .ZN(n3668) );
  OR2_X1 U3657 ( .A1(n3673), .A2(n3674), .ZN(n3667) );
  AND2_X1 U3658 ( .A1(n2195), .A2(n3664), .ZN(n3674) );
  AND2_X1 U3659 ( .A1(n3662), .A2(n3675), .ZN(n3673) );
  OR2_X1 U3660 ( .A1(n3664), .A2(n2195), .ZN(n3675) );
  OR2_X1 U3661 ( .A1(n2198), .A2(n2290), .ZN(n2195) );
  OR2_X1 U3662 ( .A1(n3676), .A2(n3677), .ZN(n3664) );
  AND2_X1 U3663 ( .A1(n3661), .A2(n3660), .ZN(n3677) );
  AND2_X1 U3664 ( .A1(n3658), .A2(n3678), .ZN(n3676) );
  OR2_X1 U3665 ( .A1(n3660), .A2(n3661), .ZN(n3678) );
  OR2_X1 U3666 ( .A1(n2292), .A2(n2198), .ZN(n3661) );
  OR2_X1 U3667 ( .A1(n3679), .A2(n3680), .ZN(n3660) );
  AND2_X1 U3668 ( .A1(n3657), .A2(n3656), .ZN(n3680) );
  AND2_X1 U3669 ( .A1(n3654), .A2(n3681), .ZN(n3679) );
  OR2_X1 U3670 ( .A1(n3656), .A2(n3657), .ZN(n3681) );
  OR2_X1 U3671 ( .A1(n2297), .A2(n2198), .ZN(n3657) );
  OR2_X1 U3672 ( .A1(n3682), .A2(n3683), .ZN(n3656) );
  AND2_X1 U3673 ( .A1(n3650), .A2(n3653), .ZN(n3683) );
  AND2_X1 U3674 ( .A1(n3684), .A2(n3652), .ZN(n3682) );
  OR2_X1 U3675 ( .A1(n3685), .A2(n3686), .ZN(n3652) );
  AND2_X1 U3676 ( .A1(n3649), .A2(n3648), .ZN(n3686) );
  AND2_X1 U3677 ( .A1(n3646), .A2(n3687), .ZN(n3685) );
  OR2_X1 U3678 ( .A1(n3648), .A2(n3649), .ZN(n3687) );
  OR2_X1 U3679 ( .A1(n2304), .A2(n2198), .ZN(n3649) );
  OR2_X1 U3680 ( .A1(n3688), .A2(n3689), .ZN(n3648) );
  AND2_X1 U3681 ( .A1(n3642), .A2(n3645), .ZN(n3689) );
  AND2_X1 U3682 ( .A1(n3690), .A2(n3644), .ZN(n3688) );
  OR2_X1 U3683 ( .A1(n3691), .A2(n3692), .ZN(n3644) );
  AND2_X1 U3684 ( .A1(n3638), .A2(n3641), .ZN(n3692) );
  AND2_X1 U3685 ( .A1(n3693), .A2(n3640), .ZN(n3691) );
  OR2_X1 U3686 ( .A1(n3694), .A2(n3695), .ZN(n3640) );
  AND2_X1 U3687 ( .A1(n3635), .A2(n3637), .ZN(n3695) );
  AND2_X1 U3688 ( .A1(n3696), .A2(n3636), .ZN(n3694) );
  OR2_X1 U3689 ( .A1(n3697), .A2(n3698), .ZN(n3636) );
  AND2_X1 U3690 ( .A1(n3630), .A2(n3633), .ZN(n3698) );
  AND2_X1 U3691 ( .A1(n3632), .A2(n3699), .ZN(n3697) );
  OR2_X1 U3692 ( .A1(n3633), .A2(n3630), .ZN(n3699) );
  OR2_X1 U3693 ( .A1(n2318), .A2(n2198), .ZN(n3630) );
  OR2_X1 U3694 ( .A1(n2755), .A2(n3700), .ZN(n3633) );
  OR2_X1 U3695 ( .A1(n2198), .A2(n2286), .ZN(n3700) );
  INV_X1 U3696 ( .A(n3701), .ZN(n3632) );
  OR2_X1 U3697 ( .A1(n3702), .A2(n3703), .ZN(n3701) );
  AND2_X1 U3698 ( .A1(b_4_), .A2(n3704), .ZN(n3703) );
  OR2_X1 U3699 ( .A1(n3705), .A2(n2043), .ZN(n3704) );
  AND2_X1 U3700 ( .A1(a_14_), .A2(n2235), .ZN(n3705) );
  AND2_X1 U3701 ( .A1(b_3_), .A2(n3706), .ZN(n3702) );
  OR2_X1 U3702 ( .A1(n3707), .A2(n2056), .ZN(n3706) );
  AND2_X1 U3703 ( .A1(a_15_), .A2(n2286), .ZN(n3707) );
  OR2_X1 U3704 ( .A1(n3637), .A2(n3635), .ZN(n3696) );
  XNOR2_X1 U3705 ( .A(n3708), .B(n3709), .ZN(n3635) );
  XNOR2_X1 U3706 ( .A(n3710), .B(n3711), .ZN(n3709) );
  OR2_X1 U3707 ( .A1(n2313), .A2(n2198), .ZN(n3637) );
  OR2_X1 U3708 ( .A1(n3641), .A2(n3638), .ZN(n3693) );
  XNOR2_X1 U3709 ( .A(n3712), .B(n3713), .ZN(n3638) );
  XNOR2_X1 U3710 ( .A(n3714), .B(n3715), .ZN(n3712) );
  OR2_X1 U3711 ( .A1(n2311), .A2(n2198), .ZN(n3641) );
  OR2_X1 U3712 ( .A1(n3645), .A2(n3642), .ZN(n3690) );
  XOR2_X1 U3713 ( .A(n3716), .B(n3717), .Z(n3642) );
  XOR2_X1 U3714 ( .A(n3718), .B(n3719), .Z(n3717) );
  OR2_X1 U3715 ( .A1(n2306), .A2(n2198), .ZN(n3645) );
  XOR2_X1 U3716 ( .A(n3720), .B(n3721), .Z(n3646) );
  XOR2_X1 U3717 ( .A(n3722), .B(n3723), .Z(n3721) );
  OR2_X1 U3718 ( .A1(n3653), .A2(n3650), .ZN(n3684) );
  XOR2_X1 U3719 ( .A(n3724), .B(n3725), .Z(n3650) );
  XOR2_X1 U3720 ( .A(n3726), .B(n3727), .Z(n3725) );
  OR2_X1 U3721 ( .A1(n2299), .A2(n2198), .ZN(n3653) );
  INV_X1 U3722 ( .A(b_5_), .ZN(n2198) );
  XOR2_X1 U3723 ( .A(n3728), .B(n3729), .Z(n3654) );
  XOR2_X1 U3724 ( .A(n3730), .B(n3731), .Z(n3729) );
  XOR2_X1 U3725 ( .A(n3732), .B(n3733), .Z(n3658) );
  XOR2_X1 U3726 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR2_X1 U3727 ( .A(n3736), .B(n3737), .Z(n3662) );
  XOR2_X1 U3728 ( .A(n3738), .B(n3739), .Z(n3737) );
  XOR2_X1 U3729 ( .A(n3740), .B(n3741), .Z(n3665) );
  XOR2_X1 U3730 ( .A(n3742), .B(n3743), .Z(n3741) );
  XNOR2_X1 U3731 ( .A(n3744), .B(n2622), .ZN(n2616) );
  XOR2_X1 U3732 ( .A(n2629), .B(n3745), .Z(n2622) );
  XOR2_X1 U3733 ( .A(n2628), .B(n2627), .Z(n3745) );
  OR2_X1 U3734 ( .A1(n2290), .A2(n2235), .ZN(n2627) );
  OR2_X1 U3735 ( .A1(n3746), .A2(n3747), .ZN(n2628) );
  AND2_X1 U3736 ( .A1(n3748), .A2(n3749), .ZN(n3747) );
  AND2_X1 U3737 ( .A1(n3750), .A2(n3751), .ZN(n3746) );
  OR2_X1 U3738 ( .A1(n3749), .A2(n3748), .ZN(n3751) );
  XOR2_X1 U3739 ( .A(n2636), .B(n3752), .Z(n2629) );
  XOR2_X1 U3740 ( .A(n2635), .B(n2634), .Z(n3752) );
  OR2_X1 U3741 ( .A1(n2279), .A2(n2292), .ZN(n2634) );
  OR2_X1 U3742 ( .A1(n3753), .A2(n3754), .ZN(n2635) );
  AND2_X1 U3743 ( .A1(n3755), .A2(n3756), .ZN(n3754) );
  AND2_X1 U3744 ( .A1(n3757), .A2(n3758), .ZN(n3753) );
  OR2_X1 U3745 ( .A1(n3756), .A2(n3755), .ZN(n3758) );
  XOR2_X1 U3746 ( .A(n2641), .B(n3759), .Z(n2636) );
  XOR2_X1 U3747 ( .A(n2642), .B(n2644), .Z(n3759) );
  OR2_X1 U3748 ( .A1(n2299), .A2(n2271), .ZN(n2644) );
  OR2_X1 U3749 ( .A1(n3760), .A2(n3761), .ZN(n2642) );
  AND2_X1 U3750 ( .A1(n3762), .A2(n3763), .ZN(n3761) );
  AND2_X1 U3751 ( .A1(n3764), .A2(n3765), .ZN(n3760) );
  OR2_X1 U3752 ( .A1(n3763), .A2(n3762), .ZN(n3764) );
  OR2_X1 U3753 ( .A1(n2275), .A2(n2297), .ZN(n2641) );
  XNOR2_X1 U3754 ( .A(n2287), .B(n2621), .ZN(n3744) );
  OR2_X1 U3755 ( .A1(n3766), .A2(n3767), .ZN(n2621) );
  AND2_X1 U3756 ( .A1(n3743), .A2(n3742), .ZN(n3767) );
  AND2_X1 U3757 ( .A1(n3740), .A2(n3768), .ZN(n3766) );
  OR2_X1 U3758 ( .A1(n3742), .A2(n3743), .ZN(n3768) );
  OR2_X1 U3759 ( .A1(n2290), .A2(n2286), .ZN(n3743) );
  OR2_X1 U3760 ( .A1(n3769), .A2(n3770), .ZN(n3742) );
  AND2_X1 U3761 ( .A1(n3739), .A2(n3738), .ZN(n3770) );
  AND2_X1 U3762 ( .A1(n3736), .A2(n3771), .ZN(n3769) );
  OR2_X1 U3763 ( .A1(n3738), .A2(n3739), .ZN(n3771) );
  OR2_X1 U3764 ( .A1(n2292), .A2(n2286), .ZN(n3739) );
  OR2_X1 U3765 ( .A1(n3772), .A2(n3773), .ZN(n3738) );
  AND2_X1 U3766 ( .A1(n3735), .A2(n3734), .ZN(n3773) );
  AND2_X1 U3767 ( .A1(n3732), .A2(n3774), .ZN(n3772) );
  OR2_X1 U3768 ( .A1(n3734), .A2(n3735), .ZN(n3774) );
  OR2_X1 U3769 ( .A1(n2297), .A2(n2286), .ZN(n3735) );
  OR2_X1 U3770 ( .A1(n3775), .A2(n3776), .ZN(n3734) );
  AND2_X1 U3771 ( .A1(n3731), .A2(n3730), .ZN(n3776) );
  AND2_X1 U3772 ( .A1(n3728), .A2(n3777), .ZN(n3775) );
  OR2_X1 U3773 ( .A1(n3730), .A2(n3731), .ZN(n3777) );
  OR2_X1 U3774 ( .A1(n2299), .A2(n2286), .ZN(n3731) );
  OR2_X1 U3775 ( .A1(n3778), .A2(n3779), .ZN(n3730) );
  AND2_X1 U3776 ( .A1(n3724), .A2(n3727), .ZN(n3779) );
  AND2_X1 U3777 ( .A1(n3780), .A2(n3726), .ZN(n3778) );
  OR2_X1 U3778 ( .A1(n3781), .A2(n3782), .ZN(n3726) );
  AND2_X1 U3779 ( .A1(n3723), .A2(n3722), .ZN(n3782) );
  AND2_X1 U3780 ( .A1(n3720), .A2(n3783), .ZN(n3781) );
  OR2_X1 U3781 ( .A1(n3722), .A2(n3723), .ZN(n3783) );
  OR2_X1 U3782 ( .A1(n2306), .A2(n2286), .ZN(n3723) );
  OR2_X1 U3783 ( .A1(n3784), .A2(n3785), .ZN(n3722) );
  AND2_X1 U3784 ( .A1(n3716), .A2(n3719), .ZN(n3785) );
  AND2_X1 U3785 ( .A1(n3786), .A2(n3718), .ZN(n3784) );
  OR2_X1 U3786 ( .A1(n3787), .A2(n3788), .ZN(n3718) );
  AND2_X1 U3787 ( .A1(n3713), .A2(n3715), .ZN(n3788) );
  AND2_X1 U3788 ( .A1(n3789), .A2(n3714), .ZN(n3787) );
  OR2_X1 U3789 ( .A1(n3790), .A2(n3791), .ZN(n3714) );
  AND2_X1 U3790 ( .A1(n3708), .A2(n3711), .ZN(n3791) );
  AND2_X1 U3791 ( .A1(n3710), .A2(n3792), .ZN(n3790) );
  OR2_X1 U3792 ( .A1(n3711), .A2(n3708), .ZN(n3792) );
  OR2_X1 U3793 ( .A1(n2318), .A2(n2286), .ZN(n3708) );
  OR2_X1 U3794 ( .A1(n2755), .A2(n3793), .ZN(n3711) );
  OR2_X1 U3795 ( .A1(n2235), .A2(n2286), .ZN(n3793) );
  INV_X1 U3796 ( .A(n3794), .ZN(n3710) );
  OR2_X1 U3797 ( .A1(n3795), .A2(n3796), .ZN(n3794) );
  AND2_X1 U3798 ( .A1(b_3_), .A2(n3797), .ZN(n3796) );
  OR2_X1 U3799 ( .A1(n3798), .A2(n2043), .ZN(n3797) );
  AND2_X1 U3800 ( .A1(a_14_), .A2(n2279), .ZN(n3798) );
  AND2_X1 U3801 ( .A1(b_2_), .A2(n3799), .ZN(n3795) );
  OR2_X1 U3802 ( .A1(n3800), .A2(n2056), .ZN(n3799) );
  AND2_X1 U3803 ( .A1(a_15_), .A2(n2235), .ZN(n3800) );
  OR2_X1 U3804 ( .A1(n3715), .A2(n3713), .ZN(n3789) );
  XNOR2_X1 U3805 ( .A(n3801), .B(n3802), .ZN(n3713) );
  XNOR2_X1 U3806 ( .A(n3803), .B(n3804), .ZN(n3802) );
  OR2_X1 U3807 ( .A1(n2313), .A2(n2286), .ZN(n3715) );
  OR2_X1 U3808 ( .A1(n3719), .A2(n3716), .ZN(n3786) );
  XNOR2_X1 U3809 ( .A(n3805), .B(n3806), .ZN(n3716) );
  XNOR2_X1 U3810 ( .A(n3807), .B(n3808), .ZN(n3805) );
  OR2_X1 U3811 ( .A1(n2311), .A2(n2286), .ZN(n3719) );
  XOR2_X1 U3812 ( .A(n3809), .B(n3810), .Z(n3720) );
  XOR2_X1 U3813 ( .A(n3811), .B(n3812), .Z(n3810) );
  OR2_X1 U3814 ( .A1(n3727), .A2(n3724), .ZN(n3780) );
  XOR2_X1 U3815 ( .A(n3813), .B(n3814), .Z(n3724) );
  XOR2_X1 U3816 ( .A(n3815), .B(n3816), .Z(n3814) );
  OR2_X1 U3817 ( .A1(n2304), .A2(n2286), .ZN(n3727) );
  INV_X1 U3818 ( .A(b_4_), .ZN(n2286) );
  XOR2_X1 U3819 ( .A(n3817), .B(n3818), .Z(n3728) );
  XOR2_X1 U3820 ( .A(n3819), .B(n3820), .Z(n3818) );
  XOR2_X1 U3821 ( .A(n3821), .B(n3822), .Z(n3732) );
  XOR2_X1 U3822 ( .A(n3823), .B(n3824), .Z(n3822) );
  XOR2_X1 U3823 ( .A(n3825), .B(n3826), .Z(n3736) );
  XOR2_X1 U3824 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR2_X1 U3825 ( .A(n3750), .B(n3829), .Z(n3740) );
  XOR2_X1 U3826 ( .A(n3749), .B(n3748), .Z(n3829) );
  OR2_X1 U3827 ( .A1(n2292), .A2(n2235), .ZN(n3748) );
  OR2_X1 U3828 ( .A1(n3830), .A2(n3831), .ZN(n3749) );
  AND2_X1 U3829 ( .A1(n3828), .A2(n3827), .ZN(n3831) );
  AND2_X1 U3830 ( .A1(n3825), .A2(n3832), .ZN(n3830) );
  OR2_X1 U3831 ( .A1(n3827), .A2(n3828), .ZN(n3832) );
  OR2_X1 U3832 ( .A1(n2297), .A2(n2235), .ZN(n3828) );
  OR2_X1 U3833 ( .A1(n3833), .A2(n3834), .ZN(n3827) );
  AND2_X1 U3834 ( .A1(n3824), .A2(n3823), .ZN(n3834) );
  AND2_X1 U3835 ( .A1(n3821), .A2(n3835), .ZN(n3833) );
  OR2_X1 U3836 ( .A1(n3823), .A2(n3824), .ZN(n3835) );
  OR2_X1 U3837 ( .A1(n2299), .A2(n2235), .ZN(n3824) );
  OR2_X1 U3838 ( .A1(n3836), .A2(n3837), .ZN(n3823) );
  AND2_X1 U3839 ( .A1(n3820), .A2(n3819), .ZN(n3837) );
  AND2_X1 U3840 ( .A1(n3817), .A2(n3838), .ZN(n3836) );
  OR2_X1 U3841 ( .A1(n3819), .A2(n3820), .ZN(n3838) );
  OR2_X1 U3842 ( .A1(n2304), .A2(n2235), .ZN(n3820) );
  OR2_X1 U3843 ( .A1(n3839), .A2(n3840), .ZN(n3819) );
  AND2_X1 U3844 ( .A1(n3813), .A2(n3816), .ZN(n3840) );
  AND2_X1 U3845 ( .A1(n3841), .A2(n3815), .ZN(n3839) );
  OR2_X1 U3846 ( .A1(n3842), .A2(n3843), .ZN(n3815) );
  AND2_X1 U3847 ( .A1(n3812), .A2(n3811), .ZN(n3843) );
  AND2_X1 U3848 ( .A1(n3809), .A2(n3844), .ZN(n3842) );
  OR2_X1 U3849 ( .A1(n3811), .A2(n3812), .ZN(n3844) );
  OR2_X1 U3850 ( .A1(n2311), .A2(n2235), .ZN(n3812) );
  OR2_X1 U3851 ( .A1(n3845), .A2(n3846), .ZN(n3811) );
  AND2_X1 U3852 ( .A1(n3806), .A2(n3808), .ZN(n3846) );
  AND2_X1 U3853 ( .A1(n3847), .A2(n3807), .ZN(n3845) );
  OR2_X1 U3854 ( .A1(n3848), .A2(n3849), .ZN(n3807) );
  AND2_X1 U3855 ( .A1(n3801), .A2(n3804), .ZN(n3849) );
  AND2_X1 U3856 ( .A1(n3803), .A2(n3850), .ZN(n3848) );
  OR2_X1 U3857 ( .A1(n3804), .A2(n3801), .ZN(n3850) );
  OR2_X1 U3858 ( .A1(n2318), .A2(n2235), .ZN(n3801) );
  OR2_X1 U3859 ( .A1(n2755), .A2(n3851), .ZN(n3804) );
  OR2_X1 U3860 ( .A1(n2279), .A2(n2235), .ZN(n3851) );
  INV_X1 U3861 ( .A(n3852), .ZN(n3803) );
  OR2_X1 U3862 ( .A1(n3853), .A2(n3854), .ZN(n3852) );
  AND2_X1 U3863 ( .A1(b_2_), .A2(n3855), .ZN(n3854) );
  OR2_X1 U3864 ( .A1(n3856), .A2(n2043), .ZN(n3855) );
  AND2_X1 U3865 ( .A1(a_14_), .A2(n2275), .ZN(n3856) );
  AND2_X1 U3866 ( .A1(b_1_), .A2(n3857), .ZN(n3853) );
  OR2_X1 U3867 ( .A1(n3858), .A2(n2056), .ZN(n3857) );
  AND2_X1 U3868 ( .A1(a_15_), .A2(n2279), .ZN(n3858) );
  OR2_X1 U3869 ( .A1(n3808), .A2(n3806), .ZN(n3847) );
  XNOR2_X1 U3870 ( .A(n3859), .B(n3860), .ZN(n3806) );
  XNOR2_X1 U3871 ( .A(n3861), .B(n3862), .ZN(n3860) );
  OR2_X1 U3872 ( .A1(n2313), .A2(n2235), .ZN(n3808) );
  XNOR2_X1 U3873 ( .A(n3863), .B(n3864), .ZN(n3809) );
  XNOR2_X1 U3874 ( .A(n3865), .B(n3866), .ZN(n3863) );
  OR2_X1 U3875 ( .A1(n3816), .A2(n3813), .ZN(n3841) );
  XOR2_X1 U3876 ( .A(n3867), .B(n3868), .Z(n3813) );
  XOR2_X1 U3877 ( .A(n3869), .B(n3870), .Z(n3868) );
  OR2_X1 U3878 ( .A1(n2306), .A2(n2235), .ZN(n3816) );
  INV_X1 U3879 ( .A(b_3_), .ZN(n2235) );
  XOR2_X1 U3880 ( .A(n3871), .B(n3872), .Z(n3817) );
  XOR2_X1 U3881 ( .A(n3873), .B(n3874), .Z(n3872) );
  XOR2_X1 U3882 ( .A(n3875), .B(n3876), .Z(n3821) );
  XOR2_X1 U3883 ( .A(n3877), .B(n3878), .Z(n3876) );
  XOR2_X1 U3884 ( .A(n3879), .B(n3880), .Z(n3825) );
  XOR2_X1 U3885 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR2_X1 U3886 ( .A(n3757), .B(n3883), .Z(n3750) );
  XOR2_X1 U3887 ( .A(n3756), .B(n3755), .Z(n3883) );
  OR2_X1 U3888 ( .A1(n2279), .A2(n2297), .ZN(n3755) );
  OR2_X1 U3889 ( .A1(n3884), .A2(n3885), .ZN(n3756) );
  AND2_X1 U3890 ( .A1(n3882), .A2(n3881), .ZN(n3885) );
  AND2_X1 U3891 ( .A1(n3879), .A2(n3886), .ZN(n3884) );
  OR2_X1 U3892 ( .A1(n3881), .A2(n3882), .ZN(n3886) );
  OR2_X1 U3893 ( .A1(n2279), .A2(n2299), .ZN(n3882) );
  OR2_X1 U3894 ( .A1(n3887), .A2(n3888), .ZN(n3881) );
  AND2_X1 U3895 ( .A1(n3878), .A2(n3877), .ZN(n3888) );
  AND2_X1 U3896 ( .A1(n3875), .A2(n3889), .ZN(n3887) );
  OR2_X1 U3897 ( .A1(n3877), .A2(n3878), .ZN(n3889) );
  OR2_X1 U3898 ( .A1(n2279), .A2(n2304), .ZN(n3878) );
  OR2_X1 U3899 ( .A1(n3890), .A2(n3891), .ZN(n3877) );
  AND2_X1 U3900 ( .A1(n3874), .A2(n3873), .ZN(n3891) );
  AND2_X1 U3901 ( .A1(n3871), .A2(n3892), .ZN(n3890) );
  OR2_X1 U3902 ( .A1(n3873), .A2(n3874), .ZN(n3892) );
  OR2_X1 U3903 ( .A1(n2279), .A2(n2306), .ZN(n3874) );
  OR2_X1 U3904 ( .A1(n3893), .A2(n3894), .ZN(n3873) );
  AND2_X1 U3905 ( .A1(n3867), .A2(n3870), .ZN(n3894) );
  AND2_X1 U3906 ( .A1(n3895), .A2(n3869), .ZN(n3893) );
  OR2_X1 U3907 ( .A1(n3896), .A2(n3897), .ZN(n3869) );
  AND2_X1 U3908 ( .A1(n3866), .A2(n3865), .ZN(n3897) );
  AND2_X1 U3909 ( .A1(n3864), .A2(n3898), .ZN(n3896) );
  OR2_X1 U3910 ( .A1(n3865), .A2(n3866), .ZN(n3898) );
  OR2_X1 U3911 ( .A1(n2279), .A2(n2313), .ZN(n3866) );
  OR2_X1 U3912 ( .A1(n3899), .A2(n3900), .ZN(n3865) );
  AND2_X1 U3913 ( .A1(n3859), .A2(n3862), .ZN(n3900) );
  AND2_X1 U3914 ( .A1(n3861), .A2(n3901), .ZN(n3899) );
  OR2_X1 U3915 ( .A1(n3862), .A2(n3859), .ZN(n3901) );
  OR2_X1 U3916 ( .A1(n2279), .A2(n2318), .ZN(n3859) );
  OR2_X1 U3917 ( .A1(n2755), .A2(n3902), .ZN(n3862) );
  OR2_X1 U3918 ( .A1(n2275), .A2(n2279), .ZN(n3902) );
  INV_X1 U3919 ( .A(n3903), .ZN(n3861) );
  OR2_X1 U3920 ( .A1(n3904), .A2(n3905), .ZN(n3903) );
  AND2_X1 U3921 ( .A1(b_1_), .A2(n3906), .ZN(n3905) );
  OR2_X1 U3922 ( .A1(n3907), .A2(n2043), .ZN(n3906) );
  AND2_X1 U3923 ( .A1(n2322), .A2(a_14_), .ZN(n2043) );
  AND2_X1 U3924 ( .A1(a_14_), .A2(n2271), .ZN(n3907) );
  AND2_X1 U3925 ( .A1(b_0_), .A2(n3908), .ZN(n3904) );
  OR2_X1 U3926 ( .A1(n3909), .A2(n2056), .ZN(n3908) );
  AND2_X1 U3927 ( .A1(n2048), .A2(a_15_), .ZN(n2056) );
  AND2_X1 U3928 ( .A1(a_15_), .A2(n2275), .ZN(n3909) );
  XNOR2_X1 U3929 ( .A(n3910), .B(n3911), .ZN(n3864) );
  OR2_X1 U3930 ( .A1(n3912), .A2(n3913), .ZN(n3910) );
  INV_X1 U3931 ( .A(n3914), .ZN(n3913) );
  AND2_X1 U3932 ( .A1(n3915), .A2(n3916), .ZN(n3912) );
  OR2_X1 U3933 ( .A1(n3870), .A2(n3867), .ZN(n3895) );
  XOR2_X1 U3934 ( .A(n3917), .B(n3918), .Z(n3867) );
  XOR2_X1 U3935 ( .A(n3919), .B(n3920), .Z(n3917) );
  OR2_X1 U3936 ( .A1(n2279), .A2(n2311), .ZN(n3870) );
  INV_X1 U3937 ( .A(b_2_), .ZN(n2279) );
  XNOR2_X1 U3938 ( .A(n3921), .B(n3922), .ZN(n3871) );
  XNOR2_X1 U3939 ( .A(n3923), .B(n3924), .ZN(n3921) );
  XNOR2_X1 U3940 ( .A(n3925), .B(n3926), .ZN(n3875) );
  XNOR2_X1 U3941 ( .A(n3927), .B(n3928), .ZN(n3925) );
  XNOR2_X1 U3942 ( .A(n3929), .B(n3930), .ZN(n3879) );
  XNOR2_X1 U3943 ( .A(n3931), .B(n3932), .ZN(n3929) );
  XOR2_X1 U3944 ( .A(n3762), .B(n3933), .Z(n3757) );
  XOR2_X1 U3945 ( .A(n3763), .B(n3765), .Z(n3933) );
  OR2_X1 U3946 ( .A1(n2304), .A2(n2271), .ZN(n3765) );
  OR2_X1 U3947 ( .A1(n3934), .A2(n3935), .ZN(n3763) );
  AND2_X1 U3948 ( .A1(n3930), .A2(n3932), .ZN(n3935) );
  AND2_X1 U3949 ( .A1(n3936), .A2(n3931), .ZN(n3934) );
  OR2_X1 U3950 ( .A1(n2306), .A2(n2271), .ZN(n3931) );
  OR2_X1 U3951 ( .A1(n3932), .A2(n3930), .ZN(n3936) );
  OR2_X1 U3952 ( .A1(n2275), .A2(n2304), .ZN(n3930) );
  OR2_X1 U3953 ( .A1(n3937), .A2(n3938), .ZN(n3932) );
  AND2_X1 U3954 ( .A1(n3926), .A2(n3928), .ZN(n3938) );
  AND2_X1 U3955 ( .A1(n3939), .A2(n3927), .ZN(n3937) );
  OR2_X1 U3956 ( .A1(n2311), .A2(n2271), .ZN(n3927) );
  OR2_X1 U3957 ( .A1(n3928), .A2(n3926), .ZN(n3939) );
  OR2_X1 U3958 ( .A1(n2275), .A2(n2306), .ZN(n3926) );
  OR2_X1 U3959 ( .A1(n3940), .A2(n3941), .ZN(n3928) );
  AND2_X1 U3960 ( .A1(n3922), .A2(n3924), .ZN(n3941) );
  AND2_X1 U3961 ( .A1(n3942), .A2(n3923), .ZN(n3940) );
  OR2_X1 U3962 ( .A1(n2313), .A2(n2271), .ZN(n3923) );
  OR2_X1 U3963 ( .A1(n3924), .A2(n3922), .ZN(n3942) );
  OR2_X1 U3964 ( .A1(n2275), .A2(n2311), .ZN(n3922) );
  OR2_X1 U3965 ( .A1(n3943), .A2(n3944), .ZN(n3924) );
  AND2_X1 U3966 ( .A1(n3918), .A2(n3920), .ZN(n3944) );
  AND2_X1 U3967 ( .A1(n3919), .A2(n3945), .ZN(n3943) );
  OR2_X1 U3968 ( .A1(n3920), .A2(n3918), .ZN(n3945) );
  OR2_X1 U3969 ( .A1(n2275), .A2(n2313), .ZN(n3918) );
  OR2_X1 U3970 ( .A1(n2318), .A2(n2271), .ZN(n3920) );
  AND2_X1 U3971 ( .A1(n3914), .A2(n3911), .ZN(n3919) );
  OR2_X1 U3972 ( .A1(n2755), .A2(n3946), .ZN(n3911) );
  OR2_X1 U3973 ( .A1(n2275), .A2(n2271), .ZN(n3946) );
  OR2_X1 U3974 ( .A1(n3916), .A2(n3915), .ZN(n3914) );
  OR2_X1 U3975 ( .A1(n2048), .A2(n2271), .ZN(n3915) );
  INV_X1 U3976 ( .A(b_0_), .ZN(n2271) );
  OR2_X1 U3977 ( .A1(n2275), .A2(n2318), .ZN(n3916) );
  OR2_X1 U3978 ( .A1(n2275), .A2(n2299), .ZN(n3762) );
  INV_X1 U3979 ( .A(b_1_), .ZN(n2275) );
  INV_X1 U3980 ( .A(n2210), .ZN(n2287) );
  AND2_X1 U3981 ( .A1(a_4_), .A2(b_4_), .ZN(n2210) );
  INV_X1 U3982 ( .A(n2034), .ZN(n1989) );
  OR2_X1 U3983 ( .A1(n3947), .A2(n3948), .ZN(n2034) );
  AND2_X1 U3984 ( .A1(b_0_), .A2(n2427), .ZN(n3948) );
  AND2_X1 U3985 ( .A1(n3949), .A2(n3950), .ZN(n3947) );
  OR2_X1 U3986 ( .A1(b_0_), .A2(n2427), .ZN(n3950) );
  INV_X1 U3987 ( .A(a_0_), .ZN(n2427) );
  AND2_X1 U3988 ( .A1(n2259), .A2(n3951), .ZN(n3949) );
  OR2_X1 U3989 ( .A1(n3952), .A2(n3953), .ZN(n3951) );
  OR2_X1 U3990 ( .A1(n2260), .A2(n3954), .ZN(n3953) );
  AND2_X1 U3991 ( .A1(b_2_), .A2(n2278), .ZN(n3954) );
  AND2_X1 U3992 ( .A1(n2274), .A2(b_1_), .ZN(n2260) );
  AND2_X1 U3993 ( .A1(n3955), .A2(n3956), .ZN(n3952) );
  OR2_X1 U3994 ( .A1(b_3_), .A2(n2283), .ZN(n3956) );
  AND2_X1 U3995 ( .A1(n3957), .A2(n3958), .ZN(n3955) );
  OR2_X1 U3996 ( .A1(n3959), .A2(n3960), .ZN(n3958) );
  OR2_X1 U3997 ( .A1(n3961), .A2(n2233), .ZN(n3960) );
  AND2_X1 U3998 ( .A1(n2283), .A2(b_3_), .ZN(n2233) );
  INV_X1 U3999 ( .A(a_3_), .ZN(n2283) );
  AND2_X1 U4000 ( .A1(n3962), .A2(n3963), .ZN(n3961) );
  OR2_X1 U4001 ( .A1(b_5_), .A2(n2290), .ZN(n3963) );
  AND2_X1 U4002 ( .A1(n3964), .A2(n3965), .ZN(n3962) );
  OR2_X1 U4003 ( .A1(n2196), .A2(n3966), .ZN(n3965) );
  OR2_X1 U4004 ( .A1(n3967), .A2(n3968), .ZN(n3966) );
  AND2_X1 U4005 ( .A1(b_6_), .A2(n2292), .ZN(n3968) );
  AND2_X1 U4006 ( .A1(n3969), .A2(n3970), .ZN(n3967) );
  OR2_X1 U4007 ( .A1(b_7_), .A2(n2297), .ZN(n3970) );
  AND2_X1 U4008 ( .A1(n3971), .A2(n3972), .ZN(n3969) );
  OR2_X1 U4009 ( .A1(n2166), .A2(n3973), .ZN(n3972) );
  OR2_X1 U4010 ( .A1(n3974), .A2(n3975), .ZN(n3973) );
  AND2_X1 U4011 ( .A1(b_8_), .A2(n2299), .ZN(n3975) );
  AND2_X1 U4012 ( .A1(n3976), .A2(n3977), .ZN(n3974) );
  OR2_X1 U4013 ( .A1(b_9_), .A2(n2304), .ZN(n3977) );
  AND2_X1 U4014 ( .A1(n3978), .A2(n3979), .ZN(n3976) );
  OR2_X1 U4015 ( .A1(n2136), .A2(n3980), .ZN(n3979) );
  OR2_X1 U4016 ( .A1(n3981), .A2(n3982), .ZN(n3980) );
  AND2_X1 U4017 ( .A1(b_10_), .A2(n2306), .ZN(n3982) );
  AND2_X1 U4018 ( .A1(n3983), .A2(n3984), .ZN(n3981) );
  OR2_X1 U4019 ( .A1(b_11_), .A2(n2311), .ZN(n3984) );
  AND2_X1 U4020 ( .A1(n3985), .A2(n3986), .ZN(n3983) );
  OR2_X1 U4021 ( .A1(n2106), .A2(n3987), .ZN(n3986) );
  OR2_X1 U4022 ( .A1(n3988), .A2(n3989), .ZN(n3987) );
  AND2_X1 U4023 ( .A1(b_12_), .A2(n2313), .ZN(n3989) );
  AND2_X1 U4024 ( .A1(n3990), .A2(n3991), .ZN(n3988) );
  OR2_X1 U4025 ( .A1(b_13_), .A2(n2318), .ZN(n3991) );
  AND2_X1 U4026 ( .A1(n3992), .A2(n3993), .ZN(n3990) );
  OR2_X1 U4027 ( .A1(n2073), .A2(n3994), .ZN(n3993) );
  OR2_X1 U4028 ( .A1(n3995), .A2(n3996), .ZN(n3994) );
  AND2_X1 U4029 ( .A1(n2322), .A2(n2048), .ZN(n3996) );
  AND2_X1 U4030 ( .A1(n3997), .A2(n3998), .ZN(n3995) );
  OR2_X1 U4031 ( .A1(b_15_), .A2(n3999), .ZN(n3998) );
  AND2_X1 U4032 ( .A1(b_14_), .A2(n2755), .ZN(n3999) );
  OR2_X1 U4033 ( .A1(n2048), .A2(n2322), .ZN(n2755) );
  INV_X1 U4034 ( .A(a_15_), .ZN(n2322) );
  INV_X1 U4035 ( .A(a_14_), .ZN(n2048) );
  INV_X1 U4036 ( .A(n2042), .ZN(n3997) );
  AND2_X1 U4037 ( .A1(n2049), .A2(a_14_), .ZN(n2042) );
  INV_X1 U4038 ( .A(b_14_), .ZN(n2049) );
  AND2_X1 U4039 ( .A1(n2318), .A2(b_13_), .ZN(n2073) );
  INV_X1 U4040 ( .A(a_13_), .ZN(n2318) );
  OR2_X1 U4041 ( .A1(b_12_), .A2(n2313), .ZN(n3992) );
  INV_X1 U4042 ( .A(a_12_), .ZN(n2313) );
  AND2_X1 U4043 ( .A1(n2311), .A2(b_11_), .ZN(n2106) );
  INV_X1 U4044 ( .A(a_11_), .ZN(n2311) );
  OR2_X1 U4045 ( .A1(b_10_), .A2(n2306), .ZN(n3985) );
  INV_X1 U4046 ( .A(a_10_), .ZN(n2306) );
  AND2_X1 U4047 ( .A1(n2304), .A2(b_9_), .ZN(n2136) );
  INV_X1 U4048 ( .A(a_9_), .ZN(n2304) );
  OR2_X1 U4049 ( .A1(b_8_), .A2(n2299), .ZN(n3978) );
  INV_X1 U4050 ( .A(a_8_), .ZN(n2299) );
  AND2_X1 U4051 ( .A1(n2297), .A2(b_7_), .ZN(n2166) );
  INV_X1 U4052 ( .A(a_7_), .ZN(n2297) );
  OR2_X1 U4053 ( .A1(b_6_), .A2(n2292), .ZN(n3971) );
  INV_X1 U4054 ( .A(a_6_), .ZN(n2292) );
  AND2_X1 U4055 ( .A1(n2290), .A2(b_5_), .ZN(n2196) );
  INV_X1 U4056 ( .A(a_5_), .ZN(n2290) );
  OR2_X1 U4057 ( .A1(b_4_), .A2(n2285), .ZN(n3964) );
  AND2_X1 U4058 ( .A1(b_4_), .A2(n2285), .ZN(n3959) );
  INV_X1 U4059 ( .A(a_4_), .ZN(n2285) );
  OR2_X1 U4060 ( .A1(b_2_), .A2(n2278), .ZN(n3957) );
  INV_X1 U4061 ( .A(a_2_), .ZN(n2278) );
  OR2_X1 U4062 ( .A1(b_1_), .A2(n2274), .ZN(n2259) );
  INV_X1 U4063 ( .A(a_1_), .ZN(n2274) );
endmodule

