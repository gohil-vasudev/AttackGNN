module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   g100, g101, g102, g103, g104, g1170, g1173, g1176, g1179, g1182,
         g1185, g1188, g1191, g1194, g1197, g1203, g18, g1960, g1961, g27, g28,
         g29, g30, g31, g41, g42, g43, g44, g45, g46, g47, g48, g5816, g82,
         g83, g84, g85, g8561, g8562, g8563, g8564, g8565, g8566, g86, g87,
         g872, g873, g88, g886, g889, g89, g892, g895, g898, g90, g901, g904,
         g907, g91, g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451,
         g95, g96, g99, test_so10, g10722, g10664, g4556, g1289, g8943, g1882,
         n1663, g255, g312, g11257, g452, g7032, g123, g6830, g207, g8920,
         g713, g4340, g1153, n1686, g4239, g1744, g6538, g1558, g8887, g695,
         g11372, g461, n1594, g8260, g940, n1712, g11391, g976, g8432, g709,
         g6088, g1092, g6478, g1574, g6795, g1864, g11320, g369, g6500, g1580,
         g5392, g1736, g10663, n1637, n3065, g6216, g1424, g1737, g10858,
         g1672, g5914, g1077, g7590, g1231, g6656, g4, g5126, g1104, n1658,
         g7290, g1304, g6841, g243, g8041, g1499, g8766, g1444, n3064, g8019,
         g6545, g1543, g256, g315, g6533, g1534, n1632, g8820, g622, n1713,
         g8941, g1927, g10859, g1660, g6922, g278, g8772, g1436, g8433, g718,
         g6526, n1669, g10793, g554, g11333, g496, n1689, g11392, g981, n1720,
         g794, g829, g6093, g1095, g8889, g704, g7302, g1265, g6525, g1786,
         g8429, g682, g7292, g1296, g6621, n1668, g7134, n3062, g260, g327,
         g6333, g1389, n1603, g6826, g1371, g1955, g1956, g10860, g1675,
         g11483, g354, g6392, g113, g7626, g639, n1692, g10866, g1684, g8193,
         g1639, g6983, g1791, n1702, g6839, g248, n1598, g4076, g1707, g4293,
         g1759, g11482, g351, g6507, g1604, g6096, g1098, g8250, g932, n1591,
         g8282, g1896, g8435, g736, g6924, g1019, g6819, n3061, g746, g745,
         g6244, g1419, n1602, g6627, n1667, g32, n1865, g6071, g1086, g8046,
         g1486, g10707, g1730, g6198, g1504, g8051, g1470, g8024, g822, g10862,
         g1678, g8050, g174, g7133, g1766, g7930, g1801, g6832, g186, g11308,
         g959, g6918, g8769, g1407, g6909, g1868, g4940, g5404, g1718, n1611,
         g11265, g396, g6930, g1015, n1650, g4891, n3059, g6224, g1415, g7586,
         g1227, g10770, g1721, n3058, n3057, g284, g11256, g426, g6824, g219,
         g1360, n3056, DFF_126_n1, g6126, g806, g8767, g1428, g6546, g1564,
         g4238, g1741, n1633, g6823, g225, g281, g11602, g1308, g9721, g611,
         n1609, g4890, n3055, DFF_136_n1, n1586, g1217, g6524, g1589, g8045,
         g1466, g6469, g1571, g6471, g1861, g6821, n3054, g11514, g1448, g4480,
         g1133, n1706, g11610, g1333, g7843, g153, g11310, g962, g11331, g486,
         n1621, g11380, g471, n1606, g6838, g1397, n1711, g8288, g1950, g755,
         g756, g4892, n3053, DFF_157_n1, g10855, g1101, g549, g10898, g105,
         g10865, g1669, g6822, g1531, n1652, g6180, g1458, n1703, g10718, g572,
         g6912, g1011, g10719, n3051, g6234, g1411, g6099, g1074, g11259, g444,
         g8039, g1474, g6059, g1080, g5396, g1713, n1610, g262, g333, g6906,
         g269, g11266, g401, g11294, g1857, n1682, g5421, g9, g8649, g664,
         g11312, g965, g6840, g1400, n1629, g254, g309, g7202, g814, g6834,
         g231, g10795, g557, g875, g869, g6831, g1383, g8060, g158, g4893,
         g627, n1701, g7244, g1023, g6026, g259, n3050, g11608, g1327, g7660,
         g654, g6911, g293, g11640, g1346, g8777, g1633, g4274, g1753, g1508,
         g7297, g1240, g11326, g538, g11269, g416, g11325, g542, g10864, g1681,
         g11290, g374, g10798, g563, g8284, g1914, g11328, g530, g10800, g575,
         g8944, g1936, n1694, g7183, n1674, g4465, g1356, g1317, g11484, g357,
         g11263, g386, g6501, g1601, g6757, g166, g11334, g501, g6042, g8384,
         g1840, g6653, n1666, g257, g318, g5849, n3048, DFF_228_n1, g6929,
         g302, g11488, g342, g7299, g1250, g4330, g1163, g1958, n3047, g7257,
         g1032, g8775, g1432, g5770, g1453, n1628, g11486, g363, g261, g330,
         g4338, g1157, g4500, n3046, g10721, n3045, DFF_242_n1, g8147, g928,
         n1604, g6038, g11337, g516, n1620, g6045, g7191, g826, g861, g8774,
         g1627, g7293, g1292, g6907, g290, g4903, n3044, g6123, g6506, g1583,
         g11376, g466, n1646, g6542, g1561, g6551, g1546, g6901, g287, g10797,
         g560, g8505, g617, n1645, n1631, g11647, g336, g11340, g456, n1641,
         g253, g305, n1681, g11625, g345, g636, g8, g6502, N599, g6049, g8945,
         g1945, n1697, g4231, g1738, n1640, g8040, g1478, n3042, DFF_275_n1,
         g6155, g1690, n1653, g8043, g1482, g5173, g1110, n1677, g6916, g296,
         g10861, g1663, g8431, g700, g4309, g1762, g11485, g360, g6334, g192,
         g10767, g1657, g8923, g722, n1693, g7189, n1673, g10799, g566, g6747,
         n3041, g6080, g1089, g3381, g5910, g1071, g11393, g986, n1722, g11349,
         g971, g6439, g143, g9266, g1814, n1608, g1212, g8940, g1918, g9269,
         g1822, n1643, g6820, g237, g8042, g1462, g6759, g178, g11487, g366,
         g802, g837, g9124, g599, n1644, g11293, g1854, g11298, g944, g8287,
         g1941, g8047, g170, g6205, g1520, n1710, g8885, g686, n1676, g11305,
         g953, g5556, n3040, g2478, g1765, g10711, g1733, g7303, g5194, g1610,
         g7541, g1796, n1626, g11607, g1324, g1540, g6827, n3038, g11332, g491,
         n1691, g4902, n3037, DFF_330_n1, g6828, g213, g6516, g1781, n1659,
         g8938, g1900, n1675, g7298, g1245, n3036, g6672, n3035, DFF_336_n1,
         g8048, g148, g798, g833, g8285, g1923, n1718, g8254, g936, n1630,
         g11604, g1314, g849, g11636, g1336, g6910, g272, g8173, g1806, g8245,
         n1716, g8281, g1887, n3034, g11314, g968, g4905, n3033, g4484, g1137,
         n1597, g8937, g1891, n1657, g7300, g1255, g6002, n1588, g874, g9110,
         g591, n1607, g8926, g731, n1696, g8631, g7632, g1218, g9150, g605,
         n1593, g6531, n1665, g6786, g182, g950, g4477, g1129, n1705, g857,
         g11258, g448, g9272, g1828, n1605, g10773, g1727, g1592, g5083, g1703,
         g8286, g1932, g8773, g1624, g6054, g11260, g440, g11338, g476, n1599,
         g5918, g119, n1613, g8922, g668, n1662, g8049, g139, g4342, g1149,
         n1685, g10720, n3031, g6755, n3030, DFF_385_n1, g6897, g263, g7709,
         g818, g4255, g1747, g5543, n1622, g6915, g275, g6513, g1524, n1649,
         g6480, g1577, g810, g11264, g391, g8973, g658, n1615, g6833, g1386,
         g5996, n1587, g4473, g1125, n1708, g5755, g201, n1619, g7295, g1280,
         n1862, g6068, g1083, g7137, g650, n1709, g8779, g1636, g853, g11270,
         g421, g5529, g11306, g956, g11291, g378, g4283, g1756, g841, g6894,
         g1027, g6902, g1003, g8765, g1403, g4498, g1145, n1617, g5148, g1107,
         n1614, g7581, g1223, g11267, g406, g10936, g1811, n1699, n3029,
         g10765, g1654, g197, n1678, g6479, g1595, g6537, g1537, g8434, g727,
         g6908, g6243, n1717, g11324, g481, g3462, n1647, g11609, g1330, g845,
         g8244, g8194, g1512, n3027, g8052, g1490, g4325, g1166, g11481, g348,
         n3026, DFF_441_n1, g7301, g1260, g6035, g8059, g131, n3025, g6015,
         g258, g11330, g521, n1698, g11605, g1318, g8921, g1872, n1616, g8883,
         g677, n1656, n3024, g6523, g1549, g947, g1834, n1655, g6481, g1598,
         g4471, g1121, n1618, g11606, g1321, g11335, g506, n1600, g10791, g546,
         g8939, g1909, g6529, g1552, g10776, g1687, g1586, g324, g4490, g1141,
         n1660, g11639, g1341, g4089, g1710, n3023, n3022, g8053, g135, g11329,
         g525, n1695, g6515, g1607, g321, g7204, n1672, g11443, g1275, g11603,
         g8770, g1615, g11292, g382, g6331, n3020, g6900, g266, g7294, g1284,
         n1864, g6829, n3019, g8428, g673, n3018, DFF_489_n1, g8054, g162,
         g11268, g411, g11262, g431, g8283, g1905, g6193, g1515, n1627, g8776,
         g1630, g7143, n1671, g6898, g991, n1871, g7291, g1300, g11478, g339,
         g6000, g4264, g1750, g8768, g1440, g10863, g1666, g1528, n1635,
         g11641, g1351, n1721, n3017, g8044, g127, n1704, g11579, g1618, g7296,
         g1235, g6923, g299, g11261, g435, n1878, g6638, n1664, g1555, g6895,
         g995, g8771, g1621, g4506, n3016, g7441, g643, g8055, g1494, g1567,
         g8430, g691, g11327, g534, g6508, g1776, n1715, g10717, g569, g4334,
         g1160, n1585, g6679, g1, g11336, g511, n1679, g10771, g1724, g5445,
         g12, g8559, g1878, g7219, g5390, n1654, n1512, n1486, n1485, n1544,
         n1530, n1420, n1855, n1239, n1566, n1567, n1479, n1858, n1480, n1546,
         n1478, n968, n1137, n1195, n1404, n1262, n1227, n1450, n916, n822,
         n958, n918, n1054, n1116, n1159, n812, n1057, n1056, n1258, n817,
         n929, n837, n804, n1016, n1380, n926, n1385, n1391, n1564, n1231,
         n1232, n1260, n1107, n1093, n1214, n931, n962, n1193, n1153, n1125,
         n1099, n917, n806, n1097, n1123, n1151, n1090, n967, n921, n898,
         n1055, n1150, n1096, n1098, n1213, n1152, n836, n838, Tg1_OUT1,
         Tg1_OUT2, Tg1_OUT3, Tg1_OUT4, Tg1_OUT5, Tg1_OUT6, Tg1_OUT7, Tg1_OUT8,
         Tg2_OUT1, Tg2_OUT2, Tg2_OUT3, Tg2_OUT4, Tg2_OUT5, Tg2_OUT6, Tg2_OUT7,
         Tg2_OUT8, test_se_NOT, Trigger_select, n2, n9, n13, n23, n34, n37,
         n38, n39, n49, n50, n55, n62, n63, n69, n80, n81, n82, n91, n99, n100,
         n101, n140, n142, n145, n147, n148, n151, n152, n154, n160, n167,
         n170, n185, n224, n228, n248, n249, n250, n275, n319, n342, n363,
         n364, n365, n366, n367, n438, n487, n497, n507, n508, n510, n523,
         n527, n2636, n2637, n2638, n2640, n2641, n2642, n2645, n2646, n2647,
         n2648, n2650, n2652, n2653, n2655, n2657, n2658, n2659, n2660, n2661,
         n2662, n2665, n2667, n2670, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2692, n2693, n2694, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2708, n2709, n2710, n2711, n2712, n2713, n2715,
         n2717, n2718, n2721, n2723, n2724, n2725, n2727, n2729, n2730, n2731,
         n2735, n2736, n2737, n2738, n2752, n2755, n2757, n2758, n2759, n2764,
         n2766, n2784, n2785, n2787, n2788, n2789, n2791, n2792, n2793, n2794,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2808, n2810,
         n2811, n2812, n2813, n2814, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2829, n2830, n2832, n2834,
         n2835, n2836, n2837, n2838, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2849, n2850, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2862, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2885,
         n2887, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2897, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3021, n3028, n3032, n3039,
         n3043, n3049, n3052, n3060, n3063, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, U1550_n1, U1551_n1, U1586_n1, U1754_n1,
         U1798_n1, U1839_n1, U1843_n1, U1877_n1, U1908_n1, U1909_n1, U1987_n1,
         U2031_n1, U2035_n1, U2418_n1, U2468_n1, U2478_n1, U2488_n1, U2533_n1,
         U2534_n1, U2639_n1, U2641_n1, U2654_n1, U2658_n1, U2683_n1, U2699_n1,
         U2846_n1, U2847_n1, U2848_n1, U2859_n1, U2860_n1, U2861_n1, U2867_n1,
         U2879_n1, U2881_n1, U2882_n1, U2883_n1, U2884_n1, U2885_n1, U2886_n1,
         U2887_n1, U2888_n1, U2889_n1, U2890_n1, U2891_n1, U2892_n1, U2893_n1,
         U2894_n1, U2895_n1, U2896_n1, U2897_n1, U2898_n1, U2899_n1, U2900_n1,
         U2901_n1, U2902_n1, U3090_n1, U3092_n1, U3094_n1, U3096_n1, U3098_n1,
         U3124_n1, U3171_n1;
  assign g11489 = 1'b0;
  assign g6280 = g100;
  assign g6281 = g101;
  assign g6282 = g102;
  assign g6283 = g103;
  assign g6284 = g104;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6285 = g28;
  assign g6253 = g29;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g8271 = g5816;
  assign g6264 = g82;
  assign g6265 = g83;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6920 = g8561;
  assign g6926 = g8562;
  assign g6932 = g8563;
  assign g6942 = g8564;
  assign g6949 = g8565;
  assign g6955 = g8566;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g5101 = g872;
  assign g8061 = g872;
  assign g5105 = g873;
  assign g8062 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g9961 = g9451;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g8984 = test_so10;

  SDFFX1 DFF_0_Q_reg ( .D(g4556), .SI(test_si1), .SE(n3069), .CLK(n3109), .Q(
        g1289), .QN(n2912) );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(n2954), .CLK(n3145), .Q(
        g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(n2986), .CLK(n3130), .Q(g312), 
        .QN(n2855) );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(n3008), .CLK(n3119), .Q(g452), .QN(n2814) );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(n3011), .CLK(n3117), .Q(g123)
         );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(n2966), .CLK(n3140), .Q(g207)
         );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(n2944), .CLK(n3151), .Q(g713), 
        .QN(n2694) );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(n2944), .CLK(n3151), .Q(g1153), .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(n2943), .CLK(n3151), .Q(
        g1744) );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(n2943), .CLK(n3151), .Q(
        g1558), .QN(n2725) );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(n3004), .CLK(n3120), .Q(
        g695), .QN(n2913) );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(n3004), .CLK(n3121), .Q(
        g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(n3066), .CLK(n3110), .Q(g940), .QN(n1712) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(n3063), .CLK(n3110), .Q(
        g976), .QN(n2880) );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(n2952), .CLK(n3147), .Q(g709) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(n3004), .CLK(n3121), .Q(
        g1092) );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(n2971), .CLK(n3137), .Q(
        g1574), .QN(n2724) );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(n2970), .CLK(n3137), .Q(
        g1864), .QN(n2899) );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(n2970), .CLK(n3137), .Q(
        g369), .QN(n2789) );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(n3003), .CLK(n3121), .Q(
        g1580) );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(n3003), .CLK(n3121), .Q(
        g1736) );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(n3003), .CLK(n3121), .Q(
        n1637) );
  SDFFX1 DFF_23_Q_reg ( .D(n69), .SI(n1637), .SE(n3002), .CLK(n3121), .Q(n3065), .QN(n5222) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(n3002), .CLK(n3121), .Q(
        g1424) );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(n3002), .CLK(n3121), .Q(
        g1737) );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(n2943), .CLK(n3151), .Q(
        g1672) );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(n3028), .CLK(n3114), .Q(
        g1077) );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(n3068), .CLK(n3109), .Q(
        g1231), .QN(n2685) );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(n3049), .CLK(n3112), .Q(g4), 
        .QN(n2757) );
  SDFFX1 DFF_30_Q_reg ( .D(n100), .SI(g4), .SE(n2984), .CLK(n3130), .Q(g4177)
         );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(n2960), .CLK(n3142), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(n3015), .CLK(n3115), .Q(
        g1304) );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(n2978), .CLK(n3134), .Q(
        g243) );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(n3039), .CLK(n3113), .Q(
        g1499), .QN(n2845) );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(n2980), .CLK(n3133), .Q(
        g1444), .QN(n2892) );
  SDFFX1 DFF_37_Q_reg ( .D(n23), .SI(g1444), .SE(n3066), .CLK(n3110), .Q(n3064), .QN(n5214) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(n2984), .CLK(n3131), .Q(
        g4180), .QN(n2920) );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(n2955), .CLK(n3145), .Q(
        g1543), .QN(n2721) );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(n2985), .CLK(n3130), .Q(g315), .QN(n2874) );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(n2999), .CLK(n3123), .Q(
        g1534), .QN(n1632) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(n2999), .CLK(n3123), .Q(
        g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(n3052), .CLK(n3112), .Q(
        g1927), .QN(n2800) );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(n2974), .CLK(n3136), .Q(
        g1660) );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(n2951), .CLK(n3147), .Q(
        g278) );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(n2950), .CLK(n3147), .Q(
        g1436), .QN(n2889) );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(n2950), .CLK(n3147), .Q(
        g718) );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(n2950), .CLK(n3147), .Q(
        g8985), .QN(n1669) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(n2950), .CLK(n3148), .Q(
        g554) );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(n2993), .CLK(n3126), .Q(
        g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(n2992), .CLK(n3126), .Q(
        g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n55), .SI(g981), .SE(n3063), .CLK(n3110), .Q(g3007)
         );
  SDFFX1 DFF_54_Q_reg ( .D(g1713), .SI(g3007), .SE(n2985), .CLK(n3130), .Q(
        test_so1), .QN(n2938) );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(n2989), .CLK(n3128), .Q(
        g829) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(n2944), .CLK(n3150), .Q(
        g1095) );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(n2944), .CLK(n3151), .Q(
        g704), .QN(n2854) );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(n3021), .CLK(n3115), .Q(
        g1265), .QN(n2805) );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(n2965), .CLK(n3140), .Q(
        g1786), .QN(n2904) );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(n3005), .CLK(n3120), .Q(
        g682), .QN(n2784) );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(n3015), .CLK(n3115), .Q(
        g1296) );
  SDFFX1 DFF_62_Q_reg ( .D(g104), .SI(g1296), .SE(n3015), .CLK(n3115), .Q(
        g2602) );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(n2988), .CLK(n3129), .Q(
        g8977), .QN(n1668) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(n2952), .CLK(n3146), .Q(
        n3062), .QN(n5226) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(n2952), .CLK(n3146), .Q(g327), .QN(n2836) );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(n2986), .CLK(n3129), .Q(
        g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(n2966), .CLK(n3139), .Q(
        g1371), .QN(n2847) );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(n2960), .CLK(n3143), .Q(
        g1956) );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(n3001), .CLK(n3122), .Q(
        g1675) );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(n3000), .CLK(n3122), .Q(
        g354) );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(n3000), .CLK(n3122), .Q(g113) );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(n3000), .CLK(n3122), .Q(g639), .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(n3000), .CLK(n3123), .Q(
        g1684) );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(n3000), .CLK(n3123), .Q(
        g1639) );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(n2964), .CLK(n3140), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(n2962), .CLK(n3141), .Q(
        g248), .QN(n1598) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(n2962), .CLK(n3141), .Q(
        g1707), .QN(n2905) );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(n2998), .CLK(n3124), .Q(
        g1759), .QN(n2887) );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(n2998), .CLK(n3124), .Q(
        g351) );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(n2998), .CLK(n3124), .Q(
        g1957) );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(n2997), .CLK(n3124), .Q(
        g1604) );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(n2997), .CLK(n3124), .Q(
        g1098) );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(n2997), .CLK(n3124), .Q(
        g932), .QN(n1591) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(n3060), .CLK(n3111), .Q(
        g1896), .QN(n2785) );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(n3005), .CLK(n3120), .Q(
        g736), .QN(n2866) );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(n2997), .CLK(n3124), .Q(
        g1019), .QN(n2792) );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(n2997), .CLK(n3124), .Q(
        n3061), .QN(n5227) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(n2996), .CLK(n3124), .Q(g745), .QN(n2684) );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(n2996), .CLK(n3124), .Q(
        g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(n2988), .CLK(n3129), .Q(
        g8979), .QN(n1667) );
  SDFFX1 DFF_92_Q_reg ( .D(n2928), .SI(g8979), .SE(n3049), .CLK(n3112), .Q(g32), .QN(n5219) );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(n3049), .CLK(n3112), .Q(n1865), .QN(n2661) );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(n3049), .CLK(n3112), .Q(
        g1086) );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(n3006), .CLK(n3120), .Q(
        g1486), .QN(n2819) );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(n2973), .CLK(n3136), .Q(
        g1730), .QN(n2647) );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(n2973), .CLK(n3136), .Q(
        g1504), .QN(n2702) );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(n2979), .CLK(n3133), .Q(
        g1470) );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(n2979), .CLK(n3133), .Q(
        g822), .QN(n2917) );
  SDFFX1 DFF_100_Q_reg ( .D(g29), .SI(g822), .SE(n2979), .CLK(n3133), .Q(g2609) );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(n2982), .CLK(n3132), .Q(
        g1678) );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(n2982), .CLK(n3132), .Q(
        g174), .QN(n2908) );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(n2976), .CLK(n3135), .Q(
        g1766), .QN(n2897) );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(n2983), .CLK(n3131), .Q(
        g1801), .QN(n2902) );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(n2983), .CLK(n3131), .Q(
        g186), .QN(n2690) );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(n2968), .CLK(n3139), .Q(
        g959), .QN(n2646) );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(n2944), .CLK(n3150), .Q(
        test_so2) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(n2959), .CLK(n3143), 
        .Q(g1407), .QN(n2705) );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(n2994), .CLK(n3126), .Q(
        g1868) );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(n2993), .CLK(n3126), .Q(
        g4173), .QN(n2924) );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(n2974), .CLK(n3135), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(n3009), .CLK(n3118), .Q(
        g396) );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(n2961), .CLK(n3142), .Q(
        g1015), .QN(n2791) );
  SDFFX1 DFF_116_Q_reg ( .D(n91), .SI(g1015), .SE(n2961), .CLK(n3142), .Q(
        n1650), .QN(n5225) );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(n2981), .CLK(n3132), .Q(
        n3059) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(n2980), .CLK(n3132), .Q(
        g1415), .QN(n2700) );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(n3068), .CLK(n3109), .Q(
        g1227), .QN(n2686) );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(n2972), .CLK(n3136), .Q(
        g1721) );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(n2972), .CLK(n3136), .Q(
        n3058), .QN(n5215) );
  SDFFX1 DFF_122_Q_reg ( .D(n2933), .SI(n3058), .SE(n2972), .CLK(n3137), .Q(
        n3057) );
  SDFFX1 DFF_123_Q_reg ( .D(n170), .SI(n3057), .SE(n2972), .CLK(n3137), .Q(
        g284), .QN(n2738) );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(n3066), .CLK(n3110), .Q(
        g426), .QN(n2873) );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(n2966), .CLK(n3139), .Q(
        g219), .QN(n2693) );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(n2961), .CLK(n3142), .Q(
        n3056), .QN(DFF_126_n1) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(n2961), .CLK(n3142), .Q(
        g806), .QN(n2918) );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(n2967), .CLK(n3139), .Q(
        g1428), .QN(n2891) );
  SDFFX1 DFF_129_Q_reg ( .D(g102), .SI(g1428), .SE(n2967), .CLK(n3139), .Q(
        g2605) );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(n2967), .CLK(n3139), .Q(
        g1564) );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(n2967), .CLK(n3139), .Q(
        g1741), .QN(n1633) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(n2967), .CLK(n3139), .Q(
        g225) );
  SDFFX1 DFF_133_Q_reg ( .D(n152), .SI(g225), .SE(n2960), .CLK(n3143), .Q(g281), .QN(n2737) );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(n2959), .CLK(n3143), .Q(
        g1308), .QN(n2660) );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(n2953), .CLK(n3146), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(n2981), .CLK(n3132), .Q(
        n3055), .QN(DFF_136_n1) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(n2981), .CLK(n3132), .Q(
        g1217) );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(n2959), .CLK(n3143), .Q(
        g1589), .QN(n2718) );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(n2979), .CLK(n3133), .Q(
        g1466), .QN(n2823) );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(n2971), .CLK(n3137), .Q(
        g1571), .QN(n2717) );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(n2994), .CLK(n3126), .Q(
        g1861), .QN(n2901) );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(n2994), .CLK(n3126), .Q(
        n3054), .QN(n5228) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(n2980), .CLK(n3132), .Q(
        g1448), .QN(n2825) );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(n2980), .CLK(n3132), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(n3068), .CLK(n3109), .Q(
        g1333), .QN(n2659) );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(n2950), .CLK(n3148), .Q(
        g153), .QN(n2842) );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(n2950), .CLK(n3148), .Q(
        g962) );
  SDFFX1 DFF_149_Q_reg ( .D(n99), .SI(g962), .SE(n2993), .CLK(n3126), .Q(g4175) );
  SDFFX1 DFF_150_Q_reg ( .D(g28), .SI(g4175), .SE(n2993), .CLK(n3126), .Q(
        g2603) );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(n2993), .CLK(n3126), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(n2963), .CLK(n3141), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(n2963), .CLK(n3141), .Q(
        g1397), .QN(n1711) );
  SDFFX1 DFF_154_Q_reg ( .D(g103), .SI(g1397), .SE(n2962), .CLK(n3141), .Q(
        g2606) );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(n3063), .CLK(n3111), .Q(
        g1950), .QN(n2868) );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(n3052), .CLK(n3111), .Q(
        g756) );
  SDFFX1 DFF_157_Q_reg ( .D(g4892), .SI(g756), .SE(n2980), .CLK(n3133), .Q(
        n3053), .QN(DFF_157_n1) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(n2959), .CLK(n3143), .Q(
        g549) );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(n3067), .CLK(n3109), .Q(
        g105) );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(n3067), .CLK(n3109), .Q(
        g1669) );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(n3067), .CLK(n3109), .Q(
        test_so3), .QN(n2846) );
  SDFFX1 DFF_164_Q_reg ( .D(n81), .SI(test_si4), .SE(n2971), .CLK(n3137), .Q(
        g1531), .QN(n1652) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(n3039), .CLK(n3113), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(n2974), .CLK(n3135), .Q(
        g572) );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(n3003), .CLK(n3121), .Q(
        g1011), .QN(n2830) );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(n3003), .CLK(n3121), .Q(
        n3051) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(n3003), .CLK(n3121), .Q(
        g1411), .QN(n2723) );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(n2961), .CLK(n3142), .Q(
        g1074) );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(n3007), .CLK(n3119), .Q(
        g444), .QN(n2812) );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(n2996), .CLK(n3125), .Q(
        g1474) );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(n2985), .CLK(n3130), .Q(
        g1080) );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(n2985), .CLK(n3130), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(n2977), .CLK(n3134), .Q(
        g333), .QN(n2857) );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(n2977), .CLK(n3134), .Q(
        g269), .QN(n2736) );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(n3008), .CLK(n3118), .Q(
        g401), .QN(n2837) );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(n3039), .CLK(n3113), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(n3032), .CLK(n3113), .Q(g9) );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(n3005), .CLK(n3120), .Q(g664), 
        .QN(n2794) );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(n2978), .CLK(n3133), .Q(
        g965) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(n2978), .CLK(n3133), .Q(
        g1400), .QN(n1629) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(n2978), .CLK(n3133), .Q(
        g309), .QN(n2638) );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(n2978), .CLK(n3134), .Q(
        g814), .QN(n2919) );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(n2978), .CLK(n3134), .Q(
        g231), .QN(n2849) );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(n2975), .CLK(n3135), .Q(
        g557) );
  SDFFX1 DFF_187_Q_reg ( .D(g103), .SI(g557), .SE(n2975), .CLK(n3135), .Q(
        g2612) );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(n2974), .CLK(n3135), .Q(
        g869), .QN(n2683) );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(n2965), .CLK(n3140), .Q(
        g1383), .QN(n2689) );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(n2981), .CLK(n3132), .Q(
        g158), .QN(n2822) );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(n2981), .CLK(n3132), .Q(
        g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(n2947), .CLK(n3149), .Q(
        g1023), .QN(n2766) );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(n2947), .CLK(n3149), .Q(
        g259) );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(n2947), .CLK(n3149), .Q(
        n3050), .QN(n5216) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(n2947), .CLK(n3149), .Q(
        g1327) );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(n3014), .CLK(n3116), .Q(
        g654) );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(n2990), .CLK(n3127), .Q(
        g293), .QN(n2735) );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(n2990), .CLK(n3128), .Q(
        g1346), .QN(n2878) );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(n2955), .CLK(n3145), .Q(
        g1633) );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(n2955), .CLK(n3145), .Q(
        g1753) );
  SDFFX1 DFF_201_Q_reg ( .D(n2930), .SI(g1753), .SE(n2955), .CLK(n3145), .Q(
        g1508) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(n3028), .CLK(n3114), .Q(
        g1240), .QN(n2871) );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(n2991), .CLK(n3127), .Q(
        g538) );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(n3008), .CLK(n3119), .Q(
        g416), .QN(n2810) );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(n2991), .CLK(n3127), .Q(
        g542), .QN(n2865) );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(n2974), .CLK(n3136), .Q(
        g1681) );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(n2970), .CLK(n3138), .Q(
        g374) );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(n2969), .CLK(n3138), .Q(
        g563) );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(n2969), .CLK(n3138), .Q(
        g1914) );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(n2991), .CLK(n3127), .Q(
        g530), .QN(n2862) );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(n2991), .CLK(n3127), .Q(
        g575) );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(n2954), .CLK(n3146), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(n2954), .CLK(n3146), .Q(
        g8978), .QN(n1674) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(n2954), .CLK(n3146), .Q(
        test_so4), .QN(n2935) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(n2946), .CLK(n3150), 
        .Q(g1317) );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(n3009), .CLK(n3118), .Q(
        g357) );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(n3009), .CLK(n3118), .Q(
        g386), .QN(n2835) );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(n2956), .CLK(n3145), .Q(
        g1601) );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(n2956), .CLK(n3145), .Q(
        g166), .QN(n2820) );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(n2992), .CLK(n3126), .Q(
        g501) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(n2977), .CLK(n3134), .Q(
        g262) );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(n2977), .CLK(n3134), .Q(
        g1840), .QN(n2867) );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(n2977), .CLK(n3134), .Q(
        g8983), .QN(n1666) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(n2963), .CLK(n3141), .Q(
        g318), .QN(n2834) );
  SDFFX1 DFF_226_Q_reg ( .D(n224), .SI(g318), .SE(n2989), .CLK(n3128), .Q(
        g1356) );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(n2989), .CLK(n3128), .Q(
        g794), .QN(n2915) );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(n2989), .CLK(n3128), .Q(
        n3048), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(n3010), .CLK(n3118), .Q(
        g302) );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(n2961), .CLK(n3142), .Q(
        g342) );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(n3021), .CLK(n3114), .Q(
        g1250) );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(n3021), .CLK(n3114), .Q(
        g1163), .QN(n5213) );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(n2998), .CLK(n3123), .Q(
        n3047), .QN(g5816) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(n3028), .CLK(n3114), .Q(
        g1032), .QN(n2764) );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(n2949), .CLK(n3148), .Q(
        g1432), .QN(n2826) );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(n3039), .CLK(n3113), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(n3002), .CLK(n3122), .Q(
        g363) );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(n3001), .CLK(n3122), .Q(g330), .QN(n2637) );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(n3001), .CLK(n3122), .Q(
        g1157), .QN(n2838) );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(n3001), .CLK(n3122), .Q(
        n3046), .QN(n5229) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(n3001), .CLK(n3122), .Q(
        n3045), .QN(DFF_242_n1) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(n3001), .CLK(n3122), .Q(
        g928), .QN(n1604) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(n2973), .CLK(n3136), .Q(
        g261) );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(n2992), .CLK(n3127), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(n2990), .CLK(n3127), .Q(
        g254) );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(n2984), .CLK(n3131), .Q(
        g4178), .QN(n2921) );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(n2948), .CLK(n3149), .Q(
        g861), .QN(n2642) );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(n2948), .CLK(n3149), .Q(
        g1627), .QN(n2755) );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(n3015), .CLK(n3115), .Q(
        g1292) );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(n2952), .CLK(n3147), .Q(
        g290) );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(n2995), .CLK(n3125), .Q(
        n3044) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(n2984), .CLK(n3130), .Q(
        g4176), .QN(n2922) );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(n3002), .CLK(n3122), .Q(
        g1583), .QN(n2715) );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(n3002), .CLK(n3122), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(n3039), .CLK(n3113), .Q(
        g1561) );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(n2971), .CLK(n3137), .Q(
        g1546), .QN(n2713) );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(n2953), .CLK(n3146), .Q(
        g287) );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(n2953), .CLK(n3146), .Q(
        g560) );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(n2953), .CLK(n3146), .Q(
        g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n2931), .SI(g617), .SE(n2952), .CLK(n3147), .Q(
        n1631) );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(n3068), .CLK(n3109), .Q(
        g336) );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(n2962), .CLK(n3142), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(n2962), .CLK(n3142), .Q(g305), .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(n3032), .CLK(n3114), .Q(
        g345) );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(n3012), .CLK(n3116), .Q(g8), 
        .QN(n2636) );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(n3012), .CLK(n3117), .Q(
        test_so5) );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(n2983), .CLK(n3131), .Q(
        g2648), .QN(n5218) );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(n2986), .CLK(n3130), .Q(
        g255) );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(n3052), .CLK(n3112), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(n3052), .CLK(n3112), .Q(
        g1738), .QN(n1640) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(n3049), .CLK(n3112), .Q(
        g1478), .QN(n2895) );
  SDFFX1 DFF_275_Q_reg ( .D(n497), .SI(g1478), .SE(n3049), .CLK(n3112), .Q(
        n3042), .QN(DFF_275_n1) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(n2962), .CLK(n3142), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(n2968), .CLK(n3139), .Q(
        g1482), .QN(n2824) );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(n2967), .CLK(n3139), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(n2946), .CLK(n3149), .Q(
        g296), .QN(n2731) );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(n2946), .CLK(n3150), .Q(
        g1663) );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(n3004), .CLK(n3120), .Q(
        g700) );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(n2945), .CLK(n3150), .Q(
        g1762), .QN(n2885) );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(n3004), .CLK(n3121), .Q(
        g360) );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(n2986), .CLK(n3129), .Q(
        g192) );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(n3012), .CLK(n3117), .Q(
        g1657) );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(n3011), .CLK(n3117), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(n3011), .CLK(n3117), .Q(
        g8980), .QN(n1673) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(n3011), .CLK(n3117), .Q(
        g566) );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(n3067), .CLK(n3110), .Q(
        n3041), .QN(n5211) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(n3067), .CLK(n3110), .Q(
        g1089) );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(n3066), .CLK(n3110), .Q(
        g2986), .QN(n2662) );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(n2947), .CLK(n3149), .Q(
        g1071) );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(n3066), .CLK(n3110), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(n3066), .CLK(n3110), .Q(
        g971), .QN(n2881) );
  SDFFX1 DFF_295_Q_reg ( .D(g83), .SI(g971), .SE(n3063), .CLK(n3110), .Q(g1955) );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(n3010), .CLK(n3117), .Q(
        g143), .QN(n2843) );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(n2977), .CLK(n3134), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(n2976), .CLK(n3134), .Q(
        g1212), .QN(n2911) );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(n3052), .CLK(n3111), .Q(
        g1918), .QN(n2853) );
  SDFFX1 DFF_301_Q_reg ( .D(n101), .SI(g1918), .SE(n2984), .CLK(n3131), .Q(
        g4179) );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(n2970), .CLK(n3137), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(n2997), .CLK(n3124), .Q(
        g237), .QN(n2850) );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(n2996), .CLK(n3124), .Q(g746), .QN(n2900) );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(n2959), .CLK(n3143), .Q(
        g1462), .QN(n2894) );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(n2958), .CLK(n3143), .Q(
        g178) );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(n2957), .CLK(n3144), .Q(
        g366) );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(n2957), .CLK(n3144), .Q(g837), .QN(n2641) );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(n3013), .CLK(n3116), .Q(
        g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(n3032), .CLK(n3113), .Q(
        g1854) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(n3063), .CLK(n3111), .Q(
        g944), .QN(n2650) );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(n3063), .CLK(n3111), .Q(
        g1941), .QN(n2799) );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(n3011), .CLK(n3117), .Q(
        g170), .QN(n2909) );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(n2996), .CLK(n3125), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(n2999), .CLK(n3123), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(n2999), .CLK(n3123), .Q(
        g953), .QN(n2648) );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(n2999), .CLK(n3123), .Q(
        g1958) );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(n2998), .CLK(n3123), .Q(
        n3040), .QN(n5224) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(n2998), .CLK(n3123), .Q(
        g1765) );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(n2972), .CLK(n3136), .Q(
        g1733) );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(n3015), .CLK(n3115), .Q(
        test_so6) );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(n2975), .CLK(n3135), 
        .Q(g1610) );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(n2964), .CLK(n3140), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(n2964), .CLK(n3141), .Q(
        g1324), .QN(n2653) );
  SDFFX1 DFF_326_Q_reg ( .D(n145), .SI(g1324), .SE(n2964), .CLK(n3141), .Q(
        g1540), .QN(n2712) );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(n2966), .CLK(n3139), .Q(
        n3038), .QN(n5230) );
  SDFFX1 DFF_328_Q_reg ( .D(n2932), .SI(n3038), .SE(n2990), .CLK(n3128), .Q(
        g3069) );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(n2993), .CLK(n3126), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(n2995), .CLK(n3125), .Q(
        n3037), .QN(DFF_330_n1) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(n2966), .CLK(n3140), .Q(
        g213), .QN(n2692) );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(n2965), .CLK(n3140), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(n3060), .CLK(n3111), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(n3028), .CLK(n3114), .Q(
        g1245) );
  SDFFX1 DFF_335_Q_reg ( .D(n9), .SI(g1245), .SE(n3021), .CLK(n3114), .Q(n3036), .QN(n5217) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(n2981), .CLK(n3132), .Q(
        n3035), .QN(DFF_336_n1) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(n3010), .CLK(n3117), .Q(
        g148), .QN(n2844) );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(n2989), .CLK(n3128), .Q(g833), .QN(n2640) );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(n2969), .CLK(n3138), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(n2969), .CLK(n3138), .Q(
        g936), .QN(n1630) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(n2969), .CLK(n3138), .Q(
        g1314) );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(n2969), .CLK(n3138), .Q(
        g849), .QN(n2926) );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(n2968), .CLK(n3138), .Q(
        g1336), .QN(n2879) );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(n2949), .CLK(n3148), .Q(
        g272), .QN(n2730) );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(n2948), .CLK(n3148), .Q(
        g1806), .QN(n2903) );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(n2948), .CLK(n3148), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(n3060), .CLK(n3111), .Q(
        g1887), .QN(n2759) );
  SDFFX1 DFF_350_Q_reg ( .D(n63), .SI(g1887), .SE(n3039), .CLK(n3113), .Q(
        n3034) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(n2948), .CLK(n3149), .Q(
        g968) );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(n2994), .CLK(n3125), .Q(
        n3033), .QN(n5234) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(n2994), .CLK(n3125), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(n2954), .CLK(n3145), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(n3021), .CLK(n3115), .Q(
        g1255), .QN(n2802) );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(n2963), .CLK(n3141), .Q(
        g257) );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(n2963), .CLK(n3141), .Q(
        g874) );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(n3013), .CLK(n3116), .Q(
        g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(n3012), .CLK(n3116), .Q(
        g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(n3012), .CLK(n3116), .Q(
        g636) );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(n3069), .CLK(n3109), .Q(
        g1218), .QN(n2687) );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(n2999), .CLK(n3123), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(n2988), .CLK(n3128), .Q(
        g8986), .QN(n1665) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(n2958), .CLK(n3143), .Q(
        g182), .QN(n2841) );
  SDFFX1 DFF_365_Q_reg ( .D(n319), .SI(g182), .SE(n2957), .CLK(n3144), .Q(g950) );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(n2957), .CLK(n3144), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(n2979), .CLK(n3133), .Q(
        g857) );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(n3007), .CLK(n3119), .Q(
        g448), .QN(n2813) );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(n2976), .CLK(n3134), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(n2976), .CLK(n3134), .Q(
        g1727), .QN(n2667) );
  SDFFX1 DFF_371_Q_reg ( .D(n363), .SI(g1727), .SE(n2976), .CLK(n3135), .Q(
        g1592), .QN(n2711) );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(n2976), .CLK(n3135), .Q(
        g1703), .QN(n2916) );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(n2970), .CLK(n3138), .Q(
        g1932), .QN(n2801) );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(n2970), .CLK(n3138), .Q(
        g1624) );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(n3068), .CLK(n3109), .Q(
        test_so7) );
  SDFFX1 DFF_377_Q_reg ( .D(g101), .SI(test_si8), .SE(n3069), .CLK(n3109), .Q(
        g2601) );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(n3007), .CLK(n3119), .Q(
        g440), .QN(n2811) );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(n2992), .CLK(n3127), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(n2991), .CLK(n3127), .Q(
        g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(n3013), .CLK(n3116), .Q(
        g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(n2947), .CLK(n3149), .Q(
        g139), .QN(n2817) );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(n2946), .CLK(n3149), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(n2946), .CLK(n3149), .Q(
        n3031) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(n2995), .CLK(n3125), .Q(
        n3030), .QN(DFF_385_n1) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(n2958), .CLK(n3143), .Q(
        g263), .QN(n2729) );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(n2958), .CLK(n3144), .Q(
        g818), .QN(n2907) );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(n2958), .CLK(n3144), .Q(
        g1747) );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(n2958), .CLK(n3144), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(n2951), .CLK(n3147), .Q(
        g275) );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(n2951), .CLK(n3147), .Q(
        g1524), .QN(n1649) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(n2951), .CLK(n3147), .Q(
        g1577), .QN(n2710) );
  SDFFX1 DFF_393_Q_reg ( .D(n140), .SI(g1577), .SE(n2987), .CLK(n3129), .Q(
        g810), .QN(n2906) );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(n3009), .CLK(n3118), .Q(
        g391), .QN(n2875) );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(n3014), .CLK(n3116), .Q(
        g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(n2983), .CLK(n3131), .Q(
        g1386), .QN(n2840) );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(n2983), .CLK(n3131), .Q(
        g253) );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(n2982), .CLK(n3131), .Q(
        g875) );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(n2982), .CLK(n3131), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(n2946), .CLK(n3150), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(n3014), .CLK(n3115), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(n3014), .CLK(n3115), .Q(
        g1083) );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(n3014), .CLK(n3116), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(n2979), .CLK(n3133), .Q(
        g1636) );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(n2957), .CLK(n3144), .Q(
        g853), .QN(n2645) );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(n3008), .CLK(n3119), .Q(
        g421), .QN(n2856) );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(n2984), .CLK(n3130), .Q(
        g4174), .QN(n2923) );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(n2987), .CLK(n3129), .Q(
        g956), .QN(n2652) );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(n2987), .CLK(n3129), .Q(
        g378), .QN(n2788) );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(n2964), .CLK(n3140), .Q(
        g1756) );
  SDFFX1 DFF_411_Q_reg ( .D(g29), .SI(g1756), .SE(n2964), .CLK(n3141), .Q(
        g2604) );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(n2960), .CLK(n3142), .Q(
        g841) );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(n3068), .CLK(n3109), .Q(
        g1027), .QN(n2910) );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(n3043), .CLK(n3112), .Q(
        g1003), .QN(n2872) );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(n3043), .CLK(n3112), .Q(
        g1403), .QN(n2827) );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(n3043), .CLK(n3112), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(n2960), .CLK(n3142), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(n2960), .CLK(n3143), .Q(
        g1223), .QN(n2688) );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(n3008), .CLK(n3118), .Q(
        g406), .QN(n2804) );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(n3043), .CLK(n3113), .Q(
        g1811), .QN(n1699) );
  SDFFX1 DFF_421_Q_reg ( .D(n366), .SI(g1811), .SE(n2975), .CLK(n3135), .Q(
        n3029), .QN(n5221) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(n2973), .CLK(n3136), .Q(
        g1654) );
  SDFFX1 DFF_424_Q_reg ( .D(n438), .SI(g1654), .SE(n2986), .CLK(n3129), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(n2949), .CLK(n3148), .Q(
        g1595), .QN(n2709) );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(n3005), .CLK(n3120), .Q(
        g1537) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(n3005), .CLK(n3120), .Q(
        g727), .QN(n2798) );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(n2943), .CLK(n3151), .Q(
        test_so8) );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(n2989), .CLK(n3128), 
        .Q(g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(n2988), .CLK(n3128), .Q(
        g481) );
  SDFFX1 DFF_431_Q_reg ( .D(g3462), .SI(g481), .SE(n2988), .CLK(n3128), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(n2948), .CLK(n3148), .Q(
        g1330), .QN(n2658) );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(n2987), .CLK(n3129), .Q(
        g845), .QN(n2927) );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(n2983), .CLK(n3131), .Q(
        g4181), .QN(n2925) );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(n2959), .CLK(n3143), .Q(
        g1512) );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(n2944), .CLK(n3150), .Q(
        n3027), .QN(n5209) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(n3006), .CLK(n3120), .Q(
        g1490), .QN(n2893) );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(n3006), .CLK(n3120), .Q(
        g1166) );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(n2985), .CLK(n3130), .Q(
        g348) );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(n2963), .CLK(n3141), .Q(
        n3026), .QN(DFF_441_n1) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(n3021), .CLK(n3115), .Q(
        g1260), .QN(n2803) );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(n3011), .CLK(n3117), .Q(
        g260) );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(n2953), .CLK(n3146), .Q(
        g131), .QN(n2816) );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(n3032), .CLK(n3113), .Q(
        n3025) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(n3032), .CLK(n3114), .Q(
        g258) );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(n3032), .CLK(n3114), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(n2965), .CLK(n3140), .Q(
        g1318), .QN(n2655) );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(n2954), .CLK(n3145), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(n3013), .CLK(n3116), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g28), .SI(g677), .SE(n3013), .CLK(n3116), .Q(g2608) );
  SDFFX1 DFF_452_Q_reg ( .D(n39), .SI(g2608), .SE(n3013), .CLK(n3116), .Q(
        n3024), .QN(n5210) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(n2995), .CLK(n3125), .Q(
        g1549), .QN(n2708) );
  SDFFX1 DFF_454_Q_reg ( .D(n342), .SI(g1549), .SE(n2995), .CLK(n3125), .Q(
        g947) );
  SDFFX1 DFF_455_Q_reg ( .D(n248), .SI(g947), .SE(n2995), .CLK(n3125), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(n2949), .CLK(n3148), .Q(
        g1598) );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(n2949), .CLK(n3148), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(n2949), .CLK(n3148), .Q(
        g1321), .QN(n2657) );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(n2992), .CLK(n3126), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(n3010), .CLK(n3117), .Q(
        g546) );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(n3060), .CLK(n3111), .Q(
        g1909), .QN(n2914) );
  SDFFX1 DFF_462_Q_reg ( .D(g83), .SI(g1909), .SE(n3052), .CLK(n3111), .Q(g755) );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(n2951), .CLK(n3147), .Q(
        g1552), .QN(n2706) );
  SDFFX1 DFF_464_Q_reg ( .D(g101), .SI(g1552), .SE(n2951), .CLK(n3147), .Q(
        g2610) );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(n3010), .CLK(n3118), .Q(
        g1687) );
  SDFFX1 DFF_466_Q_reg ( .D(n160), .SI(g1687), .SE(n3010), .CLK(n3118), .Q(
        g1586), .QN(n2704) );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(n3009), .CLK(n3118), .Q(
        g324), .QN(n2832) );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(n3009), .CLK(n3118), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(n2968), .CLK(n3138), .Q(
        g1341), .QN(n2877) );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(n2968), .CLK(n3138), .Q(
        g1710) );
  SDFFX1 DFF_472_Q_reg ( .D(n365), .SI(g1710), .SE(n2968), .CLK(n3139), .Q(
        n3023), .QN(n5220) );
  SDFFX1 DFF_473_Q_reg ( .D(n38), .SI(n3023), .SE(n3067), .CLK(n3110), .Q(
        n3022), .QN(n5231) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(n2990), .CLK(n3127), .Q(
        g135), .QN(n2818) );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(n2945), .CLK(n3150), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g104), .SI(g525), .SE(n2945), .CLK(n3150), .Q(
        g2607) );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(n2945), .CLK(n3150), .Q(
        g1607), .QN(n2703) );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(n2945), .CLK(n3150), .Q(
        g321), .QN(n2876) );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(n2945), .CLK(n3150), .Q(
        g8982), .QN(n1672) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(n3028), .CLK(n3114), .Q(
        g1275), .QN(n2869) );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(n3012), .CLK(n3117), .Q(
        test_so9), .QN(n2937) );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(n2982), .CLK(n3131), 
        .Q(g1615) );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(n2987), .CLK(n3129), .Q(
        g382) );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(n2987), .CLK(n3129), .Q(
        n3020), .QN(n5212) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(n2957), .CLK(n3144), .Q(
        g266), .QN(n2727) );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(n3014), .CLK(n3115), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(n2966), .CLK(n3140), .Q(
        n3019), .QN(n5232) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(n3005), .CLK(n3120), .Q(
        g673), .QN(n2758) );
  SDFFX1 DFF_489_Q_reg ( .D(n275), .SI(g673), .SE(n2994), .CLK(n3125), .Q(
        n3018), .QN(DFF_489_n1) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(n2982), .CLK(n3132), .Q(
        g162), .QN(n2821) );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(n3008), .CLK(n3118), .Q(
        g411), .QN(n2858) );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(n2943), .CLK(n3151), .Q(
        g431) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(n3060), .CLK(n3111), .Q(
        g1905) );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(n2996), .CLK(n3125), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(n2955), .CLK(n3145), .Q(
        g1630), .QN(n2752) );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(n2955), .CLK(n3145), .Q(
        g8976), .QN(n1671) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(n2943), .CLK(n3151), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(n3015), .CLK(n3115), .Q(
        g1300), .QN(n2808) );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(n2986), .CLK(n3130), .Q(
        g339) );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(n2985), .CLK(n3130), .Q(
        g256) );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(n2965), .CLK(n3140), .Q(
        g1750) );
  SDFFX1 DFF_502_Q_reg ( .D(g102), .SI(g1750), .SE(n2965), .CLK(n3140), .Q(
        g2611) );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(n2956), .CLK(n3144), .Q(
        g1440), .QN(n2890) );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(n2956), .CLK(n3144), .Q(
        g1666) );
  SDFFX1 DFF_505_Q_reg ( .D(n148), .SI(g1666), .SE(n2956), .CLK(n3144), .Q(
        g1528), .QN(n1635) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(n2990), .CLK(n3128), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(n367), .SI(g1351), .SE(n2975), .CLK(n3135), .Q(
        n3017), .QN(n5223) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(n2953), .CLK(n3146), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(n3043), .CLK(n3113), .Q(
        g1618) );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(n3028), .CLK(n3114), .Q(
        g1235), .QN(n2829) );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(n2956), .CLK(n3145), .Q(
        g299) );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(n3007), .CLK(n3119), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(n3007), .CLK(n3119), .Q(
        g8981), .QN(n1664) );
  SDFFX1 DFF_514_Q_reg ( .D(n185), .SI(g8981), .SE(n3007), .CLK(n3119), .Q(
        g1555), .QN(n2701) );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(n3006), .CLK(n3119), .Q(
        g995), .QN(n2870) );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(n3006), .CLK(n3119), .Q(
        g1621) );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(n3006), .CLK(n3119), .Q(
        n3016), .QN(n5233) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(n2952), .CLK(n3146), .Q(
        g643) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(n3000), .CLK(n3123), .Q(
        g1494), .QN(n2859) );
  SDFFX1 DFF_520_Q_reg ( .D(n167), .SI(g1494), .SE(n2971), .CLK(n3137), .Q(
        g1567), .QN(n2699) );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(n3004), .CLK(n3120), .Q(
        g691), .QN(n2787) );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(n2991), .CLK(n3127), .Q(
        g534) );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(n2975), .CLK(n3135), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(n2974), .CLK(n3136), .Q(
        g569) );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(n2973), .CLK(n3136), .Q(
        g1160) );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(n2973), .CLK(n3136), .Q(
        g1360) );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(n3043), .CLK(n3113), .Q(g1), .QN(n2670) );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(n2992), .CLK(n3127), .Q(g511), .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(n2972), .CLK(n3137), .Q(
        g1724), .QN(n2665) );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(n2971), .CLK(n3137), .Q(
        g12) );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(n3060), .CLK(n3111), .Q(
        g1878), .QN(n2793) );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(n2988), .CLK(n3129), .Q(
        test_so10), .QN(n2936) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(n2980), .CLK(n3133), .Q(
        g1101), .QN(n1654) );
  AND2X2 Tg1_Trojan1 ( .IN1(n38), .IN2(n39), .Q(Tg1_OUT1) );
  AND2X2 Tg1_Trojan2 ( .IN1(n37), .IN2(n151), .Q(Tg1_OUT2) );
  AND2X2 Tg1_Trojan3 ( .IN1(n2), .IN2(n1858), .Q(Tg1_OUT3) );
  AND2X2 Tg1_Trojan4 ( .IN1(g5556), .IN2(n898), .Q(Tg1_OUT4) );
  AND4X1 Tg1_Trojan1234 ( .IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), 
        .IN4(Tg1_OUT4) );
  NOR2X0 Tg1_Trojan5 ( .IN1(n1391), .IN2(n931), .QN(Tg1_OUT5) );
  NOR2X0 Tg1_Trojan6 ( .IN1(n13), .IN2(n49), .QN(Tg1_OUT6) );
  NOR2X0 Tg1_Trojan7 ( .IN1(n1239), .IN2(n1239), .QN(Tg1_OUT7) );
  NOR2X0 Tg1_Trojan8 ( .IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8) );
  AND4X1 Tg1_Trojan5678 ( .IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), 
        .IN4(Tg1_OUT8) );
  AND2X2 Tg2_Trojan1 ( .IN1(n50), .IN2(n34), .Q(Tg2_OUT1) );
  AND2X2 Tg2_Trojan2 ( .IN1(n34), .IN2(n34), .Q(Tg2_OUT2) );
  AND2X2 Tg2_Trojan3 ( .IN1(n34), .IN2(n34), .Q(Tg2_OUT3) );
  AND2X2 Tg2_Trojan4 ( .IN1(n34), .IN2(n34), .Q(Tg2_OUT4) );
  AND4X1 Tg2_Trojan1234 ( .IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), 
        .IN4(Tg2_OUT4) );
  AND2X2 Tg2_Trojan5 ( .IN1(n147), .IN2(n142), .Q(Tg2_OUT5) );
  AND2X2 Tg2_Trojan6 ( .IN1(n1116), .IN2(n80), .Q(Tg2_OUT6) );
  AND2X2 Tg2_Trojan7 ( .IN1(n82), .IN2(n1107), .Q(Tg2_OUT7) );
  AND2X2 Tg2_Trojan8 ( .IN1(n929), .IN2(n154), .Q(Tg2_OUT8) );
  AND4X1 Tg2_Trojan5678 ( .IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), 
        .IN4(Tg2_OUT8) );
  INVX0 TrojanINVtest_se ( .INP(n3069), .ZN(test_se_NOT) );
  AND2X2 Trojan_Trigger ( .IN1(1'b1), .IN2(test_se_NOT), .Q(Trigger_select) );
  MUX21X2 Trojan_Paylaod ( .IN1(g1200), .IN2(n968), .S(Trigger_select), .Q(
        g4207) );
  INVX0 U2972 ( .INP(g109), .ZN(n2939) );
  INVX0 U2973 ( .INP(g109), .ZN(n2940) );
  INVX0 U2974 ( .INP(g109), .ZN(n2941) );
  INVX0 U2975 ( .INP(g109), .ZN(n2942) );
  NBUFFX2 U2976 ( .INP(n3160), .Z(n3111) );
  NBUFFX2 U2977 ( .INP(n3160), .Z(n3110) );
  NBUFFX2 U2978 ( .INP(n3160), .Z(n3109) );
  NBUFFX2 U2979 ( .INP(n3153), .Z(n3144) );
  NBUFFX2 U2980 ( .INP(n3154), .Z(n3138) );
  NBUFFX2 U2981 ( .INP(n3156), .Z(n3127) );
  NBUFFX2 U2982 ( .INP(n3159), .Z(n3116) );
  NBUFFX2 U2983 ( .INP(n3152), .Z(n3149) );
  NBUFFX2 U2984 ( .INP(n3157), .Z(n3125) );
  NBUFFX2 U2985 ( .INP(n3158), .Z(n3118) );
  NBUFFX2 U2986 ( .INP(n3155), .Z(n3135) );
  NBUFFX2 U2987 ( .INP(n3155), .Z(n3132) );
  NBUFFX2 U2988 ( .INP(n3157), .Z(n3124) );
  NBUFFX2 U2989 ( .INP(n3154), .Z(n3141) );
  NBUFFX2 U2990 ( .INP(n3157), .Z(n3122) );
  NBUFFX2 U2991 ( .INP(n3153), .Z(n3143) );
  NBUFFX2 U2992 ( .INP(n3154), .Z(n3139) );
  NBUFFX2 U2993 ( .INP(n3153), .Z(n3146) );
  NBUFFX2 U2994 ( .INP(n3156), .Z(n3129) );
  NBUFFX2 U2995 ( .INP(n3152), .Z(n3150) );
  NBUFFX2 U2996 ( .INP(n3156), .Z(n3128) );
  NBUFFX2 U2997 ( .INP(n3157), .Z(n3126) );
  NBUFFX2 U2998 ( .INP(n3152), .Z(n3148) );
  NBUFFX2 U2999 ( .INP(n3155), .Z(n3136) );
  NBUFFX2 U3000 ( .INP(n3157), .Z(n3123) );
  NBUFFX2 U3001 ( .INP(n3156), .Z(n3131) );
  NBUFFX2 U3002 ( .INP(n3155), .Z(n3133) );
  NBUFFX2 U3003 ( .INP(n3159), .Z(n3113) );
  NBUFFX2 U3004 ( .INP(n3155), .Z(n3134) );
  NBUFFX2 U3005 ( .INP(n3159), .Z(n3115) );
  NBUFFX2 U3006 ( .INP(n3153), .Z(n3142) );
  NBUFFX2 U3007 ( .INP(n3159), .Z(n3112) );
  NBUFFX2 U3008 ( .INP(n3159), .Z(n3114) );
  NBUFFX2 U3009 ( .INP(n3154), .Z(n3137) );
  NBUFFX2 U3010 ( .INP(n3152), .Z(n3147) );
  NBUFFX2 U3011 ( .INP(n3158), .Z(n3121) );
  NBUFFX2 U3012 ( .INP(n3158), .Z(n3120) );
  NBUFFX2 U3013 ( .INP(n3154), .Z(n3140) );
  NBUFFX2 U3014 ( .INP(n3158), .Z(n3117) );
  NBUFFX2 U3015 ( .INP(n3158), .Z(n3119) );
  NBUFFX2 U3016 ( .INP(n3156), .Z(n3130) );
  NBUFFX2 U3017 ( .INP(n3153), .Z(n3145) );
  NBUFFX2 U3018 ( .INP(n3152), .Z(n3151) );
  NBUFFX2 U3019 ( .INP(n3098), .Z(n2943) );
  NBUFFX2 U3020 ( .INP(n3098), .Z(n2944) );
  NBUFFX2 U3021 ( .INP(n3097), .Z(n2945) );
  NBUFFX2 U3022 ( .INP(n3097), .Z(n2946) );
  NBUFFX2 U3023 ( .INP(n3097), .Z(n2947) );
  NBUFFX2 U3024 ( .INP(n3096), .Z(n2948) );
  NBUFFX2 U3025 ( .INP(n3096), .Z(n2949) );
  NBUFFX2 U3026 ( .INP(n3096), .Z(n2950) );
  NBUFFX2 U3027 ( .INP(n3095), .Z(n2951) );
  NBUFFX2 U3028 ( .INP(n3095), .Z(n2952) );
  NBUFFX2 U3029 ( .INP(n3095), .Z(n2953) );
  NBUFFX2 U3030 ( .INP(n3094), .Z(n2954) );
  NBUFFX2 U3031 ( .INP(n3094), .Z(n2955) );
  NBUFFX2 U3032 ( .INP(n3094), .Z(n2956) );
  NBUFFX2 U3033 ( .INP(n3093), .Z(n2957) );
  NBUFFX2 U3034 ( .INP(n3093), .Z(n2958) );
  NBUFFX2 U3035 ( .INP(n3093), .Z(n2959) );
  NBUFFX2 U3036 ( .INP(n3092), .Z(n2960) );
  NBUFFX2 U3037 ( .INP(n3092), .Z(n2961) );
  NBUFFX2 U3038 ( .INP(n3092), .Z(n2962) );
  NBUFFX2 U3039 ( .INP(n3091), .Z(n2963) );
  NBUFFX2 U3040 ( .INP(n3091), .Z(n2964) );
  NBUFFX2 U3041 ( .INP(n3091), .Z(n2965) );
  NBUFFX2 U3042 ( .INP(n3090), .Z(n2966) );
  NBUFFX2 U3043 ( .INP(n3090), .Z(n2967) );
  NBUFFX2 U3044 ( .INP(n3090), .Z(n2968) );
  NBUFFX2 U3045 ( .INP(n3089), .Z(n2969) );
  NBUFFX2 U3046 ( .INP(n3089), .Z(n2970) );
  NBUFFX2 U3047 ( .INP(n3089), .Z(n2971) );
  NBUFFX2 U3048 ( .INP(n3088), .Z(n2972) );
  NBUFFX2 U3049 ( .INP(n3088), .Z(n2973) );
  NBUFFX2 U3050 ( .INP(n3088), .Z(n2974) );
  NBUFFX2 U3051 ( .INP(n3087), .Z(n2975) );
  NBUFFX2 U3052 ( .INP(n3087), .Z(n2976) );
  NBUFFX2 U3053 ( .INP(n3087), .Z(n2977) );
  NBUFFX2 U3054 ( .INP(n3086), .Z(n2978) );
  NBUFFX2 U3055 ( .INP(n3086), .Z(n2979) );
  NBUFFX2 U3056 ( .INP(n3086), .Z(n2980) );
  NBUFFX2 U3057 ( .INP(n3085), .Z(n2981) );
  NBUFFX2 U3058 ( .INP(n3085), .Z(n2982) );
  NBUFFX2 U3059 ( .INP(n3085), .Z(n2983) );
  NBUFFX2 U3060 ( .INP(n3084), .Z(n2984) );
  NBUFFX2 U3061 ( .INP(n3084), .Z(n2985) );
  NBUFFX2 U3062 ( .INP(n3084), .Z(n2986) );
  NBUFFX2 U3063 ( .INP(n3083), .Z(n2987) );
  NBUFFX2 U3064 ( .INP(n3083), .Z(n2988) );
  NBUFFX2 U3065 ( .INP(n3083), .Z(n2989) );
  NBUFFX2 U3066 ( .INP(n3082), .Z(n2990) );
  NBUFFX2 U3067 ( .INP(n3082), .Z(n2991) );
  NBUFFX2 U3068 ( .INP(n3082), .Z(n2992) );
  NBUFFX2 U3069 ( .INP(n3081), .Z(n2993) );
  NBUFFX2 U3070 ( .INP(n3081), .Z(n2994) );
  NBUFFX2 U3071 ( .INP(n3081), .Z(n2995) );
  NBUFFX2 U3072 ( .INP(n3080), .Z(n2996) );
  NBUFFX2 U3073 ( .INP(n3080), .Z(n2997) );
  NBUFFX2 U3074 ( .INP(n3080), .Z(n2998) );
  NBUFFX2 U3075 ( .INP(n3079), .Z(n2999) );
  NBUFFX2 U3076 ( .INP(n3079), .Z(n3000) );
  NBUFFX2 U3077 ( .INP(n3079), .Z(n3001) );
  NBUFFX2 U3078 ( .INP(n3078), .Z(n3002) );
  NBUFFX2 U3079 ( .INP(n3078), .Z(n3003) );
  NBUFFX2 U3080 ( .INP(n3078), .Z(n3004) );
  NBUFFX2 U3081 ( .INP(n3077), .Z(n3005) );
  NBUFFX2 U3082 ( .INP(n3077), .Z(n3006) );
  NBUFFX2 U3083 ( .INP(n3077), .Z(n3007) );
  NBUFFX2 U3084 ( .INP(n3076), .Z(n3008) );
  NBUFFX2 U3085 ( .INP(n3076), .Z(n3009) );
  NBUFFX2 U3086 ( .INP(n3076), .Z(n3010) );
  NBUFFX2 U3087 ( .INP(n3075), .Z(n3011) );
  NBUFFX2 U3088 ( .INP(n3075), .Z(n3012) );
  NBUFFX2 U3089 ( .INP(n3075), .Z(n3013) );
  NBUFFX2 U3091 ( .INP(n3074), .Z(n3014) );
  NBUFFX2 U3093 ( .INP(n3074), .Z(n3015) );
  NBUFFX2 U3095 ( .INP(n3074), .Z(n3021) );
  NBUFFX2 U3097 ( .INP(n3073), .Z(n3028) );
  NBUFFX2 U3099 ( .INP(n3073), .Z(n3032) );
  NBUFFX2 U3100 ( .INP(n3073), .Z(n3039) );
  NBUFFX2 U3101 ( .INP(n3072), .Z(n3043) );
  NBUFFX2 U3102 ( .INP(n3072), .Z(n3049) );
  NBUFFX2 U3103 ( .INP(n3072), .Z(n3052) );
  NBUFFX2 U3104 ( .INP(n3071), .Z(n3060) );
  NBUFFX2 U3105 ( .INP(n3071), .Z(n3063) );
  NBUFFX2 U3106 ( .INP(n3071), .Z(n3066) );
  NBUFFX2 U3107 ( .INP(n3070), .Z(n3067) );
  NBUFFX2 U3108 ( .INP(n3070), .Z(n3068) );
  NBUFFX2 U3109 ( .INP(n3070), .Z(n3069) );
  NBUFFX2 U3110 ( .INP(n3108), .Z(n3070) );
  NBUFFX2 U3111 ( .INP(n3108), .Z(n3071) );
  NBUFFX2 U3112 ( .INP(n3107), .Z(n3072) );
  NBUFFX2 U3113 ( .INP(n3107), .Z(n3073) );
  NBUFFX2 U3114 ( .INP(n3107), .Z(n3074) );
  NBUFFX2 U3115 ( .INP(n3106), .Z(n3075) );
  NBUFFX2 U3116 ( .INP(n3106), .Z(n3076) );
  NBUFFX2 U3117 ( .INP(n3106), .Z(n3077) );
  NBUFFX2 U3118 ( .INP(n3105), .Z(n3078) );
  NBUFFX2 U3119 ( .INP(n3105), .Z(n3079) );
  NBUFFX2 U3120 ( .INP(n3105), .Z(n3080) );
  NBUFFX2 U3121 ( .INP(n3104), .Z(n3081) );
  NBUFFX2 U3122 ( .INP(n3104), .Z(n3082) );
  NBUFFX2 U3123 ( .INP(n3104), .Z(n3083) );
  NBUFFX2 U3125 ( .INP(n3103), .Z(n3084) );
  NBUFFX2 U3126 ( .INP(n3103), .Z(n3085) );
  NBUFFX2 U3127 ( .INP(n3103), .Z(n3086) );
  NBUFFX2 U3128 ( .INP(n3102), .Z(n3087) );
  NBUFFX2 U3129 ( .INP(n3102), .Z(n3088) );
  NBUFFX2 U3130 ( .INP(n3102), .Z(n3089) );
  NBUFFX2 U3131 ( .INP(n3101), .Z(n3090) );
  NBUFFX2 U3132 ( .INP(n3101), .Z(n3091) );
  NBUFFX2 U3133 ( .INP(n3101), .Z(n3092) );
  NBUFFX2 U3134 ( .INP(n3100), .Z(n3093) );
  NBUFFX2 U3135 ( .INP(n3100), .Z(n3094) );
  NBUFFX2 U3136 ( .INP(n3100), .Z(n3095) );
  NBUFFX2 U3137 ( .INP(n3099), .Z(n3096) );
  NBUFFX2 U3138 ( .INP(n3099), .Z(n3097) );
  NBUFFX2 U3139 ( .INP(n3099), .Z(n3098) );
  NBUFFX2 U3140 ( .INP(test_se), .Z(n3099) );
  NBUFFX2 U3141 ( .INP(n3104), .Z(n3100) );
  NBUFFX2 U3142 ( .INP(n3081), .Z(n3101) );
  NBUFFX2 U3143 ( .INP(n3082), .Z(n3102) );
  NBUFFX2 U3144 ( .INP(n3083), .Z(n3103) );
  NBUFFX2 U3145 ( .INP(test_se), .Z(n3104) );
  NBUFFX2 U3146 ( .INP(test_se), .Z(n3105) );
  NBUFFX2 U3147 ( .INP(n3098), .Z(n3106) );
  NBUFFX2 U3148 ( .INP(test_se), .Z(n3107) );
  NBUFFX2 U3149 ( .INP(n3099), .Z(n3108) );
  NBUFFX2 U3150 ( .INP(CK), .Z(n3152) );
  NBUFFX2 U3151 ( .INP(CK), .Z(n3153) );
  NBUFFX2 U3152 ( .INP(CK), .Z(n3154) );
  NBUFFX2 U3153 ( .INP(CK), .Z(n3155) );
  NBUFFX2 U3154 ( .INP(CK), .Z(n3156) );
  NBUFFX2 U3155 ( .INP(CK), .Z(n3157) );
  NBUFFX2 U3156 ( .INP(CK), .Z(n3158) );
  NBUFFX2 U3157 ( .INP(CK), .Z(n3159) );
  NBUFFX2 U3158 ( .INP(CK), .Z(n3160) );
  NOR2X0 U3160 ( .IN1(n3161), .IN2(n3162), .QN(n99) );
  INVX0 U3161 ( .INP(n3163), .ZN(n3162) );
  NOR2X0 U3162 ( .IN1(n1213), .IN2(n1193), .QN(n3163) );
  NAND2X0 U3163 ( .IN1(n3164), .IN2(n3165), .QN(n962) );
  INVX0 U3164 ( .INP(n3166), .ZN(n3165) );
  NOR2X0 U3165 ( .IN1(n49), .IN2(n1696), .QN(n3166) );
  NAND2X0 U3166 ( .IN1(n3167), .IN2(n1696), .QN(n3164) );
  INVX0 U3167 ( .INP(n3168), .ZN(n3167) );
  NAND2X0 U3168 ( .IN1(n3169), .IN2(n3170), .QN(n917) );
  INVX0 U3169 ( .INP(n3171), .ZN(n3170) );
  NOR2X0 U3170 ( .IN1(n13), .IN2(n1697), .QN(n3171) );
  NAND2X0 U3172 ( .IN1(n3172), .IN2(n1697), .QN(n3169) );
  INVX0 U3173 ( .INP(n3173), .ZN(n3172) );
  INVX0 U3174 ( .INP(n3174), .ZN(n898) );
  NOR2X0 U3175 ( .IN1(n3175), .IN2(n3176), .QN(n838) );
  INVX0 U3176 ( .INP(n3177), .ZN(n81) );
  NOR2X0 U3177 ( .IN1(n3178), .IN2(n3179), .QN(n3177) );
  NOR2X0 U3178 ( .IN1(n3180), .IN2(n1652), .QN(n3179) );
  NOR2X0 U3179 ( .IN1(n3181), .IN2(n2845), .QN(n3178) );
  NOR2X0 U3180 ( .IN1(n5222), .IN2(n364), .QN(n69) );
  INVX0 U3181 ( .INP(n3182), .ZN(n55) );
  INVX0 U3182 ( .INP(n3183), .ZN(n527) );
  NOR2X0 U3183 ( .IN1(n5212), .IN2(n2940), .QN(n438) );
  NOR2X0 U3184 ( .IN1(n5211), .IN2(n3184), .QN(n38) );
  INVX0 U3185 ( .INP(n39), .ZN(n3184) );
  NOR2X0 U3186 ( .IN1(n3185), .IN2(n3186), .QN(n39) );
  INVX0 U3187 ( .INP(g6331), .ZN(n3185) );
  NOR2X0 U3188 ( .IN1(n5223), .IN2(n364), .QN(n367) );
  NOR2X0 U3189 ( .IN1(n5221), .IN2(n364), .QN(n366) );
  NOR2X0 U3190 ( .IN1(n5220), .IN2(n364), .QN(n365) );
  INVX0 U3191 ( .INP(n3187), .ZN(n363) );
  NOR2X0 U3192 ( .IN1(n3188), .IN2(n3189), .QN(n3187) );
  NOR2X0 U3193 ( .IN1(n3180), .IN2(n2711), .QN(n3189) );
  NOR2X0 U3194 ( .IN1(n3181), .IN2(n2827), .QN(n3188) );
  NAND2X0 U3195 ( .IN1(n3190), .IN2(n3191), .QN(n342) );
  NAND2X0 U3196 ( .IN1(n1855), .IN2(g833), .QN(n3191) );
  NAND2X0 U3197 ( .IN1(n3192), .IN2(g947), .QN(n3190) );
  NAND2X0 U3198 ( .IN1(n3193), .IN2(n3194), .QN(n319) );
  NAND2X0 U3199 ( .IN1(n1855), .IN2(g837), .QN(n3194) );
  NAND2X0 U3200 ( .IN1(n3192), .IN2(g950), .QN(n3193) );
  NOR2X0 U3201 ( .IN1(n2942), .IN2(n3195), .QN(n2929) );
  INVX0 U3202 ( .INP(n3196), .ZN(n3195) );
  NAND2X0 U3203 ( .IN1(n3197), .IN2(n5214), .QN(n3196) );
  INVX0 U3204 ( .INP(n3198), .ZN(n275) );
  NOR2X0 U3205 ( .IN1(n3199), .IN2(n3200), .QN(n248) );
  INVX0 U3206 ( .INP(n3201), .ZN(n3200) );
  NOR2X0 U3207 ( .IN1(n3202), .IN2(n3203), .QN(n3201) );
  NOR2X0 U3208 ( .IN1(g1834), .IN2(n806), .QN(n3203) );
  NOR2X0 U3209 ( .IN1(n3204), .IN2(n1655), .QN(n3202) );
  NAND2X0 U3210 ( .IN1(n249), .IN2(n926), .QN(n3204) );
  NAND2X0 U3211 ( .IN1(n2867), .IN2(n3205), .QN(n249) );
  NAND2X0 U3212 ( .IN1(n250), .IN2(n3206), .QN(n3205) );
  INVX0 U3213 ( .INP(n3207), .ZN(n250) );
  INVX0 U3214 ( .INP(n3208), .ZN(n23) );
  INVX0 U3215 ( .INP(n3209), .ZN(n228) );
  NAND2X0 U3216 ( .IN1(n3210), .IN2(g109), .QN(n224) );
  NAND2X0 U3217 ( .IN1(n5217), .IN2(n3211), .QN(n3210) );
  INVX0 U3218 ( .INP(n3212), .ZN(n185) );
  NOR2X0 U3219 ( .IN1(n3213), .IN2(n3214), .QN(n3212) );
  NOR2X0 U3220 ( .IN1(n3180), .IN2(n2701), .QN(n3214) );
  NOR2X0 U3221 ( .IN1(n3181), .IN2(n2823), .QN(n3213) );
  INVX0 U3222 ( .INP(n3215), .ZN(n170) );
  NOR2X0 U3223 ( .IN1(n3216), .IN2(n3217), .QN(n3215) );
  NOR2X0 U3224 ( .IN1(n3218), .IN2(n2738), .QN(n3217) );
  NOR2X0 U3225 ( .IN1(n3219), .IN2(n2909), .QN(n3216) );
  INVX0 U3226 ( .INP(n3220), .ZN(n167) );
  NOR2X0 U3227 ( .IN1(n3221), .IN2(n3222), .QN(n3220) );
  NOR2X0 U3228 ( .IN1(n3180), .IN2(n2699), .QN(n3222) );
  NOR2X0 U3229 ( .IN1(n3181), .IN2(n2700), .QN(n3221) );
  INVX0 U3230 ( .INP(n3223), .ZN(n160) );
  NOR2X0 U3231 ( .IN1(n3224), .IN2(n3225), .QN(n3223) );
  NOR2X0 U3232 ( .IN1(n3180), .IN2(n2704), .QN(n3225) );
  NOR2X0 U3233 ( .IN1(n3181), .IN2(n2705), .QN(n3224) );
  INVX0 U3234 ( .INP(n3226), .ZN(n1588) );
  NOR2X0 U3235 ( .IN1(n3227), .IN2(n3228), .QN(n3226) );
  NAND2X0 U3236 ( .IN1(n3229), .IN2(n3230), .QN(n3227) );
  NAND2X0 U3237 ( .IN1(n3231), .IN2(n3230), .QN(n1587) );
  NAND2X0 U3238 ( .IN1(n3232), .IN2(n3231), .QN(n1586) );
  NOR2X0 U3239 ( .IN1(g46), .IN2(n3233), .QN(n3232) );
  NAND2X0 U3240 ( .IN1(n3234), .IN2(n3235), .QN(n1585) );
  NOR2X0 U3241 ( .IN1(g46), .IN2(g42), .QN(n3235) );
  NOR2X0 U3242 ( .IN1(n3233), .IN2(n3228), .QN(n3234) );
  INVX0 U3243 ( .INP(n3236), .ZN(n1546) );
  INVX0 U3244 ( .INP(n3237), .ZN(n152) );
  NOR2X0 U3245 ( .IN1(n3238), .IN2(n3239), .QN(n3237) );
  NOR2X0 U3246 ( .IN1(n3218), .IN2(n2737), .QN(n3239) );
  NOR2X0 U3247 ( .IN1(n3219), .IN2(n2908), .QN(n3238) );
  INVX0 U3248 ( .INP(n3240), .ZN(n151) );
  INVX0 U3249 ( .INP(n3241), .ZN(n148) );
  NOR2X0 U3250 ( .IN1(n3242), .IN2(n3243), .QN(n3241) );
  NOR2X0 U3251 ( .IN1(n3180), .IN2(n1635), .QN(n3243) );
  NOR2X0 U3252 ( .IN1(n3181), .IN2(n2702), .QN(n3242) );
  INVX0 U3253 ( .INP(n3244), .ZN(n145) );
  NOR2X0 U3254 ( .IN1(n3245), .IN2(n3246), .QN(n3244) );
  NOR2X0 U3255 ( .IN1(n3180), .IN2(n2712), .QN(n3246) );
  NOR2X0 U3256 ( .IN1(n3181), .IN2(n2819), .QN(n3245) );
  NOR2X0 U3257 ( .IN1(n3247), .IN2(n3248), .QN(n140) );
  INVX0 U3258 ( .INP(n3249), .ZN(n3248) );
  NOR2X0 U3259 ( .IN1(n1150), .IN2(n1123), .QN(n3249) );
  INVX0 U3260 ( .INP(n3250), .ZN(n1258) );
  NAND2X0 U3261 ( .IN1(g4173), .IN2(g4174), .QN(n1214) );
  NAND2X0 U3262 ( .IN1(n1193), .IN2(g4176), .QN(n1153) );
  NAND2X0 U3263 ( .IN1(n3251), .IN2(g806), .QN(n1151) );
  NAND2X0 U3264 ( .IN1(n1125), .IN2(g4178), .QN(n1099) );
  NAND2X0 U3265 ( .IN1(n1123), .IN2(g814), .QN(n1097) );
  NOR2X0 U3266 ( .IN1(n3161), .IN2(n3252), .QN(n101) );
  INVX0 U3267 ( .INP(n3253), .ZN(n3252) );
  NOR2X0 U3268 ( .IN1(n1098), .IN2(n1093), .QN(n3253) );
  NOR2X0 U3269 ( .IN1(n3161), .IN2(n3254), .QN(n100) );
  INVX0 U3270 ( .INP(n3255), .ZN(n3254) );
  NOR2X0 U3271 ( .IN1(n1152), .IN2(n1125), .QN(n3255) );
  NOR2X0 U3272 ( .IN1(n3256), .IN2(n3199), .QN(g9721) );
  XOR2X1 U3273 ( .IN1(n3257), .IN2(n1609), .Q(n3256) );
  NAND2X0 U3274 ( .IN1(n3258), .IN2(n3259), .QN(n3257) );
  NAND2X0 U3275 ( .IN1(n3260), .IN2(n3261), .QN(n3259) );
  NOR2X0 U3276 ( .IN1(n804), .IN2(n3262), .QN(n3260) );
  NOR2X0 U3277 ( .IN1(n3263), .IN2(n3264), .QN(n3258) );
  INVX0 U3278 ( .INP(n3265), .ZN(n3263) );
  NAND2X0 U3279 ( .IN1(n3266), .IN2(n3267), .QN(g9451) );
  NOR2X0 U3280 ( .IN1(g31), .IN2(g30), .QN(n3266) );
  NOR2X0 U3281 ( .IN1(n3199), .IN2(n3268), .QN(g9272) );
  NAND2X0 U3282 ( .IN1(n3269), .IN2(n3270), .QN(n3268) );
  NAND2X0 U3283 ( .IN1(n3271), .IN2(g1828), .QN(n3270) );
  NAND2X0 U3284 ( .IN1(n3272), .IN2(n1605), .QN(n3269) );
  NOR2X0 U3285 ( .IN1(n3273), .IN2(n3271), .QN(n3272) );
  NOR2X0 U3286 ( .IN1(n3206), .IN2(n3274), .QN(n3271) );
  NOR2X0 U3287 ( .IN1(n3275), .IN2(n3276), .QN(n3274) );
  INVX0 U3288 ( .INP(n3277), .ZN(n3275) );
  NOR2X0 U3289 ( .IN1(n3278), .IN2(n3279), .QN(n3277) );
  NOR2X0 U3290 ( .IN1(n1605), .IN2(n3280), .QN(n3278) );
  NAND2X0 U3291 ( .IN1(g1814), .IN2(g1822), .QN(n3280) );
  NOR2X0 U3292 ( .IN1(n3199), .IN2(n3281), .QN(g9269) );
  XOR2X1 U3293 ( .IN1(g1822), .IN2(n3282), .Q(n3281) );
  NAND2X0 U3294 ( .IN1(n812), .IN2(n3283), .QN(n3282) );
  NAND2X0 U3295 ( .IN1(n3284), .IN2(n3285), .QN(n3283) );
  NAND2X0 U3296 ( .IN1(n1643), .IN2(n3286), .QN(n3285) );
  NOR2X0 U3297 ( .IN1(n3276), .IN2(n3287), .QN(n3284) );
  NOR2X0 U3298 ( .IN1(n3199), .IN2(n3288), .QN(g9266) );
  XOR2X1 U3299 ( .IN1(n1608), .IN2(n3289), .Q(n3288) );
  NOR2X0 U3300 ( .IN1(n3290), .IN2(n3206), .QN(n3289) );
  INVX0 U3301 ( .INP(n812), .ZN(n3206) );
  NOR2X0 U3302 ( .IN1(n3291), .IN2(n3292), .QN(n3290) );
  NAND2X0 U3303 ( .IN1(n3293), .IN2(n3207), .QN(n3292) );
  NOR2X0 U3304 ( .IN1(n817), .IN2(g1822), .QN(n3291) );
  NOR2X0 U3305 ( .IN1(n3199), .IN2(n3294), .QN(g9150) );
  NAND2X0 U3306 ( .IN1(n3295), .IN2(n3296), .QN(n3294) );
  NAND2X0 U3307 ( .IN1(n3297), .IN2(g605), .QN(n3296) );
  NAND2X0 U3308 ( .IN1(n3298), .IN2(n1593), .QN(n3295) );
  NOR2X0 U3309 ( .IN1(n3297), .IN2(n3299), .QN(n3298) );
  INVX0 U3310 ( .INP(n3300), .ZN(n3297) );
  NAND2X0 U3311 ( .IN1(n804), .IN2(n3301), .QN(n3300) );
  NAND2X0 U3312 ( .IN1(n3302), .IN2(n3303), .QN(n3301) );
  NOR2X0 U3313 ( .IN1(n3304), .IN2(n3305), .QN(n3302) );
  NOR2X0 U3314 ( .IN1(n1644), .IN2(n3306), .QN(n3305) );
  NOR2X0 U3315 ( .IN1(n3307), .IN2(g622), .QN(n3304) );
  NOR2X0 U3316 ( .IN1(n3308), .IN2(n3199), .QN(g9124) );
  XOR2X1 U3317 ( .IN1(g599), .IN2(n836), .Q(n3308) );
  NOR2X0 U3318 ( .IN1(n3309), .IN2(n3199), .QN(g9110) );
  XOR2X1 U3319 ( .IN1(n3310), .IN2(n1607), .Q(n3309) );
  NAND2X0 U3320 ( .IN1(n837), .IN2(n3311), .QN(n3310) );
  NAND2X0 U3321 ( .IN1(n804), .IN2(n3312), .QN(n3311) );
  NAND2X0 U3322 ( .IN1(n3307), .IN2(n3313), .QN(n3312) );
  NAND2X0 U3323 ( .IN1(n3314), .IN2(n3315), .QN(n837) );
  NOR2X0 U3324 ( .IN1(g599), .IN2(n3176), .QN(n3314) );
  NAND2X0 U3325 ( .IN1(n3316), .IN2(n3317), .QN(g8973) );
  NAND2X0 U3326 ( .IN1(n3318), .IN2(n3319), .QN(n3317) );
  XOR2X1 U3327 ( .IN1(n3320), .IN2(n1615), .Q(n3318) );
  NAND2X0 U3328 ( .IN1(n3321), .IN2(n3322), .QN(n3320) );
  NAND2X0 U3329 ( .IN1(n2794), .IN2(n3323), .QN(n3322) );
  NAND2X0 U3330 ( .IN1(n3324), .IN2(n3325), .QN(g8945) );
  NAND2X0 U3331 ( .IN1(n3326), .IN2(n3327), .QN(n3325) );
  XNOR2X1 U3332 ( .IN1(n1697), .IN2(n3328), .Q(n3326) );
  NOR2X0 U3333 ( .IN1(n3329), .IN2(n3330), .QN(n3328) );
  NAND2X0 U3334 ( .IN1(n3331), .IN2(n3332), .QN(n3330) );
  NAND2X0 U3335 ( .IN1(n2868), .IN2(n3333), .QN(n3332) );
  NAND2X0 U3336 ( .IN1(n3334), .IN2(n3335), .QN(n3331) );
  INVX0 U3337 ( .INP(n3336), .ZN(n3334) );
  NAND2X0 U3338 ( .IN1(n13), .IN2(n3173), .QN(n3336) );
  NAND2X0 U3339 ( .IN1(n3337), .IN2(n3338), .QN(n3173) );
  NOR2X0 U3340 ( .IN1(g1936), .IN2(n3339), .QN(n3338) );
  NAND2X0 U3341 ( .IN1(n1675), .IN2(n3340), .QN(n3339) );
  NOR2X0 U3342 ( .IN1(g1909), .IN2(n3341), .QN(n3337) );
  NAND2X0 U3343 ( .IN1(n3342), .IN2(n921), .QN(n13) );
  NOR2X0 U3344 ( .IN1(n1694), .IN2(n3343), .QN(n3342) );
  INVX0 U3345 ( .INP(n3344), .ZN(n3343) );
  NAND2X0 U3346 ( .IN1(n3324), .IN2(n3345), .QN(g8944) );
  NAND2X0 U3347 ( .IN1(n3346), .IN2(n3327), .QN(n3345) );
  XOR2X1 U3348 ( .IN1(n3347), .IN2(n1694), .Q(n3346) );
  NAND2X0 U3349 ( .IN1(n3348), .IN2(n3349), .QN(n3347) );
  NAND2X0 U3350 ( .IN1(n3350), .IN2(n3351), .QN(n3349) );
  NAND2X0 U3351 ( .IN1(n3352), .IN2(n3353), .QN(n3351) );
  INVX0 U3352 ( .INP(n3341), .ZN(n3352) );
  NAND2X0 U3353 ( .IN1(n2800), .IN2(n2853), .QN(n3341) );
  NOR2X0 U3354 ( .IN1(n3354), .IN2(n3355), .QN(n3350) );
  NOR2X0 U3355 ( .IN1(n3333), .IN2(n3356), .QN(n3355) );
  NAND2X0 U3356 ( .IN1(n921), .IN2(n3344), .QN(n3356) );
  NOR2X0 U3357 ( .IN1(n3357), .IN2(n3358), .QN(n3344) );
  NOR2X0 U3358 ( .IN1(n2799), .IN2(n3335), .QN(n3354) );
  NAND2X0 U3359 ( .IN1(n3324), .IN2(n3359), .QN(g8943) );
  NAND2X0 U3360 ( .IN1(n3360), .IN2(n3327), .QN(n3359) );
  XOR2X1 U3361 ( .IN1(g1882), .IN2(n3361), .Q(n3360) );
  NOR2X0 U3362 ( .IN1(n3362), .IN2(n3363), .QN(n3361) );
  NAND2X0 U3363 ( .IN1(n3364), .IN2(n3365), .QN(n3363) );
  NAND2X0 U3364 ( .IN1(n2759), .IN2(n3333), .QN(n3365) );
  NAND2X0 U3365 ( .IN1(n3366), .IN2(n3335), .QN(n3364) );
  NOR2X0 U3366 ( .IN1(n1616), .IN2(n3367), .QN(n3366) );
  NAND2X0 U3367 ( .IN1(n3324), .IN2(n3368), .QN(g8941) );
  NAND2X0 U3368 ( .IN1(n3369), .IN2(n3327), .QN(n3368) );
  XNOR2X1 U3369 ( .IN1(n2800), .IN2(n3370), .Q(n3369) );
  NOR2X0 U3370 ( .IN1(n3371), .IN2(n3329), .QN(n3370) );
  NOR2X0 U3371 ( .IN1(n3372), .IN2(n3373), .QN(n3371) );
  NAND2X0 U3372 ( .IN1(n3374), .IN2(n3375), .QN(n3373) );
  INVX0 U3373 ( .INP(n3376), .ZN(n3375) );
  NOR2X0 U3374 ( .IN1(n3377), .IN2(n3357), .QN(n3376) );
  NAND2X0 U3375 ( .IN1(n3378), .IN2(g1900), .QN(n3357) );
  NOR2X0 U3376 ( .IN1(n2914), .IN2(n2853), .QN(n3378) );
  NAND2X0 U3377 ( .IN1(n3353), .IN2(n2853), .QN(n3374) );
  INVX0 U3378 ( .INP(n3379), .ZN(n3353) );
  NOR2X0 U3379 ( .IN1(n2801), .IN2(n3335), .QN(n3372) );
  NAND2X0 U3380 ( .IN1(n3324), .IN2(n3380), .QN(g8940) );
  NAND2X0 U3381 ( .IN1(n3381), .IN2(n3327), .QN(n3380) );
  XNOR2X1 U3382 ( .IN1(n2853), .IN2(n3382), .Q(n3381) );
  NOR2X0 U3383 ( .IN1(n3383), .IN2(n3329), .QN(n3382) );
  INVX0 U3384 ( .INP(n3348), .ZN(n3329) );
  NOR2X0 U3385 ( .IN1(n3384), .IN2(n3385), .QN(n3383) );
  NAND2X0 U3386 ( .IN1(n3386), .IN2(n3379), .QN(n3385) );
  NAND2X0 U3387 ( .IN1(n3387), .IN2(n3388), .QN(n3379) );
  NOR2X0 U3388 ( .IN1(g1900), .IN2(g1909), .QN(n3387) );
  NAND2X0 U3389 ( .IN1(n3389), .IN2(n3390), .QN(n3386) );
  NOR2X0 U3390 ( .IN1(n2914), .IN2(n1675), .QN(n3389) );
  NOR2X0 U3391 ( .IN1(n1718), .IN2(n3335), .QN(n3384) );
  NAND2X0 U3392 ( .IN1(n3324), .IN2(n3391), .QN(g8939) );
  NAND2X0 U3393 ( .IN1(n3392), .IN2(n3327), .QN(n3391) );
  XOR2X1 U3394 ( .IN1(n3393), .IN2(n2914), .Q(n3392) );
  NAND2X0 U3395 ( .IN1(n3394), .IN2(n3348), .QN(n3393) );
  NAND2X0 U3396 ( .IN1(n3395), .IN2(n3396), .QN(n3394) );
  NAND2X0 U3397 ( .IN1(n3333), .IN2(g1914), .QN(n3396) );
  NOR2X0 U3398 ( .IN1(n3397), .IN2(n3398), .QN(n3395) );
  NOR2X0 U3399 ( .IN1(g1900), .IN2(n3399), .QN(n3398) );
  NOR2X0 U3400 ( .IN1(n1675), .IN2(n3377), .QN(n3397) );
  NAND2X0 U3401 ( .IN1(n3324), .IN2(n3400), .QN(g8938) );
  NAND2X0 U3402 ( .IN1(n3401), .IN2(n3327), .QN(n3400) );
  XOR2X1 U3403 ( .IN1(n3402), .IN2(n1675), .Q(n3401) );
  NAND2X0 U3404 ( .IN1(n3403), .IN2(n3348), .QN(n3402) );
  NAND2X0 U3405 ( .IN1(n3404), .IN2(n3405), .QN(n3403) );
  NAND2X0 U3406 ( .IN1(n3333), .IN2(g1905), .QN(n3405) );
  NOR2X0 U3407 ( .IN1(n3390), .IN2(n3388), .QN(n3404) );
  INVX0 U3408 ( .INP(n3399), .ZN(n3388) );
  NAND2X0 U3409 ( .IN1(n3335), .IN2(n3340), .QN(n3399) );
  NOR2X0 U3410 ( .IN1(n3406), .IN2(n3407), .QN(n3340) );
  NAND2X0 U3411 ( .IN1(n3408), .IN2(n1616), .QN(n3407) );
  NAND2X0 U3412 ( .IN1(n1657), .IN2(n1663), .QN(n3406) );
  INVX0 U3413 ( .INP(n3377), .ZN(n3390) );
  NAND2X0 U3414 ( .IN1(n3409), .IN2(n3335), .QN(n3377) );
  NOR2X0 U3415 ( .IN1(n1657), .IN2(n3358), .QN(n3409) );
  NAND2X0 U3416 ( .IN1(n3410), .IN2(n3367), .QN(n3358) );
  NOR2X0 U3417 ( .IN1(n1663), .IN2(n1616), .QN(n3410) );
  NAND2X0 U3418 ( .IN1(n3324), .IN2(n3411), .QN(g8937) );
  NAND2X0 U3419 ( .IN1(n3412), .IN2(n3327), .QN(n3411) );
  XNOR2X1 U3420 ( .IN1(n1657), .IN2(n3413), .Q(n3412) );
  NOR2X0 U3421 ( .IN1(n3362), .IN2(n3414), .QN(n3413) );
  NAND2X0 U3422 ( .IN1(n3415), .IN2(n3416), .QN(n3414) );
  NAND2X0 U3423 ( .IN1(n2785), .IN2(n3333), .QN(n3416) );
  NAND2X0 U3424 ( .IN1(n3417), .IN2(n3335), .QN(n3415) );
  NAND2X0 U3425 ( .IN1(n3418), .IN2(n3419), .QN(n3417) );
  NAND2X0 U3426 ( .IN1(n1663), .IN2(g1872), .QN(n3419) );
  NAND2X0 U3427 ( .IN1(n3408), .IN2(g1882), .QN(n3418) );
  NAND2X0 U3428 ( .IN1(n3348), .IN2(n3420), .QN(n3362) );
  NAND2X0 U3429 ( .IN1(n3421), .IN2(n3335), .QN(n3420) );
  NOR2X0 U3430 ( .IN1(n3408), .IN2(g1872), .QN(n3421) );
  INVX0 U3431 ( .INP(n3367), .ZN(n3408) );
  NAND2X0 U3432 ( .IN1(n3422), .IN2(n3423), .QN(n3367) );
  NAND2X0 U3433 ( .IN1(n1643), .IN2(g1814), .QN(n3423) );
  NOR2X0 U3434 ( .IN1(n3276), .IN2(n3279), .QN(n3422) );
  NOR2X0 U3435 ( .IN1(g1828), .IN2(n3293), .QN(n3279) );
  NAND2X0 U3436 ( .IN1(n3316), .IN2(n3424), .QN(g8926) );
  NAND2X0 U3437 ( .IN1(n3425), .IN2(n3319), .QN(n3424) );
  XOR2X1 U3438 ( .IN1(n1696), .IN2(n3174), .Q(n3425) );
  NAND2X0 U3439 ( .IN1(n3426), .IN2(n3321), .QN(n3174) );
  NOR2X0 U3440 ( .IN1(n3427), .IN2(n3428), .QN(n3426) );
  NOR2X0 U3441 ( .IN1(n3323), .IN2(n3429), .QN(n3428) );
  NAND2X0 U3442 ( .IN1(n3168), .IN2(n49), .QN(n3429) );
  NAND2X0 U3443 ( .IN1(n3430), .IN2(n967), .QN(n49) );
  INVX0 U3444 ( .INP(n3431), .ZN(n3430) );
  NAND2X0 U3445 ( .IN1(g722), .IN2(n3432), .QN(n3431) );
  NAND2X0 U3446 ( .IN1(n3433), .IN2(n3434), .QN(n3168) );
  NOR2X0 U3447 ( .IN1(g722), .IN2(n3435), .QN(n3434) );
  NAND2X0 U3448 ( .IN1(n1676), .IN2(n3436), .QN(n3435) );
  NOR2X0 U3449 ( .IN1(g695), .IN2(n3437), .QN(n3433) );
  NOR2X0 U3450 ( .IN1(n3438), .IN2(g736), .QN(n3427) );
  NAND2X0 U3451 ( .IN1(n3316), .IN2(n3439), .QN(g8923) );
  NAND2X0 U3452 ( .IN1(n3440), .IN2(n3319), .QN(n3439) );
  XOR2X1 U3453 ( .IN1(n3441), .IN2(n1693), .Q(n3440) );
  NAND2X0 U3454 ( .IN1(n3321), .IN2(n3442), .QN(n3441) );
  NAND2X0 U3455 ( .IN1(n3443), .IN2(n3444), .QN(n3442) );
  NAND2X0 U3456 ( .IN1(n3445), .IN2(n3446), .QN(n3444) );
  INVX0 U3457 ( .INP(n3437), .ZN(n3445) );
  NAND2X0 U3458 ( .IN1(n2694), .IN2(n2854), .QN(n3437) );
  NOR2X0 U3459 ( .IN1(n3447), .IN2(n3448), .QN(n3443) );
  NOR2X0 U3460 ( .IN1(n3323), .IN2(n3449), .QN(n3448) );
  NAND2X0 U3461 ( .IN1(n967), .IN2(n3432), .QN(n3449) );
  NOR2X0 U3462 ( .IN1(n3450), .IN2(n3451), .QN(n3432) );
  NOR2X0 U3463 ( .IN1(n2798), .IN2(n3438), .QN(n3447) );
  NAND2X0 U3464 ( .IN1(n3316), .IN2(n3452), .QN(g8922) );
  NAND2X0 U3465 ( .IN1(n3453), .IN2(n3319), .QN(n3452) );
  XOR2X1 U3466 ( .IN1(g668), .IN2(n3454), .Q(n3453) );
  NOR2X0 U3467 ( .IN1(n3455), .IN2(n3456), .QN(n3454) );
  NAND2X0 U3468 ( .IN1(n3457), .IN2(n3458), .QN(n3456) );
  NAND2X0 U3469 ( .IN1(n2758), .IN2(n3323), .QN(n3458) );
  NAND2X0 U3470 ( .IN1(n3459), .IN2(n3438), .QN(n3457) );
  NOR2X0 U3471 ( .IN1(n1615), .IN2(n3460), .QN(n3459) );
  NAND2X0 U3472 ( .IN1(n3324), .IN2(n3461), .QN(g8921) );
  NAND2X0 U3473 ( .IN1(n3462), .IN2(n3327), .QN(n3461) );
  XOR2X1 U3474 ( .IN1(n3463), .IN2(n1616), .Q(n3462) );
  NAND2X0 U3475 ( .IN1(n3348), .IN2(n3464), .QN(n3463) );
  NAND2X0 U3476 ( .IN1(n2793), .IN2(n3333), .QN(n3464) );
  INVX0 U3477 ( .INP(n3335), .ZN(n3333) );
  NAND2X0 U3478 ( .IN1(n3335), .IN2(n918), .QN(n3348) );
  NAND2X0 U3479 ( .IN1(n3465), .IN2(n926), .QN(n918) );
  NAND2X0 U3480 ( .IN1(n3466), .IN2(n3207), .QN(n3465) );
  NAND2X0 U3481 ( .IN1(n3467), .IN2(n2867), .QN(n3207) );
  NOR2X0 U3482 ( .IN1(n1655), .IN2(n1608), .QN(n3467) );
  NAND2X0 U3483 ( .IN1(g1857), .IN2(n3468), .QN(n3466) );
  NAND2X0 U3484 ( .IN1(n1643), .IN2(n1605), .QN(n3468) );
  NOR2X0 U3485 ( .IN1(n3469), .IN2(n929), .QN(n3335) );
  NAND2X0 U3486 ( .IN1(n3470), .IN2(n3471), .QN(n3324) );
  NOR2X0 U3487 ( .IN1(n3327), .IN2(n3276), .QN(n3471) );
  INVX0 U3488 ( .INP(n3472), .ZN(n3276) );
  NOR2X0 U3489 ( .IN1(n3273), .IN2(n812), .QN(n3327) );
  NOR2X0 U3490 ( .IN1(n3273), .IN2(n3473), .QN(n3470) );
  INVX0 U3491 ( .INP(n916), .ZN(n3473) );
  NAND2X0 U3492 ( .IN1(n3316), .IN2(n3474), .QN(g8920) );
  NAND2X0 U3493 ( .IN1(n3475), .IN2(n3319), .QN(n3474) );
  XOR2X1 U3494 ( .IN1(n2694), .IN2(n931), .Q(n3475) );
  NAND2X0 U3495 ( .IN1(n3321), .IN2(n3476), .QN(n931) );
  NAND2X0 U3496 ( .IN1(n3477), .IN2(n3478), .QN(n3476) );
  NAND2X0 U3497 ( .IN1(n3323), .IN2(g718), .QN(n3478) );
  NOR2X0 U3498 ( .IN1(n3479), .IN2(n3480), .QN(n3477) );
  INVX0 U3499 ( .INP(n3481), .ZN(n3480) );
  NAND2X0 U3500 ( .IN1(n2854), .IN2(n3446), .QN(n3481) );
  NOR2X0 U3501 ( .IN1(n3450), .IN2(n3482), .QN(n3479) );
  NAND2X0 U3502 ( .IN1(n3483), .IN2(g686), .QN(n3450) );
  NOR2X0 U3503 ( .IN1(n2913), .IN2(n2854), .QN(n3483) );
  NAND2X0 U3504 ( .IN1(n3316), .IN2(n3484), .QN(g8889) );
  NAND2X0 U3505 ( .IN1(n3485), .IN2(n3319), .QN(n3484) );
  XNOR2X1 U3506 ( .IN1(n50), .IN2(n2854), .Q(n3485) );
  NOR2X0 U3507 ( .IN1(n3486), .IN2(n3487), .QN(n50) );
  INVX0 U3508 ( .INP(n3488), .ZN(n3486) );
  NAND2X0 U3509 ( .IN1(n3489), .IN2(n3490), .QN(n3488) );
  NAND2X0 U3510 ( .IN1(n3323), .IN2(g709), .QN(n3490) );
  NOR2X0 U3511 ( .IN1(n3446), .IN2(n3491), .QN(n3489) );
  NOR2X0 U3512 ( .IN1(n3482), .IN2(n3492), .QN(n3491) );
  NAND2X0 U3513 ( .IN1(g686), .IN2(g695), .QN(n3492) );
  NOR2X0 U3514 ( .IN1(n3493), .IN2(n3494), .QN(n3446) );
  NAND2X0 U3515 ( .IN1(n1676), .IN2(n2913), .QN(n3493) );
  NAND2X0 U3516 ( .IN1(n3316), .IN2(n3495), .QN(g8887) );
  NAND2X0 U3517 ( .IN1(n3496), .IN2(n3319), .QN(n3495) );
  XOR2X1 U3518 ( .IN1(n3497), .IN2(n2913), .Q(n3496) );
  NAND2X0 U3519 ( .IN1(n3498), .IN2(n3321), .QN(n3497) );
  NAND2X0 U3520 ( .IN1(n3499), .IN2(n3500), .QN(n3498) );
  NAND2X0 U3521 ( .IN1(n3323), .IN2(g700), .QN(n3500) );
  NOR2X0 U3522 ( .IN1(n3501), .IN2(n3502), .QN(n3499) );
  NOR2X0 U3523 ( .IN1(g686), .IN2(n3494), .QN(n3502) );
  NOR2X0 U3524 ( .IN1(n1676), .IN2(n3482), .QN(n3501) );
  NAND2X0 U3525 ( .IN1(n3316), .IN2(n3503), .QN(g8885) );
  NAND2X0 U3526 ( .IN1(n3504), .IN2(n3319), .QN(n3503) );
  XOR2X1 U3527 ( .IN1(g686), .IN2(n3505), .Q(n3504) );
  NOR2X0 U3528 ( .IN1(n3487), .IN2(n3506), .QN(n3505) );
  NOR2X0 U3529 ( .IN1(n3507), .IN2(n3508), .QN(n3506) );
  NAND2X0 U3530 ( .IN1(n3494), .IN2(n3482), .QN(n3508) );
  NAND2X0 U3531 ( .IN1(n3509), .IN2(n3438), .QN(n3482) );
  NOR2X0 U3532 ( .IN1(n1656), .IN2(n3451), .QN(n3509) );
  NAND2X0 U3533 ( .IN1(n3510), .IN2(n3460), .QN(n3451) );
  NOR2X0 U3534 ( .IN1(n1662), .IN2(n1615), .QN(n3510) );
  NAND2X0 U3535 ( .IN1(n3438), .IN2(n3436), .QN(n3494) );
  NOR2X0 U3536 ( .IN1(n3511), .IN2(n3512), .QN(n3436) );
  NAND2X0 U3537 ( .IN1(n3513), .IN2(n1615), .QN(n3512) );
  NAND2X0 U3538 ( .IN1(n1656), .IN2(n1662), .QN(n3511) );
  NOR2X0 U3539 ( .IN1(n2787), .IN2(n3438), .QN(n3507) );
  INVX0 U3540 ( .INP(n3321), .ZN(n3487) );
  NAND2X0 U3541 ( .IN1(n3316), .IN2(n3514), .QN(g8883) );
  NAND2X0 U3542 ( .IN1(n3515), .IN2(n3319), .QN(n3514) );
  XNOR2X1 U3543 ( .IN1(n1656), .IN2(n3516), .Q(n3515) );
  NOR2X0 U3544 ( .IN1(n3455), .IN2(n3517), .QN(n3516) );
  NAND2X0 U3545 ( .IN1(n3518), .IN2(n3519), .QN(n3517) );
  NAND2X0 U3546 ( .IN1(n2784), .IN2(n3323), .QN(n3519) );
  INVX0 U3547 ( .INP(n3438), .ZN(n3323) );
  NAND2X0 U3548 ( .IN1(n3520), .IN2(n3438), .QN(n3518) );
  NAND2X0 U3549 ( .IN1(n3521), .IN2(n3522), .QN(n3520) );
  NAND2X0 U3550 ( .IN1(n1662), .IN2(g658), .QN(n3522) );
  NAND2X0 U3551 ( .IN1(n3513), .IN2(g668), .QN(n3521) );
  NAND2X0 U3552 ( .IN1(n3321), .IN2(n3523), .QN(n3455) );
  NAND2X0 U3553 ( .IN1(n3524), .IN2(n3438), .QN(n3523) );
  NOR2X0 U3554 ( .IN1(n3513), .IN2(g658), .QN(n3524) );
  INVX0 U3555 ( .INP(n3460), .ZN(n3513) );
  NAND2X0 U3556 ( .IN1(n3303), .IN2(n3525), .QN(n3460) );
  NAND2X0 U3557 ( .IN1(n1644), .IN2(g591), .QN(n3525) );
  NOR2X0 U3558 ( .IN1(n3526), .IN2(n3527), .QN(n3303) );
  NOR2X0 U3559 ( .IN1(g605), .IN2(n3313), .QN(n3527) );
  NAND2X0 U3560 ( .IN1(n3438), .IN2(n958), .QN(n3321) );
  NAND2X0 U3561 ( .IN1(n3528), .IN2(n3529), .QN(n958) );
  NAND2X0 U3562 ( .IN1(n3530), .IN2(n3307), .QN(n3529) );
  NAND2X0 U3563 ( .IN1(g639), .IN2(n3531), .QN(n3530) );
  NAND2X0 U3564 ( .IN1(n1644), .IN2(n1593), .QN(n3531) );
  NOR2X0 U3565 ( .IN1(n3264), .IN2(n3532), .QN(n3438) );
  NAND2X0 U3566 ( .IN1(n3533), .IN2(n3534), .QN(n3316) );
  NOR2X0 U3567 ( .IN1(n3319), .IN2(n3261), .QN(n3534) );
  INVX0 U3568 ( .INP(n3307), .ZN(n3261) );
  INVX0 U3569 ( .INP(n3535), .ZN(n3319) );
  NOR2X0 U3570 ( .IN1(n3299), .IN2(n3536), .QN(n3533) );
  NAND2X0 U3571 ( .IN1(n3265), .IN2(n3537), .QN(g8820) );
  NAND2X0 U3572 ( .IN1(n3538), .IN2(g622), .QN(n3537) );
  NAND2X0 U3573 ( .IN1(n3535), .IN2(n3539), .QN(n3538) );
  NAND2X0 U3574 ( .IN1(n3540), .IN2(n3307), .QN(n3539) );
  NAND2X0 U3575 ( .IN1(n3540), .IN2(n3176), .QN(n3535) );
  NAND2X0 U3576 ( .IN1(n3541), .IN2(n1713), .QN(n3265) );
  NOR2X0 U3577 ( .IN1(n3176), .IN2(n3307), .QN(n3541) );
  NAND2X0 U3578 ( .IN1(n3542), .IN2(n1645), .QN(n3307) );
  NOR2X0 U3579 ( .IN1(n1609), .IN2(n1607), .QN(n3542) );
  INVX0 U3580 ( .INP(n804), .ZN(n3176) );
  NAND2X0 U3581 ( .IN1(n3543), .IN2(n3544), .QN(g8779) );
  NAND2X0 U3582 ( .IN1(n968), .IN2(g1636), .QN(n3544) );
  NAND2X0 U3583 ( .IN1(n3545), .IN2(n3546), .QN(n3543) );
  NAND2X0 U3584 ( .IN1(n3547), .IN2(n3548), .QN(g8777) );
  NAND2X0 U3585 ( .IN1(n968), .IN2(g1633), .QN(n3548) );
  NAND2X0 U3586 ( .IN1(n3549), .IN2(n3546), .QN(n3547) );
  NAND2X0 U3587 ( .IN1(n3550), .IN2(n3551), .QN(g8776) );
  NAND2X0 U3588 ( .IN1(n968), .IN2(g1630), .QN(n3551) );
  NAND2X0 U3589 ( .IN1(n3552), .IN2(n3546), .QN(n3550) );
  NOR2X0 U3590 ( .IN1(n2939), .IN2(n3553), .QN(g8775) );
  XOR2X1 U3591 ( .IN1(n3554), .IN2(n2889), .Q(n3553) );
  NAND2X0 U3592 ( .IN1(n3555), .IN2(n3556), .QN(g8774) );
  NAND2X0 U3593 ( .IN1(n968), .IN2(g1627), .QN(n3556) );
  NAND2X0 U3594 ( .IN1(n3554), .IN2(n3546), .QN(n3555) );
  NAND2X0 U3595 ( .IN1(n3557), .IN2(n3558), .QN(n3554) );
  NOR2X0 U3596 ( .IN1(n3559), .IN2(n3560), .QN(n3557) );
  NOR2X0 U3597 ( .IN1(g1133), .IN2(n3561), .QN(n3560) );
  NAND2X0 U3598 ( .IN1(n3562), .IN2(n3563), .QN(n3561) );
  NOR2X0 U3599 ( .IN1(n1706), .IN2(n3564), .QN(n3559) );
  NAND2X0 U3600 ( .IN1(n3565), .IN2(n3199), .QN(n3564) );
  NAND2X0 U3601 ( .IN1(n3562), .IN2(n3566), .QN(n3565) );
  NOR2X0 U3602 ( .IN1(n1614), .IN2(g1101), .QN(n3562) );
  NAND2X0 U3603 ( .IN1(n3567), .IN2(n3568), .QN(g8773) );
  NAND2X0 U3604 ( .IN1(n968), .IN2(g1624), .QN(n3568) );
  NAND2X0 U3605 ( .IN1(n3569), .IN2(n3546), .QN(n3567) );
  NOR2X0 U3606 ( .IN1(n2940), .IN2(n3570), .QN(g8772) );
  XOR2X1 U3607 ( .IN1(n3552), .IN2(n2890), .Q(n3570) );
  NAND2X0 U3608 ( .IN1(n3571), .IN2(n3572), .QN(n3552) );
  NOR2X0 U3609 ( .IN1(n3573), .IN2(n3574), .QN(n3571) );
  NOR2X0 U3610 ( .IN1(g1137), .IN2(n3575), .QN(n3574) );
  NAND2X0 U3611 ( .IN1(n3576), .IN2(n3563), .QN(n3575) );
  NOR2X0 U3612 ( .IN1(n1597), .IN2(n3577), .QN(n3573) );
  NAND2X0 U3613 ( .IN1(n3578), .IN2(n3199), .QN(n3577) );
  NAND2X0 U3614 ( .IN1(n3576), .IN2(n3566), .QN(n3578) );
  NOR2X0 U3615 ( .IN1(n1654), .IN2(n1614), .QN(n3576) );
  NAND2X0 U3616 ( .IN1(n3579), .IN2(n3580), .QN(g8771) );
  NAND2X0 U3617 ( .IN1(n968), .IN2(g1621), .QN(n3580) );
  NAND2X0 U3618 ( .IN1(n3581), .IN2(n3546), .QN(n3579) );
  NAND2X0 U3619 ( .IN1(n3582), .IN2(n3583), .QN(g8770) );
  NAND2X0 U3620 ( .IN1(n968), .IN2(g1615), .QN(n3583) );
  NAND2X0 U3621 ( .IN1(n3584), .IN2(n3546), .QN(n3582) );
  NOR2X0 U3622 ( .IN1(n2941), .IN2(n3585), .QN(g8769) );
  XOR2X1 U3623 ( .IN1(n3584), .IN2(n2891), .Q(n3585) );
  NAND2X0 U3624 ( .IN1(n3586), .IN2(n3587), .QN(n3584) );
  NOR2X0 U3625 ( .IN1(n3588), .IN2(n3589), .QN(n3586) );
  NOR2X0 U3626 ( .IN1(g1121), .IN2(n3590), .QN(n3589) );
  NAND2X0 U3627 ( .IN1(n3563), .IN2(n3591), .QN(n3590) );
  NOR2X0 U3628 ( .IN1(n3592), .IN2(g18), .QN(n3563) );
  NOR2X0 U3629 ( .IN1(n1618), .IN2(n3593), .QN(n3588) );
  NAND2X0 U3630 ( .IN1(n3594), .IN2(n3199), .QN(n3593) );
  NAND2X0 U3631 ( .IN1(n3566), .IN2(n3591), .QN(n3594) );
  INVX0 U3632 ( .INP(n3592), .ZN(n3566) );
  NOR2X0 U3633 ( .IN1(n2942), .IN2(n3595), .QN(g8768) );
  XOR2X1 U3634 ( .IN1(n3549), .IN2(n2892), .Q(n3595) );
  NAND2X0 U3635 ( .IN1(n3596), .IN2(n3597), .QN(n3549) );
  NAND2X0 U3636 ( .IN1(n3598), .IN2(n3199), .QN(n3596) );
  XOR2X1 U3637 ( .IN1(n3599), .IN2(n1660), .Q(n3598) );
  NAND2X0 U3638 ( .IN1(n3600), .IN2(n1658), .QN(n3599) );
  NOR2X0 U3639 ( .IN1(n2939), .IN2(n3601), .QN(g8767) );
  XOR2X1 U3640 ( .IN1(n3581), .IN2(n2827), .Q(n3601) );
  NAND2X0 U3641 ( .IN1(n3602), .IN2(n3603), .QN(n3581) );
  NAND2X0 U3642 ( .IN1(n3604), .IN2(n3199), .QN(n3603) );
  XOR2X1 U3643 ( .IN1(n3605), .IN2(n1708), .Q(n3604) );
  NAND2X0 U3644 ( .IN1(n3606), .IN2(n1654), .QN(n3605) );
  NOR2X0 U3645 ( .IN1(n2940), .IN2(n3607), .QN(g8766) );
  XOR2X1 U3646 ( .IN1(n3545), .IN2(n2825), .Q(n3607) );
  NAND2X0 U3647 ( .IN1(n3608), .IN2(n3609), .QN(n3545) );
  NAND2X0 U3648 ( .IN1(n3610), .IN2(n3199), .QN(n3608) );
  XOR2X1 U3649 ( .IN1(n3611), .IN2(n1617), .Q(n3610) );
  NAND2X0 U3650 ( .IN1(n3612), .IN2(g1110), .QN(n3611) );
  NOR2X0 U3651 ( .IN1(n2941), .IN2(n3613), .QN(g8765) );
  XOR2X1 U3652 ( .IN1(n3569), .IN2(n2826), .Q(n3613) );
  NAND2X0 U3653 ( .IN1(n3614), .IN2(n3615), .QN(n3569) );
  NAND2X0 U3654 ( .IN1(n3616), .IN2(n3199), .QN(n3615) );
  XOR2X1 U3655 ( .IN1(n3617), .IN2(n1705), .Q(n3616) );
  NAND2X0 U3656 ( .IN1(n3606), .IN2(g1101), .QN(n3617) );
  NOR2X0 U3657 ( .IN1(n3618), .IN2(g1110), .QN(n3606) );
  NAND2X0 U3658 ( .IN1(g1107), .IN2(n1658), .QN(n3618) );
  NAND2X0 U3659 ( .IN1(n3619), .IN2(n3620), .QN(g8649) );
  NAND2X0 U3660 ( .IN1(n1016), .IN2(g664), .QN(n3620) );
  NOR2X0 U3661 ( .IN1(n3299), .IN2(n3621), .QN(n3619) );
  NAND2X0 U3662 ( .IN1(n3622), .IN2(n3623), .QN(g8631) );
  NAND2X0 U3663 ( .IN1(n3624), .IN2(n3540), .QN(n3623) );
  NAND2X0 U3664 ( .IN1(n3625), .IN2(n3626), .QN(n3624) );
  NAND2X0 U3665 ( .IN1(n3627), .IN2(g636), .QN(n3626) );
  NAND2X0 U3666 ( .IN1(n3628), .IN2(n3629), .QN(n3627) );
  XOR2X1 U3667 ( .IN1(n3630), .IN2(n3631), .Q(n3629) );
  NAND2X0 U3668 ( .IN1(n3632), .IN2(n3633), .QN(n3631) );
  NAND2X0 U3669 ( .IN1(n3313), .IN2(g639), .QN(n3633) );
  NAND2X0 U3670 ( .IN1(n3634), .IN2(n1692), .QN(n3632) );
  NOR2X0 U3671 ( .IN1(n3315), .IN2(g611), .QN(n3634) );
  INVX0 U3672 ( .INP(n3306), .ZN(n3315) );
  NAND2X0 U3673 ( .IN1(g255), .IN2(g622), .QN(n3630) );
  NOR2X0 U3674 ( .IN1(n3635), .IN2(n3636), .QN(n3628) );
  NOR2X0 U3675 ( .IN1(n3637), .IN2(n3638), .QN(n3635) );
  NAND2X0 U3676 ( .IN1(n1609), .IN2(n1644), .QN(n3638) );
  NAND2X0 U3677 ( .IN1(n3639), .IN2(n3306), .QN(n3637) );
  NAND2X0 U3678 ( .IN1(n3526), .IN2(n1713), .QN(n3625) );
  INVX0 U3679 ( .INP(n3640), .ZN(n3526) );
  NAND2X0 U3680 ( .IN1(n3299), .IN2(n3641), .QN(n3622) );
  NAND2X0 U3681 ( .IN1(n3642), .IN2(n3643), .QN(n3641) );
  INVX0 U3682 ( .INP(n3644), .ZN(n3643) );
  NOR2X0 U3683 ( .IN1(n3645), .IN2(n3646), .QN(n3644) );
  NOR2X0 U3684 ( .IN1(n2918), .IN2(n1622), .QN(n3645) );
  NOR2X0 U3685 ( .IN1(n1716), .IN2(n3647), .QN(n3642) );
  NOR2X0 U3686 ( .IN1(n3648), .IN2(n3649), .QN(n3647) );
  NOR2X0 U3687 ( .IN1(n2907), .IN2(n2917), .QN(n3649) );
  NOR2X0 U3688 ( .IN1(n2906), .IN2(n2919), .QN(n3648) );
  NAND2X0 U3689 ( .IN1(n3650), .IN2(n3651), .QN(g8566) );
  NAND2X0 U3690 ( .IN1(n1653), .IN2(g1669), .QN(n3651) );
  NAND2X0 U3691 ( .IN1(g1690), .IN2(g1687), .QN(n3650) );
  NAND2X0 U3692 ( .IN1(n3652), .IN2(n3653), .QN(g8565) );
  NAND2X0 U3693 ( .IN1(n1653), .IN2(g1666), .QN(n3653) );
  NAND2X0 U3694 ( .IN1(g1690), .IN2(g1684), .QN(n3652) );
  NAND2X0 U3695 ( .IN1(n3654), .IN2(n3655), .QN(g8564) );
  NAND2X0 U3696 ( .IN1(n1653), .IN2(g1663), .QN(n3655) );
  NAND2X0 U3697 ( .IN1(g1690), .IN2(g1681), .QN(n3654) );
  NAND2X0 U3698 ( .IN1(n3656), .IN2(n3657), .QN(g8563) );
  NAND2X0 U3699 ( .IN1(n1653), .IN2(g1660), .QN(n3657) );
  NAND2X0 U3700 ( .IN1(g1690), .IN2(g1678), .QN(n3656) );
  NAND2X0 U3701 ( .IN1(n3658), .IN2(n3659), .QN(g8562) );
  NAND2X0 U3702 ( .IN1(n1653), .IN2(g1657), .QN(n3659) );
  NAND2X0 U3703 ( .IN1(g1690), .IN2(g1675), .QN(n3658) );
  NAND2X0 U3704 ( .IN1(n3660), .IN2(n3661), .QN(g8561) );
  NAND2X0 U3705 ( .IN1(n1653), .IN2(g1654), .QN(n3661) );
  NAND2X0 U3706 ( .IN1(g1690), .IN2(g1672), .QN(n3660) );
  NAND2X0 U3707 ( .IN1(n3662), .IN2(n3663), .QN(g8559) );
  NAND2X0 U3708 ( .IN1(n3664), .IN2(g1878), .QN(n3663) );
  NOR2X0 U3709 ( .IN1(n3273), .IN2(n3665), .QN(n3662) );
  NOR2X0 U3710 ( .IN1(n3666), .IN2(n3199), .QN(g8505) );
  XNOR2X1 U3711 ( .IN1(n3667), .IN2(n1645), .Q(n3666) );
  NOR2X0 U3712 ( .IN1(n3532), .IN2(n3621), .QN(n3667) );
  NOR2X0 U3713 ( .IN1(n1016), .IN2(n2866), .QN(n3621) );
  INVX0 U3714 ( .INP(n3668), .ZN(n3532) );
  NAND2X0 U3715 ( .IN1(n3669), .IN2(n3670), .QN(n3668) );
  NOR2X0 U3716 ( .IN1(g599), .IN2(n3262), .QN(n3670) );
  NOR2X0 U3717 ( .IN1(n3639), .IN2(g611), .QN(n3669) );
  NAND2X0 U3718 ( .IN1(n3671), .IN2(n1645), .QN(n3639) );
  NOR2X0 U3719 ( .IN1(n1607), .IN2(g605), .QN(n3671) );
  NAND2X0 U3720 ( .IN1(n3672), .IN2(n3673), .QN(g8435) );
  NAND2X0 U3721 ( .IN1(n3674), .IN2(g736), .QN(n3673) );
  NAND2X0 U3722 ( .IN1(n3675), .IN2(g727), .QN(n3672) );
  NAND2X0 U3723 ( .IN1(n3676), .IN2(n3677), .QN(g8434) );
  NAND2X0 U3724 ( .IN1(n3674), .IN2(g727), .QN(n3677) );
  NAND2X0 U3725 ( .IN1(n3675), .IN2(g718), .QN(n3676) );
  NAND2X0 U3726 ( .IN1(n3678), .IN2(n3679), .QN(g8433) );
  NAND2X0 U3727 ( .IN1(n3674), .IN2(g718), .QN(n3679) );
  NAND2X0 U3728 ( .IN1(n3675), .IN2(g709), .QN(n3678) );
  NAND2X0 U3729 ( .IN1(n3680), .IN2(n3681), .QN(g8432) );
  NAND2X0 U3730 ( .IN1(n3674), .IN2(g709), .QN(n3681) );
  NAND2X0 U3731 ( .IN1(n3675), .IN2(g700), .QN(n3680) );
  NAND2X0 U3732 ( .IN1(n3682), .IN2(n3683), .QN(g8431) );
  NAND2X0 U3733 ( .IN1(n3674), .IN2(g700), .QN(n3683) );
  NAND2X0 U3734 ( .IN1(n3675), .IN2(g691), .QN(n3682) );
  NAND2X0 U3735 ( .IN1(n3684), .IN2(n3685), .QN(g8430) );
  NAND2X0 U3736 ( .IN1(n3674), .IN2(g691), .QN(n3685) );
  NAND2X0 U3737 ( .IN1(n3675), .IN2(g682), .QN(n3684) );
  NAND2X0 U3738 ( .IN1(n3686), .IN2(n3687), .QN(g8429) );
  NAND2X0 U3739 ( .IN1(n3674), .IN2(g682), .QN(n3687) );
  NAND2X0 U3740 ( .IN1(n3675), .IN2(g673), .QN(n3686) );
  NAND2X0 U3741 ( .IN1(n3688), .IN2(n3689), .QN(g8428) );
  NAND2X0 U3742 ( .IN1(n3674), .IN2(g673), .QN(n3689) );
  NOR2X0 U3743 ( .IN1(n3675), .IN2(n3299), .QN(n3674) );
  NAND2X0 U3744 ( .IN1(n3675), .IN2(g664), .QN(n3688) );
  INVX0 U3745 ( .INP(n1016), .ZN(n3675) );
  NAND2X0 U3746 ( .IN1(n3264), .IN2(n1609), .QN(n1016) );
  NOR2X0 U3747 ( .IN1(n3262), .IN2(n1645), .QN(n3264) );
  NOR2X0 U3748 ( .IN1(n3690), .IN2(n3199), .QN(g8384) );
  XNOR2X1 U3749 ( .IN1(n2867), .IN2(n3691), .Q(n3690) );
  NOR2X0 U3750 ( .IN1(n3665), .IN2(n929), .QN(n3691) );
  NOR2X0 U3751 ( .IN1(n3692), .IN2(g1822), .QN(n929) );
  INVX0 U3752 ( .INP(n3693), .ZN(n3692) );
  NOR2X0 U3753 ( .IN1(n487), .IN2(n3694), .QN(n3693) );
  NOR2X0 U3754 ( .IN1(n3664), .IN2(n2868), .QN(n3665) );
  NAND2X0 U3755 ( .IN1(n1665), .IN2(n3695), .QN(g8352) );
  NAND2X0 U3756 ( .IN1(n1669), .IN2(n3695), .QN(g8349) );
  NAND2X0 U3757 ( .IN1(n1671), .IN2(n3695), .QN(g8347) );
  NAND2X0 U3758 ( .IN1(n2936), .IN2(n3695), .QN(g8340) );
  NAND2X0 U3759 ( .IN1(n1666), .IN2(n3695), .QN(g8335) );
  NAND2X0 U3760 ( .IN1(n1672), .IN2(n3695), .QN(g8331) );
  NAND2X0 U3761 ( .IN1(n1664), .IN2(n3695), .QN(g8328) );
  NAND2X0 U3762 ( .IN1(n1673), .IN2(n3695), .QN(g8323) );
  NAND2X0 U3763 ( .IN1(n1667), .IN2(n3695), .QN(g8318) );
  NAND2X0 U3764 ( .IN1(n1674), .IN2(n3695), .QN(g8316) );
  NAND2X0 U3765 ( .IN1(n1668), .IN2(n3695), .QN(g8313) );
  INVX0 U3766 ( .INP(g82), .ZN(n3695) );
  NAND2X0 U3767 ( .IN1(n3696), .IN2(n3697), .QN(g8288) );
  NAND2X0 U3768 ( .IN1(n3698), .IN2(g1950), .QN(n3697) );
  NAND2X0 U3769 ( .IN1(n3699), .IN2(g1941), .QN(n3696) );
  NAND2X0 U3770 ( .IN1(n3700), .IN2(n3701), .QN(g8287) );
  NAND2X0 U3771 ( .IN1(n3698), .IN2(g1941), .QN(n3701) );
  NAND2X0 U3772 ( .IN1(n3699), .IN2(g1932), .QN(n3700) );
  NAND2X0 U3773 ( .IN1(n3702), .IN2(n3703), .QN(g8286) );
  NAND2X0 U3774 ( .IN1(n3698), .IN2(g1932), .QN(n3703) );
  NAND2X0 U3775 ( .IN1(n3699), .IN2(g1923), .QN(n3702) );
  NAND2X0 U3776 ( .IN1(n3704), .IN2(n3705), .QN(g8285) );
  NAND2X0 U3777 ( .IN1(n3698), .IN2(g1923), .QN(n3705) );
  NAND2X0 U3778 ( .IN1(n3699), .IN2(g1914), .QN(n3704) );
  NAND2X0 U3779 ( .IN1(n3706), .IN2(n3707), .QN(g8284) );
  NAND2X0 U3780 ( .IN1(n3698), .IN2(g1914), .QN(n3707) );
  NAND2X0 U3781 ( .IN1(n3699), .IN2(g1905), .QN(n3706) );
  NAND2X0 U3782 ( .IN1(n3708), .IN2(n3709), .QN(g8283) );
  NAND2X0 U3783 ( .IN1(n3698), .IN2(g1905), .QN(n3709) );
  NAND2X0 U3784 ( .IN1(n3699), .IN2(g1896), .QN(n3708) );
  NAND2X0 U3785 ( .IN1(n3710), .IN2(n3711), .QN(g8282) );
  NAND2X0 U3786 ( .IN1(n3698), .IN2(g1896), .QN(n3711) );
  NAND2X0 U3787 ( .IN1(n3699), .IN2(g1887), .QN(n3710) );
  NAND2X0 U3788 ( .IN1(n3712), .IN2(n3713), .QN(g8281) );
  NAND2X0 U3789 ( .IN1(n3698), .IN2(g1887), .QN(n3713) );
  NOR2X0 U3790 ( .IN1(n3699), .IN2(n3273), .QN(n3698) );
  NAND2X0 U3791 ( .IN1(n3699), .IN2(g1878), .QN(n3712) );
  INVX0 U3792 ( .INP(n3664), .ZN(n3699) );
  NAND2X0 U3793 ( .IN1(n3469), .IN2(n1655), .QN(n3664) );
  NOR2X0 U3794 ( .IN1(n487), .IN2(n2867), .QN(n3469) );
  NOR2X0 U3795 ( .IN1(n1712), .IN2(n3714), .QN(g8260) );
  NOR2X0 U3796 ( .IN1(n1630), .IN2(n3714), .QN(g8254) );
  NOR2X0 U3797 ( .IN1(n1591), .IN2(n3714), .QN(g8250) );
  NOR2X0 U3798 ( .IN1(n3247), .IN2(n3715), .QN(g8245) );
  XOR2X1 U3799 ( .IN1(n1716), .IN2(n3716), .Q(n3715) );
  NOR2X0 U3800 ( .IN1(n2917), .IN2(n3717), .QN(n3716) );
  INVX0 U3801 ( .INP(n1090), .ZN(n3717) );
  NOR2X0 U3802 ( .IN1(n3161), .IN2(n3718), .QN(g8244) );
  NAND2X0 U3803 ( .IN1(n3719), .IN2(n3720), .QN(n3718) );
  NAND2X0 U3804 ( .IN1(n2925), .IN2(n3721), .QN(n3719) );
  NAND2X0 U3805 ( .IN1(n1093), .IN2(g4180), .QN(n3721) );
  NAND2X0 U3806 ( .IN1(n3722), .IN2(n3723), .QN(g8194) );
  NAND2X0 U3807 ( .IN1(n968), .IN2(g1512), .QN(n3723) );
  NAND2X0 U3808 ( .IN1(n3724), .IN2(n3546), .QN(n3722) );
  XOR2X1 U3809 ( .IN1(n3725), .IN2(n5233), .Q(n3724) );
  NAND2X0 U3810 ( .IN1(n3600), .IN2(g1104), .QN(n3725) );
  NOR2X0 U3811 ( .IN1(n3726), .IN2(n1677), .QN(n3600) );
  NAND2X0 U3812 ( .IN1(n3727), .IN2(n3728), .QN(g8193) );
  NAND2X0 U3813 ( .IN1(n968), .IN2(g1639), .QN(n3728) );
  NAND2X0 U3814 ( .IN1(n3729), .IN2(n3546), .QN(n3727) );
  XOR2X1 U3815 ( .IN1(test_so4), .IN2(n3730), .Q(n3729) );
  NOR2X0 U3816 ( .IN1(n3592), .IN2(n3726), .QN(n3730) );
  NAND2X0 U3817 ( .IN1(n1654), .IN2(n1614), .QN(n3726) );
  NAND2X0 U3818 ( .IN1(n1677), .IN2(g1104), .QN(n3592) );
  NOR2X0 U3819 ( .IN1(n3731), .IN2(g1713), .QN(g8173) );
  NOR2X0 U3820 ( .IN1(n3732), .IN2(n3733), .QN(n3731) );
  NOR2X0 U3821 ( .IN1(n2903), .IN2(n3734), .QN(n3733) );
  NOR2X0 U3822 ( .IN1(n1055), .IN2(n1054), .QN(n3734) );
  NOR2X0 U3823 ( .IN1(n3735), .IN2(n3736), .QN(n3732) );
  NAND2X0 U3824 ( .IN1(n1055), .IN2(g1801), .QN(n3736) );
  NAND2X0 U3825 ( .IN1(n3737), .IN2(n1057), .QN(n1055) );
  NOR2X0 U3826 ( .IN1(n3738), .IN2(n1626), .QN(n1057) );
  NOR2X0 U3827 ( .IN1(n2903), .IN2(n2902), .QN(n3737) );
  INVX0 U3828 ( .INP(n1056), .ZN(n3735) );
  NOR2X0 U3829 ( .IN1(n1604), .IN2(n3714), .QN(g8147) );
  NAND2X0 U3830 ( .IN1(n3739), .IN2(g109), .QN(n3714) );
  NAND2X0 U3831 ( .IN1(n3740), .IN2(n5209), .QN(n3739) );
  NOR2X0 U3832 ( .IN1(g881), .IN2(n3741), .QN(n3740) );
  NOR2X0 U3833 ( .IN1(n2942), .IN2(n3742), .QN(g8060) );
  XOR2X1 U3834 ( .IN1(g6002), .IN2(n2821), .Q(n3742) );
  NOR2X0 U3835 ( .IN1(n2939), .IN2(n3743), .QN(g8059) );
  XOR2X1 U3836 ( .IN1(g6042), .IN2(n2818), .Q(n3743) );
  NOR2X0 U3837 ( .IN1(n2940), .IN2(n3744), .QN(g8055) );
  XOR2X1 U3838 ( .IN1(n3745), .IN2(n2893), .Q(n3744) );
  NOR2X0 U3839 ( .IN1(n2941), .IN2(n3746), .QN(g8054) );
  XOR2X1 U3840 ( .IN1(g6015), .IN2(n2908), .Q(n3746) );
  NOR2X0 U3841 ( .IN1(n2942), .IN2(n3747), .QN(g8053) );
  XOR2X1 U3842 ( .IN1(g6045), .IN2(n2817), .Q(n3747) );
  NOR2X0 U3843 ( .IN1(n2939), .IN2(n3748), .QN(g8052) );
  XOR2X1 U3844 ( .IN1(n3749), .IN2(n2819), .Q(n3748) );
  NOR2X0 U3845 ( .IN1(n2940), .IN2(n3750), .QN(g8051) );
  XOR2X1 U3846 ( .IN1(n3751), .IN2(n2823), .Q(n3750) );
  NOR2X0 U3847 ( .IN1(n2941), .IN2(n3752), .QN(g8050) );
  XOR2X1 U3848 ( .IN1(g6026), .IN2(n2909), .Q(n3752) );
  NOR2X0 U3849 ( .IN1(n2942), .IN2(n3753), .QN(g8049) );
  XOR2X1 U3850 ( .IN1(g6049), .IN2(n2820), .Q(n3753) );
  NOR2X0 U3851 ( .IN1(n2939), .IN2(n3754), .QN(g8048) );
  XOR2X1 U3852 ( .IN1(g5996), .IN2(n2842), .Q(n3754) );
  NOR2X0 U3853 ( .IN1(n2940), .IN2(n3755), .QN(g8047) );
  XOR2X1 U3854 ( .IN1(g6035), .IN2(n1704), .Q(n3755) );
  NOR2X0 U3855 ( .IN1(n2941), .IN2(n3756), .QN(g8046) );
  XOR2X1 U3856 ( .IN1(n3757), .IN2(n2824), .Q(n3756) );
  NOR2X0 U3857 ( .IN1(n2942), .IN2(n3758), .QN(g8045) );
  XOR2X1 U3858 ( .IN1(n3759), .IN2(n2894), .Q(n3758) );
  NOR2X0 U3859 ( .IN1(n2939), .IN2(n3760), .QN(g8044) );
  XOR2X1 U3860 ( .IN1(g6038), .IN2(n2816), .Q(n3760) );
  NOR2X0 U3861 ( .IN1(n2940), .IN2(n3761), .QN(g8043) );
  XOR2X1 U3862 ( .IN1(n3762), .IN2(n2895), .Q(n3761) );
  NOR2X0 U3863 ( .IN1(n2941), .IN2(n3763), .QN(g8042) );
  XOR2X1 U3864 ( .IN1(n3764), .IN2(n1703), .Q(n3763) );
  NOR2X0 U3865 ( .IN1(n2942), .IN2(n3765), .QN(g8041) );
  XOR2X1 U3866 ( .IN1(n3766), .IN2(n2859), .Q(n3765) );
  NOR2X0 U3867 ( .IN1(n2939), .IN2(n3767), .QN(g8040) );
  XOR2X1 U3868 ( .IN1(g1474), .IN2(n3768), .Q(n3767) );
  NOR2X0 U3869 ( .IN1(n2940), .IN2(n3769), .QN(g8039) );
  XOR2X1 U3870 ( .IN1(g1470), .IN2(n3770), .Q(n3769) );
  NOR2X0 U3871 ( .IN1(n3247), .IN2(n3771), .QN(g8024) );
  XOR2X1 U3872 ( .IN1(n2917), .IN2(n1090), .Q(n3771) );
  NOR2X0 U3873 ( .IN1(n3161), .IN2(n3772), .QN(g8019) );
  XOR2X1 U3874 ( .IN1(n2920), .IN2(n1093), .Q(n3772) );
  NOR2X0 U3875 ( .IN1(g1713), .IN2(n3773), .QN(g7930) );
  XOR2X1 U3876 ( .IN1(n2902), .IN2(n1056), .Q(n3773) );
  NOR2X0 U3877 ( .IN1(n2941), .IN2(n3774), .QN(g7843) );
  XOR2X1 U3878 ( .IN1(g6000), .IN2(n2822), .Q(n3774) );
  INVX0 U3879 ( .INP(n3775), .ZN(g7709) );
  NAND2X0 U3880 ( .IN1(n3776), .IN2(n3777), .QN(n3775) );
  NOR2X0 U3881 ( .IN1(n1096), .IN2(n1090), .QN(n3777) );
  NAND2X0 U3882 ( .IN1(n3778), .IN2(n3779), .QN(g7660) );
  NAND2X0 U3883 ( .IN1(n3780), .IN2(g654), .QN(n3779) );
  NOR2X0 U3884 ( .IN1(n3528), .IN2(n3299), .QN(n3778) );
  NOR2X0 U3885 ( .IN1(n3781), .IN2(n3782), .QN(g7632) );
  NAND2X0 U3886 ( .IN1(n3783), .IN2(n3784), .QN(n3782) );
  NAND2X0 U3887 ( .IN1(n2687), .IN2(n3785), .QN(n3783) );
  NAND2X0 U3888 ( .IN1(n3786), .IN2(n3540), .QN(g7626) );
  NOR2X0 U3889 ( .IN1(n3787), .IN2(n3788), .QN(n3786) );
  NOR2X0 U3890 ( .IN1(g639), .IN2(n3789), .QN(n3788) );
  NAND2X0 U3891 ( .IN1(n3528), .IN2(n3790), .QN(n3789) );
  NAND2X0 U3892 ( .IN1(n3791), .IN2(n3175), .QN(n3790) );
  INVX0 U3893 ( .INP(n3536), .ZN(n3175) );
  NAND2X0 U3894 ( .IN1(n3640), .IN2(n3792), .QN(n3536) );
  NAND2X0 U3895 ( .IN1(n1593), .IN2(g599), .QN(n3792) );
  NAND2X0 U3896 ( .IN1(n3793), .IN2(n1644), .QN(n3640) );
  NOR2X0 U3897 ( .IN1(n1593), .IN2(g591), .QN(n3793) );
  INVX0 U3898 ( .INP(n3794), .ZN(n3791) );
  NAND2X0 U3899 ( .IN1(n3306), .IN2(n3313), .QN(n3794) );
  NAND2X0 U3900 ( .IN1(n1607), .IN2(g599), .QN(n3313) );
  NAND2X0 U3901 ( .IN1(g605), .IN2(g591), .QN(n3306) );
  NOR2X0 U3902 ( .IN1(n1692), .IN2(n3528), .QN(n3787) );
  NOR2X0 U3903 ( .IN1(n3795), .IN2(n3781), .QN(g7590) );
  NOR2X0 U3904 ( .IN1(n3796), .IN2(g1231), .QN(n3795) );
  NOR2X0 U3905 ( .IN1(n3797), .IN2(n3781), .QN(g7586) );
  NOR2X0 U3906 ( .IN1(n3798), .IN2(n1107), .QN(n3797) );
  NOR2X0 U3907 ( .IN1(n3799), .IN2(n3784), .QN(n1107) );
  INVX0 U3908 ( .INP(n3800), .ZN(n3799) );
  NOR2X0 U3909 ( .IN1(n2688), .IN2(n3801), .QN(n3800) );
  NOR2X0 U3910 ( .IN1(n2686), .IN2(n3796), .QN(n3798) );
  NOR2X0 U3911 ( .IN1(n3802), .IN2(n3784), .QN(n3796) );
  INVX0 U3912 ( .INP(n3803), .ZN(n3802) );
  NOR2X0 U3913 ( .IN1(n2688), .IN2(n2686), .QN(n3803) );
  NOR2X0 U3914 ( .IN1(n3781), .IN2(n3804), .QN(g7581) );
  XNOR2X1 U3915 ( .IN1(n2688), .IN2(n3784), .Q(n3804) );
  NAND2X0 U3916 ( .IN1(n3805), .IN2(n3806), .QN(n3784) );
  NOR2X0 U3917 ( .IN1(n2687), .IN2(n3807), .QN(n3805) );
  NAND2X0 U3918 ( .IN1(n2911), .IN2(g109), .QN(n3781) );
  NOR2X0 U3919 ( .IN1(g1713), .IN2(n3808), .QN(g7541) );
  NAND2X0 U3920 ( .IN1(n3809), .IN2(n3810), .QN(n3808) );
  NAND2X0 U3921 ( .IN1(n1056), .IN2(g1796), .QN(n3810) );
  NAND2X0 U3922 ( .IN1(n1626), .IN2(n3811), .QN(n3809) );
  INVX0 U3923 ( .INP(n1116), .ZN(n3811) );
  NAND2X0 U3924 ( .IN1(n3812), .IN2(n3813), .QN(g7441) );
  NAND2X0 U3925 ( .IN1(n1701), .IN2(g643), .QN(n3813) );
  NOR2X0 U3926 ( .IN1(n3814), .IN2(n3299), .QN(n3812) );
  INVX0 U3927 ( .INP(n3540), .ZN(n3299) );
  NAND2X0 U3928 ( .IN1(n3815), .IN2(n3816), .QN(g7303) );
  NAND2X0 U3929 ( .IN1(n3817), .IN2(test_so6), .QN(n3816) );
  NAND2X0 U3930 ( .IN1(n3806), .IN2(g1265), .QN(n3815) );
  NAND2X0 U3931 ( .IN1(n3818), .IN2(n3819), .QN(g7302) );
  NAND2X0 U3932 ( .IN1(n3817), .IN2(g1265), .QN(n3819) );
  NAND2X0 U3933 ( .IN1(n3806), .IN2(g1260), .QN(n3818) );
  NAND2X0 U3934 ( .IN1(n3820), .IN2(n3821), .QN(g7301) );
  NAND2X0 U3935 ( .IN1(n3817), .IN2(g1260), .QN(n3821) );
  NAND2X0 U3936 ( .IN1(n3806), .IN2(g1255), .QN(n3820) );
  NAND2X0 U3937 ( .IN1(n3822), .IN2(n3823), .QN(g7300) );
  NAND2X0 U3938 ( .IN1(n3817), .IN2(g1255), .QN(n3823) );
  NAND2X0 U3939 ( .IN1(n3806), .IN2(g1250), .QN(n3822) );
  NAND2X0 U3940 ( .IN1(n3824), .IN2(n3825), .QN(g7299) );
  NAND2X0 U3941 ( .IN1(n3817), .IN2(g1250), .QN(n3825) );
  NAND2X0 U3942 ( .IN1(n3806), .IN2(g1245), .QN(n3824) );
  NAND2X0 U3943 ( .IN1(n3826), .IN2(n3827), .QN(g7298) );
  NAND2X0 U3944 ( .IN1(n3817), .IN2(g1245), .QN(n3827) );
  NAND2X0 U3945 ( .IN1(n3806), .IN2(g1240), .QN(n3826) );
  NAND2X0 U3946 ( .IN1(n3828), .IN2(n3829), .QN(g7297) );
  NAND2X0 U3947 ( .IN1(n3817), .IN2(g1240), .QN(n3829) );
  NAND2X0 U3948 ( .IN1(n3806), .IN2(g1235), .QN(n3828) );
  NAND2X0 U3949 ( .IN1(n3830), .IN2(n3831), .QN(g7296) );
  NAND2X0 U3950 ( .IN1(n3817), .IN2(g1235), .QN(n3831) );
  NAND2X0 U3951 ( .IN1(n3806), .IN2(g1275), .QN(n3830) );
  NAND2X0 U3952 ( .IN1(n3832), .IN2(n3833), .QN(g7295) );
  NAND2X0 U3953 ( .IN1(n3817), .IN2(g1280), .QN(n3833) );
  NAND2X0 U3954 ( .IN1(n3806), .IN2(g1284), .QN(n3832) );
  NAND2X0 U3955 ( .IN1(n3834), .IN2(n3835), .QN(g7294) );
  NAND2X0 U3956 ( .IN1(n3817), .IN2(g1284), .QN(n3835) );
  NAND2X0 U3957 ( .IN1(n3806), .IN2(g1292), .QN(n3834) );
  NAND2X0 U3958 ( .IN1(n3836), .IN2(n3837), .QN(g7293) );
  NAND2X0 U3959 ( .IN1(n3817), .IN2(g1292), .QN(n3837) );
  NAND2X0 U3960 ( .IN1(n3806), .IN2(g1296), .QN(n3836) );
  NAND2X0 U3961 ( .IN1(n3838), .IN2(n3839), .QN(g7292) );
  NAND2X0 U3962 ( .IN1(n3817), .IN2(g1296), .QN(n3839) );
  NAND2X0 U3963 ( .IN1(n3806), .IN2(g1300), .QN(n3838) );
  NAND2X0 U3964 ( .IN1(n3840), .IN2(n3841), .QN(g7291) );
  NAND2X0 U3965 ( .IN1(n3817), .IN2(g1300), .QN(n3841) );
  NAND2X0 U3966 ( .IN1(n3806), .IN2(g1304), .QN(n3840) );
  NAND2X0 U3967 ( .IN1(n3842), .IN2(n3843), .QN(g7290) );
  NAND2X0 U3968 ( .IN1(n3817), .IN2(g1304), .QN(n3843) );
  NAND2X0 U3969 ( .IN1(n3806), .IN2(test_so6), .QN(n3842) );
  NAND2X0 U3970 ( .IN1(n3844), .IN2(n3845), .QN(g7257) );
  NAND2X0 U3971 ( .IN1(n3546), .IN2(g1077), .QN(n3845) );
  NAND2X0 U3972 ( .IN1(n968), .IN2(g1032), .QN(n3844) );
  NAND2X0 U3973 ( .IN1(n3846), .IN2(n3847), .QN(g7244) );
  NAND2X0 U3974 ( .IN1(n3546), .IN2(g1071), .QN(n3847) );
  NAND2X0 U3975 ( .IN1(n968), .IN2(g1023), .QN(n3846) );
  NAND2X0 U3976 ( .IN1(n2936), .IN2(n3848), .QN(g7219) );
  NAND2X0 U3977 ( .IN1(n1672), .IN2(n3848), .QN(g7204) );
  NOR2X0 U3978 ( .IN1(n3247), .IN2(n3849), .QN(g7202) );
  XOR2X1 U3979 ( .IN1(n2919), .IN2(n1123), .Q(n3849) );
  NOR2X0 U3980 ( .IN1(n3161), .IN2(n3850), .QN(g7191) );
  XOR2X1 U3981 ( .IN1(n2921), .IN2(n1125), .Q(n3850) );
  NAND2X0 U3982 ( .IN1(n1673), .IN2(n3848), .QN(g7189) );
  NAND2X0 U3983 ( .IN1(n1674), .IN2(n3848), .QN(g7183) );
  NAND2X0 U3984 ( .IN1(n1671), .IN2(n3848), .QN(g7143) );
  NOR2X0 U3985 ( .IN1(n3851), .IN2(n3852), .QN(g7137) );
  XOR2X1 U3986 ( .IN1(n1709), .IN2(n3853), .Q(n3851) );
  NOR2X0 U3987 ( .IN1(n3854), .IN2(n3852), .QN(g7134) );
  NAND2X0 U3988 ( .IN1(n3540), .IN2(n3262), .QN(n3852) );
  INVX0 U3989 ( .INP(n3528), .ZN(n3262) );
  NOR2X0 U3990 ( .IN1(n3780), .IN2(g654), .QN(n3528) );
  NAND2X0 U3991 ( .IN1(n1709), .IN2(n3853), .QN(n3780) );
  NOR2X0 U3992 ( .IN1(n3855), .IN2(n3853), .QN(n3854) );
  INVX0 U3993 ( .INP(n3856), .ZN(n3853) );
  NAND2X0 U3994 ( .IN1(n5226), .IN2(n3814), .QN(n3856) );
  NOR2X0 U3995 ( .IN1(n5226), .IN2(n3814), .QN(n3855) );
  NOR2X0 U3996 ( .IN1(g643), .IN2(n1701), .QN(n3814) );
  NAND2X0 U3997 ( .IN1(n1610), .IN2(n3857), .QN(g7133) );
  XOR2X1 U3998 ( .IN1(g1766), .IN2(n1054), .Q(n3857) );
  NAND2X0 U3999 ( .IN1(n3240), .IN2(n3858), .QN(g7032) );
  NAND2X0 U4000 ( .IN1(g109), .IN2(g123), .QN(n3858) );
  NAND2X0 U4001 ( .IN1(n3859), .IN2(n3860), .QN(n3240) );
  NOR2X0 U4002 ( .IN1(n3861), .IN2(n3862), .QN(n3860) );
  INVX0 U4003 ( .INP(n3863), .ZN(n3862) );
  NOR2X0 U4004 ( .IN1(n3864), .IN2(n3865), .QN(n3863) );
  NAND2X0 U4005 ( .IN1(g6786), .IN2(n1704), .QN(n3864) );
  NAND2X0 U4006 ( .IN1(n3866), .IN2(n3867), .QN(n3861) );
  NOR2X0 U4007 ( .IN1(n2909), .IN2(n2908), .QN(n3867) );
  NOR2X0 U4008 ( .IN1(n2841), .IN2(n2820), .QN(n3866) );
  NOR2X0 U4009 ( .IN1(n3868), .IN2(n3869), .QN(n3859) );
  NAND2X0 U4010 ( .IN1(n3870), .IN2(n3871), .QN(n3869) );
  NOR2X0 U4011 ( .IN1(g158), .IN2(g153), .QN(n3871) );
  NOR2X0 U4012 ( .IN1(g143), .IN2(g148), .QN(n3870) );
  NAND2X0 U4013 ( .IN1(n3872), .IN2(n3873), .QN(n3868) );
  NOR2X0 U4014 ( .IN1(g131), .IN2(g139), .QN(n3873) );
  NOR2X0 U4015 ( .IN1(g135), .IN2(g162), .QN(n3872) );
  NOR2X0 U4016 ( .IN1(n3874), .IN2(g1713), .QN(g6983) );
  NOR2X0 U4017 ( .IN1(n3875), .IN2(n3876), .QN(n3874) );
  NOR2X0 U4018 ( .IN1(n1702), .IN2(n1116), .QN(n3876) );
  NOR2X0 U4019 ( .IN1(n3738), .IN2(n1054), .QN(n1116) );
  NOR2X0 U4020 ( .IN1(n3877), .IN2(n3878), .QN(n3875) );
  NAND2X0 U4021 ( .IN1(n3738), .IN2(g1786), .QN(n3878) );
  NAND2X0 U4022 ( .IN1(n3879), .IN2(n3880), .QN(n3738) );
  NOR2X0 U4023 ( .IN1(n2904), .IN2(n1702), .QN(n3880) );
  NOR2X0 U4024 ( .IN1(n1659), .IN2(n3881), .QN(n3879) );
  NAND2X0 U4025 ( .IN1(n3882), .IN2(n3883), .QN(g6930) );
  NAND2X0 U4026 ( .IN1(n3546), .IN2(g1074), .QN(n3883) );
  INVX0 U4027 ( .INP(n3884), .ZN(n3882) );
  NOR2X0 U4028 ( .IN1(n3546), .IN2(n2791), .QN(n3884) );
  NAND2X0 U4029 ( .IN1(n3885), .IN2(n3886), .QN(g6929) );
  NAND2X0 U4030 ( .IN1(n3219), .IN2(g302), .QN(n3886) );
  NAND2X0 U4031 ( .IN1(n3218), .IN2(g143), .QN(n3885) );
  NAND2X0 U4032 ( .IN1(n3887), .IN2(n3888), .QN(g6924) );
  NAND2X0 U4033 ( .IN1(n3546), .IN2(g1098), .QN(n3888) );
  INVX0 U4034 ( .INP(n3889), .ZN(n3887) );
  NOR2X0 U4035 ( .IN1(n3546), .IN2(n2792), .QN(n3889) );
  NAND2X0 U4036 ( .IN1(n3890), .IN2(n3891), .QN(g6923) );
  NAND2X0 U4037 ( .IN1(n3219), .IN2(g299), .QN(n3891) );
  INVX0 U4038 ( .INP(n3892), .ZN(n3890) );
  NOR2X0 U4039 ( .IN1(n3219), .IN2(n2820), .QN(n3892) );
  NAND2X0 U4040 ( .IN1(n3893), .IN2(n3894), .QN(g6922) );
  NAND2X0 U4041 ( .IN1(n3219), .IN2(g278), .QN(n3894) );
  NAND2X0 U4042 ( .IN1(n3218), .IN2(g162), .QN(n3893) );
  NAND2X0 U4043 ( .IN1(n3895), .IN2(n3896), .QN(g6918) );
  NAND2X0 U4044 ( .IN1(n3546), .IN2(g1095), .QN(n3896) );
  NAND2X0 U4045 ( .IN1(test_so2), .IN2(n968), .QN(n3895) );
  NAND2X0 U4046 ( .IN1(n3897), .IN2(n3898), .QN(g6916) );
  NAND2X0 U4047 ( .IN1(n3219), .IN2(g296), .QN(n3898) );
  NAND2X0 U4048 ( .IN1(n3218), .IN2(g139), .QN(n3897) );
  NAND2X0 U4049 ( .IN1(n3899), .IN2(n3900), .QN(g6915) );
  NAND2X0 U4050 ( .IN1(n3219), .IN2(g275), .QN(n3900) );
  NAND2X0 U4051 ( .IN1(n3218), .IN2(g158), .QN(n3899) );
  NAND2X0 U4052 ( .IN1(n3901), .IN2(n3902), .QN(g6912) );
  NAND2X0 U4053 ( .IN1(n3546), .IN2(g1092), .QN(n3902) );
  NAND2X0 U4054 ( .IN1(n968), .IN2(g1011), .QN(n3901) );
  NAND2X0 U4055 ( .IN1(n3903), .IN2(n3904), .QN(g6911) );
  NAND2X0 U4056 ( .IN1(n3219), .IN2(g293), .QN(n3904) );
  NAND2X0 U4057 ( .IN1(n3218), .IN2(g135), .QN(n3903) );
  NAND2X0 U4058 ( .IN1(n3905), .IN2(n3906), .QN(g6910) );
  NAND2X0 U4059 ( .IN1(n3219), .IN2(g272), .QN(n3906) );
  NAND2X0 U4060 ( .IN1(n3218), .IN2(g153), .QN(n3905) );
  NAND2X0 U4061 ( .IN1(n3907), .IN2(n3908), .QN(g6909) );
  NAND2X0 U4062 ( .IN1(n3909), .IN2(g1868), .QN(n3908) );
  INVX0 U4063 ( .INP(n3910), .ZN(n3907) );
  NAND2X0 U4064 ( .IN1(n3911), .IN2(n3912), .QN(g6908) );
  NAND2X0 U4065 ( .IN1(n3546), .IN2(g1089), .QN(n3912) );
  NAND2X0 U4066 ( .IN1(test_so8), .IN2(n968), .QN(n3911) );
  NAND2X0 U4067 ( .IN1(n3913), .IN2(n3914), .QN(g6907) );
  NAND2X0 U4068 ( .IN1(n3219), .IN2(g290), .QN(n3914) );
  NAND2X0 U4069 ( .IN1(n3218), .IN2(g131), .QN(n3913) );
  NAND2X0 U4070 ( .IN1(n3915), .IN2(n3916), .QN(g6906) );
  NAND2X0 U4071 ( .IN1(n3219), .IN2(g269), .QN(n3916) );
  NAND2X0 U4072 ( .IN1(n3218), .IN2(g148), .QN(n3915) );
  NAND2X0 U4073 ( .IN1(n3917), .IN2(n3918), .QN(g6902) );
  NAND2X0 U4074 ( .IN1(n3546), .IN2(g1086), .QN(n3918) );
  NAND2X0 U4075 ( .IN1(n968), .IN2(g1003), .QN(n3917) );
  NAND2X0 U4076 ( .IN1(n3919), .IN2(n3920), .QN(g6901) );
  NAND2X0 U4077 ( .IN1(n3219), .IN2(g287), .QN(n3920) );
  INVX0 U4078 ( .INP(n3921), .ZN(n3919) );
  NOR2X0 U4079 ( .IN1(n3219), .IN2(n1704), .QN(n3921) );
  NAND2X0 U4080 ( .IN1(n3922), .IN2(n3923), .QN(g6900) );
  NAND2X0 U4081 ( .IN1(n3219), .IN2(g266), .QN(n3923) );
  NAND2X0 U4082 ( .IN1(n3218), .IN2(g178), .QN(n3922) );
  NAND2X0 U4083 ( .IN1(n3924), .IN2(n3925), .QN(g6898) );
  NAND2X0 U4084 ( .IN1(n3546), .IN2(g1083), .QN(n3925) );
  NAND2X0 U4085 ( .IN1(n968), .IN2(g991), .QN(n3924) );
  INVX0 U4086 ( .INP(n3926), .ZN(g6897) );
  NOR2X0 U4087 ( .IN1(n3927), .IN2(n3928), .QN(n3926) );
  NOR2X0 U4088 ( .IN1(n3218), .IN2(n2729), .QN(n3928) );
  NOR2X0 U4089 ( .IN1(n3219), .IN2(n2841), .QN(n3927) );
  INVX0 U4090 ( .INP(n3218), .ZN(n3219) );
  NAND2X0 U4091 ( .IN1(n3865), .IN2(g109), .QN(n3218) );
  NAND2X0 U4092 ( .IN1(n1137), .IN2(n1613), .QN(n3865) );
  NOR2X0 U4093 ( .IN1(n3199), .IN2(n5231), .QN(n1137) );
  NAND2X0 U4094 ( .IN1(n3929), .IN2(n3930), .QN(g6895) );
  NAND2X0 U4095 ( .IN1(n3546), .IN2(g1080), .QN(n3930) );
  INVX0 U4096 ( .INP(n3931), .ZN(n3929) );
  NOR2X0 U4097 ( .IN1(n3546), .IN2(n2870), .QN(n3931) );
  NAND2X0 U4098 ( .IN1(n3932), .IN2(n3933), .QN(g6894) );
  NAND2X0 U4099 ( .IN1(test_so7), .IN2(n3546), .QN(n3933) );
  NAND2X0 U4100 ( .IN1(n968), .IN2(g1027), .QN(n3932) );
  NOR2X0 U4101 ( .IN1(g1696), .IN2(g4089), .QN(g6842) );
  NOR2X0 U4102 ( .IN1(n1629), .IN2(n2941), .QN(g6841) );
  NOR2X0 U4103 ( .IN1(n1598), .IN2(n2942), .QN(g6840) );
  NOR2X0 U4104 ( .IN1(n1711), .IN2(n2939), .QN(g6839) );
  NOR2X0 U4105 ( .IN1(n5228), .IN2(n2940), .QN(g6834) );
  NOR2X0 U4106 ( .IN1(n5232), .IN2(n2941), .QN(g6830) );
  NOR2X0 U4107 ( .IN1(n5230), .IN2(n2942), .QN(g6828) );
  NOR2X0 U4108 ( .IN1(n5227), .IN2(n2939), .QN(g6820) );
  NOR2X0 U4109 ( .IN1(n3934), .IN2(n3910), .QN(g6795) );
  NOR2X0 U4110 ( .IN1(n3935), .IN2(n62), .QN(n3934) );
  INVX0 U4111 ( .INP(n3909), .ZN(n62) );
  NAND2X0 U4112 ( .IN1(n2899), .IN2(n3936), .QN(n3909) );
  NOR2X0 U4113 ( .IN1(n2899), .IN2(n3936), .QN(n3935) );
  NAND2X0 U4114 ( .IN1(n5234), .IN2(n3937), .QN(g6755) );
  NOR2X0 U4115 ( .IN1(n3022), .IN2(n3938), .QN(g6747) );
  NAND2X0 U4116 ( .IN1(n3939), .IN2(g109), .QN(n3938) );
  NAND2X0 U4117 ( .IN1(n5210), .IN2(n5211), .QN(n3939) );
  NAND2X0 U4118 ( .IN1(n3940), .IN2(n3941), .QN(g6679) );
  NAND2X0 U4119 ( .IN1(n142), .IN2(n82), .QN(n3941) );
  INVX0 U4120 ( .INP(n3942), .ZN(n82) );
  NAND2X0 U4121 ( .IN1(n3943), .IN2(n3944), .QN(n3942) );
  NOR2X0 U4122 ( .IN1(n3945), .IN2(n3946), .QN(n3944) );
  NAND2X0 U4123 ( .IN1(g1436), .IN2(g1440), .QN(n3946) );
  NAND2X0 U4124 ( .IN1(g1428), .IN2(g1444), .QN(n3945) );
  NOR2X0 U4125 ( .IN1(n3947), .IN2(n3948), .QN(n3943) );
  NAND2X0 U4126 ( .IN1(n2827), .IN2(n2723), .QN(n3948) );
  NAND2X0 U4127 ( .IN1(n2705), .IN2(n2700), .QN(n3947) );
  INVX0 U4128 ( .INP(n3949), .ZN(n142) );
  NAND2X0 U4129 ( .IN1(n3950), .IN2(n3951), .QN(n3949) );
  NOR2X0 U4130 ( .IN1(n3952), .IN2(n3953), .QN(n3951) );
  NAND2X0 U4131 ( .IN1(g1515), .IN2(g1520), .QN(n3953) );
  NAND2X0 U4132 ( .IN1(g1448), .IN2(g1432), .QN(n3952) );
  NOR2X0 U4133 ( .IN1(n3954), .IN2(n3955), .QN(n3950) );
  NAND2X0 U4134 ( .IN1(n1159), .IN2(g1419), .QN(n3955) );
  INVX0 U4135 ( .INP(g6234), .ZN(n3954) );
  NAND2X0 U4136 ( .IN1(g109), .IN2(g1), .QN(n3940) );
  NAND2X0 U4137 ( .IN1(n1701), .IN2(n3956), .QN(g6672) );
  NAND2X0 U4138 ( .IN1(n3957), .IN2(n3958), .QN(g6656) );
  NAND2X0 U4139 ( .IN1(n80), .IN2(n147), .QN(n3958) );
  INVX0 U4140 ( .INP(n3959), .ZN(n147) );
  NAND2X0 U4141 ( .IN1(n3960), .IN2(n3961), .QN(n3959) );
  NOR2X0 U4142 ( .IN1(n3962), .IN2(n3963), .QN(n3961) );
  NAND2X0 U4143 ( .IN1(g1508), .IN2(g1494), .QN(n3963) );
  NAND2X0 U4144 ( .IN1(g1474), .IN2(g1470), .QN(n3962) );
  NOR2X0 U4145 ( .IN1(n3964), .IN2(n3965), .QN(n3960) );
  NAND2X0 U4146 ( .IN1(n2930), .IN2(g1453), .QN(n3965) );
  NOR2X0 U4147 ( .IN1(n2942), .IN2(n2702), .QN(n2930) );
  INVX0 U4148 ( .INP(n3966), .ZN(n80) );
  NAND2X0 U4149 ( .IN1(n3967), .IN2(n3968), .QN(n3966) );
  NOR2X0 U4150 ( .IN1(n3969), .IN2(n3970), .QN(n3968) );
  NAND2X0 U4151 ( .IN1(n1703), .IN2(g1490), .QN(n3970) );
  NAND2X0 U4152 ( .IN1(g1462), .IN2(g1478), .QN(n3969) );
  NOR2X0 U4153 ( .IN1(n3971), .IN2(n3972), .QN(n3967) );
  NAND2X0 U4154 ( .IN1(n2845), .IN2(n2824), .QN(n3972) );
  NAND2X0 U4155 ( .IN1(n2823), .IN2(n2819), .QN(n3971) );
  NAND2X0 U4156 ( .IN1(g109), .IN2(g4), .QN(n3957) );
  NOR2X0 U4157 ( .IN1(n1666), .IN2(n3973), .QN(g6653) );
  NOR2X0 U4158 ( .IN1(n1664), .IN2(n3973), .QN(g6638) );
  NOR2X0 U4159 ( .IN1(n1667), .IN2(n3973), .QN(g6627) );
  NOR2X0 U4160 ( .IN1(n1668), .IN2(n3973), .QN(g6621) );
  NAND2X0 U4161 ( .IN1(n3974), .IN2(n3975), .QN(g6551) );
  NAND2X0 U4162 ( .IN1(n3181), .IN2(g1546), .QN(n3975) );
  NAND2X0 U4163 ( .IN1(n3180), .IN2(g1478), .QN(n3974) );
  NAND2X0 U4164 ( .IN1(n3976), .IN2(n3977), .QN(g6546) );
  NAND2X0 U4165 ( .IN1(n3181), .IN2(g1564), .QN(n3977) );
  NAND2X0 U4166 ( .IN1(n3180), .IN2(g1453), .QN(n3976) );
  INVX0 U4167 ( .INP(n3978), .ZN(g6545) );
  NOR2X0 U4168 ( .IN1(n3979), .IN2(n3980), .QN(n3978) );
  NOR2X0 U4169 ( .IN1(n3180), .IN2(n2721), .QN(n3980) );
  NOR2X0 U4170 ( .IN1(n3181), .IN2(n2824), .QN(n3979) );
  NAND2X0 U4171 ( .IN1(n3981), .IN2(n3982), .QN(g6542) );
  NAND2X0 U4172 ( .IN1(n3181), .IN2(g1561), .QN(n3982) );
  INVX0 U4173 ( .INP(n3983), .ZN(n3981) );
  NOR2X0 U4174 ( .IN1(n3181), .IN2(n1703), .QN(n3983) );
  NAND2X0 U4175 ( .IN1(n3984), .IN2(n3985), .QN(g6538) );
  NAND2X0 U4176 ( .IN1(n3181), .IN2(g1558), .QN(n3985) );
  NAND2X0 U4177 ( .IN1(n3180), .IN2(g1462), .QN(n3984) );
  NAND2X0 U4178 ( .IN1(n3986), .IN2(n3987), .QN(g6537) );
  NAND2X0 U4179 ( .IN1(n3181), .IN2(g1537), .QN(n3987) );
  NAND2X0 U4180 ( .IN1(n3180), .IN2(g1490), .QN(n3986) );
  NAND2X0 U4181 ( .IN1(n3988), .IN2(n3989), .QN(g6533) );
  NAND2X0 U4182 ( .IN1(n3181), .IN2(g1534), .QN(n3989) );
  NAND2X0 U4183 ( .IN1(n3180), .IN2(g1494), .QN(n3988) );
  NOR2X0 U4184 ( .IN1(n1665), .IN2(n3973), .QN(g6531) );
  NAND2X0 U4185 ( .IN1(n3990), .IN2(n3991), .QN(g6529) );
  NAND2X0 U4186 ( .IN1(n3181), .IN2(g1552), .QN(n3991) );
  NAND2X0 U4187 ( .IN1(n3180), .IN2(g1470), .QN(n3990) );
  NOR2X0 U4188 ( .IN1(n1669), .IN2(n3973), .QN(g6526) );
  NOR2X0 U4189 ( .IN1(g1713), .IN2(n3992), .QN(g6525) );
  XOR2X1 U4190 ( .IN1(g1786), .IN2(n3877), .Q(n3992) );
  NAND2X0 U4191 ( .IN1(n3993), .IN2(n3994), .QN(g6524) );
  NAND2X0 U4192 ( .IN1(n3181), .IN2(g1589), .QN(n3994) );
  NAND2X0 U4193 ( .IN1(n3180), .IN2(g1428), .QN(n3993) );
  NAND2X0 U4194 ( .IN1(n3995), .IN2(n3996), .QN(g6523) );
  NAND2X0 U4195 ( .IN1(n3181), .IN2(g1549), .QN(n3996) );
  NAND2X0 U4196 ( .IN1(n3180), .IN2(g1474), .QN(n3995) );
  NOR2X0 U4197 ( .IN1(g1713), .IN2(n3997), .QN(g6516) );
  INVX0 U4198 ( .INP(n3998), .ZN(n3997) );
  NOR2X0 U4199 ( .IN1(n3999), .IN2(n154), .QN(n3998) );
  INVX0 U4200 ( .INP(n3877), .ZN(n154) );
  NAND2X0 U4201 ( .IN1(n4000), .IN2(g1781), .QN(n3877) );
  NOR2X0 U4202 ( .IN1(g1781), .IN2(n4000), .QN(n3999) );
  NAND2X0 U4203 ( .IN1(n4001), .IN2(n4002), .QN(g6515) );
  NAND2X0 U4204 ( .IN1(n3181), .IN2(g1607), .QN(n4002) );
  NAND2X0 U4205 ( .IN1(n3180), .IN2(g1448), .QN(n4001) );
  NAND2X0 U4206 ( .IN1(n4003), .IN2(n4004), .QN(g6513) );
  NAND2X0 U4207 ( .IN1(n3181), .IN2(g1524), .QN(n4004) );
  NAND2X0 U4208 ( .IN1(n3180), .IN2(g1508), .QN(n4003) );
  NOR2X0 U4209 ( .IN1(n4005), .IN2(g1713), .QN(g6508) );
  NOR2X0 U4210 ( .IN1(n4006), .IN2(n4007), .QN(n4005) );
  NOR2X0 U4211 ( .IN1(n1715), .IN2(n4000), .QN(n4007) );
  NOR2X0 U4212 ( .IN1(n3881), .IN2(n1054), .QN(n4000) );
  NOR2X0 U4213 ( .IN1(n4008), .IN2(n4009), .QN(n4006) );
  NAND2X0 U4214 ( .IN1(test_so5), .IN2(n3881), .QN(n4009) );
  NAND2X0 U4215 ( .IN1(n4010), .IN2(n4011), .QN(g6507) );
  NAND2X0 U4216 ( .IN1(n3181), .IN2(g1604), .QN(n4011) );
  NAND2X0 U4217 ( .IN1(n3180), .IN2(g1444), .QN(n4010) );
  NAND2X0 U4218 ( .IN1(n4012), .IN2(n4013), .QN(g6506) );
  NAND2X0 U4219 ( .IN1(n3181), .IN2(g1583), .QN(n4013) );
  NAND2X0 U4220 ( .IN1(n3180), .IN2(g1424), .QN(n4012) );
  NOR2X0 U4221 ( .IN1(n4014), .IN2(g1713), .QN(g6502) );
  XOR2X1 U4222 ( .IN1(test_so5), .IN2(n4008), .Q(n4014) );
  NAND2X0 U4223 ( .IN1(n364), .IN2(g1766), .QN(n4008) );
  NAND2X0 U4224 ( .IN1(n4015), .IN2(n4016), .QN(g6501) );
  NAND2X0 U4225 ( .IN1(n3181), .IN2(g1601), .QN(n4016) );
  NAND2X0 U4226 ( .IN1(n3180), .IN2(g1440), .QN(n4015) );
  NAND2X0 U4227 ( .IN1(n4017), .IN2(n4018), .QN(g6500) );
  NAND2X0 U4228 ( .IN1(n3181), .IN2(g1580), .QN(n4018) );
  NAND2X0 U4229 ( .IN1(n3180), .IN2(g1411), .QN(n4017) );
  NAND2X0 U4230 ( .IN1(n4019), .IN2(n4020), .QN(g6481) );
  NAND2X0 U4231 ( .IN1(n3181), .IN2(g1598), .QN(n4020) );
  NAND2X0 U4232 ( .IN1(n3180), .IN2(g1436), .QN(n4019) );
  NAND2X0 U4233 ( .IN1(n4021), .IN2(n4022), .QN(g6480) );
  NAND2X0 U4234 ( .IN1(n3181), .IN2(g1577), .QN(n4022) );
  NAND2X0 U4235 ( .IN1(n3180), .IN2(g1419), .QN(n4021) );
  NAND2X0 U4236 ( .IN1(n4023), .IN2(n4024), .QN(g6479) );
  NAND2X0 U4237 ( .IN1(n3181), .IN2(g1595), .QN(n4024) );
  NAND2X0 U4238 ( .IN1(n3180), .IN2(g1432), .QN(n4023) );
  NAND2X0 U4239 ( .IN1(n4025), .IN2(n4026), .QN(g6478) );
  NAND2X0 U4240 ( .IN1(n3181), .IN2(g1574), .QN(n4026) );
  NAND2X0 U4241 ( .IN1(n3180), .IN2(g1515), .QN(n4025) );
  NOR2X0 U4242 ( .IN1(n4027), .IN2(n3910), .QN(g6471) );
  NOR2X0 U4243 ( .IN1(n4028), .IN2(n3936), .QN(n4027) );
  NOR2X0 U4244 ( .IN1(g1861), .IN2(n5234), .QN(n3936) );
  NOR2X0 U4245 ( .IN1(n2901), .IN2(n3033), .QN(n4028) );
  NAND2X0 U4246 ( .IN1(n4029), .IN2(n4030), .QN(g6469) );
  NAND2X0 U4247 ( .IN1(n3181), .IN2(g1571), .QN(n4030) );
  INVX0 U4248 ( .INP(n3180), .ZN(n3181) );
  NAND2X0 U4249 ( .IN1(n3180), .IN2(g1520), .QN(n4029) );
  NAND2X0 U4250 ( .IN1(g109), .IN2(n3964), .QN(n3180) );
  INVX0 U4251 ( .INP(n1159), .ZN(n3964) );
  NOR2X0 U4252 ( .IN1(n2939), .IN2(n4031), .QN(g6439) );
  XOR2X1 U4253 ( .IN1(n4032), .IN2(n4033), .Q(n4031) );
  XOR2X1 U4254 ( .IN1(n2844), .IN2(n2843), .Q(n4033) );
  XOR2X1 U4255 ( .IN1(n2841), .IN2(g153), .Q(n4032) );
  NOR2X0 U4256 ( .IN1(n3741), .IN2(n4034), .QN(g6392) );
  NOR2X0 U4257 ( .IN1(n2940), .IN2(n4035), .QN(n4034) );
  NOR2X0 U4258 ( .IN1(n1603), .IN2(n2940), .QN(g6334) );
  NAND2X0 U4259 ( .IN1(n4036), .IN2(n3776), .QN(g6243) );
  INVX0 U4260 ( .INP(n3247), .ZN(n3776) );
  XNOR2X1 U4261 ( .IN1(n1717), .IN2(n2915), .Q(n4036) );
  NOR2X0 U4262 ( .IN1(n1710), .IN2(n2941), .QN(g6224) );
  NOR2X0 U4263 ( .IN1(n1627), .IN2(n2942), .QN(g6205) );
  NAND2X0 U4264 ( .IN1(n4037), .IN2(n4038), .QN(g6155) );
  NAND2X0 U4265 ( .IN1(g4076), .IN2(g1690), .QN(n4038) );
  NAND2X0 U4266 ( .IN1(n4039), .IN2(n1653), .QN(n4037) );
  NOR2X0 U4267 ( .IN1(n2905), .IN2(n497), .QN(n4039) );
  NOR2X0 U4268 ( .IN1(n3247), .IN2(n4040), .QN(g6126) );
  XOR2X1 U4269 ( .IN1(n2918), .IN2(n3251), .Q(n4040) );
  NOR2X0 U4270 ( .IN1(n3161), .IN2(n4041), .QN(g6123) );
  XOR2X1 U4271 ( .IN1(n2922), .IN2(n1193), .Q(n4041) );
  NAND2X0 U4272 ( .IN1(n4042), .IN2(n4043), .QN(g6099) );
  NAND2X0 U4273 ( .IN1(n4044), .IN2(g342), .QN(n4043) );
  NAND2X0 U4274 ( .IN1(n4045), .IN2(g1074), .QN(n4042) );
  NAND2X0 U4275 ( .IN1(n4046), .IN2(n4047), .QN(g6096) );
  NAND2X0 U4276 ( .IN1(n4044), .IN2(g366), .QN(n4047) );
  NAND2X0 U4277 ( .IN1(n4045), .IN2(g1098), .QN(n4046) );
  NAND2X0 U4278 ( .IN1(n4048), .IN2(n4049), .QN(g6093) );
  NAND2X0 U4279 ( .IN1(n4044), .IN2(g363), .QN(n4049) );
  NAND2X0 U4280 ( .IN1(n4045), .IN2(g1095), .QN(n4048) );
  NAND2X0 U4281 ( .IN1(n4050), .IN2(n4051), .QN(g6088) );
  NAND2X0 U4282 ( .IN1(n4044), .IN2(g360), .QN(n4051) );
  NAND2X0 U4283 ( .IN1(n4045), .IN2(g1092), .QN(n4050) );
  NAND2X0 U4284 ( .IN1(n4052), .IN2(n4053), .QN(g6080) );
  NAND2X0 U4285 ( .IN1(n4044), .IN2(g357), .QN(n4053) );
  NAND2X0 U4286 ( .IN1(n4045), .IN2(g1089), .QN(n4052) );
  NAND2X0 U4287 ( .IN1(n4054), .IN2(n4055), .QN(g6071) );
  NAND2X0 U4288 ( .IN1(n4044), .IN2(g354), .QN(n4055) );
  NAND2X0 U4289 ( .IN1(n4045), .IN2(g1086), .QN(n4054) );
  NAND2X0 U4290 ( .IN1(n4056), .IN2(n4057), .QN(g6068) );
  NAND2X0 U4291 ( .IN1(n4044), .IN2(g351), .QN(n4057) );
  NAND2X0 U4292 ( .IN1(n4045), .IN2(g1083), .QN(n4056) );
  NAND2X0 U4293 ( .IN1(n4058), .IN2(n4059), .QN(g6059) );
  NAND2X0 U4294 ( .IN1(n4044), .IN2(g348), .QN(n4059) );
  NAND2X0 U4295 ( .IN1(n4045), .IN2(g1080), .QN(n4058) );
  NAND2X0 U4296 ( .IN1(n4060), .IN2(n4061), .QN(g6054) );
  NAND2X0 U4297 ( .IN1(n4044), .IN2(g336), .QN(n4061) );
  NAND2X0 U4298 ( .IN1(test_so7), .IN2(n4045), .QN(n4060) );
  NAND2X0 U4299 ( .IN1(n4062), .IN2(n4063), .QN(g6049) );
  NAND2X0 U4300 ( .IN1(n3199), .IN2(g549), .QN(n4062) );
  NAND2X0 U4301 ( .IN1(n4064), .IN2(n4065), .QN(g6045) );
  NAND2X0 U4302 ( .IN1(n3199), .IN2(g575), .QN(n4064) );
  NAND2X0 U4303 ( .IN1(n4066), .IN2(n4067), .QN(g6042) );
  NAND2X0 U4304 ( .IN1(n3199), .IN2(g572), .QN(n4066) );
  NAND2X0 U4305 ( .IN1(n4068), .IN2(n3609), .QN(g6038) );
  NAND2X0 U4306 ( .IN1(g18), .IN2(g237), .QN(n3609) );
  NAND2X0 U4307 ( .IN1(n3199), .IN2(g569), .QN(n4068) );
  NAND2X0 U4308 ( .IN1(n4069), .IN2(n3597), .QN(g6035) );
  NAND2X0 U4309 ( .IN1(g18), .IN2(g231), .QN(n3597) );
  NAND2X0 U4310 ( .IN1(n3199), .IN2(g566), .QN(n4069) );
  NAND2X0 U4311 ( .IN1(n3572), .IN2(n4070), .QN(g6026) );
  NAND2X0 U4312 ( .IN1(n3199), .IN2(g563), .QN(n4070) );
  NAND2X0 U4313 ( .IN1(n3558), .IN2(n4071), .QN(g6015) );
  NAND2X0 U4314 ( .IN1(n3199), .IN2(g560), .QN(n4071) );
  NAND2X0 U4315 ( .IN1(n3614), .IN2(n4072), .QN(g6002) );
  NAND2X0 U4316 ( .IN1(n3199), .IN2(g557), .QN(n4072) );
  NAND2X0 U4317 ( .IN1(n3602), .IN2(n4073), .QN(g6000) );
  NAND2X0 U4318 ( .IN1(n3199), .IN2(g554), .QN(n4073) );
  NAND2X0 U4319 ( .IN1(n3587), .IN2(n4074), .QN(g5996) );
  NAND2X0 U4320 ( .IN1(n3199), .IN2(g546), .QN(n4074) );
  NAND2X0 U4321 ( .IN1(n4075), .IN2(n4076), .QN(g5918) );
  INVX0 U4322 ( .INP(n4077), .ZN(n4076) );
  NOR2X0 U4323 ( .IN1(n2941), .IN2(n1613), .QN(n4077) );
  NAND2X0 U4324 ( .IN1(n4078), .IN2(n4079), .QN(g5914) );
  NAND2X0 U4325 ( .IN1(n4044), .IN2(g345), .QN(n4079) );
  NAND2X0 U4326 ( .IN1(n4045), .IN2(g1077), .QN(n4078) );
  NAND2X0 U4327 ( .IN1(n4080), .IN2(n4081), .QN(g5910) );
  NAND2X0 U4328 ( .IN1(n4044), .IN2(g339), .QN(n4081) );
  NAND2X0 U4329 ( .IN1(n4045), .IN2(g1071), .QN(n4080) );
  NAND2X0 U4330 ( .IN1(n4082), .IN2(n4083), .QN(g5770) );
  NAND2X0 U4331 ( .IN1(n4084), .IN2(n4085), .QN(n4083) );
  NOR2X0 U4332 ( .IN1(n2942), .IN2(g1453), .QN(n4084) );
  NAND2X0 U4333 ( .IN1(g6180), .IN2(n4086), .QN(n4082) );
  INVX0 U4334 ( .INP(n4085), .ZN(n4086) );
  XOR2X1 U4335 ( .IN1(g1508), .IN2(n4087), .Q(n4085) );
  XOR2X1 U4336 ( .IN1(n2859), .IN2(n2845), .Q(n4087) );
  NOR2X0 U4337 ( .IN1(n2939), .IN2(n1628), .QN(g6180) );
  NAND2X0 U4338 ( .IN1(n4088), .IN2(n4089), .QN(g5755) );
  NAND2X0 U4339 ( .IN1(g6333), .IN2(n4090), .QN(n4089) );
  XOR2X1 U4340 ( .IN1(n1619), .IN2(n4091), .Q(n4090) );
  NOR2X0 U4341 ( .IN1(n2940), .IN2(n1678), .QN(g6333) );
  NAND2X0 U4342 ( .IN1(n4092), .IN2(n1678), .QN(n4088) );
  NOR2X0 U4343 ( .IN1(n4093), .IN2(n4094), .QN(n4092) );
  NOR2X0 U4344 ( .IN1(g6331), .IN2(n4091), .QN(n4094) );
  INVX0 U4345 ( .INP(n4095), .ZN(n4091) );
  NOR2X0 U4346 ( .IN1(n2941), .IN2(n1619), .QN(g6331) );
  NOR2X0 U4347 ( .IN1(n4096), .IN2(n4095), .QN(n4093) );
  XOR2X1 U4348 ( .IN1(g1389), .IN2(n4097), .Q(n4095) );
  NOR2X0 U4349 ( .IN1(n37), .IN2(g1386), .QN(n4097) );
  NOR2X0 U4350 ( .IN1(g201), .IN2(n3186), .QN(n37) );
  NAND2X0 U4351 ( .IN1(n4098), .IN2(n4099), .QN(n3186) );
  NOR2X0 U4352 ( .IN1(n4100), .IN2(n4101), .QN(n4099) );
  NAND2X0 U4353 ( .IN1(n4102), .IN2(n4103), .QN(n4101) );
  NOR2X0 U4354 ( .IN1(g207), .IN2(n4104), .QN(n4103) );
  NAND2X0 U4355 ( .IN1(n2690), .IN2(n2689), .QN(n4104) );
  NOR2X0 U4356 ( .IN1(g192), .IN2(n4105), .QN(n4102) );
  NAND2X0 U4357 ( .IN1(n2693), .IN2(n2692), .QN(n4105) );
  NAND2X0 U4358 ( .IN1(n4106), .IN2(n4107), .QN(n4100) );
  NOR2X0 U4359 ( .IN1(g1389), .IN2(n4108), .QN(n4107) );
  NAND2X0 U4360 ( .IN1(n1598), .IN2(n2846), .QN(n4108) );
  NOR2X0 U4361 ( .IN1(g1397), .IN2(n4109), .QN(n4106) );
  NAND2X0 U4362 ( .IN1(n1678), .IN2(n1629), .QN(n4109) );
  NOR2X0 U4363 ( .IN1(n4110), .IN2(n4111), .QN(n4098) );
  NAND2X0 U4364 ( .IN1(n4112), .IN2(n4113), .QN(n4111) );
  NOR2X0 U4365 ( .IN1(n3054), .IN2(n4114), .QN(n4113) );
  NAND2X0 U4366 ( .IN1(n5230), .IN2(n5232), .QN(n4114) );
  INVX0 U4367 ( .INP(n4115), .ZN(n4112) );
  NAND2X0 U4368 ( .IN1(n5227), .IN2(n5212), .QN(n4115) );
  NAND2X0 U4369 ( .IN1(n4116), .IN2(n4117), .QN(n4110) );
  NOR2X0 U4370 ( .IN1(g225), .IN2(n4118), .QN(n4117) );
  NAND2X0 U4371 ( .IN1(n2847), .IN2(n2840), .QN(n4118) );
  NOR2X0 U4372 ( .IN1(g243), .IN2(n4119), .QN(n4116) );
  NAND2X0 U4373 ( .IN1(n2850), .IN2(n2849), .QN(n4119) );
  NOR2X0 U4374 ( .IN1(n2942), .IN2(g201), .QN(n4096) );
  NOR2X0 U4375 ( .IN1(n4120), .IN2(n4121), .QN(g5659) );
  NAND2X0 U4376 ( .IN1(g743), .IN2(g109), .QN(n4121) );
  INVX0 U4377 ( .INP(g744), .ZN(n4120) );
  NOR2X0 U4378 ( .IN1(n4122), .IN2(n4123), .QN(g5658) );
  NAND2X0 U4379 ( .IN1(g741), .IN2(g109), .QN(n4123) );
  INVX0 U4380 ( .INP(g742), .ZN(n4122) );
  NOR2X0 U4381 ( .IN1(n4124), .IN2(n4125), .QN(g5556) );
  NAND2X0 U4382 ( .IN1(n4126), .IN2(n4127), .QN(n4125) );
  NOR2X0 U4383 ( .IN1(n1653), .IN2(n1626), .QN(n4127) );
  NOR2X0 U4384 ( .IN1(n3881), .IN2(g1781), .QN(n4126) );
  NAND2X0 U4385 ( .IN1(n4128), .IN2(test_so5), .QN(n3881) );
  NOR2X0 U4386 ( .IN1(n2897), .IN2(n1715), .QN(n4128) );
  NAND2X0 U4387 ( .IN1(n4129), .IN2(n4130), .QN(n4124) );
  NOR2X0 U4388 ( .IN1(n2903), .IN2(n4131), .QN(n4130) );
  NAND2X0 U4389 ( .IN1(g1786), .IN2(g1707), .QN(n4131) );
  NOR2X0 U4390 ( .IN1(n2902), .IN2(n1702), .QN(n4129) );
  NOR2X0 U4391 ( .IN1(n3251), .IN2(n4132), .QN(g5543) );
  NOR2X0 U4392 ( .IN1(n4133), .IN2(n4134), .QN(n4132) );
  NOR2X0 U4393 ( .IN1(n1717), .IN2(g5849), .QN(n4134) );
  INVX0 U4394 ( .INP(n4135), .ZN(g5849) );
  NOR2X0 U4395 ( .IN1(n3247), .IN2(n2915), .QN(n4135) );
  NOR2X0 U4396 ( .IN1(n1622), .IN2(n3247), .QN(n4133) );
  NAND2X0 U4397 ( .IN1(n4136), .IN2(g109), .QN(n3247) );
  NOR2X0 U4398 ( .IN1(n2900), .IN2(n2684), .QN(n4136) );
  NOR2X0 U4399 ( .IN1(n4137), .IN2(n1622), .QN(n3251) );
  INVX0 U4400 ( .INP(n3646), .ZN(n4137) );
  NOR2X0 U4401 ( .IN1(n2915), .IN2(n1717), .QN(n3646) );
  NAND2X0 U4402 ( .IN1(n4138), .IN2(n4139), .QN(g5529) );
  NAND2X0 U4403 ( .IN1(g4940), .IN2(g4174), .QN(n4139) );
  NAND2X0 U4404 ( .IN1(n4140), .IN2(n2923), .QN(n4138) );
  NOR2X0 U4405 ( .IN1(n2924), .IN2(n3161), .QN(n4140) );
  NAND2X0 U4406 ( .IN1(n4075), .IN2(n4141), .QN(g5445) );
  NAND2X0 U4407 ( .IN1(g109), .IN2(g12), .QN(n4141) );
  NAND2X0 U4408 ( .IN1(n4075), .IN2(n4142), .QN(g5421) );
  NAND2X0 U4409 ( .IN1(g109), .IN2(g9), .QN(n4142) );
  INVX0 U4410 ( .INP(n1195), .ZN(n4075) );
  NAND2X0 U4411 ( .IN1(n4143), .IN2(n4144), .QN(g5404) );
  NAND2X0 U4412 ( .IN1(n3546), .IN2(g1713), .QN(n4144) );
  NAND2X0 U4413 ( .IN1(n968), .IN2(g1718), .QN(n4143) );
  NAND2X0 U4414 ( .IN1(n4145), .IN2(n4146), .QN(g5396) );
  NAND2X0 U4415 ( .IN1(n3546), .IN2(g1710), .QN(n4146) );
  NAND2X0 U4416 ( .IN1(n968), .IN2(g1713), .QN(n4145) );
  NOR2X0 U4417 ( .IN1(n1654), .IN2(n4147), .QN(g5390) );
  NOR2X0 U4418 ( .IN1(n1677), .IN2(n4147), .QN(g5173) );
  NOR2X0 U4419 ( .IN1(n1614), .IN2(n4147), .QN(g5148) );
  NOR2X0 U4420 ( .IN1(n1658), .IN2(n4147), .QN(g5126) );
  NAND2X0 U4421 ( .IN1(g109), .IN2(DFF_126_n1), .QN(n4147) );
  NOR2X0 U4422 ( .IN1(n3546), .IN2(n4148), .QN(g5083) );
  INVX0 U4423 ( .INP(n4149), .ZN(n4148) );
  NOR2X0 U4424 ( .IN1(n4150), .IN2(g4089), .QN(n4149) );
  NOR2X0 U4425 ( .IN1(g4173), .IN2(n3161), .QN(g4940) );
  NAND2X0 U4426 ( .IN1(g109), .IN2(n2938), .QN(n3161) );
  NOR2X0 U4427 ( .IN1(n2933), .IN2(DFF_489_n1), .QN(g4905) );
  NOR2X0 U4428 ( .IN1(n2933), .IN2(DFF_330_n1), .QN(g4903) );
  NOR2X0 U4429 ( .IN1(n2933), .IN2(DFF_385_n1), .QN(g4902) );
  NOR2X0 U4430 ( .IN1(n2931), .IN2(DFF_157_n1), .QN(g4893) );
  INVX0 U4431 ( .INP(n3636), .ZN(g4892) );
  NAND2X0 U4432 ( .IN1(n3956), .IN2(n3059), .QN(n3636) );
  INVX0 U4433 ( .INP(n2931), .ZN(n3956) );
  NOR2X0 U4434 ( .IN1(n2931), .IN2(DFF_136_n1), .QN(g4891) );
  NOR2X0 U4435 ( .IN1(n2931), .IN2(DFF_336_n1), .QN(g4890) );
  NAND2X0 U4436 ( .IN1(n3540), .IN2(n4151), .QN(n2931) );
  NAND2X0 U4437 ( .IN1(n1607), .IN2(g611), .QN(n4151) );
  NAND2X0 U4438 ( .IN1(n4152), .IN2(n4153), .QN(n3540) );
  NOR2X0 U4439 ( .IN1(g591), .IN2(g605), .QN(n4153) );
  NOR2X0 U4440 ( .IN1(g599), .IN2(g611), .QN(n4152) );
  NAND2X0 U4441 ( .IN1(n2912), .IN2(n2911), .QN(g4556) );
  NOR2X0 U4442 ( .IN1(n5233), .IN2(n2939), .QN(g4506) );
  NOR2X0 U4443 ( .IN1(n5229), .IN2(n3546), .QN(g4500) );
  NOR2X0 U4444 ( .IN1(n1617), .IN2(n2940), .QN(g4498) );
  NOR2X0 U4445 ( .IN1(n1660), .IN2(n2941), .QN(g4490) );
  NOR2X0 U4446 ( .IN1(n1597), .IN2(n2942), .QN(g4484) );
  NOR2X0 U4447 ( .IN1(n1706), .IN2(n2939), .QN(g4480) );
  NOR2X0 U4448 ( .IN1(n1705), .IN2(n2940), .QN(g4477) );
  NOR2X0 U4449 ( .IN1(n1708), .IN2(n2941), .QN(g4473) );
  NOR2X0 U4450 ( .IN1(n1618), .IN2(n2942), .QN(g4471) );
  NOR2X0 U4451 ( .IN1(n2939), .IN2(n2935), .QN(g4465) );
  NOR2X0 U4452 ( .IN1(n1685), .IN2(n2939), .QN(g4342) );
  NOR2X0 U4453 ( .IN1(n1686), .IN2(n2940), .QN(g4340) );
  NAND2X0 U4454 ( .IN1(n4154), .IN2(n4155), .QN(g4309) );
  NAND2X0 U4455 ( .IN1(n4156), .IN2(g1806), .QN(n4155) );
  NAND2X0 U4456 ( .IN1(n4157), .IN2(g1762), .QN(n4154) );
  NAND2X0 U4457 ( .IN1(n4158), .IN2(n4159), .QN(g4293) );
  NAND2X0 U4458 ( .IN1(n4156), .IN2(g1801), .QN(n4159) );
  NAND2X0 U4459 ( .IN1(n4157), .IN2(g1759), .QN(n4158) );
  NAND2X0 U4460 ( .IN1(n4160), .IN2(n4161), .QN(g4283) );
  NAND2X0 U4461 ( .IN1(n4156), .IN2(g1796), .QN(n4161) );
  NAND2X0 U4462 ( .IN1(n4157), .IN2(g1756), .QN(n4160) );
  NAND2X0 U4463 ( .IN1(n4162), .IN2(n4163), .QN(g4274) );
  NAND2X0 U4464 ( .IN1(n4156), .IN2(g1791), .QN(n4163) );
  NAND2X0 U4465 ( .IN1(n4157), .IN2(g1753), .QN(n4162) );
  NAND2X0 U4466 ( .IN1(n4164), .IN2(n4165), .QN(g4264) );
  NAND2X0 U4467 ( .IN1(n4156), .IN2(g1786), .QN(n4165) );
  NAND2X0 U4468 ( .IN1(n4157), .IN2(g1750), .QN(n4164) );
  NAND2X0 U4469 ( .IN1(n4166), .IN2(n4167), .QN(g4255) );
  NAND2X0 U4470 ( .IN1(n4156), .IN2(g1781), .QN(n4167) );
  NAND2X0 U4471 ( .IN1(n4157), .IN2(g1747), .QN(n4166) );
  NAND2X0 U4472 ( .IN1(n4168), .IN2(n4169), .QN(g4239) );
  NAND2X0 U4473 ( .IN1(n4156), .IN2(g1776), .QN(n4169) );
  NAND2X0 U4474 ( .IN1(n4157), .IN2(g1744), .QN(n4168) );
  NAND2X0 U4475 ( .IN1(n4170), .IN2(n4171), .QN(g4238) );
  NAND2X0 U4476 ( .IN1(n4156), .IN2(test_so5), .QN(n4171) );
  NAND2X0 U4477 ( .IN1(n4157), .IN2(g1741), .QN(n4170) );
  NAND2X0 U4478 ( .IN1(n4172), .IN2(n4173), .QN(g4231) );
  NAND2X0 U4479 ( .IN1(n4156), .IN2(g1766), .QN(n4173) );
  INVX0 U4480 ( .INP(n4157), .ZN(n4156) );
  NAND2X0 U4481 ( .IN1(n4157), .IN2(g1738), .QN(n4172) );
  NAND2X0 U4482 ( .IN1(g1700), .IN2(DFF_275_n1), .QN(g4089) );
  NOR2X0 U4483 ( .IN1(g1707), .IN2(n497), .QN(g4076) );
  INVX0 U4484 ( .INP(g1700), .ZN(n497) );
  NOR2X0 U4485 ( .IN1(n2900), .IN2(n4174), .QN(g3462) );
  NOR2X0 U4486 ( .IN1(n4175), .IN2(n3973), .QN(n4174) );
  NOR2X0 U4487 ( .IN1(n1647), .IN2(g750), .QN(n4175) );
  NOR2X0 U4488 ( .IN1(n4176), .IN2(n4177), .QN(g3381) );
  NAND2X0 U4489 ( .IN1(g932), .IN2(g928), .QN(n4177) );
  NAND2X0 U4490 ( .IN1(g936), .IN2(g940), .QN(n4176) );
  INVX0 U4491 ( .INP(g23), .ZN(g3327) );
  NOR2X0 U4492 ( .IN1(g1610), .IN2(g1737), .QN(g2478) );
  NAND2X0 U4493 ( .IN1(n4178), .IN2(n4179), .QN(g11647) );
  NAND2X0 U4494 ( .IN1(n3848), .IN2(g336), .QN(n4179) );
  NAND2X0 U4495 ( .IN1(n3973), .IN2(n4180), .QN(n4178) );
  NAND2X0 U4496 ( .IN1(n4181), .IN2(n4182), .QN(n4180) );
  NAND2X0 U4497 ( .IN1(n4183), .IN2(n4184), .QN(n4182) );
  NAND2X0 U4498 ( .IN1(n4185), .IN2(n4186), .QN(n4181) );
  NOR2X0 U4499 ( .IN1(n4187), .IN2(n4188), .QN(g11641) );
  NOR2X0 U4500 ( .IN1(n4189), .IN2(n4190), .QN(n4187) );
  NOR2X0 U4501 ( .IN1(n1721), .IN2(n2), .QN(n4190) );
  NOR2X0 U4502 ( .IN1(n4191), .IN2(n1227), .QN(n2) );
  NOR2X0 U4503 ( .IN1(n3209), .IN2(n4192), .QN(n4189) );
  NAND2X0 U4504 ( .IN1(n9), .IN2(n4191), .QN(n4192) );
  INVX0 U4505 ( .INP(n2932), .ZN(n4191) );
  NOR2X0 U4506 ( .IN1(n3209), .IN2(n1721), .QN(n2932) );
  NAND2X0 U4507 ( .IN1(n4193), .IN2(g1341), .QN(n3209) );
  NOR2X0 U4508 ( .IN1(n2879), .IN2(n2878), .QN(n4193) );
  NOR2X0 U4509 ( .IN1(n4194), .IN2(n4188), .QN(g11640) );
  NOR2X0 U4510 ( .IN1(n4195), .IN2(n4196), .QN(n4194) );
  INVX0 U4511 ( .INP(n4197), .ZN(n4196) );
  NAND2X0 U4512 ( .IN1(n1231), .IN2(n1232), .QN(n4197) );
  NOR2X0 U4513 ( .IN1(n2878), .IN2(n4198), .QN(n4195) );
  NOR2X0 U4514 ( .IN1(n1227), .IN2(n4199), .QN(n4198) );
  NAND2X0 U4515 ( .IN1(g1341), .IN2(g1336), .QN(n4199) );
  NOR2X0 U4516 ( .IN1(n4188), .IN2(n4200), .QN(g11639) );
  XOR2X1 U4517 ( .IN1(n2877), .IN2(n1231), .Q(n4200) );
  NOR2X0 U4518 ( .IN1(n4188), .IN2(n4201), .QN(g11636) );
  XOR2X1 U4519 ( .IN1(n2879), .IN2(n9), .Q(n4201) );
  NAND2X0 U4520 ( .IN1(n4202), .IN2(g109), .QN(n4188) );
  NAND2X0 U4521 ( .IN1(n4203), .IN2(n5217), .QN(n4202) );
  NOR2X0 U4522 ( .IN1(n2911), .IN2(n4204), .QN(n4203) );
  INVX0 U4523 ( .INP(n3211), .ZN(n4204) );
  NAND2X0 U4524 ( .IN1(n4205), .IN2(n4206), .QN(g11625) );
  NAND2X0 U4525 ( .IN1(n3848), .IN2(g345), .QN(n4206) );
  NAND2X0 U4526 ( .IN1(n3973), .IN2(n4207), .QN(n4205) );
  XOR2X1 U4527 ( .IN1(n4183), .IN2(n4186), .Q(n4207) );
  NOR2X0 U4528 ( .IN1(n4208), .IN2(n4209), .QN(n4186) );
  NOR2X0 U4529 ( .IN1(n1239), .IN2(n1681), .QN(n4209) );
  NOR2X0 U4530 ( .IN1(n4210), .IN2(n34), .QN(n4208) );
  XOR2X1 U4531 ( .IN1(n4211), .IN2(n4212), .Q(n4210) );
  NAND2X0 U4532 ( .IN1(n1594), .IN2(n4213), .QN(n4211) );
  XOR2X1 U4533 ( .IN1(n4214), .IN2(n4215), .Q(n4183) );
  XOR2X1 U4534 ( .IN1(n4216), .IN2(n4217), .Q(n4215) );
  XOR2X1 U4535 ( .IN1(n4218), .IN2(n4219), .Q(n4217) );
  XNOR2X1 U4536 ( .IN1(n4220), .IN2(n4221), .Q(n4219) );
  XNOR2X1 U4537 ( .IN1(n4222), .IN2(n4223), .Q(n4218) );
  XOR2X1 U4538 ( .IN1(n4224), .IN2(n4225), .Q(n4216) );
  XOR2X1 U4539 ( .IN1(n4226), .IN2(n4227), .Q(n4225) );
  XOR2X1 U4540 ( .IN1(n4228), .IN2(n4229), .Q(n4224) );
  NAND2X0 U4541 ( .IN1(n4230), .IN2(n4231), .QN(g11610) );
  NAND2X0 U4542 ( .IN1(n4232), .IN2(g1806), .QN(n4231) );
  NAND2X0 U4543 ( .IN1(n4233), .IN2(g1333), .QN(n4230) );
  NAND2X0 U4544 ( .IN1(n4234), .IN2(n4235), .QN(g11609) );
  NAND2X0 U4545 ( .IN1(n4232), .IN2(g1801), .QN(n4235) );
  NAND2X0 U4546 ( .IN1(n4233), .IN2(g1330), .QN(n4234) );
  NAND2X0 U4547 ( .IN1(n4236), .IN2(n4237), .QN(g11608) );
  NAND2X0 U4548 ( .IN1(n4232), .IN2(g1796), .QN(n4237) );
  NAND2X0 U4549 ( .IN1(n4233), .IN2(g1327), .QN(n4236) );
  NAND2X0 U4550 ( .IN1(n4238), .IN2(n4239), .QN(g11607) );
  NAND2X0 U4551 ( .IN1(n4232), .IN2(g1791), .QN(n4239) );
  NAND2X0 U4552 ( .IN1(n4233), .IN2(g1324), .QN(n4238) );
  NAND2X0 U4553 ( .IN1(n4240), .IN2(n4241), .QN(g11606) );
  NAND2X0 U4554 ( .IN1(n4232), .IN2(g1786), .QN(n4241) );
  NAND2X0 U4555 ( .IN1(n4233), .IN2(g1321), .QN(n4240) );
  NAND2X0 U4556 ( .IN1(n4242), .IN2(n4243), .QN(g11605) );
  NAND2X0 U4557 ( .IN1(n4232), .IN2(g1781), .QN(n4243) );
  NAND2X0 U4558 ( .IN1(n4233), .IN2(g1318), .QN(n4242) );
  NAND2X0 U4559 ( .IN1(n4244), .IN2(n4245), .QN(g11604) );
  NAND2X0 U4560 ( .IN1(n4232), .IN2(g1776), .QN(n4245) );
  NAND2X0 U4561 ( .IN1(n4233), .IN2(g1314), .QN(n4244) );
  NAND2X0 U4562 ( .IN1(n4246), .IN2(n4247), .QN(g11603) );
  NAND2X0 U4563 ( .IN1(test_so9), .IN2(n4233), .QN(n4247) );
  NAND2X0 U4564 ( .IN1(n4232), .IN2(test_so5), .QN(n4246) );
  NAND2X0 U4565 ( .IN1(n4248), .IN2(n4249), .QN(g11602) );
  NAND2X0 U4566 ( .IN1(n4232), .IN2(g1766), .QN(n4249) );
  INVX0 U4567 ( .INP(n4233), .ZN(n4232) );
  NAND2X0 U4568 ( .IN1(n4233), .IN2(g1308), .QN(n4248) );
  NAND2X0 U4569 ( .IN1(n9), .IN2(g1317), .QN(n4233) );
  INVX0 U4570 ( .INP(n1227), .ZN(n9) );
  NAND2X0 U4571 ( .IN1(n4250), .IN2(n3806), .QN(n1227) );
  NOR2X0 U4572 ( .IN1(n4251), .IN2(n4252), .QN(n4250) );
  NOR2X0 U4573 ( .IN1(n4253), .IN2(n4254), .QN(n4251) );
  NAND2X0 U4574 ( .IN1(n4255), .IN2(n4256), .QN(n4254) );
  NOR2X0 U4575 ( .IN1(n4257), .IN2(n4258), .QN(n4256) );
  NAND2X0 U4576 ( .IN1(n4259), .IN2(n4260), .QN(n4258) );
  XOR2X1 U4577 ( .IN1(n2830), .IN2(g1250), .Q(n4260) );
  XOR2X1 U4578 ( .IN1(n1871), .IN2(g1235), .Q(n4259) );
  XOR2X1 U4579 ( .IN1(n2803), .IN2(n2792), .Q(n4257) );
  NOR2X0 U4580 ( .IN1(n4261), .IN2(n4262), .QN(n4255) );
  XOR2X1 U4581 ( .IN1(n2872), .IN2(n2871), .Q(n4262) );
  XOR2X1 U4582 ( .IN1(n2870), .IN2(n2869), .Q(n4261) );
  NAND2X0 U4583 ( .IN1(n4263), .IN2(n4264), .QN(n4253) );
  NOR2X0 U4584 ( .IN1(n4265), .IN2(n4266), .QN(n4264) );
  NAND2X0 U4585 ( .IN1(n4267), .IN2(n4268), .QN(n4266) );
  XOR2X1 U4586 ( .IN1(test_so2), .IN2(n2802), .Q(n4268) );
  XNOR2X1 U4587 ( .IN1(n4269), .IN2(n4270), .Q(n4267) );
  XNOR2X1 U4588 ( .IN1(n2766), .IN2(test_so6), .Q(n4265) );
  NOR2X0 U4589 ( .IN1(n4271), .IN2(n4272), .QN(n4263) );
  XOR2X1 U4590 ( .IN1(n2805), .IN2(n2791), .Q(n4272) );
  XOR2X1 U4591 ( .IN1(test_so8), .IN2(g1245), .Q(n4271) );
  NAND2X0 U4592 ( .IN1(n4273), .IN2(n4274), .QN(g11579) );
  NAND2X0 U4593 ( .IN1(n968), .IN2(g1618), .QN(n4274) );
  NAND2X0 U4594 ( .IN1(n4275), .IN2(n3546), .QN(n4273) );
  XOR2X1 U4595 ( .IN1(g1610), .IN2(n4276), .Q(n4275) );
  NAND2X0 U4596 ( .IN1(n4277), .IN2(n4278), .QN(n4276) );
  NAND2X0 U4597 ( .IN1(n4279), .IN2(n4280), .QN(n4278) );
  NAND2X0 U4598 ( .IN1(n1262), .IN2(n3250), .QN(n4280) );
  NAND2X0 U4599 ( .IN1(n4281), .IN2(n4282), .QN(n3250) );
  INVX0 U4600 ( .INP(n4283), .ZN(n1262) );
  NOR2X0 U4601 ( .IN1(n4282), .IN2(n4281), .QN(n4283) );
  NAND2X0 U4602 ( .IN1(n4284), .IN2(n4285), .QN(n4281) );
  INVX0 U4603 ( .INP(n4286), .ZN(n4285) );
  NOR2X0 U4604 ( .IN1(n1685), .IN2(n1686), .QN(n4286) );
  NAND2X0 U4605 ( .IN1(n4287), .IN2(n1686), .QN(n4284) );
  NOR2X0 U4606 ( .IN1(n4288), .IN2(g1149), .QN(n4287) );
  NOR2X0 U4607 ( .IN1(n4289), .IN2(n4290), .QN(n4288) );
  NAND2X0 U4608 ( .IN1(n4291), .IN2(n4292), .QN(n4290) );
  NOR2X0 U4609 ( .IN1(g1166), .IN2(n4293), .QN(n4292) );
  NAND2X0 U4610 ( .IN1(n2838), .IN2(n1708), .QN(n4293) );
  NOR2X0 U4611 ( .IN1(g1160), .IN2(n4294), .QN(n4291) );
  NAND2X0 U4612 ( .IN1(n5213), .IN2(n5233), .QN(n4294) );
  NAND2X0 U4613 ( .IN1(n4295), .IN2(n4296), .QN(n4289) );
  NOR2X0 U4614 ( .IN1(n4297), .IN2(n4298), .QN(n4296) );
  NAND2X0 U4615 ( .IN1(n1618), .IN2(n1617), .QN(n4298) );
  NAND2X0 U4616 ( .IN1(n1597), .IN2(n2935), .QN(n4297) );
  NOR2X0 U4617 ( .IN1(g1133), .IN2(n4299), .QN(n4295) );
  NAND2X0 U4618 ( .IN1(n1705), .IN2(n1660), .QN(n4299) );
  NAND2X0 U4619 ( .IN1(n1677), .IN2(n3612), .QN(n4282) );
  INVX0 U4620 ( .INP(n4300), .ZN(n3612) );
  NAND2X0 U4621 ( .IN1(n1658), .IN2(n3591), .QN(n4300) );
  NOR2X0 U4622 ( .IN1(g1107), .IN2(n1654), .QN(n3591) );
  NAND2X0 U4623 ( .IN1(n1260), .IN2(n4301), .QN(n4277) );
  INVX0 U4624 ( .INP(n4279), .ZN(n4301) );
  NAND2X0 U4625 ( .IN1(n4302), .IN2(n4303), .QN(g11514) );
  NAND2X0 U4626 ( .IN1(n4304), .IN2(n4305), .QN(n4303) );
  INVX0 U4627 ( .INP(n4306), .ZN(n4305) );
  NOR2X0 U4628 ( .IN1(n2940), .IN2(g1419), .QN(n4304) );
  NAND2X0 U4629 ( .IN1(g6193), .IN2(n4306), .QN(n4302) );
  XOR2X1 U4630 ( .IN1(n4307), .IN2(n4308), .Q(n4306) );
  XOR2X1 U4631 ( .IN1(n2825), .IN2(n2700), .Q(n4308) );
  XOR2X1 U4632 ( .IN1(n4279), .IN2(n1627), .Q(n4307) );
  NAND2X0 U4633 ( .IN1(n4309), .IN2(n4310), .QN(n4279) );
  NAND2X0 U4634 ( .IN1(g18), .IN2(g201), .QN(n4310) );
  NAND2X0 U4635 ( .IN1(n4311), .IN2(n3199), .QN(n4309) );
  NAND2X0 U4636 ( .IN1(n4312), .IN2(n4313), .QN(n4311) );
  NAND2X0 U4637 ( .IN1(n4314), .IN2(n1699), .QN(n4313) );
  NAND2X0 U4638 ( .IN1(n4315), .IN2(n4316), .QN(n4312) );
  NAND2X0 U4639 ( .IN1(n4317), .IN2(n4318), .QN(n4316) );
  INVX0 U4640 ( .INP(n4314), .ZN(n4315) );
  NOR2X0 U4641 ( .IN1(n4319), .IN2(n4320), .QN(n4314) );
  NAND2X0 U4642 ( .IN1(n5223), .IN2(n5222), .QN(n4320) );
  NAND2X0 U4643 ( .IN1(n5221), .IN2(n5220), .QN(n4319) );
  NOR2X0 U4644 ( .IN1(n2941), .IN2(n1602), .QN(g6193) );
  NAND2X0 U4645 ( .IN1(n4321), .IN2(n4322), .QN(g11488) );
  NAND2X0 U4646 ( .IN1(n3848), .IN2(g342), .QN(n4322) );
  INVX0 U4647 ( .INP(n4323), .ZN(n4321) );
  NOR2X0 U4648 ( .IN1(n3848), .IN2(n4229), .QN(n4323) );
  NOR2X0 U4649 ( .IN1(n4324), .IN2(n4325), .QN(n4229) );
  NOR2X0 U4650 ( .IN1(n1239), .IN2(n2638), .QN(n4325) );
  NOR2X0 U4651 ( .IN1(n4326), .IN2(n34), .QN(n4324) );
  XOR2X1 U4652 ( .IN1(n4327), .IN2(n1620), .Q(n4326) );
  NOR2X0 U4653 ( .IN1(n4328), .IN2(n1641), .QN(n4327) );
  NAND2X0 U4654 ( .IN1(n4329), .IN2(n4330), .QN(g11487) );
  NAND2X0 U4655 ( .IN1(n3848), .IN2(g366), .QN(n4330) );
  INVX0 U4656 ( .INP(n4331), .ZN(n4329) );
  NOR2X0 U4657 ( .IN1(n3848), .IN2(n4228), .QN(n4331) );
  NOR2X0 U4658 ( .IN1(n4332), .IN2(n4333), .QN(n4228) );
  NOR2X0 U4659 ( .IN1(n1239), .IN2(n2857), .QN(n4333) );
  NOR2X0 U4660 ( .IN1(n4334), .IN2(n34), .QN(n4332) );
  XOR2X1 U4661 ( .IN1(n1679), .IN2(n4335), .Q(n4334) );
  NOR2X0 U4662 ( .IN1(n4328), .IN2(g456), .QN(n4335) );
  NAND2X0 U4663 ( .IN1(n4336), .IN2(n1594), .QN(n4328) );
  NOR2X0 U4664 ( .IN1(n1606), .IN2(g466), .QN(n4336) );
  NAND2X0 U4665 ( .IN1(n4337), .IN2(n4338), .QN(g11486) );
  NAND2X0 U4666 ( .IN1(n3848), .IN2(g363), .QN(n4338) );
  INVX0 U4667 ( .INP(n4339), .ZN(n4337) );
  NOR2X0 U4668 ( .IN1(n3848), .IN2(n4227), .QN(n4339) );
  NOR2X0 U4669 ( .IN1(n4340), .IN2(n4341), .QN(n4227) );
  NOR2X0 U4670 ( .IN1(n1239), .IN2(n2637), .QN(n4341) );
  NOR2X0 U4671 ( .IN1(n4342), .IN2(n34), .QN(n4340) );
  XOR2X1 U4672 ( .IN1(n1600), .IN2(n4343), .Q(n4342) );
  NOR2X0 U4673 ( .IN1(g471), .IN2(n4344), .QN(n4343) );
  NAND2X0 U4674 ( .IN1(n4345), .IN2(n4346), .QN(g11485) );
  NAND2X0 U4675 ( .IN1(n3848), .IN2(g360), .QN(n4346) );
  INVX0 U4676 ( .INP(n4347), .ZN(n4345) );
  NOR2X0 U4677 ( .IN1(n3848), .IN2(n4226), .QN(n4347) );
  NOR2X0 U4678 ( .IN1(n4348), .IN2(n4349), .QN(n4226) );
  NOR2X0 U4679 ( .IN1(n1239), .IN2(n2836), .QN(n4349) );
  NOR2X0 U4680 ( .IN1(n4350), .IN2(n34), .QN(n4348) );
  XOR2X1 U4681 ( .IN1(n4351), .IN2(g501), .Q(n4350) );
  NAND2X0 U4682 ( .IN1(n4352), .IN2(g461), .QN(n4351) );
  NAND2X0 U4683 ( .IN1(n4353), .IN2(n4354), .QN(g11484) );
  NAND2X0 U4684 ( .IN1(n3848), .IN2(g357), .QN(n4354) );
  NAND2X0 U4685 ( .IN1(n3973), .IN2(n4355), .QN(n4353) );
  INVX0 U4686 ( .INP(n4223), .ZN(n4355) );
  NOR2X0 U4687 ( .IN1(n4356), .IN2(n4357), .QN(n4223) );
  NOR2X0 U4688 ( .IN1(n1239), .IN2(n2832), .QN(n4357) );
  NOR2X0 U4689 ( .IN1(n4358), .IN2(n34), .QN(n4356) );
  XOR2X1 U4690 ( .IN1(n1689), .IN2(n4359), .Q(n4358) );
  NOR2X0 U4691 ( .IN1(n4360), .IN2(n4361), .QN(n4359) );
  NAND2X0 U4692 ( .IN1(n1594), .IN2(n1606), .QN(n4361) );
  NAND2X0 U4693 ( .IN1(g456), .IN2(g466), .QN(n4360) );
  NAND2X0 U4694 ( .IN1(n4362), .IN2(n4363), .QN(g11483) );
  NAND2X0 U4695 ( .IN1(n3848), .IN2(g354), .QN(n4363) );
  NAND2X0 U4696 ( .IN1(n3973), .IN2(n4222), .QN(n4362) );
  NAND2X0 U4697 ( .IN1(n4364), .IN2(n4365), .QN(n4222) );
  INVX0 U4698 ( .INP(n4366), .ZN(n4365) );
  NOR2X0 U4699 ( .IN1(n1239), .IN2(n2876), .QN(n4366) );
  NAND2X0 U4700 ( .IN1(n4367), .IN2(n1239), .QN(n4364) );
  XOR2X1 U4701 ( .IN1(n4368), .IN2(n1691), .Q(n4367) );
  NAND2X0 U4702 ( .IN1(n4352), .IN2(n1594), .QN(n4368) );
  NOR2X0 U4703 ( .IN1(n4369), .IN2(g456), .QN(n4352) );
  NAND2X0 U4704 ( .IN1(g466), .IN2(n1606), .QN(n4369) );
  NAND2X0 U4705 ( .IN1(n4370), .IN2(n4371), .QN(g11482) );
  NAND2X0 U4706 ( .IN1(n3848), .IN2(g351), .QN(n4371) );
  NAND2X0 U4707 ( .IN1(n3973), .IN2(n4214), .QN(n4370) );
  NAND2X0 U4708 ( .IN1(n4372), .IN2(n4373), .QN(n4214) );
  NAND2X0 U4709 ( .IN1(n34), .IN2(g318), .QN(n4373) );
  NAND2X0 U4710 ( .IN1(n4374), .IN2(n1239), .QN(n4372) );
  XOR2X1 U4711 ( .IN1(n4375), .IN2(n1621), .Q(n4374) );
  NAND2X0 U4712 ( .IN1(n4213), .IN2(g461), .QN(n4375) );
  NOR2X0 U4713 ( .IN1(n4376), .IN2(g466), .QN(n4213) );
  NAND2X0 U4714 ( .IN1(g456), .IN2(n1606), .QN(n4376) );
  NAND2X0 U4715 ( .IN1(n4377), .IN2(n4378), .QN(g11481) );
  NAND2X0 U4716 ( .IN1(n3848), .IN2(g348), .QN(n4378) );
  NAND2X0 U4717 ( .IN1(n3973), .IN2(n4221), .QN(n4377) );
  NAND2X0 U4718 ( .IN1(n4379), .IN2(n4380), .QN(n4221) );
  INVX0 U4719 ( .INP(n4381), .ZN(n4380) );
  NOR2X0 U4720 ( .IN1(n1239), .IN2(n2874), .QN(n4381) );
  NAND2X0 U4721 ( .IN1(n4382), .IN2(n1239), .QN(n4379) );
  XOR2X1 U4722 ( .IN1(g481), .IN2(n4383), .Q(n4382) );
  NOR2X0 U4723 ( .IN1(g471), .IN2(n4384), .QN(n4383) );
  NAND2X0 U4724 ( .IN1(n4385), .IN2(n4386), .QN(g11478) );
  NAND2X0 U4725 ( .IN1(n3848), .IN2(g339), .QN(n4386) );
  NAND2X0 U4726 ( .IN1(n3973), .IN2(n4387), .QN(n4385) );
  INVX0 U4727 ( .INP(n4220), .ZN(n4387) );
  NOR2X0 U4728 ( .IN1(n4388), .IN2(n4389), .QN(n4220) );
  NOR2X0 U4729 ( .IN1(n1239), .IN2(n2855), .QN(n4389) );
  NOR2X0 U4730 ( .IN1(n4390), .IN2(n34), .QN(n4388) );
  XOR2X1 U4731 ( .IN1(n1599), .IN2(n4391), .Q(n4390) );
  NOR2X0 U4732 ( .IN1(n1606), .IN2(n4384), .QN(n4391) );
  NAND2X0 U4733 ( .IN1(n4392), .IN2(n1641), .QN(n4384) );
  NOR2X0 U4734 ( .IN1(n1594), .IN2(g466), .QN(n4392) );
  INVX0 U4735 ( .INP(n3848), .ZN(n3973) );
  NAND2X0 U4736 ( .IN1(n1647), .IN2(g750), .QN(n3848) );
  NAND2X0 U4737 ( .IN1(n4393), .IN2(n4394), .QN(g11443) );
  NAND2X0 U4738 ( .IN1(n3817), .IN2(g1275), .QN(n4394) );
  NOR2X0 U4739 ( .IN1(n3806), .IN2(n2941), .QN(n3817) );
  NAND2X0 U4740 ( .IN1(n3806), .IN2(n4270), .QN(n4393) );
  NAND2X0 U4741 ( .IN1(n4395), .IN2(n4396), .QN(n4270) );
  NAND2X0 U4742 ( .IN1(n4269), .IN2(n4252), .QN(n4396) );
  XNOR2X1 U4743 ( .IN1(n2910), .IN2(n4397), .Q(n4269) );
  NOR2X0 U4744 ( .IN1(n4185), .IN2(n2764), .QN(n4397) );
  INVX0 U4745 ( .INP(n4184), .ZN(n4185) );
  NAND2X0 U4746 ( .IN1(n4398), .IN2(n3807), .QN(n4395) );
  INVX0 U4747 ( .INP(n4252), .ZN(n3807) );
  NAND2X0 U4748 ( .IN1(n4399), .IN2(n3801), .QN(n4252) );
  NOR2X0 U4749 ( .IN1(n2687), .IN2(n2686), .QN(n3801) );
  NOR2X0 U4750 ( .IN1(n2688), .IN2(n2685), .QN(n4399) );
  NAND2X0 U4751 ( .IN1(n4400), .IN2(n4401), .QN(n4398) );
  NAND2X0 U4752 ( .IN1(n1864), .IN2(g1280), .QN(n4401) );
  NAND2X0 U4753 ( .IN1(n1862), .IN2(n4402), .QN(n4400) );
  NAND2X0 U4754 ( .IN1(n1864), .IN2(n4403), .QN(n4402) );
  NAND2X0 U4755 ( .IN1(n4404), .IN2(n4405), .QN(n4403) );
  NOR2X0 U4756 ( .IN1(n4406), .IN2(n4407), .QN(n4405) );
  NAND2X0 U4757 ( .IN1(n4408), .IN2(n2808), .QN(n4407) );
  NOR2X0 U4758 ( .IN1(g1292), .IN2(g1296), .QN(n4408) );
  NAND2X0 U4759 ( .IN1(n4409), .IN2(n4410), .QN(n4406) );
  NOR2X0 U4760 ( .IN1(test_so6), .IN2(g1255), .QN(n4410) );
  NOR2X0 U4761 ( .IN1(g1260), .IN2(g1265), .QN(n4409) );
  NOR2X0 U4762 ( .IN1(n4411), .IN2(n4412), .QN(n4404) );
  NAND2X0 U4763 ( .IN1(n4413), .IN2(n2871), .QN(n4412) );
  NOR2X0 U4764 ( .IN1(g1250), .IN2(g1275), .QN(n4413) );
  NAND2X0 U4765 ( .IN1(n4414), .IN2(n2829), .QN(n4411) );
  NOR2X0 U4766 ( .IN1(g1304), .IN2(g1245), .QN(n4414) );
  INVX0 U4767 ( .INP(n3785), .ZN(n3806) );
  NAND2X0 U4768 ( .IN1(n4415), .IN2(n1610), .QN(n3785) );
  NOR2X0 U4769 ( .IN1(n2912), .IN2(n968), .QN(n4415) );
  NOR2X0 U4770 ( .IN1(n4416), .IN2(n4417), .QN(g11393) );
  NOR2X0 U4771 ( .IN1(n4418), .IN2(n4419), .QN(n4416) );
  NOR2X0 U4772 ( .IN1(n1722), .IN2(n4420), .QN(n4419) );
  NOR2X0 U4773 ( .IN1(n3208), .IN2(n3182), .QN(n4420) );
  NOR2X0 U4774 ( .IN1(n4421), .IN2(n4422), .QN(n4418) );
  NAND2X0 U4775 ( .IN1(n3182), .IN2(g981), .QN(n4422) );
  NAND2X0 U4776 ( .IN1(n4423), .IN2(n4424), .QN(n3182) );
  NOR2X0 U4777 ( .IN1(n2881), .IN2(n2880), .QN(n4424) );
  NOR2X0 U4778 ( .IN1(n1722), .IN2(n1720), .QN(n4423) );
  NOR2X0 U4779 ( .IN1(n4417), .IN2(n4425), .QN(g11392) );
  XOR2X1 U4780 ( .IN1(g981), .IN2(n4421), .Q(n4425) );
  NAND2X0 U4781 ( .IN1(n4426), .IN2(g976), .QN(n4421) );
  NOR2X0 U4782 ( .IN1(n4417), .IN2(n4427), .QN(g11391) );
  XOR2X1 U4783 ( .IN1(n2880), .IN2(n4426), .Q(n4427) );
  NOR2X0 U4784 ( .IN1(n4428), .IN2(n4429), .QN(g11380) );
  NOR2X0 U4785 ( .IN1(n4430), .IN2(g471), .QN(n4428) );
  NOR2X0 U4786 ( .IN1(n4431), .IN2(n4429), .QN(g11376) );
  NOR2X0 U4787 ( .IN1(n4432), .IN2(n4433), .QN(n4431) );
  NOR2X0 U4788 ( .IN1(n1646), .IN2(n4430), .QN(n4433) );
  NOR2X0 U4789 ( .IN1(n4434), .IN2(n4344), .QN(n4430) );
  INVX0 U4790 ( .INP(n4435), .ZN(n4434) );
  NOR2X0 U4791 ( .IN1(n4436), .IN2(n4437), .QN(n4432) );
  NAND2X0 U4792 ( .IN1(n4344), .IN2(g461), .QN(n4437) );
  NOR2X0 U4793 ( .IN1(n4429), .IN2(n4438), .QN(g11372) );
  XOR2X1 U4794 ( .IN1(g461), .IN2(n4436), .Q(n4438) );
  NAND2X0 U4795 ( .IN1(n4435), .IN2(g456), .QN(n4436) );
  NOR2X0 U4796 ( .IN1(n4417), .IN2(n4439), .QN(g11349) );
  NAND2X0 U4797 ( .IN1(n4440), .IN2(n4441), .QN(n4439) );
  INVX0 U4798 ( .INP(n4426), .ZN(n4441) );
  NOR2X0 U4799 ( .IN1(n3208), .IN2(n2881), .QN(n4426) );
  NAND2X0 U4800 ( .IN1(n2881), .IN2(n3208), .QN(n4440) );
  NAND2X0 U4801 ( .IN1(n4442), .IN2(n1420), .QN(n3208) );
  NOR2X0 U4802 ( .IN1(n34), .IN2(n4443), .QN(n4442) );
  NOR2X0 U4803 ( .IN1(n4444), .IN2(n4445), .QN(n4443) );
  NAND2X0 U4804 ( .IN1(n4446), .IN2(n4447), .QN(n4445) );
  NOR2X0 U4805 ( .IN1(n4448), .IN2(n4449), .QN(n4447) );
  NAND2X0 U4806 ( .IN1(n4450), .IN2(n4451), .QN(n4449) );
  XOR2X1 U4807 ( .IN1(n2836), .IN2(g401), .Q(n4451) );
  XOR2X1 U4808 ( .IN1(n2832), .IN2(g396), .Q(n4450) );
  XOR2X1 U4809 ( .IN1(n2835), .IN2(n2834), .Q(n4448) );
  NOR2X0 U4810 ( .IN1(n4452), .IN2(n4453), .QN(n4446) );
  XOR2X1 U4811 ( .IN1(n2858), .IN2(n2857), .Q(n4453) );
  XOR2X1 U4812 ( .IN1(n2856), .IN2(n2855), .Q(n4452) );
  NAND2X0 U4813 ( .IN1(n4454), .IN2(n4455), .QN(n4444) );
  NOR2X0 U4814 ( .IN1(n4456), .IN2(n4457), .QN(n4455) );
  NAND2X0 U4815 ( .IN1(n4458), .IN2(n4459), .QN(n4457) );
  XOR2X1 U4816 ( .IN1(n2638), .IN2(g416), .Q(n4459) );
  XNOR2X1 U4817 ( .IN1(n1681), .IN2(n4460), .Q(n4458) );
  XOR2X1 U4818 ( .IN1(n2804), .IN2(n2637), .Q(n4456) );
  NOR2X0 U4819 ( .IN1(n4461), .IN2(n4462), .QN(n4454) );
  XOR2X1 U4820 ( .IN1(n2876), .IN2(n2875), .Q(n4462) );
  XOR2X1 U4821 ( .IN1(n2874), .IN2(n2873), .Q(n4461) );
  NAND2X0 U4822 ( .IN1(n4463), .IN2(g109), .QN(n4417) );
  NAND2X0 U4823 ( .IN1(n4464), .IN2(n5214), .QN(n4463) );
  NOR2X0 U4824 ( .IN1(n2683), .IN2(n4465), .QN(n4464) );
  INVX0 U4825 ( .INP(n3197), .ZN(n4465) );
  NOR2X0 U4826 ( .IN1(n4429), .IN2(n4466), .QN(g11340) );
  XOR2X1 U4827 ( .IN1(n1641), .IN2(n4435), .Q(n4466) );
  NOR2X0 U4828 ( .IN1(n4467), .IN2(n34), .QN(n4435) );
  NOR2X0 U4829 ( .IN1(n4344), .IN2(n1606), .QN(n4467) );
  NAND2X0 U4830 ( .IN1(n4468), .IN2(g461), .QN(n4344) );
  NOR2X0 U4831 ( .IN1(n1646), .IN2(n1641), .QN(n4468) );
  NAND2X0 U4832 ( .IN1(g109), .IN2(DFF_441_n1), .QN(n4429) );
  NAND2X0 U4833 ( .IN1(n4469), .IN2(n4470), .QN(g11338) );
  NAND2X0 U4834 ( .IN1(n34), .IN2(g476), .QN(n4470) );
  NAND2X0 U4835 ( .IN1(n1239), .IN2(g516), .QN(n4469) );
  NAND2X0 U4836 ( .IN1(n4471), .IN2(n4472), .QN(g11337) );
  NAND2X0 U4837 ( .IN1(n34), .IN2(g516), .QN(n4472) );
  NAND2X0 U4838 ( .IN1(n1239), .IN2(g511), .QN(n4471) );
  NAND2X0 U4839 ( .IN1(n4473), .IN2(n4474), .QN(g11336) );
  NAND2X0 U4840 ( .IN1(n34), .IN2(g511), .QN(n4474) );
  NAND2X0 U4841 ( .IN1(n1239), .IN2(g506), .QN(n4473) );
  NAND2X0 U4842 ( .IN1(n4475), .IN2(n4476), .QN(g11335) );
  NAND2X0 U4843 ( .IN1(n34), .IN2(g506), .QN(n4476) );
  NAND2X0 U4844 ( .IN1(n1239), .IN2(g501), .QN(n4475) );
  NAND2X0 U4845 ( .IN1(n4477), .IN2(n4478), .QN(g11334) );
  NAND2X0 U4846 ( .IN1(n34), .IN2(g501), .QN(n4478) );
  NAND2X0 U4847 ( .IN1(n1239), .IN2(g496), .QN(n4477) );
  NAND2X0 U4848 ( .IN1(n4479), .IN2(n4480), .QN(g11333) );
  NAND2X0 U4849 ( .IN1(n34), .IN2(g496), .QN(n4480) );
  NAND2X0 U4850 ( .IN1(n1239), .IN2(g491), .QN(n4479) );
  NAND2X0 U4851 ( .IN1(n4481), .IN2(n4482), .QN(g11332) );
  NAND2X0 U4852 ( .IN1(n34), .IN2(g491), .QN(n4482) );
  NAND2X0 U4853 ( .IN1(n1239), .IN2(g486), .QN(n4481) );
  NAND2X0 U4854 ( .IN1(n4483), .IN2(n4484), .QN(g11331) );
  NAND2X0 U4855 ( .IN1(n34), .IN2(g486), .QN(n4484) );
  NAND2X0 U4856 ( .IN1(n1239), .IN2(g481), .QN(n4483) );
  NAND2X0 U4857 ( .IN1(n4485), .IN2(n4486), .QN(g11330) );
  NAND2X0 U4858 ( .IN1(n34), .IN2(g521), .QN(n4486) );
  NAND2X0 U4859 ( .IN1(n1239), .IN2(g525), .QN(n4485) );
  NAND2X0 U4860 ( .IN1(n4487), .IN2(n4488), .QN(g11329) );
  NAND2X0 U4861 ( .IN1(n34), .IN2(g525), .QN(n4488) );
  NAND2X0 U4862 ( .IN1(n1239), .IN2(g530), .QN(n4487) );
  NAND2X0 U4863 ( .IN1(n4489), .IN2(n4490), .QN(g11328) );
  NAND2X0 U4864 ( .IN1(n34), .IN2(g530), .QN(n4490) );
  NAND2X0 U4865 ( .IN1(n1239), .IN2(g534), .QN(n4489) );
  NAND2X0 U4866 ( .IN1(n4491), .IN2(n4492), .QN(g11327) );
  NAND2X0 U4867 ( .IN1(n34), .IN2(g534), .QN(n4492) );
  NAND2X0 U4868 ( .IN1(n1239), .IN2(g538), .QN(n4491) );
  NAND2X0 U4869 ( .IN1(n4493), .IN2(n4494), .QN(g11326) );
  NAND2X0 U4870 ( .IN1(n34), .IN2(g538), .QN(n4494) );
  NAND2X0 U4871 ( .IN1(n1239), .IN2(g542), .QN(n4493) );
  NAND2X0 U4872 ( .IN1(n4495), .IN2(n4496), .QN(g11325) );
  NAND2X0 U4873 ( .IN1(n34), .IN2(g542), .QN(n4496) );
  NAND2X0 U4874 ( .IN1(n1239), .IN2(g476), .QN(n4495) );
  NAND2X0 U4875 ( .IN1(n4497), .IN2(n4498), .QN(g11324) );
  NAND2X0 U4876 ( .IN1(n34), .IN2(g481), .QN(n4498) );
  NAND2X0 U4877 ( .IN1(n4212), .IN2(n1239), .QN(n4497) );
  NAND2X0 U4878 ( .IN1(n4499), .IN2(n4500), .QN(n4212) );
  NAND2X0 U4879 ( .IN1(n1695), .IN2(g521), .QN(n4500) );
  NAND2X0 U4880 ( .IN1(n1698), .IN2(n4501), .QN(n4499) );
  NAND2X0 U4881 ( .IN1(n1695), .IN2(n4502), .QN(n4501) );
  NAND2X0 U4882 ( .IN1(n4503), .IN2(n4504), .QN(n4502) );
  NOR2X0 U4883 ( .IN1(n4505), .IN2(n4506), .QN(n4504) );
  NAND2X0 U4884 ( .IN1(n4507), .IN2(n1689), .QN(n4506) );
  NOR2X0 U4885 ( .IN1(g511), .IN2(g481), .QN(n4507) );
  NAND2X0 U4886 ( .IN1(n4508), .IN2(n4509), .QN(n4505) );
  NOR2X0 U4887 ( .IN1(g476), .IN2(g506), .QN(n4509) );
  NOR2X0 U4888 ( .IN1(g516), .IN2(g486), .QN(n4508) );
  NOR2X0 U4889 ( .IN1(n4510), .IN2(n4511), .QN(n4503) );
  NAND2X0 U4890 ( .IN1(n4512), .IN2(n2865), .QN(n4511) );
  NOR2X0 U4891 ( .IN1(g534), .IN2(g538), .QN(n4512) );
  NAND2X0 U4892 ( .IN1(n4513), .IN2(n2862), .QN(n4510) );
  NOR2X0 U4893 ( .IN1(g501), .IN2(g491), .QN(n4513) );
  NOR2X0 U4894 ( .IN1(n4514), .IN2(n4515), .QN(g11320) );
  NAND2X0 U4895 ( .IN1(n4516), .IN2(n4517), .QN(n4515) );
  NAND2X0 U4896 ( .IN1(n2789), .IN2(n4518), .QN(n4516) );
  NAND2X0 U4897 ( .IN1(n4519), .IN2(n4520), .QN(g11314) );
  NAND2X0 U4898 ( .IN1(n1855), .IN2(g861), .QN(n4520) );
  NAND2X0 U4899 ( .IN1(n3192), .IN2(g968), .QN(n4519) );
  NAND2X0 U4900 ( .IN1(n4521), .IN2(n4522), .QN(g11312) );
  NAND2X0 U4901 ( .IN1(n1855), .IN2(g857), .QN(n4522) );
  NAND2X0 U4902 ( .IN1(g965), .IN2(n3192), .QN(n4521) );
  NAND2X0 U4903 ( .IN1(n4523), .IN2(n4524), .QN(g11310) );
  NAND2X0 U4904 ( .IN1(n1855), .IN2(g853), .QN(n4524) );
  NAND2X0 U4905 ( .IN1(g962), .IN2(n3192), .QN(n4523) );
  INVX0 U4906 ( .INP(n4525), .ZN(g11308) );
  NOR2X0 U4907 ( .IN1(n4526), .IN2(n4527), .QN(n4525) );
  NOR2X0 U4908 ( .IN1(n3192), .IN2(n2926), .QN(n4527) );
  NOR2X0 U4909 ( .IN1(n1855), .IN2(n2646), .QN(n4526) );
  INVX0 U4910 ( .INP(n4528), .ZN(g11306) );
  NOR2X0 U4911 ( .IN1(n4529), .IN2(n4530), .QN(n4528) );
  NOR2X0 U4912 ( .IN1(n3192), .IN2(n2927), .QN(n4530) );
  NOR2X0 U4913 ( .IN1(n1855), .IN2(n2652), .QN(n4529) );
  NAND2X0 U4914 ( .IN1(n4531), .IN2(n4532), .QN(g11305) );
  NAND2X0 U4915 ( .IN1(n1855), .IN2(g841), .QN(n4532) );
  NAND2X0 U4916 ( .IN1(n3192), .IN2(g953), .QN(n4531) );
  NAND2X0 U4917 ( .IN1(n4533), .IN2(n4534), .QN(g11298) );
  NAND2X0 U4918 ( .IN1(n3192), .IN2(g944), .QN(n4534) );
  INVX0 U4919 ( .INP(n1855), .ZN(n3192) );
  NAND2X0 U4920 ( .IN1(n1855), .IN2(g829), .QN(n4533) );
  NAND2X0 U4921 ( .IN1(n4535), .IN2(n4536), .QN(g11294) );
  NAND2X0 U4922 ( .IN1(n4537), .IN2(n3273), .QN(n4536) );
  NOR2X0 U4923 ( .IN1(n4538), .IN2(n4539), .QN(n4537) );
  NOR2X0 U4924 ( .IN1(g1690), .IN2(n4540), .QN(n4539) );
  NAND2X0 U4925 ( .IN1(n4541), .IN2(n4542), .QN(n4540) );
  NAND2X0 U4926 ( .IN1(n4543), .IN2(n4544), .QN(n4542) );
  NAND2X0 U4927 ( .IN1(g1796), .IN2(g1801), .QN(n4544) );
  NAND2X0 U4928 ( .IN1(g1791), .IN2(g1786), .QN(n4543) );
  NAND2X0 U4929 ( .IN1(n4545), .IN2(n4546), .QN(n4541) );
  NAND2X0 U4930 ( .IN1(g1781), .IN2(g1776), .QN(n4546) );
  NAND2X0 U4931 ( .IN1(test_so5), .IN2(g1766), .QN(n4545) );
  NOR2X0 U4932 ( .IN1(n1653), .IN2(n4547), .QN(n4538) );
  NAND2X0 U4933 ( .IN1(n4548), .IN2(n4549), .QN(n4547) );
  NAND2X0 U4934 ( .IN1(n4550), .IN2(n4551), .QN(n4549) );
  NAND2X0 U4935 ( .IN1(n91), .IN2(n63), .QN(n4551) );
  NAND2X0 U4936 ( .IN1(g10664), .IN2(g10663), .QN(n4550) );
  NAND2X0 U4937 ( .IN1(n4552), .IN2(n4553), .QN(n4548) );
  NAND2X0 U4938 ( .IN1(g10719), .IN2(g10720), .QN(n4553) );
  NAND2X0 U4939 ( .IN1(g10722), .IN2(g10721), .QN(n4552) );
  NOR2X0 U4940 ( .IN1(n4554), .IN2(n4555), .QN(n4535) );
  NOR2X0 U4941 ( .IN1(g1857), .IN2(n4556), .QN(n4555) );
  NAND2X0 U4942 ( .IN1(n926), .IN2(n4557), .QN(n4556) );
  NAND2X0 U4943 ( .IN1(n4558), .IN2(n4559), .QN(n4557) );
  INVX0 U4944 ( .INP(n4560), .ZN(n4559) );
  NAND2X0 U4945 ( .IN1(n3472), .IN2(n3293), .QN(n4560) );
  NOR2X0 U4946 ( .IN1(n3287), .IN2(n3286), .QN(n4558) );
  INVX0 U4947 ( .INP(n817), .ZN(n3286) );
  NAND2X0 U4948 ( .IN1(g1814), .IN2(g1828), .QN(n817) );
  INVX0 U4949 ( .INP(n822), .ZN(n3287) );
  NOR2X0 U4950 ( .IN1(n1682), .IN2(n3910), .QN(n4554) );
  NAND2X0 U4951 ( .IN1(n4561), .IN2(n487), .QN(n3910) );
  INVX0 U4952 ( .INP(n926), .ZN(n487) );
  NAND2X0 U4953 ( .IN1(n4562), .IN2(n4563), .QN(g11293) );
  NAND2X0 U4954 ( .IN1(n4564), .IN2(n4561), .QN(n4563) );
  NAND2X0 U4955 ( .IN1(n3472), .IN2(n4565), .QN(n4564) );
  NAND2X0 U4956 ( .IN1(n4566), .IN2(g1854), .QN(n4565) );
  NAND2X0 U4957 ( .IN1(n4567), .IN2(n4568), .QN(n4566) );
  NOR2X0 U4958 ( .IN1(n4569), .IN2(n4570), .QN(n4568) );
  NOR2X0 U4959 ( .IN1(n4571), .IN2(g1857), .QN(n4570) );
  XNOR2X1 U4960 ( .IN1(n1380), .IN2(n4572), .Q(n4571) );
  NOR2X0 U4961 ( .IN1(n1682), .IN2(n4573), .QN(n4569) );
  XNOR2X1 U4962 ( .IN1(n4572), .IN2(n3293), .Q(n4573) );
  NOR2X0 U4963 ( .IN1(n4574), .IN2(n3198), .QN(n4567) );
  NAND2X0 U4964 ( .IN1(n3937), .IN2(n3044), .QN(n3198) );
  INVX0 U4965 ( .INP(n2933), .ZN(n3937) );
  NAND2X0 U4966 ( .IN1(n4561), .IN2(n4575), .QN(n2933) );
  NAND2X0 U4967 ( .IN1(n1608), .IN2(g1834), .QN(n4575) );
  NOR2X0 U4968 ( .IN1(n4576), .IN2(n4577), .QN(n4574) );
  NAND2X0 U4969 ( .IN1(n1380), .IN2(n822), .QN(n4577) );
  NAND2X0 U4970 ( .IN1(n1605), .IN2(g1822), .QN(n822) );
  NAND2X0 U4971 ( .IN1(n3293), .IN2(n3694), .QN(n4576) );
  NAND2X0 U4972 ( .IN1(n4578), .IN2(n4579), .QN(n3694) );
  NOR2X0 U4973 ( .IN1(n1608), .IN2(g1828), .QN(n4579) );
  INVX0 U4974 ( .INP(n4580), .ZN(n4578) );
  NAND2X0 U4975 ( .IN1(n1655), .IN2(n2867), .QN(n4580) );
  NAND2X0 U4976 ( .IN1(n1608), .IN2(g1822), .QN(n3293) );
  NAND2X0 U4977 ( .IN1(n4581), .IN2(n1608), .QN(n3472) );
  NOR2X0 U4978 ( .IN1(n1605), .IN2(g1822), .QN(n4581) );
  NAND2X0 U4979 ( .IN1(n4582), .IN2(n3273), .QN(n4562) );
  INVX0 U4980 ( .INP(n4561), .ZN(n3273) );
  NAND2X0 U4981 ( .IN1(n4583), .IN2(n4584), .QN(n4561) );
  NOR2X0 U4982 ( .IN1(g1828), .IN2(g1834), .QN(n4584) );
  NOR2X0 U4983 ( .IN1(g1822), .IN2(g1814), .QN(n4583) );
  NAND2X0 U4984 ( .IN1(n4585), .IN2(n4586), .QN(n4582) );
  NAND2X0 U4985 ( .IN1(n4587), .IN2(g1690), .QN(n4586) );
  NAND2X0 U4986 ( .IN1(n1653), .IN2(n2903), .QN(n4585) );
  NOR2X0 U4987 ( .IN1(n4588), .IN2(n4514), .QN(g11292) );
  NOR2X0 U4988 ( .IN1(n4589), .IN2(g382), .QN(n4588) );
  NOR2X0 U4989 ( .IN1(n4590), .IN2(n4514), .QN(g11291) );
  NOR2X0 U4990 ( .IN1(n4591), .IN2(n4592), .QN(n4590) );
  NOR2X0 U4991 ( .IN1(n2788), .IN2(n4589), .QN(n4592) );
  NOR2X0 U4992 ( .IN1(n4518), .IN2(n1385), .QN(n4589) );
  NAND2X0 U4993 ( .IN1(n4593), .IN2(g374), .QN(n1385) );
  NOR2X0 U4994 ( .IN1(n4517), .IN2(n4594), .QN(n4591) );
  NAND2X0 U4995 ( .IN1(n4595), .IN2(g374), .QN(n4594) );
  INVX0 U4996 ( .INP(n4593), .ZN(n4595) );
  NOR2X0 U4997 ( .IN1(n2789), .IN2(n2788), .QN(n4593) );
  NOR2X0 U4998 ( .IN1(n4514), .IN2(n4596), .QN(g11290) );
  XOR2X1 U4999 ( .IN1(g374), .IN2(n4517), .Q(n4596) );
  INVX0 U5000 ( .INP(n4597), .ZN(n4517) );
  NOR2X0 U5001 ( .IN1(n4518), .IN2(n2789), .QN(n4597) );
  NAND2X0 U5002 ( .IN1(n1239), .IN2(n4598), .QN(n4518) );
  NAND2X0 U5003 ( .IN1(n2683), .IN2(g109), .QN(n4514) );
  NAND2X0 U5004 ( .IN1(n4599), .IN2(n4600), .QN(g11270) );
  NAND2X0 U5005 ( .IN1(n34), .IN2(g421), .QN(n4600) );
  NAND2X0 U5006 ( .IN1(n1239), .IN2(g416), .QN(n4599) );
  NAND2X0 U5007 ( .IN1(n4601), .IN2(n4602), .QN(g11269) );
  NAND2X0 U5008 ( .IN1(n34), .IN2(g416), .QN(n4602) );
  NAND2X0 U5009 ( .IN1(n1239), .IN2(g411), .QN(n4601) );
  NAND2X0 U5010 ( .IN1(n4603), .IN2(n4604), .QN(g11268) );
  NAND2X0 U5011 ( .IN1(n34), .IN2(g411), .QN(n4604) );
  NAND2X0 U5012 ( .IN1(n1239), .IN2(g406), .QN(n4603) );
  NAND2X0 U5013 ( .IN1(n4605), .IN2(n4606), .QN(g11267) );
  NAND2X0 U5014 ( .IN1(n34), .IN2(g406), .QN(n4606) );
  NAND2X0 U5015 ( .IN1(n1239), .IN2(g401), .QN(n4605) );
  NAND2X0 U5016 ( .IN1(n4607), .IN2(n4608), .QN(g11266) );
  NAND2X0 U5017 ( .IN1(n34), .IN2(g401), .QN(n4608) );
  NAND2X0 U5018 ( .IN1(n1239), .IN2(g396), .QN(n4607) );
  NAND2X0 U5019 ( .IN1(n4609), .IN2(n4610), .QN(g11265) );
  NAND2X0 U5020 ( .IN1(n34), .IN2(g396), .QN(n4610) );
  NAND2X0 U5021 ( .IN1(n1239), .IN2(g391), .QN(n4609) );
  NAND2X0 U5022 ( .IN1(n4611), .IN2(n4612), .QN(g11264) );
  NAND2X0 U5023 ( .IN1(n34), .IN2(g391), .QN(n4612) );
  NAND2X0 U5024 ( .IN1(n1239), .IN2(g386), .QN(n4611) );
  NAND2X0 U5025 ( .IN1(n4613), .IN2(n4614), .QN(g11263) );
  NAND2X0 U5026 ( .IN1(n34), .IN2(g386), .QN(n4614) );
  NAND2X0 U5027 ( .IN1(n1239), .IN2(g426), .QN(n4613) );
  NAND2X0 U5028 ( .IN1(n4615), .IN2(n4616), .QN(g11262) );
  NAND2X0 U5029 ( .IN1(n34), .IN2(g431), .QN(n4616) );
  NAND2X0 U5030 ( .IN1(n1239), .IN2(g435), .QN(n4615) );
  NAND2X0 U5031 ( .IN1(n4617), .IN2(n4618), .QN(g11261) );
  NAND2X0 U5032 ( .IN1(n34), .IN2(g435), .QN(n4618) );
  NAND2X0 U5033 ( .IN1(n1239), .IN2(g440), .QN(n4617) );
  NAND2X0 U5034 ( .IN1(n4619), .IN2(n4620), .QN(g11260) );
  NAND2X0 U5035 ( .IN1(n34), .IN2(g440), .QN(n4620) );
  NAND2X0 U5036 ( .IN1(n1239), .IN2(g444), .QN(n4619) );
  NAND2X0 U5037 ( .IN1(n4621), .IN2(n4622), .QN(g11259) );
  NAND2X0 U5038 ( .IN1(n34), .IN2(g444), .QN(n4622) );
  NAND2X0 U5039 ( .IN1(n1239), .IN2(g448), .QN(n4621) );
  NAND2X0 U5040 ( .IN1(n4623), .IN2(n4624), .QN(g11258) );
  NAND2X0 U5041 ( .IN1(n34), .IN2(g448), .QN(n4624) );
  NAND2X0 U5042 ( .IN1(n1239), .IN2(g452), .QN(n4623) );
  NAND2X0 U5043 ( .IN1(n4625), .IN2(n4626), .QN(g11257) );
  NAND2X0 U5044 ( .IN1(n34), .IN2(g452), .QN(n4626) );
  NAND2X0 U5045 ( .IN1(n1239), .IN2(g421), .QN(n4625) );
  NAND2X0 U5046 ( .IN1(n4627), .IN2(n4628), .QN(g11256) );
  NAND2X0 U5047 ( .IN1(n34), .IN2(g426), .QN(n4628) );
  INVX0 U5048 ( .INP(n1239), .ZN(n34) );
  NAND2X0 U5049 ( .IN1(n4629), .IN2(n1239), .QN(n4627) );
  NAND2X0 U5050 ( .IN1(n4630), .IN2(n4631), .QN(n1239) );
  NOR2X0 U5051 ( .IN1(n4632), .IN2(n4633), .QN(n4631) );
  NAND2X0 U5052 ( .IN1(n2642), .IN2(n2641), .QN(n4633) );
  NAND2X0 U5053 ( .IN1(n4634), .IN2(n2640), .QN(n4632) );
  NOR2X0 U5054 ( .IN1(n4635), .IN2(g829), .QN(n4634) );
  NOR2X0 U5055 ( .IN1(n4636), .IN2(n4637), .QN(n4635) );
  NAND2X0 U5056 ( .IN1(n4638), .IN2(n4639), .QN(n4637) );
  INVX0 U5057 ( .INP(n4640), .ZN(n4639) );
  NOR2X0 U5058 ( .IN1(n2942), .IN2(n4641), .QN(n4636) );
  NOR2X0 U5059 ( .IN1(n4642), .IN2(n4643), .QN(n4641) );
  NOR2X0 U5060 ( .IN1(n4644), .IN2(n4645), .QN(n4630) );
  NAND2X0 U5061 ( .IN1(n2927), .IN2(n2926), .QN(n4645) );
  NAND2X0 U5062 ( .IN1(n4646), .IN2(n2645), .QN(n4644) );
  NOR2X0 U5063 ( .IN1(g841), .IN2(g857), .QN(n4646) );
  INVX0 U5064 ( .INP(n4460), .ZN(n4629) );
  NAND2X0 U5065 ( .IN1(n4647), .IN2(n4648), .QN(n4460) );
  NAND2X0 U5066 ( .IN1(n1681), .IN2(n4598), .QN(n4648) );
  INVX0 U5067 ( .INP(n1420), .ZN(n4598) );
  NAND2X0 U5068 ( .IN1(n4649), .IN2(n1420), .QN(n4647) );
  NAND2X0 U5069 ( .IN1(n4650), .IN2(n4651), .QN(n4649) );
  NAND2X0 U5070 ( .IN1(g431), .IN2(g435), .QN(n4651) );
  NAND2X0 U5071 ( .IN1(n4652), .IN2(n1878), .QN(n4650) );
  NOR2X0 U5072 ( .IN1(n4653), .IN2(g431), .QN(n4652) );
  NOR2X0 U5073 ( .IN1(n4654), .IN2(n4655), .QN(n4653) );
  NAND2X0 U5074 ( .IN1(n4656), .IN2(n4657), .QN(n4655) );
  NOR2X0 U5075 ( .IN1(g421), .IN2(n4658), .QN(n4657) );
  NAND2X0 U5076 ( .IN1(n2837), .IN2(n2835), .QN(n4658) );
  NOR2X0 U5077 ( .IN1(g391), .IN2(n4659), .QN(n4656) );
  NAND2X0 U5078 ( .IN1(n2873), .IN2(n2858), .QN(n4659) );
  NAND2X0 U5079 ( .IN1(n4660), .IN2(n4661), .QN(n4654) );
  NOR2X0 U5080 ( .IN1(n4662), .IN2(n4663), .QN(n4661) );
  NAND2X0 U5081 ( .IN1(n2812), .IN2(n2811), .QN(n4663) );
  NAND2X0 U5082 ( .IN1(n2804), .IN2(n2810), .QN(n4662) );
  NOR2X0 U5083 ( .IN1(g396), .IN2(n4664), .QN(n4660) );
  NAND2X0 U5084 ( .IN1(n2814), .IN2(n2813), .QN(n4664) );
  NOR2X0 U5085 ( .IN1(n4665), .IN2(n4666), .QN(g11206) );
  XOR2X1 U5086 ( .IN1(n4667), .IN2(n4665), .Q(g11163) );
  NAND2X0 U5087 ( .IN1(n4668), .IN2(n4669), .QN(n4665) );
  NAND2X0 U5088 ( .IN1(n4670), .IN2(g109), .QN(n4669) );
  NAND2X0 U5089 ( .IN1(n4671), .IN2(n4672), .QN(n4670) );
  NOR2X0 U5090 ( .IN1(n4673), .IN2(n4674), .QN(n4672) );
  NOR2X0 U5091 ( .IN1(n5217), .IN2(n4638), .QN(n4674) );
  NOR2X0 U5092 ( .IN1(n4675), .IN2(n3211), .QN(n4673) );
  NAND2X0 U5093 ( .IN1(n5216), .IN2(g3069), .QN(n3211) );
  NOR2X0 U5094 ( .IN1(n4676), .IN2(n4677), .QN(n4671) );
  NOR2X0 U5095 ( .IN1(n5218), .IN2(n4678), .QN(n4677) );
  NOR2X0 U5096 ( .IN1(n4318), .IN2(g105), .QN(n4676) );
  NAND2X0 U5097 ( .IN1(g5392), .IN2(g10663), .QN(n4668) );
  NOR2X0 U5098 ( .IN1(n4157), .IN2(n2942), .QN(g5392) );
  NAND2X0 U5099 ( .IN1(g1765), .IN2(g1610), .QN(n4157) );
  NAND2X0 U5100 ( .IN1(n4679), .IN2(n4680), .QN(g10936) );
  NAND2X0 U5101 ( .IN1(n1054), .IN2(g1811), .QN(n4680) );
  NAND2X0 U5102 ( .IN1(n1391), .IN2(n364), .QN(n4679) );
  INVX0 U5103 ( .INP(n1054), .ZN(n364) );
  NAND2X0 U5104 ( .IN1(g1696), .IN2(n2916), .QN(n1054) );
  NAND2X0 U5105 ( .IN1(n4681), .IN2(n4682), .QN(n1391) );
  INVX0 U5106 ( .INP(n4683), .ZN(n4682) );
  NAND2X0 U5107 ( .IN1(n4684), .IN2(n4317), .QN(n4683) );
  NOR2X0 U5108 ( .IN1(n4643), .IN2(n4638), .QN(n4681) );
  NAND2X0 U5109 ( .IN1(n4685), .IN2(n4686), .QN(g10898) );
  NAND2X0 U5110 ( .IN1(n968), .IN2(g105), .QN(n4686) );
  NAND2X0 U5111 ( .IN1(n4687), .IN2(n3546), .QN(n4685) );
  NAND2X0 U5112 ( .IN1(n4688), .IN2(n4184), .QN(n4687) );
  NAND2X0 U5113 ( .IN1(n4317), .IN2(n4689), .QN(n4184) );
  NAND2X0 U5114 ( .IN1(n4690), .IN2(n3231), .QN(n4317) );
  NOR2X0 U5115 ( .IN1(n3228), .IN2(n3229), .QN(n3231) );
  NAND2X0 U5116 ( .IN1(n4691), .IN2(n4692), .QN(n3228) );
  NOR2X0 U5117 ( .IN1(g48), .IN2(g45), .QN(n4692) );
  NOR2X0 U5118 ( .IN1(g46), .IN2(n4693), .QN(n4690) );
  XOR2X1 U5119 ( .IN1(n4694), .IN2(n4695), .Q(n4688) );
  XOR2X1 U5120 ( .IN1(n4696), .IN2(n4697), .Q(n4695) );
  XOR2X1 U5121 ( .IN1(n4698), .IN2(n4699), .Q(n4697) );
  XNOR2X1 U5122 ( .IN1(g1023), .IN2(n1871), .Q(n4699) );
  XNOR2X1 U5123 ( .IN1(g1011), .IN2(n2791), .Q(n4698) );
  XOR2X1 U5124 ( .IN1(n4700), .IN2(n4701), .Q(n4696) );
  XOR2X1 U5125 ( .IN1(n2872), .IN2(n2870), .Q(n4701) );
  XNOR2X1 U5126 ( .IN1(test_so2), .IN2(g1027), .Q(n4700) );
  XNOR2X1 U5127 ( .IN1(n2792), .IN2(test_so8), .Q(n4694) );
  NAND2X0 U5128 ( .IN1(n4702), .IN2(n4703), .QN(g10866) );
  NAND2X0 U5129 ( .IN1(n968), .IN2(g1684), .QN(n4703) );
  NAND2X0 U5130 ( .IN1(n4704), .IN2(n4705), .QN(g10865) );
  NAND2X0 U5131 ( .IN1(n4045), .IN2(g1669), .QN(n4705) );
  NAND2X0 U5132 ( .IN1(n4706), .IN2(n4044), .QN(n4704) );
  NOR2X0 U5133 ( .IN1(n4707), .IN2(n4708), .QN(n4706) );
  NOR2X0 U5134 ( .IN1(n2939), .IN2(g10722), .QN(n4707) );
  NAND2X0 U5135 ( .IN1(n4709), .IN2(n4710), .QN(g10864) );
  NAND2X0 U5136 ( .IN1(n968), .IN2(g1681), .QN(n4710) );
  NAND2X0 U5137 ( .IN1(n4711), .IN2(n4712), .QN(g10863) );
  NAND2X0 U5138 ( .IN1(n4045), .IN2(g1666), .QN(n4712) );
  NAND2X0 U5139 ( .IN1(n4713), .IN2(n4044), .QN(n4711) );
  NOR2X0 U5140 ( .IN1(n4714), .IN2(n4715), .QN(n4713) );
  NOR2X0 U5141 ( .IN1(n4640), .IN2(g1718), .QN(n4715) );
  NAND2X0 U5142 ( .IN1(n4716), .IN2(n4717), .QN(g10862) );
  NAND2X0 U5143 ( .IN1(n968), .IN2(g1678), .QN(n4717) );
  NAND2X0 U5144 ( .IN1(n4718), .IN2(n4719), .QN(g10861) );
  NAND2X0 U5145 ( .IN1(n4045), .IN2(g1663), .QN(n4719) );
  NAND2X0 U5146 ( .IN1(n4044), .IN2(n4720), .QN(n4718) );
  NAND2X0 U5147 ( .IN1(n4721), .IN2(n4722), .QN(g10860) );
  NAND2X0 U5148 ( .IN1(n968), .IN2(g1675), .QN(n4722) );
  NAND2X0 U5149 ( .IN1(n4723), .IN2(n4724), .QN(g10859) );
  NAND2X0 U5150 ( .IN1(n4045), .IN2(g1660), .QN(n4724) );
  NAND2X0 U5151 ( .IN1(n4044), .IN2(n4725), .QN(n4723) );
  NAND2X0 U5152 ( .IN1(n4726), .IN2(n4727), .QN(g10858) );
  NAND2X0 U5153 ( .IN1(n968), .IN2(g1672), .QN(n4727) );
  NAND2X0 U5154 ( .IN1(n4728), .IN2(n4729), .QN(g10855) );
  NAND2X0 U5155 ( .IN1(n968), .IN2(g549), .QN(n4729) );
  NAND2X0 U5156 ( .IN1(n4720), .IN2(n3546), .QN(n4728) );
  NAND2X0 U5157 ( .IN1(n4730), .IN2(n1611), .QN(n4720) );
  NOR2X0 U5158 ( .IN1(n4731), .IN2(n4732), .QN(n4730) );
  INVX0 U5159 ( .INP(n4733), .ZN(n4732) );
  NAND2X0 U5160 ( .IN1(n4714), .IN2(n3764), .QN(n4733) );
  NAND2X0 U5161 ( .IN1(n4734), .IN2(n4063), .QN(n3764) );
  NAND2X0 U5162 ( .IN1(g18), .IN2(g192), .QN(n4063) );
  NAND2X0 U5163 ( .IN1(n3199), .IN2(g1512), .QN(n4734) );
  NOR2X0 U5164 ( .IN1(n4714), .IN2(n4735), .QN(n4731) );
  NAND2X0 U5165 ( .IN1(g109), .IN2(g10720), .QN(n4735) );
  NAND2X0 U5166 ( .IN1(n2934), .IN2(n4667), .QN(g10801) );
  INVX0 U5167 ( .INP(n2928), .ZN(n4667) );
  XOR2X1 U5168 ( .IN1(n4736), .IN2(n4737), .Q(n2928) );
  XOR2X1 U5169 ( .IN1(n4738), .IN2(n4739), .Q(n4737) );
  NAND2X0 U5170 ( .IN1(n5219), .IN2(n4740), .QN(n4739) );
  NAND2X0 U5171 ( .IN1(n4741), .IN2(n4642), .QN(n4738) );
  NAND2X0 U5172 ( .IN1(n4742), .IN2(n4689), .QN(n4642) );
  NOR2X0 U5173 ( .IN1(n91), .IN2(g10664), .QN(n4742) );
  NOR2X0 U5174 ( .IN1(n4743), .IN2(n4744), .QN(n4741) );
  NOR2X0 U5175 ( .IN1(g10664), .IN2(n4745), .QN(n4744) );
  NAND2X0 U5176 ( .IN1(g10663), .IN2(n91), .QN(n4745) );
  NOR2X0 U5177 ( .IN1(n4678), .IN2(n4746), .QN(n4743) );
  XOR2X1 U5178 ( .IN1(g10663), .IN2(n4318), .Q(n4746) );
  XNOR2X1 U5179 ( .IN1(n4747), .IN2(n1858), .Q(n4736) );
  XNOR2X1 U5180 ( .IN1(g10722), .IN2(g10721), .Q(n1858) );
  NAND2X0 U5181 ( .IN1(n4748), .IN2(n4643), .QN(n4747) );
  NAND2X0 U5182 ( .IN1(n4749), .IN2(n4587), .QN(n4643) );
  NOR2X0 U5183 ( .IN1(n63), .IN2(g10720), .QN(n4749) );
  NOR2X0 U5184 ( .IN1(n4750), .IN2(n4751), .QN(n4748) );
  NOR2X0 U5185 ( .IN1(g10720), .IN2(n4752), .QN(n4751) );
  NAND2X0 U5186 ( .IN1(g10719), .IN2(n63), .QN(n4752) );
  NOR2X0 U5187 ( .IN1(n4753), .IN2(n4754), .QN(n4750) );
  XOR2X1 U5188 ( .IN1(n63), .IN2(n4587), .Q(n4754) );
  INVX0 U5189 ( .INP(n4675), .ZN(n63) );
  NAND2X0 U5190 ( .IN1(n4755), .IN2(n4756), .QN(g10800) );
  NAND2X0 U5191 ( .IN1(n968), .IN2(g575), .QN(n4756) );
  NAND2X0 U5192 ( .IN1(n4725), .IN2(n3546), .QN(n4755) );
  NAND2X0 U5193 ( .IN1(n4757), .IN2(n1611), .QN(n4725) );
  NOR2X0 U5194 ( .IN1(n4758), .IN2(n4759), .QN(n4757) );
  INVX0 U5195 ( .INP(n4760), .ZN(n4759) );
  NAND2X0 U5196 ( .IN1(n4714), .IN2(n3759), .QN(n4760) );
  NAND2X0 U5197 ( .IN1(n4761), .IN2(n4065), .QN(n3759) );
  NAND2X0 U5198 ( .IN1(g18), .IN2(g248), .QN(n4065) );
  NAND2X0 U5199 ( .IN1(n3199), .IN2(g1636), .QN(n4761) );
  NOR2X0 U5200 ( .IN1(n4714), .IN2(n4762), .QN(n4758) );
  NOR2X0 U5201 ( .IN1(n2940), .IN2(g10719), .QN(n4762) );
  NAND2X0 U5202 ( .IN1(n4763), .IN2(n4764), .QN(g10799) );
  NAND2X0 U5203 ( .IN1(n968), .IN2(g566), .QN(n4764) );
  NAND2X0 U5204 ( .IN1(n4702), .IN2(n4765), .QN(g10798) );
  NAND2X0 U5205 ( .IN1(n968), .IN2(g563), .QN(n4765) );
  NAND2X0 U5206 ( .IN1(n4766), .IN2(n3546), .QN(n4702) );
  NAND2X0 U5207 ( .IN1(n4767), .IN2(n4768), .QN(n4766) );
  NAND2X0 U5208 ( .IN1(n4714), .IN2(n3762), .QN(n4768) );
  NAND2X0 U5209 ( .IN1(n3572), .IN2(n4769), .QN(n3762) );
  NAND2X0 U5210 ( .IN1(n3199), .IN2(g1624), .QN(n4769) );
  NAND2X0 U5211 ( .IN1(g18), .IN2(g225), .QN(n3572) );
  NAND2X0 U5212 ( .IN1(n1404), .IN2(n4572), .QN(n4767) );
  NAND2X0 U5213 ( .IN1(n4709), .IN2(n4770), .QN(g10797) );
  NAND2X0 U5214 ( .IN1(n968), .IN2(g560), .QN(n4770) );
  NAND2X0 U5215 ( .IN1(n4771), .IN2(n3546), .QN(n4709) );
  NAND2X0 U5216 ( .IN1(n4772), .IN2(n4773), .QN(n4771) );
  NAND2X0 U5217 ( .IN1(n4714), .IN2(n3757), .QN(n4773) );
  NAND2X0 U5218 ( .IN1(n3558), .IN2(n4774), .QN(n3757) );
  NAND2X0 U5219 ( .IN1(n3199), .IN2(g1621), .QN(n4774) );
  NAND2X0 U5220 ( .IN1(g18), .IN2(g219), .QN(n3558) );
  NAND2X0 U5221 ( .IN1(n1404), .IN2(n4775), .QN(n4772) );
  NAND2X0 U5222 ( .IN1(n4716), .IN2(n4776), .QN(g10795) );
  NAND2X0 U5223 ( .IN1(n968), .IN2(g557), .QN(n4776) );
  NAND2X0 U5224 ( .IN1(n4777), .IN2(n3546), .QN(n4716) );
  NAND2X0 U5225 ( .IN1(n4778), .IN2(n4779), .QN(n4777) );
  NAND2X0 U5226 ( .IN1(n4714), .IN2(n3749), .QN(n4779) );
  NAND2X0 U5227 ( .IN1(n3614), .IN2(n4780), .QN(n3749) );
  NAND2X0 U5228 ( .IN1(n3199), .IN2(g1615), .QN(n4780) );
  NAND2X0 U5229 ( .IN1(g18), .IN2(g213), .QN(n3614) );
  NAND2X0 U5230 ( .IN1(n1404), .IN2(n4640), .QN(n4778) );
  NAND2X0 U5231 ( .IN1(n4721), .IN2(n4781), .QN(g10793) );
  NAND2X0 U5232 ( .IN1(n968), .IN2(g554), .QN(n4781) );
  NAND2X0 U5233 ( .IN1(n4782), .IN2(n4783), .QN(n4721) );
  INVX0 U5234 ( .INP(n4784), .ZN(n4783) );
  NOR2X0 U5235 ( .IN1(n4785), .IN2(n3745), .QN(n4784) );
  NAND2X0 U5236 ( .IN1(n3602), .IN2(n4786), .QN(n3745) );
  NAND2X0 U5237 ( .IN1(n3199), .IN2(g1639), .QN(n4786) );
  NAND2X0 U5238 ( .IN1(g18), .IN2(g207), .QN(n3602) );
  NOR2X0 U5239 ( .IN1(n968), .IN2(n4787), .QN(n4782) );
  NOR2X0 U5240 ( .IN1(n4708), .IN2(n4788), .QN(n4787) );
  NAND2X0 U5241 ( .IN1(n4753), .IN2(g109), .QN(n4788) );
  NAND2X0 U5242 ( .IN1(n4726), .IN2(n4789), .QN(g10791) );
  NAND2X0 U5243 ( .IN1(n968), .IN2(g546), .QN(n4789) );
  NAND2X0 U5244 ( .IN1(n4790), .IN2(n3546), .QN(n4726) );
  NAND2X0 U5245 ( .IN1(n4791), .IN2(n4792), .QN(n4790) );
  NAND2X0 U5246 ( .IN1(n4793), .IN2(n1404), .QN(n4792) );
  NAND2X0 U5247 ( .IN1(n4714), .IN2(n3766), .QN(n4791) );
  NAND2X0 U5248 ( .IN1(n3587), .IN2(n4794), .QN(n3766) );
  NAND2X0 U5249 ( .IN1(n3199), .IN2(g1618), .QN(n4794) );
  NAND2X0 U5250 ( .IN1(g18), .IN2(g186), .QN(n3587) );
  NAND2X0 U5251 ( .IN1(n4763), .IN2(n4795), .QN(g10776) );
  NAND2X0 U5252 ( .IN1(n968), .IN2(g1687), .QN(n4795) );
  NAND2X0 U5253 ( .IN1(n4796), .IN2(n3546), .QN(n4763) );
  NAND2X0 U5254 ( .IN1(n4797), .IN2(n4798), .QN(n4796) );
  NAND2X0 U5255 ( .IN1(n1404), .IN2(n91), .QN(n4798) );
  NOR2X0 U5256 ( .IN1(n1450), .IN2(n4799), .QN(n4797) );
  NOR2X0 U5257 ( .IN1(n3768), .IN2(n4785), .QN(n4799) );
  NAND2X0 U5258 ( .IN1(n4800), .IN2(n4801), .QN(n3768) );
  NAND2X0 U5259 ( .IN1(n2755), .IN2(n3199), .QN(n4801) );
  NAND2X0 U5260 ( .IN1(g18), .IN2(n2849), .QN(n4800) );
  NAND2X0 U5261 ( .IN1(n4802), .IN2(n4803), .QN(g10773) );
  NAND2X0 U5262 ( .IN1(n4150), .IN2(n4640), .QN(n4803) );
  NAND2X0 U5263 ( .IN1(n4804), .IN2(g1727), .QN(n4802) );
  NAND2X0 U5264 ( .IN1(n4805), .IN2(n4806), .QN(g10771) );
  NAND2X0 U5265 ( .IN1(n4804), .IN2(g1724), .QN(n4806) );
  NAND2X0 U5266 ( .IN1(n4807), .IN2(n4150), .QN(n4805) );
  NOR2X0 U5267 ( .IN1(n4753), .IN2(n2939), .QN(n4807) );
  NAND2X0 U5268 ( .IN1(n4808), .IN2(n4809), .QN(g10770) );
  NAND2X0 U5269 ( .IN1(n4804), .IN2(g1721), .QN(n4809) );
  NAND2X0 U5270 ( .IN1(n4793), .IN2(n4150), .QN(n4808) );
  NOR2X0 U5271 ( .IN1(n4587), .IN2(n2940), .QN(n4793) );
  NAND2X0 U5272 ( .IN1(n4810), .IN2(n4811), .QN(g10767) );
  NAND2X0 U5273 ( .IN1(n4045), .IN2(g1657), .QN(n4811) );
  NAND2X0 U5274 ( .IN1(n4044), .IN2(n4812), .QN(n4810) );
  NAND2X0 U5275 ( .IN1(n4813), .IN2(n4814), .QN(g10765) );
  NAND2X0 U5276 ( .IN1(n4045), .IN2(g1654), .QN(n4814) );
  INVX0 U5277 ( .INP(n4044), .ZN(n4045) );
  NAND2X0 U5278 ( .IN1(n4044), .IN2(n4815), .QN(n4813) );
  NOR2X0 U5279 ( .IN1(g1696), .IN2(n2916), .QN(n4044) );
  NAND2X0 U5280 ( .IN1(n4816), .IN2(n4817), .QN(g10718) );
  NAND2X0 U5281 ( .IN1(n968), .IN2(g572), .QN(n4817) );
  NAND2X0 U5282 ( .IN1(n4812), .IN2(n3546), .QN(n4816) );
  NAND2X0 U5283 ( .IN1(n4818), .IN2(n1611), .QN(n4812) );
  NOR2X0 U5284 ( .IN1(n4819), .IN2(n4820), .QN(n4818) );
  INVX0 U5285 ( .INP(n4821), .ZN(n4820) );
  NAND2X0 U5286 ( .IN1(n4714), .IN2(n3751), .QN(n4821) );
  NAND2X0 U5287 ( .IN1(n4822), .IN2(n4067), .QN(n3751) );
  NAND2X0 U5288 ( .IN1(g18), .IN2(g243), .QN(n4067) );
  NAND2X0 U5289 ( .IN1(n3199), .IN2(g1633), .QN(n4822) );
  NOR2X0 U5290 ( .IN1(n4714), .IN2(n4823), .QN(n4819) );
  NAND2X0 U5291 ( .IN1(g109), .IN2(g10664), .QN(n4823) );
  INVX0 U5292 ( .INP(n4785), .ZN(n4714) );
  NAND2X0 U5293 ( .IN1(n4824), .IN2(n4825), .QN(g10717) );
  NAND2X0 U5294 ( .IN1(n968), .IN2(g569), .QN(n4825) );
  NAND2X0 U5295 ( .IN1(n4815), .IN2(n3546), .QN(n4824) );
  INVX0 U5296 ( .INP(n968), .ZN(n3546) );
  NAND2X0 U5297 ( .IN1(n2916), .IN2(n4826), .QN(n968) );
  NAND2X0 U5298 ( .IN1(n4827), .IN2(n4828), .QN(n4815) );
  NAND2X0 U5299 ( .IN1(n1404), .IN2(g10663), .QN(n4828) );
  INVX0 U5300 ( .INP(n4708), .ZN(n1404) );
  NAND2X0 U5301 ( .IN1(n1611), .IN2(n4785), .QN(n4708) );
  NOR2X0 U5302 ( .IN1(n1450), .IN2(n4829), .QN(n4827) );
  NOR2X0 U5303 ( .IN1(n3770), .IN2(n4785), .QN(n4829) );
  NAND2X0 U5304 ( .IN1(n5229), .IN2(n1611), .QN(n4785) );
  NAND2X0 U5305 ( .IN1(n4830), .IN2(n4831), .QN(n3770) );
  NAND2X0 U5306 ( .IN1(n2752), .IN2(n3199), .QN(n4831) );
  INVX0 U5307 ( .INP(g18), .ZN(n3199) );
  NAND2X0 U5308 ( .IN1(g18), .IN2(n2850), .QN(n4830) );
  NAND2X0 U5309 ( .IN1(n4832), .IN2(n4833), .QN(g10711) );
  NAND2X0 U5310 ( .IN1(n4804), .IN2(g1733), .QN(n4833) );
  NAND2X0 U5311 ( .IN1(n4150), .IN2(n4572), .QN(n4832) );
  NAND2X0 U5312 ( .IN1(g109), .IN2(n4675), .QN(n4572) );
  NAND2X0 U5313 ( .IN1(n4834), .IN2(n4835), .QN(g10707) );
  NAND2X0 U5314 ( .IN1(n4804), .IN2(g1730), .QN(n4835) );
  INVX0 U5315 ( .INP(n4150), .ZN(n4804) );
  NAND2X0 U5316 ( .IN1(n4150), .IN2(n4775), .QN(n4834) );
  INVX0 U5317 ( .INP(n4638), .ZN(n4775) );
  NOR2X0 U5318 ( .IN1(n4826), .IN2(n2916), .QN(n4150) );
  INVX0 U5319 ( .INP(g1696), .ZN(n4826) );
  INVX0 U5320 ( .INP(n4678), .ZN(g10664) );
  NOR2X0 U5321 ( .IN1(n4836), .IN2(n4837), .QN(n4678) );
  NAND2X0 U5322 ( .IN1(n4838), .IN2(n4839), .QN(n4837) );
  NOR2X0 U5323 ( .IN1(n4840), .IN2(n4841), .QN(n4839) );
  NOR2X0 U5324 ( .IN1(n4842), .IN2(n2937), .QN(n4841) );
  NOR2X0 U5325 ( .IN1(n2713), .IN2(n4843), .QN(n4840) );
  NOR2X0 U5326 ( .IN1(n4844), .IN2(n4845), .QN(n4838) );
  NAND2X0 U5327 ( .IN1(n4846), .IN2(n4847), .QN(n4845) );
  NAND2X0 U5328 ( .IN1(n4848), .IN2(n4849), .QN(n4847) );
  NOR2X0 U5329 ( .IN1(n4850), .IN2(n4851), .QN(n4848) );
  NAND2X0 U5330 ( .IN1(n1478), .IN2(n4852), .QN(n4851) );
  NAND2X0 U5331 ( .IN1(n4853), .IN2(n4854), .QN(n4850) );
  NOR2X0 U5332 ( .IN1(n4855), .IN2(n4856), .QN(n4853) );
  NAND2X0 U5333 ( .IN1(g1191), .IN2(n4857), .QN(n4846) );
  NOR2X0 U5334 ( .IN1(n1633), .IN2(n4858), .QN(n4844) );
  NAND2X0 U5335 ( .IN1(n4859), .IN2(n4860), .QN(n4836) );
  NOR2X0 U5336 ( .IN1(n4861), .IN2(n4862), .QN(n4860) );
  NAND2X0 U5337 ( .IN1(n4863), .IN2(n4864), .QN(n4862) );
  NAND2X0 U5338 ( .IN1(g919), .IN2(n4865), .QN(n4864) );
  NAND2X0 U5339 ( .IN1(n4866), .IN2(g947), .QN(n4863) );
  NOR2X0 U5340 ( .IN1(n2738), .IN2(n4867), .QN(n4861) );
  NOR2X0 U5341 ( .IN1(n4868), .IN2(n4869), .QN(n4859) );
  NOR2X0 U5342 ( .IN1(n2718), .IN2(n4870), .QN(n4869) );
  NOR2X0 U5343 ( .IN1(n5224), .IN2(n4871), .QN(n4868) );
  INVX0 U5344 ( .INP(n4666), .ZN(g10628) );
  NAND2X0 U5345 ( .IN1(n4872), .IN2(n4873), .QN(n4666) );
  NAND2X0 U5346 ( .IN1(n4874), .IN2(g109), .QN(n4873) );
  NAND2X0 U5347 ( .IN1(n4875), .IN2(n4876), .QN(n4874) );
  NOR2X0 U5348 ( .IN1(n4877), .IN2(n4878), .QN(n4876) );
  NOR2X0 U5349 ( .IN1(n5214), .IN2(n4638), .QN(n4878) );
  NAND2X0 U5350 ( .IN1(g10722), .IN2(g109), .QN(n4638) );
  NAND2X0 U5351 ( .IN1(n4879), .IN2(n4880), .QN(g10722) );
  NOR2X0 U5352 ( .IN1(n4881), .IN2(n4882), .QN(n4880) );
  NAND2X0 U5353 ( .IN1(n4883), .IN2(n4884), .QN(n4882) );
  NOR2X0 U5354 ( .IN1(n4885), .IN2(n4886), .QN(n4884) );
  NAND2X0 U5355 ( .IN1(n4887), .IN2(n4888), .QN(n4886) );
  NAND2X0 U5356 ( .IN1(g907), .IN2(n4865), .QN(n4888) );
  NAND2X0 U5357 ( .IN1(n4866), .IN2(g986), .QN(n4887) );
  NOR2X0 U5358 ( .IN1(n2653), .IN2(n4889), .QN(n4885) );
  NOR2X0 U5359 ( .IN1(n4890), .IN2(n4891), .QN(n4883) );
  NOR2X0 U5360 ( .IN1(n4849), .IN2(n4892), .QN(n4891) );
  INVX0 U5361 ( .INP(g1179), .ZN(n4892) );
  NOR2X0 U5362 ( .IN1(n2647), .IN2(n4858), .QN(n4890) );
  NAND2X0 U5363 ( .IN1(n4893), .IN2(n4894), .QN(n4881) );
  NOR2X0 U5364 ( .IN1(n4895), .IN2(n4896), .QN(n4894) );
  NAND2X0 U5365 ( .IN1(n4897), .IN2(n4898), .QN(n4896) );
  NAND2X0 U5366 ( .IN1(n4899), .IN2(n1631), .QN(n4897) );
  NOR2X0 U5367 ( .IN1(n2636), .IN2(n4900), .QN(n4895) );
  NOR2X0 U5368 ( .IN1(n4901), .IN2(n4902), .QN(n4893) );
  NAND2X0 U5369 ( .IN1(n4903), .IN2(n4904), .QN(n4902) );
  NAND2X0 U5370 ( .IN1(n4905), .IN2(g940), .QN(n4904) );
  NAND2X0 U5371 ( .IN1(g895), .IN2(n4906), .QN(n4903) );
  NOR2X0 U5372 ( .IN1(n2646), .IN2(n510), .QN(n4901) );
  NOR2X0 U5373 ( .IN1(n4907), .IN2(n4908), .QN(n4879) );
  NAND2X0 U5374 ( .IN1(n4909), .IN2(n4910), .QN(n4908) );
  NOR2X0 U5375 ( .IN1(n4911), .IN2(n4912), .QN(n4910) );
  NAND2X0 U5376 ( .IN1(n4913), .IN2(n4914), .QN(n4912) );
  NAND2X0 U5377 ( .IN1(n1480), .IN2(g1601), .QN(n4914) );
  NAND2X0 U5378 ( .IN1(g1203), .IN2(n1512), .QN(n4913) );
  NOR2X0 U5379 ( .IN1(n2725), .IN2(n4915), .QN(n4911) );
  NOR2X0 U5380 ( .IN1(n4916), .IN2(n4917), .QN(n4909) );
  NOR2X0 U5381 ( .IN1(n1632), .IN2(n4843), .QN(n4917) );
  NOR2X0 U5382 ( .IN1(n2710), .IN2(n4870), .QN(n4916) );
  NAND2X0 U5383 ( .IN1(n4918), .IN2(n4919), .QN(n4907) );
  NOR2X0 U5384 ( .IN1(n4920), .IN2(n4921), .QN(n4919) );
  NAND2X0 U5385 ( .IN1(n4922), .IN2(n4923), .QN(n4921) );
  INVX0 U5386 ( .INP(n4924), .ZN(n4923) );
  NOR2X0 U5387 ( .IN1(n4842), .IN2(n1721), .QN(n4924) );
  NAND2X0 U5388 ( .IN1(n4925), .IN2(g1753), .QN(n4922) );
  NOR2X0 U5389 ( .IN1(n2730), .IN2(n4867), .QN(n4920) );
  NOR2X0 U5390 ( .IN1(n4926), .IN2(n4927), .QN(n4918) );
  NOR2X0 U5391 ( .IN1(n4871), .IN2(DFF_228_n1), .QN(n4927) );
  NOR2X0 U5392 ( .IN1(n2731), .IN2(n4928), .QN(n4926) );
  NOR2X0 U5393 ( .IN1(n4675), .IN2(n3197), .QN(n4877) );
  NAND2X0 U5394 ( .IN1(n2661), .IN2(g3007), .QN(n3197) );
  NOR2X0 U5395 ( .IN1(n4929), .IN2(n4930), .QN(n4875) );
  NOR2X0 U5396 ( .IN1(n4753), .IN2(n4035), .QN(n4930) );
  INVX0 U5397 ( .INP(g881), .ZN(n4035) );
  NOR2X0 U5398 ( .IN1(n4587), .IN2(n4931), .QN(n4929) );
  INVX0 U5399 ( .INP(g877), .ZN(n4931) );
  NAND2X0 U5400 ( .IN1(n4640), .IN2(n3741), .QN(n4872) );
  INVX0 U5401 ( .INP(n4932), .ZN(n3741) );
  NAND2X0 U5402 ( .IN1(n4933), .IN2(n5215), .QN(n4932) );
  NOR2X0 U5403 ( .IN1(n2662), .IN2(n2941), .QN(n4933) );
  NOR2X0 U5404 ( .IN1(n4684), .IN2(n2942), .QN(n4640) );
  NAND2X0 U5405 ( .IN1(n2934), .IN2(n4318), .QN(g10465) );
  INVX0 U5406 ( .INP(n91), .ZN(n4318) );
  NAND2X0 U5407 ( .IN1(n4934), .IN2(n4935), .QN(n91) );
  NOR2X0 U5408 ( .IN1(n4936), .IN2(n4937), .QN(n4935) );
  NAND2X0 U5409 ( .IN1(n4938), .IN2(n4939), .QN(n4937) );
  NAND2X0 U5410 ( .IN1(n4940), .IN2(g965), .QN(n4939) );
  NOR2X0 U5411 ( .IN1(n4941), .IN2(n4942), .QN(n4938) );
  NOR2X0 U5412 ( .IN1(n2703), .IN2(n4943), .QN(n4942) );
  NOR2X0 U5413 ( .IN1(n2658), .IN2(n4889), .QN(n4941) );
  INVX0 U5414 ( .INP(n4944), .ZN(n4936) );
  NOR2X0 U5415 ( .IN1(n4945), .IN2(n4946), .QN(n4944) );
  NAND2X0 U5416 ( .IN1(n4947), .IN2(n4948), .QN(n4946) );
  NAND2X0 U5417 ( .IN1(g913), .IN2(n4865), .QN(n4948) );
  NAND2X0 U5418 ( .IN1(n4949), .IN2(n4950), .QN(n4945) );
  NAND2X0 U5419 ( .IN1(g1185), .IN2(n4857), .QN(n4950) );
  NAND2X0 U5420 ( .IN1(n4951), .IN2(g278), .QN(n4949) );
  NOR2X0 U5421 ( .IN1(n4952), .IN2(n4953), .QN(n4934) );
  NAND2X0 U5422 ( .IN1(n4954), .IN2(n4955), .QN(n4953) );
  NAND2X0 U5423 ( .IN1(n4956), .IN2(g302), .QN(n4955) );
  NOR2X0 U5424 ( .IN1(n4957), .IN2(n4958), .QN(n4954) );
  NOR2X0 U5425 ( .IN1(n2712), .IN2(n4843), .QN(n4958) );
  NOR2X0 U5426 ( .IN1(n2715), .IN2(n4870), .QN(n4957) );
  NAND2X0 U5427 ( .IN1(n4959), .IN2(n4960), .QN(n4952) );
  NAND2X0 U5428 ( .IN1(n1479), .IN2(g1564), .QN(n4960) );
  NOR2X0 U5429 ( .IN1(n4961), .IN2(n4962), .QN(n4959) );
  NOR2X0 U5430 ( .IN1(n5225), .IN2(n4871), .QN(n4962) );
  NOR2X0 U5431 ( .IN1(n2887), .IN2(n4963), .QN(n4961) );
  NAND2X0 U5432 ( .IN1(n2934), .IN2(n4675), .QN(g10463) );
  NOR2X0 U5433 ( .IN1(n4964), .IN2(n4965), .QN(n4675) );
  NAND2X0 U5434 ( .IN1(n4966), .IN2(n4967), .QN(n4965) );
  NOR2X0 U5435 ( .IN1(n4968), .IN2(n4969), .QN(n4967) );
  NAND2X0 U5436 ( .IN1(n4970), .IN2(n4971), .QN(n4969) );
  NAND2X0 U5437 ( .IN1(n4951), .IN2(g275), .QN(n4971) );
  NAND2X0 U5438 ( .IN1(n4956), .IN2(g299), .QN(n4970) );
  NAND2X0 U5439 ( .IN1(n4972), .IN2(n4973), .QN(n4968) );
  NAND2X0 U5440 ( .IN1(n1485), .IN2(g1580), .QN(n4973) );
  NAND2X0 U5441 ( .IN1(n1486), .IN2(g1537), .QN(n4972) );
  NOR2X0 U5442 ( .IN1(n4974), .IN2(n4975), .QN(n4966) );
  NAND2X0 U5443 ( .IN1(n4976), .IN2(n4977), .QN(n4975) );
  NAND2X0 U5444 ( .IN1(n4925), .IN2(g1756), .QN(n4977) );
  NAND2X0 U5445 ( .IN1(n4740), .IN2(n3034), .QN(n4976) );
  NAND2X0 U5446 ( .IN1(n4978), .IN2(n4979), .QN(n4974) );
  NAND2X0 U5447 ( .IN1(n4899), .IN2(n3057), .QN(n4979) );
  NAND2X0 U5448 ( .IN1(n4980), .IN2(n4981), .QN(n4978) );
  INVX0 U5449 ( .INP(n4982), .ZN(n4980) );
  NAND2X0 U5450 ( .IN1(n4983), .IN2(n4984), .QN(n4964) );
  NOR2X0 U5451 ( .IN1(n4985), .IN2(n4986), .QN(n4984) );
  NAND2X0 U5452 ( .IN1(n4987), .IN2(n4988), .QN(n4986) );
  NAND2X0 U5453 ( .IN1(n4989), .IN2(g1327), .QN(n4988) );
  NAND2X0 U5454 ( .IN1(g1182), .IN2(n4857), .QN(n4987) );
  NAND2X0 U5455 ( .IN1(n4990), .IN2(n4991), .QN(n4985) );
  NAND2X0 U5456 ( .IN1(n4856), .IN2(g1733), .QN(n4991) );
  NAND2X0 U5457 ( .IN1(n1480), .IN2(g1604), .QN(n4990) );
  NOR2X0 U5458 ( .IN1(n4992), .IN2(n4993), .QN(n4983) );
  NAND2X0 U5459 ( .IN1(n4994), .IN2(n4995), .QN(n4993) );
  NAND2X0 U5460 ( .IN1(n4940), .IN2(g962), .QN(n4995) );
  NAND2X0 U5461 ( .IN1(n1479), .IN2(g1561), .QN(n4994) );
  NAND2X0 U5462 ( .IN1(n4996), .IN2(n4997), .QN(n4992) );
  NAND2X0 U5463 ( .IN1(n4998), .IN2(n3025), .QN(n4997) );
  NAND2X0 U5464 ( .IN1(g910), .IN2(n4865), .QN(n4996) );
  NAND2X0 U5465 ( .IN1(n2934), .IN2(n4684), .QN(g10459) );
  INVX0 U5466 ( .INP(g10721), .ZN(n4684) );
  NAND2X0 U5467 ( .IN1(n4999), .IN2(n5000), .QN(g10721) );
  NOR2X0 U5468 ( .IN1(n5001), .IN2(n5002), .QN(n5000) );
  NAND2X0 U5469 ( .IN1(n5003), .IN2(n5004), .QN(n5002) );
  NOR2X0 U5470 ( .IN1(n5005), .IN2(n5006), .QN(n5004) );
  NAND2X0 U5471 ( .IN1(n5007), .IN2(n5008), .QN(n5006) );
  NAND2X0 U5472 ( .IN1(g904), .IN2(n4865), .QN(n5008) );
  NAND2X0 U5473 ( .IN1(n4866), .IN2(g981), .QN(n5007) );
  NOR2X0 U5474 ( .IN1(n2657), .IN2(n4889), .QN(n5005) );
  NOR2X0 U5475 ( .IN1(n5009), .IN2(n5010), .QN(n5003) );
  NOR2X0 U5476 ( .IN1(n4849), .IN2(n5011), .QN(n5010) );
  INVX0 U5477 ( .INP(g1176), .ZN(n5011) );
  NOR2X0 U5478 ( .IN1(n2667), .IN2(n4858), .QN(n5009) );
  NAND2X0 U5479 ( .IN1(n5012), .IN2(n5013), .QN(n5001) );
  NOR2X0 U5480 ( .IN1(n5014), .IN2(n5015), .QN(n5013) );
  NAND2X0 U5481 ( .IN1(n5016), .IN2(n4898), .QN(n5015) );
  NAND2X0 U5482 ( .IN1(n4899), .IN2(g9), .QN(n5016) );
  NOR2X0 U5483 ( .IN1(n2670), .IN2(n4900), .QN(n5014) );
  NOR2X0 U5484 ( .IN1(n5017), .IN2(n5018), .QN(n5012) );
  NAND2X0 U5485 ( .IN1(n5019), .IN2(n5020), .QN(n5018) );
  NAND2X0 U5486 ( .IN1(n4905), .IN2(g936), .QN(n5020) );
  NAND2X0 U5487 ( .IN1(g892), .IN2(n4906), .QN(n5019) );
  NOR2X0 U5488 ( .IN1(n2652), .IN2(n510), .QN(n5017) );
  NOR2X0 U5489 ( .IN1(n5021), .IN2(n5022), .QN(n4999) );
  NAND2X0 U5490 ( .IN1(n5023), .IN2(n5024), .QN(n5022) );
  NOR2X0 U5491 ( .IN1(n5025), .IN2(n5026), .QN(n5024) );
  NAND2X0 U5492 ( .IN1(n5027), .IN2(n5028), .QN(n5026) );
  NAND2X0 U5493 ( .IN1(n1480), .IN2(g1598), .QN(n5028) );
  INVX0 U5494 ( .INP(n4943), .ZN(n1480) );
  NAND2X0 U5495 ( .IN1(n1512), .IN2(g1200), .QN(n5027) );
  NOR2X0 U5496 ( .IN1(n2701), .IN2(n4915), .QN(n5025) );
  NOR2X0 U5497 ( .IN1(n5029), .IN2(n5030), .QN(n5023) );
  NOR2X0 U5498 ( .IN1(n1652), .IN2(n4843), .QN(n5030) );
  NOR2X0 U5499 ( .IN1(n2724), .IN2(n4870), .QN(n5029) );
  NAND2X0 U5500 ( .IN1(n5031), .IN2(n5032), .QN(n5021) );
  NOR2X0 U5501 ( .IN1(n5033), .IN2(n5034), .QN(n5032) );
  NAND2X0 U5502 ( .IN1(n5035), .IN2(n5036), .QN(n5034) );
  NAND2X0 U5503 ( .IN1(n4855), .IN2(g1346), .QN(n5036) );
  NAND2X0 U5504 ( .IN1(n4925), .IN2(g1750), .QN(n5035) );
  NOR2X0 U5505 ( .IN1(n2736), .IN2(n4867), .QN(n5033) );
  NOR2X0 U5506 ( .IN1(n5037), .IN2(n5038), .QN(n5031) );
  NOR2X0 U5507 ( .IN1(n4871), .IN2(DFF_242_n1), .QN(n5038) );
  NOR2X0 U5508 ( .IN1(n2735), .IN2(n4928), .QN(n5037) );
  INVX0 U5509 ( .INP(n4956), .ZN(n4928) );
  NAND2X0 U5510 ( .IN1(n2934), .IN2(n4753), .QN(g10457) );
  INVX0 U5511 ( .INP(g10720), .ZN(n4753) );
  NAND2X0 U5512 ( .IN1(n5039), .IN2(n5040), .QN(g10720) );
  NOR2X0 U5513 ( .IN1(n5041), .IN2(n5042), .QN(n5040) );
  NAND2X0 U5514 ( .IN1(n5043), .IN2(n5044), .QN(n5042) );
  NOR2X0 U5515 ( .IN1(n5045), .IN2(n5046), .QN(n5044) );
  NAND2X0 U5516 ( .IN1(n5047), .IN2(n5048), .QN(n5046) );
  NAND2X0 U5517 ( .IN1(g901), .IN2(n4865), .QN(n5048) );
  NAND2X0 U5518 ( .IN1(n4866), .IN2(g976), .QN(n5047) );
  INVX0 U5519 ( .INP(n5049), .ZN(n4866) );
  NOR2X0 U5520 ( .IN1(n2655), .IN2(n4889), .QN(n5045) );
  NOR2X0 U5521 ( .IN1(n5050), .IN2(n5051), .QN(n5043) );
  NOR2X0 U5522 ( .IN1(n4849), .IN2(n5052), .QN(n5051) );
  INVX0 U5523 ( .INP(g1173), .ZN(n5052) );
  NOR2X0 U5524 ( .IN1(n2665), .IN2(n4858), .QN(n5050) );
  NAND2X0 U5525 ( .IN1(n5053), .IN2(n5054), .QN(n5041) );
  NOR2X0 U5526 ( .IN1(n5055), .IN2(n5056), .QN(n5054) );
  NAND2X0 U5527 ( .IN1(n5057), .IN2(n4898), .QN(n5056) );
  NAND2X0 U5528 ( .IN1(n4899), .IN2(g12), .QN(n5057) );
  NOR2X0 U5529 ( .IN1(n2757), .IN2(n4900), .QN(n5055) );
  NOR2X0 U5530 ( .IN1(n5058), .IN2(n5059), .QN(n5053) );
  NAND2X0 U5531 ( .IN1(n5060), .IN2(n5061), .QN(n5059) );
  NAND2X0 U5532 ( .IN1(n4905), .IN2(g932), .QN(n5061) );
  NAND2X0 U5533 ( .IN1(g889), .IN2(n4906), .QN(n5060) );
  NOR2X0 U5534 ( .IN1(n2648), .IN2(n510), .QN(n5058) );
  NOR2X0 U5535 ( .IN1(n5062), .IN2(n5063), .QN(n5039) );
  NAND2X0 U5536 ( .IN1(n5064), .IN2(n5065), .QN(n5063) );
  NOR2X0 U5537 ( .IN1(n5066), .IN2(n5067), .QN(n5065) );
  NAND2X0 U5538 ( .IN1(n5068), .IN2(n5069), .QN(n5067) );
  NAND2X0 U5539 ( .IN1(g1197), .IN2(n1512), .QN(n5069) );
  NAND2X0 U5540 ( .IN1(n1530), .IN2(g925), .QN(n5068) );
  NOR2X0 U5541 ( .IN1(n2706), .IN2(n4915), .QN(n5066) );
  NOR2X0 U5542 ( .IN1(n5070), .IN2(n5071), .QN(n5064) );
  NOR2X0 U5543 ( .IN1(n1635), .IN2(n4843), .QN(n5071) );
  NOR2X0 U5544 ( .IN1(n2717), .IN2(n4870), .QN(n5070) );
  NAND2X0 U5545 ( .IN1(n5072), .IN2(n5073), .QN(n5062) );
  NOR2X0 U5546 ( .IN1(n5074), .IN2(n5075), .QN(n5073) );
  NAND2X0 U5547 ( .IN1(n5076), .IN2(n5077), .QN(n5075) );
  NAND2X0 U5548 ( .IN1(n4855), .IN2(g1341), .QN(n5077) );
  NAND2X0 U5549 ( .IN1(n4925), .IN2(g1747), .QN(n5076) );
  NOR2X0 U5550 ( .IN1(n2727), .IN2(n4867), .QN(n5074) );
  NOR2X0 U5551 ( .IN1(n5078), .IN2(n5079), .QN(n5072) );
  NAND2X0 U5552 ( .IN1(n5080), .IN2(n5081), .QN(n5079) );
  NAND2X0 U5553 ( .IN1(n4956), .IN2(g290), .QN(n5081) );
  NAND2X0 U5554 ( .IN1(n4740), .IN2(n3031), .QN(n5080) );
  NOR2X0 U5555 ( .IN1(n2709), .IN2(n4943), .QN(n5078) );
  NAND2X0 U5556 ( .IN1(n2934), .IN2(n4587), .QN(g10455) );
  INVX0 U5557 ( .INP(g10719), .ZN(n4587) );
  NAND2X0 U5558 ( .IN1(n5082), .IN2(n5083), .QN(g10719) );
  NOR2X0 U5559 ( .IN1(n5084), .IN2(n5085), .QN(n5083) );
  NAND2X0 U5560 ( .IN1(n5086), .IN2(n5087), .QN(n5085) );
  NOR2X0 U5561 ( .IN1(n5088), .IN2(n5089), .QN(n5087) );
  NAND2X0 U5562 ( .IN1(n5090), .IN2(n5091), .QN(n5089) );
  NAND2X0 U5563 ( .IN1(n4940), .IN2(g950), .QN(n5091) );
  INVX0 U5564 ( .INP(n510), .ZN(n4940) );
  NAND2X0 U5565 ( .IN1(g898), .IN2(n4865), .QN(n5090) );
  NOR2X0 U5566 ( .IN1(n2881), .IN2(n5049), .QN(n5088) );
  NOR2X0 U5567 ( .IN1(n5092), .IN2(n5093), .QN(n5086) );
  NAND2X0 U5568 ( .IN1(n5094), .IN2(n5095), .QN(n5093) );
  NAND2X0 U5569 ( .IN1(n4989), .IN2(g1314), .QN(n5095) );
  NAND2X0 U5570 ( .IN1(n4856), .IN2(g1721), .QN(n5094) );
  INVX0 U5571 ( .INP(n4858), .ZN(n4856) );
  NOR2X0 U5572 ( .IN1(n4849), .IN2(n5096), .QN(n5092) );
  INVX0 U5573 ( .INP(g1170), .ZN(n5096) );
  NAND2X0 U5574 ( .IN1(n5097), .IN2(n5098), .QN(n5084) );
  NOR2X0 U5575 ( .IN1(n5099), .IN2(n5100), .QN(n5098) );
  NAND2X0 U5576 ( .IN1(n4898), .IN2(n5101), .QN(n5100) );
  INVX0 U5577 ( .INP(n523), .ZN(n5101) );
  NAND2X0 U5578 ( .IN1(n5102), .IN2(n5103), .QN(n4898) );
  NOR2X0 U5579 ( .IN1(n1512), .IN2(n4855), .QN(n5103) );
  NOR2X0 U5580 ( .IN1(n4899), .IN2(n4982), .QN(n5102) );
  NAND2X0 U5581 ( .IN1(n5104), .IN2(n5105), .QN(n4982) );
  NOR2X0 U5582 ( .IN1(n523), .IN2(n4998), .QN(n5105) );
  NOR2X0 U5583 ( .IN1(n5106), .IN2(n3236), .QN(n5104) );
  NAND2X0 U5584 ( .IN1(n5107), .IN2(n5108), .QN(n3236) );
  NOR2X0 U5585 ( .IN1(n5109), .IN2(n5110), .QN(n5108) );
  NAND2X0 U5586 ( .IN1(n5049), .IN2(n510), .QN(n5110) );
  NAND2X0 U5587 ( .IN1(n5111), .IN2(n508), .QN(n510) );
  INVX0 U5588 ( .INP(n5112), .ZN(n5109) );
  NOR2X0 U5589 ( .IN1(n4865), .IN2(n1530), .QN(n5112) );
  NOR2X0 U5590 ( .IN1(n5113), .IN2(n5114), .QN(n5107) );
  NAND2X0 U5591 ( .IN1(n4871), .IN2(n5115), .QN(n5114) );
  INVX0 U5592 ( .INP(n5116), .ZN(n5113) );
  NOR2X0 U5593 ( .IN1(n4905), .IN2(n4906), .QN(n5116) );
  INVX0 U5594 ( .INP(n4981), .ZN(n4899) );
  NOR2X0 U5595 ( .IN1(n1613), .IN2(n4981), .QN(n5099) );
  NAND2X0 U5596 ( .IN1(n5117), .IN2(n3229), .QN(n4981) );
  NOR2X0 U5597 ( .IN1(n5118), .IN2(n5119), .QN(n5097) );
  NAND2X0 U5598 ( .IN1(n5120), .IN2(n5121), .QN(n5119) );
  NAND2X0 U5599 ( .IN1(n4998), .IN2(g123), .QN(n5121) );
  INVX0 U5600 ( .INP(n4900), .ZN(n4998) );
  NAND2X0 U5601 ( .IN1(n5117), .IN2(g42), .QN(n4900) );
  NOR2X0 U5602 ( .IN1(n5122), .IN2(n5123), .QN(n5117) );
  NAND2X0 U5603 ( .IN1(n5124), .IN2(n5125), .QN(n5122) );
  NAND2X0 U5604 ( .IN1(n4905), .IN2(g928), .QN(n5120) );
  NOR2X0 U5605 ( .IN1(n5126), .IN2(n5127), .QN(n4905) );
  NAND2X0 U5606 ( .IN1(n5128), .IN2(g44), .QN(n5126) );
  INVX0 U5607 ( .INP(n5129), .ZN(n5118) );
  NAND2X0 U5608 ( .IN1(n4906), .IN2(g886), .QN(n5129) );
  NOR2X0 U5609 ( .IN1(n5130), .IN2(n5127), .QN(n4906) );
  NAND2X0 U5610 ( .IN1(n5131), .IN2(g45), .QN(n5127) );
  NOR2X0 U5611 ( .IN1(n3229), .IN2(n5132), .QN(n5131) );
  NAND2X0 U5612 ( .IN1(n5124), .IN2(g43), .QN(n5130) );
  NOR2X0 U5613 ( .IN1(n5133), .IN2(n5134), .QN(n5082) );
  NAND2X0 U5614 ( .IN1(n5135), .IN2(n5136), .QN(n5134) );
  NOR2X0 U5615 ( .IN1(n5137), .IN2(n5138), .QN(n5136) );
  NAND2X0 U5616 ( .IN1(n5139), .IN2(n5140), .QN(n5138) );
  NAND2X0 U5617 ( .IN1(g1194), .IN2(n1512), .QN(n5140) );
  NAND2X0 U5618 ( .IN1(g922), .IN2(n1530), .QN(n5139) );
  NOR2X0 U5619 ( .IN1(n2708), .IN2(n4915), .QN(n5137) );
  NOR2X0 U5620 ( .IN1(n5141), .IN2(n5142), .QN(n5135) );
  NOR2X0 U5621 ( .IN1(n1649), .IN2(n4843), .QN(n5142) );
  NOR2X0 U5622 ( .IN1(n2699), .IN2(n4870), .QN(n5141) );
  NAND2X0 U5623 ( .IN1(n5143), .IN2(n5144), .QN(n5133) );
  NOR2X0 U5624 ( .IN1(n5145), .IN2(n5146), .QN(n5144) );
  NAND2X0 U5625 ( .IN1(n5147), .IN2(n5148), .QN(n5146) );
  NAND2X0 U5626 ( .IN1(n4855), .IN2(g1336), .QN(n5148) );
  NAND2X0 U5627 ( .IN1(n4925), .IN2(g1744), .QN(n5147) );
  NOR2X0 U5628 ( .IN1(n2729), .IN2(n4867), .QN(n5145) );
  NOR2X0 U5629 ( .IN1(n5149), .IN2(n5150), .QN(n5143) );
  NAND2X0 U5630 ( .IN1(n5151), .IN2(n5152), .QN(n5150) );
  NAND2X0 U5631 ( .IN1(n4956), .IN2(g287), .QN(n5152) );
  NAND2X0 U5632 ( .IN1(n4740), .IN2(n3051), .QN(n5151) );
  NOR2X0 U5633 ( .IN1(n2711), .IN2(n4943), .QN(n5149) );
  NAND2X0 U5634 ( .IN1(n2934), .IN2(n4689), .QN(g10377) );
  INVX0 U5635 ( .INP(g10663), .ZN(n4689) );
  NAND2X0 U5636 ( .IN1(n5153), .IN2(n5154), .QN(g10663) );
  NOR2X0 U5637 ( .IN1(n5155), .IN2(n5156), .QN(n5154) );
  NAND2X0 U5638 ( .IN1(n5157), .IN2(n5158), .QN(n5156) );
  NAND2X0 U5639 ( .IN1(g1188), .IN2(n4857), .QN(n5158) );
  INVX0 U5640 ( .INP(n4849), .ZN(n4857) );
  NOR2X0 U5641 ( .IN1(n5159), .IN2(n5160), .QN(n5157) );
  NOR2X0 U5642 ( .IN1(n1640), .IN2(n4858), .QN(n5160) );
  NOR2X0 U5643 ( .IN1(n2659), .IN2(n4889), .QN(n5159) );
  NAND2X0 U5644 ( .IN1(n5161), .IN2(n5162), .QN(n5155) );
  NOR2X0 U5645 ( .IN1(n1564), .IN2(n523), .QN(n5162) );
  NOR2X0 U5646 ( .IN1(n5163), .IN2(n5164), .QN(n523) );
  NAND2X0 U5647 ( .IN1(n3183), .IN2(n5165), .QN(n5164) );
  NOR2X0 U5648 ( .IN1(n5166), .IN2(n5124), .QN(n3183) );
  NAND2X0 U5649 ( .IN1(n3229), .IN2(n5125), .QN(n5166) );
  INVX0 U5650 ( .INP(n5167), .ZN(n5163) );
  NOR2X0 U5651 ( .IN1(n3233), .IN2(n5168), .QN(n5167) );
  NOR2X0 U5652 ( .IN1(n5169), .IN2(n5170), .QN(n5161) );
  NOR2X0 U5653 ( .IN1(n2650), .IN2(n5049), .QN(n5170) );
  NAND2X0 U5654 ( .IN1(n5171), .IN2(n508), .QN(n5049) );
  INVX0 U5655 ( .INP(n5172), .ZN(n5169) );
  NAND2X0 U5656 ( .IN1(n4865), .IN2(g916), .QN(n5172) );
  INVX0 U5657 ( .INP(n5173), .ZN(n4865) );
  NAND2X0 U5658 ( .IN1(n508), .IN2(n5174), .QN(n5173) );
  INVX0 U5659 ( .INP(n5132), .ZN(n508) );
  NAND2X0 U5660 ( .IN1(n3230), .IN2(n5165), .QN(n5132) );
  NOR2X0 U5661 ( .IN1(n5168), .IN2(n4693), .QN(n3230) );
  NOR2X0 U5662 ( .IN1(n5175), .IN2(n5176), .QN(n5153) );
  NAND2X0 U5663 ( .IN1(n5177), .IN2(n5178), .QN(n5176) );
  NOR2X0 U5664 ( .IN1(n5179), .IN2(n5180), .QN(n5178) );
  NOR2X0 U5665 ( .IN1(n4855), .IN2(n4947), .QN(n5180) );
  NAND2X0 U5666 ( .IN1(n1478), .IN2(n5181), .QN(n4947) );
  INVX0 U5667 ( .INP(n5106), .ZN(n5181) );
  NAND2X0 U5668 ( .IN1(n5182), .IN2(n5183), .QN(n5106) );
  NOR2X0 U5669 ( .IN1(n4925), .IN2(n5184), .QN(n5183) );
  NAND2X0 U5670 ( .IN1(n4852), .IN2(n4854), .QN(n5184) );
  INVX0 U5671 ( .INP(n1567), .ZN(n4854) );
  NAND2X0 U5672 ( .IN1(n4943), .IN2(n5185), .QN(n1567) );
  NAND2X0 U5673 ( .IN1(n5171), .IN2(n507), .QN(n5185) );
  NAND2X0 U5674 ( .IN1(n5111), .IN2(n507), .QN(n4943) );
  INVX0 U5675 ( .INP(n1566), .ZN(n4852) );
  NAND2X0 U5676 ( .IN1(n4915), .IN2(n5186), .QN(n1566) );
  NAND2X0 U5677 ( .IN1(n507), .IN2(n5174), .QN(n5186) );
  INVX0 U5678 ( .INP(n1479), .ZN(n4915) );
  INVX0 U5679 ( .INP(n4963), .ZN(n4925) );
  NOR2X0 U5680 ( .IN1(n4989), .IN2(n5187), .QN(n5182) );
  NAND2X0 U5681 ( .IN1(n4858), .IN2(n4849), .QN(n5187) );
  NAND2X0 U5682 ( .IN1(n1544), .IN2(n5174), .QN(n4849) );
  NOR2X0 U5683 ( .IN1(n5188), .IN2(n5124), .QN(n5174) );
  NAND2X0 U5684 ( .IN1(n5125), .IN2(g42), .QN(n5188) );
  NOR2X0 U5685 ( .IN1(n5128), .IN2(g45), .QN(n5125) );
  INVX0 U5686 ( .INP(g43), .ZN(n5128) );
  NAND2X0 U5687 ( .IN1(n5189), .IN2(g42), .QN(n4858) );
  INVX0 U5688 ( .INP(n4889), .ZN(n4989) );
  NAND2X0 U5689 ( .IN1(n5111), .IN2(n1544), .QN(n4889) );
  NOR2X0 U5690 ( .IN1(n5190), .IN2(g42), .QN(n5111) );
  INVX0 U5691 ( .INP(n4842), .ZN(n4855) );
  NOR2X0 U5692 ( .IN1(n2660), .IN2(n4842), .QN(n5179) );
  NAND2X0 U5693 ( .IN1(n5171), .IN2(n1544), .QN(n4842) );
  NOR2X0 U5694 ( .IN1(n5190), .IN2(n3229), .QN(n5171) );
  NAND2X0 U5695 ( .IN1(n4691), .IN2(g45), .QN(n5190) );
  NOR2X0 U5696 ( .IN1(g44), .IN2(g43), .QN(n4691) );
  NOR2X0 U5697 ( .IN1(n5191), .IN2(n5192), .QN(n5177) );
  NOR2X0 U5698 ( .IN1(n2721), .IN2(n4843), .QN(n5192) );
  INVX0 U5699 ( .INP(n1486), .ZN(n4843) );
  NOR2X0 U5700 ( .IN1(n2704), .IN2(n4870), .QN(n5191) );
  INVX0 U5701 ( .INP(n1485), .ZN(n4870) );
  NAND2X0 U5702 ( .IN1(n5193), .IN2(n5194), .QN(n5175) );
  NAND2X0 U5703 ( .IN1(n4740), .IN2(n1637), .QN(n5194) );
  NOR2X0 U5704 ( .IN1(n5195), .IN2(n5196), .QN(n5193) );
  NOR2X0 U5705 ( .IN1(n2737), .IN2(n4867), .QN(n5196) );
  INVX0 U5706 ( .INP(n4951), .ZN(n4867) );
  NOR2X0 U5707 ( .IN1(n5115), .IN2(n4956), .QN(n4951) );
  NOR2X0 U5708 ( .IN1(n5115), .IN2(g42), .QN(n4956) );
  NAND2X0 U5709 ( .IN1(n5197), .IN2(n5198), .QN(n5115) );
  NOR2X0 U5710 ( .IN1(g45), .IN2(g43), .QN(n5198) );
  NOR2X0 U5711 ( .IN1(n5124), .IN2(n5123), .QN(n5197) );
  INVX0 U5712 ( .INP(n507), .ZN(n5123) );
  NOR2X0 U5713 ( .IN1(n5199), .IN2(n4693), .QN(n507) );
  NAND2X0 U5714 ( .IN1(n5200), .IN2(n3267), .QN(n4693) );
  INVX0 U5715 ( .INP(g47), .ZN(n5200) );
  INVX0 U5716 ( .INP(g44), .ZN(n5124) );
  NOR2X0 U5717 ( .IN1(n2885), .IN2(n4963), .QN(n5195) );
  NAND2X0 U5718 ( .IN1(n5189), .IN2(n3229), .QN(n4963) );
  INVX0 U5719 ( .INP(g42), .ZN(n3229) );
  NOR2X0 U5720 ( .IN1(n5201), .IN2(n5202), .QN(n5189) );
  NAND2X0 U5721 ( .IN1(g43), .IN2(g44), .QN(n5202) );
  NAND2X0 U5722 ( .IN1(n1544), .IN2(g45), .QN(n5201) );
  NOR2X0 U5723 ( .IN1(n5199), .IN2(n3233), .QN(n1544) );
  NAND2X0 U5724 ( .IN1(g47), .IN2(n3267), .QN(n3233) );
  NAND2X0 U5725 ( .IN1(n5203), .IN2(n5204), .QN(n3267) );
  NAND2X0 U5726 ( .IN1(n5205), .IN2(n5206), .QN(n5204) );
  INVX0 U5727 ( .INP(g30), .ZN(n5206) );
  NOR2X0 U5728 ( .IN1(g48), .IN2(g41), .QN(n5205) );
  NAND2X0 U5729 ( .IN1(n4871), .IN2(n5165), .QN(n5203) );
  NAND2X0 U5730 ( .IN1(n5168), .IN2(n5165), .QN(n5199) );
  NOR2X0 U5731 ( .IN1(n5207), .IN2(g41), .QN(n5165) );
  INVX0 U5732 ( .INP(g46), .ZN(n5168) );
  NOR2X0 U5733 ( .IN1(n4740), .IN2(g30), .QN(n2934) );
  INVX0 U5734 ( .INP(n4871), .ZN(n4740) );
  NOR2X0 U5735 ( .IN1(n5207), .IN2(g31), .QN(n4871) );
  INVX0 U5736 ( .INP(g48), .ZN(n5207) );
  XNOR2X1 U5737 ( .IN1(test_so1), .IN2(n3720), .Q(N599) );
  NAND2X0 U5738 ( .IN1(n5208), .IN2(n1093), .QN(n3720) );
  NOR2X0 U5739 ( .IN1(n2925), .IN2(n2920), .QN(n5208) );
  NOR2X0 U1550_U2 ( .IN1(g10722), .IN2(n2934), .QN(U1550_n1) );
  INVX0 U1550_U1 ( .INP(U1550_n1), .ZN(g10461) );
  NOR2X0 U1551_U2 ( .IN1(g10664), .IN2(n2934), .QN(U1551_n1) );
  INVX0 U1551_U1 ( .INP(U1551_n1), .ZN(g10379) );
  INVX0 U1586_U2 ( .INP(n23), .ZN(U1586_n1) );
  NOR2X0 U1586_U1 ( .IN1(n2929), .IN2(U1586_n1), .QN(n1855) );
  INVX0 U1754_U2 ( .INP(n507), .ZN(U1754_n1) );
  NOR2X0 U1754_U1 ( .IN1(n527), .IN2(U1754_n1), .QN(n1479) );
  INVX0 U1798_U2 ( .INP(n1567), .ZN(U1798_n1) );
  NOR2X0 U1798_U1 ( .IN1(n1480), .IN2(U1798_n1), .QN(n1485) );
  INVX0 U1839_U2 ( .INP(n1566), .ZN(U1839_n1) );
  NOR2X0 U1839_U1 ( .IN1(n1479), .IN2(U1839_n1), .QN(n1486) );
  INVX0 U1843_U2 ( .INP(n1546), .ZN(U1843_n1) );
  NOR2X0 U1843_U1 ( .IN1(n523), .IN2(U1843_n1), .QN(n1478) );
  INVX0 U1877_U2 ( .INP(n1137), .ZN(U1877_n1) );
  NOR2X0 U1877_U1 ( .IN1(n2939), .IN2(U1877_n1), .QN(n1195) );
  INVX0 U1908_U2 ( .INP(n1544), .ZN(U1908_n1) );
  NOR2X0 U1908_U1 ( .IN1(n527), .IN2(U1908_n1), .QN(n1512) );
  INVX0 U1909_U2 ( .INP(n508), .ZN(U1909_n1) );
  NOR2X0 U1909_U1 ( .IN1(n527), .IN2(U1909_n1), .QN(n1530) );
  INVX0 U1987_U2 ( .INP(n822), .ZN(U1987_n1) );
  NOR2X0 U1987_U1 ( .IN1(n250), .IN2(U1987_n1), .QN(n916) );
  INVX0 U2031_U2 ( .INP(n1057), .ZN(U2031_n1) );
  NOR2X0 U2031_U1 ( .IN1(n1054), .IN2(U2031_n1), .QN(n1056) );
  INVX0 U2035_U2 ( .INP(n1404), .ZN(U2035_n1) );
  NOR2X0 U2035_U1 ( .IN1(g109), .IN2(U2035_n1), .QN(n1450) );
  INVX0 U2418_U2 ( .INP(g968), .ZN(U2418_n1) );
  NOR2X0 U2418_U1 ( .IN1(n510), .IN2(U2418_n1), .QN(n1564) );
  INVX0 U2468_U2 ( .INP(g1336), .ZN(U2468_n1) );
  NOR2X0 U2468_U1 ( .IN1(n1227), .IN2(U2468_n1), .QN(n1231) );
  INVX0 U2478_U2 ( .INP(g1341), .ZN(U2478_n1) );
  NOR2X0 U2478_U1 ( .IN1(n228), .IN2(U2478_n1), .QN(n1232) );
  INVX0 U2488_U2 ( .INP(n1262), .ZN(U2488_n1) );
  NOR2X0 U2488_U1 ( .IN1(n1258), .IN2(U2488_n1), .QN(n1260) );
  INVX0 U2533_U2 ( .INP(g178), .ZN(U2533_n1) );
  NOR2X0 U2533_U1 ( .IN1(n2939), .IN2(U2533_n1), .QN(g6786) );
  INVX0 U2534_U2 ( .INP(g1424), .ZN(U2534_n1) );
  NOR2X0 U2534_U1 ( .IN1(n2940), .IN2(U2534_n1), .QN(g6234) );
  INVX0 U2639_U2 ( .INP(n962), .ZN(U2639_n1) );
  NOR2X0 U2639_U1 ( .IN1(n958), .IN2(U2639_n1), .QN(n804) );
  INVX0 U2641_U2 ( .INP(n62), .ZN(U2641_n1) );
  NOR2X0 U2641_U1 ( .IN1(g1868), .IN2(U2641_n1), .QN(n926) );
  INVX0 U2654_U2 ( .INP(g746), .ZN(U2654_n1) );
  NOR2X0 U2654_U1 ( .IN1(g750), .IN2(U2654_n1), .QN(g4171) );
  INVX0 U2658_U2 ( .INP(n917), .ZN(U2658_n1) );
  NOR2X0 U2658_U1 ( .IN1(n918), .IN2(U2658_n1), .QN(n812) );
  INVX0 U2683_U2 ( .INP(g382), .ZN(U2683_n1) );
  NOR2X0 U2683_U1 ( .IN1(n1385), .IN2(U2683_n1), .QN(n1420) );
  INVX0 U2699_U2 ( .INP(n249), .ZN(U2699_n1) );
  NOR2X0 U2699_U1 ( .IN1(n487), .IN2(U2699_n1), .QN(n806) );
  INVX0 U2846_U2 ( .INP(g4175), .ZN(U2846_n1) );
  NOR2X0 U2846_U1 ( .IN1(n1214), .IN2(U2846_n1), .QN(n1193) );
  INVX0 U2847_U2 ( .INP(g4177), .ZN(U2847_n1) );
  NOR2X0 U2847_U1 ( .IN1(n1153), .IN2(U2847_n1), .QN(n1125) );
  INVX0 U2848_U2 ( .INP(g4179), .ZN(U2848_n1) );
  NOR2X0 U2848_U1 ( .IN1(n1099), .IN2(U2848_n1), .QN(n1093) );
  INVX0 U2859_U2 ( .INP(n1137), .ZN(U2859_n1) );
  NOR2X0 U2859_U1 ( .IN1(g12), .IN2(U2859_n1), .QN(n1159) );
  INVX0 U2860_U2 ( .INP(g810), .ZN(U2860_n1) );
  NOR2X0 U2860_U1 ( .IN1(n1151), .IN2(U2860_n1), .QN(n1123) );
  INVX0 U2861_U2 ( .INP(g818), .ZN(U2861_n1) );
  NOR2X0 U2861_U1 ( .IN1(n1097), .IN2(U2861_n1), .QN(n1090) );
  INVX0 U2867_U2 ( .INP(n817), .ZN(U2867_n1) );
  NOR2X0 U2867_U1 ( .IN1(g1834), .IN2(U2867_n1), .QN(n1380) );
  INVX0 U2879_U2 ( .INP(g713), .ZN(U2879_n1) );
  NOR2X0 U2879_U1 ( .IN1(n1656), .IN2(U2879_n1), .QN(n967) );
  INVX0 U2881_U2 ( .INP(g1927), .ZN(U2881_n1) );
  NOR2X0 U2881_U1 ( .IN1(n1657), .IN2(U2881_n1), .QN(n921) );
  INVX0 U2882_U2 ( .INP(g1160), .ZN(U2882_n1) );
  NOR2X0 U2882_U1 ( .IN1(n2941), .IN2(U2882_n1), .QN(g4334) );
  INVX0 U2883_U2 ( .INP(g1166), .ZN(U2883_n1) );
  NOR2X0 U2883_U1 ( .IN1(n2942), .IN2(U2883_n1), .QN(g4325) );
  INVX0 U2884_U2 ( .INP(g148), .ZN(U2884_n1) );
  NOR2X0 U2884_U1 ( .IN1(n2939), .IN2(U2884_n1), .QN(g6759) );
  INVX0 U2885_U2 ( .INP(g1157), .ZN(U2885_n1) );
  NOR2X0 U2885_U1 ( .IN1(n2940), .IN2(U2885_n1), .QN(g4338) );
  INVX0 U2886_U2 ( .INP(g1163), .ZN(U2886_n1) );
  NOR2X0 U2886_U1 ( .IN1(n2941), .IN2(U2886_n1), .QN(g4330) );
  INVX0 U2887_U2 ( .INP(g237), .ZN(U2887_n1) );
  NOR2X0 U2887_U1 ( .IN1(n2942), .IN2(U2887_n1), .QN(g6821) );
  INVX0 U2888_U2 ( .INP(g1499), .ZN(U2888_n1) );
  NOR2X0 U2888_U1 ( .IN1(n2939), .IN2(U2888_n1), .QN(g6198) );
  INVX0 U2889_U2 ( .INP(g1411), .ZN(U2889_n1) );
  NOR2X0 U2889_U1 ( .IN1(n2940), .IN2(U2889_n1), .QN(g6244) );
  INVX0 U2890_U2 ( .INP(g225), .ZN(U2890_n1) );
  NOR2X0 U2890_U1 ( .IN1(n2941), .IN2(U2890_n1), .QN(g6826) );
  INVX0 U2891_U2 ( .INP(g1407), .ZN(U2891_n1) );
  NOR2X0 U2891_U1 ( .IN1(n2942), .IN2(U2891_n1), .QN(g6216) );
  INVX0 U2892_U2 ( .INP(g213), .ZN(U2892_n1) );
  NOR2X0 U2892_U1 ( .IN1(n2939), .IN2(U2892_n1), .QN(g6829) );
  INVX0 U2893_U2 ( .INP(g186), .ZN(U2893_n1) );
  NOR2X0 U2893_U1 ( .IN1(n2940), .IN2(U2893_n1), .QN(g6833) );
  INVX0 U2894_U2 ( .INP(g219), .ZN(U2894_n1) );
  NOR2X0 U2894_U1 ( .IN1(n2941), .IN2(U2894_n1), .QN(g6827) );
  INVX0 U2895_U2 ( .INP(g143), .ZN(U2895_n1) );
  NOR2X0 U2895_U1 ( .IN1(n2942), .IN2(U2895_n1), .QN(g6757) );
  INVX0 U2896_U2 ( .INP(g207), .ZN(U2896_n1) );
  NOR2X0 U2896_U1 ( .IN1(n2939), .IN2(U2896_n1), .QN(g6831) );
  INVX0 U2897_U2 ( .INP(g231), .ZN(U2897_n1) );
  NOR2X0 U2897_U1 ( .IN1(n2940), .IN2(U2897_n1), .QN(g6822) );
  INVX0 U2898_U2 ( .INP(g192), .ZN(U2898_n1) );
  NOR2X0 U2898_U1 ( .IN1(n2941), .IN2(U2898_n1), .QN(g6838) );
  INVX0 U2899_U2 ( .INP(test_so3), .ZN(U2899_n1) );
  NOR2X0 U2899_U1 ( .IN1(n2942), .IN2(U2899_n1), .QN(g6823) );
  INVX0 U2900_U2 ( .INP(g1371), .ZN(U2900_n1) );
  NOR2X0 U2900_U1 ( .IN1(n2939), .IN2(U2900_n1), .QN(g6824) );
  INVX0 U2901_U2 ( .INP(g1383), .ZN(U2901_n1) );
  NOR2X0 U2901_U1 ( .IN1(n2940), .IN2(U2901_n1), .QN(g6832) );
  INVX0 U2902_U2 ( .INP(g243), .ZN(U2902_n1) );
  NOR2X0 U2902_U1 ( .IN1(n2941), .IN2(U2902_n1), .QN(g6819) );
  INVX0 U3090_U2 ( .INP(n1151), .ZN(U3090_n1) );
  NOR2X0 U3090_U1 ( .IN1(g810), .IN2(U3090_n1), .QN(n1150) );
  INVX0 U3092_U2 ( .INP(n1097), .ZN(U3092_n1) );
  NOR2X0 U3092_U1 ( .IN1(g818), .IN2(U3092_n1), .QN(n1096) );
  INVX0 U3094_U2 ( .INP(n1099), .ZN(U3094_n1) );
  NOR2X0 U3094_U1 ( .IN1(g4179), .IN2(U3094_n1), .QN(n1098) );
  INVX0 U3096_U2 ( .INP(n1214), .ZN(U3096_n1) );
  NOR2X0 U3096_U1 ( .IN1(g4175), .IN2(U3096_n1), .QN(n1213) );
  INVX0 U3098_U2 ( .INP(n1153), .ZN(U3098_n1) );
  NOR2X0 U3098_U1 ( .IN1(g4177), .IN2(U3098_n1), .QN(n1152) );
  INVX0 U3124_U2 ( .INP(n837), .ZN(U3124_n1) );
  NOR2X0 U3124_U1 ( .IN1(n838), .IN2(U3124_n1), .QN(n836) );
  INVX0 U3171_U2 ( .INP(g1610), .ZN(U3171_n1) );
  NOR2X0 U3171_U1 ( .IN1(n364), .IN2(U3171_n1), .QN(g5194) );
endmodule

