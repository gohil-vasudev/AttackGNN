module add_mul_mix_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        c_0_, c_1_, c_2_, c_3_, d_0_, d_1_, d_2_, d_3_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, c_0_, c_1_, c_2_, c_3_,
         d_0_, d_1_, d_2_, d_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238;

  XOR2_X1 U122 ( .A(n116), .B(n117), .Z(Result_6_) );
  NOR2_X1 U123 ( .A1(n118), .A2(n119), .ZN(n116) );
  XNOR2_X1 U124 ( .A(n120), .B(n121), .ZN(Result_5_) );
  NAND2_X1 U125 ( .A1(n122), .A2(n123), .ZN(n120) );
  XOR2_X1 U126 ( .A(n124), .B(n125), .Z(Result_4_) );
  XNOR2_X1 U127 ( .A(n126), .B(n127), .ZN(n125) );
  XOR2_X1 U128 ( .A(n128), .B(n129), .Z(Result_3_) );
  XOR2_X1 U129 ( .A(n130), .B(n131), .Z(Result_2_) );
  XOR2_X1 U130 ( .A(n132), .B(n133), .Z(Result_1_) );
  NAND2_X1 U131 ( .A1(n134), .A2(n135), .ZN(Result_0_) );
  NAND2_X1 U132 ( .A1(n133), .A2(n132), .ZN(n135) );
  NOR2_X1 U133 ( .A1(n136), .A2(n137), .ZN(n132) );
  INV_X1 U134 ( .A(n138), .ZN(n137) );
  NAND2_X1 U135 ( .A1(n139), .A2(n140), .ZN(n138) );
  NOR2_X1 U136 ( .A1(n130), .A2(n131), .ZN(n133) );
  XNOR2_X1 U137 ( .A(n141), .B(n142), .ZN(n131) );
  INV_X1 U138 ( .A(n143), .ZN(n130) );
  NOR2_X1 U139 ( .A1(n128), .A2(n129), .ZN(n143) );
  XOR2_X1 U140 ( .A(n144), .B(n145), .Z(n129) );
  NAND2_X1 U141 ( .A1(n146), .A2(n147), .ZN(n144) );
  NAND2_X1 U142 ( .A1(n148), .A2(n149), .ZN(n128) );
  NAND2_X1 U143 ( .A1(n124), .A2(n150), .ZN(n149) );
  NAND2_X1 U144 ( .A1(n127), .A2(n126), .ZN(n150) );
  XNOR2_X1 U145 ( .A(n151), .B(n152), .ZN(n124) );
  XOR2_X1 U146 ( .A(n153), .B(n154), .Z(n152) );
  NAND2_X1 U147 ( .A1(n155), .A2(n156), .ZN(n154) );
  INV_X1 U148 ( .A(n157), .ZN(n148) );
  NOR2_X1 U149 ( .A1(n126), .A2(n127), .ZN(n157) );
  NOR2_X1 U150 ( .A1(n158), .A2(n118), .ZN(n127) );
  NAND2_X1 U151 ( .A1(n122), .A2(n159), .ZN(n126) );
  NAND2_X1 U152 ( .A1(n121), .A2(n123), .ZN(n159) );
  NAND2_X1 U153 ( .A1(n160), .A2(n161), .ZN(n123) );
  NAND2_X1 U154 ( .A1(n155), .A2(n162), .ZN(n161) );
  XOR2_X1 U155 ( .A(n163), .B(n164), .Z(n121) );
  NOR2_X1 U156 ( .A1(n165), .A2(n166), .ZN(n163) );
  NAND2_X1 U157 ( .A1(n167), .A2(n155), .ZN(n122) );
  INV_X1 U158 ( .A(n160), .ZN(n167) );
  NAND2_X1 U159 ( .A1(Result_7_), .A2(n164), .ZN(n160) );
  NOR2_X1 U160 ( .A1(n168), .A2(n119), .ZN(n164) );
  NOR2_X1 U161 ( .A1(n118), .A2(n166), .ZN(Result_7_) );
  INV_X1 U162 ( .A(n162), .ZN(n118) );
  XOR2_X1 U163 ( .A(c_3_), .B(d_3_), .Z(n162) );
  NOR2_X1 U164 ( .A1(n136), .A2(n169), .ZN(n134) );
  NOR2_X1 U165 ( .A1(n170), .A2(n158), .ZN(n169) );
  NOR2_X1 U166 ( .A1(n171), .A2(n172), .ZN(n170) );
  NOR2_X1 U167 ( .A1(n173), .A2(n174), .ZN(n171) );
  NOR2_X1 U168 ( .A1(n140), .A2(n139), .ZN(n136) );
  NAND2_X1 U169 ( .A1(n175), .A2(n176), .ZN(n139) );
  NAND2_X1 U170 ( .A1(n177), .A2(n178), .ZN(n176) );
  NAND2_X1 U171 ( .A1(n179), .A2(n180), .ZN(n178) );
  NOR2_X1 U172 ( .A1(n181), .A2(n173), .ZN(n179) );
  INV_X1 U173 ( .A(n172), .ZN(n177) );
  NAND2_X1 U174 ( .A1(n180), .A2(n172), .ZN(n175) );
  NAND2_X1 U175 ( .A1(n182), .A2(n183), .ZN(n172) );
  NAND2_X1 U176 ( .A1(n155), .A2(n184), .ZN(n183) );
  NAND2_X1 U177 ( .A1(n142), .A2(n141), .ZN(n140) );
  NAND2_X1 U178 ( .A1(n146), .A2(n185), .ZN(n141) );
  NAND2_X1 U179 ( .A1(n145), .A2(n147), .ZN(n185) );
  NAND2_X1 U180 ( .A1(n186), .A2(n187), .ZN(n147) );
  NAND2_X1 U181 ( .A1(n180), .A2(n156), .ZN(n187) );
  INV_X1 U182 ( .A(n168), .ZN(n156) );
  INV_X1 U183 ( .A(n188), .ZN(n186) );
  XOR2_X1 U184 ( .A(n189), .B(n190), .Z(n145) );
  XOR2_X1 U185 ( .A(n191), .B(n174), .Z(n190) );
  INV_X1 U186 ( .A(n181), .ZN(n174) );
  NAND2_X1 U187 ( .A1(n180), .A2(n188), .ZN(n146) );
  NAND2_X1 U188 ( .A1(n192), .A2(n193), .ZN(n188) );
  NAND2_X1 U189 ( .A1(n194), .A2(n155), .ZN(n193) );
  NOR2_X1 U190 ( .A1(n195), .A2(n168), .ZN(n194) );
  NOR2_X1 U191 ( .A1(n196), .A2(n151), .ZN(n195) );
  NAND2_X1 U192 ( .A1(n196), .A2(n151), .ZN(n192) );
  XOR2_X1 U193 ( .A(n197), .B(n198), .Z(n151) );
  INV_X1 U194 ( .A(n153), .ZN(n196) );
  NAND2_X1 U195 ( .A1(n197), .A2(n117), .ZN(n153) );
  NOR2_X1 U196 ( .A1(n168), .A2(n166), .ZN(n117) );
  XOR2_X1 U197 ( .A(n199), .B(n200), .Z(n168) );
  XOR2_X1 U198 ( .A(d_2_), .B(c_2_), .Z(n200) );
  NAND2_X1 U199 ( .A1(c_3_), .A2(d_3_), .ZN(n199) );
  XNOR2_X1 U200 ( .A(n201), .B(n202), .ZN(n142) );
  NOR2_X1 U201 ( .A1(n173), .A2(n203), .ZN(n202) );
  NAND2_X1 U202 ( .A1(n182), .A2(n204), .ZN(n201) );
  NAND2_X1 U203 ( .A1(n205), .A2(n206), .ZN(n204) );
  NAND2_X1 U204 ( .A1(n207), .A2(n180), .ZN(n206) );
  INV_X1 U205 ( .A(n184), .ZN(n205) );
  NAND2_X1 U206 ( .A1(n180), .A2(n184), .ZN(n182) );
  NAND2_X1 U207 ( .A1(n208), .A2(n191), .ZN(n184) );
  NAND2_X1 U208 ( .A1(n198), .A2(n197), .ZN(n191) );
  NOR2_X1 U209 ( .A1(n165), .A2(n119), .ZN(n197) );
  NOR2_X1 U210 ( .A1(n166), .A2(n173), .ZN(n198) );
  XNOR2_X1 U211 ( .A(a_3_), .B(b_3_), .ZN(n166) );
  NAND2_X1 U212 ( .A1(n189), .A2(n181), .ZN(n208) );
  NOR2_X1 U213 ( .A1(n165), .A2(n203), .ZN(n181) );
  INV_X1 U214 ( .A(n155), .ZN(n203) );
  XOR2_X1 U215 ( .A(n209), .B(n210), .Z(n155) );
  XOR2_X1 U216 ( .A(b_1_), .B(a_1_), .Z(n210) );
  INV_X1 U217 ( .A(n207), .ZN(n165) );
  XOR2_X1 U218 ( .A(n211), .B(n212), .Z(n207) );
  XOR2_X1 U219 ( .A(d_1_), .B(c_1_), .Z(n212) );
  NOR2_X1 U220 ( .A1(n173), .A2(n119), .ZN(n189) );
  XOR2_X1 U221 ( .A(n213), .B(n214), .Z(n119) );
  XOR2_X1 U222 ( .A(b_2_), .B(a_2_), .Z(n214) );
  NAND2_X1 U223 ( .A1(a_3_), .A2(b_3_), .ZN(n213) );
  XOR2_X1 U224 ( .A(n215), .B(n216), .Z(n173) );
  XOR2_X1 U225 ( .A(d_0_), .B(c_0_), .Z(n216) );
  NAND2_X1 U226 ( .A1(n217), .A2(n218), .ZN(n215) );
  NAND2_X1 U227 ( .A1(n219), .A2(n220), .ZN(n218) );
  INV_X1 U228 ( .A(d_1_), .ZN(n220) );
  NAND2_X1 U229 ( .A1(c_1_), .A2(n211), .ZN(n219) );
  INV_X1 U230 ( .A(n221), .ZN(n217) );
  NOR2_X1 U231 ( .A1(n211), .A2(c_1_), .ZN(n221) );
  NAND2_X1 U232 ( .A1(n222), .A2(n223), .ZN(n211) );
  NAND2_X1 U233 ( .A1(n224), .A2(c_3_), .ZN(n223) );
  NOR2_X1 U234 ( .A1(n225), .A2(n226), .ZN(n224) );
  INV_X1 U235 ( .A(d_3_), .ZN(n226) );
  NOR2_X1 U236 ( .A1(c_2_), .A2(d_2_), .ZN(n225) );
  NAND2_X1 U237 ( .A1(c_2_), .A2(d_2_), .ZN(n222) );
  INV_X1 U238 ( .A(n158), .ZN(n180) );
  XOR2_X1 U239 ( .A(n227), .B(n228), .Z(n158) );
  XOR2_X1 U240 ( .A(b_0_), .B(a_0_), .Z(n228) );
  NAND2_X1 U241 ( .A1(n229), .A2(n230), .ZN(n227) );
  NAND2_X1 U242 ( .A1(n231), .A2(n232), .ZN(n230) );
  INV_X1 U243 ( .A(b_1_), .ZN(n232) );
  NAND2_X1 U244 ( .A1(a_1_), .A2(n209), .ZN(n231) );
  INV_X1 U245 ( .A(n233), .ZN(n229) );
  NOR2_X1 U246 ( .A1(n209), .A2(a_1_), .ZN(n233) );
  NAND2_X1 U247 ( .A1(n234), .A2(n235), .ZN(n209) );
  NAND2_X1 U248 ( .A1(n236), .A2(a_3_), .ZN(n235) );
  NOR2_X1 U249 ( .A1(n237), .A2(n238), .ZN(n236) );
  INV_X1 U250 ( .A(b_3_), .ZN(n238) );
  NOR2_X1 U251 ( .A1(a_2_), .A2(b_2_), .ZN(n237) );
  NAND2_X1 U252 ( .A1(a_2_), .A2(b_2_), .ZN(n234) );
endmodule

