module locked_c1355 (  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT  );
  input  G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n374_, new_n375_, new_n376_, new_n378_, new_n379_, new_n381_, new_n382_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n404_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n415_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n426_, new_n427_, new_n429_, new_n431_, new_n432_, new_n434_, new_n435_, new_n437_, new_n439_, new_n441_, new_n442_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n470_, new_n471_, new_n472_, new_n474_, new_n475_, new_n477_, new_n478_, new_n480_, new_n481_, new_n483_, new_n484_, new_n485_, new_n487_, new_n489_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n515_, new_n517_, new_n518_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n531_, new_n532_, new_n534_, new_n536_, new_n537_;
  INV_X1 g000 ( .A(G1GAT), .ZN(new_n138_) );
  XNOR2_X1 g001 ( .A(G155GAT), .B(KEYINPUT3), .ZN(new_n139_) );
  XNOR2_X1 g002 ( .A(G141GAT), .B(KEYINPUT2), .ZN(new_n140_) );
  XNOR2_X1 g003 ( .A(new_n139_), .B(new_n140_), .ZN(new_n141_) );
  XNOR2_X1 g004 ( .A(G57GAT), .B(KEYINPUT1), .ZN(new_n142_) );
  NAND2_X1 g005 ( .A1(G225GAT), .A2(G233GAT), .ZN(new_n143_) );
  XNOR2_X1 g006 ( .A(new_n142_), .B(new_n143_), .ZN(new_n144_) );
  XNOR2_X1 g007 ( .A(new_n141_), .B(new_n144_), .ZN(new_n145_) );
  XNOR2_X1 g008 ( .A(G120GAT), .B(G127GAT), .ZN(new_n146_) );
  XNOR2_X1 g009 ( .A(G113GAT), .B(KEYINPUT0), .ZN(new_n147_) );
  XNOR2_X1 g010 ( .A(new_n146_), .B(new_n147_), .ZN(new_n148_) );
  XNOR2_X1 g011 ( .A(new_n148_), .B(new_n138_), .ZN(new_n149_) );
  XNOR2_X1 g012 ( .A(new_n145_), .B(new_n149_), .ZN(new_n150_) );
  XNOR2_X1 g013 ( .A(G29GAT), .B(G134GAT), .ZN(new_n151_) );
  NAND2_X1 g014 ( .A1(new_n150_), .A2(new_n151_), .ZN(new_n152_) );
  OR2_X1 g015 ( .A1(new_n150_), .A2(new_n151_), .ZN(new_n153_) );
  NAND2_X1 g016 ( .A1(new_n153_), .A2(new_n152_), .ZN(new_n154_) );
  XOR2_X1 g017 ( .A(G85GAT), .B(G162GAT), .Z(new_n155_) );
  INV_X1 g018 ( .A(new_n155_), .ZN(new_n156_) );
  NAND2_X1 g019 ( .A1(new_n154_), .A2(new_n156_), .ZN(new_n157_) );
  NAND3_X1 g020 ( .A1(new_n153_), .A2(new_n152_), .A3(new_n155_), .ZN(new_n158_) );
  NAND2_X1 g021 ( .A1(new_n157_), .A2(new_n158_), .ZN(new_n159_) );
  XOR2_X1 g022 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(new_n160_) );
  XNOR2_X1 g023 ( .A(G148GAT), .B(KEYINPUT6), .ZN(new_n161_) );
  XNOR2_X1 g024 ( .A(new_n160_), .B(new_n161_), .ZN(new_n162_) );
  XOR2_X1 g025 ( .A(new_n159_), .B(new_n162_), .Z(new_n163_) );
  INV_X1 g026 ( .A(KEYINPUT26), .ZN(new_n164_) );
  INV_X1 g027 ( .A(new_n141_), .ZN(new_n165_) );
  INV_X1 g028 ( .A(G197GAT), .ZN(new_n166_) );
  XNOR2_X1 g029 ( .A(G211GAT), .B(G218GAT), .ZN(new_n167_) );
  XNOR2_X1 g030 ( .A(G204GAT), .B(KEYINPUT21), .ZN(new_n168_) );
  NAND2_X1 g031 ( .A1(new_n167_), .A2(new_n168_), .ZN(new_n169_) );
  OR2_X1 g032 ( .A1(new_n167_), .A2(new_n168_), .ZN(new_n170_) );
  NAND2_X1 g033 ( .A1(new_n170_), .A2(new_n169_), .ZN(new_n171_) );
  NAND2_X1 g034 ( .A1(new_n171_), .A2(new_n166_), .ZN(new_n172_) );
  NAND3_X1 g035 ( .A1(new_n170_), .A2(G197GAT), .A3(new_n169_), .ZN(new_n173_) );
  NAND3_X1 g036 ( .A1(new_n172_), .A2(new_n165_), .A3(new_n173_), .ZN(new_n174_) );
  NAND2_X1 g037 ( .A1(new_n172_), .A2(new_n173_), .ZN(new_n175_) );
  NAND2_X1 g038 ( .A1(new_n175_), .A2(new_n141_), .ZN(new_n176_) );
  NAND2_X1 g039 ( .A1(new_n176_), .A2(new_n174_), .ZN(new_n177_) );
  XOR2_X1 g040 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(new_n178_) );
  XNOR2_X1 g041 ( .A(G22GAT), .B(KEYINPUT22), .ZN(new_n179_) );
  XNOR2_X1 g042 ( .A(new_n178_), .B(new_n179_), .ZN(new_n180_) );
  OR2_X1 g043 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n181_) );
  NAND2_X1 g044 ( .A1(G78GAT), .A2(G106GAT), .ZN(new_n182_) );
  NAND2_X1 g045 ( .A1(new_n181_), .A2(new_n182_), .ZN(new_n183_) );
  NAND2_X1 g046 ( .A1(new_n183_), .A2(G148GAT), .ZN(new_n184_) );
  INV_X1 g047 ( .A(G148GAT), .ZN(new_n185_) );
  NAND3_X1 g048 ( .A1(new_n181_), .A2(new_n185_), .A3(new_n182_), .ZN(new_n186_) );
  NAND2_X1 g049 ( .A1(new_n184_), .A2(new_n186_), .ZN(new_n187_) );
  XNOR2_X1 g050 ( .A(new_n180_), .B(new_n187_), .ZN(new_n188_) );
  NAND2_X1 g051 ( .A1(new_n177_), .A2(new_n188_), .ZN(new_n189_) );
  INV_X1 g052 ( .A(new_n188_), .ZN(new_n190_) );
  NAND3_X1 g053 ( .A1(new_n190_), .A2(new_n174_), .A3(new_n176_), .ZN(new_n191_) );
  NAND2_X1 g054 ( .A1(new_n189_), .A2(new_n191_), .ZN(new_n192_) );
  XOR2_X1 g055 ( .A(G50GAT), .B(G162GAT), .Z(new_n193_) );
  INV_X1 g056 ( .A(new_n193_), .ZN(new_n194_) );
  NAND2_X1 g057 ( .A1(new_n192_), .A2(new_n194_), .ZN(new_n195_) );
  NAND3_X1 g058 ( .A1(new_n189_), .A2(new_n191_), .A3(new_n193_), .ZN(new_n196_) );
  NAND2_X1 g059 ( .A1(new_n195_), .A2(new_n196_), .ZN(new_n197_) );
  NAND2_X1 g060 ( .A1(G228GAT), .A2(G233GAT), .ZN(new_n198_) );
  NAND2_X1 g061 ( .A1(new_n197_), .A2(new_n198_), .ZN(new_n199_) );
  NAND4_X1 g062 ( .A1(new_n195_), .A2(G228GAT), .A3(G233GAT), .A4(new_n196_), .ZN(new_n200_) );
  NAND2_X1 g063 ( .A1(new_n199_), .A2(new_n200_), .ZN(new_n201_) );
  INV_X1 g064 ( .A(G15GAT), .ZN(new_n202_) );
  XNOR2_X1 g065 ( .A(new_n148_), .B(new_n202_), .ZN(new_n203_) );
  NAND2_X1 g066 ( .A1(G227GAT), .A2(G233GAT), .ZN(new_n204_) );
  NAND2_X1 g067 ( .A1(new_n203_), .A2(new_n204_), .ZN(new_n205_) );
  OR2_X1 g068 ( .A1(new_n203_), .A2(new_n204_), .ZN(new_n206_) );
  NAND2_X1 g069 ( .A1(new_n206_), .A2(new_n205_), .ZN(new_n207_) );
  XNOR2_X1 g070 ( .A(G176GAT), .B(G183GAT), .ZN(new_n208_) );
  XNOR2_X1 g071 ( .A(G71GAT), .B(KEYINPUT20), .ZN(new_n209_) );
  XOR2_X1 g072 ( .A(new_n208_), .B(new_n209_), .Z(new_n210_) );
  INV_X1 g073 ( .A(new_n210_), .ZN(new_n211_) );
  NAND2_X1 g074 ( .A1(new_n207_), .A2(new_n211_), .ZN(new_n212_) );
  NAND3_X1 g075 ( .A1(new_n206_), .A2(new_n205_), .A3(new_n210_), .ZN(new_n213_) );
  NAND2_X1 g076 ( .A1(new_n212_), .A2(new_n213_), .ZN(new_n214_) );
  XNOR2_X1 g077 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(new_n215_) );
  XNOR2_X1 g078 ( .A(G169GAT), .B(KEYINPUT19), .ZN(new_n216_) );
  XOR2_X1 g079 ( .A(new_n215_), .B(new_n216_), .Z(new_n217_) );
  XOR2_X1 g080 ( .A(G134GAT), .B(G190GAT), .Z(new_n218_) );
  XNOR2_X1 g081 ( .A(G43GAT), .B(G99GAT), .ZN(new_n219_) );
  XNOR2_X1 g082 ( .A(new_n218_), .B(new_n219_), .ZN(new_n220_) );
  XNOR2_X1 g083 ( .A(new_n217_), .B(new_n220_), .ZN(new_n221_) );
  INV_X1 g084 ( .A(new_n221_), .ZN(new_n222_) );
  NAND2_X1 g085 ( .A1(new_n214_), .A2(new_n222_), .ZN(new_n223_) );
  NAND3_X1 g086 ( .A1(new_n212_), .A2(new_n213_), .A3(new_n221_), .ZN(new_n224_) );
  NAND2_X1 g087 ( .A1(new_n223_), .A2(new_n224_), .ZN(new_n225_) );
  NAND2_X1 g088 ( .A1(new_n201_), .A2(new_n225_), .ZN(new_n226_) );
  NAND2_X1 g089 ( .A1(new_n226_), .A2(new_n164_), .ZN(new_n227_) );
  NAND3_X1 g090 ( .A1(new_n201_), .A2(new_n225_), .A3(KEYINPUT26), .ZN(new_n228_) );
  NAND2_X1 g091 ( .A1(new_n227_), .A2(new_n228_), .ZN(new_n229_) );
  INV_X1 g092 ( .A(KEYINPUT27), .ZN(new_n230_) );
  XNOR2_X1 g093 ( .A(G64GAT), .B(G176GAT), .ZN(new_n231_) );
  XNOR2_X1 g094 ( .A(new_n231_), .B(G92GAT), .ZN(new_n232_) );
  NAND2_X1 g095 ( .A1(G226GAT), .A2(G233GAT), .ZN(new_n233_) );
  XNOR2_X1 g096 ( .A(new_n232_), .B(new_n233_), .ZN(new_n234_) );
  XOR2_X1 g097 ( .A(G8GAT), .B(G183GAT), .Z(new_n235_) );
  INV_X1 g098 ( .A(new_n235_), .ZN(new_n236_) );
  NAND2_X1 g099 ( .A1(new_n234_), .A2(new_n236_), .ZN(new_n237_) );
  OR2_X1 g100 ( .A1(new_n234_), .A2(new_n236_), .ZN(new_n238_) );
  NAND2_X1 g101 ( .A1(new_n238_), .A2(new_n237_), .ZN(new_n239_) );
  XNOR2_X1 g102 ( .A(G36GAT), .B(G190GAT), .ZN(new_n240_) );
  NAND3_X1 g103 ( .A1(new_n172_), .A2(new_n173_), .A3(new_n240_), .ZN(new_n241_) );
  INV_X1 g104 ( .A(new_n240_), .ZN(new_n242_) );
  NAND2_X1 g105 ( .A1(new_n175_), .A2(new_n242_), .ZN(new_n243_) );
  NAND2_X1 g106 ( .A1(new_n243_), .A2(new_n241_), .ZN(new_n244_) );
  NAND2_X1 g107 ( .A1(new_n239_), .A2(new_n244_), .ZN(new_n245_) );
  NAND4_X1 g108 ( .A1(new_n238_), .A2(new_n237_), .A3(new_n241_), .A4(new_n243_), .ZN(new_n246_) );
  NAND2_X1 g109 ( .A1(new_n245_), .A2(new_n246_), .ZN(new_n247_) );
  NAND2_X1 g110 ( .A1(new_n247_), .A2(new_n217_), .ZN(new_n248_) );
  INV_X1 g111 ( .A(new_n217_), .ZN(new_n249_) );
  NAND3_X1 g112 ( .A1(new_n245_), .A2(new_n249_), .A3(new_n246_), .ZN(new_n250_) );
  NAND2_X1 g113 ( .A1(new_n248_), .A2(new_n250_), .ZN(new_n251_) );
  XNOR2_X1 g114 ( .A(new_n251_), .B(new_n230_), .ZN(new_n252_) );
  NAND2_X1 g115 ( .A1(new_n229_), .A2(new_n252_), .ZN(new_n253_) );
  INV_X1 g116 ( .A(KEYINPUT25), .ZN(new_n254_) );
  NAND4_X1 g117 ( .A1(new_n223_), .A2(new_n248_), .A3(new_n224_), .A4(new_n250_), .ZN(new_n255_) );
  NAND3_X1 g118 ( .A1(new_n255_), .A2(new_n199_), .A3(new_n200_), .ZN(new_n256_) );
  XNOR2_X1 g119 ( .A(new_n256_), .B(new_n254_), .ZN(new_n257_) );
  NAND2_X1 g120 ( .A1(new_n253_), .A2(new_n257_), .ZN(new_n258_) );
  NAND2_X1 g121 ( .A1(new_n258_), .A2(new_n163_), .ZN(new_n259_) );
  INV_X1 g122 ( .A(KEYINPUT28), .ZN(new_n260_) );
  XNOR2_X1 g123 ( .A(new_n201_), .B(new_n260_), .ZN(new_n261_) );
  INV_X1 g124 ( .A(new_n225_), .ZN(new_n262_) );
  NOR2_X1 g125 ( .A1(new_n163_), .A2(new_n262_), .ZN(new_n263_) );
  NAND3_X1 g126 ( .A1(new_n263_), .A2(new_n252_), .A3(new_n261_), .ZN(new_n264_) );
  NAND2_X1 g127 ( .A1(new_n259_), .A2(new_n264_), .ZN(new_n265_) );
  XNOR2_X1 g128 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(new_n266_) );
  AND2_X1 g129 ( .A1(G232GAT), .A2(G233GAT), .ZN(new_n267_) );
  OR2_X1 g130 ( .A1(new_n266_), .A2(new_n267_), .ZN(new_n268_) );
  NAND2_X1 g131 ( .A1(new_n266_), .A2(new_n267_), .ZN(new_n269_) );
  NAND2_X1 g132 ( .A1(new_n268_), .A2(new_n269_), .ZN(new_n270_) );
  NAND2_X1 g133 ( .A1(new_n270_), .A2(KEYINPUT9), .ZN(new_n271_) );
  INV_X1 g134 ( .A(KEYINPUT9), .ZN(new_n272_) );
  NAND3_X1 g135 ( .A1(new_n268_), .A2(new_n272_), .A3(new_n269_), .ZN(new_n273_) );
  NAND2_X1 g136 ( .A1(new_n271_), .A2(new_n273_), .ZN(new_n274_) );
  OR2_X1 g137 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n275_) );
  NAND2_X1 g138 ( .A1(G43GAT), .A2(KEYINPUT8), .ZN(new_n276_) );
  NAND2_X1 g139 ( .A1(new_n275_), .A2(new_n276_), .ZN(new_n277_) );
  NAND2_X1 g140 ( .A1(new_n277_), .A2(KEYINPUT7), .ZN(new_n278_) );
  INV_X1 g141 ( .A(KEYINPUT7), .ZN(new_n279_) );
  NAND3_X1 g142 ( .A1(new_n275_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_) );
  NAND2_X1 g143 ( .A1(new_n278_), .A2(new_n280_), .ZN(new_n281_) );
  XNOR2_X1 g144 ( .A(G85GAT), .B(G99GAT), .ZN(new_n282_) );
  NAND2_X1 g145 ( .A1(new_n282_), .A2(G92GAT), .ZN(new_n283_) );
  INV_X1 g146 ( .A(G92GAT), .ZN(new_n284_) );
  OR2_X1 g147 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n285_) );
  NAND2_X1 g148 ( .A1(G85GAT), .A2(G99GAT), .ZN(new_n286_) );
  NAND3_X1 g149 ( .A1(new_n285_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_) );
  NAND2_X1 g150 ( .A1(new_n283_), .A2(new_n287_), .ZN(new_n288_) );
  XNOR2_X1 g151 ( .A(new_n281_), .B(new_n288_), .ZN(new_n289_) );
  NAND2_X1 g152 ( .A1(new_n289_), .A2(new_n274_), .ZN(new_n290_) );
  NAND2_X1 g153 ( .A1(new_n281_), .A2(new_n288_), .ZN(new_n291_) );
  OR2_X1 g154 ( .A1(new_n281_), .A2(new_n288_), .ZN(new_n292_) );
  NAND4_X1 g155 ( .A1(new_n292_), .A2(new_n271_), .A3(new_n273_), .A4(new_n291_), .ZN(new_n293_) );
  NAND2_X1 g156 ( .A1(new_n290_), .A2(new_n293_), .ZN(new_n294_) );
  XNOR2_X1 g157 ( .A(G106GAT), .B(G218GAT), .ZN(new_n295_) );
  XOR2_X1 g158 ( .A(new_n151_), .B(new_n295_), .Z(new_n296_) );
  INV_X1 g159 ( .A(new_n296_), .ZN(new_n297_) );
  NAND2_X1 g160 ( .A1(new_n294_), .A2(new_n297_), .ZN(new_n298_) );
  NAND3_X1 g161 ( .A1(new_n290_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n299_) );
  NAND2_X1 g162 ( .A1(new_n298_), .A2(new_n299_), .ZN(new_n300_) );
  NAND2_X1 g163 ( .A1(new_n300_), .A2(new_n193_), .ZN(new_n301_) );
  NAND3_X1 g164 ( .A1(new_n298_), .A2(new_n194_), .A3(new_n299_), .ZN(new_n302_) );
  NAND2_X1 g165 ( .A1(new_n301_), .A2(new_n302_), .ZN(new_n303_) );
  NAND2_X1 g166 ( .A1(new_n303_), .A2(new_n240_), .ZN(new_n304_) );
  NAND3_X1 g167 ( .A1(new_n301_), .A2(new_n242_), .A3(new_n302_), .ZN(new_n305_) );
  XNOR2_X1 g168 ( .A(G57GAT), .B(G71GAT), .ZN(new_n306_) );
  XOR2_X1 g169 ( .A(new_n306_), .B(KEYINPUT13), .Z(new_n307_) );
  XNOR2_X1 g170 ( .A(G15GAT), .B(G22GAT), .ZN(new_n308_) );
  XNOR2_X1 g171 ( .A(new_n308_), .B(new_n138_), .ZN(new_n309_) );
  XNOR2_X1 g172 ( .A(new_n307_), .B(new_n309_), .ZN(new_n310_) );
  XNOR2_X1 g173 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(new_n311_) );
  XNOR2_X1 g174 ( .A(G64GAT), .B(KEYINPUT15), .ZN(new_n312_) );
  XNOR2_X1 g175 ( .A(new_n311_), .B(new_n312_), .ZN(new_n313_) );
  XNOR2_X1 g176 ( .A(G78GAT), .B(G155GAT), .ZN(new_n314_) );
  XNOR2_X1 g177 ( .A(G127GAT), .B(G211GAT), .ZN(new_n315_) );
  XNOR2_X1 g178 ( .A(new_n314_), .B(new_n315_), .ZN(new_n316_) );
  XNOR2_X1 g179 ( .A(new_n313_), .B(new_n316_), .ZN(new_n317_) );
  XNOR2_X1 g180 ( .A(new_n310_), .B(new_n317_), .ZN(new_n318_) );
  XNOR2_X1 g181 ( .A(new_n318_), .B(new_n235_), .ZN(new_n319_) );
  NAND2_X1 g182 ( .A1(G231GAT), .A2(G233GAT), .ZN(new_n320_) );
  XNOR2_X1 g183 ( .A(new_n319_), .B(new_n320_), .ZN(new_n321_) );
  NAND3_X1 g184 ( .A1(new_n321_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n322_) );
  XOR2_X1 g185 ( .A(new_n322_), .B(KEYINPUT16), .Z(new_n323_) );
  AND2_X1 g186 ( .A1(new_n265_), .A2(new_n323_), .ZN(new_n324_) );
  INV_X1 g187 ( .A(new_n231_), .ZN(new_n325_) );
  NAND2_X1 g188 ( .A1(new_n187_), .A2(new_n288_), .ZN(new_n326_) );
  NAND4_X1 g189 ( .A1(new_n184_), .A2(new_n283_), .A3(new_n186_), .A4(new_n287_), .ZN(new_n327_) );
  NAND2_X1 g190 ( .A1(new_n326_), .A2(new_n327_), .ZN(new_n328_) );
  XNOR2_X1 g191 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(new_n329_) );
  NAND2_X1 g192 ( .A1(G230GAT), .A2(G233GAT), .ZN(new_n330_) );
  INV_X1 g193 ( .A(new_n330_), .ZN(new_n331_) );
  NAND2_X1 g194 ( .A1(new_n329_), .A2(new_n331_), .ZN(new_n332_) );
  OR2_X1 g195 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n333_) );
  NAND2_X1 g196 ( .A1(KEYINPUT33), .A2(KEYINPUT31), .ZN(new_n334_) );
  NAND3_X1 g197 ( .A1(new_n333_), .A2(new_n334_), .A3(new_n330_), .ZN(new_n335_) );
  NAND2_X1 g198 ( .A1(new_n332_), .A2(new_n335_), .ZN(new_n336_) );
  NAND2_X1 g199 ( .A1(new_n336_), .A2(KEYINPUT32), .ZN(new_n337_) );
  INV_X1 g200 ( .A(KEYINPUT32), .ZN(new_n338_) );
  NAND3_X1 g201 ( .A1(new_n332_), .A2(new_n338_), .A3(new_n335_), .ZN(new_n339_) );
  NAND2_X1 g202 ( .A1(new_n337_), .A2(new_n339_), .ZN(new_n340_) );
  NAND2_X1 g203 ( .A1(new_n328_), .A2(new_n340_), .ZN(new_n341_) );
  NAND4_X1 g204 ( .A1(new_n326_), .A2(new_n337_), .A3(new_n327_), .A4(new_n339_), .ZN(new_n342_) );
  NAND2_X1 g205 ( .A1(new_n341_), .A2(new_n342_), .ZN(new_n343_) );
  NAND2_X1 g206 ( .A1(new_n343_), .A2(new_n325_), .ZN(new_n344_) );
  NAND3_X1 g207 ( .A1(new_n341_), .A2(new_n231_), .A3(new_n342_), .ZN(new_n345_) );
  NAND2_X1 g208 ( .A1(new_n344_), .A2(new_n345_), .ZN(new_n346_) );
  XNOR2_X1 g209 ( .A(G120GAT), .B(G204GAT), .ZN(new_n347_) );
  NAND2_X1 g210 ( .A1(new_n346_), .A2(new_n347_), .ZN(new_n348_) );
  INV_X1 g211 ( .A(new_n347_), .ZN(new_n349_) );
  NAND3_X1 g212 ( .A1(new_n344_), .A2(new_n345_), .A3(new_n349_), .ZN(new_n350_) );
  NAND2_X1 g213 ( .A1(new_n348_), .A2(new_n350_), .ZN(new_n351_) );
  NAND2_X1 g214 ( .A1(new_n351_), .A2(new_n307_), .ZN(new_n352_) );
  INV_X1 g215 ( .A(new_n307_), .ZN(new_n353_) );
  NAND3_X1 g216 ( .A1(new_n348_), .A2(new_n353_), .A3(new_n350_), .ZN(new_n354_) );
  NAND2_X1 g217 ( .A1(new_n352_), .A2(new_n354_), .ZN(new_n355_) );
  XOR2_X1 g218 ( .A(new_n309_), .B(new_n281_), .Z(new_n356_) );
  XNOR2_X1 g219 ( .A(G8GAT), .B(G169GAT), .ZN(new_n357_) );
  XNOR2_X1 g220 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(new_n358_) );
  XNOR2_X1 g221 ( .A(new_n357_), .B(new_n358_), .ZN(new_n359_) );
  XNOR2_X1 g222 ( .A(G113GAT), .B(G197GAT), .ZN(new_n360_) );
  XNOR2_X1 g223 ( .A(G29GAT), .B(G141GAT), .ZN(new_n361_) );
  XNOR2_X1 g224 ( .A(new_n360_), .B(new_n361_), .ZN(new_n362_) );
  XNOR2_X1 g225 ( .A(new_n359_), .B(new_n362_), .ZN(new_n363_) );
  XNOR2_X1 g226 ( .A(new_n356_), .B(new_n363_), .ZN(new_n364_) );
  XNOR2_X1 g227 ( .A(G36GAT), .B(G50GAT), .ZN(new_n365_) );
  NAND2_X1 g228 ( .A1(G229GAT), .A2(G233GAT), .ZN(new_n366_) );
  XOR2_X1 g229 ( .A(new_n365_), .B(new_n366_), .Z(new_n367_) );
  XNOR2_X1 g230 ( .A(new_n364_), .B(new_n367_), .ZN(new_n368_) );
  AND2_X1 g231 ( .A1(new_n355_), .A2(new_n368_), .ZN(new_n369_) );
  NAND2_X1 g232 ( .A1(new_n324_), .A2(new_n369_), .ZN(new_n370_) );
  NOR2_X1 g233 ( .A1(new_n370_), .A2(new_n163_), .ZN(new_n371_) );
  XNOR2_X1 g234 ( .A(new_n371_), .B(KEYINPUT34), .ZN(new_n372_) );
  XNOR2_X1 g235 ( .A(new_n372_), .B(new_n138_), .ZN(G1324GAT) );
  INV_X1 g236 ( .A(new_n251_), .ZN(new_n374_) );
  INV_X1 g237 ( .A(new_n370_), .ZN(new_n375_) );
  NAND2_X1 g238 ( .A1(new_n375_), .A2(new_n374_), .ZN(new_n376_) );
  XNOR2_X1 g239 ( .A(new_n376_), .B(G8GAT), .ZN(G1325GAT) );
  NOR2_X1 g240 ( .A1(new_n370_), .A2(new_n225_), .ZN(new_n378_) );
  XNOR2_X1 g241 ( .A(G15GAT), .B(KEYINPUT35), .ZN(new_n379_) );
  XNOR2_X1 g242 ( .A(new_n378_), .B(new_n379_), .ZN(G1326GAT) );
  INV_X1 g243 ( .A(new_n261_), .ZN(new_n381_) );
  NAND2_X1 g244 ( .A1(new_n375_), .A2(new_n381_), .ZN(new_n382_) );
  XNOR2_X1 g245 ( .A(new_n382_), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 g246 ( .A(KEYINPUT38), .ZN(new_n384_) );
  INV_X1 g247 ( .A(KEYINPUT36), .ZN(new_n385_) );
  NAND2_X1 g248 ( .A1(new_n304_), .A2(new_n305_), .ZN(new_n386_) );
  NAND2_X1 g249 ( .A1(new_n386_), .A2(new_n385_), .ZN(new_n387_) );
  NAND3_X1 g250 ( .A1(new_n304_), .A2(KEYINPUT36), .A3(new_n305_), .ZN(new_n388_) );
  NAND2_X1 g251 ( .A1(new_n387_), .A2(new_n388_), .ZN(new_n389_) );
  NOR2_X1 g252 ( .A1(new_n389_), .A2(new_n321_), .ZN(new_n390_) );
  NAND2_X1 g253 ( .A1(new_n265_), .A2(new_n390_), .ZN(new_n391_) );
  NAND2_X1 g254 ( .A1(new_n391_), .A2(KEYINPUT37), .ZN(new_n392_) );
  INV_X1 g255 ( .A(KEYINPUT37), .ZN(new_n393_) );
  NAND3_X1 g256 ( .A1(new_n265_), .A2(new_n393_), .A3(new_n390_), .ZN(new_n394_) );
  NAND2_X1 g257 ( .A1(new_n392_), .A2(new_n394_), .ZN(new_n395_) );
  NAND2_X1 g258 ( .A1(new_n395_), .A2(new_n369_), .ZN(new_n396_) );
  NAND2_X1 g259 ( .A1(new_n396_), .A2(new_n384_), .ZN(new_n397_) );
  NAND3_X1 g260 ( .A1(new_n395_), .A2(KEYINPUT38), .A3(new_n369_), .ZN(new_n398_) );
  NAND2_X1 g261 ( .A1(new_n397_), .A2(new_n398_), .ZN(new_n399_) );
  INV_X1 g262 ( .A(new_n399_), .ZN(new_n400_) );
  NOR2_X1 g263 ( .A1(new_n400_), .A2(new_n163_), .ZN(new_n401_) );
  XNOR2_X1 g264 ( .A(G29GAT), .B(KEYINPUT39), .ZN(new_n402_) );
  XNOR2_X1 g265 ( .A(new_n401_), .B(new_n402_), .ZN(G1328GAT) );
  NAND2_X1 g266 ( .A1(new_n399_), .A2(new_n374_), .ZN(new_n404_) );
  XNOR2_X1 g267 ( .A(new_n404_), .B(G36GAT), .ZN(G1329GAT) );
  INV_X1 g268 ( .A(G43GAT), .ZN(new_n406_) );
  INV_X1 g269 ( .A(KEYINPUT40), .ZN(new_n407_) );
  NAND2_X1 g270 ( .A1(new_n399_), .A2(new_n262_), .ZN(new_n408_) );
  NAND2_X1 g271 ( .A1(new_n408_), .A2(new_n407_), .ZN(new_n409_) );
  NAND3_X1 g272 ( .A1(new_n399_), .A2(KEYINPUT40), .A3(new_n262_), .ZN(new_n410_) );
  NAND2_X1 g273 ( .A1(new_n409_), .A2(new_n410_), .ZN(new_n411_) );
  NAND2_X1 g274 ( .A1(new_n411_), .A2(new_n406_), .ZN(new_n412_) );
  NAND3_X1 g275 ( .A1(new_n409_), .A2(G43GAT), .A3(new_n410_), .ZN(new_n413_) );
  NAND2_X1 g276 ( .A1(new_n412_), .A2(new_n413_), .ZN(G1330GAT) );
  NAND2_X1 g277 ( .A1(new_n399_), .A2(new_n381_), .ZN(new_n415_) );
  XNOR2_X1 g278 ( .A(new_n415_), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 g279 ( .A(KEYINPUT41), .ZN(new_n417_) );
  NAND2_X1 g280 ( .A1(new_n355_), .A2(new_n417_), .ZN(new_n418_) );
  NAND3_X1 g281 ( .A1(new_n352_), .A2(KEYINPUT41), .A3(new_n354_), .ZN(new_n419_) );
  NAND2_X1 g282 ( .A1(new_n418_), .A2(new_n419_), .ZN(new_n420_) );
  NOR2_X1 g283 ( .A1(new_n420_), .A2(new_n368_), .ZN(new_n421_) );
  NAND2_X1 g284 ( .A1(new_n324_), .A2(new_n421_), .ZN(new_n422_) );
  NOR2_X1 g285 ( .A1(new_n422_), .A2(new_n163_), .ZN(new_n423_) );
  XOR2_X1 g286 ( .A(G57GAT), .B(KEYINPUT42), .Z(new_n424_) );
  XNOR2_X1 g287 ( .A(new_n423_), .B(new_n424_), .ZN(G1332GAT) );
  INV_X1 g288 ( .A(new_n422_), .ZN(new_n426_) );
  NAND2_X1 g289 ( .A1(new_n426_), .A2(new_n374_), .ZN(new_n427_) );
  XNOR2_X1 g290 ( .A(new_n427_), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 g291 ( .A1(new_n426_), .A2(new_n262_), .ZN(new_n429_) );
  XNOR2_X1 g292 ( .A(new_n429_), .B(G71GAT), .ZN(G1334GAT) );
  NOR2_X1 g293 ( .A1(new_n422_), .A2(new_n261_), .ZN(new_n431_) );
  XNOR2_X1 g294 ( .A(G78GAT), .B(KEYINPUT43), .ZN(new_n432_) );
  XNOR2_X1 g295 ( .A(new_n431_), .B(new_n432_), .ZN(G1335GAT) );
  NAND2_X1 g296 ( .A1(new_n395_), .A2(new_n421_), .ZN(new_n434_) );
  NOR2_X1 g297 ( .A1(new_n434_), .A2(new_n163_), .ZN(new_n435_) );
  XOR2_X1 g298 ( .A(new_n435_), .B(G85GAT), .Z(G1336GAT) );
  NOR2_X1 g299 ( .A1(new_n434_), .A2(new_n251_), .ZN(new_n437_) );
  XNOR2_X1 g300 ( .A(new_n437_), .B(new_n284_), .ZN(G1337GAT) );
  NOR2_X1 g301 ( .A1(new_n434_), .A2(new_n225_), .ZN(new_n439_) );
  XOR2_X1 g302 ( .A(new_n439_), .B(G99GAT), .Z(G1338GAT) );
  NOR2_X1 g303 ( .A1(new_n434_), .A2(new_n261_), .ZN(new_n441_) );
  XNOR2_X1 g304 ( .A(new_n441_), .B(KEYINPUT44), .ZN(new_n442_) );
  XOR2_X1 g305 ( .A(new_n442_), .B(G106GAT), .Z(G1339GAT) );
  INV_X1 g306 ( .A(KEYINPUT47), .ZN(new_n444_) );
  NAND4_X1 g307 ( .A1(new_n418_), .A2(KEYINPUT46), .A3(new_n368_), .A4(new_n419_), .ZN(new_n445_) );
  INV_X1 g308 ( .A(KEYINPUT46), .ZN(new_n446_) );
  NAND3_X1 g309 ( .A1(new_n418_), .A2(new_n368_), .A3(new_n419_), .ZN(new_n447_) );
  NAND2_X1 g310 ( .A1(new_n447_), .A2(new_n446_), .ZN(new_n448_) );
  NOR2_X1 g311 ( .A1(new_n321_), .A2(new_n386_), .ZN(new_n449_) );
  NAND4_X1 g312 ( .A1(new_n448_), .A2(new_n444_), .A3(new_n445_), .A4(new_n449_), .ZN(new_n450_) );
  INV_X1 g313 ( .A(KEYINPUT45), .ZN(new_n451_) );
  NAND4_X1 g314 ( .A1(new_n387_), .A2(new_n321_), .A3(new_n451_), .A4(new_n388_), .ZN(new_n452_) );
  NAND3_X1 g315 ( .A1(new_n387_), .A2(new_n321_), .A3(new_n388_), .ZN(new_n453_) );
  NAND2_X1 g316 ( .A1(new_n453_), .A2(KEYINPUT45), .ZN(new_n454_) );
  INV_X1 g317 ( .A(new_n355_), .ZN(new_n455_) );
  NOR2_X1 g318 ( .A1(new_n455_), .A2(new_n368_), .ZN(new_n456_) );
  NAND3_X1 g319 ( .A1(new_n454_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_) );
  NAND3_X1 g320 ( .A1(new_n448_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n458_) );
  NAND2_X1 g321 ( .A1(new_n458_), .A2(KEYINPUT47), .ZN(new_n459_) );
  NAND4_X1 g322 ( .A1(new_n459_), .A2(new_n457_), .A3(KEYINPUT48), .A4(new_n450_), .ZN(new_n460_) );
  INV_X1 g323 ( .A(KEYINPUT48), .ZN(new_n461_) );
  NAND3_X1 g324 ( .A1(new_n459_), .A2(new_n450_), .A3(new_n457_), .ZN(new_n462_) );
  NAND2_X1 g325 ( .A1(new_n462_), .A2(new_n461_), .ZN(new_n463_) );
  INV_X1 g326 ( .A(new_n252_), .ZN(new_n464_) );
  NOR2_X1 g327 ( .A1(new_n163_), .A2(new_n464_), .ZN(new_n465_) );
  AND3_X1 g328 ( .A1(new_n463_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n466_) );
  AND3_X1 g329 ( .A1(new_n466_), .A2(new_n262_), .A3(new_n261_), .ZN(new_n467_) );
  NAND2_X1 g330 ( .A1(new_n467_), .A2(new_n368_), .ZN(new_n468_) );
  XNOR2_X1 g331 ( .A(new_n468_), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 g332 ( .A(new_n420_), .ZN(new_n470_) );
  NAND2_X1 g333 ( .A1(new_n467_), .A2(new_n470_), .ZN(new_n471_) );
  XOR2_X1 g334 ( .A(G120GAT), .B(KEYINPUT49), .Z(new_n472_) );
  XNOR2_X1 g335 ( .A(new_n471_), .B(new_n472_), .ZN(G1341GAT) );
  NAND2_X1 g336 ( .A1(new_n467_), .A2(new_n321_), .ZN(new_n474_) );
  XNOR2_X1 g337 ( .A(new_n474_), .B(KEYINPUT50), .ZN(new_n475_) );
  XNOR2_X1 g338 ( .A(new_n475_), .B(G127GAT), .ZN(G1342GAT) );
  NAND2_X1 g339 ( .A1(new_n467_), .A2(new_n386_), .ZN(new_n477_) );
  XOR2_X1 g340 ( .A(G134GAT), .B(KEYINPUT51), .Z(new_n478_) );
  XNOR2_X1 g341 ( .A(new_n477_), .B(new_n478_), .ZN(G1343GAT) );
  AND2_X1 g342 ( .A1(new_n466_), .A2(new_n229_), .ZN(new_n480_) );
  NAND2_X1 g343 ( .A1(new_n480_), .A2(new_n368_), .ZN(new_n481_) );
  XNOR2_X1 g344 ( .A(new_n481_), .B(G141GAT), .ZN(G1344GAT) );
  NAND2_X1 g345 ( .A1(new_n480_), .A2(new_n470_), .ZN(new_n483_) );
  XNOR2_X1 g346 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(new_n484_) );
  XNOR2_X1 g347 ( .A(new_n483_), .B(new_n484_), .ZN(new_n485_) );
  XNOR2_X1 g348 ( .A(new_n485_), .B(new_n185_), .ZN(G1345GAT) );
  NAND2_X1 g349 ( .A1(new_n480_), .A2(new_n321_), .ZN(new_n487_) );
  XNOR2_X1 g350 ( .A(new_n487_), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 g351 ( .A1(new_n480_), .A2(new_n386_), .ZN(new_n489_) );
  XNOR2_X1 g352 ( .A(new_n489_), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 g353 ( .A(new_n201_), .ZN(new_n491_) );
  NAND3_X1 g354 ( .A1(new_n463_), .A2(new_n374_), .A3(new_n460_), .ZN(new_n492_) );
  NAND2_X1 g355 ( .A1(new_n492_), .A2(KEYINPUT54), .ZN(new_n493_) );
  INV_X1 g356 ( .A(KEYINPUT54), .ZN(new_n494_) );
  NAND4_X1 g357 ( .A1(new_n463_), .A2(new_n494_), .A3(new_n374_), .A4(new_n460_), .ZN(new_n495_) );
  NAND4_X1 g358 ( .A1(new_n493_), .A2(new_n163_), .A3(new_n491_), .A4(new_n495_), .ZN(new_n496_) );
  NAND2_X1 g359 ( .A1(new_n496_), .A2(KEYINPUT55), .ZN(new_n497_) );
  INV_X1 g360 ( .A(KEYINPUT55), .ZN(new_n498_) );
  AND2_X1 g361 ( .A1(new_n495_), .A2(new_n491_), .ZN(new_n499_) );
  NAND4_X1 g362 ( .A1(new_n499_), .A2(new_n498_), .A3(new_n163_), .A4(new_n493_), .ZN(new_n500_) );
  NAND2_X1 g363 ( .A1(new_n497_), .A2(new_n500_), .ZN(new_n501_) );
  AND2_X1 g364 ( .A1(new_n501_), .A2(new_n262_), .ZN(new_n502_) );
  NAND2_X1 g365 ( .A1(new_n502_), .A2(new_n368_), .ZN(new_n503_) );
  XNOR2_X1 g366 ( .A(new_n503_), .B(G169GAT), .ZN(G1348GAT) );
  INV_X1 g367 ( .A(G176GAT), .ZN(new_n505_) );
  NAND3_X1 g368 ( .A1(new_n501_), .A2(new_n262_), .A3(new_n470_), .ZN(new_n506_) );
  XNOR2_X1 g369 ( .A(KEYINPUT57), .B(KEYINPUT56), .ZN(new_n507_) );
  NAND2_X1 g370 ( .A1(new_n506_), .A2(new_n507_), .ZN(new_n508_) );
  INV_X1 g371 ( .A(new_n507_), .ZN(new_n509_) );
  NAND4_X1 g372 ( .A1(new_n501_), .A2(new_n262_), .A3(new_n470_), .A4(new_n509_), .ZN(new_n510_) );
  NAND2_X1 g373 ( .A1(new_n508_), .A2(new_n510_), .ZN(new_n511_) );
  NAND2_X1 g374 ( .A1(new_n511_), .A2(new_n505_), .ZN(new_n512_) );
  NAND3_X1 g375 ( .A1(new_n508_), .A2(G176GAT), .A3(new_n510_), .ZN(new_n513_) );
  NAND2_X1 g376 ( .A1(new_n512_), .A2(new_n513_), .ZN(G1349GAT) );
  NAND2_X1 g377 ( .A1(new_n502_), .A2(new_n321_), .ZN(new_n515_) );
  XNOR2_X1 g378 ( .A(new_n515_), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 g379 ( .A1(new_n502_), .A2(new_n386_), .ZN(new_n517_) );
  XNOR2_X1 g380 ( .A(G190GAT), .B(KEYINPUT58), .ZN(new_n518_) );
  XNOR2_X1 g381 ( .A(new_n517_), .B(new_n518_), .ZN(G1351GAT) );
  AND2_X1 g382 ( .A1(new_n493_), .A2(new_n163_), .ZN(new_n520_) );
  AND2_X1 g383 ( .A1(new_n495_), .A2(new_n229_), .ZN(new_n521_) );
  AND2_X1 g384 ( .A1(new_n520_), .A2(new_n521_), .ZN(new_n522_) );
  NAND2_X1 g385 ( .A1(new_n522_), .A2(new_n368_), .ZN(new_n523_) );
  XNOR2_X1 g386 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(new_n524_) );
  XNOR2_X1 g387 ( .A(new_n523_), .B(new_n524_), .ZN(new_n525_) );
  NAND2_X1 g388 ( .A1(new_n525_), .A2(new_n166_), .ZN(new_n526_) );
  NAND2_X1 g389 ( .A1(new_n523_), .A2(new_n524_), .ZN(new_n527_) );
  OR2_X1 g390 ( .A1(new_n523_), .A2(new_n524_), .ZN(new_n528_) );
  NAND3_X1 g391 ( .A1(new_n528_), .A2(G197GAT), .A3(new_n527_), .ZN(new_n529_) );
  NAND2_X1 g392 ( .A1(new_n526_), .A2(new_n529_), .ZN(G1352GAT) );
  NAND2_X1 g393 ( .A1(new_n522_), .A2(new_n455_), .ZN(new_n531_) );
  XOR2_X1 g394 ( .A(G204GAT), .B(KEYINPUT61), .Z(new_n532_) );
  XNOR2_X1 g395 ( .A(new_n531_), .B(new_n532_), .ZN(G1353GAT) );
  NAND2_X1 g396 ( .A1(new_n522_), .A2(new_n321_), .ZN(new_n534_) );
  XNOR2_X1 g397 ( .A(new_n534_), .B(G211GAT), .ZN(G1354GAT) );
  NAND4_X1 g398 ( .A1(new_n520_), .A2(new_n387_), .A3(new_n388_), .A4(new_n521_), .ZN(new_n536_) );
  XNOR2_X1 g399 ( .A(new_n536_), .B(KEYINPUT62), .ZN(new_n537_) );
  XNOR2_X1 g400 ( .A(new_n537_), .B(G218GAT), .ZN(G1355GAT) );
endmodule


