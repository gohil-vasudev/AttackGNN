module s38417 ( CK, g1249, g16297, g16355, g16399, g16437, g16496, g1943, 
        g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g2637, 
        g27380, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, 
        g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, 
        g3231, g3232, g3233, g3234, g3993, g4088, g4090, g4200, g4321, g4323, 
        g4450, g4590, g51, g5388, g5437, g5472, g5511, g5549, g5555, g5595, 
        g5612, g5629, g563, g5637, g5648, g5657, g5686, g5695, g5738, g5747, 
        g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, 
        g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, 
        g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, 
        g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, 
        g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, 
        g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, 
        g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, test_se, 
        test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, test_si4, 
        test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, test_so7, 
        test_si8, test_so8, test_si9, test_so9, test_si10, test_so10, 
        test_si11, test_so11, test_si12, test_so12, test_si13, test_so13, 
        test_si14, test_so14, test_si15, test_so15, test_si16, test_so16, 
        test_si17, test_so17, test_si18, test_so18, test_si19, test_so19, 
        test_si20, test_so20, test_si21, test_so21, test_si22, test_so22, 
        test_si23, test_so23, test_si24, test_so24, test_si25, test_so25, 
        test_si26, test_so26, test_si27, test_so27, test_si28, test_so28, 
        test_si29, test_so29, test_si30, test_so30, test_si31, test_so31, 
        test_si32, test_so32, test_si33, test_so33, test_si34, test_so34, 
        test_si35, test_so35, test_si36, test_so36, test_si37, test_so37, 
        test_si38, test_so38, test_si39, test_so39, test_si40, test_so40, 
        test_si41, test_so41, test_si42, test_so42, test_si43, test_so43, 
        test_si44, test_so44, test_si45, test_so45, test_si46, test_so46, 
        test_si47, test_so47, test_si48, test_so48, test_si49, test_so49, 
        test_si50, test_so50, test_si51, test_so51, test_si52, test_so52, 
        test_si53, test_so53, test_si54, test_so54, test_si55, test_so55, 
        test_si56, test_so56, test_si57, test_so57, test_si58, test_so58, 
        test_si59, test_so59, test_si60, test_so60, test_si61, test_so61, 
        test_si62, test_so62, test_si63, test_so63, test_si64, test_so64, 
        test_si65, test_so65, test_si66, test_so66, test_si67, test_so67, 
        test_si68, test_so68, test_si69, test_so69, test_si70, test_so70, 
        test_si71, test_so71, test_si72, test_so72, test_si73, test_so73, 
        test_si74, test_so74, test_si75, test_so75, test_si76, test_so76, 
        test_si77, test_so77, test_si78, test_so78, test_si79, test_so79, 
        test_si80, test_so80, test_si81, test_so81, test_si82, test_so82, 
        test_si83, test_so83, test_si84, test_so84, test_si85, test_so85, 
        test_si86, test_so86, test_si87, test_so87, test_si88, test_so88, 
        test_si89, test_so89, test_si90, test_so90, test_si91, test_so91, 
        test_si92, test_so92, test_si93, test_so93, test_si94, test_so94, 
        test_si95, test_so95, test_si96, test_so96, test_si97, test_so97, 
        test_si98, test_so98, test_si99, test_so99, test_si100, test_so100 );
  input CK, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217,
         g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227,
         g3228, g3229, g3230, g3231, g3232, g3233, g3234, g51, g563, test_se,
         test_si1, test_si2, test_si3, test_si4, test_si5, test_si6, test_si7,
         test_si8, test_si9, test_si10, test_si11, test_si12, test_si13,
         test_si14, test_si15, test_si16, test_si17, test_si18, test_si19,
         test_si20, test_si21, test_si22, test_si23, test_si24, test_si25,
         test_si26, test_si27, test_si28, test_si29, test_si30, test_si31,
         test_si32, test_si33, test_si34, test_si35, test_si36, test_si37,
         test_si38, test_si39, test_si40, test_si41, test_si42, test_si43,
         test_si44, test_si45, test_si46, test_si47, test_si48, test_si49,
         test_si50, test_si51, test_si52, test_si53, test_si54, test_si55,
         test_si56, test_si57, test_si58, test_si59, test_si60, test_si61,
         test_si62, test_si63, test_si64, test_si65, test_si66, test_si67,
         test_si68, test_si69, test_si70, test_si71, test_si72, test_si73,
         test_si74, test_si75, test_si76, test_si77, test_si78, test_si79,
         test_si80, test_si81, test_si82, test_si83, test_si84, test_si85,
         test_si86, test_si87, test_si88, test_si89, test_si90, test_si91,
         test_si92, test_si93, test_si94, test_si95, test_si96, test_si97,
         test_si98, test_si99, test_si100;
  output g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435,
         g25442, g25489, g26104, g26135, g26149, g27380, g3993, g4088, g4090,
         g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549,
         g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738,
         g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518,
         g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944,
         g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334,
         g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012,
         g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249,
         g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266,
         g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275,
         test_so1, test_so2, test_so3, test_so4, test_so5, test_so6, test_so7,
         test_so8, test_so9, test_so10, test_so11, test_so12, test_so13,
         test_so14, test_so15, test_so16, test_so17, test_so18, test_so19,
         test_so20, test_so21, test_so22, test_so23, test_so24, test_so25,
         test_so26, test_so27, test_so28, test_so29, test_so30, test_so31,
         test_so32, test_so33, test_so34, test_so35, test_so36, test_so37,
         test_so38, test_so39, test_so40, test_so41, test_so42, test_so43,
         test_so44, test_so45, test_so46, test_so47, test_so48, test_so49,
         test_so50, test_so51, test_so52, test_so53, test_so54, test_so55,
         test_so56, test_so57, test_so58, test_so59, test_so60, test_so61,
         test_so62, test_so63, test_so64, test_so65, test_so66, test_so67,
         test_so68, test_so69, test_so70, test_so71, test_so72, test_so73,
         test_so74, test_so75, test_so76, test_so77, test_so78, test_so79,
         test_so80, test_so81, test_so82, test_so83, test_so84, test_so85,
         test_so86, test_so87, test_so88, test_so89, test_so90, test_so91,
         test_so92, test_so93, test_so94, test_so95, test_so96, test_so97,
         test_so98, test_so99, test_so100;
  wire   test_so3, test_so4, test_so5, test_so23, test_so57, test_so63,
         test_so73, test_so99, test_so100, n2230, n2217, n2231, n2374, n2361,
         n2375, DFF_2_n1, n4264, n2445, n2446, n2440, n2426, n2670, n2671,
         n2669, n2685, n2686, n2684, n2718, n2719, n2717, n2982, g2124, n2981,
         n2985, g1430, n2984, n2988, g744, n2987, n2991, g56, n2990, n3742,
         n3741, n8104, g16802, n8103, DFF_1_n1, g16823, n8102, g2950, n4423,
         n4274, g2883, n4330, g22026, g2888, g2896, n4431, g24473, g2892,
         g2903, n4305, g26037, g2900, n4291, g26798, g2908, n4355, n4273,
         g2912, n4482, g23357, g2917, n4479, g24476, g2924, n4349, g25199,
         g2920, n4280, DFF_15_n1, n4281, n8099, DFF_16_n1, n8098, DFF_18_n1,
         n4279, g2879, n4351, g2934, g2935, g2938, g2941, g2944, g2947, g2953,
         g2956, g2959, g2962, g2963, g2969, g2972, g2975, g2978, g2981, g2874,
         g18754, g1506, n4288, g18781, g1501, n4565, g18803, g1496, n4557,
         g18821, g1491, n4326, g18835, g1486, n4390, g18852, g1481, n4320,
         g18866, g1476, n4374, g18883, g1471, n4378, g21880, g2877, g19154,
         g813, n4289, g19163, g809, n4567, g19173, g805, n4559, g19184, g801,
         n4327, g20310, g797, n4391, g20343, g793, n4321, g20376, g789, n4375,
         g20417, g785, n4379, g21878, g2873, g19153, g125, n4290, g19162, g121,
         n4569, g19172, g117, n4561, g19144, g113, n4328, g19149, g109, n4392,
         g19157, g105, n4322, g19167, g101, n4376, g19178, g97, n4380, g20874,
         g2857, g18885, g2200, n4287, g18975, g2195, n4563, g18968, g2190,
         n4555, g18942, g2185, n4325, g18906, g2180, n4389, g18867, g2175,
         n4319, g18836, g2170, n4373, g18957, g2165, n4377, g21882, g2878,
         n4598, n4382, n4383, g3109, n4494, g18669, g18719, g3211, g18782,
         g3084, n4445, g17222, g3085, n4340, g17225, g3086, n4337, g17234,
         g3087, n4344, g17224, g3091, n4448, g17228, g3092, n4451, g17246,
         g3093, g17226, g3094, g17235, g3095, n4439, g17269, g3096, n4336,
         g25450, g3097, n4433, g25451, g3098, n4434, g25452, g3099, n4443,
         g28420, g3100, n4342, g28421, g28425, g3102, n4343, g29936, g3103,
         n4447, g29939, g3104, n4452, g29941, g3105, g30796, g3106, n4438,
         g30798, g3107, n4437, g30801, g3108, n4334, g17229, g3155, g17247,
         g3158, n4436, g17302, g3161, g17236, g3164, n4339, g17270, g3167,
         n4348, g17340, g3170, n4441, g17248, g3173, n4338, g17303, g3176,
         n4450, g17383, g17271, g3182, n4453, g17341, g3185, n4442, g17429,
         g3088, n4341, n8090, n8089, g3197, n8088, g3201, n4406, g3204, g3207,
         n4329, g3188, n4405, g3133, n8087, DFF_140_n1, g3128, n8086, n8084,
         g3124, n8083, DFF_146_n1, n8082, n8081, n8080, g3112, g3110, g3111,
         n8079, n8078, n8077, DFF_155_n1, n8076, DFF_156_n1, g3151, n4424,
         g3142, n4301, g185, n4384, n4318, n4512, g165, n4369, g22100, g130,
         g22122, g131, g22141, g129, g22123, g133, g22142, g134, g22161, g132,
         g22025, g142, g22027, g143, g22030, g141, g22028, g145, g22031, g146,
         g22037, g22032, g148, g22038, g149, g22047, g147, g22039, g151,
         g22048, g152, g22063, g150, g22049, g154, g22064, g155, g22079, g153,
         g22065, g157, g22080, g158, g22101, g156, g22081, g160, g22102, g161,
         g22124, g159, g22103, g22125, g164, g22143, g162, g25204, g169,
         g25206, g170, g25211, g168, g25207, g172, g25212, g173, g25218, g171,
         g25213, g175, g25219, g176, g25228, g174, g25220, g178, g25229, g179,
         g25239, g177, g30261, g186, g30267, g30275, g192, g30637, g231,
         g30640, g234, g30645, g237, g30668, g195, g30674, g198, g30680, g201,
         g30641, g240, g30646, g243, g30653, g246, g30276, g204, g30284, g207,
         g30292, g210, g30254, g249, g30257, g252, g30262, g30245, g213,
         g30246, g216, g30248, g219, g30258, g258, g30263, g261, g30268, g264,
         g30635, g222, g30636, g225, g30639, g228, g30661, g267, g30669, g270,
         g30675, g273, g25027, g92, g88, g26529, g83, g27594, g74, g28145, g70,
         g28634, g65, g29109, g61, g29353, g29579, g52, g180, g181, n4506,
         g309, n4388, g27253, g354, g27255, g343, g27258, g27256, g369, g27259,
         g358, g27265, g361, g27260, g384, g27266, g373, g27277, g376, g27267,
         g398, g27278, g388, g27293, g391, g28732, g408, g28735, g411, g28744,
         g414, g29194, g417, g29197, g420, g29201, g423, g28736, g28745, g428,
         g28754, g426, g26803, g429, g26804, g432, g26807, g435, g26805, g438,
         g26808, g441, g26812, g444, g27759, g448, g27760, g449, g27762, g447,
         g29606, g312, g29608, g313, g29611, g314, g30699, g315, g30700,
         g30702, g317, g30455, g318, g30468, g319, g30482, g320, g29167, g322,
         g29169, g323, g29172, g321, g26655, g403, g26659, g404, g26664, g402,
         g450, n8066, DFF_299_n1, g452, n8065, DFF_301_n1, g454, DFF_303_n1,
         g280, n8062, DFF_305_n1, g282, n8061, DFF_307_n1, g284, n8060,
         DFF_309_n1, g286, n8059, DFF_311_n1, g288, n8058, DFF_313_n1, g290,
         n8057, n4485, n4282, n8056, g21346, g305, n4278, n8055, DFF_328_n1,
         g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368,
         g372, g379, g380, g381, g383, g387, g394, g395, g396, g397, g324,
         g337, n4298, n4372, g550, n4313, g554, g18678, g557, n4360, g18726,
         g513, g523, g524, g455, g564, g569, g458, g570, g571, g461, g572,
         g573, g465, g574, g565, g566, g567, g471, g568, g489, n4461, g485,
         n4466, g23067, g486, g23093, g487, g23117, g488, g23385, g23399,
         g24174, g24178, g477, g24207, g478, g24216, g479, g23092, g480,
         g23000, g484, g23022, g464, g24206, g24215, g24228, g528, g535, g542,
         g13149, g543, g544, g21851, g548, g13111, g549, g499, n4541, g13160,
         g558, g559, g27261, g576, g27268, g577, g27279, g575, g27269, g579,
         g27280, g27294, g578, g27281, g582, g27295, g583, g27311, g581,
         g27296, g585, g27312, g586, g27327, g584, g24491, g587, g24498, g590,
         g24507, g593, g24499, g596, g24508, g599, g24519, g602, g28345, g614,
         g28349, g617, g28353, g28342, g605, g28344, g608, g28348, g611,
         g26541, g490, g26545, g493, g26553, g496, g506, n4570, g22578, n4571,
         g525, n8047, n8046, DFF_445_n1, n8045, DFF_446_n1, n8044, n8043, g536,
         g537, g24059, g538, n4492, n8040, n4359, g629, n4295, g16654, g630,
         g20314, g659, g20682, g640, n4404, g23136, g633, n4478, g23324, g653,
         n4422, g24426, g646, n4414, g25185, g660, n4403, g26660, g672, n4413,
         g26776, g27672, g679, n4477, g686, n4396, g28668, g692, n4418, g20875,
         g699, g20879, g700, g20891, g698, g20880, g702, g20892, g703, g20901,
         g701, g20893, g705, g20902, g706, g20921, g704, g20903, g708, g20922,
         g709, g20944, g707, g20923, g20945, g712, g20966, g710, g20946, g714,
         g20967, g715, g20989, g713, g20968, g717, g20990, g718, g21009, g716,
         g20991, g720, g21010, g721, g21031, g719, g21011, g723, g21032, g724,
         g21051, g722, g20876, g726, g20881, g20894, g725, g20924, g729,
         g20947, g730, g20969, g728, g20948, g732, g20970, g733, g20992, g731,
         g25260, g735, g25262, g736, g25266, g734, g738, g22231, g739, g22242,
         g737, n4323, n4312, g22126, g818, g22145, g819, g22162, g817, g22146,
         g821, g22163, g822, g22177, g820, g22029, g830, g22033, g831, g22040,
         g829, g22034, g833, g22041, g834, g22054, g832, g22042, g836, g22055,
         g837, g22066, g835, g22056, g22067, g840, g22087, g838, g22068, g842,
         g22088, g843, g22104, g841, g22089, g845, g22105, g846, g22127, g844,
         g22106, g848, g22128, g849, g22147, g847, g22129, g851, g22148, g852,
         g22164, g850, g25209, g857, g25214, g25221, g856, g25215, g860,
         g25222, g861, g25230, g859, g25223, g863, g25231, g864, g25240, g862,
         g25232, g866, g25241, g867, g25248, g865, g30269, g873, g30277, g876,
         g30285, g879, g30643, g918, g30648, g921, g30654, g30676, g882,
         g30681, g885, g30687, g888, g30649, g927, g30655, g930, g30662, g933,
         g30286, g891, g30293, g894, g30298, g897, g30259, g936, g30264, g939,
         g30270, g942, g30247, g900, g30249, g903, g30251, g906, g30265,
         g30271, g948, g30278, g951, g30638, g909, g30642, g912, g30647, g915,
         g30670, g954, g30677, g957, g30682, g960, g25042, g780, g25935, g776,
         g26530, g771, g27123, g767, g27603, g762, g28146, g758, g28635, g753,
         g29110, g29354, g29580, g740, g868, g869, n4363, n4364, g1088, n4381,
         g996, n4387, g27257, g1041, g27262, g1030, g27270, g1033, g27263,
         g1056, g27271, g1045, g27282, g1048, g27272, g27283, g1060, g27297,
         g1063, g27284, g1085, g27298, g1075, g27313, g1078, g28738, g1095,
         g28746, g1098, g28758, g1101, g29198, g1104, g29204, g1107, g29209,
         g1110, g28747, g1114, g28759, g1115, g28767, g1113, g26806, g1116,
         g26809, g26813, g1122, g26810, g1125, g26814, g1128, g26818, g1131,
         g27761, g1135, g27763, g1136, g27765, g1134, g29609, g999, g29612,
         g1000, g29616, g1001, g30701, g1002, g30703, g1003, g30705, g1004,
         g30470, g1005, g30485, g1006, g30500, g29170, g1009, g29173, g1010,
         g29179, g1008, g26661, g1090, g26665, g1091, g26669, g1089, g1137,
         n8027, DFF_649_n1, g1139, n8026, DFF_651_n1, g1141, n8025, DFF_653_n1,
         g967, n8024, DFF_655_n1, g969, DFF_657_n1, g971, n8021, DFF_659_n1,
         g973, n8020, DFF_661_n1, g975, n8019, DFF_663_n1, g977, n8018, n4486,
         n4283, g986, n4432, g992, n4277, n8017, g1029, g1036, g1037, g1038,
         g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067,
         g1068, g1069, g1070, g1074, g1081, g1083, g1084, g1011, g1024, n4371,
         n4316, g1236, n4300, g1240, g18707, g1243, n4353, g18763, g1196,
         n4304, g1199, g1209, g1210, g1142, g1255, g1145, g1256, g1257, g1148,
         g1258, g1259, g1152, g1260, g1251, g1155, g1252, g1253, g1158, g1254,
         g1176, n4460, n4459, g1172, n4465, g23081, g1173, g23111, g23126,
         g1175, g23392, g23406, g24179, g24181, g1164, g24213, g1165, g24223,
         g1166, g23110, g1167, g23014, g1171, g23039, g1151, g24212, g24222,
         g24235, g1214, g1221, g13155, g1229, n4549, n4361, g13124, g1235,
         g1186, n4548, g13171, g1244, g1245, g27273, g1262, g27285, g1263,
         g27299, g1261, g27286, g1265, g27300, g1266, g27314, g1264, g27301,
         g1268, g27315, g1269, g27328, g27316, g1271, g27329, g1272, g27339,
         g1270, g24501, g1273, g24510, g1276, g24521, g1279, g24511, g1282,
         g24522, g1285, g24532, g1288, g28351, g1300, g28355, g1303, g28360,
         g1306, g28346, g1291, g28350, g1294, g28354, g1297, g26547, g26557,
         g1180, g26569, g1183, g1192, n4454, g22615, n8009, DFF_783_n1,
         DFF_792_n1, g1211, n8008, n8007, DFF_795_n1, n8006, DFF_796_n1, n8005,
         n8004, n8003, g1222, g1223, g24072, g1224, n4489, n4358, g1315, n4294,
         g16671, g1316, g20333, g1345, n4428, g20717, g1326, n4402, g21969,
         g1319, n4476, g23329, g1339, n4421, g24430, g1332, n4412, g25189,
         g1346, n4401, g26666, g1358, n4411, g26781, g1352, n4469, g27678,
         g1365, n4475, g27718, g1372, n4395, g28321, g1378, n4417, g20882,
         g20896, g1386, g20910, g1384, g20897, g1388, g20911, g1389, g20925,
         g1387, g20912, g1391, g20926, g1392, g20949, g1390, g20927, g1394,
         g20950, g1395, g20972, g1393, g20951, g1397, g20973, g1398, g20993,
         g1396, g20974, g1400, g20994, g21015, g1399, g20995, g1403, g21016,
         g1404, g21033, g1402, g21017, g1406, g21034, g1407, g21052, g1405,
         g21035, g1409, g21053, g1410, g21070, g1408, g20883, g1412, g20898,
         g1413, g20913, g1411, g20952, g1415, g20975, g1416, g20996, g20976,
         g1418, g20997, g1419, g21018, g1417, g25263, g1421, g25267, g1422,
         g25270, g1420, g1424, g22247, g1425, g22263, g1423, n4317, n4515,
         g1547, n4368, g22149, g1512, g22166, g1513, g22178, g1511, g22167,
         g22179, g1516, g22191, g1514, g22035, g1524, g22043, g1525, g22057,
         g1523, g22044, g1527, g22058, g1528, g22073, g1526, g22059, g1530,
         g22074, g1531, g22090, g1529, g22075, g1533, g22091, g1534, g22112,
         g1532, g22092, g1536, g22113, g22130, g1535, g22114, g1539, g22131,
         g1540, g22150, g1538, g22132, g1542, g22151, g1543, g22168, g1541,
         g22152, g1545, g22169, g1546, g22180, g1544, g25217, g1551, g25224,
         g1552, g25233, g1550, g25225, g1554, g25234, g1555, g25242, g25235,
         g1557, g25243, g1558, g25249, g1556, g25244, g1560, g25250, g1561,
         g25255, g1559, g30279, g1567, g30287, g1570, g30294, g1573, g30651,
         g1612, g30657, g1615, g30663, g1618, g30683, g1576, g30688, g1579,
         g30692, g1582, g30658, g30664, g1624, g30671, g1627, g30295, g1585,
         g30299, g1588, g30302, g1591, g30266, g1630, g30272, g1633, g30280,
         g1636, g30250, g1594, g30252, g1597, g30255, g1600, g30273, g1639,
         g30281, g1642, g30288, g1645, g30644, g1603, g30650, g30656, g1609,
         g30678, g1648, g30684, g1651, g30689, g1654, g25056, g1466, g1462,
         g26531, g1457, g1453, g27612, g1448, g28147, g1444, g28636, g1439,
         g29111, g1435, g29355, g29581, g1426, g1562, g1563, n4518, g1690,
         n4386, g27264, g1735, g27274, g1724, g27287, g1727, g27275, g1750,
         g27288, g1739, g27302, g1742, g27289, g1765, g27303, g1754, g27317,
         g1757, g27304, g1779, g27318, g27330, g1772, g28749, g1789, g28760,
         g1792, g28771, g1795, g29205, g1798, g29212, g1801, g29218, g1804,
         g28761, g1808, g28772, g1809, g28778, g1807, g26811, g1810, g26815,
         g1813, g26820, g1816, g26816, g1819, g26821, g1822, g26824, g27764,
         g1829, g27766, g1830, g27768, g1828, g29613, g1693, g29617, g1694,
         g29620, g1695, g30704, g1696, g30706, g1697, g30708, g1698, g30487,
         g1699, g30503, g1700, g30338, g1701, g29178, g1703, g29181, g1704,
         g29184, g1702, g26667, g26670, g1785, g26675, g1783, g1831, n7988,
         DFF_999_n1, g1833, n7987, DFF_1001_n1, g1835, n7986, DFF_1003_n1,
         g1661, n7985, DFF_1005_n1, g1663, n7984, DFF_1007_n1, g1665, n7983,
         DFF_1009_n1, g1667, DFF_1011_n1, g1669, n7980, DFF_1013_n1, g1671,
         n7979, n4484, n4284, g1680, n4488, g1686, n4276, n7978, g1723, g1730,
         g1731, g1732, g1733, g1734, g1738, g1745, g1747, g1748, g1749, g1753,
         g1760, g1761, g1762, g1763, g1764, g1768, g1775, g1776, g1777, g1778,
         g1705, g1718, n4296, n4315, g1930, n4366, g1934, g18743, g1937, n4311,
         g18794, g1890, n4297, g1893, g1903, g1904, g1836, g1944, g1949, g1950,
         g1951, g1842, g1953, g1846, g1954, g1945, g1849, g1946, g1947, g1852,
         g1948, g1870, n4458, n4457, g1866, n4464, g23097, g1867, g23124,
         g1868, g23137, g1869, g23400, g23413, g24182, g24208, g1858, g24219,
         g1859, g24231, g1860, g23123, g1861, g23030, g1865, g23058, g1845,
         g24218, g24230, g24243, g1908, g1915, g1922, g13164, g1923,
         DFF_1099_n1, n7971, DFF_1100_n1, g13135, g1929, g1880, n4545, g13182,
         g1938, g1939, g27290, g1956, g27305, g1957, g27319, g1955, g27306,
         g1959, g27320, g1960, g27331, g1958, g27321, g1962, g27332, g1963,
         g27340, g1961, g27333, g27341, g1966, g27346, g1964, g24513, g1967,
         g24524, g1970, g24534, g1973, g24525, g1976, g24535, g1979, g24545,
         g1982, g28357, g1994, g28362, g1997, g28366, g2000, g28352, g1985,
         g28356, g1988, g28361, g1991, g26559, g26573, g1874, g26592, g1877,
         g1886, n4493, g22651, n7968, DFF_1133_n1, DFF_1142_n1, g1905, n7967,
         n7966, DFF_1145_n1, n7965, DFF_1146_n1, n7964, n7963, n7962, g1916,
         g1917, g24083, n7960, n4357, g2009, n4293, g16692, g2010, g20353,
         g2039, n4427, g20752, g2020, n4400, g21972, g2013, n4474, g23339,
         g2033, n4420, g24434, g2026, n4410, g25194, g2040, n4399, g26671,
         g2052, n4409, g26789, g2046, n4468, g27682, g2059, n4473, g27722,
         g28325, g2072, n4416, g20899, g2079, g20915, g2080, g20934, g2078,
         g20916, g2082, g20935, g2083, g20953, g2081, g20936, g2085, g20954,
         g2086, g20977, g2084, g20955, g2088, g20978, g2089, g20999, g2087,
         g20979, g2091, g21000, g21019, g2090, g21001, g2094, g21020, g2095,
         g21039, g2093, g21021, g2097, g21040, g2098, g21054, g2096, g21041,
         g2100, g21055, g2101, g21071, g2099, g21056, g2103, g21072, g2104,
         g21080, g2102, g20900, g2106, g20917, g20937, g2105, g20980, g2109,
         g21002, g2110, g21022, g2108, g21003, g2112, g21023, g2113, g21042,
         g2111, g25268, g2115, g25271, g2116, g25279, g2114, g2118, g22267,
         g2119, g22280, g2117, n4324, g2241, n4367, g22170, g2206, g22182,
         g2207, g22192, g2205, g22183, g2209, g22193, g2210, g22200, g2208,
         g22045, g2218, g22060, g2219, g22076, g2217, g22061, g2221, g22077,
         g2222, g22097, g2220, g22078, g2224, g22098, g22115, g2223, g22099,
         g2227, g22116, g2228, g22138, g2226, g22117, g2230, g22139, g2231,
         g22153, g2229, g22140, g2233, g22154, g2234, g22171, g2232, g22155,
         g2236, g22172, g2237, g22184, g2235, g22173, g2239, g22185, g22194,
         g2238, g25227, g2245, g25236, g2246, g25245, g2244, g25237, g2248,
         g25246, g2249, g25251, g2247, g25247, g2251, g25252, g2252, g25256,
         g2250, g25253, g2254, g25257, g2255, g25259, g2253, g30289, g2261,
         g30296, g30300, g2267, g30660, g2306, g30666, g2309, g30672, g2312,
         g30690, g2270, g30693, g2273, g30695, g2276, g30667, g2315, g30673,
         g2318, g30679, g2321, g30301, g2279, g30303, g2282, g30304, g2285,
         g30274, g2324, g30282, g30290, g2330, g30253, g2288, g30256, g2291,
         g30260, g2294, g30283, g2333, g30291, g2336, g30297, g2339, g30652,
         g2297, g30659, g2300, g30665, g2303, g30686, g2342, g30691, g2345,
         g30694, g2348, g25067, g2160, g26532, g2151, g2147, g27621, g2142,
         g28148, g2138, g28637, g2133, g29112, g2129, g29357, g29582, g2120,
         g2256, g2257, n4516, g27276, g2429, g27291, g2418, g27307, g2421,
         g27292, g2444, g27308, g2433, g27322, g2436, g27309, g2459, g27323,
         g2448, g27334, g2451, g27324, g2473, g27335, g2463, g27342, g2466,
         g28763, g2483, g28773, g2486, g28782, g29213, g2492, g29221, g2495,
         g29226, g2498, g28774, g2502, g28783, g2503, g28788, g2501, g26817,
         g2504, g26822, g2507, g26825, g2510, g26823, g2513, g26826, g2516,
         g26827, g2519, g27767, g2523, g27769, g2524, g27771, g29618, g2387,
         g29621, g2388, g29623, g2389, g30707, g2390, g30709, g2391, g30566,
         g2392, g30505, g2393, g30341, g2394, g30356, g2395, g29182, g2397,
         g29185, g2398, g29187, g2396, g26672, g2478, g26676, g2479, g26025,
         g2525, n7946, DFF_1349_n1, g2527, n7945, DFF_1351_n1, g2529, n7944,
         DFF_1353_n1, g2355, n7943, DFF_1355_n1, g2357, n7942, DFF_1357_n1,
         g2359, n7941, DFF_1359_n1, g2361, n7940, DFF_1361_n1, n7938,
         DFF_1363_n1, g2365, n7937, n4483, n4285, g2374, n4487, g30055, g2380,
         n4275, n7936, DFF_1378_n1, g2417, g2424, g2425, g2426, g2427, g2428,
         g2432, g2439, g2441, g2442, g2443, g2447, g2454, g2455, g2456, g2457,
         g2458, g2462, g2469, g2470, g2471, g2472, g2412, n4314, n4370, g2624,
         n4299, g2628, g18780, g2631, n4352, g18820, g2584, n4303, g2587,
         g2597, g2598, g2530, g2638, g2643, g2533, g2645, g2536, g2646, g2647,
         g2540, g2648, g2639, g2543, g2640, g2641, g2546, g2642, g2564, n4456,
         n4455, g2560, n4463, g23114, g2561, g23133, g2562, g21970, g23407,
         g23418, g24209, g24214, g2552, g24226, g2553, g24238, g2554, g23132,
         g2555, g23047, g2559, g23076, g2539, g24225, g24237, g24250, g2602,
         g2609, g13175, g2617, n7930, g30072, n7929, g13143, g2623, g2574,
         n4543, g13194, g2632, g2633, g27310, g2650, g27325, g2651, g27336,
         g2649, g27326, g2653, g27337, g2654, g27343, g2652, g27338, g2656,
         g27344, g27347, g2655, g27345, g2659, g27348, g2660, g27354, g2658,
         g24527, g2661, g24537, g2664, g24547, g2667, g24538, g2670, g24548,
         g2673, g24557, g2676, g28364, g2688, g28368, g2691, g28371, g2694,
         g28358, g2679, g28363, g28367, g2685, g26575, g2565, g26596, g2568,
         g26616, g2571, g2580, g22687, n7926, g30061, g2599, n7925, n7924,
         DFF_1495_n1, n7923, DFF_1496_n1, n7922, n7921, n7920, g2611, g24092,
         g2612, n4490, n7918, n4356, g2703, n4292, g16718, g2704, g20375,
         g2733, g20789, g2714, n4398, g21974, g2707, n4472, g23348, g2727,
         n4419, g24438, g2720, n4408, g25197, g2734, n4397, g26677, g2746,
         n4407, g26795, g27243, g2753, n4471, g2760, n4393, g28328, g2766,
         n4415, g20918, g2773, g20939, g2774, g20962, g2772, g20940, g2776,
         g20963, g2777, g20981, g2775, g20964, g2779, g20982, g2780, g21004,
         g2778, g20983, g2782, g21005, g2783, g21025, g21006, g2785, g21026,
         g2786, g21043, g2784, g21027, g2788, g21044, g2789, g21060, g2787,
         g21045, g2791, g21061, g2792, g21073, g2790, g21062, g2794, g21074,
         g2795, g21081, g2793, g21075, g2797, g21082, g2798, g21094, g20919,
         g2800, g20941, g2801, g20965, g2799, g21007, g2803, g21028, g2804,
         g21046, g2802, g21029, g2806, g21047, g2807, g21063, g2805, g25272,
         g2809, g25280, g2810, g25288, g2808, g2812, g22284, g2813, g22299,
         g20877, n7913, DFF_1561_n1, g20884, n7912, DFF_1562_n1,
         n4263_Tj_Payload, n4269, g3043, n4268, g3044, n4267, g3045, n4266,
         g3046, n4265, g3047, n4272, g3048, n4271, g3049, n4270, g3050, n4259,
         g3051, n4236, g3052, n4239, g3053, n4237, n4234, g3056, n4233, g3057,
         n4238, g3058, n4235, g3059, n4240, g3060, n4232, g3061, n4245, g3062,
         n4248, g3063, n4246, g3064, n4243, g3065, n4242, g3066, n4247, g3067,
         n4244, g3068, n4249, g3069, n4241, n4254, g3071, n4257, g3072, n4255,
         g3073, n4252, g3074, n4251, g3075, n4256, g3076, n4253, g3077, n4258,
         g3078, n4250, g2997, g25265, g2993, g26048, n7909, g23330, g3006,
         g24445, g3002, g25191, g3013, g26031, g26786, g3024, n4262, g3018,
         n4481, g23359, g3028, n4350, g24446, g3036, n4480, g25202, g3032,
         n7907, DFF_1612_n1, g2987, n4365, g16824, g16844, g16853, g16860,
         g16803, DFF_1618_n1, g16835, g16851, g16857, g16866, g3083, n4261,
         N995, n4577, g16845, g16854, g16861, g16880, DFF_1628_n1, g18755,
         g18804, g18837, g18868, g18907, g2990, N690, n4578, n4260, n4309,
         n4308, n4307, n4306, n4524, n4525, n4511, n4509, n4499, n4520, n3683,
         n3887, n3686, n3890, n3692, n3896, n4513, n3897, n3424, n3427, n3433,
         n4529, n4530, n4522, n4523, n4521, n3171, n3159, n3163, n3893, n3690,
         n3689, n3431, n3430, n3168, n3160, n3164, n3172, n4527, n4528, n4526,
         n3167, n3894, n3888, n3891, n2302, n2289, n2303, n2275, n4066, n4065,
         n4606, n4618, n4640, n2792, n2632, n3936, n3252, n3254, n4102, n3038,
         n3070, n3102, n3130, n3036, n3068, n3065, n3128, n2800, n2798, n2616,
         n2594, n3940, n3705, n3933, n3939, n3016, n3000, n3008, n3023, n3700,
         n4058, n4123, n4101, n4182, n4073, n3749, n3751, n3758, n3788, n4057,
         n4122, n4263, Tj_OUT1, Tj_OUT2, Tj_OUT3, Tj_OUT4, Tj_OUT1234, Tj_OUT5,
         Tj_OUT6, Tj_OUT7, Tj_OUT8, Tj_OUT5678, Tj_Trigger, n6, n7, n15, n46,
         n47, n50, n51, n53, n54, n92, n158, n276, n295, n296, n299, n307,
         n348, n477, n478, n492, n506, n521, n522, n532, n540, n541, n548,
         n549, n550, n552, n589, n614, n681, n845, n846, n854, n890, n984,
         n1149, n1152, n1159, n1194, n1290, n1421, n1456, n1457, n1458, n1464,
         n1499, n1524, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8395, n8397,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8411,
         n8412, n8413, n8415, n8416, n8418, n8419, n8420, n8421, n8422, n8423,
         n8428, n8429, n8431, n8433, n8434, n8436, n8437, n8439, n8440, n8441,
         n8443, n8445, n8447, n8449, n8451, n8452, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8471, n8473, n8475, n8477, n8478, n8480, n8481, n8482,
         n8487, n8488, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8515, n8517, n8521, n8523, n8526, n8527, n8528, n8529, n8530, n8531,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8544, n8545, n8546,
         n8547, n8548, n8554, n8558, n8559, n8560, n8561, n8562, n8563, n8566,
         n8568, n8570, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8586, n8588, n8590, n8595, n8596, n8597, n8598, n8601, n8602,
         n8604, n8609, n8610, n8611, n8612, n8613, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8630, n8631, n8632, n8633, n8637, n8640, n8642, n8643, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8675, n8676, n8678, n8679,
         n8681, n8683, n8685, n8686, n8687, n8688, n8689, n8691, n8692, n8693,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8713, n8715, n8719,
         n8721, n8723, n8726, n8728, n8730, n8732, n8733, n8734, n8736, n8737,
         n8739, n8740, n8742, n8743, n8745, n8746, n8747, n8749, n8750, n8752,
         n8753, n8755, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8774, n8776, n8777, n8779, n8785, n8787, n8789, n8790, n8792,
         n8793, n8794, n8803, n8805, n8815, n8816, n8817, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8837, n8839, n8841, n8843,
         n8850, n8853, n8856, n8859, n8862, n8865, n8867, n8870, n8872, n8875,
         n8878, n8881, n8884, n8887, n8890, n8893, n8896, n8898, n8901, n8903,
         n8906, n8908, n8913, n8915, n8919, n8924, n8926, n8929, n8931, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8943, n8946, n8950, n8951,
         n8954, n8956, n8957, n8958, n8962, n8963, n8964, n8965, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8998, n8999, n9001, n9002,
         n9004, n9005, n9007, n9008, n9010, n9011, n9013, n9015, n9016, n9018,
         n9019, n9021, n9022, n9024, n9025, n9027, n9028, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9040, n9042, n9044, n9046, n9048, n9050,
         n9052, n9054, n9056, n9058, n9061, n9063, n9065, n9067, n9070, n9072,
         n9074, n9076, n9078, n9080, n9082, n9084, n9087, n9089, n9091, n9093,
         n9095, n9097, n9099, n9101, n9103, n9105, n9106, n9108, n9110, n9112,
         n9152, n9153, n9154, n9155, n9156, n9158, n9160, n9163, n9165, n9167,
         n9169, n9171, n9174, n9176, n9178, n9180, n9182, n9183, n9200, n9202,
         n9204, n9206, n9208, n9210, n9212, n9214, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9236, n9238, n9240, n9241, n9242, n9244, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9270, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         U3772_n1, U3776_n1, U3777_n1, U3778_n1, U3779_n1, U3780_n1, U3781_n1,
         U3782_n1, U3783_n1, U3784_n1, U3785_n1, U3786_n1, U3787_n1, U3901_n1,
         U3902_n1, U4467_n1, U4904_n1, U4930_n1, U5128_n1, U5141_n1, U5749_n1,
         U5750_n1, U5751_n1, U5752_n1, U5753_n1, U5754_n1, U5755_n1, U5756_n1,
         U5757_n1, U5758_n1, U5759_n1, U5760_n1, U5761_n1, U5762_n1, U5763_n1,
         U5764_n1, U5882_n1, U5939_n1, U5940_n1, U5941_n1, U5942_n1, U6140_n1,
         U6460_n1, U6470_n1, U6562_n1, U6563_n1, U6718_n1, U7116_n1, U7118_n1,
         U7293_n1;
  assign g8251 = test_so3;
  assign g7519 = test_so4;
  assign g4450 = test_so5;
  assign g7909 = test_so23;
  assign g5612 = test_so57;
  assign g5695 = test_so63;
  assign g7084 = test_so73;
  assign g8270 = test_so99;
  assign g8258 = test_so100;

  SDFFX1 DFF_0_Q_reg ( .D(g51), .SI(test_si1), .SE(n9295), .CLK(n9482), .Q(
        n8104), .QN(n16829) );
  SDFFX1 DFF_1_Q_reg ( .D(g16802), .SI(n8104), .SE(n9295), .CLK(n9482), .Q(
        n8103), .QN(DFF_1_n1) );
  SDFFX1 DFF_2_Q_reg ( .D(g16823), .SI(n8103), .SE(n9295), .CLK(n9482), .Q(
        n8102), .QN(DFF_2_n1) );
  SDFFX1 DFF_3_Q_reg ( .D(n4264), .SI(n8102), .SE(n9295), .CLK(n9482), .Q(
        g2950), .QN(n4423) );
  SDFFX1 DFF_4_Q_reg ( .D(n4274), .SI(g2950), .SE(n9296), .CLK(n9483), .Q(
        g2883), .QN(n4330) );
  SDFFX1 DFF_5_Q_reg ( .D(g22026), .SI(g2883), .SE(n9296), .CLK(n9483), .Q(
        g2888) );
  SDFFX1 DFF_6_Q_reg ( .D(n6), .SI(g2888), .SE(n9296), .CLK(n9483), .Q(g2896), 
        .QN(n4431) );
  SDFFX1 DFF_7_Q_reg ( .D(g24473), .SI(g2896), .SE(n9296), .CLK(n9483), .Q(
        g2892) );
  SDFFX1 DFF_8_Q_reg ( .D(n7), .SI(g2892), .SE(n9296), .CLK(n9483), .Q(g2903), 
        .QN(n4305) );
  SDFFX1 DFF_9_Q_reg ( .D(g26037), .SI(g2903), .SE(n9296), .CLK(n9483), .Q(
        g2900), .QN(n4291) );
  SDFFX1 DFF_10_Q_reg ( .D(g26798), .SI(g2900), .SE(n9296), .CLK(n9483), .Q(
        g2908), .QN(n4355) );
  SDFFX1 DFF_11_Q_reg ( .D(n4273), .SI(g2908), .SE(n9296), .CLK(n9483), .Q(
        g2912), .QN(n4482) );
  SDFFX1 DFF_12_Q_reg ( .D(g23357), .SI(g2912), .SE(n9296), .CLK(n9483), .Q(
        g2917), .QN(n4479) );
  SDFFX1 DFF_13_Q_reg ( .D(g24476), .SI(g2917), .SE(n9296), .CLK(n9483), .Q(
        g2924), .QN(n4349) );
  SDFFX1 DFF_14_Q_reg ( .D(g25199), .SI(g2924), .SE(n9296), .CLK(n9483), .Q(
        g2920), .QN(n8985) );
  SDFFX1 DFF_15_Q_reg ( .D(n4280), .SI(g2920), .SE(n9296), .CLK(n9483), .Q(
        test_so1), .QN(DFF_15_n1) );
  SDFFX1 DFF_16_Q_reg ( .D(n4281), .SI(test_si2), .SE(n9293), .CLK(n9480), .Q(
        n8099), .QN(DFF_16_n1) );
  SDFFX1 DFF_17_Q_reg ( .D(g51), .SI(n8099), .SE(n9293), .CLK(n9480), .Q(g8021) );
  SDFFX1 DFF_18_Q_reg ( .D(g8021), .SI(g8021), .SE(n9293), .CLK(n9480), .Q(
        n8098), .QN(DFF_18_n1) );
  SDFFX1 DFF_19_Q_reg ( .D(n4279), .SI(n8098), .SE(n9293), .CLK(n9480), .Q(
        g2879), .QN(n4351) );
  SDFFX1 DFF_20_Q_reg ( .D(g3212), .SI(g2879), .SE(n9293), .CLK(n9480), .Q(
        g2934) );
  SDFFX1 DFF_21_Q_reg ( .D(g3228), .SI(g2934), .SE(n9293), .CLK(n9480), .Q(
        g2935), .QN(n9234) );
  SDFFX1 DFF_22_Q_reg ( .D(g3227), .SI(g2935), .SE(n9294), .CLK(n9481), .Q(
        g2938) );
  SDFFX1 DFF_23_Q_reg ( .D(g3226), .SI(g2938), .SE(n9294), .CLK(n9481), .Q(
        g2941), .QN(n9232) );
  SDFFX1 DFF_24_Q_reg ( .D(g3225), .SI(g2941), .SE(n9294), .CLK(n9481), .Q(
        g2944), .QN(n9238) );
  SDFFX1 DFF_25_Q_reg ( .D(g3224), .SI(g2944), .SE(n9294), .CLK(n9481), .Q(
        g2947), .QN(n9236) );
  SDFFX1 DFF_26_Q_reg ( .D(g3223), .SI(g2947), .SE(n9294), .CLK(n9481), .Q(
        g2953) );
  SDFFX1 DFF_27_Q_reg ( .D(g3222), .SI(g2953), .SE(n9294), .CLK(n9481), .Q(
        g2956) );
  SDFFX1 DFF_28_Q_reg ( .D(g3221), .SI(g2956), .SE(n9294), .CLK(n9481), .Q(
        g2959), .QN(n9233) );
  SDFFX1 DFF_29_Q_reg ( .D(g3232), .SI(g2959), .SE(n9294), .CLK(n9481), .Q(
        g2962), .QN(n9252) );
  SDFFX1 DFF_30_Q_reg ( .D(g3220), .SI(g2962), .SE(n9294), .CLK(n9481), .Q(
        g2963), .QN(n9242) );
  SDFFX1 DFF_31_Q_reg ( .D(g3219), .SI(g2963), .SE(n9294), .CLK(n9481), .Q(
        test_so2) );
  SDFFX1 DFF_32_Q_reg ( .D(g3218), .SI(test_si3), .SE(n9293), .CLK(n9480), .Q(
        g2969) );
  SDFFX1 DFF_33_Q_reg ( .D(g3217), .SI(g2969), .SE(n9293), .CLK(n9480), .Q(
        g2972) );
  SDFFX1 DFF_34_Q_reg ( .D(g3216), .SI(g2972), .SE(n9293), .CLK(n9480), .Q(
        g2975), .QN(n9244) );
  SDFFX1 DFF_35_Q_reg ( .D(g3215), .SI(g2975), .SE(n9293), .CLK(n9480), .Q(
        g2978), .QN(n9240) );
  SDFFX1 DFF_36_Q_reg ( .D(g3214), .SI(g2978), .SE(n9293), .CLK(n9480), .Q(
        g2981) );
  SDFFX1 DFF_37_Q_reg ( .D(g3213), .SI(g2981), .SE(n9293), .CLK(n9480), .Q(
        g2874), .QN(n9241) );
  SDFFX1 DFF_38_Q_reg ( .D(g18754), .SI(g2874), .SE(n9294), .CLK(n9481), .Q(
        g1506), .QN(n4288) );
  SDFFX1 DFF_39_Q_reg ( .D(g18781), .SI(g1506), .SE(n9294), .CLK(n9481), .Q(
        g1501), .QN(n4565) );
  SDFFX1 DFF_40_Q_reg ( .D(g18803), .SI(g1501), .SE(n9295), .CLK(n9482), .Q(
        g1496), .QN(n4557) );
  SDFFX1 DFF_41_Q_reg ( .D(g18821), .SI(g1496), .SE(n9295), .CLK(n9482), .Q(
        g1491), .QN(n4326) );
  SDFFX1 DFF_42_Q_reg ( .D(g18835), .SI(g1491), .SE(n9295), .CLK(n9482), .Q(
        g1486), .QN(n4390) );
  SDFFX1 DFF_43_Q_reg ( .D(g18852), .SI(g1486), .SE(n9295), .CLK(n9482), .Q(
        g1481), .QN(n4320) );
  SDFFX1 DFF_44_Q_reg ( .D(g18866), .SI(g1481), .SE(n9295), .CLK(n9482), .Q(
        g1476), .QN(n4374) );
  SDFFX1 DFF_45_Q_reg ( .D(g18883), .SI(g1476), .SE(n9295), .CLK(n9482), .Q(
        g1471), .QN(n4378) );
  SDFFX1 DFF_46_Q_reg ( .D(g21880), .SI(g1471), .SE(n9300), .CLK(n9487), .Q(
        g2877) );
  SDFFX1 DFF_47_Q_reg ( .D(g19154), .SI(g2877), .SE(n9301), .CLK(n9488), .Q(
        test_so3) );
  SDFFX1 DFF_48_Q_reg ( .D(test_so3), .SI(test_si4), .SE(n9301), .CLK(n9488), 
        .Q(g813), .QN(n4289) );
  SDFFX1 DFF_49_Q_reg ( .D(g19163), .SI(g813), .SE(n9301), .CLK(n9488), .Q(
        g4090) );
  SDFFX1 DFF_50_Q_reg ( .D(g4090), .SI(g4090), .SE(n9301), .CLK(n9488), .Q(
        g809), .QN(n4567) );
  SDFFX1 DFF_51_Q_reg ( .D(g19173), .SI(g809), .SE(n9301), .CLK(n9488), .Q(
        g4323) );
  SDFFX1 DFF_52_Q_reg ( .D(g4323), .SI(g4323), .SE(n9301), .CLK(n9488), .Q(
        g805), .QN(n4559) );
  SDFFX1 DFF_53_Q_reg ( .D(g19184), .SI(g805), .SE(n9301), .CLK(n9488), .Q(
        g4590) );
  SDFFX1 DFF_54_Q_reg ( .D(g4590), .SI(g4590), .SE(n9301), .CLK(n9488), .Q(
        g801), .QN(n4327) );
  SDFFX1 DFF_55_Q_reg ( .D(g20310), .SI(g801), .SE(n9301), .CLK(n9488), .Q(
        g6225) );
  SDFFX1 DFF_56_Q_reg ( .D(g6225), .SI(g6225), .SE(n9301), .CLK(n9488), .Q(
        g797), .QN(n4391) );
  SDFFX1 DFF_57_Q_reg ( .D(g20343), .SI(g797), .SE(n9301), .CLK(n9488), .Q(
        g6442) );
  SDFFX1 DFF_58_Q_reg ( .D(g6442), .SI(g6442), .SE(n9302), .CLK(n9489), .Q(
        g793), .QN(n4321) );
  SDFFX1 DFF_59_Q_reg ( .D(g20376), .SI(g793), .SE(n9302), .CLK(n9489), .Q(
        g6895) );
  SDFFX1 DFF_60_Q_reg ( .D(g6895), .SI(g6895), .SE(n9302), .CLK(n9489), .Q(
        g789), .QN(n4375) );
  SDFFX1 DFF_61_Q_reg ( .D(g20417), .SI(g789), .SE(n9302), .CLK(n9489), .Q(
        g7334) );
  SDFFX1 DFF_62_Q_reg ( .D(g7334), .SI(g7334), .SE(n9302), .CLK(n9489), .Q(
        g785), .QN(n4379) );
  SDFFX1 DFF_63_Q_reg ( .D(g21878), .SI(g785), .SE(n9302), .CLK(n9489), .Q(
        test_so4) );
  SDFFX1 DFF_64_Q_reg ( .D(test_so4), .SI(test_si5), .SE(n9303), .CLK(n9490), 
        .Q(g2873) );
  SDFFX1 DFF_65_Q_reg ( .D(g19153), .SI(g2873), .SE(n9303), .CLK(n9490), .Q(
        g8249) );
  SDFFX1 DFF_66_Q_reg ( .D(g8249), .SI(g8249), .SE(n9303), .CLK(n9490), .Q(
        g125), .QN(n4290) );
  SDFFX1 DFF_67_Q_reg ( .D(g19162), .SI(g125), .SE(n9303), .CLK(n9490), .Q(
        g4088) );
  SDFFX1 DFF_68_Q_reg ( .D(g4088), .SI(g4088), .SE(n9303), .CLK(n9490), .Q(
        g121), .QN(n4569) );
  SDFFX1 DFF_69_Q_reg ( .D(g19172), .SI(g121), .SE(n9303), .CLK(n9490), .Q(
        g4321) );
  SDFFX1 DFF_70_Q_reg ( .D(g4321), .SI(g4321), .SE(n9303), .CLK(n9490), .Q(
        g117), .QN(n4561) );
  SDFFX1 DFF_71_Q_reg ( .D(g19144), .SI(g117), .SE(n9303), .CLK(n9490), .Q(
        g8023) );
  SDFFX1 DFF_72_Q_reg ( .D(g8023), .SI(g8023), .SE(n9303), .CLK(n9490), .Q(
        g113), .QN(n4328) );
  SDFFX1 DFF_73_Q_reg ( .D(g19149), .SI(g113), .SE(n9303), .CLK(n9490), .Q(
        g8175) );
  SDFFX1 DFF_74_Q_reg ( .D(g8175), .SI(g8175), .SE(n9304), .CLK(n9491), .Q(
        g109), .QN(n4392) );
  SDFFX1 DFF_75_Q_reg ( .D(g19157), .SI(g109), .SE(n9304), .CLK(n9491), .Q(
        g3993) );
  SDFFX1 DFF_76_Q_reg ( .D(g3993), .SI(g3993), .SE(n9304), .CLK(n9491), .Q(
        g105), .QN(n4322) );
  SDFFX1 DFF_77_Q_reg ( .D(g19167), .SI(g105), .SE(n9304), .CLK(n9491), .Q(
        g4200) );
  SDFFX1 DFF_78_Q_reg ( .D(g4200), .SI(g4200), .SE(n9304), .CLK(n9491), .Q(
        g101), .QN(n4376) );
  SDFFX1 DFF_79_Q_reg ( .D(g19178), .SI(g101), .SE(n9304), .CLK(n9491), .Q(
        test_so5) );
  SDFFX1 DFF_80_Q_reg ( .D(test_so5), .SI(test_si6), .SE(n9304), .CLK(n9491), 
        .Q(g97), .QN(n4380) );
  SDFFX1 DFF_81_Q_reg ( .D(g20874), .SI(g97), .SE(n9304), .CLK(n9491), .Q(
        g8096) );
  SDFFX1 DFF_82_Q_reg ( .D(g8096), .SI(g8096), .SE(n9304), .CLK(n9491), .Q(
        g2857) );
  SDFFX1 DFF_83_Q_reg ( .D(g18885), .SI(g2857), .SE(n9304), .CLK(n9491), .Q(
        g2200), .QN(n4287) );
  SDFFX1 DFF_84_Q_reg ( .D(g18975), .SI(g2200), .SE(n9304), .CLK(n9491), .Q(
        g2195), .QN(n4563) );
  SDFFX1 DFF_85_Q_reg ( .D(g18968), .SI(g2195), .SE(n9304), .CLK(n9491), .Q(
        g2190), .QN(n4555) );
  SDFFX1 DFF_86_Q_reg ( .D(g18942), .SI(g2190), .SE(n9305), .CLK(n9492), .Q(
        g2185), .QN(n4325) );
  SDFFX1 DFF_87_Q_reg ( .D(g18906), .SI(g2185), .SE(n9305), .CLK(n9492), .Q(
        g2180), .QN(n4389) );
  SDFFX1 DFF_88_Q_reg ( .D(g18867), .SI(g2180), .SE(n9305), .CLK(n9492), .Q(
        g2175), .QN(n4319) );
  SDFFX1 DFF_89_Q_reg ( .D(g18836), .SI(g2175), .SE(n9305), .CLK(n9492), .Q(
        g2170), .QN(n4373) );
  SDFFX1 DFF_90_Q_reg ( .D(g18957), .SI(g2170), .SE(n9305), .CLK(n9492), .Q(
        g2165), .QN(n4377) );
  SDFFX1 DFF_91_Q_reg ( .D(g21882), .SI(g2165), .SE(n9321), .CLK(n9508), .Q(
        g2878) );
  SDFFX1 DFF_92_Q_reg ( .D(n4598), .SI(g2878), .SE(n9419), .CLK(n9606), .Q(
        g8106), .QN(n4382) );
  SDFFX1 DFF_93_Q_reg ( .D(g8106), .SI(g8106), .SE(n9419), .CLK(n9606), .Q(
        g8030), .QN(n4383) );
  SDFFX1 DFF_94_Q_reg ( .D(g8030), .SI(g8030), .SE(n9419), .CLK(n9606), .Q(
        g3109), .QN(n4494) );
  SDFFX1 DFF_95_Q_reg ( .D(g18669), .SI(g3109), .SE(n9420), .CLK(n9607), .Q(
        test_so6) );
  SDFFX1 DFF_96_Q_reg ( .D(g18719), .SI(test_si7), .SE(n9419), .CLK(n9606), 
        .Q(g3211) );
  SDFFX1 DFF_97_Q_reg ( .D(g18782), .SI(g3211), .SE(n9419), .CLK(n9606), .Q(
        g3084), .QN(n4445) );
  SDFFX1 DFF_98_Q_reg ( .D(g17222), .SI(g3084), .SE(n9421), .CLK(n9608), .Q(
        g3085), .QN(n4340) );
  SDFFX1 DFF_99_Q_reg ( .D(g17225), .SI(g3085), .SE(n9421), .CLK(n9608), .Q(
        g3086), .QN(n4337) );
  SDFFX1 DFF_100_Q_reg ( .D(g17234), .SI(g3086), .SE(n9421), .CLK(n9608), .Q(
        g3087), .QN(n4344) );
  SDFFX1 DFF_101_Q_reg ( .D(g17224), .SI(g3087), .SE(n9421), .CLK(n9608), .Q(
        g3091), .QN(n4448) );
  SDFFX1 DFF_102_Q_reg ( .D(g17228), .SI(g3091), .SE(n9421), .CLK(n9608), .Q(
        g3092), .QN(n4451) );
  SDFFX1 DFF_103_Q_reg ( .D(g17246), .SI(g3092), .SE(n9422), .CLK(n9609), .Q(
        g3093) );
  SDFFX1 DFF_104_Q_reg ( .D(g17226), .SI(g3093), .SE(n9422), .CLK(n9609), .Q(
        g3094) );
  SDFFX1 DFF_105_Q_reg ( .D(g17235), .SI(g3094), .SE(n9422), .CLK(n9609), .Q(
        g3095), .QN(n4439) );
  SDFFX1 DFF_106_Q_reg ( .D(g17269), .SI(g3095), .SE(n9422), .CLK(n9609), .Q(
        g3096), .QN(n4336) );
  SDFFX1 DFF_107_Q_reg ( .D(g25450), .SI(g3096), .SE(n9422), .CLK(n9609), .Q(
        g3097), .QN(n4433) );
  SDFFX1 DFF_108_Q_reg ( .D(g25451), .SI(g3097), .SE(n9422), .CLK(n9609), .Q(
        g3098), .QN(n4434) );
  SDFFX1 DFF_109_Q_reg ( .D(g25452), .SI(g3098), .SE(n9422), .CLK(n9609), .Q(
        g3099), .QN(n4443) );
  SDFFX1 DFF_110_Q_reg ( .D(g28420), .SI(g3099), .SE(n9422), .CLK(n9609), .Q(
        g3100), .QN(n4342) );
  SDFFX1 DFF_111_Q_reg ( .D(g28421), .SI(g3100), .SE(n9422), .CLK(n9609), .Q(
        test_so7), .QN(n9288) );
  SDFFX1 DFF_112_Q_reg ( .D(g28425), .SI(test_si8), .SE(n9419), .CLK(n9606), 
        .Q(g3102), .QN(n4343) );
  SDFFX1 DFF_113_Q_reg ( .D(g29936), .SI(g3102), .SE(n9420), .CLK(n9607), .Q(
        g3103), .QN(n4447) );
  SDFFX1 DFF_114_Q_reg ( .D(g29939), .SI(g3103), .SE(n9420), .CLK(n9607), .Q(
        g3104), .QN(n4452) );
  SDFFX1 DFF_115_Q_reg ( .D(g29941), .SI(g3104), .SE(n9420), .CLK(n9607), .Q(
        g3105) );
  SDFFX1 DFF_116_Q_reg ( .D(g30796), .SI(g3105), .SE(n9420), .CLK(n9607), .Q(
        g3106), .QN(n4438) );
  SDFFX1 DFF_117_Q_reg ( .D(g30798), .SI(g3106), .SE(n9420), .CLK(n9607), .Q(
        g3107), .QN(n4437) );
  SDFFX1 DFF_118_Q_reg ( .D(g30801), .SI(g3107), .SE(n9420), .CLK(n9607), .Q(
        g3108), .QN(n4334) );
  SDFFX1 DFF_119_Q_reg ( .D(g17229), .SI(g3108), .SE(n9420), .CLK(n9607), .Q(
        g3155) );
  SDFFX1 DFF_120_Q_reg ( .D(g17247), .SI(g3155), .SE(n9420), .CLK(n9607), .Q(
        g3158), .QN(n4436) );
  SDFFX1 DFF_121_Q_reg ( .D(g17302), .SI(g3158), .SE(n9421), .CLK(n9608), .Q(
        g3161) );
  SDFFX1 DFF_122_Q_reg ( .D(g17236), .SI(g3161), .SE(n9421), .CLK(n9608), .Q(
        g3164), .QN(n4339) );
  SDFFX1 DFF_123_Q_reg ( .D(g17270), .SI(g3164), .SE(n9421), .CLK(n9608), .Q(
        g3167), .QN(n4348) );
  SDFFX1 DFF_124_Q_reg ( .D(g17340), .SI(g3167), .SE(n9421), .CLK(n9608), .Q(
        g3170), .QN(n4441) );
  SDFFX1 DFF_125_Q_reg ( .D(g17248), .SI(g3170), .SE(n9421), .CLK(n9608), .Q(
        g3173), .QN(n4338) );
  SDFFX1 DFF_126_Q_reg ( .D(g17303), .SI(g3173), .SE(n9421), .CLK(n9608), .Q(
        g3176), .QN(n4450) );
  SDFFX1 DFF_127_Q_reg ( .D(g17383), .SI(g3176), .SE(n9421), .CLK(n9608), .Q(
        test_so8) );
  SDFFX1 DFF_128_Q_reg ( .D(g17271), .SI(test_si9), .SE(n9420), .CLK(n9607), 
        .Q(g3182), .QN(n4453) );
  SDFFX1 DFF_129_Q_reg ( .D(g17341), .SI(g3182), .SE(n9420), .CLK(n9607), .Q(
        g3185), .QN(n4442) );
  SDFFX1 DFF_130_Q_reg ( .D(g17429), .SI(g3185), .SE(n9420), .CLK(n9607), .Q(
        g3088), .QN(n4341) );
  SDFFX1 DFF_131_Q_reg ( .D(g24734), .SI(g3088), .SE(n9422), .CLK(n9609), .Q(
        n8090) );
  SDFFX1 DFF_132_Q_reg ( .D(g25442), .SI(n8090), .SE(n9423), .CLK(n9610), .Q(
        n8089), .QN(n16824) );
  SDFFX1 DFF_133_Q_reg ( .D(g25435), .SI(n8089), .SE(n9423), .CLK(n9610), .Q(
        g3197) );
  SDFFX1 DFF_134_Q_reg ( .D(g25420), .SI(g3197), .SE(n9423), .CLK(n9610), .Q(
        n8088) );
  SDFFX1 DFF_135_Q_reg ( .D(g26149), .SI(n8088), .SE(n9299), .CLK(n9486), .Q(
        g3201), .QN(n4406) );
  SDFFX1 DFF_136_Q_reg ( .D(g26135), .SI(g3201), .SE(n9299), .CLK(n9486), .Q(
        g3204), .QN(n9254) );
  SDFFX1 DFF_137_Q_reg ( .D(g26104), .SI(g3204), .SE(n9299), .CLK(n9486), .Q(
        g3207), .QN(n4329) );
  SDFFX1 DFF_138_Q_reg ( .D(g27380), .SI(g3207), .SE(n9298), .CLK(n9485), .Q(
        g3188), .QN(n4405) );
  SDFFX1 DFF_139_Q_reg ( .D(n92), .SI(g3188), .SE(n9298), .CLK(n9485), .Q(
        g3133), .QN(n8696) );
  SDFFX1 DFF_140_Q_reg ( .D(g26104), .SI(g3133), .SE(n9299), .CLK(n9486), .Q(
        n8087), .QN(DFF_140_n1) );
  SDFFX1 DFF_141_Q_reg ( .D(n276), .SI(n8087), .SE(n9299), .CLK(n9486), .Q(
        g3128) );
  SDFFX1 DFF_142_Q_reg ( .D(g26149), .SI(g3128), .SE(n9299), .CLK(n9486), .Q(
        n8086) );
  SDFFX1 DFF_143_Q_reg ( .D(g25420), .SI(n8086), .SE(n9422), .CLK(n9609), .Q(
        test_so9), .QN(n8595) );
  SDFFX1 DFF_144_Q_reg ( .D(n299), .SI(test_si10), .SE(n9422), .CLK(n9609), 
        .Q(n8084) );
  SDFFX1 DFF_145_Q_reg ( .D(g25442), .SI(n8084), .SE(n9299), .CLK(n9486), .Q(
        g3124), .QN(n8597) );
  SDFFX1 DFF_146_Q_reg ( .D(n307), .SI(g3124), .SE(n9299), .CLK(n9486), .Q(
        n8083), .QN(DFF_146_n1) );
  SDFFX1 DFF_147_Q_reg ( .D(g26104), .SI(n8083), .SE(n9299), .CLK(n9486), .Q(
        n8082), .QN(n16830) );
  SDFFX1 DFF_148_Q_reg ( .D(g26135), .SI(n8082), .SE(n9299), .CLK(n9486), .Q(
        n8081), .QN(n16831) );
  SDFFX1 DFF_149_Q_reg ( .D(g26149), .SI(n8081), .SE(n9299), .CLK(n9486), .Q(
        n8080) );
  SDFFX1 DFF_150_Q_reg ( .D(g25420), .SI(n8080), .SE(n9299), .CLK(n9486), .Q(
        g3112), .QN(n8596) );
  SDFFX1 DFF_151_Q_reg ( .D(g25435), .SI(g3112), .SE(n9300), .CLK(n9487), .Q(
        g3110), .QN(n8563) );
  SDFFX1 DFF_152_Q_reg ( .D(g25442), .SI(g3110), .SE(n9300), .CLK(n9487), .Q(
        g3111), .QN(n8598) );
  SDFFX1 DFF_153_Q_reg ( .D(g27380), .SI(g3111), .SE(n9300), .CLK(n9487), .Q(
        n8079), .QN(n16825) );
  SDFFX1 DFF_154_Q_reg ( .D(g26104), .SI(n8079), .SE(n9300), .CLK(n9487), .Q(
        n8078), .QN(n16832) );
  SDFFX1 DFF_155_Q_reg ( .D(g26135), .SI(n8078), .SE(n9300), .CLK(n9487), .Q(
        n8077), .QN(DFF_155_n1) );
  SDFFX1 DFF_156_Q_reg ( .D(g26149), .SI(n8077), .SE(n9300), .CLK(n9487), .Q(
        n8076), .QN(DFF_156_n1) );
  SDFFX1 DFF_157_Q_reg ( .D(g27380), .SI(n8076), .SE(n9300), .CLK(n9487), .Q(
        g3151), .QN(n4424) );
  SDFFX1 DFF_158_Q_reg ( .D(g26104), .SI(g3151), .SE(n9300), .CLK(n9487), .Q(
        g3142), .QN(n4301) );
  SDFFX1 DFF_159_Q_reg ( .D(g26135), .SI(g3142), .SE(n9300), .CLK(n9487), .Q(
        test_so10), .QN(n9287) );
  SDFFX1 DFF_160_Q_reg ( .D(n92), .SI(test_si11), .SE(n9298), .CLK(n9485), .Q(
        g185), .QN(n4384) );
  SDFFX1 DFF_161_Q_reg ( .D(g2950), .SI(g185), .SE(n9298), .CLK(n9485), .Q(
        g6231), .QN(n4318) );
  SDFFX1 DFF_162_Q_reg ( .D(g6231), .SI(g6231), .SE(n9298), .CLK(n9485), .Q(
        g6313), .QN(n4512) );
  SDFFX1 DFF_163_Q_reg ( .D(g6313), .SI(g6313), .SE(n9298), .CLK(n9485), .Q(
        g165), .QN(n4369) );
  SDFFX1 DFF_164_Q_reg ( .D(g22100), .SI(g165), .SE(n9312), .CLK(n9499), .Q(
        g130) );
  SDFFX1 DFF_165_Q_reg ( .D(g22122), .SI(g130), .SE(n9312), .CLK(n9499), .Q(
        g131), .QN(n9214) );
  SDFFX1 DFF_166_Q_reg ( .D(g22141), .SI(g131), .SE(n9312), .CLK(n9499), .Q(
        g129) );
  SDFFX1 DFF_167_Q_reg ( .D(g22123), .SI(g129), .SE(n9313), .CLK(n9500), .Q(
        g133) );
  SDFFX1 DFF_168_Q_reg ( .D(g22142), .SI(g133), .SE(n9313), .CLK(n9500), .Q(
        g134), .QN(n9212) );
  SDFFX1 DFF_169_Q_reg ( .D(g22161), .SI(g134), .SE(n9313), .CLK(n9500), .Q(
        g132) );
  SDFFX1 DFF_170_Q_reg ( .D(g22025), .SI(g132), .SE(n9313), .CLK(n9500), .Q(
        g142) );
  SDFFX1 DFF_171_Q_reg ( .D(g22027), .SI(g142), .SE(n9313), .CLK(n9500), .Q(
        g143), .QN(n9210) );
  SDFFX1 DFF_172_Q_reg ( .D(g22030), .SI(g143), .SE(n9313), .CLK(n9500), .Q(
        g141) );
  SDFFX1 DFF_173_Q_reg ( .D(g22028), .SI(g141), .SE(n9313), .CLK(n9500), .Q(
        g145) );
  SDFFX1 DFF_174_Q_reg ( .D(g22031), .SI(g145), .SE(n9313), .CLK(n9500), .Q(
        g146), .QN(n9208) );
  SDFFX1 DFF_175_Q_reg ( .D(g22037), .SI(g146), .SE(n9313), .CLK(n9500), .Q(
        test_so11) );
  SDFFX1 DFF_176_Q_reg ( .D(g22032), .SI(test_si12), .SE(n9311), .CLK(n9498), 
        .Q(g148) );
  SDFFX1 DFF_177_Q_reg ( .D(g22038), .SI(g148), .SE(n9311), .CLK(n9498), .Q(
        g149), .QN(n9206) );
  SDFFX1 DFF_178_Q_reg ( .D(g22047), .SI(g149), .SE(n9311), .CLK(n9498), .Q(
        g147) );
  SDFFX1 DFF_179_Q_reg ( .D(g22039), .SI(g147), .SE(n9312), .CLK(n9499), .Q(
        g151) );
  SDFFX1 DFF_180_Q_reg ( .D(g22048), .SI(g151), .SE(n9312), .CLK(n9499), .Q(
        g152), .QN(n9204) );
  SDFFX1 DFF_181_Q_reg ( .D(g22063), .SI(g152), .SE(n9312), .CLK(n9499), .Q(
        g150) );
  SDFFX1 DFF_182_Q_reg ( .D(g22049), .SI(g150), .SE(n9312), .CLK(n9499), .Q(
        g154) );
  SDFFX1 DFF_183_Q_reg ( .D(g22064), .SI(g154), .SE(n9312), .CLK(n9499), .Q(
        g155), .QN(n9202) );
  SDFFX1 DFF_184_Q_reg ( .D(g22079), .SI(g155), .SE(n9312), .CLK(n9499), .Q(
        g153) );
  SDFFX1 DFF_185_Q_reg ( .D(g22065), .SI(g153), .SE(n9308), .CLK(n9495), .Q(
        g157) );
  SDFFX1 DFF_186_Q_reg ( .D(g22080), .SI(g157), .SE(n9310), .CLK(n9497), .Q(
        g158), .QN(n9200) );
  SDFFX1 DFF_187_Q_reg ( .D(g22101), .SI(g158), .SE(n9310), .CLK(n9497), .Q(
        g156) );
  SDFFX1 DFF_188_Q_reg ( .D(g22081), .SI(g156), .SE(n9312), .CLK(n9499), .Q(
        g160), .QN(n8792) );
  SDFFX1 DFF_189_Q_reg ( .D(g22102), .SI(g160), .SE(n9312), .CLK(n9499), .Q(
        g161) );
  SDFFX1 DFF_190_Q_reg ( .D(g22124), .SI(g161), .SE(n9312), .CLK(n9499), .Q(
        g159), .QN(n8790) );
  SDFFX1 DFF_191_Q_reg ( .D(g22103), .SI(g159), .SE(n9313), .CLK(n9500), .Q(
        test_so12) );
  SDFFX1 DFF_192_Q_reg ( .D(g22125), .SI(test_si13), .SE(n9310), .CLK(n9497), 
        .Q(g164) );
  SDFFX1 DFF_193_Q_reg ( .D(g22143), .SI(g164), .SE(n9310), .CLK(n9497), .Q(
        g162), .QN(n8828) );
  SDFFX1 DFF_194_Q_reg ( .D(g25204), .SI(g162), .SE(n9310), .CLK(n9497), .Q(
        g169) );
  SDFFX1 DFF_195_Q_reg ( .D(g25206), .SI(g169), .SE(n9310), .CLK(n9497), .Q(
        g170), .QN(n8893) );
  SDFFX1 DFF_196_Q_reg ( .D(g25211), .SI(g170), .SE(n9310), .CLK(n9497), .Q(
        g168) );
  SDFFX1 DFF_197_Q_reg ( .D(g25207), .SI(g168), .SE(n9311), .CLK(n9498), .Q(
        g172) );
  SDFFX1 DFF_198_Q_reg ( .D(g25212), .SI(g172), .SE(n9311), .CLK(n9498), .Q(
        g173), .QN(n8890) );
  SDFFX1 DFF_199_Q_reg ( .D(g25218), .SI(g173), .SE(n9311), .CLK(n9498), .Q(
        g171) );
  SDFFX1 DFF_200_Q_reg ( .D(g25213), .SI(g171), .SE(n9311), .CLK(n9498), .Q(
        g175) );
  SDFFX1 DFF_201_Q_reg ( .D(g25219), .SI(g175), .SE(n9311), .CLK(n9498), .Q(
        g176), .QN(n8887) );
  SDFFX1 DFF_202_Q_reg ( .D(g25228), .SI(g176), .SE(n9311), .CLK(n9498), .Q(
        g174) );
  SDFFX1 DFF_203_Q_reg ( .D(g25220), .SI(g174), .SE(n9311), .CLK(n9498), .Q(
        g178) );
  SDFFX1 DFF_204_Q_reg ( .D(g25229), .SI(g178), .SE(n9311), .CLK(n9498), .Q(
        g179), .QN(n8884) );
  SDFFX1 DFF_205_Q_reg ( .D(g25239), .SI(g179), .SE(n9311), .CLK(n9498), .Q(
        g177) );
  SDFFX1 DFF_206_Q_reg ( .D(g30261), .SI(g177), .SE(n9318), .CLK(n9505), .Q(
        g186), .QN(n8482) );
  SDFFX1 DFF_207_Q_reg ( .D(g30267), .SI(g186), .SE(n9318), .CLK(n9505), .Q(
        test_so13) );
  SDFFX1 DFF_208_Q_reg ( .D(g30275), .SI(test_si14), .SE(n9319), .CLK(n9506), 
        .Q(g192), .QN(n8546) );
  SDFFX1 DFF_209_Q_reg ( .D(g30637), .SI(g192), .SE(n9319), .CLK(n9506), .Q(
        g231), .QN(n8481) );
  SDFFX1 DFF_210_Q_reg ( .D(g30640), .SI(g231), .SE(n9319), .CLK(n9506), .Q(
        g234) );
  SDFFX1 DFF_211_Q_reg ( .D(g30645), .SI(g234), .SE(n9319), .CLK(n9506), .Q(
        g237), .QN(n8429) );
  SDFFX1 DFF_212_Q_reg ( .D(g30668), .SI(g237), .SE(n9319), .CLK(n9506), .Q(
        g195), .QN(n8480) );
  SDFFX1 DFF_213_Q_reg ( .D(g30674), .SI(g195), .SE(n9319), .CLK(n9506), .Q(
        g198) );
  SDFFX1 DFF_214_Q_reg ( .D(g30680), .SI(g198), .SE(n9308), .CLK(n9495), .Q(
        g201), .QN(n8545) );
  SDFFX1 DFF_215_Q_reg ( .D(g30641), .SI(g201), .SE(n9319), .CLK(n9506), .Q(
        g240), .QN(n8478) );
  SDFFX1 DFF_216_Q_reg ( .D(g30646), .SI(g240), .SE(n9319), .CLK(n9506), .Q(
        g243) );
  SDFFX1 DFF_217_Q_reg ( .D(g30653), .SI(g243), .SE(n9319), .CLK(n9506), .Q(
        g246), .QN(n8428) );
  SDFFX1 DFF_218_Q_reg ( .D(g30276), .SI(g246), .SE(n9319), .CLK(n9506), .Q(
        g204), .QN(n8477) );
  SDFFX1 DFF_219_Q_reg ( .D(g30284), .SI(g204), .SE(n9319), .CLK(n9506), .Q(
        g207) );
  SDFFX1 DFF_220_Q_reg ( .D(g30292), .SI(g207), .SE(n9319), .CLK(n9506), .Q(
        g210), .QN(n8534) );
  SDFFX1 DFF_221_Q_reg ( .D(g30254), .SI(g210), .SE(n9320), .CLK(n9507), .Q(
        g249), .QN(n8475) );
  SDFFX1 DFF_222_Q_reg ( .D(g30257), .SI(g249), .SE(n9320), .CLK(n9507), .Q(
        g252) );
  SDFFX1 DFF_223_Q_reg ( .D(g30262), .SI(g252), .SE(n9320), .CLK(n9507), .Q(
        test_so14) );
  SDFFX1 DFF_224_Q_reg ( .D(g30245), .SI(test_si15), .SE(n9320), .CLK(n9507), 
        .Q(g213), .QN(n8473) );
  SDFFX1 DFF_225_Q_reg ( .D(g30246), .SI(g213), .SE(n9320), .CLK(n9507), .Q(
        g216) );
  SDFFX1 DFF_226_Q_reg ( .D(g30248), .SI(g216), .SE(n9320), .CLK(n9507), .Q(
        g219), .QN(n8544) );
  SDFFX1 DFF_227_Q_reg ( .D(g30258), .SI(g219), .SE(n9320), .CLK(n9507), .Q(
        g258), .QN(n8471) );
  SDFFX1 DFF_228_Q_reg ( .D(g30263), .SI(g258), .SE(n9320), .CLK(n9507), .Q(
        g261) );
  SDFFX1 DFF_229_Q_reg ( .D(g30268), .SI(g261), .SE(n9320), .CLK(n9507), .Q(
        g264), .QN(n8529) );
  SDFFX1 DFF_230_Q_reg ( .D(g30635), .SI(g264), .SE(n9320), .CLK(n9507), .Q(
        g222), .QN(n8380) );
  SDFFX1 DFF_231_Q_reg ( .D(g30636), .SI(g222), .SE(n9320), .CLK(n9507), .Q(
        g225) );
  SDFFX1 DFF_232_Q_reg ( .D(g30639), .SI(g225), .SE(n9320), .CLK(n9507), .Q(
        g228), .QN(n8386) );
  SDFFX1 DFF_233_Q_reg ( .D(g30661), .SI(g228), .SE(n9321), .CLK(n9508), .Q(
        g267), .QN(n8415) );
  SDFFX1 DFF_234_Q_reg ( .D(g30669), .SI(g267), .SE(n9321), .CLK(n9508), .Q(
        g270) );
  SDFFX1 DFF_235_Q_reg ( .D(g30675), .SI(g270), .SE(n9308), .CLK(n9495), .Q(
        g273), .QN(n8416) );
  SDFFX1 DFF_236_Q_reg ( .D(g25027), .SI(g273), .SE(n9308), .CLK(n9495), .Q(
        g92), .QN(n8984) );
  SDFFX1 DFF_237_Q_reg ( .D(n46), .SI(g92), .SE(n9308), .CLK(n9495), .Q(g88), 
        .QN(n9264) );
  SDFFX1 DFF_238_Q_reg ( .D(g26529), .SI(g88), .SE(n9308), .CLK(n9495), .Q(g83), .QN(n8983) );
  SDFFX1 DFF_239_Q_reg ( .D(n47), .SI(g83), .SE(n9308), .CLK(n9495), .Q(
        test_so15) );
  SDFFX1 DFF_240_Q_reg ( .D(g27594), .SI(test_si16), .SE(n9308), .CLK(n9495), 
        .Q(g74), .QN(n8982) );
  SDFFX1 DFF_241_Q_reg ( .D(g28145), .SI(g74), .SE(n9309), .CLK(n9496), .Q(g70), .QN(n9275) );
  SDFFX1 DFF_242_Q_reg ( .D(g28634), .SI(g70), .SE(n9309), .CLK(n9496), .Q(g65), .QN(n8981) );
  SDFFX1 DFF_243_Q_reg ( .D(g29109), .SI(g65), .SE(n9309), .CLK(n9496), .Q(g61), .QN(n9266) );
  SDFFX1 DFF_244_Q_reg ( .D(g29353), .SI(g61), .SE(n9309), .CLK(n9496), .Q(g56), .QN(n8562) );
  SDFFX1 DFF_245_Q_reg ( .D(g29579), .SI(g56), .SE(n9309), .CLK(n9496), .Q(g52), .QN(n8391) );
  SDFFX1 DFF_246_Q_reg ( .D(n15), .SI(g52), .SE(n9309), .CLK(n9496), .Q(g180)
         );
  SDFFX1 DFF_247_Q_reg ( .D(g180), .SI(g180), .SE(n9309), .CLK(n9496), .Q(
        g5549) );
  SDFFX1 DFF_248_Q_reg ( .D(g5549), .SI(g5549), .SE(n9309), .CLK(n9496), .Q(
        g181), .QN(n8991) );
  SDFFX1 DFF_251_Q_reg ( .D(g6447), .SI(g6447), .SE(n9309), .CLK(n9496), .Q(
        n4640), .QN(n4506) );
  SDFFX1 DFF_252_Q_reg ( .D(g5549), .SI(n4640), .SE(n9309), .CLK(n9496), .Q(
        g309), .QN(n4388) );
  SDFFX1 DFF_253_Q_reg ( .D(g27253), .SI(g309), .SE(n9316), .CLK(n9503), .Q(
        g354), .QN(n8935) );
  SDFFX1 DFF_254_Q_reg ( .D(g27255), .SI(g354), .SE(n9316), .CLK(n9503), .Q(
        g343) );
  SDFFX1 DFF_255_Q_reg ( .D(g27258), .SI(g343), .SE(n9316), .CLK(n9503), .Q(
        test_so16) );
  SDFFX1 DFF_256_Q_reg ( .D(g27256), .SI(test_si17), .SE(n9316), .CLK(n9503), 
        .Q(g369), .QN(n8913) );
  SDFFX1 DFF_257_Q_reg ( .D(g27259), .SI(g369), .SE(n9316), .CLK(n9503), .Q(
        g358) );
  SDFFX1 DFF_258_Q_reg ( .D(g27265), .SI(g358), .SE(n9316), .CLK(n9503), .Q(
        g361) );
  SDFFX1 DFF_259_Q_reg ( .D(g27260), .SI(g361), .SE(n9316), .CLK(n9503), .Q(
        g384), .QN(n8643) );
  SDFFX1 DFF_260_Q_reg ( .D(g27266), .SI(g384), .SE(n9316), .CLK(n9503), .Q(
        g373) );
  SDFFX1 DFF_261_Q_reg ( .D(g27277), .SI(g373), .SE(n9315), .CLK(n9502), .Q(
        g376) );
  SDFFX1 DFF_262_Q_reg ( .D(g27267), .SI(g376), .SE(n9318), .CLK(n9505), .Q(
        g398), .QN(n8924) );
  SDFFX1 DFF_263_Q_reg ( .D(g27278), .SI(g398), .SE(n9318), .CLK(n9505), .Q(
        g388) );
  SDFFX1 DFF_264_Q_reg ( .D(g27293), .SI(g388), .SE(n9314), .CLK(n9501), .Q(
        g391) );
  SDFFX1 DFF_265_Q_reg ( .D(g28732), .SI(g391), .SE(n9314), .CLK(n9501), .Q(
        g408) );
  SDFFX1 DFF_266_Q_reg ( .D(g28735), .SI(g408), .SE(n9315), .CLK(n9502), .Q(
        g411), .QN(n8743) );
  SDFFX1 DFF_267_Q_reg ( .D(g28744), .SI(g411), .SE(n9315), .CLK(n9502), .Q(
        g414), .QN(n8742) );
  SDFFX1 DFF_268_Q_reg ( .D(g29194), .SI(g414), .SE(n9315), .CLK(n9502), .Q(
        g417) );
  SDFFX1 DFF_269_Q_reg ( .D(g29197), .SI(g417), .SE(n9315), .CLK(n9502), .Q(
        g420), .QN(n8740) );
  SDFFX1 DFF_270_Q_reg ( .D(g29201), .SI(g420), .SE(n9314), .CLK(n9501), .Q(
        g423), .QN(n8739) );
  SDFFX1 DFF_271_Q_reg ( .D(g28736), .SI(g423), .SE(n9314), .CLK(n9501), .Q(
        test_so17), .QN(n9289) );
  SDFFX1 DFF_272_Q_reg ( .D(g28745), .SI(test_si18), .SE(n9314), .CLK(n9501), 
        .Q(g428) );
  SDFFX1 DFF_273_Q_reg ( .D(g28754), .SI(g428), .SE(n9314), .CLK(n9501), .Q(
        g426) );
  SDFFX1 DFF_274_Q_reg ( .D(g26803), .SI(g426), .SE(n9314), .CLK(n9501), .Q(
        g429) );
  SDFFX1 DFF_275_Q_reg ( .D(g26804), .SI(g429), .SE(n9314), .CLK(n9501), .Q(
        g432), .QN(n8737) );
  SDFFX1 DFF_276_Q_reg ( .D(g26807), .SI(g432), .SE(n9314), .CLK(n9501), .Q(
        g435), .QN(n8736) );
  SDFFX1 DFF_277_Q_reg ( .D(g26805), .SI(g435), .SE(n9315), .CLK(n9502), .Q(
        g438) );
  SDFFX1 DFF_278_Q_reg ( .D(g26808), .SI(g438), .SE(n9315), .CLK(n9502), .Q(
        g441), .QN(n8734) );
  SDFFX1 DFF_279_Q_reg ( .D(g26812), .SI(g441), .SE(n9315), .CLK(n9502), .Q(
        g444), .QN(n8733) );
  SDFFX1 DFF_280_Q_reg ( .D(g27759), .SI(g444), .SE(n9315), .CLK(n9502), .Q(
        g448), .QN(n8965) );
  SDFFX1 DFF_281_Q_reg ( .D(g27760), .SI(g448), .SE(n9315), .CLK(n9502), .Q(
        g449), .QN(n8964) );
  SDFFX1 DFF_282_Q_reg ( .D(g27762), .SI(g449), .SE(n9314), .CLK(n9501), .Q(
        g447), .QN(n8963) );
  SDFFX1 DFF_283_Q_reg ( .D(g29606), .SI(g447), .SE(n9314), .CLK(n9501), .Q(
        g312), .QN(n8526) );
  SDFFX1 DFF_284_Q_reg ( .D(g29608), .SI(g312), .SE(n9315), .CLK(n9502), .Q(
        g313) );
  SDFFX1 DFF_285_Q_reg ( .D(g29611), .SI(g313), .SE(n9313), .CLK(n9500), .Q(
        g314) );
  SDFFX1 DFF_286_Q_reg ( .D(g30699), .SI(g314), .SE(n9313), .CLK(n9500), .Q(
        g315), .QN(n8523) );
  SDFFX1 DFF_287_Q_reg ( .D(g30700), .SI(g315), .SE(n9314), .CLK(n9501), .Q(
        test_so18) );
  SDFFX1 DFF_288_Q_reg ( .D(g30702), .SI(test_si19), .SE(n9308), .CLK(n9495), 
        .Q(g317) );
  SDFFX1 DFF_289_Q_reg ( .D(g30455), .SI(g317), .SE(n9310), .CLK(n9497), .Q(
        g318), .QN(n8521) );
  SDFFX1 DFF_290_Q_reg ( .D(g30468), .SI(g318), .SE(n9310), .CLK(n9497), .Q(
        g319) );
  SDFFX1 DFF_291_Q_reg ( .D(g30482), .SI(g319), .SE(n9308), .CLK(n9495), .Q(
        g320) );
  SDFFX1 DFF_292_Q_reg ( .D(g29167), .SI(g320), .SE(n9321), .CLK(n9508), .Q(
        g322), .QN(n8558) );
  SDFFX1 DFF_293_Q_reg ( .D(g29169), .SI(g322), .SE(n9321), .CLK(n9508), .Q(
        g323) );
  SDFFX1 DFF_294_Q_reg ( .D(g29172), .SI(g323), .SE(n9308), .CLK(n9495), .Q(
        g321) );
  SDFFX1 DFF_295_Q_reg ( .D(g26655), .SI(g321), .SE(n9310), .CLK(n9497), .Q(
        g403), .QN(n8962) );
  SDFFX1 DFF_296_Q_reg ( .D(g26659), .SI(g403), .SE(n9310), .CLK(n9497), .Q(
        g404) );
  SDFFX1 DFF_297_Q_reg ( .D(g26664), .SI(g404), .SE(n9310), .CLK(n9497), .Q(
        g402) );
  SDFFX1 DFF_298_Q_reg ( .D(n4290), .SI(g402), .SE(n9321), .CLK(n9508), .Q(
        g450) );
  SDFFX1 DFF_299_Q_reg ( .D(g450), .SI(g450), .SE(n9321), .CLK(n9508), .Q(
        n8066), .QN(DFF_299_n1) );
  SDFFX1 DFF_300_Q_reg ( .D(n4569), .SI(n8066), .SE(n9321), .CLK(n9508), .Q(
        g452) );
  SDFFX1 DFF_301_Q_reg ( .D(g452), .SI(g452), .SE(n9321), .CLK(n9508), .Q(
        n8065), .QN(DFF_301_n1) );
  SDFFX1 DFF_302_Q_reg ( .D(n4561), .SI(n8065), .SE(n9321), .CLK(n9508), .Q(
        g454) );
  SDFFX1 DFF_303_Q_reg ( .D(g454), .SI(g454), .SE(n9321), .CLK(n9508), .Q(
        test_so19), .QN(DFF_303_n1) );
  SDFFX1 DFF_304_Q_reg ( .D(n4328), .SI(test_si20), .SE(n9306), .CLK(n9493), 
        .Q(g280) );
  SDFFX1 DFF_305_Q_reg ( .D(g280), .SI(g280), .SE(n9306), .CLK(n9493), .Q(
        n8062), .QN(DFF_305_n1) );
  SDFFX1 DFF_306_Q_reg ( .D(n4392), .SI(n8062), .SE(n9307), .CLK(n9494), .Q(
        g282) );
  SDFFX1 DFF_307_Q_reg ( .D(g282), .SI(g282), .SE(n9307), .CLK(n9494), .Q(
        n8061), .QN(DFF_307_n1) );
  SDFFX1 DFF_308_Q_reg ( .D(n4322), .SI(n8061), .SE(n9307), .CLK(n9494), .Q(
        g284) );
  SDFFX1 DFF_309_Q_reg ( .D(g284), .SI(g284), .SE(n9307), .CLK(n9494), .Q(
        n8060), .QN(DFF_309_n1) );
  SDFFX1 DFF_310_Q_reg ( .D(n4376), .SI(n8060), .SE(n9307), .CLK(n9494), .Q(
        g286) );
  SDFFX1 DFF_311_Q_reg ( .D(g286), .SI(g286), .SE(n9307), .CLK(n9494), .Q(
        n8059), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(n4380), .SI(n8059), .SE(n9307), .CLK(n9494), .Q(
        g288) );
  SDFFX1 DFF_313_Q_reg ( .D(g288), .SI(g288), .SE(n9307), .CLK(n9494), .Q(
        n8058), .QN(DFF_313_n1) );
  SDFFX1 DFF_314_Q_reg ( .D(g2857), .SI(n8058), .SE(n9307), .CLK(n9494), .Q(
        g290) );
  SDFFX1 DFF_315_Q_reg ( .D(g290), .SI(g290), .SE(n9307), .CLK(n9494), .Q(
        n8057), .QN(n4485) );
  SDFFX1 DFF_316_Q_reg ( .D(n4282), .SI(n8057), .SE(n9315), .CLK(n9502), .Q(
        n8056), .QN(n16833) );
  SDFFX1 DFF_317_Q_reg ( .D(g21346), .SI(n8056), .SE(n9297), .CLK(n9484), .Q(
        g305), .QN(n8699) );
  SDFFX1 DFF_328_Q_reg ( .D(n4278), .SI(g305), .SE(n9297), .CLK(n9484), .Q(
        n8055), .QN(DFF_328_n1) );
  SDFFX1 DFF_329_Q_reg ( .D(g354), .SI(n8055), .SE(n9316), .CLK(n9503), .Q(
        test_so20) );
  SDFFX1 DFF_330_Q_reg ( .D(test_so20), .SI(test_si21), .SE(n9316), .CLK(n9503), .Q(g349) );
  SDFFX1 DFF_331_Q_reg ( .D(g343), .SI(g349), .SE(n9316), .CLK(n9503), .Q(g350) );
  SDFFX1 DFF_332_Q_reg ( .D(g350), .SI(g350), .SE(n9316), .CLK(n9503), .Q(g351), .QN(n8620) );
  SDFFX1 DFF_333_Q_reg ( .D(test_so16), .SI(g351), .SE(n9317), .CLK(n9504), 
        .Q(g352) );
  SDFFX1 DFF_334_Q_reg ( .D(g352), .SI(g352), .SE(n9317), .CLK(n9504), .Q(g353), .QN(n8619) );
  SDFFX1 DFF_335_Q_reg ( .D(g369), .SI(g353), .SE(n9317), .CLK(n9504), .Q(g357) );
  SDFFX1 DFF_336_Q_reg ( .D(g357), .SI(g357), .SE(n9317), .CLK(n9504), .Q(g364) );
  SDFFX1 DFF_337_Q_reg ( .D(g358), .SI(g364), .SE(n9317), .CLK(n9504), .Q(g365) );
  SDFFX1 DFF_338_Q_reg ( .D(g365), .SI(g365), .SE(n9317), .CLK(n9504), .Q(g366), .QN(n8409) );
  SDFFX1 DFF_339_Q_reg ( .D(g361), .SI(g366), .SE(n9317), .CLK(n9504), .Q(g367) );
  SDFFX1 DFF_340_Q_reg ( .D(g367), .SI(g367), .SE(n9317), .CLK(n9504), .Q(g368), .QN(n8408) );
  SDFFX1 DFF_341_Q_reg ( .D(g384), .SI(g368), .SE(n9317), .CLK(n9504), .Q(g372) );
  SDFFX1 DFF_342_Q_reg ( .D(g372), .SI(g372), .SE(n9317), .CLK(n9504), .Q(g379) );
  SDFFX1 DFF_343_Q_reg ( .D(g373), .SI(g379), .SE(n9317), .CLK(n9504), .Q(g380) );
  SDFFX1 DFF_344_Q_reg ( .D(g380), .SI(g380), .SE(n9317), .CLK(n9504), .Q(g381), .QN(n8583) );
  SDFFX1 DFF_345_Q_reg ( .D(g376), .SI(g381), .SE(n9318), .CLK(n9505), .Q(
        test_so21) );
  SDFFX1 DFF_346_Q_reg ( .D(test_so21), .SI(test_si22), .SE(n9318), .CLK(n9505), .Q(g383), .QN(n8582) );
  SDFFX1 DFF_347_Q_reg ( .D(g398), .SI(g383), .SE(n9318), .CLK(n9505), .Q(g387) );
  SDFFX1 DFF_348_Q_reg ( .D(g387), .SI(g387), .SE(n9318), .CLK(n9505), .Q(g394), .QN(n16823) );
  SDFFX1 DFF_349_Q_reg ( .D(g388), .SI(g394), .SE(n9318), .CLK(n9505), .Q(g395) );
  SDFFX1 DFF_350_Q_reg ( .D(g395), .SI(g395), .SE(n9318), .CLK(n9505), .Q(g396) );
  SDFFX1 DFF_351_Q_reg ( .D(g391), .SI(g396), .SE(n9318), .CLK(n9505), .Q(g397) );
  SDFFX1 DFF_352_Q_reg ( .D(g397), .SI(g397), .SE(n9318), .CLK(n9505), .Q(g324), .QN(n8632) );
  SDFFX1 DFF_353_Q_reg ( .D(n4598), .SI(g324), .SE(n9324), .CLK(n9511), .Q(
        g5629), .QN(n8630) );
  SDFFX1 DFF_354_Q_reg ( .D(g5629), .SI(g5629), .SE(n9324), .CLK(n9511), .Q(
        g5648), .QN(n8633) );
  SDFFX1 DFF_355_Q_reg ( .D(g5648), .SI(g5648), .SE(n9324), .CLK(n9511), .Q(
        g337), .QN(n8631) );
  SDFFX1 DFF_356_Q_reg ( .D(n4598), .SI(g337), .SE(n9324), .CLK(n9511), .Q(
        g6485), .QN(n4298) );
  SDFFX1 DFF_357_Q_reg ( .D(g6485), .SI(g6485), .SE(n9324), .CLK(n9511), .Q(
        g6642), .QN(n4372) );
  SDFFX1 DFF_358_Q_reg ( .D(g6642), .SI(g6642), .SE(n9324), .CLK(n9511), .Q(
        g550), .QN(n4313) );
  SDFFX1 DFF_359_Q_reg ( .D(n552), .SI(g550), .SE(n9325), .CLK(n9512), .Q(g554), .QN(n9226) );
  SDFFX1 DFF_360_Q_reg ( .D(g18678), .SI(g554), .SE(n9325), .CLK(n9512), .Q(
        g557), .QN(n4360) );
  SDFFX1 DFF_361_Q_reg ( .D(g18726), .SI(g557), .SE(n9325), .CLK(n9512), .Q(
        test_so22), .QN(n9285) );
  SDFFX1 DFF_362_Q_reg ( .D(n541), .SI(test_si23), .SE(n9325), .CLK(n9512), 
        .Q(g513) );
  SDFFX1 DFF_363_Q_reg ( .D(g513), .SI(g513), .SE(n9325), .CLK(n9512), .Q(g523) );
  SDFFX1 DFF_364_Q_reg ( .D(g523), .SI(g523), .SE(n9325), .CLK(n9512), .Q(g524) );
  SDFFX1 DFF_365_Q_reg ( .D(g455), .SI(g524), .SE(n9325), .CLK(n9512), .Q(g564) );
  SDFFX1 DFF_366_Q_reg ( .D(g564), .SI(g564), .SE(n9325), .CLK(n9512), .Q(g569), .QN(n8766) );
  SDFFX1 DFF_367_Q_reg ( .D(g458), .SI(g569), .SE(n9325), .CLK(n9512), .Q(g570) );
  SDFFX1 DFF_368_Q_reg ( .D(g570), .SI(g570), .SE(n9325), .CLK(n9512), .Q(g571) );
  SDFFX1 DFF_369_Q_reg ( .D(g461), .SI(g571), .SE(n9325), .CLK(n9512), .Q(g572) );
  SDFFX1 DFF_370_Q_reg ( .D(g572), .SI(g572), .SE(n9326), .CLK(n9513), .Q(g573), .QN(n8767) );
  SDFFX1 DFF_371_Q_reg ( .D(g465), .SI(g573), .SE(n9326), .CLK(n9513), .Q(g574) );
  SDFFX1 DFF_372_Q_reg ( .D(g574), .SI(g574), .SE(n9326), .CLK(n9513), .Q(g565), .QN(n8764) );
  SDFFX1 DFF_373_Q_reg ( .D(test_so24), .SI(g565), .SE(n9326), .CLK(n9513), 
        .Q(g566) );
  SDFFX1 DFF_374_Q_reg ( .D(g566), .SI(g566), .SE(n9326), .CLK(n9513), .Q(g567) );
  SDFFX1 DFF_375_Q_reg ( .D(g471), .SI(g567), .SE(n9326), .CLK(n9513), .Q(g568) );
  SDFFX1 DFF_376_Q_reg ( .D(g568), .SI(g568), .SE(n9326), .CLK(n9513), .Q(g489), .QN(n8765) );
  SDFFX1 DFF_377_Q_reg ( .D(g2950), .SI(g489), .SE(n9326), .CLK(n9513), .Q(
        test_so23), .QN(n9286) );
  SDFFX1 DFF_378_Q_reg ( .D(test_so23), .SI(test_si24), .SE(n9326), .CLK(n9513), .Q(g7956), .QN(n4461) );
  SDFFX1 DFF_379_Q_reg ( .D(g7956), .SI(g7956), .SE(n9326), .CLK(n9513), .Q(
        g485), .QN(n4466) );
  SDFFX1 DFF_380_Q_reg ( .D(g23067), .SI(g485), .SE(n9326), .CLK(n9513), .Q(
        g486), .QN(n9021) );
  SDFFX1 DFF_381_Q_reg ( .D(g23093), .SI(g486), .SE(n9327), .CLK(n9514), .Q(
        g487) );
  SDFFX1 DFF_382_Q_reg ( .D(g23117), .SI(g487), .SE(n9327), .CLK(n9514), .Q(
        g488), .QN(n9022) );
  SDFFX1 DFF_383_Q_reg ( .D(g23385), .SI(g488), .SE(n9327), .CLK(n9514), .Q(
        g455) );
  SDFFX1 DFF_384_Q_reg ( .D(g23399), .SI(g455), .SE(n9327), .CLK(n9514), .Q(
        g458) );
  SDFFX1 DFF_385_Q_reg ( .D(g24174), .SI(g458), .SE(n9327), .CLK(n9514), .Q(
        g461) );
  SDFFX1 DFF_386_Q_reg ( .D(g24178), .SI(g461), .SE(n9327), .CLK(n9514), .Q(
        g477), .QN(n9027) );
  SDFFX1 DFF_387_Q_reg ( .D(g24207), .SI(g477), .SE(n9327), .CLK(n9514), .Q(
        g478) );
  SDFFX1 DFF_388_Q_reg ( .D(g24216), .SI(g478), .SE(n9327), .CLK(n9514), .Q(
        g479), .QN(n9028) );
  SDFFX1 DFF_389_Q_reg ( .D(g23092), .SI(g479), .SE(n9327), .CLK(n9514), .Q(
        g480), .QN(n9024) );
  SDFFX1 DFF_390_Q_reg ( .D(g23000), .SI(g480), .SE(n9327), .CLK(n9514), .Q(
        g484) );
  SDFFX1 DFF_391_Q_reg ( .D(g23022), .SI(g484), .SE(n9327), .CLK(n9514), .Q(
        g464), .QN(n9025) );
  SDFFX1 DFF_392_Q_reg ( .D(g24206), .SI(g464), .SE(n9327), .CLK(n9514), .Q(
        g465) );
  SDFFX1 DFF_393_Q_reg ( .D(g24215), .SI(g465), .SE(n9328), .CLK(n9515), .Q(
        test_so24) );
  SDFFX1 DFF_394_Q_reg ( .D(g24228), .SI(test_si25), .SE(n9326), .CLK(n9513), 
        .Q(g471) );
  SDFFX1 DFF_395_Q_reg ( .D(n540), .SI(g471), .SE(n9328), .CLK(n9515), .Q(g528) );
  SDFFX1 DFF_396_Q_reg ( .D(g528), .SI(g528), .SE(n9328), .CLK(n9515), .Q(g535) );
  SDFFX1 DFF_397_Q_reg ( .D(g535), .SI(g535), .SE(n9328), .CLK(n9515), .Q(g542) );
  SDFFX1 DFF_398_Q_reg ( .D(g13149), .SI(g542), .SE(n9328), .CLK(n9515), .Q(
        g543) );
  SDFFX1 DFF_399_Q_reg ( .D(g543), .SI(g543), .SE(n9328), .CLK(n9515), .Q(g544) );
  SDFFX1 DFF_400_Q_reg ( .D(g21851), .SI(g544), .SE(n9328), .CLK(n9515), .Q(
        g548), .QN(n8375) );
  SDFFX1 DFF_401_Q_reg ( .D(g13111), .SI(g548), .SE(n9328), .CLK(n9515), .Q(
        g549) );
  SDFFX1 DFF_402_Q_reg ( .D(g549), .SI(g549), .SE(n9328), .CLK(n9515), .Q(g499), .QN(n4541) );
  SDFFX1 DFF_403_Q_reg ( .D(g13160), .SI(g499), .SE(n9328), .CLK(n9515), .Q(
        g558) );
  SDFFX1 DFF_404_Q_reg ( .D(g558), .SI(g558), .SE(n9328), .CLK(n9515), .Q(g559) );
  SDFFX1 DFF_405_Q_reg ( .D(g27261), .SI(g559), .SE(n9358), .CLK(n9545), .Q(
        g576) );
  SDFFX1 DFF_406_Q_reg ( .D(g27268), .SI(g576), .SE(n9358), .CLK(n9545), .Q(
        g577), .QN(n8575) );
  SDFFX1 DFF_407_Q_reg ( .D(g27279), .SI(g577), .SE(n9358), .CLK(n9545), .Q(
        g575) );
  SDFFX1 DFF_408_Q_reg ( .D(g27269), .SI(g575), .SE(n9358), .CLK(n9545), .Q(
        g579) );
  SDFFX1 DFF_409_Q_reg ( .D(g27280), .SI(g579), .SE(n9358), .CLK(n9545), .Q(
        test_so25) );
  SDFFX1 DFF_410_Q_reg ( .D(g27294), .SI(test_si26), .SE(n9358), .CLK(n9545), 
        .Q(g578) );
  SDFFX1 DFF_411_Q_reg ( .D(g27281), .SI(g578), .SE(n9358), .CLK(n9545), .Q(
        g582) );
  SDFFX1 DFF_412_Q_reg ( .D(g27295), .SI(g582), .SE(n9358), .CLK(n9545), .Q(
        g583), .QN(n8401) );
  SDFFX1 DFF_413_Q_reg ( .D(g27311), .SI(g583), .SE(n9357), .CLK(n9544), .Q(
        g581) );
  SDFFX1 DFF_414_Q_reg ( .D(g27296), .SI(g581), .SE(n9357), .CLK(n9544), .Q(
        g585) );
  SDFFX1 DFF_415_Q_reg ( .D(g27312), .SI(g585), .SE(n9358), .CLK(n9545), .Q(
        g586), .QN(n8609) );
  SDFFX1 DFF_416_Q_reg ( .D(g27327), .SI(g586), .SE(n9358), .CLK(n9545), .Q(
        g584) );
  SDFFX1 DFF_417_Q_reg ( .D(g24491), .SI(g584), .SE(n9358), .CLK(n9545), .Q(
        g587), .QN(n8669) );
  SDFFX1 DFF_418_Q_reg ( .D(g24498), .SI(g587), .SE(n9358), .CLK(n9545), .Q(
        g590), .QN(n8671) );
  SDFFX1 DFF_419_Q_reg ( .D(g24507), .SI(g590), .SE(n9359), .CLK(n9546), .Q(
        g593), .QN(n8670) );
  SDFFX1 DFF_420_Q_reg ( .D(g24499), .SI(g593), .SE(n9359), .CLK(n9546), .Q(
        g596), .QN(n8657) );
  SDFFX1 DFF_421_Q_reg ( .D(g24508), .SI(g596), .SE(n9359), .CLK(n9546), .Q(
        g599), .QN(n8659) );
  SDFFX1 DFF_422_Q_reg ( .D(g24519), .SI(g599), .SE(n9359), .CLK(n9546), .Q(
        g602), .QN(n8658) );
  SDFFX1 DFF_423_Q_reg ( .D(g28345), .SI(g602), .SE(n9359), .CLK(n9546), .Q(
        g614), .QN(n8673) );
  SDFFX1 DFF_424_Q_reg ( .D(g28349), .SI(g614), .SE(n9359), .CLK(n9546), .Q(
        g617) );
  SDFFX1 DFF_425_Q_reg ( .D(g28353), .SI(g617), .SE(n9359), .CLK(n9546), .Q(
        test_so26) );
  SDFFX1 DFF_426_Q_reg ( .D(g28342), .SI(test_si27), .SE(n9359), .CLK(n9546), 
        .Q(g605), .QN(n8675) );
  SDFFX1 DFF_427_Q_reg ( .D(g28344), .SI(g605), .SE(n9359), .CLK(n9546), .Q(
        g608) );
  SDFFX1 DFF_428_Q_reg ( .D(g28348), .SI(g608), .SE(n9359), .CLK(n9546), .Q(
        g611), .QN(n8676) );
  SDFFX1 DFF_429_Q_reg ( .D(g26541), .SI(g611), .SE(n9360), .CLK(n9547), .Q(
        g490), .QN(n8746) );
  SDFFX1 DFF_430_Q_reg ( .D(g26545), .SI(g490), .SE(n9360), .CLK(n9547), .Q(
        g493) );
  SDFFX1 DFF_431_Q_reg ( .D(g26553), .SI(g493), .SE(n9360), .CLK(n9547), .Q(
        g496), .QN(n8750) );
  SDFFX1 DFF_432_Q_reg ( .D(g499), .SI(g496), .SE(n9360), .CLK(n9547), .Q(g506), .QN(n4570) );
  SDFFX1 DFF_433_Q_reg ( .D(g22578), .SI(g506), .SE(n9360), .CLK(n9547), .Q(
        n4571), .QN(n8672) );
  SDFFX1 DFF_442_Q_reg ( .D(n550), .SI(n4571), .SE(n9360), .CLK(n9547), .Q(
        g16297) );
  SDFFX1 DFF_443_Q_reg ( .D(g16297), .SI(g16297), .SE(n9361), .CLK(n9548), .Q(
        g525), .QN(n8995) );
  SDFFX1 DFF_444_Q_reg ( .D(DFF_299_n1), .SI(g525), .SE(n9361), .CLK(n9548), 
        .Q(n8047) );
  SDFFX1 DFF_445_Q_reg ( .D(DFF_301_n1), .SI(n8047), .SE(n9361), .CLK(n9548), 
        .Q(n8046), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(DFF_303_n1), .SI(n8046), .SE(n9361), .CLK(n9548), 
        .Q(n8045), .QN(DFF_446_n1) );
  SDFFX1 DFF_447_Q_reg ( .D(DFF_305_n1), .SI(n8045), .SE(n9361), .CLK(n9548), 
        .Q(n8044) );
  SDFFX1 DFF_448_Q_reg ( .D(DFF_307_n1), .SI(n8044), .SE(n9361), .CLK(n9548), 
        .Q(n8043) );
  SDFFX1 DFF_449_Q_reg ( .D(DFF_309_n1), .SI(n8043), .SE(n9361), .CLK(n9548), 
        .Q(test_so27) );
  SDFFX1 DFF_450_Q_reg ( .D(DFF_311_n1), .SI(test_si28), .SE(n9307), .CLK(
        n9494), .Q(g536) );
  SDFFX1 DFF_451_Q_reg ( .D(DFF_313_n1), .SI(g536), .SE(n9308), .CLK(n9495), 
        .Q(g537) );
  SDFFX1 DFF_452_Q_reg ( .D(g24059), .SI(g537), .SE(n9297), .CLK(n9484), .Q(
        g538), .QN(n4492) );
  SDFFX1 DFF_453_Q_reg ( .D(n4485), .SI(g538), .SE(n9307), .CLK(n9494), .Q(
        n8040), .QN(n16816) );
  SDFFX1 DFF_455_Q_reg ( .D(g6677), .SI(g6677), .SE(n9324), .CLK(n9511), .Q(
        g6911), .QN(n4359) );
  SDFFX1 DFF_456_Q_reg ( .D(g6911), .SI(g6911), .SE(n9324), .CLK(n9511), .Q(
        g629), .QN(n4295) );
  SDFFX1 DFF_457_Q_reg ( .D(g16654), .SI(g629), .SE(n9325), .CLK(n9512), .Q(
        g630), .QN(n9034) );
  SDFFX1 DFF_458_Q_reg ( .D(g20314), .SI(g630), .SE(n9330), .CLK(n9517), .Q(
        g659) );
  SDFFX1 DFF_459_Q_reg ( .D(g20682), .SI(g659), .SE(n9330), .CLK(n9517), .Q(
        g640), .QN(n4404) );
  SDFFX1 DFF_460_Q_reg ( .D(g23136), .SI(g640), .SE(n9330), .CLK(n9517), .Q(
        g633), .QN(n4478) );
  SDFFX1 DFF_461_Q_reg ( .D(g23324), .SI(g633), .SE(n9330), .CLK(n9517), .Q(
        g653), .QN(n4422) );
  SDFFX1 DFF_462_Q_reg ( .D(g24426), .SI(g653), .SE(n9330), .CLK(n9517), .Q(
        g646), .QN(n4414) );
  SDFFX1 DFF_463_Q_reg ( .D(g25185), .SI(g646), .SE(n9330), .CLK(n9517), .Q(
        g660), .QN(n4403) );
  SDFFX1 DFF_464_Q_reg ( .D(g26660), .SI(g660), .SE(n9331), .CLK(n9518), .Q(
        g672), .QN(n4413) );
  SDFFX1 DFF_465_Q_reg ( .D(g26776), .SI(g672), .SE(n9331), .CLK(n9518), .Q(
        test_so28), .QN(n9283) );
  SDFFX1 DFF_466_Q_reg ( .D(g27672), .SI(test_si29), .SE(n9331), .CLK(n9518), 
        .Q(g679), .QN(n4477) );
  SDFFX1 DFF_467_Q_reg ( .D(n614), .SI(g679), .SE(n9331), .CLK(n9518), .Q(g686), .QN(n4396) );
  SDFFX1 DFF_468_Q_reg ( .D(g28668), .SI(g686), .SE(n9331), .CLK(n9518), .Q(
        g692), .QN(n4418) );
  SDFFX1 DFF_469_Q_reg ( .D(g20875), .SI(g692), .SE(n9331), .CLK(n9518), .Q(
        g699) );
  SDFFX1 DFF_470_Q_reg ( .D(g20879), .SI(g699), .SE(n9331), .CLK(n9518), .Q(
        g700), .QN(n9112) );
  SDFFX1 DFF_471_Q_reg ( .D(g20891), .SI(g700), .SE(n9331), .CLK(n9518), .Q(
        g698) );
  SDFFX1 DFF_472_Q_reg ( .D(g20880), .SI(g698), .SE(n9331), .CLK(n9518), .Q(
        g702) );
  SDFFX1 DFF_473_Q_reg ( .D(g20892), .SI(g702), .SE(n9331), .CLK(n9518), .Q(
        g703), .QN(n9110) );
  SDFFX1 DFF_474_Q_reg ( .D(g20901), .SI(g703), .SE(n9332), .CLK(n9519), .Q(
        g701) );
  SDFFX1 DFF_475_Q_reg ( .D(g20893), .SI(g701), .SE(n9332), .CLK(n9519), .Q(
        g705) );
  SDFFX1 DFF_476_Q_reg ( .D(g20902), .SI(g705), .SE(n9332), .CLK(n9519), .Q(
        g706), .QN(n9108) );
  SDFFX1 DFF_477_Q_reg ( .D(g20921), .SI(g706), .SE(n9332), .CLK(n9519), .Q(
        g704) );
  SDFFX1 DFF_478_Q_reg ( .D(g20903), .SI(g704), .SE(n9332), .CLK(n9519), .Q(
        g708) );
  SDFFX1 DFF_479_Q_reg ( .D(g20922), .SI(g708), .SE(n9332), .CLK(n9519), .Q(
        g709), .QN(n9106) );
  SDFFX1 DFF_480_Q_reg ( .D(g20944), .SI(g709), .SE(n9332), .CLK(n9519), .Q(
        g707) );
  SDFFX1 DFF_481_Q_reg ( .D(g20923), .SI(g707), .SE(n9332), .CLK(n9519), .Q(
        test_so29) );
  SDFFX1 DFF_482_Q_reg ( .D(g20945), .SI(test_si30), .SE(n9332), .CLK(n9519), 
        .Q(g712), .QN(n9105) );
  SDFFX1 DFF_483_Q_reg ( .D(g20966), .SI(g712), .SE(n9332), .CLK(n9519), .Q(
        g710) );
  SDFFX1 DFF_484_Q_reg ( .D(g20946), .SI(g710), .SE(n9332), .CLK(n9519), .Q(
        g714) );
  SDFFX1 DFF_485_Q_reg ( .D(g20967), .SI(g714), .SE(n9332), .CLK(n9519), .Q(
        g715), .QN(n9103) );
  SDFFX1 DFF_486_Q_reg ( .D(g20989), .SI(g715), .SE(n9333), .CLK(n9520), .Q(
        g713) );
  SDFFX1 DFF_487_Q_reg ( .D(g20968), .SI(g713), .SE(n9333), .CLK(n9520), .Q(
        g717) );
  SDFFX1 DFF_488_Q_reg ( .D(g20990), .SI(g717), .SE(n9333), .CLK(n9520), .Q(
        g718), .QN(n9101) );
  SDFFX1 DFF_489_Q_reg ( .D(g21009), .SI(g718), .SE(n9333), .CLK(n9520), .Q(
        g716) );
  SDFFX1 DFF_490_Q_reg ( .D(g20991), .SI(g716), .SE(n9333), .CLK(n9520), .Q(
        g720) );
  SDFFX1 DFF_491_Q_reg ( .D(g21010), .SI(g720), .SE(n9333), .CLK(n9520), .Q(
        g721), .QN(n9099) );
  SDFFX1 DFF_492_Q_reg ( .D(g21031), .SI(g721), .SE(n9333), .CLK(n9520), .Q(
        g719) );
  SDFFX1 DFF_493_Q_reg ( .D(g21011), .SI(g719), .SE(n9333), .CLK(n9520), .Q(
        g723) );
  SDFFX1 DFF_494_Q_reg ( .D(g21032), .SI(g723), .SE(n9333), .CLK(n9520), .Q(
        g724), .QN(n9097) );
  SDFFX1 DFF_495_Q_reg ( .D(g21051), .SI(g724), .SE(n9333), .CLK(n9520), .Q(
        g722) );
  SDFFX1 DFF_496_Q_reg ( .D(g20876), .SI(g722), .SE(n9333), .CLK(n9520), .Q(
        g726) );
  SDFFX1 DFF_497_Q_reg ( .D(g20881), .SI(g726), .SE(n9353), .CLK(n9540), .Q(
        test_so30), .QN(n9292) );
  SDFFX1 DFF_498_Q_reg ( .D(g20894), .SI(test_si31), .SE(n9331), .CLK(n9518), 
        .Q(g725) );
  SDFFX1 DFF_499_Q_reg ( .D(g20924), .SI(g725), .SE(n9359), .CLK(n9546), .Q(
        g729) );
  SDFFX1 DFF_500_Q_reg ( .D(g20947), .SI(g729), .SE(n9359), .CLK(n9546), .Q(
        g730) );
  SDFFX1 DFF_501_Q_reg ( .D(g20969), .SI(g730), .SE(n9360), .CLK(n9547), .Q(
        g728), .QN(n8901) );
  SDFFX1 DFF_502_Q_reg ( .D(g20948), .SI(g728), .SE(n9360), .CLK(n9547), .Q(
        g732) );
  SDFFX1 DFF_503_Q_reg ( .D(g20970), .SI(g732), .SE(n9360), .CLK(n9547), .Q(
        g733), .QN(n8843) );
  SDFFX1 DFF_504_Q_reg ( .D(g20992), .SI(g733), .SE(n9360), .CLK(n9547), .Q(
        g731) );
  SDFFX1 DFF_505_Q_reg ( .D(g25260), .SI(g731), .SE(n9360), .CLK(n9547), .Q(
        g735) );
  SDFFX1 DFF_506_Q_reg ( .D(g25262), .SI(g735), .SE(n9360), .CLK(n9547), .Q(
        g736) );
  SDFFX1 DFF_507_Q_reg ( .D(g25266), .SI(g736), .SE(n9297), .CLK(n9484), .Q(
        g734) );
  SDFFX1 DFF_508_Q_reg ( .D(n589), .SI(g734), .SE(n9331), .CLK(n9518), .Q(g738), .QN(n9155) );
  SDFFX1 DFF_509_Q_reg ( .D(g22231), .SI(g738), .SE(n9333), .CLK(n9520), .Q(
        g739) );
  SDFFX1 DFF_510_Q_reg ( .D(g22242), .SI(g739), .SE(n9334), .CLK(n9521), .Q(
        g737), .QN(n9222) );
  SDFFX1 DFF_511_Q_reg ( .D(g2950), .SI(g737), .SE(n9334), .CLK(n9521), .Q(
        g6368), .QN(n4323) );
  SDFFX1 DFF_512_Q_reg ( .D(g6368), .SI(g6368), .SE(n9334), .CLK(n9521), .Q(
        g6518), .QN(n4312) );
  SDFFX1 DFF_513_Q_reg ( .D(g6518), .SI(g6518), .SE(n9334), .CLK(n9521), .Q(
        test_so31), .QN(n9279) );
  SDFFX1 DFF_514_Q_reg ( .D(g22126), .SI(test_si32), .SE(n9335), .CLK(n9522), 
        .Q(g818) );
  SDFFX1 DFF_515_Q_reg ( .D(g22145), .SI(g818), .SE(n9338), .CLK(n9525), .Q(
        g819) );
  SDFFX1 DFF_516_Q_reg ( .D(g22162), .SI(g819), .SE(n9338), .CLK(n9525), .Q(
        g817), .QN(n8827) );
  SDFFX1 DFF_517_Q_reg ( .D(g22146), .SI(g817), .SE(n9335), .CLK(n9522), .Q(
        g821) );
  SDFFX1 DFF_518_Q_reg ( .D(g22163), .SI(g821), .SE(n9338), .CLK(n9525), .Q(
        g822) );
  SDFFX1 DFF_519_Q_reg ( .D(g22177), .SI(g822), .SE(n9338), .CLK(n9525), .Q(
        g820), .QN(n8826) );
  SDFFX1 DFF_520_Q_reg ( .D(g22029), .SI(g820), .SE(n9338), .CLK(n9525), .Q(
        g830) );
  SDFFX1 DFF_521_Q_reg ( .D(g22033), .SI(g830), .SE(n9338), .CLK(n9525), .Q(
        g831) );
  SDFFX1 DFF_522_Q_reg ( .D(g22040), .SI(g831), .SE(n9338), .CLK(n9525), .Q(
        g829), .QN(n8825) );
  SDFFX1 DFF_523_Q_reg ( .D(g22034), .SI(g829), .SE(n9339), .CLK(n9526), .Q(
        g833) );
  SDFFX1 DFF_524_Q_reg ( .D(g22041), .SI(g833), .SE(n9339), .CLK(n9526), .Q(
        g834) );
  SDFFX1 DFF_525_Q_reg ( .D(g22054), .SI(g834), .SE(n9339), .CLK(n9526), .Q(
        g832), .QN(n8824) );
  SDFFX1 DFF_526_Q_reg ( .D(g22042), .SI(g832), .SE(n9339), .CLK(n9526), .Q(
        g836) );
  SDFFX1 DFF_527_Q_reg ( .D(g22055), .SI(g836), .SE(n9339), .CLK(n9526), .Q(
        g837) );
  SDFFX1 DFF_528_Q_reg ( .D(g22066), .SI(g837), .SE(n9339), .CLK(n9526), .Q(
        g835), .QN(n8823) );
  SDFFX1 DFF_529_Q_reg ( .D(g22056), .SI(g835), .SE(n9339), .CLK(n9526), .Q(
        test_so32) );
  SDFFX1 DFF_530_Q_reg ( .D(g22067), .SI(test_si33), .SE(n9337), .CLK(n9524), 
        .Q(g840) );
  SDFFX1 DFF_531_Q_reg ( .D(g22087), .SI(g840), .SE(n9337), .CLK(n9524), .Q(
        g838), .QN(n8822) );
  SDFFX1 DFF_532_Q_reg ( .D(g22068), .SI(g838), .SE(n9337), .CLK(n9524), .Q(
        g842) );
  SDFFX1 DFF_533_Q_reg ( .D(g22088), .SI(g842), .SE(n9337), .CLK(n9524), .Q(
        g843) );
  SDFFX1 DFF_534_Q_reg ( .D(g22104), .SI(g843), .SE(n9337), .CLK(n9524), .Q(
        g841), .QN(n8821) );
  SDFFX1 DFF_535_Q_reg ( .D(g22089), .SI(g841), .SE(n9337), .CLK(n9524), .Q(
        g845) );
  SDFFX1 DFF_536_Q_reg ( .D(g22105), .SI(g845), .SE(n9337), .CLK(n9524), .Q(
        g846) );
  SDFFX1 DFF_537_Q_reg ( .D(g22127), .SI(g846), .SE(n9337), .CLK(n9524), .Q(
        g844), .QN(n8820) );
  SDFFX1 DFF_538_Q_reg ( .D(g22106), .SI(g844), .SE(n9337), .CLK(n9524), .Q(
        g848) );
  SDFFX1 DFF_539_Q_reg ( .D(g22128), .SI(g848), .SE(n9337), .CLK(n9524), .Q(
        g849) );
  SDFFX1 DFF_540_Q_reg ( .D(g22147), .SI(g849), .SE(n9337), .CLK(n9524), .Q(
        g847), .QN(n8817) );
  SDFFX1 DFF_541_Q_reg ( .D(g22129), .SI(g847), .SE(n9338), .CLK(n9525), .Q(
        g851), .QN(n8816) );
  SDFFX1 DFF_542_Q_reg ( .D(g22148), .SI(g851), .SE(n9338), .CLK(n9525), .Q(
        g852), .QN(n8815) );
  SDFFX1 DFF_543_Q_reg ( .D(g22164), .SI(g852), .SE(n9338), .CLK(n9525), .Q(
        g850) );
  SDFFX1 DFF_544_Q_reg ( .D(g25209), .SI(g850), .SE(n9338), .CLK(n9525), .Q(
        g857) );
  SDFFX1 DFF_545_Q_reg ( .D(g25214), .SI(g857), .SE(n9338), .CLK(n9525), .Q(
        test_so33) );
  SDFFX1 DFF_546_Q_reg ( .D(g25221), .SI(test_si34), .SE(n9334), .CLK(n9521), 
        .Q(g856), .QN(n8881) );
  SDFFX1 DFF_547_Q_reg ( .D(g25215), .SI(g856), .SE(n9334), .CLK(n9521), .Q(
        g860) );
  SDFFX1 DFF_548_Q_reg ( .D(g25222), .SI(g860), .SE(n9334), .CLK(n9521), .Q(
        g861) );
  SDFFX1 DFF_549_Q_reg ( .D(g25230), .SI(g861), .SE(n9334), .CLK(n9521), .Q(
        g859), .QN(n8878) );
  SDFFX1 DFF_550_Q_reg ( .D(g25223), .SI(g859), .SE(n9334), .CLK(n9521), .Q(
        g863) );
  SDFFX1 DFF_551_Q_reg ( .D(g25231), .SI(g863), .SE(n9334), .CLK(n9521), .Q(
        g864) );
  SDFFX1 DFF_552_Q_reg ( .D(g25240), .SI(g864), .SE(n9334), .CLK(n9521), .Q(
        g862), .QN(n8875) );
  SDFFX1 DFF_553_Q_reg ( .D(g25232), .SI(g862), .SE(n9334), .CLK(n9521), .Q(
        g866) );
  SDFFX1 DFF_554_Q_reg ( .D(g25241), .SI(g866), .SE(n9335), .CLK(n9522), .Q(
        g867) );
  SDFFX1 DFF_555_Q_reg ( .D(g25248), .SI(g867), .SE(n9335), .CLK(n9522), .Q(
        g865), .QN(n8872) );
  SDFFX1 DFF_556_Q_reg ( .D(g30269), .SI(g865), .SE(n9340), .CLK(n9527), .Q(
        g873), .QN(n8469) );
  SDFFX1 DFF_557_Q_reg ( .D(g30277), .SI(g873), .SE(n9340), .CLK(n9527), .Q(
        g876), .QN(n8468) );
  SDFFX1 DFF_558_Q_reg ( .D(g30285), .SI(g876), .SE(n9340), .CLK(n9527), .Q(
        g879) );
  SDFFX1 DFF_559_Q_reg ( .D(g30643), .SI(g879), .SE(n9340), .CLK(n9527), .Q(
        g918), .QN(n8467) );
  SDFFX1 DFF_560_Q_reg ( .D(g30648), .SI(g918), .SE(n9340), .CLK(n9527), .Q(
        g921), .QN(n8488) );
  SDFFX1 DFF_561_Q_reg ( .D(g30654), .SI(g921), .SE(n9340), .CLK(n9527), .Q(
        test_so34) );
  SDFFX1 DFF_562_Q_reg ( .D(g30676), .SI(test_si35), .SE(n9335), .CLK(n9522), 
        .Q(g882), .QN(n8466) );
  SDFFX1 DFF_563_Q_reg ( .D(g30681), .SI(g882), .SE(n9335), .CLK(n9522), .Q(
        g885), .QN(n8465) );
  SDFFX1 DFF_564_Q_reg ( .D(g30687), .SI(g885), .SE(n9335), .CLK(n9522), .Q(
        g888) );
  SDFFX1 DFF_565_Q_reg ( .D(g30649), .SI(g888), .SE(n9340), .CLK(n9527), .Q(
        g927), .QN(n8464) );
  SDFFX1 DFF_566_Q_reg ( .D(g30655), .SI(g927), .SE(n9341), .CLK(n9528), .Q(
        g930), .QN(n8487) );
  SDFFX1 DFF_567_Q_reg ( .D(g30662), .SI(g930), .SE(n9341), .CLK(n9528), .Q(
        g933) );
  SDFFX1 DFF_568_Q_reg ( .D(g30286), .SI(g933), .SE(n9341), .CLK(n9528), .Q(
        g891), .QN(n8463) );
  SDFFX1 DFF_569_Q_reg ( .D(g30293), .SI(g891), .SE(n9341), .CLK(n9528), .Q(
        g894), .QN(n8462) );
  SDFFX1 DFF_570_Q_reg ( .D(g30298), .SI(g894), .SE(n9341), .CLK(n9528), .Q(
        g897) );
  SDFFX1 DFF_571_Q_reg ( .D(g30259), .SI(g897), .SE(n9341), .CLK(n9528), .Q(
        g936), .QN(n8461) );
  SDFFX1 DFF_572_Q_reg ( .D(g30264), .SI(g936), .SE(n9341), .CLK(n9528), .Q(
        g939), .QN(n8460) );
  SDFFX1 DFF_573_Q_reg ( .D(g30270), .SI(g939), .SE(n9341), .CLK(n9528), .Q(
        g942) );
  SDFFX1 DFF_574_Q_reg ( .D(g30247), .SI(g942), .SE(n9341), .CLK(n9528), .Q(
        g900), .QN(n8459) );
  SDFFX1 DFF_575_Q_reg ( .D(g30249), .SI(g900), .SE(n9341), .CLK(n9528), .Q(
        g903), .QN(n8458) );
  SDFFX1 DFF_576_Q_reg ( .D(g30251), .SI(g903), .SE(n9341), .CLK(n9528), .Q(
        g906) );
  SDFFX1 DFF_577_Q_reg ( .D(g30265), .SI(g906), .SE(n9341), .CLK(n9528), .Q(
        test_so35) );
  SDFFX1 DFF_578_Q_reg ( .D(g30271), .SI(test_si36), .SE(n9342), .CLK(n9529), 
        .Q(g948), .QN(n8457) );
  SDFFX1 DFF_579_Q_reg ( .D(g30278), .SI(g948), .SE(n9342), .CLK(n9529), .Q(
        g951) );
  SDFFX1 DFF_580_Q_reg ( .D(g30638), .SI(g951), .SE(n9342), .CLK(n9529), .Q(
        g909), .QN(n8456) );
  SDFFX1 DFF_581_Q_reg ( .D(g30642), .SI(g909), .SE(n9342), .CLK(n9529), .Q(
        g912), .QN(n8492) );
  SDFFX1 DFF_582_Q_reg ( .D(g30647), .SI(g912), .SE(n9340), .CLK(n9527), .Q(
        g915) );
  SDFFX1 DFF_583_Q_reg ( .D(g30670), .SI(g915), .SE(n9340), .CLK(n9527), .Q(
        g954), .QN(n8455) );
  SDFFX1 DFF_584_Q_reg ( .D(g30677), .SI(g954), .SE(n9340), .CLK(n9527), .Q(
        g957), .QN(n8491) );
  SDFFX1 DFF_585_Q_reg ( .D(g30682), .SI(g957), .SE(n9335), .CLK(n9522), .Q(
        g960) );
  SDFFX1 DFF_586_Q_reg ( .D(g25042), .SI(g960), .SE(n9335), .CLK(n9522), .Q(
        g780), .QN(n8980) );
  SDFFX1 DFF_587_Q_reg ( .D(g25935), .SI(g780), .SE(n9335), .CLK(n9522), .Q(
        g776), .QN(n9272) );
  SDFFX1 DFF_588_Q_reg ( .D(g26530), .SI(g776), .SE(n9335), .CLK(n9522), .Q(
        g771), .QN(n8979) );
  SDFFX1 DFF_589_Q_reg ( .D(g27123), .SI(g771), .SE(n9335), .CLK(n9522), .Q(
        g767), .QN(n9273) );
  SDFFX1 DFF_590_Q_reg ( .D(g27603), .SI(g767), .SE(n9336), .CLK(n9523), .Q(
        g762), .QN(n8978) );
  SDFFX1 DFF_591_Q_reg ( .D(g28146), .SI(g762), .SE(n9336), .CLK(n9523), .Q(
        g758), .QN(n9274) );
  SDFFX1 DFF_592_Q_reg ( .D(g28635), .SI(g758), .SE(n9336), .CLK(n9523), .Q(
        g753), .QN(n8977) );
  SDFFX1 DFF_593_Q_reg ( .D(g29110), .SI(g753), .SE(n9336), .CLK(n9523), .Q(
        test_so36) );
  SDFFX1 DFF_594_Q_reg ( .D(g29354), .SI(test_si37), .SE(n9336), .CLK(n9523), 
        .Q(g744), .QN(n8561) );
  SDFFX1 DFF_595_Q_reg ( .D(g29580), .SI(g744), .SE(n9336), .CLK(n9523), .Q(
        g740), .QN(n8390) );
  SDFFX1 DFF_596_Q_reg ( .D(n15), .SI(g740), .SE(n9336), .CLK(n9523), .Q(g868)
         );
  SDFFX1 DFF_597_Q_reg ( .D(g868), .SI(g868), .SE(n9336), .CLK(n9523), .Q(
        g5595) );
  SDFFX1 DFF_598_Q_reg ( .D(g5595), .SI(g5595), .SE(n9336), .CLK(n9523), .Q(
        g869), .QN(n8990) );
  SDFFX1 DFF_599_Q_reg ( .D(g2950), .SI(g869), .SE(n9336), .CLK(n9523), .Q(
        g5472), .QN(n4363) );
  SDFFX1 DFF_600_Q_reg ( .D(g5472), .SI(g5472), .SE(n9336), .CLK(n9523), .Q(
        g6712), .QN(n4364) );
  SDFFX1 DFF_601_Q_reg ( .D(g6712), .SI(g6712), .SE(n9336), .CLK(n9523), .Q(
        g1088), .QN(n4381) );
  SDFFX1 DFF_602_Q_reg ( .D(g5595), .SI(g1088), .SE(n9337), .CLK(n9524), .Q(
        g996), .QN(n4387) );
  SDFFX1 DFF_603_Q_reg ( .D(g27257), .SI(g996), .SE(n9345), .CLK(n9532), .Q(
        g1041) );
  SDFFX1 DFF_604_Q_reg ( .D(g27262), .SI(g1041), .SE(n9345), .CLK(n9532), .Q(
        g1030) );
  SDFFX1 DFF_605_Q_reg ( .D(g27270), .SI(g1030), .SE(n9346), .CLK(n9533), .Q(
        g1033), .QN(n8931) );
  SDFFX1 DFF_606_Q_reg ( .D(g27263), .SI(g1033), .SE(n9346), .CLK(n9533), .Q(
        g1056) );
  SDFFX1 DFF_607_Q_reg ( .D(g27271), .SI(g1056), .SE(n9346), .CLK(n9533), .Q(
        g1045) );
  SDFFX1 DFF_608_Q_reg ( .D(g27282), .SI(g1045), .SE(n9345), .CLK(n9532), .Q(
        g1048), .QN(n8908) );
  SDFFX1 DFF_609_Q_reg ( .D(g27272), .SI(g1048), .SE(n9345), .CLK(n9532), .Q(
        test_so37) );
  SDFFX1 DFF_610_Q_reg ( .D(g27283), .SI(test_si38), .SE(n9345), .CLK(n9532), 
        .Q(g1060) );
  SDFFX1 DFF_611_Q_reg ( .D(g27297), .SI(g1060), .SE(n9345), .CLK(n9532), .Q(
        g1063), .QN(n8642) );
  SDFFX1 DFF_612_Q_reg ( .D(g27284), .SI(g1063), .SE(n9346), .CLK(n9533), .Q(
        g1085) );
  SDFFX1 DFF_613_Q_reg ( .D(g27298), .SI(g1085), .SE(n9346), .CLK(n9533), .Q(
        g1075) );
  SDFFX1 DFF_614_Q_reg ( .D(g27313), .SI(g1075), .SE(n9343), .CLK(n9530), .Q(
        g1078), .QN(n8919) );
  SDFFX1 DFF_615_Q_reg ( .D(g28738), .SI(g1078), .SE(n9343), .CLK(n9530), .Q(
        g1095), .QN(n8732) );
  SDFFX1 DFF_616_Q_reg ( .D(g28746), .SI(g1095), .SE(n9345), .CLK(n9532), .Q(
        g1098), .QN(n8710) );
  SDFFX1 DFF_617_Q_reg ( .D(g28758), .SI(g1098), .SE(n9345), .CLK(n9532), .Q(
        g1101) );
  SDFFX1 DFF_618_Q_reg ( .D(g29198), .SI(g1101), .SE(n9345), .CLK(n9532), .Q(
        g1104), .QN(n8730) );
  SDFFX1 DFF_619_Q_reg ( .D(g29204), .SI(g1104), .SE(n9345), .CLK(n9532), .Q(
        g1107), .QN(n8709) );
  SDFFX1 DFF_620_Q_reg ( .D(g29209), .SI(g1107), .SE(n9343), .CLK(n9530), .Q(
        g1110) );
  SDFFX1 DFF_621_Q_reg ( .D(g28747), .SI(g1110), .SE(n9343), .CLK(n9530), .Q(
        g1114) );
  SDFFX1 DFF_622_Q_reg ( .D(g28759), .SI(g1114), .SE(n9344), .CLK(n9531), .Q(
        g1115) );
  SDFFX1 DFF_623_Q_reg ( .D(g28767), .SI(g1115), .SE(n9344), .CLK(n9531), .Q(
        g1113), .QN(n8958) );
  SDFFX1 DFF_624_Q_reg ( .D(g26806), .SI(g1113), .SE(n9344), .CLK(n9531), .Q(
        g1116), .QN(n8728) );
  SDFFX1 DFF_625_Q_reg ( .D(g26809), .SI(g1116), .SE(n9344), .CLK(n9531), .Q(
        test_so38) );
  SDFFX1 DFF_626_Q_reg ( .D(g26813), .SI(test_si39), .SE(n9344), .CLK(n9531), 
        .Q(g1122) );
  SDFFX1 DFF_627_Q_reg ( .D(g26810), .SI(g1122), .SE(n9344), .CLK(n9531), .Q(
        g1125), .QN(n8726) );
  SDFFX1 DFF_628_Q_reg ( .D(g26814), .SI(g1125), .SE(n9344), .CLK(n9531), .Q(
        g1128), .QN(n8708) );
  SDFFX1 DFF_629_Q_reg ( .D(g26818), .SI(g1128), .SE(n9344), .CLK(n9531), .Q(
        g1131) );
  SDFFX1 DFF_630_Q_reg ( .D(g27761), .SI(g1131), .SE(n9345), .CLK(n9532), .Q(
        g1135), .QN(n8957) );
  SDFFX1 DFF_631_Q_reg ( .D(g27763), .SI(g1135), .SE(n9344), .CLK(n9531), .Q(
        g1136), .QN(n8943) );
  SDFFX1 DFF_632_Q_reg ( .D(g27765), .SI(g1136), .SE(n9344), .CLK(n9531), .Q(
        g1134), .QN(n8956) );
  SDFFX1 DFF_633_Q_reg ( .D(g29609), .SI(g1134), .SE(n9344), .CLK(n9531), .Q(
        g999) );
  SDFFX1 DFF_634_Q_reg ( .D(g29612), .SI(g999), .SE(n9344), .CLK(n9531), .Q(
        g1000) );
  SDFFX1 DFF_635_Q_reg ( .D(g29616), .SI(g1000), .SE(n9340), .CLK(n9527), .Q(
        g1001), .QN(n8517) );
  SDFFX1 DFF_636_Q_reg ( .D(g30701), .SI(g1001), .SE(n9339), .CLK(n9526), .Q(
        g1002) );
  SDFFX1 DFF_637_Q_reg ( .D(g30703), .SI(g1002), .SE(n9339), .CLK(n9526), .Q(
        g1003) );
  SDFFX1 DFF_638_Q_reg ( .D(g30705), .SI(g1003), .SE(n9339), .CLK(n9526), .Q(
        g1004), .QN(n8515) );
  SDFFX1 DFF_639_Q_reg ( .D(g30470), .SI(g1004), .SE(n9339), .CLK(n9526), .Q(
        g1005) );
  SDFFX1 DFF_640_Q_reg ( .D(g30485), .SI(g1005), .SE(n9339), .CLK(n9526), .Q(
        g1006) );
  SDFFX1 DFF_641_Q_reg ( .D(g30500), .SI(g1006), .SE(n9340), .CLK(n9527), .Q(
        test_so39) );
  SDFFX1 DFF_642_Q_reg ( .D(g29170), .SI(test_si40), .SE(n9342), .CLK(n9529), 
        .Q(g1009) );
  SDFFX1 DFF_643_Q_reg ( .D(g29173), .SI(g1009), .SE(n9342), .CLK(n9529), .Q(
        g1010) );
  SDFFX1 DFF_644_Q_reg ( .D(g29179), .SI(g1010), .SE(n9342), .CLK(n9529), .Q(
        g1008), .QN(n8554) );
  SDFFX1 DFF_645_Q_reg ( .D(g26661), .SI(g1008), .SE(n9342), .CLK(n9529), .Q(
        g1090) );
  SDFFX1 DFF_646_Q_reg ( .D(g26665), .SI(g1090), .SE(n9342), .CLK(n9529), .Q(
        g1091) );
  SDFFX1 DFF_647_Q_reg ( .D(g26669), .SI(g1091), .SE(n9342), .CLK(n9529), .Q(
        g1089), .QN(n8954) );
  SDFFX1 DFF_648_Q_reg ( .D(n4289), .SI(g1089), .SE(n9342), .CLK(n9529), .Q(
        g1137) );
  SDFFX1 DFF_649_Q_reg ( .D(g1137), .SI(g1137), .SE(n9342), .CLK(n9529), .Q(
        n8027), .QN(DFF_649_n1) );
  SDFFX1 DFF_650_Q_reg ( .D(n4567), .SI(n8027), .SE(n9343), .CLK(n9530), .Q(
        g1139) );
  SDFFX1 DFF_651_Q_reg ( .D(g1139), .SI(g1139), .SE(n9343), .CLK(n9530), .Q(
        n8026), .QN(DFF_651_n1) );
  SDFFX1 DFF_652_Q_reg ( .D(n4559), .SI(n8026), .SE(n9343), .CLK(n9530), .Q(
        g1141) );
  SDFFX1 DFF_653_Q_reg ( .D(g1141), .SI(g1141), .SE(n9343), .CLK(n9530), .Q(
        n8025), .QN(DFF_653_n1) );
  SDFFX1 DFF_654_Q_reg ( .D(n4327), .SI(n8025), .SE(n9343), .CLK(n9530), .Q(
        g967) );
  SDFFX1 DFF_655_Q_reg ( .D(g967), .SI(g967), .SE(n9343), .CLK(n9530), .Q(
        n8024), .QN(DFF_655_n1) );
  SDFFX1 DFF_656_Q_reg ( .D(n4391), .SI(n8024), .SE(n9343), .CLK(n9530), .Q(
        g969) );
  SDFFX1 DFF_657_Q_reg ( .D(g969), .SI(g969), .SE(n9343), .CLK(n9530), .Q(
        test_so40), .QN(DFF_657_n1) );
  SDFFX1 DFF_658_Q_reg ( .D(n4321), .SI(test_si41), .SE(n9302), .CLK(n9489), 
        .Q(g971) );
  SDFFX1 DFF_659_Q_reg ( .D(g971), .SI(g971), .SE(n9302), .CLK(n9489), .Q(
        n8021), .QN(DFF_659_n1) );
  SDFFX1 DFF_660_Q_reg ( .D(n4375), .SI(n8021), .SE(n9302), .CLK(n9489), .Q(
        g973) );
  SDFFX1 DFF_661_Q_reg ( .D(g973), .SI(g973), .SE(n9302), .CLK(n9489), .Q(
        n8020), .QN(DFF_661_n1) );
  SDFFX1 DFF_662_Q_reg ( .D(n4379), .SI(n8020), .SE(n9302), .CLK(n9489), .Q(
        g975) );
  SDFFX1 DFF_663_Q_reg ( .D(g975), .SI(g975), .SE(n9302), .CLK(n9489), .Q(
        n8019), .QN(DFF_663_n1) );
  SDFFX1 DFF_664_Q_reg ( .D(g2873), .SI(n8019), .SE(n9303), .CLK(n9490), .Q(
        g977) );
  SDFFX1 DFF_665_Q_reg ( .D(g977), .SI(g977), .SE(n9303), .CLK(n9490), .Q(
        n8018), .QN(n4486) );
  SDFFX1 DFF_666_Q_reg ( .D(n4283), .SI(n8018), .SE(n9345), .CLK(n9532), .Q(
        g986), .QN(n4432) );
  SDFFX1 DFF_667_Q_reg ( .D(n477), .SI(g986), .SE(n9346), .CLK(n9533), .Q(g992), .QN(n8987) );
  SDFFX1 DFF_678_Q_reg ( .D(n4277), .SI(g992), .SE(n9346), .CLK(n9533), .Q(
        n8017) );
  SDFFX1 DFF_679_Q_reg ( .D(g1041), .SI(n8017), .SE(n9346), .CLK(n9533), .Q(
        g1029) );
  SDFFX1 DFF_680_Q_reg ( .D(g1029), .SI(g1029), .SE(n9346), .CLK(n9533), .Q(
        g1036) );
  SDFFX1 DFF_681_Q_reg ( .D(g1030), .SI(g1036), .SE(n9346), .CLK(n9533), .Q(
        g1037) );
  SDFFX1 DFF_682_Q_reg ( .D(g1037), .SI(g1037), .SE(n9346), .CLK(n9533), .Q(
        g1038), .QN(n8618) );
  SDFFX1 DFF_683_Q_reg ( .D(g1033), .SI(g1038), .SE(n9346), .CLK(n9533), .Q(
        test_so41) );
  SDFFX1 DFF_684_Q_reg ( .D(test_so41), .SI(test_si42), .SE(n9347), .CLK(n9534), .Q(g1040), .QN(n8617) );
  SDFFX1 DFF_685_Q_reg ( .D(g1056), .SI(g1040), .SE(n9347), .CLK(n9534), .Q(
        g1044) );
  SDFFX1 DFF_686_Q_reg ( .D(g1044), .SI(g1044), .SE(n9347), .CLK(n9534), .Q(
        g1051) );
  SDFFX1 DFF_687_Q_reg ( .D(g1045), .SI(g1051), .SE(n9347), .CLK(n9534), .Q(
        g1052) );
  SDFFX1 DFF_688_Q_reg ( .D(g1052), .SI(g1052), .SE(n9347), .CLK(n9534), .Q(
        g1053), .QN(n8407) );
  SDFFX1 DFF_689_Q_reg ( .D(g1048), .SI(g1053), .SE(n9347), .CLK(n9534), .Q(
        g1054) );
  SDFFX1 DFF_690_Q_reg ( .D(g1054), .SI(g1054), .SE(n9347), .CLK(n9534), .Q(
        g1055), .QN(n8406) );
  SDFFX1 DFF_691_Q_reg ( .D(test_so37), .SI(g1055), .SE(n9347), .CLK(n9534), 
        .Q(g1059) );
  SDFFX1 DFF_692_Q_reg ( .D(g1059), .SI(g1059), .SE(n9347), .CLK(n9534), .Q(
        g1066) );
  SDFFX1 DFF_693_Q_reg ( .D(g1060), .SI(g1066), .SE(n9347), .CLK(n9534), .Q(
        g1067) );
  SDFFX1 DFF_694_Q_reg ( .D(g1067), .SI(g1067), .SE(n9347), .CLK(n9534), .Q(
        g1068), .QN(n8581) );
  SDFFX1 DFF_695_Q_reg ( .D(g1063), .SI(g1068), .SE(n9347), .CLK(n9534), .Q(
        g1069) );
  SDFFX1 DFF_696_Q_reg ( .D(g1069), .SI(g1069), .SE(n9348), .CLK(n9535), .Q(
        g1070), .QN(n8580) );
  SDFFX1 DFF_697_Q_reg ( .D(g1085), .SI(g1070), .SE(n9348), .CLK(n9535), .Q(
        g1074) );
  SDFFX1 DFF_698_Q_reg ( .D(g1074), .SI(g1074), .SE(n9348), .CLK(n9535), .Q(
        g1081), .QN(n16822) );
  SDFFX1 DFF_699_Q_reg ( .D(g1075), .SI(g1081), .SE(n9348), .CLK(n9535), .Q(
        test_so42) );
  SDFFX1 DFF_700_Q_reg ( .D(test_so42), .SI(test_si43), .SE(n9348), .CLK(n9535), .Q(g1083) );
  SDFFX1 DFF_701_Q_reg ( .D(g1078), .SI(g1083), .SE(n9348), .CLK(n9535), .Q(
        g1084) );
  SDFFX1 DFF_702_Q_reg ( .D(g1084), .SI(g1084), .SE(n9348), .CLK(n9535), .Q(
        g1011), .QN(n8627) );
  SDFFX1 DFF_703_Q_reg ( .D(n4598), .SI(g1011), .SE(n9348), .CLK(n9535), .Q(
        g5657), .QN(n8625) );
  SDFFX1 DFF_704_Q_reg ( .D(g5657), .SI(g5657), .SE(n9348), .CLK(n9535), .Q(
        g5686), .QN(n8628) );
  SDFFX1 DFF_705_Q_reg ( .D(g5686), .SI(g5686), .SE(n9348), .CLK(n9535), .Q(
        g1024), .QN(n8626) );
  SDFFX1 DFF_706_Q_reg ( .D(n4598), .SI(g1024), .SE(n9348), .CLK(n9535), .Q(
        g6750), .QN(n4371) );
  SDFFX1 DFF_707_Q_reg ( .D(g6750), .SI(g6750), .SE(n9348), .CLK(n9535), .Q(
        g6944), .QN(n4316) );
  SDFFX1 DFF_708_Q_reg ( .D(g6944), .SI(g6944), .SE(n9349), .CLK(n9536), .Q(
        g1236), .QN(n4300) );
  SDFFX1 DFF_709_Q_reg ( .D(n854), .SI(g1236), .SE(n9349), .CLK(n9536), .Q(
        g1240), .QN(n9225) );
  SDFFX1 DFF_710_Q_reg ( .D(g18707), .SI(g1240), .SE(n9349), .CLK(n9536), .Q(
        g1243), .QN(n4353) );
  SDFFX1 DFF_711_Q_reg ( .D(g18763), .SI(g1243), .SE(n9349), .CLK(n9536), .Q(
        g1196), .QN(n4304) );
  SDFFX1 DFF_712_Q_reg ( .D(n845), .SI(g1196), .SE(n9349), .CLK(n9536), .Q(
        g1199) );
  SDFFX1 DFF_713_Q_reg ( .D(g1199), .SI(g1199), .SE(n9349), .CLK(n9536), .Q(
        g1209) );
  SDFFX1 DFF_714_Q_reg ( .D(g1209), .SI(g1209), .SE(n9349), .CLK(n9536), .Q(
        g1210) );
  SDFFX1 DFF_715_Q_reg ( .D(g1142), .SI(g1210), .SE(n9349), .CLK(n9536), .Q(
        test_so43) );
  SDFFX1 DFF_716_Q_reg ( .D(test_so43), .SI(test_si44), .SE(n9349), .CLK(n9536), .Q(g1255) );
  SDFFX1 DFF_717_Q_reg ( .D(g1145), .SI(g1255), .SE(n9349), .CLK(n9536), .Q(
        g1256) );
  SDFFX1 DFF_718_Q_reg ( .D(g1256), .SI(g1256), .SE(n9349), .CLK(n9536), .Q(
        g1257), .QN(n16827) );
  SDFFX1 DFF_719_Q_reg ( .D(g1148), .SI(g1257), .SE(n9350), .CLK(n9537), .Q(
        g1258) );
  SDFFX1 DFF_720_Q_reg ( .D(g1258), .SI(g1258), .SE(n9350), .CLK(n9537), .Q(
        g1259), .QN(n8779) );
  SDFFX1 DFF_721_Q_reg ( .D(g1152), .SI(g1259), .SE(n9350), .CLK(n9537), .Q(
        g1260) );
  SDFFX1 DFF_722_Q_reg ( .D(g1260), .SI(g1260), .SE(n9350), .CLK(n9537), .Q(
        g1251), .QN(n8776) );
  SDFFX1 DFF_723_Q_reg ( .D(g1155), .SI(g1251), .SE(n9350), .CLK(n9537), .Q(
        g1252) );
  SDFFX1 DFF_724_Q_reg ( .D(g1252), .SI(g1252), .SE(n9350), .CLK(n9537), .Q(
        g1253) );
  SDFFX1 DFF_725_Q_reg ( .D(g1158), .SI(g1253), .SE(n9350), .CLK(n9537), .Q(
        g1254) );
  SDFFX1 DFF_726_Q_reg ( .D(g1254), .SI(g1254), .SE(n9350), .CLK(n9537), .Q(
        g1176), .QN(n8777) );
  SDFFX1 DFF_727_Q_reg ( .D(g2950), .SI(g1176), .SE(n9350), .CLK(n9537), .Q(
        g7961), .QN(n4460) );
  SDFFX1 DFF_728_Q_reg ( .D(g7961), .SI(g7961), .SE(n9350), .CLK(n9537), .Q(
        g8007), .QN(n4459) );
  SDFFX1 DFF_729_Q_reg ( .D(g8007), .SI(g8007), .SE(n9350), .CLK(n9537), .Q(
        g1172), .QN(n4465) );
  SDFFX1 DFF_730_Q_reg ( .D(g23081), .SI(g1172), .SE(n9351), .CLK(n9538), .Q(
        g1173), .QN(n9013) );
  SDFFX1 DFF_731_Q_reg ( .D(g23111), .SI(g1173), .SE(n9351), .CLK(n9538), .Q(
        test_so44) );
  SDFFX1 DFF_732_Q_reg ( .D(g23126), .SI(test_si45), .SE(n9350), .CLK(n9537), 
        .Q(g1175) );
  SDFFX1 DFF_733_Q_reg ( .D(g23392), .SI(g1175), .SE(n9351), .CLK(n9538), .Q(
        g1142) );
  SDFFX1 DFF_734_Q_reg ( .D(g23406), .SI(g1142), .SE(n9351), .CLK(n9538), .Q(
        g1145) );
  SDFFX1 DFF_735_Q_reg ( .D(g24179), .SI(g1145), .SE(n9351), .CLK(n9538), .Q(
        g1148) );
  SDFFX1 DFF_736_Q_reg ( .D(g24181), .SI(g1148), .SE(n9351), .CLK(n9538), .Q(
        g1164), .QN(n9018) );
  SDFFX1 DFF_737_Q_reg ( .D(g24213), .SI(g1164), .SE(n9351), .CLK(n9538), .Q(
        g1165) );
  SDFFX1 DFF_738_Q_reg ( .D(g24223), .SI(g1165), .SE(n9351), .CLK(n9538), .Q(
        g1166), .QN(n9019) );
  SDFFX1 DFF_739_Q_reg ( .D(g23110), .SI(g1166), .SE(n9351), .CLK(n9538), .Q(
        g1167), .QN(n9015) );
  SDFFX1 DFF_740_Q_reg ( .D(g23014), .SI(g1167), .SE(n9351), .CLK(n9538), .Q(
        g1171) );
  SDFFX1 DFF_741_Q_reg ( .D(g23039), .SI(g1171), .SE(n9351), .CLK(n9538), .Q(
        g1151), .QN(n9016) );
  SDFFX1 DFF_742_Q_reg ( .D(g24212), .SI(g1151), .SE(n9352), .CLK(n9539), .Q(
        g1152) );
  SDFFX1 DFF_743_Q_reg ( .D(g24222), .SI(g1152), .SE(n9352), .CLK(n9539), .Q(
        g1155) );
  SDFFX1 DFF_744_Q_reg ( .D(g24235), .SI(g1155), .SE(n9352), .CLK(n9539), .Q(
        g1158) );
  SDFFX1 DFF_745_Q_reg ( .D(n846), .SI(g1158), .SE(n9352), .CLK(n9539), .Q(
        g1214) );
  SDFFX1 DFF_746_Q_reg ( .D(g1214), .SI(g1214), .SE(n9352), .CLK(n9539), .Q(
        g1221) );
  SDFFX1 DFF_747_Q_reg ( .D(g1221), .SI(g1221), .SE(n9352), .CLK(n9539), .Q(
        test_so45), .QN(n8654) );
  SDFFX1 DFF_748_Q_reg ( .D(g13155), .SI(test_si46), .SE(n9351), .CLK(n9538), 
        .Q(g1229) );
  SDFFX1 DFF_749_Q_reg ( .D(g1229), .SI(g1229), .SE(n9352), .CLK(n9539), .Q(
        n4549), .QN(n8373) );
  SDFFX1 DFF_750_Q_reg ( .D(n521), .SI(n4549), .SE(n9352), .CLK(n9539), .Q(
        n4361), .QN(n8374) );
  SDFFX1 DFF_751_Q_reg ( .D(g13124), .SI(n4361), .SE(n9352), .CLK(n9539), .Q(
        g1235) );
  SDFFX1 DFF_752_Q_reg ( .D(g1235), .SI(g1235), .SE(n9352), .CLK(n9539), .Q(
        g1186), .QN(n4548) );
  SDFFX1 DFF_753_Q_reg ( .D(g13171), .SI(g1186), .SE(n9352), .CLK(n9539), .Q(
        g1244) );
  SDFFX1 DFF_754_Q_reg ( .D(g1244), .SI(g1244), .SE(n9352), .CLK(n9539), .Q(
        g1245), .QN(n9037) );
  SDFFX1 DFF_755_Q_reg ( .D(g27273), .SI(g1245), .SE(n9362), .CLK(n9549), .Q(
        g1262), .QN(n8570) );
  SDFFX1 DFF_756_Q_reg ( .D(g27285), .SI(g1262), .SE(n9362), .CLK(n9549), .Q(
        g1263) );
  SDFFX1 DFF_757_Q_reg ( .D(g27299), .SI(g1263), .SE(n9362), .CLK(n9549), .Q(
        g1261) );
  SDFFX1 DFF_758_Q_reg ( .D(g27286), .SI(g1261), .SE(n9362), .CLK(n9549), .Q(
        g1265), .QN(n8590) );
  SDFFX1 DFF_759_Q_reg ( .D(g27300), .SI(g1265), .SE(n9362), .CLK(n9549), .Q(
        g1266) );
  SDFFX1 DFF_760_Q_reg ( .D(g27314), .SI(g1266), .SE(n9362), .CLK(n9549), .Q(
        g1264) );
  SDFFX1 DFF_761_Q_reg ( .D(g27301), .SI(g1264), .SE(n9362), .CLK(n9549), .Q(
        g1268), .QN(n8397) );
  SDFFX1 DFF_762_Q_reg ( .D(g27315), .SI(g1268), .SE(n9362), .CLK(n9549), .Q(
        g1269) );
  SDFFX1 DFF_763_Q_reg ( .D(g27328), .SI(g1269), .SE(n9362), .CLK(n9549), .Q(
        test_so46) );
  SDFFX1 DFF_764_Q_reg ( .D(g27316), .SI(test_si47), .SE(n9362), .CLK(n9549), 
        .Q(g1271), .QN(n8604) );
  SDFFX1 DFF_765_Q_reg ( .D(g27329), .SI(g1271), .SE(n9363), .CLK(n9550), .Q(
        g1272) );
  SDFFX1 DFF_766_Q_reg ( .D(g27339), .SI(g1272), .SE(n9361), .CLK(n9548), .Q(
        g1270) );
  SDFFX1 DFF_767_Q_reg ( .D(g24501), .SI(g1270), .SE(n9361), .CLK(n9548), .Q(
        g1273), .QN(n8666) );
  SDFFX1 DFF_768_Q_reg ( .D(g24510), .SI(g1273), .SE(n9361), .CLK(n9548), .Q(
        g1276), .QN(n8668) );
  SDFFX1 DFF_769_Q_reg ( .D(g24521), .SI(g1276), .SE(n9361), .CLK(n9548), .Q(
        g1279), .QN(n8667) );
  SDFFX1 DFF_770_Q_reg ( .D(g24511), .SI(g1279), .SE(n9361), .CLK(n9548), .Q(
        g1282), .QN(n8653) );
  SDFFX1 DFF_771_Q_reg ( .D(g24522), .SI(g1282), .SE(n9362), .CLK(n9549), .Q(
        g1285), .QN(n8656) );
  SDFFX1 DFF_772_Q_reg ( .D(g24532), .SI(g1285), .SE(n9362), .CLK(n9549), .Q(
        g1288), .QN(n8655) );
  SDFFX1 DFF_773_Q_reg ( .D(g28351), .SI(g1288), .SE(n9363), .CLK(n9550), .Q(
        g1300) );
  SDFFX1 DFF_774_Q_reg ( .D(g28355), .SI(g1300), .SE(n9363), .CLK(n9550), .Q(
        g1303), .QN(n8686) );
  SDFFX1 DFF_775_Q_reg ( .D(g28360), .SI(g1303), .SE(n9363), .CLK(n9550), .Q(
        g1306), .QN(n8685) );
  SDFFX1 DFF_776_Q_reg ( .D(g28346), .SI(g1306), .SE(n9363), .CLK(n9550), .Q(
        g1291), .QN(n8692) );
  SDFFX1 DFF_777_Q_reg ( .D(g28350), .SI(g1291), .SE(n9363), .CLK(n9550), .Q(
        g1294) );
  SDFFX1 DFF_778_Q_reg ( .D(g28354), .SI(g1294), .SE(n9363), .CLK(n9550), .Q(
        g1297), .QN(n8693) );
  SDFFX1 DFF_779_Q_reg ( .D(g26547), .SI(g1297), .SE(n9363), .CLK(n9550), .Q(
        test_so47) );
  SDFFX1 DFF_780_Q_reg ( .D(g26557), .SI(test_si48), .SE(n9363), .CLK(n9550), 
        .Q(g1180), .QN(n8753) );
  SDFFX1 DFF_781_Q_reg ( .D(g26569), .SI(g1180), .SE(n9364), .CLK(n9551), .Q(
        g1183), .QN(n8749) );
  SDFFX1 DFF_782_Q_reg ( .D(g1186), .SI(g1183), .SE(n9364), .CLK(n9551), .Q(
        g1192), .QN(n4454) );
  SDFFX1 DFF_783_Q_reg ( .D(g22615), .SI(g1192), .SE(n9364), .CLK(n9551), .Q(
        n8009), .QN(DFF_783_n1) );
  SDFFX1 DFF_792_Q_reg ( .D(n549), .SI(n8009), .SE(n9364), .CLK(n9551), .Q(
        g16355), .QN(DFF_792_n1) );
  SDFFX1 DFF_793_Q_reg ( .D(g16355), .SI(g16355), .SE(n9364), .CLK(n9551), .Q(
        g1211), .QN(n8994) );
  SDFFX1 DFF_794_Q_reg ( .D(DFF_649_n1), .SI(g1211), .SE(n9364), .CLK(n9551), 
        .Q(n8008) );
  SDFFX1 DFF_795_Q_reg ( .D(DFF_651_n1), .SI(n8008), .SE(n9364), .CLK(n9551), 
        .Q(n8007), .QN(DFF_795_n1) );
  SDFFX1 DFF_796_Q_reg ( .D(DFF_653_n1), .SI(n8007), .SE(n9364), .CLK(n9551), 
        .Q(n8006), .QN(DFF_796_n1) );
  SDFFX1 DFF_797_Q_reg ( .D(DFF_655_n1), .SI(n8006), .SE(n9364), .CLK(n9551), 
        .Q(n8005) );
  SDFFX1 DFF_798_Q_reg ( .D(DFF_657_n1), .SI(n8005), .SE(n9364), .CLK(n9551), 
        .Q(n8004) );
  SDFFX1 DFF_799_Q_reg ( .D(DFF_659_n1), .SI(n8004), .SE(n9364), .CLK(n9551), 
        .Q(n8003) );
  SDFFX1 DFF_800_Q_reg ( .D(DFF_661_n1), .SI(n8003), .SE(n9364), .CLK(n9551), 
        .Q(g1222) );
  SDFFX1 DFF_801_Q_reg ( .D(DFF_663_n1), .SI(g1222), .SE(n9365), .CLK(n9552), 
        .Q(g1223) );
  SDFFX1 DFF_802_Q_reg ( .D(g24072), .SI(g1223), .SE(n9365), .CLK(n9552), .Q(
        g1224), .QN(n4489) );
  SDFFX1 DFF_803_Q_reg ( .D(n4486), .SI(g1224), .SE(n9365), .CLK(n9552), .Q(
        test_so48), .QN(n16819) );
  SDFFX1 DFF_805_Q_reg ( .D(g6979), .SI(g6979), .SE(n9324), .CLK(n9511), .Q(
        g7161), .QN(n4358) );
  SDFFX1 DFF_806_Q_reg ( .D(g7161), .SI(g7161), .SE(n9324), .CLK(n9511), .Q(
        g1315), .QN(n4294) );
  SDFFX1 DFF_807_Q_reg ( .D(g16671), .SI(g1315), .SE(n9349), .CLK(n9536), .Q(
        g1316), .QN(n9033) );
  SDFFX1 DFF_808_Q_reg ( .D(g20333), .SI(g1316), .SE(n9353), .CLK(n9540), .Q(
        g1345), .QN(n4428) );
  SDFFX1 DFF_809_Q_reg ( .D(g20717), .SI(g1345), .SE(n9353), .CLK(n9540), .Q(
        g1326), .QN(n4402) );
  SDFFX1 DFF_810_Q_reg ( .D(g21969), .SI(g1326), .SE(n9353), .CLK(n9540), .Q(
        g1319), .QN(n4476) );
  SDFFX1 DFF_811_Q_reg ( .D(g23329), .SI(g1319), .SE(n9353), .CLK(n9540), .Q(
        g1339), .QN(n4421) );
  SDFFX1 DFF_812_Q_reg ( .D(g24430), .SI(g1339), .SE(n9353), .CLK(n9540), .Q(
        g1332), .QN(n4412) );
  SDFFX1 DFF_813_Q_reg ( .D(g25189), .SI(g1332), .SE(n9353), .CLK(n9540), .Q(
        g1346), .QN(n4401) );
  SDFFX1 DFF_814_Q_reg ( .D(g26666), .SI(g1346), .SE(n9353), .CLK(n9540), .Q(
        g1358), .QN(n4411) );
  SDFFX1 DFF_815_Q_reg ( .D(g26781), .SI(g1358), .SE(n9353), .CLK(n9540), .Q(
        g1352), .QN(n4469) );
  SDFFX1 DFF_816_Q_reg ( .D(g27678), .SI(g1352), .SE(n9353), .CLK(n9540), .Q(
        g1365), .QN(n4475) );
  SDFFX1 DFF_817_Q_reg ( .D(g27718), .SI(g1365), .SE(n9353), .CLK(n9540), .Q(
        g1372), .QN(n4395) );
  SDFFX1 DFF_818_Q_reg ( .D(g28321), .SI(g1372), .SE(n9353), .CLK(n9540), .Q(
        g1378), .QN(n4417) );
  SDFFX1 DFF_819_Q_reg ( .D(g20882), .SI(g1378), .SE(n9365), .CLK(n9552), .Q(
        test_so49) );
  SDFFX1 DFF_820_Q_reg ( .D(g20896), .SI(test_si50), .SE(n9365), .CLK(n9552), 
        .Q(g1386), .QN(n9095) );
  SDFFX1 DFF_821_Q_reg ( .D(g20910), .SI(g1386), .SE(n9365), .CLK(n9552), .Q(
        g1384) );
  SDFFX1 DFF_822_Q_reg ( .D(g20897), .SI(g1384), .SE(n9365), .CLK(n9552), .Q(
        g1388) );
  SDFFX1 DFF_823_Q_reg ( .D(g20911), .SI(g1388), .SE(n9365), .CLK(n9552), .Q(
        g1389), .QN(n9093) );
  SDFFX1 DFF_824_Q_reg ( .D(g20925), .SI(g1389), .SE(n9365), .CLK(n9552), .Q(
        g1387) );
  SDFFX1 DFF_825_Q_reg ( .D(g20912), .SI(g1387), .SE(n9365), .CLK(n9552), .Q(
        g1391) );
  SDFFX1 DFF_826_Q_reg ( .D(g20926), .SI(g1391), .SE(n9365), .CLK(n9552), .Q(
        g1392), .QN(n9091) );
  SDFFX1 DFF_827_Q_reg ( .D(g20949), .SI(g1392), .SE(n9365), .CLK(n9552), .Q(
        g1390) );
  SDFFX1 DFF_828_Q_reg ( .D(g20927), .SI(g1390), .SE(n9366), .CLK(n9553), .Q(
        g1394) );
  SDFFX1 DFF_829_Q_reg ( .D(g20950), .SI(g1394), .SE(n9366), .CLK(n9553), .Q(
        g1395), .QN(n9089) );
  SDFFX1 DFF_830_Q_reg ( .D(g20972), .SI(g1395), .SE(n9366), .CLK(n9553), .Q(
        g1393) );
  SDFFX1 DFF_831_Q_reg ( .D(g20951), .SI(g1393), .SE(n9366), .CLK(n9553), .Q(
        g1397) );
  SDFFX1 DFF_832_Q_reg ( .D(g20973), .SI(g1397), .SE(n9366), .CLK(n9553), .Q(
        g1398), .QN(n9087) );
  SDFFX1 DFF_833_Q_reg ( .D(g20993), .SI(g1398), .SE(n9366), .CLK(n9553), .Q(
        g1396) );
  SDFFX1 DFF_834_Q_reg ( .D(g20974), .SI(g1396), .SE(n9366), .CLK(n9553), .Q(
        g1400) );
  SDFFX1 DFF_835_Q_reg ( .D(g20994), .SI(g1400), .SE(n9366), .CLK(n9553), .Q(
        test_so50) );
  SDFFX1 DFF_836_Q_reg ( .D(g21015), .SI(test_si51), .SE(n9366), .CLK(n9553), 
        .Q(g1399) );
  SDFFX1 DFF_837_Q_reg ( .D(g20995), .SI(g1399), .SE(n9366), .CLK(n9553), .Q(
        g1403) );
  SDFFX1 DFF_838_Q_reg ( .D(g21016), .SI(g1403), .SE(n9366), .CLK(n9553), .Q(
        g1404), .QN(n9084) );
  SDFFX1 DFF_839_Q_reg ( .D(g21033), .SI(g1404), .SE(n9366), .CLK(n9553), .Q(
        g1402) );
  SDFFX1 DFF_840_Q_reg ( .D(g21017), .SI(g1402), .SE(n9367), .CLK(n9554), .Q(
        g1406) );
  SDFFX1 DFF_841_Q_reg ( .D(g21034), .SI(g1406), .SE(n9367), .CLK(n9554), .Q(
        g1407), .QN(n9082) );
  SDFFX1 DFF_842_Q_reg ( .D(g21052), .SI(g1407), .SE(n9367), .CLK(n9554), .Q(
        g1405) );
  SDFFX1 DFF_843_Q_reg ( .D(g21035), .SI(g1405), .SE(n9367), .CLK(n9554), .Q(
        g1409) );
  SDFFX1 DFF_844_Q_reg ( .D(g21053), .SI(g1409), .SE(n9367), .CLK(n9554), .Q(
        g1410), .QN(n9080) );
  SDFFX1 DFF_845_Q_reg ( .D(g21070), .SI(g1410), .SE(n9367), .CLK(n9554), .Q(
        g1408) );
  SDFFX1 DFF_846_Q_reg ( .D(g20883), .SI(g1408), .SE(n9367), .CLK(n9554), .Q(
        g1412) );
  SDFFX1 DFF_847_Q_reg ( .D(g20898), .SI(g1412), .SE(n9367), .CLK(n9554), .Q(
        g1413), .QN(n9078) );
  SDFFX1 DFF_848_Q_reg ( .D(g20913), .SI(g1413), .SE(n9367), .CLK(n9554), .Q(
        g1411) );
  SDFFX1 DFF_849_Q_reg ( .D(g20952), .SI(g1411), .SE(n9367), .CLK(n9554), .Q(
        g1415) );
  SDFFX1 DFF_850_Q_reg ( .D(g20975), .SI(g1415), .SE(n9367), .CLK(n9554), .Q(
        g1416) );
  SDFFX1 DFF_851_Q_reg ( .D(g20996), .SI(g1416), .SE(n9367), .CLK(n9554), .Q(
        test_so51) );
  SDFFX1 DFF_852_Q_reg ( .D(g20976), .SI(test_si52), .SE(n9363), .CLK(n9550), 
        .Q(g1418) );
  SDFFX1 DFF_853_Q_reg ( .D(g20997), .SI(g1418), .SE(n9363), .CLK(n9550), .Q(
        g1419), .QN(n8841) );
  SDFFX1 DFF_854_Q_reg ( .D(g21018), .SI(g1419), .SE(n9363), .CLK(n9550), .Q(
        g1417) );
  SDFFX1 DFF_855_Q_reg ( .D(g25263), .SI(g1417), .SE(n9368), .CLK(n9555), .Q(
        g1421) );
  SDFFX1 DFF_856_Q_reg ( .D(g25267), .SI(g1421), .SE(n9368), .CLK(n9555), .Q(
        g1422) );
  SDFFX1 DFF_857_Q_reg ( .D(g25270), .SI(g1422), .SE(n9368), .CLK(n9555), .Q(
        g1420) );
  SDFFX1 DFF_858_Q_reg ( .D(n890), .SI(g1420), .SE(n9368), .CLK(n9555), .Q(
        g1424), .QN(n9154) );
  SDFFX1 DFF_859_Q_reg ( .D(g22247), .SI(g1424), .SE(n9368), .CLK(n9555), .Q(
        g1425) );
  SDFFX1 DFF_860_Q_reg ( .D(g22263), .SI(g1425), .SE(n9368), .CLK(n9555), .Q(
        g1423), .QN(n9221) );
  SDFFX1 DFF_861_Q_reg ( .D(g2950), .SI(g1423), .SE(n9368), .CLK(n9555), .Q(
        g6573), .QN(n4317) );
  SDFFX1 DFF_862_Q_reg ( .D(g6573), .SI(g6573), .SE(n9368), .CLK(n9555), .Q(
        g6782), .QN(n4515) );
  SDFFX1 DFF_863_Q_reg ( .D(g6782), .SI(g6782), .SE(n9368), .CLK(n9555), .Q(
        g1547), .QN(n4368) );
  SDFFX1 DFF_864_Q_reg ( .D(g22149), .SI(g1547), .SE(n9369), .CLK(n9556), .Q(
        g1512) );
  SDFFX1 DFF_865_Q_reg ( .D(g22166), .SI(g1512), .SE(n9373), .CLK(n9560), .Q(
        g1513), .QN(n9183) );
  SDFFX1 DFF_866_Q_reg ( .D(g22178), .SI(g1513), .SE(n9374), .CLK(n9561), .Q(
        g1511) );
  SDFFX1 DFF_867_Q_reg ( .D(g22167), .SI(g1511), .SE(n9369), .CLK(n9556), .Q(
        test_so52) );
  SDFFX1 DFF_868_Q_reg ( .D(g22179), .SI(test_si53), .SE(n9374), .CLK(n9561), 
        .Q(g1516), .QN(n9182) );
  SDFFX1 DFF_869_Q_reg ( .D(g22191), .SI(g1516), .SE(n9374), .CLK(n9561), .Q(
        g1514) );
  SDFFX1 DFF_870_Q_reg ( .D(g22035), .SI(g1514), .SE(n9375), .CLK(n9562), .Q(
        g1524) );
  SDFFX1 DFF_871_Q_reg ( .D(g22043), .SI(g1524), .SE(n9375), .CLK(n9562), .Q(
        g1525), .QN(n9180) );
  SDFFX1 DFF_872_Q_reg ( .D(g22057), .SI(g1525), .SE(n9375), .CLK(n9562), .Q(
        g1523) );
  SDFFX1 DFF_873_Q_reg ( .D(g22044), .SI(g1523), .SE(n9375), .CLK(n9562), .Q(
        g1527) );
  SDFFX1 DFF_874_Q_reg ( .D(g22058), .SI(g1527), .SE(n9375), .CLK(n9562), .Q(
        g1528), .QN(n9178) );
  SDFFX1 DFF_875_Q_reg ( .D(g22073), .SI(g1528), .SE(n9375), .CLK(n9562), .Q(
        g1526) );
  SDFFX1 DFF_876_Q_reg ( .D(g22059), .SI(g1526), .SE(n9375), .CLK(n9562), .Q(
        g1530) );
  SDFFX1 DFF_877_Q_reg ( .D(g22074), .SI(g1530), .SE(n9375), .CLK(n9562), .Q(
        g1531), .QN(n9176) );
  SDFFX1 DFF_878_Q_reg ( .D(g22090), .SI(g1531), .SE(n9375), .CLK(n9562), .Q(
        g1529) );
  SDFFX1 DFF_879_Q_reg ( .D(g22075), .SI(g1529), .SE(n9375), .CLK(n9562), .Q(
        g1533) );
  SDFFX1 DFF_880_Q_reg ( .D(g22091), .SI(g1533), .SE(n9375), .CLK(n9562), .Q(
        g1534), .QN(n9174) );
  SDFFX1 DFF_881_Q_reg ( .D(g22112), .SI(g1534), .SE(n9375), .CLK(n9562), .Q(
        g1532) );
  SDFFX1 DFF_882_Q_reg ( .D(g22092), .SI(g1532), .SE(n9376), .CLK(n9563), .Q(
        g1536) );
  SDFFX1 DFF_883_Q_reg ( .D(g22113), .SI(g1536), .SE(n9376), .CLK(n9563), .Q(
        test_so53) );
  SDFFX1 DFF_884_Q_reg ( .D(g22130), .SI(test_si54), .SE(n9373), .CLK(n9560), 
        .Q(g1535) );
  SDFFX1 DFF_885_Q_reg ( .D(g22114), .SI(g1535), .SE(n9373), .CLK(n9560), .Q(
        g1539) );
  SDFFX1 DFF_886_Q_reg ( .D(g22131), .SI(g1539), .SE(n9373), .CLK(n9560), .Q(
        g1540), .QN(n9171) );
  SDFFX1 DFF_887_Q_reg ( .D(g22150), .SI(g1540), .SE(n9373), .CLK(n9560), .Q(
        g1538) );
  SDFFX1 DFF_888_Q_reg ( .D(g22132), .SI(g1538), .SE(n9373), .CLK(n9560), .Q(
        g1542), .QN(n8789) );
  SDFFX1 DFF_889_Q_reg ( .D(g22151), .SI(g1542), .SE(n9373), .CLK(n9560), .Q(
        g1543) );
  SDFFX1 DFF_890_Q_reg ( .D(g22168), .SI(g1543), .SE(n9373), .CLK(n9560), .Q(
        g1541), .QN(n8787) );
  SDFFX1 DFF_891_Q_reg ( .D(g22152), .SI(g1541), .SE(n9374), .CLK(n9561), .Q(
        g1545), .QN(n8805) );
  SDFFX1 DFF_892_Q_reg ( .D(g22169), .SI(g1545), .SE(n9374), .CLK(n9561), .Q(
        g1546) );
  SDFFX1 DFF_893_Q_reg ( .D(g22180), .SI(g1546), .SE(n9374), .CLK(n9561), .Q(
        g1544), .QN(n8803) );
  SDFFX1 DFF_894_Q_reg ( .D(g25217), .SI(g1544), .SE(n9374), .CLK(n9561), .Q(
        g1551) );
  SDFFX1 DFF_895_Q_reg ( .D(g25224), .SI(g1551), .SE(n9374), .CLK(n9561), .Q(
        g1552), .QN(n8870) );
  SDFFX1 DFF_896_Q_reg ( .D(g25233), .SI(g1552), .SE(n9374), .CLK(n9561), .Q(
        g1550) );
  SDFFX1 DFF_897_Q_reg ( .D(g25225), .SI(g1550), .SE(n9374), .CLK(n9561), .Q(
        g1554) );
  SDFFX1 DFF_898_Q_reg ( .D(g25234), .SI(g1554), .SE(n9374), .CLK(n9561), .Q(
        g1555), .QN(n8867) );
  SDFFX1 DFF_899_Q_reg ( .D(g25242), .SI(g1555), .SE(n9374), .CLK(n9561), .Q(
        test_so54) );
  SDFFX1 DFF_900_Q_reg ( .D(g25235), .SI(test_si55), .SE(n9368), .CLK(n9555), 
        .Q(g1557) );
  SDFFX1 DFF_901_Q_reg ( .D(g25243), .SI(g1557), .SE(n9368), .CLK(n9555), .Q(
        g1558), .QN(n8865) );
  SDFFX1 DFF_902_Q_reg ( .D(g25249), .SI(g1558), .SE(n9368), .CLK(n9555), .Q(
        g1556) );
  SDFFX1 DFF_903_Q_reg ( .D(g25244), .SI(g1556), .SE(n9369), .CLK(n9556), .Q(
        g1560) );
  SDFFX1 DFF_904_Q_reg ( .D(g25250), .SI(g1560), .SE(n9369), .CLK(n9556), .Q(
        g1561), .QN(n8862) );
  SDFFX1 DFF_905_Q_reg ( .D(g25255), .SI(g1561), .SE(n9369), .CLK(n9556), .Q(
        g1559) );
  SDFFX1 DFF_906_Q_reg ( .D(g30279), .SI(g1559), .SE(n9380), .CLK(n9567), .Q(
        g1567), .QN(n8454) );
  SDFFX1 DFF_907_Q_reg ( .D(g30287), .SI(g1567), .SE(n9380), .CLK(n9567), .Q(
        g1570) );
  SDFFX1 DFF_908_Q_reg ( .D(g30294), .SI(g1570), .SE(n9380), .CLK(n9567), .Q(
        g1573), .QN(n8540) );
  SDFFX1 DFF_909_Q_reg ( .D(g30651), .SI(g1573), .SE(n9380), .CLK(n9567), .Q(
        g1612), .QN(n8452) );
  SDFFX1 DFF_910_Q_reg ( .D(g30657), .SI(g1612), .SE(n9380), .CLK(n9567), .Q(
        g1615) );
  SDFFX1 DFF_911_Q_reg ( .D(g30663), .SI(g1615), .SE(n9380), .CLK(n9567), .Q(
        g1618), .QN(n8423) );
  SDFFX1 DFF_912_Q_reg ( .D(g30683), .SI(g1618), .SE(n9380), .CLK(n9567), .Q(
        g1576), .QN(n8451) );
  SDFFX1 DFF_913_Q_reg ( .D(g30688), .SI(g1576), .SE(n9380), .CLK(n9567), .Q(
        g1579) );
  SDFFX1 DFF_914_Q_reg ( .D(g30692), .SI(g1579), .SE(n9380), .CLK(n9567), .Q(
        g1582), .QN(n8539) );
  SDFFX1 DFF_915_Q_reg ( .D(g30658), .SI(g1582), .SE(n9380), .CLK(n9567), .Q(
        test_so55) );
  SDFFX1 DFF_916_Q_reg ( .D(g30664), .SI(test_si56), .SE(n9376), .CLK(n9563), 
        .Q(g1624) );
  SDFFX1 DFF_917_Q_reg ( .D(g30671), .SI(g1624), .SE(n9376), .CLK(n9563), .Q(
        g1627), .QN(n8422) );
  SDFFX1 DFF_918_Q_reg ( .D(g30295), .SI(g1627), .SE(n9377), .CLK(n9564), .Q(
        g1585), .QN(n8449) );
  SDFFX1 DFF_919_Q_reg ( .D(g30299), .SI(g1585), .SE(n9377), .CLK(n9564), .Q(
        g1588) );
  SDFFX1 DFF_920_Q_reg ( .D(g30302), .SI(g1588), .SE(n9369), .CLK(n9556), .Q(
        g1591), .QN(n8531) );
  SDFFX1 DFF_921_Q_reg ( .D(g30266), .SI(g1591), .SE(n9369), .CLK(n9556), .Q(
        g1630), .QN(n8447) );
  SDFFX1 DFF_922_Q_reg ( .D(g30272), .SI(g1630), .SE(n9369), .CLK(n9556), .Q(
        g1633) );
  SDFFX1 DFF_923_Q_reg ( .D(g30280), .SI(g1633), .SE(n9369), .CLK(n9556), .Q(
        g1636), .QN(n8421) );
  SDFFX1 DFF_924_Q_reg ( .D(g30250), .SI(g1636), .SE(n9376), .CLK(n9563), .Q(
        g1594), .QN(n8445) );
  SDFFX1 DFF_925_Q_reg ( .D(g30252), .SI(g1594), .SE(n9376), .CLK(n9563), .Q(
        g1597) );
  SDFFX1 DFF_926_Q_reg ( .D(g30255), .SI(g1597), .SE(n9376), .CLK(n9563), .Q(
        g1600), .QN(n8538) );
  SDFFX1 DFF_927_Q_reg ( .D(g30273), .SI(g1600), .SE(n9376), .CLK(n9563), .Q(
        g1639), .QN(n8443) );
  SDFFX1 DFF_928_Q_reg ( .D(g30281), .SI(g1639), .SE(n9376), .CLK(n9563), .Q(
        g1642) );
  SDFFX1 DFF_929_Q_reg ( .D(g30288), .SI(g1642), .SE(n9376), .CLK(n9563), .Q(
        g1645), .QN(n8528) );
  SDFFX1 DFF_930_Q_reg ( .D(g30644), .SI(g1645), .SE(n9376), .CLK(n9563), .Q(
        g1603), .QN(n8379) );
  SDFFX1 DFF_931_Q_reg ( .D(g30650), .SI(g1603), .SE(n9376), .CLK(n9563), .Q(
        test_so56) );
  SDFFX1 DFF_932_Q_reg ( .D(g30656), .SI(test_si57), .SE(n9370), .CLK(n9557), 
        .Q(g1609), .QN(n8385) );
  SDFFX1 DFF_933_Q_reg ( .D(g30678), .SI(g1609), .SE(n9370), .CLK(n9557), .Q(
        g1648), .QN(n8412) );
  SDFFX1 DFF_934_Q_reg ( .D(g30684), .SI(g1648), .SE(n9370), .CLK(n9557), .Q(
        g1651) );
  SDFFX1 DFF_935_Q_reg ( .D(g30689), .SI(g1651), .SE(n9370), .CLK(n9557), .Q(
        g1654), .QN(n8413) );
  SDFFX1 DFF_936_Q_reg ( .D(g25056), .SI(g1654), .SE(n9370), .CLK(n9557), .Q(
        g1466), .QN(n8976) );
  SDFFX1 DFF_937_Q_reg ( .D(n50), .SI(g1466), .SE(n9370), .CLK(n9557), .Q(
        g1462), .QN(n9265) );
  SDFFX1 DFF_938_Q_reg ( .D(g26531), .SI(g1462), .SE(n9370), .CLK(n9557), .Q(
        g1457), .QN(n8975) );
  SDFFX1 DFF_939_Q_reg ( .D(n51), .SI(g1457), .SE(n9370), .CLK(n9557), .Q(
        g1453), .QN(n9270) );
  SDFFX1 DFF_940_Q_reg ( .D(g27612), .SI(g1453), .SE(n9370), .CLK(n9557), .Q(
        g1448), .QN(n8974) );
  SDFFX1 DFF_941_Q_reg ( .D(g28147), .SI(g1448), .SE(n9370), .CLK(n9557), .Q(
        g1444), .QN(n9276) );
  SDFFX1 DFF_942_Q_reg ( .D(g28636), .SI(g1444), .SE(n9370), .CLK(n9557), .Q(
        g1439), .QN(n8973) );
  SDFFX1 DFF_943_Q_reg ( .D(g29111), .SI(g1439), .SE(n9370), .CLK(n9557), .Q(
        g1435), .QN(n9267) );
  SDFFX1 DFF_944_Q_reg ( .D(g29355), .SI(g1435), .SE(n9371), .CLK(n9558), .Q(
        g1430), .QN(n8560) );
  SDFFX1 DFF_945_Q_reg ( .D(g29581), .SI(g1430), .SE(n9371), .CLK(n9558), .Q(
        g1426), .QN(n8389) );
  SDFFX1 DFF_946_Q_reg ( .D(n15), .SI(g1426), .SE(n9371), .CLK(n9558), .Q(
        g1562) );
  SDFFX1 DFF_947_Q_reg ( .D(g1562), .SI(g1562), .SE(n9371), .CLK(n9558), .Q(
        test_so57) );
  SDFFX1 DFF_948_Q_reg ( .D(test_so57), .SI(test_si58), .SE(n9371), .CLK(n9558), .Q(g1563), .QN(n8989) );
  SDFFX1 DFF_949_Q_reg ( .D(g2950), .SI(g1563), .SE(n9371), .CLK(n9558), .Q(
        g5511), .QN(n4518) );
  SDFFX1 DFF_952_Q_reg ( .D(test_so57), .SI(n4618), .SE(n9371), .CLK(n9558), 
        .Q(g1690), .QN(n4386) );
  SDFFX1 DFF_953_Q_reg ( .D(g27264), .SI(g1690), .SE(n9379), .CLK(n9566), .Q(
        g1735) );
  SDFFX1 DFF_954_Q_reg ( .D(g27274), .SI(g1735), .SE(n9379), .CLK(n9566), .Q(
        g1724), .QN(n8929) );
  SDFFX1 DFF_955_Q_reg ( .D(g27287), .SI(g1724), .SE(n9379), .CLK(n9566), .Q(
        g1727) );
  SDFFX1 DFF_956_Q_reg ( .D(g27275), .SI(g1727), .SE(n9379), .CLK(n9566), .Q(
        g1750) );
  SDFFX1 DFF_957_Q_reg ( .D(g27288), .SI(g1750), .SE(n9379), .CLK(n9566), .Q(
        g1739), .QN(n8906) );
  SDFFX1 DFF_958_Q_reg ( .D(g27302), .SI(g1739), .SE(n9379), .CLK(n9566), .Q(
        g1742) );
  SDFFX1 DFF_959_Q_reg ( .D(g27289), .SI(g1742), .SE(n9379), .CLK(n9566), .Q(
        g1765) );
  SDFFX1 DFF_960_Q_reg ( .D(g27303), .SI(g1765), .SE(n9379), .CLK(n9566), .Q(
        g1754), .QN(n8640) );
  SDFFX1 DFF_961_Q_reg ( .D(g27317), .SI(g1754), .SE(n9379), .CLK(n9566), .Q(
        g1757) );
  SDFFX1 DFF_962_Q_reg ( .D(g27304), .SI(g1757), .SE(n9380), .CLK(n9567), .Q(
        g1779) );
  SDFFX1 DFF_963_Q_reg ( .D(g27318), .SI(g1779), .SE(n9380), .CLK(n9567), .Q(
        test_so58) );
  SDFFX1 DFF_964_Q_reg ( .D(g27330), .SI(test_si59), .SE(n9377), .CLK(n9564), 
        .Q(g1772) );
  SDFFX1 DFF_965_Q_reg ( .D(g28749), .SI(g1772), .SE(n9377), .CLK(n9564), .Q(
        g1789) );
  SDFFX1 DFF_966_Q_reg ( .D(g28760), .SI(g1789), .SE(n9378), .CLK(n9565), .Q(
        g1792), .QN(n8707) );
  SDFFX1 DFF_967_Q_reg ( .D(g28771), .SI(g1792), .SE(n9378), .CLK(n9565), .Q(
        g1795), .QN(n8723) );
  SDFFX1 DFF_968_Q_reg ( .D(g29205), .SI(g1795), .SE(n9379), .CLK(n9566), .Q(
        g1798) );
  SDFFX1 DFF_969_Q_reg ( .D(g29212), .SI(g1798), .SE(n9379), .CLK(n9566), .Q(
        g1801), .QN(n8706) );
  SDFFX1 DFF_970_Q_reg ( .D(g29218), .SI(g1801), .SE(n9377), .CLK(n9564), .Q(
        g1804), .QN(n8721) );
  SDFFX1 DFF_971_Q_reg ( .D(g28761), .SI(g1804), .SE(n9377), .CLK(n9564), .Q(
        g1808) );
  SDFFX1 DFF_972_Q_reg ( .D(g28772), .SI(g1808), .SE(n9377), .CLK(n9564), .Q(
        g1809), .QN(n8941) );
  SDFFX1 DFF_973_Q_reg ( .D(g28778), .SI(g1809), .SE(n9377), .CLK(n9564), .Q(
        g1807) );
  SDFFX1 DFF_974_Q_reg ( .D(g26811), .SI(g1807), .SE(n9377), .CLK(n9564), .Q(
        g1810) );
  SDFFX1 DFF_975_Q_reg ( .D(g26815), .SI(g1810), .SE(n9378), .CLK(n9565), .Q(
        g1813), .QN(n8705) );
  SDFFX1 DFF_976_Q_reg ( .D(g26820), .SI(g1813), .SE(n9378), .CLK(n9565), .Q(
        g1816), .QN(n8719) );
  SDFFX1 DFF_977_Q_reg ( .D(g26816), .SI(g1816), .SE(n9378), .CLK(n9565), .Q(
        g1819) );
  SDFFX1 DFF_978_Q_reg ( .D(g26821), .SI(g1819), .SE(n9378), .CLK(n9565), .Q(
        g1822), .QN(n8704) );
  SDFFX1 DFF_979_Q_reg ( .D(g26824), .SI(g1822), .SE(n9378), .CLK(n9565), .Q(
        test_so59) );
  SDFFX1 DFF_980_Q_reg ( .D(g27764), .SI(test_si60), .SE(n9378), .CLK(n9565), 
        .Q(g1829), .QN(n8951) );
  SDFFX1 DFF_981_Q_reg ( .D(g27766), .SI(g1829), .SE(n9378), .CLK(n9565), .Q(
        g1830), .QN(n8940) );
  SDFFX1 DFF_982_Q_reg ( .D(g27768), .SI(g1830), .SE(n9378), .CLK(n9565), .Q(
        g1828), .QN(n8950) );
  SDFFX1 DFF_983_Q_reg ( .D(g29613), .SI(g1828), .SE(n9378), .CLK(n9565), .Q(
        g1693) );
  SDFFX1 DFF_984_Q_reg ( .D(g29617), .SI(g1693), .SE(n9378), .CLK(n9565), .Q(
        g1694), .QN(n8498) );
  SDFFX1 DFF_985_Q_reg ( .D(g29620), .SI(g1694), .SE(n9377), .CLK(n9564), .Q(
        g1695) );
  SDFFX1 DFF_986_Q_reg ( .D(g30704), .SI(g1695), .SE(n9377), .CLK(n9564), .Q(
        g1696) );
  SDFFX1 DFF_987_Q_reg ( .D(g30706), .SI(g1696), .SE(n9377), .CLK(n9564), .Q(
        g1697), .QN(n8497) );
  SDFFX1 DFF_988_Q_reg ( .D(g30708), .SI(g1697), .SE(n9369), .CLK(n9556), .Q(
        g1698) );
  SDFFX1 DFF_989_Q_reg ( .D(g30487), .SI(g1698), .SE(n9371), .CLK(n9558), .Q(
        g1699) );
  SDFFX1 DFF_990_Q_reg ( .D(g30503), .SI(g1699), .SE(n9369), .CLK(n9556), .Q(
        g1700), .QN(n8496) );
  SDFFX1 DFF_991_Q_reg ( .D(g30338), .SI(g1700), .SE(n9371), .CLK(n9558), .Q(
        g1701) );
  SDFFX1 DFF_992_Q_reg ( .D(g29178), .SI(g1701), .SE(n9381), .CLK(n9568), .Q(
        g1703) );
  SDFFX1 DFF_993_Q_reg ( .D(g29181), .SI(g1703), .SE(n9381), .CLK(n9568), .Q(
        g1704), .QN(n8548) );
  SDFFX1 DFF_994_Q_reg ( .D(g29184), .SI(g1704), .SE(n9369), .CLK(n9556), .Q(
        g1702) );
  SDFFX1 DFF_995_Q_reg ( .D(g26667), .SI(g1702), .SE(n9371), .CLK(n9558), .Q(
        test_so60) );
  SDFFX1 DFF_996_Q_reg ( .D(g26670), .SI(test_si61), .SE(n9372), .CLK(n9559), 
        .Q(g1785), .QN(n8939) );
  SDFFX1 DFF_997_Q_reg ( .D(g26675), .SI(g1785), .SE(n9372), .CLK(n9559), .Q(
        g1783) );
  SDFFX1 DFF_998_Q_reg ( .D(n4288), .SI(g1783), .SE(n9372), .CLK(n9559), .Q(
        g1831) );
  SDFFX1 DFF_999_Q_reg ( .D(g1831), .SI(g1831), .SE(n9372), .CLK(n9559), .Q(
        n7988), .QN(DFF_999_n1) );
  SDFFX1 DFF_1000_Q_reg ( .D(n4565), .SI(n7988), .SE(n9372), .CLK(n9559), .Q(
        g1833) );
  SDFFX1 DFF_1001_Q_reg ( .D(g1833), .SI(g1833), .SE(n9372), .CLK(n9559), .Q(
        n7987), .QN(DFF_1001_n1) );
  SDFFX1 DFF_1002_Q_reg ( .D(n4557), .SI(n7987), .SE(n9372), .CLK(n9559), .Q(
        g1835) );
  SDFFX1 DFF_1003_Q_reg ( .D(g1835), .SI(g1835), .SE(n9372), .CLK(n9559), .Q(
        n7986), .QN(DFF_1003_n1) );
  SDFFX1 DFF_1004_Q_reg ( .D(n4326), .SI(n7986), .SE(n9372), .CLK(n9559), .Q(
        g1661) );
  SDFFX1 DFF_1005_Q_reg ( .D(g1661), .SI(g1661), .SE(n9372), .CLK(n9559), .Q(
        n7985), .QN(DFF_1005_n1) );
  SDFFX1 DFF_1006_Q_reg ( .D(n4390), .SI(n7985), .SE(n9372), .CLK(n9559), .Q(
        g1663) );
  SDFFX1 DFF_1007_Q_reg ( .D(g1663), .SI(g1663), .SE(n9372), .CLK(n9559), .Q(
        n7984), .QN(DFF_1007_n1) );
  SDFFX1 DFF_1008_Q_reg ( .D(n4320), .SI(n7984), .SE(n9373), .CLK(n9560), .Q(
        g1665) );
  SDFFX1 DFF_1009_Q_reg ( .D(g1665), .SI(g1665), .SE(n9373), .CLK(n9560), .Q(
        n7983), .QN(DFF_1009_n1) );
  SDFFX1 DFF_1010_Q_reg ( .D(n4374), .SI(n7983), .SE(n9373), .CLK(n9560), .Q(
        g1667) );
  SDFFX1 DFF_1011_Q_reg ( .D(g1667), .SI(g1667), .SE(n9373), .CLK(n9560), .Q(
        test_so61), .QN(DFF_1011_n1) );
  SDFFX1 DFF_1012_Q_reg ( .D(n4378), .SI(test_si62), .SE(n9295), .CLK(n9482), 
        .Q(g1669) );
  SDFFX1 DFF_1013_Q_reg ( .D(g1669), .SI(g1669), .SE(n9295), .CLK(n9482), .Q(
        n7980), .QN(DFF_1013_n1) );
  SDFFX1 DFF_1014_Q_reg ( .D(g2877), .SI(n7980), .SE(n9300), .CLK(n9487), .Q(
        g1671) );
  SDFFX1 DFF_1015_Q_reg ( .D(g1671), .SI(g1671), .SE(n9300), .CLK(n9487), .Q(
        n7979), .QN(n4484) );
  SDFFX1 DFF_1016_Q_reg ( .D(n4284), .SI(n7979), .SE(n9379), .CLK(n9566), .Q(
        g1680), .QN(n4488) );
  SDFFX1 DFF_1017_Q_reg ( .D(n478), .SI(g1680), .SE(n9381), .CLK(n9568), .Q(
        g1686), .QN(n8986) );
  SDFFX1 DFF_1028_Q_reg ( .D(n4276), .SI(g1686), .SE(n9381), .CLK(n9568), .Q(
        n7978) );
  SDFFX1 DFF_1029_Q_reg ( .D(g1735), .SI(n7978), .SE(n9381), .CLK(n9568), .Q(
        g1723) );
  SDFFX1 DFF_1030_Q_reg ( .D(g1723), .SI(g1723), .SE(n9381), .CLK(n9568), .Q(
        g1730) );
  SDFFX1 DFF_1031_Q_reg ( .D(g1724), .SI(g1730), .SE(n9381), .CLK(n9568), .Q(
        g1731) );
  SDFFX1 DFF_1032_Q_reg ( .D(g1731), .SI(g1731), .SE(n9381), .CLK(n9568), .Q(
        g1732), .QN(n8616) );
  SDFFX1 DFF_1033_Q_reg ( .D(g1727), .SI(g1732), .SE(n9381), .CLK(n9568), .Q(
        g1733) );
  SDFFX1 DFF_1034_Q_reg ( .D(g1733), .SI(g1733), .SE(n9381), .CLK(n9568), .Q(
        g1734), .QN(n8615) );
  SDFFX1 DFF_1035_Q_reg ( .D(g1750), .SI(g1734), .SE(n9381), .CLK(n9568), .Q(
        g1738) );
  SDFFX1 DFF_1036_Q_reg ( .D(g1738), .SI(g1738), .SE(n9381), .CLK(n9568), .Q(
        g1745) );
  SDFFX1 DFF_1037_Q_reg ( .D(g1739), .SI(g1745), .SE(n9382), .CLK(n9569), .Q(
        test_so62) );
  SDFFX1 DFF_1038_Q_reg ( .D(test_so62), .SI(test_si63), .SE(n9382), .CLK(
        n9569), .Q(g1747), .QN(n8405) );
  SDFFX1 DFF_1039_Q_reg ( .D(g1742), .SI(g1747), .SE(n9382), .CLK(n9569), .Q(
        g1748) );
  SDFFX1 DFF_1040_Q_reg ( .D(g1748), .SI(g1748), .SE(n9382), .CLK(n9569), .Q(
        g1749), .QN(n8404) );
  SDFFX1 DFF_1041_Q_reg ( .D(g1765), .SI(g1749), .SE(n9382), .CLK(n9569), .Q(
        g1753) );
  SDFFX1 DFF_1042_Q_reg ( .D(g1753), .SI(g1753), .SE(n9382), .CLK(n9569), .Q(
        g1760) );
  SDFFX1 DFF_1043_Q_reg ( .D(g1754), .SI(g1760), .SE(n9382), .CLK(n9569), .Q(
        g1761) );
  SDFFX1 DFF_1044_Q_reg ( .D(g1761), .SI(g1761), .SE(n9382), .CLK(n9569), .Q(
        g1762), .QN(n8579) );
  SDFFX1 DFF_1045_Q_reg ( .D(g1757), .SI(g1762), .SE(n9382), .CLK(n9569), .Q(
        g1763) );
  SDFFX1 DFF_1046_Q_reg ( .D(g1763), .SI(g1763), .SE(n9382), .CLK(n9569), .Q(
        g1764), .QN(n8578) );
  SDFFX1 DFF_1047_Q_reg ( .D(g1779), .SI(g1764), .SE(n9382), .CLK(n9569), .Q(
        g1768) );
  SDFFX1 DFF_1048_Q_reg ( .D(g1768), .SI(g1768), .SE(n9382), .CLK(n9569), .Q(
        g1775) );
  SDFFX1 DFF_1049_Q_reg ( .D(test_so58), .SI(g1775), .SE(n9383), .CLK(n9570), 
        .Q(g1776) );
  SDFFX1 DFF_1050_Q_reg ( .D(g1776), .SI(g1776), .SE(n9383), .CLK(n9570), .Q(
        g1777), .QN(n8624) );
  SDFFX1 DFF_1051_Q_reg ( .D(g1772), .SI(g1777), .SE(n9383), .CLK(n9570), .Q(
        g1778) );
  SDFFX1 DFF_1052_Q_reg ( .D(g1778), .SI(g1778), .SE(n9383), .CLK(n9570), .Q(
        g1705), .QN(n8622) );
  SDFFX1 DFF_1053_Q_reg ( .D(n4598), .SI(g1705), .SE(n9383), .CLK(n9570), .Q(
        test_so63) );
  SDFFX1 DFF_1054_Q_reg ( .D(test_so63), .SI(test_si64), .SE(n9383), .CLK(
        n9570), .Q(g5738), .QN(n8623) );
  SDFFX1 DFF_1055_Q_reg ( .D(g5738), .SI(g5738), .SE(n9383), .CLK(n9570), .Q(
        g1718), .QN(n8621) );
  SDFFX1 DFF_1056_Q_reg ( .D(n4598), .SI(g1718), .SE(n9383), .CLK(n9570), .Q(
        g7052), .QN(n4296) );
  SDFFX1 DFF_1057_Q_reg ( .D(g7052), .SI(g7052), .SE(n9383), .CLK(n9570), .Q(
        g7194), .QN(n4315) );
  SDFFX1 DFF_1058_Q_reg ( .D(g7194), .SI(g7194), .SE(n9383), .CLK(n9570), .Q(
        g1930), .QN(n4366) );
  SDFFX1 DFF_1059_Q_reg ( .D(n1159), .SI(g1930), .SE(n9383), .CLK(n9570), .Q(
        g1934), .QN(n9224) );
  SDFFX1 DFF_1060_Q_reg ( .D(g18743), .SI(g1934), .SE(n9383), .CLK(n9570), .Q(
        g1937), .QN(n4311) );
  SDFFX1 DFF_1061_Q_reg ( .D(g18794), .SI(g1937), .SE(n9384), .CLK(n9571), .Q(
        g1890), .QN(n4297) );
  SDFFX1 DFF_1062_Q_reg ( .D(n1152), .SI(g1890), .SE(n9385), .CLK(n9572), .Q(
        g1893) );
  SDFFX1 DFF_1063_Q_reg ( .D(g1893), .SI(g1893), .SE(n9385), .CLK(n9572), .Q(
        g1903) );
  SDFFX1 DFF_1064_Q_reg ( .D(g1903), .SI(g1903), .SE(n9385), .CLK(n9572), .Q(
        g1904) );
  SDFFX1 DFF_1065_Q_reg ( .D(g1836), .SI(g1904), .SE(n9385), .CLK(n9572), .Q(
        g1944) );
  SDFFX1 DFF_1066_Q_reg ( .D(g1944), .SI(g1944), .SE(n9385), .CLK(n9572), .Q(
        g1949), .QN(n8774) );
  SDFFX1 DFF_1067_Q_reg ( .D(test_so65), .SI(g1949), .SE(n9385), .CLK(n9572), 
        .Q(g1950) );
  SDFFX1 DFF_1068_Q_reg ( .D(g1950), .SI(g1950), .SE(n9385), .CLK(n9572), .Q(
        g1951), .QN(n16826) );
  SDFFX1 DFF_1069_Q_reg ( .D(g1842), .SI(g1951), .SE(n9385), .CLK(n9572), .Q(
        test_so64) );
  SDFFX1 DFF_1070_Q_reg ( .D(test_so64), .SI(test_si65), .SE(n9385), .CLK(
        n9572), .Q(g1953) );
  SDFFX1 DFF_1071_Q_reg ( .D(g1846), .SI(g1953), .SE(n9385), .CLK(n9572), .Q(
        g1954) );
  SDFFX1 DFF_1072_Q_reg ( .D(g1954), .SI(g1954), .SE(n9385), .CLK(n9572), .Q(
        g1945), .QN(n8772) );
  SDFFX1 DFF_1073_Q_reg ( .D(g1849), .SI(g1945), .SE(n9386), .CLK(n9573), .Q(
        g1946) );
  SDFFX1 DFF_1074_Q_reg ( .D(g1946), .SI(g1946), .SE(n9386), .CLK(n9573), .Q(
        g1947), .QN(n16828) );
  SDFFX1 DFF_1075_Q_reg ( .D(g1852), .SI(g1947), .SE(n9386), .CLK(n9573), .Q(
        g1948) );
  SDFFX1 DFF_1076_Q_reg ( .D(g1948), .SI(g1948), .SE(n9386), .CLK(n9573), .Q(
        g1870) );
  SDFFX1 DFF_1077_Q_reg ( .D(g2950), .SI(g1870), .SE(n9386), .CLK(n9573), .Q(
        g8012), .QN(n4458) );
  SDFFX1 DFF_1078_Q_reg ( .D(g8012), .SI(g8012), .SE(n9386), .CLK(n9573), .Q(
        g8082), .QN(n4457) );
  SDFFX1 DFF_1079_Q_reg ( .D(g8082), .SI(g8082), .SE(n9386), .CLK(n9573), .Q(
        g1866), .QN(n4464) );
  SDFFX1 DFF_1080_Q_reg ( .D(g23097), .SI(g1866), .SE(n9386), .CLK(n9573), .Q(
        g1867), .QN(n9004) );
  SDFFX1 DFF_1081_Q_reg ( .D(g23124), .SI(g1867), .SE(n9386), .CLK(n9573), .Q(
        g1868) );
  SDFFX1 DFF_1082_Q_reg ( .D(g23137), .SI(g1868), .SE(n9386), .CLK(n9573), .Q(
        g1869), .QN(n9005) );
  SDFFX1 DFF_1083_Q_reg ( .D(g23400), .SI(g1869), .SE(n9386), .CLK(n9573), .Q(
        g1836) );
  SDFFX1 DFF_1084_Q_reg ( .D(g23413), .SI(g1836), .SE(n9387), .CLK(n9574), .Q(
        test_so65) );
  SDFFX1 DFF_1085_Q_reg ( .D(g24182), .SI(test_si66), .SE(n9386), .CLK(n9573), 
        .Q(g1842) );
  SDFFX1 DFF_1086_Q_reg ( .D(g24208), .SI(g1842), .SE(n9387), .CLK(n9574), .Q(
        g1858), .QN(n9010) );
  SDFFX1 DFF_1087_Q_reg ( .D(g24219), .SI(g1858), .SE(n9387), .CLK(n9574), .Q(
        g1859) );
  SDFFX1 DFF_1088_Q_reg ( .D(g24231), .SI(g1859), .SE(n9387), .CLK(n9574), .Q(
        g1860), .QN(n9011) );
  SDFFX1 DFF_1089_Q_reg ( .D(g23123), .SI(g1860), .SE(n9387), .CLK(n9574), .Q(
        g1861), .QN(n9007) );
  SDFFX1 DFF_1090_Q_reg ( .D(g23030), .SI(g1861), .SE(n9387), .CLK(n9574), .Q(
        g1865) );
  SDFFX1 DFF_1091_Q_reg ( .D(g23058), .SI(g1865), .SE(n9387), .CLK(n9574), .Q(
        g1845), .QN(n9008) );
  SDFFX1 DFF_1092_Q_reg ( .D(g24218), .SI(g1845), .SE(n9387), .CLK(n9574), .Q(
        g1846) );
  SDFFX1 DFF_1093_Q_reg ( .D(g24230), .SI(g1846), .SE(n9387), .CLK(n9574), .Q(
        g1849) );
  SDFFX1 DFF_1094_Q_reg ( .D(g24243), .SI(g1849), .SE(n9387), .CLK(n9574), .Q(
        g1852) );
  SDFFX1 DFF_1095_Q_reg ( .D(n1149), .SI(g1852), .SE(n9387), .CLK(n9574), .Q(
        g1908) );
  SDFFX1 DFF_1096_Q_reg ( .D(g1908), .SI(g1908), .SE(n9387), .CLK(n9574), .Q(
        g1915) );
  SDFFX1 DFF_1097_Q_reg ( .D(g1915), .SI(g1915), .SE(n9388), .CLK(n9575), .Q(
        g1922) );
  SDFFX1 DFF_1098_Q_reg ( .D(g13164), .SI(g1922), .SE(n9388), .CLK(n9575), .Q(
        g1923) );
  SDFFX1 DFF_1099_Q_reg ( .D(g1923), .SI(g1923), .SE(n9388), .CLK(n9575), .Q(
        test_so66), .QN(DFF_1099_n1) );
  SDFFX1 DFF_1100_Q_reg ( .D(n532), .SI(test_si67), .SE(n9388), .CLK(n9575), 
        .Q(n7971), .QN(DFF_1100_n1) );
  SDFFX1 DFF_1101_Q_reg ( .D(g13135), .SI(n7971), .SE(n9388), .CLK(n9575), .Q(
        g1929) );
  SDFFX1 DFF_1102_Q_reg ( .D(g1929), .SI(g1929), .SE(n9388), .CLK(n9575), .Q(
        g1880), .QN(n4545) );
  SDFFX1 DFF_1103_Q_reg ( .D(g13182), .SI(g1880), .SE(n9388), .CLK(n9575), .Q(
        g1938) );
  SDFFX1 DFF_1104_Q_reg ( .D(g1938), .SI(g1938), .SE(n9388), .CLK(n9575), .Q(
        g1939), .QN(n9036) );
  SDFFX1 DFF_1105_Q_reg ( .D(g27290), .SI(g1939), .SE(n9389), .CLK(n9576), .Q(
        g1956) );
  SDFFX1 DFF_1106_Q_reg ( .D(g27305), .SI(g1956), .SE(n9389), .CLK(n9576), .Q(
        g1957) );
  SDFFX1 DFF_1107_Q_reg ( .D(g27319), .SI(g1957), .SE(n9389), .CLK(n9576), .Q(
        g1955), .QN(n8568) );
  SDFFX1 DFF_1108_Q_reg ( .D(g27306), .SI(g1955), .SE(n9389), .CLK(n9576), .Q(
        g1959) );
  SDFFX1 DFF_1109_Q_reg ( .D(g27320), .SI(g1959), .SE(n9389), .CLK(n9576), .Q(
        g1960) );
  SDFFX1 DFF_1110_Q_reg ( .D(g27331), .SI(g1960), .SE(n9389), .CLK(n9576), .Q(
        g1958), .QN(n8588) );
  SDFFX1 DFF_1111_Q_reg ( .D(g27321), .SI(g1958), .SE(n9389), .CLK(n9576), .Q(
        g1962) );
  SDFFX1 DFF_1112_Q_reg ( .D(g27332), .SI(g1962), .SE(n9389), .CLK(n9576), .Q(
        g1963) );
  SDFFX1 DFF_1113_Q_reg ( .D(g27340), .SI(g1963), .SE(n9389), .CLK(n9576), .Q(
        g1961), .QN(n8395) );
  SDFFX1 DFF_1114_Q_reg ( .D(g27333), .SI(g1961), .SE(n9389), .CLK(n9576), .Q(
        test_so67) );
  SDFFX1 DFF_1115_Q_reg ( .D(g27341), .SI(test_si68), .SE(n9390), .CLK(n9577), 
        .Q(g1966) );
  SDFFX1 DFF_1116_Q_reg ( .D(g27346), .SI(g1966), .SE(n9390), .CLK(n9577), .Q(
        g1964), .QN(n8602) );
  SDFFX1 DFF_1117_Q_reg ( .D(g24513), .SI(g1964), .SE(n9390), .CLK(n9577), .Q(
        g1967), .QN(n8663) );
  SDFFX1 DFF_1118_Q_reg ( .D(g24524), .SI(g1967), .SE(n9390), .CLK(n9577), .Q(
        g1970), .QN(n8665) );
  SDFFX1 DFF_1119_Q_reg ( .D(g24534), .SI(g1970), .SE(n9390), .CLK(n9577), .Q(
        g1973), .QN(n8664) );
  SDFFX1 DFF_1120_Q_reg ( .D(g24525), .SI(g1973), .SE(n9390), .CLK(n9577), .Q(
        g1976), .QN(n8650) );
  SDFFX1 DFF_1121_Q_reg ( .D(g24535), .SI(g1976), .SE(n9390), .CLK(n9577), .Q(
        g1979), .QN(n8652) );
  SDFFX1 DFF_1122_Q_reg ( .D(g24545), .SI(g1979), .SE(n9390), .CLK(n9577), .Q(
        g1982), .QN(n8651) );
  SDFFX1 DFF_1123_Q_reg ( .D(g28357), .SI(g1982), .SE(n9390), .CLK(n9577), .Q(
        g1994), .QN(n8681) );
  SDFFX1 DFF_1124_Q_reg ( .D(g28362), .SI(g1994), .SE(n9390), .CLK(n9577), .Q(
        g1997), .QN(n8683) );
  SDFFX1 DFF_1125_Q_reg ( .D(g28366), .SI(g1997), .SE(n9390), .CLK(n9577), .Q(
        g2000) );
  SDFFX1 DFF_1126_Q_reg ( .D(g28352), .SI(g2000), .SE(n9390), .CLK(n9577), .Q(
        g1985), .QN(n8689) );
  SDFFX1 DFF_1127_Q_reg ( .D(g28356), .SI(g1985), .SE(n9391), .CLK(n9578), .Q(
        g1988), .QN(n8691) );
  SDFFX1 DFF_1128_Q_reg ( .D(g28361), .SI(g1988), .SE(n9391), .CLK(n9578), .Q(
        g1991) );
  SDFFX1 DFF_1129_Q_reg ( .D(g26559), .SI(g1991), .SE(n9391), .CLK(n9578), .Q(
        test_so68) );
  SDFFX1 DFF_1130_Q_reg ( .D(g26573), .SI(test_si69), .SE(n9391), .CLK(n9578), 
        .Q(g1874), .QN(n8752) );
  SDFFX1 DFF_1131_Q_reg ( .D(g26592), .SI(g1874), .SE(n9391), .CLK(n9578), .Q(
        g1877) );
  SDFFX1 DFF_1132_Q_reg ( .D(g1880), .SI(g1877), .SE(n9391), .CLK(n9578), .Q(
        g1886), .QN(n4493) );
  SDFFX1 DFF_1133_Q_reg ( .D(g22651), .SI(g1886), .SE(n9391), .CLK(n9578), .Q(
        n7968), .QN(DFF_1133_n1) );
  SDFFX1 DFF_1142_Q_reg ( .D(n548), .SI(n7968), .SE(n9391), .CLK(n9578), .Q(
        g16399), .QN(DFF_1142_n1) );
  SDFFX1 DFF_1143_Q_reg ( .D(g16399), .SI(g16399), .SE(n9391), .CLK(n9578), 
        .Q(g1905), .QN(n8993) );
  SDFFX1 DFF_1144_Q_reg ( .D(DFF_999_n1), .SI(g1905), .SE(n9391), .CLK(n9578), 
        .Q(n7967) );
  SDFFX1 DFF_1145_Q_reg ( .D(DFF_1001_n1), .SI(n7967), .SE(n9391), .CLK(n9578), 
        .Q(n7966), .QN(DFF_1145_n1) );
  SDFFX1 DFF_1146_Q_reg ( .D(DFF_1003_n1), .SI(n7966), .SE(n9391), .CLK(n9578), 
        .Q(n7965), .QN(DFF_1146_n1) );
  SDFFX1 DFF_1147_Q_reg ( .D(DFF_1005_n1), .SI(n7965), .SE(n9392), .CLK(n9579), 
        .Q(n7964) );
  SDFFX1 DFF_1148_Q_reg ( .D(DFF_1007_n1), .SI(n7964), .SE(n9392), .CLK(n9579), 
        .Q(n7963) );
  SDFFX1 DFF_1149_Q_reg ( .D(DFF_1009_n1), .SI(n7963), .SE(n9392), .CLK(n9579), 
        .Q(n7962) );
  SDFFX1 DFF_1150_Q_reg ( .D(DFF_1011_n1), .SI(n7962), .SE(n9392), .CLK(n9579), 
        .Q(g1916) );
  SDFFX1 DFF_1151_Q_reg ( .D(DFF_1013_n1), .SI(g1916), .SE(n9392), .CLK(n9579), 
        .Q(g1917) );
  SDFFX1 DFF_1152_Q_reg ( .D(g24083), .SI(g1917), .SE(n9392), .CLK(n9579), .Q(
        test_so69) );
  SDFFX1 DFF_1153_Q_reg ( .D(n4484), .SI(test_si70), .SE(n9301), .CLK(n9488), 
        .Q(n7960), .QN(n16818) );
  SDFFX1 DFF_1155_Q_reg ( .D(g7229), .SI(g7229), .SE(n9323), .CLK(n9510), .Q(
        g7357), .QN(n4357) );
  SDFFX1 DFF_1156_Q_reg ( .D(g7357), .SI(g7357), .SE(n9323), .CLK(n9510), .Q(
        g2009), .QN(n4293) );
  SDFFX1 DFF_1157_Q_reg ( .D(g16692), .SI(g2009), .SE(n9384), .CLK(n9571), .Q(
        g2010), .QN(n9032) );
  SDFFX1 DFF_1158_Q_reg ( .D(g20353), .SI(g2010), .SE(n9384), .CLK(n9571), .Q(
        g2039), .QN(n4427) );
  SDFFX1 DFF_1159_Q_reg ( .D(g20752), .SI(g2039), .SE(n9384), .CLK(n9571), .Q(
        g2020), .QN(n4400) );
  SDFFX1 DFF_1160_Q_reg ( .D(g21972), .SI(g2020), .SE(n9384), .CLK(n9571), .Q(
        g2013), .QN(n4474) );
  SDFFX1 DFF_1161_Q_reg ( .D(g23339), .SI(g2013), .SE(n9384), .CLK(n9571), .Q(
        g2033), .QN(n4420) );
  SDFFX1 DFF_1162_Q_reg ( .D(g24434), .SI(g2033), .SE(n9384), .CLK(n9571), .Q(
        g2026), .QN(n4410) );
  SDFFX1 DFF_1163_Q_reg ( .D(g25194), .SI(g2026), .SE(n9384), .CLK(n9571), .Q(
        g2040), .QN(n4399) );
  SDFFX1 DFF_1164_Q_reg ( .D(g26671), .SI(g2040), .SE(n9384), .CLK(n9571), .Q(
        g2052), .QN(n4409) );
  SDFFX1 DFF_1165_Q_reg ( .D(g26789), .SI(g2052), .SE(n9384), .CLK(n9571), .Q(
        g2046), .QN(n4468) );
  SDFFX1 DFF_1166_Q_reg ( .D(g27682), .SI(g2046), .SE(n9384), .CLK(n9571), .Q(
        g2059), .QN(n4473) );
  SDFFX1 DFF_1167_Q_reg ( .D(g27722), .SI(g2059), .SE(n9384), .CLK(n9571), .Q(
        test_so70), .QN(n9284) );
  SDFFX1 DFF_1168_Q_reg ( .D(g28325), .SI(test_si71), .SE(n9385), .CLK(n9572), 
        .Q(g2072), .QN(n4416) );
  SDFFX1 DFF_1169_Q_reg ( .D(g20899), .SI(g2072), .SE(n9392), .CLK(n9579), .Q(
        g2079) );
  SDFFX1 DFF_1170_Q_reg ( .D(g20915), .SI(g2079), .SE(n9392), .CLK(n9579), .Q(
        g2080), .QN(n9076) );
  SDFFX1 DFF_1171_Q_reg ( .D(g20934), .SI(g2080), .SE(n9392), .CLK(n9579), .Q(
        g2078) );
  SDFFX1 DFF_1172_Q_reg ( .D(g20916), .SI(g2078), .SE(n9392), .CLK(n9579), .Q(
        g2082) );
  SDFFX1 DFF_1173_Q_reg ( .D(g20935), .SI(g2082), .SE(n9392), .CLK(n9579), .Q(
        g2083), .QN(n9074) );
  SDFFX1 DFF_1174_Q_reg ( .D(g20953), .SI(g2083), .SE(n9393), .CLK(n9580), .Q(
        g2081) );
  SDFFX1 DFF_1175_Q_reg ( .D(g20936), .SI(g2081), .SE(n9393), .CLK(n9580), .Q(
        g2085) );
  SDFFX1 DFF_1176_Q_reg ( .D(g20954), .SI(g2085), .SE(n9393), .CLK(n9580), .Q(
        g2086), .QN(n9072) );
  SDFFX1 DFF_1177_Q_reg ( .D(g20977), .SI(g2086), .SE(n9393), .CLK(n9580), .Q(
        g2084) );
  SDFFX1 DFF_1178_Q_reg ( .D(g20955), .SI(g2084), .SE(n9393), .CLK(n9580), .Q(
        g2088) );
  SDFFX1 DFF_1179_Q_reg ( .D(g20978), .SI(g2088), .SE(n9393), .CLK(n9580), .Q(
        g2089), .QN(n9070) );
  SDFFX1 DFF_1180_Q_reg ( .D(g20999), .SI(g2089), .SE(n9394), .CLK(n9581), .Q(
        g2087) );
  SDFFX1 DFF_1181_Q_reg ( .D(g20979), .SI(g2087), .SE(n9394), .CLK(n9581), .Q(
        g2091) );
  SDFFX1 DFF_1182_Q_reg ( .D(g21000), .SI(g2091), .SE(n9394), .CLK(n9581), .Q(
        test_so71), .QN(n9291) );
  SDFFX1 DFF_1183_Q_reg ( .D(g21019), .SI(test_si72), .SE(n9394), .CLK(n9581), 
        .Q(g2090) );
  SDFFX1 DFF_1184_Q_reg ( .D(g21001), .SI(g2090), .SE(n9394), .CLK(n9581), .Q(
        g2094) );
  SDFFX1 DFF_1185_Q_reg ( .D(g21020), .SI(g2094), .SE(n9394), .CLK(n9581), .Q(
        g2095), .QN(n9067) );
  SDFFX1 DFF_1186_Q_reg ( .D(g21039), .SI(g2095), .SE(n9394), .CLK(n9581), .Q(
        g2093) );
  SDFFX1 DFF_1187_Q_reg ( .D(g21021), .SI(g2093), .SE(n9394), .CLK(n9581), .Q(
        g2097) );
  SDFFX1 DFF_1188_Q_reg ( .D(g21040), .SI(g2097), .SE(n9394), .CLK(n9581), .Q(
        g2098), .QN(n9065) );
  SDFFX1 DFF_1189_Q_reg ( .D(g21054), .SI(g2098), .SE(n9394), .CLK(n9581), .Q(
        g2096) );
  SDFFX1 DFF_1190_Q_reg ( .D(g21041), .SI(g2096), .SE(n9394), .CLK(n9581), .Q(
        g2100) );
  SDFFX1 DFF_1191_Q_reg ( .D(g21055), .SI(g2100), .SE(n9394), .CLK(n9581), .Q(
        g2101), .QN(n9063) );
  SDFFX1 DFF_1192_Q_reg ( .D(g21071), .SI(g2101), .SE(n9395), .CLK(n9582), .Q(
        g2099) );
  SDFFX1 DFF_1193_Q_reg ( .D(g21056), .SI(g2099), .SE(n9395), .CLK(n9582), .Q(
        g2103) );
  SDFFX1 DFF_1194_Q_reg ( .D(g21072), .SI(g2103), .SE(n9395), .CLK(n9582), .Q(
        g2104), .QN(n9061) );
  SDFFX1 DFF_1195_Q_reg ( .D(g21080), .SI(g2104), .SE(n9395), .CLK(n9582), .Q(
        g2102) );
  SDFFX1 DFF_1196_Q_reg ( .D(g20900), .SI(g2102), .SE(n9395), .CLK(n9582), .Q(
        g2106) );
  SDFFX1 DFF_1197_Q_reg ( .D(g20917), .SI(g2106), .SE(n9395), .CLK(n9582), .Q(
        test_so72), .QN(n9290) );
  SDFFX1 DFF_1198_Q_reg ( .D(g20937), .SI(test_si73), .SE(n9392), .CLK(n9579), 
        .Q(g2105) );
  SDFFX1 DFF_1199_Q_reg ( .D(g20980), .SI(g2105), .SE(n9393), .CLK(n9580), .Q(
        g2109) );
  SDFFX1 DFF_1200_Q_reg ( .D(g21002), .SI(g2109), .SE(n9393), .CLK(n9580), .Q(
        g2110) );
  SDFFX1 DFF_1201_Q_reg ( .D(g21022), .SI(g2110), .SE(n9393), .CLK(n9580), .Q(
        g2108), .QN(n8898) );
  SDFFX1 DFF_1202_Q_reg ( .D(g21003), .SI(g2108), .SE(n9393), .CLK(n9580), .Q(
        g2112) );
  SDFFX1 DFF_1203_Q_reg ( .D(g21023), .SI(g2112), .SE(n9393), .CLK(n9580), .Q(
        g2113), .QN(n8839) );
  SDFFX1 DFF_1204_Q_reg ( .D(g21042), .SI(g2113), .SE(n9393), .CLK(n9580), .Q(
        g2111) );
  SDFFX1 DFF_1205_Q_reg ( .D(g25268), .SI(g2111), .SE(n9395), .CLK(n9582), .Q(
        g2115) );
  SDFFX1 DFF_1206_Q_reg ( .D(g25271), .SI(g2115), .SE(n9395), .CLK(n9582), .Q(
        g2116) );
  SDFFX1 DFF_1207_Q_reg ( .D(g25279), .SI(g2116), .SE(n9395), .CLK(n9582), .Q(
        g2114) );
  SDFFX1 DFF_1208_Q_reg ( .D(n1194), .SI(g2114), .SE(n9395), .CLK(n9582), .Q(
        g2118), .QN(n9153) );
  SDFFX1 DFF_1209_Q_reg ( .D(g22267), .SI(g2118), .SE(n9395), .CLK(n9582), .Q(
        g2119) );
  SDFFX1 DFF_1210_Q_reg ( .D(g22280), .SI(g2119), .SE(n9395), .CLK(n9582), .Q(
        g2117), .QN(n9220) );
  SDFFX1 DFF_1211_Q_reg ( .D(g2950), .SI(g2117), .SE(n9396), .CLK(n9583), .Q(
        g6837), .QN(n4324) );
  SDFFX1 DFF_1212_Q_reg ( .D(g6837), .SI(g6837), .SE(n9396), .CLK(n9583), .Q(
        test_so73), .QN(n9278) );
  SDFFX1 DFF_1213_Q_reg ( .D(test_so73), .SI(test_si74), .SE(n9396), .CLK(
        n9583), .Q(g2241), .QN(n4367) );
  SDFFX1 DFF_1214_Q_reg ( .D(g22170), .SI(g2241), .SE(n9396), .CLK(n9583), .Q(
        g2206) );
  SDFFX1 DFF_1215_Q_reg ( .D(g22182), .SI(g2206), .SE(n9401), .CLK(n9588), .Q(
        g2207), .QN(n9169) );
  SDFFX1 DFF_1216_Q_reg ( .D(g22192), .SI(g2207), .SE(n9401), .CLK(n9588), .Q(
        g2205) );
  SDFFX1 DFF_1217_Q_reg ( .D(g22183), .SI(g2205), .SE(n9396), .CLK(n9583), .Q(
        g2209) );
  SDFFX1 DFF_1218_Q_reg ( .D(g22193), .SI(g2209), .SE(n9402), .CLK(n9589), .Q(
        g2210), .QN(n9167) );
  SDFFX1 DFF_1219_Q_reg ( .D(g22200), .SI(g2210), .SE(n9402), .CLK(n9589), .Q(
        g2208) );
  SDFFX1 DFF_1220_Q_reg ( .D(g22045), .SI(g2208), .SE(n9402), .CLK(n9589), .Q(
        g2218) );
  SDFFX1 DFF_1221_Q_reg ( .D(g22060), .SI(g2218), .SE(n9402), .CLK(n9589), .Q(
        g2219), .QN(n9165) );
  SDFFX1 DFF_1222_Q_reg ( .D(g22076), .SI(g2219), .SE(n9402), .CLK(n9589), .Q(
        g2217) );
  SDFFX1 DFF_1223_Q_reg ( .D(g22061), .SI(g2217), .SE(n9402), .CLK(n9589), .Q(
        g2221) );
  SDFFX1 DFF_1224_Q_reg ( .D(g22077), .SI(g2221), .SE(n9402), .CLK(n9589), .Q(
        g2222), .QN(n9163) );
  SDFFX1 DFF_1225_Q_reg ( .D(g22097), .SI(g2222), .SE(n9402), .CLK(n9589), .Q(
        g2220) );
  SDFFX1 DFF_1226_Q_reg ( .D(g22078), .SI(g2220), .SE(n9402), .CLK(n9589), .Q(
        g2224) );
  SDFFX1 DFF_1227_Q_reg ( .D(g22098), .SI(g2224), .SE(n9402), .CLK(n9589), .Q(
        test_so74) );
  SDFFX1 DFF_1228_Q_reg ( .D(g22115), .SI(test_si75), .SE(n9399), .CLK(n9586), 
        .Q(g2223) );
  SDFFX1 DFF_1229_Q_reg ( .D(g22099), .SI(g2223), .SE(n9399), .CLK(n9586), .Q(
        g2227) );
  SDFFX1 DFF_1230_Q_reg ( .D(g22116), .SI(g2227), .SE(n9400), .CLK(n9587), .Q(
        g2228), .QN(n9160) );
  SDFFX1 DFF_1231_Q_reg ( .D(g22138), .SI(g2228), .SE(n9400), .CLK(n9587), .Q(
        g2226) );
  SDFFX1 DFF_1232_Q_reg ( .D(g22117), .SI(g2226), .SE(n9400), .CLK(n9587), .Q(
        g2230) );
  SDFFX1 DFF_1233_Q_reg ( .D(g22139), .SI(g2230), .SE(n9401), .CLK(n9588), .Q(
        g2231), .QN(n9158) );
  SDFFX1 DFF_1234_Q_reg ( .D(g22153), .SI(g2231), .SE(n9401), .CLK(n9588), .Q(
        g2229) );
  SDFFX1 DFF_1235_Q_reg ( .D(g22140), .SI(g2229), .SE(n9401), .CLK(n9588), .Q(
        g2233) );
  SDFFX1 DFF_1236_Q_reg ( .D(g22154), .SI(g2233), .SE(n9401), .CLK(n9588), .Q(
        g2234), .QN(n9156) );
  SDFFX1 DFF_1237_Q_reg ( .D(g22171), .SI(g2234), .SE(n9401), .CLK(n9588), .Q(
        g2232) );
  SDFFX1 DFF_1238_Q_reg ( .D(g22155), .SI(g2232), .SE(n9401), .CLK(n9588), .Q(
        g2236) );
  SDFFX1 DFF_1239_Q_reg ( .D(g22172), .SI(g2236), .SE(n9401), .CLK(n9588), .Q(
        g2237), .QN(n8785) );
  SDFFX1 DFF_1240_Q_reg ( .D(g22184), .SI(g2237), .SE(n9401), .CLK(n9588), .Q(
        g2235) );
  SDFFX1 DFF_1241_Q_reg ( .D(g22173), .SI(g2235), .SE(n9401), .CLK(n9588), .Q(
        g2239), .QN(n8794) );
  SDFFX1 DFF_1242_Q_reg ( .D(g22185), .SI(g2239), .SE(n9401), .CLK(n9588), .Q(
        test_so75) );
  SDFFX1 DFF_1243_Q_reg ( .D(g22194), .SI(test_si76), .SE(n9399), .CLK(n9586), 
        .Q(g2238), .QN(n8793) );
  SDFFX1 DFF_1244_Q_reg ( .D(g25227), .SI(g2238), .SE(n9399), .CLK(n9586), .Q(
        g2245) );
  SDFFX1 DFF_1245_Q_reg ( .D(g25236), .SI(g2245), .SE(n9399), .CLK(n9586), .Q(
        g2246), .QN(n8859) );
  SDFFX1 DFF_1246_Q_reg ( .D(g25245), .SI(g2246), .SE(n9399), .CLK(n9586), .Q(
        g2244) );
  SDFFX1 DFF_1247_Q_reg ( .D(g25237), .SI(g2244), .SE(n9400), .CLK(n9587), .Q(
        g2248) );
  SDFFX1 DFF_1248_Q_reg ( .D(g25246), .SI(g2248), .SE(n9400), .CLK(n9587), .Q(
        g2249), .QN(n8856) );
  SDFFX1 DFF_1249_Q_reg ( .D(g25251), .SI(g2249), .SE(n9400), .CLK(n9587), .Q(
        g2247) );
  SDFFX1 DFF_1250_Q_reg ( .D(g25247), .SI(g2247), .SE(n9400), .CLK(n9587), .Q(
        g2251) );
  SDFFX1 DFF_1251_Q_reg ( .D(g25252), .SI(g2251), .SE(n9400), .CLK(n9587), .Q(
        g2252), .QN(n8853) );
  SDFFX1 DFF_1252_Q_reg ( .D(g25256), .SI(g2252), .SE(n9400), .CLK(n9587), .Q(
        g2250) );
  SDFFX1 DFF_1253_Q_reg ( .D(g25253), .SI(g2250), .SE(n9400), .CLK(n9587), .Q(
        g2254) );
  SDFFX1 DFF_1254_Q_reg ( .D(g25257), .SI(g2254), .SE(n9400), .CLK(n9587), .Q(
        g2255), .QN(n8850) );
  SDFFX1 DFF_1255_Q_reg ( .D(g25259), .SI(g2255), .SE(n9400), .CLK(n9587), .Q(
        g2253) );
  SDFFX1 DFF_1256_Q_reg ( .D(g30289), .SI(g2253), .SE(n9403), .CLK(n9590), .Q(
        g2261), .QN(n8441) );
  SDFFX1 DFF_1257_Q_reg ( .D(g30296), .SI(g2261), .SE(n9403), .CLK(n9590), .Q(
        test_so76) );
  SDFFX1 DFF_1258_Q_reg ( .D(g30300), .SI(test_si77), .SE(n9403), .CLK(n9590), 
        .Q(g2267), .QN(n8537) );
  SDFFX1 DFF_1259_Q_reg ( .D(g30660), .SI(g2267), .SE(n9403), .CLK(n9590), .Q(
        g2306), .QN(n8440) );
  SDFFX1 DFF_1260_Q_reg ( .D(g30666), .SI(g2306), .SE(n9403), .CLK(n9590), .Q(
        g2309) );
  SDFFX1 DFF_1261_Q_reg ( .D(g30672), .SI(g2309), .SE(n9403), .CLK(n9590), .Q(
        g2312), .QN(n8420) );
  SDFFX1 DFF_1262_Q_reg ( .D(g30690), .SI(g2312), .SE(n9403), .CLK(n9590), .Q(
        g2270), .QN(n8439) );
  SDFFX1 DFF_1263_Q_reg ( .D(g30693), .SI(g2270), .SE(n9403), .CLK(n9590), .Q(
        g2273) );
  SDFFX1 DFF_1264_Q_reg ( .D(g30695), .SI(g2273), .SE(n9403), .CLK(n9590), .Q(
        g2276), .QN(n8536) );
  SDFFX1 DFF_1265_Q_reg ( .D(g30667), .SI(g2276), .SE(n9412), .CLK(n9599), .Q(
        g2315), .QN(n8437) );
  SDFFX1 DFF_1266_Q_reg ( .D(g30673), .SI(g2315), .SE(n9412), .CLK(n9599), .Q(
        g2318) );
  SDFFX1 DFF_1267_Q_reg ( .D(g30679), .SI(g2318), .SE(n9412), .CLK(n9599), .Q(
        g2321), .QN(n8419) );
  SDFFX1 DFF_1268_Q_reg ( .D(g30301), .SI(g2321), .SE(n9412), .CLK(n9599), .Q(
        g2279), .QN(n8436) );
  SDFFX1 DFF_1269_Q_reg ( .D(g30303), .SI(g2279), .SE(n9412), .CLK(n9599), .Q(
        g2282) );
  SDFFX1 DFF_1270_Q_reg ( .D(g30304), .SI(g2282), .SE(n9396), .CLK(n9583), .Q(
        g2285), .QN(n8530) );
  SDFFX1 DFF_1271_Q_reg ( .D(g30274), .SI(g2285), .SE(n9396), .CLK(n9583), .Q(
        g2324), .QN(n8434) );
  SDFFX1 DFF_1272_Q_reg ( .D(g30282), .SI(g2324), .SE(n9396), .CLK(n9583), .Q(
        test_so77) );
  SDFFX1 DFF_1273_Q_reg ( .D(g30290), .SI(test_si78), .SE(n9396), .CLK(n9583), 
        .Q(g2330), .QN(n8418) );
  SDFFX1 DFF_1274_Q_reg ( .D(g30253), .SI(g2330), .SE(n9396), .CLK(n9583), .Q(
        g2288), .QN(n8433) );
  SDFFX1 DFF_1275_Q_reg ( .D(g30256), .SI(g2288), .SE(n9397), .CLK(n9584), .Q(
        g2291) );
  SDFFX1 DFF_1276_Q_reg ( .D(g30260), .SI(g2291), .SE(n9397), .CLK(n9584), .Q(
        g2294), .QN(n8535) );
  SDFFX1 DFF_1277_Q_reg ( .D(g30283), .SI(g2294), .SE(n9397), .CLK(n9584), .Q(
        g2333), .QN(n8431) );
  SDFFX1 DFF_1278_Q_reg ( .D(g30291), .SI(g2333), .SE(n9397), .CLK(n9584), .Q(
        g2336) );
  SDFFX1 DFF_1279_Q_reg ( .D(g30297), .SI(g2336), .SE(n9397), .CLK(n9584), .Q(
        g2339), .QN(n8527) );
  SDFFX1 DFF_1280_Q_reg ( .D(g30652), .SI(g2339), .SE(n9397), .CLK(n9584), .Q(
        g2297), .QN(n8378) );
  SDFFX1 DFF_1281_Q_reg ( .D(g30659), .SI(g2297), .SE(n9397), .CLK(n9584), .Q(
        g2300) );
  SDFFX1 DFF_1282_Q_reg ( .D(g30665), .SI(g2300), .SE(n9396), .CLK(n9583), .Q(
        g2303), .QN(n8384) );
  SDFFX1 DFF_1283_Q_reg ( .D(g30686), .SI(g2303), .SE(n9397), .CLK(n9584), .Q(
        g2342), .QN(n8377) );
  SDFFX1 DFF_1284_Q_reg ( .D(g30691), .SI(g2342), .SE(n9397), .CLK(n9584), .Q(
        g2345) );
  SDFFX1 DFF_1285_Q_reg ( .D(g30694), .SI(g2345), .SE(n9397), .CLK(n9584), .Q(
        g2348), .QN(n8376) );
  SDFFX1 DFF_1286_Q_reg ( .D(g25067), .SI(g2348), .SE(n9397), .CLK(n9584), .Q(
        g2160), .QN(n8972) );
  SDFFX1 DFF_1287_Q_reg ( .D(n53), .SI(g2160), .SE(n9397), .CLK(n9584), .Q(
        test_so78) );
  SDFFX1 DFF_1288_Q_reg ( .D(g26532), .SI(test_si79), .SE(n9398), .CLK(n9585), 
        .Q(g2151), .QN(n8971) );
  SDFFX1 DFF_1289_Q_reg ( .D(n54), .SI(g2151), .SE(n9398), .CLK(n9585), .Q(
        g2147) );
  SDFFX1 DFF_1290_Q_reg ( .D(g27621), .SI(g2147), .SE(n9398), .CLK(n9585), .Q(
        g2142), .QN(n8970) );
  SDFFX1 DFF_1291_Q_reg ( .D(g28148), .SI(g2142), .SE(n9398), .CLK(n9585), .Q(
        g2138), .QN(n9277) );
  SDFFX1 DFF_1292_Q_reg ( .D(g28637), .SI(g2138), .SE(n9398), .CLK(n9585), .Q(
        g2133), .QN(n8969) );
  SDFFX1 DFF_1293_Q_reg ( .D(g29112), .SI(g2133), .SE(n9398), .CLK(n9585), .Q(
        g2129) );
  SDFFX1 DFF_1294_Q_reg ( .D(g29357), .SI(g2129), .SE(n9398), .CLK(n9585), .Q(
        g2124), .QN(n8559) );
  SDFFX1 DFF_1295_Q_reg ( .D(g29582), .SI(g2124), .SE(n9398), .CLK(n9585), .Q(
        g2120), .QN(n8388) );
  SDFFX1 DFF_1296_Q_reg ( .D(n15), .SI(g2120), .SE(n9398), .CLK(n9585), .Q(
        g2256) );
  SDFFX1 DFF_1297_Q_reg ( .D(g2256), .SI(g2256), .SE(n9398), .CLK(n9585), .Q(
        g5637) );
  SDFFX1 DFF_1298_Q_reg ( .D(g5637), .SI(g5637), .SE(n9398), .CLK(n9585), .Q(
        g2257), .QN(n8988) );
  SDFFX1 DFF_1299_Q_reg ( .D(g2950), .SI(g2257), .SE(n9398), .CLK(n9585), .Q(
        g5555), .QN(n4516) );
  SDFFX1 DFF_1302_Q_reg ( .D(g5637), .SI(n4606), .SE(n9399), .CLK(n9586), .Q(
        test_so79), .QN(n9281) );
  SDFFX1 DFF_1303_Q_reg ( .D(g27276), .SI(test_si80), .SE(n9406), .CLK(n9593), 
        .Q(g2429) );
  SDFFX1 DFF_1304_Q_reg ( .D(g27291), .SI(g2429), .SE(n9406), .CLK(n9593), .Q(
        g2418), .QN(n8926) );
  SDFFX1 DFF_1305_Q_reg ( .D(g27307), .SI(g2418), .SE(n9406), .CLK(n9593), .Q(
        g2421) );
  SDFFX1 DFF_1306_Q_reg ( .D(g27292), .SI(g2421), .SE(n9406), .CLK(n9593), .Q(
        g2444) );
  SDFFX1 DFF_1307_Q_reg ( .D(g27308), .SI(g2444), .SE(n9406), .CLK(n9593), .Q(
        g2433), .QN(n8903) );
  SDFFX1 DFF_1308_Q_reg ( .D(g27322), .SI(g2433), .SE(n9406), .CLK(n9593), .Q(
        g2436) );
  SDFFX1 DFF_1309_Q_reg ( .D(g27309), .SI(g2436), .SE(n9406), .CLK(n9593), .Q(
        g2459) );
  SDFFX1 DFF_1310_Q_reg ( .D(g27323), .SI(g2459), .SE(n9406), .CLK(n9593), .Q(
        g2448), .QN(n8637) );
  SDFFX1 DFF_1311_Q_reg ( .D(g27334), .SI(g2448), .SE(n9406), .CLK(n9593), .Q(
        g2451) );
  SDFFX1 DFF_1312_Q_reg ( .D(g27324), .SI(g2451), .SE(n9406), .CLK(n9593), .Q(
        g2473) );
  SDFFX1 DFF_1313_Q_reg ( .D(g27335), .SI(g2473), .SE(n9406), .CLK(n9593), .Q(
        g2463), .QN(n8915) );
  SDFFX1 DFF_1314_Q_reg ( .D(g27342), .SI(g2463), .SE(n9404), .CLK(n9591), .Q(
        g2466) );
  SDFFX1 DFF_1315_Q_reg ( .D(g28763), .SI(g2466), .SE(n9404), .CLK(n9591), .Q(
        g2483) );
  SDFFX1 DFF_1316_Q_reg ( .D(g28773), .SI(g2483), .SE(n9405), .CLK(n9592), .Q(
        g2486), .QN(n8703) );
  SDFFX1 DFF_1317_Q_reg ( .D(g28782), .SI(g2486), .SE(n9405), .CLK(n9592), .Q(
        test_so80) );
  SDFFX1 DFF_1318_Q_reg ( .D(g29213), .SI(test_si81), .SE(n9404), .CLK(n9591), 
        .Q(g2492) );
  SDFFX1 DFF_1319_Q_reg ( .D(g29221), .SI(g2492), .SE(n9404), .CLK(n9591), .Q(
        g2495), .QN(n8702) );
  SDFFX1 DFF_1320_Q_reg ( .D(g29226), .SI(g2495), .SE(n9404), .CLK(n9591), .Q(
        g2498), .QN(n8715) );
  SDFFX1 DFF_1321_Q_reg ( .D(g28774), .SI(g2498), .SE(n9404), .CLK(n9591), .Q(
        g2502) );
  SDFFX1 DFF_1322_Q_reg ( .D(g28783), .SI(g2502), .SE(n9404), .CLK(n9591), .Q(
        g2503), .QN(n8938) );
  SDFFX1 DFF_1323_Q_reg ( .D(g28788), .SI(g2503), .SE(n9404), .CLK(n9591), .Q(
        g2501) );
  SDFFX1 DFF_1324_Q_reg ( .D(g26817), .SI(g2501), .SE(n9405), .CLK(n9592), .Q(
        g2504) );
  SDFFX1 DFF_1325_Q_reg ( .D(g26822), .SI(g2504), .SE(n9405), .CLK(n9592), .Q(
        g2507), .QN(n8701) );
  SDFFX1 DFF_1326_Q_reg ( .D(g26825), .SI(g2507), .SE(n9405), .CLK(n9592), .Q(
        g2510), .QN(n8713) );
  SDFFX1 DFF_1327_Q_reg ( .D(g26823), .SI(g2510), .SE(n9405), .CLK(n9592), .Q(
        g2513) );
  SDFFX1 DFF_1328_Q_reg ( .D(g26826), .SI(g2513), .SE(n9405), .CLK(n9592), .Q(
        g2516), .QN(n8700) );
  SDFFX1 DFF_1329_Q_reg ( .D(g26827), .SI(g2516), .SE(n9405), .CLK(n9592), .Q(
        g2519), .QN(n8711) );
  SDFFX1 DFF_1330_Q_reg ( .D(g27767), .SI(g2519), .SE(n9405), .CLK(n9592), .Q(
        g2523), .QN(n8946) );
  SDFFX1 DFF_1331_Q_reg ( .D(g27769), .SI(g2523), .SE(n9405), .CLK(n9592), .Q(
        g2524), .QN(n8937) );
  SDFFX1 DFF_1332_Q_reg ( .D(g27771), .SI(g2524), .SE(n9405), .CLK(n9592), .Q(
        test_so81) );
  SDFFX1 DFF_1333_Q_reg ( .D(g29618), .SI(test_si82), .SE(n9404), .CLK(n9591), 
        .Q(g2387) );
  SDFFX1 DFF_1334_Q_reg ( .D(g29621), .SI(g2387), .SE(n9404), .CLK(n9591), .Q(
        g2388), .QN(n8495) );
  SDFFX1 DFF_1335_Q_reg ( .D(g29623), .SI(g2388), .SE(n9404), .CLK(n9591), .Q(
        g2389) );
  SDFFX1 DFF_1336_Q_reg ( .D(g30707), .SI(g2389), .SE(n9404), .CLK(n9591), .Q(
        g2390) );
  SDFFX1 DFF_1337_Q_reg ( .D(g30709), .SI(g2390), .SE(n9402), .CLK(n9589), .Q(
        g2391), .QN(n8494) );
  SDFFX1 DFF_1338_Q_reg ( .D(g30566), .SI(g2391), .SE(n9402), .CLK(n9589), .Q(
        g2392) );
  SDFFX1 DFF_1339_Q_reg ( .D(g30505), .SI(g2392), .SE(n9403), .CLK(n9590), .Q(
        g2393) );
  SDFFX1 DFF_1340_Q_reg ( .D(g30341), .SI(g2393), .SE(n9403), .CLK(n9590), .Q(
        g2394), .QN(n8493) );
  SDFFX1 DFF_1341_Q_reg ( .D(g30356), .SI(g2394), .SE(n9403), .CLK(n9590), .Q(
        g2395) );
  SDFFX1 DFF_1342_Q_reg ( .D(g29182), .SI(g2395), .SE(n9412), .CLK(n9599), .Q(
        g2397) );
  SDFFX1 DFF_1343_Q_reg ( .D(g29185), .SI(g2397), .SE(n9412), .CLK(n9599), .Q(
        g2398), .QN(n8547) );
  SDFFX1 DFF_1344_Q_reg ( .D(g29187), .SI(g2398), .SE(n9396), .CLK(n9583), .Q(
        g2396) );
  SDFFX1 DFF_1345_Q_reg ( .D(g26672), .SI(g2396), .SE(n9399), .CLK(n9586), .Q(
        g2478) );
  SDFFX1 DFF_1346_Q_reg ( .D(g26676), .SI(g2478), .SE(n9399), .CLK(n9586), .Q(
        g2479), .QN(n8936) );
  SDFFX1 DFF_1347_Q_reg ( .D(g26025), .SI(g2479), .SE(n9399), .CLK(n9586), .Q(
        test_so82) );
  SDFFX1 DFF_1348_Q_reg ( .D(n4287), .SI(test_si83), .SE(n9305), .CLK(n9492), 
        .Q(g2525) );
  SDFFX1 DFF_1349_Q_reg ( .D(g2525), .SI(g2525), .SE(n9305), .CLK(n9492), .Q(
        n7946), .QN(DFF_1349_n1) );
  SDFFX1 DFF_1350_Q_reg ( .D(n4563), .SI(n7946), .SE(n9305), .CLK(n9492), .Q(
        g2527) );
  SDFFX1 DFF_1351_Q_reg ( .D(g2527), .SI(g2527), .SE(n9305), .CLK(n9492), .Q(
        n7945), .QN(DFF_1351_n1) );
  SDFFX1 DFF_1352_Q_reg ( .D(n4555), .SI(n7945), .SE(n9305), .CLK(n9492), .Q(
        g2529) );
  SDFFX1 DFF_1353_Q_reg ( .D(g2529), .SI(g2529), .SE(n9305), .CLK(n9492), .Q(
        n7944), .QN(DFF_1353_n1) );
  SDFFX1 DFF_1354_Q_reg ( .D(n4325), .SI(n7944), .SE(n9305), .CLK(n9492), .Q(
        g2355) );
  SDFFX1 DFF_1355_Q_reg ( .D(g2355), .SI(g2355), .SE(n9306), .CLK(n9493), .Q(
        n7943), .QN(DFF_1355_n1) );
  SDFFX1 DFF_1356_Q_reg ( .D(n4389), .SI(n7943), .SE(n9306), .CLK(n9493), .Q(
        g2357) );
  SDFFX1 DFF_1357_Q_reg ( .D(g2357), .SI(g2357), .SE(n9306), .CLK(n9493), .Q(
        n7942), .QN(DFF_1357_n1) );
  SDFFX1 DFF_1358_Q_reg ( .D(n4319), .SI(n7942), .SE(n9306), .CLK(n9493), .Q(
        g2359) );
  SDFFX1 DFF_1359_Q_reg ( .D(g2359), .SI(g2359), .SE(n9306), .CLK(n9493), .Q(
        n7941), .QN(DFF_1359_n1) );
  SDFFX1 DFF_1360_Q_reg ( .D(n4373), .SI(n7941), .SE(n9306), .CLK(n9493), .Q(
        g2361) );
  SDFFX1 DFF_1361_Q_reg ( .D(g2361), .SI(g2361), .SE(n9306), .CLK(n9493), .Q(
        n7940), .QN(DFF_1361_n1) );
  SDFFX1 DFF_1362_Q_reg ( .D(n4377), .SI(n7940), .SE(n9306), .CLK(n9493), .Q(
        test_so83) );
  SDFFX1 DFF_1363_Q_reg ( .D(test_so83), .SI(test_si84), .SE(n9306), .CLK(
        n9493), .Q(n7938), .QN(DFF_1363_n1) );
  SDFFX1 DFF_1364_Q_reg ( .D(g2878), .SI(n7938), .SE(n9321), .CLK(n9508), .Q(
        g2365) );
  SDFFX1 DFF_1365_Q_reg ( .D(g2365), .SI(g2365), .SE(n9322), .CLK(n9509), .Q(
        n7937), .QN(n4483) );
  SDFFX1 DFF_1366_Q_reg ( .D(n4285), .SI(n7937), .SE(n9405), .CLK(n9592), .Q(
        g2374), .QN(n4487) );
  SDFFX1 DFF_1367_Q_reg ( .D(g30055), .SI(g2374), .SE(n9415), .CLK(n9602), .Q(
        g2380) );
  SDFFX1 DFF_1378_Q_reg ( .D(n4275), .SI(g2380), .SE(n9412), .CLK(n9599), .Q(
        n7936), .QN(DFF_1378_n1) );
  SDFFX1 DFF_1379_Q_reg ( .D(g2429), .SI(n7936), .SE(n9412), .CLK(n9599), .Q(
        g2417) );
  SDFFX1 DFF_1380_Q_reg ( .D(g2417), .SI(g2417), .SE(n9413), .CLK(n9600), .Q(
        g2424), .QN(n16820) );
  SDFFX1 DFF_1381_Q_reg ( .D(g2418), .SI(g2424), .SE(n9413), .CLK(n9600), .Q(
        g2425) );
  SDFFX1 DFF_1382_Q_reg ( .D(g2425), .SI(g2425), .SE(n9413), .CLK(n9600), .Q(
        g2426) );
  SDFFX1 DFF_1383_Q_reg ( .D(g2421), .SI(g2426), .SE(n9413), .CLK(n9600), .Q(
        g2427) );
  SDFFX1 DFF_1384_Q_reg ( .D(g2427), .SI(g2427), .SE(n9413), .CLK(n9600), .Q(
        g2428), .QN(n8612) );
  SDFFX1 DFF_1385_Q_reg ( .D(g2444), .SI(g2428), .SE(n9413), .CLK(n9600), .Q(
        g2432) );
  SDFFX1 DFF_1386_Q_reg ( .D(g2432), .SI(g2432), .SE(n9413), .CLK(n9600), .Q(
        g2439) );
  SDFFX1 DFF_1387_Q_reg ( .D(g2433), .SI(g2439), .SE(n9413), .CLK(n9600), .Q(
        test_so84) );
  SDFFX1 DFF_1388_Q_reg ( .D(test_so84), .SI(test_si85), .SE(n9413), .CLK(
        n9600), .Q(g2441), .QN(n8403) );
  SDFFX1 DFF_1389_Q_reg ( .D(g2436), .SI(g2441), .SE(n9413), .CLK(n9600), .Q(
        g2442) );
  SDFFX1 DFF_1390_Q_reg ( .D(g2442), .SI(g2442), .SE(n9413), .CLK(n9600), .Q(
        g2443), .QN(n8402) );
  SDFFX1 DFF_1391_Q_reg ( .D(g2459), .SI(g2443), .SE(n9413), .CLK(n9600), .Q(
        g2447) );
  SDFFX1 DFF_1392_Q_reg ( .D(g2447), .SI(g2447), .SE(n9414), .CLK(n9601), .Q(
        g2454) );
  SDFFX1 DFF_1393_Q_reg ( .D(g2448), .SI(g2454), .SE(n9414), .CLK(n9601), .Q(
        g2455) );
  SDFFX1 DFF_1394_Q_reg ( .D(g2455), .SI(g2455), .SE(n9414), .CLK(n9601), .Q(
        g2456), .QN(n8577) );
  SDFFX1 DFF_1395_Q_reg ( .D(g2451), .SI(g2456), .SE(n9414), .CLK(n9601), .Q(
        g2457) );
  SDFFX1 DFF_1396_Q_reg ( .D(g2457), .SI(g2457), .SE(n9414), .CLK(n9601), .Q(
        g2458), .QN(n8576) );
  SDFFX1 DFF_1397_Q_reg ( .D(g2473), .SI(g2458), .SE(n9414), .CLK(n9601), .Q(
        g2462) );
  SDFFX1 DFF_1398_Q_reg ( .D(g2462), .SI(g2462), .SE(n9414), .CLK(n9601), .Q(
        g2469), .QN(n16821) );
  SDFFX1 DFF_1399_Q_reg ( .D(g2463), .SI(g2469), .SE(n9414), .CLK(n9601), .Q(
        g2470) );
  SDFFX1 DFF_1400_Q_reg ( .D(g2470), .SI(g2470), .SE(n9414), .CLK(n9601), .Q(
        g2471), .QN(n8411) );
  SDFFX1 DFF_1401_Q_reg ( .D(g2466), .SI(g2471), .SE(n9414), .CLK(n9601), .Q(
        g2472) );
  SDFFX1 DFF_1402_Q_reg ( .D(g2472), .SI(g2472), .SE(n9414), .CLK(n9601), .Q(
        test_so85) );
  SDFFX1 DFF_1403_Q_reg ( .D(n4598), .SI(test_si86), .SE(n9328), .CLK(n9515), 
        .Q(g5747), .QN(n8610) );
  SDFFX1 DFF_1404_Q_reg ( .D(g5747), .SI(g5747), .SE(n9329), .CLK(n9516), .Q(
        g5796), .QN(n8613) );
  SDFFX1 DFF_1405_Q_reg ( .D(g5796), .SI(g5796), .SE(n9329), .CLK(n9516), .Q(
        g2412), .QN(n8611) );
  SDFFX1 DFF_1406_Q_reg ( .D(n4598), .SI(g2412), .SE(n9329), .CLK(n9516), .Q(
        g7302), .QN(n4314) );
  SDFFX1 DFF_1407_Q_reg ( .D(g7302), .SI(g7302), .SE(n9329), .CLK(n9516), .Q(
        g7390), .QN(n4370) );
  SDFFX1 DFF_1408_Q_reg ( .D(g7390), .SI(g7390), .SE(n9329), .CLK(n9516), .Q(
        g2624), .QN(n4299) );
  SDFFX1 DFF_1409_Q_reg ( .D(n1464), .SI(g2624), .SE(n9329), .CLK(n9516), .Q(
        g2628), .QN(n9223) );
  SDFFX1 DFF_1410_Q_reg ( .D(g18780), .SI(g2628), .SE(n9329), .CLK(n9516), .Q(
        g2631), .QN(n4352) );
  SDFFX1 DFF_1411_Q_reg ( .D(g18820), .SI(g2631), .SE(n9329), .CLK(n9516), .Q(
        g2584), .QN(n4303) );
  SDFFX1 DFF_1412_Q_reg ( .D(n1457), .SI(g2584), .SE(n9409), .CLK(n9596), .Q(
        g2587) );
  SDFFX1 DFF_1413_Q_reg ( .D(g2587), .SI(g2587), .SE(n9409), .CLK(n9596), .Q(
        g2597) );
  SDFFX1 DFF_1414_Q_reg ( .D(g2597), .SI(g2597), .SE(n9409), .CLK(n9596), .Q(
        g2598) );
  SDFFX1 DFF_1415_Q_reg ( .D(g2530), .SI(g2598), .SE(n9408), .CLK(n9595), .Q(
        g2638) );
  SDFFX1 DFF_1416_Q_reg ( .D(g2638), .SI(g2638), .SE(n9408), .CLK(n9595), .Q(
        g2643), .QN(n8770) );
  SDFFX1 DFF_1417_Q_reg ( .D(g2533), .SI(g2643), .SE(n9408), .CLK(n9595), .Q(
        test_so86) );
  SDFFX1 DFF_1418_Q_reg ( .D(test_so86), .SI(test_si87), .SE(n9409), .CLK(
        n9596), .Q(g2645) );
  SDFFX1 DFF_1419_Q_reg ( .D(g2536), .SI(g2645), .SE(n9409), .CLK(n9596), .Q(
        g2646) );
  SDFFX1 DFF_1420_Q_reg ( .D(g2646), .SI(g2646), .SE(n9409), .CLK(n9596), .Q(
        g2647), .QN(n8771) );
  SDFFX1 DFF_1421_Q_reg ( .D(g2540), .SI(g2647), .SE(n9407), .CLK(n9594), .Q(
        g2648) );
  SDFFX1 DFF_1422_Q_reg ( .D(g2648), .SI(g2648), .SE(n9407), .CLK(n9594), .Q(
        g2639), .QN(n8768) );
  SDFFX1 DFF_1423_Q_reg ( .D(g2543), .SI(g2639), .SE(n9407), .CLK(n9594), .Q(
        g2640) );
  SDFFX1 DFF_1424_Q_reg ( .D(g2640), .SI(g2640), .SE(n9407), .CLK(n9594), .Q(
        g2641) );
  SDFFX1 DFF_1425_Q_reg ( .D(g2546), .SI(g2641), .SE(n9407), .CLK(n9594), .Q(
        g2642) );
  SDFFX1 DFF_1426_Q_reg ( .D(g2642), .SI(g2642), .SE(n9407), .CLK(n9594), .Q(
        g2564), .QN(n8769) );
  SDFFX1 DFF_1427_Q_reg ( .D(g2950), .SI(g2564), .SE(n9407), .CLK(n9594), .Q(
        g8087), .QN(n4456) );
  SDFFX1 DFF_1428_Q_reg ( .D(g8087), .SI(g8087), .SE(n9407), .CLK(n9594), .Q(
        g8167), .QN(n4455) );
  SDFFX1 DFF_1429_Q_reg ( .D(g8167), .SI(g8167), .SE(n9408), .CLK(n9595), .Q(
        g2560), .QN(n4463) );
  SDFFX1 DFF_1430_Q_reg ( .D(g23114), .SI(g2560), .SE(n9408), .CLK(n9595), .Q(
        g2561), .QN(n8996) );
  SDFFX1 DFF_1431_Q_reg ( .D(g23133), .SI(g2561), .SE(n9408), .CLK(n9595), .Q(
        g2562) );
  SDFFX1 DFF_1432_Q_reg ( .D(g21970), .SI(g2562), .SE(n9408), .CLK(n9595), .Q(
        test_so87) );
  SDFFX1 DFF_1433_Q_reg ( .D(g23407), .SI(test_si88), .SE(n9408), .CLK(n9595), 
        .Q(g2530) );
  SDFFX1 DFF_1434_Q_reg ( .D(g23418), .SI(g2530), .SE(n9408), .CLK(n9595), .Q(
        g2533) );
  SDFFX1 DFF_1435_Q_reg ( .D(g24209), .SI(g2533), .SE(n9408), .CLK(n9595), .Q(
        g2536) );
  SDFFX1 DFF_1436_Q_reg ( .D(g24214), .SI(g2536), .SE(n9409), .CLK(n9596), .Q(
        g2552), .QN(n9001) );
  SDFFX1 DFF_1437_Q_reg ( .D(g24226), .SI(g2552), .SE(n9409), .CLK(n9596), .Q(
        g2553) );
  SDFFX1 DFF_1438_Q_reg ( .D(g24238), .SI(g2553), .SE(n9406), .CLK(n9593), .Q(
        g2554), .QN(n9002) );
  SDFFX1 DFF_1439_Q_reg ( .D(g23132), .SI(g2554), .SE(n9407), .CLK(n9594), .Q(
        g2555), .QN(n8998) );
  SDFFX1 DFF_1440_Q_reg ( .D(g23047), .SI(g2555), .SE(n9407), .CLK(n9594), .Q(
        g2559) );
  SDFFX1 DFF_1441_Q_reg ( .D(g23076), .SI(g2559), .SE(n9407), .CLK(n9594), .Q(
        g2539), .QN(n8999) );
  SDFFX1 DFF_1442_Q_reg ( .D(g24225), .SI(g2539), .SE(n9407), .CLK(n9594), .Q(
        g2540) );
  SDFFX1 DFF_1443_Q_reg ( .D(g24237), .SI(g2540), .SE(n9408), .CLK(n9595), .Q(
        g2543) );
  SDFFX1 DFF_1444_Q_reg ( .D(g24250), .SI(g2543), .SE(n9408), .CLK(n9595), .Q(
        g2546) );
  SDFFX1 DFF_1445_Q_reg ( .D(n1456), .SI(g2546), .SE(n9409), .CLK(n9596), .Q(
        g2602) );
  SDFFX1 DFF_1446_Q_reg ( .D(g2602), .SI(g2602), .SE(n9409), .CLK(n9596), .Q(
        g2609) );
  SDFFX1 DFF_1447_Q_reg ( .D(g2609), .SI(g2609), .SE(n9409), .CLK(n9596), .Q(
        test_so88), .QN(n8647) );
  SDFFX1 DFF_1448_Q_reg ( .D(g13175), .SI(test_si89), .SE(n9409), .CLK(n9596), 
        .Q(g2617) );
  SDFFX1 DFF_1449_Q_reg ( .D(g2617), .SI(g2617), .SE(n9410), .CLK(n9597), .Q(
        n7930) );
  SDFFX1 DFF_1450_Q_reg ( .D(g30072), .SI(n7930), .SE(n9410), .CLK(n9597), .Q(
        n7929) );
  SDFFX1 DFF_1451_Q_reg ( .D(g13143), .SI(n7929), .SE(n9410), .CLK(n9597), .Q(
        g2623) );
  SDFFX1 DFF_1452_Q_reg ( .D(g2623), .SI(g2623), .SE(n9410), .CLK(n9597), .Q(
        g2574), .QN(n4543) );
  SDFFX1 DFF_1453_Q_reg ( .D(g13194), .SI(g2574), .SE(n9410), .CLK(n9597), .Q(
        g2632) );
  SDFFX1 DFF_1454_Q_reg ( .D(g2632), .SI(g2632), .SE(n9410), .CLK(n9597), .Q(
        g2633), .QN(n9035) );
  SDFFX1 DFF_1455_Q_reg ( .D(g27310), .SI(g2633), .SE(n9410), .CLK(n9597), .Q(
        g2650) );
  SDFFX1 DFF_1456_Q_reg ( .D(g27325), .SI(g2650), .SE(n9411), .CLK(n9598), .Q(
        g2651), .QN(n8566) );
  SDFFX1 DFF_1457_Q_reg ( .D(g27336), .SI(g2651), .SE(n9412), .CLK(n9599), .Q(
        g2649) );
  SDFFX1 DFF_1458_Q_reg ( .D(g27326), .SI(g2649), .SE(n9412), .CLK(n9599), .Q(
        g2653) );
  SDFFX1 DFF_1459_Q_reg ( .D(g27337), .SI(g2653), .SE(n9412), .CLK(n9599), .Q(
        g2654), .QN(n8586) );
  SDFFX1 DFF_1460_Q_reg ( .D(g27343), .SI(g2654), .SE(n9410), .CLK(n9597), .Q(
        g2652) );
  SDFFX1 DFF_1461_Q_reg ( .D(g27338), .SI(g2652), .SE(n9410), .CLK(n9597), .Q(
        g2656) );
  SDFFX1 DFF_1462_Q_reg ( .D(g27344), .SI(g2656), .SE(n9410), .CLK(n9597), .Q(
        test_so89) );
  SDFFX1 DFF_1463_Q_reg ( .D(g27347), .SI(test_si90), .SE(n9410), .CLK(n9597), 
        .Q(g2655) );
  SDFFX1 DFF_1464_Q_reg ( .D(g27345), .SI(g2655), .SE(n9411), .CLK(n9598), .Q(
        g2659) );
  SDFFX1 DFF_1465_Q_reg ( .D(g27348), .SI(g2659), .SE(n9411), .CLK(n9598), .Q(
        g2660), .QN(n8601) );
  SDFFX1 DFF_1466_Q_reg ( .D(g27354), .SI(g2660), .SE(n9411), .CLK(n9598), .Q(
        g2658) );
  SDFFX1 DFF_1467_Q_reg ( .D(g24527), .SI(g2658), .SE(n9411), .CLK(n9598), .Q(
        g2661), .QN(n8660) );
  SDFFX1 DFF_1468_Q_reg ( .D(g24537), .SI(g2661), .SE(n9411), .CLK(n9598), .Q(
        g2664), .QN(n8662) );
  SDFFX1 DFF_1469_Q_reg ( .D(g24547), .SI(g2664), .SE(n9411), .CLK(n9598), .Q(
        g2667), .QN(n8661) );
  SDFFX1 DFF_1470_Q_reg ( .D(g24538), .SI(g2667), .SE(n9411), .CLK(n9598), .Q(
        g2670), .QN(n8646) );
  SDFFX1 DFF_1471_Q_reg ( .D(g24548), .SI(g2670), .SE(n9411), .CLK(n9598), .Q(
        g2673), .QN(n8649) );
  SDFFX1 DFF_1472_Q_reg ( .D(g24557), .SI(g2673), .SE(n9411), .CLK(n9598), .Q(
        g2676), .QN(n8648) );
  SDFFX1 DFF_1473_Q_reg ( .D(g28364), .SI(g2676), .SE(n9411), .CLK(n9598), .Q(
        g2688), .QN(n8678) );
  SDFFX1 DFF_1474_Q_reg ( .D(g28368), .SI(g2688), .SE(n9411), .CLK(n9598), .Q(
        g2691) );
  SDFFX1 DFF_1475_Q_reg ( .D(g28371), .SI(g2691), .SE(n9322), .CLK(n9509), .Q(
        g2694), .QN(n8679) );
  SDFFX1 DFF_1476_Q_reg ( .D(g28358), .SI(g2694), .SE(n9414), .CLK(n9601), .Q(
        g2679), .QN(n8687) );
  SDFFX1 DFF_1477_Q_reg ( .D(g28363), .SI(g2679), .SE(n9415), .CLK(n9602), .Q(
        test_so90) );
  SDFFX1 DFF_1478_Q_reg ( .D(g28367), .SI(test_si91), .SE(n9415), .CLK(n9602), 
        .Q(g2685), .QN(n8688) );
  SDFFX1 DFF_1479_Q_reg ( .D(g26575), .SI(g2685), .SE(n9415), .CLK(n9602), .Q(
        g2565), .QN(n8745) );
  SDFFX1 DFF_1480_Q_reg ( .D(g26596), .SI(g2565), .SE(n9415), .CLK(n9602), .Q(
        g2568) );
  SDFFX1 DFF_1481_Q_reg ( .D(g26616), .SI(g2568), .SE(n9322), .CLK(n9509), .Q(
        g2571), .QN(n8747) );
  SDFFX1 DFF_1482_Q_reg ( .D(g2574), .SI(g2571), .SE(n9410), .CLK(n9597), .Q(
        g2580), .QN(n8755) );
  SDFFX1 DFF_1483_Q_reg ( .D(g22687), .SI(g2580), .SE(n9322), .CLK(n9509), .Q(
        n7926) );
  SDFFX1 DFF_1492_Q_reg ( .D(g30061), .SI(n7926), .SE(n9322), .CLK(n9509), .Q(
        g16437) );
  SDFFX1 DFF_1493_Q_reg ( .D(g16437), .SI(g16437), .SE(n9322), .CLK(n9509), 
        .Q(g2599), .QN(n8992) );
  SDFFX1 DFF_1494_Q_reg ( .D(DFF_1349_n1), .SI(g2599), .SE(n9322), .CLK(n9509), 
        .Q(n7925) );
  SDFFX1 DFF_1495_Q_reg ( .D(DFF_1351_n1), .SI(n7925), .SE(n9322), .CLK(n9509), 
        .Q(n7924), .QN(DFF_1495_n1) );
  SDFFX1 DFF_1496_Q_reg ( .D(DFF_1353_n1), .SI(n7924), .SE(n9322), .CLK(n9509), 
        .Q(n7923), .QN(DFF_1496_n1) );
  SDFFX1 DFF_1497_Q_reg ( .D(DFF_1355_n1), .SI(n7923), .SE(n9323), .CLK(n9510), 
        .Q(n7922) );
  SDFFX1 DFF_1498_Q_reg ( .D(DFF_1357_n1), .SI(n7922), .SE(n9323), .CLK(n9510), 
        .Q(n7921) );
  SDFFX1 DFF_1499_Q_reg ( .D(DFF_1359_n1), .SI(n7921), .SE(n9323), .CLK(n9510), 
        .Q(n7920) );
  SDFFX1 DFF_1500_Q_reg ( .D(DFF_1361_n1), .SI(n7920), .SE(n9323), .CLK(n9510), 
        .Q(test_so91) );
  SDFFX1 DFF_1501_Q_reg ( .D(DFF_1363_n1), .SI(test_si92), .SE(n9306), .CLK(
        n9493), .Q(g2611) );
  SDFFX1 DFF_1502_Q_reg ( .D(g24092), .SI(g2611), .SE(n9415), .CLK(n9602), .Q(
        g2612), .QN(n4490) );
  SDFFX1 DFF_1503_Q_reg ( .D(n4483), .SI(g2612), .SE(n9322), .CLK(n9509), .Q(
        n7918), .QN(n16817) );
  SDFFX1 DFF_1505_Q_reg ( .D(g7425), .SI(g7425), .SE(n9329), .CLK(n9516), .Q(
        g7487), .QN(n4356) );
  SDFFX1 DFF_1506_Q_reg ( .D(g7487), .SI(g7487), .SE(n9329), .CLK(n9516), .Q(
        g2703), .QN(n4292) );
  SDFFX1 DFF_1507_Q_reg ( .D(g16718), .SI(g2703), .SE(n9329), .CLK(n9516), .Q(
        g2704), .QN(n9031) );
  SDFFX1 DFF_1508_Q_reg ( .D(g20375), .SI(g2704), .SE(n9354), .CLK(n9541), .Q(
        g2733) );
  SDFFX1 DFF_1509_Q_reg ( .D(g20789), .SI(g2733), .SE(n9354), .CLK(n9541), .Q(
        g2714), .QN(n4398) );
  SDFFX1 DFF_1510_Q_reg ( .D(g21974), .SI(g2714), .SE(n9354), .CLK(n9541), .Q(
        g2707), .QN(n4472) );
  SDFFX1 DFF_1511_Q_reg ( .D(g23348), .SI(g2707), .SE(n9354), .CLK(n9541), .Q(
        g2727), .QN(n4419) );
  SDFFX1 DFF_1512_Q_reg ( .D(g24438), .SI(g2727), .SE(n9354), .CLK(n9541), .Q(
        g2720), .QN(n4408) );
  SDFFX1 DFF_1513_Q_reg ( .D(g25197), .SI(g2720), .SE(n9354), .CLK(n9541), .Q(
        g2734), .QN(n4397) );
  SDFFX1 DFF_1514_Q_reg ( .D(g26677), .SI(g2734), .SE(n9354), .CLK(n9541), .Q(
        g2746), .QN(n4407) );
  SDFFX1 DFF_1515_Q_reg ( .D(g26795), .SI(g2746), .SE(n9354), .CLK(n9541), .Q(
        test_so92), .QN(n9282) );
  SDFFX1 DFF_1516_Q_reg ( .D(g27243), .SI(test_si93), .SE(n9354), .CLK(n9541), 
        .Q(g2753), .QN(n4471) );
  SDFFX1 DFF_1517_Q_reg ( .D(n1524), .SI(g2753), .SE(n9354), .CLK(n9541), .Q(
        g2760), .QN(n4393) );
  SDFFX1 DFF_1518_Q_reg ( .D(g28328), .SI(g2760), .SE(n9354), .CLK(n9541), .Q(
        g2766), .QN(n4415) );
  SDFFX1 DFF_1519_Q_reg ( .D(g20918), .SI(g2766), .SE(n9354), .CLK(n9541), .Q(
        g2773) );
  SDFFX1 DFF_1520_Q_reg ( .D(g20939), .SI(g2773), .SE(n9355), .CLK(n9542), .Q(
        g2774), .QN(n9058) );
  SDFFX1 DFF_1521_Q_reg ( .D(g20962), .SI(g2774), .SE(n9355), .CLK(n9542), .Q(
        g2772) );
  SDFFX1 DFF_1522_Q_reg ( .D(g20940), .SI(g2772), .SE(n9355), .CLK(n9542), .Q(
        g2776) );
  SDFFX1 DFF_1523_Q_reg ( .D(g20963), .SI(g2776), .SE(n9355), .CLK(n9542), .Q(
        g2777), .QN(n9056) );
  SDFFX1 DFF_1524_Q_reg ( .D(g20981), .SI(g2777), .SE(n9355), .CLK(n9542), .Q(
        g2775) );
  SDFFX1 DFF_1525_Q_reg ( .D(g20964), .SI(g2775), .SE(n9356), .CLK(n9543), .Q(
        g2779) );
  SDFFX1 DFF_1526_Q_reg ( .D(g20982), .SI(g2779), .SE(n9356), .CLK(n9543), .Q(
        g2780), .QN(n9054) );
  SDFFX1 DFF_1527_Q_reg ( .D(g21004), .SI(g2780), .SE(n9356), .CLK(n9543), .Q(
        g2778) );
  SDFFX1 DFF_1528_Q_reg ( .D(g20983), .SI(g2778), .SE(n9356), .CLK(n9543), .Q(
        g2782) );
  SDFFX1 DFF_1529_Q_reg ( .D(g21005), .SI(g2782), .SE(n9356), .CLK(n9543), .Q(
        g2783), .QN(n9052) );
  SDFFX1 DFF_1530_Q_reg ( .D(g21025), .SI(g2783), .SE(n9356), .CLK(n9543), .Q(
        test_so93) );
  SDFFX1 DFF_1531_Q_reg ( .D(g21006), .SI(test_si94), .SE(n9355), .CLK(n9542), 
        .Q(g2785) );
  SDFFX1 DFF_1532_Q_reg ( .D(g21026), .SI(g2785), .SE(n9356), .CLK(n9543), .Q(
        g2786), .QN(n9050) );
  SDFFX1 DFF_1533_Q_reg ( .D(g21043), .SI(g2786), .SE(n9356), .CLK(n9543), .Q(
        g2784) );
  SDFFX1 DFF_1534_Q_reg ( .D(g21027), .SI(g2784), .SE(n9356), .CLK(n9543), .Q(
        g2788) );
  SDFFX1 DFF_1535_Q_reg ( .D(g21044), .SI(g2788), .SE(n9356), .CLK(n9543), .Q(
        g2789), .QN(n9048) );
  SDFFX1 DFF_1536_Q_reg ( .D(g21060), .SI(g2789), .SE(n9356), .CLK(n9543), .Q(
        g2787) );
  SDFFX1 DFF_1537_Q_reg ( .D(g21045), .SI(g2787), .SE(n9356), .CLK(n9543), .Q(
        g2791) );
  SDFFX1 DFF_1538_Q_reg ( .D(g21061), .SI(g2791), .SE(n9357), .CLK(n9544), .Q(
        g2792), .QN(n9046) );
  SDFFX1 DFF_1539_Q_reg ( .D(g21073), .SI(g2792), .SE(n9357), .CLK(n9544), .Q(
        g2790) );
  SDFFX1 DFF_1540_Q_reg ( .D(g21062), .SI(g2790), .SE(n9357), .CLK(n9544), .Q(
        g2794) );
  SDFFX1 DFF_1541_Q_reg ( .D(g21074), .SI(g2794), .SE(n9357), .CLK(n9544), .Q(
        g2795), .QN(n9044) );
  SDFFX1 DFF_1542_Q_reg ( .D(g21081), .SI(g2795), .SE(n9357), .CLK(n9544), .Q(
        g2793) );
  SDFFX1 DFF_1543_Q_reg ( .D(g21075), .SI(g2793), .SE(n9357), .CLK(n9544), .Q(
        g2797) );
  SDFFX1 DFF_1544_Q_reg ( .D(g21082), .SI(g2797), .SE(n9357), .CLK(n9544), .Q(
        g2798), .QN(n9042) );
  SDFFX1 DFF_1545_Q_reg ( .D(g21094), .SI(g2798), .SE(n9357), .CLK(n9544), .Q(
        test_so94) );
  SDFFX1 DFF_1546_Q_reg ( .D(g20919), .SI(test_si95), .SE(n9355), .CLK(n9542), 
        .Q(g2800) );
  SDFFX1 DFF_1547_Q_reg ( .D(g20941), .SI(g2800), .SE(n9355), .CLK(n9542), .Q(
        g2801), .QN(n9040) );
  SDFFX1 DFF_1548_Q_reg ( .D(g20965), .SI(g2801), .SE(n9355), .CLK(n9542), .Q(
        g2799) );
  SDFFX1 DFF_1549_Q_reg ( .D(g21007), .SI(g2799), .SE(n9355), .CLK(n9542), .Q(
        g2803) );
  SDFFX1 DFF_1550_Q_reg ( .D(g21028), .SI(g2803), .SE(n9355), .CLK(n9542), .Q(
        g2804) );
  SDFFX1 DFF_1551_Q_reg ( .D(g21046), .SI(g2804), .SE(n9355), .CLK(n9542), .Q(
        g2802), .QN(n8896) );
  SDFFX1 DFF_1552_Q_reg ( .D(g21029), .SI(g2802), .SE(n9415), .CLK(n9602), .Q(
        g2806) );
  SDFFX1 DFF_1553_Q_reg ( .D(g21047), .SI(g2806), .SE(n9415), .CLK(n9602), .Q(
        g2807), .QN(n8837) );
  SDFFX1 DFF_1554_Q_reg ( .D(g21063), .SI(g2807), .SE(n9415), .CLK(n9602), .Q(
        g2805) );
  SDFFX1 DFF_1555_Q_reg ( .D(g25272), .SI(g2805), .SE(n9415), .CLK(n9602), .Q(
        g2809) );
  SDFFX1 DFF_1556_Q_reg ( .D(g25280), .SI(g2809), .SE(n9415), .CLK(n9602), .Q(
        g2810) );
  SDFFX1 DFF_1557_Q_reg ( .D(g25288), .SI(g2810), .SE(n9323), .CLK(n9510), .Q(
        g2808) );
  SDFFX1 DFF_1558_Q_reg ( .D(n1499), .SI(g2808), .SE(n9323), .CLK(n9510), .Q(
        g2812), .QN(n9152) );
  SDFFX1 DFF_1559_Q_reg ( .D(g22284), .SI(g2812), .SE(n9357), .CLK(n9544), .Q(
        g2813) );
  SDFFX1 DFF_1560_Q_reg ( .D(g22299), .SI(g2813), .SE(n9357), .CLK(n9544), .Q(
        test_so95) );
  SDFFX1 DFF_1561_Q_reg ( .D(g20877), .SI(test_si96), .SE(n9323), .CLK(n9510), 
        .Q(n7913), .QN(DFF_1561_n1) );
  SDFFX1 DFF_1562_Q_reg ( .D(g20884), .SI(n7913), .SE(n9323), .CLK(n9510), .Q(
        n7912), .QN(DFF_1562_n1) );
  SDFFX1 DFF_1563_Q_reg ( .D(n4263_Tj_Payload), .SI(n7912), .SE(n9323), .CLK(
        n9510), .Q(n4598), .QN(n9260) );
  SDFFX1 DFF_1564_Q_reg ( .D(n4269), .SI(n4598), .SE(n9297), .CLK(n9484), .Q(
        g3043) );
  SDFFX1 DFF_1565_Q_reg ( .D(n4268), .SI(g3043), .SE(n9297), .CLK(n9484), .Q(
        g3044) );
  SDFFX1 DFF_1566_Q_reg ( .D(n4267), .SI(g3044), .SE(n9297), .CLK(n9484), .Q(
        g3045) );
  SDFFX1 DFF_1567_Q_reg ( .D(n4266), .SI(g3045), .SE(n9297), .CLK(n9484), .Q(
        g3046) );
  SDFFX1 DFF_1568_Q_reg ( .D(n4265), .SI(g3046), .SE(n9297), .CLK(n9484), .Q(
        g3047) );
  SDFFX1 DFF_1569_Q_reg ( .D(n4272), .SI(g3047), .SE(n9297), .CLK(n9484), .Q(
        g3048) );
  SDFFX1 DFF_1570_Q_reg ( .D(n4271), .SI(g3048), .SE(n9297), .CLK(n9484), .Q(
        g3049) );
  SDFFX1 DFF_1571_Q_reg ( .D(n4270), .SI(g3049), .SE(n9297), .CLK(n9484), .Q(
        g3050) );
  SDFFX1 DFF_1572_Q_reg ( .D(n4259), .SI(g3050), .SE(n9298), .CLK(n9485), .Q(
        g3051) );
  SDFFX1 DFF_1573_Q_reg ( .D(n4236), .SI(g3051), .SE(n9298), .CLK(n9485), .Q(
        g3052) );
  SDFFX1 DFF_1574_Q_reg ( .D(n4239), .SI(g3052), .SE(n9298), .CLK(n9485), .Q(
        g3053) );
  SDFFX1 DFF_1575_Q_reg ( .D(n4237), .SI(g3053), .SE(n9298), .CLK(n9485), .Q(
        test_so96) );
  SDFFX1 DFF_1576_Q_reg ( .D(n4234), .SI(test_si97), .SE(n9388), .CLK(n9575), 
        .Q(g3056) );
  SDFFX1 DFF_1577_Q_reg ( .D(n4233), .SI(g3056), .SE(n9388), .CLK(n9575), .Q(
        g3057) );
  SDFFX1 DFF_1578_Q_reg ( .D(n4238), .SI(g3057), .SE(n9388), .CLK(n9575), .Q(
        g3058) );
  SDFFX1 DFF_1579_Q_reg ( .D(n4235), .SI(g3058), .SE(n9388), .CLK(n9575), .Q(
        g3059) );
  SDFFX1 DFF_1580_Q_reg ( .D(n4240), .SI(g3059), .SE(n9389), .CLK(n9576), .Q(
        g3060) );
  SDFFX1 DFF_1581_Q_reg ( .D(n4232), .SI(g3060), .SE(n9389), .CLK(n9576), .Q(
        g3061) );
  SDFFX1 DFF_1582_Q_reg ( .D(n4245), .SI(g3061), .SE(n9415), .CLK(n9602), .Q(
        g3062) );
  SDFFX1 DFF_1583_Q_reg ( .D(n4248), .SI(g3062), .SE(n9416), .CLK(n9603), .Q(
        g3063) );
  SDFFX1 DFF_1584_Q_reg ( .D(n4246), .SI(g3063), .SE(n9416), .CLK(n9603), .Q(
        g3064) );
  SDFFX1 DFF_1585_Q_reg ( .D(n4243), .SI(g3064), .SE(n9416), .CLK(n9603), .Q(
        g3065) );
  SDFFX1 DFF_1586_Q_reg ( .D(n4242), .SI(g3065), .SE(n9416), .CLK(n9603), .Q(
        g3066) );
  SDFFX1 DFF_1587_Q_reg ( .D(n4247), .SI(g3066), .SE(n9416), .CLK(n9603), .Q(
        g3067) );
  SDFFX1 DFF_1588_Q_reg ( .D(n4244), .SI(g3067), .SE(n9416), .CLK(n9603), .Q(
        g3068) );
  SDFFX1 DFF_1589_Q_reg ( .D(n4249), .SI(g3068), .SE(n9416), .CLK(n9603), .Q(
        g3069) );
  SDFFX1 DFF_1590_Q_reg ( .D(n4241), .SI(g3069), .SE(n9416), .CLK(n9603), .Q(
        test_so97) );
  SDFFX1 DFF_1591_Q_reg ( .D(n4254), .SI(test_si98), .SE(n9418), .CLK(n9605), 
        .Q(g3071) );
  SDFFX1 DFF_1592_Q_reg ( .D(n4257), .SI(g3071), .SE(n9418), .CLK(n9605), .Q(
        g3072) );
  SDFFX1 DFF_1593_Q_reg ( .D(n4255), .SI(g3072), .SE(n9418), .CLK(n9605), .Q(
        g3073) );
  SDFFX1 DFF_1594_Q_reg ( .D(n4252), .SI(g3073), .SE(n9418), .CLK(n9605), .Q(
        g3074) );
  SDFFX1 DFF_1595_Q_reg ( .D(n4251), .SI(g3074), .SE(n9418), .CLK(n9605), .Q(
        g3075) );
  SDFFX1 DFF_1596_Q_reg ( .D(n4256), .SI(g3075), .SE(n9418), .CLK(n9605), .Q(
        g3076) );
  SDFFX1 DFF_1597_Q_reg ( .D(n4253), .SI(g3076), .SE(n9419), .CLK(n9606), .Q(
        g3077) );
  SDFFX1 DFF_1598_Q_reg ( .D(n4258), .SI(g3077), .SE(n9419), .CLK(n9606), .Q(
        g3078) );
  SDFFX1 DFF_1599_Q_reg ( .D(n4250), .SI(g3078), .SE(n9322), .CLK(n9509), .Q(
        g2997) );
  SDFFX1 DFF_1600_Q_reg ( .D(g25265), .SI(g2997), .SE(n9322), .CLK(n9509), .Q(
        g2993), .QN(n9261) );
  SDFFX1 DFF_1601_Q_reg ( .D(g26048), .SI(g2993), .SE(n9330), .CLK(n9517), .Q(
        n7909), .QN(n16834) );
  SDFFX1 DFF_1602_Q_reg ( .D(g23330), .SI(n7909), .SE(n9330), .CLK(n9517), .Q(
        g3006), .QN(n9263) );
  SDFFX1 DFF_1603_Q_reg ( .D(g24445), .SI(g3006), .SE(n9330), .CLK(n9517), .Q(
        g3002), .QN(n9262) );
  SDFFX1 DFF_1604_Q_reg ( .D(g25191), .SI(g3002), .SE(n9330), .CLK(n9517), .Q(
        g3013) );
  SDFFX1 DFF_1605_Q_reg ( .D(g26031), .SI(g3013), .SE(n9330), .CLK(n9517), .Q(
        test_so98), .QN(n9280) );
  SDFFX1 DFF_1606_Q_reg ( .D(g26786), .SI(test_si99), .SE(n9330), .CLK(n9517), 
        .Q(g3024), .QN(n8387) );
  SDFFX1 DFF_1607_Q_reg ( .D(n4262), .SI(g3024), .SE(n9416), .CLK(n9603), .Q(
        g3018), .QN(n4481) );
  SDFFX1 DFF_1608_Q_reg ( .D(g23359), .SI(g3018), .SE(n9416), .CLK(n9603), .Q(
        g3028), .QN(n4350) );
  SDFFX1 DFF_1609_Q_reg ( .D(g24446), .SI(g3028), .SE(n9416), .CLK(n9603), .Q(
        g3036), .QN(n4480) );
  SDFFX1 DFF_1610_Q_reg ( .D(g25202), .SI(g3036), .SE(n9416), .CLK(n9603), .Q(
        g3032), .QN(n8695) );
  SDFFX1 DFF_1611_Q_reg ( .D(g3234), .SI(g3032), .SE(n9417), .CLK(n9604), .Q(
        g5388) );
  SDFFX1 DFF_1612_Q_reg ( .D(g5388), .SI(g5388), .SE(n9417), .CLK(n9604), .Q(
        n7907), .QN(DFF_1612_n1) );
  SDFFX1 DFF_1613_Q_reg ( .D(g16496), .SI(n7907), .SE(n9417), .CLK(n9604), .Q(
        g2987), .QN(n4365) );
  SDFFX1 DFF_1614_Q_reg ( .D(g16824), .SI(g2987), .SE(n9417), .CLK(n9604), .Q(
        g8275), .QN(n9247) );
  SDFFX1 DFF_1615_Q_reg ( .D(g16844), .SI(g8275), .SE(n9417), .CLK(n9604), .Q(
        g8274), .QN(n9249) );
  SDFFX1 DFF_1616_Q_reg ( .D(g16853), .SI(g8274), .SE(n9417), .CLK(n9604), .Q(
        g8273), .QN(n16835) );
  SDFFX1 DFF_1617_Q_reg ( .D(g16860), .SI(g8273), .SE(n9417), .CLK(n9604), .Q(
        g8272), .QN(n16836) );
  SDFFX1 DFF_1618_Q_reg ( .D(g16803), .SI(g8272), .SE(n9417), .CLK(n9604), .Q(
        g8268), .QN(DFF_1618_n1) );
  SDFFX1 DFF_1619_Q_reg ( .D(g16835), .SI(g8268), .SE(n9417), .CLK(n9604), .Q(
        g8269), .QN(n9250) );
  SDFFX1 DFF_1620_Q_reg ( .D(g16851), .SI(g8269), .SE(n9417), .CLK(n9604), .Q(
        test_so99) );
  SDFFX1 DFF_1621_Q_reg ( .D(g16857), .SI(test_si100), .SE(n9417), .CLK(n9604), 
        .Q(g8271), .QN(n9248) );
  SDFFX1 DFF_1622_Q_reg ( .D(g16866), .SI(g8271), .SE(n9417), .CLK(n9604), .Q(
        g3083), .QN(n9253) );
  SDFFX1 DFF_1623_Q_reg ( .D(n4261), .SI(g3083), .SE(n9418), .CLK(n9605), .Q(
        g8267) );
  SDFFX1 DFF_1624_Q_reg ( .D(N995), .SI(g8267), .SE(n9418), .CLK(n9605), .Q(
        n4577), .QN(n8698) );
  SDFFX1 DFF_1625_Q_reg ( .D(g16845), .SI(n4577), .SE(n9418), .CLK(n9605), .Q(
        g8266), .QN(n16837) );
  SDFFX1 DFF_1626_Q_reg ( .D(g16854), .SI(g8266), .SE(n9418), .CLK(n9605), .Q(
        g8265), .QN(n16838) );
  SDFFX1 DFF_1627_Q_reg ( .D(g16861), .SI(g8265), .SE(n9298), .CLK(n9485), .Q(
        g8264), .QN(n9230) );
  SDFFX1 DFF_1628_Q_reg ( .D(g16880), .SI(g8264), .SE(n9418), .CLK(n9605), .Q(
        g8262), .QN(DFF_1628_n1) );
  SDFFX1 DFF_1629_Q_reg ( .D(g18755), .SI(g8262), .SE(n9418), .CLK(n9605), .Q(
        g8263), .QN(n9231) );
  SDFFX1 DFF_1630_Q_reg ( .D(g18804), .SI(g8263), .SE(n9419), .CLK(n9606), .Q(
        g8260), .QN(n9227) );
  SDFFX1 DFF_1631_Q_reg ( .D(g18837), .SI(g8260), .SE(n9419), .CLK(n9606), .Q(
        g8261), .QN(n9228) );
  SDFFX1 DFF_1632_Q_reg ( .D(g18868), .SI(g8261), .SE(n9419), .CLK(n9606), .Q(
        g8259), .QN(n9229) );
  SDFFX1 DFF_1633_Q_reg ( .D(g18907), .SI(g8259), .SE(n9419), .CLK(n9606), .Q(
        g2990), .QN(n9251) );
  SDFFX1 DFF_1634_Q_reg ( .D(N690), .SI(g2990), .SE(n9298), .CLK(n9485), .Q(
        n4578), .QN(n8697) );
  SDFFX1 DFF_1635_Q_reg ( .D(n4260), .SI(n4578), .SE(n9423), .CLK(n9610), .Q(
        test_so100) );
  SDFFX1 DFF_454_Q_reg ( .D(n4598), .SI(n8040), .SE(n9324), .CLK(n9511), .Q(
        g6677), .QN(n4309) );
  SDFFX1 DFF_804_Q_reg ( .D(n4598), .SI(test_si49), .SE(n9324), .CLK(n9511), 
        .Q(g6979), .QN(n4308) );
  SDFFX1 DFF_1154_Q_reg ( .D(n4598), .SI(n7960), .SE(n9323), .CLK(n9510), .Q(
        g7229), .QN(n4307) );
  SDFFX1 DFF_1504_Q_reg ( .D(n4598), .SI(n7918), .SE(n9329), .CLK(n9516), .Q(
        g7425), .QN(n4306) );
  SDFFX1 DFF_1300_Q_reg ( .D(g5555), .SI(g5555), .SE(n9399), .CLK(n9586), .Q(
        g7264), .QN(n4524) );
  SDFFX1 DFF_950_Q_reg ( .D(g5511), .SI(g5511), .SE(n9371), .CLK(n9558), .Q(
        g7014), .QN(n4525) );
  SDFFX1 DFF_951_Q_reg ( .D(g7014), .SI(g7014), .SE(n9371), .CLK(n9558), .Q(
        n4618), .QN(n4511) );
  SDFFX1 DFF_1301_Q_reg ( .D(g7264), .SI(g7264), .SE(n9399), .CLK(n9586), .Q(
        n4606), .QN(n4509) );
  SDFFX1 DFF_250_Q_reg ( .D(g5437), .SI(g5437), .SE(n9309), .CLK(n9496), .Q(
        g6447), .QN(n4499) );
  SDFFX1 DFF_249_Q_reg ( .D(g2950), .SI(g181), .SE(n9309), .CLK(n9496), .Q(
        g5437), .QN(n4520) );
  NOR2X0 Trojan1 ( .IN1(n3065), .IN2(n3016), .QN(Tj_OUT1) );
  NOR2X0 Trojan2 ( .IN1(n3023), .IN2(n3000), .QN(Tj_OUT2) );
  NOR2X0 Trojan3 ( .IN1(n3008), .IN2(n3068), .QN(Tj_OUT3) );
  NOR2X0 Trojan4 ( .IN1(n3128), .IN2(n3036), .QN(Tj_OUT4) );
  AND4X1 Trojan1234_NOT ( .IN1(Tj_OUT1), .IN2(Tj_OUT2), .IN3(Tj_OUT3), .IN4(
        Tj_OUT4), .Q(Tj_OUT1234) );
  NOR2X0 Trojan5 ( .IN1(n3758), .IN2(n3788), .QN(Tj_OUT5) );
  NOR2X0 Trojan6 ( .IN1(n3751), .IN2(n3749), .QN(Tj_OUT6) );
  NOR2X0 Trojan7 ( .IN1(n2792), .IN2(n2632), .QN(Tj_OUT7) );
  NOR2X0 Trojan8 ( .IN1(n1458), .IN2(n506), .QN(Tj_OUT8) );
  AND4X1 Trojan5678_NOT ( .IN1(Tj_OUT5), .IN2(Tj_OUT6), .IN3(Tj_OUT7), .IN4(
        Tj_OUT8), .Q(Tj_OUT5678) );
  AND2X1 Trojan_CLK_NOT ( .IN1(Tj_OUT1234), .IN2(Tj_OUT5678), .Q(Tj_Trigger)
         );
  OR2X1 Trojan_Payload ( .IN1(Tj_Trigger), .IN2(n4263), .Q(n4263_Tj_Payload)
         );
  NBUFFX2 U9102 ( .INP(n9467), .Z(n9294) );
  NBUFFX2 U9103 ( .INP(n9467), .Z(n9293) );
  NBUFFX2 U9104 ( .INP(n9426), .Z(n9417) );
  NBUFFX2 U9105 ( .INP(n9425), .Z(n9418) );
  NBUFFX2 U9106 ( .INP(n9426), .Z(n9416) );
  NBUFFX2 U9107 ( .INP(n9446), .Z(n9356) );
  NBUFFX2 U9108 ( .INP(n9446), .Z(n9355) );
  NBUFFX2 U9109 ( .INP(n9447), .Z(n9354) );
  NBUFFX2 U9110 ( .INP(n9428), .Z(n9411) );
  NBUFFX2 U9111 ( .INP(n9428), .Z(n9410) );
  NBUFFX2 U9112 ( .INP(n9429), .Z(n9407) );
  NBUFFX2 U9113 ( .INP(n9429), .Z(n9408) );
  NBUFFX2 U9114 ( .INP(n9428), .Z(n9409) );
  NBUFFX2 U9115 ( .INP(n9455), .Z(n9329) );
  NBUFFX2 U9116 ( .INP(n9427), .Z(n9414) );
  NBUFFX2 U9117 ( .INP(n9427), .Z(n9413) );
  NBUFFX2 U9118 ( .INP(n9426), .Z(n9415) );
  NBUFFX2 U9119 ( .INP(n9457), .Z(n9322) );
  NBUFFX2 U9120 ( .INP(n9430), .Z(n9405) );
  NBUFFX2 U9121 ( .INP(n9430), .Z(n9404) );
  NBUFFX2 U9122 ( .INP(n9429), .Z(n9406) );
  NBUFFX2 U9123 ( .INP(n9432), .Z(n9398) );
  NBUFFX2 U9124 ( .INP(n9432), .Z(n9397) );
  NBUFFX2 U9125 ( .INP(n9427), .Z(n9412) );
  NBUFFX2 U9126 ( .INP(n9430), .Z(n9403) );
  NBUFFX2 U9127 ( .INP(n9431), .Z(n9400) );
  NBUFFX2 U9128 ( .INP(n9432), .Z(n9399) );
  NBUFFX2 U9129 ( .INP(n9431), .Z(n9402) );
  NBUFFX2 U9130 ( .INP(n9431), .Z(n9401) );
  NBUFFX2 U9131 ( .INP(n9433), .Z(n9396) );
  NBUFFX2 U9132 ( .INP(n9433), .Z(n9395) );
  NBUFFX2 U9133 ( .INP(n9433), .Z(n9394) );
  NBUFFX2 U9134 ( .INP(n9434), .Z(n9393) );
  NBUFFX2 U9135 ( .INP(n9457), .Z(n9323) );
  NBUFFX2 U9136 ( .INP(n9434), .Z(n9392) );
  NBUFFX2 U9137 ( .INP(n9434), .Z(n9391) );
  NBUFFX2 U9138 ( .INP(n9435), .Z(n9390) );
  NBUFFX2 U9139 ( .INP(n9435), .Z(n9389) );
  NBUFFX2 U9140 ( .INP(n9435), .Z(n9388) );
  NBUFFX2 U9141 ( .INP(n9436), .Z(n9387) );
  NBUFFX2 U9142 ( .INP(n9436), .Z(n9386) );
  NBUFFX2 U9143 ( .INP(n9436), .Z(n9385) );
  NBUFFX2 U9144 ( .INP(n9437), .Z(n9384) );
  NBUFFX2 U9145 ( .INP(n9437), .Z(n9383) );
  NBUFFX2 U9146 ( .INP(n9437), .Z(n9382) );
  NBUFFX2 U9147 ( .INP(n9441), .Z(n9372) );
  NBUFFX2 U9148 ( .INP(n9438), .Z(n9381) );
  NBUFFX2 U9149 ( .INP(n9439), .Z(n9378) );
  NBUFFX2 U9150 ( .INP(n9438), .Z(n9379) );
  NBUFFX2 U9151 ( .INP(n9441), .Z(n9371) );
  NBUFFX2 U9152 ( .INP(n9441), .Z(n9370) );
  NBUFFX2 U9153 ( .INP(n9439), .Z(n9377) );
  NBUFFX2 U9154 ( .INP(n9438), .Z(n9380) );
  NBUFFX2 U9155 ( .INP(n9439), .Z(n9376) );
  NBUFFX2 U9156 ( .INP(n9440), .Z(n9375) );
  NBUFFX2 U9157 ( .INP(n9440), .Z(n9374) );
  NBUFFX2 U9158 ( .INP(n9440), .Z(n9373) );
  NBUFFX2 U9159 ( .INP(n9442), .Z(n9369) );
  NBUFFX2 U9160 ( .INP(n9442), .Z(n9368) );
  NBUFFX2 U9161 ( .INP(n9442), .Z(n9367) );
  NBUFFX2 U9162 ( .INP(n9443), .Z(n9366) );
  NBUFFX2 U9163 ( .INP(n9443), .Z(n9365) );
  NBUFFX2 U9164 ( .INP(n9443), .Z(n9364) );
  NBUFFX2 U9165 ( .INP(n9444), .Z(n9363) );
  NBUFFX2 U9166 ( .INP(n9444), .Z(n9362) );
  NBUFFX2 U9167 ( .INP(n9447), .Z(n9352) );
  NBUFFX2 U9168 ( .INP(n9448), .Z(n9351) );
  NBUFFX2 U9169 ( .INP(n9448), .Z(n9350) );
  NBUFFX2 U9170 ( .INP(n9448), .Z(n9349) );
  NBUFFX2 U9171 ( .INP(n9449), .Z(n9348) );
  NBUFFX2 U9172 ( .INP(n9449), .Z(n9347) );
  NBUFFX2 U9173 ( .INP(n9450), .Z(n9344) );
  NBUFFX2 U9174 ( .INP(n9450), .Z(n9343) );
  NBUFFX2 U9175 ( .INP(n9449), .Z(n9346) );
  NBUFFX2 U9176 ( .INP(n9450), .Z(n9345) );
  NBUFFX2 U9177 ( .INP(n9453), .Z(n9336) );
  NBUFFX2 U9178 ( .INP(n9451), .Z(n9342) );
  NBUFFX2 U9179 ( .INP(n9451), .Z(n9341) );
  NBUFFX2 U9180 ( .INP(n9451), .Z(n9340) );
  NBUFFX2 U9181 ( .INP(n9452), .Z(n9337) );
  NBUFFX2 U9182 ( .INP(n9452), .Z(n9339) );
  NBUFFX2 U9183 ( .INP(n9452), .Z(n9338) );
  NBUFFX2 U9184 ( .INP(n9453), .Z(n9335) );
  NBUFFX2 U9185 ( .INP(n9453), .Z(n9334) );
  NBUFFX2 U9186 ( .INP(n9447), .Z(n9353) );
  NBUFFX2 U9187 ( .INP(n9454), .Z(n9333) );
  NBUFFX2 U9188 ( .INP(n9454), .Z(n9332) );
  NBUFFX2 U9189 ( .INP(n9454), .Z(n9331) );
  NBUFFX2 U9190 ( .INP(n9455), .Z(n9330) );
  NBUFFX2 U9191 ( .INP(n9444), .Z(n9361) );
  NBUFFX2 U9192 ( .INP(n9445), .Z(n9360) );
  NBUFFX2 U9193 ( .INP(n9445), .Z(n9359) );
  NBUFFX2 U9194 ( .INP(n9446), .Z(n9357) );
  NBUFFX2 U9195 ( .INP(n9445), .Z(n9358) );
  NBUFFX2 U9196 ( .INP(n9455), .Z(n9328) );
  NBUFFX2 U9197 ( .INP(n9456), .Z(n9327) );
  NBUFFX2 U9198 ( .INP(n9456), .Z(n9326) );
  NBUFFX2 U9199 ( .INP(n9456), .Z(n9325) );
  NBUFFX2 U9200 ( .INP(n9457), .Z(n9324) );
  NBUFFX2 U9201 ( .INP(n9459), .Z(n9317) );
  NBUFFX2 U9202 ( .INP(n9466), .Z(n9297) );
  NBUFFX2 U9203 ( .INP(n9462), .Z(n9307) );
  NBUFFX2 U9204 ( .INP(n9463), .Z(n9306) );
  NBUFFX2 U9205 ( .INP(n9460), .Z(n9314) );
  NBUFFX2 U9206 ( .INP(n9460), .Z(n9315) );
  NBUFFX2 U9207 ( .INP(n9459), .Z(n9316) );
  NBUFFX2 U9208 ( .INP(n9462), .Z(n9309) );
  NBUFFX2 U9209 ( .INP(n9458), .Z(n9320) );
  NBUFFX2 U9210 ( .INP(n9458), .Z(n9319) );
  NBUFFX2 U9211 ( .INP(n9459), .Z(n9318) );
  NBUFFX2 U9212 ( .INP(n9461), .Z(n9310) );
  NBUFFX2 U9213 ( .INP(n9462), .Z(n9308) );
  NBUFFX2 U9214 ( .INP(n9461), .Z(n9311) );
  NBUFFX2 U9215 ( .INP(n9460), .Z(n9313) );
  NBUFFX2 U9216 ( .INP(n9461), .Z(n9312) );
  NBUFFX2 U9217 ( .INP(n9465), .Z(n9298) );
  NBUFFX2 U9218 ( .INP(n9465), .Z(n9299) );
  NBUFFX2 U9219 ( .INP(n9424), .Z(n9422) );
  NBUFFX2 U9220 ( .INP(n9424), .Z(n9421) );
  NBUFFX2 U9221 ( .INP(n9425), .Z(n9420) );
  NBUFFX2 U9222 ( .INP(n9425), .Z(n9419) );
  NBUFFX2 U9223 ( .INP(n9458), .Z(n9321) );
  NBUFFX2 U9224 ( .INP(n9463), .Z(n9305) );
  NBUFFX2 U9225 ( .INP(n9463), .Z(n9304) );
  NBUFFX2 U9226 ( .INP(n9464), .Z(n9303) );
  NBUFFX2 U9227 ( .INP(n9464), .Z(n9302) );
  NBUFFX2 U9228 ( .INP(n9464), .Z(n9301) );
  NBUFFX2 U9229 ( .INP(n9465), .Z(n9300) );
  NBUFFX2 U9230 ( .INP(n9466), .Z(n9296) );
  NBUFFX2 U9231 ( .INP(n9466), .Z(n9295) );
  NBUFFX2 U9232 ( .INP(n9654), .Z(n9481) );
  NBUFFX2 U9233 ( .INP(n9654), .Z(n9480) );
  NBUFFX2 U9234 ( .INP(n9613), .Z(n9604) );
  NBUFFX2 U9235 ( .INP(n9612), .Z(n9605) );
  NBUFFX2 U9236 ( .INP(n9613), .Z(n9603) );
  NBUFFX2 U9237 ( .INP(n9633), .Z(n9543) );
  NBUFFX2 U9238 ( .INP(n9633), .Z(n9542) );
  NBUFFX2 U9239 ( .INP(n9634), .Z(n9541) );
  NBUFFX2 U9240 ( .INP(n9615), .Z(n9598) );
  NBUFFX2 U9241 ( .INP(n9615), .Z(n9597) );
  NBUFFX2 U9242 ( .INP(n9616), .Z(n9594) );
  NBUFFX2 U9243 ( .INP(n9616), .Z(n9595) );
  NBUFFX2 U9244 ( .INP(n9615), .Z(n9596) );
  NBUFFX2 U9245 ( .INP(n9642), .Z(n9516) );
  NBUFFX2 U9246 ( .INP(n9614), .Z(n9601) );
  NBUFFX2 U9247 ( .INP(n9614), .Z(n9600) );
  NBUFFX2 U9248 ( .INP(n9613), .Z(n9602) );
  NBUFFX2 U9249 ( .INP(n9644), .Z(n9509) );
  NBUFFX2 U9250 ( .INP(n9617), .Z(n9592) );
  NBUFFX2 U9251 ( .INP(n9617), .Z(n9591) );
  NBUFFX2 U9252 ( .INP(n9616), .Z(n9593) );
  NBUFFX2 U9253 ( .INP(n9619), .Z(n9585) );
  NBUFFX2 U9254 ( .INP(n9619), .Z(n9584) );
  NBUFFX2 U9255 ( .INP(n9614), .Z(n9599) );
  NBUFFX2 U9256 ( .INP(n9617), .Z(n9590) );
  NBUFFX2 U9257 ( .INP(n9618), .Z(n9587) );
  NBUFFX2 U9258 ( .INP(n9619), .Z(n9586) );
  NBUFFX2 U9259 ( .INP(n9618), .Z(n9589) );
  NBUFFX2 U9260 ( .INP(n9618), .Z(n9588) );
  NBUFFX2 U9261 ( .INP(n9620), .Z(n9583) );
  NBUFFX2 U9262 ( .INP(n9620), .Z(n9582) );
  NBUFFX2 U9263 ( .INP(n9620), .Z(n9581) );
  NBUFFX2 U9264 ( .INP(n9621), .Z(n9580) );
  NBUFFX2 U9265 ( .INP(n9644), .Z(n9510) );
  NBUFFX2 U9266 ( .INP(n9621), .Z(n9579) );
  NBUFFX2 U9267 ( .INP(n9621), .Z(n9578) );
  NBUFFX2 U9268 ( .INP(n9622), .Z(n9577) );
  NBUFFX2 U9269 ( .INP(n9622), .Z(n9576) );
  NBUFFX2 U9270 ( .INP(n9622), .Z(n9575) );
  NBUFFX2 U9271 ( .INP(n9623), .Z(n9574) );
  NBUFFX2 U9272 ( .INP(n9623), .Z(n9573) );
  NBUFFX2 U9273 ( .INP(n9623), .Z(n9572) );
  NBUFFX2 U9274 ( .INP(n9624), .Z(n9571) );
  NBUFFX2 U9275 ( .INP(n9624), .Z(n9570) );
  NBUFFX2 U9276 ( .INP(n9624), .Z(n9569) );
  NBUFFX2 U9277 ( .INP(n9628), .Z(n9559) );
  NBUFFX2 U9278 ( .INP(n9625), .Z(n9568) );
  NBUFFX2 U9279 ( .INP(n9626), .Z(n9565) );
  NBUFFX2 U9280 ( .INP(n9625), .Z(n9566) );
  NBUFFX2 U9281 ( .INP(n9628), .Z(n9558) );
  NBUFFX2 U9282 ( .INP(n9628), .Z(n9557) );
  NBUFFX2 U9283 ( .INP(n9626), .Z(n9564) );
  NBUFFX2 U9284 ( .INP(n9625), .Z(n9567) );
  NBUFFX2 U9285 ( .INP(n9626), .Z(n9563) );
  NBUFFX2 U9286 ( .INP(n9627), .Z(n9562) );
  NBUFFX2 U9287 ( .INP(n9627), .Z(n9561) );
  NBUFFX2 U9288 ( .INP(n9627), .Z(n9560) );
  NBUFFX2 U9289 ( .INP(n9629), .Z(n9556) );
  NBUFFX2 U9290 ( .INP(n9629), .Z(n9555) );
  NBUFFX2 U9291 ( .INP(n9629), .Z(n9554) );
  NBUFFX2 U9292 ( .INP(n9630), .Z(n9553) );
  NBUFFX2 U9293 ( .INP(n9630), .Z(n9552) );
  NBUFFX2 U9294 ( .INP(n9630), .Z(n9551) );
  NBUFFX2 U9295 ( .INP(n9631), .Z(n9550) );
  NBUFFX2 U9296 ( .INP(n9631), .Z(n9549) );
  NBUFFX2 U9297 ( .INP(n9634), .Z(n9539) );
  NBUFFX2 U9298 ( .INP(n9635), .Z(n9538) );
  NBUFFX2 U9299 ( .INP(n9635), .Z(n9537) );
  NBUFFX2 U9300 ( .INP(n9635), .Z(n9536) );
  NBUFFX2 U9301 ( .INP(n9636), .Z(n9535) );
  NBUFFX2 U9302 ( .INP(n9636), .Z(n9534) );
  NBUFFX2 U9303 ( .INP(n9637), .Z(n9531) );
  NBUFFX2 U9304 ( .INP(n9637), .Z(n9530) );
  NBUFFX2 U9305 ( .INP(n9636), .Z(n9533) );
  NBUFFX2 U9306 ( .INP(n9637), .Z(n9532) );
  NBUFFX2 U9307 ( .INP(n9640), .Z(n9523) );
  NBUFFX2 U9308 ( .INP(n9638), .Z(n9529) );
  NBUFFX2 U9309 ( .INP(n9638), .Z(n9528) );
  NBUFFX2 U9310 ( .INP(n9638), .Z(n9527) );
  NBUFFX2 U9311 ( .INP(n9639), .Z(n9524) );
  NBUFFX2 U9312 ( .INP(n9639), .Z(n9526) );
  NBUFFX2 U9313 ( .INP(n9639), .Z(n9525) );
  NBUFFX2 U9314 ( .INP(n9640), .Z(n9522) );
  NBUFFX2 U9315 ( .INP(n9640), .Z(n9521) );
  NBUFFX2 U9316 ( .INP(n9634), .Z(n9540) );
  NBUFFX2 U9317 ( .INP(n9641), .Z(n9520) );
  NBUFFX2 U9318 ( .INP(n9641), .Z(n9519) );
  NBUFFX2 U9319 ( .INP(n9641), .Z(n9518) );
  NBUFFX2 U9320 ( .INP(n9642), .Z(n9517) );
  NBUFFX2 U9321 ( .INP(n9631), .Z(n9548) );
  NBUFFX2 U9322 ( .INP(n9632), .Z(n9547) );
  NBUFFX2 U9323 ( .INP(n9632), .Z(n9546) );
  NBUFFX2 U9324 ( .INP(n9633), .Z(n9544) );
  NBUFFX2 U9325 ( .INP(n9632), .Z(n9545) );
  NBUFFX2 U9326 ( .INP(n9642), .Z(n9515) );
  NBUFFX2 U9327 ( .INP(n9643), .Z(n9514) );
  NBUFFX2 U9328 ( .INP(n9643), .Z(n9513) );
  NBUFFX2 U9329 ( .INP(n9643), .Z(n9512) );
  NBUFFX2 U9330 ( .INP(n9644), .Z(n9511) );
  NBUFFX2 U9331 ( .INP(n9646), .Z(n9504) );
  NBUFFX2 U9332 ( .INP(n9653), .Z(n9484) );
  NBUFFX2 U9333 ( .INP(n9649), .Z(n9494) );
  NBUFFX2 U9334 ( .INP(n9650), .Z(n9493) );
  NBUFFX2 U9335 ( .INP(n9647), .Z(n9501) );
  NBUFFX2 U9336 ( .INP(n9647), .Z(n9502) );
  NBUFFX2 U9337 ( .INP(n9646), .Z(n9503) );
  NBUFFX2 U9338 ( .INP(n9649), .Z(n9496) );
  NBUFFX2 U9339 ( .INP(n9645), .Z(n9507) );
  NBUFFX2 U9340 ( .INP(n9645), .Z(n9506) );
  NBUFFX2 U9341 ( .INP(n9646), .Z(n9505) );
  NBUFFX2 U9342 ( .INP(n9648), .Z(n9497) );
  NBUFFX2 U9343 ( .INP(n9649), .Z(n9495) );
  NBUFFX2 U9344 ( .INP(n9648), .Z(n9498) );
  NBUFFX2 U9345 ( .INP(n9647), .Z(n9500) );
  NBUFFX2 U9346 ( .INP(n9648), .Z(n9499) );
  NBUFFX2 U9347 ( .INP(n9652), .Z(n9485) );
  NBUFFX2 U9348 ( .INP(n9652), .Z(n9486) );
  NBUFFX2 U9349 ( .INP(n9611), .Z(n9609) );
  NBUFFX2 U9350 ( .INP(n9611), .Z(n9608) );
  NBUFFX2 U9351 ( .INP(n9612), .Z(n9607) );
  NBUFFX2 U9352 ( .INP(n9612), .Z(n9606) );
  NBUFFX2 U9353 ( .INP(n9645), .Z(n9508) );
  NBUFFX2 U9354 ( .INP(n9650), .Z(n9492) );
  NBUFFX2 U9355 ( .INP(n9650), .Z(n9491) );
  NBUFFX2 U9356 ( .INP(n9651), .Z(n9490) );
  NBUFFX2 U9357 ( .INP(n9651), .Z(n9489) );
  NBUFFX2 U9358 ( .INP(n9651), .Z(n9488) );
  NBUFFX2 U9359 ( .INP(n9652), .Z(n9487) );
  NBUFFX2 U9360 ( .INP(n9653), .Z(n9483) );
  NBUFFX2 U9361 ( .INP(n9653), .Z(n9482) );
  NBUFFX2 U9362 ( .INP(n9424), .Z(n9423) );
  NBUFFX2 U9363 ( .INP(n9611), .Z(n9610) );
  NBUFFX2 U9364 ( .INP(n9663), .Z(n9613) );
  NBUFFX2 U9365 ( .INP(n9476), .Z(n9426) );
  NBUFFX2 U9366 ( .INP(n9663), .Z(n9614) );
  NBUFFX2 U9367 ( .INP(n9476), .Z(n9427) );
  NBUFFX2 U9368 ( .INP(n9663), .Z(n9611) );
  NBUFFX2 U9369 ( .INP(n9476), .Z(n9424) );
  NBUFFX2 U9370 ( .INP(n9663), .Z(n9612) );
  NBUFFX2 U9371 ( .INP(n9476), .Z(n9425) );
  NBUFFX2 U9372 ( .INP(n9662), .Z(n9615) );
  NBUFFX2 U9373 ( .INP(n9475), .Z(n9428) );
  NBUFFX2 U9374 ( .INP(n9662), .Z(n9616) );
  NBUFFX2 U9375 ( .INP(n9475), .Z(n9429) );
  NBUFFX2 U9376 ( .INP(n9662), .Z(n9617) );
  NBUFFX2 U9377 ( .INP(n9475), .Z(n9430) );
  NBUFFX2 U9378 ( .INP(n9662), .Z(n9619) );
  NBUFFX2 U9379 ( .INP(n9475), .Z(n9432) );
  NBUFFX2 U9380 ( .INP(n9662), .Z(n9618) );
  NBUFFX2 U9381 ( .INP(n9475), .Z(n9431) );
  NBUFFX2 U9382 ( .INP(n9661), .Z(n9620) );
  NBUFFX2 U9383 ( .INP(n9474), .Z(n9433) );
  NBUFFX2 U9384 ( .INP(n9661), .Z(n9621) );
  NBUFFX2 U9385 ( .INP(n9474), .Z(n9434) );
  NBUFFX2 U9386 ( .INP(n9661), .Z(n9622) );
  NBUFFX2 U9387 ( .INP(n9474), .Z(n9435) );
  NBUFFX2 U9388 ( .INP(n9661), .Z(n9623) );
  NBUFFX2 U9389 ( .INP(n9474), .Z(n9436) );
  NBUFFX2 U9390 ( .INP(n9661), .Z(n9624) );
  NBUFFX2 U9391 ( .INP(n9474), .Z(n9437) );
  NBUFFX2 U9392 ( .INP(n9660), .Z(n9628) );
  NBUFFX2 U9393 ( .INP(n9473), .Z(n9441) );
  NBUFFX2 U9394 ( .INP(n9660), .Z(n9625) );
  NBUFFX2 U9395 ( .INP(n9473), .Z(n9438) );
  NBUFFX2 U9396 ( .INP(n9660), .Z(n9626) );
  NBUFFX2 U9397 ( .INP(n9473), .Z(n9439) );
  NBUFFX2 U9398 ( .INP(n9660), .Z(n9627) );
  NBUFFX2 U9399 ( .INP(n9473), .Z(n9440) );
  NBUFFX2 U9400 ( .INP(n9660), .Z(n9629) );
  NBUFFX2 U9401 ( .INP(n9473), .Z(n9442) );
  NBUFFX2 U9402 ( .INP(n9659), .Z(n9630) );
  NBUFFX2 U9403 ( .INP(n9472), .Z(n9443) );
  NBUFFX2 U9404 ( .INP(n9658), .Z(n9635) );
  NBUFFX2 U9405 ( .INP(n9471), .Z(n9448) );
  NBUFFX2 U9406 ( .INP(n9658), .Z(n9636) );
  NBUFFX2 U9407 ( .INP(n9471), .Z(n9449) );
  NBUFFX2 U9408 ( .INP(n9658), .Z(n9637) );
  NBUFFX2 U9409 ( .INP(n9471), .Z(n9450) );
  NBUFFX2 U9410 ( .INP(n9658), .Z(n9638) );
  NBUFFX2 U9411 ( .INP(n9471), .Z(n9451) );
  NBUFFX2 U9412 ( .INP(n9658), .Z(n9639) );
  NBUFFX2 U9413 ( .INP(n9471), .Z(n9452) );
  NBUFFX2 U9414 ( .INP(n9657), .Z(n9640) );
  NBUFFX2 U9415 ( .INP(n9470), .Z(n9453) );
  NBUFFX2 U9416 ( .INP(n9659), .Z(n9634) );
  NBUFFX2 U9417 ( .INP(n9472), .Z(n9447) );
  NBUFFX2 U9418 ( .INP(n9657), .Z(n9641) );
  NBUFFX2 U9419 ( .INP(n9470), .Z(n9454) );
  NBUFFX2 U9420 ( .INP(n9659), .Z(n9631) );
  NBUFFX2 U9421 ( .INP(n9472), .Z(n9444) );
  NBUFFX2 U9422 ( .INP(n9659), .Z(n9633) );
  NBUFFX2 U9423 ( .INP(n9472), .Z(n9446) );
  NBUFFX2 U9424 ( .INP(n9659), .Z(n9632) );
  NBUFFX2 U9425 ( .INP(n9472), .Z(n9445) );
  NBUFFX2 U9426 ( .INP(n9657), .Z(n9642) );
  NBUFFX2 U9427 ( .INP(n9470), .Z(n9455) );
  NBUFFX2 U9428 ( .INP(n9657), .Z(n9643) );
  NBUFFX2 U9429 ( .INP(n9470), .Z(n9456) );
  NBUFFX2 U9430 ( .INP(n9657), .Z(n9644) );
  NBUFFX2 U9431 ( .INP(n9470), .Z(n9457) );
  NBUFFX2 U9432 ( .INP(n9656), .Z(n9646) );
  NBUFFX2 U9433 ( .INP(n9469), .Z(n9459) );
  NBUFFX2 U9434 ( .INP(n9656), .Z(n9649) );
  NBUFFX2 U9435 ( .INP(n9469), .Z(n9462) );
  NBUFFX2 U9436 ( .INP(n9656), .Z(n9647) );
  NBUFFX2 U9437 ( .INP(n9469), .Z(n9460) );
  NBUFFX2 U9438 ( .INP(n9656), .Z(n9648) );
  NBUFFX2 U9439 ( .INP(n9469), .Z(n9461) );
  NBUFFX2 U9440 ( .INP(n9656), .Z(n9645) );
  NBUFFX2 U9441 ( .INP(n9469), .Z(n9458) );
  NBUFFX2 U9442 ( .INP(n9655), .Z(n9650) );
  NBUFFX2 U9443 ( .INP(n9468), .Z(n9463) );
  NBUFFX2 U9444 ( .INP(n9655), .Z(n9651) );
  NBUFFX2 U9445 ( .INP(n9468), .Z(n9464) );
  NBUFFX2 U9446 ( .INP(n9655), .Z(n9652) );
  NBUFFX2 U9447 ( .INP(n9468), .Z(n9465) );
  NBUFFX2 U9448 ( .INP(n9655), .Z(n9653) );
  NBUFFX2 U9449 ( .INP(n9468), .Z(n9466) );
  NBUFFX2 U9450 ( .INP(n9655), .Z(n9654) );
  NBUFFX2 U9451 ( .INP(n9468), .Z(n9467) );
  NBUFFX2 U9452 ( .INP(n9479), .Z(n9468) );
  NBUFFX2 U9453 ( .INP(n9479), .Z(n9469) );
  NBUFFX2 U9454 ( .INP(n9479), .Z(n9470) );
  NBUFFX2 U9455 ( .INP(n9478), .Z(n9471) );
  NBUFFX2 U9456 ( .INP(n9478), .Z(n9472) );
  NBUFFX2 U9457 ( .INP(n9478), .Z(n9473) );
  NBUFFX2 U9458 ( .INP(n9477), .Z(n9474) );
  NBUFFX2 U9459 ( .INP(n9477), .Z(n9475) );
  NBUFFX2 U9460 ( .INP(n9477), .Z(n9476) );
  NBUFFX2 U9461 ( .INP(test_se), .Z(n9477) );
  NBUFFX2 U9462 ( .INP(test_se), .Z(n9478) );
  NBUFFX2 U9463 ( .INP(test_se), .Z(n9479) );
  NBUFFX2 U9464 ( .INP(n9666), .Z(n9655) );
  NBUFFX2 U9465 ( .INP(n9666), .Z(n9656) );
  NBUFFX2 U9466 ( .INP(n9666), .Z(n9657) );
  NBUFFX2 U9467 ( .INP(n9665), .Z(n9658) );
  NBUFFX2 U9468 ( .INP(n9665), .Z(n9659) );
  NBUFFX2 U9469 ( .INP(n9665), .Z(n9660) );
  NBUFFX2 U9470 ( .INP(n9664), .Z(n9661) );
  NBUFFX2 U9471 ( .INP(n9664), .Z(n9662) );
  NBUFFX2 U9472 ( .INP(n9664), .Z(n9663) );
  NBUFFX2 U9473 ( .INP(CK), .Z(n9664) );
  NBUFFX2 U9474 ( .INP(CK), .Z(n9665) );
  NBUFFX2 U9475 ( .INP(CK), .Z(n9666) );
  INVX0 U9476 ( .INP(n9667), .ZN(n984) );
  INVX0 U9477 ( .INP(g27380), .ZN(n92) );
  INVX0 U9478 ( .INP(n9668), .ZN(n890) );
  NAND2X0 U9479 ( .IN1(n9669), .IN2(n9670), .QN(n9668) );
  NAND2X0 U9480 ( .IN1(n9671), .IN2(n9154), .QN(n9670) );
  INVX0 U9481 ( .INP(n9672), .ZN(n854) );
  NOR2X0 U9482 ( .IN1(n9673), .IN2(n9674), .QN(n9672) );
  NOR2X0 U9483 ( .IN1(g1236), .IN2(n9225), .QN(n9674) );
  INVX0 U9484 ( .INP(n9675), .ZN(n846) );
  INVX0 U9485 ( .INP(n9676), .ZN(n7) );
  NAND2X0 U9486 ( .IN1(n9677), .IN2(n9678), .QN(n9676) );
  NOR2X0 U9487 ( .IN1(n4057), .IN2(n9679), .QN(n9678) );
  INVX0 U9488 ( .INP(n9680), .ZN(n681) );
  INVX0 U9489 ( .INP(n9681), .ZN(n614) );
  NAND2X0 U9490 ( .IN1(n9682), .IN2(n9683), .QN(n9681) );
  NOR2X0 U9491 ( .IN1(n9684), .IN2(n9685), .QN(n9683) );
  NAND2X0 U9492 ( .IN1(n9686), .IN2(n4396), .QN(n9682) );
  INVX0 U9493 ( .INP(n9687), .ZN(n6) );
  NAND2X0 U9494 ( .IN1(n9677), .IN2(n9688), .QN(n9687) );
  NOR2X0 U9495 ( .IN1(n4122), .IN2(n9689), .QN(n9688) );
  INVX0 U9496 ( .INP(n9690), .ZN(n589) );
  NAND2X0 U9497 ( .IN1(n9691), .IN2(n9692), .QN(n9690) );
  NAND2X0 U9498 ( .IN1(n9693), .IN2(n9155), .QN(n9692) );
  INVX0 U9499 ( .INP(n9694), .ZN(n552) );
  NOR2X0 U9500 ( .IN1(n9695), .IN2(n9696), .QN(n9694) );
  NOR2X0 U9501 ( .IN1(g550), .IN2(n9226), .QN(n9696) );
  INVX0 U9502 ( .INP(n9697), .ZN(n550) );
  INVX0 U9503 ( .INP(n9698), .ZN(n549) );
  INVX0 U9504 ( .INP(n9699), .ZN(n54) );
  NAND2X0 U9505 ( .IN1(n4522), .IN2(n9700), .QN(n9699) );
  NOR2X0 U9506 ( .IN1(n9701), .IN2(n9702), .QN(n9700) );
  NOR2X0 U9507 ( .IN1(g2147), .IN2(n3683), .QN(n9701) );
  INVX0 U9508 ( .INP(n9703), .ZN(n53) );
  NAND2X0 U9509 ( .IN1(n4526), .IN2(n9704), .QN(n9703) );
  NOR2X0 U9510 ( .IN1(n9705), .IN2(n9702), .QN(n9704) );
  NOR2X0 U9511 ( .IN1(test_so78), .IN2(n3887), .QN(n9705) );
  INVX0 U9512 ( .INP(n9706), .ZN(n522) );
  INVX0 U9513 ( .INP(n9707), .ZN(n51) );
  NAND2X0 U9514 ( .IN1(n4523), .IN2(n9708), .QN(n9707) );
  NOR2X0 U9515 ( .IN1(n9709), .IN2(n9710), .QN(n9708) );
  NOR2X0 U9516 ( .IN1(g1453), .IN2(n3686), .QN(n9709) );
  INVX0 U9517 ( .INP(n9711), .ZN(n50) );
  NAND2X0 U9518 ( .IN1(n4527), .IN2(n9712), .QN(n9711) );
  NOR2X0 U9519 ( .IN1(n9713), .IN2(n9710), .QN(n9712) );
  NOR2X0 U9520 ( .IN1(g1462), .IN2(n3890), .QN(n9713) );
  INVX0 U9521 ( .INP(n9714), .ZN(n492) );
  INVX0 U9522 ( .INP(n9715), .ZN(n477) );
  INVX0 U9523 ( .INP(n9716), .ZN(n47) );
  NAND2X0 U9524 ( .IN1(n4521), .IN2(n9717), .QN(n9716) );
  NOR2X0 U9525 ( .IN1(n9718), .IN2(n9719), .QN(n9717) );
  NOR2X0 U9526 ( .IN1(test_so15), .IN2(n3692), .QN(n9718) );
  INVX0 U9527 ( .INP(n9720), .ZN(n46) );
  NAND2X0 U9528 ( .IN1(n4528), .IN2(n9721), .QN(n9720) );
  NOR2X0 U9529 ( .IN1(n9722), .IN2(n9719), .QN(n9721) );
  NOR2X0 U9530 ( .IN1(g88), .IN2(n3896), .QN(n9722) );
  XOR2X1 U9531 ( .IN1(n9252), .IN2(n9723), .Q(n4281) );
  XOR2X1 U9532 ( .IN1(g2934), .IN2(n9724), .Q(n4280) );
  NAND2X0 U9533 ( .IN1(g2879), .IN2(n9725), .QN(n4279) );
  NAND2X0 U9534 ( .IN1(DFF_18_n1), .IN2(g8021), .QN(n9725) );
  NOR2X0 U9535 ( .IN1(n9726), .IN2(n9727), .QN(n4278) );
  NOR2X0 U9536 ( .IN1(n9728), .IN2(n9729), .QN(n9727) );
  NOR2X0 U9537 ( .IN1(n9730), .IN2(n9731), .QN(n9726) );
  NAND2X0 U9538 ( .IN1(n9732), .IN2(n9733), .QN(n9731) );
  NOR2X0 U9539 ( .IN1(n9734), .IN2(n9735), .QN(n9733) );
  NAND2X0 U9540 ( .IN1(n9736), .IN2(n9737), .QN(n9735) );
  XNOR2X1 U9541 ( .IN1(n9738), .IN2(n8981), .Q(n9737) );
  XNOR2X1 U9542 ( .IN1(n9739), .IN2(n9264), .Q(n9736) );
  XNOR2X1 U9543 ( .IN1(n9266), .IN2(n9740), .Q(n9734) );
  NOR2X0 U9544 ( .IN1(n9741), .IN2(n9742), .QN(n9732) );
  NAND2X0 U9545 ( .IN1(n9743), .IN2(n9744), .QN(n9742) );
  XNOR2X1 U9546 ( .IN1(n9745), .IN2(n8983), .Q(n9744) );
  XNOR2X1 U9547 ( .IN1(n9746), .IN2(n8562), .Q(n9743) );
  XNOR2X1 U9548 ( .IN1(n8982), .IN2(n9747), .Q(n9741) );
  NAND2X0 U9549 ( .IN1(n9748), .IN2(n9749), .QN(n9730) );
  NOR2X0 U9550 ( .IN1(n9750), .IN2(n9751), .QN(n9749) );
  NAND2X0 U9551 ( .IN1(n9752), .IN2(n9753), .QN(n9751) );
  XNOR2X1 U9552 ( .IN1(n9754), .IN2(test_so15), .Q(n9750) );
  NOR2X0 U9553 ( .IN1(n9755), .IN2(n9756), .QN(n9748) );
  NAND2X0 U9554 ( .IN1(n9757), .IN2(n9758), .QN(n9756) );
  XNOR2X1 U9555 ( .IN1(n9759), .IN2(n8391), .Q(n9758) );
  XNOR2X1 U9556 ( .IN1(n4513), .IN2(n8984), .Q(n9757) );
  XNOR2X1 U9557 ( .IN1(n9275), .IN2(n9760), .Q(n9755) );
  NOR2X0 U9558 ( .IN1(n9761), .IN2(n9762), .QN(n4277) );
  NOR2X0 U9559 ( .IN1(n9763), .IN2(n9764), .QN(n9762) );
  NOR2X0 U9560 ( .IN1(n9765), .IN2(n9766), .QN(n9761) );
  NAND2X0 U9561 ( .IN1(n9767), .IN2(n9768), .QN(n9766) );
  NOR2X0 U9562 ( .IN1(n9769), .IN2(n9770), .QN(n9768) );
  NAND2X0 U9563 ( .IN1(n9771), .IN2(n9772), .QN(n9770) );
  XNOR2X1 U9564 ( .IN1(n9773), .IN2(n8977), .Q(n9772) );
  XNOR2X1 U9565 ( .IN1(n9774), .IN2(n9274), .Q(n9771) );
  XNOR2X1 U9566 ( .IN1(n8978), .IN2(n9775), .Q(n9769) );
  NOR2X0 U9567 ( .IN1(n9776), .IN2(n9777), .QN(n9767) );
  NAND2X0 U9568 ( .IN1(n9778), .IN2(n9779), .QN(n9777) );
  XOR2X1 U9569 ( .IN1(n9780), .IN2(n8980), .Q(n9779) );
  XNOR2X1 U9570 ( .IN1(n9781), .IN2(n9272), .Q(n9778) );
  XNOR2X1 U9571 ( .IN1(n9273), .IN2(n9782), .Q(n9776) );
  NAND2X0 U9572 ( .IN1(n9783), .IN2(n9784), .QN(n9765) );
  NOR2X0 U9573 ( .IN1(n9785), .IN2(n9786), .QN(n9784) );
  NAND2X0 U9574 ( .IN1(n9787), .IN2(n9753), .QN(n9786) );
  XNOR2X1 U9575 ( .IN1(n9788), .IN2(test_so36), .Q(n9785) );
  NOR2X0 U9576 ( .IN1(n9789), .IN2(n9790), .QN(n9783) );
  NAND2X0 U9577 ( .IN1(n9791), .IN2(n9792), .QN(n9790) );
  XOR2X1 U9578 ( .IN1(n9793), .IN2(n8390), .Q(n9792) );
  XNOR2X1 U9579 ( .IN1(n9794), .IN2(n8979), .Q(n9791) );
  XNOR2X1 U9580 ( .IN1(n8561), .IN2(n9795), .Q(n9789) );
  NOR2X0 U9581 ( .IN1(n9796), .IN2(n9797), .QN(n4276) );
  NOR2X0 U9582 ( .IN1(n9798), .IN2(n9799), .QN(n9797) );
  NOR2X0 U9583 ( .IN1(n9800), .IN2(n9801), .QN(n9796) );
  NAND2X0 U9584 ( .IN1(n9802), .IN2(n9803), .QN(n9801) );
  NOR2X0 U9585 ( .IN1(n9804), .IN2(n9805), .QN(n9803) );
  NAND2X0 U9586 ( .IN1(n9806), .IN2(n9807), .QN(n9805) );
  XNOR2X1 U9587 ( .IN1(n9808), .IN2(n8973), .Q(n9807) );
  XNOR2X1 U9588 ( .IN1(n9809), .IN2(n9267), .Q(n9806) );
  XNOR2X1 U9589 ( .IN1(n8976), .IN2(n9810), .Q(n9804) );
  NOR2X0 U9590 ( .IN1(n9811), .IN2(n9812), .QN(n9802) );
  NAND2X0 U9591 ( .IN1(n9813), .IN2(n9814), .QN(n9812) );
  XNOR2X1 U9592 ( .IN1(n9815), .IN2(n8975), .Q(n9814) );
  XNOR2X1 U9593 ( .IN1(n9816), .IN2(n8560), .Q(n9813) );
  XNOR2X1 U9594 ( .IN1(n8974), .IN2(n9817), .Q(n9811) );
  NAND2X0 U9595 ( .IN1(n9818), .IN2(n9819), .QN(n9800) );
  NOR2X0 U9596 ( .IN1(n9820), .IN2(n9821), .QN(n9819) );
  NAND2X0 U9597 ( .IN1(n9822), .IN2(n9753), .QN(n9821) );
  XNOR2X1 U9598 ( .IN1(n9270), .IN2(n9823), .Q(n9820) );
  NOR2X0 U9599 ( .IN1(n9824), .IN2(n9825), .QN(n9818) );
  NAND2X0 U9600 ( .IN1(n9826), .IN2(n9827), .QN(n9825) );
  XNOR2X1 U9601 ( .IN1(n9828), .IN2(n9265), .Q(n9827) );
  XNOR2X1 U9602 ( .IN1(n9829), .IN2(n9276), .Q(n9826) );
  XNOR2X1 U9603 ( .IN1(n8389), .IN2(n9830), .Q(n9824) );
  NOR2X0 U9604 ( .IN1(n9831), .IN2(n9832), .QN(n4275) );
  NOR2X0 U9605 ( .IN1(n9833), .IN2(n9834), .QN(n9832) );
  NOR2X0 U9606 ( .IN1(n9835), .IN2(n9836), .QN(n9831) );
  NAND2X0 U9607 ( .IN1(n9837), .IN2(n9838), .QN(n9836) );
  NOR2X0 U9608 ( .IN1(n9839), .IN2(n9840), .QN(n9838) );
  NAND2X0 U9609 ( .IN1(n9841), .IN2(n9842), .QN(n9840) );
  XNOR2X1 U9610 ( .IN1(n9843), .IN2(n8969), .Q(n9842) );
  XNOR2X1 U9611 ( .IN1(n9844), .IN2(g2129), .Q(n9841) );
  XNOR2X1 U9612 ( .IN1(n8972), .IN2(n9845), .Q(n9839) );
  NOR2X0 U9613 ( .IN1(n9846), .IN2(n9847), .QN(n9837) );
  NAND2X0 U9614 ( .IN1(n9848), .IN2(n9849), .QN(n9847) );
  XNOR2X1 U9615 ( .IN1(n9850), .IN2(n8971), .Q(n9849) );
  XNOR2X1 U9616 ( .IN1(n9851), .IN2(n8559), .Q(n9848) );
  XNOR2X1 U9617 ( .IN1(n8970), .IN2(n9852), .Q(n9846) );
  NAND2X0 U9618 ( .IN1(n9853), .IN2(n9854), .QN(n9835) );
  NOR2X0 U9619 ( .IN1(n9855), .IN2(n9856), .QN(n9854) );
  NAND2X0 U9620 ( .IN1(n9857), .IN2(n9753), .QN(n9856) );
  XNOR2X1 U9621 ( .IN1(n9858), .IN2(test_so78), .Q(n9855) );
  NOR2X0 U9622 ( .IN1(n9859), .IN2(n9860), .QN(n9853) );
  NAND2X0 U9623 ( .IN1(n9861), .IN2(n9862), .QN(n9860) );
  XNOR2X1 U9624 ( .IN1(n9863), .IN2(n8388), .Q(n9862) );
  XNOR2X1 U9625 ( .IN1(n9864), .IN2(g2147), .Q(n9861) );
  XNOR2X1 U9626 ( .IN1(n9277), .IN2(n9865), .Q(n9859) );
  NAND2X0 U9627 ( .IN1(n9866), .IN2(n9677), .QN(n4274) );
  INVX0 U9628 ( .INP(n9867), .ZN(n9677) );
  XOR2X1 U9629 ( .IN1(n4330), .IN2(g2950), .Q(n9866) );
  NAND2X0 U9630 ( .IN1(n9868), .IN2(n9869), .QN(n4273) );
  NAND2X0 U9631 ( .IN1(n9870), .IN2(n9871), .QN(n9869) );
  NAND2X0 U9632 ( .IN1(n4482), .IN2(n9872), .QN(n9870) );
  NAND2X0 U9633 ( .IN1(n2426), .IN2(n9873), .QN(n4272) );
  NAND2X0 U9634 ( .IN1(n9874), .IN2(n9875), .QN(n9873) );
  NOR2X0 U9635 ( .IN1(n9876), .IN2(n9877), .QN(n9874) );
  NOR2X0 U9636 ( .IN1(test_so27), .IN2(n9878), .QN(n9877) );
  NOR2X0 U9637 ( .IN1(n9879), .IN2(n9880), .QN(n9876) );
  NAND2X0 U9638 ( .IN1(n9881), .IN2(n9882), .QN(n4271) );
  NAND2X0 U9639 ( .IN1(n2446), .IN2(n9883), .QN(n9882) );
  NAND2X0 U9640 ( .IN1(n9884), .IN2(n9875), .QN(n9881) );
  NOR2X0 U9641 ( .IN1(n9885), .IN2(n9886), .QN(n9884) );
  NOR2X0 U9642 ( .IN1(n9878), .IN2(g536), .QN(n9886) );
  NOR2X0 U9643 ( .IN1(n9879), .IN2(n9887), .QN(n9885) );
  NAND2X0 U9644 ( .IN1(n9888), .IN2(n9889), .QN(n4270) );
  NAND2X0 U9645 ( .IN1(n2446), .IN2(n9890), .QN(n9889) );
  NAND2X0 U9646 ( .IN1(n9891), .IN2(n9875), .QN(n9888) );
  NOR2X0 U9647 ( .IN1(n9892), .IN2(n9893), .QN(n9891) );
  NOR2X0 U9648 ( .IN1(n9878), .IN2(g537), .QN(n9893) );
  NOR2X0 U9649 ( .IN1(n9879), .IN2(n9894), .QN(n9892) );
  NAND2X0 U9650 ( .IN1(n9895), .IN2(n9896), .QN(n4269) );
  NAND2X0 U9651 ( .IN1(n9897), .IN2(n9875), .QN(n9896) );
  NOR2X0 U9652 ( .IN1(n9898), .IN2(n9899), .QN(n9897) );
  NOR2X0 U9653 ( .IN1(n9878), .IN2(n8047), .QN(n9899) );
  NOR2X0 U9654 ( .IN1(n9879), .IN2(n9900), .QN(n9898) );
  NAND2X0 U9655 ( .IN1(n9901), .IN2(n2440), .QN(n4268) );
  NOR2X0 U9656 ( .IN1(n9902), .IN2(n9903), .QN(n9901) );
  NOR2X0 U9657 ( .IN1(n9904), .IN2(n9905), .QN(n9902) );
  NAND2X0 U9658 ( .IN1(n9906), .IN2(n9907), .QN(n9905) );
  NAND2X0 U9659 ( .IN1(n9908), .IN2(n9909), .QN(n9907) );
  INVX0 U9660 ( .INP(n9910), .ZN(n9908) );
  NAND2X0 U9661 ( .IN1(n9911), .IN2(DFF_445_n1), .QN(n9906) );
  NAND2X0 U9662 ( .IN1(n9912), .IN2(n2440), .QN(n4267) );
  NOR2X0 U9663 ( .IN1(n9913), .IN2(n9903), .QN(n9912) );
  NOR2X0 U9664 ( .IN1(n9904), .IN2(n9914), .QN(n9913) );
  NAND2X0 U9665 ( .IN1(n9915), .IN2(n9916), .QN(n9914) );
  INVX0 U9666 ( .INP(n9917), .ZN(n9916) );
  NOR2X0 U9667 ( .IN1(n9918), .IN2(n9879), .QN(n9917) );
  NAND2X0 U9668 ( .IN1(n9911), .IN2(DFF_446_n1), .QN(n9915) );
  NAND2X0 U9669 ( .IN1(n9895), .IN2(n9919), .QN(n4266) );
  NAND2X0 U9670 ( .IN1(n9920), .IN2(n9875), .QN(n9919) );
  NOR2X0 U9671 ( .IN1(n9921), .IN2(n9922), .QN(n9920) );
  NOR2X0 U9672 ( .IN1(n9878), .IN2(n8044), .QN(n9922) );
  NOR2X0 U9673 ( .IN1(n9879), .IN2(n9923), .QN(n9921) );
  NOR2X0 U9674 ( .IN1(n9903), .IN2(n9924), .QN(n9895) );
  INVX0 U9675 ( .INP(n9925), .ZN(n9924) );
  NAND2X0 U9676 ( .IN1(n2446), .IN2(n2445), .QN(n9925) );
  INVX0 U9677 ( .INP(n2426), .ZN(n9903) );
  NAND2X0 U9678 ( .IN1(n2426), .IN2(n9926), .QN(n4265) );
  NAND2X0 U9679 ( .IN1(n9927), .IN2(n9875), .QN(n9926) );
  NOR2X0 U9680 ( .IN1(n9928), .IN2(n9929), .QN(n9927) );
  NOR2X0 U9681 ( .IN1(n9878), .IN2(n8043), .QN(n9929) );
  INVX0 U9682 ( .INP(n9911), .ZN(n9878) );
  NOR2X0 U9683 ( .IN1(n9879), .IN2(n9930), .QN(n9928) );
  INVX0 U9684 ( .INP(n9909), .ZN(n9879) );
  NAND2X0 U9685 ( .IN1(DFF_1562_n1), .IN2(n9931), .QN(n4263) );
  NAND2X0 U9686 ( .IN1(n9932), .IN2(n9933), .QN(n4262) );
  XNOR2X1 U9687 ( .IN1(n4481), .IN2(n9934), .Q(n9932) );
  XNOR2X1 U9688 ( .IN1(n9935), .IN2(n9936), .Q(n4261) );
  INVX0 U9689 ( .INP(n9937), .ZN(n9936) );
  XNOR2X1 U9690 ( .IN1(n9938), .IN2(n9935), .Q(n4260) );
  NOR2X0 U9691 ( .IN1(g3231), .IN2(n16832), .QN(n9935) );
  NAND2X0 U9692 ( .IN1(n9939), .IN2(n9940), .QN(n4259) );
  NAND2X0 U9693 ( .IN1(test_so22), .IN2(n9941), .QN(n9940) );
  XOR2X1 U9694 ( .IN1(n9942), .IN2(n9943), .Q(n9941) );
  XOR2X1 U9695 ( .IN1(n9944), .IN2(n9945), .Q(n9943) );
  XOR2X1 U9696 ( .IN1(n9923), .IN2(n9930), .Q(n9945) );
  NAND2X0 U9697 ( .IN1(n9946), .IN2(n9947), .QN(n9930) );
  NOR2X0 U9698 ( .IN1(n9948), .IN2(n9949), .QN(n9946) );
  NOR2X0 U9699 ( .IN1(n9950), .IN2(n9951), .QN(n9949) );
  NOR2X0 U9700 ( .IN1(n9952), .IN2(n9953), .QN(n9948) );
  NAND2X0 U9701 ( .IN1(n9954), .IN2(n9955), .QN(n9923) );
  NOR2X0 U9702 ( .IN1(n9956), .IN2(n9957), .QN(n9954) );
  NOR2X0 U9703 ( .IN1(n9958), .IN2(n9959), .QN(n9957) );
  INVX0 U9704 ( .INP(n9960), .ZN(n9958) );
  NOR2X0 U9705 ( .IN1(n9961), .IN2(n9960), .QN(n9956) );
  XOR2X1 U9706 ( .IN1(n9910), .IN2(n9918), .Q(n9944) );
  NAND2X0 U9707 ( .IN1(n9962), .IN2(n9955), .QN(n9918) );
  NOR2X0 U9708 ( .IN1(n9963), .IN2(n9964), .QN(n9962) );
  NOR2X0 U9709 ( .IN1(n9965), .IN2(n9951), .QN(n9964) );
  NOR2X0 U9710 ( .IN1(n9952), .IN2(n9966), .QN(n9963) );
  NAND2X0 U9711 ( .IN1(n9967), .IN2(n9955), .QN(n9910) );
  NOR2X0 U9712 ( .IN1(n9968), .IN2(n9969), .QN(n9967) );
  NOR2X0 U9713 ( .IN1(n9970), .IN2(n9959), .QN(n9969) );
  NOR2X0 U9714 ( .IN1(n9961), .IN2(n9971), .QN(n9968) );
  XOR2X1 U9715 ( .IN1(n9972), .IN2(n9973), .Q(n9942) );
  XOR2X1 U9716 ( .IN1(n9894), .IN2(n9900), .Q(n9973) );
  NAND2X0 U9717 ( .IN1(n9974), .IN2(n9955), .QN(n9900) );
  NOR2X0 U9718 ( .IN1(n9975), .IN2(n9976), .QN(n9974) );
  NOR2X0 U9719 ( .IN1(n9977), .IN2(n9951), .QN(n9976) );
  NOR2X0 U9720 ( .IN1(n9952), .IN2(n9978), .QN(n9975) );
  NAND2X0 U9721 ( .IN1(n9979), .IN2(n9955), .QN(n9894) );
  NOR2X0 U9722 ( .IN1(n9980), .IN2(n9981), .QN(n9979) );
  NOR2X0 U9723 ( .IN1(n9982), .IN2(n9959), .QN(n9981) );
  INVX0 U9724 ( .INP(n9983), .ZN(n9982) );
  NOR2X0 U9725 ( .IN1(n9961), .IN2(n9983), .QN(n9980) );
  XOR2X1 U9726 ( .IN1(n9880), .IN2(n9887), .Q(n9972) );
  NAND2X0 U9727 ( .IN1(n9984), .IN2(n9947), .QN(n9887) );
  NOR2X0 U9728 ( .IN1(n9985), .IN2(n9986), .QN(n9984) );
  NOR2X0 U9729 ( .IN1(n9987), .IN2(n9951), .QN(n9986) );
  NOR2X0 U9730 ( .IN1(n9952), .IN2(n9988), .QN(n9985) );
  NAND2X0 U9731 ( .IN1(n9989), .IN2(n9990), .QN(n9880) );
  NOR2X0 U9732 ( .IN1(n9991), .IN2(n9992), .QN(n9989) );
  NOR2X0 U9733 ( .IN1(n9993), .IN2(n9959), .QN(n9992) );
  NOR2X0 U9734 ( .IN1(n9961), .IN2(n9994), .QN(n9991) );
  NOR2X0 U9735 ( .IN1(n9995), .IN2(n9996), .QN(n9939) );
  NOR2X0 U9736 ( .IN1(n4360), .IN2(n9997), .QN(n9996) );
  XNOR2X1 U9737 ( .IN1(n9890), .IN2(n9883), .Q(n9997) );
  NAND2X0 U9738 ( .IN1(n9998), .IN2(n9947), .QN(n9883) );
  INVX0 U9739 ( .INP(n9999), .ZN(n9947) );
  NAND2X0 U9740 ( .IN1(n9955), .IN2(n506), .QN(n9999) );
  NAND2X0 U9741 ( .IN1(n10000), .IN2(n10001), .QN(n506) );
  NOR2X0 U9742 ( .IN1(n10002), .IN2(n10003), .QN(n9998) );
  NOR2X0 U9743 ( .IN1(n10004), .IN2(n9951), .QN(n10003) );
  NAND2X0 U9744 ( .IN1(n9952), .IN2(n10005), .QN(n9951) );
  NOR2X0 U9745 ( .IN1(n9952), .IN2(n10006), .QN(n10002) );
  NAND2X0 U9746 ( .IN1(n10007), .IN2(n9990), .QN(n9890) );
  INVX0 U9747 ( .INP(n10008), .ZN(n9990) );
  NAND2X0 U9748 ( .IN1(n9955), .IN2(n10009), .QN(n10008) );
  NAND2X0 U9749 ( .IN1(n10000), .IN2(n10010), .QN(n10009) );
  NOR2X0 U9750 ( .IN1(n9714), .IN2(n4541), .QN(n9955) );
  NOR2X0 U9751 ( .IN1(n10011), .IN2(n10012), .QN(n10007) );
  NOR2X0 U9752 ( .IN1(n10013), .IN2(n9959), .QN(n10012) );
  NAND2X0 U9753 ( .IN1(n9961), .IN2(n10005), .QN(n9959) );
  NOR2X0 U9754 ( .IN1(n9961), .IN2(n10014), .QN(n10011) );
  NOR2X0 U9755 ( .IN1(n10015), .IN2(n10016), .QN(n9995) );
  NAND2X0 U9756 ( .IN1(n9875), .IN2(n9911), .QN(n10016) );
  NOR2X0 U9757 ( .IN1(n9909), .IN2(n9714), .QN(n9911) );
  NAND2X0 U9758 ( .IN1(n10017), .IN2(n10018), .QN(n9714) );
  NOR2X0 U9759 ( .IN1(g563), .IN2(n10019), .QN(n10018) );
  NOR2X0 U9760 ( .IN1(n4298), .IN2(g499), .QN(n10019) );
  NOR2X0 U9761 ( .IN1(g559), .IN2(g21851), .QN(n10017) );
  NAND2X0 U9762 ( .IN1(n10020), .IN2(n10021), .QN(n10015) );
  NAND2X0 U9763 ( .IN1(n16816), .IN2(n10022), .QN(n10021) );
  NAND2X0 U9764 ( .IN1(n4492), .IN2(g3229), .QN(n10020) );
  NAND2X0 U9765 ( .IN1(n10023), .IN2(n10024), .QN(n4258) );
  NAND2X0 U9766 ( .IN1(n2361), .IN2(n10025), .QN(n10024) );
  NAND2X0 U9767 ( .IN1(n10026), .IN2(n10027), .QN(n10023) );
  NOR2X0 U9768 ( .IN1(n10028), .IN2(n10029), .QN(n10026) );
  NOR2X0 U9769 ( .IN1(n10030), .IN2(g2611), .QN(n10029) );
  NOR2X0 U9770 ( .IN1(n10031), .IN2(n10032), .QN(n10028) );
  NAND2X0 U9771 ( .IN1(n10033), .IN2(n2375), .QN(n4257) );
  NOR2X0 U9772 ( .IN1(n10034), .IN2(n10035), .QN(n10033) );
  NOR2X0 U9773 ( .IN1(n10036), .IN2(n10037), .QN(n10035) );
  NAND2X0 U9774 ( .IN1(n10038), .IN2(n10039), .QN(n10037) );
  NAND2X0 U9775 ( .IN1(n10040), .IN2(n10041), .QN(n10039) );
  NAND2X0 U9776 ( .IN1(n10042), .IN2(DFF_1495_n1), .QN(n10038) );
  NAND2X0 U9777 ( .IN1(n10043), .IN2(n10044), .QN(n4256) );
  NAND2X0 U9778 ( .IN1(n10045), .IN2(n10027), .QN(n10044) );
  NOR2X0 U9779 ( .IN1(n10046), .IN2(n10047), .QN(n10045) );
  NOR2X0 U9780 ( .IN1(n10030), .IN2(n7920), .QN(n10047) );
  NOR2X0 U9781 ( .IN1(n10031), .IN2(n10048), .QN(n10046) );
  NAND2X0 U9782 ( .IN1(n10049), .IN2(n2375), .QN(n4255) );
  NOR2X0 U9783 ( .IN1(n10034), .IN2(n10050), .QN(n10049) );
  NOR2X0 U9784 ( .IN1(n10036), .IN2(n10051), .QN(n10050) );
  NAND2X0 U9785 ( .IN1(n10052), .IN2(n10053), .QN(n10051) );
  NAND2X0 U9786 ( .IN1(n10054), .IN2(n10041), .QN(n10053) );
  INVX0 U9787 ( .INP(n10055), .ZN(n10054) );
  NAND2X0 U9788 ( .IN1(n10042), .IN2(DFF_1496_n1), .QN(n10052) );
  NAND2X0 U9789 ( .IN1(n10056), .IN2(n10057), .QN(n4254) );
  NAND2X0 U9790 ( .IN1(n10058), .IN2(n10027), .QN(n10057) );
  NOR2X0 U9791 ( .IN1(n10059), .IN2(n10060), .QN(n10058) );
  NOR2X0 U9792 ( .IN1(n10030), .IN2(n7925), .QN(n10060) );
  NOR2X0 U9793 ( .IN1(n10031), .IN2(n10061), .QN(n10059) );
  NAND2X0 U9794 ( .IN1(n10062), .IN2(n10063), .QN(n4253) );
  NAND2X0 U9795 ( .IN1(n2361), .IN2(n10064), .QN(n10063) );
  NAND2X0 U9796 ( .IN1(n10065), .IN2(n10027), .QN(n10062) );
  NOR2X0 U9797 ( .IN1(n10066), .IN2(n10067), .QN(n10065) );
  NOR2X0 U9798 ( .IN1(test_so91), .IN2(n10030), .QN(n10067) );
  NOR2X0 U9799 ( .IN1(n10031), .IN2(n10068), .QN(n10066) );
  NAND2X0 U9800 ( .IN1(n10056), .IN2(n10069), .QN(n4252) );
  NAND2X0 U9801 ( .IN1(n10070), .IN2(n10027), .QN(n10069) );
  NOR2X0 U9802 ( .IN1(n10071), .IN2(n10072), .QN(n10070) );
  NOR2X0 U9803 ( .IN1(n10030), .IN2(n7922), .QN(n10072) );
  NOR2X0 U9804 ( .IN1(n10031), .IN2(n10073), .QN(n10071) );
  NOR2X0 U9805 ( .IN1(n10034), .IN2(n10074), .QN(n10056) );
  INVX0 U9806 ( .INP(n10075), .ZN(n10074) );
  NAND2X0 U9807 ( .IN1(n2361), .IN2(n2374), .QN(n10075) );
  INVX0 U9808 ( .INP(n10043), .ZN(n10034) );
  NAND2X0 U9809 ( .IN1(n10043), .IN2(n10076), .QN(n4251) );
  NAND2X0 U9810 ( .IN1(n10077), .IN2(n10027), .QN(n10076) );
  NOR2X0 U9811 ( .IN1(n10078), .IN2(n10079), .QN(n10077) );
  NOR2X0 U9812 ( .IN1(n10030), .IN2(n7921), .QN(n10079) );
  INVX0 U9813 ( .INP(n10042), .ZN(n10030) );
  NOR2X0 U9814 ( .IN1(n10031), .IN2(n10080), .QN(n10078) );
  INVX0 U9815 ( .INP(n10041), .ZN(n10031) );
  NAND2X0 U9816 ( .IN1(n2361), .IN2(n10081), .QN(n10043) );
  NAND2X0 U9817 ( .IN1(n10082), .IN2(n10083), .QN(n4250) );
  NAND2X0 U9818 ( .IN1(n10084), .IN2(g2631), .QN(n10083) );
  XOR2X1 U9819 ( .IN1(n10025), .IN2(n10064), .Q(n10084) );
  NAND2X0 U9820 ( .IN1(n10085), .IN2(n10086), .QN(n10064) );
  NOR2X0 U9821 ( .IN1(n10087), .IN2(n10088), .QN(n10085) );
  NOR2X0 U9822 ( .IN1(n10089), .IN2(n10090), .QN(n10088) );
  NOR2X0 U9823 ( .IN1(n10091), .IN2(n10092), .QN(n10087) );
  NAND2X0 U9824 ( .IN1(n10093), .IN2(n10094), .QN(n10025) );
  NOR2X0 U9825 ( .IN1(n10095), .IN2(n10096), .QN(n10093) );
  NOR2X0 U9826 ( .IN1(n10097), .IN2(n10098), .QN(n10096) );
  INVX0 U9827 ( .INP(n10099), .ZN(n10097) );
  NOR2X0 U9828 ( .IN1(n10100), .IN2(n10099), .QN(n10095) );
  NOR2X0 U9829 ( .IN1(n10101), .IN2(n10102), .QN(n10082) );
  NOR2X0 U9830 ( .IN1(n4303), .IN2(n10103), .QN(n10102) );
  XOR2X1 U9831 ( .IN1(n10104), .IN2(n10105), .Q(n10103) );
  XOR2X1 U9832 ( .IN1(n10106), .IN2(n10107), .Q(n10105) );
  XNOR2X1 U9833 ( .IN1(n10080), .IN2(n10073), .Q(n10107) );
  NAND2X0 U9834 ( .IN1(n10108), .IN2(n10109), .QN(n10073) );
  NOR2X0 U9835 ( .IN1(n10110), .IN2(n10111), .QN(n10108) );
  NOR2X0 U9836 ( .IN1(n10112), .IN2(n10098), .QN(n10111) );
  INVX0 U9837 ( .INP(n10113), .ZN(n10112) );
  NOR2X0 U9838 ( .IN1(n10100), .IN2(n10113), .QN(n10110) );
  NAND2X0 U9839 ( .IN1(n10114), .IN2(n10086), .QN(n10080) );
  NOR2X0 U9840 ( .IN1(n10115), .IN2(n10116), .QN(n10114) );
  NOR2X0 U9841 ( .IN1(n10117), .IN2(n10090), .QN(n10116) );
  NOR2X0 U9842 ( .IN1(n10091), .IN2(n10118), .QN(n10115) );
  XNOR2X1 U9843 ( .IN1(n10068), .IN2(n10061), .Q(n10106) );
  NAND2X0 U9844 ( .IN1(n10119), .IN2(n10109), .QN(n10061) );
  NOR2X0 U9845 ( .IN1(n10120), .IN2(n10121), .QN(n10119) );
  NOR2X0 U9846 ( .IN1(n10122), .IN2(n10090), .QN(n10121) );
  NOR2X0 U9847 ( .IN1(n10091), .IN2(n10123), .QN(n10120) );
  NAND2X0 U9848 ( .IN1(n10124), .IN2(n10086), .QN(n10068) );
  INVX0 U9849 ( .INP(n10125), .ZN(n10086) );
  NAND2X0 U9850 ( .IN1(n10109), .IN2(n1458), .QN(n10125) );
  NOR2X0 U9851 ( .IN1(n10126), .IN2(n10127), .QN(n10124) );
  NOR2X0 U9852 ( .IN1(n10128), .IN2(n10090), .QN(n10127) );
  NOR2X0 U9853 ( .IN1(n10091), .IN2(n10129), .QN(n10126) );
  XOR2X1 U9854 ( .IN1(n10130), .IN2(n10131), .Q(n10104) );
  XNOR2X1 U9855 ( .IN1(n10032), .IN2(n10040), .Q(n10131) );
  INVX0 U9856 ( .INP(n10132), .ZN(n10040) );
  NAND2X0 U9857 ( .IN1(n10133), .IN2(n10109), .QN(n10132) );
  NOR2X0 U9858 ( .IN1(n10134), .IN2(n10135), .QN(n10133) );
  NOR2X0 U9859 ( .IN1(n10136), .IN2(n10098), .QN(n10135) );
  NOR2X0 U9860 ( .IN1(n10100), .IN2(n10137), .QN(n10134) );
  NAND2X0 U9861 ( .IN1(n10138), .IN2(n10109), .QN(n10032) );
  NOR2X0 U9862 ( .IN1(n10139), .IN2(n10140), .QN(n10138) );
  NOR2X0 U9863 ( .IN1(n10141), .IN2(n10098), .QN(n10140) );
  INVX0 U9864 ( .INP(n10142), .ZN(n10141) );
  NOR2X0 U9865 ( .IN1(n10100), .IN2(n10142), .QN(n10139) );
  XNOR2X1 U9866 ( .IN1(n10048), .IN2(n10055), .Q(n10130) );
  NAND2X0 U9867 ( .IN1(n10143), .IN2(n10109), .QN(n10055) );
  NOR2X0 U9868 ( .IN1(n10144), .IN2(n10145), .QN(n10143) );
  NOR2X0 U9869 ( .IN1(n10146), .IN2(n10090), .QN(n10145) );
  NAND2X0 U9870 ( .IN1(n10091), .IN2(n10147), .QN(n10090) );
  NOR2X0 U9871 ( .IN1(n10091), .IN2(n10148), .QN(n10144) );
  NAND2X0 U9872 ( .IN1(n10149), .IN2(n10094), .QN(n10048) );
  INVX0 U9873 ( .INP(n10150), .ZN(n10094) );
  NAND2X0 U9874 ( .IN1(n10109), .IN2(n10151), .QN(n10150) );
  NAND2X0 U9875 ( .IN1(n10152), .IN2(n10153), .QN(n10151) );
  NOR2X0 U9876 ( .IN1(n10081), .IN2(n4543), .QN(n10109) );
  NOR2X0 U9877 ( .IN1(n10154), .IN2(n10155), .QN(n10149) );
  NOR2X0 U9878 ( .IN1(n10156), .IN2(n10098), .QN(n10155) );
  NAND2X0 U9879 ( .IN1(n10100), .IN2(n10147), .QN(n10098) );
  NOR2X0 U9880 ( .IN1(n10100), .IN2(n10157), .QN(n10154) );
  NOR2X0 U9881 ( .IN1(n10158), .IN2(n10159), .QN(n10101) );
  NAND2X0 U9882 ( .IN1(n10027), .IN2(n10042), .QN(n10159) );
  NOR2X0 U9883 ( .IN1(n10081), .IN2(n10041), .QN(n10042) );
  NAND2X0 U9884 ( .IN1(n10160), .IN2(n9035), .QN(n10081) );
  NOR2X0 U9885 ( .IN1(g2637), .IN2(g30072), .QN(n10160) );
  NAND2X0 U9886 ( .IN1(n10161), .IN2(n10162), .QN(n10158) );
  NAND2X0 U9887 ( .IN1(n16817), .IN2(n10022), .QN(n10162) );
  NAND2X0 U9888 ( .IN1(n4490), .IN2(g3229), .QN(n10161) );
  NAND2X0 U9889 ( .IN1(n10163), .IN2(n10164), .QN(n4249) );
  NAND2X0 U9890 ( .IN1(n2289), .IN2(n10165), .QN(n10164) );
  NAND2X0 U9891 ( .IN1(n10166), .IN2(n10167), .QN(n10163) );
  NOR2X0 U9892 ( .IN1(n10168), .IN2(n10169), .QN(n10166) );
  NOR2X0 U9893 ( .IN1(n10170), .IN2(g1917), .QN(n10169) );
  NOR2X0 U9894 ( .IN1(n10171), .IN2(n10172), .QN(n10168) );
  NAND2X0 U9895 ( .IN1(n10173), .IN2(n2303), .QN(n4248) );
  NOR2X0 U9896 ( .IN1(n10174), .IN2(n10175), .QN(n10173) );
  NOR2X0 U9897 ( .IN1(n10176), .IN2(n10177), .QN(n10174) );
  NAND2X0 U9898 ( .IN1(n10178), .IN2(n10179), .QN(n10177) );
  NAND2X0 U9899 ( .IN1(n10180), .IN2(n10181), .QN(n10179) );
  NAND2X0 U9900 ( .IN1(n10182), .IN2(DFF_1145_n1), .QN(n10178) );
  NAND2X0 U9901 ( .IN1(n2275), .IN2(n10183), .QN(n4247) );
  NAND2X0 U9902 ( .IN1(n10184), .IN2(n10167), .QN(n10183) );
  NOR2X0 U9903 ( .IN1(n10185), .IN2(n10186), .QN(n10184) );
  NOR2X0 U9904 ( .IN1(n10170), .IN2(n7962), .QN(n10186) );
  NOR2X0 U9905 ( .IN1(n10171), .IN2(n10187), .QN(n10185) );
  NAND2X0 U9906 ( .IN1(n10188), .IN2(n2303), .QN(n4246) );
  NOR2X0 U9907 ( .IN1(n10189), .IN2(n10175), .QN(n10188) );
  NOR2X0 U9908 ( .IN1(n10176), .IN2(n10190), .QN(n10189) );
  NAND2X0 U9909 ( .IN1(n10191), .IN2(n10192), .QN(n10190) );
  NAND2X0 U9910 ( .IN1(n10193), .IN2(n10181), .QN(n10192) );
  INVX0 U9911 ( .INP(n10194), .ZN(n10193) );
  NAND2X0 U9912 ( .IN1(n10182), .IN2(DFF_1146_n1), .QN(n10191) );
  NAND2X0 U9913 ( .IN1(n10195), .IN2(n10196), .QN(n4245) );
  NAND2X0 U9914 ( .IN1(n10197), .IN2(n10167), .QN(n10196) );
  NOR2X0 U9915 ( .IN1(n10198), .IN2(n10199), .QN(n10197) );
  NOR2X0 U9916 ( .IN1(n10170), .IN2(n7967), .QN(n10199) );
  NOR2X0 U9917 ( .IN1(n10171), .IN2(n10200), .QN(n10198) );
  NAND2X0 U9918 ( .IN1(n10201), .IN2(n10202), .QN(n4244) );
  NAND2X0 U9919 ( .IN1(n2289), .IN2(n10203), .QN(n10202) );
  NAND2X0 U9920 ( .IN1(n10204), .IN2(n10167), .QN(n10201) );
  NOR2X0 U9921 ( .IN1(n10205), .IN2(n10206), .QN(n10204) );
  NOR2X0 U9922 ( .IN1(n10170), .IN2(g1916), .QN(n10206) );
  NOR2X0 U9923 ( .IN1(n10171), .IN2(n10207), .QN(n10205) );
  NAND2X0 U9924 ( .IN1(n10195), .IN2(n10208), .QN(n4243) );
  NAND2X0 U9925 ( .IN1(n10209), .IN2(n10167), .QN(n10208) );
  NOR2X0 U9926 ( .IN1(n10210), .IN2(n10211), .QN(n10209) );
  NOR2X0 U9927 ( .IN1(n10170), .IN2(n7964), .QN(n10211) );
  NOR2X0 U9928 ( .IN1(n10171), .IN2(n10212), .QN(n10210) );
  NOR2X0 U9929 ( .IN1(n10175), .IN2(n10213), .QN(n10195) );
  INVX0 U9930 ( .INP(n10214), .ZN(n10213) );
  NAND2X0 U9931 ( .IN1(n2289), .IN2(n2302), .QN(n10214) );
  INVX0 U9932 ( .INP(n2275), .ZN(n10175) );
  NAND2X0 U9933 ( .IN1(n2275), .IN2(n10215), .QN(n4242) );
  NAND2X0 U9934 ( .IN1(n10216), .IN2(n10167), .QN(n10215) );
  NOR2X0 U9935 ( .IN1(n10217), .IN2(n10218), .QN(n10216) );
  NOR2X0 U9936 ( .IN1(n10170), .IN2(n7963), .QN(n10218) );
  INVX0 U9937 ( .INP(n10182), .ZN(n10170) );
  NOR2X0 U9938 ( .IN1(n10171), .IN2(n10219), .QN(n10217) );
  INVX0 U9939 ( .INP(n10181), .ZN(n10171) );
  NAND2X0 U9940 ( .IN1(n10220), .IN2(n10221), .QN(n4241) );
  NAND2X0 U9941 ( .IN1(n10222), .IN2(g1937), .QN(n10221) );
  XOR2X1 U9942 ( .IN1(n10165), .IN2(n10203), .Q(n10222) );
  NAND2X0 U9943 ( .IN1(n10223), .IN2(n10224), .QN(n10203) );
  NOR2X0 U9944 ( .IN1(n10225), .IN2(n10226), .QN(n10223) );
  NOR2X0 U9945 ( .IN1(n10227), .IN2(n10228), .QN(n10226) );
  NOR2X0 U9946 ( .IN1(n10229), .IN2(n10230), .QN(n10225) );
  NAND2X0 U9947 ( .IN1(n10231), .IN2(n10232), .QN(n10165) );
  NOR2X0 U9948 ( .IN1(n10233), .IN2(n10234), .QN(n10231) );
  NOR2X0 U9949 ( .IN1(n10235), .IN2(n10236), .QN(n10234) );
  NOR2X0 U9950 ( .IN1(n10237), .IN2(n10238), .QN(n10233) );
  NOR2X0 U9951 ( .IN1(n10239), .IN2(n10240), .QN(n10220) );
  NOR2X0 U9952 ( .IN1(n4297), .IN2(n10241), .QN(n10240) );
  XOR2X1 U9953 ( .IN1(n10242), .IN2(n10243), .Q(n10241) );
  XOR2X1 U9954 ( .IN1(n10244), .IN2(n10245), .Q(n10243) );
  XNOR2X1 U9955 ( .IN1(n10219), .IN2(n10212), .Q(n10245) );
  NAND2X0 U9956 ( .IN1(n10246), .IN2(n10247), .QN(n10212) );
  NOR2X0 U9957 ( .IN1(n10248), .IN2(n10249), .QN(n10246) );
  NOR2X0 U9958 ( .IN1(n10250), .IN2(n10236), .QN(n10249) );
  NOR2X0 U9959 ( .IN1(n10237), .IN2(n10251), .QN(n10248) );
  NAND2X0 U9960 ( .IN1(n10252), .IN2(n10224), .QN(n10219) );
  NOR2X0 U9961 ( .IN1(n10253), .IN2(n10254), .QN(n10252) );
  NOR2X0 U9962 ( .IN1(n10255), .IN2(n10228), .QN(n10254) );
  NOR2X0 U9963 ( .IN1(n10229), .IN2(n10256), .QN(n10253) );
  XNOR2X1 U9964 ( .IN1(n10207), .IN2(n10200), .Q(n10244) );
  NAND2X0 U9965 ( .IN1(n10257), .IN2(n10247), .QN(n10200) );
  NOR2X0 U9966 ( .IN1(n10258), .IN2(n10259), .QN(n10257) );
  NOR2X0 U9967 ( .IN1(n10260), .IN2(n10228), .QN(n10259) );
  INVX0 U9968 ( .INP(n10261), .ZN(n10260) );
  NOR2X0 U9969 ( .IN1(n10229), .IN2(n10261), .QN(n10258) );
  NAND2X0 U9970 ( .IN1(n10262), .IN2(n10224), .QN(n10207) );
  INVX0 U9971 ( .INP(n10263), .ZN(n10224) );
  NAND2X0 U9972 ( .IN1(n10247), .IN2(n10264), .QN(n10263) );
  NAND2X0 U9973 ( .IN1(n10265), .IN2(n10266), .QN(n10264) );
  NOR2X0 U9974 ( .IN1(n10267), .IN2(n10268), .QN(n10262) );
  NOR2X0 U9975 ( .IN1(n10269), .IN2(n10228), .QN(n10268) );
  NOR2X0 U9976 ( .IN1(n10229), .IN2(n10270), .QN(n10267) );
  XOR2X1 U9977 ( .IN1(n10271), .IN2(n10272), .Q(n10242) );
  XNOR2X1 U9978 ( .IN1(n10172), .IN2(n10180), .Q(n10272) );
  INVX0 U9979 ( .INP(n10273), .ZN(n10180) );
  NAND2X0 U9980 ( .IN1(n10274), .IN2(n10247), .QN(n10273) );
  NOR2X0 U9981 ( .IN1(n10275), .IN2(n10276), .QN(n10274) );
  NOR2X0 U9982 ( .IN1(n10277), .IN2(n10236), .QN(n10276) );
  INVX0 U9983 ( .INP(n10278), .ZN(n10277) );
  NOR2X0 U9984 ( .IN1(n10237), .IN2(n10278), .QN(n10275) );
  NAND2X0 U9985 ( .IN1(n10279), .IN2(n10247), .QN(n10172) );
  NOR2X0 U9986 ( .IN1(n10280), .IN2(n10281), .QN(n10279) );
  NOR2X0 U9987 ( .IN1(n10282), .IN2(n10236), .QN(n10281) );
  NOR2X0 U9988 ( .IN1(n10237), .IN2(n10283), .QN(n10280) );
  XNOR2X1 U9989 ( .IN1(n10187), .IN2(n10194), .Q(n10271) );
  NAND2X0 U9990 ( .IN1(n10284), .IN2(n10247), .QN(n10194) );
  NOR2X0 U9991 ( .IN1(n10285), .IN2(n10286), .QN(n10284) );
  NOR2X0 U9992 ( .IN1(n10287), .IN2(n10228), .QN(n10286) );
  NAND2X0 U9993 ( .IN1(n10229), .IN2(n10288), .QN(n10228) );
  INVX0 U9994 ( .INP(n10289), .ZN(n10287) );
  NOR2X0 U9995 ( .IN1(n10229), .IN2(n10289), .QN(n10285) );
  NAND2X0 U9996 ( .IN1(n10290), .IN2(n10232), .QN(n10187) );
  INVX0 U9997 ( .INP(n10291), .ZN(n10232) );
  NAND2X0 U9998 ( .IN1(n10247), .IN2(n10292), .QN(n10291) );
  NAND2X0 U9999 ( .IN1(n10265), .IN2(n10293), .QN(n10292) );
  NOR2X0 U10000 ( .IN1(n9706), .IN2(n4545), .QN(n10247) );
  NOR2X0 U10001 ( .IN1(n10294), .IN2(n10295), .QN(n10290) );
  NOR2X0 U10002 ( .IN1(n10296), .IN2(n10236), .QN(n10295) );
  NAND2X0 U10003 ( .IN1(n10237), .IN2(n10288), .QN(n10236) );
  NOR2X0 U10004 ( .IN1(n10237), .IN2(n10297), .QN(n10294) );
  NOR2X0 U10005 ( .IN1(n10298), .IN2(n10299), .QN(n10239) );
  NAND2X0 U10006 ( .IN1(n10167), .IN2(n10182), .QN(n10299) );
  NOR2X0 U10007 ( .IN1(n9706), .IN2(n10181), .QN(n10182) );
  NAND2X0 U10008 ( .IN1(n10300), .IN2(n9036), .QN(n9706) );
  NOR2X0 U10009 ( .IN1(g1943), .IN2(n532), .QN(n10300) );
  NAND2X0 U10010 ( .IN1(n10301), .IN2(n10302), .QN(n10298) );
  INVX0 U10011 ( .INP(n10303), .ZN(n10302) );
  NOR2X0 U10012 ( .IN1(n10022), .IN2(test_so69), .QN(n10303) );
  NAND2X0 U10013 ( .IN1(n16818), .IN2(n10022), .QN(n10301) );
  NAND2X0 U10014 ( .IN1(n10304), .IN2(n10305), .QN(n4240) );
  NAND2X0 U10015 ( .IN1(n2217), .IN2(n10306), .QN(n10305) );
  NAND2X0 U10016 ( .IN1(n10307), .IN2(n10308), .QN(n10304) );
  NOR2X0 U10017 ( .IN1(n10309), .IN2(n10310), .QN(n10307) );
  NOR2X0 U10018 ( .IN1(n10311), .IN2(g1223), .QN(n10310) );
  NOR2X0 U10019 ( .IN1(n10312), .IN2(n10313), .QN(n10309) );
  NAND2X0 U10020 ( .IN1(n10314), .IN2(n2231), .QN(n4239) );
  NOR2X0 U10021 ( .IN1(n10315), .IN2(n10316), .QN(n10314) );
  NOR2X0 U10022 ( .IN1(n10317), .IN2(n10318), .QN(n10316) );
  NAND2X0 U10023 ( .IN1(n10319), .IN2(n10320), .QN(n10318) );
  NAND2X0 U10024 ( .IN1(n10321), .IN2(n10322), .QN(n10320) );
  NAND2X0 U10025 ( .IN1(n10323), .IN2(DFF_795_n1), .QN(n10319) );
  NAND2X0 U10026 ( .IN1(n10324), .IN2(n10325), .QN(n4238) );
  NAND2X0 U10027 ( .IN1(n10326), .IN2(n10308), .QN(n10325) );
  NOR2X0 U10028 ( .IN1(n10327), .IN2(n10328), .QN(n10326) );
  NOR2X0 U10029 ( .IN1(n10311), .IN2(n8003), .QN(n10328) );
  NOR2X0 U10030 ( .IN1(n10312), .IN2(n10329), .QN(n10327) );
  NAND2X0 U10031 ( .IN1(n10330), .IN2(n2231), .QN(n4237) );
  NOR2X0 U10032 ( .IN1(n10315), .IN2(n10331), .QN(n10330) );
  NOR2X0 U10033 ( .IN1(n10317), .IN2(n10332), .QN(n10331) );
  NAND2X0 U10034 ( .IN1(n10333), .IN2(n10334), .QN(n10332) );
  NAND2X0 U10035 ( .IN1(n10335), .IN2(n10322), .QN(n10334) );
  INVX0 U10036 ( .INP(n10336), .ZN(n10335) );
  NAND2X0 U10037 ( .IN1(n10323), .IN2(DFF_796_n1), .QN(n10333) );
  NAND2X0 U10038 ( .IN1(n10337), .IN2(n10338), .QN(n4236) );
  NAND2X0 U10039 ( .IN1(n10339), .IN2(n10308), .QN(n10338) );
  NOR2X0 U10040 ( .IN1(n10340), .IN2(n10341), .QN(n10339) );
  NOR2X0 U10041 ( .IN1(n10311), .IN2(n8008), .QN(n10341) );
  NOR2X0 U10042 ( .IN1(n10312), .IN2(n10342), .QN(n10340) );
  NAND2X0 U10043 ( .IN1(n10343), .IN2(n10344), .QN(n4235) );
  NAND2X0 U10044 ( .IN1(n2217), .IN2(n10345), .QN(n10344) );
  NAND2X0 U10045 ( .IN1(n10346), .IN2(n10308), .QN(n10343) );
  NOR2X0 U10046 ( .IN1(n10347), .IN2(n10348), .QN(n10346) );
  NOR2X0 U10047 ( .IN1(n10311), .IN2(g1222), .QN(n10348) );
  NOR2X0 U10048 ( .IN1(n10312), .IN2(n10349), .QN(n10347) );
  NAND2X0 U10049 ( .IN1(n10337), .IN2(n10350), .QN(n4234) );
  NAND2X0 U10050 ( .IN1(n10351), .IN2(n10308), .QN(n10350) );
  NOR2X0 U10051 ( .IN1(n10352), .IN2(n10353), .QN(n10351) );
  NOR2X0 U10052 ( .IN1(n10311), .IN2(n8005), .QN(n10353) );
  NOR2X0 U10053 ( .IN1(n10312), .IN2(n10354), .QN(n10352) );
  NOR2X0 U10054 ( .IN1(n10315), .IN2(n10355), .QN(n10337) );
  INVX0 U10055 ( .INP(n10356), .ZN(n10355) );
  NAND2X0 U10056 ( .IN1(n2217), .IN2(n2230), .QN(n10356) );
  INVX0 U10057 ( .INP(n10324), .ZN(n10315) );
  NAND2X0 U10058 ( .IN1(n10324), .IN2(n10357), .QN(n4233) );
  NAND2X0 U10059 ( .IN1(n10358), .IN2(n10308), .QN(n10357) );
  NOR2X0 U10060 ( .IN1(n10359), .IN2(n10360), .QN(n10358) );
  NOR2X0 U10061 ( .IN1(n10311), .IN2(n8004), .QN(n10360) );
  INVX0 U10062 ( .INP(n10323), .ZN(n10311) );
  NOR2X0 U10063 ( .IN1(n10312), .IN2(n10361), .QN(n10359) );
  INVX0 U10064 ( .INP(n10322), .ZN(n10312) );
  NAND2X0 U10065 ( .IN1(n2217), .IN2(n10362), .QN(n10324) );
  NAND2X0 U10066 ( .IN1(n10363), .IN2(n10364), .QN(n4232) );
  NAND2X0 U10067 ( .IN1(n10365), .IN2(g1243), .QN(n10364) );
  XOR2X1 U10068 ( .IN1(n10306), .IN2(n10345), .Q(n10365) );
  NAND2X0 U10069 ( .IN1(n10366), .IN2(n10367), .QN(n10345) );
  NOR2X0 U10070 ( .IN1(n10368), .IN2(n10369), .QN(n10366) );
  NOR2X0 U10071 ( .IN1(n10370), .IN2(n10371), .QN(n10369) );
  NOR2X0 U10072 ( .IN1(n10372), .IN2(n10373), .QN(n10368) );
  NAND2X0 U10073 ( .IN1(n10374), .IN2(n10375), .QN(n10306) );
  NOR2X0 U10074 ( .IN1(n10376), .IN2(n10377), .QN(n10374) );
  NOR2X0 U10075 ( .IN1(n10378), .IN2(n10379), .QN(n10377) );
  NOR2X0 U10076 ( .IN1(n10380), .IN2(n10381), .QN(n10376) );
  NOR2X0 U10077 ( .IN1(n10382), .IN2(n10383), .QN(n10363) );
  NOR2X0 U10078 ( .IN1(n4304), .IN2(n10384), .QN(n10383) );
  XOR2X1 U10079 ( .IN1(n10385), .IN2(n10386), .Q(n10384) );
  XOR2X1 U10080 ( .IN1(n10387), .IN2(n10388), .Q(n10386) );
  XNOR2X1 U10081 ( .IN1(n10361), .IN2(n10354), .Q(n10388) );
  NAND2X0 U10082 ( .IN1(n10389), .IN2(n10390), .QN(n10354) );
  NOR2X0 U10083 ( .IN1(n10391), .IN2(n10392), .QN(n10389) );
  NOR2X0 U10084 ( .IN1(n10393), .IN2(n10379), .QN(n10392) );
  NOR2X0 U10085 ( .IN1(n10380), .IN2(n10394), .QN(n10391) );
  NAND2X0 U10086 ( .IN1(n10395), .IN2(n10367), .QN(n10361) );
  NOR2X0 U10087 ( .IN1(n10396), .IN2(n10397), .QN(n10395) );
  NOR2X0 U10088 ( .IN1(n10398), .IN2(n10371), .QN(n10397) );
  NOR2X0 U10089 ( .IN1(n10372), .IN2(n10399), .QN(n10396) );
  XNOR2X1 U10090 ( .IN1(n10349), .IN2(n10342), .Q(n10387) );
  NAND2X0 U10091 ( .IN1(n10400), .IN2(n10390), .QN(n10342) );
  NOR2X0 U10092 ( .IN1(n10401), .IN2(n10402), .QN(n10400) );
  NOR2X0 U10093 ( .IN1(n10403), .IN2(n10371), .QN(n10402) );
  INVX0 U10094 ( .INP(n10404), .ZN(n10403) );
  NOR2X0 U10095 ( .IN1(n10372), .IN2(n10404), .QN(n10401) );
  NAND2X0 U10096 ( .IN1(n10405), .IN2(n10367), .QN(n10349) );
  INVX0 U10097 ( .INP(n10406), .ZN(n10367) );
  NAND2X0 U10098 ( .IN1(n10390), .IN2(n10407), .QN(n10406) );
  NAND2X0 U10099 ( .IN1(n10408), .IN2(n10409), .QN(n10407) );
  NOR2X0 U10100 ( .IN1(n10410), .IN2(n10411), .QN(n10405) );
  NOR2X0 U10101 ( .IN1(n10412), .IN2(n10371), .QN(n10411) );
  NOR2X0 U10102 ( .IN1(n10372), .IN2(n10413), .QN(n10410) );
  XOR2X1 U10103 ( .IN1(n10414), .IN2(n10415), .Q(n10385) );
  XNOR2X1 U10104 ( .IN1(n10313), .IN2(n10321), .Q(n10415) );
  INVX0 U10105 ( .INP(n10416), .ZN(n10321) );
  NAND2X0 U10106 ( .IN1(n10417), .IN2(n10390), .QN(n10416) );
  NOR2X0 U10107 ( .IN1(n10418), .IN2(n10419), .QN(n10417) );
  NOR2X0 U10108 ( .IN1(n10420), .IN2(n10379), .QN(n10419) );
  INVX0 U10109 ( .INP(n10421), .ZN(n10420) );
  NOR2X0 U10110 ( .IN1(n10380), .IN2(n10421), .QN(n10418) );
  NAND2X0 U10111 ( .IN1(n10422), .IN2(n10390), .QN(n10313) );
  NOR2X0 U10112 ( .IN1(n10423), .IN2(n10424), .QN(n10422) );
  NOR2X0 U10113 ( .IN1(n10425), .IN2(n10379), .QN(n10424) );
  NOR2X0 U10114 ( .IN1(n10380), .IN2(n10426), .QN(n10423) );
  XNOR2X1 U10115 ( .IN1(n10329), .IN2(n10336), .Q(n10414) );
  NAND2X0 U10116 ( .IN1(n10427), .IN2(n10390), .QN(n10336) );
  NOR2X0 U10117 ( .IN1(n10428), .IN2(n10429), .QN(n10427) );
  NOR2X0 U10118 ( .IN1(n10430), .IN2(n10371), .QN(n10429) );
  NAND2X0 U10119 ( .IN1(n10372), .IN2(n10431), .QN(n10371) );
  NOR2X0 U10120 ( .IN1(n10372), .IN2(n10432), .QN(n10428) );
  NAND2X0 U10121 ( .IN1(n10433), .IN2(n10375), .QN(n10329) );
  INVX0 U10122 ( .INP(n10434), .ZN(n10375) );
  NAND2X0 U10123 ( .IN1(n10390), .IN2(n10435), .QN(n10434) );
  NAND2X0 U10124 ( .IN1(n10408), .IN2(n10436), .QN(n10435) );
  NOR2X0 U10125 ( .IN1(n10362), .IN2(n4548), .QN(n10390) );
  NOR2X0 U10126 ( .IN1(n10437), .IN2(n10438), .QN(n10433) );
  NOR2X0 U10127 ( .IN1(n10439), .IN2(n10379), .QN(n10438) );
  NAND2X0 U10128 ( .IN1(n10380), .IN2(n10431), .QN(n10379) );
  NOR2X0 U10129 ( .IN1(n10380), .IN2(n10440), .QN(n10437) );
  NOR2X0 U10130 ( .IN1(n10441), .IN2(n10442), .QN(n10382) );
  NAND2X0 U10131 ( .IN1(n10308), .IN2(n10323), .QN(n10442) );
  NOR2X0 U10132 ( .IN1(n10362), .IN2(n10322), .QN(n10323) );
  NAND2X0 U10133 ( .IN1(n10443), .IN2(n9037), .QN(n10362) );
  NOR2X0 U10134 ( .IN1(g1249), .IN2(n521), .QN(n10443) );
  NAND2X0 U10135 ( .IN1(n10444), .IN2(n10445), .QN(n10441) );
  NAND2X0 U10136 ( .IN1(n4489), .IN2(g3229), .QN(n10445) );
  NAND2X0 U10137 ( .IN1(n10022), .IN2(n16819), .QN(n10444) );
  INVX0 U10138 ( .INP(n10446), .ZN(n3788) );
  INVX0 U10139 ( .INP(n10447), .ZN(n3758) );
  INVX0 U10140 ( .INP(n10448), .ZN(n3751) );
  NAND2X0 U10141 ( .IN1(n3896), .IN2(g88), .QN(n4528) );
  NAND2X0 U10142 ( .IN1(n3890), .IN2(g1462), .QN(n4527) );
  NAND2X0 U10143 ( .IN1(n3887), .IN2(test_so78), .QN(n4526) );
  INVX0 U10144 ( .INP(n10449), .ZN(n348) );
  NAND2X0 U10145 ( .IN1(n3692), .IN2(test_so15), .QN(n4521) );
  NAND2X0 U10146 ( .IN1(n3686), .IN2(g1453), .QN(n4523) );
  NAND2X0 U10147 ( .IN1(n3683), .IN2(g2147), .QN(n4522) );
  NAND2X0 U10148 ( .IN1(n10450), .IN2(n10451), .QN(n3254) );
  INVX0 U10149 ( .INP(n10452), .ZN(n10450) );
  NOR2X0 U10150 ( .IN1(n10453), .IN2(n10454), .QN(n10452) );
  INVX0 U10151 ( .INP(n10455), .ZN(n3128) );
  INVX0 U10152 ( .INP(g24734), .ZN(n307) );
  INVX0 U10153 ( .INP(n10456), .ZN(n3068) );
  NAND2X0 U10154 ( .IN1(n10457), .IN2(n10458), .QN(n3023) );
  NOR2X0 U10155 ( .IN1(n4388), .IN2(n10459), .QN(n10458) );
  NOR2X0 U10156 ( .IN1(n10460), .IN2(n10461), .QN(n10457) );
  NAND2X0 U10157 ( .IN1(n10462), .IN2(n10463), .QN(n3016) );
  NOR2X0 U10158 ( .IN1(n10464), .IN2(n10465), .QN(n10463) );
  NAND2X0 U10159 ( .IN1(n10466), .IN2(g996), .QN(n10465) );
  NOR2X0 U10160 ( .IN1(n10467), .IN2(n10468), .QN(n10462) );
  NAND2X0 U10161 ( .IN1(n10469), .IN2(n10470), .QN(n3008) );
  NOR2X0 U10162 ( .IN1(n4386), .IN2(n10471), .QN(n10470) );
  NOR2X0 U10163 ( .IN1(n10472), .IN2(n10473), .QN(n10469) );
  NAND2X0 U10164 ( .IN1(n10474), .IN2(n10475), .QN(n3000) );
  NOR2X0 U10165 ( .IN1(n10476), .IN2(n10477), .QN(n10475) );
  NAND2X0 U10166 ( .IN1(test_so79), .IN2(n10478), .QN(n10477) );
  NOR2X0 U10167 ( .IN1(n10479), .IN2(n10480), .QN(n10474) );
  INVX0 U10168 ( .INP(g25435), .ZN(n299) );
  INVX0 U10169 ( .INP(n10481), .ZN(n295) );
  XNOR2X1 U10170 ( .IN1(n10482), .IN2(n10483), .Q(n2800) );
  NAND2X0 U10171 ( .IN1(n10484), .IN2(n10485), .QN(n10482) );
  NAND2X0 U10172 ( .IN1(n10486), .IN2(n10487), .QN(n10485) );
  NAND2X0 U10173 ( .IN1(n10488), .IN2(n10489), .QN(n10487) );
  NOR2X0 U10174 ( .IN1(n10490), .IN2(n10491), .QN(n10488) );
  NOR2X0 U10175 ( .IN1(n10492), .IN2(n10493), .QN(n10491) );
  NAND2X0 U10176 ( .IN1(n10494), .IN2(g996), .QN(n10493) );
  NOR2X0 U10177 ( .IN1(n10495), .IN2(n10496), .QN(n10490) );
  NAND2X0 U10178 ( .IN1(n10497), .IN2(n10498), .QN(n10484) );
  INVX0 U10179 ( .INP(n10499), .ZN(n10497) );
  INVX0 U10180 ( .INP(g26135), .ZN(n276) );
  XNOR2X1 U10181 ( .IN1(n10500), .IN2(n10501), .Q(n2719) );
  XNOR2X1 U10182 ( .IN1(n10502), .IN2(n4530), .Q(n2686) );
  XNOR2X1 U10183 ( .IN1(n9851), .IN2(n10503), .Q(n2671) );
  XNOR2X1 U10184 ( .IN1(n10492), .IN2(n10504), .Q(n2616) );
  NOR2X0 U10185 ( .IN1(n10505), .IN2(n10506), .QN(n10504) );
  NOR2X0 U10186 ( .IN1(n10507), .IN2(n10508), .QN(n10506) );
  NOR2X0 U10187 ( .IN1(n10509), .IN2(n10510), .QN(n10508) );
  NOR2X0 U10188 ( .IN1(n10492), .IN2(n10511), .QN(n10510) );
  NOR2X0 U10189 ( .IN1(n10512), .IN2(n10513), .QN(n10511) );
  NOR2X0 U10190 ( .IN1(n10483), .IN2(n10514), .QN(n10513) );
  NAND2X0 U10191 ( .IN1(n10515), .IN2(n10496), .QN(n10514) );
  NOR2X0 U10192 ( .IN1(n10516), .IN2(n10517), .QN(n10496) );
  NOR2X0 U10193 ( .IN1(n10518), .IN2(n10519), .QN(n10517) );
  NOR2X0 U10194 ( .IN1(n10520), .IN2(n10521), .QN(n10515) );
  NOR2X0 U10195 ( .IN1(n10522), .IN2(n10519), .QN(n10521) );
  INVX0 U10196 ( .INP(n10523), .ZN(n10522) );
  NOR2X0 U10197 ( .IN1(n2632), .IN2(n10524), .QN(n10520) );
  NOR2X0 U10198 ( .IN1(n10486), .IN2(n10525), .QN(n10512) );
  NAND2X0 U10199 ( .IN1(n2632), .IN2(n10467), .QN(n10525) );
  NOR2X0 U10200 ( .IN1(n10495), .IN2(n10526), .QN(n10509) );
  NOR2X0 U10201 ( .IN1(n10527), .IN2(n10519), .QN(n10526) );
  NOR2X0 U10202 ( .IN1(n10528), .IN2(n10524), .QN(n10527) );
  NOR2X0 U10203 ( .IN1(n10523), .IN2(n10529), .QN(n10528) );
  NAND2X0 U10204 ( .IN1(n10486), .IN2(n10518), .QN(n10529) );
  NOR2X0 U10205 ( .IN1(n10530), .IN2(n10489), .QN(n10505) );
  NOR2X0 U10206 ( .IN1(n10483), .IN2(n10492), .QN(n10530) );
  NOR2X0 U10207 ( .IN1(n9909), .IN2(n9875), .QN(n2446) );
  INVX0 U10208 ( .INP(n9904), .ZN(n9875) );
  NAND2X0 U10209 ( .IN1(n4360), .IN2(n10531), .QN(n9904) );
  NAND2X0 U10210 ( .IN1(n8995), .IN2(n9285), .QN(n10531) );
  NAND2X0 U10211 ( .IN1(n9285), .IN2(n10532), .QN(n9909) );
  NAND2X0 U10212 ( .IN1(n4360), .IN2(n8995), .QN(n10532) );
  NAND2X0 U10213 ( .IN1(g499), .IN2(n10533), .QN(n2445) );
  NAND2X0 U10214 ( .IN1(n10534), .IN2(n10535), .QN(n10533) );
  NOR2X0 U10215 ( .IN1(n10000), .IN2(n10536), .QN(n10535) );
  NOR2X0 U10216 ( .IN1(n4295), .IN2(g734), .QN(n10536) );
  INVX0 U10217 ( .INP(n10005), .ZN(n10000) );
  NAND2X0 U10218 ( .IN1(n10537), .IN2(n10538), .QN(n10005) );
  NOR2X0 U10219 ( .IN1(n10539), .IN2(n10540), .QN(n10538) );
  NAND2X0 U10220 ( .IN1(n10541), .IN2(n9994), .QN(n10540) );
  NOR2X0 U10221 ( .IN1(n10004), .IN2(n9987), .QN(n10541) );
  INVX0 U10222 ( .INP(n10006), .ZN(n10004) );
  INVX0 U10223 ( .INP(n10542), .ZN(n10539) );
  NOR2X0 U10224 ( .IN1(n10543), .IN2(n10013), .QN(n10542) );
  INVX0 U10225 ( .INP(n10014), .ZN(n10013) );
  NAND2X0 U10226 ( .IN1(n10544), .IN2(n9953), .QN(n10543) );
  NOR2X0 U10227 ( .IN1(n10545), .IN2(n10546), .QN(n10537) );
  NAND2X0 U10228 ( .IN1(n10547), .IN2(n9965), .QN(n10546) );
  NOR2X0 U10229 ( .IN1(n9960), .IN2(n9971), .QN(n10547) );
  NAND2X0 U10230 ( .IN1(n10548), .IN2(n9977), .QN(n10545) );
  NOR2X0 U10231 ( .IN1(n10549), .IN2(n9983), .QN(n10548) );
  NOR2X0 U10232 ( .IN1(n10550), .IN2(n10551), .QN(n10549) );
  NAND2X0 U10233 ( .IN1(n10552), .IN2(n10553), .QN(n10551) );
  NAND2X0 U10234 ( .IN1(n9222), .IN2(g629), .QN(n10553) );
  NAND2X0 U10235 ( .IN1(n9155), .IN2(g6677), .QN(n10552) );
  NOR2X0 U10236 ( .IN1(n4359), .IN2(g739), .QN(n10550) );
  NOR2X0 U10237 ( .IN1(n10554), .IN2(n10555), .QN(n10534) );
  NOR2X0 U10238 ( .IN1(n4359), .IN2(g736), .QN(n10555) );
  NOR2X0 U10239 ( .IN1(n4309), .IN2(g735), .QN(n10554) );
  NAND2X0 U10240 ( .IN1(g2574), .IN2(n10556), .QN(n2374) );
  NAND2X0 U10241 ( .IN1(n10557), .IN2(n10558), .QN(n10556) );
  NOR2X0 U10242 ( .IN1(n10152), .IN2(n10559), .QN(n10558) );
  NOR2X0 U10243 ( .IN1(n4292), .IN2(g2808), .QN(n10559) );
  NOR2X0 U10244 ( .IN1(n10560), .IN2(n10561), .QN(n10557) );
  NOR2X0 U10245 ( .IN1(n4356), .IN2(g2810), .QN(n10561) );
  NOR2X0 U10246 ( .IN1(n4306), .IN2(g2809), .QN(n10560) );
  NOR2X0 U10247 ( .IN1(n10041), .IN2(n10027), .QN(n2361) );
  INVX0 U10248 ( .INP(n10036), .ZN(n10027) );
  NAND2X0 U10249 ( .IN1(n4352), .IN2(n10562), .QN(n10036) );
  NAND2X0 U10250 ( .IN1(n4303), .IN2(n8992), .QN(n10562) );
  NAND2X0 U10251 ( .IN1(n4303), .IN2(n10563), .QN(n10041) );
  NAND2X0 U10252 ( .IN1(n8992), .IN2(n4352), .QN(n10563) );
  NAND2X0 U10253 ( .IN1(g1880), .IN2(n10564), .QN(n2302) );
  NAND2X0 U10254 ( .IN1(n10565), .IN2(n10566), .QN(n10564) );
  NOR2X0 U10255 ( .IN1(n10265), .IN2(n10567), .QN(n10566) );
  NOR2X0 U10256 ( .IN1(n4293), .IN2(g2114), .QN(n10567) );
  INVX0 U10257 ( .INP(n10288), .ZN(n10265) );
  NAND2X0 U10258 ( .IN1(n10568), .IN2(n10569), .QN(n10288) );
  NOR2X0 U10259 ( .IN1(n10570), .IN2(n10571), .QN(n10569) );
  NAND2X0 U10260 ( .IN1(n10572), .IN2(n10297), .QN(n10571) );
  NOR2X0 U10261 ( .IN1(n10227), .IN2(n10269), .QN(n10572) );
  INVX0 U10262 ( .INP(n10230), .ZN(n10227) );
  INVX0 U10263 ( .INP(n10573), .ZN(n10570) );
  NOR2X0 U10264 ( .IN1(n10574), .IN2(n10255), .QN(n10573) );
  NAND2X0 U10265 ( .IN1(n10238), .IN2(n10575), .QN(n10574) );
  NOR2X0 U10266 ( .IN1(n10576), .IN2(n10577), .QN(n10568) );
  NAND2X0 U10267 ( .IN1(n10578), .IN2(n10282), .QN(n10577) );
  NOR2X0 U10268 ( .IN1(n10278), .IN2(n10289), .QN(n10578) );
  NAND2X0 U10269 ( .IN1(n10579), .IN2(n10250), .QN(n10576) );
  INVX0 U10270 ( .INP(n10251), .ZN(n10250) );
  NOR2X0 U10271 ( .IN1(n10580), .IN2(n10261), .QN(n10579) );
  NOR2X0 U10272 ( .IN1(n10581), .IN2(n10582), .QN(n10580) );
  NAND2X0 U10273 ( .IN1(n10583), .IN2(n10584), .QN(n10582) );
  NAND2X0 U10274 ( .IN1(n9220), .IN2(g2009), .QN(n10584) );
  NAND2X0 U10275 ( .IN1(n9153), .IN2(g7229), .QN(n10583) );
  NOR2X0 U10276 ( .IN1(n4357), .IN2(g2119), .QN(n10581) );
  NOR2X0 U10277 ( .IN1(n10585), .IN2(n10586), .QN(n10565) );
  NOR2X0 U10278 ( .IN1(n4357), .IN2(g2116), .QN(n10586) );
  NOR2X0 U10279 ( .IN1(n4307), .IN2(g2115), .QN(n10585) );
  NOR2X0 U10280 ( .IN1(n10181), .IN2(n10167), .QN(n2289) );
  INVX0 U10281 ( .INP(n10176), .ZN(n10167) );
  NAND2X0 U10282 ( .IN1(n4311), .IN2(n10587), .QN(n10176) );
  NAND2X0 U10283 ( .IN1(n4297), .IN2(n8993), .QN(n10587) );
  NAND2X0 U10284 ( .IN1(n4297), .IN2(n10588), .QN(n10181) );
  NAND2X0 U10285 ( .IN1(n8993), .IN2(n4311), .QN(n10588) );
  NAND2X0 U10286 ( .IN1(g1186), .IN2(n10589), .QN(n2230) );
  NAND2X0 U10287 ( .IN1(n10590), .IN2(n10591), .QN(n10589) );
  NOR2X0 U10288 ( .IN1(n10408), .IN2(n10592), .QN(n10591) );
  NOR2X0 U10289 ( .IN1(n4294), .IN2(g1420), .QN(n10592) );
  INVX0 U10290 ( .INP(n10431), .ZN(n10408) );
  NAND2X0 U10291 ( .IN1(n10593), .IN2(n10594), .QN(n10431) );
  NOR2X0 U10292 ( .IN1(n10595), .IN2(n10596), .QN(n10594) );
  NAND2X0 U10293 ( .IN1(n10597), .IN2(n10440), .QN(n10596) );
  NOR2X0 U10294 ( .IN1(n10370), .IN2(n10412), .QN(n10597) );
  INVX0 U10295 ( .INP(n10373), .ZN(n10370) );
  INVX0 U10296 ( .INP(n10598), .ZN(n10595) );
  NOR2X0 U10297 ( .IN1(n10599), .IN2(n10398), .QN(n10598) );
  NAND2X0 U10298 ( .IN1(n10381), .IN2(n10600), .QN(n10599) );
  NOR2X0 U10299 ( .IN1(n10601), .IN2(n10602), .QN(n10593) );
  NAND2X0 U10300 ( .IN1(n10603), .IN2(n10425), .QN(n10602) );
  NOR2X0 U10301 ( .IN1(n10421), .IN2(n10432), .QN(n10603) );
  NAND2X0 U10302 ( .IN1(n10604), .IN2(n10393), .QN(n10601) );
  NOR2X0 U10303 ( .IN1(n10605), .IN2(n10404), .QN(n10604) );
  NOR2X0 U10304 ( .IN1(n10606), .IN2(n10607), .QN(n10605) );
  NAND2X0 U10305 ( .IN1(n10608), .IN2(n10609), .QN(n10607) );
  NAND2X0 U10306 ( .IN1(n9221), .IN2(g1315), .QN(n10609) );
  NAND2X0 U10307 ( .IN1(n9154), .IN2(g6979), .QN(n10608) );
  NOR2X0 U10308 ( .IN1(n4358), .IN2(g1425), .QN(n10606) );
  NOR2X0 U10309 ( .IN1(n10610), .IN2(n10611), .QN(n10590) );
  NOR2X0 U10310 ( .IN1(n4358), .IN2(g1422), .QN(n10611) );
  NOR2X0 U10311 ( .IN1(n4308), .IN2(g1421), .QN(n10610) );
  NOR2X0 U10312 ( .IN1(n10322), .IN2(n10308), .QN(n2217) );
  INVX0 U10313 ( .INP(n10317), .ZN(n10308) );
  NAND2X0 U10314 ( .IN1(n4353), .IN2(n10612), .QN(n10317) );
  NAND2X0 U10315 ( .IN1(n4304), .IN2(n8994), .QN(n10612) );
  NAND2X0 U10316 ( .IN1(n4304), .IN2(n10613), .QN(n10322) );
  NAND2X0 U10317 ( .IN1(n8994), .IN2(n4353), .QN(n10613) );
  INVX0 U10318 ( .INP(n10614), .ZN(n1524) );
  NAND2X0 U10319 ( .IN1(n10615), .IN2(n10616), .QN(n10614) );
  NOR2X0 U10320 ( .IN1(n10617), .IN2(n10618), .QN(n10616) );
  NAND2X0 U10321 ( .IN1(n10619), .IN2(n4393), .QN(n10615) );
  INVX0 U10322 ( .INP(n10620), .ZN(n15) );
  INVX0 U10323 ( .INP(n10621), .ZN(n1499) );
  NAND2X0 U10324 ( .IN1(n10622), .IN2(n10623), .QN(n10621) );
  NAND2X0 U10325 ( .IN1(n10624), .IN2(n9152), .QN(n10623) );
  INVX0 U10326 ( .INP(n10625), .ZN(n1464) );
  NOR2X0 U10327 ( .IN1(n10626), .IN2(n10627), .QN(n10625) );
  NOR2X0 U10328 ( .IN1(g2624), .IN2(n9223), .QN(n10627) );
  NAND2X0 U10329 ( .IN1(n10152), .IN2(n10628), .QN(n1458) );
  INVX0 U10330 ( .INP(n10147), .ZN(n10152) );
  NAND2X0 U10331 ( .IN1(n10629), .IN2(n10630), .QN(n10147) );
  NOR2X0 U10332 ( .IN1(n10631), .IN2(n10632), .QN(n10630) );
  NAND2X0 U10333 ( .IN1(n10633), .IN2(n10157), .QN(n10632) );
  NOR2X0 U10334 ( .IN1(n10089), .IN2(n10128), .QN(n10633) );
  INVX0 U10335 ( .INP(n10634), .ZN(n10631) );
  NOR2X0 U10336 ( .IN1(n10635), .IN2(n10117), .QN(n10634) );
  NAND2X0 U10337 ( .IN1(n10099), .IN2(n10636), .QN(n10635) );
  NOR2X0 U10338 ( .IN1(n10637), .IN2(n10638), .QN(n10629) );
  NAND2X0 U10339 ( .IN1(n10639), .IN2(n10146), .QN(n10638) );
  NOR2X0 U10340 ( .IN1(n10113), .IN2(n10137), .QN(n10639) );
  NAND2X0 U10341 ( .IN1(n10640), .IN2(n10122), .QN(n10637) );
  NOR2X0 U10342 ( .IN1(n10641), .IN2(n10142), .QN(n10640) );
  NOR2X0 U10343 ( .IN1(n10642), .IN2(n10643), .QN(n10641) );
  NAND2X0 U10344 ( .IN1(n10644), .IN2(n10645), .QN(n10643) );
  INVX0 U10345 ( .INP(n10646), .ZN(n10645) );
  NOR2X0 U10346 ( .IN1(n4292), .IN2(test_so95), .QN(n10646) );
  NAND2X0 U10347 ( .IN1(n9152), .IN2(g7425), .QN(n10644) );
  NOR2X0 U10348 ( .IN1(n4356), .IN2(g2813), .QN(n10642) );
  INVX0 U10349 ( .INP(n10647), .ZN(n1456) );
  INVX0 U10350 ( .INP(n10648), .ZN(n1290) );
  INVX0 U10351 ( .INP(n10649), .ZN(n1194) );
  NAND2X0 U10352 ( .IN1(n10650), .IN2(n10651), .QN(n10649) );
  NAND2X0 U10353 ( .IN1(n10652), .IN2(n9153), .QN(n10651) );
  INVX0 U10354 ( .INP(n10653), .ZN(n1159) );
  NOR2X0 U10355 ( .IN1(n10654), .IN2(n10655), .QN(n10653) );
  NOR2X0 U10356 ( .IN1(g1930), .IN2(n9224), .QN(n10655) );
  NAND2X0 U10357 ( .IN1(n10656), .IN2(n10657), .QN(g30801) );
  INVX0 U10358 ( .INP(n10658), .ZN(n10657) );
  NOR2X0 U10359 ( .IN1(g3109), .IN2(n4334), .QN(n10658) );
  NAND2X0 U10360 ( .IN1(g30072), .IN2(g3109), .QN(n10656) );
  NAND2X0 U10361 ( .IN1(n10659), .IN2(n10660), .QN(g30798) );
  INVX0 U10362 ( .INP(n10661), .ZN(n10660) );
  NOR2X0 U10363 ( .IN1(g8030), .IN2(n4437), .QN(n10661) );
  NAND2X0 U10364 ( .IN1(g30072), .IN2(g8030), .QN(n10659) );
  NAND2X0 U10365 ( .IN1(n10662), .IN2(n10663), .QN(g30796) );
  INVX0 U10366 ( .INP(n10664), .ZN(n10663) );
  NOR2X0 U10367 ( .IN1(g8106), .IN2(n4438), .QN(n10664) );
  NAND2X0 U10368 ( .IN1(g30072), .IN2(g8106), .QN(n10662) );
  NAND2X0 U10369 ( .IN1(n10665), .IN2(n10666), .QN(g30709) );
  NAND2X0 U10370 ( .IN1(n10667), .IN2(g7264), .QN(n10666) );
  INVX0 U10371 ( .INP(n10668), .ZN(n10665) );
  NOR2X0 U10372 ( .IN1(n10669), .IN2(n8494), .QN(n10668) );
  NAND2X0 U10373 ( .IN1(n10670), .IN2(n10671), .QN(g30708) );
  NAND2X0 U10374 ( .IN1(n10672), .IN2(n4618), .QN(n10671) );
  NAND2X0 U10375 ( .IN1(n4511), .IN2(g1698), .QN(n10670) );
  NAND2X0 U10376 ( .IN1(n10673), .IN2(n10674), .QN(g30707) );
  NAND2X0 U10377 ( .IN1(n10667), .IN2(g5555), .QN(n10674) );
  NAND2X0 U10378 ( .IN1(n4516), .IN2(g2390), .QN(n10673) );
  NAND2X0 U10379 ( .IN1(n10675), .IN2(n10676), .QN(g30706) );
  NAND2X0 U10380 ( .IN1(n10672), .IN2(g7014), .QN(n10676) );
  INVX0 U10381 ( .INP(n10677), .ZN(n10675) );
  NOR2X0 U10382 ( .IN1(n10678), .IN2(n8497), .QN(n10677) );
  NAND2X0 U10383 ( .IN1(n10679), .IN2(n10680), .QN(g30705) );
  INVX0 U10384 ( .INP(n10681), .ZN(n10680) );
  NOR2X0 U10385 ( .IN1(g1088), .IN2(n8515), .QN(n10681) );
  NAND2X0 U10386 ( .IN1(n2594), .IN2(g1088), .QN(n10679) );
  NAND2X0 U10387 ( .IN1(n10682), .IN2(n10683), .QN(g30704) );
  NAND2X0 U10388 ( .IN1(n10672), .IN2(g5511), .QN(n10683) );
  NOR2X0 U10389 ( .IN1(n10684), .IN2(n10685), .QN(n10672) );
  XNOR2X1 U10390 ( .IN1(n10686), .IN2(n10687), .Q(n10684) );
  NOR2X0 U10391 ( .IN1(n10688), .IN2(n10689), .QN(n10687) );
  NOR2X0 U10392 ( .IN1(n10690), .IN2(n10691), .QN(n10689) );
  NAND2X0 U10393 ( .IN1(n10692), .IN2(n10693), .QN(n10691) );
  NAND2X0 U10394 ( .IN1(n10694), .IN2(n10686), .QN(n10693) );
  NOR2X0 U10395 ( .IN1(n10695), .IN2(n10696), .QN(n10692) );
  NOR2X0 U10396 ( .IN1(n10697), .IN2(n10698), .QN(n10696) );
  NOR2X0 U10397 ( .IN1(n10699), .IN2(n10700), .QN(n10697) );
  NOR2X0 U10398 ( .IN1(n10701), .IN2(n10702), .QN(n10695) );
  NOR2X0 U10399 ( .IN1(n10703), .IN2(n10704), .QN(n10701) );
  NOR2X0 U10400 ( .IN1(n10686), .IN2(n10699), .QN(n10704) );
  NOR2X0 U10401 ( .IN1(n10705), .IN2(n10700), .QN(n10703) );
  XNOR2X1 U10402 ( .IN1(n10706), .IN2(n10707), .Q(n10705) );
  NAND2X0 U10403 ( .IN1(n10708), .IN2(n10709), .QN(n10706) );
  NOR2X0 U10404 ( .IN1(n10710), .IN2(n10711), .QN(n10688) );
  NAND2X0 U10405 ( .IN1(n4518), .IN2(g1696), .QN(n10682) );
  NAND2X0 U10406 ( .IN1(n10712), .IN2(n10713), .QN(g30703) );
  NAND2X0 U10407 ( .IN1(n4364), .IN2(g1003), .QN(n10713) );
  NAND2X0 U10408 ( .IN1(n2594), .IN2(g6712), .QN(n10712) );
  NAND2X0 U10409 ( .IN1(n10714), .IN2(n10715), .QN(g30702) );
  NAND2X0 U10410 ( .IN1(n10716), .IN2(n4640), .QN(n10715) );
  NAND2X0 U10411 ( .IN1(n4506), .IN2(g317), .QN(n10714) );
  NAND2X0 U10412 ( .IN1(n10717), .IN2(n10718), .QN(g30701) );
  NAND2X0 U10413 ( .IN1(n4363), .IN2(g1002), .QN(n10718) );
  NAND2X0 U10414 ( .IN1(n2594), .IN2(g5472), .QN(n10717) );
  NAND2X0 U10415 ( .IN1(n10719), .IN2(n10720), .QN(g30700) );
  NAND2X0 U10416 ( .IN1(n10716), .IN2(g6447), .QN(n10720) );
  NAND2X0 U10417 ( .IN1(test_so18), .IN2(n4499), .QN(n10719) );
  NAND2X0 U10418 ( .IN1(n10721), .IN2(n10722), .QN(g30699) );
  NAND2X0 U10419 ( .IN1(n10716), .IN2(g5437), .QN(n10722) );
  NOR2X0 U10420 ( .IN1(n10723), .IN2(n10724), .QN(n10716) );
  XNOR2X1 U10421 ( .IN1(n10725), .IN2(n10726), .Q(n10723) );
  NOR2X0 U10422 ( .IN1(n10727), .IN2(n10728), .QN(n10726) );
  NOR2X0 U10423 ( .IN1(n10729), .IN2(n10730), .QN(n10728) );
  NAND2X0 U10424 ( .IN1(n10731), .IN2(n10732), .QN(n10730) );
  NAND2X0 U10425 ( .IN1(n10733), .IN2(n10725), .QN(n10732) );
  NOR2X0 U10426 ( .IN1(n10734), .IN2(n10735), .QN(n10731) );
  NOR2X0 U10427 ( .IN1(n10736), .IN2(n10737), .QN(n10735) );
  NOR2X0 U10428 ( .IN1(n10738), .IN2(n10739), .QN(n10736) );
  NOR2X0 U10429 ( .IN1(n10740), .IN2(n10741), .QN(n10734) );
  NOR2X0 U10430 ( .IN1(n10742), .IN2(n10743), .QN(n10740) );
  NOR2X0 U10431 ( .IN1(n10725), .IN2(n10738), .QN(n10743) );
  NOR2X0 U10432 ( .IN1(n10744), .IN2(n10739), .QN(n10742) );
  XNOR2X1 U10433 ( .IN1(n10745), .IN2(n10746), .Q(n10744) );
  NAND2X0 U10434 ( .IN1(n10747), .IN2(n10748), .QN(n10745) );
  NOR2X0 U10435 ( .IN1(n10749), .IN2(n10750), .QN(n10727) );
  INVX0 U10436 ( .INP(n10751), .ZN(n10721) );
  NOR2X0 U10437 ( .IN1(n10752), .IN2(n8523), .QN(n10751) );
  NAND2X0 U10438 ( .IN1(n10753), .IN2(n10754), .QN(g30695) );
  INVX0 U10439 ( .INP(n10755), .ZN(n10754) );
  NOR2X0 U10440 ( .IN1(g2241), .IN2(n8536), .QN(n10755) );
  NAND2X0 U10441 ( .IN1(n10756), .IN2(g2241), .QN(n10753) );
  NAND2X0 U10442 ( .IN1(n10757), .IN2(n10758), .QN(g30694) );
  INVX0 U10443 ( .INP(n10759), .ZN(n10758) );
  NOR2X0 U10444 ( .IN1(g2241), .IN2(n8376), .QN(n10759) );
  NAND2X0 U10445 ( .IN1(n10760), .IN2(g2241), .QN(n10757) );
  NAND2X0 U10446 ( .IN1(n10761), .IN2(n10762), .QN(g30693) );
  NAND2X0 U10447 ( .IN1(g2273), .IN2(n9278), .QN(n10762) );
  NAND2X0 U10448 ( .IN1(test_so73), .IN2(n10756), .QN(n10761) );
  NAND2X0 U10449 ( .IN1(n10763), .IN2(n10764), .QN(g30692) );
  INVX0 U10450 ( .INP(n10765), .ZN(n10764) );
  NOR2X0 U10451 ( .IN1(g1547), .IN2(n8539), .QN(n10765) );
  NAND2X0 U10452 ( .IN1(n10766), .IN2(g1547), .QN(n10763) );
  NAND2X0 U10453 ( .IN1(n10767), .IN2(n10768), .QN(g30691) );
  NAND2X0 U10454 ( .IN1(g2345), .IN2(n9278), .QN(n10768) );
  NAND2X0 U10455 ( .IN1(n10760), .IN2(test_so73), .QN(n10767) );
  NAND2X0 U10456 ( .IN1(n10769), .IN2(n10770), .QN(g30690) );
  INVX0 U10457 ( .INP(n10771), .ZN(n10770) );
  NOR2X0 U10458 ( .IN1(g6837), .IN2(n8439), .QN(n10771) );
  NAND2X0 U10459 ( .IN1(n10756), .IN2(g6837), .QN(n10769) );
  NAND2X0 U10460 ( .IN1(n10772), .IN2(n10773), .QN(n10756) );
  NOR2X0 U10461 ( .IN1(n10774), .IN2(n10775), .QN(n10772) );
  NOR2X0 U10462 ( .IN1(n4319), .IN2(n10776), .QN(n10775) );
  NOR2X0 U10463 ( .IN1(n10777), .IN2(n10778), .QN(n10774) );
  XNOR2X1 U10464 ( .IN1(n9850), .IN2(n10779), .Q(n10778) );
  NAND2X0 U10465 ( .IN1(n10780), .IN2(n10781), .QN(g30689) );
  INVX0 U10466 ( .INP(n10782), .ZN(n10781) );
  NOR2X0 U10467 ( .IN1(g1547), .IN2(n8413), .QN(n10782) );
  NAND2X0 U10468 ( .IN1(n10783), .IN2(g1547), .QN(n10780) );
  NAND2X0 U10469 ( .IN1(n10784), .IN2(n10785), .QN(g30688) );
  NAND2X0 U10470 ( .IN1(n4515), .IN2(g1579), .QN(n10785) );
  NAND2X0 U10471 ( .IN1(n10766), .IN2(g6782), .QN(n10784) );
  NAND2X0 U10472 ( .IN1(n10786), .IN2(n10787), .QN(g30687) );
  NAND2X0 U10473 ( .IN1(g888), .IN2(n9279), .QN(n10787) );
  NAND2X0 U10474 ( .IN1(test_so31), .IN2(n10788), .QN(n10786) );
  NAND2X0 U10475 ( .IN1(n10789), .IN2(n10790), .QN(g30686) );
  INVX0 U10476 ( .INP(n10791), .ZN(n10790) );
  NOR2X0 U10477 ( .IN1(g6837), .IN2(n8377), .QN(n10791) );
  NAND2X0 U10478 ( .IN1(n10760), .IN2(g6837), .QN(n10789) );
  INVX0 U10479 ( .INP(n10792), .ZN(n10760) );
  NAND2X0 U10480 ( .IN1(n10793), .IN2(n10794), .QN(n10792) );
  NAND2X0 U10481 ( .IN1(n10795), .IN2(n10796), .QN(n10794) );
  NOR2X0 U10482 ( .IN1(n10797), .IN2(n10798), .QN(n10793) );
  NOR2X0 U10483 ( .IN1(n10777), .IN2(n10799), .QN(n10798) );
  XNOR2X1 U10484 ( .IN1(n2669), .IN2(n10800), .Q(n10799) );
  NAND2X0 U10485 ( .IN1(n10801), .IN2(n10802), .QN(g30684) );
  NAND2X0 U10486 ( .IN1(n4515), .IN2(g1651), .QN(n10802) );
  NAND2X0 U10487 ( .IN1(n10783), .IN2(g6782), .QN(n10801) );
  NAND2X0 U10488 ( .IN1(n10803), .IN2(n10804), .QN(g30683) );
  INVX0 U10489 ( .INP(n10805), .ZN(n10804) );
  NOR2X0 U10490 ( .IN1(g6573), .IN2(n8451), .QN(n10805) );
  NAND2X0 U10491 ( .IN1(n10766), .IN2(g6573), .QN(n10803) );
  NAND2X0 U10492 ( .IN1(n10806), .IN2(n10807), .QN(n10766) );
  NOR2X0 U10493 ( .IN1(n10808), .IN2(n10809), .QN(n10806) );
  NOR2X0 U10494 ( .IN1(n4320), .IN2(n10810), .QN(n10809) );
  NOR2X0 U10495 ( .IN1(n10811), .IN2(n10812), .QN(n10808) );
  XNOR2X1 U10496 ( .IN1(n9815), .IN2(n10813), .Q(n10812) );
  NAND2X0 U10497 ( .IN1(n10814), .IN2(n10815), .QN(g30682) );
  NAND2X0 U10498 ( .IN1(g960), .IN2(n9279), .QN(n10815) );
  NAND2X0 U10499 ( .IN1(n10816), .IN2(test_so31), .QN(n10814) );
  NAND2X0 U10500 ( .IN1(n10817), .IN2(n10818), .QN(g30681) );
  INVX0 U10501 ( .INP(n10819), .ZN(n10818) );
  NOR2X0 U10502 ( .IN1(g6518), .IN2(n8465), .QN(n10819) );
  NAND2X0 U10503 ( .IN1(n10788), .IN2(g6518), .QN(n10817) );
  NAND2X0 U10504 ( .IN1(n10820), .IN2(n10821), .QN(g30680) );
  INVX0 U10505 ( .INP(n10822), .ZN(n10821) );
  NOR2X0 U10506 ( .IN1(g165), .IN2(n8545), .QN(n10822) );
  NAND2X0 U10507 ( .IN1(n10823), .IN2(g165), .QN(n10820) );
  NAND2X0 U10508 ( .IN1(n10824), .IN2(n10825), .QN(g30679) );
  INVX0 U10509 ( .INP(n10826), .ZN(n10825) );
  NOR2X0 U10510 ( .IN1(g2241), .IN2(n8419), .QN(n10826) );
  NAND2X0 U10511 ( .IN1(n10827), .IN2(g2241), .QN(n10824) );
  NAND2X0 U10512 ( .IN1(n10828), .IN2(n10829), .QN(g30678) );
  INVX0 U10513 ( .INP(n10830), .ZN(n10829) );
  NOR2X0 U10514 ( .IN1(g6573), .IN2(n8412), .QN(n10830) );
  NAND2X0 U10515 ( .IN1(n10783), .IN2(g6573), .QN(n10828) );
  INVX0 U10516 ( .INP(n10831), .ZN(n10783) );
  NAND2X0 U10517 ( .IN1(n10832), .IN2(n10833), .QN(n10831) );
  NAND2X0 U10518 ( .IN1(n10834), .IN2(n10835), .QN(n10833) );
  NOR2X0 U10519 ( .IN1(n10836), .IN2(n10837), .QN(n10832) );
  NOR2X0 U10520 ( .IN1(n10811), .IN2(n10838), .QN(n10837) );
  XNOR2X1 U10521 ( .IN1(n2684), .IN2(n9830), .Q(n10838) );
  NAND2X0 U10522 ( .IN1(n10839), .IN2(n10840), .QN(g30677) );
  INVX0 U10523 ( .INP(n10841), .ZN(n10840) );
  NOR2X0 U10524 ( .IN1(g6518), .IN2(n8491), .QN(n10841) );
  NAND2X0 U10525 ( .IN1(n10816), .IN2(g6518), .QN(n10839) );
  NAND2X0 U10526 ( .IN1(n10842), .IN2(n10843), .QN(g30676) );
  INVX0 U10527 ( .INP(n10844), .ZN(n10843) );
  NOR2X0 U10528 ( .IN1(g6368), .IN2(n8466), .QN(n10844) );
  NAND2X0 U10529 ( .IN1(n10788), .IN2(g6368), .QN(n10842) );
  NAND2X0 U10530 ( .IN1(n10845), .IN2(n10846), .QN(n10788) );
  NOR2X0 U10531 ( .IN1(n10847), .IN2(n10848), .QN(n10845) );
  NOR2X0 U10532 ( .IN1(n4321), .IN2(n10849), .QN(n10848) );
  NOR2X0 U10533 ( .IN1(n10850), .IN2(n10851), .QN(n10847) );
  XNOR2X1 U10534 ( .IN1(n9794), .IN2(n10852), .Q(n10851) );
  NAND2X0 U10535 ( .IN1(n10853), .IN2(n10854), .QN(g30675) );
  INVX0 U10536 ( .INP(n10855), .ZN(n10854) );
  NOR2X0 U10537 ( .IN1(g165), .IN2(n8416), .QN(n10855) );
  NAND2X0 U10538 ( .IN1(n10856), .IN2(g165), .QN(n10853) );
  NAND2X0 U10539 ( .IN1(n10857), .IN2(n10858), .QN(g30674) );
  NAND2X0 U10540 ( .IN1(n4512), .IN2(g198), .QN(n10858) );
  NAND2X0 U10541 ( .IN1(n10823), .IN2(g6313), .QN(n10857) );
  NAND2X0 U10542 ( .IN1(n10859), .IN2(n10860), .QN(g30673) );
  NAND2X0 U10543 ( .IN1(g2318), .IN2(n9278), .QN(n10860) );
  NAND2X0 U10544 ( .IN1(n10827), .IN2(test_so73), .QN(n10859) );
  NAND2X0 U10545 ( .IN1(n10861), .IN2(n10862), .QN(g30672) );
  INVX0 U10546 ( .INP(n10863), .ZN(n10862) );
  NOR2X0 U10547 ( .IN1(g2241), .IN2(n8420), .QN(n10863) );
  NAND2X0 U10548 ( .IN1(n10864), .IN2(g2241), .QN(n10861) );
  NAND2X0 U10549 ( .IN1(n10865), .IN2(n10866), .QN(g30671) );
  INVX0 U10550 ( .INP(n10867), .ZN(n10866) );
  NOR2X0 U10551 ( .IN1(g1547), .IN2(n8422), .QN(n10867) );
  NAND2X0 U10552 ( .IN1(n10868), .IN2(g1547), .QN(n10865) );
  NAND2X0 U10553 ( .IN1(n10869), .IN2(n10870), .QN(g30670) );
  INVX0 U10554 ( .INP(n10871), .ZN(n10870) );
  NOR2X0 U10555 ( .IN1(g6368), .IN2(n8455), .QN(n10871) );
  NAND2X0 U10556 ( .IN1(n10816), .IN2(g6368), .QN(n10869) );
  INVX0 U10557 ( .INP(n10872), .ZN(n10816) );
  NAND2X0 U10558 ( .IN1(n10873), .IN2(n10874), .QN(n10872) );
  NAND2X0 U10559 ( .IN1(n10875), .IN2(n10876), .QN(n10874) );
  NOR2X0 U10560 ( .IN1(n10877), .IN2(n10878), .QN(n10873) );
  NOR2X0 U10561 ( .IN1(n10879), .IN2(n10850), .QN(n10878) );
  XNOR2X1 U10562 ( .IN1(n10880), .IN2(n9793), .Q(n10879) );
  NAND2X0 U10563 ( .IN1(n10881), .IN2(n10882), .QN(n10880) );
  XNOR2X1 U10564 ( .IN1(n9795), .IN2(n10883), .Q(n10882) );
  NAND2X0 U10565 ( .IN1(n10884), .IN2(n10885), .QN(g30669) );
  NAND2X0 U10566 ( .IN1(n4512), .IN2(g270), .QN(n10885) );
  NAND2X0 U10567 ( .IN1(n10856), .IN2(g6313), .QN(n10884) );
  NAND2X0 U10568 ( .IN1(n10886), .IN2(n10887), .QN(g30668) );
  INVX0 U10569 ( .INP(n10888), .ZN(n10887) );
  NOR2X0 U10570 ( .IN1(g6231), .IN2(n8480), .QN(n10888) );
  NAND2X0 U10571 ( .IN1(n10823), .IN2(g6231), .QN(n10886) );
  NAND2X0 U10572 ( .IN1(n10889), .IN2(n10890), .QN(n10823) );
  NOR2X0 U10573 ( .IN1(n10891), .IN2(n10892), .QN(n10889) );
  NOR2X0 U10574 ( .IN1(n4322), .IN2(n10893), .QN(n10892) );
  NOR2X0 U10575 ( .IN1(n10894), .IN2(n10895), .QN(n10891) );
  XNOR2X1 U10576 ( .IN1(n9745), .IN2(n10896), .Q(n10895) );
  NAND2X0 U10577 ( .IN1(n10897), .IN2(n10898), .QN(g30667) );
  INVX0 U10578 ( .INP(n10899), .ZN(n10898) );
  NOR2X0 U10579 ( .IN1(g6837), .IN2(n8437), .QN(n10899) );
  NAND2X0 U10580 ( .IN1(n10827), .IN2(g6837), .QN(n10897) );
  INVX0 U10581 ( .INP(n10900), .ZN(n10827) );
  NAND2X0 U10582 ( .IN1(n10901), .IN2(n10902), .QN(n10900) );
  NAND2X0 U10583 ( .IN1(n10795), .IN2(n4389), .QN(n10902) );
  NOR2X0 U10584 ( .IN1(n10797), .IN2(n10903), .QN(n10901) );
  NOR2X0 U10585 ( .IN1(n10904), .IN2(n10777), .QN(n10903) );
  XOR2X1 U10586 ( .IN1(n9864), .IN2(n10905), .Q(n10904) );
  NAND2X0 U10587 ( .IN1(n10906), .IN2(n10907), .QN(g30666) );
  NAND2X0 U10588 ( .IN1(g2309), .IN2(n9278), .QN(n10907) );
  NAND2X0 U10589 ( .IN1(n10864), .IN2(test_so73), .QN(n10906) );
  NAND2X0 U10590 ( .IN1(n10908), .IN2(n10909), .QN(g30665) );
  INVX0 U10591 ( .INP(n10910), .ZN(n10909) );
  NOR2X0 U10592 ( .IN1(g2241), .IN2(n8384), .QN(n10910) );
  NAND2X0 U10593 ( .IN1(n10911), .IN2(g2241), .QN(n10908) );
  NAND2X0 U10594 ( .IN1(n10912), .IN2(n10913), .QN(g30664) );
  NAND2X0 U10595 ( .IN1(n4515), .IN2(g1624), .QN(n10913) );
  NAND2X0 U10596 ( .IN1(n10868), .IN2(g6782), .QN(n10912) );
  NAND2X0 U10597 ( .IN1(n10914), .IN2(n10915), .QN(g30663) );
  INVX0 U10598 ( .INP(n10916), .ZN(n10915) );
  NOR2X0 U10599 ( .IN1(g1547), .IN2(n8423), .QN(n10916) );
  NAND2X0 U10600 ( .IN1(n10917), .IN2(g1547), .QN(n10914) );
  NAND2X0 U10601 ( .IN1(n10918), .IN2(n10919), .QN(g30662) );
  NAND2X0 U10602 ( .IN1(g933), .IN2(n9279), .QN(n10919) );
  NAND2X0 U10603 ( .IN1(n10920), .IN2(test_so31), .QN(n10918) );
  NAND2X0 U10604 ( .IN1(n10921), .IN2(n10922), .QN(g30661) );
  INVX0 U10605 ( .INP(n10923), .ZN(n10922) );
  NOR2X0 U10606 ( .IN1(g6231), .IN2(n8415), .QN(n10923) );
  NAND2X0 U10607 ( .IN1(n10856), .IN2(g6231), .QN(n10921) );
  INVX0 U10608 ( .INP(n10924), .ZN(n10856) );
  NAND2X0 U10609 ( .IN1(n10925), .IN2(n10926), .QN(n10924) );
  NAND2X0 U10610 ( .IN1(n10927), .IN2(n10928), .QN(n10926) );
  NOR2X0 U10611 ( .IN1(n10929), .IN2(n10930), .QN(n10925) );
  NOR2X0 U10612 ( .IN1(n10894), .IN2(n10931), .QN(n10930) );
  XNOR2X1 U10613 ( .IN1(n2717), .IN2(n10932), .Q(n10931) );
  NAND2X0 U10614 ( .IN1(n10933), .IN2(n10934), .QN(g30660) );
  INVX0 U10615 ( .INP(n10935), .ZN(n10934) );
  NOR2X0 U10616 ( .IN1(g6837), .IN2(n8440), .QN(n10935) );
  NAND2X0 U10617 ( .IN1(n10864), .IN2(g6837), .QN(n10933) );
  INVX0 U10618 ( .INP(n10936), .ZN(n10864) );
  NAND2X0 U10619 ( .IN1(n10937), .IN2(n10938), .QN(n10936) );
  NAND2X0 U10620 ( .IN1(n10795), .IN2(n4373), .QN(n10938) );
  NOR2X0 U10621 ( .IN1(n10797), .IN2(n10939), .QN(n10937) );
  NOR2X0 U10622 ( .IN1(n10940), .IN2(n10777), .QN(n10939) );
  XNOR2X1 U10623 ( .IN1(n9858), .IN2(n10941), .Q(n10940) );
  NOR2X0 U10624 ( .IN1(n10942), .IN2(n10503), .QN(n10797) );
  INVX0 U10625 ( .INP(n10943), .ZN(n10942) );
  NAND2X0 U10626 ( .IN1(n10944), .IN2(n10945), .QN(g30659) );
  NAND2X0 U10627 ( .IN1(g2300), .IN2(n9278), .QN(n10945) );
  NAND2X0 U10628 ( .IN1(test_so73), .IN2(n10911), .QN(n10944) );
  NAND2X0 U10629 ( .IN1(n10946), .IN2(n10947), .QN(g30658) );
  NAND2X0 U10630 ( .IN1(n10868), .IN2(g6573), .QN(n10947) );
  INVX0 U10631 ( .INP(n10948), .ZN(n10868) );
  NAND2X0 U10632 ( .IN1(n10949), .IN2(n10950), .QN(n10948) );
  NAND2X0 U10633 ( .IN1(n10834), .IN2(n4390), .QN(n10950) );
  NOR2X0 U10634 ( .IN1(n10836), .IN2(n10951), .QN(n10949) );
  NOR2X0 U10635 ( .IN1(n10952), .IN2(n10811), .QN(n10951) );
  XNOR2X1 U10636 ( .IN1(n10953), .IN2(n10954), .Q(n10952) );
  NAND2X0 U10637 ( .IN1(test_so55), .IN2(n4317), .QN(n10946) );
  NAND2X0 U10638 ( .IN1(n10955), .IN2(n10956), .QN(g30657) );
  NAND2X0 U10639 ( .IN1(n4515), .IN2(g1615), .QN(n10956) );
  NAND2X0 U10640 ( .IN1(n10917), .IN2(g6782), .QN(n10955) );
  NAND2X0 U10641 ( .IN1(n10957), .IN2(n10958), .QN(g30656) );
  INVX0 U10642 ( .INP(n10959), .ZN(n10958) );
  NOR2X0 U10643 ( .IN1(g1547), .IN2(n8385), .QN(n10959) );
  NAND2X0 U10644 ( .IN1(n10960), .IN2(g1547), .QN(n10957) );
  NAND2X0 U10645 ( .IN1(n10961), .IN2(n10962), .QN(g30655) );
  INVX0 U10646 ( .INP(n10963), .ZN(n10962) );
  NOR2X0 U10647 ( .IN1(g6518), .IN2(n8487), .QN(n10963) );
  NAND2X0 U10648 ( .IN1(n10920), .IN2(g6518), .QN(n10961) );
  NAND2X0 U10649 ( .IN1(n10964), .IN2(n10965), .QN(g30654) );
  NAND2X0 U10650 ( .IN1(test_so34), .IN2(n9279), .QN(n10965) );
  NAND2X0 U10651 ( .IN1(n10966), .IN2(test_so31), .QN(n10964) );
  NAND2X0 U10652 ( .IN1(n10967), .IN2(n10968), .QN(g30653) );
  INVX0 U10653 ( .INP(n10969), .ZN(n10968) );
  NOR2X0 U10654 ( .IN1(g165), .IN2(n8428), .QN(n10969) );
  NAND2X0 U10655 ( .IN1(n10970), .IN2(g165), .QN(n10967) );
  NAND2X0 U10656 ( .IN1(n10971), .IN2(n10972), .QN(g30652) );
  INVX0 U10657 ( .INP(n10973), .ZN(n10972) );
  NOR2X0 U10658 ( .IN1(g6837), .IN2(n8378), .QN(n10973) );
  NAND2X0 U10659 ( .IN1(n10911), .IN2(g6837), .QN(n10971) );
  NAND2X0 U10660 ( .IN1(n10974), .IN2(n10773), .QN(n10911) );
  NAND2X0 U10661 ( .IN1(n10943), .IN2(n10975), .QN(n10773) );
  NOR2X0 U10662 ( .IN1(n10976), .IN2(n10977), .QN(n10974) );
  NOR2X0 U10663 ( .IN1(n10978), .IN2(n10776), .QN(n10977) );
  INVX0 U10664 ( .INP(n10795), .ZN(n10776) );
  NOR2X0 U10665 ( .IN1(n10777), .IN2(n10979), .QN(n10976) );
  XNOR2X1 U10666 ( .IN1(n9851), .IN2(n2670), .Q(n10979) );
  NAND2X0 U10667 ( .IN1(n10980), .IN2(n10981), .QN(n2670) );
  XNOR2X1 U10668 ( .IN1(n9844), .IN2(n4529), .Q(n10981) );
  NAND2X0 U10669 ( .IN1(n10982), .IN2(n10983), .QN(g30651) );
  INVX0 U10670 ( .INP(n10984), .ZN(n10983) );
  NOR2X0 U10671 ( .IN1(g6573), .IN2(n8452), .QN(n10984) );
  NAND2X0 U10672 ( .IN1(n10917), .IN2(g6573), .QN(n10982) );
  INVX0 U10673 ( .INP(n10985), .ZN(n10917) );
  NAND2X0 U10674 ( .IN1(n10986), .IN2(n10987), .QN(n10985) );
  NAND2X0 U10675 ( .IN1(n10834), .IN2(n4374), .QN(n10987) );
  NOR2X0 U10676 ( .IN1(n10836), .IN2(n10988), .QN(n10986) );
  NOR2X0 U10677 ( .IN1(n10989), .IN2(n10811), .QN(n10988) );
  XNOR2X1 U10678 ( .IN1(n9828), .IN2(n10990), .Q(n10989) );
  NOR2X0 U10679 ( .IN1(n10991), .IN2(n10992), .QN(n10836) );
  INVX0 U10680 ( .INP(n10993), .ZN(n10991) );
  NAND2X0 U10681 ( .IN1(n10994), .IN2(n10995), .QN(g30650) );
  NAND2X0 U10682 ( .IN1(test_so56), .IN2(n4515), .QN(n10995) );
  NAND2X0 U10683 ( .IN1(n10960), .IN2(g6782), .QN(n10994) );
  NAND2X0 U10684 ( .IN1(n10996), .IN2(n10997), .QN(g30649) );
  INVX0 U10685 ( .INP(n10998), .ZN(n10997) );
  NOR2X0 U10686 ( .IN1(g6368), .IN2(n8464), .QN(n10998) );
  NAND2X0 U10687 ( .IN1(n10920), .IN2(g6368), .QN(n10996) );
  INVX0 U10688 ( .INP(n10999), .ZN(n10920) );
  NAND2X0 U10689 ( .IN1(n11000), .IN2(n11001), .QN(n10999) );
  NAND2X0 U10690 ( .IN1(n10875), .IN2(n4391), .QN(n11001) );
  NOR2X0 U10691 ( .IN1(n10877), .IN2(n11002), .QN(n11000) );
  NOR2X0 U10692 ( .IN1(n11003), .IN2(n10850), .QN(n11002) );
  XNOR2X1 U10693 ( .IN1(n11004), .IN2(n11005), .Q(n11003) );
  NAND2X0 U10694 ( .IN1(n11006), .IN2(n11007), .QN(g30648) );
  INVX0 U10695 ( .INP(n11008), .ZN(n11007) );
  NOR2X0 U10696 ( .IN1(g6518), .IN2(n8488), .QN(n11008) );
  NAND2X0 U10697 ( .IN1(n10966), .IN2(g6518), .QN(n11006) );
  NAND2X0 U10698 ( .IN1(n11009), .IN2(n11010), .QN(g30647) );
  NAND2X0 U10699 ( .IN1(g915), .IN2(n9279), .QN(n11010) );
  NAND2X0 U10700 ( .IN1(test_so31), .IN2(n11011), .QN(n11009) );
  NAND2X0 U10701 ( .IN1(n11012), .IN2(n11013), .QN(g30646) );
  NAND2X0 U10702 ( .IN1(n4512), .IN2(g243), .QN(n11013) );
  NAND2X0 U10703 ( .IN1(n10970), .IN2(g6313), .QN(n11012) );
  NAND2X0 U10704 ( .IN1(n11014), .IN2(n11015), .QN(g30645) );
  INVX0 U10705 ( .INP(n11016), .ZN(n11015) );
  NOR2X0 U10706 ( .IN1(g165), .IN2(n8429), .QN(n11016) );
  NAND2X0 U10707 ( .IN1(n11017), .IN2(g165), .QN(n11014) );
  NAND2X0 U10708 ( .IN1(n11018), .IN2(n11019), .QN(g30644) );
  INVX0 U10709 ( .INP(n11020), .ZN(n11019) );
  NOR2X0 U10710 ( .IN1(g6573), .IN2(n8379), .QN(n11020) );
  NAND2X0 U10711 ( .IN1(n10960), .IN2(g6573), .QN(n11018) );
  NAND2X0 U10712 ( .IN1(n11021), .IN2(n10807), .QN(n10960) );
  NAND2X0 U10713 ( .IN1(n10993), .IN2(n11022), .QN(n10807) );
  NOR2X0 U10714 ( .IN1(n11023), .IN2(n11024), .QN(n11021) );
  NOR2X0 U10715 ( .IN1(n11025), .IN2(n10810), .QN(n11024) );
  INVX0 U10716 ( .INP(n10834), .ZN(n10810) );
  NOR2X0 U10717 ( .IN1(n10811), .IN2(n11026), .QN(n11023) );
  XNOR2X1 U10718 ( .IN1(n9816), .IN2(n2685), .Q(n11026) );
  NAND2X0 U10719 ( .IN1(n11027), .IN2(n11028), .QN(n2685) );
  XNOR2X1 U10720 ( .IN1(n11029), .IN2(n4530), .Q(n11028) );
  NAND2X0 U10721 ( .IN1(n11030), .IN2(n11031), .QN(g30643) );
  INVX0 U10722 ( .INP(n11032), .ZN(n11031) );
  NOR2X0 U10723 ( .IN1(g6368), .IN2(n8467), .QN(n11032) );
  NAND2X0 U10724 ( .IN1(n10966), .IN2(g6368), .QN(n11030) );
  INVX0 U10725 ( .INP(n11033), .ZN(n10966) );
  NAND2X0 U10726 ( .IN1(n11034), .IN2(n11035), .QN(n11033) );
  NAND2X0 U10727 ( .IN1(n10875), .IN2(n4375), .QN(n11035) );
  NOR2X0 U10728 ( .IN1(n10877), .IN2(n11036), .QN(n11034) );
  NOR2X0 U10729 ( .IN1(n11037), .IN2(n10850), .QN(n11036) );
  XNOR2X1 U10730 ( .IN1(n9781), .IN2(n11038), .Q(n11037) );
  NOR2X0 U10731 ( .IN1(n11039), .IN2(n11040), .QN(n10877) );
  INVX0 U10732 ( .INP(n11041), .ZN(n11039) );
  NAND2X0 U10733 ( .IN1(n11042), .IN2(n11043), .QN(g30642) );
  INVX0 U10734 ( .INP(n11044), .ZN(n11043) );
  NOR2X0 U10735 ( .IN1(g6518), .IN2(n8492), .QN(n11044) );
  NAND2X0 U10736 ( .IN1(n11011), .IN2(g6518), .QN(n11042) );
  NAND2X0 U10737 ( .IN1(n11045), .IN2(n11046), .QN(g30641) );
  INVX0 U10738 ( .INP(n11047), .ZN(n11046) );
  NOR2X0 U10739 ( .IN1(g6231), .IN2(n8478), .QN(n11047) );
  NAND2X0 U10740 ( .IN1(n10970), .IN2(g6231), .QN(n11045) );
  INVX0 U10741 ( .INP(n11048), .ZN(n10970) );
  NAND2X0 U10742 ( .IN1(n11049), .IN2(n11050), .QN(n11048) );
  NAND2X0 U10743 ( .IN1(n10927), .IN2(n4392), .QN(n11050) );
  NOR2X0 U10744 ( .IN1(n10929), .IN2(n11051), .QN(n11049) );
  NOR2X0 U10745 ( .IN1(n11052), .IN2(n10894), .QN(n11051) );
  XNOR2X1 U10746 ( .IN1(n9754), .IN2(n11053), .Q(n11052) );
  NAND2X0 U10747 ( .IN1(n11054), .IN2(n11055), .QN(g30640) );
  NAND2X0 U10748 ( .IN1(n4512), .IN2(g234), .QN(n11055) );
  NAND2X0 U10749 ( .IN1(n11017), .IN2(g6313), .QN(n11054) );
  NAND2X0 U10750 ( .IN1(n11056), .IN2(n11057), .QN(g30639) );
  INVX0 U10751 ( .INP(n11058), .ZN(n11057) );
  NOR2X0 U10752 ( .IN1(g165), .IN2(n8386), .QN(n11058) );
  NAND2X0 U10753 ( .IN1(n11059), .IN2(g165), .QN(n11056) );
  NAND2X0 U10754 ( .IN1(n11060), .IN2(n11061), .QN(g30638) );
  INVX0 U10755 ( .INP(n11062), .ZN(n11061) );
  NOR2X0 U10756 ( .IN1(g6368), .IN2(n8456), .QN(n11062) );
  NAND2X0 U10757 ( .IN1(n11011), .IN2(g6368), .QN(n11060) );
  NAND2X0 U10758 ( .IN1(n11063), .IN2(n10846), .QN(n11011) );
  NAND2X0 U10759 ( .IN1(n11041), .IN2(n11040), .QN(n10846) );
  NOR2X0 U10760 ( .IN1(n11064), .IN2(n11065), .QN(n11063) );
  NOR2X0 U10761 ( .IN1(n11066), .IN2(n10849), .QN(n11065) );
  INVX0 U10762 ( .INP(n10875), .ZN(n10849) );
  NOR2X0 U10763 ( .IN1(n10850), .IN2(n11067), .QN(n11064) );
  XNOR2X1 U10764 ( .IN1(n10881), .IN2(n9795), .Q(n11067) );
  INVX0 U10765 ( .INP(n11068), .ZN(n10881) );
  NAND2X0 U10766 ( .IN1(n11069), .IN2(n11070), .QN(n11068) );
  XNOR2X1 U10767 ( .IN1(n11071), .IN2(n10883), .Q(n11070) );
  INVX0 U10768 ( .INP(n11072), .ZN(n10850) );
  NAND2X0 U10769 ( .IN1(n11073), .IN2(n11074), .QN(g30637) );
  INVX0 U10770 ( .INP(n11075), .ZN(n11074) );
  NOR2X0 U10771 ( .IN1(g6231), .IN2(n8481), .QN(n11075) );
  NAND2X0 U10772 ( .IN1(n11017), .IN2(g6231), .QN(n11073) );
  INVX0 U10773 ( .INP(n11076), .ZN(n11017) );
  NAND2X0 U10774 ( .IN1(n11077), .IN2(n11078), .QN(n11076) );
  NAND2X0 U10775 ( .IN1(n10927), .IN2(n4376), .QN(n11078) );
  NOR2X0 U10776 ( .IN1(n10929), .IN2(n11079), .QN(n11077) );
  NOR2X0 U10777 ( .IN1(n11080), .IN2(n10894), .QN(n11079) );
  XNOR2X1 U10778 ( .IN1(n9739), .IN2(n11081), .Q(n11080) );
  NOR2X0 U10779 ( .IN1(n11082), .IN2(n11083), .QN(n10929) );
  INVX0 U10780 ( .INP(n11084), .ZN(n11082) );
  NAND2X0 U10781 ( .IN1(n11085), .IN2(n11086), .QN(g30636) );
  NAND2X0 U10782 ( .IN1(n4512), .IN2(g225), .QN(n11086) );
  NAND2X0 U10783 ( .IN1(n11059), .IN2(g6313), .QN(n11085) );
  NAND2X0 U10784 ( .IN1(n11087), .IN2(n11088), .QN(g30635) );
  INVX0 U10785 ( .INP(n11089), .ZN(n11088) );
  NOR2X0 U10786 ( .IN1(g6231), .IN2(n8380), .QN(n11089) );
  NAND2X0 U10787 ( .IN1(n11059), .IN2(g6231), .QN(n11087) );
  NAND2X0 U10788 ( .IN1(n11090), .IN2(n10890), .QN(n11059) );
  NAND2X0 U10789 ( .IN1(n11084), .IN2(n11083), .QN(n10890) );
  NOR2X0 U10790 ( .IN1(n11091), .IN2(n11092), .QN(n11090) );
  NOR2X0 U10791 ( .IN1(n11093), .IN2(n10893), .QN(n11092) );
  INVX0 U10792 ( .INP(n10927), .ZN(n10893) );
  NOR2X0 U10793 ( .IN1(n10894), .IN2(n11094), .QN(n11091) );
  XNOR2X1 U10794 ( .IN1(n9746), .IN2(n2718), .Q(n11094) );
  NAND2X0 U10795 ( .IN1(n11095), .IN2(n11096), .QN(n2718) );
  XNOR2X1 U10796 ( .IN1(n9740), .IN2(n10501), .Q(n11096) );
  INVX0 U10797 ( .INP(n11097), .ZN(n10894) );
  NAND2X0 U10798 ( .IN1(n11098), .IN2(n11099), .QN(g30566) );
  NAND2X0 U10799 ( .IN1(n10667), .IN2(n4606), .QN(n11099) );
  NOR2X0 U10800 ( .IN1(n11100), .IN2(n11101), .QN(n10667) );
  XNOR2X1 U10801 ( .IN1(n11102), .IN2(n11103), .Q(n11100) );
  NOR2X0 U10802 ( .IN1(n11104), .IN2(n11105), .QN(n11103) );
  NOR2X0 U10803 ( .IN1(n11106), .IN2(n11107), .QN(n11105) );
  NOR2X0 U10804 ( .IN1(n11108), .IN2(n11109), .QN(n11107) );
  NOR2X0 U10805 ( .IN1(n11110), .IN2(n11111), .QN(n11109) );
  NOR2X0 U10806 ( .IN1(n11112), .IN2(n11113), .QN(n11111) );
  NOR2X0 U10807 ( .IN1(n11114), .IN2(n11115), .QN(n11113) );
  NAND2X0 U10808 ( .IN1(n11116), .IN2(n11117), .QN(n11115) );
  NOR2X0 U10809 ( .IN1(n11118), .IN2(n11119), .QN(n11116) );
  NOR2X0 U10810 ( .IN1(n2792), .IN2(n11120), .QN(n11119) );
  INVX0 U10811 ( .INP(n11121), .ZN(n11120) );
  INVX0 U10812 ( .INP(n11122), .ZN(n11118) );
  NOR2X0 U10813 ( .IN1(n11123), .IN2(n11124), .QN(n11112) );
  NAND2X0 U10814 ( .IN1(n2792), .IN2(n10479), .QN(n11124) );
  NOR2X0 U10815 ( .IN1(n11102), .IN2(n11125), .QN(n11108) );
  NOR2X0 U10816 ( .IN1(n11126), .IN2(n11127), .QN(n11125) );
  NOR2X0 U10817 ( .IN1(n11128), .IN2(n11129), .QN(n11126) );
  NOR2X0 U10818 ( .IN1(n11114), .IN2(n11130), .QN(n11128) );
  NAND2X0 U10819 ( .IN1(n11131), .IN2(n11122), .QN(n11130) );
  NOR2X0 U10820 ( .IN1(n11132), .IN2(n11133), .QN(n11104) );
  NAND2X0 U10821 ( .IN1(n4509), .IN2(g2392), .QN(n11098) );
  NAND2X0 U10822 ( .IN1(n11134), .IN2(n11135), .QN(g30505) );
  NAND2X0 U10823 ( .IN1(n11136), .IN2(g5555), .QN(n11135) );
  NAND2X0 U10824 ( .IN1(n4516), .IN2(g2393), .QN(n11134) );
  NAND2X0 U10825 ( .IN1(n11137), .IN2(n11138), .QN(g30503) );
  NAND2X0 U10826 ( .IN1(n11139), .IN2(g7014), .QN(n11138) );
  INVX0 U10827 ( .INP(n11140), .ZN(n11137) );
  NOR2X0 U10828 ( .IN1(n10678), .IN2(n8496), .QN(n11140) );
  NAND2X0 U10829 ( .IN1(n11141), .IN2(n11142), .QN(g30500) );
  NAND2X0 U10830 ( .IN1(n2798), .IN2(g1088), .QN(n11142) );
  NAND2X0 U10831 ( .IN1(test_so39), .IN2(n4381), .QN(n11141) );
  NAND2X0 U10832 ( .IN1(n11143), .IN2(n11144), .QN(g30487) );
  NAND2X0 U10833 ( .IN1(n11139), .IN2(g5511), .QN(n11144) );
  NAND2X0 U10834 ( .IN1(n4518), .IN2(g1699), .QN(n11143) );
  NAND2X0 U10835 ( .IN1(n11145), .IN2(n11146), .QN(g30485) );
  NAND2X0 U10836 ( .IN1(n4364), .IN2(g1006), .QN(n11146) );
  NAND2X0 U10837 ( .IN1(n2798), .IN2(g6712), .QN(n11145) );
  NAND2X0 U10838 ( .IN1(n11147), .IN2(n11148), .QN(g30482) );
  NAND2X0 U10839 ( .IN1(n11149), .IN2(n4640), .QN(n11148) );
  NAND2X0 U10840 ( .IN1(n4506), .IN2(g320), .QN(n11147) );
  NAND2X0 U10841 ( .IN1(n11150), .IN2(n11151), .QN(g30470) );
  NAND2X0 U10842 ( .IN1(n4363), .IN2(g1005), .QN(n11151) );
  NAND2X0 U10843 ( .IN1(n2798), .IN2(g5472), .QN(n11150) );
  NAND2X0 U10844 ( .IN1(n11152), .IN2(n11153), .QN(g30468) );
  NAND2X0 U10845 ( .IN1(n11149), .IN2(g6447), .QN(n11153) );
  NAND2X0 U10846 ( .IN1(n4499), .IN2(g319), .QN(n11152) );
  NAND2X0 U10847 ( .IN1(n11154), .IN2(n11155), .QN(g30455) );
  NAND2X0 U10848 ( .IN1(n11149), .IN2(g5437), .QN(n11155) );
  NOR2X0 U10849 ( .IN1(n11156), .IN2(n10724), .QN(n11149) );
  XNOR2X1 U10850 ( .IN1(n11157), .IN2(n11158), .Q(n11156) );
  NAND2X0 U10851 ( .IN1(n11159), .IN2(n11160), .QN(n11157) );
  NAND2X0 U10852 ( .IN1(n11158), .IN2(n11161), .QN(n11160) );
  NAND2X0 U10853 ( .IN1(n11162), .IN2(n10750), .QN(n11161) );
  NOR2X0 U10854 ( .IN1(n11163), .IN2(n11164), .QN(n11162) );
  NOR2X0 U10855 ( .IN1(n10746), .IN2(n11165), .QN(n11164) );
  NAND2X0 U10856 ( .IN1(n11166), .IN2(g309), .QN(n11165) );
  NOR2X0 U10857 ( .IN1(n10725), .IN2(n11167), .QN(n11163) );
  NOR2X0 U10858 ( .IN1(n11168), .IN2(n10733), .QN(n11167) );
  NOR2X0 U10859 ( .IN1(n10741), .IN2(n10748), .QN(n11168) );
  NAND2X0 U10860 ( .IN1(n11169), .IN2(n10739), .QN(n11159) );
  NOR2X0 U10861 ( .IN1(n11170), .IN2(n11171), .QN(n11169) );
  NAND2X0 U10862 ( .IN1(n10750), .IN2(n10746), .QN(n11170) );
  INVX0 U10863 ( .INP(n11172), .ZN(n11154) );
  NOR2X0 U10864 ( .IN1(n10752), .IN2(n8521), .QN(n11172) );
  NAND2X0 U10865 ( .IN1(n11173), .IN2(n11174), .QN(g30356) );
  NAND2X0 U10866 ( .IN1(n11136), .IN2(n4606), .QN(n11174) );
  NAND2X0 U10867 ( .IN1(n4509), .IN2(g2395), .QN(n11173) );
  NAND2X0 U10868 ( .IN1(n11175), .IN2(n11176), .QN(g30341) );
  NAND2X0 U10869 ( .IN1(n11136), .IN2(g7264), .QN(n11176) );
  NOR2X0 U10870 ( .IN1(n11177), .IN2(n11101), .QN(n11136) );
  XNOR2X1 U10871 ( .IN1(n11178), .IN2(n11123), .Q(n11177) );
  NAND2X0 U10872 ( .IN1(n11179), .IN2(n11180), .QN(n11178) );
  NAND2X0 U10873 ( .IN1(n11123), .IN2(n11181), .QN(n11180) );
  NAND2X0 U10874 ( .IN1(n11182), .IN2(n11133), .QN(n11181) );
  NOR2X0 U10875 ( .IN1(n11183), .IN2(n11184), .QN(n11182) );
  NOR2X0 U10876 ( .IN1(n11110), .IN2(n11185), .QN(n11184) );
  INVX0 U10877 ( .INP(n11186), .ZN(n11185) );
  NOR2X0 U10878 ( .IN1(n11187), .IN2(n9281), .QN(n11186) );
  NOR2X0 U10879 ( .IN1(n11102), .IN2(n11117), .QN(n11183) );
  NOR2X0 U10880 ( .IN1(n11188), .IN2(n11189), .QN(n11117) );
  NOR2X0 U10881 ( .IN1(n11131), .IN2(n11127), .QN(n11189) );
  NAND2X0 U10882 ( .IN1(n11190), .IN2(n11114), .QN(n11179) );
  NOR2X0 U10883 ( .IN1(n11191), .IN2(n11192), .QN(n11190) );
  NAND2X0 U10884 ( .IN1(n11133), .IN2(n11110), .QN(n11191) );
  INVX0 U10885 ( .INP(n11193), .ZN(n11175) );
  NOR2X0 U10886 ( .IN1(n10669), .IN2(n8493), .QN(n11193) );
  NAND2X0 U10887 ( .IN1(n11194), .IN2(n11195), .QN(g30338) );
  NAND2X0 U10888 ( .IN1(n11139), .IN2(n4618), .QN(n11195) );
  NOR2X0 U10889 ( .IN1(n11196), .IN2(n10685), .QN(n11139) );
  XNOR2X1 U10890 ( .IN1(n11197), .IN2(n11198), .Q(n11196) );
  NAND2X0 U10891 ( .IN1(n11199), .IN2(n11200), .QN(n11197) );
  NAND2X0 U10892 ( .IN1(n11198), .IN2(n11201), .QN(n11200) );
  NAND2X0 U10893 ( .IN1(n11202), .IN2(n10711), .QN(n11201) );
  NOR2X0 U10894 ( .IN1(n11203), .IN2(n11204), .QN(n11202) );
  NOR2X0 U10895 ( .IN1(n10707), .IN2(n11205), .QN(n11204) );
  NAND2X0 U10896 ( .IN1(n11206), .IN2(g1690), .QN(n11205) );
  NOR2X0 U10897 ( .IN1(n10686), .IN2(n11207), .QN(n11203) );
  NOR2X0 U10898 ( .IN1(n11208), .IN2(n10694), .QN(n11207) );
  NOR2X0 U10899 ( .IN1(n10702), .IN2(n10709), .QN(n11208) );
  NAND2X0 U10900 ( .IN1(n11209), .IN2(n10700), .QN(n11199) );
  NOR2X0 U10901 ( .IN1(n11210), .IN2(n11211), .QN(n11209) );
  NAND2X0 U10902 ( .IN1(n10711), .IN2(n10707), .QN(n11210) );
  NAND2X0 U10903 ( .IN1(n4511), .IN2(g1701), .QN(n11194) );
  NAND2X0 U10904 ( .IN1(n11212), .IN2(n11213), .QN(g30304) );
  INVX0 U10905 ( .INP(n11214), .ZN(n11213) );
  NOR2X0 U10906 ( .IN1(g2241), .IN2(n8530), .QN(n11214) );
  NAND2X0 U10907 ( .IN1(n11215), .IN2(g2241), .QN(n11212) );
  NAND2X0 U10908 ( .IN1(n11216), .IN2(n11217), .QN(g30303) );
  NAND2X0 U10909 ( .IN1(g2282), .IN2(n9278), .QN(n11217) );
  NAND2X0 U10910 ( .IN1(test_so73), .IN2(n11215), .QN(n11216) );
  NAND2X0 U10911 ( .IN1(n11218), .IN2(n11219), .QN(g30302) );
  INVX0 U10912 ( .INP(n11220), .ZN(n11219) );
  NOR2X0 U10913 ( .IN1(g1547), .IN2(n8531), .QN(n11220) );
  NAND2X0 U10914 ( .IN1(n11221), .IN2(g1547), .QN(n11218) );
  NAND2X0 U10915 ( .IN1(n11222), .IN2(n11223), .QN(g30301) );
  INVX0 U10916 ( .INP(n11224), .ZN(n11223) );
  NOR2X0 U10917 ( .IN1(g6837), .IN2(n8436), .QN(n11224) );
  NAND2X0 U10918 ( .IN1(n11215), .IN2(g6837), .QN(n11222) );
  NAND2X0 U10919 ( .IN1(n11225), .IN2(n11226), .QN(n11215) );
  NAND2X0 U10920 ( .IN1(n11227), .IN2(n11228), .QN(n11226) );
  XNOR2X1 U10921 ( .IN1(n11229), .IN2(n9852), .Q(n11227) );
  NAND2X0 U10922 ( .IN1(n10795), .IN2(g2185), .QN(n11225) );
  NAND2X0 U10923 ( .IN1(n11230), .IN2(n11231), .QN(g30300) );
  INVX0 U10924 ( .INP(n11232), .ZN(n11231) );
  NOR2X0 U10925 ( .IN1(g2241), .IN2(n8537), .QN(n11232) );
  NAND2X0 U10926 ( .IN1(n11233), .IN2(g2241), .QN(n11230) );
  NAND2X0 U10927 ( .IN1(n11234), .IN2(n11235), .QN(g30299) );
  NAND2X0 U10928 ( .IN1(n4515), .IN2(g1588), .QN(n11235) );
  NAND2X0 U10929 ( .IN1(n11221), .IN2(g6782), .QN(n11234) );
  NAND2X0 U10930 ( .IN1(n11236), .IN2(n11237), .QN(g30298) );
  NAND2X0 U10931 ( .IN1(g897), .IN2(n9279), .QN(n11237) );
  NAND2X0 U10932 ( .IN1(test_so31), .IN2(n11238), .QN(n11236) );
  NAND2X0 U10933 ( .IN1(n11239), .IN2(n11240), .QN(g30297) );
  INVX0 U10934 ( .INP(n11241), .ZN(n11240) );
  NOR2X0 U10935 ( .IN1(g2241), .IN2(n8527), .QN(n11241) );
  NAND2X0 U10936 ( .IN1(n11242), .IN2(g2241), .QN(n11239) );
  NAND2X0 U10937 ( .IN1(n11243), .IN2(n11244), .QN(g30296) );
  NAND2X0 U10938 ( .IN1(test_so76), .IN2(n9278), .QN(n11244) );
  NAND2X0 U10939 ( .IN1(test_so73), .IN2(n11233), .QN(n11243) );
  NAND2X0 U10940 ( .IN1(n11245), .IN2(n11246), .QN(g30295) );
  INVX0 U10941 ( .INP(n11247), .ZN(n11246) );
  NOR2X0 U10942 ( .IN1(g6573), .IN2(n8449), .QN(n11247) );
  NAND2X0 U10943 ( .IN1(n11221), .IN2(g6573), .QN(n11245) );
  NAND2X0 U10944 ( .IN1(n11248), .IN2(n11249), .QN(n11221) );
  NAND2X0 U10945 ( .IN1(n11250), .IN2(n11251), .QN(n11249) );
  XNOR2X1 U10946 ( .IN1(n11252), .IN2(n9817), .Q(n11250) );
  NAND2X0 U10947 ( .IN1(n10834), .IN2(g1491), .QN(n11248) );
  NAND2X0 U10948 ( .IN1(n11253), .IN2(n11254), .QN(g30294) );
  INVX0 U10949 ( .INP(n11255), .ZN(n11254) );
  NOR2X0 U10950 ( .IN1(g1547), .IN2(n8540), .QN(n11255) );
  NAND2X0 U10951 ( .IN1(n11256), .IN2(g1547), .QN(n11253) );
  NAND2X0 U10952 ( .IN1(n11257), .IN2(n11258), .QN(g30293) );
  INVX0 U10953 ( .INP(n11259), .ZN(n11258) );
  NOR2X0 U10954 ( .IN1(g6518), .IN2(n8462), .QN(n11259) );
  NAND2X0 U10955 ( .IN1(n11238), .IN2(g6518), .QN(n11257) );
  NAND2X0 U10956 ( .IN1(n11260), .IN2(n11261), .QN(g30292) );
  INVX0 U10957 ( .INP(n11262), .ZN(n11261) );
  NOR2X0 U10958 ( .IN1(g165), .IN2(n8534), .QN(n11262) );
  NAND2X0 U10959 ( .IN1(n11263), .IN2(g165), .QN(n11260) );
  NAND2X0 U10960 ( .IN1(n11264), .IN2(n11265), .QN(g30291) );
  NAND2X0 U10961 ( .IN1(g2336), .IN2(n9278), .QN(n11265) );
  NAND2X0 U10962 ( .IN1(test_so73), .IN2(n11242), .QN(n11264) );
  NAND2X0 U10963 ( .IN1(n11266), .IN2(n11267), .QN(g30290) );
  INVX0 U10964 ( .INP(n11268), .ZN(n11267) );
  NOR2X0 U10965 ( .IN1(g2241), .IN2(n8418), .QN(n11268) );
  NAND2X0 U10966 ( .IN1(n11269), .IN2(g2241), .QN(n11266) );
  NAND2X0 U10967 ( .IN1(n11270), .IN2(n11271), .QN(g30289) );
  INVX0 U10968 ( .INP(n11272), .ZN(n11271) );
  NOR2X0 U10969 ( .IN1(g6837), .IN2(n8441), .QN(n11272) );
  NAND2X0 U10970 ( .IN1(n11233), .IN2(g6837), .QN(n11270) );
  NAND2X0 U10971 ( .IN1(n11273), .IN2(n11274), .QN(n11233) );
  NAND2X0 U10972 ( .IN1(n11228), .IN2(n11275), .QN(n11274) );
  XNOR2X1 U10973 ( .IN1(n11276), .IN2(n9845), .Q(n11275) );
  NAND2X0 U10974 ( .IN1(n10795), .IN2(g2165), .QN(n11273) );
  NAND2X0 U10975 ( .IN1(n11277), .IN2(n11278), .QN(g30288) );
  INVX0 U10976 ( .INP(n11279), .ZN(n11278) );
  NOR2X0 U10977 ( .IN1(g1547), .IN2(n8528), .QN(n11279) );
  NAND2X0 U10978 ( .IN1(n11280), .IN2(g1547), .QN(n11277) );
  NAND2X0 U10979 ( .IN1(n11281), .IN2(n11282), .QN(g30287) );
  NAND2X0 U10980 ( .IN1(n4515), .IN2(g1570), .QN(n11282) );
  NAND2X0 U10981 ( .IN1(n11256), .IN2(g6782), .QN(n11281) );
  NAND2X0 U10982 ( .IN1(n11283), .IN2(n11284), .QN(g30286) );
  INVX0 U10983 ( .INP(n11285), .ZN(n11284) );
  NOR2X0 U10984 ( .IN1(g6368), .IN2(n8463), .QN(n11285) );
  NAND2X0 U10985 ( .IN1(n11238), .IN2(g6368), .QN(n11283) );
  NAND2X0 U10986 ( .IN1(n11286), .IN2(n11287), .QN(n11238) );
  NAND2X0 U10987 ( .IN1(n11288), .IN2(n11072), .QN(n11287) );
  XNOR2X1 U10988 ( .IN1(n11289), .IN2(n9775), .Q(n11288) );
  NAND2X0 U10989 ( .IN1(n10875), .IN2(g801), .QN(n11286) );
  NAND2X0 U10990 ( .IN1(n11290), .IN2(n11291), .QN(g30285) );
  NAND2X0 U10991 ( .IN1(g879), .IN2(n9279), .QN(n11291) );
  NAND2X0 U10992 ( .IN1(test_so31), .IN2(n11292), .QN(n11290) );
  NAND2X0 U10993 ( .IN1(n11293), .IN2(n11294), .QN(g30284) );
  NAND2X0 U10994 ( .IN1(n4512), .IN2(g207), .QN(n11294) );
  NAND2X0 U10995 ( .IN1(n11263), .IN2(g6313), .QN(n11293) );
  NAND2X0 U10996 ( .IN1(n11295), .IN2(n11296), .QN(g30283) );
  INVX0 U10997 ( .INP(n11297), .ZN(n11296) );
  NOR2X0 U10998 ( .IN1(g6837), .IN2(n8431), .QN(n11297) );
  NAND2X0 U10999 ( .IN1(n11242), .IN2(g6837), .QN(n11295) );
  NAND2X0 U11000 ( .IN1(n11298), .IN2(n11299), .QN(n11242) );
  NAND2X0 U11001 ( .IN1(n11300), .IN2(n11301), .QN(n11299) );
  XOR2X1 U11002 ( .IN1(n10980), .IN2(n9844), .Q(n11301) );
  NOR2X0 U11003 ( .IN1(n11302), .IN2(n11303), .QN(n10980) );
  XNOR2X1 U11004 ( .IN1(n11304), .IN2(n10503), .Q(n11303) );
  NAND2X0 U11005 ( .IN1(n10795), .IN2(g2200), .QN(n11298) );
  NAND2X0 U11006 ( .IN1(n11305), .IN2(n11306), .QN(g30282) );
  NAND2X0 U11007 ( .IN1(test_so77), .IN2(n9278), .QN(n11306) );
  NAND2X0 U11008 ( .IN1(test_so73), .IN2(n11269), .QN(n11305) );
  NAND2X0 U11009 ( .IN1(n11307), .IN2(n11308), .QN(g30281) );
  NAND2X0 U11010 ( .IN1(n4515), .IN2(g1642), .QN(n11308) );
  NAND2X0 U11011 ( .IN1(n11280), .IN2(g6782), .QN(n11307) );
  NAND2X0 U11012 ( .IN1(n11309), .IN2(n11310), .QN(g30280) );
  INVX0 U11013 ( .INP(n11311), .ZN(n11310) );
  NOR2X0 U11014 ( .IN1(g1547), .IN2(n8421), .QN(n11311) );
  NAND2X0 U11015 ( .IN1(n11312), .IN2(g1547), .QN(n11309) );
  NAND2X0 U11016 ( .IN1(n11313), .IN2(n11314), .QN(g30279) );
  INVX0 U11017 ( .INP(n11315), .ZN(n11314) );
  NOR2X0 U11018 ( .IN1(g6573), .IN2(n8454), .QN(n11315) );
  NAND2X0 U11019 ( .IN1(n11256), .IN2(g6573), .QN(n11313) );
  NAND2X0 U11020 ( .IN1(n11316), .IN2(n11317), .QN(n11256) );
  NAND2X0 U11021 ( .IN1(n11251), .IN2(n11318), .QN(n11317) );
  XNOR2X1 U11022 ( .IN1(n11319), .IN2(n11320), .Q(n11318) );
  NAND2X0 U11023 ( .IN1(n10834), .IN2(g1471), .QN(n11316) );
  NAND2X0 U11024 ( .IN1(n11321), .IN2(n11322), .QN(g30278) );
  NAND2X0 U11025 ( .IN1(g951), .IN2(n9279), .QN(n11322) );
  NAND2X0 U11026 ( .IN1(test_so31), .IN2(n11323), .QN(n11321) );
  NAND2X0 U11027 ( .IN1(n11324), .IN2(n11325), .QN(g30277) );
  INVX0 U11028 ( .INP(n11326), .ZN(n11325) );
  NOR2X0 U11029 ( .IN1(g6518), .IN2(n8468), .QN(n11326) );
  NAND2X0 U11030 ( .IN1(n11292), .IN2(g6518), .QN(n11324) );
  NAND2X0 U11031 ( .IN1(n11327), .IN2(n11328), .QN(g30276) );
  INVX0 U11032 ( .INP(n11329), .ZN(n11328) );
  NOR2X0 U11033 ( .IN1(g6231), .IN2(n8477), .QN(n11329) );
  NAND2X0 U11034 ( .IN1(n11263), .IN2(g6231), .QN(n11327) );
  NAND2X0 U11035 ( .IN1(n11330), .IN2(n11331), .QN(n11263) );
  NAND2X0 U11036 ( .IN1(n11332), .IN2(n11097), .QN(n11331) );
  XNOR2X1 U11037 ( .IN1(n11333), .IN2(n9747), .Q(n11332) );
  NAND2X0 U11038 ( .IN1(n10927), .IN2(g113), .QN(n11330) );
  NAND2X0 U11039 ( .IN1(n11334), .IN2(n11335), .QN(g30275) );
  INVX0 U11040 ( .INP(n11336), .ZN(n11335) );
  NOR2X0 U11041 ( .IN1(g165), .IN2(n8546), .QN(n11336) );
  NAND2X0 U11042 ( .IN1(n11337), .IN2(g165), .QN(n11334) );
  NAND2X0 U11043 ( .IN1(n11338), .IN2(n11339), .QN(g30274) );
  INVX0 U11044 ( .INP(n11340), .ZN(n11339) );
  NOR2X0 U11045 ( .IN1(g6837), .IN2(n8434), .QN(n11340) );
  NAND2X0 U11046 ( .IN1(n11269), .IN2(g6837), .QN(n11338) );
  NAND2X0 U11047 ( .IN1(n11341), .IN2(n11342), .QN(n11269) );
  NAND2X0 U11048 ( .IN1(n11300), .IN2(n11343), .QN(n11342) );
  XNOR2X1 U11049 ( .IN1(n11344), .IN2(n9865), .Q(n11343) );
  NAND2X0 U11050 ( .IN1(n11345), .IN2(n11346), .QN(n11344) );
  NAND2X0 U11051 ( .IN1(n10503), .IN2(n9852), .QN(n11346) );
  NOR2X0 U11052 ( .IN1(n10943), .IN2(n10777), .QN(n11300) );
  INVX0 U11053 ( .INP(n11228), .ZN(n10777) );
  NAND2X0 U11054 ( .IN1(n10795), .IN2(g2190), .QN(n11341) );
  NAND2X0 U11055 ( .IN1(n11347), .IN2(n11348), .QN(g30273) );
  INVX0 U11056 ( .INP(n11349), .ZN(n11348) );
  NOR2X0 U11057 ( .IN1(g6573), .IN2(n8443), .QN(n11349) );
  NAND2X0 U11058 ( .IN1(n11280), .IN2(g6573), .QN(n11347) );
  NAND2X0 U11059 ( .IN1(n11350), .IN2(n11351), .QN(n11280) );
  NAND2X0 U11060 ( .IN1(n11352), .IN2(n11353), .QN(n11351) );
  XNOR2X1 U11061 ( .IN1(n9809), .IN2(n11027), .Q(n11353) );
  NOR2X0 U11062 ( .IN1(n11354), .IN2(n11355), .QN(n11027) );
  XNOR2X1 U11063 ( .IN1(n9808), .IN2(n4530), .Q(n11355) );
  NAND2X0 U11064 ( .IN1(n10834), .IN2(g1506), .QN(n11350) );
  NAND2X0 U11065 ( .IN1(n11356), .IN2(n11357), .QN(g30272) );
  NAND2X0 U11066 ( .IN1(n4515), .IN2(g1633), .QN(n11357) );
  NAND2X0 U11067 ( .IN1(n11312), .IN2(g6782), .QN(n11356) );
  NAND2X0 U11068 ( .IN1(n11358), .IN2(n11359), .QN(g30271) );
  INVX0 U11069 ( .INP(n11360), .ZN(n11359) );
  NOR2X0 U11070 ( .IN1(g6518), .IN2(n8457), .QN(n11360) );
  NAND2X0 U11071 ( .IN1(n11323), .IN2(g6518), .QN(n11358) );
  NAND2X0 U11072 ( .IN1(n11361), .IN2(n11362), .QN(g30270) );
  NAND2X0 U11073 ( .IN1(g942), .IN2(n9279), .QN(n11362) );
  NAND2X0 U11074 ( .IN1(test_so31), .IN2(n11363), .QN(n11361) );
  NAND2X0 U11075 ( .IN1(n11364), .IN2(n11365), .QN(g30269) );
  INVX0 U11076 ( .INP(n11366), .ZN(n11365) );
  NOR2X0 U11077 ( .IN1(g6368), .IN2(n8469), .QN(n11366) );
  NAND2X0 U11078 ( .IN1(n11292), .IN2(g6368), .QN(n11364) );
  NAND2X0 U11079 ( .IN1(n11367), .IN2(n11368), .QN(n11292) );
  NAND2X0 U11080 ( .IN1(n11072), .IN2(n11369), .QN(n11368) );
  XNOR2X1 U11081 ( .IN1(n11370), .IN2(n9780), .Q(n11369) );
  NAND2X0 U11082 ( .IN1(n10875), .IN2(g785), .QN(n11367) );
  NAND2X0 U11083 ( .IN1(n11371), .IN2(n11372), .QN(g30268) );
  INVX0 U11084 ( .INP(n11373), .ZN(n11372) );
  NOR2X0 U11085 ( .IN1(g165), .IN2(n8529), .QN(n11373) );
  NAND2X0 U11086 ( .IN1(n11374), .IN2(g165), .QN(n11371) );
  NAND2X0 U11087 ( .IN1(n11375), .IN2(n11376), .QN(g30267) );
  NAND2X0 U11088 ( .IN1(test_so13), .IN2(n4512), .QN(n11376) );
  NAND2X0 U11089 ( .IN1(n11337), .IN2(g6313), .QN(n11375) );
  NAND2X0 U11090 ( .IN1(n11377), .IN2(n11378), .QN(g30266) );
  INVX0 U11091 ( .INP(n11379), .ZN(n11378) );
  NOR2X0 U11092 ( .IN1(g6573), .IN2(n8447), .QN(n11379) );
  NAND2X0 U11093 ( .IN1(n11312), .IN2(g6573), .QN(n11377) );
  NAND2X0 U11094 ( .IN1(n11380), .IN2(n11381), .QN(n11312) );
  NAND2X0 U11095 ( .IN1(n11352), .IN2(n11382), .QN(n11381) );
  XNOR2X1 U11096 ( .IN1(n11383), .IN2(n11384), .Q(n11382) );
  NAND2X0 U11097 ( .IN1(n11385), .IN2(n11386), .QN(n11383) );
  NAND2X0 U11098 ( .IN1(n10992), .IN2(n9817), .QN(n11386) );
  NOR2X0 U11099 ( .IN1(n10993), .IN2(n10811), .QN(n11352) );
  INVX0 U11100 ( .INP(n11251), .ZN(n10811) );
  NAND2X0 U11101 ( .IN1(n10834), .IN2(g1496), .QN(n11380) );
  NAND2X0 U11102 ( .IN1(n11387), .IN2(n11388), .QN(g30265) );
  NAND2X0 U11103 ( .IN1(test_so35), .IN2(n4323), .QN(n11388) );
  NAND2X0 U11104 ( .IN1(n11323), .IN2(g6368), .QN(n11387) );
  NAND2X0 U11105 ( .IN1(n11389), .IN2(n11390), .QN(n11323) );
  NAND2X0 U11106 ( .IN1(n11391), .IN2(n11072), .QN(n11390) );
  XNOR2X1 U11107 ( .IN1(n9788), .IN2(n11069), .Q(n11391) );
  NOR2X0 U11108 ( .IN1(n11392), .IN2(n11393), .QN(n11069) );
  XNOR2X1 U11109 ( .IN1(n9773), .IN2(n10883), .Q(n11393) );
  NAND2X0 U11110 ( .IN1(n10875), .IN2(g813), .QN(n11389) );
  NAND2X0 U11111 ( .IN1(n11394), .IN2(n11395), .QN(g30264) );
  INVX0 U11112 ( .INP(n11396), .ZN(n11395) );
  NOR2X0 U11113 ( .IN1(g6518), .IN2(n8460), .QN(n11396) );
  NAND2X0 U11114 ( .IN1(n11363), .IN2(g6518), .QN(n11394) );
  NAND2X0 U11115 ( .IN1(n11397), .IN2(n11398), .QN(g30263) );
  NAND2X0 U11116 ( .IN1(n4512), .IN2(g261), .QN(n11398) );
  NAND2X0 U11117 ( .IN1(n11374), .IN2(g6313), .QN(n11397) );
  NAND2X0 U11118 ( .IN1(n11399), .IN2(n11400), .QN(g30262) );
  NAND2X0 U11119 ( .IN1(n4369), .IN2(test_so14), .QN(n11400) );
  NAND2X0 U11120 ( .IN1(n11401), .IN2(g165), .QN(n11399) );
  NAND2X0 U11121 ( .IN1(n11402), .IN2(n11403), .QN(g30261) );
  INVX0 U11122 ( .INP(n11404), .ZN(n11403) );
  NOR2X0 U11123 ( .IN1(g6231), .IN2(n8482), .QN(n11404) );
  NAND2X0 U11124 ( .IN1(n11337), .IN2(g6231), .QN(n11402) );
  NAND2X0 U11125 ( .IN1(n11405), .IN2(n11406), .QN(n11337) );
  NAND2X0 U11126 ( .IN1(n11097), .IN2(n11407), .QN(n11406) );
  XNOR2X1 U11127 ( .IN1(n11408), .IN2(n4513), .Q(n11407) );
  NAND2X0 U11128 ( .IN1(n10927), .IN2(g97), .QN(n11405) );
  NAND2X0 U11129 ( .IN1(n11409), .IN2(n11410), .QN(g30260) );
  INVX0 U11130 ( .INP(n11411), .ZN(n11410) );
  NOR2X0 U11131 ( .IN1(g2241), .IN2(n8535), .QN(n11411) );
  NAND2X0 U11132 ( .IN1(n11412), .IN2(g2241), .QN(n11409) );
  NAND2X0 U11133 ( .IN1(n11413), .IN2(n11414), .QN(g30259) );
  INVX0 U11134 ( .INP(n11415), .ZN(n11414) );
  NOR2X0 U11135 ( .IN1(g6368), .IN2(n8461), .QN(n11415) );
  NAND2X0 U11136 ( .IN1(n11363), .IN2(g6368), .QN(n11413) );
  NAND2X0 U11137 ( .IN1(n11416), .IN2(n11417), .QN(n11363) );
  NAND2X0 U11138 ( .IN1(n11418), .IN2(n11072), .QN(n11417) );
  XNOR2X1 U11139 ( .IN1(n11419), .IN2(n11420), .Q(n11418) );
  NAND2X0 U11140 ( .IN1(n11421), .IN2(n11422), .QN(n11419) );
  NAND2X0 U11141 ( .IN1(n11040), .IN2(n9775), .QN(n11422) );
  NAND2X0 U11142 ( .IN1(n10875), .IN2(g805), .QN(n11416) );
  NAND2X0 U11143 ( .IN1(n11423), .IN2(n11424), .QN(g30258) );
  INVX0 U11144 ( .INP(n11425), .ZN(n11424) );
  NOR2X0 U11145 ( .IN1(g6231), .IN2(n8471), .QN(n11425) );
  NAND2X0 U11146 ( .IN1(n11374), .IN2(g6231), .QN(n11423) );
  NAND2X0 U11147 ( .IN1(n11426), .IN2(n11427), .QN(n11374) );
  NAND2X0 U11148 ( .IN1(n11428), .IN2(n11097), .QN(n11427) );
  XOR2X1 U11149 ( .IN1(n9740), .IN2(n11095), .Q(n11428) );
  NOR2X0 U11150 ( .IN1(n11429), .IN2(n11430), .QN(n11095) );
  XNOR2X1 U11151 ( .IN1(n9738), .IN2(n10501), .Q(n11430) );
  NAND2X0 U11152 ( .IN1(n10927), .IN2(g125), .QN(n11426) );
  NAND2X0 U11153 ( .IN1(n11431), .IN2(n11432), .QN(g30257) );
  NAND2X0 U11154 ( .IN1(n4512), .IN2(g252), .QN(n11432) );
  NAND2X0 U11155 ( .IN1(n11401), .IN2(g6313), .QN(n11431) );
  NAND2X0 U11156 ( .IN1(n11433), .IN2(n11434), .QN(g30256) );
  NAND2X0 U11157 ( .IN1(g2291), .IN2(n9278), .QN(n11434) );
  NAND2X0 U11158 ( .IN1(test_so73), .IN2(n11412), .QN(n11433) );
  NAND2X0 U11159 ( .IN1(n11435), .IN2(n11436), .QN(g30255) );
  INVX0 U11160 ( .INP(n11437), .ZN(n11436) );
  NOR2X0 U11161 ( .IN1(g1547), .IN2(n8538), .QN(n11437) );
  NAND2X0 U11162 ( .IN1(n11438), .IN2(g1547), .QN(n11435) );
  NAND2X0 U11163 ( .IN1(n11439), .IN2(n11440), .QN(g30254) );
  INVX0 U11164 ( .INP(n11441), .ZN(n11440) );
  NOR2X0 U11165 ( .IN1(g6231), .IN2(n8475), .QN(n11441) );
  NAND2X0 U11166 ( .IN1(n11401), .IN2(g6231), .QN(n11439) );
  NAND2X0 U11167 ( .IN1(n11442), .IN2(n11443), .QN(n11401) );
  NAND2X0 U11168 ( .IN1(n11444), .IN2(n11097), .QN(n11443) );
  XNOR2X1 U11169 ( .IN1(n11445), .IN2(n9760), .Q(n11444) );
  NAND2X0 U11170 ( .IN1(n11446), .IN2(n11447), .QN(n11445) );
  NAND2X0 U11171 ( .IN1(n11083), .IN2(n9747), .QN(n11447) );
  NAND2X0 U11172 ( .IN1(n10927), .IN2(g117), .QN(n11442) );
  NAND2X0 U11173 ( .IN1(n11448), .IN2(n11449), .QN(g30253) );
  INVX0 U11174 ( .INP(n11450), .ZN(n11449) );
  NOR2X0 U11175 ( .IN1(g6837), .IN2(n8433), .QN(n11450) );
  NAND2X0 U11176 ( .IN1(n11412), .IN2(g6837), .QN(n11448) );
  NAND2X0 U11177 ( .IN1(n11451), .IN2(n11452), .QN(n11412) );
  NAND2X0 U11178 ( .IN1(n11453), .IN2(n11228), .QN(n11452) );
  XNOR2X1 U11179 ( .IN1(n11302), .IN2(n11304), .Q(n11453) );
  NAND2X0 U11180 ( .IN1(n11454), .IN2(n11345), .QN(n11302) );
  NOR2X0 U11181 ( .IN1(n11229), .IN2(n11455), .QN(n11345) );
  NOR2X0 U11182 ( .IN1(n10503), .IN2(n9852), .QN(n11455) );
  NAND2X0 U11183 ( .IN1(n10905), .IN2(n11456), .QN(n11229) );
  XNOR2X1 U11184 ( .IN1(n9864), .IN2(n4529), .Q(n11456) );
  NOR2X0 U11185 ( .IN1(n10779), .IN2(n11457), .QN(n10905) );
  XNOR2X1 U11186 ( .IN1(n11458), .IN2(n10503), .Q(n11457) );
  NAND2X0 U11187 ( .IN1(n10941), .IN2(n11459), .QN(n10779) );
  XNOR2X1 U11188 ( .IN1(n9858), .IN2(n10503), .Q(n11459) );
  NOR2X0 U11189 ( .IN1(n11460), .IN2(n11276), .QN(n10941) );
  XNOR2X1 U11190 ( .IN1(n9845), .IN2(n10503), .Q(n11460) );
  NOR2X0 U11191 ( .IN1(n11461), .IN2(n11462), .QN(n11454) );
  NOR2X0 U11192 ( .IN1(n11463), .IN2(n4529), .QN(n11462) );
  NOR2X0 U11193 ( .IN1(n11464), .IN2(n9865), .QN(n11461) );
  NAND2X0 U11194 ( .IN1(n10795), .IN2(g2195), .QN(n11451) );
  NOR2X0 U11195 ( .IN1(n10943), .IN2(n11228), .QN(n10795) );
  NOR2X0 U11196 ( .IN1(n11465), .IN2(n11466), .QN(n11228) );
  NOR2X0 U11197 ( .IN1(n11467), .IN2(n11276), .QN(n11466) );
  NOR2X0 U11198 ( .IN1(n11468), .IN2(n11469), .QN(n11467) );
  NOR2X0 U11199 ( .IN1(n9833), .IN2(n4529), .QN(n11469) );
  INVX0 U11200 ( .INP(n11470), .ZN(n11468) );
  NOR2X0 U11201 ( .IN1(n11471), .IN2(n11465), .QN(n10943) );
  NAND2X0 U11202 ( .IN1(n11472), .IN2(n11473), .QN(n11465) );
  NAND2X0 U11203 ( .IN1(n11188), .IN2(n11133), .QN(n11473) );
  NOR2X0 U11204 ( .IN1(n11101), .IN2(n11474), .QN(n11472) );
  NOR2X0 U11205 ( .IN1(n2792), .IN2(n11475), .QN(n11474) );
  NOR2X0 U11206 ( .IN1(n11476), .IN2(n11477), .QN(n11475) );
  NOR2X0 U11207 ( .IN1(n11187), .IN2(n11478), .QN(n11476) );
  NAND2X0 U11208 ( .IN1(n11102), .IN2(n11133), .QN(n11478) );
  NAND2X0 U11209 ( .IN1(n11479), .IN2(n11480), .QN(n2792) );
  NAND2X0 U11210 ( .IN1(n11481), .IN2(n11482), .QN(n11480) );
  NAND2X0 U11211 ( .IN1(n8547), .IN2(n10669), .QN(n11482) );
  NOR2X0 U11212 ( .IN1(n11483), .IN2(n11484), .QN(n11481) );
  NOR2X0 U11213 ( .IN1(n4516), .IN2(g2397), .QN(n11484) );
  NOR2X0 U11214 ( .IN1(n4509), .IN2(g2396), .QN(n11483) );
  NAND2X0 U11215 ( .IN1(n11485), .IN2(n11486), .QN(n11471) );
  NAND2X0 U11216 ( .IN1(n9833), .IN2(n11470), .QN(n11486) );
  NAND2X0 U11217 ( .IN1(n11487), .IN2(n11488), .QN(n11470) );
  NOR2X0 U11218 ( .IN1(n11489), .IN2(n11490), .QN(n11488) );
  NAND2X0 U11219 ( .IN1(n10800), .IN2(n11491), .QN(n11490) );
  NAND2X0 U11220 ( .IN1(n11492), .IN2(n11458), .QN(n11489) );
  NOR2X0 U11221 ( .IN1(n10975), .IN2(n11493), .QN(n11487) );
  NAND2X0 U11222 ( .IN1(n11494), .IN2(n9864), .QN(n11493) );
  INVX0 U11223 ( .INP(n11495), .ZN(n11494) );
  INVX0 U11224 ( .INP(n4529), .ZN(n10975) );
  NAND2X0 U11225 ( .IN1(n11496), .IN2(n11497), .QN(n9833) );
  NOR2X0 U11226 ( .IN1(n9864), .IN2(n11498), .QN(n11497) );
  NAND2X0 U11227 ( .IN1(n9863), .IN2(n9858), .QN(n11498) );
  NOR2X0 U11228 ( .IN1(n11495), .IN2(n11499), .QN(n11496) );
  NAND2X0 U11229 ( .IN1(n9851), .IN2(n9850), .QN(n11499) );
  NAND2X0 U11230 ( .IN1(n11500), .IN2(n11501), .QN(n11495) );
  NOR2X0 U11231 ( .IN1(n9844), .IN2(n11502), .QN(n11501) );
  NAND2X0 U11232 ( .IN1(n9843), .IN2(n11463), .QN(n11502) );
  NOR2X0 U11233 ( .IN1(n9845), .IN2(n9852), .QN(n11500) );
  INVX0 U11234 ( .INP(n11276), .ZN(n11485) );
  NOR2X0 U11235 ( .IN1(n4529), .IN2(n11503), .QN(n11276) );
  NAND2X0 U11236 ( .IN1(n11504), .IN2(n11505), .QN(g30252) );
  NAND2X0 U11237 ( .IN1(n4515), .IN2(g1597), .QN(n11505) );
  NAND2X0 U11238 ( .IN1(n11438), .IN2(g6782), .QN(n11504) );
  NAND2X0 U11239 ( .IN1(n11506), .IN2(n11507), .QN(g30251) );
  NAND2X0 U11240 ( .IN1(g906), .IN2(n9279), .QN(n11507) );
  NAND2X0 U11241 ( .IN1(test_so31), .IN2(n11508), .QN(n11506) );
  NAND2X0 U11242 ( .IN1(n11509), .IN2(n11510), .QN(g30250) );
  INVX0 U11243 ( .INP(n11511), .ZN(n11510) );
  NOR2X0 U11244 ( .IN1(g6573), .IN2(n8445), .QN(n11511) );
  NAND2X0 U11245 ( .IN1(n11438), .IN2(g6573), .QN(n11509) );
  NAND2X0 U11246 ( .IN1(n11512), .IN2(n11513), .QN(n11438) );
  NAND2X0 U11247 ( .IN1(n11514), .IN2(n11251), .QN(n11513) );
  XNOR2X1 U11248 ( .IN1(n11354), .IN2(n11515), .Q(n11514) );
  NAND2X0 U11249 ( .IN1(n11516), .IN2(n11385), .QN(n11354) );
  NOR2X0 U11250 ( .IN1(n11252), .IN2(n11517), .QN(n11385) );
  NOR2X0 U11251 ( .IN1(n10992), .IN2(n9817), .QN(n11517) );
  NAND2X0 U11252 ( .IN1(n10954), .IN2(n11518), .QN(n11252) );
  XNOR2X1 U11253 ( .IN1(n9823), .IN2(n4530), .Q(n11518) );
  NOR2X0 U11254 ( .IN1(n10813), .IN2(n11519), .QN(n10954) );
  XNOR2X1 U11255 ( .IN1(n9815), .IN2(n4530), .Q(n11519) );
  NAND2X0 U11256 ( .IN1(n10990), .IN2(n11520), .QN(n10813) );
  XNOR2X1 U11257 ( .IN1(n11521), .IN2(n4530), .Q(n11520) );
  NOR2X0 U11258 ( .IN1(n11522), .IN2(n11523), .QN(n10990) );
  XNOR2X1 U11259 ( .IN1(n11320), .IN2(n4530), .Q(n11522) );
  NOR2X0 U11260 ( .IN1(n11524), .IN2(n11525), .QN(n11516) );
  NOR2X0 U11261 ( .IN1(n9829), .IN2(n4530), .QN(n11525) );
  NOR2X0 U11262 ( .IN1(n11526), .IN2(n11384), .QN(n11524) );
  NAND2X0 U11263 ( .IN1(n10834), .IN2(g1501), .QN(n11512) );
  NOR2X0 U11264 ( .IN1(n10993), .IN2(n11251), .QN(n10834) );
  NOR2X0 U11265 ( .IN1(n11527), .IN2(n11528), .QN(n11251) );
  NOR2X0 U11266 ( .IN1(n11529), .IN2(n11523), .QN(n11528) );
  NOR2X0 U11267 ( .IN1(n11530), .IN2(n11531), .QN(n11529) );
  NOR2X0 U11268 ( .IN1(n9798), .IN2(n4530), .QN(n11531) );
  INVX0 U11269 ( .INP(n11532), .ZN(n11530) );
  NOR2X0 U11270 ( .IN1(n11533), .IN2(n11527), .QN(n10993) );
  NAND2X0 U11271 ( .IN1(n11534), .IN2(n11535), .QN(n11527) );
  NAND2X0 U11272 ( .IN1(n11536), .IN2(n10456), .QN(n11535) );
  NOR2X0 U11273 ( .IN1(n10685), .IN2(n11537), .QN(n11534) );
  NOR2X0 U11274 ( .IN1(n10690), .IN2(n11538), .QN(n11537) );
  NOR2X0 U11275 ( .IN1(n11539), .IN2(n10694), .QN(n11538) );
  NOR2X0 U11276 ( .IN1(n11540), .IN2(n10698), .QN(n11539) );
  INVX0 U11277 ( .INP(n11541), .ZN(n10698) );
  NOR2X0 U11278 ( .IN1(n11542), .IN2(n11543), .QN(n11541) );
  NAND2X0 U11279 ( .IN1(n11536), .IN2(n10686), .QN(n11542) );
  NAND2X0 U11280 ( .IN1(n11544), .IN2(n11545), .QN(n11536) );
  NAND2X0 U11281 ( .IN1(n8548), .IN2(n10678), .QN(n11545) );
  NOR2X0 U11282 ( .IN1(n11546), .IN2(n11547), .QN(n11544) );
  NOR2X0 U11283 ( .IN1(n4518), .IN2(g1703), .QN(n11547) );
  NOR2X0 U11284 ( .IN1(n4511), .IN2(g1702), .QN(n11546) );
  NAND2X0 U11285 ( .IN1(n11319), .IN2(n11548), .QN(n11533) );
  NAND2X0 U11286 ( .IN1(n9798), .IN2(n11532), .QN(n11548) );
  NAND2X0 U11287 ( .IN1(n11549), .IN2(n11550), .QN(n11532) );
  NOR2X0 U11288 ( .IN1(n11551), .IN2(n11552), .QN(n11550) );
  NAND2X0 U11289 ( .IN1(n9830), .IN2(n11521), .QN(n11552) );
  NAND2X0 U11290 ( .IN1(n10502), .IN2(n11553), .QN(n11551) );
  NOR2X0 U11291 ( .IN1(n11022), .IN2(n11554), .QN(n11549) );
  NAND2X0 U11292 ( .IN1(n11555), .IN2(n9823), .QN(n11554) );
  INVX0 U11293 ( .INP(n11556), .ZN(n11555) );
  INVX0 U11294 ( .INP(n4530), .ZN(n11022) );
  NAND2X0 U11295 ( .IN1(n11557), .IN2(n11558), .QN(n9798) );
  NOR2X0 U11296 ( .IN1(n9830), .IN2(n11559), .QN(n11558) );
  NAND2X0 U11297 ( .IN1(n9828), .IN2(n10953), .QN(n11559) );
  INVX0 U11298 ( .INP(n9823), .ZN(n10953) );
  NOR2X0 U11299 ( .IN1(n11556), .IN2(n11560), .QN(n11557) );
  NAND2X0 U11300 ( .IN1(n9816), .IN2(n9815), .QN(n11560) );
  NAND2X0 U11301 ( .IN1(n11561), .IN2(n11562), .QN(n11556) );
  NOR2X0 U11302 ( .IN1(n11029), .IN2(n11563), .QN(n11562) );
  NAND2X0 U11303 ( .IN1(n9808), .IN2(n9829), .QN(n11563) );
  NOR2X0 U11304 ( .IN1(n9810), .IN2(n9817), .QN(n11561) );
  INVX0 U11305 ( .INP(n11523), .ZN(n11319) );
  NOR2X0 U11306 ( .IN1(n4530), .IN2(n11564), .QN(n11523) );
  NAND2X0 U11307 ( .IN1(n11565), .IN2(n11566), .QN(g30249) );
  INVX0 U11308 ( .INP(n11567), .ZN(n11566) );
  NOR2X0 U11309 ( .IN1(g6518), .IN2(n8458), .QN(n11567) );
  NAND2X0 U11310 ( .IN1(n11508), .IN2(g6518), .QN(n11565) );
  NAND2X0 U11311 ( .IN1(n11568), .IN2(n11569), .QN(g30248) );
  INVX0 U11312 ( .INP(n11570), .ZN(n11569) );
  NOR2X0 U11313 ( .IN1(g165), .IN2(n8544), .QN(n11570) );
  NAND2X0 U11314 ( .IN1(n11571), .IN2(g165), .QN(n11568) );
  NAND2X0 U11315 ( .IN1(n11572), .IN2(n11573), .QN(g30247) );
  INVX0 U11316 ( .INP(n11574), .ZN(n11573) );
  NOR2X0 U11317 ( .IN1(g6368), .IN2(n8459), .QN(n11574) );
  NAND2X0 U11318 ( .IN1(n11508), .IN2(g6368), .QN(n11572) );
  NAND2X0 U11319 ( .IN1(n11575), .IN2(n11576), .QN(n11508) );
  NAND2X0 U11320 ( .IN1(n11577), .IN2(n11072), .QN(n11576) );
  XNOR2X1 U11321 ( .IN1(n11392), .IN2(n11578), .Q(n11577) );
  NAND2X0 U11322 ( .IN1(n11579), .IN2(n11421), .QN(n11392) );
  NOR2X0 U11323 ( .IN1(n11289), .IN2(n11580), .QN(n11421) );
  NOR2X0 U11324 ( .IN1(n11040), .IN2(n9775), .QN(n11580) );
  NAND2X0 U11325 ( .IN1(n11005), .IN2(n11581), .QN(n11289) );
  XNOR2X1 U11326 ( .IN1(n9782), .IN2(n10883), .Q(n11581) );
  NOR2X0 U11327 ( .IN1(n10852), .IN2(n11582), .QN(n11005) );
  XNOR2X1 U11328 ( .IN1(n9794), .IN2(n10883), .Q(n11582) );
  NAND2X0 U11329 ( .IN1(n11038), .IN2(n11583), .QN(n10852) );
  XNOR2X1 U11330 ( .IN1(n11584), .IN2(n10883), .Q(n11583) );
  NOR2X0 U11331 ( .IN1(n11585), .IN2(n11370), .QN(n11038) );
  XNOR2X1 U11332 ( .IN1(n9780), .IN2(n11040), .Q(n11585) );
  NOR2X0 U11333 ( .IN1(n11586), .IN2(n11587), .QN(n11579) );
  NOR2X0 U11334 ( .IN1(n9774), .IN2(n10883), .QN(n11587) );
  NOR2X0 U11335 ( .IN1(n11588), .IN2(n11420), .QN(n11586) );
  NAND2X0 U11336 ( .IN1(n10875), .IN2(g809), .QN(n11575) );
  NOR2X0 U11337 ( .IN1(n11041), .IN2(n11072), .QN(n10875) );
  NOR2X0 U11338 ( .IN1(n11589), .IN2(n11590), .QN(n11072) );
  NOR2X0 U11339 ( .IN1(n11591), .IN2(n11370), .QN(n11590) );
  NOR2X0 U11340 ( .IN1(n11592), .IN2(n11593), .QN(n11591) );
  NOR2X0 U11341 ( .IN1(n9763), .IN2(n10883), .QN(n11593) );
  INVX0 U11342 ( .INP(n11594), .ZN(n11592) );
  NOR2X0 U11343 ( .IN1(n11595), .IN2(n11589), .QN(n11041) );
  NAND2X0 U11344 ( .IN1(n11596), .IN2(n11597), .QN(n11589) );
  NAND2X0 U11345 ( .IN1(n10516), .IN2(n10489), .QN(n11597) );
  NOR2X0 U11346 ( .IN1(n158), .IN2(n11598), .QN(n11596) );
  NOR2X0 U11347 ( .IN1(n2632), .IN2(n11599), .QN(n11598) );
  NOR2X0 U11348 ( .IN1(n11600), .IN2(n11601), .QN(n11599) );
  NOR2X0 U11349 ( .IN1(n10492), .IN2(n11602), .QN(n11600) );
  NAND2X0 U11350 ( .IN1(n10489), .IN2(n10494), .QN(n11602) );
  NAND2X0 U11351 ( .IN1(n11603), .IN2(n11604), .QN(n2632) );
  NAND2X0 U11352 ( .IN1(n11605), .IN2(n11606), .QN(n11604) );
  NAND2X0 U11353 ( .IN1(n8554), .IN2(g1088), .QN(n11606) );
  NOR2X0 U11354 ( .IN1(n11607), .IN2(n11608), .QN(n11605) );
  NOR2X0 U11355 ( .IN1(n4364), .IN2(g1010), .QN(n11608) );
  NOR2X0 U11356 ( .IN1(n4363), .IN2(g1009), .QN(n11607) );
  NAND2X0 U11357 ( .IN1(n11609), .IN2(n11610), .QN(n11595) );
  NAND2X0 U11358 ( .IN1(n9763), .IN2(n11594), .QN(n11610) );
  NAND2X0 U11359 ( .IN1(n11611), .IN2(n11612), .QN(n11594) );
  NOR2X0 U11360 ( .IN1(n11613), .IN2(n11614), .QN(n11612) );
  NAND2X0 U11361 ( .IN1(n9795), .IN2(n9793), .QN(n11614) );
  NAND2X0 U11362 ( .IN1(n11584), .IN2(n9782), .QN(n11613) );
  NOR2X0 U11363 ( .IN1(n11040), .IN2(n11615), .QN(n11611) );
  NAND2X0 U11364 ( .IN1(n11616), .IN2(n11617), .QN(n11615) );
  INVX0 U11365 ( .INP(n11618), .ZN(n11616) );
  NAND2X0 U11366 ( .IN1(n11619), .IN2(n11620), .QN(n9763) );
  NOR2X0 U11367 ( .IN1(n9795), .IN2(n11621), .QN(n11620) );
  INVX0 U11368 ( .INP(n11622), .ZN(n11621) );
  NOR2X0 U11369 ( .IN1(n11617), .IN2(n9793), .QN(n11622) );
  NOR2X0 U11370 ( .IN1(n11618), .IN2(n11623), .QN(n11619) );
  NAND2X0 U11371 ( .IN1(n11004), .IN2(n9781), .QN(n11623) );
  NAND2X0 U11372 ( .IN1(n11624), .IN2(n11625), .QN(n11618) );
  NOR2X0 U11373 ( .IN1(n11420), .IN2(n11626), .QN(n11625) );
  NAND2X0 U11374 ( .IN1(n9773), .IN2(n9788), .QN(n11626) );
  NOR2X0 U11375 ( .IN1(n9775), .IN2(n9780), .QN(n11624) );
  INVX0 U11376 ( .INP(n11370), .ZN(n11609) );
  NOR2X0 U11377 ( .IN1(n10883), .IN2(n11627), .QN(n11370) );
  NAND2X0 U11378 ( .IN1(n11628), .IN2(n11629), .QN(g30246) );
  NAND2X0 U11379 ( .IN1(n4512), .IN2(g216), .QN(n11629) );
  NAND2X0 U11380 ( .IN1(n11571), .IN2(g6313), .QN(n11628) );
  NAND2X0 U11381 ( .IN1(n11630), .IN2(n11631), .QN(g30245) );
  INVX0 U11382 ( .INP(n11632), .ZN(n11631) );
  NOR2X0 U11383 ( .IN1(g6231), .IN2(n8473), .QN(n11632) );
  NAND2X0 U11384 ( .IN1(n11571), .IN2(g6231), .QN(n11630) );
  NAND2X0 U11385 ( .IN1(n11633), .IN2(n11634), .QN(n11571) );
  NAND2X0 U11386 ( .IN1(n11635), .IN2(n11097), .QN(n11634) );
  XNOR2X1 U11387 ( .IN1(n11429), .IN2(n11636), .Q(n11635) );
  NAND2X0 U11388 ( .IN1(n11637), .IN2(n11446), .QN(n11429) );
  NOR2X0 U11389 ( .IN1(n11333), .IN2(n11638), .QN(n11446) );
  NOR2X0 U11390 ( .IN1(n11083), .IN2(n9747), .QN(n11638) );
  NAND2X0 U11391 ( .IN1(n11053), .IN2(n11639), .QN(n11333) );
  XNOR2X1 U11392 ( .IN1(n11640), .IN2(n10501), .Q(n11639) );
  NOR2X0 U11393 ( .IN1(n10896), .IN2(n11641), .QN(n11053) );
  XNOR2X1 U11394 ( .IN1(n9745), .IN2(n10501), .Q(n11641) );
  NAND2X0 U11395 ( .IN1(n11081), .IN2(n11642), .QN(n10896) );
  XNOR2X1 U11396 ( .IN1(n11643), .IN2(n10501), .Q(n11642) );
  NOR2X0 U11397 ( .IN1(n11644), .IN2(n11645), .QN(n11081) );
  XNOR2X1 U11398 ( .IN1(n4513), .IN2(n10501), .Q(n11644) );
  INVX0 U11399 ( .INP(n11646), .ZN(n4513) );
  NAND2X0 U11400 ( .IN1(n11647), .IN2(n11648), .QN(n11646) );
  NAND2X0 U11401 ( .IN1(test_so13), .IN2(g6313), .QN(n11648) );
  NOR2X0 U11402 ( .IN1(n11649), .IN2(n11650), .QN(n11647) );
  NOR2X0 U11403 ( .IN1(n8546), .IN2(n4369), .QN(n11650) );
  NOR2X0 U11404 ( .IN1(n8482), .IN2(n4318), .QN(n11649) );
  NOR2X0 U11405 ( .IN1(n11651), .IN2(n11652), .QN(n11637) );
  NOR2X0 U11406 ( .IN1(n11653), .IN2(n10501), .QN(n11652) );
  NOR2X0 U11407 ( .IN1(n11654), .IN2(n9760), .QN(n11651) );
  NAND2X0 U11408 ( .IN1(n10927), .IN2(g121), .QN(n11633) );
  NOR2X0 U11409 ( .IN1(n11084), .IN2(n11097), .QN(n10927) );
  NOR2X0 U11410 ( .IN1(n11655), .IN2(n11656), .QN(n11097) );
  NOR2X0 U11411 ( .IN1(n11657), .IN2(n11645), .QN(n11656) );
  NOR2X0 U11412 ( .IN1(n11658), .IN2(n11659), .QN(n11657) );
  NOR2X0 U11413 ( .IN1(n9728), .IN2(n10501), .QN(n11659) );
  INVX0 U11414 ( .INP(n11660), .ZN(n11658) );
  NOR2X0 U11415 ( .IN1(n11661), .IN2(n11655), .QN(n11084) );
  NAND2X0 U11416 ( .IN1(n11662), .IN2(n11663), .QN(n11655) );
  NAND2X0 U11417 ( .IN1(n11664), .IN2(n10455), .QN(n11663) );
  NOR2X0 U11418 ( .IN1(n10724), .IN2(n11665), .QN(n11662) );
  NOR2X0 U11419 ( .IN1(n10729), .IN2(n11666), .QN(n11665) );
  NOR2X0 U11420 ( .IN1(n11667), .IN2(n10733), .QN(n11666) );
  NOR2X0 U11421 ( .IN1(n11668), .IN2(n10737), .QN(n11667) );
  INVX0 U11422 ( .INP(n11669), .ZN(n10737) );
  NOR2X0 U11423 ( .IN1(n11670), .IN2(n11671), .QN(n11669) );
  NAND2X0 U11424 ( .IN1(n11664), .IN2(n10725), .QN(n11670) );
  NAND2X0 U11425 ( .IN1(n11672), .IN2(n11673), .QN(n11664) );
  NAND2X0 U11426 ( .IN1(n8558), .IN2(n10752), .QN(n11673) );
  NOR2X0 U11427 ( .IN1(n11674), .IN2(n11675), .QN(n11672) );
  NOR2X0 U11428 ( .IN1(n4506), .IN2(g321), .QN(n11675) );
  NOR2X0 U11429 ( .IN1(n4499), .IN2(g323), .QN(n11674) );
  NAND2X0 U11430 ( .IN1(n11408), .IN2(n11676), .QN(n11661) );
  NAND2X0 U11431 ( .IN1(n9728), .IN2(n11660), .QN(n11676) );
  NAND2X0 U11432 ( .IN1(n11677), .IN2(n11678), .QN(n11660) );
  NOR2X0 U11433 ( .IN1(n11679), .IN2(n11680), .QN(n11678) );
  NAND2X0 U11434 ( .IN1(n10932), .IN2(n11643), .QN(n11680) );
  NAND2X0 U11435 ( .IN1(n10500), .IN2(n11681), .QN(n11679) );
  INVX0 U11436 ( .INP(n11682), .ZN(n11677) );
  NAND2X0 U11437 ( .IN1(n10501), .IN2(n11683), .QN(n11682) );
  NOR2X0 U11438 ( .IN1(n11684), .IN2(n9754), .QN(n11683) );
  NAND2X0 U11439 ( .IN1(n11685), .IN2(n11686), .QN(n9728) );
  NOR2X0 U11440 ( .IN1(n11643), .IN2(n11687), .QN(n11686) );
  NAND2X0 U11441 ( .IN1(n9759), .IN2(n9754), .QN(n11687) );
  NOR2X0 U11442 ( .IN1(n11684), .IN2(n11688), .QN(n11685) );
  NAND2X0 U11443 ( .IN1(n9746), .IN2(n9745), .QN(n11688) );
  NAND2X0 U11444 ( .IN1(n11689), .IN2(n11690), .QN(n11684) );
  NOR2X0 U11445 ( .IN1(n9740), .IN2(n11691), .QN(n11690) );
  NAND2X0 U11446 ( .IN1(n9738), .IN2(n11653), .QN(n11691) );
  INVX0 U11447 ( .INP(n11636), .ZN(n9738) );
  NOR2X0 U11448 ( .IN1(n9747), .IN2(n11692), .QN(n11689) );
  INVX0 U11449 ( .INP(n11645), .ZN(n11408) );
  NOR2X0 U11450 ( .IN1(n10501), .IN2(n11693), .QN(n11645) );
  NAND2X0 U11451 ( .IN1(n11694), .IN2(n11695), .QN(g30072) );
  NAND2X0 U11452 ( .IN1(g2574), .IN2(n7930), .QN(n11695) );
  NAND2X0 U11453 ( .IN1(n4543), .IN2(n11696), .QN(n11694) );
  NAND2X0 U11454 ( .IN1(n11697), .IN2(n11698), .QN(n11696) );
  NAND2X0 U11455 ( .IN1(n532), .IN2(n11699), .QN(n11698) );
  NAND2X0 U11456 ( .IN1(n11700), .IN2(n7929), .QN(n11697) );
  NAND2X0 U11457 ( .IN1(n11701), .IN2(n11702), .QN(g30061) );
  NAND2X0 U11458 ( .IN1(g2580), .IN2(n7926), .QN(n11702) );
  NAND2X0 U11459 ( .IN1(n8755), .IN2(n11703), .QN(n11701) );
  NAND2X0 U11460 ( .IN1(n11704), .IN2(n11705), .QN(n11703) );
  NAND2X0 U11461 ( .IN1(n4370), .IN2(g16437), .QN(n11705) );
  NAND2X0 U11462 ( .IN1(n548), .IN2(g7390), .QN(n11704) );
  INVX0 U11463 ( .INP(n11706), .ZN(n548) );
  NAND2X0 U11464 ( .IN1(n11707), .IN2(n11708), .QN(n11706) );
  NAND2X0 U11465 ( .IN1(g1886), .IN2(DFF_1133_n1), .QN(n11708) );
  NAND2X0 U11466 ( .IN1(n4493), .IN2(n11709), .QN(n11707) );
  NAND2X0 U11467 ( .IN1(n11710), .IN2(n11711), .QN(n11709) );
  NAND2X0 U11468 ( .IN1(n4315), .IN2(DFF_1142_n1), .QN(n11711) );
  NAND2X0 U11469 ( .IN1(n9698), .IN2(g7194), .QN(n11710) );
  NAND2X0 U11470 ( .IN1(n11712), .IN2(n11713), .QN(n9698) );
  NAND2X0 U11471 ( .IN1(g1192), .IN2(DFF_783_n1), .QN(n11713) );
  NAND2X0 U11472 ( .IN1(n4454), .IN2(n11714), .QN(n11712) );
  NAND2X0 U11473 ( .IN1(n11715), .IN2(n11716), .QN(n11714) );
  NAND2X0 U11474 ( .IN1(n4316), .IN2(DFF_792_n1), .QN(n11716) );
  NAND2X0 U11475 ( .IN1(n9697), .IN2(g6944), .QN(n11715) );
  NAND2X0 U11476 ( .IN1(n11717), .IN2(n11718), .QN(n9697) );
  NAND2X0 U11477 ( .IN1(n8672), .IN2(g506), .QN(n11718) );
  NAND2X0 U11478 ( .IN1(n11719), .IN2(n4570), .QN(n11717) );
  NOR2X0 U11479 ( .IN1(g6642), .IN2(g16297), .QN(n11719) );
  NAND2X0 U11480 ( .IN1(n11720), .IN2(n11721), .QN(g30055) );
  NAND2X0 U11481 ( .IN1(n4487), .IN2(DFF_1378_n1), .QN(n11721) );
  NAND2X0 U11482 ( .IN1(n11722), .IN2(g2374), .QN(n11720) );
  NAND2X0 U11483 ( .IN1(n11723), .IN2(n11724), .QN(n11722) );
  NAND2X0 U11484 ( .IN1(n478), .IN2(g7264), .QN(n11724) );
  INVX0 U11485 ( .INP(n11725), .ZN(n478) );
  NAND2X0 U11486 ( .IN1(n11726), .IN2(n11727), .QN(n11725) );
  NAND2X0 U11487 ( .IN1(n4488), .IN2(n7978), .QN(n11727) );
  NAND2X0 U11488 ( .IN1(n11728), .IN2(g1680), .QN(n11726) );
  NOR2X0 U11489 ( .IN1(n11729), .IN2(n11730), .QN(n11728) );
  NOR2X0 U11490 ( .IN1(n8986), .IN2(n10678), .QN(n11730) );
  NOR2X0 U11491 ( .IN1(n9715), .IN2(n11731), .QN(n11729) );
  NAND2X0 U11492 ( .IN1(n11732), .IN2(n11733), .QN(n9715) );
  NAND2X0 U11493 ( .IN1(n4432), .IN2(n8017), .QN(n11733) );
  NAND2X0 U11494 ( .IN1(n11734), .IN2(g986), .QN(n11732) );
  NAND2X0 U11495 ( .IN1(n11735), .IN2(n11736), .QN(n11734) );
  NAND2X0 U11496 ( .IN1(n4364), .IN2(n8987), .QN(n11736) );
  INVX0 U11497 ( .INP(n11737), .ZN(n11735) );
  NOR2X0 U11498 ( .IN1(g21346), .IN2(n4364), .QN(n11737) );
  NAND2X0 U11499 ( .IN1(n4524), .IN2(g2380), .QN(n11723) );
  NAND2X0 U11500 ( .IN1(n11738), .IN2(n11739), .QN(g29941) );
  NAND2X0 U11501 ( .IN1(n4494), .IN2(g3105), .QN(n11739) );
  NAND2X0 U11502 ( .IN1(n532), .IN2(g3109), .QN(n11738) );
  NAND2X0 U11503 ( .IN1(n11740), .IN2(n11741), .QN(g29939) );
  INVX0 U11504 ( .INP(n11742), .ZN(n11741) );
  NOR2X0 U11505 ( .IN1(g8030), .IN2(n4452), .QN(n11742) );
  NAND2X0 U11506 ( .IN1(n532), .IN2(g8030), .QN(n11740) );
  NAND2X0 U11507 ( .IN1(n11743), .IN2(n11744), .QN(g29936) );
  INVX0 U11508 ( .INP(n11745), .ZN(n11744) );
  NOR2X0 U11509 ( .IN1(g8106), .IN2(n4447), .QN(n11745) );
  NAND2X0 U11510 ( .IN1(n532), .IN2(g8106), .QN(n11743) );
  INVX0 U11511 ( .INP(n11746), .ZN(n532) );
  NAND2X0 U11512 ( .IN1(n11747), .IN2(n11748), .QN(n11746) );
  NAND2X0 U11513 ( .IN1(g1880), .IN2(DFF_1099_n1), .QN(n11748) );
  NAND2X0 U11514 ( .IN1(n11749), .IN2(n4545), .QN(n11747) );
  NOR2X0 U11515 ( .IN1(n11750), .IN2(n11751), .QN(n11749) );
  NOR2X0 U11516 ( .IN1(g7052), .IN2(DFF_1100_n1), .QN(n11751) );
  NOR2X0 U11517 ( .IN1(n4296), .IN2(n11752), .QN(n11750) );
  NAND2X0 U11518 ( .IN1(n11753), .IN2(n11754), .QN(g29623) );
  NAND2X0 U11519 ( .IN1(n11755), .IN2(n4606), .QN(n11754) );
  NAND2X0 U11520 ( .IN1(n4509), .IN2(g2389), .QN(n11753) );
  NAND2X0 U11521 ( .IN1(n11756), .IN2(n11757), .QN(g29621) );
  NAND2X0 U11522 ( .IN1(n11755), .IN2(g7264), .QN(n11757) );
  INVX0 U11523 ( .INP(n11758), .ZN(n11756) );
  NOR2X0 U11524 ( .IN1(n10669), .IN2(n8495), .QN(n11758) );
  NAND2X0 U11525 ( .IN1(n11759), .IN2(n11760), .QN(g29620) );
  NAND2X0 U11526 ( .IN1(n11761), .IN2(n4618), .QN(n11760) );
  NAND2X0 U11527 ( .IN1(n4511), .IN2(g1695), .QN(n11759) );
  NAND2X0 U11528 ( .IN1(n11762), .IN2(n11763), .QN(g29618) );
  NAND2X0 U11529 ( .IN1(n11755), .IN2(g5555), .QN(n11763) );
  NOR2X0 U11530 ( .IN1(n11764), .IN2(n11101), .QN(n11755) );
  INVX0 U11531 ( .INP(n11765), .ZN(n11101) );
  NAND2X0 U11532 ( .IN1(n11479), .IN2(n11766), .QN(n11765) );
  NOR2X0 U11533 ( .IN1(n4529), .IN2(n11767), .QN(n11764) );
  NOR2X0 U11534 ( .IN1(n11768), .IN2(n11477), .QN(n11767) );
  NAND2X0 U11535 ( .IN1(n11187), .IN2(n11133), .QN(n11768) );
  INVX0 U11536 ( .INP(n10503), .ZN(n4529) );
  NAND2X0 U11537 ( .IN1(n11769), .IN2(n11123), .QN(n10503) );
  NOR2X0 U11538 ( .IN1(n11102), .IN2(n11133), .QN(n11769) );
  NAND2X0 U11539 ( .IN1(n4516), .IN2(g2387), .QN(n11762) );
  NAND2X0 U11540 ( .IN1(n11770), .IN2(n11771), .QN(g29617) );
  NAND2X0 U11541 ( .IN1(n11761), .IN2(g7014), .QN(n11771) );
  INVX0 U11542 ( .INP(n11772), .ZN(n11770) );
  NOR2X0 U11543 ( .IN1(n10678), .IN2(n8498), .QN(n11772) );
  NAND2X0 U11544 ( .IN1(n11773), .IN2(n11774), .QN(g29616) );
  INVX0 U11545 ( .INP(n11775), .ZN(n11774) );
  NOR2X0 U11546 ( .IN1(g1088), .IN2(n8517), .QN(n11775) );
  NAND2X0 U11547 ( .IN1(n11776), .IN2(g1088), .QN(n11773) );
  NAND2X0 U11548 ( .IN1(n11777), .IN2(n11778), .QN(g29613) );
  NAND2X0 U11549 ( .IN1(n11761), .IN2(g5511), .QN(n11778) );
  NOR2X0 U11550 ( .IN1(n11779), .IN2(n10685), .QN(n11761) );
  NOR2X0 U11551 ( .IN1(n11543), .IN2(n11780), .QN(n10685) );
  INVX0 U11552 ( .INP(n11781), .ZN(n11780) );
  NOR2X0 U11553 ( .IN1(n4530), .IN2(n11782), .QN(n11779) );
  NOR2X0 U11554 ( .IN1(n11783), .IN2(n11206), .QN(n11782) );
  NAND2X0 U11555 ( .IN1(n10711), .IN2(n11784), .QN(n11783) );
  INVX0 U11556 ( .INP(n10992), .ZN(n4530) );
  NAND2X0 U11557 ( .IN1(n11785), .IN2(n11198), .QN(n10992) );
  NOR2X0 U11558 ( .IN1(n10686), .IN2(n10711), .QN(n11785) );
  NAND2X0 U11559 ( .IN1(n4518), .IN2(g1693), .QN(n11777) );
  NAND2X0 U11560 ( .IN1(n11786), .IN2(n11787), .QN(g29612) );
  NAND2X0 U11561 ( .IN1(n4364), .IN2(g1000), .QN(n11787) );
  NAND2X0 U11562 ( .IN1(n11776), .IN2(g6712), .QN(n11786) );
  NAND2X0 U11563 ( .IN1(n11788), .IN2(n11789), .QN(g29611) );
  NAND2X0 U11564 ( .IN1(n11790), .IN2(n4640), .QN(n11789) );
  NAND2X0 U11565 ( .IN1(n4506), .IN2(g314), .QN(n11788) );
  NAND2X0 U11566 ( .IN1(n11791), .IN2(n11792), .QN(g29609) );
  NAND2X0 U11567 ( .IN1(n4363), .IN2(g999), .QN(n11792) );
  NAND2X0 U11568 ( .IN1(n11776), .IN2(g5472), .QN(n11791) );
  NOR2X0 U11569 ( .IN1(n11793), .IN2(n158), .QN(n11776) );
  INVX0 U11570 ( .INP(n11794), .ZN(n158) );
  NAND2X0 U11571 ( .IN1(n11603), .IN2(n11795), .QN(n11794) );
  NOR2X0 U11572 ( .IN1(n10883), .IN2(n11796), .QN(n11793) );
  NOR2X0 U11573 ( .IN1(n11797), .IN2(n10494), .QN(n11796) );
  NAND2X0 U11574 ( .IN1(n10489), .IN2(n11798), .QN(n11797) );
  INVX0 U11575 ( .INP(n11040), .ZN(n10883) );
  NAND2X0 U11576 ( .IN1(n11799), .IN2(n10486), .QN(n11040) );
  NOR2X0 U11577 ( .IN1(n10495), .IN2(n10489), .QN(n11799) );
  NAND2X0 U11578 ( .IN1(n11800), .IN2(n11801), .QN(g29608) );
  NAND2X0 U11579 ( .IN1(n11790), .IN2(g6447), .QN(n11801) );
  NAND2X0 U11580 ( .IN1(n4499), .IN2(g313), .QN(n11800) );
  NAND2X0 U11581 ( .IN1(n11802), .IN2(n11803), .QN(g29606) );
  NAND2X0 U11582 ( .IN1(n11790), .IN2(g5437), .QN(n11803) );
  NOR2X0 U11583 ( .IN1(n11804), .IN2(n10724), .QN(n11790) );
  NOR2X0 U11584 ( .IN1(n11671), .IN2(n11805), .QN(n10724) );
  INVX0 U11585 ( .INP(n11806), .ZN(n11805) );
  NOR2X0 U11586 ( .IN1(n10501), .IN2(n11807), .QN(n11804) );
  NOR2X0 U11587 ( .IN1(n11808), .IN2(n11166), .QN(n11807) );
  NAND2X0 U11588 ( .IN1(n10750), .IN2(n11809), .QN(n11808) );
  INVX0 U11589 ( .INP(n11083), .ZN(n10501) );
  NAND2X0 U11590 ( .IN1(n11810), .IN2(n11158), .QN(n11083) );
  NOR2X0 U11591 ( .IN1(n10725), .IN2(n10750), .QN(n11810) );
  INVX0 U11592 ( .INP(n11811), .ZN(n11802) );
  NOR2X0 U11593 ( .IN1(n10752), .IN2(n8526), .QN(n11811) );
  NOR2X0 U11594 ( .IN1(n9702), .IN2(n11812), .QN(g29582) );
  XNOR2X1 U11595 ( .IN1(n8388), .IN2(n2981), .Q(n11812) );
  NOR2X0 U11596 ( .IN1(n9710), .IN2(n11813), .QN(g29581) );
  XNOR2X1 U11597 ( .IN1(n8389), .IN2(n2984), .Q(n11813) );
  NOR2X0 U11598 ( .IN1(n11814), .IN2(n11815), .QN(g29580) );
  XNOR2X1 U11599 ( .IN1(n8390), .IN2(n2987), .Q(n11815) );
  NOR2X0 U11600 ( .IN1(n9719), .IN2(n11816), .QN(g29579) );
  XNOR2X1 U11601 ( .IN1(n8391), .IN2(n2990), .Q(n11816) );
  NAND2X0 U11602 ( .IN1(n11817), .IN2(n11818), .QN(g29357) );
  INVX0 U11603 ( .INP(n11819), .ZN(n11818) );
  NOR2X0 U11604 ( .IN1(n11820), .IN2(n8559), .QN(n11819) );
  NAND2X0 U11605 ( .IN1(n11821), .IN2(n8559), .QN(n11817) );
  NOR2X0 U11606 ( .IN1(n9702), .IN2(n2982), .QN(n11821) );
  NAND2X0 U11607 ( .IN1(n11822), .IN2(n11823), .QN(g29355) );
  INVX0 U11608 ( .INP(n11824), .ZN(n11823) );
  NOR2X0 U11609 ( .IN1(n11825), .IN2(n8560), .QN(n11824) );
  NAND2X0 U11610 ( .IN1(n11826), .IN2(n8560), .QN(n11822) );
  NOR2X0 U11611 ( .IN1(n9710), .IN2(n2985), .QN(n11826) );
  NAND2X0 U11612 ( .IN1(n11827), .IN2(n11828), .QN(g29354) );
  INVX0 U11613 ( .INP(n11829), .ZN(n11828) );
  NOR2X0 U11614 ( .IN1(n11830), .IN2(n8561), .QN(n11829) );
  NAND2X0 U11615 ( .IN1(n11831), .IN2(n8561), .QN(n11827) );
  NOR2X0 U11616 ( .IN1(n11814), .IN2(n2988), .QN(n11831) );
  NAND2X0 U11617 ( .IN1(n11832), .IN2(n11833), .QN(g29353) );
  INVX0 U11618 ( .INP(n11834), .ZN(n11833) );
  NOR2X0 U11619 ( .IN1(n11835), .IN2(n8562), .QN(n11834) );
  NAND2X0 U11620 ( .IN1(n11836), .IN2(n8562), .QN(n11832) );
  NOR2X0 U11621 ( .IN1(n9719), .IN2(n2991), .QN(n11836) );
  NAND2X0 U11622 ( .IN1(n11837), .IN2(n11838), .QN(g29226) );
  NAND2X0 U11623 ( .IN1(n11839), .IN2(n4606), .QN(n11838) );
  INVX0 U11624 ( .INP(n11840), .ZN(n11837) );
  NOR2X0 U11625 ( .IN1(n11841), .IN2(n8715), .QN(n11840) );
  NAND2X0 U11626 ( .IN1(n11842), .IN2(n11843), .QN(g29221) );
  NAND2X0 U11627 ( .IN1(n11839), .IN2(g7264), .QN(n11843) );
  INVX0 U11628 ( .INP(n11844), .ZN(n11842) );
  NOR2X0 U11629 ( .IN1(n10669), .IN2(n8702), .QN(n11844) );
  NAND2X0 U11630 ( .IN1(n11845), .IN2(n11846), .QN(g29218) );
  NAND2X0 U11631 ( .IN1(n11847), .IN2(n4618), .QN(n11846) );
  INVX0 U11632 ( .INP(n11848), .ZN(n11845) );
  NOR2X0 U11633 ( .IN1(n11849), .IN2(n8721), .QN(n11848) );
  NAND2X0 U11634 ( .IN1(n11850), .IN2(n11851), .QN(g29213) );
  NAND2X0 U11635 ( .IN1(n11839), .IN2(g5555), .QN(n11851) );
  XNOR2X1 U11636 ( .IN1(n10478), .IN2(n11852), .Q(n11839) );
  NOR2X0 U11637 ( .IN1(n9281), .IN2(n11853), .QN(n11852) );
  NAND2X0 U11638 ( .IN1(n11854), .IN2(n11855), .QN(n11853) );
  NAND2X0 U11639 ( .IN1(n11856), .IN2(n4285), .QN(n11855) );
  NAND2X0 U11640 ( .IN1(n11857), .IN2(n11858), .QN(n11856) );
  NOR2X0 U11641 ( .IN1(n11859), .IN2(n11860), .QN(n11857) );
  NAND2X0 U11642 ( .IN1(n11861), .IN2(n10478), .QN(n11854) );
  NAND2X0 U11643 ( .IN1(n11859), .IN2(n11862), .QN(n11861) );
  NAND2X0 U11644 ( .IN1(n10479), .IN2(n11863), .QN(n11862) );
  NAND2X0 U11645 ( .IN1(n11858), .IN2(n10476), .QN(n11863) );
  INVX0 U11646 ( .INP(n11188), .ZN(n10479) );
  NAND2X0 U11647 ( .IN1(n4516), .IN2(g2492), .QN(n11850) );
  NAND2X0 U11648 ( .IN1(n11864), .IN2(n11865), .QN(g29212) );
  NAND2X0 U11649 ( .IN1(n11847), .IN2(g7014), .QN(n11865) );
  INVX0 U11650 ( .INP(n11866), .ZN(n11864) );
  NOR2X0 U11651 ( .IN1(n10678), .IN2(n8706), .QN(n11866) );
  NAND2X0 U11652 ( .IN1(n11867), .IN2(n11868), .QN(g29209) );
  NAND2X0 U11653 ( .IN1(n4381), .IN2(g1110), .QN(n11868) );
  NAND2X0 U11654 ( .IN1(n11869), .IN2(g1088), .QN(n11867) );
  NAND2X0 U11655 ( .IN1(n11870), .IN2(n11871), .QN(g29205) );
  NAND2X0 U11656 ( .IN1(n11847), .IN2(g5511), .QN(n11871) );
  XNOR2X1 U11657 ( .IN1(n11872), .IN2(n11873), .Q(n11847) );
  NOR2X0 U11658 ( .IN1(n11874), .IN2(n11875), .QN(n11873) );
  NAND2X0 U11659 ( .IN1(n11876), .IN2(g1690), .QN(n11875) );
  NAND2X0 U11660 ( .IN1(n11877), .IN2(n10471), .QN(n11876) );
  NAND2X0 U11661 ( .IN1(n10694), .IN2(n11872), .QN(n10471) );
  NAND2X0 U11662 ( .IN1(n11878), .IN2(n10472), .QN(n11877) );
  XNOR2X1 U11663 ( .IN1(n10473), .IN2(n11872), .Q(n11874) );
  NAND2X0 U11664 ( .IN1(n4518), .IN2(g1798), .QN(n11870) );
  NAND2X0 U11665 ( .IN1(n11879), .IN2(n11880), .QN(g29204) );
  INVX0 U11666 ( .INP(n11881), .ZN(n11880) );
  NOR2X0 U11667 ( .IN1(g6712), .IN2(n8709), .QN(n11881) );
  NAND2X0 U11668 ( .IN1(n11869), .IN2(g6712), .QN(n11879) );
  NAND2X0 U11669 ( .IN1(n11882), .IN2(n11883), .QN(g29201) );
  NAND2X0 U11670 ( .IN1(n11884), .IN2(n4640), .QN(n11883) );
  INVX0 U11671 ( .INP(n11885), .ZN(n11882) );
  NOR2X0 U11672 ( .IN1(n11886), .IN2(n8739), .QN(n11885) );
  NAND2X0 U11673 ( .IN1(n11887), .IN2(n11888), .QN(g29198) );
  INVX0 U11674 ( .INP(n11889), .ZN(n11888) );
  NOR2X0 U11675 ( .IN1(g5472), .IN2(n8730), .QN(n11889) );
  NAND2X0 U11676 ( .IN1(n11869), .IN2(g5472), .QN(n11887) );
  XNOR2X1 U11677 ( .IN1(n10466), .IN2(n11890), .Q(n11869) );
  NOR2X0 U11678 ( .IN1(n4387), .IN2(n11891), .QN(n11890) );
  NAND2X0 U11679 ( .IN1(n11892), .IN2(n11893), .QN(n11891) );
  NAND2X0 U11680 ( .IN1(n11894), .IN2(n4283), .QN(n11893) );
  NAND2X0 U11681 ( .IN1(n11895), .IN2(n11896), .QN(n11894) );
  NOR2X0 U11682 ( .IN1(n11897), .IN2(n11898), .QN(n11895) );
  NAND2X0 U11683 ( .IN1(n11899), .IN2(n10466), .QN(n11892) );
  NAND2X0 U11684 ( .IN1(n11897), .IN2(n11900), .QN(n11899) );
  NAND2X0 U11685 ( .IN1(n10467), .IN2(n11901), .QN(n11900) );
  NAND2X0 U11686 ( .IN1(n11896), .IN2(n10464), .QN(n11901) );
  INVX0 U11687 ( .INP(n10516), .ZN(n10467) );
  NAND2X0 U11688 ( .IN1(n11902), .IN2(n11903), .QN(g29197) );
  NAND2X0 U11689 ( .IN1(n11884), .IN2(g6447), .QN(n11903) );
  INVX0 U11690 ( .INP(n11904), .ZN(n11902) );
  NOR2X0 U11691 ( .IN1(n11905), .IN2(n8740), .QN(n11904) );
  NAND2X0 U11692 ( .IN1(n11906), .IN2(n11907), .QN(g29194) );
  NAND2X0 U11693 ( .IN1(n11884), .IN2(g5437), .QN(n11907) );
  XNOR2X1 U11694 ( .IN1(n11908), .IN2(n11909), .Q(n11884) );
  NOR2X0 U11695 ( .IN1(n11910), .IN2(n11911), .QN(n11909) );
  NAND2X0 U11696 ( .IN1(n11912), .IN2(g309), .QN(n11911) );
  NAND2X0 U11697 ( .IN1(n11913), .IN2(n10459), .QN(n11912) );
  NAND2X0 U11698 ( .IN1(n10733), .IN2(n11908), .QN(n10459) );
  NAND2X0 U11699 ( .IN1(n11914), .IN2(n10460), .QN(n11913) );
  XNOR2X1 U11700 ( .IN1(n10461), .IN2(n11908), .Q(n11910) );
  NAND2X0 U11701 ( .IN1(n4520), .IN2(g417), .QN(n11906) );
  NAND2X0 U11702 ( .IN1(n11915), .IN2(n11916), .QN(g29187) );
  NAND2X0 U11703 ( .IN1(n11917), .IN2(g2396), .QN(n11916) );
  NAND2X0 U11704 ( .IN1(n11918), .IN2(n11841), .QN(n11917) );
  NAND2X0 U11705 ( .IN1(n11919), .IN2(n11841), .QN(n11915) );
  NAND2X0 U11706 ( .IN1(n11920), .IN2(n11921), .QN(g29185) );
  NAND2X0 U11707 ( .IN1(n11922), .IN2(g2398), .QN(n11921) );
  NAND2X0 U11708 ( .IN1(n11918), .IN2(n10669), .QN(n11922) );
  NAND2X0 U11709 ( .IN1(n11919), .IN2(n10669), .QN(n11920) );
  NAND2X0 U11710 ( .IN1(n11923), .IN2(n11924), .QN(g29184) );
  NAND2X0 U11711 ( .IN1(n11925), .IN2(g1702), .QN(n11924) );
  NAND2X0 U11712 ( .IN1(n11926), .IN2(n11849), .QN(n11925) );
  NAND2X0 U11713 ( .IN1(n11927), .IN2(n11849), .QN(n11923) );
  NAND2X0 U11714 ( .IN1(n11928), .IN2(n11929), .QN(g29182) );
  NAND2X0 U11715 ( .IN1(n11930), .IN2(g2397), .QN(n11929) );
  NAND2X0 U11716 ( .IN1(n11918), .IN2(n11931), .QN(n11930) );
  NAND2X0 U11717 ( .IN1(n11919), .IN2(n11931), .QN(n11928) );
  NOR2X0 U11718 ( .IN1(n11932), .IN2(n11918), .QN(n11919) );
  NOR2X0 U11719 ( .IN1(n11932), .IN2(n11933), .QN(n11918) );
  INVX0 U11720 ( .INP(n11934), .ZN(n11933) );
  NAND2X0 U11721 ( .IN1(n3036), .IN2(n11935), .QN(n11934) );
  NAND2X0 U11722 ( .IN1(n11936), .IN2(n11937), .QN(n11935) );
  NOR2X0 U11723 ( .IN1(n11106), .IN2(n11114), .QN(n11937) );
  NOR2X0 U11724 ( .IN1(n11938), .IN2(n11187), .QN(n11936) );
  NAND2X0 U11725 ( .IN1(n11121), .IN2(n11122), .QN(n11187) );
  NAND2X0 U11726 ( .IN1(n3038), .IN2(n11939), .QN(n11122) );
  NAND2X0 U11727 ( .IN1(n11940), .IN2(n11941), .QN(n11939) );
  NAND2X0 U11728 ( .IN1(n11942), .IN2(n11943), .QN(n11941) );
  NOR2X0 U11729 ( .IN1(n11944), .IN2(n11945), .QN(n11942) );
  NOR2X0 U11730 ( .IN1(n11946), .IN2(n11947), .QN(n11945) );
  INVX0 U11731 ( .INP(n11948), .ZN(n11947) );
  NOR2X0 U11732 ( .IN1(n11949), .IN2(n11950), .QN(n11944) );
  NOR2X0 U11733 ( .IN1(n11951), .IN2(n11952), .QN(n11940) );
  NOR2X0 U11734 ( .IN1(n11953), .IN2(n11954), .QN(n11952) );
  NAND2X0 U11735 ( .IN1(n11955), .IN2(n11956), .QN(n11954) );
  NAND2X0 U11736 ( .IN1(n11957), .IN2(n11958), .QN(n11956) );
  NAND2X0 U11737 ( .IN1(n11959), .IN2(n11948), .QN(n11955) );
  NOR2X0 U11738 ( .IN1(n11959), .IN2(n11960), .QN(n11951) );
  NAND2X0 U11739 ( .IN1(n11961), .IN2(n11962), .QN(n11960) );
  NAND2X0 U11740 ( .IN1(n11958), .IN2(n11953), .QN(n11962) );
  INVX0 U11741 ( .INP(n11946), .ZN(n11953) );
  INVX0 U11742 ( .INP(n11949), .ZN(n11958) );
  NAND2X0 U11743 ( .IN1(n11957), .IN2(n11948), .QN(n11961) );
  NAND2X0 U11744 ( .IN1(n3038), .IN2(n11129), .QN(n11121) );
  NAND2X0 U11745 ( .IN1(n11963), .IN2(n11964), .QN(n11129) );
  NAND2X0 U11746 ( .IN1(n11965), .IN2(n11966), .QN(n11964) );
  NOR2X0 U11747 ( .IN1(n11967), .IN2(n11968), .QN(n11965) );
  NOR2X0 U11748 ( .IN1(n11969), .IN2(n11970), .QN(n11968) );
  NOR2X0 U11749 ( .IN1(n11971), .IN2(n11972), .QN(n11967) );
  INVX0 U11750 ( .INP(n11973), .ZN(n11972) );
  NOR2X0 U11751 ( .IN1(n11974), .IN2(n11975), .QN(n11963) );
  NOR2X0 U11752 ( .IN1(n11973), .IN2(n11976), .QN(n11975) );
  NAND2X0 U11753 ( .IN1(n11977), .IN2(n11978), .QN(n11976) );
  NAND2X0 U11754 ( .IN1(n11979), .IN2(n11980), .QN(n11978) );
  NAND2X0 U11755 ( .IN1(n11981), .IN2(n11982), .QN(n11977) );
  NOR2X0 U11756 ( .IN1(n11979), .IN2(n11983), .QN(n11974) );
  NAND2X0 U11757 ( .IN1(n11984), .IN2(n11985), .QN(n11983) );
  NAND2X0 U11758 ( .IN1(n11981), .IN2(n11973), .QN(n11985) );
  NAND2X0 U11759 ( .IN1(n11982), .IN2(n11980), .QN(n11984) );
  INVX0 U11760 ( .INP(n11971), .ZN(n11980) );
  INVX0 U11761 ( .INP(n11966), .ZN(n11982) );
  NAND2X0 U11762 ( .IN1(n11477), .IN2(n11479), .QN(n3036) );
  INVX0 U11763 ( .INP(n11938), .ZN(n11479) );
  NOR2X0 U11764 ( .IN1(n11986), .IN2(n11987), .QN(n11932) );
  NOR2X0 U11765 ( .IN1(n11192), .IN2(n11477), .QN(n11987) );
  NAND2X0 U11766 ( .IN1(n11131), .IN2(n3038), .QN(n11192) );
  NAND2X0 U11767 ( .IN1(n11988), .IN2(n11989), .QN(n11131) );
  NOR2X0 U11768 ( .IN1(n11990), .IN2(n11991), .QN(n11989) );
  NAND2X0 U11769 ( .IN1(n11959), .IN2(n11957), .QN(n11991) );
  INVX0 U11770 ( .INP(n11943), .ZN(n11957) );
  XNOR2X1 U11771 ( .IN1(n11463), .IN2(g2190), .Q(n11943) );
  INVX0 U11772 ( .INP(n9865), .ZN(n11463) );
  NAND2X0 U11773 ( .IN1(n11992), .IN2(n11993), .QN(n9865) );
  NAND2X0 U11774 ( .IN1(test_so77), .IN2(test_so73), .QN(n11993) );
  NOR2X0 U11775 ( .IN1(n11994), .IN2(n11995), .QN(n11992) );
  NOR2X0 U11776 ( .IN1(n8418), .IN2(n4367), .QN(n11995) );
  NOR2X0 U11777 ( .IN1(n8434), .IN2(n4324), .QN(n11994) );
  INVX0 U11778 ( .INP(n11950), .ZN(n11959) );
  XNOR2X1 U11779 ( .IN1(n9863), .IN2(n11996), .Q(n11950) );
  INVX0 U11780 ( .INP(n10800), .ZN(n9863) );
  NAND2X0 U11781 ( .IN1(n11997), .IN2(n11998), .QN(n10800) );
  NAND2X0 U11782 ( .IN1(test_so73), .IN2(g2345), .QN(n11998) );
  NOR2X0 U11783 ( .IN1(n11999), .IN2(n12000), .QN(n11997) );
  NOR2X0 U11784 ( .IN1(n8376), .IN2(n4367), .QN(n12000) );
  NOR2X0 U11785 ( .IN1(n8377), .IN2(n4324), .QN(n11999) );
  NAND2X0 U11786 ( .IN1(n12001), .IN2(n11948), .QN(n11990) );
  XNOR2X1 U11787 ( .IN1(n9844), .IN2(g2200), .Q(n11948) );
  NAND2X0 U11788 ( .IN1(n12002), .IN2(n12003), .QN(n9844) );
  NAND2X0 U11789 ( .IN1(test_so73), .IN2(g2336), .QN(n12003) );
  NOR2X0 U11790 ( .IN1(n12004), .IN2(n12005), .QN(n12002) );
  NOR2X0 U11791 ( .IN1(n8527), .IN2(n4367), .QN(n12005) );
  NOR2X0 U11792 ( .IN1(n8431), .IN2(n4324), .QN(n12004) );
  NOR2X0 U11793 ( .IN1(n11946), .IN2(n11949), .QN(n12001) );
  XOR2X1 U11794 ( .IN1(n9864), .IN2(g2180), .Q(n11949) );
  NAND2X0 U11795 ( .IN1(n12006), .IN2(n12007), .QN(n9864) );
  NAND2X0 U11796 ( .IN1(test_so73), .IN2(g2318), .QN(n12007) );
  NOR2X0 U11797 ( .IN1(n12008), .IN2(n12009), .QN(n12006) );
  NOR2X0 U11798 ( .IN1(n8419), .IN2(n4367), .QN(n12009) );
  NOR2X0 U11799 ( .IN1(n8437), .IN2(n4324), .QN(n12008) );
  XNOR2X1 U11800 ( .IN1(n9858), .IN2(g2170), .Q(n11946) );
  INVX0 U11801 ( .INP(n11491), .ZN(n9858) );
  NAND2X0 U11802 ( .IN1(n12010), .IN2(n12011), .QN(n11491) );
  NAND2X0 U11803 ( .IN1(test_so73), .IN2(g2309), .QN(n12011) );
  NOR2X0 U11804 ( .IN1(n12012), .IN2(n12013), .QN(n12010) );
  NOR2X0 U11805 ( .IN1(n8420), .IN2(n4367), .QN(n12013) );
  NOR2X0 U11806 ( .IN1(n8440), .IN2(n4324), .QN(n12012) );
  NOR2X0 U11807 ( .IN1(n12014), .IN2(n12015), .QN(n11988) );
  NAND2X0 U11808 ( .IN1(n11979), .IN2(n11981), .QN(n12015) );
  INVX0 U11809 ( .INP(n11969), .ZN(n11981) );
  XNOR2X1 U11810 ( .IN1(n9850), .IN2(g2175), .Q(n11969) );
  INVX0 U11811 ( .INP(n11458), .ZN(n9850) );
  NAND2X0 U11812 ( .IN1(n12016), .IN2(n12017), .QN(n11458) );
  NAND2X0 U11813 ( .IN1(test_so73), .IN2(g2273), .QN(n12017) );
  NOR2X0 U11814 ( .IN1(n12018), .IN2(n12019), .QN(n12016) );
  NOR2X0 U11815 ( .IN1(n8536), .IN2(n4367), .QN(n12019) );
  NOR2X0 U11816 ( .IN1(n8439), .IN2(n4324), .QN(n12018) );
  INVX0 U11817 ( .INP(n11970), .ZN(n11979) );
  XNOR2X1 U11818 ( .IN1(n9851), .IN2(n12020), .Q(n11970) );
  INVX0 U11819 ( .INP(n11492), .ZN(n9851) );
  NAND2X0 U11820 ( .IN1(n12021), .IN2(n12022), .QN(n11492) );
  NAND2X0 U11821 ( .IN1(test_so73), .IN2(g2300), .QN(n12022) );
  NOR2X0 U11822 ( .IN1(n12023), .IN2(n12024), .QN(n12021) );
  NOR2X0 U11823 ( .IN1(n8384), .IN2(n4367), .QN(n12024) );
  NOR2X0 U11824 ( .IN1(n8378), .IN2(n4324), .QN(n12023) );
  NAND2X0 U11825 ( .IN1(n12025), .IN2(n11973), .QN(n12014) );
  XNOR2X1 U11826 ( .IN1(n9845), .IN2(g2165), .Q(n11973) );
  NAND2X0 U11827 ( .IN1(n12026), .IN2(n12027), .QN(n9845) );
  NAND2X0 U11828 ( .IN1(test_so76), .IN2(test_so73), .QN(n12027) );
  NOR2X0 U11829 ( .IN1(n12028), .IN2(n12029), .QN(n12026) );
  NOR2X0 U11830 ( .IN1(n8537), .IN2(n4367), .QN(n12029) );
  NOR2X0 U11831 ( .IN1(n8441), .IN2(n4324), .QN(n12028) );
  NOR2X0 U11832 ( .IN1(n11971), .IN2(n11966), .QN(n12025) );
  XNOR2X1 U11833 ( .IN1(n11464), .IN2(g2185), .Q(n11966) );
  INVX0 U11834 ( .INP(n9852), .ZN(n11464) );
  NAND2X0 U11835 ( .IN1(n12030), .IN2(n12031), .QN(n9852) );
  NAND2X0 U11836 ( .IN1(test_so73), .IN2(g2282), .QN(n12031) );
  NOR2X0 U11837 ( .IN1(n12032), .IN2(n12033), .QN(n12030) );
  NOR2X0 U11838 ( .IN1(n8530), .IN2(n4367), .QN(n12033) );
  NOR2X0 U11839 ( .IN1(n8436), .IN2(n4324), .QN(n12032) );
  XNOR2X1 U11840 ( .IN1(n9843), .IN2(g2195), .Q(n11971) );
  INVX0 U11841 ( .INP(n11304), .ZN(n9843) );
  NAND2X0 U11842 ( .IN1(n12034), .IN2(n12035), .QN(n11304) );
  NAND2X0 U11843 ( .IN1(test_so73), .IN2(g2291), .QN(n12035) );
  NOR2X0 U11844 ( .IN1(n12036), .IN2(n12037), .QN(n12034) );
  NOR2X0 U11845 ( .IN1(n8535), .IN2(n4367), .QN(n12037) );
  NOR2X0 U11846 ( .IN1(n8433), .IN2(n4324), .QN(n12036) );
  NOR2X0 U11847 ( .IN1(n12038), .IN2(n9281), .QN(n11986) );
  NAND2X0 U11848 ( .IN1(n12039), .IN2(n12040), .QN(g29181) );
  NAND2X0 U11849 ( .IN1(n12041), .IN2(g1704), .QN(n12040) );
  NAND2X0 U11850 ( .IN1(n11926), .IN2(n10678), .QN(n12041) );
  NAND2X0 U11851 ( .IN1(n11927), .IN2(n10678), .QN(n12039) );
  NAND2X0 U11852 ( .IN1(n12042), .IN2(n12043), .QN(g29179) );
  NAND2X0 U11853 ( .IN1(n12044), .IN2(g1008), .QN(n12043) );
  NAND2X0 U11854 ( .IN1(n12045), .IN2(g1088), .QN(n12044) );
  NAND2X0 U11855 ( .IN1(n12046), .IN2(g1088), .QN(n12042) );
  NAND2X0 U11856 ( .IN1(n12047), .IN2(n12048), .QN(g29178) );
  NAND2X0 U11857 ( .IN1(n12049), .IN2(g1703), .QN(n12048) );
  NAND2X0 U11858 ( .IN1(n11926), .IN2(n12050), .QN(n12049) );
  NAND2X0 U11859 ( .IN1(n11927), .IN2(n12050), .QN(n12047) );
  NOR2X0 U11860 ( .IN1(n12051), .IN2(n11926), .QN(n11927) );
  NOR2X0 U11861 ( .IN1(n12051), .IN2(n12052), .QN(n11926) );
  NOR2X0 U11862 ( .IN1(n10456), .IN2(n12053), .QN(n12052) );
  INVX0 U11863 ( .INP(n12054), .ZN(n12053) );
  NAND2X0 U11864 ( .IN1(n12055), .IN2(n12056), .QN(n12054) );
  NOR2X0 U11865 ( .IN1(n11540), .IN2(n10690), .QN(n12056) );
  INVX0 U11866 ( .INP(n11206), .ZN(n11540) );
  NAND2X0 U11867 ( .IN1(n3070), .IN2(n12057), .QN(n11206) );
  NAND2X0 U11868 ( .IN1(n10699), .IN2(n10708), .QN(n12057) );
  INVX0 U11869 ( .INP(n12058), .ZN(n10708) );
  NAND2X0 U11870 ( .IN1(n12059), .IN2(n12060), .QN(n12058) );
  NAND2X0 U11871 ( .IN1(n12061), .IN2(n12062), .QN(n12060) );
  NOR2X0 U11872 ( .IN1(n12063), .IN2(n12064), .QN(n12061) );
  INVX0 U11873 ( .INP(n12065), .ZN(n12063) );
  NAND2X0 U11874 ( .IN1(n12066), .IN2(n12067), .QN(n12065) );
  NOR2X0 U11875 ( .IN1(n12068), .IN2(n12069), .QN(n12059) );
  NOR2X0 U11876 ( .IN1(n12070), .IN2(n12071), .QN(n12069) );
  NAND2X0 U11877 ( .IN1(n12072), .IN2(n12073), .QN(n12071) );
  NAND2X0 U11878 ( .IN1(n12074), .IN2(n12066), .QN(n12073) );
  NAND2X0 U11879 ( .IN1(n12067), .IN2(n12075), .QN(n12072) );
  NOR2X0 U11880 ( .IN1(n12067), .IN2(n12076), .QN(n12068) );
  NAND2X0 U11881 ( .IN1(n12077), .IN2(n12078), .QN(n12076) );
  NAND2X0 U11882 ( .IN1(n12066), .IN2(n12070), .QN(n12078) );
  INVX0 U11883 ( .INP(n12079), .ZN(n12070) );
  NAND2X0 U11884 ( .IN1(n12074), .IN2(n12075), .QN(n12077) );
  INVX0 U11885 ( .INP(n12080), .ZN(n12075) );
  INVX0 U11886 ( .INP(n12081), .ZN(n10699) );
  NAND2X0 U11887 ( .IN1(n12082), .IN2(n12083), .QN(n12081) );
  NAND2X0 U11888 ( .IN1(n12084), .IN2(n12085), .QN(n12083) );
  NOR2X0 U11889 ( .IN1(n12086), .IN2(n12087), .QN(n12084) );
  NOR2X0 U11890 ( .IN1(n12088), .IN2(n12089), .QN(n12087) );
  NOR2X0 U11891 ( .IN1(n12090), .IN2(n12091), .QN(n12086) );
  NOR2X0 U11892 ( .IN1(n12092), .IN2(n12093), .QN(n12082) );
  NOR2X0 U11893 ( .IN1(n12094), .IN2(n12095), .QN(n12093) );
  NAND2X0 U11894 ( .IN1(n12096), .IN2(n12097), .QN(n12095) );
  NAND2X0 U11895 ( .IN1(n12098), .IN2(n12099), .QN(n12097) );
  NAND2X0 U11896 ( .IN1(n12100), .IN2(n12101), .QN(n12096) );
  NOR2X0 U11897 ( .IN1(n12098), .IN2(n12102), .QN(n12092) );
  NAND2X0 U11898 ( .IN1(n12103), .IN2(n12104), .QN(n12102) );
  NAND2X0 U11899 ( .IN1(n12094), .IN2(n12101), .QN(n12104) );
  INVX0 U11900 ( .INP(n12088), .ZN(n12101) );
  NAND2X0 U11901 ( .IN1(n12099), .IN2(n12100), .QN(n12103) );
  INVX0 U11902 ( .INP(n12085), .ZN(n12100) );
  NOR2X0 U11903 ( .IN1(n10700), .IN2(n11543), .QN(n12055) );
  NOR2X0 U11904 ( .IN1(n11784), .IN2(n11543), .QN(n10456) );
  NOR2X0 U11905 ( .IN1(n12105), .IN2(n12106), .QN(n12051) );
  NOR2X0 U11906 ( .IN1(n11784), .IN2(n4386), .QN(n12106) );
  NOR2X0 U11907 ( .IN1(n11211), .IN2(n12107), .QN(n12105) );
  NAND2X0 U11908 ( .IN1(n10709), .IN2(n3070), .QN(n11211) );
  NAND2X0 U11909 ( .IN1(n12108), .IN2(n12109), .QN(n10709) );
  NOR2X0 U11910 ( .IN1(n12110), .IN2(n12111), .QN(n12109) );
  NAND2X0 U11911 ( .IN1(n12098), .IN2(n12094), .QN(n12111) );
  INVX0 U11912 ( .INP(n12091), .ZN(n12094) );
  XNOR2X1 U11913 ( .IN1(n11320), .IN2(g1471), .Q(n12091) );
  INVX0 U11914 ( .INP(n9810), .ZN(n11320) );
  NAND2X0 U11915 ( .IN1(n12112), .IN2(n12113), .QN(n9810) );
  NAND2X0 U11916 ( .IN1(g6782), .IN2(g1570), .QN(n12113) );
  NOR2X0 U11917 ( .IN1(n12114), .IN2(n12115), .QN(n12112) );
  NOR2X0 U11918 ( .IN1(n8540), .IN2(n4368), .QN(n12115) );
  NOR2X0 U11919 ( .IN1(n8454), .IN2(n4317), .QN(n12114) );
  INVX0 U11920 ( .INP(n12089), .ZN(n12098) );
  XNOR2X1 U11921 ( .IN1(n9816), .IN2(n12116), .Q(n12089) );
  INVX0 U11922 ( .INP(n10502), .ZN(n9816) );
  NAND2X0 U11923 ( .IN1(n12117), .IN2(n12118), .QN(n10502) );
  NAND2X0 U11924 ( .IN1(test_so56), .IN2(g6782), .QN(n12118) );
  NOR2X0 U11925 ( .IN1(n12119), .IN2(n12120), .QN(n12117) );
  NOR2X0 U11926 ( .IN1(n8385), .IN2(n4368), .QN(n12120) );
  NOR2X0 U11927 ( .IN1(n8379), .IN2(n4317), .QN(n12119) );
  NAND2X0 U11928 ( .IN1(n12121), .IN2(n12099), .QN(n12110) );
  INVX0 U11929 ( .INP(n12090), .ZN(n12099) );
  XNOR2X1 U11930 ( .IN1(n9808), .IN2(g1501), .Q(n12090) );
  INVX0 U11931 ( .INP(n11515), .ZN(n9808) );
  NAND2X0 U11932 ( .IN1(n12122), .IN2(n12123), .QN(n11515) );
  NAND2X0 U11933 ( .IN1(g6782), .IN2(g1597), .QN(n12123) );
  NOR2X0 U11934 ( .IN1(n12124), .IN2(n12125), .QN(n12122) );
  NOR2X0 U11935 ( .IN1(n8538), .IN2(n4368), .QN(n12125) );
  NOR2X0 U11936 ( .IN1(n8445), .IN2(n4317), .QN(n12124) );
  NOR2X0 U11937 ( .IN1(n12088), .IN2(n12085), .QN(n12121) );
  XNOR2X1 U11938 ( .IN1(n11526), .IN2(g1491), .Q(n12085) );
  INVX0 U11939 ( .INP(n9817), .ZN(n11526) );
  NAND2X0 U11940 ( .IN1(n12126), .IN2(n12127), .QN(n9817) );
  NAND2X0 U11941 ( .IN1(g6782), .IN2(g1588), .QN(n12127) );
  NOR2X0 U11942 ( .IN1(n12128), .IN2(n12129), .QN(n12126) );
  NOR2X0 U11943 ( .IN1(n8531), .IN2(n4368), .QN(n12129) );
  NOR2X0 U11944 ( .IN1(n8449), .IN2(n4317), .QN(n12128) );
  XNOR2X1 U11945 ( .IN1(n9815), .IN2(g1481), .Q(n12088) );
  INVX0 U11946 ( .INP(n11553), .ZN(n9815) );
  NAND2X0 U11947 ( .IN1(n12130), .IN2(n12131), .QN(n11553) );
  NAND2X0 U11948 ( .IN1(g6782), .IN2(g1579), .QN(n12131) );
  NOR2X0 U11949 ( .IN1(n12132), .IN2(n12133), .QN(n12130) );
  NOR2X0 U11950 ( .IN1(n8539), .IN2(n4368), .QN(n12133) );
  NOR2X0 U11951 ( .IN1(n8451), .IN2(n4317), .QN(n12132) );
  NOR2X0 U11952 ( .IN1(n12134), .IN2(n12135), .QN(n12108) );
  NAND2X0 U11953 ( .IN1(n12067), .IN2(n12074), .QN(n12135) );
  INVX0 U11954 ( .INP(n12062), .ZN(n12074) );
  XNOR2X1 U11955 ( .IN1(n9829), .IN2(g1496), .Q(n12062) );
  INVX0 U11956 ( .INP(n11384), .ZN(n9829) );
  NAND2X0 U11957 ( .IN1(n12136), .IN2(n12137), .QN(n11384) );
  NAND2X0 U11958 ( .IN1(g6782), .IN2(g1633), .QN(n12137) );
  NOR2X0 U11959 ( .IN1(n12138), .IN2(n12139), .QN(n12136) );
  NOR2X0 U11960 ( .IN1(n8421), .IN2(n4368), .QN(n12139) );
  NOR2X0 U11961 ( .IN1(n8447), .IN2(n4317), .QN(n12138) );
  XOR2X1 U11962 ( .IN1(n10835), .IN2(n9830), .Q(n12067) );
  NAND2X0 U11963 ( .IN1(n12140), .IN2(n12141), .QN(n9830) );
  NAND2X0 U11964 ( .IN1(g6782), .IN2(g1651), .QN(n12141) );
  NOR2X0 U11965 ( .IN1(n12142), .IN2(n12143), .QN(n12140) );
  NOR2X0 U11966 ( .IN1(n8413), .IN2(n4368), .QN(n12143) );
  NOR2X0 U11967 ( .IN1(n8412), .IN2(n4317), .QN(n12142) );
  NAND2X0 U11968 ( .IN1(n12064), .IN2(n12066), .QN(n12134) );
  XNOR2X1 U11969 ( .IN1(n9823), .IN2(g1486), .Q(n12066) );
  NAND2X0 U11970 ( .IN1(n12144), .IN2(n12145), .QN(n9823) );
  NAND2X0 U11971 ( .IN1(g6782), .IN2(g1624), .QN(n12145) );
  NOR2X0 U11972 ( .IN1(n12146), .IN2(n12147), .QN(n12144) );
  NOR2X0 U11973 ( .IN1(n8422), .IN2(n4368), .QN(n12147) );
  INVX0 U11974 ( .INP(n12148), .ZN(n12146) );
  NAND2X0 U11975 ( .IN1(g6573), .IN2(test_so55), .QN(n12148) );
  NOR2X0 U11976 ( .IN1(n12080), .IN2(n12079), .QN(n12064) );
  XNOR2X1 U11977 ( .IN1(n9828), .IN2(g1476), .Q(n12079) );
  INVX0 U11978 ( .INP(n11521), .ZN(n9828) );
  NAND2X0 U11979 ( .IN1(n12149), .IN2(n12150), .QN(n11521) );
  NAND2X0 U11980 ( .IN1(g6782), .IN2(g1615), .QN(n12150) );
  NOR2X0 U11981 ( .IN1(n12151), .IN2(n12152), .QN(n12149) );
  NOR2X0 U11982 ( .IN1(n8423), .IN2(n4368), .QN(n12152) );
  NOR2X0 U11983 ( .IN1(n8452), .IN2(n4317), .QN(n12151) );
  XNOR2X1 U11984 ( .IN1(n9809), .IN2(g1506), .Q(n12080) );
  INVX0 U11985 ( .INP(n11029), .ZN(n9809) );
  NAND2X0 U11986 ( .IN1(n12153), .IN2(n12154), .QN(n11029) );
  NAND2X0 U11987 ( .IN1(g6782), .IN2(g1642), .QN(n12154) );
  NOR2X0 U11988 ( .IN1(n12155), .IN2(n12156), .QN(n12153) );
  NOR2X0 U11989 ( .IN1(n8528), .IN2(n4368), .QN(n12156) );
  NOR2X0 U11990 ( .IN1(n8443), .IN2(n4317), .QN(n12155) );
  NAND2X0 U11991 ( .IN1(n12157), .IN2(n12158), .QN(g29173) );
  NAND2X0 U11992 ( .IN1(n12159), .IN2(g1010), .QN(n12158) );
  NAND2X0 U11993 ( .IN1(n12045), .IN2(g6712), .QN(n12159) );
  NAND2X0 U11994 ( .IN1(n12046), .IN2(g6712), .QN(n12157) );
  NAND2X0 U11995 ( .IN1(n12160), .IN2(n12161), .QN(g29172) );
  NAND2X0 U11996 ( .IN1(n12162), .IN2(g321), .QN(n12161) );
  NAND2X0 U11997 ( .IN1(n12163), .IN2(n11886), .QN(n12162) );
  NAND2X0 U11998 ( .IN1(n12164), .IN2(n11886), .QN(n12160) );
  NAND2X0 U11999 ( .IN1(n12165), .IN2(n12166), .QN(g29170) );
  NAND2X0 U12000 ( .IN1(n12167), .IN2(g1009), .QN(n12166) );
  NAND2X0 U12001 ( .IN1(n12045), .IN2(g5472), .QN(n12167) );
  NAND2X0 U12002 ( .IN1(n12046), .IN2(g5472), .QN(n12165) );
  NOR2X0 U12003 ( .IN1(n12168), .IN2(n12045), .QN(n12046) );
  INVX0 U12004 ( .INP(n3065), .ZN(n12045) );
  NAND2X0 U12005 ( .IN1(n12169), .IN2(n11603), .QN(n3065) );
  NOR2X0 U12006 ( .IN1(n12170), .IN2(n12171), .QN(n12169) );
  NOR2X0 U12007 ( .IN1(n11601), .IN2(n12172), .QN(n12171) );
  NOR2X0 U12008 ( .IN1(n10499), .IN2(n12173), .QN(n12172) );
  NAND2X0 U12009 ( .IN1(n10486), .IN2(n10494), .QN(n12173) );
  NAND2X0 U12010 ( .IN1(n3102), .IN2(n12174), .QN(n10494) );
  INVX0 U12011 ( .INP(n12175), .ZN(n12174) );
  NOR2X0 U12012 ( .IN1(n10523), .IN2(n10524), .QN(n12175) );
  NAND2X0 U12013 ( .IN1(n12176), .IN2(n12177), .QN(n10524) );
  NAND2X0 U12014 ( .IN1(n12178), .IN2(n12179), .QN(n12177) );
  NOR2X0 U12015 ( .IN1(n12180), .IN2(n12181), .QN(n12178) );
  NOR2X0 U12016 ( .IN1(n12182), .IN2(n12183), .QN(n12181) );
  NOR2X0 U12017 ( .IN1(n12184), .IN2(n12185), .QN(n12180) );
  NOR2X0 U12018 ( .IN1(n12186), .IN2(n12187), .QN(n12176) );
  NOR2X0 U12019 ( .IN1(n12188), .IN2(n12189), .QN(n12187) );
  NAND2X0 U12020 ( .IN1(n12190), .IN2(n12191), .QN(n12189) );
  NAND2X0 U12021 ( .IN1(n12192), .IN2(n12193), .QN(n12191) );
  NOR2X0 U12022 ( .IN1(n12194), .IN2(n12195), .QN(n12186) );
  NAND2X0 U12023 ( .IN1(n12196), .IN2(n12197), .QN(n12195) );
  NAND2X0 U12024 ( .IN1(n12188), .IN2(n12193), .QN(n12197) );
  INVX0 U12025 ( .INP(n12184), .ZN(n12193) );
  NAND2X0 U12026 ( .IN1(n12198), .IN2(n12192), .QN(n12196) );
  NAND2X0 U12027 ( .IN1(n12199), .IN2(n12200), .QN(n10523) );
  NAND2X0 U12028 ( .IN1(n12201), .IN2(n12202), .QN(n12200) );
  NOR2X0 U12029 ( .IN1(n12203), .IN2(n12204), .QN(n12201) );
  NOR2X0 U12030 ( .IN1(n12205), .IN2(n12206), .QN(n12204) );
  INVX0 U12031 ( .INP(n12207), .ZN(n12203) );
  NOR2X0 U12032 ( .IN1(n12208), .IN2(n12209), .QN(n12199) );
  NOR2X0 U12033 ( .IN1(n12210), .IN2(n12211), .QN(n12209) );
  NAND2X0 U12034 ( .IN1(n12212), .IN2(n12213), .QN(n12211) );
  NAND2X0 U12035 ( .IN1(n12214), .IN2(n12215), .QN(n12213) );
  NAND2X0 U12036 ( .IN1(n12216), .IN2(n12217), .QN(n12212) );
  NOR2X0 U12037 ( .IN1(n12214), .IN2(n12218), .QN(n12208) );
  NAND2X0 U12038 ( .IN1(n12219), .IN2(n12220), .QN(n12218) );
  NAND2X0 U12039 ( .IN1(n12217), .IN2(n12215), .QN(n12220) );
  INVX0 U12040 ( .INP(n12205), .ZN(n12215) );
  INVX0 U12041 ( .INP(n12202), .ZN(n12217) );
  NAND2X0 U12042 ( .IN1(n12216), .IN2(n12210), .QN(n12219) );
  NAND2X0 U12043 ( .IN1(n12221), .IN2(n3102), .QN(n10499) );
  NOR2X0 U12044 ( .IN1(n10507), .IN2(n12222), .QN(n12221) );
  INVX0 U12045 ( .INP(n12223), .ZN(n12168) );
  NOR2X0 U12046 ( .IN1(n12170), .IN2(n12224), .QN(n12223) );
  NOR2X0 U12047 ( .IN1(n11601), .IN2(n12225), .QN(n12224) );
  NOR2X0 U12048 ( .IN1(n12222), .IN2(n10519), .QN(n12225) );
  INVX0 U12049 ( .INP(n10518), .ZN(n12222) );
  NAND2X0 U12050 ( .IN1(n12226), .IN2(n12227), .QN(n10518) );
  NOR2X0 U12051 ( .IN1(n12228), .IN2(n12207), .QN(n12227) );
  NAND2X0 U12052 ( .IN1(n12216), .IN2(n12214), .QN(n12207) );
  XOR2X1 U12053 ( .IN1(n9793), .IN2(n10876), .Q(n12214) );
  NAND2X0 U12054 ( .IN1(n12229), .IN2(n12230), .QN(n9793) );
  NAND2X0 U12055 ( .IN1(test_so31), .IN2(g960), .QN(n12230) );
  NOR2X0 U12056 ( .IN1(n12231), .IN2(n12232), .QN(n12229) );
  NOR2X0 U12057 ( .IN1(n8455), .IN2(n4323), .QN(n12232) );
  NOR2X0 U12058 ( .IN1(n8491), .IN2(n4312), .QN(n12231) );
  XNOR2X1 U12059 ( .IN1(n11004), .IN2(n4391), .Q(n12216) );
  INVX0 U12060 ( .INP(n9782), .ZN(n11004) );
  NAND2X0 U12061 ( .IN1(n12233), .IN2(n12234), .QN(n9782) );
  NAND2X0 U12062 ( .IN1(test_so31), .IN2(g933), .QN(n12234) );
  NOR2X0 U12063 ( .IN1(n12235), .IN2(n12236), .QN(n12233) );
  NOR2X0 U12064 ( .IN1(n8464), .IN2(n4323), .QN(n12236) );
  NOR2X0 U12065 ( .IN1(n8487), .IN2(n4312), .QN(n12235) );
  NAND2X0 U12066 ( .IN1(n12237), .IN2(n12210), .QN(n12228) );
  INVX0 U12067 ( .INP(n12206), .ZN(n12210) );
  XNOR2X1 U12068 ( .IN1(n9781), .IN2(g789), .Q(n12206) );
  INVX0 U12069 ( .INP(n11584), .ZN(n9781) );
  NAND2X0 U12070 ( .IN1(n12238), .IN2(n12239), .QN(n11584) );
  NAND2X0 U12071 ( .IN1(test_so34), .IN2(test_so31), .QN(n12239) );
  NOR2X0 U12072 ( .IN1(n12240), .IN2(n12241), .QN(n12238) );
  NOR2X0 U12073 ( .IN1(n8467), .IN2(n4323), .QN(n12241) );
  NOR2X0 U12074 ( .IN1(n8488), .IN2(n4312), .QN(n12240) );
  NOR2X0 U12075 ( .IN1(n12205), .IN2(n12202), .QN(n12237) );
  XNOR2X1 U12076 ( .IN1(n9774), .IN2(g805), .Q(n12202) );
  INVX0 U12077 ( .INP(n11420), .ZN(n9774) );
  NAND2X0 U12078 ( .IN1(n12242), .IN2(n12243), .QN(n11420) );
  NAND2X0 U12079 ( .IN1(test_so31), .IN2(g942), .QN(n12243) );
  NOR2X0 U12080 ( .IN1(n12244), .IN2(n12245), .QN(n12242) );
  NOR2X0 U12081 ( .IN1(n8461), .IN2(n4323), .QN(n12245) );
  NOR2X0 U12082 ( .IN1(n8460), .IN2(n4312), .QN(n12244) );
  XNOR2X1 U12083 ( .IN1(n9788), .IN2(g813), .Q(n12205) );
  INVX0 U12084 ( .INP(n11071), .ZN(n9788) );
  NAND2X0 U12085 ( .IN1(n12246), .IN2(n12247), .QN(n11071) );
  NAND2X0 U12086 ( .IN1(test_so31), .IN2(g951), .QN(n12247) );
  NOR2X0 U12087 ( .IN1(n12248), .IN2(n12249), .QN(n12246) );
  INVX0 U12088 ( .INP(n12250), .ZN(n12249) );
  NAND2X0 U12089 ( .IN1(g6368), .IN2(test_so35), .QN(n12250) );
  NOR2X0 U12090 ( .IN1(n8457), .IN2(n4312), .QN(n12248) );
  NOR2X0 U12091 ( .IN1(n12251), .IN2(n12190), .QN(n12226) );
  NAND2X0 U12092 ( .IN1(n12194), .IN2(n12198), .QN(n12190) );
  INVX0 U12093 ( .INP(n12183), .ZN(n12198) );
  XNOR2X1 U12094 ( .IN1(n9773), .IN2(g809), .Q(n12183) );
  INVX0 U12095 ( .INP(n11578), .ZN(n9773) );
  NAND2X0 U12096 ( .IN1(n12252), .IN2(n12253), .QN(n11578) );
  NAND2X0 U12097 ( .IN1(test_so31), .IN2(g906), .QN(n12253) );
  NOR2X0 U12098 ( .IN1(n12254), .IN2(n12255), .QN(n12252) );
  NOR2X0 U12099 ( .IN1(n8459), .IN2(n4323), .QN(n12255) );
  NOR2X0 U12100 ( .IN1(n8458), .IN2(n4312), .QN(n12254) );
  INVX0 U12101 ( .INP(n12185), .ZN(n12194) );
  XNOR2X1 U12102 ( .IN1(n12256), .IN2(n12257), .Q(n12185) );
  INVX0 U12103 ( .INP(n9795), .ZN(n12256) );
  NAND2X0 U12104 ( .IN1(n12258), .IN2(n12259), .QN(n9795) );
  NAND2X0 U12105 ( .IN1(test_so31), .IN2(g915), .QN(n12259) );
  NOR2X0 U12106 ( .IN1(n12260), .IN2(n12261), .QN(n12258) );
  NOR2X0 U12107 ( .IN1(n8456), .IN2(n4323), .QN(n12261) );
  NOR2X0 U12108 ( .IN1(n8492), .IN2(n4312), .QN(n12260) );
  NAND2X0 U12109 ( .IN1(n12262), .IN2(n12192), .QN(n12251) );
  INVX0 U12110 ( .INP(n12179), .ZN(n12192) );
  XNOR2X1 U12111 ( .IN1(n11588), .IN2(g801), .Q(n12179) );
  INVX0 U12112 ( .INP(n9775), .ZN(n11588) );
  NAND2X0 U12113 ( .IN1(n12263), .IN2(n12264), .QN(n9775) );
  NAND2X0 U12114 ( .IN1(test_so31), .IN2(g897), .QN(n12264) );
  NOR2X0 U12115 ( .IN1(n12265), .IN2(n12266), .QN(n12263) );
  NOR2X0 U12116 ( .IN1(n8463), .IN2(n4323), .QN(n12266) );
  NOR2X0 U12117 ( .IN1(n8462), .IN2(n4312), .QN(n12265) );
  NOR2X0 U12118 ( .IN1(n12184), .IN2(n12182), .QN(n12262) );
  INVX0 U12119 ( .INP(n12188), .ZN(n12182) );
  XOR2X1 U12120 ( .IN1(n9780), .IN2(n4379), .Q(n12188) );
  NAND2X0 U12121 ( .IN1(n12267), .IN2(n12268), .QN(n9780) );
  NAND2X0 U12122 ( .IN1(test_so31), .IN2(g879), .QN(n12268) );
  NOR2X0 U12123 ( .IN1(n12269), .IN2(n12270), .QN(n12267) );
  NOR2X0 U12124 ( .IN1(n8469), .IN2(n4323), .QN(n12270) );
  NOR2X0 U12125 ( .IN1(n8468), .IN2(n4312), .QN(n12269) );
  XNOR2X1 U12126 ( .IN1(n9794), .IN2(g793), .Q(n12184) );
  INVX0 U12127 ( .INP(n11617), .ZN(n9794) );
  NAND2X0 U12128 ( .IN1(n12271), .IN2(n12272), .QN(n11617) );
  NAND2X0 U12129 ( .IN1(test_so31), .IN2(g888), .QN(n12272) );
  NOR2X0 U12130 ( .IN1(n12273), .IN2(n12274), .QN(n12271) );
  NOR2X0 U12131 ( .IN1(n8466), .IN2(n4323), .QN(n12274) );
  NOR2X0 U12132 ( .IN1(n8465), .IN2(n4312), .QN(n12273) );
  NOR2X0 U12133 ( .IN1(n11798), .IN2(g996), .QN(n12170) );
  NAND2X0 U12134 ( .IN1(n12275), .IN2(n12276), .QN(g29169) );
  NAND2X0 U12135 ( .IN1(n12277), .IN2(g323), .QN(n12276) );
  NAND2X0 U12136 ( .IN1(n12163), .IN2(n11905), .QN(n12277) );
  NAND2X0 U12137 ( .IN1(n12164), .IN2(n11905), .QN(n12275) );
  NAND2X0 U12138 ( .IN1(n12278), .IN2(n12279), .QN(g29167) );
  NAND2X0 U12139 ( .IN1(n12280), .IN2(g322), .QN(n12279) );
  NAND2X0 U12140 ( .IN1(n12163), .IN2(n10752), .QN(n12280) );
  NAND2X0 U12141 ( .IN1(n12164), .IN2(n10752), .QN(n12278) );
  NOR2X0 U12142 ( .IN1(n12281), .IN2(n12163), .QN(n12164) );
  NOR2X0 U12143 ( .IN1(n12281), .IN2(n12282), .QN(n12163) );
  NOR2X0 U12144 ( .IN1(n10455), .IN2(n12283), .QN(n12282) );
  INVX0 U12145 ( .INP(n12284), .ZN(n12283) );
  NAND2X0 U12146 ( .IN1(n12285), .IN2(n12286), .QN(n12284) );
  NOR2X0 U12147 ( .IN1(n11668), .IN2(n10729), .QN(n12286) );
  INVX0 U12148 ( .INP(n11166), .ZN(n11668) );
  NAND2X0 U12149 ( .IN1(n3130), .IN2(n12287), .QN(n11166) );
  NAND2X0 U12150 ( .IN1(n10738), .IN2(n10747), .QN(n12287) );
  INVX0 U12151 ( .INP(n12288), .ZN(n10747) );
  NAND2X0 U12152 ( .IN1(n12289), .IN2(n12290), .QN(n12288) );
  NAND2X0 U12153 ( .IN1(n12291), .IN2(n12292), .QN(n12290) );
  NOR2X0 U12154 ( .IN1(n12293), .IN2(n12294), .QN(n12291) );
  NOR2X0 U12155 ( .IN1(n12295), .IN2(n12296), .QN(n12293) );
  NOR2X0 U12156 ( .IN1(n12297), .IN2(n12298), .QN(n12289) );
  NOR2X0 U12157 ( .IN1(n12299), .IN2(n12300), .QN(n12298) );
  NAND2X0 U12158 ( .IN1(n12301), .IN2(n12302), .QN(n12300) );
  NAND2X0 U12159 ( .IN1(n12303), .IN2(n12304), .QN(n12302) );
  NAND2X0 U12160 ( .IN1(n12305), .IN2(n12306), .QN(n12301) );
  NOR2X0 U12161 ( .IN1(n12305), .IN2(n12307), .QN(n12297) );
  NAND2X0 U12162 ( .IN1(n12308), .IN2(n12309), .QN(n12307) );
  NAND2X0 U12163 ( .IN1(n12304), .IN2(n12299), .QN(n12309) );
  INVX0 U12164 ( .INP(n12310), .ZN(n12299) );
  NAND2X0 U12165 ( .IN1(n12303), .IN2(n12306), .QN(n12308) );
  INVX0 U12166 ( .INP(n12311), .ZN(n12306) );
  INVX0 U12167 ( .INP(n12312), .ZN(n10738) );
  NAND2X0 U12168 ( .IN1(n12313), .IN2(n12314), .QN(n12312) );
  NAND2X0 U12169 ( .IN1(n12315), .IN2(n12316), .QN(n12314) );
  NOR2X0 U12170 ( .IN1(n12317), .IN2(n12318), .QN(n12315) );
  NOR2X0 U12171 ( .IN1(n12319), .IN2(n12320), .QN(n12318) );
  INVX0 U12172 ( .INP(n12321), .ZN(n12317) );
  NAND2X0 U12173 ( .IN1(n12322), .IN2(n12323), .QN(n12321) );
  NOR2X0 U12174 ( .IN1(n12324), .IN2(n12325), .QN(n12313) );
  NOR2X0 U12175 ( .IN1(n12323), .IN2(n12326), .QN(n12325) );
  NAND2X0 U12176 ( .IN1(n12327), .IN2(n12328), .QN(n12326) );
  NAND2X0 U12177 ( .IN1(n12329), .IN2(n12322), .QN(n12328) );
  NAND2X0 U12178 ( .IN1(n12330), .IN2(n12331), .QN(n12327) );
  NOR2X0 U12179 ( .IN1(n12329), .IN2(n12332), .QN(n12324) );
  NAND2X0 U12180 ( .IN1(n12333), .IN2(n12334), .QN(n12332) );
  NAND2X0 U12181 ( .IN1(n12323), .IN2(n12331), .QN(n12334) );
  INVX0 U12182 ( .INP(n12319), .ZN(n12331) );
  NAND2X0 U12183 ( .IN1(n12322), .IN2(n12330), .QN(n12333) );
  INVX0 U12184 ( .INP(n12316), .ZN(n12330) );
  NOR2X0 U12185 ( .IN1(n10739), .IN2(n11671), .QN(n12285) );
  NOR2X0 U12186 ( .IN1(n11809), .IN2(n11671), .QN(n10455) );
  NOR2X0 U12187 ( .IN1(n12335), .IN2(n12336), .QN(n12281) );
  NOR2X0 U12188 ( .IN1(n11809), .IN2(n4388), .QN(n12336) );
  NOR2X0 U12189 ( .IN1(n11171), .IN2(n12337), .QN(n12335) );
  NAND2X0 U12190 ( .IN1(n10748), .IN2(n3130), .QN(n11171) );
  NAND2X0 U12191 ( .IN1(n12338), .IN2(n12339), .QN(n10748) );
  NOR2X0 U12192 ( .IN1(n12340), .IN2(n12341), .QN(n12339) );
  NAND2X0 U12193 ( .IN1(n12329), .IN2(n12323), .QN(n12341) );
  XNOR2X1 U12194 ( .IN1(n11692), .IN2(g97), .Q(n12323) );
  INVX0 U12195 ( .INP(n4513), .ZN(n11692) );
  INVX0 U12196 ( .INP(n12320), .ZN(n12329) );
  XNOR2X1 U12197 ( .IN1(n9746), .IN2(n12342), .Q(n12320) );
  INVX0 U12198 ( .INP(n10500), .ZN(n9746) );
  NAND2X0 U12199 ( .IN1(n12343), .IN2(n12344), .QN(n10500) );
  NAND2X0 U12200 ( .IN1(g6313), .IN2(g225), .QN(n12344) );
  NOR2X0 U12201 ( .IN1(n12345), .IN2(n12346), .QN(n12343) );
  NOR2X0 U12202 ( .IN1(n8386), .IN2(n4369), .QN(n12346) );
  NOR2X0 U12203 ( .IN1(n8380), .IN2(n4318), .QN(n12345) );
  NAND2X0 U12204 ( .IN1(n12347), .IN2(n12322), .QN(n12340) );
  XNOR2X1 U12205 ( .IN1(n11636), .IN2(g121), .Q(n12322) );
  NAND2X0 U12206 ( .IN1(n12348), .IN2(n12349), .QN(n11636) );
  NAND2X0 U12207 ( .IN1(g6313), .IN2(g216), .QN(n12349) );
  NOR2X0 U12208 ( .IN1(n12350), .IN2(n12351), .QN(n12348) );
  NOR2X0 U12209 ( .IN1(n8544), .IN2(n4369), .QN(n12351) );
  NOR2X0 U12210 ( .IN1(n8473), .IN2(n4318), .QN(n12350) );
  NOR2X0 U12211 ( .IN1(n12319), .IN2(n12316), .QN(n12347) );
  XNOR2X1 U12212 ( .IN1(n11654), .IN2(g113), .Q(n12316) );
  INVX0 U12213 ( .INP(n9747), .ZN(n11654) );
  NAND2X0 U12214 ( .IN1(n12352), .IN2(n12353), .QN(n9747) );
  NAND2X0 U12215 ( .IN1(g6313), .IN2(g207), .QN(n12353) );
  NOR2X0 U12216 ( .IN1(n12354), .IN2(n12355), .QN(n12352) );
  NOR2X0 U12217 ( .IN1(n8534), .IN2(n4369), .QN(n12355) );
  NOR2X0 U12218 ( .IN1(n8477), .IN2(n4318), .QN(n12354) );
  XOR2X1 U12219 ( .IN1(n9745), .IN2(n4322), .Q(n12319) );
  INVX0 U12220 ( .INP(n11681), .ZN(n9745) );
  NAND2X0 U12221 ( .IN1(n12356), .IN2(n12357), .QN(n11681) );
  NAND2X0 U12222 ( .IN1(g6313), .IN2(g198), .QN(n12357) );
  NOR2X0 U12223 ( .IN1(n12358), .IN2(n12359), .QN(n12356) );
  NOR2X0 U12224 ( .IN1(n8545), .IN2(n4369), .QN(n12359) );
  NOR2X0 U12225 ( .IN1(n8480), .IN2(n4318), .QN(n12358) );
  NOR2X0 U12226 ( .IN1(n12360), .IN2(n12361), .QN(n12338) );
  NAND2X0 U12227 ( .IN1(n12305), .IN2(n12303), .QN(n12361) );
  INVX0 U12228 ( .INP(n12292), .ZN(n12303) );
  XNOR2X1 U12229 ( .IN1(n11653), .IN2(g117), .Q(n12292) );
  INVX0 U12230 ( .INP(n9760), .ZN(n11653) );
  NAND2X0 U12231 ( .IN1(n12362), .IN2(n12363), .QN(n9760) );
  NAND2X0 U12232 ( .IN1(g6313), .IN2(g252), .QN(n12363) );
  NOR2X0 U12233 ( .IN1(n12364), .IN2(n12365), .QN(n12362) );
  INVX0 U12234 ( .INP(n12366), .ZN(n12365) );
  NAND2X0 U12235 ( .IN1(g165), .IN2(test_so14), .QN(n12366) );
  NOR2X0 U12236 ( .IN1(n8475), .IN2(n4318), .QN(n12364) );
  INVX0 U12237 ( .INP(n12296), .ZN(n12305) );
  XNOR2X1 U12238 ( .IN1(n9759), .IN2(n12367), .Q(n12296) );
  INVX0 U12239 ( .INP(n10932), .ZN(n9759) );
  NAND2X0 U12240 ( .IN1(n12368), .IN2(n12369), .QN(n10932) );
  NAND2X0 U12241 ( .IN1(g6313), .IN2(g270), .QN(n12369) );
  NOR2X0 U12242 ( .IN1(n12370), .IN2(n12371), .QN(n12368) );
  NOR2X0 U12243 ( .IN1(n8416), .IN2(n4369), .QN(n12371) );
  NOR2X0 U12244 ( .IN1(n8415), .IN2(n4318), .QN(n12370) );
  NAND2X0 U12245 ( .IN1(n12294), .IN2(n12304), .QN(n12360) );
  INVX0 U12246 ( .INP(n12295), .ZN(n12304) );
  XNOR2X1 U12247 ( .IN1(n9754), .IN2(g109), .Q(n12295) );
  INVX0 U12248 ( .INP(n11640), .ZN(n9754) );
  NAND2X0 U12249 ( .IN1(n12372), .IN2(n12373), .QN(n11640) );
  NAND2X0 U12250 ( .IN1(g6313), .IN2(g243), .QN(n12373) );
  NOR2X0 U12251 ( .IN1(n12374), .IN2(n12375), .QN(n12372) );
  NOR2X0 U12252 ( .IN1(n8428), .IN2(n4369), .QN(n12375) );
  NOR2X0 U12253 ( .IN1(n8478), .IN2(n4318), .QN(n12374) );
  NOR2X0 U12254 ( .IN1(n12311), .IN2(n12310), .QN(n12294) );
  XOR2X1 U12255 ( .IN1(n9739), .IN2(n4376), .Q(n12310) );
  INVX0 U12256 ( .INP(n11643), .ZN(n9739) );
  NAND2X0 U12257 ( .IN1(n12376), .IN2(n12377), .QN(n11643) );
  NAND2X0 U12258 ( .IN1(g6313), .IN2(g234), .QN(n12377) );
  NOR2X0 U12259 ( .IN1(n12378), .IN2(n12379), .QN(n12376) );
  NOR2X0 U12260 ( .IN1(n8429), .IN2(n4369), .QN(n12379) );
  NOR2X0 U12261 ( .IN1(n8481), .IN2(n4318), .QN(n12378) );
  XOR2X1 U12262 ( .IN1(n9740), .IN2(g125), .Q(n12311) );
  NAND2X0 U12263 ( .IN1(n12380), .IN2(n12381), .QN(n9740) );
  NAND2X0 U12264 ( .IN1(g6313), .IN2(g261), .QN(n12381) );
  NOR2X0 U12265 ( .IN1(n12382), .IN2(n12383), .QN(n12380) );
  NOR2X0 U12266 ( .IN1(n8529), .IN2(n4369), .QN(n12383) );
  NOR2X0 U12267 ( .IN1(n8471), .IN2(n4318), .QN(n12382) );
  NOR2X0 U12268 ( .IN1(n12384), .IN2(n11820), .QN(g29112) );
  NAND2X0 U12269 ( .IN1(n2982), .IN2(n12385), .QN(n11820) );
  NAND2X0 U12270 ( .IN1(n3159), .IN2(g2129), .QN(n2982) );
  NOR2X0 U12271 ( .IN1(n3159), .IN2(g2129), .QN(n12384) );
  NOR2X0 U12272 ( .IN1(n12386), .IN2(n11825), .QN(g29111) );
  NAND2X0 U12273 ( .IN1(n2985), .IN2(n12387), .QN(n11825) );
  NAND2X0 U12274 ( .IN1(n3163), .IN2(g1435), .QN(n2985) );
  NOR2X0 U12275 ( .IN1(n3163), .IN2(g1435), .QN(n12386) );
  NOR2X0 U12276 ( .IN1(n12388), .IN2(n11830), .QN(g29110) );
  NAND2X0 U12277 ( .IN1(n2988), .IN2(n12389), .QN(n11830) );
  NAND2X0 U12278 ( .IN1(n3167), .IN2(test_so36), .QN(n2988) );
  NOR2X0 U12279 ( .IN1(n3167), .IN2(test_so36), .QN(n12388) );
  NOR2X0 U12280 ( .IN1(n12390), .IN2(n11835), .QN(g29109) );
  NAND2X0 U12281 ( .IN1(n2991), .IN2(n12391), .QN(n11835) );
  NAND2X0 U12282 ( .IN1(n3171), .IN2(g61), .QN(n2991) );
  NOR2X0 U12283 ( .IN1(n3171), .IN2(g61), .QN(n12390) );
  NAND2X0 U12284 ( .IN1(n12392), .IN2(n12393), .QN(g28788) );
  NAND2X0 U12285 ( .IN1(n12394), .IN2(g2501), .QN(n12393) );
  NAND2X0 U12286 ( .IN1(n12395), .IN2(n11841), .QN(n12394) );
  NAND2X0 U12287 ( .IN1(n12396), .IN2(n11841), .QN(n12392) );
  NAND2X0 U12288 ( .IN1(n12397), .IN2(n12398), .QN(g28783) );
  NAND2X0 U12289 ( .IN1(n12399), .IN2(g2503), .QN(n12398) );
  NAND2X0 U12290 ( .IN1(n12395), .IN2(n10669), .QN(n12399) );
  NAND2X0 U12291 ( .IN1(n12396), .IN2(n10669), .QN(n12397) );
  NAND2X0 U12292 ( .IN1(n12400), .IN2(n12401), .QN(g28782) );
  NAND2X0 U12293 ( .IN1(n4606), .IN2(n12402), .QN(n12401) );
  NAND2X0 U12294 ( .IN1(n4509), .IN2(test_so80), .QN(n12400) );
  NAND2X0 U12295 ( .IN1(n12403), .IN2(n12404), .QN(g28778) );
  NAND2X0 U12296 ( .IN1(n12405), .IN2(g1807), .QN(n12404) );
  NAND2X0 U12297 ( .IN1(n12406), .IN2(n11849), .QN(n12405) );
  NAND2X0 U12298 ( .IN1(n12407), .IN2(n11849), .QN(n12403) );
  NAND2X0 U12299 ( .IN1(n12408), .IN2(n12409), .QN(g28774) );
  NAND2X0 U12300 ( .IN1(n12410), .IN2(g2502), .QN(n12409) );
  NAND2X0 U12301 ( .IN1(n12395), .IN2(n11931), .QN(n12410) );
  NOR2X0 U12302 ( .IN1(n12411), .IN2(n11858), .QN(n12395) );
  NAND2X0 U12303 ( .IN1(n12396), .IN2(n11931), .QN(n12408) );
  NAND2X0 U12304 ( .IN1(n12412), .IN2(n12413), .QN(g28773) );
  NAND2X0 U12305 ( .IN1(g7264), .IN2(n12402), .QN(n12413) );
  INVX0 U12306 ( .INP(n12414), .ZN(n12412) );
  NOR2X0 U12307 ( .IN1(n10669), .IN2(n8703), .QN(n12414) );
  NAND2X0 U12308 ( .IN1(n12415), .IN2(n12416), .QN(g28772) );
  NAND2X0 U12309 ( .IN1(n12417), .IN2(g1809), .QN(n12416) );
  NAND2X0 U12310 ( .IN1(n12406), .IN2(n10678), .QN(n12417) );
  NAND2X0 U12311 ( .IN1(n12407), .IN2(n10678), .QN(n12415) );
  NAND2X0 U12312 ( .IN1(n12418), .IN2(n12419), .QN(g28771) );
  NAND2X0 U12313 ( .IN1(n4618), .IN2(n12420), .QN(n12419) );
  INVX0 U12314 ( .INP(n12421), .ZN(n12418) );
  NOR2X0 U12315 ( .IN1(n11849), .IN2(n8723), .QN(n12421) );
  NAND2X0 U12316 ( .IN1(n12422), .IN2(n12423), .QN(g28767) );
  NAND2X0 U12317 ( .IN1(n12424), .IN2(g1113), .QN(n12423) );
  NAND2X0 U12318 ( .IN1(n12425), .IN2(g1088), .QN(n12424) );
  NAND2X0 U12319 ( .IN1(n12426), .IN2(g1088), .QN(n12422) );
  NAND2X0 U12320 ( .IN1(n12427), .IN2(n12428), .QN(g28763) );
  NAND2X0 U12321 ( .IN1(g5555), .IN2(n12402), .QN(n12428) );
  INVX0 U12322 ( .INP(n12429), .ZN(n12402) );
  NOR2X0 U12323 ( .IN1(n12396), .IN2(n12430), .QN(n12429) );
  NOR2X0 U12324 ( .IN1(n12431), .IN2(n11860), .QN(n12430) );
  INVX0 U12325 ( .INP(n10476), .ZN(n11860) );
  NOR2X0 U12326 ( .IN1(n9281), .IN2(n12432), .QN(n12431) );
  NOR2X0 U12327 ( .IN1(n11858), .IN2(n12433), .QN(n12432) );
  INVX0 U12328 ( .INP(n12434), .ZN(n12433) );
  NAND2X0 U12329 ( .IN1(n12435), .IN2(n12436), .QN(n11858) );
  NAND2X0 U12330 ( .IN1(n8938), .IN2(n10669), .QN(n12436) );
  NOR2X0 U12331 ( .IN1(n12437), .IN2(n12438), .QN(n12435) );
  NOR2X0 U12332 ( .IN1(n4516), .IN2(g2502), .QN(n12438) );
  NOR2X0 U12333 ( .IN1(n4509), .IN2(g2501), .QN(n12437) );
  NOR2X0 U12334 ( .IN1(n12411), .IN2(n10476), .QN(n12396) );
  NAND2X0 U12335 ( .IN1(n12439), .IN2(n12440), .QN(n10476) );
  NAND2X0 U12336 ( .IN1(g5555), .IN2(g2483), .QN(n12440) );
  NOR2X0 U12337 ( .IN1(n12441), .IN2(n12442), .QN(n12439) );
  NOR2X0 U12338 ( .IN1(n8703), .IN2(n12443), .QN(n12442) );
  INVX0 U12339 ( .INP(n12444), .ZN(n12441) );
  NAND2X0 U12340 ( .IN1(n4606), .IN2(test_so80), .QN(n12444) );
  NAND2X0 U12341 ( .IN1(n12434), .IN2(test_so79), .QN(n12411) );
  NAND2X0 U12342 ( .IN1(n12445), .IN2(n12446), .QN(n12434) );
  NAND2X0 U12343 ( .IN1(n4285), .IN2(n10480), .QN(n12446) );
  NAND2X0 U12344 ( .IN1(n12447), .IN2(n11859), .QN(n12445) );
  INVX0 U12345 ( .INP(n10480), .ZN(n11859) );
  NAND2X0 U12346 ( .IN1(n12448), .IN2(n12449), .QN(n10480) );
  NOR2X0 U12347 ( .IN1(n10978), .IN2(n10796), .QN(n12448) );
  NOR2X0 U12348 ( .IN1(n11188), .IN2(n4285), .QN(n12447) );
  NOR2X0 U12349 ( .IN1(n10648), .IN2(n8988), .QN(n11188) );
  NAND2X0 U12350 ( .IN1(n12450), .IN2(n12451), .QN(n10648) );
  NAND2X0 U12351 ( .IN1(n8859), .IN2(test_so73), .QN(n12451) );
  NOR2X0 U12352 ( .IN1(n12452), .IN2(n12453), .QN(n12450) );
  NOR2X0 U12353 ( .IN1(n4367), .IN2(g2244), .QN(n12453) );
  NOR2X0 U12354 ( .IN1(n4324), .IN2(g2245), .QN(n12452) );
  NAND2X0 U12355 ( .IN1(n4516), .IN2(g2483), .QN(n12427) );
  NAND2X0 U12356 ( .IN1(n12454), .IN2(n12455), .QN(g28761) );
  NAND2X0 U12357 ( .IN1(n12456), .IN2(g1808), .QN(n12455) );
  NAND2X0 U12358 ( .IN1(n12406), .IN2(n12050), .QN(n12456) );
  NOR2X0 U12359 ( .IN1(n12457), .IN2(n11878), .QN(n12406) );
  NAND2X0 U12360 ( .IN1(n12407), .IN2(n12050), .QN(n12454) );
  NAND2X0 U12361 ( .IN1(n12458), .IN2(n12459), .QN(g28760) );
  NAND2X0 U12362 ( .IN1(g7014), .IN2(n12420), .QN(n12459) );
  INVX0 U12363 ( .INP(n12460), .ZN(n12458) );
  NOR2X0 U12364 ( .IN1(n10678), .IN2(n8707), .QN(n12460) );
  NAND2X0 U12365 ( .IN1(n12461), .IN2(n12462), .QN(g28759) );
  NAND2X0 U12366 ( .IN1(n12463), .IN2(g1115), .QN(n12462) );
  NAND2X0 U12367 ( .IN1(n12425), .IN2(g6712), .QN(n12463) );
  NAND2X0 U12368 ( .IN1(n12426), .IN2(g6712), .QN(n12461) );
  NAND2X0 U12369 ( .IN1(n12464), .IN2(n12465), .QN(g28758) );
  NAND2X0 U12370 ( .IN1(n4381), .IN2(g1101), .QN(n12465) );
  NAND2X0 U12371 ( .IN1(n12466), .IN2(g1088), .QN(n12464) );
  NAND2X0 U12372 ( .IN1(n12467), .IN2(n12468), .QN(g28754) );
  NAND2X0 U12373 ( .IN1(n12469), .IN2(g426), .QN(n12468) );
  NAND2X0 U12374 ( .IN1(n12470), .IN2(n11886), .QN(n12469) );
  NAND2X0 U12375 ( .IN1(n12471), .IN2(n11886), .QN(n12467) );
  NAND2X0 U12376 ( .IN1(n12472), .IN2(n12473), .QN(g28749) );
  NAND2X0 U12377 ( .IN1(g5511), .IN2(n12420), .QN(n12473) );
  NAND2X0 U12378 ( .IN1(n12474), .IN2(n12475), .QN(n12420) );
  NAND2X0 U12379 ( .IN1(n12476), .IN2(n10472), .QN(n12475) );
  NAND2X0 U12380 ( .IN1(g1690), .IN2(n12477), .QN(n12476) );
  NAND2X0 U12381 ( .IN1(n12478), .IN2(n12479), .QN(n12477) );
  INVX0 U12382 ( .INP(n11878), .ZN(n12478) );
  NAND2X0 U12383 ( .IN1(n12480), .IN2(n12481), .QN(n11878) );
  NAND2X0 U12384 ( .IN1(n8941), .IN2(n10678), .QN(n12481) );
  NOR2X0 U12385 ( .IN1(n12482), .IN2(n12483), .QN(n12480) );
  NOR2X0 U12386 ( .IN1(n4518), .IN2(g1808), .QN(n12483) );
  NOR2X0 U12387 ( .IN1(n4511), .IN2(g1807), .QN(n12482) );
  INVX0 U12388 ( .INP(n12407), .ZN(n12474) );
  NOR2X0 U12389 ( .IN1(n12457), .IN2(n10472), .QN(n12407) );
  NAND2X0 U12390 ( .IN1(n12484), .IN2(n12485), .QN(n10472) );
  NAND2X0 U12391 ( .IN1(g5511), .IN2(g1789), .QN(n12485) );
  NOR2X0 U12392 ( .IN1(n12486), .IN2(n12487), .QN(n12484) );
  NOR2X0 U12393 ( .IN1(n8707), .IN2(n11731), .QN(n12487) );
  NOR2X0 U12394 ( .IN1(n8723), .IN2(n12488), .QN(n12486) );
  NAND2X0 U12395 ( .IN1(g1690), .IN2(n12479), .QN(n12457) );
  NAND2X0 U12396 ( .IN1(n12489), .IN2(n12490), .QN(n12479) );
  NAND2X0 U12397 ( .IN1(n4284), .IN2(n10473), .QN(n12490) );
  NAND2X0 U12398 ( .IN1(n12491), .IN2(n12492), .QN(n12489) );
  INVX0 U12399 ( .INP(n10473), .ZN(n12492) );
  NAND2X0 U12400 ( .IN1(n12493), .IN2(n12494), .QN(n10473) );
  NOR2X0 U12401 ( .IN1(n11025), .IN2(n10835), .QN(n12493) );
  NOR2X0 U12402 ( .IN1(n10694), .IN2(n4284), .QN(n12491) );
  NOR2X0 U12403 ( .IN1(n9667), .IN2(n8989), .QN(n10694) );
  NAND2X0 U12404 ( .IN1(n12495), .IN2(n12496), .QN(n9667) );
  NAND2X0 U12405 ( .IN1(n8870), .IN2(g6782), .QN(n12496) );
  NOR2X0 U12406 ( .IN1(n12497), .IN2(n12498), .QN(n12495) );
  NOR2X0 U12407 ( .IN1(n4368), .IN2(g1550), .QN(n12498) );
  NOR2X0 U12408 ( .IN1(n4317), .IN2(g1551), .QN(n12497) );
  NAND2X0 U12409 ( .IN1(n4518), .IN2(g1789), .QN(n12472) );
  NAND2X0 U12410 ( .IN1(n12499), .IN2(n12500), .QN(g28747) );
  NAND2X0 U12411 ( .IN1(n12501), .IN2(g1114), .QN(n12500) );
  NAND2X0 U12412 ( .IN1(n12425), .IN2(g5472), .QN(n12501) );
  NOR2X0 U12413 ( .IN1(n12502), .IN2(n11896), .QN(n12425) );
  NAND2X0 U12414 ( .IN1(n12426), .IN2(g5472), .QN(n12499) );
  NAND2X0 U12415 ( .IN1(n12503), .IN2(n12504), .QN(g28746) );
  INVX0 U12416 ( .INP(n12505), .ZN(n12504) );
  NOR2X0 U12417 ( .IN1(g6712), .IN2(n8710), .QN(n12505) );
  NAND2X0 U12418 ( .IN1(n12466), .IN2(g6712), .QN(n12503) );
  NAND2X0 U12419 ( .IN1(n12506), .IN2(n12507), .QN(g28745) );
  NAND2X0 U12420 ( .IN1(n12508), .IN2(g428), .QN(n12507) );
  NAND2X0 U12421 ( .IN1(n12470), .IN2(n11905), .QN(n12508) );
  NAND2X0 U12422 ( .IN1(n12471), .IN2(n11905), .QN(n12506) );
  NAND2X0 U12423 ( .IN1(n12509), .IN2(n12510), .QN(g28744) );
  NAND2X0 U12424 ( .IN1(n4640), .IN2(n12511), .QN(n12510) );
  INVX0 U12425 ( .INP(n12512), .ZN(n12509) );
  NOR2X0 U12426 ( .IN1(n11886), .IN2(n8742), .QN(n12512) );
  NAND2X0 U12427 ( .IN1(n12513), .IN2(n12514), .QN(g28738) );
  INVX0 U12428 ( .INP(n12515), .ZN(n12514) );
  NOR2X0 U12429 ( .IN1(g5472), .IN2(n8732), .QN(n12515) );
  NAND2X0 U12430 ( .IN1(n12466), .IN2(g5472), .QN(n12513) );
  INVX0 U12431 ( .INP(n12516), .ZN(n12466) );
  NOR2X0 U12432 ( .IN1(n12426), .IN2(n12517), .QN(n12516) );
  NOR2X0 U12433 ( .IN1(n12518), .IN2(n11898), .QN(n12517) );
  INVX0 U12434 ( .INP(n10464), .ZN(n11898) );
  NOR2X0 U12435 ( .IN1(n4387), .IN2(n12519), .QN(n12518) );
  NOR2X0 U12436 ( .IN1(n11896), .IN2(n12520), .QN(n12519) );
  INVX0 U12437 ( .INP(n12521), .ZN(n12520) );
  NAND2X0 U12438 ( .IN1(n12522), .IN2(n12523), .QN(n11896) );
  NAND2X0 U12439 ( .IN1(n8958), .IN2(g1088), .QN(n12523) );
  NOR2X0 U12440 ( .IN1(n12524), .IN2(n12525), .QN(n12522) );
  NOR2X0 U12441 ( .IN1(n4364), .IN2(g1115), .QN(n12525) );
  NOR2X0 U12442 ( .IN1(n4363), .IN2(g1114), .QN(n12524) );
  NOR2X0 U12443 ( .IN1(n12502), .IN2(n10464), .QN(n12426) );
  NAND2X0 U12444 ( .IN1(n12526), .IN2(n12527), .QN(n10464) );
  NAND2X0 U12445 ( .IN1(g1088), .IN2(g1101), .QN(n12527) );
  NOR2X0 U12446 ( .IN1(n12528), .IN2(n12529), .QN(n12526) );
  NOR2X0 U12447 ( .IN1(n8710), .IN2(n4364), .QN(n12529) );
  NOR2X0 U12448 ( .IN1(n8732), .IN2(n4363), .QN(n12528) );
  NAND2X0 U12449 ( .IN1(g996), .IN2(n12521), .QN(n12502) );
  NAND2X0 U12450 ( .IN1(n12530), .IN2(n12531), .QN(n12521) );
  NAND2X0 U12451 ( .IN1(n4283), .IN2(n10468), .QN(n12531) );
  NAND2X0 U12452 ( .IN1(n12532), .IN2(n11897), .QN(n12530) );
  INVX0 U12453 ( .INP(n10468), .ZN(n11897) );
  NAND2X0 U12454 ( .IN1(n12533), .IN2(n12534), .QN(n10468) );
  NOR2X0 U12455 ( .IN1(n11066), .IN2(n10876), .QN(n12533) );
  NOR2X0 U12456 ( .IN1(n10516), .IN2(n4283), .QN(n12532) );
  NOR2X0 U12457 ( .IN1(n9680), .IN2(n8990), .QN(n10516) );
  NAND2X0 U12458 ( .IN1(n12535), .IN2(n12536), .QN(n9680) );
  NAND2X0 U12459 ( .IN1(test_so31), .IN2(n8881), .QN(n12536) );
  NOR2X0 U12460 ( .IN1(n12537), .IN2(n12538), .QN(n12535) );
  NOR2X0 U12461 ( .IN1(n4323), .IN2(g857), .QN(n12538) );
  NOR2X0 U12462 ( .IN1(test_so33), .IN2(n4312), .QN(n12537) );
  NAND2X0 U12463 ( .IN1(n12539), .IN2(n12540), .QN(g28736) );
  NAND2X0 U12464 ( .IN1(test_so17), .IN2(n12541), .QN(n12540) );
  NAND2X0 U12465 ( .IN1(n12470), .IN2(n10752), .QN(n12541) );
  NOR2X0 U12466 ( .IN1(n12542), .IN2(n11914), .QN(n12470) );
  NAND2X0 U12467 ( .IN1(n12471), .IN2(n10752), .QN(n12539) );
  NAND2X0 U12468 ( .IN1(n12543), .IN2(n12544), .QN(g28735) );
  NAND2X0 U12469 ( .IN1(g6447), .IN2(n12511), .QN(n12544) );
  INVX0 U12470 ( .INP(n12545), .ZN(n12543) );
  NOR2X0 U12471 ( .IN1(n11905), .IN2(n8743), .QN(n12545) );
  NAND2X0 U12472 ( .IN1(n12546), .IN2(n12547), .QN(g28732) );
  NAND2X0 U12473 ( .IN1(g5437), .IN2(n12511), .QN(n12547) );
  NAND2X0 U12474 ( .IN1(n12548), .IN2(n12549), .QN(n12511) );
  NAND2X0 U12475 ( .IN1(n12550), .IN2(n10460), .QN(n12549) );
  NAND2X0 U12476 ( .IN1(g309), .IN2(n12551), .QN(n12550) );
  NAND2X0 U12477 ( .IN1(n12552), .IN2(n12553), .QN(n12551) );
  INVX0 U12478 ( .INP(n11914), .ZN(n12552) );
  NAND2X0 U12479 ( .IN1(n12554), .IN2(n12555), .QN(n11914) );
  NAND2X0 U12480 ( .IN1(n10752), .IN2(n9289), .QN(n12555) );
  NOR2X0 U12481 ( .IN1(n12556), .IN2(n12557), .QN(n12554) );
  NOR2X0 U12482 ( .IN1(n4506), .IN2(g426), .QN(n12557) );
  NOR2X0 U12483 ( .IN1(n4499), .IN2(g428), .QN(n12556) );
  INVX0 U12484 ( .INP(n12471), .ZN(n12548) );
  NOR2X0 U12485 ( .IN1(n12542), .IN2(n10460), .QN(n12471) );
  NAND2X0 U12486 ( .IN1(n12558), .IN2(n12559), .QN(n10460) );
  NAND2X0 U12487 ( .IN1(g5437), .IN2(g408), .QN(n12559) );
  NOR2X0 U12488 ( .IN1(n12560), .IN2(n12561), .QN(n12558) );
  NOR2X0 U12489 ( .IN1(n8743), .IN2(n12562), .QN(n12561) );
  NOR2X0 U12490 ( .IN1(n8742), .IN2(n12563), .QN(n12560) );
  NAND2X0 U12491 ( .IN1(g309), .IN2(n12553), .QN(n12542) );
  NAND2X0 U12492 ( .IN1(n12564), .IN2(n12565), .QN(n12553) );
  NAND2X0 U12493 ( .IN1(n4282), .IN2(n10461), .QN(n12565) );
  NAND2X0 U12494 ( .IN1(n12566), .IN2(n12567), .QN(n12564) );
  INVX0 U12495 ( .INP(n10461), .ZN(n12567) );
  NAND2X0 U12496 ( .IN1(n12568), .IN2(n12569), .QN(n10461) );
  NOR2X0 U12497 ( .IN1(n11093), .IN2(n10928), .QN(n12568) );
  NOR2X0 U12498 ( .IN1(n10733), .IN2(n4282), .QN(n12566) );
  NOR2X0 U12499 ( .IN1(n10449), .IN2(n8991), .QN(n10733) );
  NAND2X0 U12500 ( .IN1(n12570), .IN2(n12571), .QN(n10449) );
  NAND2X0 U12501 ( .IN1(n8893), .IN2(g6313), .QN(n12571) );
  NOR2X0 U12502 ( .IN1(n12572), .IN2(n12573), .QN(n12570) );
  NOR2X0 U12503 ( .IN1(n4369), .IN2(g168), .QN(n12573) );
  NOR2X0 U12504 ( .IN1(n4318), .IN2(g169), .QN(n12572) );
  NAND2X0 U12505 ( .IN1(n4520), .IN2(g408), .QN(n12546) );
  NOR2X0 U12506 ( .IN1(n9684), .IN2(n12574), .QN(g28668) );
  XOR2X1 U12507 ( .IN1(n4418), .IN2(n9685), .Q(n12574) );
  NOR2X0 U12508 ( .IN1(n9686), .IN2(n4396), .QN(n9685) );
  NAND2X0 U12509 ( .IN1(n12575), .IN2(n12576), .QN(g28637) );
  INVX0 U12510 ( .INP(n12577), .ZN(n12576) );
  NOR2X0 U12511 ( .IN1(n12578), .IN2(n8969), .QN(n12577) );
  NAND2X0 U12512 ( .IN1(n12579), .IN2(n8969), .QN(n12575) );
  NOR2X0 U12513 ( .IN1(n9702), .IN2(n3160), .QN(n12579) );
  NAND2X0 U12514 ( .IN1(n12580), .IN2(n12581), .QN(g28636) );
  INVX0 U12515 ( .INP(n12582), .ZN(n12581) );
  NOR2X0 U12516 ( .IN1(n12583), .IN2(n8973), .QN(n12582) );
  NAND2X0 U12517 ( .IN1(n12584), .IN2(n8973), .QN(n12580) );
  NOR2X0 U12518 ( .IN1(n9710), .IN2(n3164), .QN(n12584) );
  NAND2X0 U12519 ( .IN1(n12585), .IN2(n12586), .QN(g28635) );
  INVX0 U12520 ( .INP(n12587), .ZN(n12586) );
  NOR2X0 U12521 ( .IN1(n12588), .IN2(n8977), .QN(n12587) );
  NAND2X0 U12522 ( .IN1(n12589), .IN2(n8977), .QN(n12585) );
  NOR2X0 U12523 ( .IN1(n11814), .IN2(n3168), .QN(n12589) );
  NAND2X0 U12524 ( .IN1(n12590), .IN2(n12591), .QN(g28634) );
  INVX0 U12525 ( .INP(n12592), .ZN(n12591) );
  NOR2X0 U12526 ( .IN1(n12593), .IN2(n8981), .QN(n12592) );
  NAND2X0 U12527 ( .IN1(n12594), .IN2(n8981), .QN(n12590) );
  NOR2X0 U12528 ( .IN1(n9719), .IN2(n3172), .QN(n12594) );
  NAND2X0 U12529 ( .IN1(n12595), .IN2(n12596), .QN(g28425) );
  INVX0 U12530 ( .INP(n12597), .ZN(n12596) );
  NOR2X0 U12531 ( .IN1(g3109), .IN2(n4343), .QN(n12597) );
  NAND2X0 U12532 ( .IN1(n521), .IN2(g3109), .QN(n12595) );
  NAND2X0 U12533 ( .IN1(n12598), .IN2(n12599), .QN(g28421) );
  NAND2X0 U12534 ( .IN1(n4383), .IN2(test_so7), .QN(n12599) );
  NAND2X0 U12535 ( .IN1(n521), .IN2(g8030), .QN(n12598) );
  NAND2X0 U12536 ( .IN1(n12600), .IN2(n12601), .QN(g28420) );
  INVX0 U12537 ( .INP(n12602), .ZN(n12601) );
  NOR2X0 U12538 ( .IN1(g8106), .IN2(n4342), .QN(n12602) );
  NAND2X0 U12539 ( .IN1(n521), .IN2(g8106), .QN(n12600) );
  INVX0 U12540 ( .INP(n11752), .ZN(n521) );
  NAND2X0 U12541 ( .IN1(n12603), .IN2(n12604), .QN(n11752) );
  NAND2X0 U12542 ( .IN1(n8373), .IN2(g1186), .QN(n12604) );
  NAND2X0 U12543 ( .IN1(n12605), .IN2(n4548), .QN(n12603) );
  NOR2X0 U12544 ( .IN1(n12606), .IN2(n12607), .QN(n12605) );
  NOR2X0 U12545 ( .IN1(n8374), .IN2(n12608), .QN(n12607) );
  INVX0 U12546 ( .INP(n12609), .ZN(n12606) );
  NAND2X0 U12547 ( .IN1(g21851), .IN2(g6750), .QN(n12609) );
  NAND2X0 U12548 ( .IN1(n12610), .IN2(n12611), .QN(g28371) );
  INVX0 U12549 ( .INP(n12612), .ZN(n12611) );
  NOR2X0 U12550 ( .IN1(g2624), .IN2(n8679), .QN(n12612) );
  NAND2X0 U12551 ( .IN1(n12613), .IN2(g2624), .QN(n12610) );
  NAND2X0 U12552 ( .IN1(n12614), .IN2(n12615), .QN(g28368) );
  NAND2X0 U12553 ( .IN1(n4370), .IN2(g2691), .QN(n12615) );
  NAND2X0 U12554 ( .IN1(n12613), .IN2(g7390), .QN(n12614) );
  NAND2X0 U12555 ( .IN1(n12616), .IN2(n12617), .QN(g28367) );
  INVX0 U12556 ( .INP(n12618), .ZN(n12617) );
  NOR2X0 U12557 ( .IN1(g2624), .IN2(n8688), .QN(n12618) );
  NAND2X0 U12558 ( .IN1(n12619), .IN2(g2624), .QN(n12616) );
  NAND2X0 U12559 ( .IN1(n12620), .IN2(n12621), .QN(g28366) );
  NAND2X0 U12560 ( .IN1(n4366), .IN2(g2000), .QN(n12621) );
  NAND2X0 U12561 ( .IN1(n12622), .IN2(g1930), .QN(n12620) );
  NAND2X0 U12562 ( .IN1(n12623), .IN2(n12624), .QN(g28364) );
  INVX0 U12563 ( .INP(n12625), .ZN(n12624) );
  NOR2X0 U12564 ( .IN1(n11699), .IN2(n8678), .QN(n12625) );
  NAND2X0 U12565 ( .IN1(n12613), .IN2(n11699), .QN(n12623) );
  NAND2X0 U12566 ( .IN1(n12626), .IN2(n12627), .QN(n12613) );
  NAND2X0 U12567 ( .IN1(n3252), .IN2(n12628), .QN(n12627) );
  NAND2X0 U12568 ( .IN1(n10153), .IN2(n12629), .QN(n12626) );
  NAND2X0 U12569 ( .IN1(n12630), .IN2(n12631), .QN(g28363) );
  NAND2X0 U12570 ( .IN1(n12619), .IN2(g7390), .QN(n12631) );
  NAND2X0 U12571 ( .IN1(n4370), .IN2(test_so90), .QN(n12630) );
  NAND2X0 U12572 ( .IN1(n12632), .IN2(n12633), .QN(g28362) );
  INVX0 U12573 ( .INP(n12634), .ZN(n12633) );
  NOR2X0 U12574 ( .IN1(g7194), .IN2(n8683), .QN(n12634) );
  NAND2X0 U12575 ( .IN1(n12622), .IN2(g7194), .QN(n12632) );
  NAND2X0 U12576 ( .IN1(n12635), .IN2(n12636), .QN(g28361) );
  NAND2X0 U12577 ( .IN1(n4366), .IN2(g1991), .QN(n12636) );
  NAND2X0 U12578 ( .IN1(n12637), .IN2(g1930), .QN(n12635) );
  NAND2X0 U12579 ( .IN1(n12638), .IN2(n12639), .QN(g28360) );
  INVX0 U12580 ( .INP(n12640), .ZN(n12639) );
  NOR2X0 U12581 ( .IN1(g1236), .IN2(n8685), .QN(n12640) );
  NAND2X0 U12582 ( .IN1(n12641), .IN2(g1236), .QN(n12638) );
  NAND2X0 U12583 ( .IN1(n12642), .IN2(n12643), .QN(g28358) );
  NAND2X0 U12584 ( .IN1(g7302), .IN2(n12619), .QN(n12643) );
  NAND2X0 U12585 ( .IN1(n12644), .IN2(n12645), .QN(n12619) );
  NAND2X0 U12586 ( .IN1(n10628), .IN2(n12629), .QN(n12645) );
  NAND2X0 U12587 ( .IN1(n12646), .IN2(n12628), .QN(n12644) );
  NOR2X0 U12588 ( .IN1(n12647), .IN2(n10454), .QN(n12646) );
  NAND2X0 U12589 ( .IN1(n12648), .IN2(n12649), .QN(n10454) );
  NOR2X0 U12590 ( .IN1(n12650), .IN2(n12651), .QN(n12649) );
  NOR2X0 U12591 ( .IN1(n12652), .IN2(n12653), .QN(n12651) );
  NAND2X0 U12592 ( .IN1(n12654), .IN2(n12655), .QN(n12653) );
  NAND2X0 U12593 ( .IN1(n12656), .IN2(n12657), .QN(n12655) );
  NAND2X0 U12594 ( .IN1(n12658), .IN2(n12659), .QN(n12657) );
  NOR2X0 U12595 ( .IN1(n12660), .IN2(n12661), .QN(n12650) );
  NOR2X0 U12596 ( .IN1(n12662), .IN2(n12663), .QN(n12660) );
  INVX0 U12597 ( .INP(n12664), .ZN(n12663) );
  NAND2X0 U12598 ( .IN1(n12658), .IN2(n12665), .QN(n12664) );
  NAND2X0 U12599 ( .IN1(n12666), .IN2(n12667), .QN(n12658) );
  NAND2X0 U12600 ( .IN1(n12668), .IN2(n12669), .QN(n12667) );
  NOR2X0 U12601 ( .IN1(n12656), .IN2(n12670), .QN(n12662) );
  INVX0 U12602 ( .INP(n12671), .ZN(n12656) );
  NAND2X0 U12603 ( .IN1(n12672), .IN2(n12673), .QN(n12671) );
  NAND2X0 U12604 ( .IN1(n12674), .IN2(n12675), .QN(n12673) );
  NAND2X0 U12605 ( .IN1(n12676), .IN2(n12669), .QN(n12672) );
  NOR2X0 U12606 ( .IN1(n12677), .IN2(n12678), .QN(n12648) );
  NOR2X0 U12607 ( .IN1(n12675), .IN2(n12679), .QN(n12678) );
  NAND2X0 U12608 ( .IN1(n12680), .IN2(n12681), .QN(n12679) );
  NAND2X0 U12609 ( .IN1(n12682), .IN2(n12683), .QN(n12680) );
  NAND2X0 U12610 ( .IN1(n12684), .IN2(n12685), .QN(n12683) );
  NAND2X0 U12611 ( .IN1(n12654), .IN2(n12676), .QN(n12685) );
  NOR2X0 U12612 ( .IN1(n12686), .IN2(n12669), .QN(n12677) );
  NOR2X0 U12613 ( .IN1(n12687), .IN2(n12688), .QN(n12686) );
  NOR2X0 U12614 ( .IN1(n12668), .IN2(n12689), .QN(n12688) );
  NOR2X0 U12615 ( .IN1(n12690), .IN2(n12684), .QN(n12689) );
  NOR2X0 U12616 ( .IN1(n12652), .IN2(n12665), .QN(n12690) );
  NOR2X0 U12617 ( .IN1(n12691), .IN2(n12692), .QN(n12687) );
  NAND2X0 U12618 ( .IN1(n12684), .IN2(n12674), .QN(n12692) );
  NAND2X0 U12619 ( .IN1(n12666), .IN2(n12693), .QN(n12691) );
  NAND2X0 U12620 ( .IN1(n12694), .IN2(n10451), .QN(n12647) );
  NAND2X0 U12621 ( .IN1(n10453), .IN2(n12695), .QN(n10451) );
  NAND2X0 U12622 ( .IN1(n1421), .IN2(n12696), .QN(n12694) );
  INVX0 U12623 ( .INP(n12697), .ZN(n1421) );
  NAND2X0 U12624 ( .IN1(n12698), .IN2(n12699), .QN(n12697) );
  NAND2X0 U12625 ( .IN1(n12700), .IN2(n12661), .QN(n12699) );
  NAND2X0 U12626 ( .IN1(n12701), .IN2(n12702), .QN(n12700) );
  NAND2X0 U12627 ( .IN1(n12703), .IN2(n12665), .QN(n12702) );
  NAND2X0 U12628 ( .IN1(n12675), .IN2(n12704), .QN(n12701) );
  NAND2X0 U12629 ( .IN1(n12705), .IN2(n12706), .QN(n12704) );
  NAND2X0 U12630 ( .IN1(n12684), .IN2(n12681), .QN(n12706) );
  NOR2X0 U12631 ( .IN1(n12707), .IN2(n12708), .QN(n12705) );
  NOR2X0 U12632 ( .IN1(n12670), .IN2(n12709), .QN(n12708) );
  INVX0 U12633 ( .INP(n12710), .ZN(n12709) );
  NOR2X0 U12634 ( .IN1(n12665), .IN2(n12711), .QN(n12707) );
  NAND2X0 U12635 ( .IN1(n12676), .IN2(n12693), .QN(n12711) );
  NOR2X0 U12636 ( .IN1(n12712), .IN2(n12713), .QN(n12698) );
  NOR2X0 U12637 ( .IN1(n12675), .IN2(n12714), .QN(n12713) );
  NOR2X0 U12638 ( .IN1(n12715), .IN2(n12716), .QN(n12714) );
  NOR2X0 U12639 ( .IN1(n12717), .IN2(n12661), .QN(n12716) );
  NOR2X0 U12640 ( .IN1(n12718), .IN2(n12719), .QN(n12717) );
  NAND2X0 U12641 ( .IN1(n12720), .IN2(n12721), .QN(n12719) );
  NAND2X0 U12642 ( .IN1(n12710), .IN2(n12684), .QN(n12721) );
  INVX0 U12643 ( .INP(n12659), .ZN(n12684) );
  INVX0 U12644 ( .INP(n12722), .ZN(n12720) );
  NOR2X0 U12645 ( .IN1(n12682), .IN2(n12681), .QN(n12722) );
  NAND2X0 U12646 ( .IN1(n12723), .IN2(n12666), .QN(n12682) );
  NOR2X0 U12647 ( .IN1(n12654), .IN2(n12665), .QN(n12723) );
  INVX0 U12648 ( .INP(n12724), .ZN(n12665) );
  NAND2X0 U12649 ( .IN1(n12725), .IN2(n12726), .QN(n12724) );
  NAND2X0 U12650 ( .IN1(test_so85), .IN2(g2412), .QN(n12726) );
  NOR2X0 U12651 ( .IN1(n12727), .IN2(n12728), .QN(n12725) );
  NOR2X0 U12652 ( .IN1(n16821), .IN2(n8610), .QN(n12728) );
  NOR2X0 U12653 ( .IN1(n8613), .IN2(n8411), .QN(n12727) );
  INVX0 U12654 ( .INP(n12693), .ZN(n12654) );
  NOR2X0 U12655 ( .IN1(n12666), .IN2(n12693), .QN(n12718) );
  NOR2X0 U12656 ( .IN1(n12668), .IN2(n12670), .QN(n12715) );
  NAND2X0 U12657 ( .IN1(n12659), .IN2(n12693), .QN(n12670) );
  NOR2X0 U12658 ( .IN1(n12693), .IN2(n12729), .QN(n12712) );
  NAND2X0 U12659 ( .IN1(n12730), .IN2(n12681), .QN(n12729) );
  NAND2X0 U12660 ( .IN1(n12731), .IN2(n12732), .QN(n12730) );
  NAND2X0 U12661 ( .IN1(n12675), .IN2(n12666), .QN(n12732) );
  INVX0 U12662 ( .INP(n12669), .ZN(n12675) );
  NAND2X0 U12663 ( .IN1(n12733), .IN2(n12734), .QN(n12669) );
  NAND2X0 U12664 ( .IN1(g5796), .IN2(g2426), .QN(n12734) );
  NOR2X0 U12665 ( .IN1(n12735), .IN2(n12736), .QN(n12733) );
  NOR2X0 U12666 ( .IN1(n8612), .IN2(n8611), .QN(n12736) );
  NOR2X0 U12667 ( .IN1(n16820), .IN2(n8610), .QN(n12735) );
  NAND2X0 U12668 ( .IN1(n12652), .IN2(n12659), .QN(n12731) );
  NAND2X0 U12669 ( .IN1(n12737), .IN2(n12738), .QN(n12659) );
  NAND2X0 U12670 ( .IN1(g5747), .IN2(g2454), .QN(n12738) );
  NOR2X0 U12671 ( .IN1(n12739), .IN2(n12740), .QN(n12737) );
  NOR2X0 U12672 ( .IN1(n8613), .IN2(n8577), .QN(n12740) );
  NOR2X0 U12673 ( .IN1(n8611), .IN2(n8576), .QN(n12739) );
  NAND2X0 U12674 ( .IN1(n12741), .IN2(n12742), .QN(n12693) );
  NAND2X0 U12675 ( .IN1(g5747), .IN2(g2439), .QN(n12742) );
  NOR2X0 U12676 ( .IN1(n12743), .IN2(n12744), .QN(n12741) );
  NOR2X0 U12677 ( .IN1(n8613), .IN2(n8403), .QN(n12744) );
  NOR2X0 U12678 ( .IN1(n8611), .IN2(n8402), .QN(n12743) );
  INVX0 U12679 ( .INP(n12745), .ZN(n12642) );
  NOR2X0 U12680 ( .IN1(n11699), .IN2(n8687), .QN(n12745) );
  NAND2X0 U12681 ( .IN1(n12746), .IN2(n12747), .QN(g28357) );
  INVX0 U12682 ( .INP(n12748), .ZN(n12747) );
  NOR2X0 U12683 ( .IN1(n12749), .IN2(n8681), .QN(n12748) );
  NAND2X0 U12684 ( .IN1(n12622), .IN2(n12749), .QN(n12746) );
  NAND2X0 U12685 ( .IN1(n12750), .IN2(n12751), .QN(n12622) );
  NAND2X0 U12686 ( .IN1(n10293), .IN2(n12629), .QN(n12751) );
  NAND2X0 U12687 ( .IN1(n12752), .IN2(n12628), .QN(n12750) );
  NOR2X0 U12688 ( .IN1(n12753), .IN2(n12754), .QN(n12752) );
  NAND2X0 U12689 ( .IN1(n12755), .IN2(n12756), .QN(n12753) );
  INVX0 U12690 ( .INP(n12757), .ZN(n12755) );
  NOR2X0 U12691 ( .IN1(n12758), .IN2(n12759), .QN(n12757) );
  NAND2X0 U12692 ( .IN1(n12760), .IN2(n12761), .QN(g28356) );
  INVX0 U12693 ( .INP(n12762), .ZN(n12761) );
  NOR2X0 U12694 ( .IN1(g7194), .IN2(n8691), .QN(n12762) );
  NAND2X0 U12695 ( .IN1(n12637), .IN2(g7194), .QN(n12760) );
  NAND2X0 U12696 ( .IN1(n12763), .IN2(n12764), .QN(g28355) );
  INVX0 U12697 ( .INP(n12765), .ZN(n12764) );
  NOR2X0 U12698 ( .IN1(g6944), .IN2(n8686), .QN(n12765) );
  NAND2X0 U12699 ( .IN1(n12641), .IN2(g6944), .QN(n12763) );
  NAND2X0 U12700 ( .IN1(n12766), .IN2(n12767), .QN(g28354) );
  INVX0 U12701 ( .INP(n12768), .ZN(n12767) );
  NOR2X0 U12702 ( .IN1(g1236), .IN2(n8693), .QN(n12768) );
  NAND2X0 U12703 ( .IN1(n12769), .IN2(g1236), .QN(n12766) );
  NAND2X0 U12704 ( .IN1(n12770), .IN2(n12771), .QN(g28353) );
  NAND2X0 U12705 ( .IN1(n12772), .IN2(g550), .QN(n12771) );
  NAND2X0 U12706 ( .IN1(test_so26), .IN2(n4313), .QN(n12770) );
  NAND2X0 U12707 ( .IN1(n12773), .IN2(n12774), .QN(g28352) );
  NAND2X0 U12708 ( .IN1(g7052), .IN2(n12637), .QN(n12774) );
  NAND2X0 U12709 ( .IN1(n12775), .IN2(n12776), .QN(n12637) );
  NAND2X0 U12710 ( .IN1(n10266), .IN2(n12629), .QN(n12776) );
  NAND2X0 U12711 ( .IN1(n12777), .IN2(n12628), .QN(n12775) );
  NOR2X0 U12712 ( .IN1(n12778), .IN2(n12759), .QN(n12777) );
  NAND2X0 U12713 ( .IN1(n12779), .IN2(n12780), .QN(n12759) );
  NOR2X0 U12714 ( .IN1(n12781), .IN2(n12782), .QN(n12780) );
  NOR2X0 U12715 ( .IN1(n12783), .IN2(n12784), .QN(n12782) );
  NAND2X0 U12716 ( .IN1(n12785), .IN2(n12786), .QN(n12784) );
  NAND2X0 U12717 ( .IN1(n12787), .IN2(n12788), .QN(n12786) );
  NAND2X0 U12718 ( .IN1(n12789), .IN2(n12790), .QN(n12788) );
  NOR2X0 U12719 ( .IN1(n12791), .IN2(n12792), .QN(n12781) );
  NOR2X0 U12720 ( .IN1(n12793), .IN2(n12794), .QN(n12791) );
  INVX0 U12721 ( .INP(n12795), .ZN(n12794) );
  NAND2X0 U12722 ( .IN1(n12789), .IN2(n12796), .QN(n12795) );
  NAND2X0 U12723 ( .IN1(n12797), .IN2(n12798), .QN(n12789) );
  NAND2X0 U12724 ( .IN1(n12799), .IN2(n12800), .QN(n12798) );
  NOR2X0 U12725 ( .IN1(n12787), .IN2(n12801), .QN(n12793) );
  INVX0 U12726 ( .INP(n12802), .ZN(n12787) );
  NAND2X0 U12727 ( .IN1(n12803), .IN2(n12804), .QN(n12802) );
  NAND2X0 U12728 ( .IN1(n12805), .IN2(n12806), .QN(n12804) );
  NAND2X0 U12729 ( .IN1(n12807), .IN2(n12800), .QN(n12803) );
  NOR2X0 U12730 ( .IN1(n12808), .IN2(n12809), .QN(n12779) );
  NOR2X0 U12731 ( .IN1(n12806), .IN2(n12810), .QN(n12809) );
  NAND2X0 U12732 ( .IN1(n12811), .IN2(n12812), .QN(n12810) );
  NAND2X0 U12733 ( .IN1(n12813), .IN2(n12814), .QN(n12811) );
  NAND2X0 U12734 ( .IN1(n12815), .IN2(n12816), .QN(n12814) );
  NAND2X0 U12735 ( .IN1(n12785), .IN2(n12807), .QN(n12816) );
  NOR2X0 U12736 ( .IN1(n12817), .IN2(n12800), .QN(n12808) );
  NOR2X0 U12737 ( .IN1(n12818), .IN2(n12819), .QN(n12817) );
  NOR2X0 U12738 ( .IN1(n12799), .IN2(n12820), .QN(n12819) );
  NOR2X0 U12739 ( .IN1(n12821), .IN2(n12815), .QN(n12820) );
  NOR2X0 U12740 ( .IN1(n12783), .IN2(n12796), .QN(n12821) );
  NOR2X0 U12741 ( .IN1(n12822), .IN2(n12823), .QN(n12818) );
  NAND2X0 U12742 ( .IN1(n12815), .IN2(n12805), .QN(n12823) );
  NAND2X0 U12743 ( .IN1(n12797), .IN2(n12824), .QN(n12822) );
  NAND2X0 U12744 ( .IN1(n12756), .IN2(n12825), .QN(n12778) );
  INVX0 U12745 ( .INP(n12826), .ZN(n12825) );
  NOR2X0 U12746 ( .IN1(n12827), .IN2(n12754), .QN(n12826) );
  NAND2X0 U12747 ( .IN1(n12828), .IN2(n12829), .QN(n12754) );
  NAND2X0 U12748 ( .IN1(n12830), .IN2(n12792), .QN(n12829) );
  NAND2X0 U12749 ( .IN1(n12831), .IN2(n12832), .QN(n12830) );
  NAND2X0 U12750 ( .IN1(n12833), .IN2(n12796), .QN(n12832) );
  NAND2X0 U12751 ( .IN1(n12806), .IN2(n12834), .QN(n12831) );
  NAND2X0 U12752 ( .IN1(n12835), .IN2(n12836), .QN(n12834) );
  NAND2X0 U12753 ( .IN1(n12815), .IN2(n12812), .QN(n12836) );
  NOR2X0 U12754 ( .IN1(n12837), .IN2(n12838), .QN(n12835) );
  NOR2X0 U12755 ( .IN1(n12801), .IN2(n12839), .QN(n12838) );
  INVX0 U12756 ( .INP(n12840), .ZN(n12839) );
  NOR2X0 U12757 ( .IN1(n12796), .IN2(n12841), .QN(n12837) );
  NAND2X0 U12758 ( .IN1(n12807), .IN2(n12824), .QN(n12841) );
  NOR2X0 U12759 ( .IN1(n12842), .IN2(n12843), .QN(n12828) );
  NOR2X0 U12760 ( .IN1(n12806), .IN2(n12844), .QN(n12843) );
  NOR2X0 U12761 ( .IN1(n12845), .IN2(n12846), .QN(n12844) );
  NOR2X0 U12762 ( .IN1(n12847), .IN2(n12792), .QN(n12846) );
  NOR2X0 U12763 ( .IN1(n12848), .IN2(n12849), .QN(n12847) );
  NAND2X0 U12764 ( .IN1(n12850), .IN2(n12851), .QN(n12849) );
  NAND2X0 U12765 ( .IN1(n12840), .IN2(n12815), .QN(n12851) );
  INVX0 U12766 ( .INP(n12790), .ZN(n12815) );
  INVX0 U12767 ( .INP(n12852), .ZN(n12850) );
  NOR2X0 U12768 ( .IN1(n12813), .IN2(n12812), .QN(n12852) );
  NAND2X0 U12769 ( .IN1(n12853), .IN2(n12797), .QN(n12813) );
  NOR2X0 U12770 ( .IN1(n12785), .IN2(n12796), .QN(n12853) );
  INVX0 U12771 ( .INP(n12854), .ZN(n12796) );
  NAND2X0 U12772 ( .IN1(n12855), .IN2(n12856), .QN(n12854) );
  NAND2X0 U12773 ( .IN1(test_so63), .IN2(g1775), .QN(n12856) );
  NOR2X0 U12774 ( .IN1(n12857), .IN2(n12858), .QN(n12855) );
  NOR2X0 U12775 ( .IN1(n8624), .IN2(n8623), .QN(n12858) );
  NOR2X0 U12776 ( .IN1(n8622), .IN2(n8621), .QN(n12857) );
  INVX0 U12777 ( .INP(n12824), .ZN(n12785) );
  NOR2X0 U12778 ( .IN1(n12797), .IN2(n12824), .QN(n12848) );
  NOR2X0 U12779 ( .IN1(n12799), .IN2(n12801), .QN(n12845) );
  NAND2X0 U12780 ( .IN1(n12790), .IN2(n12824), .QN(n12801) );
  NOR2X0 U12781 ( .IN1(n12824), .IN2(n12859), .QN(n12842) );
  NAND2X0 U12782 ( .IN1(n12860), .IN2(n12812), .QN(n12859) );
  NAND2X0 U12783 ( .IN1(n12861), .IN2(n12862), .QN(n12860) );
  NAND2X0 U12784 ( .IN1(n12806), .IN2(n12797), .QN(n12862) );
  INVX0 U12785 ( .INP(n12800), .ZN(n12806) );
  NAND2X0 U12786 ( .IN1(n12863), .IN2(n12864), .QN(n12800) );
  NAND2X0 U12787 ( .IN1(test_so63), .IN2(g1730), .QN(n12864) );
  NOR2X0 U12788 ( .IN1(n12865), .IN2(n12866), .QN(n12863) );
  NOR2X0 U12789 ( .IN1(n8623), .IN2(n8616), .QN(n12866) );
  NOR2X0 U12790 ( .IN1(n8621), .IN2(n8615), .QN(n12865) );
  NAND2X0 U12791 ( .IN1(n12783), .IN2(n12790), .QN(n12861) );
  NAND2X0 U12792 ( .IN1(n12867), .IN2(n12868), .QN(n12790) );
  NAND2X0 U12793 ( .IN1(test_so63), .IN2(g1760), .QN(n12868) );
  NOR2X0 U12794 ( .IN1(n12869), .IN2(n12870), .QN(n12867) );
  NOR2X0 U12795 ( .IN1(n8623), .IN2(n8579), .QN(n12870) );
  NOR2X0 U12796 ( .IN1(n8621), .IN2(n8578), .QN(n12869) );
  NAND2X0 U12797 ( .IN1(n12871), .IN2(n12872), .QN(n12824) );
  NAND2X0 U12798 ( .IN1(test_so63), .IN2(g1745), .QN(n12872) );
  NOR2X0 U12799 ( .IN1(n12873), .IN2(n12874), .QN(n12871) );
  NOR2X0 U12800 ( .IN1(n8623), .IN2(n8405), .QN(n12874) );
  NOR2X0 U12801 ( .IN1(n8621), .IN2(n8404), .QN(n12873) );
  NAND2X0 U12802 ( .IN1(n12758), .IN2(n12827), .QN(n12756) );
  INVX0 U12803 ( .INP(n12875), .ZN(n12773) );
  NOR2X0 U12804 ( .IN1(n12749), .IN2(n8689), .QN(n12875) );
  NAND2X0 U12805 ( .IN1(n12876), .IN2(n12877), .QN(g28351) );
  NAND2X0 U12806 ( .IN1(n4371), .IN2(g1300), .QN(n12877) );
  NAND2X0 U12807 ( .IN1(n12641), .IN2(n12608), .QN(n12876) );
  NAND2X0 U12808 ( .IN1(n12878), .IN2(n12879), .QN(n12641) );
  NAND2X0 U12809 ( .IN1(n10436), .IN2(n12629), .QN(n12879) );
  NAND2X0 U12810 ( .IN1(n12880), .IN2(n12628), .QN(n12878) );
  NOR2X0 U12811 ( .IN1(n12881), .IN2(n12882), .QN(n12880) );
  NAND2X0 U12812 ( .IN1(n12883), .IN2(n12884), .QN(n12881) );
  INVX0 U12813 ( .INP(n12885), .ZN(n12883) );
  NOR2X0 U12814 ( .IN1(n12886), .IN2(n12887), .QN(n12885) );
  NAND2X0 U12815 ( .IN1(n12888), .IN2(n12889), .QN(g28350) );
  NAND2X0 U12816 ( .IN1(n4316), .IN2(g1294), .QN(n12889) );
  NAND2X0 U12817 ( .IN1(n12769), .IN2(g6944), .QN(n12888) );
  NAND2X0 U12818 ( .IN1(n12890), .IN2(n12891), .QN(g28349) );
  NAND2X0 U12819 ( .IN1(n4372), .IN2(g617), .QN(n12891) );
  NAND2X0 U12820 ( .IN1(n12772), .IN2(g6642), .QN(n12890) );
  NAND2X0 U12821 ( .IN1(n12892), .IN2(n12893), .QN(g28348) );
  INVX0 U12822 ( .INP(n12894), .ZN(n12893) );
  NOR2X0 U12823 ( .IN1(g550), .IN2(n8676), .QN(n12894) );
  NAND2X0 U12824 ( .IN1(n12895), .IN2(g550), .QN(n12892) );
  NAND2X0 U12825 ( .IN1(n12896), .IN2(n12897), .QN(g28346) );
  NAND2X0 U12826 ( .IN1(g6750), .IN2(n12769), .QN(n12897) );
  NAND2X0 U12827 ( .IN1(n12898), .IN2(n12899), .QN(n12769) );
  NAND2X0 U12828 ( .IN1(n10409), .IN2(n12629), .QN(n12899) );
  NAND2X0 U12829 ( .IN1(n12900), .IN2(n12628), .QN(n12898) );
  NOR2X0 U12830 ( .IN1(n12901), .IN2(n12887), .QN(n12900) );
  NAND2X0 U12831 ( .IN1(n12902), .IN2(n12903), .QN(n12887) );
  NOR2X0 U12832 ( .IN1(n12904), .IN2(n12905), .QN(n12903) );
  NOR2X0 U12833 ( .IN1(n12906), .IN2(n12907), .QN(n12905) );
  NAND2X0 U12834 ( .IN1(n12908), .IN2(n12909), .QN(n12907) );
  NAND2X0 U12835 ( .IN1(n12910), .IN2(n12911), .QN(n12909) );
  NAND2X0 U12836 ( .IN1(n12912), .IN2(n12913), .QN(n12911) );
  NOR2X0 U12837 ( .IN1(n12914), .IN2(n12915), .QN(n12904) );
  NOR2X0 U12838 ( .IN1(n12916), .IN2(n12917), .QN(n12914) );
  INVX0 U12839 ( .INP(n12918), .ZN(n12917) );
  NAND2X0 U12840 ( .IN1(n12912), .IN2(n12919), .QN(n12918) );
  NAND2X0 U12841 ( .IN1(n12920), .IN2(n12921), .QN(n12912) );
  NAND2X0 U12842 ( .IN1(n12922), .IN2(n12923), .QN(n12921) );
  NOR2X0 U12843 ( .IN1(n12910), .IN2(n12924), .QN(n12916) );
  INVX0 U12844 ( .INP(n12925), .ZN(n12910) );
  NAND2X0 U12845 ( .IN1(n12926), .IN2(n12927), .QN(n12925) );
  NAND2X0 U12846 ( .IN1(n12928), .IN2(n12929), .QN(n12927) );
  NAND2X0 U12847 ( .IN1(n12930), .IN2(n12923), .QN(n12926) );
  NOR2X0 U12848 ( .IN1(n12931), .IN2(n12932), .QN(n12902) );
  NOR2X0 U12849 ( .IN1(n12929), .IN2(n12933), .QN(n12932) );
  NAND2X0 U12850 ( .IN1(n12934), .IN2(n12935), .QN(n12933) );
  NAND2X0 U12851 ( .IN1(n12936), .IN2(n12937), .QN(n12934) );
  NAND2X0 U12852 ( .IN1(n12938), .IN2(n12939), .QN(n12937) );
  NAND2X0 U12853 ( .IN1(n12908), .IN2(n12930), .QN(n12939) );
  NOR2X0 U12854 ( .IN1(n12940), .IN2(n12923), .QN(n12931) );
  NOR2X0 U12855 ( .IN1(n12941), .IN2(n12942), .QN(n12940) );
  NOR2X0 U12856 ( .IN1(n12922), .IN2(n12943), .QN(n12942) );
  NOR2X0 U12857 ( .IN1(n12944), .IN2(n12938), .QN(n12943) );
  NOR2X0 U12858 ( .IN1(n12906), .IN2(n12919), .QN(n12944) );
  NOR2X0 U12859 ( .IN1(n12945), .IN2(n12946), .QN(n12941) );
  NAND2X0 U12860 ( .IN1(n12938), .IN2(n12928), .QN(n12946) );
  NAND2X0 U12861 ( .IN1(n12920), .IN2(n12947), .QN(n12945) );
  NAND2X0 U12862 ( .IN1(n12884), .IN2(n12948), .QN(n12901) );
  INVX0 U12863 ( .INP(n12949), .ZN(n12948) );
  NOR2X0 U12864 ( .IN1(n12950), .IN2(n12882), .QN(n12949) );
  NAND2X0 U12865 ( .IN1(n12951), .IN2(n12952), .QN(n12882) );
  NAND2X0 U12866 ( .IN1(n12953), .IN2(n12915), .QN(n12952) );
  NAND2X0 U12867 ( .IN1(n12954), .IN2(n12955), .QN(n12953) );
  NAND2X0 U12868 ( .IN1(n12956), .IN2(n12919), .QN(n12955) );
  NAND2X0 U12869 ( .IN1(n12929), .IN2(n12957), .QN(n12954) );
  NAND2X0 U12870 ( .IN1(n12958), .IN2(n12959), .QN(n12957) );
  NAND2X0 U12871 ( .IN1(n12938), .IN2(n12935), .QN(n12959) );
  NOR2X0 U12872 ( .IN1(n12960), .IN2(n12961), .QN(n12958) );
  NOR2X0 U12873 ( .IN1(n12924), .IN2(n12962), .QN(n12961) );
  INVX0 U12874 ( .INP(n12963), .ZN(n12962) );
  NOR2X0 U12875 ( .IN1(n12919), .IN2(n12964), .QN(n12960) );
  NAND2X0 U12876 ( .IN1(n12930), .IN2(n12947), .QN(n12964) );
  NOR2X0 U12877 ( .IN1(n12965), .IN2(n12966), .QN(n12951) );
  NOR2X0 U12878 ( .IN1(n12929), .IN2(n12967), .QN(n12966) );
  NOR2X0 U12879 ( .IN1(n12968), .IN2(n12969), .QN(n12967) );
  NOR2X0 U12880 ( .IN1(n12970), .IN2(n12915), .QN(n12969) );
  NOR2X0 U12881 ( .IN1(n12971), .IN2(n12972), .QN(n12970) );
  NAND2X0 U12882 ( .IN1(n12973), .IN2(n12974), .QN(n12972) );
  NAND2X0 U12883 ( .IN1(n12963), .IN2(n12938), .QN(n12974) );
  INVX0 U12884 ( .INP(n12913), .ZN(n12938) );
  INVX0 U12885 ( .INP(n12975), .ZN(n12973) );
  NOR2X0 U12886 ( .IN1(n12936), .IN2(n12935), .QN(n12975) );
  NAND2X0 U12887 ( .IN1(n12976), .IN2(n12920), .QN(n12936) );
  NOR2X0 U12888 ( .IN1(n12908), .IN2(n12919), .QN(n12976) );
  INVX0 U12889 ( .INP(n12977), .ZN(n12919) );
  NAND2X0 U12890 ( .IN1(n12978), .IN2(n12979), .QN(n12977) );
  NAND2X0 U12891 ( .IN1(g5686), .IN2(g1083), .QN(n12979) );
  NOR2X0 U12892 ( .IN1(n12980), .IN2(n12981), .QN(n12978) );
  NOR2X0 U12893 ( .IN1(n8627), .IN2(n8626), .QN(n12981) );
  NOR2X0 U12894 ( .IN1(n16822), .IN2(n8625), .QN(n12980) );
  INVX0 U12895 ( .INP(n12947), .ZN(n12908) );
  NOR2X0 U12896 ( .IN1(n12920), .IN2(n12947), .QN(n12971) );
  NOR2X0 U12897 ( .IN1(n12922), .IN2(n12924), .QN(n12968) );
  NAND2X0 U12898 ( .IN1(n12913), .IN2(n12947), .QN(n12924) );
  NOR2X0 U12899 ( .IN1(n12947), .IN2(n12982), .QN(n12965) );
  NAND2X0 U12900 ( .IN1(n12983), .IN2(n12935), .QN(n12982) );
  NAND2X0 U12901 ( .IN1(n12984), .IN2(n12985), .QN(n12983) );
  NAND2X0 U12902 ( .IN1(n12929), .IN2(n12920), .QN(n12985) );
  INVX0 U12903 ( .INP(n12923), .ZN(n12929) );
  NAND2X0 U12904 ( .IN1(n12986), .IN2(n12987), .QN(n12923) );
  NAND2X0 U12905 ( .IN1(g5657), .IN2(g1036), .QN(n12987) );
  NOR2X0 U12906 ( .IN1(n12988), .IN2(n12989), .QN(n12986) );
  NOR2X0 U12907 ( .IN1(n8628), .IN2(n8618), .QN(n12989) );
  NOR2X0 U12908 ( .IN1(n8626), .IN2(n8617), .QN(n12988) );
  NAND2X0 U12909 ( .IN1(n12906), .IN2(n12913), .QN(n12984) );
  NAND2X0 U12910 ( .IN1(n12990), .IN2(n12991), .QN(n12913) );
  NAND2X0 U12911 ( .IN1(g5657), .IN2(g1066), .QN(n12991) );
  NOR2X0 U12912 ( .IN1(n12992), .IN2(n12993), .QN(n12990) );
  NOR2X0 U12913 ( .IN1(n8628), .IN2(n8581), .QN(n12993) );
  NOR2X0 U12914 ( .IN1(n8626), .IN2(n8580), .QN(n12992) );
  NAND2X0 U12915 ( .IN1(n12994), .IN2(n12995), .QN(n12947) );
  NAND2X0 U12916 ( .IN1(g5657), .IN2(g1051), .QN(n12995) );
  NOR2X0 U12917 ( .IN1(n12996), .IN2(n12997), .QN(n12994) );
  NOR2X0 U12918 ( .IN1(n8628), .IN2(n8407), .QN(n12997) );
  NOR2X0 U12919 ( .IN1(n8626), .IN2(n8406), .QN(n12996) );
  NAND2X0 U12920 ( .IN1(n12886), .IN2(n12950), .QN(n12884) );
  INVX0 U12921 ( .INP(n12998), .ZN(n12896) );
  NOR2X0 U12922 ( .IN1(n12608), .IN2(n8692), .QN(n12998) );
  NAND2X0 U12923 ( .IN1(n12999), .IN2(n13000), .QN(g28345) );
  INVX0 U12924 ( .INP(n13001), .ZN(n13000) );
  NOR2X0 U12925 ( .IN1(n13002), .IN2(n8673), .QN(n13001) );
  NAND2X0 U12926 ( .IN1(n12772), .IN2(n13002), .QN(n12999) );
  NAND2X0 U12927 ( .IN1(n13003), .IN2(n13004), .QN(n12772) );
  NAND2X0 U12928 ( .IN1(n10010), .IN2(n12629), .QN(n13004) );
  NAND2X0 U12929 ( .IN1(n13005), .IN2(n12628), .QN(n13003) );
  NOR2X0 U12930 ( .IN1(n13006), .IN2(n13007), .QN(n13005) );
  NAND2X0 U12931 ( .IN1(n13008), .IN2(n13009), .QN(n13006) );
  INVX0 U12932 ( .INP(n13010), .ZN(n13008) );
  NOR2X0 U12933 ( .IN1(n13011), .IN2(n13012), .QN(n13010) );
  NAND2X0 U12934 ( .IN1(n13013), .IN2(n13014), .QN(g28344) );
  NAND2X0 U12935 ( .IN1(n4372), .IN2(g608), .QN(n13014) );
  NAND2X0 U12936 ( .IN1(n12895), .IN2(g6642), .QN(n13013) );
  NAND2X0 U12937 ( .IN1(n13015), .IN2(n13016), .QN(g28342) );
  NAND2X0 U12938 ( .IN1(g6485), .IN2(n12895), .QN(n13016) );
  NAND2X0 U12939 ( .IN1(n13017), .IN2(n13018), .QN(n12895) );
  NAND2X0 U12940 ( .IN1(n10001), .IN2(n12629), .QN(n13018) );
  INVX0 U12941 ( .INP(n12628), .ZN(n12629) );
  NAND2X0 U12942 ( .IN1(n13019), .IN2(n12628), .QN(n13017) );
  NOR2X0 U12943 ( .IN1(n13020), .IN2(n13012), .QN(n13019) );
  NAND2X0 U12944 ( .IN1(n13021), .IN2(n13022), .QN(n13012) );
  NOR2X0 U12945 ( .IN1(n13023), .IN2(n13024), .QN(n13022) );
  NOR2X0 U12946 ( .IN1(n13025), .IN2(n13026), .QN(n13024) );
  NAND2X0 U12947 ( .IN1(n13027), .IN2(n13028), .QN(n13026) );
  NAND2X0 U12948 ( .IN1(n13029), .IN2(n13030), .QN(n13028) );
  NAND2X0 U12949 ( .IN1(n13031), .IN2(n13032), .QN(n13030) );
  NOR2X0 U12950 ( .IN1(n13033), .IN2(n13034), .QN(n13023) );
  NOR2X0 U12951 ( .IN1(n13035), .IN2(n13036), .QN(n13033) );
  INVX0 U12952 ( .INP(n13037), .ZN(n13036) );
  NAND2X0 U12953 ( .IN1(n13031), .IN2(n13038), .QN(n13037) );
  NAND2X0 U12954 ( .IN1(n13039), .IN2(n13040), .QN(n13031) );
  NAND2X0 U12955 ( .IN1(n13041), .IN2(n13042), .QN(n13040) );
  NOR2X0 U12956 ( .IN1(n13029), .IN2(n13043), .QN(n13035) );
  INVX0 U12957 ( .INP(n13044), .ZN(n13029) );
  NAND2X0 U12958 ( .IN1(n13045), .IN2(n13046), .QN(n13044) );
  NAND2X0 U12959 ( .IN1(n13047), .IN2(n13048), .QN(n13046) );
  NAND2X0 U12960 ( .IN1(n13049), .IN2(n13042), .QN(n13045) );
  NOR2X0 U12961 ( .IN1(n13050), .IN2(n13051), .QN(n13021) );
  NOR2X0 U12962 ( .IN1(n13048), .IN2(n13052), .QN(n13051) );
  NAND2X0 U12963 ( .IN1(n13053), .IN2(n13054), .QN(n13052) );
  NAND2X0 U12964 ( .IN1(n13055), .IN2(n13056), .QN(n13053) );
  NAND2X0 U12965 ( .IN1(n13057), .IN2(n13058), .QN(n13056) );
  NAND2X0 U12966 ( .IN1(n13027), .IN2(n13049), .QN(n13058) );
  NOR2X0 U12967 ( .IN1(n13059), .IN2(n13042), .QN(n13050) );
  NOR2X0 U12968 ( .IN1(n13060), .IN2(n13061), .QN(n13059) );
  NOR2X0 U12969 ( .IN1(n13041), .IN2(n13062), .QN(n13061) );
  NOR2X0 U12970 ( .IN1(n13063), .IN2(n13057), .QN(n13062) );
  NOR2X0 U12971 ( .IN1(n13025), .IN2(n13038), .QN(n13063) );
  NOR2X0 U12972 ( .IN1(n13064), .IN2(n13065), .QN(n13060) );
  NAND2X0 U12973 ( .IN1(n13057), .IN2(n13047), .QN(n13065) );
  NAND2X0 U12974 ( .IN1(n13039), .IN2(n13066), .QN(n13064) );
  NAND2X0 U12975 ( .IN1(n13009), .IN2(n13067), .QN(n13020) );
  INVX0 U12976 ( .INP(n13068), .ZN(n13067) );
  NOR2X0 U12977 ( .IN1(n13069), .IN2(n13007), .QN(n13068) );
  NAND2X0 U12978 ( .IN1(n13070), .IN2(n13071), .QN(n13007) );
  NAND2X0 U12979 ( .IN1(n13072), .IN2(n13034), .QN(n13071) );
  NAND2X0 U12980 ( .IN1(n13073), .IN2(n13074), .QN(n13072) );
  NAND2X0 U12981 ( .IN1(n13075), .IN2(n13038), .QN(n13074) );
  NAND2X0 U12982 ( .IN1(n13048), .IN2(n13076), .QN(n13073) );
  NAND2X0 U12983 ( .IN1(n13077), .IN2(n13078), .QN(n13076) );
  NAND2X0 U12984 ( .IN1(n13057), .IN2(n13054), .QN(n13078) );
  NOR2X0 U12985 ( .IN1(n13079), .IN2(n13080), .QN(n13077) );
  NOR2X0 U12986 ( .IN1(n13043), .IN2(n13081), .QN(n13080) );
  INVX0 U12987 ( .INP(n13082), .ZN(n13081) );
  NOR2X0 U12988 ( .IN1(n13038), .IN2(n13083), .QN(n13079) );
  NAND2X0 U12989 ( .IN1(n13049), .IN2(n13066), .QN(n13083) );
  NOR2X0 U12990 ( .IN1(n13084), .IN2(n13085), .QN(n13070) );
  NOR2X0 U12991 ( .IN1(n13048), .IN2(n13086), .QN(n13085) );
  NOR2X0 U12992 ( .IN1(n13087), .IN2(n13088), .QN(n13086) );
  NOR2X0 U12993 ( .IN1(n13089), .IN2(n13034), .QN(n13088) );
  NOR2X0 U12994 ( .IN1(n13090), .IN2(n13091), .QN(n13089) );
  NAND2X0 U12995 ( .IN1(n13092), .IN2(n13093), .QN(n13091) );
  NAND2X0 U12996 ( .IN1(n13082), .IN2(n13057), .QN(n13093) );
  INVX0 U12997 ( .INP(n13032), .ZN(n13057) );
  INVX0 U12998 ( .INP(n13094), .ZN(n13092) );
  NOR2X0 U12999 ( .IN1(n13055), .IN2(n13054), .QN(n13094) );
  NAND2X0 U13000 ( .IN1(n13095), .IN2(n13039), .QN(n13055) );
  NOR2X0 U13001 ( .IN1(n13027), .IN2(n13038), .QN(n13095) );
  INVX0 U13002 ( .INP(n13096), .ZN(n13038) );
  NAND2X0 U13003 ( .IN1(n13097), .IN2(n13098), .QN(n13096) );
  NAND2X0 U13004 ( .IN1(g5648), .IN2(g396), .QN(n13098) );
  NOR2X0 U13005 ( .IN1(n13099), .IN2(n13100), .QN(n13097) );
  NOR2X0 U13006 ( .IN1(n8632), .IN2(n8631), .QN(n13100) );
  NOR2X0 U13007 ( .IN1(n16823), .IN2(n8630), .QN(n13099) );
  INVX0 U13008 ( .INP(n13066), .ZN(n13027) );
  NOR2X0 U13009 ( .IN1(n13039), .IN2(n13066), .QN(n13090) );
  NOR2X0 U13010 ( .IN1(n13041), .IN2(n13043), .QN(n13087) );
  NAND2X0 U13011 ( .IN1(n13032), .IN2(n13066), .QN(n13043) );
  NOR2X0 U13012 ( .IN1(n13066), .IN2(n13101), .QN(n13084) );
  NAND2X0 U13013 ( .IN1(n13102), .IN2(n13054), .QN(n13101) );
  NAND2X0 U13014 ( .IN1(n13103), .IN2(n13104), .QN(n13102) );
  NAND2X0 U13015 ( .IN1(n13048), .IN2(n13039), .QN(n13104) );
  INVX0 U13016 ( .INP(n13042), .ZN(n13048) );
  NAND2X0 U13017 ( .IN1(n13105), .IN2(n13106), .QN(n13042) );
  NAND2X0 U13018 ( .IN1(g5629), .IN2(g349), .QN(n13106) );
  NOR2X0 U13019 ( .IN1(n13107), .IN2(n13108), .QN(n13105) );
  NOR2X0 U13020 ( .IN1(n8633), .IN2(n8620), .QN(n13108) );
  NOR2X0 U13021 ( .IN1(n8631), .IN2(n8619), .QN(n13107) );
  NAND2X0 U13022 ( .IN1(n13025), .IN2(n13032), .QN(n13103) );
  NAND2X0 U13023 ( .IN1(n13109), .IN2(n13110), .QN(n13032) );
  NAND2X0 U13024 ( .IN1(g5629), .IN2(g379), .QN(n13110) );
  NOR2X0 U13025 ( .IN1(n13111), .IN2(n13112), .QN(n13109) );
  NOR2X0 U13026 ( .IN1(n8633), .IN2(n8583), .QN(n13112) );
  NOR2X0 U13027 ( .IN1(n8631), .IN2(n8582), .QN(n13111) );
  NAND2X0 U13028 ( .IN1(n13113), .IN2(n13114), .QN(n13066) );
  NAND2X0 U13029 ( .IN1(g5629), .IN2(g364), .QN(n13114) );
  NOR2X0 U13030 ( .IN1(n13115), .IN2(n13116), .QN(n13113) );
  NOR2X0 U13031 ( .IN1(n8633), .IN2(n8409), .QN(n13116) );
  NOR2X0 U13032 ( .IN1(n8631), .IN2(n8408), .QN(n13115) );
  NAND2X0 U13033 ( .IN1(n13011), .IN2(n13069), .QN(n13009) );
  INVX0 U13034 ( .INP(n13117), .ZN(n13015) );
  NOR2X0 U13035 ( .IN1(n13002), .IN2(n8675), .QN(n13117) );
  NOR2X0 U13036 ( .IN1(n10617), .IN2(n13118), .QN(g28328) );
  XOR2X1 U13037 ( .IN1(n4415), .IN2(n10618), .Q(n13118) );
  NOR2X0 U13038 ( .IN1(n10619), .IN2(n4393), .QN(n10618) );
  NAND2X0 U13039 ( .IN1(n13119), .IN2(n13120), .QN(g28325) );
  INVX0 U13040 ( .INP(n13121), .ZN(n13120) );
  NOR2X0 U13041 ( .IN1(n13122), .IN2(n4416), .QN(n13121) );
  NAND2X0 U13042 ( .IN1(n13123), .IN2(n4416), .QN(n13119) );
  NOR2X0 U13043 ( .IN1(n9284), .IN2(n13124), .QN(n13123) );
  NAND2X0 U13044 ( .IN1(n13125), .IN2(n13126), .QN(n13124) );
  NAND2X0 U13045 ( .IN1(n13127), .IN2(n13128), .QN(g28321) );
  INVX0 U13046 ( .INP(n13129), .ZN(n13128) );
  NOR2X0 U13047 ( .IN1(n13130), .IN2(n4417), .QN(n13129) );
  NAND2X0 U13048 ( .IN1(n13131), .IN2(n4417), .QN(n13127) );
  NOR2X0 U13049 ( .IN1(n13132), .IN2(n13133), .QN(n13131) );
  NAND2X0 U13050 ( .IN1(n13134), .IN2(g1372), .QN(n13133) );
  NOR2X0 U13051 ( .IN1(n13135), .IN2(n12578), .QN(g28148) );
  NAND2X0 U13052 ( .IN1(n3160), .IN2(n12385), .QN(n12578) );
  INVX0 U13053 ( .INP(n9702), .ZN(n12385) );
  NAND2X0 U13054 ( .IN1(n3424), .IN2(g2138), .QN(n3160) );
  NOR2X0 U13055 ( .IN1(n3424), .IN2(g2138), .QN(n13135) );
  NOR2X0 U13056 ( .IN1(n13136), .IN2(n12583), .QN(g28147) );
  NAND2X0 U13057 ( .IN1(n3164), .IN2(n12387), .QN(n12583) );
  INVX0 U13058 ( .INP(n9710), .ZN(n12387) );
  NAND2X0 U13059 ( .IN1(n3427), .IN2(g1444), .QN(n3164) );
  NOR2X0 U13060 ( .IN1(n3427), .IN2(g1444), .QN(n13136) );
  NOR2X0 U13061 ( .IN1(n13137), .IN2(n12588), .QN(g28146) );
  NAND2X0 U13062 ( .IN1(n3168), .IN2(n12389), .QN(n12588) );
  NAND2X0 U13063 ( .IN1(n3430), .IN2(g758), .QN(n3168) );
  NOR2X0 U13064 ( .IN1(n3430), .IN2(g758), .QN(n13137) );
  NOR2X0 U13065 ( .IN1(n13138), .IN2(n12593), .QN(g28145) );
  NAND2X0 U13066 ( .IN1(n3172), .IN2(n12391), .QN(n12593) );
  INVX0 U13067 ( .INP(n9719), .ZN(n12391) );
  NAND2X0 U13068 ( .IN1(n3433), .IN2(g70), .QN(n3172) );
  NOR2X0 U13069 ( .IN1(n3433), .IN2(g70), .QN(n13138) );
  NAND2X0 U13070 ( .IN1(n13139), .IN2(n13140), .QN(g27771) );
  NAND2X0 U13071 ( .IN1(test_so81), .IN2(n13141), .QN(n13140) );
  NAND2X0 U13072 ( .IN1(n13142), .IN2(n11841), .QN(n13141) );
  NAND2X0 U13073 ( .IN1(n13143), .IN2(n11841), .QN(n13139) );
  NAND2X0 U13074 ( .IN1(n13144), .IN2(n13145), .QN(g27769) );
  NAND2X0 U13075 ( .IN1(n13146), .IN2(g2524), .QN(n13145) );
  NAND2X0 U13076 ( .IN1(n13142), .IN2(n10669), .QN(n13146) );
  NAND2X0 U13077 ( .IN1(n13143), .IN2(n10669), .QN(n13144) );
  NAND2X0 U13078 ( .IN1(n13147), .IN2(n13148), .QN(g27768) );
  NAND2X0 U13079 ( .IN1(n13149), .IN2(g1828), .QN(n13148) );
  NAND2X0 U13080 ( .IN1(n13150), .IN2(n11849), .QN(n13149) );
  NAND2X0 U13081 ( .IN1(n13151), .IN2(n11849), .QN(n13147) );
  NAND2X0 U13082 ( .IN1(n13152), .IN2(n13153), .QN(g27767) );
  NAND2X0 U13083 ( .IN1(n13154), .IN2(g2523), .QN(n13153) );
  NAND2X0 U13084 ( .IN1(n13142), .IN2(n11931), .QN(n13154) );
  INVX0 U13085 ( .INP(n13155), .ZN(n13142) );
  NAND2X0 U13086 ( .IN1(n13156), .IN2(n13157), .QN(n13155) );
  NOR2X0 U13087 ( .IN1(n13158), .IN2(n13159), .QN(n13157) );
  NOR2X0 U13088 ( .IN1(n9281), .IN2(n13160), .QN(n13156) );
  NAND2X0 U13089 ( .IN1(n13143), .IN2(n11931), .QN(n13152) );
  NOR2X0 U13090 ( .IN1(n13161), .IN2(n9281), .QN(n13143) );
  INVX0 U13091 ( .INP(n13162), .ZN(n13161) );
  NOR2X0 U13092 ( .IN1(n13163), .IN2(n13164), .QN(n13162) );
  NOR2X0 U13093 ( .IN1(n13165), .IN2(n13166), .QN(n13164) );
  NOR2X0 U13094 ( .IN1(n13167), .IN2(n13168), .QN(n13165) );
  NOR2X0 U13095 ( .IN1(n13169), .IN2(n13170), .QN(n13163) );
  NOR2X0 U13096 ( .IN1(n13171), .IN2(n13172), .QN(n13170) );
  NAND2X0 U13097 ( .IN1(n13173), .IN2(n13174), .QN(g27766) );
  NAND2X0 U13098 ( .IN1(n13175), .IN2(g1830), .QN(n13174) );
  NAND2X0 U13099 ( .IN1(n13150), .IN2(n10678), .QN(n13175) );
  NAND2X0 U13100 ( .IN1(n13151), .IN2(n10678), .QN(n13173) );
  NAND2X0 U13101 ( .IN1(n13176), .IN2(n13177), .QN(g27765) );
  NAND2X0 U13102 ( .IN1(n13178), .IN2(g1134), .QN(n13177) );
  NAND2X0 U13103 ( .IN1(n13179), .IN2(g1088), .QN(n13178) );
  NAND2X0 U13104 ( .IN1(n13180), .IN2(g1088), .QN(n13176) );
  NAND2X0 U13105 ( .IN1(n13181), .IN2(n13182), .QN(g27764) );
  NAND2X0 U13106 ( .IN1(n13183), .IN2(g1829), .QN(n13182) );
  NAND2X0 U13107 ( .IN1(n13150), .IN2(n12050), .QN(n13183) );
  NOR2X0 U13108 ( .IN1(n13184), .IN2(n13185), .QN(n13150) );
  NAND2X0 U13109 ( .IN1(n13186), .IN2(n13187), .QN(n13184) );
  NAND2X0 U13110 ( .IN1(n13151), .IN2(n12050), .QN(n13181) );
  NAND2X0 U13111 ( .IN1(n13188), .IN2(n13189), .QN(n13151) );
  NAND2X0 U13112 ( .IN1(n13190), .IN2(n13191), .QN(n13189) );
  NAND2X0 U13113 ( .IN1(n13192), .IN2(n13193), .QN(n13188) );
  NAND2X0 U13114 ( .IN1(n13194), .IN2(n13195), .QN(g27763) );
  NAND2X0 U13115 ( .IN1(n13196), .IN2(g1136), .QN(n13195) );
  NAND2X0 U13116 ( .IN1(n13179), .IN2(g6712), .QN(n13196) );
  NAND2X0 U13117 ( .IN1(n13180), .IN2(g6712), .QN(n13194) );
  NAND2X0 U13118 ( .IN1(n13197), .IN2(n13198), .QN(g27762) );
  NAND2X0 U13119 ( .IN1(n13199), .IN2(g447), .QN(n13198) );
  NAND2X0 U13120 ( .IN1(n13200), .IN2(n11886), .QN(n13199) );
  NAND2X0 U13121 ( .IN1(n13201), .IN2(n11886), .QN(n13197) );
  NAND2X0 U13122 ( .IN1(n13202), .IN2(n13203), .QN(g27761) );
  NAND2X0 U13123 ( .IN1(n13204), .IN2(g1135), .QN(n13203) );
  NAND2X0 U13124 ( .IN1(n13179), .IN2(g5472), .QN(n13204) );
  NOR2X0 U13125 ( .IN1(n13205), .IN2(n13206), .QN(n13179) );
  NAND2X0 U13126 ( .IN1(n13207), .IN2(n13208), .QN(n13205) );
  NAND2X0 U13127 ( .IN1(n13180), .IN2(g5472), .QN(n13202) );
  NAND2X0 U13128 ( .IN1(n13209), .IN2(n13210), .QN(n13180) );
  NAND2X0 U13129 ( .IN1(n13211), .IN2(n13212), .QN(n13210) );
  NAND2X0 U13130 ( .IN1(n13213), .IN2(n13214), .QN(n13209) );
  NAND2X0 U13131 ( .IN1(n13215), .IN2(n13216), .QN(g27760) );
  NAND2X0 U13132 ( .IN1(n13217), .IN2(g449), .QN(n13216) );
  NAND2X0 U13133 ( .IN1(n13200), .IN2(n11905), .QN(n13217) );
  NAND2X0 U13134 ( .IN1(n13201), .IN2(n11905), .QN(n13215) );
  NAND2X0 U13135 ( .IN1(n13218), .IN2(n13219), .QN(g27759) );
  NAND2X0 U13136 ( .IN1(n13220), .IN2(g448), .QN(n13219) );
  NAND2X0 U13137 ( .IN1(n13200), .IN2(n10752), .QN(n13220) );
  NOR2X0 U13138 ( .IN1(n13221), .IN2(n13222), .QN(n13200) );
  NAND2X0 U13139 ( .IN1(n13223), .IN2(n13224), .QN(n13221) );
  NAND2X0 U13140 ( .IN1(n13201), .IN2(n10752), .QN(n13218) );
  NAND2X0 U13141 ( .IN1(n13225), .IN2(n13226), .QN(n13201) );
  NAND2X0 U13142 ( .IN1(n13227), .IN2(n13228), .QN(n13226) );
  NAND2X0 U13143 ( .IN1(n13229), .IN2(n13230), .QN(n13225) );
  NOR2X0 U13144 ( .IN1(n13231), .IN2(n13122), .QN(g27722) );
  NAND2X0 U13145 ( .IN1(n13126), .IN2(n13232), .QN(n13122) );
  NAND2X0 U13146 ( .IN1(test_so70), .IN2(n13125), .QN(n13232) );
  NOR2X0 U13147 ( .IN1(n13125), .IN2(test_so70), .QN(n13231) );
  INVX0 U13148 ( .INP(n13233), .ZN(n13125) );
  NOR2X0 U13149 ( .IN1(n13234), .IN2(n13130), .QN(g27718) );
  NAND2X0 U13150 ( .IN1(n13134), .IN2(n13235), .QN(n13130) );
  NAND2X0 U13151 ( .IN1(n13236), .IN2(g1372), .QN(n13235) );
  NOR2X0 U13152 ( .IN1(n13236), .IN2(g1372), .QN(n13234) );
  INVX0 U13153 ( .INP(n13132), .ZN(n13236) );
  NOR2X0 U13154 ( .IN1(n13237), .IN2(n13238), .QN(g27682) );
  NAND2X0 U13155 ( .IN1(n13233), .IN2(n13126), .QN(n13238) );
  NAND2X0 U13156 ( .IN1(n13239), .IN2(n13240), .QN(n13233) );
  NOR2X0 U13157 ( .IN1(n4473), .IN2(n4468), .QN(n13239) );
  NOR2X0 U13158 ( .IN1(n13241), .IN2(g2059), .QN(n13237) );
  NOR2X0 U13159 ( .IN1(n4468), .IN2(n13242), .QN(n13241) );
  NOR2X0 U13160 ( .IN1(n13243), .IN2(n13244), .QN(g27678) );
  NAND2X0 U13161 ( .IN1(n13132), .IN2(n13134), .QN(n13244) );
  NAND2X0 U13162 ( .IN1(n13245), .IN2(n13246), .QN(n13132) );
  NOR2X0 U13163 ( .IN1(n4475), .IN2(n4469), .QN(n13245) );
  NOR2X0 U13164 ( .IN1(n13247), .IN2(g1365), .QN(n13243) );
  NOR2X0 U13165 ( .IN1(n4469), .IN2(n13248), .QN(n13247) );
  NOR2X0 U13166 ( .IN1(n13249), .IN2(n13250), .QN(g27672) );
  NAND2X0 U13167 ( .IN1(n13251), .IN2(n9686), .QN(n13250) );
  NAND2X0 U13168 ( .IN1(n13252), .IN2(test_so28), .QN(n9686) );
  NOR2X0 U13169 ( .IN1(n4477), .IN2(n13253), .QN(n13252) );
  NOR2X0 U13170 ( .IN1(n13254), .IN2(g679), .QN(n13249) );
  NOR2X0 U13171 ( .IN1(n13253), .IN2(n9283), .QN(n13254) );
  NOR2X0 U13172 ( .IN1(n9702), .IN2(n13255), .QN(g27621) );
  XNOR2X1 U13173 ( .IN1(n4522), .IN2(n8970), .Q(n13255) );
  NOR2X0 U13174 ( .IN1(n9710), .IN2(n13256), .QN(g27612) );
  XNOR2X1 U13175 ( .IN1(n4523), .IN2(n8974), .Q(n13256) );
  NAND2X0 U13176 ( .IN1(n13257), .IN2(n13258), .QN(g27603) );
  INVX0 U13177 ( .INP(n13259), .ZN(n13258) );
  NOR2X0 U13178 ( .IN1(n13260), .IN2(n8978), .QN(n13259) );
  NAND2X0 U13179 ( .IN1(n13261), .IN2(n8978), .QN(n13257) );
  NOR2X0 U13180 ( .IN1(n11814), .IN2(n3431), .QN(n13261) );
  NOR2X0 U13181 ( .IN1(n9719), .IN2(n13262), .QN(g27594) );
  XNOR2X1 U13182 ( .IN1(n4521), .IN2(n8982), .Q(n13262) );
  NAND2X0 U13183 ( .IN1(n13263), .IN2(n13264), .QN(g27380) );
  NOR2X0 U13184 ( .IN1(n13265), .IN2(n13266), .QN(n13264) );
  NAND2X0 U13185 ( .IN1(n13267), .IN2(n13268), .QN(n13266) );
  NAND2X0 U13186 ( .IN1(n13269), .IN2(n13270), .QN(n13268) );
  NAND2X0 U13187 ( .IN1(n13271), .IN2(n13272), .QN(n13270) );
  NAND2X0 U13188 ( .IN1(n13273), .IN2(n4384), .QN(n13272) );
  NOR2X0 U13189 ( .IN1(n4405), .IN2(n13274), .QN(n13273) );
  INVX0 U13190 ( .INP(n13275), .ZN(n13267) );
  NOR2X0 U13191 ( .IN1(n13276), .IN2(n4424), .QN(n13275) );
  NAND2X0 U13192 ( .IN1(n13277), .IN2(n13278), .QN(n13265) );
  NAND2X0 U13193 ( .IN1(n13279), .IN2(n13280), .QN(n13277) );
  NOR2X0 U13194 ( .IN1(n13281), .IN2(n13282), .QN(n13280) );
  NOR2X0 U13195 ( .IN1(n16830), .IN2(n13283), .QN(n13282) );
  NOR2X0 U13196 ( .IN1(n16831), .IN2(n13284), .QN(n13281) );
  INVX0 U13197 ( .INP(n13285), .ZN(n13284) );
  NOR2X0 U13198 ( .IN1(n13286), .IN2(n13274), .QN(n13279) );
  NOR2X0 U13199 ( .IN1(n13287), .IN2(n13288), .QN(n13263) );
  NAND2X0 U13200 ( .IN1(n13289), .IN2(n13290), .QN(n13288) );
  INVX0 U13201 ( .INP(n13291), .ZN(n13290) );
  NOR2X0 U13202 ( .IN1(n13292), .IN2(n16825), .QN(n13291) );
  NAND2X0 U13203 ( .IN1(n8696), .IN2(n13293), .QN(n13289) );
  INVX0 U13204 ( .INP(n3700), .ZN(n13287) );
  NAND2X0 U13205 ( .IN1(n13294), .IN2(n13295), .QN(g27354) );
  NAND2X0 U13206 ( .IN1(n13296), .IN2(g2658), .QN(n13295) );
  NAND2X0 U13207 ( .IN1(n13297), .IN2(n13298), .QN(n13294) );
  NAND2X0 U13208 ( .IN1(n13299), .IN2(n13300), .QN(g27348) );
  NAND2X0 U13209 ( .IN1(n13301), .IN2(n13298), .QN(n13300) );
  INVX0 U13210 ( .INP(n13302), .ZN(n13299) );
  NOR2X0 U13211 ( .IN1(n13301), .IN2(n8601), .QN(n13302) );
  NAND2X0 U13212 ( .IN1(n13303), .IN2(n13304), .QN(g27347) );
  NAND2X0 U13213 ( .IN1(n13296), .IN2(g2655), .QN(n13304) );
  NAND2X0 U13214 ( .IN1(n13297), .IN2(n13305), .QN(n13303) );
  NAND2X0 U13215 ( .IN1(n13306), .IN2(n13307), .QN(g27346) );
  INVX0 U13216 ( .INP(n13308), .ZN(n13307) );
  NOR2X0 U13217 ( .IN1(n13309), .IN2(n8602), .QN(n13308) );
  NAND2X0 U13218 ( .IN1(n13309), .IN2(n13310), .QN(n13306) );
  NAND2X0 U13219 ( .IN1(n13311), .IN2(n13312), .QN(g27345) );
  NAND2X0 U13220 ( .IN1(n13313), .IN2(n13298), .QN(n13312) );
  NAND2X0 U13221 ( .IN1(n12703), .IN2(n13314), .QN(n13298) );
  NOR2X0 U13222 ( .IN1(n12676), .IN2(n12681), .QN(n12703) );
  NAND2X0 U13223 ( .IN1(n13315), .IN2(g2659), .QN(n13311) );
  NAND2X0 U13224 ( .IN1(n13316), .IN2(n13317), .QN(g27344) );
  NAND2X0 U13225 ( .IN1(test_so89), .IN2(n13318), .QN(n13317) );
  NAND2X0 U13226 ( .IN1(n13301), .IN2(n13305), .QN(n13316) );
  NAND2X0 U13227 ( .IN1(n13319), .IN2(n13320), .QN(g27343) );
  NAND2X0 U13228 ( .IN1(n13296), .IN2(g2652), .QN(n13320) );
  NAND2X0 U13229 ( .IN1(n13321), .IN2(n13297), .QN(n13319) );
  NAND2X0 U13230 ( .IN1(n13322), .IN2(n13323), .QN(g27342) );
  NAND2X0 U13231 ( .IN1(n13324), .IN2(g2466), .QN(n13323) );
  NAND2X0 U13232 ( .IN1(n13325), .IN2(n13326), .QN(n13322) );
  NAND2X0 U13233 ( .IN1(n13327), .IN2(n13328), .QN(g27341) );
  NAND2X0 U13234 ( .IN1(n13329), .IN2(g1966), .QN(n13328) );
  NAND2X0 U13235 ( .IN1(n13330), .IN2(n13310), .QN(n13327) );
  NAND2X0 U13236 ( .IN1(n13331), .IN2(n13332), .QN(g27340) );
  INVX0 U13237 ( .INP(n13333), .ZN(n13332) );
  NOR2X0 U13238 ( .IN1(n13309), .IN2(n8395), .QN(n13333) );
  NAND2X0 U13239 ( .IN1(n13309), .IN2(n13334), .QN(n13331) );
  NAND2X0 U13240 ( .IN1(n13335), .IN2(n13336), .QN(g27339) );
  NAND2X0 U13241 ( .IN1(n13337), .IN2(g1270), .QN(n13336) );
  NAND2X0 U13242 ( .IN1(n13338), .IN2(n13339), .QN(n13335) );
  NAND2X0 U13243 ( .IN1(n13340), .IN2(n13341), .QN(g27338) );
  NAND2X0 U13244 ( .IN1(n13315), .IN2(g2656), .QN(n13341) );
  NAND2X0 U13245 ( .IN1(n13313), .IN2(n13305), .QN(n13340) );
  INVX0 U13246 ( .INP(n13342), .ZN(n13305) );
  NAND2X0 U13247 ( .IN1(n13343), .IN2(n13344), .QN(n13342) );
  NAND2X0 U13248 ( .IN1(n12710), .IN2(n13345), .QN(n13344) );
  NOR2X0 U13249 ( .IN1(n12681), .IN2(n13346), .QN(n12710) );
  NAND2X0 U13250 ( .IN1(n13314), .IN2(n12681), .QN(n13343) );
  NAND2X0 U13251 ( .IN1(n13347), .IN2(n13348), .QN(g27337) );
  INVX0 U13252 ( .INP(n13349), .ZN(n13348) );
  NOR2X0 U13253 ( .IN1(n13301), .IN2(n8586), .QN(n13349) );
  NAND2X0 U13254 ( .IN1(n13321), .IN2(n13301), .QN(n13347) );
  NAND2X0 U13255 ( .IN1(n13350), .IN2(n13351), .QN(g27336) );
  NAND2X0 U13256 ( .IN1(n13296), .IN2(g2649), .QN(n13351) );
  NAND2X0 U13257 ( .IN1(n13352), .IN2(n13297), .QN(n13350) );
  INVX0 U13258 ( .INP(n13296), .ZN(n13297) );
  NAND2X0 U13259 ( .IN1(g2624), .IN2(g22687), .QN(n13296) );
  NAND2X0 U13260 ( .IN1(n13353), .IN2(n13354), .QN(g27335) );
  NAND2X0 U13261 ( .IN1(n13355), .IN2(n13326), .QN(n13354) );
  INVX0 U13262 ( .INP(n13356), .ZN(n13353) );
  NOR2X0 U13263 ( .IN1(n13355), .IN2(n8915), .QN(n13356) );
  NAND2X0 U13264 ( .IN1(n13357), .IN2(n13358), .QN(g27334) );
  NAND2X0 U13265 ( .IN1(n13324), .IN2(g2451), .QN(n13358) );
  NAND2X0 U13266 ( .IN1(n13325), .IN2(n13359), .QN(n13357) );
  NAND2X0 U13267 ( .IN1(n13360), .IN2(n13361), .QN(g27333) );
  NAND2X0 U13268 ( .IN1(n13362), .IN2(n13310), .QN(n13361) );
  NAND2X0 U13269 ( .IN1(n12833), .IN2(n13363), .QN(n13310) );
  NOR2X0 U13270 ( .IN1(n12807), .IN2(n12812), .QN(n12833) );
  NAND2X0 U13271 ( .IN1(test_so67), .IN2(n13364), .QN(n13360) );
  NAND2X0 U13272 ( .IN1(n13365), .IN2(n13366), .QN(g27332) );
  NAND2X0 U13273 ( .IN1(n13329), .IN2(g1963), .QN(n13366) );
  NAND2X0 U13274 ( .IN1(n13330), .IN2(n13334), .QN(n13365) );
  NAND2X0 U13275 ( .IN1(n13367), .IN2(n13368), .QN(g27331) );
  INVX0 U13276 ( .INP(n13369), .ZN(n13368) );
  NOR2X0 U13277 ( .IN1(n13309), .IN2(n8588), .QN(n13369) );
  NAND2X0 U13278 ( .IN1(n13370), .IN2(n13309), .QN(n13367) );
  NAND2X0 U13279 ( .IN1(n13371), .IN2(n13372), .QN(g27330) );
  NAND2X0 U13280 ( .IN1(n13373), .IN2(g1772), .QN(n13372) );
  NAND2X0 U13281 ( .IN1(n13374), .IN2(n13375), .QN(n13371) );
  NAND2X0 U13282 ( .IN1(n13376), .IN2(n13377), .QN(g27329) );
  NAND2X0 U13283 ( .IN1(n13378), .IN2(g1272), .QN(n13377) );
  NAND2X0 U13284 ( .IN1(n13379), .IN2(n13339), .QN(n13376) );
  NAND2X0 U13285 ( .IN1(n13380), .IN2(n13381), .QN(g27328) );
  NAND2X0 U13286 ( .IN1(test_so46), .IN2(n13337), .QN(n13381) );
  NAND2X0 U13287 ( .IN1(n13338), .IN2(n13382), .QN(n13380) );
  NAND2X0 U13288 ( .IN1(n13383), .IN2(n13384), .QN(g27327) );
  NAND2X0 U13289 ( .IN1(n13385), .IN2(g584), .QN(n13384) );
  NAND2X0 U13290 ( .IN1(n13386), .IN2(n13387), .QN(n13383) );
  NAND2X0 U13291 ( .IN1(n13388), .IN2(n13389), .QN(g27326) );
  NAND2X0 U13292 ( .IN1(n13315), .IN2(g2653), .QN(n13389) );
  NAND2X0 U13293 ( .IN1(n13321), .IN2(n13313), .QN(n13388) );
  NOR2X0 U13294 ( .IN1(n13390), .IN2(n13391), .QN(n13321) );
  NOR2X0 U13295 ( .IN1(n13314), .IN2(n12666), .QN(n13391) );
  INVX0 U13296 ( .INP(n13345), .ZN(n13314) );
  XNOR2X1 U13297 ( .IN1(n12652), .IN2(n10022), .Q(n13345) );
  INVX0 U13298 ( .INP(n12661), .ZN(n12652) );
  NAND2X0 U13299 ( .IN1(n13392), .IN2(n13393), .QN(g27325) );
  INVX0 U13300 ( .INP(n13394), .ZN(n13393) );
  NOR2X0 U13301 ( .IN1(n13301), .IN2(n8566), .QN(n13394) );
  NAND2X0 U13302 ( .IN1(n13352), .IN2(n13301), .QN(n13392) );
  INVX0 U13303 ( .INP(n13318), .ZN(n13301) );
  NAND2X0 U13304 ( .IN1(g7390), .IN2(g22687), .QN(n13318) );
  NAND2X0 U13305 ( .IN1(n13395), .IN2(n13396), .QN(g27324) );
  NAND2X0 U13306 ( .IN1(n13397), .IN2(n13326), .QN(n13396) );
  NAND2X0 U13307 ( .IN1(n13398), .IN2(n13399), .QN(n13326) );
  NOR2X0 U13308 ( .IN1(n13400), .IN2(n13401), .QN(n13398) );
  NAND2X0 U13309 ( .IN1(n13402), .IN2(g2473), .QN(n13395) );
  NAND2X0 U13310 ( .IN1(n13403), .IN2(n13404), .QN(g27323) );
  INVX0 U13311 ( .INP(n13405), .ZN(n13404) );
  NOR2X0 U13312 ( .IN1(n13355), .IN2(n8637), .QN(n13405) );
  NAND2X0 U13313 ( .IN1(n13355), .IN2(n13359), .QN(n13403) );
  NAND2X0 U13314 ( .IN1(n13406), .IN2(n13407), .QN(g27322) );
  NAND2X0 U13315 ( .IN1(n13408), .IN2(n13325), .QN(n13407) );
  NAND2X0 U13316 ( .IN1(n13324), .IN2(g2436), .QN(n13406) );
  NAND2X0 U13317 ( .IN1(n13409), .IN2(n13410), .QN(g27321) );
  NAND2X0 U13318 ( .IN1(n13364), .IN2(g1962), .QN(n13410) );
  NAND2X0 U13319 ( .IN1(n13362), .IN2(n13334), .QN(n13409) );
  INVX0 U13320 ( .INP(n13411), .ZN(n13334) );
  NAND2X0 U13321 ( .IN1(n13412), .IN2(n13413), .QN(n13411) );
  NAND2X0 U13322 ( .IN1(n12840), .IN2(n13414), .QN(n13413) );
  NOR2X0 U13323 ( .IN1(n12812), .IN2(n13415), .QN(n12840) );
  NAND2X0 U13324 ( .IN1(n13363), .IN2(n12812), .QN(n13412) );
  NAND2X0 U13325 ( .IN1(n13416), .IN2(n13417), .QN(g27320) );
  NAND2X0 U13326 ( .IN1(n13329), .IN2(g1960), .QN(n13417) );
  NAND2X0 U13327 ( .IN1(n13370), .IN2(n13330), .QN(n13416) );
  NAND2X0 U13328 ( .IN1(n13418), .IN2(n13419), .QN(g27319) );
  INVX0 U13329 ( .INP(n13420), .ZN(n13419) );
  NOR2X0 U13330 ( .IN1(n13309), .IN2(n8568), .QN(n13420) );
  NAND2X0 U13331 ( .IN1(n13421), .IN2(n13309), .QN(n13418) );
  NOR2X0 U13332 ( .IN1(n13422), .IN2(n4366), .QN(n13309) );
  INVX0 U13333 ( .INP(g22651), .ZN(n13422) );
  NAND2X0 U13334 ( .IN1(n13423), .IN2(n13424), .QN(g27318) );
  NAND2X0 U13335 ( .IN1(n13425), .IN2(n13375), .QN(n13424) );
  NAND2X0 U13336 ( .IN1(test_so58), .IN2(n13426), .QN(n13423) );
  NAND2X0 U13337 ( .IN1(n13427), .IN2(n13428), .QN(g27317) );
  NAND2X0 U13338 ( .IN1(n13373), .IN2(g1757), .QN(n13428) );
  NAND2X0 U13339 ( .IN1(n13374), .IN2(n13429), .QN(n13427) );
  NAND2X0 U13340 ( .IN1(n13430), .IN2(n13431), .QN(g27316) );
  NAND2X0 U13341 ( .IN1(n13432), .IN2(n13339), .QN(n13431) );
  NAND2X0 U13342 ( .IN1(n12956), .IN2(n13433), .QN(n13339) );
  NOR2X0 U13343 ( .IN1(n12930), .IN2(n12935), .QN(n12956) );
  INVX0 U13344 ( .INP(n13434), .ZN(n13430) );
  NOR2X0 U13345 ( .IN1(n13432), .IN2(n8604), .QN(n13434) );
  NAND2X0 U13346 ( .IN1(n13435), .IN2(n13436), .QN(g27315) );
  NAND2X0 U13347 ( .IN1(n13378), .IN2(g1269), .QN(n13436) );
  NAND2X0 U13348 ( .IN1(n13379), .IN2(n13382), .QN(n13435) );
  NAND2X0 U13349 ( .IN1(n13437), .IN2(n13438), .QN(g27314) );
  NAND2X0 U13350 ( .IN1(n13337), .IN2(g1264), .QN(n13438) );
  NAND2X0 U13351 ( .IN1(n13439), .IN2(n13338), .QN(n13437) );
  NAND2X0 U13352 ( .IN1(n13440), .IN2(n13441), .QN(g27313) );
  INVX0 U13353 ( .INP(n13442), .ZN(n13441) );
  NOR2X0 U13354 ( .IN1(n13443), .IN2(n8919), .QN(n13442) );
  NAND2X0 U13355 ( .IN1(n13443), .IN2(n13444), .QN(n13440) );
  NAND2X0 U13356 ( .IN1(n13445), .IN2(n13446), .QN(g27312) );
  NAND2X0 U13357 ( .IN1(n13447), .IN2(n13387), .QN(n13446) );
  INVX0 U13358 ( .INP(n13448), .ZN(n13445) );
  NOR2X0 U13359 ( .IN1(n13447), .IN2(n8609), .QN(n13448) );
  NAND2X0 U13360 ( .IN1(n13449), .IN2(n13450), .QN(g27311) );
  NAND2X0 U13361 ( .IN1(n13385), .IN2(g581), .QN(n13450) );
  NAND2X0 U13362 ( .IN1(n13386), .IN2(n13451), .QN(n13449) );
  NAND2X0 U13363 ( .IN1(n13452), .IN2(n13453), .QN(g27310) );
  NAND2X0 U13364 ( .IN1(n13315), .IN2(g2650), .QN(n13453) );
  NAND2X0 U13365 ( .IN1(n13352), .IN2(n13313), .QN(n13452) );
  INVX0 U13366 ( .INP(n13315), .ZN(n13313) );
  NAND2X0 U13367 ( .IN1(g7302), .IN2(g22687), .QN(n13315) );
  INVX0 U13368 ( .INP(n13454), .ZN(n13352) );
  NAND2X0 U13369 ( .IN1(n13455), .IN2(n13456), .QN(n13454) );
  NAND2X0 U13370 ( .IN1(g3229), .IN2(n13346), .QN(n13456) );
  NOR2X0 U13371 ( .IN1(n13457), .IN2(n13458), .QN(n13455) );
  NOR2X0 U13372 ( .IN1(n13390), .IN2(n13459), .QN(n13458) );
  NAND2X0 U13373 ( .IN1(n12668), .IN2(n12661), .QN(n13459) );
  NAND2X0 U13374 ( .IN1(n13460), .IN2(n13461), .QN(n12661) );
  NAND2X0 U13375 ( .IN1(n8566), .IN2(g7390), .QN(n13461) );
  NOR2X0 U13376 ( .IN1(n13462), .IN2(n13463), .QN(n13460) );
  NOR2X0 U13377 ( .IN1(n4314), .IN2(g2650), .QN(n13463) );
  NOR2X0 U13378 ( .IN1(n4299), .IN2(g2649), .QN(n13462) );
  INVX0 U13379 ( .INP(n13346), .ZN(n12668) );
  NAND2X0 U13380 ( .IN1(n13464), .IN2(n13465), .QN(n13346) );
  NAND2X0 U13381 ( .IN1(n8601), .IN2(g7390), .QN(n13465) );
  NOR2X0 U13382 ( .IN1(n13466), .IN2(n13467), .QN(n13464) );
  NOR2X0 U13383 ( .IN1(n4314), .IN2(g2659), .QN(n13467) );
  NOR2X0 U13384 ( .IN1(n4299), .IN2(g2658), .QN(n13466) );
  INVX0 U13385 ( .INP(n13468), .ZN(n13457) );
  NAND2X0 U13386 ( .IN1(n10022), .IN2(n13390), .QN(n13468) );
  NOR2X0 U13387 ( .IN1(n12676), .IN2(n12674), .QN(n13390) );
  INVX0 U13388 ( .INP(n12681), .ZN(n12674) );
  NAND2X0 U13389 ( .IN1(n13469), .IN2(n13470), .QN(n12681) );
  NAND2X0 U13390 ( .IN1(n8586), .IN2(g7390), .QN(n13470) );
  NOR2X0 U13391 ( .IN1(n13471), .IN2(n13472), .QN(n13469) );
  NOR2X0 U13392 ( .IN1(n4314), .IN2(g2653), .QN(n13472) );
  NOR2X0 U13393 ( .IN1(n4299), .IN2(g2652), .QN(n13471) );
  INVX0 U13394 ( .INP(n12666), .ZN(n12676) );
  NOR2X0 U13395 ( .IN1(n13473), .IN2(n13474), .QN(n12666) );
  NOR2X0 U13396 ( .IN1(n4370), .IN2(test_so89), .QN(n13474) );
  INVX0 U13397 ( .INP(n13475), .ZN(n13473) );
  NOR2X0 U13398 ( .IN1(n13476), .IN2(n13477), .QN(n13475) );
  NOR2X0 U13399 ( .IN1(n4314), .IN2(g2656), .QN(n13477) );
  NOR2X0 U13400 ( .IN1(n4299), .IN2(g2655), .QN(n13476) );
  NAND2X0 U13401 ( .IN1(n13478), .IN2(n13479), .QN(g27309) );
  NAND2X0 U13402 ( .IN1(n13402), .IN2(g2459), .QN(n13479) );
  NAND2X0 U13403 ( .IN1(n13397), .IN2(n13359), .QN(n13478) );
  INVX0 U13404 ( .INP(n13480), .ZN(n13359) );
  NAND2X0 U13405 ( .IN1(n13481), .IN2(n13482), .QN(n13480) );
  NAND2X0 U13406 ( .IN1(n13483), .IN2(n13400), .QN(n13482) );
  NAND2X0 U13407 ( .IN1(n13484), .IN2(n13485), .QN(n13481) );
  NOR2X0 U13408 ( .IN1(n13483), .IN2(n13486), .QN(n13484) );
  INVX0 U13409 ( .INP(n13401), .ZN(n13483) );
  XNOR2X1 U13410 ( .IN1(n13487), .IN2(n10022), .Q(n13401) );
  NAND2X0 U13411 ( .IN1(n13488), .IN2(n13489), .QN(g27308) );
  NAND2X0 U13412 ( .IN1(n13408), .IN2(n13355), .QN(n13489) );
  INVX0 U13413 ( .INP(n13490), .ZN(n13488) );
  NOR2X0 U13414 ( .IN1(n13355), .IN2(n8903), .QN(n13490) );
  NAND2X0 U13415 ( .IN1(n13491), .IN2(n13492), .QN(g27307) );
  NAND2X0 U13416 ( .IN1(n13324), .IN2(g2421), .QN(n13492) );
  INVX0 U13417 ( .INP(n13325), .ZN(n13324) );
  NAND2X0 U13418 ( .IN1(n13493), .IN2(n13325), .QN(n13491) );
  NOR2X0 U13419 ( .IN1(n13494), .IN2(n4509), .QN(n13325) );
  NAND2X0 U13420 ( .IN1(n13495), .IN2(n13496), .QN(g27306) );
  NAND2X0 U13421 ( .IN1(n13364), .IN2(g1959), .QN(n13496) );
  NAND2X0 U13422 ( .IN1(n13370), .IN2(n13362), .QN(n13495) );
  NOR2X0 U13423 ( .IN1(n13497), .IN2(n13498), .QN(n13370) );
  NOR2X0 U13424 ( .IN1(n13363), .IN2(n12797), .QN(n13498) );
  INVX0 U13425 ( .INP(n12807), .ZN(n12797) );
  INVX0 U13426 ( .INP(n13414), .ZN(n13363) );
  XNOR2X1 U13427 ( .IN1(n12783), .IN2(n10022), .Q(n13414) );
  INVX0 U13428 ( .INP(n12792), .ZN(n12783) );
  NAND2X0 U13429 ( .IN1(n13499), .IN2(n13500), .QN(g27305) );
  NAND2X0 U13430 ( .IN1(n13329), .IN2(g1957), .QN(n13500) );
  NAND2X0 U13431 ( .IN1(n13421), .IN2(n13330), .QN(n13499) );
  INVX0 U13432 ( .INP(n13329), .ZN(n13330) );
  NAND2X0 U13433 ( .IN1(g22651), .IN2(g7194), .QN(n13329) );
  NAND2X0 U13434 ( .IN1(n13501), .IN2(n13502), .QN(g27304) );
  NAND2X0 U13435 ( .IN1(n13503), .IN2(n13375), .QN(n13502) );
  NAND2X0 U13436 ( .IN1(n13504), .IN2(n13505), .QN(n13375) );
  NOR2X0 U13437 ( .IN1(n13506), .IN2(n13507), .QN(n13504) );
  NAND2X0 U13438 ( .IN1(n13508), .IN2(g1779), .QN(n13501) );
  NAND2X0 U13439 ( .IN1(n13509), .IN2(n13510), .QN(g27303) );
  INVX0 U13440 ( .INP(n13511), .ZN(n13510) );
  NOR2X0 U13441 ( .IN1(n13425), .IN2(n8640), .QN(n13511) );
  NAND2X0 U13442 ( .IN1(n13425), .IN2(n13429), .QN(n13509) );
  NAND2X0 U13443 ( .IN1(n13512), .IN2(n13513), .QN(g27302) );
  NAND2X0 U13444 ( .IN1(n13514), .IN2(n13374), .QN(n13513) );
  NAND2X0 U13445 ( .IN1(n13373), .IN2(g1742), .QN(n13512) );
  NAND2X0 U13446 ( .IN1(n13515), .IN2(n13516), .QN(g27301) );
  INVX0 U13447 ( .INP(n13517), .ZN(n13516) );
  NOR2X0 U13448 ( .IN1(n13432), .IN2(n8397), .QN(n13517) );
  NAND2X0 U13449 ( .IN1(n13432), .IN2(n13382), .QN(n13515) );
  INVX0 U13450 ( .INP(n13518), .ZN(n13382) );
  NAND2X0 U13451 ( .IN1(n13519), .IN2(n13520), .QN(n13518) );
  NAND2X0 U13452 ( .IN1(n12963), .IN2(n13521), .QN(n13520) );
  NOR2X0 U13453 ( .IN1(n12935), .IN2(n13522), .QN(n12963) );
  NAND2X0 U13454 ( .IN1(n13433), .IN2(n12935), .QN(n13519) );
  NAND2X0 U13455 ( .IN1(n13523), .IN2(n13524), .QN(g27300) );
  NAND2X0 U13456 ( .IN1(n13378), .IN2(g1266), .QN(n13524) );
  NAND2X0 U13457 ( .IN1(n13439), .IN2(n13379), .QN(n13523) );
  NAND2X0 U13458 ( .IN1(n13525), .IN2(n13526), .QN(g27299) );
  NAND2X0 U13459 ( .IN1(n13337), .IN2(g1261), .QN(n13526) );
  INVX0 U13460 ( .INP(n13338), .ZN(n13337) );
  NAND2X0 U13461 ( .IN1(n13527), .IN2(n13338), .QN(n13525) );
  NOR2X0 U13462 ( .IN1(n13528), .IN2(n4300), .QN(n13338) );
  NAND2X0 U13463 ( .IN1(n13529), .IN2(n13530), .QN(g27298) );
  NAND2X0 U13464 ( .IN1(n13531), .IN2(n13444), .QN(n13530) );
  NAND2X0 U13465 ( .IN1(n13532), .IN2(g1075), .QN(n13529) );
  NAND2X0 U13466 ( .IN1(n13533), .IN2(n13534), .QN(g27297) );
  INVX0 U13467 ( .INP(n13535), .ZN(n13534) );
  NOR2X0 U13468 ( .IN1(n13443), .IN2(n8642), .QN(n13535) );
  NAND2X0 U13469 ( .IN1(n13443), .IN2(n13536), .QN(n13533) );
  NAND2X0 U13470 ( .IN1(n13537), .IN2(n13538), .QN(g27296) );
  NAND2X0 U13471 ( .IN1(n13539), .IN2(n13387), .QN(n13538) );
  NAND2X0 U13472 ( .IN1(n13075), .IN2(n13540), .QN(n13387) );
  NOR2X0 U13473 ( .IN1(n13049), .IN2(n13054), .QN(n13075) );
  NAND2X0 U13474 ( .IN1(n13541), .IN2(g585), .QN(n13537) );
  NAND2X0 U13475 ( .IN1(n13542), .IN2(n13543), .QN(g27295) );
  INVX0 U13476 ( .INP(n13544), .ZN(n13543) );
  NOR2X0 U13477 ( .IN1(n13447), .IN2(n8401), .QN(n13544) );
  NAND2X0 U13478 ( .IN1(n13447), .IN2(n13451), .QN(n13542) );
  NAND2X0 U13479 ( .IN1(n13545), .IN2(n13546), .QN(g27294) );
  NAND2X0 U13480 ( .IN1(n13385), .IN2(g578), .QN(n13546) );
  NAND2X0 U13481 ( .IN1(n13547), .IN2(n13386), .QN(n13545) );
  NAND2X0 U13482 ( .IN1(n13548), .IN2(n13549), .QN(g27293) );
  NAND2X0 U13483 ( .IN1(n13550), .IN2(g391), .QN(n13549) );
  NAND2X0 U13484 ( .IN1(n13551), .IN2(n13552), .QN(n13548) );
  NAND2X0 U13485 ( .IN1(n13553), .IN2(n13554), .QN(g27292) );
  NAND2X0 U13486 ( .IN1(n13408), .IN2(n13397), .QN(n13554) );
  INVX0 U13487 ( .INP(n13555), .ZN(n13408) );
  NAND2X0 U13488 ( .IN1(n13556), .IN2(n13557), .QN(n13555) );
  NAND2X0 U13489 ( .IN1(n13558), .IN2(n13487), .QN(n13557) );
  INVX0 U13490 ( .INP(n13559), .ZN(n13487) );
  NOR2X0 U13491 ( .IN1(g3229), .IN2(n13399), .QN(n13558) );
  INVX0 U13492 ( .INP(n13560), .ZN(n13399) );
  NOR2X0 U13493 ( .IN1(n13561), .IN2(n13562), .QN(n13556) );
  NAND2X0 U13494 ( .IN1(n13402), .IN2(g2444), .QN(n13553) );
  NAND2X0 U13495 ( .IN1(n13563), .IN2(n13564), .QN(g27291) );
  INVX0 U13496 ( .INP(n13565), .ZN(n13564) );
  NOR2X0 U13497 ( .IN1(n13355), .IN2(n8926), .QN(n13565) );
  NAND2X0 U13498 ( .IN1(n13493), .IN2(n13355), .QN(n13563) );
  NOR2X0 U13499 ( .IN1(n13494), .IN2(n12443), .QN(n13355) );
  INVX0 U13500 ( .INP(n13566), .ZN(n13494) );
  NAND2X0 U13501 ( .IN1(n13567), .IN2(n13568), .QN(g27290) );
  NAND2X0 U13502 ( .IN1(n13364), .IN2(g1956), .QN(n13568) );
  NAND2X0 U13503 ( .IN1(n13421), .IN2(n13362), .QN(n13567) );
  INVX0 U13504 ( .INP(n13364), .ZN(n13362) );
  NAND2X0 U13505 ( .IN1(g7052), .IN2(g22651), .QN(n13364) );
  INVX0 U13506 ( .INP(n13569), .ZN(n13421) );
  NAND2X0 U13507 ( .IN1(n13570), .IN2(n13571), .QN(n13569) );
  NAND2X0 U13508 ( .IN1(g3229), .IN2(n13415), .QN(n13571) );
  NOR2X0 U13509 ( .IN1(n13572), .IN2(n13573), .QN(n13570) );
  NOR2X0 U13510 ( .IN1(n13497), .IN2(n13574), .QN(n13573) );
  NAND2X0 U13511 ( .IN1(n12799), .IN2(n12792), .QN(n13574) );
  NAND2X0 U13512 ( .IN1(n13575), .IN2(n13576), .QN(n12792) );
  NAND2X0 U13513 ( .IN1(n8568), .IN2(g1930), .QN(n13576) );
  NOR2X0 U13514 ( .IN1(n13577), .IN2(n13578), .QN(n13575) );
  NOR2X0 U13515 ( .IN1(n4315), .IN2(g1957), .QN(n13578) );
  NOR2X0 U13516 ( .IN1(n4296), .IN2(g1956), .QN(n13577) );
  INVX0 U13517 ( .INP(n13415), .ZN(n12799) );
  NAND2X0 U13518 ( .IN1(n13579), .IN2(n13580), .QN(n13415) );
  NAND2X0 U13519 ( .IN1(n8602), .IN2(g1930), .QN(n13580) );
  NOR2X0 U13520 ( .IN1(n13581), .IN2(n13582), .QN(n13579) );
  NOR2X0 U13521 ( .IN1(n4315), .IN2(g1966), .QN(n13582) );
  NOR2X0 U13522 ( .IN1(test_so67), .IN2(n4296), .QN(n13581) );
  INVX0 U13523 ( .INP(n13583), .ZN(n13572) );
  NAND2X0 U13524 ( .IN1(n10022), .IN2(n13497), .QN(n13583) );
  NOR2X0 U13525 ( .IN1(n12807), .IN2(n12805), .QN(n13497) );
  INVX0 U13526 ( .INP(n12812), .ZN(n12805) );
  NAND2X0 U13527 ( .IN1(n13584), .IN2(n13585), .QN(n12812) );
  NAND2X0 U13528 ( .IN1(n8588), .IN2(g1930), .QN(n13585) );
  NOR2X0 U13529 ( .IN1(n13586), .IN2(n13587), .QN(n13584) );
  NOR2X0 U13530 ( .IN1(n4315), .IN2(g1960), .QN(n13587) );
  NOR2X0 U13531 ( .IN1(n4296), .IN2(g1959), .QN(n13586) );
  NAND2X0 U13532 ( .IN1(n13588), .IN2(n13589), .QN(n12807) );
  NAND2X0 U13533 ( .IN1(n8395), .IN2(g1930), .QN(n13589) );
  NOR2X0 U13534 ( .IN1(n13590), .IN2(n13591), .QN(n13588) );
  NOR2X0 U13535 ( .IN1(n4315), .IN2(g1963), .QN(n13591) );
  NOR2X0 U13536 ( .IN1(n4296), .IN2(g1962), .QN(n13590) );
  NAND2X0 U13537 ( .IN1(n13592), .IN2(n13593), .QN(g27289) );
  NAND2X0 U13538 ( .IN1(n13508), .IN2(g1765), .QN(n13593) );
  NAND2X0 U13539 ( .IN1(n13503), .IN2(n13429), .QN(n13592) );
  INVX0 U13540 ( .INP(n13594), .ZN(n13429) );
  NAND2X0 U13541 ( .IN1(n13595), .IN2(n13596), .QN(n13594) );
  NAND2X0 U13542 ( .IN1(n13597), .IN2(n13506), .QN(n13596) );
  NAND2X0 U13543 ( .IN1(n13598), .IN2(n13599), .QN(n13595) );
  NOR2X0 U13544 ( .IN1(n13597), .IN2(n13600), .QN(n13598) );
  INVX0 U13545 ( .INP(n13507), .ZN(n13597) );
  XNOR2X1 U13546 ( .IN1(n13601), .IN2(n10022), .Q(n13507) );
  NAND2X0 U13547 ( .IN1(n13602), .IN2(n13603), .QN(g27288) );
  NAND2X0 U13548 ( .IN1(n13514), .IN2(n13425), .QN(n13603) );
  INVX0 U13549 ( .INP(n13604), .ZN(n13602) );
  NOR2X0 U13550 ( .IN1(n13425), .IN2(n8906), .QN(n13604) );
  NAND2X0 U13551 ( .IN1(n13605), .IN2(n13606), .QN(g27287) );
  NAND2X0 U13552 ( .IN1(n13373), .IN2(g1727), .QN(n13606) );
  NAND2X0 U13553 ( .IN1(n13607), .IN2(n13374), .QN(n13605) );
  INVX0 U13554 ( .INP(n13373), .ZN(n13374) );
  NAND2X0 U13555 ( .IN1(n13608), .IN2(n11849), .QN(n13373) );
  NAND2X0 U13556 ( .IN1(n13609), .IN2(n13610), .QN(g27286) );
  INVX0 U13557 ( .INP(n13611), .ZN(n13610) );
  NOR2X0 U13558 ( .IN1(n13432), .IN2(n8590), .QN(n13611) );
  NAND2X0 U13559 ( .IN1(n13439), .IN2(n13432), .QN(n13609) );
  NOR2X0 U13560 ( .IN1(n13612), .IN2(n13613), .QN(n13439) );
  NOR2X0 U13561 ( .IN1(n13433), .IN2(n12920), .QN(n13613) );
  INVX0 U13562 ( .INP(n12930), .ZN(n12920) );
  INVX0 U13563 ( .INP(n13521), .ZN(n13433) );
  XNOR2X1 U13564 ( .IN1(n12906), .IN2(n10022), .Q(n13521) );
  INVX0 U13565 ( .INP(n12915), .ZN(n12906) );
  NAND2X0 U13566 ( .IN1(n13614), .IN2(n13615), .QN(g27285) );
  NAND2X0 U13567 ( .IN1(n13378), .IN2(g1263), .QN(n13615) );
  INVX0 U13568 ( .INP(n13379), .ZN(n13378) );
  NAND2X0 U13569 ( .IN1(n13527), .IN2(n13379), .QN(n13614) );
  NOR2X0 U13570 ( .IN1(n13528), .IN2(n4316), .QN(n13379) );
  NAND2X0 U13571 ( .IN1(n13616), .IN2(n13617), .QN(g27284) );
  NAND2X0 U13572 ( .IN1(n13618), .IN2(n13444), .QN(n13617) );
  NAND2X0 U13573 ( .IN1(n13619), .IN2(n13620), .QN(n13444) );
  NOR2X0 U13574 ( .IN1(n13621), .IN2(n13622), .QN(n13619) );
  NAND2X0 U13575 ( .IN1(n13623), .IN2(g1085), .QN(n13616) );
  NAND2X0 U13576 ( .IN1(n13624), .IN2(n13625), .QN(g27283) );
  NAND2X0 U13577 ( .IN1(n13532), .IN2(g1060), .QN(n13625) );
  NAND2X0 U13578 ( .IN1(n13531), .IN2(n13536), .QN(n13624) );
  NAND2X0 U13579 ( .IN1(n13626), .IN2(n13627), .QN(g27282) );
  NAND2X0 U13580 ( .IN1(n13628), .IN2(n13443), .QN(n13627) );
  INVX0 U13581 ( .INP(n13629), .ZN(n13626) );
  NOR2X0 U13582 ( .IN1(n13443), .IN2(n8908), .QN(n13629) );
  NAND2X0 U13583 ( .IN1(n13630), .IN2(n13631), .QN(g27281) );
  NAND2X0 U13584 ( .IN1(n13541), .IN2(g582), .QN(n13631) );
  NAND2X0 U13585 ( .IN1(n13539), .IN2(n13451), .QN(n13630) );
  INVX0 U13586 ( .INP(n13632), .ZN(n13451) );
  NAND2X0 U13587 ( .IN1(n13633), .IN2(n13634), .QN(n13632) );
  NAND2X0 U13588 ( .IN1(n13082), .IN2(n13635), .QN(n13634) );
  NOR2X0 U13589 ( .IN1(n13054), .IN2(n13636), .QN(n13082) );
  NAND2X0 U13590 ( .IN1(n13540), .IN2(n13054), .QN(n13633) );
  INVX0 U13591 ( .INP(n13047), .ZN(n13054) );
  NAND2X0 U13592 ( .IN1(n13637), .IN2(n13638), .QN(g27280) );
  NAND2X0 U13593 ( .IN1(test_so25), .IN2(n13639), .QN(n13638) );
  NAND2X0 U13594 ( .IN1(n13547), .IN2(n13447), .QN(n13637) );
  NAND2X0 U13595 ( .IN1(n13640), .IN2(n13641), .QN(g27279) );
  NAND2X0 U13596 ( .IN1(n13385), .IN2(g575), .QN(n13641) );
  NAND2X0 U13597 ( .IN1(n13642), .IN2(n13386), .QN(n13640) );
  INVX0 U13598 ( .INP(n13385), .ZN(n13386) );
  NAND2X0 U13599 ( .IN1(g550), .IN2(g22578), .QN(n13385) );
  NAND2X0 U13600 ( .IN1(n13643), .IN2(n13644), .QN(g27278) );
  NAND2X0 U13601 ( .IN1(n13645), .IN2(n13552), .QN(n13644) );
  NAND2X0 U13602 ( .IN1(n13646), .IN2(g388), .QN(n13643) );
  NAND2X0 U13603 ( .IN1(n13647), .IN2(n13648), .QN(g27277) );
  NAND2X0 U13604 ( .IN1(n13550), .IN2(g376), .QN(n13648) );
  NAND2X0 U13605 ( .IN1(n13551), .IN2(n13649), .QN(n13647) );
  NAND2X0 U13606 ( .IN1(n13650), .IN2(n13651), .QN(g27276) );
  NAND2X0 U13607 ( .IN1(n13402), .IN2(g2429), .QN(n13651) );
  NAND2X0 U13608 ( .IN1(n13493), .IN2(n13397), .QN(n13650) );
  INVX0 U13609 ( .INP(n13402), .ZN(n13397) );
  NAND2X0 U13610 ( .IN1(n13566), .IN2(g5555), .QN(n13402) );
  NOR2X0 U13611 ( .IN1(n13652), .IN2(n13653), .QN(n13566) );
  NOR2X0 U13612 ( .IN1(n9753), .IN2(n11503), .QN(n13653) );
  NOR2X0 U13613 ( .IN1(n13654), .IN2(n13655), .QN(n13493) );
  NAND2X0 U13614 ( .IN1(n13656), .IN2(n13657), .QN(n13655) );
  NAND2X0 U13615 ( .IN1(n10022), .IN2(n13561), .QN(n13657) );
  NOR2X0 U13616 ( .IN1(n13560), .IN2(n13485), .QN(n13561) );
  INVX0 U13617 ( .INP(n13400), .ZN(n13485) );
  NAND2X0 U13618 ( .IN1(n13486), .IN2(g3229), .QN(n13656) );
  INVX0 U13619 ( .INP(n13658), .ZN(n13654) );
  NOR2X0 U13620 ( .IN1(n13562), .IN2(n13659), .QN(n13658) );
  NOR2X0 U13621 ( .IN1(n13486), .IN2(n13660), .QN(n13659) );
  NAND2X0 U13622 ( .IN1(n13661), .IN2(n13559), .QN(n13660) );
  NAND2X0 U13623 ( .IN1(g3229), .IN2(n13400), .QN(n13661) );
  NAND2X0 U13624 ( .IN1(n13662), .IN2(n13663), .QN(n13400) );
  NAND2X0 U13625 ( .IN1(n8903), .IN2(n10669), .QN(n13663) );
  NOR2X0 U13626 ( .IN1(n13664), .IN2(n13665), .QN(n13662) );
  NOR2X0 U13627 ( .IN1(n4516), .IN2(g2444), .QN(n13665) );
  NOR2X0 U13628 ( .IN1(n4509), .IN2(g2436), .QN(n13664) );
  NAND2X0 U13629 ( .IN1(n13666), .IN2(n13667), .QN(n13486) );
  NAND2X0 U13630 ( .IN1(n8915), .IN2(n10669), .QN(n13667) );
  NOR2X0 U13631 ( .IN1(n13668), .IN2(n13669), .QN(n13666) );
  NOR2X0 U13632 ( .IN1(n4516), .IN2(g2473), .QN(n13669) );
  NOR2X0 U13633 ( .IN1(n4509), .IN2(g2466), .QN(n13668) );
  NOR2X0 U13634 ( .IN1(n13670), .IN2(n10022), .QN(n13562) );
  NAND2X0 U13635 ( .IN1(n13560), .IN2(n13559), .QN(n13670) );
  NAND2X0 U13636 ( .IN1(n13671), .IN2(n13672), .QN(n13559) );
  NAND2X0 U13637 ( .IN1(n8926), .IN2(n10669), .QN(n13672) );
  NOR2X0 U13638 ( .IN1(n13673), .IN2(n13674), .QN(n13671) );
  NOR2X0 U13639 ( .IN1(n4516), .IN2(g2429), .QN(n13674) );
  NOR2X0 U13640 ( .IN1(n4509), .IN2(g2421), .QN(n13673) );
  NAND2X0 U13641 ( .IN1(n13675), .IN2(n13676), .QN(n13560) );
  NAND2X0 U13642 ( .IN1(n8637), .IN2(n10669), .QN(n13676) );
  NOR2X0 U13643 ( .IN1(n13677), .IN2(n13678), .QN(n13675) );
  NOR2X0 U13644 ( .IN1(n4516), .IN2(g2459), .QN(n13678) );
  NOR2X0 U13645 ( .IN1(n4509), .IN2(g2451), .QN(n13677) );
  NAND2X0 U13646 ( .IN1(n13679), .IN2(n13680), .QN(g27275) );
  NAND2X0 U13647 ( .IN1(n13514), .IN2(n13503), .QN(n13680) );
  INVX0 U13648 ( .INP(n13681), .ZN(n13514) );
  NAND2X0 U13649 ( .IN1(n13682), .IN2(n13683), .QN(n13681) );
  NAND2X0 U13650 ( .IN1(n13684), .IN2(n13601), .QN(n13683) );
  INVX0 U13651 ( .INP(n13685), .ZN(n13601) );
  NOR2X0 U13652 ( .IN1(g3229), .IN2(n13505), .QN(n13684) );
  INVX0 U13653 ( .INP(n13686), .ZN(n13505) );
  NOR2X0 U13654 ( .IN1(n13687), .IN2(n13688), .QN(n13682) );
  NAND2X0 U13655 ( .IN1(n13508), .IN2(g1750), .QN(n13679) );
  NAND2X0 U13656 ( .IN1(n13689), .IN2(n13690), .QN(g27274) );
  INVX0 U13657 ( .INP(n13691), .ZN(n13690) );
  NOR2X0 U13658 ( .IN1(n13425), .IN2(n8929), .QN(n13691) );
  NAND2X0 U13659 ( .IN1(n13607), .IN2(n13425), .QN(n13689) );
  INVX0 U13660 ( .INP(n13426), .ZN(n13425) );
  NAND2X0 U13661 ( .IN1(n13608), .IN2(g7014), .QN(n13426) );
  NAND2X0 U13662 ( .IN1(n13692), .IN2(n13693), .QN(g27273) );
  INVX0 U13663 ( .INP(n13694), .ZN(n13693) );
  NOR2X0 U13664 ( .IN1(n13432), .IN2(n8570), .QN(n13694) );
  NAND2X0 U13665 ( .IN1(n13527), .IN2(n13432), .QN(n13692) );
  NOR2X0 U13666 ( .IN1(n13695), .IN2(n13528), .QN(n13432) );
  INVX0 U13667 ( .INP(g22615), .ZN(n13528) );
  INVX0 U13668 ( .INP(n13696), .ZN(n13527) );
  NAND2X0 U13669 ( .IN1(n13697), .IN2(n13698), .QN(n13696) );
  NAND2X0 U13670 ( .IN1(g3229), .IN2(n13522), .QN(n13698) );
  NOR2X0 U13671 ( .IN1(n13699), .IN2(n13700), .QN(n13697) );
  NOR2X0 U13672 ( .IN1(n13612), .IN2(n13701), .QN(n13700) );
  NAND2X0 U13673 ( .IN1(n12922), .IN2(n12915), .QN(n13701) );
  NAND2X0 U13674 ( .IN1(n13702), .IN2(n13703), .QN(n12915) );
  NAND2X0 U13675 ( .IN1(n8570), .IN2(n12608), .QN(n13703) );
  NOR2X0 U13676 ( .IN1(n13704), .IN2(n13705), .QN(n13702) );
  NOR2X0 U13677 ( .IN1(n4316), .IN2(g1263), .QN(n13705) );
  NOR2X0 U13678 ( .IN1(n4300), .IN2(g1261), .QN(n13704) );
  INVX0 U13679 ( .INP(n13522), .ZN(n12922) );
  NAND2X0 U13680 ( .IN1(n13706), .IN2(n13707), .QN(n13522) );
  NAND2X0 U13681 ( .IN1(n8604), .IN2(n12608), .QN(n13707) );
  NOR2X0 U13682 ( .IN1(n13708), .IN2(n13709), .QN(n13706) );
  NOR2X0 U13683 ( .IN1(n4316), .IN2(g1272), .QN(n13709) );
  NOR2X0 U13684 ( .IN1(n4300), .IN2(g1270), .QN(n13708) );
  INVX0 U13685 ( .INP(n13710), .ZN(n13699) );
  NAND2X0 U13686 ( .IN1(n10022), .IN2(n13612), .QN(n13710) );
  NOR2X0 U13687 ( .IN1(n12930), .IN2(n12928), .QN(n13612) );
  INVX0 U13688 ( .INP(n12935), .ZN(n12928) );
  NAND2X0 U13689 ( .IN1(n13711), .IN2(n13712), .QN(n12935) );
  NAND2X0 U13690 ( .IN1(n8590), .IN2(n12608), .QN(n13712) );
  NOR2X0 U13691 ( .IN1(n13713), .IN2(n13714), .QN(n13711) );
  NOR2X0 U13692 ( .IN1(n4316), .IN2(g1266), .QN(n13714) );
  NOR2X0 U13693 ( .IN1(n4300), .IN2(g1264), .QN(n13713) );
  NAND2X0 U13694 ( .IN1(n13715), .IN2(n13716), .QN(n12930) );
  NAND2X0 U13695 ( .IN1(n8397), .IN2(n12608), .QN(n13716) );
  NOR2X0 U13696 ( .IN1(n13717), .IN2(n13718), .QN(n13715) );
  NOR2X0 U13697 ( .IN1(n4316), .IN2(g1269), .QN(n13718) );
  NOR2X0 U13698 ( .IN1(test_so46), .IN2(n4300), .QN(n13717) );
  NAND2X0 U13699 ( .IN1(n13719), .IN2(n13720), .QN(g27272) );
  NAND2X0 U13700 ( .IN1(test_so37), .IN2(n13623), .QN(n13720) );
  NAND2X0 U13701 ( .IN1(n13618), .IN2(n13536), .QN(n13719) );
  INVX0 U13702 ( .INP(n13721), .ZN(n13536) );
  NAND2X0 U13703 ( .IN1(n13722), .IN2(n13723), .QN(n13721) );
  NAND2X0 U13704 ( .IN1(n13724), .IN2(n13621), .QN(n13723) );
  NAND2X0 U13705 ( .IN1(n13725), .IN2(n13726), .QN(n13722) );
  NOR2X0 U13706 ( .IN1(n13724), .IN2(n13727), .QN(n13725) );
  INVX0 U13707 ( .INP(n13622), .ZN(n13724) );
  XNOR2X1 U13708 ( .IN1(n13728), .IN2(n10022), .Q(n13622) );
  NAND2X0 U13709 ( .IN1(n13729), .IN2(n13730), .QN(g27271) );
  NAND2X0 U13710 ( .IN1(n13628), .IN2(n13531), .QN(n13730) );
  NAND2X0 U13711 ( .IN1(n13532), .IN2(g1045), .QN(n13729) );
  NAND2X0 U13712 ( .IN1(n13731), .IN2(n13732), .QN(g27270) );
  INVX0 U13713 ( .INP(n13733), .ZN(n13732) );
  NOR2X0 U13714 ( .IN1(n13443), .IN2(n8931), .QN(n13733) );
  NAND2X0 U13715 ( .IN1(n13734), .IN2(n13443), .QN(n13731) );
  NOR2X0 U13716 ( .IN1(n13735), .IN2(n4381), .QN(n13443) );
  NAND2X0 U13717 ( .IN1(n13736), .IN2(n13737), .QN(g27269) );
  NAND2X0 U13718 ( .IN1(n13541), .IN2(g579), .QN(n13737) );
  NAND2X0 U13719 ( .IN1(n13547), .IN2(n13539), .QN(n13736) );
  NOR2X0 U13720 ( .IN1(n13738), .IN2(n13739), .QN(n13547) );
  NOR2X0 U13721 ( .IN1(n13540), .IN2(n13039), .QN(n13739) );
  INVX0 U13722 ( .INP(n13049), .ZN(n13039) );
  INVX0 U13723 ( .INP(n13635), .ZN(n13540) );
  XNOR2X1 U13724 ( .IN1(n13025), .IN2(n10022), .Q(n13635) );
  INVX0 U13725 ( .INP(n13034), .ZN(n13025) );
  NAND2X0 U13726 ( .IN1(n13740), .IN2(n13741), .QN(g27268) );
  INVX0 U13727 ( .INP(n13742), .ZN(n13741) );
  NOR2X0 U13728 ( .IN1(n13447), .IN2(n8575), .QN(n13742) );
  NAND2X0 U13729 ( .IN1(n13642), .IN2(n13447), .QN(n13740) );
  INVX0 U13730 ( .INP(n13639), .ZN(n13447) );
  NAND2X0 U13731 ( .IN1(g6642), .IN2(g22578), .QN(n13639) );
  NAND2X0 U13732 ( .IN1(n13743), .IN2(n13744), .QN(g27267) );
  NAND2X0 U13733 ( .IN1(n13745), .IN2(n13552), .QN(n13744) );
  NAND2X0 U13734 ( .IN1(n13746), .IN2(n13747), .QN(n13552) );
  NOR2X0 U13735 ( .IN1(n13748), .IN2(n13749), .QN(n13746) );
  INVX0 U13736 ( .INP(n13750), .ZN(n13743) );
  NOR2X0 U13737 ( .IN1(n13745), .IN2(n8924), .QN(n13750) );
  NAND2X0 U13738 ( .IN1(n13751), .IN2(n13752), .QN(g27266) );
  NAND2X0 U13739 ( .IN1(n13646), .IN2(g373), .QN(n13752) );
  NAND2X0 U13740 ( .IN1(n13645), .IN2(n13649), .QN(n13751) );
  NAND2X0 U13741 ( .IN1(n13753), .IN2(n13754), .QN(g27265) );
  NAND2X0 U13742 ( .IN1(n13755), .IN2(n13551), .QN(n13754) );
  NAND2X0 U13743 ( .IN1(n13550), .IN2(g361), .QN(n13753) );
  NAND2X0 U13744 ( .IN1(n13756), .IN2(n13757), .QN(g27264) );
  NAND2X0 U13745 ( .IN1(n13508), .IN2(g1735), .QN(n13757) );
  NAND2X0 U13746 ( .IN1(n13607), .IN2(n13503), .QN(n13756) );
  INVX0 U13747 ( .INP(n13508), .ZN(n13503) );
  NAND2X0 U13748 ( .IN1(n13608), .IN2(g5511), .QN(n13508) );
  NOR2X0 U13749 ( .IN1(n13758), .IN2(n13759), .QN(n13608) );
  NOR2X0 U13750 ( .IN1(n9753), .IN2(n11564), .QN(n13759) );
  INVX0 U13751 ( .INP(n13760), .ZN(n13607) );
  NAND2X0 U13752 ( .IN1(n13761), .IN2(n13762), .QN(n13760) );
  NOR2X0 U13753 ( .IN1(n13763), .IN2(n13764), .QN(n13762) );
  INVX0 U13754 ( .INP(n13765), .ZN(n13764) );
  NAND2X0 U13755 ( .IN1(n10022), .IN2(n13687), .QN(n13765) );
  NOR2X0 U13756 ( .IN1(n13686), .IN2(n13599), .QN(n13687) );
  INVX0 U13757 ( .INP(n13506), .ZN(n13599) );
  NOR2X0 U13758 ( .IN1(n13766), .IN2(n10022), .QN(n13763) );
  NOR2X0 U13759 ( .IN1(n13688), .IN2(n13767), .QN(n13761) );
  NOR2X0 U13760 ( .IN1(n13600), .IN2(n13768), .QN(n13767) );
  NAND2X0 U13761 ( .IN1(n13769), .IN2(n13685), .QN(n13768) );
  NAND2X0 U13762 ( .IN1(g3229), .IN2(n13506), .QN(n13769) );
  NAND2X0 U13763 ( .IN1(n13770), .IN2(n13771), .QN(n13506) );
  NAND2X0 U13764 ( .IN1(n8906), .IN2(n10678), .QN(n13771) );
  NOR2X0 U13765 ( .IN1(n13772), .IN2(n13773), .QN(n13770) );
  NOR2X0 U13766 ( .IN1(n4518), .IN2(g1750), .QN(n13773) );
  NOR2X0 U13767 ( .IN1(n4511), .IN2(g1742), .QN(n13772) );
  INVX0 U13768 ( .INP(n13766), .ZN(n13600) );
  NOR2X0 U13769 ( .IN1(n13774), .IN2(n13775), .QN(n13766) );
  NOR2X0 U13770 ( .IN1(n4525), .IN2(test_so58), .QN(n13775) );
  INVX0 U13771 ( .INP(n13776), .ZN(n13774) );
  NOR2X0 U13772 ( .IN1(n13777), .IN2(n13778), .QN(n13776) );
  NOR2X0 U13773 ( .IN1(n4518), .IN2(g1779), .QN(n13778) );
  NOR2X0 U13774 ( .IN1(n4511), .IN2(g1772), .QN(n13777) );
  NOR2X0 U13775 ( .IN1(n13779), .IN2(n10022), .QN(n13688) );
  NAND2X0 U13776 ( .IN1(n13686), .IN2(n13685), .QN(n13779) );
  NAND2X0 U13777 ( .IN1(n13780), .IN2(n13781), .QN(n13685) );
  NAND2X0 U13778 ( .IN1(n8929), .IN2(n10678), .QN(n13781) );
  NOR2X0 U13779 ( .IN1(n13782), .IN2(n13783), .QN(n13780) );
  NOR2X0 U13780 ( .IN1(n4518), .IN2(g1735), .QN(n13783) );
  NOR2X0 U13781 ( .IN1(n4511), .IN2(g1727), .QN(n13782) );
  NAND2X0 U13782 ( .IN1(n13784), .IN2(n13785), .QN(n13686) );
  NAND2X0 U13783 ( .IN1(n8640), .IN2(n10678), .QN(n13785) );
  NOR2X0 U13784 ( .IN1(n13786), .IN2(n13787), .QN(n13784) );
  NOR2X0 U13785 ( .IN1(n4518), .IN2(g1765), .QN(n13787) );
  NOR2X0 U13786 ( .IN1(n4511), .IN2(g1757), .QN(n13786) );
  NAND2X0 U13787 ( .IN1(n13788), .IN2(n13789), .QN(g27263) );
  NAND2X0 U13788 ( .IN1(n13628), .IN2(n13618), .QN(n13789) );
  INVX0 U13789 ( .INP(n13790), .ZN(n13628) );
  NAND2X0 U13790 ( .IN1(n13791), .IN2(n13792), .QN(n13790) );
  NAND2X0 U13791 ( .IN1(n13793), .IN2(n13728), .QN(n13792) );
  INVX0 U13792 ( .INP(n13794), .ZN(n13728) );
  NOR2X0 U13793 ( .IN1(g3229), .IN2(n13620), .QN(n13793) );
  INVX0 U13794 ( .INP(n13795), .ZN(n13620) );
  NOR2X0 U13795 ( .IN1(n13796), .IN2(n13797), .QN(n13791) );
  NAND2X0 U13796 ( .IN1(n13623), .IN2(g1056), .QN(n13788) );
  NAND2X0 U13797 ( .IN1(n13798), .IN2(n13799), .QN(g27262) );
  NAND2X0 U13798 ( .IN1(n13532), .IN2(g1030), .QN(n13799) );
  INVX0 U13799 ( .INP(n13531), .ZN(n13532) );
  NAND2X0 U13800 ( .IN1(n13734), .IN2(n13531), .QN(n13798) );
  NOR2X0 U13801 ( .IN1(n13735), .IN2(n4364), .QN(n13531) );
  NAND2X0 U13802 ( .IN1(n13800), .IN2(n13801), .QN(g27261) );
  NAND2X0 U13803 ( .IN1(n13541), .IN2(g576), .QN(n13801) );
  NAND2X0 U13804 ( .IN1(n13642), .IN2(n13539), .QN(n13800) );
  INVX0 U13805 ( .INP(n13541), .ZN(n13539) );
  NAND2X0 U13806 ( .IN1(g6485), .IN2(g22578), .QN(n13541) );
  INVX0 U13807 ( .INP(n13802), .ZN(n13642) );
  NAND2X0 U13808 ( .IN1(n13803), .IN2(n13804), .QN(n13802) );
  NAND2X0 U13809 ( .IN1(g3229), .IN2(n13636), .QN(n13804) );
  NOR2X0 U13810 ( .IN1(n13805), .IN2(n13806), .QN(n13803) );
  NOR2X0 U13811 ( .IN1(n13738), .IN2(n13807), .QN(n13806) );
  NAND2X0 U13812 ( .IN1(n13041), .IN2(n13034), .QN(n13807) );
  NAND2X0 U13813 ( .IN1(n13808), .IN2(n13809), .QN(n13034) );
  NAND2X0 U13814 ( .IN1(n8575), .IN2(g6642), .QN(n13809) );
  NOR2X0 U13815 ( .IN1(n13810), .IN2(n13811), .QN(n13808) );
  NOR2X0 U13816 ( .IN1(n4313), .IN2(g575), .QN(n13811) );
  NOR2X0 U13817 ( .IN1(n4298), .IN2(g576), .QN(n13810) );
  INVX0 U13818 ( .INP(n13636), .ZN(n13041) );
  NAND2X0 U13819 ( .IN1(n13812), .IN2(n13813), .QN(n13636) );
  NAND2X0 U13820 ( .IN1(n8609), .IN2(g6642), .QN(n13813) );
  NOR2X0 U13821 ( .IN1(n13814), .IN2(n13815), .QN(n13812) );
  NOR2X0 U13822 ( .IN1(n4313), .IN2(g584), .QN(n13815) );
  NOR2X0 U13823 ( .IN1(n4298), .IN2(g585), .QN(n13814) );
  INVX0 U13824 ( .INP(n13816), .ZN(n13805) );
  NAND2X0 U13825 ( .IN1(n10022), .IN2(n13738), .QN(n13816) );
  NOR2X0 U13826 ( .IN1(n13049), .IN2(n13047), .QN(n13738) );
  NOR2X0 U13827 ( .IN1(n13817), .IN2(n13818), .QN(n13047) );
  NOR2X0 U13828 ( .IN1(n4372), .IN2(test_so25), .QN(n13818) );
  INVX0 U13829 ( .INP(n13819), .ZN(n13817) );
  NOR2X0 U13830 ( .IN1(n13820), .IN2(n13821), .QN(n13819) );
  NOR2X0 U13831 ( .IN1(n4313), .IN2(g578), .QN(n13821) );
  NOR2X0 U13832 ( .IN1(n4298), .IN2(g579), .QN(n13820) );
  NAND2X0 U13833 ( .IN1(n13822), .IN2(n13823), .QN(n13049) );
  NAND2X0 U13834 ( .IN1(n8401), .IN2(g6642), .QN(n13823) );
  NOR2X0 U13835 ( .IN1(n13824), .IN2(n13825), .QN(n13822) );
  NOR2X0 U13836 ( .IN1(n4313), .IN2(g581), .QN(n13825) );
  NOR2X0 U13837 ( .IN1(n4298), .IN2(g582), .QN(n13824) );
  NAND2X0 U13838 ( .IN1(n13826), .IN2(n13827), .QN(g27260) );
  INVX0 U13839 ( .INP(n13828), .ZN(n13827) );
  NOR2X0 U13840 ( .IN1(n13745), .IN2(n8643), .QN(n13828) );
  NAND2X0 U13841 ( .IN1(n13745), .IN2(n13649), .QN(n13826) );
  INVX0 U13842 ( .INP(n13829), .ZN(n13649) );
  NAND2X0 U13843 ( .IN1(n13830), .IN2(n13831), .QN(n13829) );
  NAND2X0 U13844 ( .IN1(n13832), .IN2(n13748), .QN(n13831) );
  NAND2X0 U13845 ( .IN1(n13833), .IN2(n13834), .QN(n13830) );
  NOR2X0 U13846 ( .IN1(n13832), .IN2(n13835), .QN(n13833) );
  INVX0 U13847 ( .INP(n13749), .ZN(n13832) );
  XNOR2X1 U13848 ( .IN1(n13836), .IN2(n10022), .Q(n13749) );
  NAND2X0 U13849 ( .IN1(n13837), .IN2(n13838), .QN(g27259) );
  NAND2X0 U13850 ( .IN1(n13755), .IN2(n13645), .QN(n13838) );
  NAND2X0 U13851 ( .IN1(n13646), .IN2(g358), .QN(n13837) );
  NAND2X0 U13852 ( .IN1(n13839), .IN2(n13840), .QN(g27258) );
  NAND2X0 U13853 ( .IN1(test_so16), .IN2(n13550), .QN(n13840) );
  NAND2X0 U13854 ( .IN1(n13841), .IN2(n13551), .QN(n13839) );
  INVX0 U13855 ( .INP(n13550), .ZN(n13551) );
  NAND2X0 U13856 ( .IN1(n13842), .IN2(n11886), .QN(n13550) );
  NAND2X0 U13857 ( .IN1(n13843), .IN2(n13844), .QN(g27257) );
  NAND2X0 U13858 ( .IN1(n13623), .IN2(g1041), .QN(n13844) );
  INVX0 U13859 ( .INP(n13618), .ZN(n13623) );
  NAND2X0 U13860 ( .IN1(n13734), .IN2(n13618), .QN(n13843) );
  NOR2X0 U13861 ( .IN1(n13735), .IN2(n4363), .QN(n13618) );
  NAND2X0 U13862 ( .IN1(n9787), .IN2(n13845), .QN(n13735) );
  NAND2X0 U13863 ( .IN1(n13846), .IN2(n9764), .QN(n13845) );
  NOR2X0 U13864 ( .IN1(n13847), .IN2(n13848), .QN(n13734) );
  NAND2X0 U13865 ( .IN1(n13849), .IN2(n13850), .QN(n13848) );
  NAND2X0 U13866 ( .IN1(n10022), .IN2(n13796), .QN(n13850) );
  NOR2X0 U13867 ( .IN1(n13795), .IN2(n13726), .QN(n13796) );
  INVX0 U13868 ( .INP(n13621), .ZN(n13726) );
  NAND2X0 U13869 ( .IN1(n13727), .IN2(g3229), .QN(n13849) );
  INVX0 U13870 ( .INP(n13851), .ZN(n13847) );
  NOR2X0 U13871 ( .IN1(n13797), .IN2(n13852), .QN(n13851) );
  NOR2X0 U13872 ( .IN1(n13727), .IN2(n13853), .QN(n13852) );
  NAND2X0 U13873 ( .IN1(n13854), .IN2(n13794), .QN(n13853) );
  NAND2X0 U13874 ( .IN1(g3229), .IN2(n13621), .QN(n13854) );
  NAND2X0 U13875 ( .IN1(n13855), .IN2(n13856), .QN(n13621) );
  NAND2X0 U13876 ( .IN1(n8908), .IN2(g1088), .QN(n13856) );
  NOR2X0 U13877 ( .IN1(n13857), .IN2(n13858), .QN(n13855) );
  NOR2X0 U13878 ( .IN1(n4364), .IN2(g1045), .QN(n13858) );
  NOR2X0 U13879 ( .IN1(n4363), .IN2(g1056), .QN(n13857) );
  NAND2X0 U13880 ( .IN1(n13859), .IN2(n13860), .QN(n13727) );
  NAND2X0 U13881 ( .IN1(n8919), .IN2(g1088), .QN(n13860) );
  NOR2X0 U13882 ( .IN1(n13861), .IN2(n13862), .QN(n13859) );
  NOR2X0 U13883 ( .IN1(n4364), .IN2(g1075), .QN(n13862) );
  NOR2X0 U13884 ( .IN1(n4363), .IN2(g1085), .QN(n13861) );
  NOR2X0 U13885 ( .IN1(n13863), .IN2(n10022), .QN(n13797) );
  NAND2X0 U13886 ( .IN1(n13795), .IN2(n13794), .QN(n13863) );
  NAND2X0 U13887 ( .IN1(n13864), .IN2(n13865), .QN(n13794) );
  NAND2X0 U13888 ( .IN1(n8931), .IN2(g1088), .QN(n13865) );
  NOR2X0 U13889 ( .IN1(n13866), .IN2(n13867), .QN(n13864) );
  NOR2X0 U13890 ( .IN1(n4364), .IN2(g1030), .QN(n13867) );
  NOR2X0 U13891 ( .IN1(n4363), .IN2(g1041), .QN(n13866) );
  NAND2X0 U13892 ( .IN1(n13868), .IN2(n13869), .QN(n13795) );
  NAND2X0 U13893 ( .IN1(n8642), .IN2(g1088), .QN(n13869) );
  NOR2X0 U13894 ( .IN1(n13870), .IN2(n13871), .QN(n13868) );
  NOR2X0 U13895 ( .IN1(n4364), .IN2(g1060), .QN(n13871) );
  NOR2X0 U13896 ( .IN1(test_so37), .IN2(n4363), .QN(n13870) );
  NAND2X0 U13897 ( .IN1(n13872), .IN2(n13873), .QN(g27256) );
  NAND2X0 U13898 ( .IN1(n13755), .IN2(n13745), .QN(n13873) );
  INVX0 U13899 ( .INP(n13874), .ZN(n13755) );
  NAND2X0 U13900 ( .IN1(n13875), .IN2(n13876), .QN(n13874) );
  NAND2X0 U13901 ( .IN1(n13877), .IN2(n13836), .QN(n13876) );
  INVX0 U13902 ( .INP(n13878), .ZN(n13836) );
  NOR2X0 U13903 ( .IN1(g3229), .IN2(n13747), .QN(n13877) );
  INVX0 U13904 ( .INP(n13879), .ZN(n13747) );
  NOR2X0 U13905 ( .IN1(n13880), .IN2(n13881), .QN(n13875) );
  INVX0 U13906 ( .INP(n13882), .ZN(n13872) );
  NOR2X0 U13907 ( .IN1(n13745), .IN2(n8913), .QN(n13882) );
  NAND2X0 U13908 ( .IN1(n13883), .IN2(n13884), .QN(g27255) );
  NAND2X0 U13909 ( .IN1(n13646), .IN2(g343), .QN(n13884) );
  NAND2X0 U13910 ( .IN1(n13841), .IN2(n13645), .QN(n13883) );
  INVX0 U13911 ( .INP(n13646), .ZN(n13645) );
  NAND2X0 U13912 ( .IN1(n13842), .IN2(g6447), .QN(n13646) );
  NAND2X0 U13913 ( .IN1(n13885), .IN2(n13886), .QN(g27253) );
  INVX0 U13914 ( .INP(n13887), .ZN(n13886) );
  NOR2X0 U13915 ( .IN1(n13745), .IN2(n8935), .QN(n13887) );
  NAND2X0 U13916 ( .IN1(n13841), .IN2(n13745), .QN(n13885) );
  INVX0 U13917 ( .INP(n13888), .ZN(n13745) );
  NAND2X0 U13918 ( .IN1(n13842), .IN2(g5437), .QN(n13888) );
  NOR2X0 U13919 ( .IN1(n13889), .IN2(n13890), .QN(n13842) );
  NOR2X0 U13920 ( .IN1(n9753), .IN2(n11693), .QN(n13890) );
  NOR2X0 U13921 ( .IN1(n13891), .IN2(n13892), .QN(n13841) );
  NAND2X0 U13922 ( .IN1(n13893), .IN2(n13894), .QN(n13892) );
  NAND2X0 U13923 ( .IN1(n10022), .IN2(n13880), .QN(n13894) );
  NOR2X0 U13924 ( .IN1(n13879), .IN2(n13834), .QN(n13880) );
  INVX0 U13925 ( .INP(n13748), .ZN(n13834) );
  NAND2X0 U13926 ( .IN1(n13835), .IN2(g3229), .QN(n13893) );
  INVX0 U13927 ( .INP(n13895), .ZN(n13891) );
  NOR2X0 U13928 ( .IN1(n13881), .IN2(n13896), .QN(n13895) );
  NOR2X0 U13929 ( .IN1(n13835), .IN2(n13897), .QN(n13896) );
  NAND2X0 U13930 ( .IN1(n13898), .IN2(n13878), .QN(n13897) );
  NAND2X0 U13931 ( .IN1(g3229), .IN2(n13748), .QN(n13898) );
  NAND2X0 U13932 ( .IN1(n13899), .IN2(n13900), .QN(n13748) );
  NAND2X0 U13933 ( .IN1(n8913), .IN2(n10752), .QN(n13900) );
  NOR2X0 U13934 ( .IN1(n13901), .IN2(n13902), .QN(n13899) );
  NOR2X0 U13935 ( .IN1(n4506), .IN2(g361), .QN(n13902) );
  NOR2X0 U13936 ( .IN1(n4499), .IN2(g358), .QN(n13901) );
  NAND2X0 U13937 ( .IN1(n13903), .IN2(n13904), .QN(n13835) );
  NAND2X0 U13938 ( .IN1(n8924), .IN2(n10752), .QN(n13904) );
  NOR2X0 U13939 ( .IN1(n13905), .IN2(n13906), .QN(n13903) );
  NOR2X0 U13940 ( .IN1(n4506), .IN2(g391), .QN(n13906) );
  NOR2X0 U13941 ( .IN1(n4499), .IN2(g388), .QN(n13905) );
  NOR2X0 U13942 ( .IN1(n13907), .IN2(n10022), .QN(n13881) );
  NAND2X0 U13943 ( .IN1(n13879), .IN2(n13878), .QN(n13907) );
  NAND2X0 U13944 ( .IN1(n13908), .IN2(n13909), .QN(n13878) );
  NAND2X0 U13945 ( .IN1(n8935), .IN2(n10752), .QN(n13909) );
  NOR2X0 U13946 ( .IN1(n13910), .IN2(n13911), .QN(n13908) );
  NOR2X0 U13947 ( .IN1(test_so16), .IN2(n4506), .QN(n13911) );
  NOR2X0 U13948 ( .IN1(n4499), .IN2(g343), .QN(n13910) );
  NAND2X0 U13949 ( .IN1(n13912), .IN2(n13913), .QN(n13879) );
  NAND2X0 U13950 ( .IN1(n8643), .IN2(n10752), .QN(n13913) );
  NOR2X0 U13951 ( .IN1(n13914), .IN2(n13915), .QN(n13912) );
  NOR2X0 U13952 ( .IN1(n4506), .IN2(g376), .QN(n13915) );
  NOR2X0 U13953 ( .IN1(n4499), .IN2(g373), .QN(n13914) );
  NOR2X0 U13954 ( .IN1(n13916), .IN2(n13917), .QN(g27243) );
  NAND2X0 U13955 ( .IN1(n13918), .IN2(n10619), .QN(n13917) );
  NAND2X0 U13956 ( .IN1(n13919), .IN2(test_so92), .QN(n10619) );
  NOR2X0 U13957 ( .IN1(n4471), .IN2(n13920), .QN(n13919) );
  NOR2X0 U13958 ( .IN1(n13921), .IN2(g2753), .QN(n13916) );
  NOR2X0 U13959 ( .IN1(n13920), .IN2(n9282), .QN(n13921) );
  NOR2X0 U13960 ( .IN1(n13922), .IN2(n13260), .QN(g27123) );
  NAND2X0 U13961 ( .IN1(n3431), .IN2(n12389), .QN(n13260) );
  NAND2X0 U13962 ( .IN1(n3689), .IN2(g767), .QN(n3431) );
  NOR2X0 U13963 ( .IN1(n3689), .IN2(g767), .QN(n13922) );
  NAND2X0 U13964 ( .IN1(n13923), .IN2(n13924), .QN(g26827) );
  NAND2X0 U13965 ( .IN1(n13925), .IN2(n4606), .QN(n13924) );
  INVX0 U13966 ( .INP(n13926), .ZN(n13923) );
  NOR2X0 U13967 ( .IN1(n11841), .IN2(n8711), .QN(n13926) );
  NAND2X0 U13968 ( .IN1(n13927), .IN2(n13928), .QN(g26826) );
  NAND2X0 U13969 ( .IN1(n13925), .IN2(g7264), .QN(n13928) );
  INVX0 U13970 ( .INP(n13929), .ZN(n13927) );
  NOR2X0 U13971 ( .IN1(n10669), .IN2(n8700), .QN(n13929) );
  NAND2X0 U13972 ( .IN1(n13930), .IN2(n13931), .QN(g26825) );
  NAND2X0 U13973 ( .IN1(n4606), .IN2(n13932), .QN(n13931) );
  INVX0 U13974 ( .INP(n13933), .ZN(n13930) );
  NOR2X0 U13975 ( .IN1(n11841), .IN2(n8713), .QN(n13933) );
  NAND2X0 U13976 ( .IN1(n13934), .IN2(n13935), .QN(g26824) );
  NAND2X0 U13977 ( .IN1(n13936), .IN2(n4618), .QN(n13935) );
  NAND2X0 U13978 ( .IN1(test_so59), .IN2(n4511), .QN(n13934) );
  NAND2X0 U13979 ( .IN1(n13937), .IN2(n13938), .QN(g26823) );
  NAND2X0 U13980 ( .IN1(n13925), .IN2(g5555), .QN(n13938) );
  XNOR2X1 U13981 ( .IN1(n13939), .IN2(n13166), .Q(n13925) );
  NAND2X0 U13982 ( .IN1(n13940), .IN2(test_so79), .QN(n13939) );
  NOR2X0 U13983 ( .IN1(n13941), .IN2(n13159), .QN(n13940) );
  INVX0 U13984 ( .INP(n13942), .ZN(n13159) );
  NAND2X0 U13985 ( .IN1(n13943), .IN2(n13944), .QN(n13942) );
  NAND2X0 U13986 ( .IN1(n13945), .IN2(n13167), .QN(n13944) );
  NOR2X0 U13987 ( .IN1(n13169), .IN2(n13168), .QN(n13945) );
  INVX0 U13988 ( .INP(n13166), .ZN(n13169) );
  NAND2X0 U13989 ( .IN1(n13946), .IN2(n13171), .QN(n13943) );
  NOR2X0 U13990 ( .IN1(n13172), .IN2(n13166), .QN(n13946) );
  INVX0 U13991 ( .INP(n13168), .ZN(n13172) );
  NOR2X0 U13992 ( .IN1(n13158), .IN2(n13160), .QN(n13941) );
  NAND2X0 U13993 ( .IN1(n13947), .IN2(n13948), .QN(n13160) );
  NAND2X0 U13994 ( .IN1(n8946), .IN2(n11931), .QN(n13948) );
  NAND2X0 U13995 ( .IN1(n8937), .IN2(n10669), .QN(n13947) );
  NOR2X0 U13996 ( .IN1(n4509), .IN2(test_so81), .QN(n13158) );
  NAND2X0 U13997 ( .IN1(n4516), .IN2(g2513), .QN(n13937) );
  NAND2X0 U13998 ( .IN1(n13949), .IN2(n13950), .QN(g26822) );
  NAND2X0 U13999 ( .IN1(g7264), .IN2(n13932), .QN(n13950) );
  INVX0 U14000 ( .INP(n13951), .ZN(n13949) );
  NOR2X0 U14001 ( .IN1(n10669), .IN2(n8701), .QN(n13951) );
  NAND2X0 U14002 ( .IN1(n13952), .IN2(n13953), .QN(g26821) );
  NAND2X0 U14003 ( .IN1(n13936), .IN2(g7014), .QN(n13953) );
  INVX0 U14004 ( .INP(n13954), .ZN(n13952) );
  NOR2X0 U14005 ( .IN1(n10678), .IN2(n8704), .QN(n13954) );
  NAND2X0 U14006 ( .IN1(n13955), .IN2(n13956), .QN(g26820) );
  NAND2X0 U14007 ( .IN1(n4618), .IN2(n13957), .QN(n13956) );
  INVX0 U14008 ( .INP(n13958), .ZN(n13955) );
  NOR2X0 U14009 ( .IN1(n11849), .IN2(n8719), .QN(n13958) );
  NAND2X0 U14010 ( .IN1(n13959), .IN2(n13960), .QN(g26818) );
  NAND2X0 U14011 ( .IN1(n4381), .IN2(g1131), .QN(n13960) );
  NAND2X0 U14012 ( .IN1(n13961), .IN2(g1088), .QN(n13959) );
  NAND2X0 U14013 ( .IN1(n13962), .IN2(n13963), .QN(g26817) );
  NAND2X0 U14014 ( .IN1(g5555), .IN2(n13932), .QN(n13963) );
  NAND2X0 U14015 ( .IN1(n13964), .IN2(n13965), .QN(n13932) );
  NAND2X0 U14016 ( .IN1(n13171), .IN2(test_so79), .QN(n13965) );
  INVX0 U14017 ( .INP(n13167), .ZN(n13171) );
  NAND2X0 U14018 ( .IN1(n12449), .IN2(n13966), .QN(n13167) );
  NAND2X0 U14019 ( .IN1(n13967), .IN2(n13968), .QN(n13966) );
  NAND2X0 U14020 ( .IN1(n8850), .IN2(test_so73), .QN(n13968) );
  NOR2X0 U14021 ( .IN1(n13969), .IN2(n13970), .QN(n13967) );
  NOR2X0 U14022 ( .IN1(n4367), .IN2(g2253), .QN(n13970) );
  NOR2X0 U14023 ( .IN1(n4324), .IN2(g2254), .QN(n13969) );
  INVX0 U14024 ( .INP(n13971), .ZN(n12449) );
  NAND2X0 U14025 ( .IN1(n13168), .IN2(n9281), .QN(n13964) );
  NAND2X0 U14026 ( .IN1(n13972), .IN2(n13973), .QN(n13168) );
  NAND2X0 U14027 ( .IN1(g5555), .IN2(g2504), .QN(n13973) );
  NOR2X0 U14028 ( .IN1(n13974), .IN2(n13975), .QN(n13972) );
  NOR2X0 U14029 ( .IN1(n8701), .IN2(n12443), .QN(n13975) );
  NOR2X0 U14030 ( .IN1(n8713), .IN2(n13976), .QN(n13974) );
  NAND2X0 U14031 ( .IN1(n4516), .IN2(g2504), .QN(n13962) );
  NAND2X0 U14032 ( .IN1(n13977), .IN2(n13978), .QN(g26816) );
  NAND2X0 U14033 ( .IN1(n13936), .IN2(g5511), .QN(n13978) );
  XNOR2X1 U14034 ( .IN1(n13979), .IN2(n13980), .Q(n13936) );
  NAND2X0 U14035 ( .IN1(n13187), .IN2(n13981), .QN(n13979) );
  NAND2X0 U14036 ( .IN1(n13982), .IN2(n13186), .QN(n13981) );
  NAND2X0 U14037 ( .IN1(n8940), .IN2(n10678), .QN(n13186) );
  INVX0 U14038 ( .INP(n13185), .ZN(n13982) );
  NAND2X0 U14039 ( .IN1(n13983), .IN2(n13984), .QN(n13185) );
  NAND2X0 U14040 ( .IN1(n8950), .IN2(n11849), .QN(n13984) );
  NAND2X0 U14041 ( .IN1(n8951), .IN2(n12050), .QN(n13983) );
  NAND2X0 U14042 ( .IN1(n13985), .IN2(n13986), .QN(n13187) );
  NAND2X0 U14043 ( .IN1(n13192), .IN2(n13191), .QN(n13986) );
  NOR2X0 U14044 ( .IN1(n13987), .IN2(n13988), .QN(n13192) );
  NAND2X0 U14045 ( .IN1(g1690), .IN2(n13989), .QN(n13987) );
  NAND2X0 U14046 ( .IN1(n13190), .IN2(n13193), .QN(n13985) );
  INVX0 U14047 ( .INP(n13191), .ZN(n13193) );
  NOR2X0 U14048 ( .IN1(n13989), .IN2(n13990), .QN(n13190) );
  NAND2X0 U14049 ( .IN1(n13988), .IN2(g1690), .QN(n13990) );
  INVX0 U14050 ( .INP(n13980), .ZN(n13989) );
  NAND2X0 U14051 ( .IN1(n4518), .IN2(g1819), .QN(n13977) );
  NAND2X0 U14052 ( .IN1(n13991), .IN2(n13992), .QN(g26815) );
  NAND2X0 U14053 ( .IN1(g7014), .IN2(n13957), .QN(n13992) );
  INVX0 U14054 ( .INP(n13993), .ZN(n13991) );
  NOR2X0 U14055 ( .IN1(n10678), .IN2(n8705), .QN(n13993) );
  NAND2X0 U14056 ( .IN1(n13994), .IN2(n13995), .QN(g26814) );
  INVX0 U14057 ( .INP(n13996), .ZN(n13995) );
  NOR2X0 U14058 ( .IN1(g6712), .IN2(n8708), .QN(n13996) );
  NAND2X0 U14059 ( .IN1(n13961), .IN2(g6712), .QN(n13994) );
  NAND2X0 U14060 ( .IN1(n13997), .IN2(n13998), .QN(g26813) );
  NAND2X0 U14061 ( .IN1(n4381), .IN2(g1122), .QN(n13998) );
  NAND2X0 U14062 ( .IN1(n13999), .IN2(g1088), .QN(n13997) );
  NAND2X0 U14063 ( .IN1(n14000), .IN2(n14001), .QN(g26812) );
  NAND2X0 U14064 ( .IN1(n14002), .IN2(n4640), .QN(n14001) );
  INVX0 U14065 ( .INP(n14003), .ZN(n14000) );
  NOR2X0 U14066 ( .IN1(n11886), .IN2(n8733), .QN(n14003) );
  NAND2X0 U14067 ( .IN1(n14004), .IN2(n14005), .QN(g26811) );
  NAND2X0 U14068 ( .IN1(g5511), .IN2(n13957), .QN(n14005) );
  NAND2X0 U14069 ( .IN1(n14006), .IN2(n14007), .QN(n13957) );
  INVX0 U14070 ( .INP(n14008), .ZN(n14007) );
  NOR2X0 U14071 ( .IN1(n13988), .IN2(n4386), .QN(n14008) );
  NAND2X0 U14072 ( .IN1(n12494), .IN2(n14009), .QN(n13988) );
  NAND2X0 U14073 ( .IN1(n14010), .IN2(n14011), .QN(n14009) );
  NAND2X0 U14074 ( .IN1(n8862), .IN2(g6782), .QN(n14011) );
  NOR2X0 U14075 ( .IN1(n14012), .IN2(n14013), .QN(n14010) );
  NOR2X0 U14076 ( .IN1(n4368), .IN2(g1559), .QN(n14013) );
  NOR2X0 U14077 ( .IN1(n4317), .IN2(g1560), .QN(n14012) );
  INVX0 U14078 ( .INP(n14014), .ZN(n12494) );
  NAND2X0 U14079 ( .IN1(n4386), .IN2(n13191), .QN(n14006) );
  NAND2X0 U14080 ( .IN1(n14015), .IN2(n14016), .QN(n13191) );
  NAND2X0 U14081 ( .IN1(g5511), .IN2(g1810), .QN(n14016) );
  NOR2X0 U14082 ( .IN1(n14017), .IN2(n14018), .QN(n14015) );
  NOR2X0 U14083 ( .IN1(n8705), .IN2(n11731), .QN(n14018) );
  NOR2X0 U14084 ( .IN1(n8719), .IN2(n12488), .QN(n14017) );
  NAND2X0 U14085 ( .IN1(n4518), .IN2(g1810), .QN(n14004) );
  NAND2X0 U14086 ( .IN1(n14019), .IN2(n14020), .QN(g26810) );
  INVX0 U14087 ( .INP(n14021), .ZN(n14020) );
  NOR2X0 U14088 ( .IN1(g5472), .IN2(n8726), .QN(n14021) );
  NAND2X0 U14089 ( .IN1(n13961), .IN2(g5472), .QN(n14019) );
  XNOR2X1 U14090 ( .IN1(n14022), .IN2(n14023), .Q(n13961) );
  NAND2X0 U14091 ( .IN1(n13208), .IN2(n14024), .QN(n14022) );
  NAND2X0 U14092 ( .IN1(n14025), .IN2(n13207), .QN(n14024) );
  NAND2X0 U14093 ( .IN1(n8943), .IN2(g6712), .QN(n13207) );
  INVX0 U14094 ( .INP(n13206), .ZN(n14025) );
  NAND2X0 U14095 ( .IN1(n14026), .IN2(n14027), .QN(n13206) );
  NAND2X0 U14096 ( .IN1(n8957), .IN2(g5472), .QN(n14027) );
  NAND2X0 U14097 ( .IN1(n8956), .IN2(g1088), .QN(n14026) );
  NAND2X0 U14098 ( .IN1(n14028), .IN2(n14029), .QN(n13208) );
  NAND2X0 U14099 ( .IN1(n13213), .IN2(n13212), .QN(n14029) );
  NOR2X0 U14100 ( .IN1(n14030), .IN2(n14031), .QN(n13213) );
  NAND2X0 U14101 ( .IN1(g996), .IN2(n14032), .QN(n14030) );
  NAND2X0 U14102 ( .IN1(n13211), .IN2(n13214), .QN(n14028) );
  INVX0 U14103 ( .INP(n13212), .ZN(n13214) );
  NOR2X0 U14104 ( .IN1(n14032), .IN2(n14033), .QN(n13211) );
  NAND2X0 U14105 ( .IN1(n14031), .IN2(g996), .QN(n14033) );
  INVX0 U14106 ( .INP(n14023), .ZN(n14032) );
  NAND2X0 U14107 ( .IN1(n14034), .IN2(n14035), .QN(g26809) );
  NAND2X0 U14108 ( .IN1(n13999), .IN2(g6712), .QN(n14035) );
  NAND2X0 U14109 ( .IN1(n4364), .IN2(test_so38), .QN(n14034) );
  NAND2X0 U14110 ( .IN1(n14036), .IN2(n14037), .QN(g26808) );
  NAND2X0 U14111 ( .IN1(n14002), .IN2(g6447), .QN(n14037) );
  INVX0 U14112 ( .INP(n14038), .ZN(n14036) );
  NOR2X0 U14113 ( .IN1(n11905), .IN2(n8734), .QN(n14038) );
  NAND2X0 U14114 ( .IN1(n14039), .IN2(n14040), .QN(g26807) );
  NAND2X0 U14115 ( .IN1(n4640), .IN2(n14041), .QN(n14040) );
  INVX0 U14116 ( .INP(n14042), .ZN(n14039) );
  NOR2X0 U14117 ( .IN1(n11886), .IN2(n8736), .QN(n14042) );
  NAND2X0 U14118 ( .IN1(n14043), .IN2(n14044), .QN(g26806) );
  INVX0 U14119 ( .INP(n14045), .ZN(n14044) );
  NOR2X0 U14120 ( .IN1(g5472), .IN2(n8728), .QN(n14045) );
  NAND2X0 U14121 ( .IN1(n13999), .IN2(g5472), .QN(n14043) );
  NAND2X0 U14122 ( .IN1(n14046), .IN2(n14047), .QN(n13999) );
  INVX0 U14123 ( .INP(n14048), .ZN(n14047) );
  NOR2X0 U14124 ( .IN1(n14031), .IN2(n4387), .QN(n14048) );
  NAND2X0 U14125 ( .IN1(n12534), .IN2(n14049), .QN(n14031) );
  NAND2X0 U14126 ( .IN1(n14050), .IN2(n14051), .QN(n14049) );
  NAND2X0 U14127 ( .IN1(n8872), .IN2(test_so31), .QN(n14051) );
  NOR2X0 U14128 ( .IN1(n14052), .IN2(n14053), .QN(n14050) );
  NOR2X0 U14129 ( .IN1(n4323), .IN2(g866), .QN(n14053) );
  NOR2X0 U14130 ( .IN1(n4312), .IN2(g867), .QN(n14052) );
  INVX0 U14131 ( .INP(n14054), .ZN(n12534) );
  NAND2X0 U14132 ( .IN1(n4387), .IN2(n13212), .QN(n14046) );
  NAND2X0 U14133 ( .IN1(n14055), .IN2(n14056), .QN(n13212) );
  NAND2X0 U14134 ( .IN1(g1088), .IN2(g1122), .QN(n14056) );
  NOR2X0 U14135 ( .IN1(n14057), .IN2(n14058), .QN(n14055) );
  INVX0 U14136 ( .INP(n14059), .ZN(n14058) );
  NAND2X0 U14137 ( .IN1(g6712), .IN2(test_so38), .QN(n14059) );
  NOR2X0 U14138 ( .IN1(n8728), .IN2(n4363), .QN(n14057) );
  NAND2X0 U14139 ( .IN1(n14060), .IN2(n14061), .QN(g26805) );
  NAND2X0 U14140 ( .IN1(n14002), .IN2(g5437), .QN(n14061) );
  XNOR2X1 U14141 ( .IN1(n14062), .IN2(n14063), .Q(n14002) );
  NAND2X0 U14142 ( .IN1(n13224), .IN2(n14064), .QN(n14062) );
  NAND2X0 U14143 ( .IN1(n14065), .IN2(n13223), .QN(n14064) );
  NAND2X0 U14144 ( .IN1(n8963), .IN2(n11886), .QN(n13223) );
  INVX0 U14145 ( .INP(n13222), .ZN(n14065) );
  NAND2X0 U14146 ( .IN1(n14066), .IN2(n14067), .QN(n13222) );
  NAND2X0 U14147 ( .IN1(n8964), .IN2(n11905), .QN(n14067) );
  NAND2X0 U14148 ( .IN1(n8965), .IN2(n10752), .QN(n14066) );
  NAND2X0 U14149 ( .IN1(n14068), .IN2(n14069), .QN(n13224) );
  NAND2X0 U14150 ( .IN1(n13229), .IN2(n13228), .QN(n14069) );
  NOR2X0 U14151 ( .IN1(n14070), .IN2(n14071), .QN(n13229) );
  NAND2X0 U14152 ( .IN1(g309), .IN2(n14072), .QN(n14070) );
  NAND2X0 U14153 ( .IN1(n13227), .IN2(n13230), .QN(n14068) );
  INVX0 U14154 ( .INP(n13228), .ZN(n13230) );
  NOR2X0 U14155 ( .IN1(n14072), .IN2(n14073), .QN(n13227) );
  NAND2X0 U14156 ( .IN1(n14071), .IN2(g309), .QN(n14073) );
  INVX0 U14157 ( .INP(n14063), .ZN(n14072) );
  NAND2X0 U14158 ( .IN1(n4520), .IN2(g438), .QN(n14060) );
  NAND2X0 U14159 ( .IN1(n14074), .IN2(n14075), .QN(g26804) );
  NAND2X0 U14160 ( .IN1(g6447), .IN2(n14041), .QN(n14075) );
  INVX0 U14161 ( .INP(n14076), .ZN(n14074) );
  NOR2X0 U14162 ( .IN1(n11905), .IN2(n8737), .QN(n14076) );
  NAND2X0 U14163 ( .IN1(n14077), .IN2(n14078), .QN(g26803) );
  NAND2X0 U14164 ( .IN1(g5437), .IN2(n14041), .QN(n14078) );
  NAND2X0 U14165 ( .IN1(n14079), .IN2(n14080), .QN(n14041) );
  INVX0 U14166 ( .INP(n14081), .ZN(n14080) );
  NOR2X0 U14167 ( .IN1(n14071), .IN2(n4388), .QN(n14081) );
  NAND2X0 U14168 ( .IN1(n12569), .IN2(n14082), .QN(n14071) );
  NAND2X0 U14169 ( .IN1(n14083), .IN2(n14084), .QN(n14082) );
  NAND2X0 U14170 ( .IN1(n8884), .IN2(g6313), .QN(n14084) );
  NOR2X0 U14171 ( .IN1(n14085), .IN2(n14086), .QN(n14083) );
  NOR2X0 U14172 ( .IN1(n4369), .IN2(g177), .QN(n14086) );
  NOR2X0 U14173 ( .IN1(n4318), .IN2(g178), .QN(n14085) );
  NAND2X0 U14174 ( .IN1(n4388), .IN2(n13228), .QN(n14079) );
  NAND2X0 U14175 ( .IN1(n14087), .IN2(n14088), .QN(n13228) );
  NAND2X0 U14176 ( .IN1(g5437), .IN2(g429), .QN(n14088) );
  NOR2X0 U14177 ( .IN1(n14089), .IN2(n14090), .QN(n14087) );
  NOR2X0 U14178 ( .IN1(n8737), .IN2(n12562), .QN(n14090) );
  NOR2X0 U14179 ( .IN1(n8736), .IN2(n12563), .QN(n14089) );
  NAND2X0 U14180 ( .IN1(n4520), .IN2(g429), .QN(n14077) );
  NOR2X0 U14181 ( .IN1(n9867), .IN2(n14091), .QN(g26798) );
  XNOR2X1 U14182 ( .IN1(n4355), .IN2(n14092), .Q(n14091) );
  NAND2X0 U14183 ( .IN1(n9679), .IN2(g2900), .QN(n14092) );
  NOR2X0 U14184 ( .IN1(n10617), .IN2(n14093), .QN(g26795) );
  XNOR2X1 U14185 ( .IN1(n13920), .IN2(n9282), .Q(n14093) );
  NOR2X0 U14186 ( .IN1(n14094), .IN2(n14095), .QN(g26789) );
  XOR2X1 U14187 ( .IN1(n4468), .IN2(n13240), .Q(n14095) );
  INVX0 U14188 ( .INP(n13242), .ZN(n13240) );
  NOR2X0 U14189 ( .IN1(n14096), .IN2(n14097), .QN(g26786) );
  XNOR2X1 U14190 ( .IN1(n8387), .IN2(n3741), .Q(n14096) );
  NOR2X0 U14191 ( .IN1(n14098), .IN2(n14099), .QN(g26781) );
  XNOR2X1 U14192 ( .IN1(n4469), .IN2(n13248), .Q(n14099) );
  NOR2X0 U14193 ( .IN1(n9684), .IN2(n14100), .QN(g26776) );
  XNOR2X1 U14194 ( .IN1(n13253), .IN2(n9283), .Q(n14100) );
  NOR2X0 U14195 ( .IN1(n14101), .IN2(n14102), .QN(g26677) );
  NAND2X0 U14196 ( .IN1(n13920), .IN2(n13918), .QN(n14102) );
  NAND2X0 U14197 ( .IN1(n14103), .IN2(n14104), .QN(n13920) );
  NOR2X0 U14198 ( .IN1(n4407), .IN2(n4397), .QN(n14103) );
  NOR2X0 U14199 ( .IN1(n14105), .IN2(g2746), .QN(n14101) );
  NOR2X0 U14200 ( .IN1(n4397), .IN2(n14106), .QN(n14105) );
  NAND2X0 U14201 ( .IN1(n14107), .IN2(n14108), .QN(g26676) );
  NAND2X0 U14202 ( .IN1(n14109), .IN2(g2479), .QN(n14108) );
  NAND2X0 U14203 ( .IN1(n14110), .IN2(n10669), .QN(n14109) );
  NAND2X0 U14204 ( .IN1(n14111), .IN2(n10669), .QN(n14107) );
  NAND2X0 U14205 ( .IN1(n14112), .IN2(n14113), .QN(g26675) );
  NAND2X0 U14206 ( .IN1(n14114), .IN2(g1783), .QN(n14113) );
  NAND2X0 U14207 ( .IN1(n10448), .IN2(n11849), .QN(n14114) );
  NAND2X0 U14208 ( .IN1(n14115), .IN2(n11849), .QN(n14112) );
  INVX0 U14209 ( .INP(n4511), .ZN(n11849) );
  NAND2X0 U14210 ( .IN1(n14116), .IN2(n14117), .QN(g26672) );
  NAND2X0 U14211 ( .IN1(n14118), .IN2(g2478), .QN(n14117) );
  NAND2X0 U14212 ( .IN1(n14110), .IN2(n11931), .QN(n14118) );
  NAND2X0 U14213 ( .IN1(n14111), .IN2(n11931), .QN(n14116) );
  INVX0 U14214 ( .INP(n4516), .ZN(n11931) );
  NOR2X0 U14215 ( .IN1(n14119), .IN2(n14120), .QN(g26671) );
  NAND2X0 U14216 ( .IN1(n13242), .IN2(n13126), .QN(n14120) );
  NAND2X0 U14217 ( .IN1(n14121), .IN2(n14122), .QN(n13242) );
  INVX0 U14218 ( .INP(n14123), .ZN(n14122) );
  NOR2X0 U14219 ( .IN1(n4409), .IN2(n4399), .QN(n14121) );
  NOR2X0 U14220 ( .IN1(n14124), .IN2(g2052), .QN(n14119) );
  NOR2X0 U14221 ( .IN1(n4399), .IN2(n14123), .QN(n14124) );
  NAND2X0 U14222 ( .IN1(n14125), .IN2(n14126), .QN(g26670) );
  NAND2X0 U14223 ( .IN1(n14127), .IN2(g1785), .QN(n14126) );
  NAND2X0 U14224 ( .IN1(n10448), .IN2(n10678), .QN(n14127) );
  NAND2X0 U14225 ( .IN1(n14115), .IN2(n10678), .QN(n14125) );
  NAND2X0 U14226 ( .IN1(n14128), .IN2(n14129), .QN(g26669) );
  NAND2X0 U14227 ( .IN1(n14130), .IN2(g1089), .QN(n14129) );
  NAND2X0 U14228 ( .IN1(n10447), .IN2(g1088), .QN(n14130) );
  NAND2X0 U14229 ( .IN1(n14131), .IN2(g1088), .QN(n14128) );
  NAND2X0 U14230 ( .IN1(n14132), .IN2(n14133), .QN(g26667) );
  NAND2X0 U14231 ( .IN1(test_so60), .IN2(n14134), .QN(n14133) );
  NAND2X0 U14232 ( .IN1(n10448), .IN2(n12050), .QN(n14134) );
  NAND2X0 U14233 ( .IN1(n14115), .IN2(n12050), .QN(n14132) );
  INVX0 U14234 ( .INP(n4518), .ZN(n12050) );
  NOR2X0 U14235 ( .IN1(n10448), .IN2(n4386), .QN(n14115) );
  NOR2X0 U14236 ( .IN1(n14135), .IN2(n11781), .QN(n10448) );
  NAND2X0 U14237 ( .IN1(n14136), .IN2(n14137), .QN(n11781) );
  NAND2X0 U14238 ( .IN1(n8939), .IN2(n10678), .QN(n14137) );
  NOR2X0 U14239 ( .IN1(n14138), .IN2(n14139), .QN(n14136) );
  NOR2X0 U14240 ( .IN1(test_so60), .IN2(n4518), .QN(n14139) );
  NOR2X0 U14241 ( .IN1(n4511), .IN2(g1783), .QN(n14138) );
  NAND2X0 U14242 ( .IN1(g1690), .IN2(n14140), .QN(n14135) );
  INVX0 U14243 ( .INP(n11543), .ZN(n14140) );
  NAND2X0 U14244 ( .IN1(n14141), .IN2(n14142), .QN(n11543) );
  NOR2X0 U14245 ( .IN1(n14143), .IN2(n14144), .QN(n14142) );
  NAND2X0 U14246 ( .IN1(n14145), .IN2(n14146), .QN(n14144) );
  XNOR2X1 U14247 ( .IN1(n10835), .IN2(n14147), .Q(n14146) );
  NOR2X0 U14248 ( .IN1(n14148), .IN2(n14149), .QN(n14147) );
  NAND2X0 U14249 ( .IN1(n14150), .IN2(n14151), .QN(n14149) );
  NAND2X0 U14250 ( .IN1(n8805), .IN2(g6573), .QN(n14151) );
  NAND2X0 U14251 ( .IN1(n8803), .IN2(g1547), .QN(n14150) );
  NOR2X0 U14252 ( .IN1(n4515), .IN2(g1546), .QN(n14148) );
  NOR2X0 U14253 ( .IN1(n14152), .IN2(n14153), .QN(n14145) );
  XNOR2X1 U14254 ( .IN1(n4378), .IN2(n14154), .Q(n14153) );
  NAND2X0 U14255 ( .IN1(n14155), .IN2(n14156), .QN(n14154) );
  NAND2X0 U14256 ( .IN1(n9183), .IN2(g6782), .QN(n14156) );
  NOR2X0 U14257 ( .IN1(n14157), .IN2(n14158), .QN(n14155) );
  NOR2X0 U14258 ( .IN1(n4368), .IN2(g1511), .QN(n14158) );
  NOR2X0 U14259 ( .IN1(n4317), .IN2(g1512), .QN(n14157) );
  XNOR2X1 U14260 ( .IN1(n4320), .IN2(n14159), .Q(n14152) );
  NAND2X0 U14261 ( .IN1(n14160), .IN2(n14161), .QN(n14159) );
  NAND2X0 U14262 ( .IN1(n9180), .IN2(g6782), .QN(n14161) );
  NOR2X0 U14263 ( .IN1(n14162), .IN2(n14163), .QN(n14160) );
  NOR2X0 U14264 ( .IN1(n4368), .IN2(g1523), .QN(n14163) );
  NOR2X0 U14265 ( .IN1(n4317), .IN2(g1524), .QN(n14162) );
  NAND2X0 U14266 ( .IN1(n14164), .IN2(n14165), .QN(n14143) );
  XNOR2X1 U14267 ( .IN1(n11025), .IN2(n14166), .Q(n14165) );
  NOR2X0 U14268 ( .IN1(n14167), .IN2(n14168), .QN(n14166) );
  NAND2X0 U14269 ( .IN1(n14169), .IN2(n14170), .QN(n14168) );
  NAND2X0 U14270 ( .IN1(n8789), .IN2(g6573), .QN(n14170) );
  NAND2X0 U14271 ( .IN1(n8787), .IN2(g1547), .QN(n14169) );
  NOR2X0 U14272 ( .IN1(n4515), .IN2(g1543), .QN(n14167) );
  NOR2X0 U14273 ( .IN1(n10702), .IN2(n14171), .QN(n14164) );
  XNOR2X1 U14274 ( .IN1(n4374), .IN2(n14172), .Q(n14171) );
  NAND2X0 U14275 ( .IN1(n14173), .IN2(n14174), .QN(n14172) );
  NAND2X0 U14276 ( .IN1(n9182), .IN2(g6782), .QN(n14174) );
  NOR2X0 U14277 ( .IN1(n14175), .IN2(n14176), .QN(n14173) );
  NOR2X0 U14278 ( .IN1(n4368), .IN2(g1514), .QN(n14176) );
  NOR2X0 U14279 ( .IN1(test_so52), .IN2(n4317), .QN(n14175) );
  INVX0 U14280 ( .INP(n3070), .ZN(n10702) );
  NOR2X0 U14281 ( .IN1(n14177), .IN2(n14178), .QN(n14141) );
  NAND2X0 U14282 ( .IN1(n14179), .IN2(n14180), .QN(n14178) );
  XNOR2X1 U14283 ( .IN1(n14181), .IN2(g1501), .Q(n14180) );
  NAND2X0 U14284 ( .IN1(n14182), .IN2(n14183), .QN(n14181) );
  INVX0 U14285 ( .INP(n14184), .ZN(n14183) );
  NOR2X0 U14286 ( .IN1(n4515), .IN2(test_so53), .QN(n14184) );
  NOR2X0 U14287 ( .IN1(n14185), .IN2(n14186), .QN(n14182) );
  NOR2X0 U14288 ( .IN1(n4368), .IN2(g1535), .QN(n14186) );
  NOR2X0 U14289 ( .IN1(n4317), .IN2(g1536), .QN(n14185) );
  XNOR2X1 U14290 ( .IN1(n14187), .IN2(g1486), .Q(n14179) );
  NAND2X0 U14291 ( .IN1(n14188), .IN2(n14189), .QN(n14187) );
  NAND2X0 U14292 ( .IN1(n9178), .IN2(g6782), .QN(n14189) );
  NOR2X0 U14293 ( .IN1(n14190), .IN2(n14191), .QN(n14188) );
  NOR2X0 U14294 ( .IN1(n4368), .IN2(g1526), .QN(n14191) );
  NOR2X0 U14295 ( .IN1(n4317), .IN2(g1527), .QN(n14190) );
  NAND2X0 U14296 ( .IN1(n14192), .IN2(n14193), .QN(n14177) );
  XNOR2X1 U14297 ( .IN1(n14194), .IN2(g1491), .Q(n14193) );
  NAND2X0 U14298 ( .IN1(n14195), .IN2(n14196), .QN(n14194) );
  NAND2X0 U14299 ( .IN1(n9176), .IN2(g6782), .QN(n14196) );
  NOR2X0 U14300 ( .IN1(n14197), .IN2(n14198), .QN(n14195) );
  NOR2X0 U14301 ( .IN1(n4368), .IN2(g1529), .QN(n14198) );
  NOR2X0 U14302 ( .IN1(n4317), .IN2(g1530), .QN(n14197) );
  NOR2X0 U14303 ( .IN1(n14199), .IN2(n14200), .QN(n14192) );
  XNOR2X1 U14304 ( .IN1(n4288), .IN2(n14201), .Q(n14200) );
  NAND2X0 U14305 ( .IN1(n14202), .IN2(n14203), .QN(n14201) );
  NAND2X0 U14306 ( .IN1(n9171), .IN2(g6782), .QN(n14203) );
  NOR2X0 U14307 ( .IN1(n14204), .IN2(n14205), .QN(n14202) );
  NOR2X0 U14308 ( .IN1(n4368), .IN2(g1538), .QN(n14205) );
  NOR2X0 U14309 ( .IN1(n4317), .IN2(g1539), .QN(n14204) );
  XNOR2X1 U14310 ( .IN1(n4557), .IN2(n14206), .Q(n14199) );
  NAND2X0 U14311 ( .IN1(n14207), .IN2(n14208), .QN(n14206) );
  NAND2X0 U14312 ( .IN1(n9174), .IN2(g6782), .QN(n14208) );
  NOR2X0 U14313 ( .IN1(n14209), .IN2(n14210), .QN(n14207) );
  NOR2X0 U14314 ( .IN1(n4368), .IN2(g1532), .QN(n14210) );
  NOR2X0 U14315 ( .IN1(n4317), .IN2(g1533), .QN(n14209) );
  NOR2X0 U14316 ( .IN1(n14211), .IN2(n14212), .QN(g26666) );
  NAND2X0 U14317 ( .IN1(n13248), .IN2(n13134), .QN(n14212) );
  INVX0 U14318 ( .INP(n13246), .ZN(n13248) );
  NOR2X0 U14319 ( .IN1(n14213), .IN2(n14214), .QN(n13246) );
  NAND2X0 U14320 ( .IN1(g1358), .IN2(g1346), .QN(n14213) );
  NOR2X0 U14321 ( .IN1(n14215), .IN2(g1358), .QN(n14211) );
  NOR2X0 U14322 ( .IN1(n4401), .IN2(n14214), .QN(n14215) );
  NAND2X0 U14323 ( .IN1(n14216), .IN2(n14217), .QN(g26665) );
  NAND2X0 U14324 ( .IN1(n14218), .IN2(g1091), .QN(n14217) );
  NAND2X0 U14325 ( .IN1(n10447), .IN2(g6712), .QN(n14218) );
  NAND2X0 U14326 ( .IN1(n14131), .IN2(g6712), .QN(n14216) );
  NAND2X0 U14327 ( .IN1(n14219), .IN2(n14220), .QN(g26664) );
  NAND2X0 U14328 ( .IN1(n14221), .IN2(g402), .QN(n14220) );
  NAND2X0 U14329 ( .IN1(n10446), .IN2(n11886), .QN(n14221) );
  NAND2X0 U14330 ( .IN1(n14222), .IN2(n11886), .QN(n14219) );
  INVX0 U14331 ( .INP(n4506), .ZN(n11886) );
  NAND2X0 U14332 ( .IN1(n14223), .IN2(n14224), .QN(g26661) );
  NAND2X0 U14333 ( .IN1(n14225), .IN2(g1090), .QN(n14224) );
  NAND2X0 U14334 ( .IN1(n10447), .IN2(g5472), .QN(n14225) );
  NAND2X0 U14335 ( .IN1(n14131), .IN2(g5472), .QN(n14223) );
  NOR2X0 U14336 ( .IN1(n10447), .IN2(n4387), .QN(n14131) );
  NOR2X0 U14337 ( .IN1(n14226), .IN2(n11795), .QN(n10447) );
  NAND2X0 U14338 ( .IN1(n14227), .IN2(n14228), .QN(n11795) );
  NAND2X0 U14339 ( .IN1(n8954), .IN2(g1088), .QN(n14228) );
  NOR2X0 U14340 ( .IN1(n14229), .IN2(n14230), .QN(n14227) );
  NOR2X0 U14341 ( .IN1(n4364), .IN2(g1091), .QN(n14230) );
  NOR2X0 U14342 ( .IN1(n4363), .IN2(g1090), .QN(n14229) );
  NAND2X0 U14343 ( .IN1(g996), .IN2(n11603), .QN(n14226) );
  INVX0 U14344 ( .INP(n14231), .ZN(n11603) );
  NAND2X0 U14345 ( .IN1(n14232), .IN2(n14233), .QN(n14231) );
  NOR2X0 U14346 ( .IN1(n14234), .IN2(n14235), .QN(n14233) );
  NAND2X0 U14347 ( .IN1(n14236), .IN2(n14237), .QN(n14235) );
  XOR2X1 U14348 ( .IN1(n14238), .IN2(n4379), .Q(n14237) );
  NAND2X0 U14349 ( .IN1(n14239), .IN2(n14240), .QN(n14238) );
  NAND2X0 U14350 ( .IN1(n8827), .IN2(test_so31), .QN(n14240) );
  NOR2X0 U14351 ( .IN1(n14241), .IN2(n14242), .QN(n14239) );
  NOR2X0 U14352 ( .IN1(n4323), .IN2(g818), .QN(n14242) );
  NOR2X0 U14353 ( .IN1(n4312), .IN2(g819), .QN(n14241) );
  NOR2X0 U14354 ( .IN1(n14243), .IN2(n14244), .QN(n14236) );
  XNOR2X1 U14355 ( .IN1(n4375), .IN2(n14245), .Q(n14244) );
  NAND2X0 U14356 ( .IN1(n14246), .IN2(n14247), .QN(n14245) );
  NAND2X0 U14357 ( .IN1(n8826), .IN2(test_so31), .QN(n14247) );
  NOR2X0 U14358 ( .IN1(n14248), .IN2(n14249), .QN(n14246) );
  NOR2X0 U14359 ( .IN1(n4323), .IN2(g821), .QN(n14249) );
  NOR2X0 U14360 ( .IN1(n4312), .IN2(g822), .QN(n14248) );
  XNOR2X1 U14361 ( .IN1(n4321), .IN2(n14250), .Q(n14243) );
  NAND2X0 U14362 ( .IN1(n14251), .IN2(n14252), .QN(n14250) );
  NAND2X0 U14363 ( .IN1(n8825), .IN2(test_so31), .QN(n14252) );
  NOR2X0 U14364 ( .IN1(n14253), .IN2(n14254), .QN(n14251) );
  NOR2X0 U14365 ( .IN1(n4323), .IN2(g830), .QN(n14254) );
  NOR2X0 U14366 ( .IN1(n4312), .IN2(g831), .QN(n14253) );
  NAND2X0 U14367 ( .IN1(n14255), .IN2(n14256), .QN(n14234) );
  XNOR2X1 U14368 ( .IN1(n10876), .IN2(n14257), .Q(n14256) );
  NOR2X0 U14369 ( .IN1(n14258), .IN2(n14259), .QN(n14257) );
  NAND2X0 U14370 ( .IN1(n14260), .IN2(n14261), .QN(n14259) );
  NAND2X0 U14371 ( .IN1(n8815), .IN2(g6518), .QN(n14261) );
  NAND2X0 U14372 ( .IN1(n8816), .IN2(g6368), .QN(n14260) );
  NOR2X0 U14373 ( .IN1(n9279), .IN2(g850), .QN(n14258) );
  NOR2X0 U14374 ( .IN1(n10519), .IN2(n14262), .QN(n14255) );
  XNOR2X1 U14375 ( .IN1(n11066), .IN2(n14263), .Q(n14262) );
  NAND2X0 U14376 ( .IN1(n14264), .IN2(n14265), .QN(n14263) );
  NAND2X0 U14377 ( .IN1(n8817), .IN2(test_so31), .QN(n14265) );
  NOR2X0 U14378 ( .IN1(n14266), .IN2(n14267), .QN(n14264) );
  NOR2X0 U14379 ( .IN1(n4323), .IN2(g848), .QN(n14267) );
  NOR2X0 U14380 ( .IN1(n4312), .IN2(g849), .QN(n14266) );
  INVX0 U14381 ( .INP(n3102), .ZN(n10519) );
  NOR2X0 U14382 ( .IN1(n14268), .IN2(n14269), .QN(n14232) );
  NAND2X0 U14383 ( .IN1(n14270), .IN2(n14271), .QN(n14269) );
  XNOR2X1 U14384 ( .IN1(n14272), .IN2(g809), .Q(n14271) );
  NAND2X0 U14385 ( .IN1(n14273), .IN2(n14274), .QN(n14272) );
  NAND2X0 U14386 ( .IN1(n8821), .IN2(test_so31), .QN(n14274) );
  NOR2X0 U14387 ( .IN1(n14275), .IN2(n14276), .QN(n14273) );
  NOR2X0 U14388 ( .IN1(n4323), .IN2(g842), .QN(n14276) );
  NOR2X0 U14389 ( .IN1(n4312), .IN2(g843), .QN(n14275) );
  XOR2X1 U14390 ( .IN1(n14277), .IN2(n4391), .Q(n14270) );
  NAND2X0 U14391 ( .IN1(n14278), .IN2(n14279), .QN(n14277) );
  NAND2X0 U14392 ( .IN1(n8824), .IN2(test_so31), .QN(n14279) );
  NOR2X0 U14393 ( .IN1(n14280), .IN2(n14281), .QN(n14278) );
  NOR2X0 U14394 ( .IN1(n4323), .IN2(g833), .QN(n14281) );
  NOR2X0 U14395 ( .IN1(n4312), .IN2(g834), .QN(n14280) );
  NAND2X0 U14396 ( .IN1(n14282), .IN2(n14283), .QN(n14268) );
  XNOR2X1 U14397 ( .IN1(n14284), .IN2(g801), .Q(n14283) );
  NAND2X0 U14398 ( .IN1(n14285), .IN2(n14286), .QN(n14284) );
  NAND2X0 U14399 ( .IN1(n8823), .IN2(test_so31), .QN(n14286) );
  NOR2X0 U14400 ( .IN1(n14287), .IN2(n14288), .QN(n14285) );
  NOR2X0 U14401 ( .IN1(n4323), .IN2(g836), .QN(n14288) );
  NOR2X0 U14402 ( .IN1(n4312), .IN2(g837), .QN(n14287) );
  NOR2X0 U14403 ( .IN1(n14289), .IN2(n14290), .QN(n14282) );
  XNOR2X1 U14404 ( .IN1(n4289), .IN2(n14291), .Q(n14290) );
  NAND2X0 U14405 ( .IN1(n14292), .IN2(n14293), .QN(n14291) );
  NAND2X0 U14406 ( .IN1(n8820), .IN2(test_so31), .QN(n14293) );
  NOR2X0 U14407 ( .IN1(n14294), .IN2(n14295), .QN(n14292) );
  NOR2X0 U14408 ( .IN1(n4323), .IN2(g845), .QN(n14295) );
  NOR2X0 U14409 ( .IN1(n4312), .IN2(g846), .QN(n14294) );
  XNOR2X1 U14410 ( .IN1(n4559), .IN2(n14296), .Q(n14289) );
  NAND2X0 U14411 ( .IN1(n14297), .IN2(n14298), .QN(n14296) );
  NAND2X0 U14412 ( .IN1(n8822), .IN2(test_so31), .QN(n14298) );
  NOR2X0 U14413 ( .IN1(n14299), .IN2(n14300), .QN(n14297) );
  NOR2X0 U14414 ( .IN1(test_so32), .IN2(n4323), .QN(n14300) );
  NOR2X0 U14415 ( .IN1(n4312), .IN2(g840), .QN(n14299) );
  NOR2X0 U14416 ( .IN1(n14301), .IN2(n14302), .QN(g26660) );
  NAND2X0 U14417 ( .IN1(n13253), .IN2(n13251), .QN(n14302) );
  NAND2X0 U14418 ( .IN1(n14303), .IN2(n14304), .QN(n13253) );
  NOR2X0 U14419 ( .IN1(n4413), .IN2(n4403), .QN(n14303) );
  NOR2X0 U14420 ( .IN1(n14305), .IN2(g672), .QN(n14301) );
  NOR2X0 U14421 ( .IN1(n4403), .IN2(n14306), .QN(n14305) );
  NAND2X0 U14422 ( .IN1(n14307), .IN2(n14308), .QN(g26659) );
  NAND2X0 U14423 ( .IN1(n14309), .IN2(g404), .QN(n14308) );
  NAND2X0 U14424 ( .IN1(n10446), .IN2(n11905), .QN(n14309) );
  NAND2X0 U14425 ( .IN1(n14222), .IN2(n11905), .QN(n14307) );
  INVX0 U14426 ( .INP(n4499), .ZN(n11905) );
  NAND2X0 U14427 ( .IN1(n14310), .IN2(n14311), .QN(g26655) );
  NAND2X0 U14428 ( .IN1(n14312), .IN2(g403), .QN(n14311) );
  NAND2X0 U14429 ( .IN1(n10446), .IN2(n10752), .QN(n14312) );
  NAND2X0 U14430 ( .IN1(n14222), .IN2(n10752), .QN(n14310) );
  NOR2X0 U14431 ( .IN1(n10446), .IN2(n4388), .QN(n14222) );
  NOR2X0 U14432 ( .IN1(n14313), .IN2(n11806), .QN(n10446) );
  NAND2X0 U14433 ( .IN1(n14314), .IN2(n14315), .QN(n11806) );
  NAND2X0 U14434 ( .IN1(n8962), .IN2(n10752), .QN(n14315) );
  NOR2X0 U14435 ( .IN1(n14316), .IN2(n14317), .QN(n14314) );
  NOR2X0 U14436 ( .IN1(n4506), .IN2(g402), .QN(n14317) );
  NOR2X0 U14437 ( .IN1(n4499), .IN2(g404), .QN(n14316) );
  NAND2X0 U14438 ( .IN1(g309), .IN2(n14318), .QN(n14313) );
  INVX0 U14439 ( .INP(n11671), .ZN(n14318) );
  NAND2X0 U14440 ( .IN1(n14319), .IN2(n14320), .QN(n11671) );
  NOR2X0 U14441 ( .IN1(n14321), .IN2(n14322), .QN(n14320) );
  NAND2X0 U14442 ( .IN1(n14323), .IN2(n14324), .QN(n14322) );
  XNOR2X1 U14443 ( .IN1(n10928), .IN2(n14325), .Q(n14324) );
  NOR2X0 U14444 ( .IN1(n14326), .IN2(n14327), .QN(n14325) );
  NAND2X0 U14445 ( .IN1(n14328), .IN2(n14329), .QN(n14327) );
  INVX0 U14446 ( .INP(n14330), .ZN(n14329) );
  NOR2X0 U14447 ( .IN1(n4318), .IN2(test_so12), .QN(n14330) );
  NAND2X0 U14448 ( .IN1(n8828), .IN2(g165), .QN(n14328) );
  NOR2X0 U14449 ( .IN1(n4512), .IN2(g164), .QN(n14326) );
  NOR2X0 U14450 ( .IN1(n14331), .IN2(n14332), .QN(n14323) );
  XNOR2X1 U14451 ( .IN1(n4380), .IN2(n14333), .Q(n14332) );
  NAND2X0 U14452 ( .IN1(n14334), .IN2(n14335), .QN(n14333) );
  NAND2X0 U14453 ( .IN1(n9214), .IN2(g6313), .QN(n14335) );
  NOR2X0 U14454 ( .IN1(n14336), .IN2(n14337), .QN(n14334) );
  NOR2X0 U14455 ( .IN1(n4369), .IN2(g129), .QN(n14337) );
  NOR2X0 U14456 ( .IN1(n4318), .IN2(g130), .QN(n14336) );
  XNOR2X1 U14457 ( .IN1(n4322), .IN2(n14338), .Q(n14331) );
  NAND2X0 U14458 ( .IN1(n14339), .IN2(n14340), .QN(n14338) );
  NAND2X0 U14459 ( .IN1(n9210), .IN2(g6313), .QN(n14340) );
  NOR2X0 U14460 ( .IN1(n14341), .IN2(n14342), .QN(n14339) );
  NOR2X0 U14461 ( .IN1(n4369), .IN2(g141), .QN(n14342) );
  NOR2X0 U14462 ( .IN1(n4318), .IN2(g142), .QN(n14341) );
  NAND2X0 U14463 ( .IN1(n14343), .IN2(n14344), .QN(n14321) );
  XNOR2X1 U14464 ( .IN1(n11093), .IN2(n14345), .Q(n14344) );
  NOR2X0 U14465 ( .IN1(n14346), .IN2(n14347), .QN(n14345) );
  NAND2X0 U14466 ( .IN1(n14348), .IN2(n14349), .QN(n14347) );
  NAND2X0 U14467 ( .IN1(n8792), .IN2(g6231), .QN(n14349) );
  NAND2X0 U14468 ( .IN1(n8790), .IN2(g165), .QN(n14348) );
  NOR2X0 U14469 ( .IN1(n4512), .IN2(g161), .QN(n14346) );
  NOR2X0 U14470 ( .IN1(n10741), .IN2(n14350), .QN(n14343) );
  XNOR2X1 U14471 ( .IN1(n4376), .IN2(n14351), .Q(n14350) );
  NAND2X0 U14472 ( .IN1(n14352), .IN2(n14353), .QN(n14351) );
  NAND2X0 U14473 ( .IN1(n9212), .IN2(g6313), .QN(n14353) );
  NOR2X0 U14474 ( .IN1(n14354), .IN2(n14355), .QN(n14352) );
  NOR2X0 U14475 ( .IN1(n4369), .IN2(g132), .QN(n14355) );
  NOR2X0 U14476 ( .IN1(n4318), .IN2(g133), .QN(n14354) );
  INVX0 U14477 ( .INP(n3130), .ZN(n10741) );
  NOR2X0 U14478 ( .IN1(n14356), .IN2(n14357), .QN(n14319) );
  NAND2X0 U14479 ( .IN1(n14358), .IN2(n14359), .QN(n14357) );
  XNOR2X1 U14480 ( .IN1(n14360), .IN2(g121), .Q(n14359) );
  NAND2X0 U14481 ( .IN1(n14361), .IN2(n14362), .QN(n14360) );
  NAND2X0 U14482 ( .IN1(n9202), .IN2(g6313), .QN(n14362) );
  NOR2X0 U14483 ( .IN1(n14363), .IN2(n14364), .QN(n14361) );
  NOR2X0 U14484 ( .IN1(n4369), .IN2(g153), .QN(n14364) );
  NOR2X0 U14485 ( .IN1(n4318), .IN2(g154), .QN(n14363) );
  XNOR2X1 U14486 ( .IN1(n14365), .IN2(g109), .Q(n14358) );
  NAND2X0 U14487 ( .IN1(n14366), .IN2(n14367), .QN(n14365) );
  NAND2X0 U14488 ( .IN1(n9208), .IN2(g6313), .QN(n14367) );
  NOR2X0 U14489 ( .IN1(n14368), .IN2(n14369), .QN(n14366) );
  NOR2X0 U14490 ( .IN1(test_so11), .IN2(n4369), .QN(n14369) );
  NOR2X0 U14491 ( .IN1(n4318), .IN2(g145), .QN(n14368) );
  NAND2X0 U14492 ( .IN1(n14370), .IN2(n14371), .QN(n14356) );
  XNOR2X1 U14493 ( .IN1(n14372), .IN2(g113), .Q(n14371) );
  NAND2X0 U14494 ( .IN1(n14373), .IN2(n14374), .QN(n14372) );
  NAND2X0 U14495 ( .IN1(n9206), .IN2(g6313), .QN(n14374) );
  NOR2X0 U14496 ( .IN1(n14375), .IN2(n14376), .QN(n14373) );
  NOR2X0 U14497 ( .IN1(n4369), .IN2(g147), .QN(n14376) );
  NOR2X0 U14498 ( .IN1(n4318), .IN2(g148), .QN(n14375) );
  NOR2X0 U14499 ( .IN1(n14377), .IN2(n14378), .QN(n14370) );
  XNOR2X1 U14500 ( .IN1(n4290), .IN2(n14379), .Q(n14378) );
  NAND2X0 U14501 ( .IN1(n14380), .IN2(n14381), .QN(n14379) );
  NAND2X0 U14502 ( .IN1(n9200), .IN2(g6313), .QN(n14381) );
  NOR2X0 U14503 ( .IN1(n14382), .IN2(n14383), .QN(n14380) );
  NOR2X0 U14504 ( .IN1(n4369), .IN2(g156), .QN(n14383) );
  NOR2X0 U14505 ( .IN1(n4318), .IN2(g157), .QN(n14382) );
  XNOR2X1 U14506 ( .IN1(n4561), .IN2(n14384), .Q(n14377) );
  NAND2X0 U14507 ( .IN1(n14385), .IN2(n14386), .QN(n14384) );
  NAND2X0 U14508 ( .IN1(n9204), .IN2(g6313), .QN(n14386) );
  NOR2X0 U14509 ( .IN1(n14387), .IN2(n14388), .QN(n14385) );
  NOR2X0 U14510 ( .IN1(n4369), .IN2(g150), .QN(n14388) );
  NOR2X0 U14511 ( .IN1(n4318), .IN2(g151), .QN(n14387) );
  NAND2X0 U14512 ( .IN1(n14389), .IN2(n14390), .QN(g26616) );
  INVX0 U14513 ( .INP(n14391), .ZN(n14390) );
  NOR2X0 U14514 ( .IN1(g2624), .IN2(n8747), .QN(n14391) );
  NAND2X0 U14515 ( .IN1(n14392), .IN2(g2624), .QN(n14389) );
  NAND2X0 U14516 ( .IN1(n14393), .IN2(n14394), .QN(g26596) );
  NAND2X0 U14517 ( .IN1(n4370), .IN2(g2568), .QN(n14394) );
  NAND2X0 U14518 ( .IN1(n14392), .IN2(g7390), .QN(n14393) );
  NAND2X0 U14519 ( .IN1(n14395), .IN2(n14396), .QN(g26592) );
  NAND2X0 U14520 ( .IN1(n4366), .IN2(g1877), .QN(n14396) );
  NAND2X0 U14521 ( .IN1(n14397), .IN2(g1930), .QN(n14395) );
  NAND2X0 U14522 ( .IN1(n14398), .IN2(n14399), .QN(g26575) );
  INVX0 U14523 ( .INP(n14400), .ZN(n14399) );
  NOR2X0 U14524 ( .IN1(n11699), .IN2(n8745), .QN(n14400) );
  NAND2X0 U14525 ( .IN1(n14392), .IN2(n11699), .QN(n14398) );
  NOR2X0 U14526 ( .IN1(n14401), .IN2(n14402), .QN(n14392) );
  NAND2X0 U14527 ( .IN1(g2584), .IN2(n10100), .QN(n14401) );
  NAND2X0 U14528 ( .IN1(n14403), .IN2(n14404), .QN(g26573) );
  INVX0 U14529 ( .INP(n14405), .ZN(n14404) );
  NOR2X0 U14530 ( .IN1(g7194), .IN2(n8752), .QN(n14405) );
  NAND2X0 U14531 ( .IN1(n14397), .IN2(g7194), .QN(n14403) );
  NAND2X0 U14532 ( .IN1(n14406), .IN2(n14407), .QN(g26569) );
  INVX0 U14533 ( .INP(n14408), .ZN(n14407) );
  NOR2X0 U14534 ( .IN1(g1236), .IN2(n8749), .QN(n14408) );
  NAND2X0 U14535 ( .IN1(n14409), .IN2(g1236), .QN(n14406) );
  NAND2X0 U14536 ( .IN1(n14410), .IN2(n14411), .QN(g26559) );
  NAND2X0 U14537 ( .IN1(n14397), .IN2(n12749), .QN(n14411) );
  NOR2X0 U14538 ( .IN1(n14412), .IN2(n14413), .QN(n14397) );
  NAND2X0 U14539 ( .IN1(g1890), .IN2(n10237), .QN(n14412) );
  NAND2X0 U14540 ( .IN1(test_so68), .IN2(n4296), .QN(n14410) );
  NAND2X0 U14541 ( .IN1(n14414), .IN2(n14415), .QN(g26557) );
  INVX0 U14542 ( .INP(n14416), .ZN(n14415) );
  NOR2X0 U14543 ( .IN1(g6944), .IN2(n8753), .QN(n14416) );
  NAND2X0 U14544 ( .IN1(n14409), .IN2(g6944), .QN(n14414) );
  NAND2X0 U14545 ( .IN1(n14417), .IN2(n14418), .QN(g26553) );
  INVX0 U14546 ( .INP(n14419), .ZN(n14418) );
  NOR2X0 U14547 ( .IN1(g550), .IN2(n8750), .QN(n14419) );
  NAND2X0 U14548 ( .IN1(n14420), .IN2(g550), .QN(n14417) );
  NAND2X0 U14549 ( .IN1(n14421), .IN2(n14422), .QN(g26547) );
  NAND2X0 U14550 ( .IN1(n14409), .IN2(n12608), .QN(n14422) );
  NOR2X0 U14551 ( .IN1(n14423), .IN2(n14424), .QN(n14409) );
  NAND2X0 U14552 ( .IN1(g1196), .IN2(n10380), .QN(n14423) );
  NAND2X0 U14553 ( .IN1(test_so47), .IN2(n4371), .QN(n14421) );
  NAND2X0 U14554 ( .IN1(n14425), .IN2(n14426), .QN(g26545) );
  NAND2X0 U14555 ( .IN1(n4372), .IN2(g493), .QN(n14426) );
  NAND2X0 U14556 ( .IN1(n14420), .IN2(g6642), .QN(n14425) );
  NAND2X0 U14557 ( .IN1(n14427), .IN2(n14428), .QN(g26541) );
  INVX0 U14558 ( .INP(n14429), .ZN(n14428) );
  NOR2X0 U14559 ( .IN1(n13002), .IN2(n8746), .QN(n14429) );
  NAND2X0 U14560 ( .IN1(n14420), .IN2(n13002), .QN(n14427) );
  NOR2X0 U14561 ( .IN1(n14430), .IN2(n14431), .QN(n14420) );
  NAND2X0 U14562 ( .IN1(n9961), .IN2(test_so22), .QN(n14430) );
  NOR2X0 U14563 ( .IN1(n9702), .IN2(n14432), .QN(g26532) );
  XNOR2X1 U14564 ( .IN1(n4526), .IN2(n8971), .Q(n14432) );
  NOR2X0 U14565 ( .IN1(n9710), .IN2(n14433), .QN(g26531) );
  XNOR2X1 U14566 ( .IN1(n4527), .IN2(n8975), .Q(n14433) );
  NAND2X0 U14567 ( .IN1(n14434), .IN2(n14435), .QN(g26530) );
  INVX0 U14568 ( .INP(n14436), .ZN(n14435) );
  NOR2X0 U14569 ( .IN1(n14437), .IN2(n8979), .QN(n14436) );
  NAND2X0 U14570 ( .IN1(n14438), .IN2(n8979), .QN(n14434) );
  NOR2X0 U14571 ( .IN1(n11814), .IN2(n3690), .QN(n14438) );
  NOR2X0 U14572 ( .IN1(n9719), .IN2(n14439), .QN(g26529) );
  XNOR2X1 U14573 ( .IN1(n4528), .IN2(n8983), .Q(n14439) );
  NAND2X0 U14574 ( .IN1(n14440), .IN2(n14441), .QN(g26149) );
  NOR2X0 U14575 ( .IN1(n14442), .IN2(n14443), .QN(n14441) );
  NAND2X0 U14576 ( .IN1(n14444), .IN2(n14445), .QN(n14443) );
  NAND2X0 U14577 ( .IN1(n14446), .IN2(g3161), .QN(n14445) );
  NOR2X0 U14578 ( .IN1(n14447), .IN2(n14448), .QN(n14444) );
  NOR2X0 U14579 ( .IN1(n4338), .IN2(n14449), .QN(n14448) );
  NOR2X0 U14580 ( .IN1(n4441), .IN2(n14450), .QN(n14447) );
  NAND2X0 U14581 ( .IN1(n14451), .IN2(n14452), .QN(n14442) );
  NAND2X0 U14582 ( .IN1(n3936), .IN2(n14453), .QN(n14452) );
  NAND2X0 U14583 ( .IN1(n14454), .IN2(n14455), .QN(n14453) );
  NOR2X0 U14584 ( .IN1(n14456), .IN2(n14457), .QN(n14455) );
  NOR2X0 U14585 ( .IN1(n4339), .IN2(n14458), .QN(n14457) );
  NOR2X0 U14586 ( .IN1(n4341), .IN2(n14459), .QN(n14456) );
  NOR2X0 U14587 ( .IN1(n14460), .IN2(n14461), .QN(n14454) );
  NOR2X0 U14588 ( .IN1(n4453), .IN2(n14462), .QN(n14461) );
  NOR2X0 U14589 ( .IN1(n4436), .IN2(n14463), .QN(n14460) );
  NOR2X0 U14590 ( .IN1(n14464), .IN2(n14465), .QN(n14451) );
  NOR2X0 U14591 ( .IN1(n14466), .IN2(n14467), .QN(n14465) );
  NOR2X0 U14592 ( .IN1(n14468), .IN2(n14469), .QN(n14466) );
  NAND2X0 U14593 ( .IN1(n14470), .IN2(n14471), .QN(n14469) );
  NAND2X0 U14594 ( .IN1(test_so8), .IN2(n14472), .QN(n14471) );
  NAND2X0 U14595 ( .IN1(n14473), .IN2(g3155), .QN(n14470) );
  NOR2X0 U14596 ( .IN1(n4442), .IN2(n14474), .QN(n14468) );
  NOR2X0 U14597 ( .IN1(n4348), .IN2(n14475), .QN(n14464) );
  NOR2X0 U14598 ( .IN1(n14476), .IN2(n14477), .QN(n14440) );
  NAND2X0 U14599 ( .IN1(n3700), .IN2(n14478), .QN(n14477) );
  NAND2X0 U14600 ( .IN1(n13293), .IN2(n8086), .QN(n14478) );
  NAND2X0 U14601 ( .IN1(n14479), .IN2(n14480), .QN(n14476) );
  NAND2X0 U14602 ( .IN1(n14481), .IN2(n8080), .QN(n14480) );
  INVX0 U14603 ( .INP(n14482), .ZN(n14481) );
  NOR2X0 U14604 ( .IN1(n14483), .IN2(n14484), .QN(n14479) );
  NOR2X0 U14605 ( .IN1(n4450), .IN2(n14485), .QN(n14484) );
  NOR2X0 U14606 ( .IN1(n13292), .IN2(DFF_156_n1), .QN(n14483) );
  NAND2X0 U14607 ( .IN1(n14486), .IN2(n14487), .QN(g26135) );
  NOR2X0 U14608 ( .IN1(n14488), .IN2(n14489), .QN(n14487) );
  NAND2X0 U14609 ( .IN1(n14490), .IN2(n14491), .QN(n14489) );
  NAND2X0 U14610 ( .IN1(n14492), .IN2(n13285), .QN(n14491) );
  NOR2X0 U14611 ( .IN1(n14493), .IN2(n14494), .QN(n14490) );
  NOR2X0 U14612 ( .IN1(n14475), .IN2(n9288), .QN(n14494) );
  NOR2X0 U14613 ( .IN1(n14495), .IN2(g3128), .QN(n14493) );
  NAND2X0 U14614 ( .IN1(n14496), .IN2(n14497), .QN(n14488) );
  NOR2X0 U14615 ( .IN1(n14498), .IN2(n14499), .QN(n14497) );
  NOR2X0 U14616 ( .IN1(n13292), .IN2(DFF_155_n1), .QN(n14499) );
  NOR2X0 U14617 ( .IN1(n4443), .IN2(n14500), .QN(n14498) );
  NOR2X0 U14618 ( .IN1(n14501), .IN2(n14502), .QN(n14496) );
  NOR2X0 U14619 ( .IN1(n16831), .IN2(n14482), .QN(n14502) );
  NOR2X0 U14620 ( .IN1(n4452), .IN2(n14485), .QN(n14501) );
  NOR2X0 U14621 ( .IN1(n14503), .IN2(n14504), .QN(n14486) );
  NAND2X0 U14622 ( .IN1(n14505), .IN2(n3700), .QN(n14504) );
  NOR2X0 U14623 ( .IN1(n14506), .IN2(n14507), .QN(n14505) );
  NOR2X0 U14624 ( .IN1(n4447), .IN2(n14449), .QN(n14507) );
  NOR2X0 U14625 ( .IN1(n4343), .IN2(n14450), .QN(n14506) );
  NAND2X0 U14626 ( .IN1(n14508), .IN2(n14509), .QN(n14503) );
  NAND2X0 U14627 ( .IN1(n3936), .IN2(n14510), .QN(n14509) );
  NAND2X0 U14628 ( .IN1(n14511), .IN2(n14512), .QN(n14510) );
  NOR2X0 U14629 ( .IN1(n14513), .IN2(n14514), .QN(n14512) );
  NOR2X0 U14630 ( .IN1(n4342), .IN2(n14458), .QN(n14514) );
  NOR2X0 U14631 ( .IN1(n4334), .IN2(n14459), .QN(n14513) );
  NOR2X0 U14632 ( .IN1(n14515), .IN2(n14516), .QN(n14511) );
  NOR2X0 U14633 ( .IN1(n4438), .IN2(n14462), .QN(n14516) );
  NOR2X0 U14634 ( .IN1(n4434), .IN2(n14463), .QN(n14515) );
  NOR2X0 U14635 ( .IN1(n14517), .IN2(n14518), .QN(n14508) );
  NOR2X0 U14636 ( .IN1(n14519), .IN2(n14467), .QN(n14518) );
  NOR2X0 U14637 ( .IN1(n14520), .IN2(n14521), .QN(n14519) );
  NAND2X0 U14638 ( .IN1(n14522), .IN2(n14523), .QN(n14521) );
  NAND2X0 U14639 ( .IN1(n14472), .IN2(g3105), .QN(n14523) );
  NAND2X0 U14640 ( .IN1(n14473), .IN2(g3097), .QN(n14522) );
  NOR2X0 U14641 ( .IN1(n4437), .IN2(n14474), .QN(n14520) );
  NOR2X0 U14642 ( .IN1(n13276), .IN2(n9287), .QN(n14517) );
  NAND2X0 U14643 ( .IN1(n14524), .IN2(n14525), .QN(g26104) );
  NOR2X0 U14644 ( .IN1(n14526), .IN2(n14527), .QN(n14525) );
  NAND2X0 U14645 ( .IN1(n14528), .IN2(n14529), .QN(n14527) );
  INVX0 U14646 ( .INP(n14530), .ZN(n14529) );
  NOR2X0 U14647 ( .IN1(n14449), .IN2(n4448), .QN(n14530) );
  NAND2X0 U14648 ( .IN1(n14531), .IN2(n3933), .QN(n14449) );
  NOR2X0 U14649 ( .IN1(g3201), .IN2(n13274), .QN(n14531) );
  NOR2X0 U14650 ( .IN1(n14532), .IN2(n14533), .QN(n14528) );
  NOR2X0 U14651 ( .IN1(n4344), .IN2(n14450), .QN(n14533) );
  NAND2X0 U14652 ( .IN1(n14534), .IN2(n4329), .QN(n14450) );
  NOR2X0 U14653 ( .IN1(n14535), .IN2(n14536), .QN(n14532) );
  INVX0 U14654 ( .INP(n3936), .ZN(n14536) );
  NOR2X0 U14655 ( .IN1(n14537), .IN2(n14538), .QN(n14535) );
  NAND2X0 U14656 ( .IN1(n14539), .IN2(n14540), .QN(n14538) );
  NAND2X0 U14657 ( .IN1(n14541), .IN2(g3211), .QN(n14540) );
  NAND2X0 U14658 ( .IN1(n13269), .IN2(g3094), .QN(n14539) );
  INVX0 U14659 ( .INP(n14542), .ZN(n14537) );
  NOR2X0 U14660 ( .IN1(n14543), .IN2(n14544), .QN(n14542) );
  NOR2X0 U14661 ( .IN1(n14459), .IN2(n4336), .QN(n14544) );
  NAND2X0 U14662 ( .IN1(g3207), .IN2(g3201), .QN(n14459) );
  NOR2X0 U14663 ( .IN1(n14458), .IN2(n4340), .QN(n14543) );
  NAND2X0 U14664 ( .IN1(n4406), .IN2(g3207), .QN(n14458) );
  NAND2X0 U14665 ( .IN1(n14545), .IN2(n14546), .QN(n14526) );
  NOR2X0 U14666 ( .IN1(n14547), .IN2(n14548), .QN(n14546) );
  NOR2X0 U14667 ( .IN1(n13283), .IN2(n13278), .QN(n14548) );
  INVX0 U14668 ( .INP(n14492), .ZN(n13278) );
  NOR2X0 U14669 ( .IN1(n13271), .IN2(n14549), .QN(n14492) );
  INVX0 U14670 ( .INP(n14550), .ZN(n13283) );
  NOR2X0 U14671 ( .IN1(n4337), .IN2(n14475), .QN(n14547) );
  NAND2X0 U14672 ( .IN1(n14551), .IN2(n14473), .QN(n14475) );
  NOR2X0 U14673 ( .IN1(n14552), .IN2(n14553), .QN(n14545) );
  NOR2X0 U14674 ( .IN1(n14554), .IN2(n14467), .QN(n14553) );
  NOR2X0 U14675 ( .IN1(n14555), .IN2(n14556), .QN(n14554) );
  NAND2X0 U14676 ( .IN1(n14557), .IN2(n14558), .QN(n14556) );
  NAND2X0 U14677 ( .IN1(n14472), .IN2(g3093), .QN(n14558) );
  NAND2X0 U14678 ( .IN1(test_so6), .IN2(n14473), .QN(n14557) );
  NOR2X0 U14679 ( .IN1(n4439), .IN2(n14474), .QN(n14555) );
  NOR2X0 U14680 ( .IN1(n4301), .IN2(n13276), .QN(n14552) );
  NAND2X0 U14681 ( .IN1(n14559), .IN2(n4073), .QN(n13276) );
  NOR2X0 U14682 ( .IN1(n9254), .IN2(n14474), .QN(n14559) );
  NOR2X0 U14683 ( .IN1(n14560), .IN2(n14561), .QN(n14524) );
  NAND2X0 U14684 ( .IN1(n14562), .IN2(n3700), .QN(n14561) );
  NOR2X0 U14685 ( .IN1(n14563), .IN2(n14564), .QN(n14562) );
  NOR2X0 U14686 ( .IN1(n14495), .IN2(DFF_140_n1), .QN(n14564) );
  NOR2X0 U14687 ( .IN1(n16830), .IN2(n14482), .QN(n14563) );
  NAND2X0 U14688 ( .IN1(n14565), .IN2(n14566), .QN(n14560) );
  INVX0 U14689 ( .INP(n14567), .ZN(n14566) );
  NOR2X0 U14690 ( .IN1(n14485), .IN2(n4451), .QN(n14567) );
  NAND2X0 U14691 ( .IN1(n14534), .IN2(g3207), .QN(n14485) );
  NOR2X0 U14692 ( .IN1(n14568), .IN2(n13274), .QN(n14534) );
  INVX0 U14693 ( .INP(n14551), .ZN(n13274) );
  NOR2X0 U14694 ( .IN1(n10481), .IN2(n9254), .QN(n14551) );
  NAND2X0 U14695 ( .IN1(n296), .IN2(g3197), .QN(n10481) );
  INVX0 U14696 ( .INP(n14569), .ZN(n296) );
  NAND2X0 U14697 ( .IN1(n14570), .IN2(n16824), .QN(n14569) );
  NOR2X0 U14698 ( .IN1(n8088), .IN2(n8090), .QN(n14570) );
  NAND2X0 U14699 ( .IN1(g3188), .IN2(n4406), .QN(n14568) );
  NOR2X0 U14700 ( .IN1(n14571), .IN2(n14572), .QN(n14565) );
  NOR2X0 U14701 ( .IN1(n16832), .IN2(n13292), .QN(n14572) );
  NAND2X0 U14702 ( .IN1(n14573), .IN2(n4073), .QN(n13292) );
  NOR2X0 U14703 ( .IN1(n9254), .IN2(n13286), .QN(n14573) );
  INVX0 U14704 ( .INP(n14472), .ZN(n13286) );
  NOR2X0 U14705 ( .IN1(n14462), .IN2(g3188), .QN(n14472) );
  INVX0 U14706 ( .INP(n13269), .ZN(n14462) );
  NOR2X0 U14707 ( .IN1(g3207), .IN2(n4406), .QN(n13269) );
  NOR2X0 U14708 ( .IN1(n4445), .IN2(n14500), .QN(n14571) );
  INVX0 U14709 ( .INP(n14446), .ZN(n14500) );
  NOR2X0 U14710 ( .IN1(n14574), .IN2(n14467), .QN(n14446) );
  INVX0 U14711 ( .INP(n3939), .ZN(n14467) );
  NAND2X0 U14712 ( .IN1(n4406), .IN2(n3933), .QN(n14574) );
  NOR2X0 U14713 ( .IN1(g3188), .IN2(n4329), .QN(n3933) );
  NAND2X0 U14714 ( .IN1(n9931), .IN2(n14575), .QN(g26048) );
  NAND2X0 U14715 ( .IN1(n14576), .IN2(n14577), .QN(n14575) );
  XNOR2X1 U14716 ( .IN1(n16834), .IN2(n14578), .Q(n14576) );
  NOR2X0 U14717 ( .IN1(n9867), .IN2(n14579), .QN(g26037) );
  XNOR2X1 U14718 ( .IN1(g2900), .IN2(n9679), .Q(n14579) );
  NOR2X0 U14719 ( .IN1(n4058), .IN2(n4305), .QN(n9679) );
  NAND2X0 U14720 ( .IN1(n9689), .IN2(g2892), .QN(n4058) );
  NOR2X0 U14721 ( .IN1(n14580), .IN2(n14097), .QN(g26031) );
  XNOR2X1 U14722 ( .IN1(n9280), .IN2(n3742), .Q(n14580) );
  NAND2X0 U14723 ( .IN1(n4065), .IN2(g3013), .QN(n3742) );
  NAND2X0 U14724 ( .IN1(n14581), .IN2(n14582), .QN(g26025) );
  NAND2X0 U14725 ( .IN1(test_so82), .IN2(n14583), .QN(n14582) );
  NAND2X0 U14726 ( .IN1(n14110), .IN2(n11841), .QN(n14583) );
  NAND2X0 U14727 ( .IN1(n14111), .IN2(n11841), .QN(n14581) );
  INVX0 U14728 ( .INP(n4509), .ZN(n11841) );
  NOR2X0 U14729 ( .IN1(n9281), .IN2(n14110), .QN(n14111) );
  INVX0 U14730 ( .INP(n3749), .ZN(n14110) );
  NAND2X0 U14731 ( .IN1(n14584), .IN2(test_so79), .QN(n3749) );
  NOR2X0 U14732 ( .IN1(n11938), .IN2(n11766), .QN(n14584) );
  NAND2X0 U14733 ( .IN1(n14585), .IN2(n14586), .QN(n11766) );
  NAND2X0 U14734 ( .IN1(n8936), .IN2(n10669), .QN(n14586) );
  NOR2X0 U14735 ( .IN1(n14587), .IN2(n14588), .QN(n14585) );
  NOR2X0 U14736 ( .IN1(n4516), .IN2(g2478), .QN(n14588) );
  NOR2X0 U14737 ( .IN1(test_so82), .IN2(n4509), .QN(n14587) );
  NAND2X0 U14738 ( .IN1(n14589), .IN2(n14590), .QN(n11938) );
  NOR2X0 U14739 ( .IN1(n14591), .IN2(n14592), .QN(n14590) );
  NAND2X0 U14740 ( .IN1(n14593), .IN2(n14594), .QN(n14592) );
  XNOR2X1 U14741 ( .IN1(n14595), .IN2(g2165), .Q(n14594) );
  NAND2X0 U14742 ( .IN1(n14596), .IN2(n14597), .QN(n14595) );
  NAND2X0 U14743 ( .IN1(n9169), .IN2(test_so73), .QN(n14597) );
  NOR2X0 U14744 ( .IN1(n14598), .IN2(n14599), .QN(n14596) );
  NOR2X0 U14745 ( .IN1(n4367), .IN2(g2205), .QN(n14599) );
  NOR2X0 U14746 ( .IN1(n4324), .IN2(g2206), .QN(n14598) );
  NOR2X0 U14747 ( .IN1(n14600), .IN2(n14601), .QN(n14593) );
  XNOR2X1 U14748 ( .IN1(n4373), .IN2(n14602), .Q(n14601) );
  NAND2X0 U14749 ( .IN1(n14603), .IN2(n14604), .QN(n14602) );
  NAND2X0 U14750 ( .IN1(n9167), .IN2(test_so73), .QN(n14604) );
  NOR2X0 U14751 ( .IN1(n14605), .IN2(n14606), .QN(n14603) );
  NOR2X0 U14752 ( .IN1(n4367), .IN2(g2208), .QN(n14606) );
  NOR2X0 U14753 ( .IN1(n4324), .IN2(g2209), .QN(n14605) );
  XNOR2X1 U14754 ( .IN1(n4319), .IN2(n14607), .Q(n14600) );
  NAND2X0 U14755 ( .IN1(n14608), .IN2(n14609), .QN(n14607) );
  NAND2X0 U14756 ( .IN1(n9165), .IN2(test_so73), .QN(n14609) );
  NOR2X0 U14757 ( .IN1(n14610), .IN2(n14611), .QN(n14608) );
  NOR2X0 U14758 ( .IN1(n4367), .IN2(g2217), .QN(n14611) );
  NOR2X0 U14759 ( .IN1(n4324), .IN2(g2218), .QN(n14610) );
  NAND2X0 U14760 ( .IN1(n14612), .IN2(n14613), .QN(n14591) );
  XNOR2X1 U14761 ( .IN1(n10796), .IN2(n14614), .Q(n14613) );
  NOR2X0 U14762 ( .IN1(n14615), .IN2(n14616), .QN(n14614) );
  NAND2X0 U14763 ( .IN1(n14617), .IN2(n14618), .QN(n14616) );
  NAND2X0 U14764 ( .IN1(n8794), .IN2(g6837), .QN(n14618) );
  NAND2X0 U14765 ( .IN1(n8793), .IN2(g2241), .QN(n14617) );
  NOR2X0 U14766 ( .IN1(test_so75), .IN2(n9278), .QN(n14615) );
  NOR2X0 U14767 ( .IN1(n11127), .IN2(n14619), .QN(n14612) );
  XNOR2X1 U14768 ( .IN1(n10978), .IN2(n14620), .Q(n14619) );
  NAND2X0 U14769 ( .IN1(n14621), .IN2(n14622), .QN(n14620) );
  NAND2X0 U14770 ( .IN1(n8785), .IN2(test_so73), .QN(n14622) );
  NOR2X0 U14771 ( .IN1(n14623), .IN2(n14624), .QN(n14621) );
  NOR2X0 U14772 ( .IN1(n4367), .IN2(g2235), .QN(n14624) );
  NOR2X0 U14773 ( .IN1(n4324), .IN2(g2236), .QN(n14623) );
  INVX0 U14774 ( .INP(n3038), .ZN(n11127) );
  NOR2X0 U14775 ( .IN1(n14625), .IN2(n14626), .QN(n14589) );
  NAND2X0 U14776 ( .IN1(n14627), .IN2(n14628), .QN(n14626) );
  XNOR2X1 U14777 ( .IN1(n14629), .IN2(g2195), .Q(n14628) );
  NAND2X0 U14778 ( .IN1(n14630), .IN2(n14631), .QN(n14629) );
  NAND2X0 U14779 ( .IN1(n9158), .IN2(test_so73), .QN(n14631) );
  NOR2X0 U14780 ( .IN1(n14632), .IN2(n14633), .QN(n14630) );
  NOR2X0 U14781 ( .IN1(n4367), .IN2(g2229), .QN(n14633) );
  NOR2X0 U14782 ( .IN1(n4324), .IN2(g2230), .QN(n14632) );
  XNOR2X1 U14783 ( .IN1(n14634), .IN2(g2180), .Q(n14627) );
  NAND2X0 U14784 ( .IN1(n14635), .IN2(n14636), .QN(n14634) );
  NAND2X0 U14785 ( .IN1(n9163), .IN2(test_so73), .QN(n14636) );
  NOR2X0 U14786 ( .IN1(n14637), .IN2(n14638), .QN(n14635) );
  NOR2X0 U14787 ( .IN1(n4367), .IN2(g2220), .QN(n14638) );
  NOR2X0 U14788 ( .IN1(n4324), .IN2(g2221), .QN(n14637) );
  NAND2X0 U14789 ( .IN1(n14639), .IN2(n14640), .QN(n14625) );
  XNOR2X1 U14790 ( .IN1(n14641), .IN2(g2185), .Q(n14640) );
  NAND2X0 U14791 ( .IN1(n14642), .IN2(n14643), .QN(n14641) );
  INVX0 U14792 ( .INP(n14644), .ZN(n14643) );
  NOR2X0 U14793 ( .IN1(n9278), .IN2(test_so74), .QN(n14644) );
  NOR2X0 U14794 ( .IN1(n14645), .IN2(n14646), .QN(n14642) );
  NOR2X0 U14795 ( .IN1(n4367), .IN2(g2223), .QN(n14646) );
  NOR2X0 U14796 ( .IN1(n4324), .IN2(g2224), .QN(n14645) );
  NOR2X0 U14797 ( .IN1(n14647), .IN2(n14648), .QN(n14639) );
  XNOR2X1 U14798 ( .IN1(n4287), .IN2(n14649), .Q(n14648) );
  NAND2X0 U14799 ( .IN1(n14650), .IN2(n14651), .QN(n14649) );
  NAND2X0 U14800 ( .IN1(n9156), .IN2(test_so73), .QN(n14651) );
  NOR2X0 U14801 ( .IN1(n14652), .IN2(n14653), .QN(n14650) );
  NOR2X0 U14802 ( .IN1(n4367), .IN2(g2232), .QN(n14653) );
  NOR2X0 U14803 ( .IN1(n4324), .IN2(g2233), .QN(n14652) );
  XNOR2X1 U14804 ( .IN1(n4555), .IN2(n14654), .Q(n14647) );
  NAND2X0 U14805 ( .IN1(n14655), .IN2(n14656), .QN(n14654) );
  NAND2X0 U14806 ( .IN1(n9160), .IN2(test_so73), .QN(n14656) );
  NOR2X0 U14807 ( .IN1(n14657), .IN2(n14658), .QN(n14655) );
  NOR2X0 U14808 ( .IN1(n4367), .IN2(g2226), .QN(n14658) );
  NOR2X0 U14809 ( .IN1(n4324), .IN2(g2227), .QN(n14657) );
  NOR2X0 U14810 ( .IN1(n14659), .IN2(n14437), .QN(g25935) );
  NAND2X0 U14811 ( .IN1(n3690), .IN2(n12389), .QN(n14437) );
  INVX0 U14812 ( .INP(n11814), .ZN(n12389) );
  NAND2X0 U14813 ( .IN1(n3893), .IN2(g776), .QN(n3690) );
  NOR2X0 U14814 ( .IN1(n3893), .IN2(g776), .QN(n14659) );
  NAND2X0 U14815 ( .IN1(n14660), .IN2(n14661), .QN(g25489) );
  NAND2X0 U14816 ( .IN1(n14662), .IN2(n14663), .QN(n14661) );
  NOR2X0 U14817 ( .IN1(n4433), .IN2(n4424), .QN(n14663) );
  NOR2X0 U14818 ( .IN1(n4301), .IN2(n14664), .QN(n14662) );
  NAND2X0 U14819 ( .IN1(n14665), .IN2(n9287), .QN(n14660) );
  NAND2X0 U14820 ( .IN1(n14664), .IN2(n14666), .QN(n14665) );
  NAND2X0 U14821 ( .IN1(n4301), .IN2(n14550), .QN(n14666) );
  NAND2X0 U14822 ( .IN1(DFF_15_n1), .IN2(DFF_16_n1), .QN(n14550) );
  NOR2X0 U14823 ( .IN1(test_so10), .IN2(n14667), .QN(n14664) );
  INVX0 U14824 ( .INP(n14668), .ZN(n14667) );
  NAND2X0 U14825 ( .IN1(n4424), .IN2(n14669), .QN(n14668) );
  INVX0 U14826 ( .INP(n14670), .ZN(n14669) );
  NOR2X0 U14827 ( .IN1(n13285), .IN2(n4301), .QN(n14670) );
  NAND2X0 U14828 ( .IN1(n8698), .IN2(n8697), .QN(n13285) );
  NAND2X0 U14829 ( .IN1(n14671), .IN2(n14672), .QN(g25452) );
  INVX0 U14830 ( .INP(n14673), .ZN(n14672) );
  NOR2X0 U14831 ( .IN1(g3109), .IN2(n4443), .QN(n14673) );
  NAND2X0 U14832 ( .IN1(g21851), .IN2(g3109), .QN(n14671) );
  NAND2X0 U14833 ( .IN1(n14674), .IN2(n14675), .QN(g25451) );
  INVX0 U14834 ( .INP(n14676), .ZN(n14675) );
  NOR2X0 U14835 ( .IN1(g8030), .IN2(n4434), .QN(n14676) );
  NAND2X0 U14836 ( .IN1(g21851), .IN2(g8030), .QN(n14674) );
  NAND2X0 U14837 ( .IN1(n14677), .IN2(n14678), .QN(g25450) );
  NAND2X0 U14838 ( .IN1(n4382), .IN2(g3097), .QN(n14678) );
  NAND2X0 U14839 ( .IN1(g21851), .IN2(g8106), .QN(n14677) );
  NAND2X0 U14840 ( .IN1(n14679), .IN2(n3700), .QN(g25442) );
  NOR2X0 U14841 ( .IN1(n14680), .IN2(n14681), .QN(n14679) );
  NOR2X0 U14842 ( .IN1(n8597), .IN2(n14495), .QN(n14681) );
  NOR2X0 U14843 ( .IN1(n8598), .IN2(n14482), .QN(n14680) );
  NAND2X0 U14844 ( .IN1(n14682), .IN2(n3700), .QN(g25435) );
  NOR2X0 U14845 ( .IN1(n14683), .IN2(n14684), .QN(n14682) );
  NOR2X0 U14846 ( .IN1(n14495), .IN2(n8084), .QN(n14684) );
  NOR2X0 U14847 ( .IN1(n8563), .IN2(n14482), .QN(n14683) );
  NAND2X0 U14848 ( .IN1(n14685), .IN2(n3700), .QN(g25420) );
  NOR2X0 U14849 ( .IN1(n14686), .IN2(n14687), .QN(n14685) );
  NOR2X0 U14850 ( .IN1(n14495), .IN2(n8595), .QN(n14687) );
  INVX0 U14851 ( .INP(n13293), .ZN(n14495) );
  NOR2X0 U14852 ( .IN1(n8596), .IN2(n14482), .QN(n14686) );
  NAND2X0 U14853 ( .IN1(n14688), .IN2(n4073), .QN(n14482) );
  NOR2X0 U14854 ( .IN1(n9254), .IN2(n14549), .QN(n14688) );
  INVX0 U14855 ( .INP(n14473), .ZN(n14549) );
  NOR2X0 U14856 ( .IN1(g3188), .IN2(n14463), .QN(n14473) );
  INVX0 U14857 ( .INP(n14541), .ZN(n14463) );
  NOR2X0 U14858 ( .IN1(g3201), .IN2(g3207), .QN(n14541) );
  NAND2X0 U14859 ( .IN1(n14689), .IN2(n14690), .QN(g25288) );
  NAND2X0 U14860 ( .IN1(n14691), .IN2(g2808), .QN(n14690) );
  NAND2X0 U14861 ( .IN1(n14692), .IN2(n14693), .QN(n14689) );
  NAND2X0 U14862 ( .IN1(n14694), .IN2(n14695), .QN(g25280) );
  NAND2X0 U14863 ( .IN1(n14696), .IN2(g2810), .QN(n14695) );
  NAND2X0 U14864 ( .IN1(n14697), .IN2(n14692), .QN(n14694) );
  NAND2X0 U14865 ( .IN1(n14698), .IN2(n14699), .QN(g25279) );
  NAND2X0 U14866 ( .IN1(n14700), .IN2(g2114), .QN(n14699) );
  NAND2X0 U14867 ( .IN1(n14701), .IN2(n14702), .QN(n14698) );
  NAND2X0 U14868 ( .IN1(n14703), .IN2(n14704), .QN(g25272) );
  NAND2X0 U14869 ( .IN1(n10624), .IN2(g2809), .QN(n14704) );
  NAND2X0 U14870 ( .IN1(n14705), .IN2(n14692), .QN(n14703) );
  INVX0 U14871 ( .INP(n14706), .ZN(n14692) );
  NAND2X0 U14872 ( .IN1(n14707), .IN2(n14708), .QN(n14706) );
  NOR2X0 U14873 ( .IN1(n14709), .IN2(n14710), .QN(n14708) );
  NAND2X0 U14874 ( .IN1(n14711), .IN2(n14712), .QN(n14710) );
  NAND2X0 U14875 ( .IN1(n14713), .IN2(n14714), .QN(n14712) );
  NOR2X0 U14876 ( .IN1(n14715), .IN2(n14716), .QN(n14714) );
  NAND2X0 U14877 ( .IN1(n14717), .IN2(n14718), .QN(n14716) );
  XNOR2X1 U14878 ( .IN1(n10117), .IN2(n4408), .Q(n14718) );
  INVX0 U14879 ( .INP(n10118), .ZN(n10117) );
  NAND2X0 U14880 ( .IN1(n14719), .IN2(n14720), .QN(n10118) );
  NAND2X0 U14881 ( .IN1(n9052), .IN2(g7487), .QN(n14720) );
  NOR2X0 U14882 ( .IN1(n14721), .IN2(n14722), .QN(n14719) );
  NOR2X0 U14883 ( .IN1(n4306), .IN2(g2782), .QN(n14722) );
  NOR2X0 U14884 ( .IN1(test_so93), .IN2(n4292), .QN(n14721) );
  XNOR2X1 U14885 ( .IN1(n10146), .IN2(n4407), .Q(n14717) );
  INVX0 U14886 ( .INP(n10148), .ZN(n10146) );
  NAND2X0 U14887 ( .IN1(n14723), .IN2(n14724), .QN(n10148) );
  NAND2X0 U14888 ( .IN1(n9048), .IN2(g7487), .QN(n14724) );
  NOR2X0 U14889 ( .IN1(n14725), .IN2(n14726), .QN(n14723) );
  NOR2X0 U14890 ( .IN1(n4306), .IN2(g2788), .QN(n14726) );
  NOR2X0 U14891 ( .IN1(n4292), .IN2(g2787), .QN(n14725) );
  NAND2X0 U14892 ( .IN1(n14727), .IN2(n14728), .QN(n14715) );
  XNOR2X1 U14893 ( .IN1(n10089), .IN2(n4415), .Q(n14728) );
  INVX0 U14894 ( .INP(n10092), .ZN(n10089) );
  NAND2X0 U14895 ( .IN1(n14729), .IN2(n14730), .QN(n10092) );
  NAND2X0 U14896 ( .IN1(n9040), .IN2(g7487), .QN(n14730) );
  NOR2X0 U14897 ( .IN1(n14731), .IN2(n14732), .QN(n14729) );
  NOR2X0 U14898 ( .IN1(n4306), .IN2(g2800), .QN(n14732) );
  NOR2X0 U14899 ( .IN1(n4292), .IN2(g2799), .QN(n14731) );
  NOR2X0 U14900 ( .IN1(n14733), .IN2(n14734), .QN(n14727) );
  XNOR2X1 U14901 ( .IN1(n4393), .IN2(n10099), .Q(n14734) );
  NAND2X0 U14902 ( .IN1(n14735), .IN2(n14736), .QN(n10099) );
  NAND2X0 U14903 ( .IN1(n9042), .IN2(g7487), .QN(n14736) );
  NOR2X0 U14904 ( .IN1(n14737), .IN2(n14738), .QN(n14735) );
  NOR2X0 U14905 ( .IN1(n4306), .IN2(g2797), .QN(n14738) );
  NOR2X0 U14906 ( .IN1(test_so94), .IN2(n4292), .QN(n14737) );
  XNOR2X1 U14907 ( .IN1(n10136), .IN2(test_so92), .Q(n14733) );
  INVX0 U14908 ( .INP(n10137), .ZN(n10136) );
  NAND2X0 U14909 ( .IN1(n14739), .IN2(n14740), .QN(n10137) );
  NAND2X0 U14910 ( .IN1(n9046), .IN2(g7487), .QN(n14740) );
  NOR2X0 U14911 ( .IN1(n14741), .IN2(n14742), .QN(n14739) );
  NOR2X0 U14912 ( .IN1(n4306), .IN2(g2791), .QN(n14742) );
  NOR2X0 U14913 ( .IN1(n4292), .IN2(g2790), .QN(n14741) );
  NOR2X0 U14914 ( .IN1(n14743), .IN2(n14744), .QN(n14713) );
  NAND2X0 U14915 ( .IN1(n14745), .IN2(n14746), .QN(n14744) );
  XNOR2X1 U14916 ( .IN1(n10156), .IN2(n4419), .Q(n14746) );
  INVX0 U14917 ( .INP(n10157), .ZN(n10156) );
  NAND2X0 U14918 ( .IN1(n14747), .IN2(n14748), .QN(n10157) );
  NAND2X0 U14919 ( .IN1(n9054), .IN2(g7487), .QN(n14748) );
  NOR2X0 U14920 ( .IN1(n14749), .IN2(n14750), .QN(n14747) );
  NOR2X0 U14921 ( .IN1(n4306), .IN2(g2779), .QN(n14750) );
  NOR2X0 U14922 ( .IN1(n4292), .IN2(g2778), .QN(n14749) );
  XNOR2X1 U14923 ( .IN1(n10128), .IN2(n4472), .Q(n14745) );
  INVX0 U14924 ( .INP(n10129), .ZN(n10128) );
  NAND2X0 U14925 ( .IN1(n14751), .IN2(n14752), .QN(n10129) );
  NAND2X0 U14926 ( .IN1(n9056), .IN2(g7487), .QN(n14752) );
  NOR2X0 U14927 ( .IN1(n14753), .IN2(n14754), .QN(n14751) );
  NOR2X0 U14928 ( .IN1(n4306), .IN2(g2776), .QN(n14754) );
  NOR2X0 U14929 ( .IN1(n4292), .IN2(g2775), .QN(n14753) );
  NAND2X0 U14930 ( .IN1(n14755), .IN2(n14756), .QN(n14743) );
  XNOR2X1 U14931 ( .IN1(n10122), .IN2(n4471), .Q(n14756) );
  INVX0 U14932 ( .INP(n10123), .ZN(n10122) );
  NAND2X0 U14933 ( .IN1(n14757), .IN2(n14758), .QN(n10123) );
  NAND2X0 U14934 ( .IN1(n9044), .IN2(g7487), .QN(n14758) );
  NOR2X0 U14935 ( .IN1(n14759), .IN2(n14760), .QN(n14757) );
  NOR2X0 U14936 ( .IN1(n4306), .IN2(g2794), .QN(n14760) );
  NOR2X0 U14937 ( .IN1(n4292), .IN2(g2793), .QN(n14759) );
  NOR2X0 U14938 ( .IN1(n14761), .IN2(n14762), .QN(n14755) );
  XNOR2X1 U14939 ( .IN1(n4398), .IN2(n10142), .Q(n14762) );
  NAND2X0 U14940 ( .IN1(n14763), .IN2(n14764), .QN(n10142) );
  NAND2X0 U14941 ( .IN1(n9058), .IN2(g7487), .QN(n14764) );
  NOR2X0 U14942 ( .IN1(n14765), .IN2(n14766), .QN(n14763) );
  NOR2X0 U14943 ( .IN1(n4306), .IN2(g2773), .QN(n14766) );
  NOR2X0 U14944 ( .IN1(n4292), .IN2(g2772), .QN(n14765) );
  XNOR2X1 U14945 ( .IN1(n4397), .IN2(n10113), .Q(n14761) );
  NAND2X0 U14946 ( .IN1(n14767), .IN2(n14768), .QN(n10113) );
  NAND2X0 U14947 ( .IN1(n9050), .IN2(g7487), .QN(n14768) );
  NOR2X0 U14948 ( .IN1(n14769), .IN2(n14770), .QN(n14767) );
  NOR2X0 U14949 ( .IN1(n4306), .IN2(g2785), .QN(n14770) );
  NOR2X0 U14950 ( .IN1(n4292), .IN2(g2784), .QN(n14769) );
  NAND2X0 U14951 ( .IN1(n8896), .IN2(g2703), .QN(n14711) );
  NOR2X0 U14952 ( .IN1(n4306), .IN2(g2803), .QN(n14709) );
  NOR2X0 U14953 ( .IN1(n14771), .IN2(n10636), .QN(n14707) );
  NAND2X0 U14954 ( .IN1(n14772), .IN2(n14773), .QN(n10636) );
  NAND2X0 U14955 ( .IN1(n8837), .IN2(g7487), .QN(n14773) );
  NOR2X0 U14956 ( .IN1(n14774), .IN2(n14775), .QN(n14772) );
  NOR2X0 U14957 ( .IN1(n4306), .IN2(g2806), .QN(n14775) );
  NOR2X0 U14958 ( .IN1(n4292), .IN2(g2805), .QN(n14774) );
  NOR2X0 U14959 ( .IN1(n4356), .IN2(g2804), .QN(n14771) );
  NAND2X0 U14960 ( .IN1(n14776), .IN2(n14777), .QN(g25271) );
  NAND2X0 U14961 ( .IN1(n14778), .IN2(n14701), .QN(n14777) );
  NAND2X0 U14962 ( .IN1(n14779), .IN2(g2116), .QN(n14776) );
  NAND2X0 U14963 ( .IN1(n14780), .IN2(n14781), .QN(g25270) );
  NAND2X0 U14964 ( .IN1(n14782), .IN2(g1420), .QN(n14781) );
  NAND2X0 U14965 ( .IN1(n14783), .IN2(n14784), .QN(n14780) );
  NAND2X0 U14966 ( .IN1(n14785), .IN2(n14786), .QN(g25268) );
  NAND2X0 U14967 ( .IN1(n10652), .IN2(g2115), .QN(n14786) );
  NAND2X0 U14968 ( .IN1(n14787), .IN2(n14701), .QN(n14785) );
  INVX0 U14969 ( .INP(n14788), .ZN(n14701) );
  NAND2X0 U14970 ( .IN1(n14789), .IN2(n14790), .QN(n14788) );
  NOR2X0 U14971 ( .IN1(n14791), .IN2(n14792), .QN(n14790) );
  NAND2X0 U14972 ( .IN1(n14793), .IN2(n14794), .QN(n14792) );
  NAND2X0 U14973 ( .IN1(n14795), .IN2(n14796), .QN(n14794) );
  NOR2X0 U14974 ( .IN1(n14797), .IN2(n14798), .QN(n14796) );
  NAND2X0 U14975 ( .IN1(n14799), .IN2(n14800), .QN(n14798) );
  XNOR2X1 U14976 ( .IN1(n10282), .IN2(n4400), .Q(n14800) );
  INVX0 U14977 ( .INP(n10283), .ZN(n10282) );
  NAND2X0 U14978 ( .IN1(n14801), .IN2(n14802), .QN(n10283) );
  NAND2X0 U14979 ( .IN1(n9076), .IN2(g7357), .QN(n14802) );
  NOR2X0 U14980 ( .IN1(n14803), .IN2(n14804), .QN(n14801) );
  NOR2X0 U14981 ( .IN1(n4307), .IN2(g2079), .QN(n14804) );
  NOR2X0 U14982 ( .IN1(n4293), .IN2(g2078), .QN(n14803) );
  XNOR2X1 U14983 ( .IN1(n10255), .IN2(n4410), .Q(n14799) );
  INVX0 U14984 ( .INP(n10256), .ZN(n10255) );
  NAND2X0 U14985 ( .IN1(n14805), .IN2(n14806), .QN(n10256) );
  NAND2X0 U14986 ( .IN1(n9070), .IN2(g7357), .QN(n14806) );
  NOR2X0 U14987 ( .IN1(n14807), .IN2(n14808), .QN(n14805) );
  NOR2X0 U14988 ( .IN1(n4307), .IN2(g2088), .QN(n14808) );
  NOR2X0 U14989 ( .IN1(n4293), .IN2(g2087), .QN(n14807) );
  NAND2X0 U14990 ( .IN1(n14809), .IN2(n14810), .QN(n14797) );
  XOR2X1 U14991 ( .IN1(n10230), .IN2(n4416), .Q(n14810) );
  NAND2X0 U14992 ( .IN1(n14811), .IN2(n14812), .QN(n10230) );
  NAND2X0 U14993 ( .IN1(g7357), .IN2(n9290), .QN(n14812) );
  NOR2X0 U14994 ( .IN1(n14813), .IN2(n14814), .QN(n14811) );
  NOR2X0 U14995 ( .IN1(n4307), .IN2(g2106), .QN(n14814) );
  NOR2X0 U14996 ( .IN1(n4293), .IN2(g2105), .QN(n14813) );
  NOR2X0 U14997 ( .IN1(n14815), .IN2(n14816), .QN(n14809) );
  XNOR2X1 U14998 ( .IN1(n4409), .IN2(n10289), .Q(n14816) );
  NAND2X0 U14999 ( .IN1(n14817), .IN2(n14818), .QN(n10289) );
  NAND2X0 U15000 ( .IN1(n9067), .IN2(g7357), .QN(n14818) );
  NOR2X0 U15001 ( .IN1(n14819), .IN2(n14820), .QN(n14817) );
  NOR2X0 U15002 ( .IN1(n4307), .IN2(g2094), .QN(n14820) );
  NOR2X0 U15003 ( .IN1(n4293), .IN2(g2093), .QN(n14819) );
  XNOR2X1 U15004 ( .IN1(n10235), .IN2(test_so70), .Q(n14815) );
  INVX0 U15005 ( .INP(n10238), .ZN(n10235) );
  NAND2X0 U15006 ( .IN1(n14821), .IN2(n14822), .QN(n10238) );
  NAND2X0 U15007 ( .IN1(n9061), .IN2(g7357), .QN(n14822) );
  NOR2X0 U15008 ( .IN1(n14823), .IN2(n14824), .QN(n14821) );
  NOR2X0 U15009 ( .IN1(n4307), .IN2(g2103), .QN(n14824) );
  NOR2X0 U15010 ( .IN1(n4293), .IN2(g2102), .QN(n14823) );
  NOR2X0 U15011 ( .IN1(n14825), .IN2(n14826), .QN(n14795) );
  NAND2X0 U15012 ( .IN1(n14827), .IN2(n14828), .QN(n14826) );
  XNOR2X1 U15013 ( .IN1(n10296), .IN2(n4420), .Q(n14828) );
  INVX0 U15014 ( .INP(n10297), .ZN(n10296) );
  NAND2X0 U15015 ( .IN1(n14829), .IN2(n14830), .QN(n10297) );
  NAND2X0 U15016 ( .IN1(n9072), .IN2(g7357), .QN(n14830) );
  NOR2X0 U15017 ( .IN1(n14831), .IN2(n14832), .QN(n14829) );
  NOR2X0 U15018 ( .IN1(n4307), .IN2(g2085), .QN(n14832) );
  NOR2X0 U15019 ( .IN1(n4293), .IN2(g2084), .QN(n14831) );
  XNOR2X1 U15020 ( .IN1(n10269), .IN2(n4474), .Q(n14827) );
  INVX0 U15021 ( .INP(n10270), .ZN(n10269) );
  NAND2X0 U15022 ( .IN1(n14833), .IN2(n14834), .QN(n10270) );
  NAND2X0 U15023 ( .IN1(n9074), .IN2(g7357), .QN(n14834) );
  NOR2X0 U15024 ( .IN1(n14835), .IN2(n14836), .QN(n14833) );
  NOR2X0 U15025 ( .IN1(n4307), .IN2(g2082), .QN(n14836) );
  NOR2X0 U15026 ( .IN1(n4293), .IN2(g2081), .QN(n14835) );
  NAND2X0 U15027 ( .IN1(n14837), .IN2(n14838), .QN(n14825) );
  XOR2X1 U15028 ( .IN1(n10251), .IN2(n4399), .Q(n14838) );
  NAND2X0 U15029 ( .IN1(n14839), .IN2(n14840), .QN(n10251) );
  NAND2X0 U15030 ( .IN1(g7357), .IN2(n9291), .QN(n14840) );
  NOR2X0 U15031 ( .IN1(n14841), .IN2(n14842), .QN(n14839) );
  NOR2X0 U15032 ( .IN1(n4307), .IN2(g2091), .QN(n14842) );
  NOR2X0 U15033 ( .IN1(n4293), .IN2(g2090), .QN(n14841) );
  NOR2X0 U15034 ( .IN1(n14843), .IN2(n14844), .QN(n14837) );
  XNOR2X1 U15035 ( .IN1(n4473), .IN2(n10261), .Q(n14844) );
  NAND2X0 U15036 ( .IN1(n14845), .IN2(n14846), .QN(n10261) );
  NAND2X0 U15037 ( .IN1(n9063), .IN2(g7357), .QN(n14846) );
  NOR2X0 U15038 ( .IN1(n14847), .IN2(n14848), .QN(n14845) );
  NOR2X0 U15039 ( .IN1(n4307), .IN2(g2100), .QN(n14848) );
  NOR2X0 U15040 ( .IN1(n4293), .IN2(g2099), .QN(n14847) );
  XNOR2X1 U15041 ( .IN1(n4468), .IN2(n10278), .Q(n14843) );
  NAND2X0 U15042 ( .IN1(n14849), .IN2(n14850), .QN(n10278) );
  NAND2X0 U15043 ( .IN1(n9065), .IN2(g7357), .QN(n14850) );
  NOR2X0 U15044 ( .IN1(n14851), .IN2(n14852), .QN(n14849) );
  NOR2X0 U15045 ( .IN1(n4307), .IN2(g2097), .QN(n14852) );
  NOR2X0 U15046 ( .IN1(n4293), .IN2(g2096), .QN(n14851) );
  NAND2X0 U15047 ( .IN1(n8898), .IN2(g2009), .QN(n14793) );
  NOR2X0 U15048 ( .IN1(n4307), .IN2(g2109), .QN(n14791) );
  NOR2X0 U15049 ( .IN1(n14853), .IN2(n10575), .QN(n14789) );
  NAND2X0 U15050 ( .IN1(n14854), .IN2(n14855), .QN(n10575) );
  NAND2X0 U15051 ( .IN1(n8839), .IN2(g7357), .QN(n14855) );
  NOR2X0 U15052 ( .IN1(n14856), .IN2(n14857), .QN(n14854) );
  NOR2X0 U15053 ( .IN1(n4307), .IN2(g2112), .QN(n14857) );
  NOR2X0 U15054 ( .IN1(n4293), .IN2(g2111), .QN(n14856) );
  NOR2X0 U15055 ( .IN1(n4357), .IN2(g2110), .QN(n14853) );
  NAND2X0 U15056 ( .IN1(n14858), .IN2(n14859), .QN(g25267) );
  NAND2X0 U15057 ( .IN1(n14860), .IN2(g1422), .QN(n14859) );
  NAND2X0 U15058 ( .IN1(n14861), .IN2(n14783), .QN(n14858) );
  NAND2X0 U15059 ( .IN1(n14862), .IN2(n14863), .QN(g25266) );
  NAND2X0 U15060 ( .IN1(n14864), .IN2(g734), .QN(n14863) );
  NAND2X0 U15061 ( .IN1(n14865), .IN2(n14866), .QN(n14862) );
  NAND2X0 U15062 ( .IN1(n14867), .IN2(n14868), .QN(g25265) );
  NAND2X0 U15063 ( .IN1(n14097), .IN2(n9931), .QN(n14868) );
  NAND2X0 U15064 ( .IN1(n14869), .IN2(n14577), .QN(n14867) );
  XOR2X1 U15065 ( .IN1(n9261), .IN2(n9260), .Q(n14869) );
  NAND2X0 U15066 ( .IN1(n14870), .IN2(n14871), .QN(g25263) );
  NAND2X0 U15067 ( .IN1(n9671), .IN2(g1421), .QN(n14871) );
  NAND2X0 U15068 ( .IN1(n14872), .IN2(n14783), .QN(n14870) );
  INVX0 U15069 ( .INP(n14873), .ZN(n14783) );
  NAND2X0 U15070 ( .IN1(n14874), .IN2(n14875), .QN(n14873) );
  NOR2X0 U15071 ( .IN1(n14876), .IN2(n14877), .QN(n14875) );
  NAND2X0 U15072 ( .IN1(n14878), .IN2(n14879), .QN(n14877) );
  NAND2X0 U15073 ( .IN1(n14880), .IN2(n14881), .QN(n14879) );
  NOR2X0 U15074 ( .IN1(n14882), .IN2(n14883), .QN(n14881) );
  NAND2X0 U15075 ( .IN1(n14884), .IN2(n14885), .QN(n14883) );
  XNOR2X1 U15076 ( .IN1(n10425), .IN2(n4402), .Q(n14885) );
  INVX0 U15077 ( .INP(n10426), .ZN(n10425) );
  NAND2X0 U15078 ( .IN1(n14886), .IN2(n14887), .QN(n10426) );
  NAND2X0 U15079 ( .IN1(n9095), .IN2(g7161), .QN(n14887) );
  NOR2X0 U15080 ( .IN1(n14888), .IN2(n14889), .QN(n14886) );
  NOR2X0 U15081 ( .IN1(test_so49), .IN2(n4308), .QN(n14889) );
  NOR2X0 U15082 ( .IN1(n4294), .IN2(g1384), .QN(n14888) );
  XNOR2X1 U15083 ( .IN1(n10398), .IN2(n4412), .Q(n14884) );
  INVX0 U15084 ( .INP(n10399), .ZN(n10398) );
  NAND2X0 U15085 ( .IN1(n14890), .IN2(n14891), .QN(n10399) );
  NAND2X0 U15086 ( .IN1(n9089), .IN2(g7161), .QN(n14891) );
  NOR2X0 U15087 ( .IN1(n14892), .IN2(n14893), .QN(n14890) );
  NOR2X0 U15088 ( .IN1(n4308), .IN2(g1394), .QN(n14893) );
  NOR2X0 U15089 ( .IN1(n4294), .IN2(g1393), .QN(n14892) );
  NAND2X0 U15090 ( .IN1(n14894), .IN2(n14895), .QN(n14882) );
  XNOR2X1 U15091 ( .IN1(n10378), .IN2(n4395), .Q(n14895) );
  INVX0 U15092 ( .INP(n10381), .ZN(n10378) );
  NAND2X0 U15093 ( .IN1(n14896), .IN2(n14897), .QN(n10381) );
  NAND2X0 U15094 ( .IN1(n9080), .IN2(g7161), .QN(n14897) );
  NOR2X0 U15095 ( .IN1(n14898), .IN2(n14899), .QN(n14896) );
  NOR2X0 U15096 ( .IN1(n4308), .IN2(g1409), .QN(n14899) );
  NOR2X0 U15097 ( .IN1(n4294), .IN2(g1408), .QN(n14898) );
  NOR2X0 U15098 ( .IN1(n14900), .IN2(n14901), .QN(n14894) );
  XNOR2X1 U15099 ( .IN1(n4417), .IN2(n10373), .Q(n14901) );
  NAND2X0 U15100 ( .IN1(n14902), .IN2(n14903), .QN(n10373) );
  NAND2X0 U15101 ( .IN1(n9078), .IN2(g7161), .QN(n14903) );
  NOR2X0 U15102 ( .IN1(n14904), .IN2(n14905), .QN(n14902) );
  NOR2X0 U15103 ( .IN1(n4308), .IN2(g1412), .QN(n14905) );
  NOR2X0 U15104 ( .IN1(n4294), .IN2(g1411), .QN(n14904) );
  XNOR2X1 U15105 ( .IN1(n4411), .IN2(n10432), .Q(n14900) );
  INVX0 U15106 ( .INP(n10430), .ZN(n10432) );
  NOR2X0 U15107 ( .IN1(n14906), .IN2(n14907), .QN(n10430) );
  NOR2X0 U15108 ( .IN1(n4358), .IN2(test_so50), .QN(n14907) );
  INVX0 U15109 ( .INP(n14908), .ZN(n14906) );
  NOR2X0 U15110 ( .IN1(n14909), .IN2(n14910), .QN(n14908) );
  NOR2X0 U15111 ( .IN1(n4308), .IN2(g1400), .QN(n14910) );
  NOR2X0 U15112 ( .IN1(n4294), .IN2(g1399), .QN(n14909) );
  NOR2X0 U15113 ( .IN1(n14911), .IN2(n14912), .QN(n14880) );
  NAND2X0 U15114 ( .IN1(n14913), .IN2(n14914), .QN(n14912) );
  XNOR2X1 U15115 ( .IN1(n10439), .IN2(n4421), .Q(n14914) );
  INVX0 U15116 ( .INP(n10440), .ZN(n10439) );
  NAND2X0 U15117 ( .IN1(n14915), .IN2(n14916), .QN(n10440) );
  NAND2X0 U15118 ( .IN1(n9091), .IN2(g7161), .QN(n14916) );
  NOR2X0 U15119 ( .IN1(n14917), .IN2(n14918), .QN(n14915) );
  NOR2X0 U15120 ( .IN1(n4308), .IN2(g1391), .QN(n14918) );
  NOR2X0 U15121 ( .IN1(n4294), .IN2(g1390), .QN(n14917) );
  XNOR2X1 U15122 ( .IN1(n10412), .IN2(n4476), .Q(n14913) );
  INVX0 U15123 ( .INP(n10413), .ZN(n10412) );
  NAND2X0 U15124 ( .IN1(n14919), .IN2(n14920), .QN(n10413) );
  NAND2X0 U15125 ( .IN1(n9093), .IN2(g7161), .QN(n14920) );
  NOR2X0 U15126 ( .IN1(n14921), .IN2(n14922), .QN(n14919) );
  NOR2X0 U15127 ( .IN1(n4308), .IN2(g1388), .QN(n14922) );
  NOR2X0 U15128 ( .IN1(n4294), .IN2(g1387), .QN(n14921) );
  NAND2X0 U15129 ( .IN1(n14923), .IN2(n14924), .QN(n14911) );
  XNOR2X1 U15130 ( .IN1(n10393), .IN2(n4401), .Q(n14924) );
  INVX0 U15131 ( .INP(n10394), .ZN(n10393) );
  NAND2X0 U15132 ( .IN1(n14925), .IN2(n14926), .QN(n10394) );
  NAND2X0 U15133 ( .IN1(n9087), .IN2(g7161), .QN(n14926) );
  NOR2X0 U15134 ( .IN1(n14927), .IN2(n14928), .QN(n14925) );
  NOR2X0 U15135 ( .IN1(n4308), .IN2(g1397), .QN(n14928) );
  NOR2X0 U15136 ( .IN1(n4294), .IN2(g1396), .QN(n14927) );
  NOR2X0 U15137 ( .IN1(n14929), .IN2(n14930), .QN(n14923) );
  XNOR2X1 U15138 ( .IN1(n4475), .IN2(n10404), .Q(n14930) );
  NAND2X0 U15139 ( .IN1(n14931), .IN2(n14932), .QN(n10404) );
  NAND2X0 U15140 ( .IN1(n9082), .IN2(g7161), .QN(n14932) );
  NOR2X0 U15141 ( .IN1(n14933), .IN2(n14934), .QN(n14931) );
  NOR2X0 U15142 ( .IN1(n4308), .IN2(g1406), .QN(n14934) );
  NOR2X0 U15143 ( .IN1(n4294), .IN2(g1405), .QN(n14933) );
  XNOR2X1 U15144 ( .IN1(n4469), .IN2(n10421), .Q(n14929) );
  NAND2X0 U15145 ( .IN1(n14935), .IN2(n14936), .QN(n10421) );
  NAND2X0 U15146 ( .IN1(n9084), .IN2(g7161), .QN(n14936) );
  NOR2X0 U15147 ( .IN1(n14937), .IN2(n14938), .QN(n14935) );
  NOR2X0 U15148 ( .IN1(n4308), .IN2(g1403), .QN(n14938) );
  NOR2X0 U15149 ( .IN1(n4294), .IN2(g1402), .QN(n14937) );
  INVX0 U15150 ( .INP(n14939), .ZN(n14878) );
  NOR2X0 U15151 ( .IN1(n4294), .IN2(test_so51), .QN(n14939) );
  NOR2X0 U15152 ( .IN1(n4308), .IN2(g1415), .QN(n14876) );
  NOR2X0 U15153 ( .IN1(n14940), .IN2(n10600), .QN(n14874) );
  NAND2X0 U15154 ( .IN1(n14941), .IN2(n14942), .QN(n10600) );
  NAND2X0 U15155 ( .IN1(n8841), .IN2(g7161), .QN(n14942) );
  NOR2X0 U15156 ( .IN1(n14943), .IN2(n14944), .QN(n14941) );
  NOR2X0 U15157 ( .IN1(n4308), .IN2(g1418), .QN(n14944) );
  NOR2X0 U15158 ( .IN1(n4294), .IN2(g1417), .QN(n14943) );
  NOR2X0 U15159 ( .IN1(n4358), .IN2(g1416), .QN(n14940) );
  NAND2X0 U15160 ( .IN1(n14945), .IN2(n14946), .QN(g25262) );
  NAND2X0 U15161 ( .IN1(n14947), .IN2(g736), .QN(n14946) );
  NAND2X0 U15162 ( .IN1(n14948), .IN2(n14865), .QN(n14945) );
  NAND2X0 U15163 ( .IN1(n14949), .IN2(n14950), .QN(g25260) );
  NAND2X0 U15164 ( .IN1(n9693), .IN2(g735), .QN(n14950) );
  NAND2X0 U15165 ( .IN1(n14951), .IN2(n14865), .QN(n14949) );
  INVX0 U15166 ( .INP(n14952), .ZN(n14865) );
  NAND2X0 U15167 ( .IN1(n14953), .IN2(n14954), .QN(n14952) );
  NOR2X0 U15168 ( .IN1(n14955), .IN2(n14956), .QN(n14954) );
  NAND2X0 U15169 ( .IN1(n14957), .IN2(n14958), .QN(n14956) );
  NAND2X0 U15170 ( .IN1(n14959), .IN2(n14960), .QN(n14958) );
  NOR2X0 U15171 ( .IN1(n14961), .IN2(n14962), .QN(n14960) );
  NAND2X0 U15172 ( .IN1(n14963), .IN2(n14964), .QN(n14962) );
  XNOR2X1 U15173 ( .IN1(n9950), .IN2(n4414), .Q(n14964) );
  INVX0 U15174 ( .INP(n9953), .ZN(n9950) );
  NAND2X0 U15175 ( .IN1(n14965), .IN2(n14966), .QN(n9953) );
  NAND2X0 U15176 ( .IN1(n9106), .IN2(g6911), .QN(n14966) );
  NOR2X0 U15177 ( .IN1(n14967), .IN2(n14968), .QN(n14965) );
  NOR2X0 U15178 ( .IN1(n4309), .IN2(g708), .QN(n14968) );
  NOR2X0 U15179 ( .IN1(n4295), .IN2(g707), .QN(n14967) );
  XNOR2X1 U15180 ( .IN1(n9965), .IN2(n4413), .Q(n14963) );
  INVX0 U15181 ( .INP(n9966), .ZN(n9965) );
  NAND2X0 U15182 ( .IN1(n14969), .IN2(n14970), .QN(n9966) );
  NAND2X0 U15183 ( .IN1(n9103), .IN2(g6911), .QN(n14970) );
  NOR2X0 U15184 ( .IN1(n14971), .IN2(n14972), .QN(n14969) );
  NOR2X0 U15185 ( .IN1(n4309), .IN2(g714), .QN(n14972) );
  NOR2X0 U15186 ( .IN1(n4295), .IN2(g713), .QN(n14971) );
  NAND2X0 U15187 ( .IN1(n14973), .IN2(n14974), .QN(n14961) );
  XOR2X1 U15188 ( .IN1(n10006), .IN2(n4418), .Q(n14974) );
  NAND2X0 U15189 ( .IN1(n14975), .IN2(n14976), .QN(n10006) );
  NAND2X0 U15190 ( .IN1(g6911), .IN2(n9292), .QN(n14976) );
  NOR2X0 U15191 ( .IN1(n14977), .IN2(n14978), .QN(n14975) );
  NOR2X0 U15192 ( .IN1(n4309), .IN2(g726), .QN(n14978) );
  NOR2X0 U15193 ( .IN1(n4295), .IN2(g725), .QN(n14977) );
  NOR2X0 U15194 ( .IN1(n14979), .IN2(n14980), .QN(n14973) );
  XNOR2X1 U15195 ( .IN1(n4396), .IN2(n10014), .Q(n14980) );
  NAND2X0 U15196 ( .IN1(n14981), .IN2(n14982), .QN(n10014) );
  NAND2X0 U15197 ( .IN1(n9097), .IN2(g6911), .QN(n14982) );
  NOR2X0 U15198 ( .IN1(n14983), .IN2(n14984), .QN(n14981) );
  NOR2X0 U15199 ( .IN1(n4309), .IN2(g723), .QN(n14984) );
  NOR2X0 U15200 ( .IN1(n4295), .IN2(g722), .QN(n14983) );
  XNOR2X1 U15201 ( .IN1(n9970), .IN2(test_so28), .Q(n14979) );
  INVX0 U15202 ( .INP(n9971), .ZN(n9970) );
  NAND2X0 U15203 ( .IN1(n14985), .IN2(n14986), .QN(n9971) );
  NAND2X0 U15204 ( .IN1(n9101), .IN2(g6911), .QN(n14986) );
  NOR2X0 U15205 ( .IN1(n14987), .IN2(n14988), .QN(n14985) );
  NOR2X0 U15206 ( .IN1(n4309), .IN2(g717), .QN(n14988) );
  NOR2X0 U15207 ( .IN1(n4295), .IN2(g716), .QN(n14987) );
  NOR2X0 U15208 ( .IN1(n14989), .IN2(n14990), .QN(n14959) );
  NAND2X0 U15209 ( .IN1(n14991), .IN2(n14992), .QN(n14990) );
  XNOR2X1 U15210 ( .IN1(n9993), .IN2(n4422), .Q(n14992) );
  INVX0 U15211 ( .INP(n9994), .ZN(n9993) );
  NAND2X0 U15212 ( .IN1(n14993), .IN2(n14994), .QN(n9994) );
  NAND2X0 U15213 ( .IN1(n9108), .IN2(g6911), .QN(n14994) );
  NOR2X0 U15214 ( .IN1(n14995), .IN2(n14996), .QN(n14993) );
  NOR2X0 U15215 ( .IN1(n4309), .IN2(g705), .QN(n14996) );
  NOR2X0 U15216 ( .IN1(n4295), .IN2(g704), .QN(n14995) );
  XNOR2X1 U15217 ( .IN1(n9987), .IN2(n4478), .Q(n14991) );
  INVX0 U15218 ( .INP(n9988), .ZN(n9987) );
  NAND2X0 U15219 ( .IN1(n14997), .IN2(n14998), .QN(n9988) );
  NAND2X0 U15220 ( .IN1(n9110), .IN2(g6911), .QN(n14998) );
  NOR2X0 U15221 ( .IN1(n14999), .IN2(n15000), .QN(n14997) );
  NOR2X0 U15222 ( .IN1(n4309), .IN2(g702), .QN(n15000) );
  NOR2X0 U15223 ( .IN1(n4295), .IN2(g701), .QN(n14999) );
  NAND2X0 U15224 ( .IN1(n15001), .IN2(n15002), .QN(n14989) );
  XNOR2X1 U15225 ( .IN1(n9977), .IN2(n4477), .Q(n15002) );
  INVX0 U15226 ( .INP(n9978), .ZN(n9977) );
  NAND2X0 U15227 ( .IN1(n15003), .IN2(n15004), .QN(n9978) );
  NAND2X0 U15228 ( .IN1(n9099), .IN2(g6911), .QN(n15004) );
  NOR2X0 U15229 ( .IN1(n15005), .IN2(n15006), .QN(n15003) );
  NOR2X0 U15230 ( .IN1(n4309), .IN2(g720), .QN(n15006) );
  NOR2X0 U15231 ( .IN1(n4295), .IN2(g719), .QN(n15005) );
  NOR2X0 U15232 ( .IN1(n15007), .IN2(n15008), .QN(n15001) );
  XNOR2X1 U15233 ( .IN1(n4404), .IN2(n9983), .Q(n15008) );
  NAND2X0 U15234 ( .IN1(n15009), .IN2(n15010), .QN(n9983) );
  NAND2X0 U15235 ( .IN1(n9112), .IN2(g6911), .QN(n15010) );
  NOR2X0 U15236 ( .IN1(n15011), .IN2(n15012), .QN(n15009) );
  NOR2X0 U15237 ( .IN1(n4309), .IN2(g699), .QN(n15012) );
  NOR2X0 U15238 ( .IN1(n4295), .IN2(g698), .QN(n15011) );
  XNOR2X1 U15239 ( .IN1(n4403), .IN2(n9960), .Q(n15007) );
  NAND2X0 U15240 ( .IN1(n15013), .IN2(n15014), .QN(n9960) );
  NAND2X0 U15241 ( .IN1(n9105), .IN2(g6911), .QN(n15014) );
  NOR2X0 U15242 ( .IN1(n15015), .IN2(n15016), .QN(n15013) );
  NOR2X0 U15243 ( .IN1(test_so29), .IN2(n4309), .QN(n15016) );
  NOR2X0 U15244 ( .IN1(n4295), .IN2(g710), .QN(n15015) );
  NAND2X0 U15245 ( .IN1(n8901), .IN2(g629), .QN(n14957) );
  NOR2X0 U15246 ( .IN1(n4309), .IN2(g729), .QN(n14955) );
  NOR2X0 U15247 ( .IN1(n15017), .IN2(n10544), .QN(n14953) );
  NAND2X0 U15248 ( .IN1(n15018), .IN2(n15019), .QN(n10544) );
  NAND2X0 U15249 ( .IN1(n8843), .IN2(g6911), .QN(n15019) );
  NOR2X0 U15250 ( .IN1(n15020), .IN2(n15021), .QN(n15018) );
  NOR2X0 U15251 ( .IN1(n4309), .IN2(g732), .QN(n15021) );
  NOR2X0 U15252 ( .IN1(n4295), .IN2(g731), .QN(n15020) );
  NOR2X0 U15253 ( .IN1(n4359), .IN2(g730), .QN(n15017) );
  NAND2X0 U15254 ( .IN1(n15022), .IN2(n15023), .QN(g25259) );
  NAND2X0 U15255 ( .IN1(n15024), .IN2(g2253), .QN(n15023) );
  NAND2X0 U15256 ( .IN1(n15025), .IN2(n13971), .QN(n15022) );
  NAND2X0 U15257 ( .IN1(n15026), .IN2(n15027), .QN(g25257) );
  INVX0 U15258 ( .INP(n15028), .ZN(n15027) );
  NOR2X0 U15259 ( .IN1(n15029), .IN2(n8850), .QN(n15028) );
  NAND2X0 U15260 ( .IN1(n15029), .IN2(n13971), .QN(n15026) );
  NAND2X0 U15261 ( .IN1(n15030), .IN2(n15031), .QN(g25256) );
  NAND2X0 U15262 ( .IN1(n15025), .IN2(n4377), .QN(n15031) );
  NAND2X0 U15263 ( .IN1(n15024), .IN2(g2250), .QN(n15030) );
  NAND2X0 U15264 ( .IN1(n15032), .IN2(n15033), .QN(g25255) );
  NAND2X0 U15265 ( .IN1(n15034), .IN2(g1559), .QN(n15033) );
  NAND2X0 U15266 ( .IN1(n15035), .IN2(n14014), .QN(n15032) );
  NAND2X0 U15267 ( .IN1(n15036), .IN2(n15037), .QN(g25253) );
  NAND2X0 U15268 ( .IN1(n15038), .IN2(g2254), .QN(n15037) );
  NAND2X0 U15269 ( .IN1(n15039), .IN2(n13971), .QN(n15036) );
  NAND2X0 U15270 ( .IN1(n15040), .IN2(n15041), .QN(n13971) );
  NOR2X0 U15271 ( .IN1(n15042), .IN2(n15043), .QN(n15041) );
  NAND2X0 U15272 ( .IN1(g2165), .IN2(g2180), .QN(n15043) );
  NAND2X0 U15273 ( .IN1(g2190), .IN2(g2195), .QN(n15042) );
  NOR2X0 U15274 ( .IN1(n15044), .IN2(n15045), .QN(n15040) );
  NAND2X0 U15275 ( .IN1(g2200), .IN2(g2175), .QN(n15045) );
  NAND2X0 U15276 ( .IN1(g2185), .IN2(g2170), .QN(n15044) );
  NAND2X0 U15277 ( .IN1(n15046), .IN2(n15047), .QN(g25252) );
  NAND2X0 U15278 ( .IN1(n15029), .IN2(n4377), .QN(n15047) );
  INVX0 U15279 ( .INP(n15048), .ZN(n15046) );
  NOR2X0 U15280 ( .IN1(n15029), .IN2(n8853), .QN(n15048) );
  NAND2X0 U15281 ( .IN1(n15049), .IN2(n15050), .QN(g25251) );
  NAND2X0 U15282 ( .IN1(n15025), .IN2(n4373), .QN(n15050) );
  NAND2X0 U15283 ( .IN1(n15024), .IN2(g2247), .QN(n15049) );
  NAND2X0 U15284 ( .IN1(n15051), .IN2(n15052), .QN(g25250) );
  INVX0 U15285 ( .INP(n15053), .ZN(n15052) );
  NOR2X0 U15286 ( .IN1(n15054), .IN2(n8862), .QN(n15053) );
  NAND2X0 U15287 ( .IN1(n15054), .IN2(n14014), .QN(n15051) );
  NAND2X0 U15288 ( .IN1(n15055), .IN2(n15056), .QN(g25249) );
  NAND2X0 U15289 ( .IN1(n15035), .IN2(n4378), .QN(n15056) );
  NAND2X0 U15290 ( .IN1(n15034), .IN2(g1556), .QN(n15055) );
  NAND2X0 U15291 ( .IN1(n15057), .IN2(n15058), .QN(g25248) );
  INVX0 U15292 ( .INP(n15059), .ZN(n15058) );
  NOR2X0 U15293 ( .IN1(n15060), .IN2(n8872), .QN(n15059) );
  NAND2X0 U15294 ( .IN1(n15060), .IN2(n14054), .QN(n15057) );
  NAND2X0 U15295 ( .IN1(n15061), .IN2(n15062), .QN(g25247) );
  NAND2X0 U15296 ( .IN1(n15039), .IN2(n4377), .QN(n15062) );
  NAND2X0 U15297 ( .IN1(n15038), .IN2(g2251), .QN(n15061) );
  NAND2X0 U15298 ( .IN1(n15063), .IN2(n15064), .QN(g25246) );
  NAND2X0 U15299 ( .IN1(n15029), .IN2(n4373), .QN(n15064) );
  INVX0 U15300 ( .INP(n15065), .ZN(n15063) );
  NOR2X0 U15301 ( .IN1(n15029), .IN2(n8856), .QN(n15065) );
  NAND2X0 U15302 ( .IN1(n15066), .IN2(n15067), .QN(g25245) );
  NAND2X0 U15303 ( .IN1(n15024), .IN2(g2244), .QN(n15067) );
  INVX0 U15304 ( .INP(n15025), .ZN(n15024) );
  NAND2X0 U15305 ( .IN1(n15068), .IN2(n15025), .QN(n15066) );
  NOR2X0 U15306 ( .IN1(n10620), .IN2(n4367), .QN(n15025) );
  NAND2X0 U15307 ( .IN1(n15069), .IN2(n15070), .QN(g25244) );
  NAND2X0 U15308 ( .IN1(n15071), .IN2(g1560), .QN(n15070) );
  NAND2X0 U15309 ( .IN1(n15072), .IN2(n14014), .QN(n15069) );
  NAND2X0 U15310 ( .IN1(n15073), .IN2(n15074), .QN(n14014) );
  NOR2X0 U15311 ( .IN1(n15075), .IN2(n15076), .QN(n15074) );
  NAND2X0 U15312 ( .IN1(g1471), .IN2(g1486), .QN(n15076) );
  NAND2X0 U15313 ( .IN1(g1496), .IN2(g1501), .QN(n15075) );
  NOR2X0 U15314 ( .IN1(n15077), .IN2(n15078), .QN(n15073) );
  NAND2X0 U15315 ( .IN1(g1506), .IN2(g1481), .QN(n15078) );
  NAND2X0 U15316 ( .IN1(g1491), .IN2(g1476), .QN(n15077) );
  NAND2X0 U15317 ( .IN1(n15079), .IN2(n15080), .QN(g25243) );
  NAND2X0 U15318 ( .IN1(n15054), .IN2(n4378), .QN(n15080) );
  INVX0 U15319 ( .INP(n15081), .ZN(n15079) );
  NOR2X0 U15320 ( .IN1(n15054), .IN2(n8865), .QN(n15081) );
  NAND2X0 U15321 ( .IN1(n15082), .IN2(n15083), .QN(g25242) );
  NAND2X0 U15322 ( .IN1(test_so54), .IN2(n15034), .QN(n15083) );
  NAND2X0 U15323 ( .IN1(n15035), .IN2(n4374), .QN(n15082) );
  NAND2X0 U15324 ( .IN1(n15084), .IN2(n15085), .QN(g25241) );
  NAND2X0 U15325 ( .IN1(n15086), .IN2(g867), .QN(n15085) );
  NAND2X0 U15326 ( .IN1(n15087), .IN2(n14054), .QN(n15084) );
  NAND2X0 U15327 ( .IN1(n15088), .IN2(n15089), .QN(g25240) );
  NAND2X0 U15328 ( .IN1(n4379), .IN2(n15060), .QN(n15089) );
  INVX0 U15329 ( .INP(n15090), .ZN(n15088) );
  NOR2X0 U15330 ( .IN1(n15060), .IN2(n8875), .QN(n15090) );
  NAND2X0 U15331 ( .IN1(n15091), .IN2(n15092), .QN(g25239) );
  NAND2X0 U15332 ( .IN1(n15093), .IN2(g177), .QN(n15092) );
  NAND2X0 U15333 ( .IN1(n15094), .IN2(n15095), .QN(n15091) );
  NAND2X0 U15334 ( .IN1(n15096), .IN2(n15097), .QN(g25237) );
  NAND2X0 U15335 ( .IN1(n15039), .IN2(n4373), .QN(n15097) );
  NAND2X0 U15336 ( .IN1(n15038), .IN2(g2248), .QN(n15096) );
  NAND2X0 U15337 ( .IN1(n15098), .IN2(n15099), .QN(g25236) );
  INVX0 U15338 ( .INP(n15100), .ZN(n15099) );
  NOR2X0 U15339 ( .IN1(n15029), .IN2(n8859), .QN(n15100) );
  NAND2X0 U15340 ( .IN1(n15068), .IN2(n15029), .QN(n15098) );
  NOR2X0 U15341 ( .IN1(n10620), .IN2(n9278), .QN(n15029) );
  NAND2X0 U15342 ( .IN1(n15101), .IN2(n15102), .QN(g25235) );
  NAND2X0 U15343 ( .IN1(n15072), .IN2(n4378), .QN(n15102) );
  NAND2X0 U15344 ( .IN1(n15071), .IN2(g1557), .QN(n15101) );
  NAND2X0 U15345 ( .IN1(n15103), .IN2(n15104), .QN(g25234) );
  NAND2X0 U15346 ( .IN1(n15054), .IN2(n4374), .QN(n15104) );
  INVX0 U15347 ( .INP(n15105), .ZN(n15103) );
  NOR2X0 U15348 ( .IN1(n15054), .IN2(n8867), .QN(n15105) );
  NAND2X0 U15349 ( .IN1(n15106), .IN2(n15107), .QN(g25233) );
  NAND2X0 U15350 ( .IN1(n15034), .IN2(g1550), .QN(n15107) );
  INVX0 U15351 ( .INP(n15035), .ZN(n15034) );
  NAND2X0 U15352 ( .IN1(n15108), .IN2(n15035), .QN(n15106) );
  NOR2X0 U15353 ( .IN1(n10620), .IN2(n4368), .QN(n15035) );
  NAND2X0 U15354 ( .IN1(n15109), .IN2(n15110), .QN(g25232) );
  NAND2X0 U15355 ( .IN1(n15111), .IN2(g866), .QN(n15110) );
  NAND2X0 U15356 ( .IN1(n15112), .IN2(n14054), .QN(n15109) );
  NAND2X0 U15357 ( .IN1(n15113), .IN2(n15114), .QN(n14054) );
  NOR2X0 U15358 ( .IN1(n15115), .IN2(n15116), .QN(n15114) );
  NAND2X0 U15359 ( .IN1(g785), .IN2(g797), .QN(n15116) );
  NAND2X0 U15360 ( .IN1(g805), .IN2(g809), .QN(n15115) );
  NOR2X0 U15361 ( .IN1(n15117), .IN2(n15118), .QN(n15113) );
  NAND2X0 U15362 ( .IN1(g813), .IN2(g793), .QN(n15118) );
  NAND2X0 U15363 ( .IN1(g801), .IN2(g789), .QN(n15117) );
  NAND2X0 U15364 ( .IN1(n15119), .IN2(n15120), .QN(g25231) );
  NAND2X0 U15365 ( .IN1(n4379), .IN2(n15087), .QN(n15120) );
  NAND2X0 U15366 ( .IN1(n15086), .IN2(g864), .QN(n15119) );
  NAND2X0 U15367 ( .IN1(n15121), .IN2(n15122), .QN(g25230) );
  NAND2X0 U15368 ( .IN1(n15060), .IN2(n4375), .QN(n15122) );
  INVX0 U15369 ( .INP(n15123), .ZN(n15121) );
  NOR2X0 U15370 ( .IN1(n15060), .IN2(n8878), .QN(n15123) );
  NAND2X0 U15371 ( .IN1(n15124), .IN2(n15125), .QN(g25229) );
  INVX0 U15372 ( .INP(n15126), .ZN(n15125) );
  NOR2X0 U15373 ( .IN1(n15127), .IN2(n8884), .QN(n15126) );
  NAND2X0 U15374 ( .IN1(n15127), .IN2(n15095), .QN(n15124) );
  NAND2X0 U15375 ( .IN1(n15128), .IN2(n15129), .QN(g25228) );
  NAND2X0 U15376 ( .IN1(n4380), .IN2(n15094), .QN(n15129) );
  NAND2X0 U15377 ( .IN1(n15093), .IN2(g174), .QN(n15128) );
  NAND2X0 U15378 ( .IN1(n15130), .IN2(n15131), .QN(g25227) );
  NAND2X0 U15379 ( .IN1(n15038), .IN2(g2245), .QN(n15131) );
  INVX0 U15380 ( .INP(n15039), .ZN(n15038) );
  NAND2X0 U15381 ( .IN1(n15068), .IN2(n15039), .QN(n15130) );
  NOR2X0 U15382 ( .IN1(n10620), .IN2(n4324), .QN(n15039) );
  INVX0 U15383 ( .INP(n15132), .ZN(n15068) );
  NAND2X0 U15384 ( .IN1(n15133), .IN2(n15134), .QN(n15132) );
  NOR2X0 U15385 ( .IN1(n4325), .IN2(n4287), .QN(n15134) );
  NOR2X0 U15386 ( .IN1(g2190), .IN2(g2195), .QN(n15133) );
  NAND2X0 U15387 ( .IN1(n15135), .IN2(n15136), .QN(g25225) );
  NAND2X0 U15388 ( .IN1(n15072), .IN2(n4374), .QN(n15136) );
  NAND2X0 U15389 ( .IN1(n15071), .IN2(g1554), .QN(n15135) );
  NAND2X0 U15390 ( .IN1(n15137), .IN2(n15138), .QN(g25224) );
  INVX0 U15391 ( .INP(n15139), .ZN(n15138) );
  NOR2X0 U15392 ( .IN1(n15054), .IN2(n8870), .QN(n15139) );
  NAND2X0 U15393 ( .IN1(n15108), .IN2(n15054), .QN(n15137) );
  NOR2X0 U15394 ( .IN1(n10620), .IN2(n4515), .QN(n15054) );
  NAND2X0 U15395 ( .IN1(n15140), .IN2(n15141), .QN(g25223) );
  NAND2X0 U15396 ( .IN1(n15112), .IN2(n4379), .QN(n15141) );
  NAND2X0 U15397 ( .IN1(n15111), .IN2(g863), .QN(n15140) );
  NAND2X0 U15398 ( .IN1(n15142), .IN2(n15143), .QN(g25222) );
  NAND2X0 U15399 ( .IN1(n15087), .IN2(n4375), .QN(n15143) );
  NAND2X0 U15400 ( .IN1(n15086), .IN2(g861), .QN(n15142) );
  NAND2X0 U15401 ( .IN1(n15144), .IN2(n15145), .QN(g25221) );
  INVX0 U15402 ( .INP(n15146), .ZN(n15145) );
  NOR2X0 U15403 ( .IN1(n15060), .IN2(n8881), .QN(n15146) );
  NAND2X0 U15404 ( .IN1(n15147), .IN2(n15060), .QN(n15144) );
  NOR2X0 U15405 ( .IN1(n10620), .IN2(n9279), .QN(n15060) );
  NAND2X0 U15406 ( .IN1(n15148), .IN2(n15149), .QN(g25220) );
  NAND2X0 U15407 ( .IN1(n15150), .IN2(g178), .QN(n15149) );
  NAND2X0 U15408 ( .IN1(n15151), .IN2(n15095), .QN(n15148) );
  INVX0 U15409 ( .INP(n12569), .ZN(n15095) );
  NOR2X0 U15410 ( .IN1(n15152), .IN2(n15153), .QN(n12569) );
  INVX0 U15411 ( .INP(n15154), .ZN(n15153) );
  NOR2X0 U15412 ( .IN1(n15155), .IN2(n15156), .QN(n15154) );
  NAND2X0 U15413 ( .IN1(g97), .IN2(g109), .QN(n15156) );
  NAND2X0 U15414 ( .IN1(g117), .IN2(g121), .QN(n15155) );
  NAND2X0 U15415 ( .IN1(n15157), .IN2(n15158), .QN(n15152) );
  NOR2X0 U15416 ( .IN1(n4290), .IN2(n4322), .QN(n15158) );
  NOR2X0 U15417 ( .IN1(n4328), .IN2(n4376), .QN(n15157) );
  NAND2X0 U15418 ( .IN1(n15159), .IN2(n15160), .QN(g25219) );
  NAND2X0 U15419 ( .IN1(n4380), .IN2(n15127), .QN(n15160) );
  INVX0 U15420 ( .INP(n15161), .ZN(n15159) );
  NOR2X0 U15421 ( .IN1(n15127), .IN2(n8887), .QN(n15161) );
  NAND2X0 U15422 ( .IN1(n15162), .IN2(n15163), .QN(g25218) );
  NAND2X0 U15423 ( .IN1(n15094), .IN2(n4376), .QN(n15163) );
  NAND2X0 U15424 ( .IN1(n15093), .IN2(g171), .QN(n15162) );
  NAND2X0 U15425 ( .IN1(n15164), .IN2(n15165), .QN(g25217) );
  NAND2X0 U15426 ( .IN1(n15071), .IN2(g1551), .QN(n15165) );
  INVX0 U15427 ( .INP(n15072), .ZN(n15071) );
  NAND2X0 U15428 ( .IN1(n15108), .IN2(n15072), .QN(n15164) );
  NOR2X0 U15429 ( .IN1(n10620), .IN2(n4317), .QN(n15072) );
  INVX0 U15430 ( .INP(n15166), .ZN(n15108) );
  NAND2X0 U15431 ( .IN1(n15167), .IN2(n15168), .QN(n15166) );
  NOR2X0 U15432 ( .IN1(n4326), .IN2(n4288), .QN(n15168) );
  NOR2X0 U15433 ( .IN1(g1496), .IN2(g1501), .QN(n15167) );
  NAND2X0 U15434 ( .IN1(n15169), .IN2(n15170), .QN(g25215) );
  NAND2X0 U15435 ( .IN1(n15112), .IN2(n4375), .QN(n15170) );
  NAND2X0 U15436 ( .IN1(n15111), .IN2(g860), .QN(n15169) );
  NAND2X0 U15437 ( .IN1(n15171), .IN2(n15172), .QN(g25214) );
  NAND2X0 U15438 ( .IN1(test_so33), .IN2(n15086), .QN(n15172) );
  INVX0 U15439 ( .INP(n15087), .ZN(n15086) );
  NAND2X0 U15440 ( .IN1(n15147), .IN2(n15087), .QN(n15171) );
  NOR2X0 U15441 ( .IN1(n10620), .IN2(n4312), .QN(n15087) );
  NAND2X0 U15442 ( .IN1(n15173), .IN2(n15174), .QN(g25213) );
  NAND2X0 U15443 ( .IN1(n15151), .IN2(n4380), .QN(n15174) );
  NAND2X0 U15444 ( .IN1(n15150), .IN2(g175), .QN(n15173) );
  NAND2X0 U15445 ( .IN1(n15175), .IN2(n15176), .QN(g25212) );
  NAND2X0 U15446 ( .IN1(n15127), .IN2(n4376), .QN(n15176) );
  INVX0 U15447 ( .INP(n15177), .ZN(n15175) );
  NOR2X0 U15448 ( .IN1(n15127), .IN2(n8890), .QN(n15177) );
  NAND2X0 U15449 ( .IN1(n15178), .IN2(n15179), .QN(g25211) );
  NAND2X0 U15450 ( .IN1(n15093), .IN2(g168), .QN(n15179) );
  INVX0 U15451 ( .INP(n15094), .ZN(n15093) );
  NAND2X0 U15452 ( .IN1(n15180), .IN2(n15094), .QN(n15178) );
  NOR2X0 U15453 ( .IN1(n10620), .IN2(n4369), .QN(n15094) );
  NAND2X0 U15454 ( .IN1(n15181), .IN2(n15182), .QN(g25209) );
  NAND2X0 U15455 ( .IN1(n15111), .IN2(g857), .QN(n15182) );
  INVX0 U15456 ( .INP(n15112), .ZN(n15111) );
  NAND2X0 U15457 ( .IN1(n15147), .IN2(n15112), .QN(n15181) );
  NOR2X0 U15458 ( .IN1(n10620), .IN2(n4323), .QN(n15112) );
  INVX0 U15459 ( .INP(n15183), .ZN(n15147) );
  NAND2X0 U15460 ( .IN1(n15184), .IN2(n15185), .QN(n15183) );
  NOR2X0 U15461 ( .IN1(n4327), .IN2(n4289), .QN(n15185) );
  NOR2X0 U15462 ( .IN1(g805), .IN2(g809), .QN(n15184) );
  NAND2X0 U15463 ( .IN1(n15186), .IN2(n15187), .QN(g25207) );
  NAND2X0 U15464 ( .IN1(n15151), .IN2(n4376), .QN(n15187) );
  NAND2X0 U15465 ( .IN1(n15150), .IN2(g172), .QN(n15186) );
  NAND2X0 U15466 ( .IN1(n15188), .IN2(n15189), .QN(g25206) );
  INVX0 U15467 ( .INP(n15190), .ZN(n15189) );
  NOR2X0 U15468 ( .IN1(n15127), .IN2(n8893), .QN(n15190) );
  NAND2X0 U15469 ( .IN1(n15180), .IN2(n15127), .QN(n15188) );
  NOR2X0 U15470 ( .IN1(n10620), .IN2(n4512), .QN(n15127) );
  NAND2X0 U15471 ( .IN1(n15191), .IN2(n15192), .QN(g25204) );
  NAND2X0 U15472 ( .IN1(n15150), .IN2(g169), .QN(n15192) );
  INVX0 U15473 ( .INP(n15151), .ZN(n15150) );
  NAND2X0 U15474 ( .IN1(n15180), .IN2(n15151), .QN(n15191) );
  NOR2X0 U15475 ( .IN1(n10620), .IN2(n4318), .QN(n15151) );
  NAND2X0 U15476 ( .IN1(n15193), .IN2(n15194), .QN(n10620) );
  NOR2X0 U15477 ( .IN1(n15195), .IN2(n15196), .QN(n15194) );
  NAND2X0 U15478 ( .IN1(n4482), .IN2(n13846), .QN(n15196) );
  INVX0 U15479 ( .INP(n9753), .ZN(n13846) );
  INVX0 U15480 ( .INP(n15197), .ZN(n15195) );
  NOR2X0 U15481 ( .IN1(n4330), .IN2(n4349), .QN(n15197) );
  NOR2X0 U15482 ( .IN1(g2888), .IN2(n15198), .QN(n15193) );
  NAND2X0 U15483 ( .IN1(n8985), .IN2(n4479), .QN(n15198) );
  INVX0 U15484 ( .INP(n15199), .ZN(n15180) );
  NAND2X0 U15485 ( .IN1(n15200), .IN2(n15201), .QN(n15199) );
  NOR2X0 U15486 ( .IN1(n4328), .IN2(n4290), .QN(n15201) );
  NOR2X0 U15487 ( .IN1(g117), .IN2(g121), .QN(n15200) );
  NOR2X0 U15488 ( .IN1(n15202), .IN2(n15203), .QN(g25202) );
  XOR2X1 U15489 ( .IN1(n8695), .IN2(n15204), .Q(n15203) );
  NOR2X0 U15490 ( .IN1(n15205), .IN2(n15206), .QN(g25199) );
  XNOR2X1 U15491 ( .IN1(n8985), .IN2(n15207), .Q(n15206) );
  NOR2X0 U15492 ( .IN1(n10617), .IN2(n15208), .QN(g25197) );
  XNOR2X1 U15493 ( .IN1(n4397), .IN2(n14106), .Q(n15208) );
  NOR2X0 U15494 ( .IN1(n14094), .IN2(n15209), .QN(g25194) );
  XNOR2X1 U15495 ( .IN1(n4399), .IN2(n14123), .Q(n15209) );
  NOR2X0 U15496 ( .IN1(n14097), .IN2(n15210), .QN(g25191) );
  XNOR2X1 U15497 ( .IN1(g3013), .IN2(n4065), .Q(n15210) );
  NOR2X0 U15498 ( .IN1(n14098), .IN2(n15211), .QN(g25189) );
  XOR2X1 U15499 ( .IN1(g1346), .IN2(n14214), .Q(n15211) );
  NOR2X0 U15500 ( .IN1(n9684), .IN2(n15212), .QN(g25185) );
  XNOR2X1 U15501 ( .IN1(n4403), .IN2(n14306), .Q(n15212) );
  NOR2X0 U15502 ( .IN1(n9702), .IN2(n15213), .QN(g25067) );
  XNOR2X1 U15503 ( .IN1(n8972), .IN2(n3888), .Q(n15213) );
  NAND2X0 U15504 ( .IN1(g2241), .IN2(n9753), .QN(n3888) );
  NOR2X0 U15505 ( .IN1(n15214), .IN2(n9753), .QN(n9702) );
  NOR2X0 U15506 ( .IN1(n9710), .IN2(n15215), .QN(g25056) );
  XNOR2X1 U15507 ( .IN1(n8976), .IN2(n3891), .Q(n15215) );
  NAND2X0 U15508 ( .IN1(g1547), .IN2(n9753), .QN(n3891) );
  NOR2X0 U15509 ( .IN1(n15216), .IN2(n9753), .QN(n9710) );
  NOR2X0 U15510 ( .IN1(n11814), .IN2(n15217), .QN(g25042) );
  XNOR2X1 U15511 ( .IN1(n8980), .IN2(n3894), .Q(n15217) );
  NAND2X0 U15512 ( .IN1(test_so31), .IN2(n9753), .QN(n3894) );
  NOR2X0 U15513 ( .IN1(n15218), .IN2(n9753), .QN(n11814) );
  NOR2X0 U15514 ( .IN1(n9719), .IN2(n15219), .QN(g25027) );
  XNOR2X1 U15515 ( .IN1(n8984), .IN2(n3897), .Q(n15219) );
  NAND2X0 U15516 ( .IN1(g165), .IN2(n9753), .QN(n3897) );
  NOR2X0 U15517 ( .IN1(n15220), .IN2(n9753), .QN(n9719) );
  NAND2X0 U15518 ( .IN1(n15221), .IN2(n15222), .QN(n9753) );
  NOR2X0 U15519 ( .IN1(g2903), .IN2(n15223), .QN(n15222) );
  NAND2X0 U15520 ( .IN1(n4431), .IN2(n4291), .QN(n15223) );
  NOR2X0 U15521 ( .IN1(g2908), .IN2(g2892), .QN(n15221) );
  NAND2X0 U15522 ( .IN1(n3700), .IN2(n15224), .QN(g24734) );
  NAND2X0 U15523 ( .IN1(n13293), .IN2(DFF_146_n1), .QN(n15224) );
  NOR2X0 U15524 ( .IN1(n14474), .IN2(n13271), .QN(n13293) );
  INVX0 U15525 ( .INP(n3705), .ZN(n13271) );
  INVX0 U15526 ( .INP(n3940), .ZN(n14474) );
  NAND2X0 U15527 ( .IN1(n15225), .IN2(n15226), .QN(g24557) );
  NAND2X0 U15528 ( .IN1(n10626), .IN2(n10453), .QN(n15226) );
  INVX0 U15529 ( .INP(n15227), .ZN(n15225) );
  NOR2X0 U15530 ( .IN1(g2624), .IN2(n8648), .QN(n15227) );
  NAND2X0 U15531 ( .IN1(n15228), .IN2(n15229), .QN(g24548) );
  INVX0 U15532 ( .INP(n15230), .ZN(n15229) );
  NOR2X0 U15533 ( .IN1(g7390), .IN2(n8649), .QN(n15230) );
  NAND2X0 U15534 ( .IN1(n15231), .IN2(g7390), .QN(n15228) );
  NAND2X0 U15535 ( .IN1(n15232), .IN2(n15233), .QN(g24547) );
  NAND2X0 U15536 ( .IN1(n10626), .IN2(n12695), .QN(n15233) );
  NOR2X0 U15537 ( .IN1(n12628), .IN2(n4299), .QN(n10626) );
  INVX0 U15538 ( .INP(n15234), .ZN(n15232) );
  NOR2X0 U15539 ( .IN1(g2624), .IN2(n8661), .QN(n15234) );
  NAND2X0 U15540 ( .IN1(n15235), .IN2(n15236), .QN(g24545) );
  NAND2X0 U15541 ( .IN1(n10654), .IN2(n12758), .QN(n15236) );
  INVX0 U15542 ( .INP(n15237), .ZN(n15235) );
  NOR2X0 U15543 ( .IN1(g1930), .IN2(n8651), .QN(n15237) );
  NAND2X0 U15544 ( .IN1(n15238), .IN2(n15239), .QN(g24538) );
  NAND2X0 U15545 ( .IN1(n15231), .IN2(g7302), .QN(n15239) );
  NOR2X0 U15546 ( .IN1(n12628), .IN2(n15240), .QN(n15231) );
  INVX0 U15547 ( .INP(n10453), .ZN(n15240) );
  NAND2X0 U15548 ( .IN1(n15241), .IN2(n15242), .QN(n10453) );
  NOR2X0 U15549 ( .IN1(n15243), .IN2(n15244), .QN(n15242) );
  NOR2X0 U15550 ( .IN1(n8648), .IN2(n4299), .QN(n15244) );
  NOR2X0 U15551 ( .IN1(n8647), .IN2(n15245), .QN(n15243) );
  NAND2X0 U15552 ( .IN1(n10647), .IN2(g185), .QN(n15245) );
  NAND2X0 U15553 ( .IN1(n15246), .IN2(n15247), .QN(n10647) );
  NAND2X0 U15554 ( .IN1(g7390), .IN2(g2641), .QN(n15247) );
  NOR2X0 U15555 ( .IN1(n15248), .IN2(n15249), .QN(n15246) );
  NOR2X0 U15556 ( .IN1(n8768), .IN2(n4314), .QN(n15249) );
  NOR2X0 U15557 ( .IN1(n8769), .IN2(n4299), .QN(n15248) );
  NOR2X0 U15558 ( .IN1(n15250), .IN2(n15251), .QN(n15241) );
  NOR2X0 U15559 ( .IN1(n8649), .IN2(n4370), .QN(n15251) );
  NOR2X0 U15560 ( .IN1(n8646), .IN2(n4314), .QN(n15250) );
  INVX0 U15561 ( .INP(n15252), .ZN(n15238) );
  NOR2X0 U15562 ( .IN1(n11699), .IN2(n8646), .QN(n15252) );
  NAND2X0 U15563 ( .IN1(n15253), .IN2(n15254), .QN(g24537) );
  INVX0 U15564 ( .INP(n15255), .ZN(n15254) );
  NOR2X0 U15565 ( .IN1(g7390), .IN2(n8662), .QN(n15255) );
  NAND2X0 U15566 ( .IN1(n15256), .IN2(g7390), .QN(n15253) );
  NAND2X0 U15567 ( .IN1(n15257), .IN2(n15258), .QN(g24535) );
  INVX0 U15568 ( .INP(n15259), .ZN(n15258) );
  NOR2X0 U15569 ( .IN1(g7194), .IN2(n8652), .QN(n15259) );
  NAND2X0 U15570 ( .IN1(n15260), .IN2(g7194), .QN(n15257) );
  NAND2X0 U15571 ( .IN1(n15261), .IN2(n15262), .QN(g24534) );
  NAND2X0 U15572 ( .IN1(n10654), .IN2(n12827), .QN(n15262) );
  NOR2X0 U15573 ( .IN1(n12628), .IN2(n4366), .QN(n10654) );
  INVX0 U15574 ( .INP(n15263), .ZN(n15261) );
  NOR2X0 U15575 ( .IN1(g1930), .IN2(n8664), .QN(n15263) );
  NAND2X0 U15576 ( .IN1(n15264), .IN2(n15265), .QN(g24532) );
  NAND2X0 U15577 ( .IN1(n9673), .IN2(n12886), .QN(n15265) );
  INVX0 U15578 ( .INP(n15266), .ZN(n15264) );
  NOR2X0 U15579 ( .IN1(g1236), .IN2(n8655), .QN(n15266) );
  NAND2X0 U15580 ( .IN1(n15267), .IN2(n15268), .QN(g24527) );
  INVX0 U15581 ( .INP(n15269), .ZN(n15268) );
  NOR2X0 U15582 ( .IN1(n11699), .IN2(n8660), .QN(n15269) );
  NAND2X0 U15583 ( .IN1(n15256), .IN2(n11699), .QN(n15267) );
  NOR2X0 U15584 ( .IN1(n12628), .IN2(n12696), .QN(n15256) );
  INVX0 U15585 ( .INP(n12695), .ZN(n12696) );
  NAND2X0 U15586 ( .IN1(n15270), .IN2(n15271), .QN(n12695) );
  NOR2X0 U15587 ( .IN1(n15272), .IN2(n15273), .QN(n15271) );
  NOR2X0 U15588 ( .IN1(n8660), .IN2(n11700), .QN(n15273) );
  NOR2X0 U15589 ( .IN1(n1457), .IN2(n15274), .QN(n15272) );
  NAND2X0 U15590 ( .IN1(g185), .IN2(g2598), .QN(n15274) );
  INVX0 U15591 ( .INP(n15275), .ZN(n1457) );
  NAND2X0 U15592 ( .IN1(n15276), .IN2(n15277), .QN(n15275) );
  NAND2X0 U15593 ( .IN1(g7390), .IN2(g2645), .QN(n15277) );
  NOR2X0 U15594 ( .IN1(n15278), .IN2(n15279), .QN(n15276) );
  NOR2X0 U15595 ( .IN1(n8771), .IN2(n4299), .QN(n15279) );
  NOR2X0 U15596 ( .IN1(n8770), .IN2(n11700), .QN(n15278) );
  NOR2X0 U15597 ( .IN1(n15280), .IN2(n15281), .QN(n15270) );
  NOR2X0 U15598 ( .IN1(n8662), .IN2(n4370), .QN(n15281) );
  NOR2X0 U15599 ( .IN1(n8661), .IN2(n4299), .QN(n15280) );
  NAND2X0 U15600 ( .IN1(n15282), .IN2(n15283), .QN(g24525) );
  NAND2X0 U15601 ( .IN1(n15260), .IN2(g7052), .QN(n15283) );
  NOR2X0 U15602 ( .IN1(n12628), .IN2(n15284), .QN(n15260) );
  INVX0 U15603 ( .INP(n12758), .ZN(n15284) );
  NAND2X0 U15604 ( .IN1(n15285), .IN2(n15286), .QN(n12758) );
  NOR2X0 U15605 ( .IN1(n15287), .IN2(n15288), .QN(n15286) );
  NOR2X0 U15606 ( .IN1(n8650), .IN2(n4296), .QN(n15288) );
  NOR2X0 U15607 ( .IN1(n1149), .IN2(n15289), .QN(n15287) );
  NAND2X0 U15608 ( .IN1(g185), .IN2(g1922), .QN(n15289) );
  INVX0 U15609 ( .INP(n15290), .ZN(n1149) );
  NAND2X0 U15610 ( .IN1(n15291), .IN2(n15292), .QN(n15290) );
  NAND2X0 U15611 ( .IN1(g1930), .IN2(g1870), .QN(n15292) );
  NOR2X0 U15612 ( .IN1(n15293), .IN2(n15294), .QN(n15291) );
  NOR2X0 U15613 ( .IN1(n16828), .IN2(n4315), .QN(n15294) );
  NOR2X0 U15614 ( .IN1(n8772), .IN2(n4296), .QN(n15293) );
  NOR2X0 U15615 ( .IN1(n15295), .IN2(n15296), .QN(n15285) );
  NOR2X0 U15616 ( .IN1(n8651), .IN2(n4366), .QN(n15296) );
  NOR2X0 U15617 ( .IN1(n8652), .IN2(n4315), .QN(n15295) );
  INVX0 U15618 ( .INP(n15297), .ZN(n15282) );
  NOR2X0 U15619 ( .IN1(n12749), .IN2(n8650), .QN(n15297) );
  NAND2X0 U15620 ( .IN1(n15298), .IN2(n15299), .QN(g24524) );
  INVX0 U15621 ( .INP(n15300), .ZN(n15299) );
  NOR2X0 U15622 ( .IN1(g7194), .IN2(n8665), .QN(n15300) );
  NAND2X0 U15623 ( .IN1(n15301), .IN2(g7194), .QN(n15298) );
  NAND2X0 U15624 ( .IN1(n15302), .IN2(n15303), .QN(g24522) );
  INVX0 U15625 ( .INP(n15304), .ZN(n15303) );
  NOR2X0 U15626 ( .IN1(g6944), .IN2(n8656), .QN(n15304) );
  NAND2X0 U15627 ( .IN1(n15305), .IN2(g6944), .QN(n15302) );
  NAND2X0 U15628 ( .IN1(n15306), .IN2(n15307), .QN(g24521) );
  NAND2X0 U15629 ( .IN1(n9673), .IN2(n12950), .QN(n15307) );
  NOR2X0 U15630 ( .IN1(n12628), .IN2(n4300), .QN(n9673) );
  INVX0 U15631 ( .INP(n15308), .ZN(n15306) );
  NOR2X0 U15632 ( .IN1(g1236), .IN2(n8667), .QN(n15308) );
  NAND2X0 U15633 ( .IN1(n15309), .IN2(n15310), .QN(g24519) );
  NAND2X0 U15634 ( .IN1(n9695), .IN2(n13011), .QN(n15310) );
  INVX0 U15635 ( .INP(n15311), .ZN(n15309) );
  NOR2X0 U15636 ( .IN1(g550), .IN2(n8658), .QN(n15311) );
  NAND2X0 U15637 ( .IN1(n15312), .IN2(n15313), .QN(g24513) );
  INVX0 U15638 ( .INP(n15314), .ZN(n15313) );
  NOR2X0 U15639 ( .IN1(n12749), .IN2(n8663), .QN(n15314) );
  NAND2X0 U15640 ( .IN1(n15301), .IN2(n12749), .QN(n15312) );
  NOR2X0 U15641 ( .IN1(n12628), .IN2(n15315), .QN(n15301) );
  INVX0 U15642 ( .INP(n12827), .ZN(n15315) );
  NAND2X0 U15643 ( .IN1(n15316), .IN2(n15317), .QN(n12827) );
  NOR2X0 U15644 ( .IN1(n15318), .IN2(n15319), .QN(n15317) );
  NOR2X0 U15645 ( .IN1(n8663), .IN2(n15320), .QN(n15319) );
  NOR2X0 U15646 ( .IN1(n1152), .IN2(n15321), .QN(n15318) );
  NAND2X0 U15647 ( .IN1(g185), .IN2(g1904), .QN(n15321) );
  INVX0 U15648 ( .INP(n15322), .ZN(n1152) );
  NAND2X0 U15649 ( .IN1(n15323), .IN2(n15324), .QN(n15322) );
  NAND2X0 U15650 ( .IN1(g1930), .IN2(g1953), .QN(n15324) );
  NOR2X0 U15651 ( .IN1(n15325), .IN2(n15326), .QN(n15323) );
  NOR2X0 U15652 ( .IN1(n16826), .IN2(n4315), .QN(n15326) );
  NOR2X0 U15653 ( .IN1(n8774), .IN2(n15320), .QN(n15325) );
  NOR2X0 U15654 ( .IN1(n15327), .IN2(n15328), .QN(n15316) );
  NOR2X0 U15655 ( .IN1(n8664), .IN2(n4366), .QN(n15328) );
  NOR2X0 U15656 ( .IN1(n8665), .IN2(n4315), .QN(n15327) );
  NAND2X0 U15657 ( .IN1(n15329), .IN2(n15330), .QN(g24511) );
  NAND2X0 U15658 ( .IN1(n15305), .IN2(g6750), .QN(n15330) );
  NOR2X0 U15659 ( .IN1(n12628), .IN2(n15331), .QN(n15305) );
  INVX0 U15660 ( .INP(n12886), .ZN(n15331) );
  NAND2X0 U15661 ( .IN1(n15332), .IN2(n15333), .QN(n12886) );
  NOR2X0 U15662 ( .IN1(n15334), .IN2(n15335), .QN(n15333) );
  NOR2X0 U15663 ( .IN1(n8655), .IN2(n4300), .QN(n15335) );
  NOR2X0 U15664 ( .IN1(n8654), .IN2(n15336), .QN(n15334) );
  NAND2X0 U15665 ( .IN1(n9675), .IN2(g185), .QN(n15336) );
  NAND2X0 U15666 ( .IN1(n15337), .IN2(n15338), .QN(n9675) );
  NAND2X0 U15667 ( .IN1(g6944), .IN2(g1253), .QN(n15338) );
  NOR2X0 U15668 ( .IN1(n15339), .IN2(n15340), .QN(n15337) );
  NOR2X0 U15669 ( .IN1(n8777), .IN2(n4300), .QN(n15340) );
  NOR2X0 U15670 ( .IN1(n8776), .IN2(n13695), .QN(n15339) );
  NOR2X0 U15671 ( .IN1(n15341), .IN2(n15342), .QN(n15332) );
  NOR2X0 U15672 ( .IN1(n8653), .IN2(n4371), .QN(n15342) );
  NOR2X0 U15673 ( .IN1(n8656), .IN2(n4316), .QN(n15341) );
  INVX0 U15674 ( .INP(n15343), .ZN(n15329) );
  NOR2X0 U15675 ( .IN1(n12608), .IN2(n8653), .QN(n15343) );
  NAND2X0 U15676 ( .IN1(n15344), .IN2(n15345), .QN(g24510) );
  INVX0 U15677 ( .INP(n15346), .ZN(n15345) );
  NOR2X0 U15678 ( .IN1(g6944), .IN2(n8668), .QN(n15346) );
  NAND2X0 U15679 ( .IN1(n15347), .IN2(g6944), .QN(n15344) );
  NAND2X0 U15680 ( .IN1(n15348), .IN2(n15349), .QN(g24508) );
  INVX0 U15681 ( .INP(n15350), .ZN(n15349) );
  NOR2X0 U15682 ( .IN1(g6642), .IN2(n8659), .QN(n15350) );
  NAND2X0 U15683 ( .IN1(n15351), .IN2(g6642), .QN(n15348) );
  NAND2X0 U15684 ( .IN1(n15352), .IN2(n15353), .QN(g24507) );
  NAND2X0 U15685 ( .IN1(n9695), .IN2(n13069), .QN(n15353) );
  NOR2X0 U15686 ( .IN1(n12628), .IN2(n4313), .QN(n9695) );
  INVX0 U15687 ( .INP(n15354), .ZN(n15352) );
  NOR2X0 U15688 ( .IN1(g550), .IN2(n8670), .QN(n15354) );
  NAND2X0 U15689 ( .IN1(n15355), .IN2(n15356), .QN(g24501) );
  INVX0 U15690 ( .INP(n15357), .ZN(n15356) );
  NOR2X0 U15691 ( .IN1(n12608), .IN2(n8666), .QN(n15357) );
  NAND2X0 U15692 ( .IN1(n15347), .IN2(n12608), .QN(n15355) );
  NOR2X0 U15693 ( .IN1(n12628), .IN2(n15358), .QN(n15347) );
  INVX0 U15694 ( .INP(n12950), .ZN(n15358) );
  NAND2X0 U15695 ( .IN1(n15359), .IN2(n15360), .QN(n12950) );
  NOR2X0 U15696 ( .IN1(n15361), .IN2(n15362), .QN(n15360) );
  NOR2X0 U15697 ( .IN1(n8666), .IN2(n13695), .QN(n15362) );
  NOR2X0 U15698 ( .IN1(n845), .IN2(n15363), .QN(n15361) );
  NAND2X0 U15699 ( .IN1(g185), .IN2(g1210), .QN(n15363) );
  INVX0 U15700 ( .INP(n15364), .ZN(n845) );
  NAND2X0 U15701 ( .IN1(n15365), .IN2(n15366), .QN(n15364) );
  NAND2X0 U15702 ( .IN1(n12608), .IN2(g1255), .QN(n15366) );
  NOR2X0 U15703 ( .IN1(n15367), .IN2(n15368), .QN(n15365) );
  NOR2X0 U15704 ( .IN1(n16827), .IN2(n4316), .QN(n15368) );
  NOR2X0 U15705 ( .IN1(n8779), .IN2(n4300), .QN(n15367) );
  NOR2X0 U15706 ( .IN1(n15369), .IN2(n15370), .QN(n15359) );
  NOR2X0 U15707 ( .IN1(n8668), .IN2(n4316), .QN(n15370) );
  NOR2X0 U15708 ( .IN1(n8667), .IN2(n4300), .QN(n15369) );
  NAND2X0 U15709 ( .IN1(n15371), .IN2(n15372), .QN(g24499) );
  NAND2X0 U15710 ( .IN1(n15351), .IN2(g6485), .QN(n15372) );
  NOR2X0 U15711 ( .IN1(n12628), .IN2(n15373), .QN(n15351) );
  INVX0 U15712 ( .INP(n13011), .ZN(n15373) );
  NAND2X0 U15713 ( .IN1(n15374), .IN2(n15375), .QN(n13011) );
  NOR2X0 U15714 ( .IN1(n15376), .IN2(n15377), .QN(n15375) );
  NOR2X0 U15715 ( .IN1(n8657), .IN2(n15378), .QN(n15377) );
  NOR2X0 U15716 ( .IN1(n540), .IN2(n15379), .QN(n15376) );
  NAND2X0 U15717 ( .IN1(g185), .IN2(g542), .QN(n15379) );
  INVX0 U15718 ( .INP(n15380), .ZN(n540) );
  NAND2X0 U15719 ( .IN1(n15381), .IN2(n15382), .QN(n15380) );
  NAND2X0 U15720 ( .IN1(g6642), .IN2(g567), .QN(n15382) );
  NOR2X0 U15721 ( .IN1(n15383), .IN2(n15384), .QN(n15381) );
  NOR2X0 U15722 ( .IN1(n8765), .IN2(n4313), .QN(n15384) );
  NOR2X0 U15723 ( .IN1(n8764), .IN2(n4298), .QN(n15383) );
  NOR2X0 U15724 ( .IN1(n15385), .IN2(n15386), .QN(n15374) );
  NOR2X0 U15725 ( .IN1(n8659), .IN2(n4372), .QN(n15386) );
  NOR2X0 U15726 ( .IN1(n8658), .IN2(n4313), .QN(n15385) );
  INVX0 U15727 ( .INP(n15387), .ZN(n15371) );
  NOR2X0 U15728 ( .IN1(n13002), .IN2(n8657), .QN(n15387) );
  NAND2X0 U15729 ( .IN1(n15388), .IN2(n15389), .QN(g24498) );
  INVX0 U15730 ( .INP(n15390), .ZN(n15389) );
  NOR2X0 U15731 ( .IN1(g6642), .IN2(n8671), .QN(n15390) );
  NAND2X0 U15732 ( .IN1(n15391), .IN2(g6642), .QN(n15388) );
  NAND2X0 U15733 ( .IN1(n15392), .IN2(n15393), .QN(g24491) );
  INVX0 U15734 ( .INP(n15394), .ZN(n15393) );
  NOR2X0 U15735 ( .IN1(n13002), .IN2(n8669), .QN(n15394) );
  NAND2X0 U15736 ( .IN1(n15391), .IN2(n13002), .QN(n15392) );
  NOR2X0 U15737 ( .IN1(n12628), .IN2(n15395), .QN(n15391) );
  INVX0 U15738 ( .INP(n13069), .ZN(n15395) );
  NAND2X0 U15739 ( .IN1(n15396), .IN2(n15397), .QN(n13069) );
  NOR2X0 U15740 ( .IN1(n15398), .IN2(n15399), .QN(n15397) );
  NOR2X0 U15741 ( .IN1(n8669), .IN2(n4298), .QN(n15399) );
  NOR2X0 U15742 ( .IN1(n541), .IN2(n15400), .QN(n15398) );
  NAND2X0 U15743 ( .IN1(g185), .IN2(g524), .QN(n15400) );
  INVX0 U15744 ( .INP(n15401), .ZN(n541) );
  NAND2X0 U15745 ( .IN1(n15402), .IN2(n15403), .QN(n15401) );
  NAND2X0 U15746 ( .IN1(g6642), .IN2(g571), .QN(n15403) );
  NOR2X0 U15747 ( .IN1(n15404), .IN2(n15405), .QN(n15402) );
  NOR2X0 U15748 ( .IN1(n8767), .IN2(n4313), .QN(n15405) );
  NOR2X0 U15749 ( .IN1(n8766), .IN2(n15378), .QN(n15404) );
  NOR2X0 U15750 ( .IN1(n15406), .IN2(n15407), .QN(n15396) );
  NOR2X0 U15751 ( .IN1(n8671), .IN2(n4372), .QN(n15407) );
  NOR2X0 U15752 ( .IN1(n8670), .IN2(n4313), .QN(n15406) );
  NOR2X0 U15753 ( .IN1(n15408), .IN2(n15409), .QN(n12628) );
  NAND2X0 U15754 ( .IN1(n15410), .IN2(n15411), .QN(n15409) );
  NOR2X0 U15755 ( .IN1(n4350), .IN2(n4481), .QN(n15411) );
  INVX0 U15756 ( .INP(n15412), .ZN(n15410) );
  NAND2X0 U15757 ( .IN1(n4480), .IN2(n8695), .QN(n15408) );
  NOR2X0 U15758 ( .IN1(n15413), .IN2(n15414), .QN(g24476) );
  NAND2X0 U15759 ( .IN1(n15207), .IN2(n9868), .QN(n15414) );
  NAND2X0 U15760 ( .IN1(n15415), .IN2(n15416), .QN(n15207) );
  NOR2X0 U15761 ( .IN1(n4479), .IN2(n4349), .QN(n15415) );
  NOR2X0 U15762 ( .IN1(n15417), .IN2(g2924), .QN(n15413) );
  NOR2X0 U15763 ( .IN1(n4479), .IN2(n9871), .QN(n15417) );
  NOR2X0 U15764 ( .IN1(n9867), .IN2(n15418), .QN(g24473) );
  XNOR2X1 U15765 ( .IN1(g2892), .IN2(n9689), .Q(n15418) );
  NOR2X0 U15766 ( .IN1(n4123), .IN2(n4431), .QN(n9689) );
  NAND2X0 U15767 ( .IN1(n15419), .IN2(g2888), .QN(n4123) );
  INVX0 U15768 ( .INP(n15420), .ZN(g24446) );
  NAND2X0 U15769 ( .IN1(n9933), .IN2(n15421), .QN(n15420) );
  NOR2X0 U15770 ( .IN1(n15204), .IN2(n4101), .QN(n15421) );
  NOR2X0 U15771 ( .IN1(n4102), .IN2(n4480), .QN(n15204) );
  NAND2X0 U15772 ( .IN1(n15422), .IN2(g3028), .QN(n4102) );
  NOR2X0 U15773 ( .IN1(n14097), .IN2(n15423), .QN(g24445) );
  XNOR2X1 U15774 ( .IN1(n9262), .IN2(n4066), .Q(n15423) );
  NOR2X0 U15775 ( .IN1(n15424), .IN2(n15425), .QN(g24438) );
  NAND2X0 U15776 ( .IN1(n13918), .IN2(n14106), .QN(n15425) );
  INVX0 U15777 ( .INP(n14104), .ZN(n14106) );
  NOR2X0 U15778 ( .IN1(n15426), .IN2(n15427), .QN(n14104) );
  NAND2X0 U15779 ( .IN1(g2727), .IN2(g2720), .QN(n15426) );
  NOR2X0 U15780 ( .IN1(n15428), .IN2(g2720), .QN(n15424) );
  NOR2X0 U15781 ( .IN1(n4419), .IN2(n15427), .QN(n15428) );
  NOR2X0 U15782 ( .IN1(n15429), .IN2(n15430), .QN(g24434) );
  NAND2X0 U15783 ( .IN1(n14123), .IN2(n13126), .QN(n15430) );
  NAND2X0 U15784 ( .IN1(n15431), .IN2(n15432), .QN(n14123) );
  NOR2X0 U15785 ( .IN1(n4420), .IN2(n4410), .QN(n15431) );
  NOR2X0 U15786 ( .IN1(n15433), .IN2(g2026), .QN(n15429) );
  NOR2X0 U15787 ( .IN1(n4420), .IN2(n15434), .QN(n15433) );
  NOR2X0 U15788 ( .IN1(n15435), .IN2(n15436), .QN(g24430) );
  NAND2X0 U15789 ( .IN1(n14214), .IN2(n13134), .QN(n15436) );
  NAND2X0 U15790 ( .IN1(n15437), .IN2(n15438), .QN(n14214) );
  NOR2X0 U15791 ( .IN1(n4421), .IN2(n4412), .QN(n15437) );
  NOR2X0 U15792 ( .IN1(n15439), .IN2(g1332), .QN(n15435) );
  NOR2X0 U15793 ( .IN1(n4421), .IN2(n15440), .QN(n15439) );
  NOR2X0 U15794 ( .IN1(n15441), .IN2(n15442), .QN(g24426) );
  NAND2X0 U15795 ( .IN1(n13251), .IN2(n14306), .QN(n15442) );
  INVX0 U15796 ( .INP(n14304), .ZN(n14306) );
  NOR2X0 U15797 ( .IN1(n15443), .IN2(n15444), .QN(n14304) );
  NAND2X0 U15798 ( .IN1(g653), .IN2(g646), .QN(n15443) );
  NOR2X0 U15799 ( .IN1(n15445), .IN2(g646), .QN(n15441) );
  NOR2X0 U15800 ( .IN1(n4422), .IN2(n15444), .QN(n15445) );
  NAND2X0 U15801 ( .IN1(n15446), .IN2(n15447), .QN(g24250) );
  NAND2X0 U15802 ( .IN1(n4463), .IN2(g2546), .QN(n15447) );
  NAND2X0 U15803 ( .IN1(n11503), .IN2(g2560), .QN(n15446) );
  NAND2X0 U15804 ( .IN1(n15448), .IN2(n15449), .QN(g24243) );
  NAND2X0 U15805 ( .IN1(n4464), .IN2(g1852), .QN(n15449) );
  NAND2X0 U15806 ( .IN1(n11564), .IN2(g1866), .QN(n15448) );
  NAND2X0 U15807 ( .IN1(n15450), .IN2(n15451), .QN(g24238) );
  INVX0 U15808 ( .INP(n15452), .ZN(n15451) );
  NOR2X0 U15809 ( .IN1(g2560), .IN2(n9002), .QN(n15452) );
  NAND2X0 U15810 ( .IN1(n11477), .IN2(g2560), .QN(n15450) );
  NAND2X0 U15811 ( .IN1(n15453), .IN2(n15454), .QN(g24237) );
  NAND2X0 U15812 ( .IN1(n4455), .IN2(g2543), .QN(n15454) );
  NAND2X0 U15813 ( .IN1(n11503), .IN2(g8167), .QN(n15453) );
  NAND2X0 U15814 ( .IN1(n15455), .IN2(n15456), .QN(g24235) );
  NAND2X0 U15815 ( .IN1(n4465), .IN2(g1158), .QN(n15456) );
  NAND2X0 U15816 ( .IN1(n11627), .IN2(g1172), .QN(n15455) );
  NAND2X0 U15817 ( .IN1(n15457), .IN2(n15458), .QN(g24231) );
  INVX0 U15818 ( .INP(n15459), .ZN(n15458) );
  NOR2X0 U15819 ( .IN1(g1866), .IN2(n9011), .QN(n15459) );
  NAND2X0 U15820 ( .IN1(n12107), .IN2(g1866), .QN(n15457) );
  NAND2X0 U15821 ( .IN1(n15460), .IN2(n15461), .QN(g24230) );
  NAND2X0 U15822 ( .IN1(n4457), .IN2(g1849), .QN(n15461) );
  NAND2X0 U15823 ( .IN1(n11564), .IN2(g8082), .QN(n15460) );
  NAND2X0 U15824 ( .IN1(n15462), .IN2(n15463), .QN(g24228) );
  NAND2X0 U15825 ( .IN1(n4466), .IN2(g471), .QN(n15463) );
  NAND2X0 U15826 ( .IN1(n11693), .IN2(g485), .QN(n15462) );
  NAND2X0 U15827 ( .IN1(n15464), .IN2(n15465), .QN(g24226) );
  NAND2X0 U15828 ( .IN1(n4455), .IN2(g2553), .QN(n15465) );
  NAND2X0 U15829 ( .IN1(n11477), .IN2(g8167), .QN(n15464) );
  NAND2X0 U15830 ( .IN1(n15466), .IN2(n15467), .QN(g24225) );
  NAND2X0 U15831 ( .IN1(n4456), .IN2(g2540), .QN(n15467) );
  NAND2X0 U15832 ( .IN1(n11503), .IN2(g8087), .QN(n15466) );
  INVX0 U15833 ( .INP(n9834), .ZN(n11503) );
  NAND2X0 U15834 ( .IN1(n11132), .IN2(n11106), .QN(n9834) );
  NOR2X0 U15835 ( .IN1(n11110), .IN2(n11114), .QN(n11132) );
  NAND2X0 U15836 ( .IN1(n15468), .IN2(n15469), .QN(g24223) );
  INVX0 U15837 ( .INP(n15470), .ZN(n15469) );
  NOR2X0 U15838 ( .IN1(g1172), .IN2(n9019), .QN(n15470) );
  NAND2X0 U15839 ( .IN1(n11601), .IN2(g1172), .QN(n15468) );
  NAND2X0 U15840 ( .IN1(n15471), .IN2(n15472), .QN(g24222) );
  NAND2X0 U15841 ( .IN1(n4459), .IN2(g1155), .QN(n15472) );
  NAND2X0 U15842 ( .IN1(n11627), .IN2(g8007), .QN(n15471) );
  NAND2X0 U15843 ( .IN1(n15473), .IN2(n15474), .QN(g24219) );
  NAND2X0 U15844 ( .IN1(n4457), .IN2(g1859), .QN(n15474) );
  NAND2X0 U15845 ( .IN1(n12107), .IN2(g8082), .QN(n15473) );
  NAND2X0 U15846 ( .IN1(n15475), .IN2(n15476), .QN(g24218) );
  NAND2X0 U15847 ( .IN1(n4458), .IN2(g1846), .QN(n15476) );
  NAND2X0 U15848 ( .IN1(n11564), .IN2(g8012), .QN(n15475) );
  INVX0 U15849 ( .INP(n9799), .ZN(n11564) );
  NAND2X0 U15850 ( .IN1(n10710), .IN2(n10690), .QN(n9799) );
  NOR2X0 U15851 ( .IN1(n10707), .IN2(n10700), .QN(n10710) );
  NAND2X0 U15852 ( .IN1(n15477), .IN2(n15478), .QN(g24216) );
  INVX0 U15853 ( .INP(n15479), .ZN(n15478) );
  NOR2X0 U15854 ( .IN1(g485), .IN2(n9028), .QN(n15479) );
  NAND2X0 U15855 ( .IN1(n12337), .IN2(g485), .QN(n15477) );
  NAND2X0 U15856 ( .IN1(n15480), .IN2(n15481), .QN(g24215) );
  NAND2X0 U15857 ( .IN1(n11693), .IN2(g7956), .QN(n15481) );
  NAND2X0 U15858 ( .IN1(test_so24), .IN2(n4461), .QN(n15480) );
  NAND2X0 U15859 ( .IN1(n15482), .IN2(n15483), .QN(g24214) );
  INVX0 U15860 ( .INP(n15484), .ZN(n15483) );
  NOR2X0 U15861 ( .IN1(g8087), .IN2(n9001), .QN(n15484) );
  NAND2X0 U15862 ( .IN1(n11477), .IN2(g8087), .QN(n15482) );
  INVX0 U15863 ( .INP(n12038), .ZN(n11477) );
  NAND2X0 U15864 ( .IN1(n15485), .IN2(n11102), .QN(n12038) );
  NOR2X0 U15865 ( .IN1(n11123), .IN2(n11106), .QN(n15485) );
  NAND2X0 U15866 ( .IN1(n15486), .IN2(n15487), .QN(g24213) );
  NAND2X0 U15867 ( .IN1(n4459), .IN2(g1165), .QN(n15487) );
  NAND2X0 U15868 ( .IN1(n11601), .IN2(g8007), .QN(n15486) );
  NAND2X0 U15869 ( .IN1(n15488), .IN2(n15489), .QN(g24212) );
  NAND2X0 U15870 ( .IN1(n4460), .IN2(g1152), .QN(n15489) );
  NAND2X0 U15871 ( .IN1(n11627), .IN2(g7961), .QN(n15488) );
  INVX0 U15872 ( .INP(n9764), .ZN(n11627) );
  NAND2X0 U15873 ( .IN1(n15490), .IN2(n10495), .QN(n9764) );
  NOR2X0 U15874 ( .IN1(n10489), .IN2(n10483), .QN(n15490) );
  INVX0 U15875 ( .INP(n10486), .ZN(n10483) );
  NAND2X0 U15876 ( .IN1(n15491), .IN2(n15492), .QN(g24209) );
  NAND2X0 U15877 ( .IN1(n4463), .IN2(g2536), .QN(n15492) );
  NAND2X0 U15878 ( .IN1(n13652), .IN2(g2560), .QN(n15491) );
  NAND2X0 U15879 ( .IN1(n15493), .IN2(n15494), .QN(g24208) );
  INVX0 U15880 ( .INP(n15495), .ZN(n15494) );
  NOR2X0 U15881 ( .IN1(g8012), .IN2(n9010), .QN(n15495) );
  NAND2X0 U15882 ( .IN1(n12107), .IN2(g8012), .QN(n15493) );
  INVX0 U15883 ( .INP(n11784), .ZN(n12107) );
  NAND2X0 U15884 ( .IN1(n15496), .IN2(n10686), .QN(n11784) );
  NOR2X0 U15885 ( .IN1(n11198), .IN2(n10690), .QN(n15496) );
  NAND2X0 U15886 ( .IN1(n15497), .IN2(n15498), .QN(g24207) );
  NAND2X0 U15887 ( .IN1(n4461), .IN2(g478), .QN(n15498) );
  NAND2X0 U15888 ( .IN1(n12337), .IN2(g7956), .QN(n15497) );
  NAND2X0 U15889 ( .IN1(n15499), .IN2(n15500), .QN(g24206) );
  NAND2X0 U15890 ( .IN1(g465), .IN2(n9286), .QN(n15500) );
  NAND2X0 U15891 ( .IN1(test_so23), .IN2(n11693), .QN(n15499) );
  INVX0 U15892 ( .INP(n9729), .ZN(n11693) );
  NAND2X0 U15893 ( .IN1(n10749), .IN2(n10729), .QN(n9729) );
  NOR2X0 U15894 ( .IN1(n10746), .IN2(n10739), .QN(n10749) );
  NAND2X0 U15895 ( .IN1(n15501), .IN2(n15502), .QN(g24182) );
  NAND2X0 U15896 ( .IN1(n4464), .IN2(g1842), .QN(n15502) );
  NAND2X0 U15897 ( .IN1(n13758), .IN2(g1866), .QN(n15501) );
  NAND2X0 U15898 ( .IN1(n15503), .IN2(n15504), .QN(g24181) );
  INVX0 U15899 ( .INP(n15505), .ZN(n15504) );
  NOR2X0 U15900 ( .IN1(g7961), .IN2(n9018), .QN(n15505) );
  NAND2X0 U15901 ( .IN1(n11601), .IN2(g7961), .QN(n15503) );
  INVX0 U15902 ( .INP(n11798), .ZN(n11601) );
  NAND2X0 U15903 ( .IN1(n15506), .IN2(n10495), .QN(n11798) );
  NOR2X0 U15904 ( .IN1(n10507), .IN2(n10486), .QN(n15506) );
  NAND2X0 U15905 ( .IN1(n15507), .IN2(n15508), .QN(g24179) );
  NAND2X0 U15906 ( .IN1(n4465), .IN2(g1148), .QN(n15508) );
  NAND2X0 U15907 ( .IN1(n15509), .IN2(g1172), .QN(n15507) );
  NAND2X0 U15908 ( .IN1(n15510), .IN2(n15511), .QN(g24178) );
  INVX0 U15909 ( .INP(n15512), .ZN(n15511) );
  NOR2X0 U15910 ( .IN1(n9027), .IN2(test_so23), .QN(n15512) );
  NAND2X0 U15911 ( .IN1(test_so23), .IN2(n12337), .QN(n15510) );
  INVX0 U15912 ( .INP(n11809), .ZN(n12337) );
  NAND2X0 U15913 ( .IN1(n15513), .IN2(n10725), .QN(n11809) );
  NOR2X0 U15914 ( .IN1(n11158), .IN2(n10729), .QN(n15513) );
  NAND2X0 U15915 ( .IN1(n15514), .IN2(n15515), .QN(g24174) );
  NAND2X0 U15916 ( .IN1(n4466), .IN2(g461), .QN(n15515) );
  NAND2X0 U15917 ( .IN1(n13889), .IN2(g485), .QN(n15514) );
  NAND2X0 U15918 ( .IN1(n15516), .IN2(n15517), .QN(g24092) );
  NAND2X0 U15919 ( .IN1(g3229), .IN2(n4483), .QN(n15517) );
  NAND2X0 U15920 ( .IN1(n10022), .IN2(g2380), .QN(n15516) );
  INVX0 U15921 ( .INP(g3229), .ZN(n10022) );
  NAND2X0 U15922 ( .IN1(n15518), .IN2(n15519), .QN(g24083) );
  NAND2X0 U15923 ( .IN1(g3229), .IN2(n4484), .QN(n15519) );
  INVX0 U15924 ( .INP(n15520), .ZN(n15518) );
  NOR2X0 U15925 ( .IN1(g3229), .IN2(n8986), .QN(n15520) );
  NAND2X0 U15926 ( .IN1(n15521), .IN2(n15522), .QN(g24072) );
  NAND2X0 U15927 ( .IN1(g3229), .IN2(n4486), .QN(n15522) );
  INVX0 U15928 ( .INP(n15523), .ZN(n15521) );
  NOR2X0 U15929 ( .IN1(g3229), .IN2(n8987), .QN(n15523) );
  NAND2X0 U15930 ( .IN1(n15524), .IN2(n15525), .QN(g24059) );
  NAND2X0 U15931 ( .IN1(g3229), .IN2(n4485), .QN(n15525) );
  INVX0 U15932 ( .INP(n15526), .ZN(n15524) );
  NOR2X0 U15933 ( .IN1(g3229), .IN2(n8699), .QN(n15526) );
  NAND2X0 U15934 ( .IN1(n15527), .IN2(n15528), .QN(g23418) );
  NAND2X0 U15935 ( .IN1(n4455), .IN2(g2533), .QN(n15528) );
  NAND2X0 U15936 ( .IN1(n13652), .IN2(g8167), .QN(n15527) );
  NAND2X0 U15937 ( .IN1(n15529), .IN2(n15530), .QN(g23413) );
  NAND2X0 U15938 ( .IN1(n13758), .IN2(g8082), .QN(n15530) );
  NAND2X0 U15939 ( .IN1(test_so65), .IN2(n4457), .QN(n15529) );
  NAND2X0 U15940 ( .IN1(n15531), .IN2(n15532), .QN(g23407) );
  NAND2X0 U15941 ( .IN1(n4456), .IN2(g2530), .QN(n15532) );
  NAND2X0 U15942 ( .IN1(n13652), .IN2(g8087), .QN(n15531) );
  INVX0 U15943 ( .INP(n9857), .ZN(n13652) );
  NAND2X0 U15944 ( .IN1(n15533), .IN2(n11106), .QN(n9857) );
  INVX0 U15945 ( .INP(n11133), .ZN(n11106) );
  NAND2X0 U15946 ( .IN1(n15534), .IN2(n15535), .QN(n11133) );
  NAND2X0 U15947 ( .IN1(n8495), .IN2(n10669), .QN(n15535) );
  NOR2X0 U15948 ( .IN1(n15536), .IN2(n15537), .QN(n15534) );
  NOR2X0 U15949 ( .IN1(n4516), .IN2(g2387), .QN(n15537) );
  NOR2X0 U15950 ( .IN1(n4509), .IN2(g2389), .QN(n15536) );
  NOR2X0 U15951 ( .IN1(n11102), .IN2(n11123), .QN(n15533) );
  INVX0 U15952 ( .INP(n11114), .ZN(n11123) );
  NAND2X0 U15953 ( .IN1(n15538), .IN2(n15539), .QN(n11114) );
  NAND2X0 U15954 ( .IN1(n8493), .IN2(n10669), .QN(n15539) );
  NOR2X0 U15955 ( .IN1(n15540), .IN2(n15541), .QN(n15538) );
  NOR2X0 U15956 ( .IN1(n4516), .IN2(g2393), .QN(n15541) );
  NOR2X0 U15957 ( .IN1(n4509), .IN2(g2395), .QN(n15540) );
  INVX0 U15958 ( .INP(n11110), .ZN(n11102) );
  NAND2X0 U15959 ( .IN1(n15542), .IN2(n15543), .QN(n11110) );
  NAND2X0 U15960 ( .IN1(n8494), .IN2(n10669), .QN(n15543) );
  INVX0 U15961 ( .INP(n4524), .ZN(n10669) );
  NOR2X0 U15962 ( .IN1(n15544), .IN2(n15545), .QN(n15542) );
  NOR2X0 U15963 ( .IN1(n4516), .IN2(g2390), .QN(n15545) );
  NOR2X0 U15964 ( .IN1(n4509), .IN2(g2392), .QN(n15544) );
  NAND2X0 U15965 ( .IN1(n15546), .IN2(n15547), .QN(g23406) );
  NAND2X0 U15966 ( .IN1(n4459), .IN2(g1145), .QN(n15547) );
  NAND2X0 U15967 ( .IN1(n15509), .IN2(g8007), .QN(n15546) );
  NAND2X0 U15968 ( .IN1(n15548), .IN2(n15549), .QN(g23400) );
  NAND2X0 U15969 ( .IN1(n4458), .IN2(g1836), .QN(n15549) );
  NAND2X0 U15970 ( .IN1(n13758), .IN2(g8012), .QN(n15548) );
  INVX0 U15971 ( .INP(n9822), .ZN(n13758) );
  NAND2X0 U15972 ( .IN1(n15550), .IN2(n10690), .QN(n9822) );
  INVX0 U15973 ( .INP(n10711), .ZN(n10690) );
  NAND2X0 U15974 ( .IN1(n15551), .IN2(n15552), .QN(n10711) );
  NAND2X0 U15975 ( .IN1(n8498), .IN2(n10678), .QN(n15552) );
  NOR2X0 U15976 ( .IN1(n15553), .IN2(n15554), .QN(n15551) );
  NOR2X0 U15977 ( .IN1(n4518), .IN2(g1693), .QN(n15554) );
  NOR2X0 U15978 ( .IN1(n4511), .IN2(g1695), .QN(n15553) );
  NOR2X0 U15979 ( .IN1(n10686), .IN2(n11198), .QN(n15550) );
  INVX0 U15980 ( .INP(n10700), .ZN(n11198) );
  NAND2X0 U15981 ( .IN1(n15555), .IN2(n15556), .QN(n10700) );
  NAND2X0 U15982 ( .IN1(n8496), .IN2(n10678), .QN(n15556) );
  NOR2X0 U15983 ( .IN1(n15557), .IN2(n15558), .QN(n15555) );
  NOR2X0 U15984 ( .IN1(n4518), .IN2(g1699), .QN(n15558) );
  NOR2X0 U15985 ( .IN1(n4511), .IN2(g1701), .QN(n15557) );
  INVX0 U15986 ( .INP(n10707), .ZN(n10686) );
  NAND2X0 U15987 ( .IN1(n15559), .IN2(n15560), .QN(n10707) );
  NAND2X0 U15988 ( .IN1(n8497), .IN2(n10678), .QN(n15560) );
  INVX0 U15989 ( .INP(n4525), .ZN(n10678) );
  NOR2X0 U15990 ( .IN1(n15561), .IN2(n15562), .QN(n15559) );
  NOR2X0 U15991 ( .IN1(n4518), .IN2(g1696), .QN(n15562) );
  NOR2X0 U15992 ( .IN1(n4511), .IN2(g1698), .QN(n15561) );
  NAND2X0 U15993 ( .IN1(n15563), .IN2(n15564), .QN(g23399) );
  NAND2X0 U15994 ( .IN1(n4461), .IN2(g458), .QN(n15564) );
  NAND2X0 U15995 ( .IN1(n13889), .IN2(g7956), .QN(n15563) );
  NAND2X0 U15996 ( .IN1(n15565), .IN2(n15566), .QN(g23392) );
  NAND2X0 U15997 ( .IN1(n4460), .IN2(g1142), .QN(n15566) );
  NAND2X0 U15998 ( .IN1(n15509), .IN2(g7961), .QN(n15565) );
  INVX0 U15999 ( .INP(n9787), .ZN(n15509) );
  NAND2X0 U16000 ( .IN1(n10507), .IN2(n10498), .QN(n9787) );
  NOR2X0 U16001 ( .IN1(n10495), .IN2(n10486), .QN(n10498) );
  NOR2X0 U16002 ( .IN1(n15567), .IN2(n15568), .QN(n10486) );
  NOR2X0 U16003 ( .IN1(n4381), .IN2(test_so39), .QN(n15568) );
  INVX0 U16004 ( .INP(n15569), .ZN(n15567) );
  NOR2X0 U16005 ( .IN1(n15570), .IN2(n15571), .QN(n15569) );
  NOR2X0 U16006 ( .IN1(n4364), .IN2(g1006), .QN(n15571) );
  NOR2X0 U16007 ( .IN1(n4363), .IN2(g1005), .QN(n15570) );
  INVX0 U16008 ( .INP(n10492), .ZN(n10495) );
  NAND2X0 U16009 ( .IN1(n15572), .IN2(n15573), .QN(n10492) );
  NAND2X0 U16010 ( .IN1(n8515), .IN2(g1088), .QN(n15573) );
  NOR2X0 U16011 ( .IN1(n15574), .IN2(n15575), .QN(n15572) );
  NOR2X0 U16012 ( .IN1(n4364), .IN2(g1003), .QN(n15575) );
  NOR2X0 U16013 ( .IN1(n4363), .IN2(g1002), .QN(n15574) );
  INVX0 U16014 ( .INP(n10489), .ZN(n10507) );
  NAND2X0 U16015 ( .IN1(n15576), .IN2(n15577), .QN(n10489) );
  NAND2X0 U16016 ( .IN1(n8517), .IN2(g1088), .QN(n15577) );
  NOR2X0 U16017 ( .IN1(n15578), .IN2(n15579), .QN(n15576) );
  NOR2X0 U16018 ( .IN1(n4364), .IN2(g1000), .QN(n15579) );
  NOR2X0 U16019 ( .IN1(n4363), .IN2(g999), .QN(n15578) );
  NAND2X0 U16020 ( .IN1(n15580), .IN2(n15581), .QN(g23385) );
  NAND2X0 U16021 ( .IN1(g455), .IN2(n9286), .QN(n15581) );
  NAND2X0 U16022 ( .IN1(n13889), .IN2(test_so23), .QN(n15580) );
  INVX0 U16023 ( .INP(n9752), .ZN(n13889) );
  NAND2X0 U16024 ( .IN1(n15582), .IN2(n10729), .QN(n9752) );
  INVX0 U16025 ( .INP(n10750), .ZN(n10729) );
  NAND2X0 U16026 ( .IN1(n15583), .IN2(n15584), .QN(n10750) );
  NAND2X0 U16027 ( .IN1(n8526), .IN2(n10752), .QN(n15584) );
  NOR2X0 U16028 ( .IN1(n15585), .IN2(n15586), .QN(n15583) );
  NOR2X0 U16029 ( .IN1(n4506), .IN2(g314), .QN(n15586) );
  NOR2X0 U16030 ( .IN1(n4499), .IN2(g313), .QN(n15585) );
  NOR2X0 U16031 ( .IN1(n10725), .IN2(n11158), .QN(n15582) );
  INVX0 U16032 ( .INP(n10739), .ZN(n11158) );
  NAND2X0 U16033 ( .IN1(n15587), .IN2(n15588), .QN(n10739) );
  NAND2X0 U16034 ( .IN1(n8521), .IN2(n10752), .QN(n15588) );
  NOR2X0 U16035 ( .IN1(n15589), .IN2(n15590), .QN(n15587) );
  NOR2X0 U16036 ( .IN1(n4506), .IN2(g320), .QN(n15590) );
  NOR2X0 U16037 ( .IN1(n4499), .IN2(g319), .QN(n15589) );
  INVX0 U16038 ( .INP(n10746), .ZN(n10725) );
  NAND2X0 U16039 ( .IN1(n15591), .IN2(n15592), .QN(n10746) );
  NAND2X0 U16040 ( .IN1(n8523), .IN2(n10752), .QN(n15592) );
  INVX0 U16041 ( .INP(n4520), .ZN(n10752) );
  NOR2X0 U16042 ( .IN1(n15593), .IN2(n15594), .QN(n15591) );
  NOR2X0 U16043 ( .IN1(n4506), .IN2(g317), .QN(n15594) );
  NOR2X0 U16044 ( .IN1(test_so18), .IN2(n4499), .QN(n15593) );
  NOR2X0 U16045 ( .IN1(n15202), .IN2(n15595), .QN(g23359) );
  XNOR2X1 U16046 ( .IN1(g3028), .IN2(n15422), .Q(n15595) );
  NOR2X0 U16047 ( .IN1(n9934), .IN2(n4481), .QN(n15422) );
  INVX0 U16048 ( .INP(n15596), .ZN(n9934) );
  INVX0 U16049 ( .INP(n9933), .ZN(n15202) );
  NAND2X0 U16050 ( .IN1(n14097), .IN2(n15597), .QN(n9933) );
  NAND2X0 U16051 ( .IN1(n15598), .IN2(n9931), .QN(n15597) );
  INVX0 U16052 ( .INP(g3234), .ZN(n9931) );
  NAND2X0 U16053 ( .IN1(n15599), .IN2(n15600), .QN(n15598) );
  NOR2X0 U16054 ( .IN1(n8695), .IN2(n4481), .QN(n15600) );
  NOR2X0 U16055 ( .IN1(g3036), .IN2(g3028), .QN(n15599) );
  NOR2X0 U16056 ( .IN1(n15205), .IN2(n15601), .QN(g23357) );
  XNOR2X1 U16057 ( .IN1(n4479), .IN2(n9871), .Q(n15601) );
  INVX0 U16058 ( .INP(n15416), .ZN(n9871) );
  NOR2X0 U16059 ( .IN1(n9872), .IN2(n4482), .QN(n15416) );
  INVX0 U16060 ( .INP(n9868), .ZN(n15205) );
  NAND2X0 U16061 ( .IN1(n9867), .IN2(n15602), .QN(n9868) );
  NAND2X0 U16062 ( .IN1(n16829), .IN2(n15603), .QN(n15602) );
  NAND2X0 U16063 ( .IN1(n15604), .IN2(n15605), .QN(n15603) );
  NOR2X0 U16064 ( .IN1(n8985), .IN2(n4482), .QN(n15605) );
  NOR2X0 U16065 ( .IN1(g2924), .IN2(g2917), .QN(n15604) );
  NOR2X0 U16066 ( .IN1(n10617), .IN2(n15606), .QN(g23348) );
  XOR2X1 U16067 ( .IN1(g2727), .IN2(n15427), .Q(n15606) );
  NOR2X0 U16068 ( .IN1(n14094), .IN2(n15607), .QN(g23339) );
  XNOR2X1 U16069 ( .IN1(n4420), .IN2(n15434), .Q(n15607) );
  NOR2X0 U16070 ( .IN1(n14097), .IN2(n15608), .QN(g23330) );
  NAND2X0 U16071 ( .IN1(n15609), .IN2(n4066), .QN(n15608) );
  NAND2X0 U16072 ( .IN1(n15610), .IN2(n14578), .QN(n4066) );
  NOR2X0 U16073 ( .IN1(n16834), .IN2(n9263), .QN(n15610) );
  NAND2X0 U16074 ( .IN1(n9263), .IN2(n15611), .QN(n15609) );
  NAND2X0 U16075 ( .IN1(n14578), .IN2(n7909), .QN(n15611) );
  NOR2X0 U16076 ( .IN1(n9261), .IN2(n9260), .QN(n14578) );
  INVX0 U16077 ( .INP(n14577), .ZN(n14097) );
  NOR2X0 U16078 ( .IN1(g3234), .IN2(n15596), .QN(n14577) );
  NOR2X0 U16079 ( .IN1(n15412), .IN2(n9260), .QN(n15596) );
  NAND2X0 U16080 ( .IN1(n15612), .IN2(n15613), .QN(n15412) );
  NOR2X0 U16081 ( .IN1(n15614), .IN2(n15615), .QN(n15613) );
  NAND2X0 U16082 ( .IN1(g3002), .IN2(g3013), .QN(n15615) );
  NAND2X0 U16083 ( .IN1(n7909), .IN2(n9280), .QN(n15614) );
  NOR2X0 U16084 ( .IN1(g3006), .IN2(n15616), .QN(n15612) );
  NAND2X0 U16085 ( .IN1(n9261), .IN2(g3024), .QN(n15616) );
  NOR2X0 U16086 ( .IN1(n14098), .IN2(n15617), .QN(g23329) );
  XNOR2X1 U16087 ( .IN1(n4421), .IN2(n15440), .Q(n15617) );
  NOR2X0 U16088 ( .IN1(n9684), .IN2(n15618), .QN(g23324) );
  XOR2X1 U16089 ( .IN1(g653), .IN2(n15444), .Q(n15618) );
  NAND2X0 U16090 ( .IN1(n15619), .IN2(n15620), .QN(g23137) );
  INVX0 U16091 ( .INP(n15621), .ZN(n15620) );
  NOR2X0 U16092 ( .IN1(g1866), .IN2(n9005), .QN(n15621) );
  NAND2X0 U16093 ( .IN1(n13980), .IN2(g1866), .QN(n15619) );
  NOR2X0 U16094 ( .IN1(n15622), .IN2(n15623), .QN(g23136) );
  NAND2X0 U16095 ( .IN1(n15444), .IN2(n13251), .QN(n15623) );
  NAND2X0 U16096 ( .IN1(n15624), .IN2(n15625), .QN(n15444) );
  NOR2X0 U16097 ( .IN1(n4478), .IN2(n4404), .QN(n15624) );
  NOR2X0 U16098 ( .IN1(n15626), .IN2(g633), .QN(n15622) );
  NOR2X0 U16099 ( .IN1(n4404), .IN2(n15627), .QN(n15626) );
  NAND2X0 U16100 ( .IN1(n15628), .IN2(n15629), .QN(g23133) );
  NAND2X0 U16101 ( .IN1(n4455), .IN2(g2562), .QN(n15629) );
  NAND2X0 U16102 ( .IN1(n13166), .IN2(g8167), .QN(n15628) );
  NAND2X0 U16103 ( .IN1(n15630), .IN2(n15631), .QN(g23132) );
  INVX0 U16104 ( .INP(n15632), .ZN(n15631) );
  NOR2X0 U16105 ( .IN1(g8087), .IN2(n8998), .QN(n15632) );
  NAND2X0 U16106 ( .IN1(n10478), .IN2(g8087), .QN(n15630) );
  NAND2X0 U16107 ( .IN1(n15633), .IN2(n15634), .QN(g23126) );
  NAND2X0 U16108 ( .IN1(n4465), .IN2(g1175), .QN(n15634) );
  NAND2X0 U16109 ( .IN1(n14023), .IN2(g1172), .QN(n15633) );
  NAND2X0 U16110 ( .IN1(n15635), .IN2(n15636), .QN(g23124) );
  NAND2X0 U16111 ( .IN1(n4457), .IN2(g1868), .QN(n15636) );
  NAND2X0 U16112 ( .IN1(n13980), .IN2(g8082), .QN(n15635) );
  NAND2X0 U16113 ( .IN1(n15637), .IN2(n15638), .QN(g23123) );
  INVX0 U16114 ( .INP(n15639), .ZN(n15638) );
  NOR2X0 U16115 ( .IN1(g8012), .IN2(n9007), .QN(n15639) );
  NAND2X0 U16116 ( .IN1(n11872), .IN2(g8012), .QN(n15637) );
  NAND2X0 U16117 ( .IN1(n15640), .IN2(n15641), .QN(g23117) );
  INVX0 U16118 ( .INP(n15642), .ZN(n15641) );
  NOR2X0 U16119 ( .IN1(g485), .IN2(n9022), .QN(n15642) );
  NAND2X0 U16120 ( .IN1(n14063), .IN2(g485), .QN(n15640) );
  NAND2X0 U16121 ( .IN1(n15643), .IN2(n15644), .QN(g23114) );
  INVX0 U16122 ( .INP(n15645), .ZN(n15644) );
  NOR2X0 U16123 ( .IN1(g8087), .IN2(n8996), .QN(n15645) );
  NAND2X0 U16124 ( .IN1(n13166), .IN2(g8087), .QN(n15643) );
  NAND2X0 U16125 ( .IN1(n15646), .IN2(n15647), .QN(g23111) );
  NAND2X0 U16126 ( .IN1(test_so44), .IN2(n4459), .QN(n15647) );
  NAND2X0 U16127 ( .IN1(n14023), .IN2(g8007), .QN(n15646) );
  NAND2X0 U16128 ( .IN1(n15648), .IN2(n15649), .QN(g23110) );
  INVX0 U16129 ( .INP(n15650), .ZN(n15649) );
  NOR2X0 U16130 ( .IN1(g7961), .IN2(n9015), .QN(n15650) );
  NAND2X0 U16131 ( .IN1(n10466), .IN2(g7961), .QN(n15648) );
  NAND2X0 U16132 ( .IN1(n15651), .IN2(n15652), .QN(g23097) );
  INVX0 U16133 ( .INP(n15653), .ZN(n15652) );
  NOR2X0 U16134 ( .IN1(g8012), .IN2(n9004), .QN(n15653) );
  NAND2X0 U16135 ( .IN1(n13980), .IN2(g8012), .QN(n15651) );
  NAND2X0 U16136 ( .IN1(n15654), .IN2(n15655), .QN(n13980) );
  NAND2X0 U16137 ( .IN1(g5511), .IN2(g1819), .QN(n15655) );
  NOR2X0 U16138 ( .IN1(n15656), .IN2(n15657), .QN(n15654) );
  NOR2X0 U16139 ( .IN1(n8704), .IN2(n11731), .QN(n15657) );
  INVX0 U16140 ( .INP(n15658), .ZN(n15656) );
  NAND2X0 U16141 ( .IN1(n4618), .IN2(test_so59), .QN(n15658) );
  NAND2X0 U16142 ( .IN1(n15659), .IN2(n15660), .QN(g23093) );
  NAND2X0 U16143 ( .IN1(n4461), .IN2(g487), .QN(n15660) );
  NAND2X0 U16144 ( .IN1(n14063), .IN2(g7956), .QN(n15659) );
  NAND2X0 U16145 ( .IN1(n15661), .IN2(n15662), .QN(g23092) );
  INVX0 U16146 ( .INP(n15663), .ZN(n15662) );
  NOR2X0 U16147 ( .IN1(n9024), .IN2(test_so23), .QN(n15663) );
  NAND2X0 U16148 ( .IN1(test_so23), .IN2(n11908), .QN(n15661) );
  NAND2X0 U16149 ( .IN1(n15664), .IN2(n15665), .QN(g23081) );
  INVX0 U16150 ( .INP(n15666), .ZN(n15665) );
  NOR2X0 U16151 ( .IN1(g7961), .IN2(n9013), .QN(n15666) );
  NAND2X0 U16152 ( .IN1(n14023), .IN2(g7961), .QN(n15664) );
  NAND2X0 U16153 ( .IN1(n15667), .IN2(n15668), .QN(n14023) );
  NAND2X0 U16154 ( .IN1(g1088), .IN2(g1131), .QN(n15668) );
  NOR2X0 U16155 ( .IN1(n15669), .IN2(n15670), .QN(n15667) );
  NOR2X0 U16156 ( .IN1(n8708), .IN2(n4364), .QN(n15670) );
  NOR2X0 U16157 ( .IN1(n8726), .IN2(n4363), .QN(n15669) );
  NAND2X0 U16158 ( .IN1(n15671), .IN2(n15672), .QN(g23076) );
  INVX0 U16159 ( .INP(n15673), .ZN(n15672) );
  NOR2X0 U16160 ( .IN1(g2560), .IN2(n8999), .QN(n15673) );
  NAND2X0 U16161 ( .IN1(n10478), .IN2(g2560), .QN(n15671) );
  NAND2X0 U16162 ( .IN1(n15674), .IN2(n15675), .QN(g23067) );
  INVX0 U16163 ( .INP(n15676), .ZN(n15675) );
  NOR2X0 U16164 ( .IN1(n9021), .IN2(test_so23), .QN(n15676) );
  NAND2X0 U16165 ( .IN1(test_so23), .IN2(n14063), .QN(n15674) );
  NAND2X0 U16166 ( .IN1(n15677), .IN2(n15678), .QN(n14063) );
  NAND2X0 U16167 ( .IN1(g5437), .IN2(g438), .QN(n15678) );
  NOR2X0 U16168 ( .IN1(n15679), .IN2(n15680), .QN(n15677) );
  NOR2X0 U16169 ( .IN1(n8734), .IN2(n12562), .QN(n15680) );
  NOR2X0 U16170 ( .IN1(n8733), .IN2(n12563), .QN(n15679) );
  NAND2X0 U16171 ( .IN1(n15681), .IN2(n15682), .QN(g23058) );
  INVX0 U16172 ( .INP(n15683), .ZN(n15682) );
  NOR2X0 U16173 ( .IN1(g1866), .IN2(n9008), .QN(n15683) );
  NAND2X0 U16174 ( .IN1(n11872), .IN2(g1866), .QN(n15681) );
  NAND2X0 U16175 ( .IN1(n15684), .IN2(n15685), .QN(g23047) );
  NAND2X0 U16176 ( .IN1(n4455), .IN2(g2559), .QN(n15685) );
  NAND2X0 U16177 ( .IN1(n10478), .IN2(g8167), .QN(n15684) );
  INVX0 U16178 ( .INP(n4285), .ZN(n10478) );
  NAND2X0 U16179 ( .IN1(n15686), .IN2(n15687), .QN(n4285) );
  NAND2X0 U16180 ( .IN1(g5555), .IN2(g2492), .QN(n15687) );
  NOR2X0 U16181 ( .IN1(n15688), .IN2(n15689), .QN(n15686) );
  NOR2X0 U16182 ( .IN1(n8702), .IN2(n12443), .QN(n15689) );
  NOR2X0 U16183 ( .IN1(n8715), .IN2(n13976), .QN(n15688) );
  NAND2X0 U16184 ( .IN1(n15690), .IN2(n15691), .QN(g23039) );
  INVX0 U16185 ( .INP(n15692), .ZN(n15691) );
  NOR2X0 U16186 ( .IN1(g1172), .IN2(n9016), .QN(n15692) );
  NAND2X0 U16187 ( .IN1(n10466), .IN2(g1172), .QN(n15690) );
  NAND2X0 U16188 ( .IN1(n15693), .IN2(n15694), .QN(g23030) );
  NAND2X0 U16189 ( .IN1(n4457), .IN2(g1865), .QN(n15694) );
  NAND2X0 U16190 ( .IN1(n11872), .IN2(g8082), .QN(n15693) );
  INVX0 U16191 ( .INP(n4284), .ZN(n11872) );
  NAND2X0 U16192 ( .IN1(n15695), .IN2(n15696), .QN(n4284) );
  NAND2X0 U16193 ( .IN1(g5511), .IN2(g1798), .QN(n15696) );
  NOR2X0 U16194 ( .IN1(n15697), .IN2(n15698), .QN(n15695) );
  NOR2X0 U16195 ( .IN1(n8706), .IN2(n11731), .QN(n15698) );
  INVX0 U16196 ( .INP(g7014), .ZN(n11731) );
  NOR2X0 U16197 ( .IN1(n8721), .IN2(n12488), .QN(n15697) );
  INVX0 U16198 ( .INP(n4618), .ZN(n12488) );
  NAND2X0 U16199 ( .IN1(n15699), .IN2(n15700), .QN(g23022) );
  INVX0 U16200 ( .INP(n15701), .ZN(n15700) );
  NOR2X0 U16201 ( .IN1(g485), .IN2(n9025), .QN(n15701) );
  NAND2X0 U16202 ( .IN1(n11908), .IN2(g485), .QN(n15699) );
  NAND2X0 U16203 ( .IN1(n15702), .IN2(n15703), .QN(g23014) );
  NAND2X0 U16204 ( .IN1(n4459), .IN2(g1171), .QN(n15703) );
  NAND2X0 U16205 ( .IN1(n10466), .IN2(g8007), .QN(n15702) );
  INVX0 U16206 ( .INP(n4283), .ZN(n10466) );
  NAND2X0 U16207 ( .IN1(n15704), .IN2(n15705), .QN(n4283) );
  NAND2X0 U16208 ( .IN1(g1088), .IN2(g1110), .QN(n15705) );
  NOR2X0 U16209 ( .IN1(n15706), .IN2(n15707), .QN(n15704) );
  NOR2X0 U16210 ( .IN1(n8709), .IN2(n4364), .QN(n15707) );
  NOR2X0 U16211 ( .IN1(n8730), .IN2(n4363), .QN(n15706) );
  NAND2X0 U16212 ( .IN1(n15708), .IN2(n15709), .QN(g23000) );
  NAND2X0 U16213 ( .IN1(n4461), .IN2(g484), .QN(n15709) );
  NAND2X0 U16214 ( .IN1(n11908), .IN2(g7956), .QN(n15708) );
  INVX0 U16215 ( .INP(n4282), .ZN(n11908) );
  NAND2X0 U16216 ( .IN1(n15710), .IN2(n15711), .QN(n4282) );
  NAND2X0 U16217 ( .IN1(g5437), .IN2(g417), .QN(n15711) );
  NOR2X0 U16218 ( .IN1(n15712), .IN2(n15713), .QN(n15710) );
  NOR2X0 U16219 ( .IN1(n8740), .IN2(n12562), .QN(n15713) );
  INVX0 U16220 ( .INP(g6447), .ZN(n12562) );
  NOR2X0 U16221 ( .IN1(n8739), .IN2(n12563), .QN(n15712) );
  INVX0 U16222 ( .INP(n4640), .ZN(n12563) );
  NAND2X0 U16223 ( .IN1(n15714), .IN2(n15715), .QN(g22687) );
  NAND2X0 U16224 ( .IN1(n15716), .IN2(n15717), .QN(n15715) );
  INVX0 U16225 ( .INP(n14402), .ZN(n15717) );
  NOR2X0 U16226 ( .IN1(n4303), .IN2(n10100), .QN(n15716) );
  NAND2X0 U16227 ( .IN1(n15718), .IN2(n15719), .QN(n15714) );
  NAND2X0 U16228 ( .IN1(n10628), .IN2(n14402), .QN(n15718) );
  NAND2X0 U16229 ( .IN1(n15720), .IN2(n15721), .QN(n14402) );
  NAND2X0 U16230 ( .IN1(g7390), .IN2(g2568), .QN(n15721) );
  NOR2X0 U16231 ( .IN1(n15722), .IN2(n15723), .QN(n15720) );
  NOR2X0 U16232 ( .IN1(n8745), .IN2(n4314), .QN(n15723) );
  NOR2X0 U16233 ( .IN1(n8747), .IN2(n4299), .QN(n15722) );
  NAND2X0 U16234 ( .IN1(n15724), .IN2(n15725), .QN(g22651) );
  NAND2X0 U16235 ( .IN1(n15726), .IN2(n15727), .QN(n15725) );
  INVX0 U16236 ( .INP(n14413), .ZN(n15727) );
  NOR2X0 U16237 ( .IN1(n4297), .IN2(n10237), .QN(n15726) );
  NAND2X0 U16238 ( .IN1(n15728), .IN2(n15719), .QN(n15724) );
  NAND2X0 U16239 ( .IN1(n10266), .IN2(n14413), .QN(n15728) );
  NAND2X0 U16240 ( .IN1(n15729), .IN2(n15730), .QN(n14413) );
  NAND2X0 U16241 ( .IN1(g1930), .IN2(g1877), .QN(n15730) );
  NOR2X0 U16242 ( .IN1(n15731), .IN2(n15732), .QN(n15729) );
  NOR2X0 U16243 ( .IN1(n8752), .IN2(n4315), .QN(n15732) );
  INVX0 U16244 ( .INP(n15733), .ZN(n15731) );
  NAND2X0 U16245 ( .IN1(n12749), .IN2(test_so68), .QN(n15733) );
  NAND2X0 U16246 ( .IN1(n15734), .IN2(n15735), .QN(g22615) );
  NAND2X0 U16247 ( .IN1(n15736), .IN2(n15737), .QN(n15735) );
  INVX0 U16248 ( .INP(n14424), .ZN(n15737) );
  NOR2X0 U16249 ( .IN1(n4304), .IN2(n10380), .QN(n15736) );
  NAND2X0 U16250 ( .IN1(n15738), .IN2(n15719), .QN(n15734) );
  NAND2X0 U16251 ( .IN1(n10409), .IN2(n14424), .QN(n15738) );
  NAND2X0 U16252 ( .IN1(n15739), .IN2(n15740), .QN(n14424) );
  NAND2X0 U16253 ( .IN1(test_so47), .IN2(n12608), .QN(n15740) );
  NOR2X0 U16254 ( .IN1(n15741), .IN2(n15742), .QN(n15739) );
  NOR2X0 U16255 ( .IN1(n8753), .IN2(n4316), .QN(n15742) );
  NOR2X0 U16256 ( .IN1(n8749), .IN2(n4300), .QN(n15741) );
  NAND2X0 U16257 ( .IN1(n15743), .IN2(n15744), .QN(g22578) );
  NAND2X0 U16258 ( .IN1(n15745), .IN2(n15746), .QN(n15744) );
  INVX0 U16259 ( .INP(n14431), .ZN(n15746) );
  NOR2X0 U16260 ( .IN1(n9961), .IN2(n9285), .QN(n15745) );
  NAND2X0 U16261 ( .IN1(n15747), .IN2(n15719), .QN(n15743) );
  NAND2X0 U16262 ( .IN1(n10001), .IN2(n14431), .QN(n15747) );
  NAND2X0 U16263 ( .IN1(n15748), .IN2(n15749), .QN(n14431) );
  NAND2X0 U16264 ( .IN1(g6642), .IN2(g493), .QN(n15749) );
  NOR2X0 U16265 ( .IN1(n15750), .IN2(n15751), .QN(n15748) );
  NOR2X0 U16266 ( .IN1(n8750), .IN2(n4313), .QN(n15751) );
  NOR2X0 U16267 ( .IN1(n8746), .IN2(n15378), .QN(n15750) );
  NOR2X0 U16268 ( .IN1(n15752), .IN2(n15753), .QN(g22299) );
  NOR2X0 U16269 ( .IN1(n14693), .IN2(test_so95), .QN(n15753) );
  NOR2X0 U16270 ( .IN1(n10617), .IN2(n15754), .QN(g22284) );
  NOR2X0 U16271 ( .IN1(n14697), .IN2(g2813), .QN(n15754) );
  NOR2X0 U16272 ( .IN1(n15755), .IN2(n15756), .QN(g22280) );
  INVX0 U16273 ( .INP(n15757), .ZN(n15756) );
  NAND2X0 U16274 ( .IN1(n14700), .IN2(n9220), .QN(n15757) );
  NOR2X0 U16275 ( .IN1(n14094), .IN2(n15758), .QN(g22267) );
  NOR2X0 U16276 ( .IN1(n14778), .IN2(g2119), .QN(n15758) );
  INVX0 U16277 ( .INP(n15759), .ZN(g22263) );
  NAND2X0 U16278 ( .IN1(n15760), .IN2(n15761), .QN(n15759) );
  NAND2X0 U16279 ( .IN1(n14782), .IN2(n9221), .QN(n15761) );
  NOR2X0 U16280 ( .IN1(n14098), .IN2(n15762), .QN(g22247) );
  NOR2X0 U16281 ( .IN1(n14861), .IN2(g1425), .QN(n15762) );
  NOR2X0 U16282 ( .IN1(n15763), .IN2(n15764), .QN(g22242) );
  INVX0 U16283 ( .INP(n15765), .ZN(n15764) );
  NAND2X0 U16284 ( .IN1(n14864), .IN2(n9222), .QN(n15765) );
  NOR2X0 U16285 ( .IN1(n9684), .IN2(n15766), .QN(g22231) );
  NOR2X0 U16286 ( .IN1(n14948), .IN2(g739), .QN(n15766) );
  NAND2X0 U16287 ( .IN1(n15767), .IN2(n15768), .QN(g22200) );
  NAND2X0 U16288 ( .IN1(n4373), .IN2(n15769), .QN(n15768) );
  NAND2X0 U16289 ( .IN1(n15214), .IN2(g2208), .QN(n15767) );
  NAND2X0 U16290 ( .IN1(n15770), .IN2(n15771), .QN(g22194) );
  INVX0 U16291 ( .INP(n15772), .ZN(n15771) );
  NOR2X0 U16292 ( .IN1(n15769), .IN2(n8793), .QN(n15772) );
  NAND2X0 U16293 ( .IN1(n10796), .IN2(n15769), .QN(n15770) );
  NAND2X0 U16294 ( .IN1(n15773), .IN2(n15774), .QN(g22193) );
  NAND2X0 U16295 ( .IN1(n15775), .IN2(n4373), .QN(n15774) );
  INVX0 U16296 ( .INP(n15776), .ZN(n15773) );
  NOR2X0 U16297 ( .IN1(n15775), .IN2(n9167), .QN(n15776) );
  NAND2X0 U16298 ( .IN1(n15777), .IN2(n15778), .QN(g22192) );
  NAND2X0 U16299 ( .IN1(n4377), .IN2(n15769), .QN(n15778) );
  NAND2X0 U16300 ( .IN1(n15214), .IN2(g2205), .QN(n15777) );
  NAND2X0 U16301 ( .IN1(n15779), .IN2(n15780), .QN(g22191) );
  NAND2X0 U16302 ( .IN1(n4374), .IN2(n15781), .QN(n15780) );
  NAND2X0 U16303 ( .IN1(n15216), .IN2(g1514), .QN(n15779) );
  NAND2X0 U16304 ( .IN1(n15782), .IN2(n15783), .QN(g22185) );
  NAND2X0 U16305 ( .IN1(test_so75), .IN2(n15784), .QN(n15783) );
  NAND2X0 U16306 ( .IN1(n15775), .IN2(n10796), .QN(n15782) );
  NAND2X0 U16307 ( .IN1(n15785), .IN2(n15786), .QN(g22184) );
  NAND2X0 U16308 ( .IN1(n15214), .IN2(g2235), .QN(n15786) );
  NAND2X0 U16309 ( .IN1(n10978), .IN2(n15769), .QN(n15785) );
  NAND2X0 U16310 ( .IN1(n15787), .IN2(n15788), .QN(g22183) );
  NAND2X0 U16311 ( .IN1(n15789), .IN2(n4373), .QN(n15788) );
  NAND2X0 U16312 ( .IN1(n15790), .IN2(g2209), .QN(n15787) );
  NAND2X0 U16313 ( .IN1(n15791), .IN2(n15792), .QN(g22182) );
  NAND2X0 U16314 ( .IN1(n15775), .IN2(n4377), .QN(n15792) );
  INVX0 U16315 ( .INP(n15793), .ZN(n15791) );
  NOR2X0 U16316 ( .IN1(n15775), .IN2(n9169), .QN(n15793) );
  NAND2X0 U16317 ( .IN1(n15794), .IN2(n15795), .QN(g22180) );
  INVX0 U16318 ( .INP(n15796), .ZN(n15795) );
  NOR2X0 U16319 ( .IN1(n15781), .IN2(n8803), .QN(n15796) );
  NAND2X0 U16320 ( .IN1(n10835), .IN2(n15781), .QN(n15794) );
  NAND2X0 U16321 ( .IN1(n15797), .IN2(n15798), .QN(g22179) );
  NAND2X0 U16322 ( .IN1(n15799), .IN2(n4374), .QN(n15798) );
  INVX0 U16323 ( .INP(n15800), .ZN(n15797) );
  NOR2X0 U16324 ( .IN1(n15799), .IN2(n9182), .QN(n15800) );
  NAND2X0 U16325 ( .IN1(n15801), .IN2(n15802), .QN(g22178) );
  NAND2X0 U16326 ( .IN1(n4378), .IN2(n15781), .QN(n15802) );
  NAND2X0 U16327 ( .IN1(n15216), .IN2(g1511), .QN(n15801) );
  NAND2X0 U16328 ( .IN1(n15803), .IN2(n15804), .QN(g22177) );
  NAND2X0 U16329 ( .IN1(n15805), .IN2(n4375), .QN(n15804) );
  INVX0 U16330 ( .INP(n15806), .ZN(n15803) );
  NOR2X0 U16331 ( .IN1(n15805), .IN2(n8826), .QN(n15806) );
  NAND2X0 U16332 ( .IN1(n15807), .IN2(n15808), .QN(g22173) );
  INVX0 U16333 ( .INP(n15809), .ZN(n15808) );
  NOR2X0 U16334 ( .IN1(n15789), .IN2(n8794), .QN(n15809) );
  NAND2X0 U16335 ( .IN1(n15789), .IN2(n10796), .QN(n15807) );
  INVX0 U16336 ( .INP(n11996), .ZN(n10796) );
  NAND2X0 U16337 ( .IN1(n15810), .IN2(n15811), .QN(n11996) );
  NAND2X0 U16338 ( .IN1(n8856), .IN2(test_so73), .QN(n15811) );
  NOR2X0 U16339 ( .IN1(n15812), .IN2(n15813), .QN(n15810) );
  NOR2X0 U16340 ( .IN1(n4367), .IN2(g2247), .QN(n15813) );
  NOR2X0 U16341 ( .IN1(n4324), .IN2(g2248), .QN(n15812) );
  NAND2X0 U16342 ( .IN1(n15814), .IN2(n15815), .QN(g22172) );
  INVX0 U16343 ( .INP(n15816), .ZN(n15815) );
  NOR2X0 U16344 ( .IN1(n15775), .IN2(n8785), .QN(n15816) );
  NAND2X0 U16345 ( .IN1(n10978), .IN2(n15775), .QN(n15814) );
  NAND2X0 U16346 ( .IN1(n15817), .IN2(n15818), .QN(g22171) );
  NAND2X0 U16347 ( .IN1(n4287), .IN2(n15769), .QN(n15818) );
  NAND2X0 U16348 ( .IN1(n15214), .IN2(g2232), .QN(n15817) );
  NAND2X0 U16349 ( .IN1(n15819), .IN2(n15820), .QN(g22170) );
  NAND2X0 U16350 ( .IN1(n15789), .IN2(n4377), .QN(n15820) );
  NAND2X0 U16351 ( .IN1(n15790), .IN2(g2206), .QN(n15819) );
  NAND2X0 U16352 ( .IN1(n15821), .IN2(n15822), .QN(g22169) );
  NAND2X0 U16353 ( .IN1(n15823), .IN2(g1546), .QN(n15822) );
  NAND2X0 U16354 ( .IN1(n15799), .IN2(n10835), .QN(n15821) );
  NAND2X0 U16355 ( .IN1(n15824), .IN2(n15825), .QN(g22168) );
  INVX0 U16356 ( .INP(n15826), .ZN(n15825) );
  NOR2X0 U16357 ( .IN1(n15781), .IN2(n8787), .QN(n15826) );
  NAND2X0 U16358 ( .IN1(n11025), .IN2(n15781), .QN(n15824) );
  NAND2X0 U16359 ( .IN1(n15827), .IN2(n15828), .QN(g22167) );
  NAND2X0 U16360 ( .IN1(test_so52), .IN2(n15829), .QN(n15828) );
  NAND2X0 U16361 ( .IN1(n15830), .IN2(n4374), .QN(n15827) );
  NAND2X0 U16362 ( .IN1(n15831), .IN2(n15832), .QN(g22166) );
  NAND2X0 U16363 ( .IN1(n15799), .IN2(n4378), .QN(n15832) );
  INVX0 U16364 ( .INP(n15833), .ZN(n15831) );
  NOR2X0 U16365 ( .IN1(n15799), .IN2(n9183), .QN(n15833) );
  NAND2X0 U16366 ( .IN1(n15834), .IN2(n15835), .QN(g22164) );
  NAND2X0 U16367 ( .IN1(n15218), .IN2(g850), .QN(n15835) );
  INVX0 U16368 ( .INP(n15805), .ZN(n15218) );
  NAND2X0 U16369 ( .IN1(n15805), .IN2(n10876), .QN(n15834) );
  NAND2X0 U16370 ( .IN1(n15836), .IN2(n15837), .QN(g22163) );
  NAND2X0 U16371 ( .IN1(n15838), .IN2(n4375), .QN(n15837) );
  NAND2X0 U16372 ( .IN1(n15839), .IN2(g822), .QN(n15836) );
  NAND2X0 U16373 ( .IN1(n15840), .IN2(n15841), .QN(g22162) );
  NAND2X0 U16374 ( .IN1(n4379), .IN2(n15805), .QN(n15841) );
  INVX0 U16375 ( .INP(n15842), .ZN(n15840) );
  NOR2X0 U16376 ( .IN1(n15805), .IN2(n8827), .QN(n15842) );
  NAND2X0 U16377 ( .IN1(n15843), .IN2(n15844), .QN(g22161) );
  NAND2X0 U16378 ( .IN1(n4376), .IN2(n15845), .QN(n15844) );
  NAND2X0 U16379 ( .IN1(n15220), .IN2(g132), .QN(n15843) );
  NAND2X0 U16380 ( .IN1(n15846), .IN2(n15847), .QN(g22155) );
  NAND2X0 U16381 ( .IN1(n15790), .IN2(g2236), .QN(n15847) );
  NAND2X0 U16382 ( .IN1(n15789), .IN2(n10978), .QN(n15846) );
  INVX0 U16383 ( .INP(n12020), .ZN(n10978) );
  NAND2X0 U16384 ( .IN1(n15848), .IN2(n15849), .QN(n12020) );
  NAND2X0 U16385 ( .IN1(n8853), .IN2(test_so73), .QN(n15849) );
  NOR2X0 U16386 ( .IN1(n15850), .IN2(n15851), .QN(n15848) );
  NOR2X0 U16387 ( .IN1(n4367), .IN2(g2250), .QN(n15851) );
  NOR2X0 U16388 ( .IN1(n4324), .IN2(g2251), .QN(n15850) );
  NAND2X0 U16389 ( .IN1(n15852), .IN2(n15853), .QN(g22154) );
  NAND2X0 U16390 ( .IN1(n15775), .IN2(n4287), .QN(n15853) );
  INVX0 U16391 ( .INP(n15854), .ZN(n15852) );
  NOR2X0 U16392 ( .IN1(n15775), .IN2(n9156), .QN(n15854) );
  NAND2X0 U16393 ( .IN1(n15855), .IN2(n15856), .QN(g22153) );
  NAND2X0 U16394 ( .IN1(n4563), .IN2(n15769), .QN(n15856) );
  NAND2X0 U16395 ( .IN1(n15214), .IN2(g2229), .QN(n15855) );
  NAND2X0 U16396 ( .IN1(n15857), .IN2(n15858), .QN(g22152) );
  INVX0 U16397 ( .INP(n15859), .ZN(n15858) );
  NOR2X0 U16398 ( .IN1(n15830), .IN2(n8805), .QN(n15859) );
  NAND2X0 U16399 ( .IN1(n15830), .IN2(n10835), .QN(n15857) );
  INVX0 U16400 ( .INP(n15860), .ZN(n10835) );
  NAND2X0 U16401 ( .IN1(n15861), .IN2(n15862), .QN(n15860) );
  NAND2X0 U16402 ( .IN1(n8867), .IN2(g6782), .QN(n15862) );
  NOR2X0 U16403 ( .IN1(n15863), .IN2(n15864), .QN(n15861) );
  NOR2X0 U16404 ( .IN1(test_so54), .IN2(n4368), .QN(n15864) );
  NOR2X0 U16405 ( .IN1(n4317), .IN2(g1554), .QN(n15863) );
  NAND2X0 U16406 ( .IN1(n15865), .IN2(n15866), .QN(g22151) );
  NAND2X0 U16407 ( .IN1(n15823), .IN2(g1543), .QN(n15866) );
  NAND2X0 U16408 ( .IN1(n11025), .IN2(n15799), .QN(n15865) );
  NAND2X0 U16409 ( .IN1(n15867), .IN2(n15868), .QN(g22150) );
  NAND2X0 U16410 ( .IN1(n4288), .IN2(n15781), .QN(n15868) );
  NAND2X0 U16411 ( .IN1(n15216), .IN2(g1538), .QN(n15867) );
  NAND2X0 U16412 ( .IN1(n15869), .IN2(n15870), .QN(g22149) );
  NAND2X0 U16413 ( .IN1(n15830), .IN2(n4378), .QN(n15870) );
  NAND2X0 U16414 ( .IN1(n15829), .IN2(g1512), .QN(n15869) );
  NAND2X0 U16415 ( .IN1(n15871), .IN2(n15872), .QN(g22148) );
  INVX0 U16416 ( .INP(n15873), .ZN(n15872) );
  NOR2X0 U16417 ( .IN1(n15838), .IN2(n8815), .QN(n15873) );
  NAND2X0 U16418 ( .IN1(n15838), .IN2(n10876), .QN(n15871) );
  NAND2X0 U16419 ( .IN1(n15874), .IN2(n15875), .QN(g22147) );
  INVX0 U16420 ( .INP(n15876), .ZN(n15875) );
  NOR2X0 U16421 ( .IN1(n15805), .IN2(n8817), .QN(n15876) );
  NAND2X0 U16422 ( .IN1(n11066), .IN2(n15805), .QN(n15874) );
  NAND2X0 U16423 ( .IN1(n15877), .IN2(n15878), .QN(g22146) );
  NAND2X0 U16424 ( .IN1(n15879), .IN2(n4375), .QN(n15878) );
  NAND2X0 U16425 ( .IN1(n15880), .IN2(g821), .QN(n15877) );
  NAND2X0 U16426 ( .IN1(n15881), .IN2(n15882), .QN(g22145) );
  NAND2X0 U16427 ( .IN1(n15838), .IN2(n4379), .QN(n15882) );
  NAND2X0 U16428 ( .IN1(n15839), .IN2(g819), .QN(n15881) );
  NAND2X0 U16429 ( .IN1(n15883), .IN2(n15884), .QN(g22143) );
  INVX0 U16430 ( .INP(n15885), .ZN(n15884) );
  NOR2X0 U16431 ( .IN1(n15845), .IN2(n8828), .QN(n15885) );
  NAND2X0 U16432 ( .IN1(n10928), .IN2(n15845), .QN(n15883) );
  NAND2X0 U16433 ( .IN1(n15886), .IN2(n15887), .QN(g22142) );
  NAND2X0 U16434 ( .IN1(n15888), .IN2(n4376), .QN(n15887) );
  INVX0 U16435 ( .INP(n15889), .ZN(n15886) );
  NOR2X0 U16436 ( .IN1(n15888), .IN2(n9212), .QN(n15889) );
  NAND2X0 U16437 ( .IN1(n15890), .IN2(n15891), .QN(g22141) );
  NAND2X0 U16438 ( .IN1(n4380), .IN2(n15845), .QN(n15891) );
  NAND2X0 U16439 ( .IN1(n15220), .IN2(g129), .QN(n15890) );
  NAND2X0 U16440 ( .IN1(n15892), .IN2(n15893), .QN(g22140) );
  NAND2X0 U16441 ( .IN1(n15789), .IN2(n4287), .QN(n15893) );
  NAND2X0 U16442 ( .IN1(n15790), .IN2(g2233), .QN(n15892) );
  NAND2X0 U16443 ( .IN1(n15894), .IN2(n15895), .QN(g22139) );
  NAND2X0 U16444 ( .IN1(n15775), .IN2(n4563), .QN(n15895) );
  INVX0 U16445 ( .INP(n15896), .ZN(n15894) );
  NOR2X0 U16446 ( .IN1(n15775), .IN2(n9158), .QN(n15896) );
  NAND2X0 U16447 ( .IN1(n15897), .IN2(n15898), .QN(g22138) );
  NAND2X0 U16448 ( .IN1(n4555), .IN2(n15769), .QN(n15898) );
  NAND2X0 U16449 ( .IN1(n15214), .IN2(g2226), .QN(n15897) );
  NAND2X0 U16450 ( .IN1(n15899), .IN2(n15900), .QN(g22132) );
  INVX0 U16451 ( .INP(n15901), .ZN(n15900) );
  NOR2X0 U16452 ( .IN1(n15830), .IN2(n8789), .QN(n15901) );
  NAND2X0 U16453 ( .IN1(n15830), .IN2(n11025), .QN(n15899) );
  INVX0 U16454 ( .INP(n12116), .ZN(n11025) );
  NAND2X0 U16455 ( .IN1(n15902), .IN2(n15903), .QN(n12116) );
  NAND2X0 U16456 ( .IN1(n8865), .IN2(g6782), .QN(n15903) );
  NOR2X0 U16457 ( .IN1(n15904), .IN2(n15905), .QN(n15902) );
  NOR2X0 U16458 ( .IN1(n4368), .IN2(g1556), .QN(n15905) );
  NOR2X0 U16459 ( .IN1(n4317), .IN2(g1557), .QN(n15904) );
  NAND2X0 U16460 ( .IN1(n15906), .IN2(n15907), .QN(g22131) );
  NAND2X0 U16461 ( .IN1(n15799), .IN2(n4288), .QN(n15907) );
  INVX0 U16462 ( .INP(n15908), .ZN(n15906) );
  NOR2X0 U16463 ( .IN1(n15799), .IN2(n9171), .QN(n15908) );
  NAND2X0 U16464 ( .IN1(n15909), .IN2(n15910), .QN(g22130) );
  NAND2X0 U16465 ( .IN1(n4565), .IN2(n15781), .QN(n15910) );
  NAND2X0 U16466 ( .IN1(n15216), .IN2(g1535), .QN(n15909) );
  NAND2X0 U16467 ( .IN1(n15911), .IN2(n15912), .QN(g22129) );
  INVX0 U16468 ( .INP(n15913), .ZN(n15912) );
  NOR2X0 U16469 ( .IN1(n15879), .IN2(n8816), .QN(n15913) );
  NAND2X0 U16470 ( .IN1(n15879), .IN2(n10876), .QN(n15911) );
  INVX0 U16471 ( .INP(n15914), .ZN(n10876) );
  NAND2X0 U16472 ( .IN1(n15915), .IN2(n15916), .QN(n15914) );
  NAND2X0 U16473 ( .IN1(n8878), .IN2(test_so31), .QN(n15916) );
  NOR2X0 U16474 ( .IN1(n15917), .IN2(n15918), .QN(n15915) );
  NOR2X0 U16475 ( .IN1(n4323), .IN2(g860), .QN(n15918) );
  NOR2X0 U16476 ( .IN1(n4312), .IN2(g861), .QN(n15917) );
  NAND2X0 U16477 ( .IN1(n15919), .IN2(n15920), .QN(g22128) );
  NAND2X0 U16478 ( .IN1(n15839), .IN2(g849), .QN(n15920) );
  NAND2X0 U16479 ( .IN1(n11066), .IN2(n15838), .QN(n15919) );
  NAND2X0 U16480 ( .IN1(n15921), .IN2(n15922), .QN(g22127) );
  NAND2X0 U16481 ( .IN1(n4289), .IN2(n15805), .QN(n15922) );
  INVX0 U16482 ( .INP(n15923), .ZN(n15921) );
  NOR2X0 U16483 ( .IN1(n15805), .IN2(n8820), .QN(n15923) );
  NAND2X0 U16484 ( .IN1(n15924), .IN2(n15925), .QN(g22126) );
  NAND2X0 U16485 ( .IN1(n15879), .IN2(n4379), .QN(n15925) );
  NAND2X0 U16486 ( .IN1(n15880), .IN2(g818), .QN(n15924) );
  NAND2X0 U16487 ( .IN1(n15926), .IN2(n15927), .QN(g22125) );
  NAND2X0 U16488 ( .IN1(n15928), .IN2(g164), .QN(n15927) );
  NAND2X0 U16489 ( .IN1(n15888), .IN2(n10928), .QN(n15926) );
  NAND2X0 U16490 ( .IN1(n15929), .IN2(n15930), .QN(g22124) );
  INVX0 U16491 ( .INP(n15931), .ZN(n15930) );
  NOR2X0 U16492 ( .IN1(n15845), .IN2(n8790), .QN(n15931) );
  NAND2X0 U16493 ( .IN1(n11093), .IN2(n15845), .QN(n15929) );
  NAND2X0 U16494 ( .IN1(n15932), .IN2(n15933), .QN(g22123) );
  NAND2X0 U16495 ( .IN1(n15934), .IN2(n4376), .QN(n15933) );
  NAND2X0 U16496 ( .IN1(n15935), .IN2(g133), .QN(n15932) );
  NAND2X0 U16497 ( .IN1(n15936), .IN2(n15937), .QN(g22122) );
  NAND2X0 U16498 ( .IN1(n15888), .IN2(n4380), .QN(n15937) );
  INVX0 U16499 ( .INP(n15938), .ZN(n15936) );
  NOR2X0 U16500 ( .IN1(n15888), .IN2(n9214), .QN(n15938) );
  NAND2X0 U16501 ( .IN1(n15939), .IN2(n15940), .QN(g22117) );
  NAND2X0 U16502 ( .IN1(n15789), .IN2(n4563), .QN(n15940) );
  NAND2X0 U16503 ( .IN1(n15790), .IN2(g2230), .QN(n15939) );
  NAND2X0 U16504 ( .IN1(n15941), .IN2(n15942), .QN(g22116) );
  NAND2X0 U16505 ( .IN1(n15775), .IN2(n4555), .QN(n15942) );
  INVX0 U16506 ( .INP(n15943), .ZN(n15941) );
  NOR2X0 U16507 ( .IN1(n15775), .IN2(n9160), .QN(n15943) );
  NAND2X0 U16508 ( .IN1(n15944), .IN2(n15945), .QN(g22115) );
  NAND2X0 U16509 ( .IN1(n4325), .IN2(n15769), .QN(n15945) );
  NAND2X0 U16510 ( .IN1(n15214), .IN2(g2223), .QN(n15944) );
  NAND2X0 U16511 ( .IN1(n15946), .IN2(n15947), .QN(g22114) );
  NAND2X0 U16512 ( .IN1(n15830), .IN2(n4288), .QN(n15947) );
  NAND2X0 U16513 ( .IN1(n15829), .IN2(g1539), .QN(n15946) );
  NAND2X0 U16514 ( .IN1(n15948), .IN2(n15949), .QN(g22113) );
  NAND2X0 U16515 ( .IN1(test_so53), .IN2(n15823), .QN(n15949) );
  INVX0 U16516 ( .INP(n15799), .ZN(n15823) );
  NAND2X0 U16517 ( .IN1(n15799), .IN2(n4565), .QN(n15948) );
  NAND2X0 U16518 ( .IN1(n15950), .IN2(n15951), .QN(g22112) );
  NAND2X0 U16519 ( .IN1(n4557), .IN2(n15781), .QN(n15951) );
  NAND2X0 U16520 ( .IN1(n15216), .IN2(g1532), .QN(n15950) );
  NAND2X0 U16521 ( .IN1(n15952), .IN2(n15953), .QN(g22106) );
  NAND2X0 U16522 ( .IN1(n15880), .IN2(g848), .QN(n15953) );
  NAND2X0 U16523 ( .IN1(n15879), .IN2(n11066), .QN(n15952) );
  INVX0 U16524 ( .INP(n12257), .ZN(n11066) );
  NAND2X0 U16525 ( .IN1(n15954), .IN2(n15955), .QN(n12257) );
  NAND2X0 U16526 ( .IN1(n8875), .IN2(test_so31), .QN(n15955) );
  NOR2X0 U16527 ( .IN1(n15956), .IN2(n15957), .QN(n15954) );
  NOR2X0 U16528 ( .IN1(n4323), .IN2(g863), .QN(n15957) );
  NOR2X0 U16529 ( .IN1(n4312), .IN2(g864), .QN(n15956) );
  NAND2X0 U16530 ( .IN1(n15958), .IN2(n15959), .QN(g22105) );
  NAND2X0 U16531 ( .IN1(n4289), .IN2(n15838), .QN(n15959) );
  NAND2X0 U16532 ( .IN1(n15839), .IN2(g846), .QN(n15958) );
  NAND2X0 U16533 ( .IN1(n15960), .IN2(n15961), .QN(g22104) );
  NAND2X0 U16534 ( .IN1(n15805), .IN2(n4567), .QN(n15961) );
  INVX0 U16535 ( .INP(n15962), .ZN(n15960) );
  NOR2X0 U16536 ( .IN1(n15805), .IN2(n8821), .QN(n15962) );
  NAND2X0 U16537 ( .IN1(n15963), .IN2(n15964), .QN(g22103) );
  NAND2X0 U16538 ( .IN1(test_so12), .IN2(n15935), .QN(n15964) );
  NAND2X0 U16539 ( .IN1(n15934), .IN2(n10928), .QN(n15963) );
  INVX0 U16540 ( .INP(n12367), .ZN(n10928) );
  NAND2X0 U16541 ( .IN1(n15965), .IN2(n15966), .QN(n12367) );
  NAND2X0 U16542 ( .IN1(n8890), .IN2(g6313), .QN(n15966) );
  NOR2X0 U16543 ( .IN1(n15967), .IN2(n15968), .QN(n15965) );
  NOR2X0 U16544 ( .IN1(n4369), .IN2(g171), .QN(n15968) );
  NOR2X0 U16545 ( .IN1(n4318), .IN2(g172), .QN(n15967) );
  NAND2X0 U16546 ( .IN1(n15969), .IN2(n15970), .QN(g22102) );
  NAND2X0 U16547 ( .IN1(n15928), .IN2(g161), .QN(n15970) );
  INVX0 U16548 ( .INP(n15888), .ZN(n15928) );
  NAND2X0 U16549 ( .IN1(n11093), .IN2(n15888), .QN(n15969) );
  NAND2X0 U16550 ( .IN1(n15971), .IN2(n15972), .QN(g22101) );
  NAND2X0 U16551 ( .IN1(n4290), .IN2(n15845), .QN(n15972) );
  NAND2X0 U16552 ( .IN1(n15220), .IN2(g156), .QN(n15971) );
  NAND2X0 U16553 ( .IN1(n15973), .IN2(n15974), .QN(g22100) );
  NAND2X0 U16554 ( .IN1(n15934), .IN2(n4380), .QN(n15974) );
  NAND2X0 U16555 ( .IN1(n15935), .IN2(g130), .QN(n15973) );
  NAND2X0 U16556 ( .IN1(n15975), .IN2(n15976), .QN(g22099) );
  NAND2X0 U16557 ( .IN1(n15789), .IN2(n4555), .QN(n15976) );
  NAND2X0 U16558 ( .IN1(n15790), .IN2(g2227), .QN(n15975) );
  NAND2X0 U16559 ( .IN1(n15977), .IN2(n15978), .QN(g22098) );
  NAND2X0 U16560 ( .IN1(test_so74), .IN2(n15784), .QN(n15978) );
  INVX0 U16561 ( .INP(n15775), .ZN(n15784) );
  NAND2X0 U16562 ( .IN1(n15775), .IN2(n4325), .QN(n15977) );
  NAND2X0 U16563 ( .IN1(n15979), .IN2(n15980), .QN(g22097) );
  NAND2X0 U16564 ( .IN1(n4389), .IN2(n15769), .QN(n15980) );
  NAND2X0 U16565 ( .IN1(n15214), .IN2(g2220), .QN(n15979) );
  NAND2X0 U16566 ( .IN1(n15981), .IN2(n15982), .QN(g22092) );
  NAND2X0 U16567 ( .IN1(n15830), .IN2(n4565), .QN(n15982) );
  NAND2X0 U16568 ( .IN1(n15829), .IN2(g1536), .QN(n15981) );
  NAND2X0 U16569 ( .IN1(n15983), .IN2(n15984), .QN(g22091) );
  NAND2X0 U16570 ( .IN1(n15799), .IN2(n4557), .QN(n15984) );
  INVX0 U16571 ( .INP(n15985), .ZN(n15983) );
  NOR2X0 U16572 ( .IN1(n15799), .IN2(n9174), .QN(n15985) );
  NAND2X0 U16573 ( .IN1(n15986), .IN2(n15987), .QN(g22090) );
  NAND2X0 U16574 ( .IN1(n4326), .IN2(n15781), .QN(n15987) );
  NAND2X0 U16575 ( .IN1(n15216), .IN2(g1529), .QN(n15986) );
  NAND2X0 U16576 ( .IN1(n15988), .IN2(n15989), .QN(g22089) );
  NAND2X0 U16577 ( .IN1(n4289), .IN2(n15879), .QN(n15989) );
  NAND2X0 U16578 ( .IN1(n15880), .IN2(g845), .QN(n15988) );
  NAND2X0 U16579 ( .IN1(n15990), .IN2(n15991), .QN(g22088) );
  NAND2X0 U16580 ( .IN1(n15838), .IN2(n4567), .QN(n15991) );
  NAND2X0 U16581 ( .IN1(n15839), .IN2(g843), .QN(n15990) );
  NAND2X0 U16582 ( .IN1(n15992), .IN2(n15993), .QN(g22087) );
  NAND2X0 U16583 ( .IN1(n15805), .IN2(n4559), .QN(n15993) );
  INVX0 U16584 ( .INP(n15994), .ZN(n15992) );
  NOR2X0 U16585 ( .IN1(n15805), .IN2(n8822), .QN(n15994) );
  NAND2X0 U16586 ( .IN1(n15995), .IN2(n15996), .QN(g22081) );
  INVX0 U16587 ( .INP(n15997), .ZN(n15996) );
  NOR2X0 U16588 ( .IN1(n15934), .IN2(n8792), .QN(n15997) );
  NAND2X0 U16589 ( .IN1(n15934), .IN2(n11093), .QN(n15995) );
  INVX0 U16590 ( .INP(n12342), .ZN(n11093) );
  NAND2X0 U16591 ( .IN1(n15998), .IN2(n15999), .QN(n12342) );
  NAND2X0 U16592 ( .IN1(n8887), .IN2(g6313), .QN(n15999) );
  NOR2X0 U16593 ( .IN1(n16000), .IN2(n16001), .QN(n15998) );
  NOR2X0 U16594 ( .IN1(n4369), .IN2(g174), .QN(n16001) );
  NOR2X0 U16595 ( .IN1(n4318), .IN2(g175), .QN(n16000) );
  NAND2X0 U16596 ( .IN1(n16002), .IN2(n16003), .QN(g22080) );
  NAND2X0 U16597 ( .IN1(n4290), .IN2(n15888), .QN(n16003) );
  INVX0 U16598 ( .INP(n16004), .ZN(n16002) );
  NOR2X0 U16599 ( .IN1(n15888), .IN2(n9200), .QN(n16004) );
  NAND2X0 U16600 ( .IN1(n16005), .IN2(n16006), .QN(g22079) );
  NAND2X0 U16601 ( .IN1(n4569), .IN2(n15845), .QN(n16006) );
  NAND2X0 U16602 ( .IN1(n15220), .IN2(g153), .QN(n16005) );
  NAND2X0 U16603 ( .IN1(n16007), .IN2(n16008), .QN(g22078) );
  NAND2X0 U16604 ( .IN1(n15789), .IN2(n4325), .QN(n16008) );
  NAND2X0 U16605 ( .IN1(n15790), .IN2(g2224), .QN(n16007) );
  NAND2X0 U16606 ( .IN1(n16009), .IN2(n16010), .QN(g22077) );
  NAND2X0 U16607 ( .IN1(n15775), .IN2(n4389), .QN(n16010) );
  INVX0 U16608 ( .INP(n16011), .ZN(n16009) );
  NOR2X0 U16609 ( .IN1(n15775), .IN2(n9163), .QN(n16011) );
  NAND2X0 U16610 ( .IN1(n16012), .IN2(n16013), .QN(g22076) );
  NAND2X0 U16611 ( .IN1(n4319), .IN2(n15769), .QN(n16013) );
  NAND2X0 U16612 ( .IN1(n15214), .IN2(g2217), .QN(n16012) );
  INVX0 U16613 ( .INP(n15769), .ZN(n15214) );
  NOR2X0 U16614 ( .IN1(n4367), .IN2(n8988), .QN(n15769) );
  NAND2X0 U16615 ( .IN1(n16014), .IN2(n16015), .QN(g22075) );
  NAND2X0 U16616 ( .IN1(n15830), .IN2(n4557), .QN(n16015) );
  NAND2X0 U16617 ( .IN1(n15829), .IN2(g1533), .QN(n16014) );
  NAND2X0 U16618 ( .IN1(n16016), .IN2(n16017), .QN(g22074) );
  NAND2X0 U16619 ( .IN1(n15799), .IN2(n4326), .QN(n16017) );
  INVX0 U16620 ( .INP(n16018), .ZN(n16016) );
  NOR2X0 U16621 ( .IN1(n15799), .IN2(n9176), .QN(n16018) );
  NAND2X0 U16622 ( .IN1(n16019), .IN2(n16020), .QN(g22073) );
  NAND2X0 U16623 ( .IN1(n4390), .IN2(n15781), .QN(n16020) );
  NAND2X0 U16624 ( .IN1(n15216), .IN2(g1526), .QN(n16019) );
  NAND2X0 U16625 ( .IN1(n16021), .IN2(n16022), .QN(g22068) );
  NAND2X0 U16626 ( .IN1(n15879), .IN2(n4567), .QN(n16022) );
  NAND2X0 U16627 ( .IN1(n15880), .IN2(g842), .QN(n16021) );
  NAND2X0 U16628 ( .IN1(n16023), .IN2(n16024), .QN(g22067) );
  NAND2X0 U16629 ( .IN1(n15838), .IN2(n4559), .QN(n16024) );
  NAND2X0 U16630 ( .IN1(n15839), .IN2(g840), .QN(n16023) );
  NAND2X0 U16631 ( .IN1(n16025), .IN2(n16026), .QN(g22066) );
  NAND2X0 U16632 ( .IN1(n4327), .IN2(n15805), .QN(n16026) );
  INVX0 U16633 ( .INP(n16027), .ZN(n16025) );
  NOR2X0 U16634 ( .IN1(n15805), .IN2(n8823), .QN(n16027) );
  NAND2X0 U16635 ( .IN1(n16028), .IN2(n16029), .QN(g22065) );
  NAND2X0 U16636 ( .IN1(n4290), .IN2(n15934), .QN(n16029) );
  NAND2X0 U16637 ( .IN1(n15935), .IN2(g157), .QN(n16028) );
  NAND2X0 U16638 ( .IN1(n16030), .IN2(n16031), .QN(g22064) );
  NAND2X0 U16639 ( .IN1(n15888), .IN2(n4569), .QN(n16031) );
  INVX0 U16640 ( .INP(n16032), .ZN(n16030) );
  NOR2X0 U16641 ( .IN1(n15888), .IN2(n9202), .QN(n16032) );
  NAND2X0 U16642 ( .IN1(n16033), .IN2(n16034), .QN(g22063) );
  NAND2X0 U16643 ( .IN1(n4561), .IN2(n15845), .QN(n16034) );
  NAND2X0 U16644 ( .IN1(n15220), .IN2(g150), .QN(n16033) );
  NAND2X0 U16645 ( .IN1(n16035), .IN2(n16036), .QN(g22061) );
  NAND2X0 U16646 ( .IN1(n15789), .IN2(n4389), .QN(n16036) );
  NAND2X0 U16647 ( .IN1(n15790), .IN2(g2221), .QN(n16035) );
  NAND2X0 U16648 ( .IN1(n16037), .IN2(n16038), .QN(g22060) );
  NAND2X0 U16649 ( .IN1(n15775), .IN2(n4319), .QN(n16038) );
  INVX0 U16650 ( .INP(n16039), .ZN(n16037) );
  NOR2X0 U16651 ( .IN1(n15775), .IN2(n9165), .QN(n16039) );
  NOR2X0 U16652 ( .IN1(n9278), .IN2(n8988), .QN(n15775) );
  NAND2X0 U16653 ( .IN1(n16040), .IN2(n16041), .QN(g22059) );
  NAND2X0 U16654 ( .IN1(n15830), .IN2(n4326), .QN(n16041) );
  NAND2X0 U16655 ( .IN1(n15829), .IN2(g1530), .QN(n16040) );
  NAND2X0 U16656 ( .IN1(n16042), .IN2(n16043), .QN(g22058) );
  NAND2X0 U16657 ( .IN1(n15799), .IN2(n4390), .QN(n16043) );
  INVX0 U16658 ( .INP(n16044), .ZN(n16042) );
  NOR2X0 U16659 ( .IN1(n15799), .IN2(n9178), .QN(n16044) );
  NAND2X0 U16660 ( .IN1(n16045), .IN2(n16046), .QN(g22057) );
  NAND2X0 U16661 ( .IN1(n4320), .IN2(n15781), .QN(n16046) );
  NAND2X0 U16662 ( .IN1(n15216), .IN2(g1523), .QN(n16045) );
  INVX0 U16663 ( .INP(n15781), .ZN(n15216) );
  NOR2X0 U16664 ( .IN1(n4368), .IN2(n8989), .QN(n15781) );
  NAND2X0 U16665 ( .IN1(n16047), .IN2(n16048), .QN(g22056) );
  NAND2X0 U16666 ( .IN1(test_so32), .IN2(n15880), .QN(n16048) );
  NAND2X0 U16667 ( .IN1(n15879), .IN2(n4559), .QN(n16047) );
  NAND2X0 U16668 ( .IN1(n16049), .IN2(n16050), .QN(g22055) );
  NAND2X0 U16669 ( .IN1(n4327), .IN2(n15838), .QN(n16050) );
  NAND2X0 U16670 ( .IN1(n15839), .IN2(g837), .QN(n16049) );
  NAND2X0 U16671 ( .IN1(n16051), .IN2(n16052), .QN(g22054) );
  NAND2X0 U16672 ( .IN1(n15805), .IN2(n4391), .QN(n16052) );
  INVX0 U16673 ( .INP(n16053), .ZN(n16051) );
  NOR2X0 U16674 ( .IN1(n15805), .IN2(n8824), .QN(n16053) );
  NAND2X0 U16675 ( .IN1(n16054), .IN2(n16055), .QN(g22049) );
  NAND2X0 U16676 ( .IN1(n15934), .IN2(n4569), .QN(n16055) );
  NAND2X0 U16677 ( .IN1(n15935), .IN2(g154), .QN(n16054) );
  NAND2X0 U16678 ( .IN1(n16056), .IN2(n16057), .QN(g22048) );
  NAND2X0 U16679 ( .IN1(n15888), .IN2(n4561), .QN(n16057) );
  INVX0 U16680 ( .INP(n16058), .ZN(n16056) );
  NOR2X0 U16681 ( .IN1(n15888), .IN2(n9204), .QN(n16058) );
  NAND2X0 U16682 ( .IN1(n16059), .IN2(n16060), .QN(g22047) );
  NAND2X0 U16683 ( .IN1(n4328), .IN2(n15845), .QN(n16060) );
  NAND2X0 U16684 ( .IN1(n15220), .IN2(g147), .QN(n16059) );
  NAND2X0 U16685 ( .IN1(n16061), .IN2(n16062), .QN(g22045) );
  NAND2X0 U16686 ( .IN1(n15789), .IN2(n4319), .QN(n16062) );
  NAND2X0 U16687 ( .IN1(n15790), .IN2(g2218), .QN(n16061) );
  INVX0 U16688 ( .INP(n15789), .ZN(n15790) );
  NOR2X0 U16689 ( .IN1(n4324), .IN2(n8988), .QN(n15789) );
  NAND2X0 U16690 ( .IN1(n16063), .IN2(n16064), .QN(g22044) );
  NAND2X0 U16691 ( .IN1(n15830), .IN2(n4390), .QN(n16064) );
  NAND2X0 U16692 ( .IN1(n15829), .IN2(g1527), .QN(n16063) );
  NAND2X0 U16693 ( .IN1(n16065), .IN2(n16066), .QN(g22043) );
  NAND2X0 U16694 ( .IN1(n15799), .IN2(n4320), .QN(n16066) );
  INVX0 U16695 ( .INP(n16067), .ZN(n16065) );
  NOR2X0 U16696 ( .IN1(n15799), .IN2(n9180), .QN(n16067) );
  NOR2X0 U16697 ( .IN1(n4515), .IN2(n8989), .QN(n15799) );
  NAND2X0 U16698 ( .IN1(n16068), .IN2(n16069), .QN(g22042) );
  NAND2X0 U16699 ( .IN1(n4327), .IN2(n15879), .QN(n16069) );
  NAND2X0 U16700 ( .IN1(n15880), .IN2(g836), .QN(n16068) );
  NAND2X0 U16701 ( .IN1(n16070), .IN2(n16071), .QN(g22041) );
  NAND2X0 U16702 ( .IN1(n15838), .IN2(n4391), .QN(n16071) );
  NAND2X0 U16703 ( .IN1(n15839), .IN2(g834), .QN(n16070) );
  NAND2X0 U16704 ( .IN1(n16072), .IN2(n16073), .QN(g22040) );
  NAND2X0 U16705 ( .IN1(n4321), .IN2(n15805), .QN(n16073) );
  INVX0 U16706 ( .INP(n16074), .ZN(n16072) );
  NOR2X0 U16707 ( .IN1(n15805), .IN2(n8825), .QN(n16074) );
  NOR2X0 U16708 ( .IN1(n9279), .IN2(n8990), .QN(n15805) );
  NAND2X0 U16709 ( .IN1(n16075), .IN2(n16076), .QN(g22039) );
  NAND2X0 U16710 ( .IN1(n15934), .IN2(n4561), .QN(n16076) );
  NAND2X0 U16711 ( .IN1(n15935), .IN2(g151), .QN(n16075) );
  NAND2X0 U16712 ( .IN1(n16077), .IN2(n16078), .QN(g22038) );
  NAND2X0 U16713 ( .IN1(n4328), .IN2(n15888), .QN(n16078) );
  INVX0 U16714 ( .INP(n16079), .ZN(n16077) );
  NOR2X0 U16715 ( .IN1(n15888), .IN2(n9206), .QN(n16079) );
  NAND2X0 U16716 ( .IN1(n16080), .IN2(n16081), .QN(g22037) );
  NAND2X0 U16717 ( .IN1(test_so11), .IN2(n15220), .QN(n16081) );
  NAND2X0 U16718 ( .IN1(n4392), .IN2(n15845), .QN(n16080) );
  NAND2X0 U16719 ( .IN1(n16082), .IN2(n16083), .QN(g22035) );
  NAND2X0 U16720 ( .IN1(n15830), .IN2(n4320), .QN(n16083) );
  NAND2X0 U16721 ( .IN1(n15829), .IN2(g1524), .QN(n16082) );
  INVX0 U16722 ( .INP(n15830), .ZN(n15829) );
  NOR2X0 U16723 ( .IN1(n4317), .IN2(n8989), .QN(n15830) );
  NAND2X0 U16724 ( .IN1(n16084), .IN2(n16085), .QN(g22034) );
  NAND2X0 U16725 ( .IN1(n15879), .IN2(n4391), .QN(n16085) );
  NAND2X0 U16726 ( .IN1(n15880), .IN2(g833), .QN(n16084) );
  NAND2X0 U16727 ( .IN1(n16086), .IN2(n16087), .QN(g22033) );
  NAND2X0 U16728 ( .IN1(n4321), .IN2(n15838), .QN(n16087) );
  NAND2X0 U16729 ( .IN1(n15839), .IN2(g831), .QN(n16086) );
  INVX0 U16730 ( .INP(n15838), .ZN(n15839) );
  NOR2X0 U16731 ( .IN1(n4312), .IN2(n8990), .QN(n15838) );
  NAND2X0 U16732 ( .IN1(n16088), .IN2(n16089), .QN(g22032) );
  NAND2X0 U16733 ( .IN1(n4328), .IN2(n15934), .QN(n16089) );
  NAND2X0 U16734 ( .IN1(n15935), .IN2(g148), .QN(n16088) );
  NAND2X0 U16735 ( .IN1(n16090), .IN2(n16091), .QN(g22031) );
  NAND2X0 U16736 ( .IN1(n15888), .IN2(n4392), .QN(n16091) );
  INVX0 U16737 ( .INP(n16092), .ZN(n16090) );
  NOR2X0 U16738 ( .IN1(n15888), .IN2(n9208), .QN(n16092) );
  NAND2X0 U16739 ( .IN1(n16093), .IN2(n16094), .QN(g22030) );
  NAND2X0 U16740 ( .IN1(n4322), .IN2(n15845), .QN(n16094) );
  NAND2X0 U16741 ( .IN1(n15220), .IN2(g141), .QN(n16093) );
  INVX0 U16742 ( .INP(n15845), .ZN(n15220) );
  NOR2X0 U16743 ( .IN1(n4369), .IN2(n8991), .QN(n15845) );
  NAND2X0 U16744 ( .IN1(n16095), .IN2(n16096), .QN(g22029) );
  NAND2X0 U16745 ( .IN1(n4321), .IN2(n15879), .QN(n16096) );
  NAND2X0 U16746 ( .IN1(n15880), .IN2(g830), .QN(n16095) );
  INVX0 U16747 ( .INP(n15879), .ZN(n15880) );
  NOR2X0 U16748 ( .IN1(n4323), .IN2(n8990), .QN(n15879) );
  NAND2X0 U16749 ( .IN1(n16097), .IN2(n16098), .QN(g22028) );
  NAND2X0 U16750 ( .IN1(n15934), .IN2(n4392), .QN(n16098) );
  NAND2X0 U16751 ( .IN1(n15935), .IN2(g145), .QN(n16097) );
  NAND2X0 U16752 ( .IN1(n16099), .IN2(n16100), .QN(g22027) );
  NAND2X0 U16753 ( .IN1(n4322), .IN2(n15888), .QN(n16100) );
  INVX0 U16754 ( .INP(n16101), .ZN(n16099) );
  NOR2X0 U16755 ( .IN1(n15888), .IN2(n9210), .QN(n16101) );
  NOR2X0 U16756 ( .IN1(n4512), .IN2(n8991), .QN(n15888) );
  NOR2X0 U16757 ( .IN1(n9867), .IN2(n16102), .QN(g22026) );
  XNOR2X1 U16758 ( .IN1(g2888), .IN2(n15419), .Q(n16102) );
  NOR2X0 U16759 ( .IN1(n4423), .IN2(n4330), .QN(n15419) );
  NAND2X0 U16760 ( .IN1(n16829), .IN2(n9872), .QN(n9867) );
  NAND2X0 U16761 ( .IN1(n16103), .IN2(n16104), .QN(n9872) );
  NOR2X0 U16762 ( .IN1(n16105), .IN2(n16106), .QN(n16104) );
  NAND2X0 U16763 ( .IN1(n4182), .IN2(g2908), .QN(n16106) );
  NAND2X0 U16764 ( .IN1(g2950), .IN2(g2888), .QN(n16105) );
  NOR2X0 U16765 ( .IN1(g2896), .IN2(n16107), .QN(n16103) );
  NAND2X0 U16766 ( .IN1(n4330), .IN2(n4291), .QN(n16107) );
  NAND2X0 U16767 ( .IN1(n16108), .IN2(n16109), .QN(g22025) );
  NAND2X0 U16768 ( .IN1(n4322), .IN2(n15934), .QN(n16109) );
  NAND2X0 U16769 ( .IN1(n15935), .IN2(g142), .QN(n16108) );
  INVX0 U16770 ( .INP(n15934), .ZN(n15935) );
  NOR2X0 U16771 ( .IN1(n4318), .IN2(n8991), .QN(n15934) );
  NOR2X0 U16772 ( .IN1(n16110), .IN2(n16111), .QN(g21974) );
  NAND2X0 U16773 ( .IN1(n15427), .IN2(n13918), .QN(n16111) );
  NAND2X0 U16774 ( .IN1(n16112), .IN2(n16113), .QN(n15427) );
  NOR2X0 U16775 ( .IN1(n4472), .IN2(n4398), .QN(n16112) );
  NOR2X0 U16776 ( .IN1(n16114), .IN2(g2707), .QN(n16110) );
  NOR2X0 U16777 ( .IN1(n4398), .IN2(n16115), .QN(n16114) );
  NOR2X0 U16778 ( .IN1(n16116), .IN2(n16117), .QN(g21972) );
  NAND2X0 U16779 ( .IN1(n15434), .IN2(n13126), .QN(n16117) );
  INVX0 U16780 ( .INP(n15432), .ZN(n15434) );
  NOR2X0 U16781 ( .IN1(n16118), .IN2(n16119), .QN(n15432) );
  NAND2X0 U16782 ( .IN1(g2013), .IN2(g2020), .QN(n16118) );
  NOR2X0 U16783 ( .IN1(n16120), .IN2(g2013), .QN(n16116) );
  NOR2X0 U16784 ( .IN1(n4400), .IN2(n16119), .QN(n16120) );
  NAND2X0 U16785 ( .IN1(n16121), .IN2(n16122), .QN(g21970) );
  NAND2X0 U16786 ( .IN1(test_so87), .IN2(n4463), .QN(n16122) );
  NAND2X0 U16787 ( .IN1(n13166), .IN2(g2560), .QN(n16121) );
  NAND2X0 U16788 ( .IN1(n16123), .IN2(n16124), .QN(n13166) );
  NAND2X0 U16789 ( .IN1(g5555), .IN2(g2513), .QN(n16124) );
  NOR2X0 U16790 ( .IN1(n16125), .IN2(n16126), .QN(n16123) );
  NOR2X0 U16791 ( .IN1(n8700), .IN2(n12443), .QN(n16126) );
  INVX0 U16792 ( .INP(g7264), .ZN(n12443) );
  NOR2X0 U16793 ( .IN1(n8711), .IN2(n13976), .QN(n16125) );
  INVX0 U16794 ( .INP(n4606), .ZN(n13976) );
  NOR2X0 U16795 ( .IN1(n16127), .IN2(n16128), .QN(g21969) );
  NAND2X0 U16796 ( .IN1(n15440), .IN2(n13134), .QN(n16128) );
  INVX0 U16797 ( .INP(n15438), .ZN(n15440) );
  NOR2X0 U16798 ( .IN1(n16129), .IN2(n16130), .QN(n15438) );
  NAND2X0 U16799 ( .IN1(g1319), .IN2(g1326), .QN(n16129) );
  NOR2X0 U16800 ( .IN1(n16131), .IN2(g1319), .QN(n16127) );
  NOR2X0 U16801 ( .IN1(n4402), .IN2(n16130), .QN(n16131) );
  NAND2X0 U16802 ( .IN1(n16132), .IN2(n16133), .QN(g21882) );
  NAND2X0 U16803 ( .IN1(n4351), .IN2(g2878), .QN(n16133) );
  NAND2X0 U16804 ( .IN1(n16134), .IN2(g2879), .QN(n16132) );
  NAND2X0 U16805 ( .IN1(n16135), .IN2(n16136), .QN(g21880) );
  NAND2X0 U16806 ( .IN1(n4351), .IN2(g2877), .QN(n16136) );
  NAND2X0 U16807 ( .IN1(n16137), .IN2(g2879), .QN(n16135) );
  NAND2X0 U16808 ( .IN1(n16138), .IN2(n16139), .QN(g21878) );
  NAND2X0 U16809 ( .IN1(test_so4), .IN2(g2879), .QN(n16139) );
  NAND2X0 U16810 ( .IN1(n16134), .IN2(n4351), .QN(n16138) );
  XOR2X1 U16811 ( .IN1(n16140), .IN2(n9723), .Q(n16134) );
  XNOR2X1 U16812 ( .IN1(n16141), .IN2(n16142), .Q(n9723) );
  XOR2X1 U16813 ( .IN1(n16143), .IN2(n16144), .Q(n16142) );
  XNOR2X1 U16814 ( .IN1(g2969), .IN2(n9244), .Q(n16144) );
  XNOR2X1 U16815 ( .IN1(test_so2), .IN2(g2981), .Q(n16143) );
  XOR2X1 U16816 ( .IN1(n16145), .IN2(n16146), .Q(n16141) );
  XNOR2X1 U16817 ( .IN1(g2972), .IN2(n9242), .Q(n16146) );
  XNOR2X1 U16818 ( .IN1(n9240), .IN2(n9241), .Q(n16145) );
  NAND2X0 U16819 ( .IN1(n16147), .IN2(n16148), .QN(g21851) );
  NAND2X0 U16820 ( .IN1(g499), .IN2(g544), .QN(n16148) );
  NAND2X0 U16821 ( .IN1(n16149), .IN2(n4541), .QN(n16147) );
  NOR2X0 U16822 ( .IN1(n8375), .IN2(n13002), .QN(n16149) );
  NAND2X0 U16823 ( .IN1(n16150), .IN2(n16151), .QN(g21346) );
  NAND2X0 U16824 ( .IN1(n16833), .IN2(DFF_328_n1), .QN(n16151) );
  NAND2X0 U16825 ( .IN1(n16152), .IN2(n8056), .QN(n16150) );
  NOR2X0 U16826 ( .IN1(n8699), .IN2(g6447), .QN(n16152) );
  NAND2X0 U16827 ( .IN1(n16153), .IN2(n16154), .QN(g21094) );
  NAND2X0 U16828 ( .IN1(test_so94), .IN2(n14691), .QN(n16154) );
  NAND2X0 U16829 ( .IN1(n14693), .IN2(n4393), .QN(n16153) );
  NAND2X0 U16830 ( .IN1(n16155), .IN2(n16156), .QN(g21082) );
  NAND2X0 U16831 ( .IN1(n14697), .IN2(n4393), .QN(n16156) );
  INVX0 U16832 ( .INP(n16157), .ZN(n16155) );
  NOR2X0 U16833 ( .IN1(n14697), .IN2(n9042), .QN(n16157) );
  NAND2X0 U16834 ( .IN1(n16158), .IN2(n16159), .QN(g21081) );
  NAND2X0 U16835 ( .IN1(n14693), .IN2(n4471), .QN(n16159) );
  NAND2X0 U16836 ( .IN1(n14691), .IN2(g2793), .QN(n16158) );
  NAND2X0 U16837 ( .IN1(n16160), .IN2(n16161), .QN(g21080) );
  NAND2X0 U16838 ( .IN1(n14702), .IN2(n9284), .QN(n16161) );
  NAND2X0 U16839 ( .IN1(n14700), .IN2(g2102), .QN(n16160) );
  NAND2X0 U16840 ( .IN1(n16162), .IN2(n16163), .QN(g21075) );
  NAND2X0 U16841 ( .IN1(n14705), .IN2(n4393), .QN(n16163) );
  NAND2X0 U16842 ( .IN1(n10624), .IN2(g2797), .QN(n16162) );
  NAND2X0 U16843 ( .IN1(n16164), .IN2(n16165), .QN(g21074) );
  NAND2X0 U16844 ( .IN1(n14697), .IN2(n4471), .QN(n16165) );
  INVX0 U16845 ( .INP(n16166), .ZN(n16164) );
  NOR2X0 U16846 ( .IN1(n14697), .IN2(n9044), .QN(n16166) );
  NAND2X0 U16847 ( .IN1(n16167), .IN2(n16168), .QN(g21073) );
  NAND2X0 U16848 ( .IN1(n14693), .IN2(n9282), .QN(n16168) );
  NAND2X0 U16849 ( .IN1(n14691), .IN2(g2790), .QN(n16167) );
  NAND2X0 U16850 ( .IN1(n16169), .IN2(n16170), .QN(g21072) );
  NAND2X0 U16851 ( .IN1(n14778), .IN2(n9284), .QN(n16170) );
  INVX0 U16852 ( .INP(n16171), .ZN(n16169) );
  NOR2X0 U16853 ( .IN1(n14778), .IN2(n9061), .QN(n16171) );
  NAND2X0 U16854 ( .IN1(n16172), .IN2(n16173), .QN(g21071) );
  NAND2X0 U16855 ( .IN1(n14702), .IN2(n4473), .QN(n16173) );
  NAND2X0 U16856 ( .IN1(n14700), .IN2(g2099), .QN(n16172) );
  NAND2X0 U16857 ( .IN1(n16174), .IN2(n16175), .QN(g21070) );
  NAND2X0 U16858 ( .IN1(n14784), .IN2(n4395), .QN(n16175) );
  NAND2X0 U16859 ( .IN1(n14782), .IN2(g1408), .QN(n16174) );
  NAND2X0 U16860 ( .IN1(n16176), .IN2(n16177), .QN(g21063) );
  NAND2X0 U16861 ( .IN1(n16178), .IN2(g2805), .QN(n16177) );
  INVX0 U16862 ( .INP(n15752), .ZN(n16178) );
  NAND2X0 U16863 ( .IN1(n15752), .IN2(n10091), .QN(n16176) );
  NAND2X0 U16864 ( .IN1(n16179), .IN2(n16180), .QN(g21062) );
  NAND2X0 U16865 ( .IN1(n14705), .IN2(n4471), .QN(n16180) );
  NAND2X0 U16866 ( .IN1(n10624), .IN2(g2794), .QN(n16179) );
  NAND2X0 U16867 ( .IN1(n16181), .IN2(n16182), .QN(g21061) );
  NAND2X0 U16868 ( .IN1(n14697), .IN2(n9282), .QN(n16182) );
  INVX0 U16869 ( .INP(n16183), .ZN(n16181) );
  NOR2X0 U16870 ( .IN1(n14697), .IN2(n9046), .QN(n16183) );
  NAND2X0 U16871 ( .IN1(n16184), .IN2(n16185), .QN(g21060) );
  NAND2X0 U16872 ( .IN1(n14693), .IN2(n4407), .QN(n16185) );
  NAND2X0 U16873 ( .IN1(n14691), .IN2(g2787), .QN(n16184) );
  NAND2X0 U16874 ( .IN1(n16186), .IN2(n16187), .QN(g21056) );
  NAND2X0 U16875 ( .IN1(n14787), .IN2(n9284), .QN(n16187) );
  NAND2X0 U16876 ( .IN1(n10652), .IN2(g2103), .QN(n16186) );
  NAND2X0 U16877 ( .IN1(n16188), .IN2(n16189), .QN(g21055) );
  NAND2X0 U16878 ( .IN1(n14778), .IN2(n4473), .QN(n16189) );
  INVX0 U16879 ( .INP(n16190), .ZN(n16188) );
  NOR2X0 U16880 ( .IN1(n14778), .IN2(n9063), .QN(n16190) );
  NAND2X0 U16881 ( .IN1(n16191), .IN2(n16192), .QN(g21054) );
  NAND2X0 U16882 ( .IN1(n4468), .IN2(n14702), .QN(n16192) );
  NAND2X0 U16883 ( .IN1(n14700), .IN2(g2096), .QN(n16191) );
  NAND2X0 U16884 ( .IN1(n16193), .IN2(n16194), .QN(g21053) );
  NAND2X0 U16885 ( .IN1(n14861), .IN2(n4395), .QN(n16194) );
  INVX0 U16886 ( .INP(n16195), .ZN(n16193) );
  NOR2X0 U16887 ( .IN1(n14861), .IN2(n9080), .QN(n16195) );
  NAND2X0 U16888 ( .IN1(n16196), .IN2(n16197), .QN(g21052) );
  NAND2X0 U16889 ( .IN1(n14784), .IN2(n4475), .QN(n16197) );
  NAND2X0 U16890 ( .IN1(n14782), .IN2(g1405), .QN(n16196) );
  NAND2X0 U16891 ( .IN1(n16198), .IN2(n16199), .QN(g21051) );
  NAND2X0 U16892 ( .IN1(n14866), .IN2(n4396), .QN(n16199) );
  NAND2X0 U16893 ( .IN1(n14864), .IN2(g722), .QN(n16198) );
  NAND2X0 U16894 ( .IN1(n16200), .IN2(n16201), .QN(g21047) );
  NAND2X0 U16895 ( .IN1(n10617), .IN2(n10091), .QN(n16201) );
  INVX0 U16896 ( .INP(n16202), .ZN(n16200) );
  NOR2X0 U16897 ( .IN1(n10617), .IN2(n8837), .QN(n16202) );
  NAND2X0 U16898 ( .IN1(n16203), .IN2(n16204), .QN(g21046) );
  INVX0 U16899 ( .INP(n16205), .ZN(n16204) );
  NOR2X0 U16900 ( .IN1(n15752), .IN2(n8896), .QN(n16205) );
  NAND2X0 U16901 ( .IN1(n15752), .IN2(n10100), .QN(n16203) );
  NOR2X0 U16902 ( .IN1(n4292), .IN2(n9031), .QN(n15752) );
  NAND2X0 U16903 ( .IN1(n16206), .IN2(n16207), .QN(g21045) );
  NAND2X0 U16904 ( .IN1(n14705), .IN2(n9282), .QN(n16207) );
  NAND2X0 U16905 ( .IN1(n10624), .IN2(g2791), .QN(n16206) );
  NAND2X0 U16906 ( .IN1(n16208), .IN2(n16209), .QN(g21044) );
  NAND2X0 U16907 ( .IN1(n14697), .IN2(n4407), .QN(n16209) );
  INVX0 U16908 ( .INP(n16210), .ZN(n16208) );
  NOR2X0 U16909 ( .IN1(n14697), .IN2(n9048), .QN(n16210) );
  NAND2X0 U16910 ( .IN1(n16211), .IN2(n16212), .QN(g21043) );
  NAND2X0 U16911 ( .IN1(n4397), .IN2(n14693), .QN(n16212) );
  NAND2X0 U16912 ( .IN1(n14691), .IN2(g2784), .QN(n16211) );
  NAND2X0 U16913 ( .IN1(n16213), .IN2(n16214), .QN(g21042) );
  NAND2X0 U16914 ( .IN1(n16215), .IN2(g2111), .QN(n16214) );
  INVX0 U16915 ( .INP(n15755), .ZN(n16215) );
  NAND2X0 U16916 ( .IN1(n15755), .IN2(n10229), .QN(n16213) );
  NAND2X0 U16917 ( .IN1(n16216), .IN2(n16217), .QN(g21041) );
  NAND2X0 U16918 ( .IN1(n14787), .IN2(n4473), .QN(n16217) );
  NAND2X0 U16919 ( .IN1(n10652), .IN2(g2100), .QN(n16216) );
  NAND2X0 U16920 ( .IN1(n16218), .IN2(n16219), .QN(g21040) );
  NAND2X0 U16921 ( .IN1(n4468), .IN2(n14778), .QN(n16219) );
  INVX0 U16922 ( .INP(n16220), .ZN(n16218) );
  NOR2X0 U16923 ( .IN1(n14778), .IN2(n9065), .QN(n16220) );
  NAND2X0 U16924 ( .IN1(n16221), .IN2(n16222), .QN(g21039) );
  NAND2X0 U16925 ( .IN1(n14702), .IN2(n4409), .QN(n16222) );
  NAND2X0 U16926 ( .IN1(n14700), .IN2(g2093), .QN(n16221) );
  NAND2X0 U16927 ( .IN1(n16223), .IN2(n16224), .QN(g21035) );
  NAND2X0 U16928 ( .IN1(n14872), .IN2(n4395), .QN(n16224) );
  NAND2X0 U16929 ( .IN1(n9671), .IN2(g1409), .QN(n16223) );
  NAND2X0 U16930 ( .IN1(n16225), .IN2(n16226), .QN(g21034) );
  NAND2X0 U16931 ( .IN1(n14861), .IN2(n4475), .QN(n16226) );
  INVX0 U16932 ( .INP(n16227), .ZN(n16225) );
  NOR2X0 U16933 ( .IN1(n14861), .IN2(n9082), .QN(n16227) );
  NAND2X0 U16934 ( .IN1(n16228), .IN2(n16229), .QN(g21033) );
  NAND2X0 U16935 ( .IN1(n4469), .IN2(n14784), .QN(n16229) );
  NAND2X0 U16936 ( .IN1(n14782), .IN2(g1402), .QN(n16228) );
  NAND2X0 U16937 ( .IN1(n16230), .IN2(n16231), .QN(g21032) );
  NAND2X0 U16938 ( .IN1(n14948), .IN2(n4396), .QN(n16231) );
  INVX0 U16939 ( .INP(n16232), .ZN(n16230) );
  NOR2X0 U16940 ( .IN1(n14948), .IN2(n9097), .QN(n16232) );
  NAND2X0 U16941 ( .IN1(n16233), .IN2(n16234), .QN(g21031) );
  NAND2X0 U16942 ( .IN1(n14866), .IN2(n4477), .QN(n16234) );
  NAND2X0 U16943 ( .IN1(n14864), .IN2(g719), .QN(n16233) );
  NAND2X0 U16944 ( .IN1(n16235), .IN2(n16236), .QN(g21029) );
  NAND2X0 U16945 ( .IN1(n10622), .IN2(g2806), .QN(n16236) );
  NAND2X0 U16946 ( .IN1(n16237), .IN2(n10091), .QN(n16235) );
  INVX0 U16947 ( .INP(n10628), .ZN(n10091) );
  NAND2X0 U16948 ( .IN1(n16238), .IN2(n16239), .QN(n10628) );
  NAND2X0 U16949 ( .IN1(test_so90), .IN2(g7390), .QN(n16239) );
  NOR2X0 U16950 ( .IN1(n16240), .IN2(n16241), .QN(n16238) );
  NOR2X0 U16951 ( .IN1(n8688), .IN2(n4299), .QN(n16241) );
  NOR2X0 U16952 ( .IN1(n8687), .IN2(n11700), .QN(n16240) );
  INVX0 U16953 ( .INP(g7302), .ZN(n11700) );
  NAND2X0 U16954 ( .IN1(n16242), .IN2(n16243), .QN(g21028) );
  NAND2X0 U16955 ( .IN1(n10617), .IN2(n10100), .QN(n16243) );
  NAND2X0 U16956 ( .IN1(n13918), .IN2(g2804), .QN(n16242) );
  INVX0 U16957 ( .INP(n10617), .ZN(n13918) );
  NAND2X0 U16958 ( .IN1(n16244), .IN2(n16245), .QN(g21027) );
  NAND2X0 U16959 ( .IN1(n14705), .IN2(n4407), .QN(n16245) );
  NAND2X0 U16960 ( .IN1(n10624), .IN2(g2788), .QN(n16244) );
  NAND2X0 U16961 ( .IN1(n16246), .IN2(n16247), .QN(g21026) );
  NAND2X0 U16962 ( .IN1(n4397), .IN2(n14697), .QN(n16247) );
  INVX0 U16963 ( .INP(n16248), .ZN(n16246) );
  NOR2X0 U16964 ( .IN1(n14697), .IN2(n9050), .QN(n16248) );
  NAND2X0 U16965 ( .IN1(n16249), .IN2(n16250), .QN(g21025) );
  NAND2X0 U16966 ( .IN1(test_so93), .IN2(n14691), .QN(n16250) );
  NAND2X0 U16967 ( .IN1(n14693), .IN2(n4408), .QN(n16249) );
  NAND2X0 U16968 ( .IN1(n16251), .IN2(n16252), .QN(g21023) );
  INVX0 U16969 ( .INP(n16253), .ZN(n16252) );
  NOR2X0 U16970 ( .IN1(n14094), .IN2(n8839), .QN(n16253) );
  NAND2X0 U16971 ( .IN1(n14094), .IN2(n10229), .QN(n16251) );
  NAND2X0 U16972 ( .IN1(n16254), .IN2(n16255), .QN(g21022) );
  INVX0 U16973 ( .INP(n16256), .ZN(n16255) );
  NOR2X0 U16974 ( .IN1(n15755), .IN2(n8898), .QN(n16256) );
  NAND2X0 U16975 ( .IN1(n15755), .IN2(n10237), .QN(n16254) );
  NOR2X0 U16976 ( .IN1(n4293), .IN2(n9032), .QN(n15755) );
  NAND2X0 U16977 ( .IN1(n16257), .IN2(n16258), .QN(g21021) );
  NAND2X0 U16978 ( .IN1(n4468), .IN2(n14787), .QN(n16258) );
  NAND2X0 U16979 ( .IN1(n10652), .IN2(g2097), .QN(n16257) );
  NAND2X0 U16980 ( .IN1(n16259), .IN2(n16260), .QN(g21020) );
  NAND2X0 U16981 ( .IN1(n14778), .IN2(n4409), .QN(n16260) );
  INVX0 U16982 ( .INP(n16261), .ZN(n16259) );
  NOR2X0 U16983 ( .IN1(n14778), .IN2(n9067), .QN(n16261) );
  NAND2X0 U16984 ( .IN1(n16262), .IN2(n16263), .QN(g21019) );
  NAND2X0 U16985 ( .IN1(n4399), .IN2(n14702), .QN(n16263) );
  NAND2X0 U16986 ( .IN1(n14700), .IN2(g2090), .QN(n16262) );
  NAND2X0 U16987 ( .IN1(n16264), .IN2(n16265), .QN(g21018) );
  NAND2X0 U16988 ( .IN1(n15760), .IN2(g1417), .QN(n16265) );
  NAND2X0 U16989 ( .IN1(n16266), .IN2(n10372), .QN(n16264) );
  NAND2X0 U16990 ( .IN1(n16267), .IN2(n16268), .QN(g21017) );
  NAND2X0 U16991 ( .IN1(n14872), .IN2(n4475), .QN(n16268) );
  NAND2X0 U16992 ( .IN1(n9671), .IN2(g1406), .QN(n16267) );
  NAND2X0 U16993 ( .IN1(n16269), .IN2(n16270), .QN(g21016) );
  NAND2X0 U16994 ( .IN1(n4469), .IN2(n14861), .QN(n16270) );
  INVX0 U16995 ( .INP(n16271), .ZN(n16269) );
  NOR2X0 U16996 ( .IN1(n14861), .IN2(n9084), .QN(n16271) );
  NAND2X0 U16997 ( .IN1(n16272), .IN2(n16273), .QN(g21015) );
  NAND2X0 U16998 ( .IN1(n14784), .IN2(n4411), .QN(n16273) );
  NAND2X0 U16999 ( .IN1(n14782), .IN2(g1399), .QN(n16272) );
  NAND2X0 U17000 ( .IN1(n16274), .IN2(n16275), .QN(g21011) );
  NAND2X0 U17001 ( .IN1(n14951), .IN2(n4396), .QN(n16275) );
  NAND2X0 U17002 ( .IN1(n9693), .IN2(g723), .QN(n16274) );
  NAND2X0 U17003 ( .IN1(n16276), .IN2(n16277), .QN(g21010) );
  NAND2X0 U17004 ( .IN1(n14948), .IN2(n4477), .QN(n16277) );
  INVX0 U17005 ( .INP(n16278), .ZN(n16276) );
  NOR2X0 U17006 ( .IN1(n14948), .IN2(n9099), .QN(n16278) );
  NAND2X0 U17007 ( .IN1(n16279), .IN2(n16280), .QN(g21009) );
  NAND2X0 U17008 ( .IN1(n14866), .IN2(n9283), .QN(n16280) );
  NAND2X0 U17009 ( .IN1(n14864), .IN2(g716), .QN(n16279) );
  NAND2X0 U17010 ( .IN1(n16281), .IN2(n16282), .QN(g21007) );
  NAND2X0 U17011 ( .IN1(n10622), .IN2(g2803), .QN(n16282) );
  INVX0 U17012 ( .INP(n16237), .ZN(n10622) );
  NAND2X0 U17013 ( .IN1(n16237), .IN2(n10100), .QN(n16281) );
  INVX0 U17014 ( .INP(n10153), .ZN(n10100) );
  NAND2X0 U17015 ( .IN1(n16283), .IN2(n16284), .QN(n10153) );
  NAND2X0 U17016 ( .IN1(g7390), .IN2(g2691), .QN(n16284) );
  NOR2X0 U17017 ( .IN1(n16285), .IN2(n16286), .QN(n16283) );
  NOR2X0 U17018 ( .IN1(n8678), .IN2(n4314), .QN(n16286) );
  NOR2X0 U17019 ( .IN1(n8679), .IN2(n4299), .QN(n16285) );
  NOR2X0 U17020 ( .IN1(n4306), .IN2(n9031), .QN(n16237) );
  NAND2X0 U17021 ( .IN1(n16287), .IN2(n16288), .QN(g21006) );
  NAND2X0 U17022 ( .IN1(n4397), .IN2(n14705), .QN(n16288) );
  NAND2X0 U17023 ( .IN1(n10624), .IN2(g2785), .QN(n16287) );
  NAND2X0 U17024 ( .IN1(n16289), .IN2(n16290), .QN(g21005) );
  NAND2X0 U17025 ( .IN1(n14697), .IN2(n4408), .QN(n16290) );
  INVX0 U17026 ( .INP(n16291), .ZN(n16289) );
  NOR2X0 U17027 ( .IN1(n14697), .IN2(n9052), .QN(n16291) );
  NAND2X0 U17028 ( .IN1(n16292), .IN2(n16293), .QN(g21004) );
  NAND2X0 U17029 ( .IN1(n4419), .IN2(n14693), .QN(n16293) );
  NAND2X0 U17030 ( .IN1(n14691), .IN2(g2778), .QN(n16292) );
  NAND2X0 U17031 ( .IN1(n16294), .IN2(n16295), .QN(g21003) );
  NAND2X0 U17032 ( .IN1(n10650), .IN2(g2112), .QN(n16295) );
  NAND2X0 U17033 ( .IN1(n16296), .IN2(n10229), .QN(n16294) );
  INVX0 U17034 ( .INP(n10266), .ZN(n10229) );
  NAND2X0 U17035 ( .IN1(n16297), .IN2(n16298), .QN(n10266) );
  NAND2X0 U17036 ( .IN1(g1930), .IN2(g1991), .QN(n16298) );
  NOR2X0 U17037 ( .IN1(n16299), .IN2(n16300), .QN(n16297) );
  NOR2X0 U17038 ( .IN1(n8691), .IN2(n4315), .QN(n16300) );
  NOR2X0 U17039 ( .IN1(n8689), .IN2(n15320), .QN(n16299) );
  INVX0 U17040 ( .INP(g7052), .ZN(n15320) );
  NAND2X0 U17041 ( .IN1(n16301), .IN2(n16302), .QN(g21002) );
  NAND2X0 U17042 ( .IN1(n13126), .IN2(g2110), .QN(n16302) );
  INVX0 U17043 ( .INP(n14094), .ZN(n13126) );
  NAND2X0 U17044 ( .IN1(n14094), .IN2(n10237), .QN(n16301) );
  NAND2X0 U17045 ( .IN1(n16303), .IN2(n16304), .QN(g21001) );
  NAND2X0 U17046 ( .IN1(n14787), .IN2(n4409), .QN(n16304) );
  NAND2X0 U17047 ( .IN1(n10652), .IN2(g2094), .QN(n16303) );
  NAND2X0 U17048 ( .IN1(n16305), .IN2(n16306), .QN(g21000) );
  NAND2X0 U17049 ( .IN1(test_so71), .IN2(n14779), .QN(n16306) );
  NAND2X0 U17050 ( .IN1(n4399), .IN2(n14778), .QN(n16305) );
  NAND2X0 U17051 ( .IN1(n16307), .IN2(n16308), .QN(g20999) );
  NAND2X0 U17052 ( .IN1(n14702), .IN2(n4410), .QN(n16308) );
  NAND2X0 U17053 ( .IN1(n14700), .IN2(g2087), .QN(n16307) );
  NAND2X0 U17054 ( .IN1(n16309), .IN2(n16310), .QN(g20997) );
  INVX0 U17055 ( .INP(n16311), .ZN(n16310) );
  NOR2X0 U17056 ( .IN1(n14098), .IN2(n8841), .QN(n16311) );
  NAND2X0 U17057 ( .IN1(n14098), .IN2(n10372), .QN(n16309) );
  NAND2X0 U17058 ( .IN1(n16312), .IN2(n16313), .QN(g20996) );
  NAND2X0 U17059 ( .IN1(test_so51), .IN2(n15760), .QN(n16313) );
  INVX0 U17060 ( .INP(n16266), .ZN(n15760) );
  NAND2X0 U17061 ( .IN1(n16266), .IN2(n10380), .QN(n16312) );
  NOR2X0 U17062 ( .IN1(n4294), .IN2(n9033), .QN(n16266) );
  NAND2X0 U17063 ( .IN1(n16314), .IN2(n16315), .QN(g20995) );
  NAND2X0 U17064 ( .IN1(n4469), .IN2(n14872), .QN(n16315) );
  NAND2X0 U17065 ( .IN1(n9671), .IN2(g1403), .QN(n16314) );
  NAND2X0 U17066 ( .IN1(n16316), .IN2(n16317), .QN(g20994) );
  NAND2X0 U17067 ( .IN1(test_so50), .IN2(n14860), .QN(n16317) );
  NAND2X0 U17068 ( .IN1(n14861), .IN2(n4411), .QN(n16316) );
  NAND2X0 U17069 ( .IN1(n16318), .IN2(n16319), .QN(g20993) );
  NAND2X0 U17070 ( .IN1(n4401), .IN2(n14784), .QN(n16319) );
  NAND2X0 U17071 ( .IN1(n14782), .IN2(g1396), .QN(n16318) );
  NAND2X0 U17072 ( .IN1(n16320), .IN2(n16321), .QN(g20992) );
  NAND2X0 U17073 ( .IN1(n16322), .IN2(g731), .QN(n16321) );
  INVX0 U17074 ( .INP(n15763), .ZN(n16322) );
  NAND2X0 U17075 ( .IN1(n15763), .IN2(n9952), .QN(n16320) );
  NAND2X0 U17076 ( .IN1(n16323), .IN2(n16324), .QN(g20991) );
  NAND2X0 U17077 ( .IN1(n14951), .IN2(n4477), .QN(n16324) );
  NAND2X0 U17078 ( .IN1(n9693), .IN2(g720), .QN(n16323) );
  NAND2X0 U17079 ( .IN1(n16325), .IN2(n16326), .QN(g20990) );
  NAND2X0 U17080 ( .IN1(n14948), .IN2(n9283), .QN(n16326) );
  INVX0 U17081 ( .INP(n16327), .ZN(n16325) );
  NOR2X0 U17082 ( .IN1(n14948), .IN2(n9101), .QN(n16327) );
  NAND2X0 U17083 ( .IN1(n16328), .IN2(n16329), .QN(g20989) );
  NAND2X0 U17084 ( .IN1(n14866), .IN2(n4413), .QN(n16329) );
  NAND2X0 U17085 ( .IN1(n14864), .IN2(g713), .QN(n16328) );
  NAND2X0 U17086 ( .IN1(n16330), .IN2(n16331), .QN(g20983) );
  NAND2X0 U17087 ( .IN1(n14705), .IN2(n4408), .QN(n16331) );
  NAND2X0 U17088 ( .IN1(n10624), .IN2(g2782), .QN(n16330) );
  NAND2X0 U17089 ( .IN1(n16332), .IN2(n16333), .QN(g20982) );
  NAND2X0 U17090 ( .IN1(n4419), .IN2(n14697), .QN(n16333) );
  INVX0 U17091 ( .INP(n16334), .ZN(n16332) );
  NOR2X0 U17092 ( .IN1(n14697), .IN2(n9054), .QN(n16334) );
  NAND2X0 U17093 ( .IN1(n16335), .IN2(n16336), .QN(g20981) );
  NAND2X0 U17094 ( .IN1(n14693), .IN2(n4472), .QN(n16336) );
  NAND2X0 U17095 ( .IN1(n14691), .IN2(g2775), .QN(n16335) );
  NAND2X0 U17096 ( .IN1(n16337), .IN2(n16338), .QN(g20980) );
  NAND2X0 U17097 ( .IN1(n10650), .IN2(g2109), .QN(n16338) );
  INVX0 U17098 ( .INP(n16296), .ZN(n10650) );
  NAND2X0 U17099 ( .IN1(n16296), .IN2(n10237), .QN(n16337) );
  INVX0 U17100 ( .INP(n10293), .ZN(n10237) );
  NAND2X0 U17101 ( .IN1(n16339), .IN2(n16340), .QN(n10293) );
  NAND2X0 U17102 ( .IN1(g1930), .IN2(g2000), .QN(n16340) );
  NOR2X0 U17103 ( .IN1(n16341), .IN2(n16342), .QN(n16339) );
  NOR2X0 U17104 ( .IN1(n8683), .IN2(n4315), .QN(n16342) );
  NOR2X0 U17105 ( .IN1(n8681), .IN2(n4296), .QN(n16341) );
  NOR2X0 U17106 ( .IN1(n4307), .IN2(n9032), .QN(n16296) );
  NAND2X0 U17107 ( .IN1(n16343), .IN2(n16344), .QN(g20979) );
  NAND2X0 U17108 ( .IN1(n4399), .IN2(n14787), .QN(n16344) );
  NAND2X0 U17109 ( .IN1(n10652), .IN2(g2091), .QN(n16343) );
  NAND2X0 U17110 ( .IN1(n16345), .IN2(n16346), .QN(g20978) );
  NAND2X0 U17111 ( .IN1(n14778), .IN2(n4410), .QN(n16346) );
  INVX0 U17112 ( .INP(n16347), .ZN(n16345) );
  NOR2X0 U17113 ( .IN1(n14778), .IN2(n9070), .QN(n16347) );
  NAND2X0 U17114 ( .IN1(n16348), .IN2(n16349), .QN(g20977) );
  NAND2X0 U17115 ( .IN1(n4420), .IN2(n14702), .QN(n16349) );
  NAND2X0 U17116 ( .IN1(n14700), .IN2(g2084), .QN(n16348) );
  NAND2X0 U17117 ( .IN1(n16350), .IN2(n16351), .QN(g20976) );
  NAND2X0 U17118 ( .IN1(n9669), .IN2(g1418), .QN(n16351) );
  NAND2X0 U17119 ( .IN1(n16352), .IN2(n10372), .QN(n16350) );
  INVX0 U17120 ( .INP(n10409), .ZN(n10372) );
  NAND2X0 U17121 ( .IN1(n16353), .IN2(n16354), .QN(n10409) );
  NAND2X0 U17122 ( .IN1(g6944), .IN2(g1294), .QN(n16354) );
  NOR2X0 U17123 ( .IN1(n16355), .IN2(n16356), .QN(n16353) );
  NOR2X0 U17124 ( .IN1(n8693), .IN2(n4300), .QN(n16356) );
  NOR2X0 U17125 ( .IN1(n8692), .IN2(n13695), .QN(n16355) );
  INVX0 U17126 ( .INP(g6750), .ZN(n13695) );
  NAND2X0 U17127 ( .IN1(n16357), .IN2(n16358), .QN(g20975) );
  NAND2X0 U17128 ( .IN1(n13134), .IN2(g1416), .QN(n16358) );
  INVX0 U17129 ( .INP(n14098), .ZN(n13134) );
  NAND2X0 U17130 ( .IN1(n14098), .IN2(n10380), .QN(n16357) );
  NAND2X0 U17131 ( .IN1(n16359), .IN2(n16360), .QN(g20974) );
  NAND2X0 U17132 ( .IN1(n14872), .IN2(n4411), .QN(n16360) );
  NAND2X0 U17133 ( .IN1(n9671), .IN2(g1400), .QN(n16359) );
  NAND2X0 U17134 ( .IN1(n16361), .IN2(n16362), .QN(g20973) );
  NAND2X0 U17135 ( .IN1(n4401), .IN2(n14861), .QN(n16362) );
  INVX0 U17136 ( .INP(n16363), .ZN(n16361) );
  NOR2X0 U17137 ( .IN1(n14861), .IN2(n9087), .QN(n16363) );
  NAND2X0 U17138 ( .IN1(n16364), .IN2(n16365), .QN(g20972) );
  NAND2X0 U17139 ( .IN1(n14784), .IN2(n4412), .QN(n16365) );
  NAND2X0 U17140 ( .IN1(n14782), .IN2(g1393), .QN(n16364) );
  NAND2X0 U17141 ( .IN1(n16366), .IN2(n16367), .QN(g20970) );
  INVX0 U17142 ( .INP(n16368), .ZN(n16367) );
  NOR2X0 U17143 ( .IN1(n9684), .IN2(n8843), .QN(n16368) );
  NAND2X0 U17144 ( .IN1(n9684), .IN2(n9952), .QN(n16366) );
  NAND2X0 U17145 ( .IN1(n16369), .IN2(n16370), .QN(g20969) );
  INVX0 U17146 ( .INP(n16371), .ZN(n16370) );
  NOR2X0 U17147 ( .IN1(n15763), .IN2(n8901), .QN(n16371) );
  NAND2X0 U17148 ( .IN1(n15763), .IN2(n9961), .QN(n16369) );
  NOR2X0 U17149 ( .IN1(n4295), .IN2(n9034), .QN(n15763) );
  NAND2X0 U17150 ( .IN1(n16372), .IN2(n16373), .QN(g20968) );
  NAND2X0 U17151 ( .IN1(n14951), .IN2(n9283), .QN(n16373) );
  NAND2X0 U17152 ( .IN1(n9693), .IN2(g717), .QN(n16372) );
  NAND2X0 U17153 ( .IN1(n16374), .IN2(n16375), .QN(g20967) );
  NAND2X0 U17154 ( .IN1(n14948), .IN2(n4413), .QN(n16375) );
  INVX0 U17155 ( .INP(n16376), .ZN(n16374) );
  NOR2X0 U17156 ( .IN1(n14948), .IN2(n9103), .QN(n16376) );
  NAND2X0 U17157 ( .IN1(n16377), .IN2(n16378), .QN(g20966) );
  NAND2X0 U17158 ( .IN1(n4403), .IN2(n14866), .QN(n16378) );
  NAND2X0 U17159 ( .IN1(n14864), .IN2(g710), .QN(n16377) );
  NAND2X0 U17160 ( .IN1(n16379), .IN2(n16380), .QN(g20965) );
  NAND2X0 U17161 ( .IN1(n4415), .IN2(n14693), .QN(n16380) );
  NAND2X0 U17162 ( .IN1(n14691), .IN2(g2799), .QN(n16379) );
  NAND2X0 U17163 ( .IN1(n16381), .IN2(n16382), .QN(g20964) );
  NAND2X0 U17164 ( .IN1(n4419), .IN2(n14705), .QN(n16382) );
  NAND2X0 U17165 ( .IN1(n10624), .IN2(g2779), .QN(n16381) );
  NAND2X0 U17166 ( .IN1(n16383), .IN2(n16384), .QN(g20963) );
  NAND2X0 U17167 ( .IN1(n14697), .IN2(n4472), .QN(n16384) );
  INVX0 U17168 ( .INP(n16385), .ZN(n16383) );
  NOR2X0 U17169 ( .IN1(n14697), .IN2(n9056), .QN(n16385) );
  NAND2X0 U17170 ( .IN1(n16386), .IN2(n16387), .QN(g20962) );
  NAND2X0 U17171 ( .IN1(n4398), .IN2(n14693), .QN(n16387) );
  INVX0 U17172 ( .INP(n14691), .ZN(n14693) );
  NAND2X0 U17173 ( .IN1(n14691), .IN2(g2772), .QN(n16386) );
  NAND2X0 U17174 ( .IN1(n16388), .IN2(n16113), .QN(n14691) );
  NAND2X0 U17175 ( .IN1(n16389), .IN2(n16390), .QN(g20955) );
  NAND2X0 U17176 ( .IN1(n14787), .IN2(n4410), .QN(n16390) );
  NAND2X0 U17177 ( .IN1(n10652), .IN2(g2088), .QN(n16389) );
  NAND2X0 U17178 ( .IN1(n16391), .IN2(n16392), .QN(g20954) );
  NAND2X0 U17179 ( .IN1(n4420), .IN2(n14778), .QN(n16392) );
  INVX0 U17180 ( .INP(n16393), .ZN(n16391) );
  NOR2X0 U17181 ( .IN1(n14778), .IN2(n9072), .QN(n16393) );
  NAND2X0 U17182 ( .IN1(n16394), .IN2(n16395), .QN(g20953) );
  NAND2X0 U17183 ( .IN1(n14702), .IN2(n4474), .QN(n16395) );
  NAND2X0 U17184 ( .IN1(n14700), .IN2(g2081), .QN(n16394) );
  NAND2X0 U17185 ( .IN1(n16396), .IN2(n16397), .QN(g20952) );
  NAND2X0 U17186 ( .IN1(n9669), .IN2(g1415), .QN(n16397) );
  INVX0 U17187 ( .INP(n16352), .ZN(n9669) );
  NAND2X0 U17188 ( .IN1(n16352), .IN2(n10380), .QN(n16396) );
  INVX0 U17189 ( .INP(n10436), .ZN(n10380) );
  NAND2X0 U17190 ( .IN1(n16398), .IN2(n16399), .QN(n10436) );
  NAND2X0 U17191 ( .IN1(n12608), .IN2(g1300), .QN(n16399) );
  NOR2X0 U17192 ( .IN1(n16400), .IN2(n16401), .QN(n16398) );
  NOR2X0 U17193 ( .IN1(n8686), .IN2(n4316), .QN(n16401) );
  NOR2X0 U17194 ( .IN1(n8685), .IN2(n4300), .QN(n16400) );
  NOR2X0 U17195 ( .IN1(n4308), .IN2(n9033), .QN(n16352) );
  NAND2X0 U17196 ( .IN1(n16402), .IN2(n16403), .QN(g20951) );
  NAND2X0 U17197 ( .IN1(n4401), .IN2(n14872), .QN(n16403) );
  NAND2X0 U17198 ( .IN1(n9671), .IN2(g1397), .QN(n16402) );
  NAND2X0 U17199 ( .IN1(n16404), .IN2(n16405), .QN(g20950) );
  NAND2X0 U17200 ( .IN1(n14861), .IN2(n4412), .QN(n16405) );
  INVX0 U17201 ( .INP(n16406), .ZN(n16404) );
  NOR2X0 U17202 ( .IN1(n14861), .IN2(n9089), .QN(n16406) );
  NAND2X0 U17203 ( .IN1(n16407), .IN2(n16408), .QN(g20949) );
  NAND2X0 U17204 ( .IN1(n4421), .IN2(n14784), .QN(n16408) );
  NAND2X0 U17205 ( .IN1(n14782), .IN2(g1390), .QN(n16407) );
  NAND2X0 U17206 ( .IN1(n16409), .IN2(n16410), .QN(g20948) );
  NAND2X0 U17207 ( .IN1(n9691), .IN2(g732), .QN(n16410) );
  NAND2X0 U17208 ( .IN1(n16411), .IN2(n9952), .QN(n16409) );
  INVX0 U17209 ( .INP(n10001), .ZN(n9952) );
  NAND2X0 U17210 ( .IN1(n16412), .IN2(n16413), .QN(n10001) );
  NAND2X0 U17211 ( .IN1(g6642), .IN2(g608), .QN(n16413) );
  NOR2X0 U17212 ( .IN1(n16414), .IN2(n16415), .QN(n16412) );
  NOR2X0 U17213 ( .IN1(n8676), .IN2(n4313), .QN(n16415) );
  NOR2X0 U17214 ( .IN1(n8675), .IN2(n4298), .QN(n16414) );
  NAND2X0 U17215 ( .IN1(n16416), .IN2(n16417), .QN(g20947) );
  NAND2X0 U17216 ( .IN1(n13251), .IN2(g730), .QN(n16417) );
  INVX0 U17217 ( .INP(n9684), .ZN(n13251) );
  NAND2X0 U17218 ( .IN1(n9684), .IN2(n9961), .QN(n16416) );
  NAND2X0 U17219 ( .IN1(n16418), .IN2(n16419), .QN(g20946) );
  NAND2X0 U17220 ( .IN1(n14951), .IN2(n4413), .QN(n16419) );
  NAND2X0 U17221 ( .IN1(n9693), .IN2(g714), .QN(n16418) );
  NAND2X0 U17222 ( .IN1(n16420), .IN2(n16421), .QN(g20945) );
  NAND2X0 U17223 ( .IN1(n4403), .IN2(n14948), .QN(n16421) );
  INVX0 U17224 ( .INP(n16422), .ZN(n16420) );
  NOR2X0 U17225 ( .IN1(n14948), .IN2(n9105), .QN(n16422) );
  NAND2X0 U17226 ( .IN1(n16423), .IN2(n16424), .QN(g20944) );
  NAND2X0 U17227 ( .IN1(n14866), .IN2(n4414), .QN(n16424) );
  NAND2X0 U17228 ( .IN1(n14864), .IN2(g707), .QN(n16423) );
  NAND2X0 U17229 ( .IN1(n16425), .IN2(n16426), .QN(g20941) );
  NAND2X0 U17230 ( .IN1(n4415), .IN2(n14697), .QN(n16426) );
  INVX0 U17231 ( .INP(n16427), .ZN(n16425) );
  NOR2X0 U17232 ( .IN1(n14697), .IN2(n9040), .QN(n16427) );
  NAND2X0 U17233 ( .IN1(n16428), .IN2(n16429), .QN(g20940) );
  NAND2X0 U17234 ( .IN1(n14705), .IN2(n4472), .QN(n16429) );
  NAND2X0 U17235 ( .IN1(n10624), .IN2(g2776), .QN(n16428) );
  NAND2X0 U17236 ( .IN1(n16430), .IN2(n16431), .QN(g20939) );
  NAND2X0 U17237 ( .IN1(n4398), .IN2(n14697), .QN(n16431) );
  INVX0 U17238 ( .INP(n16432), .ZN(n16430) );
  NOR2X0 U17239 ( .IN1(n14697), .IN2(n9058), .QN(n16432) );
  INVX0 U17240 ( .INP(n14696), .ZN(n14697) );
  NAND2X0 U17241 ( .IN1(n16433), .IN2(n16388), .QN(n14696) );
  NOR2X0 U17242 ( .IN1(n4356), .IN2(g2733), .QN(n16433) );
  NAND2X0 U17243 ( .IN1(n16434), .IN2(n16435), .QN(g20937) );
  NAND2X0 U17244 ( .IN1(n14702), .IN2(n4416), .QN(n16435) );
  NAND2X0 U17245 ( .IN1(n14700), .IN2(g2105), .QN(n16434) );
  NAND2X0 U17246 ( .IN1(n16436), .IN2(n16437), .QN(g20936) );
  NAND2X0 U17247 ( .IN1(n4420), .IN2(n14787), .QN(n16437) );
  NAND2X0 U17248 ( .IN1(n10652), .IN2(g2085), .QN(n16436) );
  NAND2X0 U17249 ( .IN1(n16438), .IN2(n16439), .QN(g20935) );
  NAND2X0 U17250 ( .IN1(n14778), .IN2(n4474), .QN(n16439) );
  INVX0 U17251 ( .INP(n16440), .ZN(n16438) );
  NOR2X0 U17252 ( .IN1(n14778), .IN2(n9074), .QN(n16440) );
  NAND2X0 U17253 ( .IN1(n16441), .IN2(n16442), .QN(g20934) );
  NAND2X0 U17254 ( .IN1(n4400), .IN2(n14702), .QN(n16442) );
  NAND2X0 U17255 ( .IN1(n14700), .IN2(g2078), .QN(n16441) );
  INVX0 U17256 ( .INP(n14702), .ZN(n14700) );
  NOR2X0 U17257 ( .IN1(n16443), .IN2(n4293), .QN(n14702) );
  NAND2X0 U17258 ( .IN1(n16444), .IN2(n16445), .QN(g20927) );
  NAND2X0 U17259 ( .IN1(n14872), .IN2(n4412), .QN(n16445) );
  NAND2X0 U17260 ( .IN1(n9671), .IN2(g1394), .QN(n16444) );
  NAND2X0 U17261 ( .IN1(n16446), .IN2(n16447), .QN(g20926) );
  NAND2X0 U17262 ( .IN1(n4421), .IN2(n14861), .QN(n16447) );
  INVX0 U17263 ( .INP(n16448), .ZN(n16446) );
  NOR2X0 U17264 ( .IN1(n14861), .IN2(n9091), .QN(n16448) );
  NAND2X0 U17265 ( .IN1(n16449), .IN2(n16450), .QN(g20925) );
  NAND2X0 U17266 ( .IN1(n14784), .IN2(n4476), .QN(n16450) );
  NAND2X0 U17267 ( .IN1(n14782), .IN2(g1387), .QN(n16449) );
  NAND2X0 U17268 ( .IN1(n16451), .IN2(n16452), .QN(g20924) );
  NAND2X0 U17269 ( .IN1(n9691), .IN2(g729), .QN(n16452) );
  INVX0 U17270 ( .INP(n16411), .ZN(n9691) );
  NAND2X0 U17271 ( .IN1(n16411), .IN2(n9961), .QN(n16451) );
  INVX0 U17272 ( .INP(n10010), .ZN(n9961) );
  NAND2X0 U17273 ( .IN1(n16453), .IN2(n16454), .QN(n10010) );
  NAND2X0 U17274 ( .IN1(g6642), .IN2(g617), .QN(n16454) );
  NOR2X0 U17275 ( .IN1(n16455), .IN2(n16456), .QN(n16453) );
  INVX0 U17276 ( .INP(n16457), .ZN(n16456) );
  NAND2X0 U17277 ( .IN1(g550), .IN2(test_so26), .QN(n16457) );
  NOR2X0 U17278 ( .IN1(n8673), .IN2(n15378), .QN(n16455) );
  INVX0 U17279 ( .INP(g6485), .ZN(n15378) );
  NOR2X0 U17280 ( .IN1(n4309), .IN2(n9034), .QN(n16411) );
  NAND2X0 U17281 ( .IN1(n16458), .IN2(n16459), .QN(g20923) );
  NAND2X0 U17282 ( .IN1(test_so29), .IN2(n9693), .QN(n16459) );
  NAND2X0 U17283 ( .IN1(n4403), .IN2(n14951), .QN(n16458) );
  NAND2X0 U17284 ( .IN1(n16460), .IN2(n16461), .QN(g20922) );
  NAND2X0 U17285 ( .IN1(n14948), .IN2(n4414), .QN(n16461) );
  INVX0 U17286 ( .INP(n16462), .ZN(n16460) );
  NOR2X0 U17287 ( .IN1(n14948), .IN2(n9106), .QN(n16462) );
  NAND2X0 U17288 ( .IN1(n16463), .IN2(n16464), .QN(g20921) );
  NAND2X0 U17289 ( .IN1(n4422), .IN2(n14866), .QN(n16464) );
  NAND2X0 U17290 ( .IN1(n14864), .IN2(g704), .QN(n16463) );
  NAND2X0 U17291 ( .IN1(n16465), .IN2(n16466), .QN(g20919) );
  NAND2X0 U17292 ( .IN1(n4415), .IN2(n14705), .QN(n16466) );
  NAND2X0 U17293 ( .IN1(n10624), .IN2(g2800), .QN(n16465) );
  NAND2X0 U17294 ( .IN1(n16467), .IN2(n16468), .QN(g20918) );
  NAND2X0 U17295 ( .IN1(n4398), .IN2(n14705), .QN(n16468) );
  INVX0 U17296 ( .INP(n10624), .ZN(n14705) );
  NAND2X0 U17297 ( .IN1(n10624), .IN2(g2773), .QN(n16467) );
  NAND2X0 U17298 ( .IN1(n16469), .IN2(n16388), .QN(n10624) );
  NOR2X0 U17299 ( .IN1(n4490), .IN2(n8992), .QN(n16388) );
  NOR2X0 U17300 ( .IN1(n4306), .IN2(g2733), .QN(n16469) );
  NAND2X0 U17301 ( .IN1(n16470), .IN2(n16471), .QN(g20917) );
  NAND2X0 U17302 ( .IN1(test_so72), .IN2(n14779), .QN(n16471) );
  INVX0 U17303 ( .INP(n14778), .ZN(n14779) );
  NAND2X0 U17304 ( .IN1(n14778), .IN2(n4416), .QN(n16470) );
  NAND2X0 U17305 ( .IN1(n16472), .IN2(n16473), .QN(g20916) );
  NAND2X0 U17306 ( .IN1(n14787), .IN2(n4474), .QN(n16473) );
  NAND2X0 U17307 ( .IN1(n10652), .IN2(g2082), .QN(n16472) );
  NAND2X0 U17308 ( .IN1(n16474), .IN2(n16475), .QN(g20915) );
  NAND2X0 U17309 ( .IN1(n4400), .IN2(n14778), .QN(n16475) );
  INVX0 U17310 ( .INP(n16476), .ZN(n16474) );
  NOR2X0 U17311 ( .IN1(n14778), .IN2(n9076), .QN(n16476) );
  NOR2X0 U17312 ( .IN1(n16443), .IN2(n4357), .QN(n14778) );
  NAND2X0 U17313 ( .IN1(n16477), .IN2(n16478), .QN(g20913) );
  NAND2X0 U17314 ( .IN1(n14784), .IN2(n4417), .QN(n16478) );
  NAND2X0 U17315 ( .IN1(n14782), .IN2(g1411), .QN(n16477) );
  NAND2X0 U17316 ( .IN1(n16479), .IN2(n16480), .QN(g20912) );
  NAND2X0 U17317 ( .IN1(n4421), .IN2(n14872), .QN(n16480) );
  NAND2X0 U17318 ( .IN1(n9671), .IN2(g1391), .QN(n16479) );
  NAND2X0 U17319 ( .IN1(n16481), .IN2(n16482), .QN(g20911) );
  NAND2X0 U17320 ( .IN1(n14861), .IN2(n4476), .QN(n16482) );
  INVX0 U17321 ( .INP(n16483), .ZN(n16481) );
  NOR2X0 U17322 ( .IN1(n14861), .IN2(n9093), .QN(n16483) );
  NAND2X0 U17323 ( .IN1(n16484), .IN2(n16485), .QN(g20910) );
  NAND2X0 U17324 ( .IN1(n4402), .IN2(n14784), .QN(n16485) );
  NAND2X0 U17325 ( .IN1(n14782), .IN2(g1384), .QN(n16484) );
  INVX0 U17326 ( .INP(n14784), .ZN(n14782) );
  NOR2X0 U17327 ( .IN1(n16130), .IN2(n16486), .QN(n14784) );
  NAND2X0 U17328 ( .IN1(n16487), .IN2(n16488), .QN(g20903) );
  NAND2X0 U17329 ( .IN1(n14951), .IN2(n4414), .QN(n16488) );
  NAND2X0 U17330 ( .IN1(n9693), .IN2(g708), .QN(n16487) );
  NAND2X0 U17331 ( .IN1(n16489), .IN2(n16490), .QN(g20902) );
  NAND2X0 U17332 ( .IN1(n4422), .IN2(n14948), .QN(n16490) );
  INVX0 U17333 ( .INP(n16491), .ZN(n16489) );
  NOR2X0 U17334 ( .IN1(n14948), .IN2(n9108), .QN(n16491) );
  NAND2X0 U17335 ( .IN1(n16492), .IN2(n16493), .QN(g20901) );
  NAND2X0 U17336 ( .IN1(n14866), .IN2(n4478), .QN(n16493) );
  NAND2X0 U17337 ( .IN1(n14864), .IN2(g701), .QN(n16492) );
  NAND2X0 U17338 ( .IN1(n16494), .IN2(n16495), .QN(g20900) );
  NAND2X0 U17339 ( .IN1(n14787), .IN2(n4416), .QN(n16495) );
  NAND2X0 U17340 ( .IN1(n10652), .IN2(g2106), .QN(n16494) );
  NAND2X0 U17341 ( .IN1(n16496), .IN2(n16497), .QN(g20899) );
  NAND2X0 U17342 ( .IN1(n4400), .IN2(n14787), .QN(n16497) );
  NAND2X0 U17343 ( .IN1(n10652), .IN2(g2079), .QN(n16496) );
  INVX0 U17344 ( .INP(n14787), .ZN(n10652) );
  NOR2X0 U17345 ( .IN1(n16443), .IN2(n4307), .QN(n14787) );
  NAND2X0 U17346 ( .IN1(n16498), .IN2(test_so69), .QN(n16443) );
  NOR2X0 U17347 ( .IN1(n8993), .IN2(g2039), .QN(n16498) );
  NAND2X0 U17348 ( .IN1(n16499), .IN2(n16500), .QN(g20898) );
  NAND2X0 U17349 ( .IN1(n14861), .IN2(n4417), .QN(n16500) );
  INVX0 U17350 ( .INP(n16501), .ZN(n16499) );
  NOR2X0 U17351 ( .IN1(n14861), .IN2(n9078), .QN(n16501) );
  NAND2X0 U17352 ( .IN1(n16502), .IN2(n16503), .QN(g20897) );
  NAND2X0 U17353 ( .IN1(n14872), .IN2(n4476), .QN(n16503) );
  NAND2X0 U17354 ( .IN1(n9671), .IN2(g1388), .QN(n16502) );
  NAND2X0 U17355 ( .IN1(n16504), .IN2(n16505), .QN(g20896) );
  NAND2X0 U17356 ( .IN1(n4402), .IN2(n14861), .QN(n16505) );
  INVX0 U17357 ( .INP(n16506), .ZN(n16504) );
  NOR2X0 U17358 ( .IN1(n14861), .IN2(n9095), .QN(n16506) );
  INVX0 U17359 ( .INP(n14860), .ZN(n14861) );
  NAND2X0 U17360 ( .IN1(n16507), .IN2(n4428), .QN(n14860) );
  NOR2X0 U17361 ( .IN1(n4358), .IN2(n16486), .QN(n16507) );
  NAND2X0 U17362 ( .IN1(n16508), .IN2(n16509), .QN(g20894) );
  NAND2X0 U17363 ( .IN1(n4418), .IN2(n14866), .QN(n16509) );
  NAND2X0 U17364 ( .IN1(n14864), .IN2(g725), .QN(n16508) );
  NAND2X0 U17365 ( .IN1(n16510), .IN2(n16511), .QN(g20893) );
  NAND2X0 U17366 ( .IN1(n4422), .IN2(n14951), .QN(n16511) );
  NAND2X0 U17367 ( .IN1(n9693), .IN2(g705), .QN(n16510) );
  NAND2X0 U17368 ( .IN1(n16512), .IN2(n16513), .QN(g20892) );
  NAND2X0 U17369 ( .IN1(n14948), .IN2(n4478), .QN(n16513) );
  INVX0 U17370 ( .INP(n16514), .ZN(n16512) );
  NOR2X0 U17371 ( .IN1(n14948), .IN2(n9110), .QN(n16514) );
  NAND2X0 U17372 ( .IN1(n16515), .IN2(n16516), .QN(g20891) );
  NAND2X0 U17373 ( .IN1(n4404), .IN2(n14866), .QN(n16516) );
  INVX0 U17374 ( .INP(n14864), .ZN(n14866) );
  NAND2X0 U17375 ( .IN1(n14864), .IN2(g698), .QN(n16515) );
  NAND2X0 U17376 ( .IN1(n16517), .IN2(n15625), .QN(n14864) );
  NOR2X0 U17377 ( .IN1(g3234), .IN2(DFF_1561_n1), .QN(g20884) );
  NAND2X0 U17378 ( .IN1(n16518), .IN2(n16519), .QN(g20883) );
  NAND2X0 U17379 ( .IN1(n14872), .IN2(n4417), .QN(n16519) );
  NAND2X0 U17380 ( .IN1(n9671), .IN2(g1412), .QN(n16518) );
  NAND2X0 U17381 ( .IN1(n16520), .IN2(n16521), .QN(g20882) );
  NAND2X0 U17382 ( .IN1(test_so49), .IN2(n9671), .QN(n16521) );
  NAND2X0 U17383 ( .IN1(n4402), .IN2(n14872), .QN(n16520) );
  INVX0 U17384 ( .INP(n9671), .ZN(n14872) );
  NAND2X0 U17385 ( .IN1(n16522), .IN2(n4428), .QN(n9671) );
  NOR2X0 U17386 ( .IN1(n4308), .IN2(n16486), .QN(n16522) );
  INVX0 U17387 ( .INP(n16523), .ZN(n16486) );
  NOR2X0 U17388 ( .IN1(n4489), .IN2(n8994), .QN(n16523) );
  NAND2X0 U17389 ( .IN1(n16524), .IN2(n16525), .QN(g20881) );
  NAND2X0 U17390 ( .IN1(test_so30), .IN2(n14947), .QN(n16525) );
  NAND2X0 U17391 ( .IN1(n4418), .IN2(n14948), .QN(n16524) );
  NAND2X0 U17392 ( .IN1(n16526), .IN2(n16527), .QN(g20880) );
  NAND2X0 U17393 ( .IN1(n14951), .IN2(n4478), .QN(n16527) );
  NAND2X0 U17394 ( .IN1(n9693), .IN2(g702), .QN(n16526) );
  NAND2X0 U17395 ( .IN1(n16528), .IN2(n16529), .QN(g20879) );
  NAND2X0 U17396 ( .IN1(n4404), .IN2(n14948), .QN(n16529) );
  INVX0 U17397 ( .INP(n16530), .ZN(n16528) );
  NOR2X0 U17398 ( .IN1(n14948), .IN2(n9112), .QN(n16530) );
  INVX0 U17399 ( .INP(n14947), .ZN(n14948) );
  NAND2X0 U17400 ( .IN1(n16531), .IN2(n16517), .QN(n14947) );
  NOR2X0 U17401 ( .IN1(n4359), .IN2(g659), .QN(n16531) );
  NAND2X0 U17402 ( .IN1(n16532), .IN2(n16533), .QN(g20876) );
  NAND2X0 U17403 ( .IN1(n4418), .IN2(n14951), .QN(n16533) );
  NAND2X0 U17404 ( .IN1(n9693), .IN2(g726), .QN(n16532) );
  NAND2X0 U17405 ( .IN1(n16534), .IN2(n16535), .QN(g20875) );
  NAND2X0 U17406 ( .IN1(n4404), .IN2(n14951), .QN(n16535) );
  INVX0 U17407 ( .INP(n9693), .ZN(n14951) );
  NAND2X0 U17408 ( .IN1(n9693), .IN2(g699), .QN(n16534) );
  NAND2X0 U17409 ( .IN1(n16536), .IN2(n16517), .QN(n9693) );
  NOR2X0 U17410 ( .IN1(n4492), .IN2(n8995), .QN(n16517) );
  NOR2X0 U17411 ( .IN1(n4309), .IN2(g659), .QN(n16536) );
  NAND2X0 U17412 ( .IN1(n16537), .IN2(n16538), .QN(g20874) );
  NAND2X0 U17413 ( .IN1(g2879), .IN2(g8096), .QN(n16538) );
  NAND2X0 U17414 ( .IN1(n4351), .IN2(n16137), .QN(n16537) );
  XNOR2X1 U17415 ( .IN1(n16140), .IN2(n9724), .Q(n16137) );
  XNOR2X1 U17416 ( .IN1(n16539), .IN2(n16540), .Q(n9724) );
  XOR2X1 U17417 ( .IN1(n16541), .IN2(n16542), .Q(n16540) );
  XNOR2X1 U17418 ( .IN1(g2953), .IN2(n9236), .Q(n16542) );
  XNOR2X1 U17419 ( .IN1(g2956), .IN2(n9238), .Q(n16541) );
  XOR2X1 U17420 ( .IN1(n16543), .IN2(n16544), .Q(n16539) );
  XNOR2X1 U17421 ( .IN1(g2938), .IN2(n9234), .Q(n16544) );
  XNOR2X1 U17422 ( .IN1(n9232), .IN2(n9233), .Q(n16543) );
  NOR2X0 U17423 ( .IN1(n16825), .IN2(g3231), .QN(n16140) );
  NOR2X0 U17424 ( .IN1(n10617), .IN2(n16545), .QN(g20789) );
  XNOR2X1 U17425 ( .IN1(n4398), .IN2(n16115), .Q(n16545) );
  INVX0 U17426 ( .INP(n16113), .ZN(n16115) );
  NOR2X0 U17427 ( .IN1(g2733), .IN2(n4292), .QN(n16113) );
  NOR2X0 U17428 ( .IN1(n9031), .IN2(n4356), .QN(n10617) );
  NOR2X0 U17429 ( .IN1(n14094), .IN2(n16546), .QN(g20752) );
  XOR2X1 U17430 ( .IN1(g2020), .IN2(n16119), .Q(n16546) );
  NAND2X0 U17431 ( .IN1(n4427), .IN2(g2009), .QN(n16119) );
  NOR2X0 U17432 ( .IN1(n4357), .IN2(n9032), .QN(n14094) );
  NOR2X0 U17433 ( .IN1(n14098), .IN2(n16547), .QN(g20717) );
  XOR2X1 U17434 ( .IN1(g1326), .IN2(n16130), .Q(n16547) );
  NAND2X0 U17435 ( .IN1(n4428), .IN2(g1315), .QN(n16130) );
  NOR2X0 U17436 ( .IN1(n4358), .IN2(n9033), .QN(n14098) );
  NOR2X0 U17437 ( .IN1(n9684), .IN2(n16548), .QN(g20682) );
  XNOR2X1 U17438 ( .IN1(n4404), .IN2(n15627), .Q(n16548) );
  INVX0 U17439 ( .INP(n15625), .ZN(n15627) );
  NOR2X0 U17440 ( .IN1(g659), .IN2(n4295), .QN(n15625) );
  NOR2X0 U17441 ( .IN1(n9034), .IN2(n4359), .QN(n9684) );
  NAND2X0 U17442 ( .IN1(n16549), .IN2(n16550), .QN(g20417) );
  NAND2X0 U17443 ( .IN1(n4351), .IN2(g2963), .QN(n16550) );
  NAND2X0 U17444 ( .IN1(g2879), .IN2(g7334), .QN(n16549) );
  NAND2X0 U17445 ( .IN1(n16551), .IN2(n16552), .QN(g20376) );
  NAND2X0 U17446 ( .IN1(test_so2), .IN2(n4351), .QN(n16552) );
  NAND2X0 U17447 ( .IN1(g2879), .IN2(g6895), .QN(n16551) );
  NAND2X0 U17448 ( .IN1(n16553), .IN2(n16554), .QN(g20375) );
  NAND2X0 U17449 ( .IN1(n4292), .IN2(g2733), .QN(n16554) );
  NAND2X0 U17450 ( .IN1(n16555), .IN2(g2703), .QN(n16553) );
  NAND2X0 U17451 ( .IN1(n16556), .IN2(n16557), .QN(g20353) );
  NAND2X0 U17452 ( .IN1(n4293), .IN2(g2039), .QN(n16557) );
  NAND2X0 U17453 ( .IN1(n16555), .IN2(g2009), .QN(n16556) );
  NAND2X0 U17454 ( .IN1(n16558), .IN2(n16559), .QN(g20343) );
  NAND2X0 U17455 ( .IN1(n4351), .IN2(g2969), .QN(n16559) );
  NAND2X0 U17456 ( .IN1(g2879), .IN2(g6442), .QN(n16558) );
  NAND2X0 U17457 ( .IN1(n16560), .IN2(n16561), .QN(g20333) );
  INVX0 U17458 ( .INP(n16562), .ZN(n16561) );
  NOR2X0 U17459 ( .IN1(g1315), .IN2(n4428), .QN(n16562) );
  NAND2X0 U17460 ( .IN1(n16555), .IN2(g1315), .QN(n16560) );
  NAND2X0 U17461 ( .IN1(n16563), .IN2(n16564), .QN(g20314) );
  NAND2X0 U17462 ( .IN1(n4295), .IN2(g659), .QN(n16564) );
  NAND2X0 U17463 ( .IN1(n16555), .IN2(g629), .QN(n16563) );
  INVX0 U17464 ( .INP(n15719), .ZN(n16555) );
  NAND2X0 U17465 ( .IN1(n16565), .IN2(n16566), .QN(n15719) );
  NOR2X0 U17466 ( .IN1(g3024), .IN2(n16567), .QN(n16566) );
  NAND2X0 U17467 ( .IN1(n9263), .IN2(n9280), .QN(n16567) );
  NOR2X0 U17468 ( .IN1(g3002), .IN2(g3013), .QN(n16565) );
  NAND2X0 U17469 ( .IN1(n16568), .IN2(n16569), .QN(g20310) );
  NAND2X0 U17470 ( .IN1(n4351), .IN2(g2972), .QN(n16569) );
  NAND2X0 U17471 ( .IN1(g2879), .IN2(g6225), .QN(n16568) );
  NAND2X0 U17472 ( .IN1(n16570), .IN2(n16571), .QN(g19184) );
  NAND2X0 U17473 ( .IN1(n4351), .IN2(g2975), .QN(n16571) );
  NAND2X0 U17474 ( .IN1(g2879), .IN2(g4590), .QN(n16570) );
  NAND2X0 U17475 ( .IN1(n16572), .IN2(n16573), .QN(g19178) );
  NAND2X0 U17476 ( .IN1(n4351), .IN2(g2935), .QN(n16573) );
  NAND2X0 U17477 ( .IN1(test_so5), .IN2(g2879), .QN(n16572) );
  NAND2X0 U17478 ( .IN1(n16574), .IN2(n16575), .QN(g19173) );
  NAND2X0 U17479 ( .IN1(n4351), .IN2(g2978), .QN(n16575) );
  NAND2X0 U17480 ( .IN1(g2879), .IN2(g4323), .QN(n16574) );
  NAND2X0 U17481 ( .IN1(n16576), .IN2(n16577), .QN(g19172) );
  NAND2X0 U17482 ( .IN1(n4351), .IN2(g2953), .QN(n16577) );
  NAND2X0 U17483 ( .IN1(g2879), .IN2(g4321), .QN(n16576) );
  NAND2X0 U17484 ( .IN1(n16578), .IN2(n16579), .QN(g19167) );
  NAND2X0 U17485 ( .IN1(n4351), .IN2(g2938), .QN(n16579) );
  NAND2X0 U17486 ( .IN1(g2879), .IN2(g4200), .QN(n16578) );
  NAND2X0 U17487 ( .IN1(n16580), .IN2(n16581), .QN(g19163) );
  NAND2X0 U17488 ( .IN1(n4351), .IN2(g2981), .QN(n16581) );
  NAND2X0 U17489 ( .IN1(g2879), .IN2(g4090), .QN(n16580) );
  NAND2X0 U17490 ( .IN1(n16582), .IN2(n16583), .QN(g19162) );
  NAND2X0 U17491 ( .IN1(n4351), .IN2(g2956), .QN(n16583) );
  NAND2X0 U17492 ( .IN1(g2879), .IN2(g4088), .QN(n16582) );
  NAND2X0 U17493 ( .IN1(n16584), .IN2(n16585), .QN(g19157) );
  NAND2X0 U17494 ( .IN1(n4351), .IN2(g2941), .QN(n16585) );
  NAND2X0 U17495 ( .IN1(g2879), .IN2(g3993), .QN(n16584) );
  NAND2X0 U17496 ( .IN1(n16586), .IN2(n16587), .QN(g19154) );
  NAND2X0 U17497 ( .IN1(n4351), .IN2(g2874), .QN(n16587) );
  NAND2X0 U17498 ( .IN1(test_so3), .IN2(g2879), .QN(n16586) );
  NAND2X0 U17499 ( .IN1(n16588), .IN2(n16589), .QN(g19153) );
  NAND2X0 U17500 ( .IN1(n4351), .IN2(g2959), .QN(n16589) );
  NAND2X0 U17501 ( .IN1(g2879), .IN2(g8249), .QN(n16588) );
  NAND2X0 U17502 ( .IN1(n16590), .IN2(n16591), .QN(g19149) );
  NAND2X0 U17503 ( .IN1(n4351), .IN2(g2944), .QN(n16591) );
  NAND2X0 U17504 ( .IN1(g2879), .IN2(g8175), .QN(n16590) );
  NAND2X0 U17505 ( .IN1(n16592), .IN2(n16593), .QN(g19144) );
  NAND2X0 U17506 ( .IN1(n4351), .IN2(g2947), .QN(n16593) );
  NAND2X0 U17507 ( .IN1(g2879), .IN2(g8023), .QN(n16592) );
  NAND2X0 U17508 ( .IN1(n16594), .IN2(n16595), .QN(g18975) );
  NAND2X0 U17509 ( .IN1(n4351), .IN2(g2195), .QN(n16595) );
  NAND2X0 U17510 ( .IN1(g2879), .IN2(g2981), .QN(n16594) );
  NAND2X0 U17511 ( .IN1(n16596), .IN2(n16597), .QN(g18968) );
  NAND2X0 U17512 ( .IN1(n4351), .IN2(g2190), .QN(n16597) );
  NAND2X0 U17513 ( .IN1(g2879), .IN2(g2978), .QN(n16596) );
  NAND2X0 U17514 ( .IN1(n16598), .IN2(n16599), .QN(g18957) );
  NAND2X0 U17515 ( .IN1(n4351), .IN2(g2165), .QN(n16599) );
  NAND2X0 U17516 ( .IN1(g2879), .IN2(g2963), .QN(n16598) );
  NAND2X0 U17517 ( .IN1(n16600), .IN2(n16601), .QN(g18942) );
  NAND2X0 U17518 ( .IN1(g2879), .IN2(g2975), .QN(n16601) );
  NAND2X0 U17519 ( .IN1(n4351), .IN2(g2185), .QN(n16600) );
  NAND2X0 U17520 ( .IN1(n16602), .IN2(n16603), .QN(g18907) );
  NAND2X0 U17521 ( .IN1(n4365), .IN2(g3061), .QN(n16603) );
  NAND2X0 U17522 ( .IN1(g2987), .IN2(g2997), .QN(n16602) );
  NAND2X0 U17523 ( .IN1(n16604), .IN2(n16605), .QN(g18906) );
  NAND2X0 U17524 ( .IN1(n4351), .IN2(g2180), .QN(n16605) );
  NAND2X0 U17525 ( .IN1(g2879), .IN2(g2972), .QN(n16604) );
  NAND2X0 U17526 ( .IN1(n16606), .IN2(n16607), .QN(g18885) );
  NAND2X0 U17527 ( .IN1(g2879), .IN2(g2874), .QN(n16607) );
  NAND2X0 U17528 ( .IN1(n4351), .IN2(g2200), .QN(n16606) );
  NAND2X0 U17529 ( .IN1(n16608), .IN2(n16609), .QN(g18883) );
  NAND2X0 U17530 ( .IN1(n4351), .IN2(g1471), .QN(n16609) );
  NAND2X0 U17531 ( .IN1(g2879), .IN2(g2935), .QN(n16608) );
  NAND2X0 U17532 ( .IN1(n16610), .IN2(n16611), .QN(g18868) );
  NAND2X0 U17533 ( .IN1(n4365), .IN2(g3060), .QN(n16611) );
  NAND2X0 U17534 ( .IN1(g2987), .IN2(g3078), .QN(n16610) );
  NAND2X0 U17535 ( .IN1(n16612), .IN2(n16613), .QN(g18867) );
  NAND2X0 U17536 ( .IN1(g2879), .IN2(g2969), .QN(n16613) );
  NAND2X0 U17537 ( .IN1(n4351), .IN2(g2175), .QN(n16612) );
  NAND2X0 U17538 ( .IN1(n16614), .IN2(n16615), .QN(g18866) );
  NAND2X0 U17539 ( .IN1(n4351), .IN2(g1476), .QN(n16615) );
  NAND2X0 U17540 ( .IN1(g2879), .IN2(g2938), .QN(n16614) );
  NAND2X0 U17541 ( .IN1(n16616), .IN2(n16617), .QN(g18852) );
  NAND2X0 U17542 ( .IN1(g2879), .IN2(g2941), .QN(n16617) );
  NAND2X0 U17543 ( .IN1(n4351), .IN2(g1481), .QN(n16616) );
  NAND2X0 U17544 ( .IN1(n16618), .IN2(n16619), .QN(g18837) );
  NAND2X0 U17545 ( .IN1(n4365), .IN2(g3059), .QN(n16619) );
  NAND2X0 U17546 ( .IN1(g2987), .IN2(g3077), .QN(n16618) );
  NAND2X0 U17547 ( .IN1(n16620), .IN2(n16621), .QN(g18836) );
  NAND2X0 U17548 ( .IN1(n4351), .IN2(g2170), .QN(n16621) );
  NAND2X0 U17549 ( .IN1(test_so2), .IN2(g2879), .QN(n16620) );
  NAND2X0 U17550 ( .IN1(n16622), .IN2(n16623), .QN(g18835) );
  NAND2X0 U17551 ( .IN1(n4351), .IN2(g1486), .QN(n16623) );
  NAND2X0 U17552 ( .IN1(g2879), .IN2(g2944), .QN(n16622) );
  NAND2X0 U17553 ( .IN1(n16624), .IN2(n16625), .QN(g18821) );
  NAND2X0 U17554 ( .IN1(g2879), .IN2(g2947), .QN(n16625) );
  NAND2X0 U17555 ( .IN1(n4351), .IN2(g1491), .QN(n16624) );
  NAND2X0 U17556 ( .IN1(n16626), .IN2(n16627), .QN(g18820) );
  NAND2X0 U17557 ( .IN1(n4299), .IN2(g2584), .QN(n16627) );
  NAND2X0 U17558 ( .IN1(g2624), .IN2(g2631), .QN(n16626) );
  NAND2X0 U17559 ( .IN1(n16628), .IN2(n16629), .QN(g18804) );
  NAND2X0 U17560 ( .IN1(n4365), .IN2(g3058), .QN(n16629) );
  NAND2X0 U17561 ( .IN1(g2987), .IN2(g3076), .QN(n16628) );
  NAND2X0 U17562 ( .IN1(n16630), .IN2(n16631), .QN(g18803) );
  NAND2X0 U17563 ( .IN1(n4351), .IN2(g1496), .QN(n16631) );
  NAND2X0 U17564 ( .IN1(g2879), .IN2(g2953), .QN(n16630) );
  NAND2X0 U17565 ( .IN1(n16632), .IN2(n16633), .QN(g18794) );
  NAND2X0 U17566 ( .IN1(g1937), .IN2(g1930), .QN(n16633) );
  NAND2X0 U17567 ( .IN1(n4366), .IN2(g1890), .QN(n16632) );
  NAND2X0 U17568 ( .IN1(n16634), .IN2(n16635), .QN(g18782) );
  NAND2X0 U17569 ( .IN1(g3109), .IN2(g559), .QN(n16635) );
  INVX0 U17570 ( .INP(n16636), .ZN(n16634) );
  NOR2X0 U17571 ( .IN1(g3109), .IN2(n4445), .QN(n16636) );
  NAND2X0 U17572 ( .IN1(n16637), .IN2(n16638), .QN(g18781) );
  NAND2X0 U17573 ( .IN1(n4351), .IN2(g1501), .QN(n16638) );
  NAND2X0 U17574 ( .IN1(g2879), .IN2(g2956), .QN(n16637) );
  NAND2X0 U17575 ( .IN1(n16639), .IN2(n16640), .QN(g18780) );
  NAND2X0 U17576 ( .IN1(n4299), .IN2(g2631), .QN(n16640) );
  NAND2X0 U17577 ( .IN1(n9223), .IN2(g2624), .QN(n16639) );
  NAND2X0 U17578 ( .IN1(n16641), .IN2(n16642), .QN(g18763) );
  NAND2X0 U17579 ( .IN1(n4300), .IN2(g1196), .QN(n16642) );
  NAND2X0 U17580 ( .IN1(g1236), .IN2(g1243), .QN(n16641) );
  NAND2X0 U17581 ( .IN1(n16643), .IN2(n16644), .QN(g18755) );
  NAND2X0 U17582 ( .IN1(n4365), .IN2(g3057), .QN(n16644) );
  NAND2X0 U17583 ( .IN1(g2987), .IN2(g3075), .QN(n16643) );
  NAND2X0 U17584 ( .IN1(n16645), .IN2(n16646), .QN(g18754) );
  NAND2X0 U17585 ( .IN1(g2879), .IN2(g2959), .QN(n16646) );
  NAND2X0 U17586 ( .IN1(n4351), .IN2(g1506), .QN(n16645) );
  NAND2X0 U17587 ( .IN1(n16647), .IN2(n16648), .QN(g18743) );
  NAND2X0 U17588 ( .IN1(n9224), .IN2(g1930), .QN(n16648) );
  NAND2X0 U17589 ( .IN1(n4366), .IN2(g1937), .QN(n16647) );
  NAND2X0 U17590 ( .IN1(n16649), .IN2(n16650), .QN(g18726) );
  NAND2X0 U17591 ( .IN1(test_so22), .IN2(n4313), .QN(n16650) );
  NAND2X0 U17592 ( .IN1(g550), .IN2(g557), .QN(n16649) );
  NAND2X0 U17593 ( .IN1(n16651), .IN2(n16652), .QN(g18719) );
  NAND2X0 U17594 ( .IN1(n4383), .IN2(g3211), .QN(n16652) );
  NAND2X0 U17595 ( .IN1(g8030), .IN2(g559), .QN(n16651) );
  NAND2X0 U17596 ( .IN1(n16653), .IN2(n16654), .QN(g18707) );
  NAND2X0 U17597 ( .IN1(n4300), .IN2(g1243), .QN(n16654) );
  NAND2X0 U17598 ( .IN1(n9225), .IN2(g1236), .QN(n16653) );
  NAND2X0 U17599 ( .IN1(n16655), .IN2(n16656), .QN(g18678) );
  NAND2X0 U17600 ( .IN1(n4313), .IN2(g557), .QN(n16656) );
  NAND2X0 U17601 ( .IN1(n9226), .IN2(g550), .QN(n16655) );
  NAND2X0 U17602 ( .IN1(n16657), .IN2(n16658), .QN(g18669) );
  NAND2X0 U17603 ( .IN1(n4382), .IN2(test_so6), .QN(n16658) );
  NAND2X0 U17604 ( .IN1(g8106), .IN2(g559), .QN(n16657) );
  NAND2X0 U17605 ( .IN1(n16659), .IN2(n16660), .QN(g17429) );
  NAND2X0 U17606 ( .IN1(g3109), .IN2(g2574), .QN(n16660) );
  INVX0 U17607 ( .INP(n16661), .ZN(n16659) );
  NOR2X0 U17608 ( .IN1(g3109), .IN2(n4341), .QN(n16661) );
  NAND2X0 U17609 ( .IN1(n16662), .IN2(n16663), .QN(g17383) );
  NAND2X0 U17610 ( .IN1(n4494), .IN2(test_so8), .QN(n16663) );
  NAND2X0 U17611 ( .IN1(g3109), .IN2(g1880), .QN(n16662) );
  NAND2X0 U17612 ( .IN1(n16664), .IN2(n16665), .QN(g17341) );
  INVX0 U17613 ( .INP(n16666), .ZN(n16665) );
  NOR2X0 U17614 ( .IN1(g8030), .IN2(n4442), .QN(n16666) );
  NAND2X0 U17615 ( .IN1(g8030), .IN2(g2574), .QN(n16664) );
  NAND2X0 U17616 ( .IN1(n16667), .IN2(n16668), .QN(g17340) );
  NAND2X0 U17617 ( .IN1(g3109), .IN2(g1186), .QN(n16668) );
  INVX0 U17618 ( .INP(n16669), .ZN(n16667) );
  NOR2X0 U17619 ( .IN1(g3109), .IN2(n4441), .QN(n16669) );
  NAND2X0 U17620 ( .IN1(n16670), .IN2(n16671), .QN(g17303) );
  INVX0 U17621 ( .INP(n16672), .ZN(n16671) );
  NOR2X0 U17622 ( .IN1(g8030), .IN2(n4450), .QN(n16672) );
  NAND2X0 U17623 ( .IN1(g8030), .IN2(g1880), .QN(n16670) );
  NAND2X0 U17624 ( .IN1(n16673), .IN2(n16674), .QN(g17302) );
  NAND2X0 U17625 ( .IN1(g3109), .IN2(g499), .QN(n16674) );
  NAND2X0 U17626 ( .IN1(n4494), .IN2(g3161), .QN(n16673) );
  NAND2X0 U17627 ( .IN1(n16675), .IN2(n16676), .QN(g17271) );
  INVX0 U17628 ( .INP(n16677), .ZN(n16676) );
  NOR2X0 U17629 ( .IN1(g8106), .IN2(n4453), .QN(n16677) );
  NAND2X0 U17630 ( .IN1(g8106), .IN2(g2574), .QN(n16675) );
  NAND2X0 U17631 ( .IN1(n16678), .IN2(n16679), .QN(g17270) );
  NAND2X0 U17632 ( .IN1(g8030), .IN2(g1186), .QN(n16679) );
  INVX0 U17633 ( .INP(n16680), .ZN(n16678) );
  NOR2X0 U17634 ( .IN1(g8030), .IN2(n4348), .QN(n16680) );
  NAND2X0 U17635 ( .IN1(n16681), .IN2(n16682), .QN(g17269) );
  NAND2X0 U17636 ( .IN1(g3109), .IN2(g2633), .QN(n16682) );
  NAND2X0 U17637 ( .IN1(n4494), .IN2(g3096), .QN(n16681) );
  NAND2X0 U17638 ( .IN1(n16683), .IN2(n16684), .QN(g17248) );
  NAND2X0 U17639 ( .IN1(g8106), .IN2(g1880), .QN(n16684) );
  INVX0 U17640 ( .INP(n16685), .ZN(n16683) );
  NOR2X0 U17641 ( .IN1(g8106), .IN2(n4338), .QN(n16685) );
  NAND2X0 U17642 ( .IN1(n16686), .IN2(n16687), .QN(g17247) );
  INVX0 U17643 ( .INP(n16688), .ZN(n16687) );
  NOR2X0 U17644 ( .IN1(g8030), .IN2(n4436), .QN(n16688) );
  NAND2X0 U17645 ( .IN1(g8030), .IN2(g499), .QN(n16686) );
  NAND2X0 U17646 ( .IN1(n16689), .IN2(n16690), .QN(g17246) );
  NAND2X0 U17647 ( .IN1(g3109), .IN2(g1939), .QN(n16690) );
  NAND2X0 U17648 ( .IN1(n4494), .IN2(g3093), .QN(n16689) );
  NAND2X0 U17649 ( .IN1(n16691), .IN2(n16692), .QN(g17236) );
  NAND2X0 U17650 ( .IN1(g8106), .IN2(g1186), .QN(n16692) );
  INVX0 U17651 ( .INP(n16693), .ZN(n16691) );
  NOR2X0 U17652 ( .IN1(g8106), .IN2(n4339), .QN(n16693) );
  NAND2X0 U17653 ( .IN1(n16694), .IN2(n16695), .QN(g17235) );
  INVX0 U17654 ( .INP(n16696), .ZN(n16695) );
  NOR2X0 U17655 ( .IN1(g8030), .IN2(n4439), .QN(n16696) );
  NAND2X0 U17656 ( .IN1(g8030), .IN2(g2633), .QN(n16694) );
  NAND2X0 U17657 ( .IN1(n16697), .IN2(n16698), .QN(g17234) );
  NAND2X0 U17658 ( .IN1(g3109), .IN2(g1245), .QN(n16698) );
  INVX0 U17659 ( .INP(n16699), .ZN(n16697) );
  NOR2X0 U17660 ( .IN1(g3109), .IN2(n4344), .QN(n16699) );
  NAND2X0 U17661 ( .IN1(n16700), .IN2(n16701), .QN(g17229) );
  NAND2X0 U17662 ( .IN1(n4382), .IN2(g3155), .QN(n16701) );
  NAND2X0 U17663 ( .IN1(g8106), .IN2(g499), .QN(n16700) );
  NAND2X0 U17664 ( .IN1(n16702), .IN2(n16703), .QN(g17228) );
  INVX0 U17665 ( .INP(n16704), .ZN(n16703) );
  NOR2X0 U17666 ( .IN1(g8030), .IN2(n4451), .QN(n16704) );
  NAND2X0 U17667 ( .IN1(g8030), .IN2(g1939), .QN(n16702) );
  NAND2X0 U17668 ( .IN1(n16705), .IN2(n16706), .QN(g17226) );
  NAND2X0 U17669 ( .IN1(n4382), .IN2(g3094), .QN(n16706) );
  NAND2X0 U17670 ( .IN1(g8106), .IN2(g2633), .QN(n16705) );
  NAND2X0 U17671 ( .IN1(n16707), .IN2(n16708), .QN(g17225) );
  NAND2X0 U17672 ( .IN1(g8030), .IN2(g1245), .QN(n16708) );
  INVX0 U17673 ( .INP(n16709), .ZN(n16707) );
  NOR2X0 U17674 ( .IN1(g8030), .IN2(n4337), .QN(n16709) );
  NAND2X0 U17675 ( .IN1(n16710), .IN2(n16711), .QN(g17224) );
  INVX0 U17676 ( .INP(n16712), .ZN(n16711) );
  NOR2X0 U17677 ( .IN1(g8106), .IN2(n4448), .QN(n16712) );
  NAND2X0 U17678 ( .IN1(g8106), .IN2(g1939), .QN(n16710) );
  NAND2X0 U17679 ( .IN1(n16713), .IN2(n16714), .QN(g17222) );
  NAND2X0 U17680 ( .IN1(g8106), .IN2(g1245), .QN(n16714) );
  NAND2X0 U17681 ( .IN1(n4382), .IN2(g3085), .QN(n16713) );
  NAND2X0 U17682 ( .IN1(n16715), .IN2(n16716), .QN(g16880) );
  NAND2X0 U17683 ( .IN1(n4365), .IN2(g3056), .QN(n16716) );
  NAND2X0 U17684 ( .IN1(g2987), .IN2(g3074), .QN(n16715) );
  NAND2X0 U17685 ( .IN1(n16717), .IN2(n16718), .QN(g16866) );
  NAND2X0 U17686 ( .IN1(n4365), .IN2(g3051), .QN(n16718) );
  NAND2X0 U17687 ( .IN1(test_so97), .IN2(g2987), .QN(n16717) );
  NAND2X0 U17688 ( .IN1(n16719), .IN2(n16720), .QN(g16861) );
  NAND2X0 U17689 ( .IN1(test_so96), .IN2(n4365), .QN(n16720) );
  NAND2X0 U17690 ( .IN1(g2987), .IN2(g3073), .QN(n16719) );
  NAND2X0 U17691 ( .IN1(n16721), .IN2(n16722), .QN(g16860) );
  NAND2X0 U17692 ( .IN1(n4365), .IN2(g3046), .QN(n16722) );
  NAND2X0 U17693 ( .IN1(g2987), .IN2(g3065), .QN(n16721) );
  NAND2X0 U17694 ( .IN1(n16723), .IN2(n16724), .QN(g16857) );
  NAND2X0 U17695 ( .IN1(n4365), .IN2(g3050), .QN(n16724) );
  NAND2X0 U17696 ( .IN1(g2987), .IN2(g3069), .QN(n16723) );
  NAND2X0 U17697 ( .IN1(n16725), .IN2(n16726), .QN(g16854) );
  NAND2X0 U17698 ( .IN1(n4365), .IN2(g3053), .QN(n16726) );
  NAND2X0 U17699 ( .IN1(g2987), .IN2(g3072), .QN(n16725) );
  NAND2X0 U17700 ( .IN1(n16727), .IN2(n16728), .QN(g16853) );
  NAND2X0 U17701 ( .IN1(n4365), .IN2(g3045), .QN(n16728) );
  NAND2X0 U17702 ( .IN1(g2987), .IN2(g3064), .QN(n16727) );
  NAND2X0 U17703 ( .IN1(n16729), .IN2(n16730), .QN(g16851) );
  NAND2X0 U17704 ( .IN1(n4365), .IN2(g3049), .QN(n16730) );
  NAND2X0 U17705 ( .IN1(g2987), .IN2(g3068), .QN(n16729) );
  NAND2X0 U17706 ( .IN1(n16731), .IN2(n16732), .QN(g16845) );
  NAND2X0 U17707 ( .IN1(n4365), .IN2(g3052), .QN(n16732) );
  NAND2X0 U17708 ( .IN1(g2987), .IN2(g3071), .QN(n16731) );
  NAND2X0 U17709 ( .IN1(n16733), .IN2(n16734), .QN(g16844) );
  NAND2X0 U17710 ( .IN1(n4365), .IN2(g3044), .QN(n16734) );
  NAND2X0 U17711 ( .IN1(g2987), .IN2(g3063), .QN(n16733) );
  NAND2X0 U17712 ( .IN1(n16735), .IN2(n16736), .QN(g16835) );
  NAND2X0 U17713 ( .IN1(n4365), .IN2(g3048), .QN(n16736) );
  NAND2X0 U17714 ( .IN1(g2987), .IN2(g3067), .QN(n16735) );
  NAND2X0 U17715 ( .IN1(n16737), .IN2(n16738), .QN(g16824) );
  NAND2X0 U17716 ( .IN1(n4365), .IN2(g3043), .QN(n16738) );
  NAND2X0 U17717 ( .IN1(g2987), .IN2(g3062), .QN(n16737) );
  NOR2X0 U17718 ( .IN1(g51), .IN2(DFF_1_n1), .QN(g16823) );
  NAND2X0 U17719 ( .IN1(n16739), .IN2(n16740), .QN(g16803) );
  NAND2X0 U17720 ( .IN1(n4365), .IN2(g3047), .QN(n16740) );
  NAND2X0 U17721 ( .IN1(g2987), .IN2(g3066), .QN(n16739) );
  NOR2X0 U17722 ( .IN1(n4423), .IN2(g51), .QN(g16802) );
  NAND2X0 U17723 ( .IN1(n16741), .IN2(n16742), .QN(g16718) );
  INVX0 U17724 ( .INP(n16743), .ZN(n16742) );
  NOR2X0 U17725 ( .IN1(g2703), .IN2(n9031), .QN(n16743) );
  NAND2X0 U17726 ( .IN1(g2703), .IN2(g2584), .QN(n16741) );
  NAND2X0 U17727 ( .IN1(n16744), .IN2(n16745), .QN(g16692) );
  INVX0 U17728 ( .INP(n16746), .ZN(n16745) );
  NOR2X0 U17729 ( .IN1(g2009), .IN2(n9032), .QN(n16746) );
  NAND2X0 U17730 ( .IN1(g2009), .IN2(g1890), .QN(n16744) );
  NAND2X0 U17731 ( .IN1(n16747), .IN2(n16748), .QN(g16671) );
  INVX0 U17732 ( .INP(n16749), .ZN(n16748) );
  NOR2X0 U17733 ( .IN1(g1315), .IN2(n9033), .QN(n16749) );
  NAND2X0 U17734 ( .IN1(g1315), .IN2(g1196), .QN(n16747) );
  NAND2X0 U17735 ( .IN1(n16750), .IN2(n16751), .QN(g16654) );
  INVX0 U17736 ( .INP(n16752), .ZN(n16751) );
  NOR2X0 U17737 ( .IN1(g629), .IN2(n9034), .QN(n16752) );
  NAND2X0 U17738 ( .IN1(test_so22), .IN2(g629), .QN(n16750) );
  NAND2X0 U17739 ( .IN1(n16753), .IN2(g2987), .QN(g16496) );
  NAND2X0 U17740 ( .IN1(DFF_1612_n1), .IN2(g5388), .QN(n16753) );
  NOR2X0 U17741 ( .IN1(n16754), .IN2(n16755), .QN(g13194) );
  NAND2X0 U17742 ( .IN1(n16756), .IN2(n16757), .QN(n16755) );
  INVX0 U17743 ( .INP(n16758), .ZN(n16757) );
  NOR2X0 U17744 ( .IN1(n4314), .IN2(test_so87), .QN(n16758) );
  NAND2X0 U17745 ( .IN1(n8996), .IN2(g7390), .QN(n16756) );
  NOR2X0 U17746 ( .IN1(n4299), .IN2(g2562), .QN(n16754) );
  NOR2X0 U17747 ( .IN1(n16759), .IN2(n16760), .QN(g13182) );
  NAND2X0 U17748 ( .IN1(n16761), .IN2(n16762), .QN(n16760) );
  NAND2X0 U17749 ( .IN1(n9005), .IN2(n12749), .QN(n16762) );
  NAND2X0 U17750 ( .IN1(n9004), .IN2(g7194), .QN(n16761) );
  NOR2X0 U17751 ( .IN1(n4366), .IN2(g1868), .QN(n16759) );
  NOR2X0 U17752 ( .IN1(n16763), .IN2(n16764), .QN(g13175) );
  NAND2X0 U17753 ( .IN1(n16765), .IN2(n16766), .QN(n16764) );
  NAND2X0 U17754 ( .IN1(n9002), .IN2(n11699), .QN(n16766) );
  NAND2X0 U17755 ( .IN1(n9001), .IN2(g7390), .QN(n16765) );
  NOR2X0 U17756 ( .IN1(n4299), .IN2(g2553), .QN(n16763) );
  NOR2X0 U17757 ( .IN1(n16767), .IN2(n16768), .QN(g13171) );
  NAND2X0 U17758 ( .IN1(n16769), .IN2(n16770), .QN(n16768) );
  INVX0 U17759 ( .INP(n16771), .ZN(n16770) );
  NOR2X0 U17760 ( .IN1(n4300), .IN2(test_so44), .QN(n16771) );
  NAND2X0 U17761 ( .IN1(n9013), .IN2(g6944), .QN(n16769) );
  NOR2X0 U17762 ( .IN1(n4371), .IN2(g1175), .QN(n16767) );
  NOR2X0 U17763 ( .IN1(n16772), .IN2(n16773), .QN(g13164) );
  NAND2X0 U17764 ( .IN1(n16774), .IN2(n16775), .QN(n16773) );
  NAND2X0 U17765 ( .IN1(n9011), .IN2(n12749), .QN(n16775) );
  NAND2X0 U17766 ( .IN1(n9010), .IN2(g7194), .QN(n16774) );
  NOR2X0 U17767 ( .IN1(n4366), .IN2(g1859), .QN(n16772) );
  NOR2X0 U17768 ( .IN1(n16776), .IN2(n16777), .QN(g13160) );
  NAND2X0 U17769 ( .IN1(n16778), .IN2(n16779), .QN(n16777) );
  NAND2X0 U17770 ( .IN1(n9022), .IN2(n13002), .QN(n16779) );
  NAND2X0 U17771 ( .IN1(n9021), .IN2(g6642), .QN(n16778) );
  NOR2X0 U17772 ( .IN1(n4313), .IN2(g487), .QN(n16776) );
  NOR2X0 U17773 ( .IN1(n16780), .IN2(n16781), .QN(g13155) );
  NAND2X0 U17774 ( .IN1(n16782), .IN2(n16783), .QN(n16781) );
  NAND2X0 U17775 ( .IN1(n9018), .IN2(g6944), .QN(n16783) );
  NAND2X0 U17776 ( .IN1(n9019), .IN2(n12608), .QN(n16782) );
  NOR2X0 U17777 ( .IN1(n4300), .IN2(g1165), .QN(n16780) );
  NOR2X0 U17778 ( .IN1(n16784), .IN2(n16785), .QN(g13149) );
  NAND2X0 U17779 ( .IN1(n16786), .IN2(n16787), .QN(n16785) );
  NAND2X0 U17780 ( .IN1(n9028), .IN2(n13002), .QN(n16787) );
  NAND2X0 U17781 ( .IN1(n9027), .IN2(g6642), .QN(n16786) );
  NOR2X0 U17782 ( .IN1(n4313), .IN2(g478), .QN(n16784) );
  NOR2X0 U17783 ( .IN1(n16788), .IN2(n16789), .QN(g13143) );
  NAND2X0 U17784 ( .IN1(n16790), .IN2(n16791), .QN(n16789) );
  NAND2X0 U17785 ( .IN1(n8999), .IN2(n11699), .QN(n16791) );
  INVX0 U17786 ( .INP(n4314), .ZN(n11699) );
  NAND2X0 U17787 ( .IN1(n8998), .IN2(g7390), .QN(n16790) );
  NOR2X0 U17788 ( .IN1(n4299), .IN2(g2559), .QN(n16788) );
  NOR2X0 U17789 ( .IN1(n16792), .IN2(n16793), .QN(g13135) );
  NAND2X0 U17790 ( .IN1(n16794), .IN2(n16795), .QN(n16793) );
  NAND2X0 U17791 ( .IN1(n9008), .IN2(n12749), .QN(n16795) );
  INVX0 U17792 ( .INP(n4296), .ZN(n12749) );
  NAND2X0 U17793 ( .IN1(n9007), .IN2(g7194), .QN(n16794) );
  NOR2X0 U17794 ( .IN1(n4366), .IN2(g1865), .QN(n16792) );
  NOR2X0 U17795 ( .IN1(n16796), .IN2(n16797), .QN(g13124) );
  NAND2X0 U17796 ( .IN1(n16798), .IN2(n16799), .QN(n16797) );
  NAND2X0 U17797 ( .IN1(n9015), .IN2(g6944), .QN(n16799) );
  NAND2X0 U17798 ( .IN1(n9016), .IN2(n12608), .QN(n16798) );
  INVX0 U17799 ( .INP(n4371), .ZN(n12608) );
  NOR2X0 U17800 ( .IN1(n4300), .IN2(g1171), .QN(n16796) );
  NOR2X0 U17801 ( .IN1(n16800), .IN2(n16801), .QN(g13111) );
  NAND2X0 U17802 ( .IN1(n16802), .IN2(n16803), .QN(n16801) );
  NAND2X0 U17803 ( .IN1(n9025), .IN2(n13002), .QN(n16803) );
  INVX0 U17804 ( .INP(n4298), .ZN(n13002) );
  NAND2X0 U17805 ( .IN1(n9024), .IN2(g6642), .QN(n16802) );
  NOR2X0 U17806 ( .IN1(n4313), .IN2(g484), .QN(n16800) );
  XNOR2X1 U17807 ( .IN1(n9937), .IN2(n9253), .Q(N995) );
  XNOR2X1 U17808 ( .IN1(n16804), .IN2(n16805), .Q(n9937) );
  XOR2X1 U17809 ( .IN1(n16806), .IN2(n16807), .Q(n16805) );
  XOR2X1 U17810 ( .IN1(n16836), .IN2(n9250), .Q(n16807) );
  XOR2X1 U17811 ( .IN1(test_so99), .IN2(n16835), .Q(n16806) );
  XOR2X1 U17812 ( .IN1(n16808), .IN2(n16809), .Q(n16804) );
  XOR2X1 U17813 ( .IN1(n9249), .IN2(n9248), .Q(n16809) );
  XOR2X1 U17814 ( .IN1(DFF_1618_n1), .IN2(n9247), .Q(n16808) );
  XOR2X1 U17815 ( .IN1(n9251), .IN2(n9938), .Q(N690) );
  XNOR2X1 U17816 ( .IN1(n16810), .IN2(n16811), .Q(n9938) );
  XOR2X1 U17817 ( .IN1(n16812), .IN2(n16813), .Q(n16811) );
  XOR2X1 U17818 ( .IN1(n9231), .IN2(n9230), .Q(n16813) );
  XOR2X1 U17819 ( .IN1(n16837), .IN2(n16838), .Q(n16812) );
  XOR2X1 U17820 ( .IN1(n16814), .IN2(n16815), .Q(n16810) );
  XOR2X1 U17821 ( .IN1(n9229), .IN2(n9228), .Q(n16815) );
  XOR2X1 U17822 ( .IN1(DFF_1628_n1), .IN2(n9227), .Q(n16814) );
  NOR2X0 U3772_U2 ( .IN1(n2230), .IN2(n2217), .QN(U3772_n1) );
  INVX0 U3772_U1 ( .INP(U3772_n1), .ZN(n2231) );
  NOR2X0 U3776_U2 ( .IN1(n2374), .IN2(n2361), .QN(U3776_n1) );
  INVX0 U3776_U1 ( .INP(U3776_n1), .ZN(n2375) );
  NOR2X0 U3777_U2 ( .IN1(g51), .IN2(DFF_2_n1), .QN(U3777_n1) );
  INVX0 U3777_U1 ( .INP(U3777_n1), .ZN(n4264) );
  NOR2X0 U3778_U2 ( .IN1(n2445), .IN2(n2446), .QN(U3778_n1) );
  INVX0 U3778_U1 ( .INP(U3778_n1), .ZN(n2440) );
  NOR2X0 U3779_U2 ( .IN1(n492), .IN2(n2446), .QN(U3779_n1) );
  INVX0 U3779_U1 ( .INP(U3779_n1), .ZN(n2426) );
  NOR2X0 U3780_U2 ( .IN1(n2670), .IN2(n2671), .QN(U3780_n1) );
  INVX0 U3780_U1 ( .INP(U3780_n1), .ZN(n2669) );
  NOR2X0 U3781_U2 ( .IN1(n2685), .IN2(n2686), .QN(U3781_n1) );
  INVX0 U3781_U1 ( .INP(U3781_n1), .ZN(n2684) );
  NOR2X0 U3782_U2 ( .IN1(n2718), .IN2(n2719), .QN(U3782_n1) );
  INVX0 U3782_U1 ( .INP(U3782_n1), .ZN(n2717) );
  NOR2X0 U3783_U2 ( .IN1(n2982), .IN2(g2124), .QN(U3783_n1) );
  INVX0 U3783_U1 ( .INP(U3783_n1), .ZN(n2981) );
  NOR2X0 U3784_U2 ( .IN1(n2985), .IN2(g1430), .QN(U3784_n1) );
  INVX0 U3784_U1 ( .INP(U3784_n1), .ZN(n2984) );
  NOR2X0 U3785_U2 ( .IN1(n2988), .IN2(g744), .QN(U3785_n1) );
  INVX0 U3785_U1 ( .INP(U3785_n1), .ZN(n2987) );
  NOR2X0 U3786_U2 ( .IN1(n2991), .IN2(g56), .QN(U3786_n1) );
  INVX0 U3786_U1 ( .INP(U3786_n1), .ZN(n2990) );
  NOR2X0 U3787_U2 ( .IN1(n3742), .IN2(test_so98), .QN(U3787_n1) );
  INVX0 U3787_U1 ( .INP(U3787_n1), .ZN(n3741) );
  NOR2X0 U3901_U2 ( .IN1(n2302), .IN2(n2289), .QN(U3901_n1) );
  INVX0 U3901_U1 ( .INP(U3901_n1), .ZN(n2303) );
  NOR2X0 U3902_U2 ( .IN1(n522), .IN2(n2289), .QN(U3902_n1) );
  INVX0 U3902_U1 ( .INP(U3902_n1), .ZN(n2275) );
  INVX0 U4467_U2 ( .INP(n1421), .ZN(U4467_n1) );
  NOR2X0 U4467_U1 ( .IN1(n3254), .IN2(U4467_n1), .QN(n3252) );
  INVX0 U4904_U2 ( .INP(n2800), .ZN(U4904_n1) );
  NOR2X0 U4904_U1 ( .IN1(n158), .IN2(U4904_n1), .QN(n2798) );
  INVX0 U4930_U2 ( .INP(n2616), .ZN(U4930_n1) );
  NOR2X0 U4930_U1 ( .IN1(n158), .IN2(U4930_n1), .QN(n2594) );
  INVX0 U5128_U2 ( .INP(n3933), .ZN(U5128_n1) );
  NOR2X0 U5128_U1 ( .IN1(n4406), .IN2(U5128_n1), .QN(n3940) );
  INVX0 U5141_U2 ( .INP(n3939), .ZN(U5141_n1) );
  NOR2X0 U5141_U1 ( .IN1(n4405), .IN2(U5141_n1), .QN(n3936) );
  INVX0 U5749_U2 ( .INP(g2133), .ZN(U5749_n1) );
  NOR2X0 U5749_U1 ( .IN1(n3160), .IN2(U5749_n1), .QN(n3159) );
  INVX0 U5750_U2 ( .INP(g1439), .ZN(U5750_n1) );
  NOR2X0 U5750_U1 ( .IN1(n3164), .IN2(U5750_n1), .QN(n3163) );
  INVX0 U5751_U2 ( .INP(g753), .ZN(U5751_n1) );
  NOR2X0 U5751_U1 ( .IN1(n3168), .IN2(U5751_n1), .QN(n3167) );
  INVX0 U5752_U2 ( .INP(g65), .ZN(U5752_n1) );
  NOR2X0 U5752_U1 ( .IN1(n3172), .IN2(U5752_n1), .QN(n3171) );
  INVX0 U5753_U2 ( .INP(g2142), .ZN(U5753_n1) );
  NOR2X0 U5753_U1 ( .IN1(n4522), .IN2(U5753_n1), .QN(n3424) );
  INVX0 U5754_U2 ( .INP(g2151), .ZN(U5754_n1) );
  NOR2X0 U5754_U1 ( .IN1(n4526), .IN2(U5754_n1), .QN(n3683) );
  INVX0 U5755_U2 ( .INP(g2160), .ZN(U5755_n1) );
  NOR2X0 U5755_U1 ( .IN1(n3888), .IN2(U5755_n1), .QN(n3887) );
  INVX0 U5756_U2 ( .INP(g1448), .ZN(U5756_n1) );
  NOR2X0 U5756_U1 ( .IN1(n4523), .IN2(U5756_n1), .QN(n3427) );
  INVX0 U5757_U2 ( .INP(g1457), .ZN(U5757_n1) );
  NOR2X0 U5757_U1 ( .IN1(n4527), .IN2(U5757_n1), .QN(n3686) );
  INVX0 U5758_U2 ( .INP(g1466), .ZN(U5758_n1) );
  NOR2X0 U5758_U1 ( .IN1(n3891), .IN2(U5758_n1), .QN(n3890) );
  INVX0 U5759_U2 ( .INP(g762), .ZN(U5759_n1) );
  NOR2X0 U5759_U1 ( .IN1(n3431), .IN2(U5759_n1), .QN(n3430) );
  INVX0 U5760_U2 ( .INP(g771), .ZN(U5760_n1) );
  NOR2X0 U5760_U1 ( .IN1(n3690), .IN2(U5760_n1), .QN(n3689) );
  INVX0 U5761_U2 ( .INP(g780), .ZN(U5761_n1) );
  NOR2X0 U5761_U1 ( .IN1(n3894), .IN2(U5761_n1), .QN(n3893) );
  INVX0 U5762_U2 ( .INP(g74), .ZN(U5762_n1) );
  NOR2X0 U5762_U1 ( .IN1(n4521), .IN2(U5762_n1), .QN(n3433) );
  INVX0 U5763_U2 ( .INP(g83), .ZN(U5763_n1) );
  NOR2X0 U5763_U1 ( .IN1(n4528), .IN2(U5763_n1), .QN(n3692) );
  INVX0 U5764_U2 ( .INP(g92), .ZN(U5764_n1) );
  NOR2X0 U5764_U1 ( .IN1(n3897), .IN2(U5764_n1), .QN(n3896) );
  INVX0 U5882_U2 ( .INP(n4102), .ZN(U5882_n1) );
  NOR2X0 U5882_U1 ( .IN1(g3036), .IN2(U5882_n1), .QN(n4101) );
  INVX0 U5939_U2 ( .INP(g2257), .ZN(U5939_n1) );
  NOR2X0 U5939_U1 ( .IN1(n1290), .IN2(U5939_n1), .QN(n3038) );
  INVX0 U5940_U2 ( .INP(g1563), .ZN(U5940_n1) );
  NOR2X0 U5940_U1 ( .IN1(n984), .IN2(U5940_n1), .QN(n3070) );
  INVX0 U5941_U2 ( .INP(g869), .ZN(U5941_n1) );
  NOR2X0 U5941_U1 ( .IN1(n681), .IN2(U5941_n1), .QN(n3102) );
  INVX0 U5942_U2 ( .INP(g181), .ZN(U5942_n1) );
  NOR2X0 U5942_U1 ( .IN1(n348), .IN2(U5942_n1), .QN(n3130) );
  INVX0 U6140_U2 ( .INP(g3002), .ZN(U6140_n1) );
  NOR2X0 U6140_U1 ( .IN1(n4066), .IN2(U6140_n1), .QN(n4065) );
  INVX0 U6460_U2 ( .INP(g3233), .ZN(U6460_n1) );
  NOR2X0 U6460_U1 ( .IN1(g3230), .IN2(U6460_n1), .QN(n3700) );
  INVX0 U6470_U2 ( .INP(g2892), .ZN(U6470_n1) );
  NOR2X0 U6470_U1 ( .IN1(n4305), .IN2(U6470_n1), .QN(n4182) );
  INVX0 U6562_U2 ( .INP(n295), .ZN(U6562_n1) );
  NOR2X0 U6562_U1 ( .IN1(g3204), .IN2(U6562_n1), .QN(n3939) );
  INVX0 U6563_U2 ( .INP(n4073), .ZN(U6563_n1) );
  NOR2X0 U6563_U1 ( .IN1(g3204), .IN2(U6563_n1), .QN(n3705) );
  INVX0 U6718_U2 ( .INP(n296), .ZN(U6718_n1) );
  NOR2X0 U6718_U1 ( .IN1(g3197), .IN2(U6718_n1), .QN(n4073) );
  INVX0 U7116_U2 ( .INP(n4058), .ZN(U7116_n1) );
  NOR2X0 U7116_U1 ( .IN1(g2903), .IN2(U7116_n1), .QN(n4057) );
  INVX0 U7118_U2 ( .INP(n4123), .ZN(U7118_n1) );
  NOR2X0 U7118_U1 ( .IN1(g2896), .IN2(U7118_n1), .QN(n4122) );
  INVX0 U7293_U2 ( .INP(n4598), .ZN(U7293_n1) );
  NOR2X0 U7293_U1 ( .IN1(g3234), .IN2(U7293_n1), .QN(g20877) );
endmodule

