module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n445_, new_n236_, new_n238_, new_n479_, new_n250_, new_n501_, new_n288_, new_n421_, new_n368_, new_n439_, new_n283_, new_n223_, new_n390_, new_n366_, new_n241_, new_n186_, new_n365_, new_n339_, new_n197_, new_n386_, new_n401_, new_n389_, new_n514_, new_n456_, new_n246_, new_n170_, new_n266_, new_n173_, new_n220_, new_n419_, new_n214_, new_n489_, new_n424_, new_n114_, new_n188_, new_n240_, new_n413_, new_n442_, new_n211_, new_n123_, new_n127_, new_n342_, new_n462_, new_n500_, new_n344_, new_n287_, new_n504_, new_n427_, new_n234_, new_n472_, new_n393_, new_n418_, new_n292_, new_n215_, new_n152_, new_n157_, new_n153_, new_n133_, new_n257_, new_n481_, new_n212_, new_n364_, new_n449_, new_n484_, new_n272_, new_n282_, new_n201_, new_n192_, new_n414_, new_n110_, new_n315_, new_n124_, new_n164_, new_n230_, new_n281_, new_n248_, new_n117_, new_n167_, new_n385_, new_n478_, new_n461_, new_n297_, new_n361_, new_n150_, new_n108_, new_n137_, new_n183_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n180_, new_n318_, new_n321_, new_n443_, new_n324_, new_n158_, new_n486_, new_n491_, new_n466_, new_n262_, new_n271_, new_n274_, new_n218_, new_n497_, new_n305_, new_n420_, new_n498_, new_n205_, new_n492_, new_n141_, new_n206_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n506_, new_n256_, new_n452_, new_n381_, new_n388_, new_n508_, new_n194_, new_n483_, new_n394_, new_n116_, new_n299_, new_n142_, new_n139_, new_n314_, new_n118_, new_n363_, new_n165_, new_n441_, new_n216_, new_n280_, new_n426_, new_n235_, new_n398_, new_n301_, new_n169_, new_n395_, new_n383_, new_n210_, new_n458_, new_n447_, new_n207_, new_n267_, new_n473_, new_n140_, new_n187_, new_n311_, new_n263_, new_n331_, new_n341_, new_n378_, new_n349_, new_n244_, new_n172_, new_n488_, new_n277_, new_n402_, new_n286_, new_n335_, new_n347_, new_n346_, new_n396_, new_n198_, new_n438_, new_n208_, new_n179_, new_n436_, new_n397_, new_n399_, new_n233_, new_n469_, new_n391_, new_n178_, new_n295_, new_n359_, new_n132_, new_n166_, new_n162_, new_n409_, new_n457_, new_n161_, new_n333_, new_n290_, new_n448_, new_n276_, new_n155_, new_n384_, new_n410_, new_n113_, new_n509_, new_n454_, new_n202_, new_n296_, new_n232_, new_n258_, new_n176_, new_n156_, new_n494_, new_n291_, new_n261_, new_n309_, new_n323_, new_n259_, new_n227_, new_n416_, new_n222_, new_n400_, new_n328_, new_n130_, new_n505_, new_n471_, new_n268_, new_n374_, new_n376_, new_n380_, new_n138_, new_n310_, new_n144_, new_n275_, new_n352_, new_n485_, new_n126_, new_n177_, new_n493_, new_n264_, new_n379_, new_n273_, new_n224_, new_n270_, new_n143_, new_n520_, new_n125_, new_n145_, new_n253_, new_n403_, new_n475_, new_n237_, new_n149_, new_n260_, new_n251_, new_n189_, new_n300_, new_n106_, new_n411_, new_n507_, new_n107_, new_n182_, new_n407_, new_n480_, new_n151_, new_n513_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n428_, new_n199_, new_n146_, new_n302_, new_n191_, new_n225_, new_n387_, new_n476_, new_n112_, new_n121_, new_n415_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n131_, new_n255_, new_n459_, new_n174_, new_n468_, new_n354_, new_n392_, new_n518_, new_n340_, new_n147_, new_n285_, new_n209_, new_n337_, new_n446_, new_n203_, new_n316_, new_n417_, new_n515_, new_n332_, new_n453_, new_n163_, new_n519_, new_n148_, new_n440_, new_n122_, new_n111_, new_n252_, new_n160_, new_n312_, new_n372_, new_n242_, new_n503_, new_n115_, new_n307_, new_n190_, new_n408_, new_n213_, new_n134_, new_n433_, new_n435_, new_n109_, new_n265_, new_n370_, new_n278_, new_n304_, new_n217_, new_n269_, new_n512_, new_n129_, new_n412_, new_n327_, new_n495_, new_n431_, new_n196_, new_n319_, new_n338_, new_n377_, new_n247_, new_n330_, new_n375_, new_n294_, new_n195_, new_n357_, new_n320_, new_n245_, new_n474_, new_n467_, new_n404_, new_n193_, new_n490_, new_n128_, new_n348_, new_n159_, new_n322_, new_n228_, new_n289_, new_n425_, new_n175_, new_n226_, new_n185_, new_n171_, new_n434_, new_n200_, new_n422_, new_n329_, new_n249_, new_n136_, new_n284_, new_n119_, new_n293_, new_n168_, new_n279_, new_n455_, new_n120_, new_n406_, new_n229_, new_n464_, new_n204_, new_n181_, new_n135_, new_n405_;

xnor g000 ( new_n106_, N65, N69 );
xnor g001 ( new_n107_, N73, N77 );
xnor g002 ( new_n108_, new_n106_, new_n107_ );
xnor g003 ( new_n109_, N81, N85 );
xnor g004 ( new_n110_, N89, N93 );
xnor g005 ( new_n111_, new_n109_, new_n110_ );
xnor g006 ( new_n112_, new_n108_, new_n111_ );
nand g007 ( new_n113_, N129, N137 );
xnor g008 ( new_n114_, new_n112_, new_n113_ );
xor g009 ( new_n115_, N1, N17 );
xnor g010 ( new_n116_, N33, N49 );
xnor g011 ( new_n117_, new_n115_, new_n116_ );
xnor g012 ( new_n118_, new_n117_, keyIn_0_9 );
xnor g013 ( new_n119_, new_n114_, new_n118_ );
not g014 ( new_n120_, new_n119_ );
xnor g015 ( new_n121_, N97, N101 );
xnor g016 ( new_n122_, new_n121_, keyIn_0_3 );
xnor g017 ( new_n123_, N105, N109 );
xnor g018 ( new_n124_, new_n122_, new_n123_ );
xnor g019 ( new_n125_, N121, N125 );
xnor g020 ( new_n126_, new_n125_, keyIn_0_4 );
xnor g021 ( new_n127_, N113, N117 );
xnor g022 ( new_n128_, new_n126_, new_n127_ );
xor g023 ( new_n129_, new_n124_, new_n128_ );
nand g024 ( new_n130_, N130, N137 );
nand g025 ( new_n131_, new_n129_, new_n130_ );
xnor g026 ( new_n132_, new_n124_, new_n128_ );
nand g027 ( new_n133_, new_n132_, N130, N137 );
nand g028 ( new_n134_, new_n131_, new_n133_ );
xnor g029 ( new_n135_, N5, N21 );
xnor g030 ( new_n136_, N37, N53 );
xnor g031 ( new_n137_, new_n135_, new_n136_ );
not g032 ( new_n138_, new_n137_ );
nand g033 ( new_n139_, new_n134_, new_n138_ );
nand g034 ( new_n140_, new_n131_, new_n133_, new_n137_ );
nand g035 ( new_n141_, new_n139_, new_n140_ );
xnor g036 ( new_n142_, new_n124_, new_n108_ );
nand g037 ( new_n143_, new_n142_, N131, N137 );
not g038 ( new_n144_, new_n108_ );
xnor g039 ( new_n145_, new_n124_, new_n144_ );
nand g040 ( new_n146_, N131, N137 );
nand g041 ( new_n147_, new_n145_, new_n146_ );
nand g042 ( new_n148_, new_n143_, new_n147_ );
xor g043 ( new_n149_, N41, N57 );
xnor g044 ( new_n150_, new_n149_, keyIn_0_6 );
xor g045 ( new_n151_, N9, N25 );
xnor g046 ( new_n152_, new_n150_, new_n151_ );
not g047 ( new_n153_, new_n152_ );
nand g048 ( new_n154_, new_n148_, new_n153_ );
nand g049 ( new_n155_, new_n143_, new_n147_, new_n152_ );
nand g050 ( new_n156_, new_n154_, new_n155_ );
not g051 ( new_n157_, new_n156_ );
nand g052 ( new_n158_, new_n157_, new_n141_, keyIn_0_12 );
nand g053 ( new_n159_, new_n154_, keyIn_0_12, new_n155_ );
nand g054 ( new_n160_, new_n159_, new_n139_, new_n140_ );
nand g055 ( new_n161_, new_n158_, new_n120_, new_n160_ );
nand g056 ( new_n162_, new_n141_, keyIn_0_13 );
not g057 ( new_n163_, keyIn_0_13 );
nand g058 ( new_n164_, new_n139_, new_n163_, new_n140_ );
nand g059 ( new_n165_, new_n162_, new_n164_ );
nand g060 ( new_n166_, new_n156_, new_n119_ );
not g061 ( new_n167_, new_n166_ );
nand g062 ( new_n168_, new_n165_, new_n167_ );
nand g063 ( new_n169_, new_n168_, new_n161_ );
not g064 ( new_n170_, new_n111_ );
xnor g065 ( new_n171_, new_n128_, new_n170_ );
nand g066 ( new_n172_, N132, N137 );
xnor g067 ( new_n173_, new_n171_, new_n172_ );
xnor g068 ( new_n174_, N13, N29 );
xnor g069 ( new_n175_, N45, N61 );
xnor g070 ( new_n176_, new_n174_, new_n175_ );
not g071 ( new_n177_, new_n176_ );
xnor g072 ( new_n178_, new_n173_, new_n177_ );
not g073 ( new_n179_, new_n178_ );
nand g074 ( new_n180_, new_n169_, new_n179_ );
not g075 ( new_n181_, new_n141_ );
not g076 ( new_n182_, keyIn_0_11 );
xnor g077 ( new_n183_, new_n119_, new_n182_ );
nand g078 ( new_n184_, new_n183_, new_n181_, new_n156_, new_n178_ );
xnor g079 ( new_n185_, new_n184_, keyIn_0_19 );
nand g080 ( new_n186_, new_n185_, new_n180_ );
not g081 ( new_n187_, keyIn_0_8 );
nand g082 ( new_n188_, N33, N37 );
not g083 ( new_n189_, N33 );
not g084 ( new_n190_, N37 );
nand g085 ( new_n191_, new_n189_, new_n190_ );
nand g086 ( new_n192_, new_n191_, new_n188_ );
nand g087 ( new_n193_, new_n192_, keyIn_0_1 );
not g088 ( new_n194_, keyIn_0_1 );
nand g089 ( new_n195_, new_n191_, new_n194_, new_n188_ );
xnor g090 ( new_n196_, N41, N45 );
nand g091 ( new_n197_, new_n196_, keyIn_0_2 );
not g092 ( new_n198_, keyIn_0_2 );
nand g093 ( new_n199_, N41, N45 );
not g094 ( new_n200_, N41 );
not g095 ( new_n201_, N45 );
nand g096 ( new_n202_, new_n200_, new_n201_ );
nand g097 ( new_n203_, new_n202_, new_n198_, new_n199_ );
nand g098 ( new_n204_, new_n193_, new_n197_, new_n195_, new_n203_ );
nand g099 ( new_n205_, new_n193_, new_n195_ );
nand g100 ( new_n206_, new_n197_, new_n203_ );
nand g101 ( new_n207_, new_n205_, new_n206_ );
nand g102 ( new_n208_, new_n207_, new_n204_ );
nand g103 ( new_n209_, new_n208_, new_n187_ );
nand g104 ( new_n210_, new_n207_, keyIn_0_8, new_n204_ );
nand g105 ( new_n211_, new_n209_, new_n210_ );
xnor g106 ( new_n212_, N49, N53 );
xnor g107 ( new_n213_, N57, N61 );
xnor g108 ( new_n214_, new_n212_, new_n213_ );
not g109 ( new_n215_, new_n214_ );
nand g110 ( new_n216_, new_n211_, new_n215_ );
nand g111 ( new_n217_, new_n209_, new_n210_, new_n214_ );
nand g112 ( new_n218_, new_n216_, new_n217_ );
nand g113 ( new_n219_, N134, N137 );
nand g114 ( new_n220_, new_n218_, new_n219_ );
nand g115 ( new_n221_, new_n216_, N134, N137, new_n217_ );
nand g116 ( new_n222_, new_n220_, new_n221_ );
xnor g117 ( new_n223_, N69, N85 );
xnor g118 ( new_n224_, N101, N117 );
xnor g119 ( new_n225_, new_n223_, new_n224_ );
nand g120 ( new_n226_, new_n222_, new_n225_ );
not g121 ( new_n227_, new_n225_ );
nand g122 ( new_n228_, new_n220_, new_n221_, new_n227_ );
nand g123 ( new_n229_, new_n226_, new_n228_ );
not g124 ( new_n230_, new_n229_ );
nand g125 ( new_n231_, new_n230_, keyIn_0_14 );
not g126 ( new_n232_, keyIn_0_14 );
nand g127 ( new_n233_, new_n229_, new_n232_ );
xnor g128 ( new_n234_, N1, N5 );
xnor g129 ( new_n235_, N9, N13 );
xnor g130 ( new_n236_, new_n234_, new_n235_ );
xor g131 ( new_n237_, N17, N21 );
nand g132 ( new_n238_, N25, N29 );
not g133 ( new_n239_, N25 );
not g134 ( new_n240_, N29 );
nand g135 ( new_n241_, new_n239_, new_n240_ );
nand g136 ( new_n242_, new_n241_, new_n238_ );
nand g137 ( new_n243_, new_n242_, keyIn_0_0 );
not g138 ( new_n244_, keyIn_0_0 );
nand g139 ( new_n245_, new_n241_, new_n244_, new_n238_ );
nand g140 ( new_n246_, new_n243_, new_n237_, new_n245_ );
not g141 ( new_n247_, new_n237_ );
nand g142 ( new_n248_, new_n243_, new_n245_ );
nand g143 ( new_n249_, new_n248_, new_n247_ );
nand g144 ( new_n250_, new_n249_, new_n246_ );
xnor g145 ( new_n251_, new_n250_, new_n236_ );
nand g146 ( new_n252_, N133, N137 );
xnor g147 ( new_n253_, new_n251_, new_n252_ );
xnor g148 ( new_n254_, N65, N81 );
xnor g149 ( new_n255_, N97, N113 );
xnor g150 ( new_n256_, new_n254_, new_n255_ );
xnor g151 ( new_n257_, new_n253_, new_n256_ );
not g152 ( new_n258_, new_n257_ );
nand g153 ( new_n259_, new_n231_, new_n233_, new_n258_ );
nand g154 ( new_n260_, new_n250_, new_n215_ );
nand g155 ( new_n261_, new_n249_, new_n214_, new_n246_ );
nand g156 ( new_n262_, new_n260_, new_n261_ );
nand g157 ( new_n263_, N136, N137 );
nand g158 ( new_n264_, new_n262_, new_n263_ );
nand g159 ( new_n265_, new_n260_, N136, N137, new_n261_ );
nand g160 ( new_n266_, new_n264_, new_n265_ );
nand g161 ( new_n267_, new_n266_, keyIn_0_10 );
not g162 ( new_n268_, keyIn_0_10 );
nand g163 ( new_n269_, new_n264_, new_n268_, new_n265_ );
nand g164 ( new_n270_, new_n267_, new_n269_ );
xnor g165 ( new_n271_, N77, N93 );
xnor g166 ( new_n272_, N109, N125 );
xnor g167 ( new_n273_, new_n271_, new_n272_ );
not g168 ( new_n274_, new_n273_ );
nand g169 ( new_n275_, new_n270_, new_n274_ );
nand g170 ( new_n276_, new_n267_, new_n269_, new_n273_ );
nand g171 ( new_n277_, new_n275_, new_n276_ );
xnor g172 ( new_n278_, new_n277_, keyIn_0_15 );
not g173 ( new_n279_, keyIn_0_5 );
not g174 ( new_n280_, new_n236_ );
nand g175 ( new_n281_, new_n211_, new_n280_ );
nand g176 ( new_n282_, new_n209_, new_n210_, new_n236_ );
nand g177 ( new_n283_, new_n281_, new_n279_, new_n282_ );
nand g178 ( new_n284_, new_n281_, new_n282_ );
nand g179 ( new_n285_, new_n284_, keyIn_0_5 );
nand g180 ( new_n286_, new_n285_, N135, N137, new_n283_ );
nand g181 ( new_n287_, N135, N137 );
nand g182 ( new_n288_, new_n285_, new_n283_ );
nand g183 ( new_n289_, new_n288_, new_n287_ );
xor g184 ( new_n290_, N105, N121 );
xnor g185 ( new_n291_, new_n290_, keyIn_0_7 );
xnor g186 ( new_n292_, N73, N89 );
xnor g187 ( new_n293_, new_n291_, new_n292_ );
not g188 ( new_n294_, new_n293_ );
nand g189 ( new_n295_, new_n289_, new_n286_, new_n294_ );
nand g190 ( new_n296_, new_n289_, new_n286_ );
nand g191 ( new_n297_, new_n296_, new_n293_ );
nand g192 ( new_n298_, new_n297_, new_n295_ );
nor g193 ( new_n299_, new_n259_, new_n278_, new_n298_ );
nand g194 ( new_n300_, new_n186_, new_n299_ );
nand g195 ( new_n301_, new_n300_, keyIn_0_24 );
not g196 ( new_n302_, keyIn_0_24 );
nand g197 ( new_n303_, new_n186_, new_n302_, new_n299_ );
nand g198 ( new_n304_, new_n301_, new_n303_ );
nand g199 ( new_n305_, new_n304_, new_n119_ );
xnor g200 ( N724, new_n305_, N1 );
nand g201 ( new_n307_, new_n304_, new_n141_ );
xnor g202 ( N725, new_n307_, N5 );
nand g203 ( new_n309_, new_n304_, new_n157_ );
nand g204 ( new_n310_, new_n309_, N9 );
not g205 ( new_n311_, N9 );
nand g206 ( new_n312_, new_n304_, new_n311_, new_n157_ );
nand g207 ( new_n313_, new_n310_, new_n312_ );
nand g208 ( new_n314_, new_n313_, keyIn_0_30 );
not g209 ( new_n315_, keyIn_0_30 );
nand g210 ( new_n316_, new_n310_, new_n315_, new_n312_ );
nand g211 ( N726, new_n314_, new_n316_ );
nand g212 ( new_n318_, new_n304_, new_n178_ );
nand g213 ( new_n319_, new_n318_, N13 );
not g214 ( new_n320_, N13 );
nand g215 ( new_n321_, new_n304_, new_n320_, new_n178_ );
nand g216 ( new_n322_, new_n319_, new_n321_ );
nand g217 ( new_n323_, new_n322_, keyIn_0_31 );
not g218 ( new_n324_, keyIn_0_31 );
nand g219 ( new_n325_, new_n319_, new_n324_, new_n321_ );
nand g220 ( N727, new_n323_, new_n325_ );
nand g221 ( new_n327_, new_n186_, new_n277_ );
not g222 ( new_n328_, new_n327_ );
nand g223 ( new_n329_, new_n298_, new_n229_, new_n258_ );
not g224 ( new_n330_, new_n329_ );
nand g225 ( new_n331_, new_n328_, new_n330_ );
not g226 ( new_n332_, new_n331_ );
nand g227 ( new_n333_, new_n332_, new_n119_ );
xnor g228 ( N728, new_n333_, N17 );
nand g229 ( new_n335_, new_n332_, new_n141_ );
xnor g230 ( N729, new_n335_, N21 );
nand g231 ( new_n337_, new_n328_, new_n157_, new_n330_ );
xnor g232 ( new_n338_, new_n337_, keyIn_0_25 );
nand g233 ( new_n339_, new_n338_, new_n239_ );
not g234 ( new_n340_, keyIn_0_25 );
xnor g235 ( new_n341_, new_n337_, new_n340_ );
nand g236 ( new_n342_, new_n341_, N25 );
nand g237 ( N730, new_n339_, new_n342_ );
nand g238 ( new_n344_, new_n328_, new_n178_, new_n330_ );
xnor g239 ( new_n345_, new_n344_, keyIn_0_26 );
nand g240 ( new_n346_, new_n345_, N29 );
not g241 ( new_n347_, keyIn_0_26 );
xnor g242 ( new_n348_, new_n344_, new_n347_ );
nand g243 ( new_n349_, new_n348_, new_n240_ );
nand g244 ( N731, new_n346_, new_n349_ );
xor g245 ( new_n351_, new_n257_, keyIn_0_16 );
nor g246 ( new_n352_, new_n351_, new_n229_, new_n298_, new_n277_ );
nand g247 ( new_n353_, new_n186_, new_n352_ );
not g248 ( new_n354_, new_n353_ );
nand g249 ( new_n355_, new_n354_, new_n119_ );
xnor g250 ( N732, new_n355_, N33 );
nand g251 ( new_n357_, new_n354_, new_n141_ );
xnor g252 ( N733, new_n357_, N37 );
nand g253 ( new_n359_, new_n354_, new_n157_ );
xnor g254 ( N734, new_n359_, N41 );
nand g255 ( new_n361_, new_n354_, new_n178_ );
xnor g256 ( N735, new_n361_, N45 );
xor g257 ( new_n363_, new_n257_, keyIn_0_17 );
nand g258 ( new_n364_, new_n328_, new_n230_, new_n298_, new_n363_ );
not g259 ( new_n365_, new_n364_ );
nand g260 ( new_n366_, new_n365_, new_n119_ );
xnor g261 ( N736, new_n366_, N49 );
nand g262 ( new_n368_, new_n365_, new_n141_ );
xnor g263 ( N737, new_n368_, N53 );
nand g264 ( new_n370_, new_n365_, new_n157_ );
xnor g265 ( N738, new_n370_, N57 );
nand g266 ( new_n372_, new_n365_, new_n178_ );
xnor g267 ( N739, new_n372_, N61 );
not g268 ( new_n374_, N65 );
xnor g269 ( new_n375_, new_n270_, new_n273_ );
nand g270 ( new_n376_, new_n375_, new_n257_ );
not g271 ( new_n377_, new_n376_ );
nand g272 ( new_n378_, new_n377_, new_n230_, new_n298_ );
nand g273 ( new_n379_, new_n378_, keyIn_0_22 );
not g274 ( new_n380_, keyIn_0_22 );
nand g275 ( new_n381_, new_n377_, new_n380_, new_n298_, new_n230_ );
nand g276 ( new_n382_, new_n298_, new_n230_ );
nand g277 ( new_n383_, new_n382_, keyIn_0_22 );
nand g278 ( new_n384_, new_n379_, new_n381_, new_n383_ );
nand g279 ( new_n385_, new_n277_, new_n257_ );
not g280 ( new_n386_, new_n385_ );
nand g281 ( new_n387_, new_n298_, new_n229_, new_n386_ );
xnor g282 ( new_n388_, new_n387_, keyIn_0_20 );
nand g283 ( new_n389_, new_n229_, new_n257_ );
not g284 ( new_n390_, new_n389_ );
nand g285 ( new_n391_, new_n390_, new_n375_, new_n295_, new_n297_ );
nand g286 ( new_n392_, new_n391_, keyIn_0_21 );
not g287 ( new_n393_, keyIn_0_21 );
xnor g288 ( new_n394_, new_n296_, new_n294_ );
nand g289 ( new_n395_, new_n394_, new_n393_, new_n375_, new_n390_ );
nand g290 ( new_n396_, new_n392_, new_n395_ );
not g291 ( new_n397_, keyIn_0_23 );
not g292 ( new_n398_, keyIn_0_18 );
nand g293 ( new_n399_, new_n297_, new_n398_, new_n295_ );
nand g294 ( new_n400_, new_n298_, keyIn_0_18 );
nand g295 ( new_n401_, new_n400_, new_n399_ );
nor g296 ( new_n402_, new_n230_, new_n257_, new_n277_ );
nand g297 ( new_n403_, new_n401_, new_n402_ );
nand g298 ( new_n404_, new_n403_, new_n397_ );
not g299 ( new_n405_, new_n404_ );
nand g300 ( new_n406_, new_n405_, new_n384_, new_n388_, new_n396_ );
nand g301 ( new_n407_, new_n379_, new_n381_ );
nand g302 ( new_n408_, new_n387_, keyIn_0_20 );
not g303 ( new_n409_, keyIn_0_20 );
nand g304 ( new_n410_, new_n298_, new_n390_, new_n409_, new_n277_ );
nand g305 ( new_n411_, new_n408_, new_n410_ );
nand g306 ( new_n412_, new_n407_, new_n411_, new_n396_, new_n403_ );
nand g307 ( new_n413_, new_n412_, keyIn_0_23 );
nand g308 ( new_n414_, new_n406_, new_n413_ );
nand g309 ( new_n415_, new_n414_, new_n258_ );
not g310 ( new_n416_, new_n415_ );
nand g311 ( new_n417_, new_n179_, new_n157_ );
nand g312 ( new_n418_, new_n181_, new_n119_ );
nor g313 ( new_n419_, new_n417_, new_n418_ );
nand g314 ( new_n420_, new_n416_, new_n374_, new_n419_ );
nand g315 ( new_n421_, new_n416_, new_n419_ );
nand g316 ( new_n422_, new_n421_, N65 );
nand g317 ( N740, new_n422_, new_n420_ );
not g318 ( new_n424_, N69 );
nand g319 ( new_n425_, new_n414_, new_n230_ );
not g320 ( new_n426_, new_n425_ );
nand g321 ( new_n427_, new_n426_, new_n424_, new_n419_ );
nand g322 ( new_n428_, new_n426_, new_n419_ );
nand g323 ( new_n429_, new_n428_, N69 );
nand g324 ( N741, new_n429_, new_n427_ );
not g325 ( new_n431_, N73 );
nand g326 ( new_n432_, new_n414_, new_n394_ );
not g327 ( new_n433_, new_n432_ );
nand g328 ( new_n434_, new_n433_, new_n431_, new_n419_ );
nand g329 ( new_n435_, new_n433_, new_n419_ );
nand g330 ( new_n436_, new_n435_, N73 );
nand g331 ( N742, new_n436_, new_n434_ );
not g332 ( new_n438_, N77 );
nand g333 ( new_n439_, new_n414_, new_n277_ );
not g334 ( new_n440_, new_n439_ );
nand g335 ( new_n441_, new_n440_, new_n438_, new_n419_ );
nand g336 ( new_n442_, new_n440_, new_n419_ );
nand g337 ( new_n443_, new_n442_, N77 );
nand g338 ( N743, new_n443_, new_n441_ );
not g339 ( new_n445_, N81 );
nand g340 ( new_n446_, new_n178_, new_n156_ );
nor g341 ( new_n447_, new_n418_, new_n446_ );
nand g342 ( new_n448_, new_n416_, new_n445_, new_n447_ );
nand g343 ( new_n449_, new_n416_, new_n447_ );
nand g344 ( new_n450_, new_n449_, N81 );
nand g345 ( N744, new_n450_, new_n448_ );
nand g346 ( new_n452_, new_n414_, new_n230_, new_n447_ );
nand g347 ( new_n453_, new_n452_, keyIn_0_27 );
not g348 ( new_n454_, keyIn_0_27 );
nand g349 ( new_n455_, new_n414_, new_n454_, new_n230_, new_n447_ );
nand g350 ( new_n456_, new_n453_, new_n455_ );
nand g351 ( new_n457_, new_n456_, N85 );
not g352 ( new_n458_, N85 );
nand g353 ( new_n459_, new_n453_, new_n458_, new_n455_ );
nand g354 ( N745, new_n457_, new_n459_ );
not g355 ( new_n461_, N89 );
nand g356 ( new_n462_, new_n433_, new_n461_, new_n447_ );
nand g357 ( new_n463_, new_n433_, new_n447_ );
nand g358 ( new_n464_, new_n463_, N89 );
nand g359 ( N746, new_n464_, new_n462_ );
nand g360 ( new_n466_, new_n440_, new_n447_ );
nand g361 ( new_n467_, new_n466_, N93 );
not g362 ( new_n468_, N93 );
nand g363 ( new_n469_, new_n440_, new_n468_, new_n447_ );
nand g364 ( N747, new_n467_, new_n469_ );
not g365 ( new_n471_, N97 );
nand g366 ( new_n472_, new_n141_, new_n120_ );
nor g367 ( new_n473_, new_n417_, new_n472_ );
nand g368 ( new_n474_, new_n416_, new_n471_, new_n473_ );
nand g369 ( new_n475_, new_n416_, new_n473_ );
nand g370 ( new_n476_, new_n475_, N97 );
nand g371 ( N748, new_n476_, new_n474_ );
nand g372 ( new_n478_, new_n426_, new_n473_ );
nand g373 ( new_n479_, new_n478_, N101 );
not g374 ( new_n480_, N101 );
nand g375 ( new_n481_, new_n426_, new_n480_, new_n473_ );
nand g376 ( N749, new_n479_, new_n481_ );
not g377 ( new_n483_, N105 );
nand g378 ( new_n484_, new_n433_, new_n483_, new_n473_ );
nand g379 ( new_n485_, new_n433_, new_n473_ );
nand g380 ( new_n486_, new_n485_, N105 );
nand g381 ( N750, new_n486_, new_n484_ );
not g382 ( new_n488_, keyIn_0_28 );
nand g383 ( new_n489_, new_n414_, new_n277_, new_n473_ );
nand g384 ( new_n490_, new_n489_, new_n488_ );
nand g385 ( new_n491_, new_n414_, keyIn_0_28, new_n277_, new_n473_ );
nand g386 ( new_n492_, new_n490_, new_n491_ );
nand g387 ( new_n493_, new_n492_, N109 );
not g388 ( new_n494_, N109 );
nand g389 ( new_n495_, new_n490_, new_n494_, new_n491_ );
nand g390 ( N751, new_n493_, new_n495_ );
not g391 ( new_n497_, N113 );
nor g392 ( new_n498_, new_n446_, new_n472_ );
nand g393 ( new_n499_, new_n416_, new_n497_, new_n498_ );
nand g394 ( new_n500_, new_n416_, new_n498_ );
nand g395 ( new_n501_, new_n500_, N113 );
nand g396 ( N752, new_n501_, new_n499_ );
not g397 ( new_n503_, N117 );
not g398 ( new_n504_, keyIn_0_29 );
nand g399 ( new_n505_, new_n414_, new_n230_, new_n498_ );
nand g400 ( new_n506_, new_n505_, new_n504_ );
nand g401 ( new_n507_, new_n414_, keyIn_0_29, new_n230_, new_n498_ );
nand g402 ( new_n508_, new_n506_, new_n507_ );
nand g403 ( new_n509_, new_n508_, new_n503_ );
nand g404 ( new_n510_, new_n506_, N117, new_n507_ );
nand g405 ( N753, new_n509_, new_n510_ );
not g406 ( new_n512_, N121 );
nand g407 ( new_n513_, new_n433_, new_n512_, new_n498_ );
nand g408 ( new_n514_, new_n433_, new_n498_ );
nand g409 ( new_n515_, new_n514_, N121 );
nand g410 ( N754, new_n515_, new_n513_ );
nand g411 ( new_n517_, new_n440_, new_n498_ );
nand g412 ( new_n518_, new_n517_, N125 );
not g413 ( new_n519_, N125 );
nand g414 ( new_n520_, new_n440_, new_n519_, new_n498_ );
nand g415 ( N755, new_n518_, new_n520_ );
endmodule