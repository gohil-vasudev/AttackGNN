module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n359_, new_n368_, new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n381_, new_n382_, new_n385_, new_n386_, new_n388_, new_n390_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n401_, new_n402_, new_n403_, new_n404_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n520_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n571_, new_n572_, new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_;
  XOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .Z(new_n359_) );
  INV_X1 g001 ( .A(new_n359_), .ZN(G218) );
  INV_X1 g002 ( .A(G132), .ZN(G219) );
  INV_X1 g003 ( .A(G82), .ZN(G220) );
  INV_X1 g004 ( .A(G96), .ZN(G221) );
  INV_X1 g005 ( .A(G69), .ZN(G235) );
  INV_X1 g006 ( .A(G120), .ZN(G236) );
  INV_X1 g007 ( .A(G57), .ZN(G237) );
  INV_X1 g008 ( .A(G108), .ZN(G238) );
  INV_X1 g009 ( .A(KEYINPUT20), .ZN(new_n368_) );
  AND2_X1 g010 ( .A1(G2078), .A2(G2084), .ZN(new_n369_) );
  AND2_X1 g011 ( .A1(new_n369_), .A2(new_n368_), .ZN(new_n370_) );
  INV_X1 g012 ( .A(new_n370_), .ZN(new_n371_) );
  OR2_X1 g013 ( .A1(new_n369_), .A2(new_n368_), .ZN(new_n372_) );
  AND2_X1 g014 ( .A1(new_n372_), .A2(G2090), .ZN(new_n373_) );
  AND2_X1 g015 ( .A1(new_n373_), .A2(new_n371_), .ZN(new_n374_) );
  AND2_X1 g016 ( .A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n375_) );
  INV_X1 g017 ( .A(new_n375_), .ZN(new_n376_) );
  OR2_X1 g018 ( .A1(new_n374_), .A2(KEYINPUT21), .ZN(new_n377_) );
  AND2_X1 g019 ( .A1(new_n377_), .A2(G2072), .ZN(new_n378_) );
  AND2_X1 g020 ( .A1(new_n378_), .A2(new_n376_), .ZN(new_n379_) );
  INV_X1 g021 ( .A(new_n379_), .ZN(G158) );
  AND2_X1 g022 ( .A1(G2), .A2(G15), .ZN(new_n381_) );
  AND2_X1 g023 ( .A1(new_n381_), .A2(G661), .ZN(new_n382_) );
  INV_X1 g024 ( .A(new_n382_), .ZN(G259) );
  AND2_X1 g025 ( .A1(G94), .A2(G452), .ZN(G173) );
  AND2_X1 g026 ( .A1(G7), .A2(G661), .ZN(new_n385_) );
  XNOR2_X1 g027 ( .A(new_n385_), .B(KEYINPUT10), .ZN(new_n386_) );
  INV_X1 g028 ( .A(new_n386_), .ZN(G223) );
  AND2_X1 g029 ( .A1(new_n386_), .A2(G567), .ZN(new_n388_) );
  XNOR2_X1 g030 ( .A(new_n388_), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 g031 ( .A(G2106), .ZN(new_n390_) );
  OR2_X1 g032 ( .A1(G223), .A2(new_n390_), .ZN(G217) );
  AND2_X1 g033 ( .A1(new_n359_), .A2(G96), .ZN(new_n392_) );
  AND2_X1 g034 ( .A1(G82), .A2(G132), .ZN(new_n393_) );
  XNOR2_X1 g035 ( .A(new_n393_), .B(KEYINPUT22), .ZN(new_n394_) );
  AND2_X1 g036 ( .A1(new_n392_), .A2(new_n394_), .ZN(new_n395_) );
  AND2_X1 g037 ( .A1(G57), .A2(G69), .ZN(new_n396_) );
  AND2_X1 g038 ( .A1(G108), .A2(G120), .ZN(new_n397_) );
  AND2_X1 g039 ( .A1(new_n396_), .A2(new_n397_), .ZN(new_n398_) );
  AND2_X1 g040 ( .A1(new_n395_), .A2(new_n398_), .ZN(G325) );
  INV_X1 g041 ( .A(G325), .ZN(G261) );
  OR2_X1 g042 ( .A1(new_n395_), .A2(new_n390_), .ZN(new_n401_) );
  INV_X1 g043 ( .A(new_n398_), .ZN(new_n402_) );
  AND2_X1 g044 ( .A1(new_n402_), .A2(G567), .ZN(new_n403_) );
  INV_X1 g045 ( .A(new_n403_), .ZN(new_n404_) );
  AND2_X1 g046 ( .A1(new_n401_), .A2(new_n404_), .ZN(G319) );
  INV_X1 g047 ( .A(G2105), .ZN(new_n406_) );
  AND2_X1 g048 ( .A1(G101), .A2(G2104), .ZN(new_n407_) );
  AND2_X1 g049 ( .A1(new_n407_), .A2(new_n406_), .ZN(new_n408_) );
  XNOR2_X1 g050 ( .A(new_n408_), .B(KEYINPUT23), .ZN(new_n409_) );
  INV_X1 g051 ( .A(G137), .ZN(new_n410_) );
  OR2_X1 g052 ( .A1(G2104), .A2(G2105), .ZN(new_n411_) );
  XNOR2_X1 g053 ( .A(new_n411_), .B(KEYINPUT17), .ZN(new_n412_) );
  INV_X1 g054 ( .A(new_n412_), .ZN(new_n413_) );
  OR2_X1 g055 ( .A1(new_n413_), .A2(new_n410_), .ZN(new_n414_) );
  AND2_X1 g056 ( .A1(new_n414_), .A2(new_n409_), .ZN(new_n415_) );
  INV_X1 g057 ( .A(G125), .ZN(new_n416_) );
  OR2_X1 g058 ( .A1(new_n416_), .A2(G2104), .ZN(new_n417_) );
  OR2_X1 g059 ( .A1(new_n417_), .A2(new_n406_), .ZN(new_n418_) );
  AND2_X1 g060 ( .A1(G113), .A2(G2104), .ZN(new_n419_) );
  AND2_X1 g061 ( .A1(new_n419_), .A2(G2105), .ZN(new_n420_) );
  INV_X1 g062 ( .A(new_n420_), .ZN(new_n421_) );
  AND2_X1 g063 ( .A1(new_n418_), .A2(new_n421_), .ZN(new_n422_) );
  AND2_X1 g064 ( .A1(new_n415_), .A2(new_n422_), .ZN(G160) );
  INV_X1 g065 ( .A(G136), .ZN(new_n424_) );
  OR2_X1 g066 ( .A1(new_n413_), .A2(new_n424_), .ZN(new_n425_) );
  INV_X1 g067 ( .A(G2104), .ZN(new_n426_) );
  AND2_X1 g068 ( .A1(new_n426_), .A2(G2105), .ZN(new_n427_) );
  AND2_X1 g069 ( .A1(new_n427_), .A2(G124), .ZN(new_n428_) );
  OR2_X1 g070 ( .A1(new_n428_), .A2(KEYINPUT44), .ZN(new_n429_) );
  INV_X1 g071 ( .A(KEYINPUT44), .ZN(new_n430_) );
  INV_X1 g072 ( .A(new_n428_), .ZN(new_n431_) );
  OR2_X1 g073 ( .A1(new_n431_), .A2(new_n430_), .ZN(new_n432_) );
  AND2_X1 g074 ( .A1(G2104), .A2(G2105), .ZN(new_n433_) );
  AND2_X1 g075 ( .A1(new_n433_), .A2(G112), .ZN(new_n434_) );
  INV_X1 g076 ( .A(new_n434_), .ZN(new_n435_) );
  INV_X1 g077 ( .A(G100), .ZN(new_n436_) );
  AND2_X1 g078 ( .A1(new_n406_), .A2(G2104), .ZN(new_n437_) );
  INV_X1 g079 ( .A(new_n437_), .ZN(new_n438_) );
  OR2_X1 g080 ( .A1(new_n438_), .A2(new_n436_), .ZN(new_n439_) );
  AND2_X1 g081 ( .A1(new_n439_), .A2(new_n435_), .ZN(new_n440_) );
  AND2_X1 g082 ( .A1(new_n432_), .A2(new_n440_), .ZN(new_n441_) );
  AND2_X1 g083 ( .A1(new_n441_), .A2(new_n429_), .ZN(new_n442_) );
  AND2_X1 g084 ( .A1(new_n442_), .A2(new_n425_), .ZN(G162) );
  AND2_X1 g085 ( .A1(new_n412_), .A2(G138), .ZN(new_n444_) );
  AND2_X1 g086 ( .A1(new_n433_), .A2(G114), .ZN(new_n445_) );
  AND2_X1 g087 ( .A1(G102), .A2(G2104), .ZN(new_n446_) );
  AND2_X1 g088 ( .A1(new_n446_), .A2(new_n406_), .ZN(new_n447_) );
  AND2_X1 g089 ( .A1(new_n427_), .A2(G126), .ZN(new_n448_) );
  OR2_X1 g090 ( .A1(new_n448_), .A2(new_n447_), .ZN(new_n449_) );
  OR2_X1 g091 ( .A1(new_n449_), .A2(new_n445_), .ZN(new_n450_) );
  OR2_X1 g092 ( .A1(new_n450_), .A2(new_n444_), .ZN(new_n451_) );
  INV_X1 g093 ( .A(new_n451_), .ZN(G164) );
  OR2_X1 g094 ( .A1(G543), .A2(G651), .ZN(new_n453_) );
  INV_X1 g095 ( .A(new_n453_), .ZN(new_n454_) );
  AND2_X1 g096 ( .A1(new_n454_), .A2(G88), .ZN(new_n455_) );
  XNOR2_X1 g097 ( .A(G543), .B(KEYINPUT0), .ZN(new_n456_) );
  AND2_X1 g098 ( .A1(new_n456_), .A2(G651), .ZN(new_n457_) );
  AND2_X1 g099 ( .A1(new_n457_), .A2(G75), .ZN(new_n458_) );
  OR2_X1 g100 ( .A1(new_n458_), .A2(new_n455_), .ZN(new_n459_) );
  INV_X1 g101 ( .A(G543), .ZN(new_n460_) );
  AND2_X1 g102 ( .A1(new_n460_), .A2(G651), .ZN(new_n461_) );
  XNOR2_X1 g103 ( .A(new_n461_), .B(KEYINPUT1), .ZN(new_n462_) );
  INV_X1 g104 ( .A(new_n462_), .ZN(new_n463_) );
  AND2_X1 g105 ( .A1(new_n463_), .A2(G62), .ZN(new_n464_) );
  INV_X1 g106 ( .A(G651), .ZN(new_n465_) );
  AND2_X1 g107 ( .A1(new_n456_), .A2(new_n465_), .ZN(new_n466_) );
  AND2_X1 g108 ( .A1(new_n466_), .A2(G50), .ZN(new_n467_) );
  OR2_X1 g109 ( .A1(new_n464_), .A2(new_n467_), .ZN(new_n468_) );
  OR2_X1 g110 ( .A1(new_n468_), .A2(new_n459_), .ZN(G303) );
  INV_X1 g111 ( .A(G303), .ZN(G166) );
  AND2_X1 g112 ( .A1(new_n466_), .A2(G51), .ZN(new_n471_) );
  AND2_X1 g113 ( .A1(new_n463_), .A2(G63), .ZN(new_n472_) );
  OR2_X1 g114 ( .A1(new_n472_), .A2(new_n471_), .ZN(new_n473_) );
  XOR2_X1 g115 ( .A(new_n473_), .B(KEYINPUT6), .Z(new_n474_) );
  AND2_X1 g116 ( .A1(new_n457_), .A2(G76), .ZN(new_n475_) );
  AND2_X1 g117 ( .A1(new_n454_), .A2(G89), .ZN(new_n476_) );
  XNOR2_X1 g118 ( .A(new_n476_), .B(KEYINPUT4), .ZN(new_n477_) );
  OR2_X1 g119 ( .A1(new_n477_), .A2(new_n475_), .ZN(new_n478_) );
  XNOR2_X1 g120 ( .A(new_n478_), .B(KEYINPUT5), .ZN(new_n479_) );
  AND2_X1 g121 ( .A1(new_n474_), .A2(new_n479_), .ZN(new_n480_) );
  XOR2_X1 g122 ( .A(new_n480_), .B(KEYINPUT7), .Z(G168) );
  AND2_X1 g123 ( .A1(new_n457_), .A2(G77), .ZN(new_n482_) );
  AND2_X1 g124 ( .A1(new_n454_), .A2(G90), .ZN(new_n483_) );
  OR2_X1 g125 ( .A1(new_n482_), .A2(new_n483_), .ZN(new_n484_) );
  INV_X1 g126 ( .A(new_n484_), .ZN(new_n485_) );
  AND2_X1 g127 ( .A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n486_) );
  INV_X1 g128 ( .A(new_n486_), .ZN(new_n487_) );
  OR2_X1 g129 ( .A1(new_n485_), .A2(KEYINPUT9), .ZN(new_n488_) );
  AND2_X1 g130 ( .A1(new_n466_), .A2(G52), .ZN(new_n489_) );
  AND2_X1 g131 ( .A1(new_n463_), .A2(G64), .ZN(new_n490_) );
  OR2_X1 g132 ( .A1(new_n490_), .A2(new_n489_), .ZN(new_n491_) );
  INV_X1 g133 ( .A(new_n491_), .ZN(new_n492_) );
  AND2_X1 g134 ( .A1(new_n488_), .A2(new_n492_), .ZN(new_n493_) );
  AND2_X1 g135 ( .A1(new_n493_), .A2(new_n487_), .ZN(G171) );
  INV_X1 g136 ( .A(G860), .ZN(new_n495_) );
  AND2_X1 g137 ( .A1(new_n457_), .A2(G68), .ZN(new_n496_) );
  AND2_X1 g138 ( .A1(new_n454_), .A2(G81), .ZN(new_n497_) );
  XNOR2_X1 g139 ( .A(new_n497_), .B(KEYINPUT12), .ZN(new_n498_) );
  OR2_X1 g140 ( .A1(new_n498_), .A2(new_n496_), .ZN(new_n499_) );
  XNOR2_X1 g141 ( .A(new_n499_), .B(KEYINPUT13), .ZN(new_n500_) );
  INV_X1 g142 ( .A(KEYINPUT14), .ZN(new_n501_) );
  INV_X1 g143 ( .A(G56), .ZN(new_n502_) );
  OR2_X1 g144 ( .A1(new_n462_), .A2(new_n502_), .ZN(new_n503_) );
  AND2_X1 g145 ( .A1(new_n503_), .A2(new_n501_), .ZN(new_n504_) );
  INV_X1 g146 ( .A(new_n504_), .ZN(new_n505_) );
  OR2_X1 g147 ( .A1(new_n503_), .A2(new_n501_), .ZN(new_n506_) );
  AND2_X1 g148 ( .A1(new_n466_), .A2(G43), .ZN(new_n507_) );
  INV_X1 g149 ( .A(new_n507_), .ZN(new_n508_) );
  AND2_X1 g150 ( .A1(new_n506_), .A2(new_n508_), .ZN(new_n509_) );
  AND2_X1 g151 ( .A1(new_n509_), .A2(new_n505_), .ZN(new_n510_) );
  AND2_X1 g152 ( .A1(new_n510_), .A2(new_n500_), .ZN(new_n511_) );
  INV_X1 g153 ( .A(new_n511_), .ZN(new_n512_) );
  OR2_X1 g154 ( .A1(new_n512_), .A2(new_n495_), .ZN(G153) );
  INV_X1 g155 ( .A(G36), .ZN(new_n514_) );
  INV_X1 g156 ( .A(G319), .ZN(new_n515_) );
  AND2_X1 g157 ( .A1(G483), .A2(G661), .ZN(new_n516_) );
  INV_X1 g158 ( .A(new_n516_), .ZN(new_n517_) );
  OR2_X1 g159 ( .A1(new_n515_), .A2(new_n517_), .ZN(new_n518_) );
  OR2_X1 g160 ( .A1(new_n518_), .A2(new_n514_), .ZN(G176) );
  AND2_X1 g161 ( .A1(G1), .A2(G3), .ZN(new_n520_) );
  OR2_X1 g162 ( .A1(new_n518_), .A2(new_n520_), .ZN(G188) );
  AND2_X1 g163 ( .A1(new_n454_), .A2(G91), .ZN(new_n522_) );
  AND2_X1 g164 ( .A1(new_n457_), .A2(G78), .ZN(new_n523_) );
  OR2_X1 g165 ( .A1(new_n523_), .A2(new_n522_), .ZN(new_n524_) );
  AND2_X1 g166 ( .A1(new_n463_), .A2(G65), .ZN(new_n525_) );
  AND2_X1 g167 ( .A1(new_n466_), .A2(G53), .ZN(new_n526_) );
  OR2_X1 g168 ( .A1(new_n525_), .A2(new_n526_), .ZN(new_n527_) );
  OR2_X1 g169 ( .A1(new_n527_), .A2(new_n524_), .ZN(G299) );
  INV_X1 g170 ( .A(G171), .ZN(G301) );
  XOR2_X1 g171 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 g172 ( .A1(new_n466_), .A2(G49), .ZN(new_n531_) );
  INV_X1 g173 ( .A(new_n456_), .ZN(new_n532_) );
  AND2_X1 g174 ( .A1(new_n532_), .A2(G87), .ZN(new_n533_) );
  AND2_X1 g175 ( .A1(G74), .A2(G651), .ZN(new_n534_) );
  OR2_X1 g176 ( .A1(new_n463_), .A2(new_n534_), .ZN(new_n535_) );
  OR2_X1 g177 ( .A1(new_n535_), .A2(new_n533_), .ZN(new_n536_) );
  OR2_X1 g178 ( .A1(new_n536_), .A2(new_n531_), .ZN(G288) );
  AND2_X1 g179 ( .A1(new_n463_), .A2(G61), .ZN(new_n538_) );
  AND2_X1 g180 ( .A1(new_n454_), .A2(G86), .ZN(new_n539_) );
  AND2_X1 g181 ( .A1(new_n466_), .A2(G48), .ZN(new_n540_) );
  OR2_X1 g182 ( .A1(new_n540_), .A2(new_n539_), .ZN(new_n541_) );
  OR2_X1 g183 ( .A1(new_n541_), .A2(new_n538_), .ZN(new_n542_) );
  INV_X1 g184 ( .A(new_n542_), .ZN(new_n543_) );
  AND2_X1 g185 ( .A1(new_n457_), .A2(G73), .ZN(new_n544_) );
  XOR2_X1 g186 ( .A(new_n544_), .B(KEYINPUT2), .Z(new_n545_) );
  AND2_X1 g187 ( .A1(new_n543_), .A2(new_n545_), .ZN(new_n546_) );
  INV_X1 g188 ( .A(new_n546_), .ZN(G305) );
  AND2_X1 g189 ( .A1(new_n454_), .A2(G85), .ZN(new_n548_) );
  AND2_X1 g190 ( .A1(new_n457_), .A2(G72), .ZN(new_n549_) );
  OR2_X1 g191 ( .A1(new_n549_), .A2(new_n548_), .ZN(new_n550_) );
  AND2_X1 g192 ( .A1(new_n463_), .A2(G60), .ZN(new_n551_) );
  AND2_X1 g193 ( .A1(new_n466_), .A2(G47), .ZN(new_n552_) );
  OR2_X1 g194 ( .A1(new_n551_), .A2(new_n552_), .ZN(new_n553_) );
  OR2_X1 g195 ( .A1(new_n553_), .A2(new_n550_), .ZN(G290) );
  AND2_X1 g196 ( .A1(G301), .A2(G868), .ZN(new_n555_) );
  INV_X1 g197 ( .A(G868), .ZN(new_n556_) );
  INV_X1 g198 ( .A(G92), .ZN(new_n557_) );
  OR2_X1 g199 ( .A1(new_n453_), .A2(new_n557_), .ZN(new_n558_) );
  AND2_X1 g200 ( .A1(new_n466_), .A2(G54), .ZN(new_n559_) );
  INV_X1 g201 ( .A(new_n559_), .ZN(new_n560_) );
  AND2_X1 g202 ( .A1(new_n560_), .A2(new_n558_), .ZN(new_n561_) );
  INV_X1 g203 ( .A(G66), .ZN(new_n562_) );
  OR2_X1 g204 ( .A1(new_n462_), .A2(new_n562_), .ZN(new_n563_) );
  AND2_X1 g205 ( .A1(new_n457_), .A2(G79), .ZN(new_n564_) );
  INV_X1 g206 ( .A(new_n564_), .ZN(new_n565_) );
  AND2_X1 g207 ( .A1(new_n565_), .A2(new_n563_), .ZN(new_n566_) );
  AND2_X1 g208 ( .A1(new_n566_), .A2(new_n561_), .ZN(new_n567_) );
  XNOR2_X1 g209 ( .A(new_n567_), .B(KEYINPUT15), .ZN(new_n568_) );
  AND2_X1 g210 ( .A1(new_n568_), .A2(new_n556_), .ZN(new_n569_) );
  OR2_X1 g211 ( .A1(new_n555_), .A2(new_n569_), .ZN(G284) );
  OR2_X1 g212 ( .A1(G286), .A2(new_n556_), .ZN(new_n571_) );
  OR2_X1 g213 ( .A1(G299), .A2(G868), .ZN(new_n572_) );
  AND2_X1 g214 ( .A1(new_n571_), .A2(new_n572_), .ZN(G297) );
  AND2_X1 g215 ( .A1(new_n495_), .A2(G559), .ZN(new_n574_) );
  OR2_X1 g216 ( .A1(new_n568_), .A2(new_n574_), .ZN(new_n575_) );
  XNOR2_X1 g217 ( .A(new_n575_), .B(KEYINPUT16), .ZN(G148) );
  OR2_X1 g218 ( .A1(new_n556_), .A2(G559), .ZN(new_n577_) );
  OR2_X1 g219 ( .A1(new_n568_), .A2(new_n577_), .ZN(new_n578_) );
  OR2_X1 g220 ( .A1(new_n512_), .A2(G868), .ZN(new_n579_) );
  AND2_X1 g221 ( .A1(new_n579_), .A2(new_n578_), .ZN(G282) );
  INV_X1 g222 ( .A(G2096), .ZN(new_n581_) );
  AND2_X1 g223 ( .A1(new_n412_), .A2(G135), .ZN(new_n582_) );
  INV_X1 g224 ( .A(new_n582_), .ZN(new_n583_) );
  AND2_X1 g225 ( .A1(new_n427_), .A2(G123), .ZN(new_n584_) );
  AND2_X1 g226 ( .A1(new_n584_), .A2(KEYINPUT18), .ZN(new_n585_) );
  INV_X1 g227 ( .A(new_n585_), .ZN(new_n586_) );
  OR2_X1 g228 ( .A1(new_n584_), .A2(KEYINPUT18), .ZN(new_n587_) );
  AND2_X1 g229 ( .A1(new_n437_), .A2(G99), .ZN(new_n588_) );
  AND2_X1 g230 ( .A1(new_n433_), .A2(G111), .ZN(new_n589_) );
  OR2_X1 g231 ( .A1(new_n588_), .A2(new_n589_), .ZN(new_n590_) );
  INV_X1 g232 ( .A(new_n590_), .ZN(new_n591_) );
  AND2_X1 g233 ( .A1(new_n591_), .A2(new_n587_), .ZN(new_n592_) );
  AND2_X1 g234 ( .A1(new_n592_), .A2(new_n586_), .ZN(new_n593_) );
  AND2_X1 g235 ( .A1(new_n593_), .A2(new_n583_), .ZN(new_n594_) );
  AND2_X1 g236 ( .A1(new_n594_), .A2(new_n581_), .ZN(new_n595_) );
  INV_X1 g237 ( .A(new_n594_), .ZN(new_n596_) );
  AND2_X1 g238 ( .A1(new_n596_), .A2(G2096), .ZN(new_n597_) );
  OR2_X1 g239 ( .A1(new_n597_), .A2(G2100), .ZN(new_n598_) );
  OR2_X1 g240 ( .A1(new_n598_), .A2(new_n595_), .ZN(G156) );
  XNOR2_X1 g241 ( .A(G1341), .B(G1348), .ZN(new_n600_) );
  XNOR2_X1 g242 ( .A(G2430), .B(G2454), .ZN(new_n601_) );
  XNOR2_X1 g243 ( .A(new_n600_), .B(new_n601_), .ZN(new_n602_) );
  XOR2_X1 g244 ( .A(G2435), .B(G2438), .Z(new_n603_) );
  XNOR2_X1 g245 ( .A(new_n602_), .B(new_n603_), .ZN(new_n604_) );
  INV_X1 g246 ( .A(new_n604_), .ZN(new_n605_) );
  XNOR2_X1 g247 ( .A(G2446), .B(G2451), .ZN(new_n606_) );
  XNOR2_X1 g248 ( .A(G2427), .B(G2443), .ZN(new_n607_) );
  XNOR2_X1 g249 ( .A(new_n606_), .B(new_n607_), .ZN(new_n608_) );
  INV_X1 g250 ( .A(new_n608_), .ZN(new_n609_) );
  AND2_X1 g251 ( .A1(new_n605_), .A2(new_n609_), .ZN(new_n610_) );
  INV_X1 g252 ( .A(new_n610_), .ZN(new_n611_) );
  AND2_X1 g253 ( .A1(new_n604_), .A2(new_n608_), .ZN(new_n612_) );
  INV_X1 g254 ( .A(new_n612_), .ZN(new_n613_) );
  AND2_X1 g255 ( .A1(new_n613_), .A2(G14), .ZN(new_n614_) );
  AND2_X1 g256 ( .A1(new_n614_), .A2(new_n611_), .ZN(G401) );
  XNOR2_X1 g257 ( .A(G2096), .B(G2100), .ZN(new_n616_) );
  XNOR2_X1 g258 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n617_) );
  XNOR2_X1 g259 ( .A(new_n616_), .B(new_n617_), .ZN(new_n618_) );
  XNOR2_X1 g260 ( .A(G2067), .B(G2072), .ZN(new_n619_) );
  XNOR2_X1 g261 ( .A(G2090), .B(KEYINPUT42), .ZN(new_n620_) );
  XNOR2_X1 g262 ( .A(new_n619_), .B(new_n620_), .ZN(new_n621_) );
  XNOR2_X1 g263 ( .A(new_n618_), .B(new_n621_), .ZN(new_n622_) );
  XOR2_X1 g264 ( .A(G2078), .B(G2084), .Z(new_n623_) );
  XOR2_X1 g265 ( .A(new_n622_), .B(new_n623_), .Z(new_n624_) );
  INV_X1 g266 ( .A(new_n624_), .ZN(G227) );
  XNOR2_X1 g267 ( .A(G1956), .B(G1966), .ZN(new_n626_) );
  XNOR2_X1 g268 ( .A(G1976), .B(G1981), .ZN(new_n627_) );
  XOR2_X1 g269 ( .A(new_n626_), .B(new_n627_), .Z(new_n628_) );
  XNOR2_X1 g270 ( .A(new_n628_), .B(G2474), .ZN(new_n629_) );
  XNOR2_X1 g271 ( .A(G1991), .B(G1996), .ZN(new_n630_) );
  XNOR2_X1 g272 ( .A(new_n629_), .B(new_n630_), .ZN(new_n631_) );
  XNOR2_X1 g273 ( .A(G1971), .B(KEYINPUT41), .ZN(new_n632_) );
  XNOR2_X1 g274 ( .A(G1961), .B(G1986), .ZN(new_n633_) );
  XNOR2_X1 g275 ( .A(new_n632_), .B(new_n633_), .ZN(new_n634_) );
  XOR2_X1 g276 ( .A(new_n631_), .B(new_n634_), .Z(new_n635_) );
  INV_X1 g277 ( .A(new_n635_), .ZN(G229) );
  INV_X1 g278 ( .A(G29), .ZN(new_n637_) );
  INV_X1 g279 ( .A(KEYINPUT55), .ZN(new_n638_) );
  INV_X1 g280 ( .A(G2090), .ZN(new_n639_) );
  XNOR2_X1 g281 ( .A(G162), .B(new_n639_), .ZN(new_n640_) );
  INV_X1 g282 ( .A(G1996), .ZN(new_n641_) );
  AND2_X1 g283 ( .A1(new_n412_), .A2(G141), .ZN(new_n642_) );
  INV_X1 g284 ( .A(new_n642_), .ZN(new_n643_) );
  AND2_X1 g285 ( .A1(new_n437_), .A2(G105), .ZN(new_n644_) );
  AND2_X1 g286 ( .A1(new_n644_), .A2(KEYINPUT38), .ZN(new_n645_) );
  INV_X1 g287 ( .A(new_n645_), .ZN(new_n646_) );
  OR2_X1 g288 ( .A1(new_n644_), .A2(KEYINPUT38), .ZN(new_n647_) );
  AND2_X1 g289 ( .A1(new_n433_), .A2(G117), .ZN(new_n648_) );
  AND2_X1 g290 ( .A1(new_n427_), .A2(G129), .ZN(new_n649_) );
  OR2_X1 g291 ( .A1(new_n649_), .A2(new_n648_), .ZN(new_n650_) );
  INV_X1 g292 ( .A(new_n650_), .ZN(new_n651_) );
  AND2_X1 g293 ( .A1(new_n651_), .A2(new_n647_), .ZN(new_n652_) );
  AND2_X1 g294 ( .A1(new_n652_), .A2(new_n646_), .ZN(new_n653_) );
  AND2_X1 g295 ( .A1(new_n653_), .A2(new_n643_), .ZN(new_n654_) );
  AND2_X1 g296 ( .A1(new_n654_), .A2(new_n641_), .ZN(new_n655_) );
  OR2_X1 g297 ( .A1(new_n640_), .A2(new_n655_), .ZN(new_n656_) );
  INV_X1 g298 ( .A(new_n656_), .ZN(new_n657_) );
  OR2_X1 g299 ( .A1(new_n657_), .A2(KEYINPUT51), .ZN(new_n658_) );
  INV_X1 g300 ( .A(KEYINPUT50), .ZN(new_n659_) );
  XNOR2_X1 g301 ( .A(new_n451_), .B(G2078), .ZN(new_n660_) );
  INV_X1 g302 ( .A(new_n660_), .ZN(new_n661_) );
  AND2_X1 g303 ( .A1(new_n427_), .A2(G127), .ZN(new_n662_) );
  AND2_X1 g304 ( .A1(new_n433_), .A2(G115), .ZN(new_n663_) );
  OR2_X1 g305 ( .A1(new_n662_), .A2(new_n663_), .ZN(new_n664_) );
  INV_X1 g306 ( .A(new_n664_), .ZN(new_n665_) );
  OR2_X1 g307 ( .A1(new_n665_), .A2(KEYINPUT47), .ZN(new_n666_) );
  INV_X1 g308 ( .A(G103), .ZN(new_n667_) );
  OR2_X1 g309 ( .A1(new_n438_), .A2(new_n667_), .ZN(new_n668_) );
  AND2_X1 g310 ( .A1(new_n666_), .A2(new_n668_), .ZN(new_n669_) );
  INV_X1 g311 ( .A(KEYINPUT47), .ZN(new_n670_) );
  OR2_X1 g312 ( .A1(new_n664_), .A2(new_n670_), .ZN(new_n671_) );
  INV_X1 g313 ( .A(G139), .ZN(new_n672_) );
  OR2_X1 g314 ( .A1(new_n413_), .A2(new_n672_), .ZN(new_n673_) );
  AND2_X1 g315 ( .A1(new_n671_), .A2(new_n673_), .ZN(new_n674_) );
  AND2_X1 g316 ( .A1(new_n669_), .A2(new_n674_), .ZN(new_n675_) );
  XNOR2_X1 g317 ( .A(new_n675_), .B(G2072), .ZN(new_n676_) );
  AND2_X1 g318 ( .A1(new_n676_), .A2(new_n661_), .ZN(new_n677_) );
  OR2_X1 g319 ( .A1(new_n677_), .A2(new_n659_), .ZN(new_n678_) );
  INV_X1 g320 ( .A(KEYINPUT51), .ZN(new_n679_) );
  OR2_X1 g321 ( .A1(new_n656_), .A2(new_n679_), .ZN(new_n680_) );
  AND2_X1 g322 ( .A1(new_n680_), .A2(new_n678_), .ZN(new_n681_) );
  AND2_X1 g323 ( .A1(new_n681_), .A2(new_n658_), .ZN(new_n682_) );
  AND2_X1 g324 ( .A1(new_n412_), .A2(G140), .ZN(new_n683_) );
  AND2_X1 g325 ( .A1(new_n437_), .A2(G104), .ZN(new_n684_) );
  OR2_X1 g326 ( .A1(new_n683_), .A2(new_n684_), .ZN(new_n685_) );
  OR2_X1 g327 ( .A1(new_n685_), .A2(KEYINPUT34), .ZN(new_n686_) );
  INV_X1 g328 ( .A(KEYINPUT34), .ZN(new_n687_) );
  INV_X1 g329 ( .A(new_n685_), .ZN(new_n688_) );
  OR2_X1 g330 ( .A1(new_n688_), .A2(new_n687_), .ZN(new_n689_) );
  AND2_X1 g331 ( .A1(new_n427_), .A2(G128), .ZN(new_n690_) );
  AND2_X1 g332 ( .A1(new_n433_), .A2(G116), .ZN(new_n691_) );
  OR2_X1 g333 ( .A1(new_n690_), .A2(new_n691_), .ZN(new_n692_) );
  XNOR2_X1 g334 ( .A(new_n692_), .B(KEYINPUT35), .ZN(new_n693_) );
  AND2_X1 g335 ( .A1(new_n689_), .A2(new_n693_), .ZN(new_n694_) );
  AND2_X1 g336 ( .A1(new_n694_), .A2(new_n686_), .ZN(new_n695_) );
  XOR2_X1 g337 ( .A(new_n695_), .B(KEYINPUT36), .Z(new_n696_) );
  INV_X1 g338 ( .A(new_n696_), .ZN(new_n697_) );
  XOR2_X1 g339 ( .A(G2067), .B(KEYINPUT37), .Z(new_n698_) );
  INV_X1 g340 ( .A(new_n698_), .ZN(new_n699_) );
  AND2_X1 g341 ( .A1(new_n697_), .A2(new_n699_), .ZN(new_n700_) );
  INV_X1 g342 ( .A(new_n700_), .ZN(new_n701_) );
  OR2_X1 g343 ( .A1(new_n697_), .A2(new_n699_), .ZN(new_n702_) );
  INV_X1 g344 ( .A(new_n677_), .ZN(new_n703_) );
  OR2_X1 g345 ( .A1(new_n703_), .A2(KEYINPUT50), .ZN(new_n704_) );
  INV_X1 g346 ( .A(new_n654_), .ZN(new_n705_) );
  AND2_X1 g347 ( .A1(new_n705_), .A2(G1996), .ZN(new_n706_) );
  AND2_X1 g348 ( .A1(new_n412_), .A2(G131), .ZN(new_n707_) );
  AND2_X1 g349 ( .A1(new_n437_), .A2(G95), .ZN(new_n708_) );
  AND2_X1 g350 ( .A1(new_n433_), .A2(G107), .ZN(new_n709_) );
  AND2_X1 g351 ( .A1(new_n427_), .A2(G119), .ZN(new_n710_) );
  OR2_X1 g352 ( .A1(new_n710_), .A2(new_n709_), .ZN(new_n711_) );
  OR2_X1 g353 ( .A1(new_n711_), .A2(new_n708_), .ZN(new_n712_) );
  OR2_X1 g354 ( .A1(new_n712_), .A2(new_n707_), .ZN(new_n713_) );
  AND2_X1 g355 ( .A1(new_n713_), .A2(G1991), .ZN(new_n714_) );
  OR2_X1 g356 ( .A1(new_n706_), .A2(new_n714_), .ZN(new_n715_) );
  INV_X1 g357 ( .A(new_n715_), .ZN(new_n716_) );
  XNOR2_X1 g358 ( .A(G160), .B(G2084), .ZN(new_n717_) );
  OR2_X1 g359 ( .A1(new_n713_), .A2(G1991), .ZN(new_n718_) );
  AND2_X1 g360 ( .A1(new_n596_), .A2(new_n718_), .ZN(new_n719_) );
  AND2_X1 g361 ( .A1(new_n719_), .A2(new_n717_), .ZN(new_n720_) );
  AND2_X1 g362 ( .A1(new_n716_), .A2(new_n720_), .ZN(new_n721_) );
  AND2_X1 g363 ( .A1(new_n704_), .A2(new_n721_), .ZN(new_n722_) );
  AND2_X1 g364 ( .A1(new_n722_), .A2(new_n702_), .ZN(new_n723_) );
  AND2_X1 g365 ( .A1(new_n723_), .A2(new_n701_), .ZN(new_n724_) );
  AND2_X1 g366 ( .A1(new_n724_), .A2(new_n682_), .ZN(new_n725_) );
  XNOR2_X1 g367 ( .A(new_n725_), .B(KEYINPUT52), .ZN(new_n726_) );
  AND2_X1 g368 ( .A1(new_n726_), .A2(new_n638_), .ZN(new_n727_) );
  OR2_X1 g369 ( .A1(new_n727_), .A2(new_n637_), .ZN(new_n728_) );
  INV_X1 g370 ( .A(G168), .ZN(new_n729_) );
  OR2_X1 g371 ( .A1(new_n729_), .A2(G1966), .ZN(new_n730_) );
  XNOR2_X1 g372 ( .A(new_n546_), .B(G1981), .ZN(new_n731_) );
  INV_X1 g373 ( .A(G1966), .ZN(new_n732_) );
  OR2_X1 g374 ( .A1(G168), .A2(new_n732_), .ZN(new_n733_) );
  AND2_X1 g375 ( .A1(new_n733_), .A2(new_n731_), .ZN(new_n734_) );
  AND2_X1 g376 ( .A1(new_n734_), .A2(new_n730_), .ZN(new_n735_) );
  XOR2_X1 g377 ( .A(new_n735_), .B(KEYINPUT57), .Z(new_n736_) );
  XNOR2_X1 g378 ( .A(new_n511_), .B(G1341), .ZN(new_n737_) );
  INV_X1 g379 ( .A(G1956), .ZN(new_n738_) );
  XNOR2_X1 g380 ( .A(G299), .B(new_n738_), .ZN(new_n739_) );
  INV_X1 g381 ( .A(G1976), .ZN(new_n740_) );
  INV_X1 g382 ( .A(G288), .ZN(new_n741_) );
  OR2_X1 g383 ( .A1(new_n741_), .A2(new_n740_), .ZN(new_n742_) );
  INV_X1 g384 ( .A(G1971), .ZN(new_n743_) );
  OR2_X1 g385 ( .A1(G166), .A2(new_n743_), .ZN(new_n744_) );
  AND2_X1 g386 ( .A1(new_n742_), .A2(new_n744_), .ZN(new_n745_) );
  AND2_X1 g387 ( .A1(new_n745_), .A2(new_n739_), .ZN(new_n746_) );
  AND2_X1 g388 ( .A1(new_n741_), .A2(new_n740_), .ZN(new_n747_) );
  AND2_X1 g389 ( .A1(G166), .A2(new_n743_), .ZN(new_n748_) );
  OR2_X1 g390 ( .A1(new_n747_), .A2(new_n748_), .ZN(new_n749_) );
  INV_X1 g391 ( .A(new_n749_), .ZN(new_n750_) );
  XOR2_X1 g392 ( .A(G290), .B(G1986), .Z(new_n751_) );
  AND2_X1 g393 ( .A1(new_n750_), .A2(new_n751_), .ZN(new_n752_) );
  AND2_X1 g394 ( .A1(new_n752_), .A2(new_n746_), .ZN(new_n753_) );
  AND2_X1 g395 ( .A1(new_n753_), .A2(new_n737_), .ZN(new_n754_) );
  XNOR2_X1 g396 ( .A(G171), .B(G1961), .ZN(new_n755_) );
  INV_X1 g397 ( .A(G1348), .ZN(new_n756_) );
  XNOR2_X1 g398 ( .A(new_n568_), .B(new_n756_), .ZN(new_n757_) );
  AND2_X1 g399 ( .A1(new_n755_), .A2(new_n757_), .ZN(new_n758_) );
  AND2_X1 g400 ( .A1(new_n754_), .A2(new_n758_), .ZN(new_n759_) );
  AND2_X1 g401 ( .A1(new_n736_), .A2(new_n759_), .ZN(new_n760_) );
  XOR2_X1 g402 ( .A(G16), .B(KEYINPUT56), .Z(new_n761_) );
  OR2_X1 g403 ( .A1(new_n760_), .A2(new_n761_), .ZN(new_n762_) );
  INV_X1 g404 ( .A(KEYINPUT53), .ZN(new_n763_) );
  XOR2_X1 g405 ( .A(G25), .B(G1991), .Z(new_n764_) );
  OR2_X1 g406 ( .A1(G33), .A2(G2072), .ZN(new_n765_) );
  AND2_X1 g407 ( .A1(new_n765_), .A2(G28), .ZN(new_n766_) );
  XOR2_X1 g408 ( .A(G32), .B(G1996), .Z(new_n767_) );
  AND2_X1 g409 ( .A1(new_n766_), .A2(new_n767_), .ZN(new_n768_) );
  AND2_X1 g410 ( .A1(new_n768_), .A2(new_n764_), .ZN(new_n769_) );
  XOR2_X1 g411 ( .A(G2078), .B(KEYINPUT25), .Z(new_n770_) );
  AND2_X1 g412 ( .A1(new_n770_), .A2(G27), .ZN(new_n771_) );
  INV_X1 g413 ( .A(new_n771_), .ZN(new_n772_) );
  OR2_X1 g414 ( .A1(new_n770_), .A2(G27), .ZN(new_n773_) );
  AND2_X1 g415 ( .A1(G33), .A2(G2072), .ZN(new_n774_) );
  INV_X1 g416 ( .A(new_n774_), .ZN(new_n775_) );
  XOR2_X1 g417 ( .A(G26), .B(G2067), .Z(new_n776_) );
  AND2_X1 g418 ( .A1(new_n776_), .A2(new_n775_), .ZN(new_n777_) );
  AND2_X1 g419 ( .A1(new_n773_), .A2(new_n777_), .ZN(new_n778_) );
  AND2_X1 g420 ( .A1(new_n778_), .A2(new_n772_), .ZN(new_n779_) );
  AND2_X1 g421 ( .A1(new_n779_), .A2(new_n769_), .ZN(new_n780_) );
  INV_X1 g422 ( .A(new_n780_), .ZN(new_n781_) );
  AND2_X1 g423 ( .A1(new_n781_), .A2(new_n763_), .ZN(new_n782_) );
  AND2_X1 g424 ( .A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n783_) );
  XNOR2_X1 g425 ( .A(G35), .B(G2090), .ZN(new_n784_) );
  XNOR2_X1 g426 ( .A(G2084), .B(KEYINPUT54), .ZN(new_n785_) );
  XNOR2_X1 g427 ( .A(new_n785_), .B(G34), .ZN(new_n786_) );
  OR2_X1 g428 ( .A1(new_n786_), .A2(new_n784_), .ZN(new_n787_) );
  OR2_X1 g429 ( .A1(new_n783_), .A2(new_n787_), .ZN(new_n788_) );
  OR2_X1 g430 ( .A1(new_n788_), .A2(new_n782_), .ZN(new_n789_) );
  INV_X1 g431 ( .A(new_n789_), .ZN(new_n790_) );
  AND2_X1 g432 ( .A1(new_n790_), .A2(new_n638_), .ZN(new_n791_) );
  AND2_X1 g433 ( .A1(new_n789_), .A2(KEYINPUT55), .ZN(new_n792_) );
  OR2_X1 g434 ( .A1(new_n792_), .A2(G29), .ZN(new_n793_) );
  OR2_X1 g435 ( .A1(new_n793_), .A2(new_n791_), .ZN(new_n794_) );
  INV_X1 g436 ( .A(KEYINPUT61), .ZN(new_n795_) );
  INV_X1 g437 ( .A(KEYINPUT58), .ZN(new_n796_) );
  XNOR2_X1 g438 ( .A(G24), .B(G1986), .ZN(new_n797_) );
  INV_X1 g439 ( .A(new_n797_), .ZN(new_n798_) );
  OR2_X1 g440 ( .A1(G23), .A2(G1976), .ZN(new_n799_) );
  OR2_X1 g441 ( .A1(G22), .A2(G1971), .ZN(new_n800_) );
  AND2_X1 g442 ( .A1(new_n799_), .A2(new_n800_), .ZN(new_n801_) );
  AND2_X1 g443 ( .A1(G22), .A2(G1971), .ZN(new_n802_) );
  AND2_X1 g444 ( .A1(G23), .A2(G1976), .ZN(new_n803_) );
  OR2_X1 g445 ( .A1(new_n802_), .A2(new_n803_), .ZN(new_n804_) );
  INV_X1 g446 ( .A(new_n804_), .ZN(new_n805_) );
  AND2_X1 g447 ( .A1(new_n805_), .A2(new_n801_), .ZN(new_n806_) );
  AND2_X1 g448 ( .A1(new_n806_), .A2(new_n798_), .ZN(new_n807_) );
  OR2_X1 g449 ( .A1(new_n807_), .A2(new_n796_), .ZN(new_n808_) );
  AND2_X1 g450 ( .A1(new_n807_), .A2(new_n796_), .ZN(new_n809_) );
  INV_X1 g451 ( .A(new_n809_), .ZN(new_n810_) );
  OR2_X1 g452 ( .A1(G21), .A2(G1966), .ZN(new_n811_) );
  OR2_X1 g453 ( .A1(G5), .A2(G1961), .ZN(new_n812_) );
  AND2_X1 g454 ( .A1(new_n811_), .A2(new_n812_), .ZN(new_n813_) );
  AND2_X1 g455 ( .A1(G5), .A2(G1961), .ZN(new_n814_) );
  AND2_X1 g456 ( .A1(G21), .A2(G1966), .ZN(new_n815_) );
  OR2_X1 g457 ( .A1(new_n814_), .A2(new_n815_), .ZN(new_n816_) );
  INV_X1 g458 ( .A(new_n816_), .ZN(new_n817_) );
  AND2_X1 g459 ( .A1(new_n817_), .A2(new_n813_), .ZN(new_n818_) );
  AND2_X1 g460 ( .A1(new_n810_), .A2(new_n818_), .ZN(new_n819_) );
  AND2_X1 g461 ( .A1(new_n819_), .A2(new_n808_), .ZN(new_n820_) );
  XNOR2_X1 g462 ( .A(G1348), .B(KEYINPUT59), .ZN(new_n821_) );
  XNOR2_X1 g463 ( .A(new_n821_), .B(G4), .ZN(new_n822_) );
  XOR2_X1 g464 ( .A(G20), .B(G1956), .Z(new_n823_) );
  XOR2_X1 g465 ( .A(G6), .B(G1981), .Z(new_n824_) );
  XOR2_X1 g466 ( .A(G19), .B(G1341), .Z(new_n825_) );
  AND2_X1 g467 ( .A1(new_n824_), .A2(new_n825_), .ZN(new_n826_) );
  AND2_X1 g468 ( .A1(new_n826_), .A2(new_n823_), .ZN(new_n827_) );
  AND2_X1 g469 ( .A1(new_n827_), .A2(new_n822_), .ZN(new_n828_) );
  XNOR2_X1 g470 ( .A(new_n828_), .B(KEYINPUT60), .ZN(new_n829_) );
  AND2_X1 g471 ( .A1(new_n820_), .A2(new_n829_), .ZN(new_n830_) );
  AND2_X1 g472 ( .A1(new_n830_), .A2(new_n795_), .ZN(new_n831_) );
  INV_X1 g473 ( .A(new_n830_), .ZN(new_n832_) );
  AND2_X1 g474 ( .A1(new_n832_), .A2(KEYINPUT61), .ZN(new_n833_) );
  OR2_X1 g475 ( .A1(new_n833_), .A2(G16), .ZN(new_n834_) );
  OR2_X1 g476 ( .A1(new_n834_), .A2(new_n831_), .ZN(new_n835_) );
  AND2_X1 g477 ( .A1(new_n835_), .A2(G11), .ZN(new_n836_) );
  AND2_X1 g478 ( .A1(new_n836_), .A2(new_n794_), .ZN(new_n837_) );
  AND2_X1 g479 ( .A1(new_n762_), .A2(new_n837_), .ZN(new_n838_) );
  AND2_X1 g480 ( .A1(new_n728_), .A2(new_n838_), .ZN(new_n839_) );
  XOR2_X1 g481 ( .A(new_n839_), .B(KEYINPUT62), .Z(G150) );
  INV_X1 g482 ( .A(G150), .ZN(G311) );
  INV_X1 g483 ( .A(new_n568_), .ZN(new_n842_) );
  AND2_X1 g484 ( .A1(new_n842_), .A2(G559), .ZN(new_n843_) );
  INV_X1 g485 ( .A(new_n843_), .ZN(new_n844_) );
  AND2_X1 g486 ( .A1(new_n844_), .A2(new_n512_), .ZN(new_n845_) );
  AND2_X1 g487 ( .A1(new_n843_), .A2(new_n511_), .ZN(new_n846_) );
  OR2_X1 g488 ( .A1(new_n846_), .A2(G860), .ZN(new_n847_) );
  OR2_X1 g489 ( .A1(new_n847_), .A2(new_n845_), .ZN(new_n848_) );
  AND2_X1 g490 ( .A1(new_n454_), .A2(G93), .ZN(new_n849_) );
  AND2_X1 g491 ( .A1(new_n457_), .A2(G80), .ZN(new_n850_) );
  OR2_X1 g492 ( .A1(new_n850_), .A2(new_n849_), .ZN(new_n851_) );
  AND2_X1 g493 ( .A1(new_n463_), .A2(G67), .ZN(new_n852_) );
  AND2_X1 g494 ( .A1(new_n466_), .A2(G55), .ZN(new_n853_) );
  OR2_X1 g495 ( .A1(new_n852_), .A2(new_n853_), .ZN(new_n854_) );
  OR2_X1 g496 ( .A1(new_n854_), .A2(new_n851_), .ZN(new_n855_) );
  XNOR2_X1 g497 ( .A(new_n848_), .B(new_n855_), .ZN(G145) );
  INV_X1 g498 ( .A(KEYINPUT45), .ZN(new_n857_) );
  AND2_X1 g499 ( .A1(new_n412_), .A2(G142), .ZN(new_n858_) );
  AND2_X1 g500 ( .A1(new_n437_), .A2(G106), .ZN(new_n859_) );
  OR2_X1 g501 ( .A1(new_n858_), .A2(new_n859_), .ZN(new_n860_) );
  AND2_X1 g502 ( .A1(new_n860_), .A2(new_n857_), .ZN(new_n861_) );
  INV_X1 g503 ( .A(new_n860_), .ZN(new_n862_) );
  AND2_X1 g504 ( .A1(new_n862_), .A2(KEYINPUT45), .ZN(new_n863_) );
  AND2_X1 g505 ( .A1(new_n433_), .A2(G118), .ZN(new_n864_) );
  AND2_X1 g506 ( .A1(new_n427_), .A2(G130), .ZN(new_n865_) );
  OR2_X1 g507 ( .A1(new_n865_), .A2(new_n864_), .ZN(new_n866_) );
  OR2_X1 g508 ( .A1(new_n863_), .A2(new_n866_), .ZN(new_n867_) );
  OR2_X1 g509 ( .A1(new_n867_), .A2(new_n861_), .ZN(new_n868_) );
  XNOR2_X1 g510 ( .A(new_n868_), .B(new_n654_), .ZN(new_n869_) );
  XNOR2_X1 g511 ( .A(new_n869_), .B(G162), .ZN(new_n870_) );
  XNOR2_X1 g512 ( .A(new_n675_), .B(G160), .ZN(new_n871_) );
  XNOR2_X1 g513 ( .A(new_n696_), .B(new_n871_), .ZN(new_n872_) );
  XOR2_X1 g514 ( .A(new_n872_), .B(new_n870_), .Z(new_n873_) );
  INV_X1 g515 ( .A(new_n873_), .ZN(new_n874_) );
  XNOR2_X1 g516 ( .A(new_n594_), .B(new_n713_), .ZN(new_n875_) );
  XOR2_X1 g517 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(new_n876_) );
  XNOR2_X1 g518 ( .A(new_n875_), .B(new_n876_), .ZN(new_n877_) );
  XNOR2_X1 g519 ( .A(new_n877_), .B(new_n451_), .ZN(new_n878_) );
  INV_X1 g520 ( .A(new_n878_), .ZN(new_n879_) );
  AND2_X1 g521 ( .A1(new_n874_), .A2(new_n879_), .ZN(new_n880_) );
  AND2_X1 g522 ( .A1(new_n873_), .A2(new_n878_), .ZN(new_n881_) );
  OR2_X1 g523 ( .A1(new_n881_), .A2(G37), .ZN(new_n882_) );
  OR2_X1 g524 ( .A1(new_n882_), .A2(new_n880_), .ZN(new_n883_) );
  INV_X1 g525 ( .A(new_n883_), .ZN(G395) );
  XNOR2_X1 g526 ( .A(new_n511_), .B(G290), .ZN(new_n885_) );
  XNOR2_X1 g527 ( .A(new_n885_), .B(new_n741_), .ZN(new_n886_) );
  XNOR2_X1 g528 ( .A(G299), .B(KEYINPUT19), .ZN(new_n887_) );
  XNOR2_X1 g529 ( .A(new_n887_), .B(G305), .ZN(new_n888_) );
  XNOR2_X1 g530 ( .A(new_n886_), .B(new_n888_), .ZN(new_n889_) );
  XOR2_X1 g531 ( .A(G303), .B(new_n855_), .Z(new_n890_) );
  XNOR2_X1 g532 ( .A(new_n889_), .B(new_n890_), .ZN(new_n891_) );
  XNOR2_X1 g533 ( .A(new_n891_), .B(new_n844_), .ZN(new_n892_) );
  AND2_X1 g534 ( .A1(new_n892_), .A2(G868), .ZN(new_n893_) );
  AND2_X1 g535 ( .A1(new_n855_), .A2(new_n556_), .ZN(new_n894_) );
  OR2_X1 g536 ( .A1(new_n893_), .A2(new_n894_), .ZN(G295) );
  XNOR2_X1 g537 ( .A(G286), .B(new_n842_), .ZN(new_n896_) );
  XNOR2_X1 g538 ( .A(new_n891_), .B(new_n896_), .ZN(new_n897_) );
  AND2_X1 g539 ( .A1(new_n897_), .A2(G301), .ZN(new_n898_) );
  INV_X1 g540 ( .A(new_n898_), .ZN(new_n899_) );
  INV_X1 g541 ( .A(G37), .ZN(new_n900_) );
  OR2_X1 g542 ( .A1(new_n897_), .A2(G301), .ZN(new_n901_) );
  AND2_X1 g543 ( .A1(new_n901_), .A2(new_n900_), .ZN(new_n902_) );
  AND2_X1 g544 ( .A1(new_n902_), .A2(new_n899_), .ZN(G397) );
  INV_X1 g545 ( .A(KEYINPUT32), .ZN(new_n904_) );
  INV_X1 g546 ( .A(KEYINPUT26), .ZN(new_n905_) );
  AND2_X1 g547 ( .A1(new_n418_), .A2(G40), .ZN(new_n906_) );
  AND2_X1 g548 ( .A1(new_n906_), .A2(new_n421_), .ZN(new_n907_) );
  AND2_X1 g549 ( .A1(new_n415_), .A2(new_n907_), .ZN(new_n908_) );
  INV_X1 g550 ( .A(G1384), .ZN(new_n909_) );
  AND2_X1 g551 ( .A1(new_n451_), .A2(new_n909_), .ZN(new_n910_) );
  AND2_X1 g552 ( .A1(new_n910_), .A2(new_n908_), .ZN(new_n911_) );
  AND2_X1 g553 ( .A1(new_n911_), .A2(G1996), .ZN(new_n912_) );
  XNOR2_X1 g554 ( .A(new_n912_), .B(new_n905_), .ZN(new_n913_) );
  INV_X1 g555 ( .A(G1341), .ZN(new_n914_) );
  OR2_X1 g556 ( .A1(new_n911_), .A2(new_n914_), .ZN(new_n915_) );
  AND2_X1 g557 ( .A1(new_n915_), .A2(new_n511_), .ZN(new_n916_) );
  AND2_X1 g558 ( .A1(new_n913_), .A2(new_n916_), .ZN(new_n917_) );
  AND2_X1 g559 ( .A1(new_n917_), .A2(new_n842_), .ZN(new_n918_) );
  INV_X1 g560 ( .A(G2067), .ZN(new_n919_) );
  INV_X1 g561 ( .A(new_n911_), .ZN(new_n920_) );
  OR2_X1 g562 ( .A1(new_n920_), .A2(new_n919_), .ZN(new_n921_) );
  OR2_X1 g563 ( .A1(new_n911_), .A2(new_n756_), .ZN(new_n922_) );
  AND2_X1 g564 ( .A1(new_n921_), .A2(new_n922_), .ZN(new_n923_) );
  OR2_X1 g565 ( .A1(new_n918_), .A2(new_n923_), .ZN(new_n924_) );
  OR2_X1 g566 ( .A1(new_n917_), .A2(new_n842_), .ZN(new_n925_) );
  AND2_X1 g567 ( .A1(new_n924_), .A2(new_n925_), .ZN(new_n926_) );
  INV_X1 g568 ( .A(G299), .ZN(new_n927_) );
  AND2_X1 g569 ( .A1(new_n911_), .A2(G2072), .ZN(new_n928_) );
  INV_X1 g570 ( .A(new_n928_), .ZN(new_n929_) );
  OR2_X1 g571 ( .A1(new_n929_), .A2(KEYINPUT27), .ZN(new_n930_) );
  OR2_X1 g572 ( .A1(new_n911_), .A2(new_n738_), .ZN(new_n931_) );
  INV_X1 g573 ( .A(KEYINPUT27), .ZN(new_n932_) );
  OR2_X1 g574 ( .A1(new_n928_), .A2(new_n932_), .ZN(new_n933_) );
  AND2_X1 g575 ( .A1(new_n933_), .A2(new_n931_), .ZN(new_n934_) );
  AND2_X1 g576 ( .A1(new_n934_), .A2(new_n930_), .ZN(new_n935_) );
  AND2_X1 g577 ( .A1(new_n935_), .A2(new_n927_), .ZN(new_n936_) );
  OR2_X1 g578 ( .A1(new_n926_), .A2(new_n936_), .ZN(new_n937_) );
  OR2_X1 g579 ( .A1(new_n935_), .A2(new_n927_), .ZN(new_n938_) );
  XNOR2_X1 g580 ( .A(new_n938_), .B(KEYINPUT28), .ZN(new_n939_) );
  AND2_X1 g581 ( .A1(new_n937_), .A2(new_n939_), .ZN(new_n940_) );
  XNOR2_X1 g582 ( .A(new_n940_), .B(KEYINPUT29), .ZN(new_n941_) );
  OR2_X1 g583 ( .A1(new_n920_), .A2(new_n770_), .ZN(new_n942_) );
  OR2_X1 g584 ( .A1(new_n911_), .A2(G1961), .ZN(new_n943_) );
  AND2_X1 g585 ( .A1(new_n942_), .A2(new_n943_), .ZN(new_n944_) );
  OR2_X1 g586 ( .A1(new_n944_), .A2(G301), .ZN(new_n945_) );
  AND2_X1 g587 ( .A1(new_n941_), .A2(new_n945_), .ZN(new_n946_) );
  AND2_X1 g588 ( .A1(new_n920_), .A2(G8), .ZN(new_n947_) );
  AND2_X1 g589 ( .A1(new_n947_), .A2(new_n732_), .ZN(new_n948_) );
  INV_X1 g590 ( .A(new_n948_), .ZN(new_n949_) );
  OR2_X1 g591 ( .A1(new_n920_), .A2(G2084), .ZN(new_n950_) );
  AND2_X1 g592 ( .A1(new_n950_), .A2(G8), .ZN(new_n951_) );
  AND2_X1 g593 ( .A1(new_n949_), .A2(new_n951_), .ZN(new_n952_) );
  INV_X1 g594 ( .A(new_n952_), .ZN(new_n953_) );
  OR2_X1 g595 ( .A1(new_n953_), .A2(KEYINPUT30), .ZN(new_n954_) );
  INV_X1 g596 ( .A(KEYINPUT30), .ZN(new_n955_) );
  OR2_X1 g597 ( .A1(new_n952_), .A2(new_n955_), .ZN(new_n956_) );
  AND2_X1 g598 ( .A1(new_n956_), .A2(new_n729_), .ZN(new_n957_) );
  AND2_X1 g599 ( .A1(new_n957_), .A2(new_n954_), .ZN(new_n958_) );
  AND2_X1 g600 ( .A1(new_n944_), .A2(G301), .ZN(new_n959_) );
  OR2_X1 g601 ( .A1(new_n958_), .A2(new_n959_), .ZN(new_n960_) );
  XOR2_X1 g602 ( .A(new_n960_), .B(KEYINPUT31), .Z(new_n961_) );
  OR2_X1 g603 ( .A1(new_n946_), .A2(new_n961_), .ZN(new_n962_) );
  AND2_X1 g604 ( .A1(new_n962_), .A2(G286), .ZN(new_n963_) );
  AND2_X1 g605 ( .A1(new_n947_), .A2(new_n743_), .ZN(new_n964_) );
  AND2_X1 g606 ( .A1(new_n911_), .A2(new_n639_), .ZN(new_n965_) );
  OR2_X1 g607 ( .A1(new_n965_), .A2(G166), .ZN(new_n966_) );
  OR2_X1 g608 ( .A1(new_n964_), .A2(new_n966_), .ZN(new_n967_) );
  INV_X1 g609 ( .A(new_n967_), .ZN(new_n968_) );
  OR2_X1 g610 ( .A1(new_n963_), .A2(new_n968_), .ZN(new_n969_) );
  AND2_X1 g611 ( .A1(new_n969_), .A2(G8), .ZN(new_n970_) );
  INV_X1 g612 ( .A(new_n970_), .ZN(new_n971_) );
  OR2_X1 g613 ( .A1(new_n971_), .A2(new_n904_), .ZN(new_n972_) );
  INV_X1 g614 ( .A(new_n962_), .ZN(new_n973_) );
  INV_X1 g615 ( .A(new_n950_), .ZN(new_n974_) );
  AND2_X1 g616 ( .A1(new_n974_), .A2(G8), .ZN(new_n975_) );
  OR2_X1 g617 ( .A1(new_n975_), .A2(new_n948_), .ZN(new_n976_) );
  OR2_X1 g618 ( .A1(new_n973_), .A2(new_n976_), .ZN(new_n977_) );
  OR2_X1 g619 ( .A1(new_n970_), .A2(KEYINPUT32), .ZN(new_n978_) );
  AND2_X1 g620 ( .A1(new_n978_), .A2(new_n977_), .ZN(new_n979_) );
  AND2_X1 g621 ( .A1(new_n979_), .A2(new_n972_), .ZN(new_n980_) );
  OR2_X1 g622 ( .A1(new_n980_), .A2(new_n749_), .ZN(new_n981_) );
  AND2_X1 g623 ( .A1(new_n947_), .A2(new_n742_), .ZN(new_n982_) );
  AND2_X1 g624 ( .A1(new_n981_), .A2(new_n982_), .ZN(new_n983_) );
  OR2_X1 g625 ( .A1(new_n983_), .A2(KEYINPUT33), .ZN(new_n984_) );
  INV_X1 g626 ( .A(new_n947_), .ZN(new_n985_) );
  AND2_X1 g627 ( .A1(new_n747_), .A2(KEYINPUT33), .ZN(new_n986_) );
  INV_X1 g628 ( .A(new_n986_), .ZN(new_n987_) );
  OR2_X1 g629 ( .A1(new_n987_), .A2(new_n985_), .ZN(new_n988_) );
  AND2_X1 g630 ( .A1(new_n988_), .A2(new_n731_), .ZN(new_n989_) );
  AND2_X1 g631 ( .A1(new_n984_), .A2(new_n989_), .ZN(new_n990_) );
  AND2_X1 g632 ( .A1(new_n639_), .A2(G8), .ZN(new_n991_) );
  AND2_X1 g633 ( .A1(G166), .A2(new_n991_), .ZN(new_n992_) );
  OR2_X1 g634 ( .A1(new_n980_), .A2(new_n992_), .ZN(new_n993_) );
  AND2_X1 g635 ( .A1(new_n993_), .A2(new_n985_), .ZN(new_n994_) );
  INV_X1 g636 ( .A(G1981), .ZN(new_n995_) );
  AND2_X1 g637 ( .A1(new_n546_), .A2(new_n995_), .ZN(new_n996_) );
  INV_X1 g638 ( .A(new_n996_), .ZN(new_n997_) );
  OR2_X1 g639 ( .A1(new_n997_), .A2(KEYINPUT24), .ZN(new_n998_) );
  INV_X1 g640 ( .A(KEYINPUT24), .ZN(new_n999_) );
  OR2_X1 g641 ( .A1(new_n996_), .A2(new_n999_), .ZN(new_n1000_) );
  AND2_X1 g642 ( .A1(new_n1000_), .A2(new_n947_), .ZN(new_n1001_) );
  AND2_X1 g643 ( .A1(new_n1001_), .A2(new_n998_), .ZN(new_n1002_) );
  OR2_X1 g644 ( .A1(new_n994_), .A2(new_n1002_), .ZN(new_n1003_) );
  OR2_X1 g645 ( .A1(new_n990_), .A2(new_n1003_), .ZN(new_n1004_) );
  INV_X1 g646 ( .A(new_n910_), .ZN(new_n1005_) );
  AND2_X1 g647 ( .A1(new_n1005_), .A2(new_n908_), .ZN(new_n1006_) );
  INV_X1 g648 ( .A(new_n1006_), .ZN(new_n1007_) );
  OR2_X1 g649 ( .A1(new_n702_), .A2(new_n1007_), .ZN(new_n1008_) );
  AND2_X1 g650 ( .A1(new_n715_), .A2(new_n1006_), .ZN(new_n1009_) );
  INV_X1 g651 ( .A(new_n1009_), .ZN(new_n1010_) );
  OR2_X1 g652 ( .A1(new_n751_), .A2(new_n1007_), .ZN(new_n1011_) );
  AND2_X1 g653 ( .A1(new_n1010_), .A2(new_n1011_), .ZN(new_n1012_) );
  AND2_X1 g654 ( .A1(new_n1008_), .A2(new_n1012_), .ZN(new_n1013_) );
  AND2_X1 g655 ( .A1(new_n1004_), .A2(new_n1013_), .ZN(new_n1014_) );
  INV_X1 g656 ( .A(new_n655_), .ZN(new_n1015_) );
  OR2_X1 g657 ( .A1(G290), .A2(G1986), .ZN(new_n1016_) );
  AND2_X1 g658 ( .A1(new_n1016_), .A2(new_n718_), .ZN(new_n1017_) );
  OR2_X1 g659 ( .A1(new_n1009_), .A2(new_n1017_), .ZN(new_n1018_) );
  AND2_X1 g660 ( .A1(new_n1018_), .A2(new_n1015_), .ZN(new_n1019_) );
  INV_X1 g661 ( .A(new_n1019_), .ZN(new_n1020_) );
  OR2_X1 g662 ( .A1(new_n1020_), .A2(KEYINPUT39), .ZN(new_n1021_) );
  INV_X1 g663 ( .A(KEYINPUT39), .ZN(new_n1022_) );
  OR2_X1 g664 ( .A1(new_n1019_), .A2(new_n1022_), .ZN(new_n1023_) );
  AND2_X1 g665 ( .A1(new_n1023_), .A2(new_n1008_), .ZN(new_n1024_) );
  AND2_X1 g666 ( .A1(new_n1024_), .A2(new_n1021_), .ZN(new_n1025_) );
  OR2_X1 g667 ( .A1(new_n1025_), .A2(new_n700_), .ZN(new_n1026_) );
  AND2_X1 g668 ( .A1(new_n1026_), .A2(new_n1006_), .ZN(new_n1027_) );
  OR2_X1 g669 ( .A1(new_n1014_), .A2(new_n1027_), .ZN(new_n1028_) );
  XNOR2_X1 g670 ( .A(new_n1028_), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 g671 ( .A(G397), .ZN(new_n1031_) );
  AND2_X1 g672 ( .A1(new_n635_), .A2(new_n624_), .ZN(new_n1032_) );
  AND2_X1 g673 ( .A1(new_n1032_), .A2(KEYINPUT49), .ZN(new_n1033_) );
  INV_X1 g674 ( .A(new_n1033_), .ZN(new_n1034_) );
  OR2_X1 g675 ( .A1(new_n1032_), .A2(KEYINPUT49), .ZN(new_n1035_) );
  OR2_X1 g676 ( .A1(G401), .A2(new_n515_), .ZN(new_n1036_) );
  INV_X1 g677 ( .A(new_n1036_), .ZN(new_n1037_) );
  AND2_X1 g678 ( .A1(new_n1035_), .A2(new_n1037_), .ZN(new_n1038_) );
  AND2_X1 g679 ( .A1(new_n1038_), .A2(new_n1034_), .ZN(new_n1039_) );
  AND2_X1 g680 ( .A1(new_n883_), .A2(new_n1039_), .ZN(new_n1040_) );
  AND2_X1 g681 ( .A1(new_n1031_), .A2(new_n1040_), .ZN(G308) );
  INV_X1 g682 ( .A(G308), .ZN(G225) );
  assign   G231 = 1'b0;
  BUF_X1 g683 ( .A(G452), .Z(G350) );
  BUF_X1 g684 ( .A(G452), .Z(G335) );
  BUF_X1 g685 ( .A(G452), .Z(G409) );
  BUF_X1 g686 ( .A(G1083), .Z(G369) );
  BUF_X1 g687 ( .A(G1083), .Z(G367) );
  BUF_X1 g688 ( .A(G2066), .Z(G411) );
  BUF_X1 g689 ( .A(G2066), .Z(G337) );
  BUF_X1 g690 ( .A(G2066), .Z(G384) );
  BUF_X1 g691 ( .A(G452), .Z(G391) );
  OR2_X1 g692 ( .A1(new_n555_), .A2(new_n569_), .ZN(G321) );
  AND2_X1 g693 ( .A1(new_n571_), .A2(new_n572_), .ZN(G280) );
  AND2_X1 g694 ( .A1(new_n579_), .A2(new_n578_), .ZN(G323) );
  OR2_X1 g695 ( .A1(new_n893_), .A2(new_n894_), .ZN(G331) );
endmodule


