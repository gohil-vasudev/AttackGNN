module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n955_, new_n608_, new_n847_, new_n250_, new_n888_, new_n501_, new_n288_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n481_, new_n212_, new_n1073_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n903_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n1083_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n351_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n1028_, new_n508_, new_n714_, new_n194_, new_n483_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n398_, new_n301_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n473_, new_n140_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n996_, new_n621_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1084_, new_n1061_, new_n333_, new_n1002_, new_n290_, new_n834_, new_n369_, new_n448_, new_n867_, new_n1032_, new_n901_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n410_, new_n985_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n809_, new_n654_, new_n713_, new_n880_, new_n604_, new_n227_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n310_, new_n144_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n931_, new_n575_, new_n839_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n1001_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n936_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1074_, new_n748_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n730_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n408_, new_n470_, new_n213_, new_n769_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n627_, new_n704_, new_n195_, new_n567_, new_n576_, new_n1033_, new_n791_, new_n357_, new_n320_, new_n780_, new_n984_, new_n245_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1011_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n757_, new_n618_, new_n521_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_;

not g000 ( new_n138_, N1 );
not g001 ( new_n139_, keyIn_0_41 );
not g002 ( new_n140_, N77 );
and g003 ( new_n141_, new_n140_, N73 );
not g004 ( new_n142_, N73 );
and g005 ( new_n143_, new_n142_, N77 );
or g006 ( new_n144_, new_n141_, new_n143_ );
and g007 ( new_n145_, new_n144_, keyIn_0_6 );
not g008 ( new_n146_, new_n145_ );
or g009 ( new_n147_, new_n144_, keyIn_0_6 );
and g010 ( new_n148_, new_n146_, new_n147_ );
not g011 ( new_n149_, new_n148_ );
not g012 ( new_n150_, keyIn_0_5 );
not g013 ( new_n151_, N69 );
and g014 ( new_n152_, new_n151_, N65 );
not g015 ( new_n153_, N65 );
and g016 ( new_n154_, new_n153_, N69 );
or g017 ( new_n155_, new_n152_, new_n154_ );
and g018 ( new_n156_, new_n155_, new_n150_ );
not g019 ( new_n157_, new_n156_ );
or g020 ( new_n158_, new_n155_, new_n150_ );
and g021 ( new_n159_, new_n157_, new_n158_ );
not g022 ( new_n160_, new_n159_ );
and g023 ( new_n161_, new_n149_, new_n160_ );
and g024 ( new_n162_, new_n148_, new_n159_ );
or g025 ( new_n163_, new_n161_, new_n162_ );
not g026 ( new_n164_, new_n163_ );
not g027 ( new_n165_, N85 );
and g028 ( new_n166_, new_n165_, N81 );
not g029 ( new_n167_, N81 );
and g030 ( new_n168_, new_n167_, N85 );
or g031 ( new_n169_, new_n166_, new_n168_ );
not g032 ( new_n170_, new_n169_ );
not g033 ( new_n171_, N93 );
and g034 ( new_n172_, new_n171_, N89 );
not g035 ( new_n173_, N89 );
and g036 ( new_n174_, new_n173_, N93 );
or g037 ( new_n175_, new_n172_, new_n174_ );
and g038 ( new_n176_, new_n170_, new_n175_ );
not g039 ( new_n177_, new_n176_ );
or g040 ( new_n178_, new_n170_, new_n175_ );
and g041 ( new_n179_, new_n177_, new_n178_ );
not g042 ( new_n180_, new_n179_ );
and g043 ( new_n181_, new_n164_, new_n180_ );
and g044 ( new_n182_, new_n163_, new_n179_ );
or g045 ( new_n183_, new_n181_, new_n182_ );
and g046 ( new_n184_, N129, N137 );
not g047 ( new_n185_, new_n184_ );
and g048 ( new_n186_, new_n183_, new_n185_ );
not g049 ( new_n187_, new_n186_ );
or g050 ( new_n188_, new_n183_, new_n185_ );
and g051 ( new_n189_, new_n187_, new_n188_ );
not g052 ( new_n190_, N17 );
and g053 ( new_n191_, new_n190_, N1 );
and g054 ( new_n192_, new_n138_, N17 );
or g055 ( new_n193_, new_n191_, new_n192_ );
not g056 ( new_n194_, new_n193_ );
not g057 ( new_n195_, N49 );
and g058 ( new_n196_, new_n195_, N33 );
not g059 ( new_n197_, N33 );
and g060 ( new_n198_, new_n197_, N49 );
or g061 ( new_n199_, new_n196_, new_n198_ );
and g062 ( new_n200_, new_n194_, new_n199_ );
not g063 ( new_n201_, new_n200_ );
or g064 ( new_n202_, new_n194_, new_n199_ );
and g065 ( new_n203_, new_n201_, new_n202_ );
not g066 ( new_n204_, new_n203_ );
and g067 ( new_n205_, new_n189_, new_n204_ );
not g068 ( new_n206_, new_n205_ );
or g069 ( new_n207_, new_n189_, new_n204_ );
and g070 ( new_n208_, new_n206_, new_n207_ );
not g071 ( new_n209_, new_n208_ );
not g072 ( new_n210_, keyIn_0_7 );
not g073 ( new_n211_, N125 );
and g074 ( new_n212_, new_n211_, N121 );
not g075 ( new_n213_, N121 );
and g076 ( new_n214_, new_n213_, N125 );
or g077 ( new_n215_, new_n212_, new_n214_ );
and g078 ( new_n216_, new_n215_, new_n210_ );
not g079 ( new_n217_, new_n216_ );
or g080 ( new_n218_, new_n215_, new_n210_ );
and g081 ( new_n219_, new_n217_, new_n218_ );
not g082 ( new_n220_, N117 );
and g083 ( new_n221_, new_n220_, N113 );
not g084 ( new_n222_, N113 );
and g085 ( new_n223_, new_n222_, N117 );
or g086 ( new_n224_, new_n221_, new_n223_ );
not g087 ( new_n225_, new_n224_ );
and g088 ( new_n226_, new_n219_, new_n225_ );
not g089 ( new_n227_, new_n226_ );
or g090 ( new_n228_, new_n219_, new_n225_ );
and g091 ( new_n229_, new_n227_, new_n228_ );
not g092 ( new_n230_, new_n229_ );
and g093 ( new_n231_, new_n230_, keyIn_0_19 );
not g094 ( new_n232_, new_n231_ );
or g095 ( new_n233_, new_n230_, keyIn_0_19 );
and g096 ( new_n234_, new_n232_, new_n233_ );
not g097 ( new_n235_, keyIn_0_18 );
not g098 ( new_n236_, N109 );
and g099 ( new_n237_, new_n236_, N105 );
not g100 ( new_n238_, N105 );
and g101 ( new_n239_, new_n238_, N109 );
or g102 ( new_n240_, new_n237_, new_n239_ );
not g103 ( new_n241_, new_n240_ );
not g104 ( new_n242_, N101 );
and g105 ( new_n243_, new_n242_, N97 );
not g106 ( new_n244_, N97 );
and g107 ( new_n245_, new_n244_, N101 );
or g108 ( new_n246_, new_n243_, new_n245_ );
and g109 ( new_n247_, new_n241_, new_n246_ );
not g110 ( new_n248_, new_n247_ );
or g111 ( new_n249_, new_n241_, new_n246_ );
and g112 ( new_n250_, new_n248_, new_n249_ );
not g113 ( new_n251_, new_n250_ );
and g114 ( new_n252_, new_n251_, new_n235_ );
and g115 ( new_n253_, new_n250_, keyIn_0_18 );
or g116 ( new_n254_, new_n252_, new_n253_ );
not g117 ( new_n255_, new_n254_ );
or g118 ( new_n256_, new_n234_, new_n255_ );
and g119 ( new_n257_, new_n234_, new_n255_ );
not g120 ( new_n258_, new_n257_ );
and g121 ( new_n259_, new_n258_, new_n256_ );
and g122 ( new_n260_, new_n259_, keyIn_0_22 );
not g123 ( new_n261_, keyIn_0_22 );
not g124 ( new_n262_, new_n259_ );
and g125 ( new_n263_, new_n262_, new_n261_ );
or g126 ( new_n264_, new_n263_, new_n260_ );
and g127 ( new_n265_, new_n264_, keyIn_0_8 );
not g128 ( new_n266_, keyIn_0_8 );
not g129 ( new_n267_, new_n260_ );
or g130 ( new_n268_, new_n259_, keyIn_0_22 );
and g131 ( new_n269_, new_n267_, new_n268_ );
and g132 ( new_n270_, new_n269_, new_n266_ );
or g133 ( new_n271_, new_n265_, new_n270_ );
and g134 ( new_n272_, N130, N137 );
not g135 ( new_n273_, new_n272_ );
and g136 ( new_n274_, new_n271_, new_n273_ );
or g137 ( new_n275_, new_n269_, new_n266_ );
or g138 ( new_n276_, new_n264_, keyIn_0_8 );
and g139 ( new_n277_, new_n276_, new_n275_ );
and g140 ( new_n278_, new_n277_, new_n272_ );
or g141 ( new_n279_, new_n274_, new_n278_ );
not g142 ( new_n280_, N21 );
and g143 ( new_n281_, new_n280_, N5 );
not g144 ( new_n282_, N5 );
and g145 ( new_n283_, new_n282_, N21 );
or g146 ( new_n284_, new_n281_, new_n283_ );
and g147 ( new_n285_, new_n284_, keyIn_0_12 );
not g148 ( new_n286_, new_n285_ );
or g149 ( new_n287_, new_n284_, keyIn_0_12 );
and g150 ( new_n288_, new_n286_, new_n287_ );
not g151 ( new_n289_, new_n288_ );
not g152 ( new_n290_, N53 );
and g153 ( new_n291_, new_n290_, N37 );
not g154 ( new_n292_, N37 );
and g155 ( new_n293_, new_n292_, N53 );
or g156 ( new_n294_, new_n291_, new_n293_ );
and g157 ( new_n295_, new_n294_, keyIn_0_13 );
not g158 ( new_n296_, new_n295_ );
or g159 ( new_n297_, new_n294_, keyIn_0_13 );
and g160 ( new_n298_, new_n296_, new_n297_ );
and g161 ( new_n299_, new_n289_, new_n298_ );
not g162 ( new_n300_, new_n299_ );
or g163 ( new_n301_, new_n289_, new_n298_ );
and g164 ( new_n302_, new_n300_, new_n301_ );
or g165 ( new_n303_, new_n279_, new_n302_ );
or g166 ( new_n304_, new_n277_, new_n272_ );
or g167 ( new_n305_, new_n271_, new_n273_ );
and g168 ( new_n306_, new_n305_, new_n304_ );
not g169 ( new_n307_, new_n302_ );
or g170 ( new_n308_, new_n306_, new_n307_ );
and g171 ( new_n309_, new_n303_, new_n308_ );
and g172 ( new_n310_, new_n309_, new_n209_ );
not g173 ( new_n311_, keyIn_0_23 );
and g174 ( new_n312_, N132, N137 );
not g175 ( new_n313_, keyIn_0_9 );
or g176 ( new_n314_, new_n234_, new_n179_ );
and g177 ( new_n315_, new_n234_, new_n179_ );
not g178 ( new_n316_, new_n315_ );
and g179 ( new_n317_, new_n316_, new_n314_ );
or g180 ( new_n318_, new_n317_, new_n313_ );
and g181 ( new_n319_, new_n317_, new_n313_ );
not g182 ( new_n320_, new_n319_ );
and g183 ( new_n321_, new_n320_, new_n318_ );
and g184 ( new_n322_, new_n321_, new_n312_ );
not g185 ( new_n323_, new_n312_ );
not g186 ( new_n324_, new_n317_ );
and g187 ( new_n325_, new_n324_, keyIn_0_9 );
or g188 ( new_n326_, new_n325_, new_n319_ );
and g189 ( new_n327_, new_n326_, new_n323_ );
or g190 ( new_n328_, new_n327_, new_n322_ );
and g191 ( new_n329_, new_n328_, new_n311_ );
or g192 ( new_n330_, new_n326_, new_n323_ );
or g193 ( new_n331_, new_n321_, new_n312_ );
and g194 ( new_n332_, new_n330_, new_n331_ );
and g195 ( new_n333_, new_n332_, keyIn_0_23 );
or g196 ( new_n334_, new_n329_, new_n333_ );
not g197 ( new_n335_, N29 );
and g198 ( new_n336_, new_n335_, N13 );
not g199 ( new_n337_, N13 );
and g200 ( new_n338_, new_n337_, N29 );
or g201 ( new_n339_, new_n336_, new_n338_ );
and g202 ( new_n340_, new_n339_, keyIn_0_14 );
not g203 ( new_n341_, new_n340_ );
or g204 ( new_n342_, new_n339_, keyIn_0_14 );
and g205 ( new_n343_, new_n341_, new_n342_ );
not g206 ( new_n344_, new_n343_ );
not g207 ( new_n345_, N61 );
and g208 ( new_n346_, new_n345_, N45 );
not g209 ( new_n347_, N45 );
and g210 ( new_n348_, new_n347_, N61 );
or g211 ( new_n349_, new_n346_, new_n348_ );
not g212 ( new_n350_, new_n349_ );
and g213 ( new_n351_, new_n344_, new_n350_ );
and g214 ( new_n352_, new_n343_, new_n349_ );
or g215 ( new_n353_, new_n351_, new_n352_ );
not g216 ( new_n354_, new_n353_ );
or g217 ( new_n355_, new_n334_, new_n354_ );
or g218 ( new_n356_, new_n332_, keyIn_0_23 );
or g219 ( new_n357_, new_n328_, new_n311_ );
and g220 ( new_n358_, new_n357_, new_n356_ );
or g221 ( new_n359_, new_n358_, new_n353_ );
and g222 ( new_n360_, new_n355_, new_n359_ );
and g223 ( new_n361_, new_n255_, new_n163_ );
and g224 ( new_n362_, new_n164_, new_n254_ );
or g225 ( new_n363_, new_n361_, new_n362_ );
and g226 ( new_n364_, N131, N137 );
not g227 ( new_n365_, new_n364_ );
and g228 ( new_n366_, new_n363_, new_n365_ );
not g229 ( new_n367_, new_n366_ );
or g230 ( new_n368_, new_n363_, new_n365_ );
and g231 ( new_n369_, new_n367_, new_n368_ );
not g232 ( new_n370_, N25 );
and g233 ( new_n371_, new_n370_, N9 );
not g234 ( new_n372_, N9 );
and g235 ( new_n373_, new_n372_, N25 );
or g236 ( new_n374_, new_n371_, new_n373_ );
not g237 ( new_n375_, new_n374_ );
not g238 ( new_n376_, N57 );
and g239 ( new_n377_, new_n376_, N41 );
not g240 ( new_n378_, N41 );
and g241 ( new_n379_, new_n378_, N57 );
or g242 ( new_n380_, new_n377_, new_n379_ );
and g243 ( new_n381_, new_n375_, new_n380_ );
not g244 ( new_n382_, new_n381_ );
or g245 ( new_n383_, new_n375_, new_n380_ );
and g246 ( new_n384_, new_n382_, new_n383_ );
not g247 ( new_n385_, new_n384_ );
and g248 ( new_n386_, new_n369_, new_n385_ );
not g249 ( new_n387_, new_n386_ );
or g250 ( new_n388_, new_n369_, new_n385_ );
and g251 ( new_n389_, new_n387_, new_n388_ );
and g252 ( new_n390_, new_n389_, keyIn_0_24 );
not g253 ( new_n391_, new_n390_ );
or g254 ( new_n392_, new_n389_, keyIn_0_24 );
and g255 ( new_n393_, new_n391_, new_n392_ );
and g256 ( new_n394_, new_n393_, keyIn_0_26 );
not g257 ( new_n395_, new_n394_ );
or g258 ( new_n396_, new_n393_, keyIn_0_26 );
and g259 ( new_n397_, new_n395_, new_n396_ );
and g260 ( new_n398_, new_n360_, new_n397_ );
and g261 ( new_n399_, new_n398_, new_n310_ );
and g262 ( new_n400_, new_n399_, keyIn_0_36 );
not g263 ( new_n401_, new_n400_ );
or g264 ( new_n402_, new_n399_, keyIn_0_36 );
and g265 ( new_n403_, new_n401_, new_n402_ );
and g266 ( new_n404_, new_n306_, new_n307_ );
and g267 ( new_n405_, new_n279_, new_n302_ );
or g268 ( new_n406_, new_n405_, new_n404_ );
and g269 ( new_n407_, new_n393_, new_n208_ );
and g270 ( new_n408_, new_n406_, new_n407_ );
and g271 ( new_n409_, new_n209_, keyIn_0_25 );
not g272 ( new_n410_, new_n409_ );
or g273 ( new_n411_, new_n209_, keyIn_0_25 );
and g274 ( new_n412_, new_n410_, new_n411_ );
or g275 ( new_n413_, new_n412_, new_n393_ );
not g276 ( new_n414_, new_n413_ );
and g277 ( new_n415_, new_n309_, new_n414_ );
or g278 ( new_n416_, new_n408_, new_n415_ );
and g279 ( new_n417_, new_n416_, new_n360_ );
and g280 ( new_n418_, new_n358_, new_n353_ );
and g281 ( new_n419_, new_n334_, new_n354_ );
or g282 ( new_n420_, new_n419_, new_n418_ );
and g283 ( new_n421_, new_n309_, new_n407_ );
and g284 ( new_n422_, new_n421_, new_n420_ );
or g285 ( new_n423_, new_n417_, new_n422_ );
or g286 ( new_n424_, new_n403_, new_n423_ );
not g287 ( new_n425_, keyIn_0_17 );
not g288 ( new_n426_, keyIn_0_2 );
and g289 ( new_n427_, new_n292_, N33 );
and g290 ( new_n428_, new_n197_, N37 );
or g291 ( new_n429_, new_n427_, new_n428_ );
and g292 ( new_n430_, new_n429_, new_n426_ );
or g293 ( new_n431_, new_n197_, N37 );
or g294 ( new_n432_, new_n292_, N33 );
and g295 ( new_n433_, new_n431_, new_n432_ );
and g296 ( new_n434_, new_n433_, keyIn_0_2 );
or g297 ( new_n435_, new_n430_, new_n434_ );
and g298 ( new_n436_, new_n347_, N41 );
and g299 ( new_n437_, new_n378_, N45 );
or g300 ( new_n438_, new_n436_, new_n437_ );
or g301 ( new_n439_, new_n438_, keyIn_0_3 );
not g302 ( new_n440_, keyIn_0_3 );
or g303 ( new_n441_, new_n378_, N45 );
or g304 ( new_n442_, new_n347_, N41 );
and g305 ( new_n443_, new_n441_, new_n442_ );
or g306 ( new_n444_, new_n443_, new_n440_ );
and g307 ( new_n445_, new_n439_, new_n444_ );
and g308 ( new_n446_, new_n435_, new_n445_ );
or g309 ( new_n447_, new_n433_, keyIn_0_2 );
or g310 ( new_n448_, new_n429_, new_n426_ );
and g311 ( new_n449_, new_n448_, new_n447_ );
and g312 ( new_n450_, new_n443_, new_n440_ );
and g313 ( new_n451_, new_n438_, keyIn_0_3 );
or g314 ( new_n452_, new_n451_, new_n450_ );
and g315 ( new_n453_, new_n452_, new_n449_ );
or g316 ( new_n454_, new_n446_, new_n453_ );
and g317 ( new_n455_, new_n454_, new_n425_ );
or g318 ( new_n456_, new_n452_, new_n449_ );
or g319 ( new_n457_, new_n435_, new_n445_ );
and g320 ( new_n458_, new_n456_, new_n457_ );
and g321 ( new_n459_, new_n458_, keyIn_0_17 );
or g322 ( new_n460_, new_n455_, new_n459_ );
and g323 ( new_n461_, new_n337_, N9 );
and g324 ( new_n462_, new_n372_, N13 );
or g325 ( new_n463_, new_n461_, new_n462_ );
not g326 ( new_n464_, new_n463_ );
and g327 ( new_n465_, new_n282_, N1 );
and g328 ( new_n466_, new_n138_, N5 );
or g329 ( new_n467_, new_n465_, new_n466_ );
and g330 ( new_n468_, new_n464_, new_n467_ );
not g331 ( new_n469_, new_n468_ );
or g332 ( new_n470_, new_n464_, new_n467_ );
and g333 ( new_n471_, new_n469_, new_n470_ );
not g334 ( new_n472_, new_n471_ );
and g335 ( new_n473_, new_n472_, keyIn_0_16 );
not g336 ( new_n474_, new_n473_ );
or g337 ( new_n475_, new_n472_, keyIn_0_16 );
and g338 ( new_n476_, new_n474_, new_n475_ );
and g339 ( new_n477_, new_n460_, new_n476_ );
or g340 ( new_n478_, new_n458_, keyIn_0_17 );
or g341 ( new_n479_, new_n454_, new_n425_ );
and g342 ( new_n480_, new_n478_, new_n479_ );
not g343 ( new_n481_, new_n476_ );
and g344 ( new_n482_, new_n480_, new_n481_ );
or g345 ( new_n483_, new_n477_, new_n482_ );
and g346 ( new_n484_, new_n483_, keyIn_0_21 );
not g347 ( new_n485_, keyIn_0_21 );
or g348 ( new_n486_, new_n480_, new_n481_ );
or g349 ( new_n487_, new_n460_, new_n476_ );
and g350 ( new_n488_, new_n487_, new_n486_ );
and g351 ( new_n489_, new_n488_, new_n485_ );
or g352 ( new_n490_, new_n484_, new_n489_ );
and g353 ( new_n491_, new_n490_, keyIn_0_10 );
not g354 ( new_n492_, keyIn_0_10 );
or g355 ( new_n493_, new_n488_, new_n485_ );
or g356 ( new_n494_, new_n483_, keyIn_0_21 );
and g357 ( new_n495_, new_n494_, new_n493_ );
and g358 ( new_n496_, new_n495_, new_n492_ );
or g359 ( new_n497_, new_n491_, new_n496_ );
and g360 ( new_n498_, N135, N137 );
not g361 ( new_n499_, new_n498_ );
and g362 ( new_n500_, new_n497_, new_n499_ );
or g363 ( new_n501_, new_n495_, new_n492_ );
or g364 ( new_n502_, new_n490_, keyIn_0_10 );
and g365 ( new_n503_, new_n502_, new_n501_ );
and g366 ( new_n504_, new_n503_, new_n498_ );
or g367 ( new_n505_, new_n500_, new_n504_ );
and g368 ( new_n506_, new_n173_, N73 );
and g369 ( new_n507_, new_n142_, N89 );
or g370 ( new_n508_, new_n506_, new_n507_ );
not g371 ( new_n509_, new_n508_ );
and g372 ( new_n510_, new_n213_, N105 );
and g373 ( new_n511_, new_n238_, N121 );
or g374 ( new_n512_, new_n510_, new_n511_ );
and g375 ( new_n513_, new_n509_, new_n512_ );
not g376 ( new_n514_, new_n513_ );
or g377 ( new_n515_, new_n509_, new_n512_ );
and g378 ( new_n516_, new_n514_, new_n515_ );
not g379 ( new_n517_, new_n516_ );
and g380 ( new_n518_, new_n517_, keyIn_0_20 );
not g381 ( new_n519_, new_n518_ );
or g382 ( new_n520_, new_n517_, keyIn_0_20 );
and g383 ( new_n521_, new_n519_, new_n520_ );
not g384 ( new_n522_, new_n521_ );
and g385 ( new_n523_, new_n505_, new_n522_ );
or g386 ( new_n524_, new_n503_, new_n498_ );
or g387 ( new_n525_, new_n497_, new_n499_ );
and g388 ( new_n526_, new_n525_, new_n524_ );
and g389 ( new_n527_, new_n526_, new_n521_ );
or g390 ( new_n528_, new_n523_, new_n527_ );
and g391 ( new_n529_, new_n424_, new_n528_ );
and g392 ( new_n530_, new_n335_, N25 );
and g393 ( new_n531_, new_n370_, N29 );
or g394 ( new_n532_, new_n530_, new_n531_ );
and g395 ( new_n533_, new_n532_, keyIn_0_1 );
not g396 ( new_n534_, new_n533_ );
or g397 ( new_n535_, new_n532_, keyIn_0_1 );
and g398 ( new_n536_, new_n534_, new_n535_ );
not g399 ( new_n537_, new_n536_ );
not g400 ( new_n538_, keyIn_0_0 );
and g401 ( new_n539_, new_n280_, N17 );
and g402 ( new_n540_, new_n190_, N21 );
or g403 ( new_n541_, new_n539_, new_n540_ );
and g404 ( new_n542_, new_n541_, new_n538_ );
not g405 ( new_n543_, new_n542_ );
or g406 ( new_n544_, new_n541_, new_n538_ );
and g407 ( new_n545_, new_n543_, new_n544_ );
and g408 ( new_n546_, new_n537_, new_n545_ );
not g409 ( new_n547_, new_n546_ );
or g410 ( new_n548_, new_n537_, new_n545_ );
and g411 ( new_n549_, new_n547_, new_n548_ );
and g412 ( new_n550_, new_n345_, N57 );
and g413 ( new_n551_, new_n376_, N61 );
or g414 ( new_n552_, new_n550_, new_n551_ );
and g415 ( new_n553_, new_n552_, keyIn_0_4 );
not g416 ( new_n554_, new_n553_ );
or g417 ( new_n555_, new_n552_, keyIn_0_4 );
and g418 ( new_n556_, new_n554_, new_n555_ );
and g419 ( new_n557_, new_n290_, N49 );
and g420 ( new_n558_, new_n195_, N53 );
or g421 ( new_n559_, new_n557_, new_n558_ );
and g422 ( new_n560_, new_n556_, new_n559_ );
not g423 ( new_n561_, new_n560_ );
or g424 ( new_n562_, new_n556_, new_n559_ );
and g425 ( new_n563_, new_n561_, new_n562_ );
not g426 ( new_n564_, new_n563_ );
and g427 ( new_n565_, new_n549_, new_n564_ );
not g428 ( new_n566_, new_n549_ );
and g429 ( new_n567_, new_n566_, new_n563_ );
or g430 ( new_n568_, new_n567_, new_n565_ );
or g431 ( new_n569_, new_n568_, keyIn_0_11 );
and g432 ( new_n570_, new_n568_, keyIn_0_11 );
not g433 ( new_n571_, new_n570_ );
and g434 ( new_n572_, new_n571_, new_n569_ );
and g435 ( new_n573_, N136, N137 );
and g436 ( new_n574_, new_n572_, new_n573_ );
not g437 ( new_n575_, new_n574_ );
or g438 ( new_n576_, new_n572_, new_n573_ );
and g439 ( new_n577_, new_n575_, new_n576_ );
and g440 ( new_n578_, new_n171_, N77 );
and g441 ( new_n579_, new_n140_, N93 );
or g442 ( new_n580_, new_n578_, new_n579_ );
not g443 ( new_n581_, new_n580_ );
and g444 ( new_n582_, new_n211_, N109 );
and g445 ( new_n583_, new_n236_, N125 );
or g446 ( new_n584_, new_n582_, new_n583_ );
and g447 ( new_n585_, new_n581_, new_n584_ );
not g448 ( new_n586_, new_n585_ );
or g449 ( new_n587_, new_n581_, new_n584_ );
and g450 ( new_n588_, new_n586_, new_n587_ );
or g451 ( new_n589_, new_n577_, new_n588_ );
not g452 ( new_n590_, new_n569_ );
or g453 ( new_n591_, new_n590_, new_n570_ );
not g454 ( new_n592_, new_n573_ );
and g455 ( new_n593_, new_n591_, new_n592_ );
or g456 ( new_n594_, new_n593_, new_n574_ );
not g457 ( new_n595_, new_n588_ );
or g458 ( new_n596_, new_n594_, new_n595_ );
and g459 ( new_n597_, new_n589_, new_n596_ );
and g460 ( new_n598_, new_n460_, new_n563_ );
and g461 ( new_n599_, new_n480_, new_n564_ );
or g462 ( new_n600_, new_n598_, new_n599_ );
and g463 ( new_n601_, N134, N137 );
not g464 ( new_n602_, new_n601_ );
and g465 ( new_n603_, new_n600_, new_n602_ );
not g466 ( new_n604_, new_n603_ );
or g467 ( new_n605_, new_n600_, new_n602_ );
and g468 ( new_n606_, new_n604_, new_n605_ );
and g469 ( new_n607_, new_n165_, N69 );
and g470 ( new_n608_, new_n151_, N85 );
or g471 ( new_n609_, new_n607_, new_n608_ );
not g472 ( new_n610_, new_n609_ );
and g473 ( new_n611_, new_n220_, N101 );
and g474 ( new_n612_, new_n242_, N117 );
or g475 ( new_n613_, new_n611_, new_n612_ );
and g476 ( new_n614_, new_n610_, new_n613_ );
not g477 ( new_n615_, new_n614_ );
or g478 ( new_n616_, new_n610_, new_n613_ );
and g479 ( new_n617_, new_n615_, new_n616_ );
not g480 ( new_n618_, new_n617_ );
and g481 ( new_n619_, new_n606_, new_n618_ );
not g482 ( new_n620_, new_n619_ );
or g483 ( new_n621_, new_n606_, new_n618_ );
and g484 ( new_n622_, new_n620_, new_n621_ );
and g485 ( new_n623_, new_n481_, new_n549_ );
and g486 ( new_n624_, new_n566_, new_n476_ );
or g487 ( new_n625_, new_n623_, new_n624_ );
and g488 ( new_n626_, N133, N137 );
not g489 ( new_n627_, new_n626_ );
and g490 ( new_n628_, new_n625_, new_n627_ );
or g491 ( new_n629_, new_n566_, new_n476_ );
not g492 ( new_n630_, new_n624_ );
and g493 ( new_n631_, new_n630_, new_n629_ );
and g494 ( new_n632_, new_n631_, new_n626_ );
or g495 ( new_n633_, new_n628_, new_n632_ );
not g496 ( new_n634_, keyIn_0_15 );
and g497 ( new_n635_, new_n222_, N97 );
and g498 ( new_n636_, new_n244_, N113 );
or g499 ( new_n637_, new_n635_, new_n636_ );
and g500 ( new_n638_, new_n637_, new_n634_ );
not g501 ( new_n639_, new_n638_ );
or g502 ( new_n640_, new_n637_, new_n634_ );
and g503 ( new_n641_, new_n639_, new_n640_ );
and g504 ( new_n642_, new_n167_, N65 );
and g505 ( new_n643_, new_n153_, N81 );
or g506 ( new_n644_, new_n642_, new_n643_ );
not g507 ( new_n645_, new_n644_ );
and g508 ( new_n646_, new_n641_, new_n645_ );
not g509 ( new_n647_, new_n646_ );
or g510 ( new_n648_, new_n641_, new_n645_ );
and g511 ( new_n649_, new_n647_, new_n648_ );
and g512 ( new_n650_, new_n633_, new_n649_ );
or g513 ( new_n651_, new_n631_, new_n626_ );
or g514 ( new_n652_, new_n625_, new_n627_ );
and g515 ( new_n653_, new_n652_, new_n651_ );
not g516 ( new_n654_, new_n649_ );
and g517 ( new_n655_, new_n653_, new_n654_ );
or g518 ( new_n656_, new_n650_, new_n655_ );
and g519 ( new_n657_, new_n622_, new_n656_ );
and g520 ( new_n658_, new_n597_, new_n657_ );
and g521 ( new_n659_, new_n529_, new_n658_ );
and g522 ( new_n660_, new_n659_, new_n209_ );
not g523 ( new_n661_, new_n660_ );
and g524 ( new_n662_, new_n661_, new_n139_ );
and g525 ( new_n663_, new_n660_, keyIn_0_41 );
or g526 ( new_n664_, new_n662_, new_n663_ );
not g527 ( new_n665_, new_n664_ );
and g528 ( new_n666_, new_n665_, new_n138_ );
and g529 ( new_n667_, new_n664_, N1 );
or g530 ( N724, new_n666_, new_n667_ );
and g531 ( new_n669_, new_n659_, new_n406_ );
not g532 ( new_n670_, new_n669_ );
and g533 ( new_n671_, new_n670_, keyIn_0_42 );
not g534 ( new_n672_, new_n671_ );
or g535 ( new_n673_, new_n670_, keyIn_0_42 );
and g536 ( new_n674_, new_n672_, new_n673_ );
not g537 ( new_n675_, new_n674_ );
and g538 ( new_n676_, new_n675_, N5 );
and g539 ( new_n677_, new_n674_, new_n282_ );
or g540 ( N725, new_n676_, new_n677_ );
not g541 ( new_n679_, new_n393_ );
and g542 ( new_n680_, new_n659_, new_n679_ );
not g543 ( new_n681_, new_n680_ );
and g544 ( new_n682_, new_n681_, N9 );
and g545 ( new_n683_, new_n680_, new_n372_ );
or g546 ( N726, new_n682_, new_n683_ );
and g547 ( new_n685_, new_n659_, new_n420_ );
not g548 ( new_n686_, new_n685_ );
and g549 ( new_n687_, new_n686_, N13 );
and g550 ( new_n688_, new_n685_, new_n337_ );
or g551 ( N727, new_n687_, new_n688_ );
or g552 ( new_n690_, new_n526_, new_n521_ );
or g553 ( new_n691_, new_n505_, new_n522_ );
and g554 ( new_n692_, new_n691_, new_n690_ );
and g555 ( new_n693_, new_n594_, new_n595_ );
and g556 ( new_n694_, new_n577_, new_n588_ );
or g557 ( new_n695_, new_n694_, new_n693_ );
and g558 ( new_n696_, new_n695_, new_n657_ );
and g559 ( new_n697_, new_n692_, new_n696_ );
and g560 ( new_n698_, new_n424_, new_n697_ );
and g561 ( new_n699_, new_n698_, new_n209_ );
not g562 ( new_n700_, new_n699_ );
and g563 ( new_n701_, new_n700_, N17 );
and g564 ( new_n702_, new_n699_, new_n190_ );
or g565 ( new_n703_, new_n701_, new_n702_ );
not g566 ( new_n704_, new_n703_ );
or g567 ( new_n705_, new_n704_, keyIn_0_54 );
not g568 ( new_n706_, keyIn_0_54 );
or g569 ( new_n707_, new_n703_, new_n706_ );
and g570 ( N728, new_n705_, new_n707_ );
and g571 ( new_n709_, new_n698_, new_n406_ );
not g572 ( new_n710_, new_n709_ );
and g573 ( new_n711_, new_n710_, N21 );
and g574 ( new_n712_, new_n709_, new_n280_ );
or g575 ( new_n713_, new_n711_, new_n712_ );
not g576 ( new_n714_, new_n713_ );
or g577 ( new_n715_, new_n714_, keyIn_0_55 );
not g578 ( new_n716_, keyIn_0_55 );
or g579 ( new_n717_, new_n713_, new_n716_ );
and g580 ( N729, new_n715_, new_n717_ );
and g581 ( new_n719_, new_n698_, new_n679_ );
not g582 ( new_n720_, new_n719_ );
and g583 ( new_n721_, new_n720_, N25 );
and g584 ( new_n722_, new_n719_, new_n370_ );
or g585 ( N730, new_n721_, new_n722_ );
and g586 ( new_n724_, new_n698_, new_n420_ );
not g587 ( new_n725_, new_n724_ );
and g588 ( new_n726_, new_n725_, keyIn_0_43 );
not g589 ( new_n727_, new_n726_ );
or g590 ( new_n728_, new_n725_, keyIn_0_43 );
and g591 ( new_n729_, new_n727_, new_n728_ );
not g592 ( new_n730_, new_n729_ );
and g593 ( new_n731_, new_n730_, new_n335_ );
and g594 ( new_n732_, new_n729_, N29 );
or g595 ( N731, new_n731_, new_n732_ );
not g596 ( new_n734_, new_n622_ );
or g597 ( new_n735_, new_n653_, new_n654_ );
or g598 ( new_n736_, new_n633_, new_n649_ );
and g599 ( new_n737_, new_n736_, new_n735_ );
and g600 ( new_n738_, new_n597_, new_n737_ );
and g601 ( new_n739_, new_n738_, new_n734_ );
and g602 ( new_n740_, new_n529_, new_n739_ );
and g603 ( new_n741_, new_n740_, new_n209_ );
not g604 ( new_n742_, new_n741_ );
and g605 ( new_n743_, new_n742_, N33 );
and g606 ( new_n744_, new_n741_, new_n197_ );
or g607 ( new_n745_, new_n743_, new_n744_ );
not g608 ( new_n746_, new_n745_ );
or g609 ( new_n747_, new_n746_, keyIn_0_56 );
not g610 ( new_n748_, keyIn_0_56 );
or g611 ( new_n749_, new_n745_, new_n748_ );
and g612 ( N732, new_n747_, new_n749_ );
and g613 ( new_n751_, new_n740_, new_n406_ );
not g614 ( new_n752_, new_n751_ );
and g615 ( new_n753_, new_n752_, N37 );
and g616 ( new_n754_, new_n751_, new_n292_ );
or g617 ( new_n755_, new_n753_, new_n754_ );
not g618 ( new_n756_, new_n755_ );
and g619 ( new_n757_, new_n756_, keyIn_0_57 );
not g620 ( new_n758_, keyIn_0_57 );
and g621 ( new_n759_, new_n755_, new_n758_ );
or g622 ( N733, new_n757_, new_n759_ );
and g623 ( new_n761_, new_n740_, new_n679_ );
not g624 ( new_n762_, new_n761_ );
and g625 ( new_n763_, new_n762_, keyIn_0_44 );
not g626 ( new_n764_, new_n763_ );
or g627 ( new_n765_, new_n762_, keyIn_0_44 );
and g628 ( new_n766_, new_n764_, new_n765_ );
not g629 ( new_n767_, new_n766_ );
and g630 ( new_n768_, new_n767_, new_n378_ );
and g631 ( new_n769_, new_n766_, N41 );
or g632 ( N734, new_n768_, new_n769_ );
not g633 ( new_n771_, keyIn_0_58 );
not g634 ( new_n772_, keyIn_0_45 );
not g635 ( new_n773_, keyIn_0_36 );
or g636 ( new_n774_, new_n406_, new_n208_ );
not g637 ( new_n775_, new_n397_ );
or g638 ( new_n776_, new_n420_, new_n775_ );
or g639 ( new_n777_, new_n774_, new_n776_ );
and g640 ( new_n778_, new_n777_, new_n773_ );
or g641 ( new_n779_, new_n778_, new_n400_ );
not g642 ( new_n780_, new_n407_ );
or g643 ( new_n781_, new_n309_, new_n780_ );
or g644 ( new_n782_, new_n406_, new_n413_ );
and g645 ( new_n783_, new_n782_, new_n781_ );
or g646 ( new_n784_, new_n783_, new_n420_ );
not g647 ( new_n785_, new_n422_ );
and g648 ( new_n786_, new_n784_, new_n785_ );
and g649 ( new_n787_, new_n779_, new_n786_ );
or g650 ( new_n788_, new_n787_, new_n692_ );
not g651 ( new_n789_, new_n739_ );
or g652 ( new_n790_, new_n788_, new_n789_ );
or g653 ( new_n791_, new_n790_, new_n360_ );
and g654 ( new_n792_, new_n791_, new_n772_ );
and g655 ( new_n793_, new_n740_, new_n420_ );
and g656 ( new_n794_, new_n793_, keyIn_0_45 );
or g657 ( new_n795_, new_n792_, new_n794_ );
or g658 ( new_n796_, new_n795_, new_n347_ );
or g659 ( new_n797_, new_n793_, keyIn_0_45 );
or g660 ( new_n798_, new_n791_, new_n772_ );
and g661 ( new_n799_, new_n798_, new_n797_ );
or g662 ( new_n800_, new_n799_, N45 );
and g663 ( new_n801_, new_n796_, new_n800_ );
or g664 ( new_n802_, new_n801_, new_n771_ );
and g665 ( new_n803_, new_n799_, N45 );
and g666 ( new_n804_, new_n795_, new_n347_ );
or g667 ( new_n805_, new_n803_, new_n804_ );
or g668 ( new_n806_, new_n805_, keyIn_0_58 );
and g669 ( N735, new_n806_, new_n802_ );
not g670 ( new_n808_, keyIn_0_39 );
and g671 ( new_n809_, new_n528_, keyIn_0_27 );
not g672 ( new_n810_, new_n809_ );
or g673 ( new_n811_, new_n528_, keyIn_0_27 );
and g674 ( new_n812_, new_n810_, new_n811_ );
not g675 ( new_n813_, new_n812_ );
and g676 ( new_n814_, new_n695_, new_n737_ );
and g677 ( new_n815_, new_n814_, new_n734_ );
and g678 ( new_n816_, new_n813_, new_n815_ );
and g679 ( new_n817_, new_n424_, new_n816_ );
not g680 ( new_n818_, new_n817_ );
and g681 ( new_n819_, new_n818_, new_n808_ );
and g682 ( new_n820_, new_n817_, keyIn_0_39 );
or g683 ( new_n821_, new_n819_, new_n820_ );
and g684 ( new_n822_, new_n821_, new_n209_ );
or g685 ( new_n823_, new_n822_, new_n195_ );
and g686 ( new_n824_, new_n822_, new_n195_ );
not g687 ( new_n825_, new_n824_ );
and g688 ( new_n826_, new_n825_, new_n823_ );
not g689 ( new_n827_, new_n826_ );
and g690 ( new_n828_, new_n827_, keyIn_0_59 );
not g691 ( new_n829_, keyIn_0_59 );
and g692 ( new_n830_, new_n826_, new_n829_ );
or g693 ( N736, new_n828_, new_n830_ );
not g694 ( new_n832_, keyIn_0_46 );
and g695 ( new_n833_, new_n821_, new_n406_ );
or g696 ( new_n834_, new_n833_, new_n832_ );
and g697 ( new_n835_, new_n833_, new_n832_ );
not g698 ( new_n836_, new_n835_ );
and g699 ( new_n837_, new_n836_, new_n834_ );
not g700 ( new_n838_, new_n837_ );
and g701 ( new_n839_, new_n838_, N53 );
and g702 ( new_n840_, new_n837_, new_n290_ );
or g703 ( N737, new_n839_, new_n840_ );
and g704 ( new_n842_, new_n821_, new_n679_ );
not g705 ( new_n843_, new_n842_ );
and g706 ( new_n844_, new_n843_, N57 );
and g707 ( new_n845_, new_n842_, new_n376_ );
or g708 ( N738, new_n844_, new_n845_ );
and g709 ( new_n847_, new_n821_, new_n420_ );
not g710 ( new_n848_, new_n847_ );
and g711 ( new_n849_, new_n848_, N61 );
and g712 ( new_n850_, new_n847_, new_n345_ );
or g713 ( N739, new_n849_, new_n850_ );
not g714 ( new_n852_, keyIn_0_37 );
not g715 ( new_n853_, keyIn_0_31 );
and g716 ( new_n854_, new_n692_, new_n853_ );
not g717 ( new_n855_, new_n854_ );
or g718 ( new_n856_, new_n692_, new_n853_ );
and g719 ( new_n857_, new_n856_, new_n739_ );
and g720 ( new_n858_, new_n857_, new_n855_ );
and g721 ( new_n859_, new_n858_, new_n852_ );
and g722 ( new_n860_, new_n528_, keyIn_0_31 );
or g723 ( new_n861_, new_n860_, new_n789_ );
or g724 ( new_n862_, new_n861_, new_n854_ );
and g725 ( new_n863_, new_n862_, keyIn_0_37 );
and g726 ( new_n864_, new_n692_, keyIn_0_32 );
not g727 ( new_n865_, keyIn_0_32 );
and g728 ( new_n866_, new_n528_, new_n865_ );
or g729 ( new_n867_, new_n866_, new_n864_ );
not g730 ( new_n868_, keyIn_0_33 );
and g731 ( new_n869_, new_n597_, new_n868_ );
and g732 ( new_n870_, new_n695_, keyIn_0_33 );
or g733 ( new_n871_, new_n870_, new_n869_ );
and g734 ( new_n872_, new_n871_, new_n657_ );
and g735 ( new_n873_, new_n867_, new_n872_ );
not g736 ( new_n874_, keyIn_0_30 );
and g737 ( new_n875_, new_n597_, new_n874_ );
not g738 ( new_n876_, new_n875_ );
or g739 ( new_n877_, new_n597_, new_n874_ );
and g740 ( new_n878_, new_n737_, keyIn_0_29 );
not g741 ( new_n879_, keyIn_0_29 );
and g742 ( new_n880_, new_n656_, new_n879_ );
or g743 ( new_n881_, new_n880_, new_n878_ );
and g744 ( new_n882_, new_n881_, new_n622_ );
and g745 ( new_n883_, new_n877_, new_n882_ );
and g746 ( new_n884_, new_n883_, new_n876_ );
and g747 ( new_n885_, new_n884_, new_n528_ );
and g748 ( new_n886_, new_n734_, keyIn_0_28 );
not g749 ( new_n887_, keyIn_0_28 );
and g750 ( new_n888_, new_n622_, new_n887_ );
or g751 ( new_n889_, new_n886_, new_n888_ );
and g752 ( new_n890_, new_n889_, new_n814_ );
and g753 ( new_n891_, new_n692_, new_n890_ );
or g754 ( new_n892_, new_n885_, new_n891_ );
or g755 ( new_n893_, new_n873_, new_n892_ );
or g756 ( new_n894_, new_n893_, new_n863_ );
or g757 ( new_n895_, new_n894_, new_n859_ );
and g758 ( new_n896_, new_n895_, keyIn_0_38 );
not g759 ( new_n897_, keyIn_0_38 );
not g760 ( new_n898_, new_n859_ );
or g761 ( new_n899_, new_n858_, new_n852_ );
or g762 ( new_n900_, new_n528_, new_n865_ );
or g763 ( new_n901_, new_n692_, keyIn_0_32 );
and g764 ( new_n902_, new_n900_, new_n901_ );
not g765 ( new_n903_, new_n872_ );
or g766 ( new_n904_, new_n902_, new_n903_ );
not g767 ( new_n905_, new_n892_ );
and g768 ( new_n906_, new_n905_, new_n904_ );
and g769 ( new_n907_, new_n906_, new_n899_ );
and g770 ( new_n908_, new_n907_, new_n898_ );
and g771 ( new_n909_, new_n908_, new_n897_ );
or g772 ( new_n910_, new_n896_, new_n909_ );
and g773 ( new_n911_, new_n360_, new_n679_ );
and g774 ( new_n912_, new_n310_, new_n911_ );
not g775 ( new_n913_, new_n912_ );
or g776 ( new_n914_, new_n910_, new_n913_ );
or g777 ( new_n915_, new_n914_, keyIn_0_40 );
not g778 ( new_n916_, keyIn_0_40 );
or g779 ( new_n917_, new_n908_, new_n897_ );
or g780 ( new_n918_, new_n895_, keyIn_0_38 );
and g781 ( new_n919_, new_n918_, new_n917_ );
and g782 ( new_n920_, new_n919_, new_n912_ );
or g783 ( new_n921_, new_n920_, new_n916_ );
and g784 ( new_n922_, new_n915_, new_n921_ );
or g785 ( new_n923_, new_n922_, new_n737_ );
and g786 ( new_n924_, new_n923_, keyIn_0_47 );
not g787 ( new_n925_, keyIn_0_47 );
and g788 ( new_n926_, new_n920_, new_n916_ );
and g789 ( new_n927_, new_n914_, keyIn_0_40 );
or g790 ( new_n928_, new_n927_, new_n926_ );
and g791 ( new_n929_, new_n928_, new_n656_ );
and g792 ( new_n930_, new_n929_, new_n925_ );
or g793 ( new_n931_, new_n924_, new_n930_ );
and g794 ( new_n932_, new_n931_, new_n153_ );
or g795 ( new_n933_, new_n929_, new_n925_ );
or g796 ( new_n934_, new_n923_, keyIn_0_47 );
and g797 ( new_n935_, new_n934_, new_n933_ );
and g798 ( new_n936_, new_n935_, N65 );
or g799 ( N740, new_n932_, new_n936_ );
or g800 ( new_n938_, new_n922_, new_n622_ );
and g801 ( new_n939_, new_n938_, keyIn_0_48 );
not g802 ( new_n940_, keyIn_0_48 );
and g803 ( new_n941_, new_n928_, new_n734_ );
and g804 ( new_n942_, new_n941_, new_n940_ );
or g805 ( new_n943_, new_n939_, new_n942_ );
and g806 ( new_n944_, new_n943_, new_n151_ );
or g807 ( new_n945_, new_n941_, new_n940_ );
or g808 ( new_n946_, new_n938_, keyIn_0_48 );
and g809 ( new_n947_, new_n946_, new_n945_ );
and g810 ( new_n948_, new_n947_, N69 );
or g811 ( N741, new_n944_, new_n948_ );
and g812 ( new_n950_, new_n928_, new_n528_ );
not g813 ( new_n951_, new_n950_ );
and g814 ( new_n952_, new_n951_, N73 );
and g815 ( new_n953_, new_n950_, new_n142_ );
or g816 ( N742, new_n952_, new_n953_ );
not g817 ( new_n955_, keyIn_0_60 );
or g818 ( new_n956_, new_n922_, new_n597_ );
and g819 ( new_n957_, new_n956_, N77 );
and g820 ( new_n958_, new_n928_, new_n695_ );
and g821 ( new_n959_, new_n958_, new_n140_ );
or g822 ( new_n960_, new_n957_, new_n959_ );
or g823 ( new_n961_, new_n960_, new_n955_ );
or g824 ( new_n962_, new_n958_, new_n140_ );
or g825 ( new_n963_, new_n956_, N77 );
and g826 ( new_n964_, new_n963_, new_n962_ );
or g827 ( new_n965_, new_n964_, keyIn_0_60 );
and g828 ( N743, new_n961_, new_n965_ );
not g829 ( new_n967_, keyIn_0_34 );
and g830 ( new_n968_, new_n406_, new_n967_ );
and g831 ( new_n969_, new_n309_, keyIn_0_34 );
or g832 ( new_n970_, new_n968_, new_n969_ );
and g833 ( new_n971_, new_n393_, new_n209_ );
and g834 ( new_n972_, new_n420_, new_n971_ );
and g835 ( new_n973_, new_n970_, new_n972_ );
and g836 ( new_n974_, new_n919_, new_n973_ );
and g837 ( new_n975_, new_n974_, new_n656_ );
not g838 ( new_n976_, new_n975_ );
and g839 ( new_n977_, new_n976_, N81 );
and g840 ( new_n978_, new_n975_, new_n167_ );
or g841 ( N744, new_n977_, new_n978_ );
not g842 ( new_n980_, keyIn_0_49 );
and g843 ( new_n981_, new_n974_, new_n734_ );
and g844 ( new_n982_, new_n981_, new_n980_ );
not g845 ( new_n983_, new_n982_ );
or g846 ( new_n984_, new_n981_, new_n980_ );
and g847 ( new_n985_, new_n983_, new_n984_ );
not g848 ( new_n986_, new_n985_ );
and g849 ( new_n987_, new_n986_, N85 );
and g850 ( new_n988_, new_n985_, new_n165_ );
or g851 ( N745, new_n987_, new_n988_ );
and g852 ( new_n990_, new_n974_, new_n528_ );
and g853 ( new_n991_, new_n990_, new_n173_ );
not g854 ( new_n992_, new_n991_ );
or g855 ( new_n993_, new_n990_, new_n173_ );
and g856 ( new_n994_, new_n992_, new_n993_ );
not g857 ( new_n995_, new_n994_ );
and g858 ( new_n996_, new_n995_, keyIn_0_61 );
not g859 ( new_n997_, keyIn_0_61 );
and g860 ( new_n998_, new_n994_, new_n997_ );
or g861 ( N746, new_n996_, new_n998_ );
and g862 ( new_n1000_, new_n974_, new_n695_ );
not g863 ( new_n1001_, new_n1000_ );
and g864 ( new_n1002_, new_n1001_, N93 );
and g865 ( new_n1003_, new_n1000_, new_n171_ );
or g866 ( N747, new_n1002_, new_n1003_ );
and g867 ( new_n1005_, new_n208_, keyIn_0_35 );
not g868 ( new_n1006_, new_n1005_ );
or g869 ( new_n1007_, new_n208_, keyIn_0_35 );
and g870 ( new_n1008_, new_n1006_, new_n1007_ );
and g871 ( new_n1009_, new_n406_, new_n1008_ );
and g872 ( new_n1010_, new_n1009_, new_n911_ );
and g873 ( new_n1011_, new_n919_, new_n1010_ );
and g874 ( new_n1012_, new_n1011_, new_n656_ );
not g875 ( new_n1013_, new_n1012_ );
and g876 ( new_n1014_, new_n1013_, N97 );
and g877 ( new_n1015_, new_n1012_, new_n244_ );
or g878 ( N748, new_n1014_, new_n1015_ );
and g879 ( new_n1017_, new_n1011_, new_n734_ );
and g880 ( new_n1018_, new_n1017_, keyIn_0_50 );
not g881 ( new_n1019_, new_n1018_ );
or g882 ( new_n1020_, new_n1017_, keyIn_0_50 );
and g883 ( new_n1021_, new_n1019_, new_n1020_ );
not g884 ( new_n1022_, new_n1021_ );
and g885 ( new_n1023_, new_n1022_, new_n242_ );
and g886 ( new_n1024_, new_n1021_, N101 );
or g887 ( N749, new_n1023_, new_n1024_ );
and g888 ( new_n1026_, new_n1011_, new_n528_ );
not g889 ( new_n1027_, new_n1026_ );
and g890 ( new_n1028_, new_n1027_, N105 );
and g891 ( new_n1029_, new_n1026_, new_n238_ );
or g892 ( N750, new_n1028_, new_n1029_ );
and g893 ( new_n1031_, new_n1011_, new_n695_ );
not g894 ( new_n1032_, new_n1031_ );
and g895 ( new_n1033_, new_n1032_, N109 );
and g896 ( new_n1034_, new_n1031_, new_n236_ );
or g897 ( N751, new_n1033_, new_n1034_ );
and g898 ( new_n1036_, new_n408_, new_n420_ );
and g899 ( new_n1037_, new_n919_, new_n1036_ );
and g900 ( new_n1038_, new_n1037_, new_n656_ );
not g901 ( new_n1039_, new_n1038_ );
and g902 ( new_n1040_, new_n1039_, N113 );
and g903 ( new_n1041_, new_n1038_, new_n222_ );
or g904 ( N752, new_n1040_, new_n1041_ );
and g905 ( new_n1043_, new_n1037_, new_n734_ );
and g906 ( new_n1044_, new_n1043_, keyIn_0_51 );
not g907 ( new_n1045_, new_n1044_ );
or g908 ( new_n1046_, new_n1043_, keyIn_0_51 );
and g909 ( new_n1047_, new_n1045_, new_n1046_ );
not g910 ( new_n1048_, new_n1047_ );
and g911 ( new_n1049_, new_n1048_, N117 );
and g912 ( new_n1050_, new_n1047_, new_n220_ );
or g913 ( N753, new_n1049_, new_n1050_ );
not g914 ( new_n1052_, keyIn_0_62 );
not g915 ( new_n1053_, keyIn_0_52 );
not g916 ( new_n1054_, new_n1036_ );
or g917 ( new_n1055_, new_n910_, new_n1054_ );
or g918 ( new_n1056_, new_n1055_, new_n692_ );
and g919 ( new_n1057_, new_n1056_, new_n1053_ );
and g920 ( new_n1058_, new_n1037_, new_n528_ );
and g921 ( new_n1059_, new_n1058_, keyIn_0_52 );
or g922 ( new_n1060_, new_n1057_, new_n1059_ );
and g923 ( new_n1061_, new_n1060_, N121 );
or g924 ( new_n1062_, new_n1058_, keyIn_0_52 );
or g925 ( new_n1063_, new_n1056_, new_n1053_ );
and g926 ( new_n1064_, new_n1063_, new_n1062_ );
and g927 ( new_n1065_, new_n1064_, new_n213_ );
or g928 ( new_n1066_, new_n1061_, new_n1065_ );
and g929 ( new_n1067_, new_n1066_, new_n1052_ );
or g930 ( new_n1068_, new_n1064_, new_n213_ );
or g931 ( new_n1069_, new_n1060_, N121 );
and g932 ( new_n1070_, new_n1068_, new_n1069_ );
and g933 ( new_n1071_, new_n1070_, keyIn_0_62 );
or g934 ( N754, new_n1067_, new_n1071_ );
or g935 ( new_n1073_, new_n1055_, new_n597_ );
and g936 ( new_n1074_, new_n1073_, keyIn_0_53 );
not g937 ( new_n1075_, keyIn_0_53 );
and g938 ( new_n1076_, new_n1037_, new_n695_ );
and g939 ( new_n1077_, new_n1076_, new_n1075_ );
or g940 ( new_n1078_, new_n1074_, new_n1077_ );
and g941 ( new_n1079_, new_n1078_, N125 );
or g942 ( new_n1080_, new_n1076_, new_n1075_ );
or g943 ( new_n1081_, new_n1073_, keyIn_0_53 );
and g944 ( new_n1082_, new_n1081_, new_n1080_ );
and g945 ( new_n1083_, new_n1082_, new_n211_ );
or g946 ( new_n1084_, new_n1079_, new_n1083_ );
or g947 ( new_n1085_, new_n1084_, keyIn_0_63 );
not g948 ( new_n1086_, keyIn_0_63 );
or g949 ( new_n1087_, new_n1082_, new_n211_ );
or g950 ( new_n1088_, new_n1078_, N125 );
and g951 ( new_n1089_, new_n1087_, new_n1088_ );
or g952 ( new_n1090_, new_n1089_, new_n1086_ );
and g953 ( N755, new_n1085_, new_n1090_ );
endmodule