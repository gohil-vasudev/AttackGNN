module add_mul_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, 
        a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, 
        a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, 
        b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, 
        b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, 
        b_28_, b_29_, b_30_, b_31_, operation, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984;

  OR2_X1 U7472 ( .A1(n7948), .A2(n7450), .ZN(n7408) );
  INV_X1 U7473 ( .A(n7408), .ZN(n7409) );
  INV_X4 U7474 ( .A(operation), .ZN(n7410) );
  INV_X2 U7475 ( .A(b_0_), .ZN(n14788) );
  INV_X2 U7476 ( .A(b_28_), .ZN(n7949) );
  INV_X2 U7477 ( .A(b_22_), .ZN(n9881) );
  INV_X2 U7478 ( .A(a_1_), .ZN(n7872) );
  INV_X2 U7479 ( .A(a_20_), .ZN(n7957) );
  INV_X2 U7480 ( .A(a_24_), .ZN(n7954) );
  INV_X2 U7481 ( .A(a_25_), .ZN(n7952) );
  INV_X2 U7482 ( .A(a_23_), .ZN(n7955) );
  INV_X2 U7483 ( .A(a_17_), .ZN(n7645) );
  INV_X2 U7484 ( .A(a_18_), .ZN(n7960) );
  INV_X2 U7485 ( .A(a_21_), .ZN(n7578) );
  NAND2_X2 U7486 ( .A1(a_30_), .A2(n7948), .ZN(n7445) );
  NAND2_X2 U7487 ( .A1(a_31_), .A2(n7450), .ZN(n7441) );
  INV_X2 U7488 ( .A(a_29_), .ZN(n7460) );
  NOR2_X1 U7489 ( .A1(n7410), .A2(n7411), .ZN(Result_9_) );
  XOR2_X1 U7490 ( .A(n7412), .B(n7413), .Z(n7411) );
  NAND2_X1 U7491 ( .A1(n7414), .A2(n7415), .ZN(n7413) );
  NOR2_X1 U7492 ( .A1(n7410), .A2(n7416), .ZN(Result_8_) );
  XOR2_X1 U7493 ( .A(n7417), .B(n7418), .Z(n7416) );
  NAND2_X1 U7494 ( .A1(n7419), .A2(n7420), .ZN(n7418) );
  NOR2_X1 U7495 ( .A1(n7410), .A2(n7421), .ZN(Result_7_) );
  XOR2_X1 U7496 ( .A(n7422), .B(n7423), .Z(n7421) );
  NAND2_X1 U7497 ( .A1(n7424), .A2(n7425), .ZN(n7423) );
  NOR2_X1 U7498 ( .A1(n7410), .A2(n7426), .ZN(Result_6_) );
  XOR2_X1 U7499 ( .A(n7427), .B(n7428), .Z(n7426) );
  NAND2_X1 U7500 ( .A1(n7429), .A2(n7430), .ZN(n7428) );
  NAND2_X1 U7501 ( .A1(n7431), .A2(n7432), .ZN(Result_63_) );
  NAND2_X1 U7502 ( .A1(n7433), .A2(n7410), .ZN(n7432) );
  XOR2_X1 U7503 ( .A(b_31_), .B(a_31_), .Z(n7433) );
  NAND2_X1 U7504 ( .A1(n7434), .A2(operation), .ZN(n7431) );
  NAND2_X1 U7505 ( .A1(n7435), .A2(n7436), .ZN(Result_62_) );
  NAND2_X1 U7506 ( .A1(operation), .A2(n7437), .ZN(n7436) );
  NAND2_X1 U7507 ( .A1(n7438), .A2(n7439), .ZN(n7437) );
  NAND2_X1 U7508 ( .A1(b_30_), .A2(n7440), .ZN(n7439) );
  NAND2_X1 U7509 ( .A1(n7441), .A2(n7442), .ZN(n7440) );
  NAND2_X1 U7510 ( .A1(a_31_), .A2(n7443), .ZN(n7442) );
  NAND2_X1 U7511 ( .A1(b_31_), .A2(n7444), .ZN(n7438) );
  NAND2_X1 U7512 ( .A1(n7445), .A2(n7446), .ZN(n7444) );
  NAND2_X1 U7513 ( .A1(a_30_), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U7514 ( .A1(n7448), .A2(n7410), .ZN(n7435) );
  XNOR2_X1 U7515 ( .A(n7434), .B(n7449), .ZN(n7448) );
  XOR2_X1 U7516 ( .A(n7450), .B(b_30_), .Z(n7449) );
  NAND2_X1 U7517 ( .A1(n7451), .A2(n7452), .ZN(Result_61_) );
  NAND2_X1 U7518 ( .A1(n7453), .A2(n7410), .ZN(n7452) );
  NAND3_X1 U7519 ( .A1(n7454), .A2(n7455), .A3(n7456), .ZN(n7453) );
  NAND2_X1 U7520 ( .A1(n7457), .A2(n7458), .ZN(n7456) );
  NAND3_X1 U7521 ( .A1(n7459), .A2(n7460), .A3(b_29_), .ZN(n7455) );
  NAND2_X1 U7522 ( .A1(n7461), .A2(n7462), .ZN(n7454) );
  XOR2_X1 U7523 ( .A(n7460), .B(n7459), .Z(n7461) );
  INV_X1 U7524 ( .A(n7458), .ZN(n7459) );
  NAND2_X1 U7525 ( .A1(n7463), .A2(operation), .ZN(n7451) );
  XOR2_X1 U7526 ( .A(n7464), .B(n7465), .Z(n7463) );
  NOR2_X1 U7527 ( .A1(n7460), .A2(n7443), .ZN(n7465) );
  XOR2_X1 U7528 ( .A(n7466), .B(n7467), .Z(n7464) );
  NAND2_X1 U7529 ( .A1(n7468), .A2(n7469), .ZN(Result_60_) );
  NAND2_X1 U7530 ( .A1(n7470), .A2(n7410), .ZN(n7469) );
  XNOR2_X1 U7531 ( .A(n7471), .B(n7472), .ZN(n7470) );
  NAND2_X1 U7532 ( .A1(n7473), .A2(n7474), .ZN(n7471) );
  NAND2_X1 U7533 ( .A1(n7475), .A2(operation), .ZN(n7468) );
  XOR2_X1 U7534 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR2_X1 U7535 ( .A(n7478), .B(n7479), .Z(n7477) );
  NOR2_X1 U7536 ( .A1(n7480), .A2(n7443), .ZN(n7479) );
  NOR2_X1 U7537 ( .A1(n7410), .A2(n7481), .ZN(Result_5_) );
  XOR2_X1 U7538 ( .A(n7482), .B(n7483), .Z(n7481) );
  NAND2_X1 U7539 ( .A1(n7484), .A2(n7485), .ZN(n7483) );
  NAND2_X1 U7540 ( .A1(n7486), .A2(n7487), .ZN(Result_59_) );
  NAND2_X1 U7541 ( .A1(n7488), .A2(n7410), .ZN(n7487) );
  NAND3_X1 U7542 ( .A1(n7489), .A2(n7490), .A3(n7491), .ZN(n7488) );
  NAND2_X1 U7543 ( .A1(n7492), .A2(n7493), .ZN(n7491) );
  OR3_X1 U7544 ( .A1(n7493), .A2(a_27_), .A3(n7494), .ZN(n7490) );
  NAND2_X1 U7545 ( .A1(n7495), .A2(n7494), .ZN(n7489) );
  XOR2_X1 U7546 ( .A(n7493), .B(a_27_), .Z(n7495) );
  NAND2_X1 U7547 ( .A1(n7496), .A2(operation), .ZN(n7486) );
  XNOR2_X1 U7548 ( .A(n7497), .B(n7498), .ZN(n7496) );
  NAND2_X1 U7549 ( .A1(n7499), .A2(n7500), .ZN(n7497) );
  NAND2_X1 U7550 ( .A1(n7501), .A2(n7502), .ZN(Result_58_) );
  NAND2_X1 U7551 ( .A1(n7503), .A2(n7410), .ZN(n7502) );
  XOR2_X1 U7552 ( .A(n7504), .B(n7505), .Z(n7503) );
  AND2_X1 U7553 ( .A1(n7506), .A2(n7507), .ZN(n7505) );
  NAND2_X1 U7554 ( .A1(n7508), .A2(operation), .ZN(n7501) );
  XOR2_X1 U7555 ( .A(n7509), .B(n7510), .Z(n7508) );
  XOR2_X1 U7556 ( .A(n7511), .B(n7512), .Z(n7509) );
  NOR2_X1 U7557 ( .A1(n7513), .A2(n7443), .ZN(n7512) );
  NAND2_X1 U7558 ( .A1(n7514), .A2(n7515), .ZN(Result_57_) );
  NAND2_X1 U7559 ( .A1(n7516), .A2(n7410), .ZN(n7515) );
  NAND3_X1 U7560 ( .A1(n7517), .A2(n7518), .A3(n7519), .ZN(n7516) );
  NAND2_X1 U7561 ( .A1(n7520), .A2(n7521), .ZN(n7519) );
  OR3_X1 U7562 ( .A1(n7521), .A2(a_25_), .A3(n7522), .ZN(n7518) );
  NAND2_X1 U7563 ( .A1(n7523), .A2(n7522), .ZN(n7517) );
  XOR2_X1 U7564 ( .A(n7521), .B(a_25_), .Z(n7523) );
  NAND2_X1 U7565 ( .A1(n7524), .A2(operation), .ZN(n7514) );
  XNOR2_X1 U7566 ( .A(n7525), .B(n7526), .ZN(n7524) );
  NAND2_X1 U7567 ( .A1(n7527), .A2(n7528), .ZN(n7525) );
  NAND2_X1 U7568 ( .A1(n7529), .A2(n7530), .ZN(Result_56_) );
  NAND2_X1 U7569 ( .A1(n7531), .A2(n7410), .ZN(n7530) );
  XOR2_X1 U7570 ( .A(n7532), .B(n7533), .Z(n7531) );
  AND2_X1 U7571 ( .A1(n7534), .A2(n7535), .ZN(n7533) );
  NAND2_X1 U7572 ( .A1(n7536), .A2(operation), .ZN(n7529) );
  XOR2_X1 U7573 ( .A(n7537), .B(n7538), .Z(n7536) );
  XNOR2_X1 U7574 ( .A(n7539), .B(n7540), .ZN(n7538) );
  NAND2_X1 U7575 ( .A1(b_31_), .A2(a_24_), .ZN(n7539) );
  NAND2_X1 U7576 ( .A1(n7541), .A2(n7542), .ZN(Result_55_) );
  NAND2_X1 U7577 ( .A1(n7543), .A2(n7410), .ZN(n7542) );
  NAND3_X1 U7578 ( .A1(n7544), .A2(n7545), .A3(n7546), .ZN(n7543) );
  NAND2_X1 U7579 ( .A1(n7547), .A2(n7548), .ZN(n7546) );
  OR3_X1 U7580 ( .A1(n7548), .A2(a_23_), .A3(n7549), .ZN(n7545) );
  NAND2_X1 U7581 ( .A1(n7550), .A2(n7549), .ZN(n7544) );
  XOR2_X1 U7582 ( .A(n7548), .B(a_23_), .Z(n7550) );
  NAND2_X1 U7583 ( .A1(n7551), .A2(operation), .ZN(n7541) );
  XNOR2_X1 U7584 ( .A(n7552), .B(n7553), .ZN(n7551) );
  NAND2_X1 U7585 ( .A1(n7554), .A2(n7555), .ZN(n7552) );
  NAND2_X1 U7586 ( .A1(n7556), .A2(n7557), .ZN(Result_54_) );
  NAND2_X1 U7587 ( .A1(n7558), .A2(n7410), .ZN(n7557) );
  XNOR2_X1 U7588 ( .A(n7559), .B(n7560), .ZN(n7558) );
  NOR2_X1 U7589 ( .A1(n7561), .A2(n7562), .ZN(n7560) );
  NAND2_X1 U7590 ( .A1(n7563), .A2(operation), .ZN(n7556) );
  XOR2_X1 U7591 ( .A(n7564), .B(n7565), .Z(n7563) );
  XOR2_X1 U7592 ( .A(n7566), .B(n7567), .Z(n7565) );
  NOR2_X1 U7593 ( .A1(n7568), .A2(n7443), .ZN(n7567) );
  NAND2_X1 U7594 ( .A1(n7569), .A2(n7570), .ZN(Result_53_) );
  NAND2_X1 U7595 ( .A1(n7571), .A2(n7410), .ZN(n7570) );
  NAND3_X1 U7596 ( .A1(n7572), .A2(n7573), .A3(n7574), .ZN(n7571) );
  NAND2_X1 U7597 ( .A1(n7575), .A2(n7576), .ZN(n7574) );
  NAND3_X1 U7598 ( .A1(n7577), .A2(n7578), .A3(b_21_), .ZN(n7573) );
  NAND2_X1 U7599 ( .A1(n7579), .A2(n7580), .ZN(n7572) );
  XOR2_X1 U7600 ( .A(n7576), .B(a_21_), .Z(n7579) );
  NAND2_X1 U7601 ( .A1(n7581), .A2(operation), .ZN(n7569) );
  XOR2_X1 U7602 ( .A(n7582), .B(n7583), .Z(n7581) );
  XNOR2_X1 U7603 ( .A(n7584), .B(n7585), .ZN(n7583) );
  NAND2_X1 U7604 ( .A1(b_31_), .A2(a_21_), .ZN(n7585) );
  NAND2_X1 U7605 ( .A1(n7586), .A2(n7587), .ZN(Result_52_) );
  NAND2_X1 U7606 ( .A1(n7588), .A2(n7410), .ZN(n7587) );
  XOR2_X1 U7607 ( .A(n7589), .B(n7590), .Z(n7588) );
  AND2_X1 U7608 ( .A1(n7591), .A2(n7592), .ZN(n7590) );
  NAND2_X1 U7609 ( .A1(n7593), .A2(operation), .ZN(n7586) );
  XOR2_X1 U7610 ( .A(n7594), .B(n7595), .Z(n7593) );
  XNOR2_X1 U7611 ( .A(n7596), .B(n7597), .ZN(n7595) );
  NAND2_X1 U7612 ( .A1(b_31_), .A2(a_20_), .ZN(n7597) );
  NAND2_X1 U7613 ( .A1(n7598), .A2(n7599), .ZN(Result_51_) );
  NAND2_X1 U7614 ( .A1(n7600), .A2(n7410), .ZN(n7599) );
  NAND3_X1 U7615 ( .A1(n7601), .A2(n7602), .A3(n7603), .ZN(n7600) );
  NAND2_X1 U7616 ( .A1(n7604), .A2(n7605), .ZN(n7603) );
  OR3_X1 U7617 ( .A1(n7605), .A2(a_19_), .A3(n7606), .ZN(n7602) );
  NAND2_X1 U7618 ( .A1(n7607), .A2(n7606), .ZN(n7601) );
  XOR2_X1 U7619 ( .A(n7605), .B(a_19_), .Z(n7607) );
  NAND2_X1 U7620 ( .A1(n7608), .A2(operation), .ZN(n7598) );
  XNOR2_X1 U7621 ( .A(n7609), .B(n7610), .ZN(n7608) );
  XOR2_X1 U7622 ( .A(n7611), .B(n7612), .Z(n7610) );
  NAND2_X1 U7623 ( .A1(b_31_), .A2(a_19_), .ZN(n7612) );
  NAND2_X1 U7624 ( .A1(n7613), .A2(n7614), .ZN(Result_50_) );
  NAND2_X1 U7625 ( .A1(n7615), .A2(n7410), .ZN(n7614) );
  XOR2_X1 U7626 ( .A(n7616), .B(n7617), .Z(n7615) );
  AND2_X1 U7627 ( .A1(n7618), .A2(n7619), .ZN(n7617) );
  NAND2_X1 U7628 ( .A1(n7620), .A2(operation), .ZN(n7613) );
  XOR2_X1 U7629 ( .A(n7621), .B(n7622), .Z(n7620) );
  XNOR2_X1 U7630 ( .A(n7623), .B(n7624), .ZN(n7622) );
  NAND2_X1 U7631 ( .A1(b_31_), .A2(a_18_), .ZN(n7624) );
  NOR2_X1 U7632 ( .A1(n7410), .A2(n7625), .ZN(Result_4_) );
  XOR2_X1 U7633 ( .A(n7626), .B(n7627), .Z(n7625) );
  NAND2_X1 U7634 ( .A1(n7628), .A2(n7629), .ZN(n7627) );
  NAND2_X1 U7635 ( .A1(n7630), .A2(n7631), .ZN(Result_49_) );
  NAND2_X1 U7636 ( .A1(n7632), .A2(n7410), .ZN(n7631) );
  NAND3_X1 U7637 ( .A1(n7633), .A2(n7634), .A3(n7635), .ZN(n7632) );
  NAND2_X1 U7638 ( .A1(n7636), .A2(n7637), .ZN(n7635) );
  OR3_X1 U7639 ( .A1(n7637), .A2(a_17_), .A3(n7638), .ZN(n7634) );
  NAND2_X1 U7640 ( .A1(n7639), .A2(n7638), .ZN(n7633) );
  XOR2_X1 U7641 ( .A(n7637), .B(a_17_), .Z(n7639) );
  NAND2_X1 U7642 ( .A1(n7640), .A2(operation), .ZN(n7630) );
  XOR2_X1 U7643 ( .A(n7641), .B(n7642), .Z(n7640) );
  XOR2_X1 U7644 ( .A(n7643), .B(n7644), .Z(n7641) );
  NOR2_X1 U7645 ( .A1(n7645), .A2(n7443), .ZN(n7644) );
  NAND2_X1 U7646 ( .A1(n7646), .A2(n7647), .ZN(Result_48_) );
  NAND2_X1 U7647 ( .A1(n7648), .A2(n7410), .ZN(n7647) );
  XNOR2_X1 U7648 ( .A(n7649), .B(n7650), .ZN(n7648) );
  NOR2_X1 U7649 ( .A1(n7651), .A2(n7652), .ZN(n7650) );
  NAND2_X1 U7650 ( .A1(n7653), .A2(operation), .ZN(n7646) );
  XOR2_X1 U7651 ( .A(n7654), .B(n7655), .Z(n7653) );
  XNOR2_X1 U7652 ( .A(n7656), .B(n7657), .ZN(n7655) );
  NAND2_X1 U7653 ( .A1(b_31_), .A2(a_16_), .ZN(n7657) );
  NAND2_X1 U7654 ( .A1(n7658), .A2(n7659), .ZN(Result_47_) );
  NAND2_X1 U7655 ( .A1(n7660), .A2(n7410), .ZN(n7659) );
  NAND3_X1 U7656 ( .A1(n7661), .A2(n7662), .A3(n7663), .ZN(n7660) );
  NAND2_X1 U7657 ( .A1(n7664), .A2(n7665), .ZN(n7663) );
  NAND3_X1 U7658 ( .A1(n7666), .A2(n7667), .A3(b_15_), .ZN(n7662) );
  NAND2_X1 U7659 ( .A1(n7668), .A2(n7669), .ZN(n7661) );
  XOR2_X1 U7660 ( .A(n7665), .B(a_15_), .Z(n7668) );
  NAND2_X1 U7661 ( .A1(n7670), .A2(operation), .ZN(n7658) );
  XOR2_X1 U7662 ( .A(n7671), .B(n7672), .Z(n7670) );
  XOR2_X1 U7663 ( .A(n7673), .B(n7674), .Z(n7671) );
  NOR2_X1 U7664 ( .A1(n7667), .A2(n7443), .ZN(n7674) );
  NAND2_X1 U7665 ( .A1(n7675), .A2(n7676), .ZN(Result_46_) );
  NAND2_X1 U7666 ( .A1(n7677), .A2(n7410), .ZN(n7676) );
  XOR2_X1 U7667 ( .A(n7678), .B(n7679), .Z(n7677) );
  AND2_X1 U7668 ( .A1(n7680), .A2(n7681), .ZN(n7679) );
  NAND2_X1 U7669 ( .A1(n7682), .A2(operation), .ZN(n7675) );
  XOR2_X1 U7670 ( .A(n7683), .B(n7684), .Z(n7682) );
  XNOR2_X1 U7671 ( .A(n7685), .B(n7686), .ZN(n7684) );
  NAND2_X1 U7672 ( .A1(b_31_), .A2(a_14_), .ZN(n7686) );
  NAND2_X1 U7673 ( .A1(n7687), .A2(n7688), .ZN(Result_45_) );
  NAND2_X1 U7674 ( .A1(n7689), .A2(n7410), .ZN(n7688) );
  NAND3_X1 U7675 ( .A1(n7690), .A2(n7691), .A3(n7692), .ZN(n7689) );
  NAND2_X1 U7676 ( .A1(n7693), .A2(n7694), .ZN(n7692) );
  OR3_X1 U7677 ( .A1(n7694), .A2(a_13_), .A3(n7695), .ZN(n7691) );
  NAND2_X1 U7678 ( .A1(n7696), .A2(n7695), .ZN(n7690) );
  XOR2_X1 U7679 ( .A(n7694), .B(a_13_), .Z(n7696) );
  NAND2_X1 U7680 ( .A1(n7697), .A2(operation), .ZN(n7687) );
  XOR2_X1 U7681 ( .A(n7698), .B(n7699), .Z(n7697) );
  XOR2_X1 U7682 ( .A(n7700), .B(n7701), .Z(n7698) );
  NOR2_X1 U7683 ( .A1(n7702), .A2(n7443), .ZN(n7701) );
  NAND2_X1 U7684 ( .A1(n7703), .A2(n7704), .ZN(Result_44_) );
  NAND2_X1 U7685 ( .A1(n7705), .A2(n7410), .ZN(n7704) );
  XNOR2_X1 U7686 ( .A(n7706), .B(n7707), .ZN(n7705) );
  NOR2_X1 U7687 ( .A1(n7708), .A2(n7709), .ZN(n7707) );
  NAND2_X1 U7688 ( .A1(n7710), .A2(operation), .ZN(n7703) );
  XOR2_X1 U7689 ( .A(n7711), .B(n7712), .Z(n7710) );
  XNOR2_X1 U7690 ( .A(n7713), .B(n7714), .ZN(n7712) );
  NAND2_X1 U7691 ( .A1(b_31_), .A2(a_12_), .ZN(n7714) );
  NAND2_X1 U7692 ( .A1(n7715), .A2(n7716), .ZN(Result_43_) );
  NAND2_X1 U7693 ( .A1(n7717), .A2(n7410), .ZN(n7716) );
  NAND3_X1 U7694 ( .A1(n7718), .A2(n7719), .A3(n7720), .ZN(n7717) );
  NAND2_X1 U7695 ( .A1(n7721), .A2(n7722), .ZN(n7720) );
  NAND3_X1 U7696 ( .A1(n7723), .A2(n7724), .A3(b_11_), .ZN(n7719) );
  NAND2_X1 U7697 ( .A1(n7725), .A2(n7726), .ZN(n7718) );
  XOR2_X1 U7698 ( .A(n7722), .B(a_11_), .Z(n7725) );
  NAND2_X1 U7699 ( .A1(n7727), .A2(operation), .ZN(n7715) );
  XNOR2_X1 U7700 ( .A(n7728), .B(n7729), .ZN(n7727) );
  XOR2_X1 U7701 ( .A(n7730), .B(n7731), .Z(n7729) );
  NAND2_X1 U7702 ( .A1(b_31_), .A2(a_11_), .ZN(n7731) );
  NAND2_X1 U7703 ( .A1(n7732), .A2(n7733), .ZN(Result_42_) );
  NAND2_X1 U7704 ( .A1(n7734), .A2(n7410), .ZN(n7733) );
  XNOR2_X1 U7705 ( .A(n7735), .B(n7736), .ZN(n7734) );
  NOR2_X1 U7706 ( .A1(n7737), .A2(n7738), .ZN(n7736) );
  NAND2_X1 U7707 ( .A1(n7739), .A2(operation), .ZN(n7732) );
  XOR2_X1 U7708 ( .A(n7740), .B(n7741), .Z(n7739) );
  XNOR2_X1 U7709 ( .A(n7742), .B(n7743), .ZN(n7741) );
  NAND2_X1 U7710 ( .A1(b_31_), .A2(a_10_), .ZN(n7743) );
  NAND2_X1 U7711 ( .A1(n7744), .A2(n7745), .ZN(Result_41_) );
  NAND2_X1 U7712 ( .A1(n7746), .A2(n7410), .ZN(n7745) );
  NAND3_X1 U7713 ( .A1(n7747), .A2(n7748), .A3(n7749), .ZN(n7746) );
  NAND2_X1 U7714 ( .A1(n7750), .A2(n7751), .ZN(n7749) );
  NAND3_X1 U7715 ( .A1(n7752), .A2(n7753), .A3(b_9_), .ZN(n7748) );
  NAND2_X1 U7716 ( .A1(n7754), .A2(n7755), .ZN(n7747) );
  XOR2_X1 U7717 ( .A(n7751), .B(a_9_), .Z(n7754) );
  NAND2_X1 U7718 ( .A1(n7756), .A2(operation), .ZN(n7744) );
  XOR2_X1 U7719 ( .A(n7757), .B(n7758), .Z(n7756) );
  XNOR2_X1 U7720 ( .A(n7759), .B(n7760), .ZN(n7758) );
  NAND2_X1 U7721 ( .A1(b_31_), .A2(a_9_), .ZN(n7760) );
  NAND2_X1 U7722 ( .A1(n7761), .A2(n7762), .ZN(Result_40_) );
  NAND2_X1 U7723 ( .A1(n7763), .A2(n7410), .ZN(n7762) );
  XNOR2_X1 U7724 ( .A(n7764), .B(n7765), .ZN(n7763) );
  NOR2_X1 U7725 ( .A1(n7766), .A2(n7767), .ZN(n7765) );
  NAND2_X1 U7726 ( .A1(n7768), .A2(operation), .ZN(n7761) );
  XOR2_X1 U7727 ( .A(n7769), .B(n7770), .Z(n7768) );
  XNOR2_X1 U7728 ( .A(n7771), .B(n7772), .ZN(n7770) );
  NAND2_X1 U7729 ( .A1(b_31_), .A2(a_8_), .ZN(n7772) );
  NOR2_X1 U7730 ( .A1(n7410), .A2(n7773), .ZN(Result_3_) );
  XOR2_X1 U7731 ( .A(n7774), .B(n7775), .Z(n7773) );
  NAND2_X1 U7732 ( .A1(n7776), .A2(n7777), .ZN(n7775) );
  NAND2_X1 U7733 ( .A1(n7778), .A2(n7779), .ZN(Result_39_) );
  NAND2_X1 U7734 ( .A1(n7780), .A2(n7410), .ZN(n7779) );
  NAND3_X1 U7735 ( .A1(n7781), .A2(n7782), .A3(n7783), .ZN(n7780) );
  NAND2_X1 U7736 ( .A1(n7784), .A2(n7785), .ZN(n7783) );
  NAND3_X1 U7737 ( .A1(n7786), .A2(n7787), .A3(b_7_), .ZN(n7782) );
  NAND2_X1 U7738 ( .A1(n7788), .A2(n7789), .ZN(n7781) );
  XOR2_X1 U7739 ( .A(n7785), .B(a_7_), .Z(n7788) );
  NAND2_X1 U7740 ( .A1(n7790), .A2(operation), .ZN(n7778) );
  XNOR2_X1 U7741 ( .A(n7791), .B(n7792), .ZN(n7790) );
  XOR2_X1 U7742 ( .A(n7793), .B(n7794), .Z(n7792) );
  NAND2_X1 U7743 ( .A1(b_31_), .A2(a_7_), .ZN(n7794) );
  NAND2_X1 U7744 ( .A1(n7795), .A2(n7796), .ZN(Result_38_) );
  NAND2_X1 U7745 ( .A1(n7797), .A2(n7410), .ZN(n7796) );
  XOR2_X1 U7746 ( .A(n7798), .B(n7799), .Z(n7797) );
  AND2_X1 U7747 ( .A1(n7800), .A2(n7801), .ZN(n7799) );
  NAND2_X1 U7748 ( .A1(n7802), .A2(operation), .ZN(n7795) );
  XOR2_X1 U7749 ( .A(n7803), .B(n7804), .Z(n7802) );
  XOR2_X1 U7750 ( .A(n7805), .B(n7806), .Z(n7803) );
  NOR2_X1 U7751 ( .A1(n7807), .A2(n7443), .ZN(n7806) );
  NAND2_X1 U7752 ( .A1(n7808), .A2(n7809), .ZN(Result_37_) );
  NAND2_X1 U7753 ( .A1(n7810), .A2(n7410), .ZN(n7809) );
  NAND3_X1 U7754 ( .A1(n7811), .A2(n7812), .A3(n7813), .ZN(n7810) );
  NAND2_X1 U7755 ( .A1(n7814), .A2(n7815), .ZN(n7813) );
  OR3_X1 U7756 ( .A1(n7815), .A2(a_5_), .A3(n7816), .ZN(n7812) );
  NAND2_X1 U7757 ( .A1(n7817), .A2(n7816), .ZN(n7811) );
  XOR2_X1 U7758 ( .A(n7815), .B(a_5_), .Z(n7817) );
  NAND2_X1 U7759 ( .A1(n7818), .A2(operation), .ZN(n7808) );
  XOR2_X1 U7760 ( .A(n7819), .B(n7820), .Z(n7818) );
  XOR2_X1 U7761 ( .A(n7821), .B(n7822), .Z(n7819) );
  NOR2_X1 U7762 ( .A1(n7823), .A2(n7443), .ZN(n7822) );
  NAND2_X1 U7763 ( .A1(n7824), .A2(n7825), .ZN(Result_36_) );
  NAND2_X1 U7764 ( .A1(n7826), .A2(n7410), .ZN(n7825) );
  XOR2_X1 U7765 ( .A(n7827), .B(n7828), .Z(n7826) );
  AND2_X1 U7766 ( .A1(n7829), .A2(n7830), .ZN(n7828) );
  NAND2_X1 U7767 ( .A1(n7831), .A2(operation), .ZN(n7824) );
  XOR2_X1 U7768 ( .A(n7832), .B(n7833), .Z(n7831) );
  XOR2_X1 U7769 ( .A(n7834), .B(n7835), .Z(n7832) );
  NOR2_X1 U7770 ( .A1(n7836), .A2(n7443), .ZN(n7835) );
  NAND2_X1 U7771 ( .A1(n7837), .A2(n7838), .ZN(Result_35_) );
  NAND2_X1 U7772 ( .A1(n7839), .A2(n7410), .ZN(n7838) );
  NAND3_X1 U7773 ( .A1(n7840), .A2(n7841), .A3(n7842), .ZN(n7839) );
  NAND2_X1 U7774 ( .A1(n7843), .A2(n7844), .ZN(n7842) );
  OR3_X1 U7775 ( .A1(n7844), .A2(a_3_), .A3(n7845), .ZN(n7841) );
  NAND2_X1 U7776 ( .A1(n7846), .A2(n7845), .ZN(n7840) );
  XOR2_X1 U7777 ( .A(n7844), .B(a_3_), .Z(n7846) );
  NAND2_X1 U7778 ( .A1(n7847), .A2(operation), .ZN(n7837) );
  XOR2_X1 U7779 ( .A(n7848), .B(n7849), .Z(n7847) );
  XOR2_X1 U7780 ( .A(n7850), .B(n7851), .Z(n7848) );
  NOR2_X1 U7781 ( .A1(n7852), .A2(n7443), .ZN(n7851) );
  NAND2_X1 U7782 ( .A1(n7853), .A2(n7854), .ZN(Result_34_) );
  NAND2_X1 U7783 ( .A1(n7855), .A2(n7410), .ZN(n7854) );
  XOR2_X1 U7784 ( .A(n7856), .B(n7857), .Z(n7855) );
  AND2_X1 U7785 ( .A1(n7858), .A2(n7859), .ZN(n7857) );
  NAND2_X1 U7786 ( .A1(n7860), .A2(operation), .ZN(n7853) );
  XOR2_X1 U7787 ( .A(n7861), .B(n7862), .Z(n7860) );
  XNOR2_X1 U7788 ( .A(n7863), .B(n7864), .ZN(n7862) );
  NAND2_X1 U7789 ( .A1(b_31_), .A2(a_2_), .ZN(n7864) );
  NAND2_X1 U7790 ( .A1(n7865), .A2(n7866), .ZN(Result_33_) );
  NAND2_X1 U7791 ( .A1(n7867), .A2(operation), .ZN(n7866) );
  XOR2_X1 U7792 ( .A(n7868), .B(n7869), .Z(n7867) );
  XOR2_X1 U7793 ( .A(n7870), .B(n7871), .Z(n7868) );
  NOR2_X1 U7794 ( .A1(n7872), .A2(n7443), .ZN(n7871) );
  NAND2_X1 U7795 ( .A1(n7873), .A2(n7410), .ZN(n7865) );
  NAND2_X1 U7796 ( .A1(n7874), .A2(n7875), .ZN(n7873) );
  NAND2_X1 U7797 ( .A1(n7876), .A2(n7877), .ZN(n7875) );
  OR2_X1 U7798 ( .A1(n7878), .A2(n7879), .ZN(n7876) );
  NAND2_X1 U7799 ( .A1(n7880), .A2(n7881), .ZN(n7874) );
  INV_X1 U7800 ( .A(n7877), .ZN(n7881) );
  XOR2_X1 U7801 ( .A(b_1_), .B(a_1_), .Z(n7880) );
  NAND2_X1 U7802 ( .A1(n7882), .A2(n7883), .ZN(Result_32_) );
  NAND2_X1 U7803 ( .A1(n7884), .A2(n7410), .ZN(n7883) );
  XOR2_X1 U7804 ( .A(n7885), .B(n7886), .Z(n7884) );
  NOR2_X1 U7805 ( .A1(n7887), .A2(n7888), .ZN(n7886) );
  NOR2_X1 U7806 ( .A1(b_0_), .A2(a_0_), .ZN(n7887) );
  NOR2_X1 U7807 ( .A1(n7879), .A2(n7889), .ZN(n7885) );
  NOR2_X1 U7808 ( .A1(n7878), .A2(n7877), .ZN(n7889) );
  NAND2_X1 U7809 ( .A1(n7859), .A2(n7890), .ZN(n7877) );
  NAND2_X1 U7810 ( .A1(n7858), .A2(n7856), .ZN(n7890) );
  NAND2_X1 U7811 ( .A1(n7891), .A2(n7892), .ZN(n7856) );
  NAND2_X1 U7812 ( .A1(n7893), .A2(n7844), .ZN(n7892) );
  NAND2_X1 U7813 ( .A1(n7830), .A2(n7894), .ZN(n7844) );
  NAND2_X1 U7814 ( .A1(n7829), .A2(n7827), .ZN(n7894) );
  NAND2_X1 U7815 ( .A1(n7895), .A2(n7896), .ZN(n7827) );
  NAND2_X1 U7816 ( .A1(n7897), .A2(n7815), .ZN(n7896) );
  NAND2_X1 U7817 ( .A1(n7801), .A2(n7898), .ZN(n7815) );
  NAND2_X1 U7818 ( .A1(n7800), .A2(n7798), .ZN(n7898) );
  NAND2_X1 U7819 ( .A1(n7899), .A2(n7900), .ZN(n7798) );
  NAND2_X1 U7820 ( .A1(n7901), .A2(n7785), .ZN(n7900) );
  INV_X1 U7821 ( .A(n7786), .ZN(n7785) );
  NOR2_X1 U7822 ( .A1(n7767), .A2(n7902), .ZN(n7786) );
  NOR2_X1 U7823 ( .A1(n7766), .A2(n7764), .ZN(n7902) );
  AND2_X1 U7824 ( .A1(n7903), .A2(n7904), .ZN(n7764) );
  NAND2_X1 U7825 ( .A1(n7905), .A2(n7751), .ZN(n7904) );
  INV_X1 U7826 ( .A(n7752), .ZN(n7751) );
  NOR2_X1 U7827 ( .A1(n7738), .A2(n7906), .ZN(n7752) );
  NOR2_X1 U7828 ( .A1(n7737), .A2(n7735), .ZN(n7906) );
  AND2_X1 U7829 ( .A1(n7907), .A2(n7908), .ZN(n7735) );
  NAND2_X1 U7830 ( .A1(n7909), .A2(n7722), .ZN(n7908) );
  INV_X1 U7831 ( .A(n7723), .ZN(n7722) );
  NOR2_X1 U7832 ( .A1(n7709), .A2(n7910), .ZN(n7723) );
  NOR2_X1 U7833 ( .A1(n7708), .A2(n7706), .ZN(n7910) );
  AND2_X1 U7834 ( .A1(n7911), .A2(n7912), .ZN(n7706) );
  NAND2_X1 U7835 ( .A1(n7913), .A2(n7694), .ZN(n7912) );
  NAND2_X1 U7836 ( .A1(n7681), .A2(n7914), .ZN(n7694) );
  NAND2_X1 U7837 ( .A1(n7680), .A2(n7678), .ZN(n7914) );
  NAND2_X1 U7838 ( .A1(n7915), .A2(n7916), .ZN(n7678) );
  NAND2_X1 U7839 ( .A1(n7917), .A2(n7665), .ZN(n7916) );
  INV_X1 U7840 ( .A(n7666), .ZN(n7665) );
  NOR2_X1 U7841 ( .A1(n7652), .A2(n7918), .ZN(n7666) );
  NOR2_X1 U7842 ( .A1(n7651), .A2(n7649), .ZN(n7918) );
  AND2_X1 U7843 ( .A1(n7919), .A2(n7920), .ZN(n7649) );
  NAND2_X1 U7844 ( .A1(n7921), .A2(n7637), .ZN(n7920) );
  NAND2_X1 U7845 ( .A1(n7619), .A2(n7922), .ZN(n7637) );
  NAND2_X1 U7846 ( .A1(n7618), .A2(n7616), .ZN(n7922) );
  NAND2_X1 U7847 ( .A1(n7923), .A2(n7924), .ZN(n7616) );
  NAND2_X1 U7848 ( .A1(n7925), .A2(n7605), .ZN(n7924) );
  NAND2_X1 U7849 ( .A1(n7592), .A2(n7926), .ZN(n7605) );
  NAND2_X1 U7850 ( .A1(n7591), .A2(n7589), .ZN(n7926) );
  NAND2_X1 U7851 ( .A1(n7927), .A2(n7928), .ZN(n7589) );
  NAND2_X1 U7852 ( .A1(n7929), .A2(n7576), .ZN(n7928) );
  INV_X1 U7853 ( .A(n7577), .ZN(n7576) );
  NOR2_X1 U7854 ( .A1(n7562), .A2(n7930), .ZN(n7577) );
  NOR2_X1 U7855 ( .A1(n7561), .A2(n7559), .ZN(n7930) );
  NOR2_X1 U7856 ( .A1(n7547), .A2(n7931), .ZN(n7559) );
  AND2_X1 U7857 ( .A1(n7932), .A2(n7548), .ZN(n7931) );
  NAND2_X1 U7858 ( .A1(n7535), .A2(n7933), .ZN(n7548) );
  NAND2_X1 U7859 ( .A1(n7534), .A2(n7532), .ZN(n7933) );
  NAND2_X1 U7860 ( .A1(n7934), .A2(n7935), .ZN(n7532) );
  NAND2_X1 U7861 ( .A1(n7936), .A2(n7521), .ZN(n7935) );
  NAND2_X1 U7862 ( .A1(n7507), .A2(n7937), .ZN(n7521) );
  NAND2_X1 U7863 ( .A1(n7506), .A2(n7504), .ZN(n7937) );
  NAND2_X1 U7864 ( .A1(n7938), .A2(n7939), .ZN(n7504) );
  NAND2_X1 U7865 ( .A1(n7940), .A2(n7493), .ZN(n7939) );
  NAND2_X1 U7866 ( .A1(n7473), .A2(n7941), .ZN(n7493) );
  NAND2_X1 U7867 ( .A1(n7474), .A2(n7472), .ZN(n7941) );
  NAND2_X1 U7868 ( .A1(n7942), .A2(n7943), .ZN(n7472) );
  NAND2_X1 U7869 ( .A1(n7944), .A2(n7458), .ZN(n7943) );
  NAND2_X1 U7870 ( .A1(n7945), .A2(n7946), .ZN(n7458) );
  NAND2_X1 U7871 ( .A1(b_30_), .A2(n7947), .ZN(n7946) );
  OR2_X1 U7872 ( .A1(a_30_), .A2(n7434), .ZN(n7947) );
  NOR2_X1 U7873 ( .A1(n7443), .A2(n7948), .ZN(n7434) );
  INV_X1 U7874 ( .A(b_31_), .ZN(n7443) );
  NAND2_X1 U7875 ( .A1(b_31_), .A2(n7409), .ZN(n7945) );
  NAND2_X1 U7876 ( .A1(n7462), .A2(n7460), .ZN(n7944) );
  NAND2_X1 U7877 ( .A1(n7949), .A2(n7480), .ZN(n7474) );
  NAND2_X1 U7878 ( .A1(n7494), .A2(n7950), .ZN(n7940) );
  NAND2_X1 U7879 ( .A1(n7951), .A2(n7513), .ZN(n7506) );
  INV_X1 U7880 ( .A(a_26_), .ZN(n7513) );
  NAND2_X1 U7881 ( .A1(n7522), .A2(n7952), .ZN(n7936) );
  NAND2_X1 U7882 ( .A1(n7953), .A2(n7954), .ZN(n7534) );
  NAND2_X1 U7883 ( .A1(n7549), .A2(n7955), .ZN(n7932) );
  NOR2_X1 U7884 ( .A1(b_22_), .A2(a_22_), .ZN(n7561) );
  NAND2_X1 U7885 ( .A1(n7580), .A2(n7578), .ZN(n7929) );
  NAND2_X1 U7886 ( .A1(n7956), .A2(n7957), .ZN(n7591) );
  NAND2_X1 U7887 ( .A1(n7606), .A2(n7958), .ZN(n7925) );
  NAND2_X1 U7888 ( .A1(n7959), .A2(n7960), .ZN(n7618) );
  NAND2_X1 U7889 ( .A1(n7638), .A2(n7645), .ZN(n7921) );
  NOR2_X1 U7890 ( .A1(b_16_), .A2(a_16_), .ZN(n7651) );
  NAND2_X1 U7891 ( .A1(n7669), .A2(n7667), .ZN(n7917) );
  NAND2_X1 U7892 ( .A1(n7961), .A2(n7962), .ZN(n7680) );
  NAND2_X1 U7893 ( .A1(n7695), .A2(n7702), .ZN(n7913) );
  NOR2_X1 U7894 ( .A1(b_12_), .A2(a_12_), .ZN(n7708) );
  NAND2_X1 U7895 ( .A1(n7726), .A2(n7724), .ZN(n7909) );
  NOR2_X1 U7896 ( .A1(b_10_), .A2(a_10_), .ZN(n7737) );
  NAND2_X1 U7897 ( .A1(n7755), .A2(n7753), .ZN(n7905) );
  NOR2_X1 U7898 ( .A1(b_8_), .A2(a_8_), .ZN(n7766) );
  NAND2_X1 U7899 ( .A1(n7789), .A2(n7787), .ZN(n7901) );
  NAND2_X1 U7900 ( .A1(n7963), .A2(n7807), .ZN(n7800) );
  NAND2_X1 U7901 ( .A1(n7816), .A2(n7823), .ZN(n7897) );
  NAND2_X1 U7902 ( .A1(n7964), .A2(n7836), .ZN(n7829) );
  NAND2_X1 U7903 ( .A1(n7845), .A2(n7852), .ZN(n7893) );
  NAND2_X1 U7904 ( .A1(n7965), .A2(n7966), .ZN(n7858) );
  NOR2_X1 U7905 ( .A1(b_1_), .A2(a_1_), .ZN(n7879) );
  NAND2_X1 U7906 ( .A1(n7967), .A2(operation), .ZN(n7882) );
  XOR2_X1 U7907 ( .A(n7968), .B(n7969), .Z(n7967) );
  XNOR2_X1 U7908 ( .A(n7970), .B(n7971), .ZN(n7969) );
  NAND2_X1 U7909 ( .A1(b_31_), .A2(a_0_), .ZN(n7971) );
  NOR2_X1 U7910 ( .A1(n7972), .A2(n7410), .ZN(Result_31_) );
  XNOR2_X1 U7911 ( .A(n7973), .B(n7974), .ZN(n7972) );
  NOR3_X1 U7912 ( .A1(n7410), .A2(n7975), .A3(n7976), .ZN(Result_30_) );
  NOR2_X1 U7913 ( .A1(n7977), .A2(n7978), .ZN(n7976) );
  AND2_X1 U7914 ( .A1(n7974), .A2(n7973), .ZN(n7977) );
  NOR2_X1 U7915 ( .A1(n7410), .A2(n7979), .ZN(Result_2_) );
  XOR2_X1 U7916 ( .A(n7980), .B(n7981), .Z(n7979) );
  NAND2_X1 U7917 ( .A1(n7982), .A2(n7983), .ZN(n7981) );
  NOR2_X1 U7918 ( .A1(n7984), .A2(n7410), .ZN(Result_29_) );
  XNOR2_X1 U7919 ( .A(n7975), .B(n7985), .ZN(n7984) );
  AND2_X1 U7920 ( .A1(n7986), .A2(n7987), .ZN(n7985) );
  NOR2_X1 U7921 ( .A1(n7410), .A2(n7988), .ZN(Result_28_) );
  XOR2_X1 U7922 ( .A(n7989), .B(n7990), .Z(n7988) );
  NOR2_X1 U7923 ( .A1(n7991), .A2(n7992), .ZN(n7990) );
  NOR2_X1 U7924 ( .A1(n7410), .A2(n7993), .ZN(Result_27_) );
  XOR2_X1 U7925 ( .A(n7994), .B(n7995), .Z(n7993) );
  NOR2_X1 U7926 ( .A1(n7996), .A2(n7997), .ZN(n7995) );
  NOR2_X1 U7927 ( .A1(n7410), .A2(n7998), .ZN(Result_26_) );
  XOR2_X1 U7928 ( .A(n7999), .B(n8000), .Z(n7998) );
  NAND2_X1 U7929 ( .A1(n8001), .A2(n8002), .ZN(n7999) );
  NOR2_X1 U7930 ( .A1(n7410), .A2(n8003), .ZN(Result_25_) );
  XOR2_X1 U7931 ( .A(n8004), .B(n8005), .Z(n8003) );
  NAND2_X1 U7932 ( .A1(n8006), .A2(n8007), .ZN(n8005) );
  NOR2_X1 U7933 ( .A1(n7410), .A2(n8008), .ZN(Result_24_) );
  XOR2_X1 U7934 ( .A(n8009), .B(n8010), .Z(n8008) );
  NAND2_X1 U7935 ( .A1(n8011), .A2(n8012), .ZN(n8010) );
  NOR2_X1 U7936 ( .A1(n7410), .A2(n8013), .ZN(Result_23_) );
  XOR2_X1 U7937 ( .A(n8014), .B(n8015), .Z(n8013) );
  NAND2_X1 U7938 ( .A1(n8016), .A2(n8017), .ZN(n8015) );
  NOR2_X1 U7939 ( .A1(n7410), .A2(n8018), .ZN(Result_22_) );
  XOR2_X1 U7940 ( .A(n8019), .B(n8020), .Z(n8018) );
  NAND2_X1 U7941 ( .A1(n8021), .A2(n8022), .ZN(n8020) );
  NOR2_X1 U7942 ( .A1(n7410), .A2(n8023), .ZN(Result_21_) );
  XOR2_X1 U7943 ( .A(n8024), .B(n8025), .Z(n8023) );
  NAND2_X1 U7944 ( .A1(n8026), .A2(n8027), .ZN(n8025) );
  NOR2_X1 U7945 ( .A1(n7410), .A2(n8028), .ZN(Result_20_) );
  XOR2_X1 U7946 ( .A(n8029), .B(n8030), .Z(n8028) );
  NAND2_X1 U7947 ( .A1(n8031), .A2(n8032), .ZN(n8030) );
  NOR2_X1 U7948 ( .A1(n7410), .A2(n8033), .ZN(Result_1_) );
  XOR2_X1 U7949 ( .A(n8034), .B(n8035), .Z(n8033) );
  NAND2_X1 U7950 ( .A1(n8036), .A2(n8037), .ZN(n8035) );
  NOR2_X1 U7951 ( .A1(n7410), .A2(n8038), .ZN(Result_19_) );
  XOR2_X1 U7952 ( .A(n8039), .B(n8040), .Z(n8038) );
  NAND2_X1 U7953 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
  NOR2_X1 U7954 ( .A1(n7410), .A2(n8043), .ZN(Result_18_) );
  XOR2_X1 U7955 ( .A(n8044), .B(n8045), .Z(n8043) );
  NAND2_X1 U7956 ( .A1(n8046), .A2(n8047), .ZN(n8045) );
  NOR2_X1 U7957 ( .A1(n7410), .A2(n8048), .ZN(Result_17_) );
  XOR2_X1 U7958 ( .A(n8049), .B(n8050), .Z(n8048) );
  NAND2_X1 U7959 ( .A1(n8051), .A2(n8052), .ZN(n8050) );
  NOR2_X1 U7960 ( .A1(n7410), .A2(n8053), .ZN(Result_16_) );
  XOR2_X1 U7961 ( .A(n8054), .B(n8055), .Z(n8053) );
  NAND2_X1 U7962 ( .A1(n8056), .A2(n8057), .ZN(n8055) );
  NOR2_X1 U7963 ( .A1(n7410), .A2(n8058), .ZN(Result_15_) );
  XOR2_X1 U7964 ( .A(n8059), .B(n8060), .Z(n8058) );
  NAND2_X1 U7965 ( .A1(n8061), .A2(n8062), .ZN(n8060) );
  NOR2_X1 U7966 ( .A1(n7410), .A2(n8063), .ZN(Result_14_) );
  XOR2_X1 U7967 ( .A(n8064), .B(n8065), .Z(n8063) );
  NAND2_X1 U7968 ( .A1(n8066), .A2(n8067), .ZN(n8065) );
  NOR2_X1 U7969 ( .A1(n7410), .A2(n8068), .ZN(Result_13_) );
  XOR2_X1 U7970 ( .A(n8069), .B(n8070), .Z(n8068) );
  NAND2_X1 U7971 ( .A1(n8071), .A2(n8072), .ZN(n8070) );
  NOR2_X1 U7972 ( .A1(n7410), .A2(n8073), .ZN(Result_12_) );
  XOR2_X1 U7973 ( .A(n8074), .B(n8075), .Z(n8073) );
  NAND2_X1 U7974 ( .A1(n8076), .A2(n8077), .ZN(n8075) );
  NOR2_X1 U7975 ( .A1(n7410), .A2(n8078), .ZN(Result_11_) );
  XOR2_X1 U7976 ( .A(n8079), .B(n8080), .Z(n8078) );
  NAND2_X1 U7977 ( .A1(n8081), .A2(n8082), .ZN(n8080) );
  NOR2_X1 U7978 ( .A1(n7410), .A2(n8083), .ZN(Result_10_) );
  XOR2_X1 U7979 ( .A(n8084), .B(n8085), .Z(n8083) );
  NAND2_X1 U7980 ( .A1(n8086), .A2(n8087), .ZN(n8085) );
  NOR2_X1 U7981 ( .A1(n8088), .A2(n7410), .ZN(Result_0_) );
  NOR3_X1 U7982 ( .A1(n8089), .A2(n8090), .A3(n8091), .ZN(n8088) );
  AND2_X1 U7983 ( .A1(n8034), .A2(n8036), .ZN(n8091) );
  NAND2_X1 U7984 ( .A1(n8092), .A2(n8093), .ZN(n8036) );
  NAND2_X1 U7985 ( .A1(n8094), .A2(n8095), .ZN(n8093) );
  XOR2_X1 U7986 ( .A(n7888), .B(n8096), .Z(n8092) );
  NAND2_X1 U7987 ( .A1(n7982), .A2(n8097), .ZN(n8034) );
  NAND2_X1 U7988 ( .A1(n7983), .A2(n7980), .ZN(n8097) );
  NAND2_X1 U7989 ( .A1(n7776), .A2(n8098), .ZN(n7980) );
  NAND2_X1 U7990 ( .A1(n7777), .A2(n7774), .ZN(n8098) );
  NAND2_X1 U7991 ( .A1(n7628), .A2(n8099), .ZN(n7774) );
  NAND2_X1 U7992 ( .A1(n7629), .A2(n7626), .ZN(n8099) );
  NAND2_X1 U7993 ( .A1(n7484), .A2(n8100), .ZN(n7626) );
  NAND2_X1 U7994 ( .A1(n7485), .A2(n7482), .ZN(n8100) );
  NAND2_X1 U7995 ( .A1(n7429), .A2(n8101), .ZN(n7482) );
  NAND2_X1 U7996 ( .A1(n7430), .A2(n7427), .ZN(n8101) );
  NAND2_X1 U7997 ( .A1(n7424), .A2(n8102), .ZN(n7427) );
  NAND2_X1 U7998 ( .A1(n7425), .A2(n7422), .ZN(n8102) );
  NAND2_X1 U7999 ( .A1(n7419), .A2(n8103), .ZN(n7422) );
  NAND2_X1 U8000 ( .A1(n7420), .A2(n7417), .ZN(n8103) );
  NAND2_X1 U8001 ( .A1(n7414), .A2(n8104), .ZN(n7417) );
  NAND2_X1 U8002 ( .A1(n7415), .A2(n7412), .ZN(n8104) );
  NAND2_X1 U8003 ( .A1(n8086), .A2(n8105), .ZN(n7412) );
  NAND2_X1 U8004 ( .A1(n8084), .A2(n8087), .ZN(n8105) );
  NAND2_X1 U8005 ( .A1(n8106), .A2(n8107), .ZN(n8087) );
  XNOR2_X1 U8006 ( .A(n8108), .B(n8109), .ZN(n8106) );
  NAND2_X1 U8007 ( .A1(n8081), .A2(n8110), .ZN(n8084) );
  NAND2_X1 U8008 ( .A1(n8079), .A2(n8082), .ZN(n8110) );
  NAND2_X1 U8009 ( .A1(n8111), .A2(n8112), .ZN(n8082) );
  NAND2_X1 U8010 ( .A1(n8113), .A2(n8107), .ZN(n8112) );
  NAND2_X1 U8011 ( .A1(n8114), .A2(n8115), .ZN(n8111) );
  NAND2_X1 U8012 ( .A1(n8076), .A2(n8116), .ZN(n8079) );
  NAND2_X1 U8013 ( .A1(n8074), .A2(n8077), .ZN(n8116) );
  NAND2_X1 U8014 ( .A1(n8117), .A2(n8118), .ZN(n8077) );
  XNOR2_X1 U8015 ( .A(n8115), .B(n8114), .ZN(n8117) );
  NAND2_X1 U8016 ( .A1(n8071), .A2(n8119), .ZN(n8074) );
  NAND2_X1 U8017 ( .A1(n8069), .A2(n8072), .ZN(n8119) );
  NAND2_X1 U8018 ( .A1(n8120), .A2(n8121), .ZN(n8072) );
  NAND2_X1 U8019 ( .A1(n8122), .A2(n8118), .ZN(n8121) );
  NAND2_X1 U8020 ( .A1(n8123), .A2(n8124), .ZN(n8120) );
  NAND2_X1 U8021 ( .A1(n8066), .A2(n8125), .ZN(n8069) );
  NAND2_X1 U8022 ( .A1(n8067), .A2(n8064), .ZN(n8125) );
  NAND2_X1 U8023 ( .A1(n8061), .A2(n8126), .ZN(n8064) );
  NAND2_X1 U8024 ( .A1(n8062), .A2(n8059), .ZN(n8126) );
  NAND2_X1 U8025 ( .A1(n8056), .A2(n8127), .ZN(n8059) );
  NAND2_X1 U8026 ( .A1(n8054), .A2(n8057), .ZN(n8127) );
  NAND2_X1 U8027 ( .A1(n8128), .A2(n8129), .ZN(n8057) );
  NAND2_X1 U8028 ( .A1(n8130), .A2(n8131), .ZN(n8129) );
  XNOR2_X1 U8029 ( .A(n8132), .B(n8133), .ZN(n8128) );
  NAND2_X1 U8030 ( .A1(n8051), .A2(n8134), .ZN(n8054) );
  NAND2_X1 U8031 ( .A1(n8052), .A2(n8049), .ZN(n8134) );
  NAND2_X1 U8032 ( .A1(n8046), .A2(n8135), .ZN(n8049) );
  NAND2_X1 U8033 ( .A1(n8044), .A2(n8047), .ZN(n8135) );
  NAND2_X1 U8034 ( .A1(n8136), .A2(n8137), .ZN(n8047) );
  NAND2_X1 U8035 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
  XNOR2_X1 U8036 ( .A(n8140), .B(n8141), .ZN(n8136) );
  NAND2_X1 U8037 ( .A1(n8041), .A2(n8142), .ZN(n8044) );
  NAND2_X1 U8038 ( .A1(n8039), .A2(n8042), .ZN(n8142) );
  NAND2_X1 U8039 ( .A1(n8143), .A2(n8144), .ZN(n8042) );
  NAND2_X1 U8040 ( .A1(n8145), .A2(n8146), .ZN(n8144) );
  XNOR2_X1 U8041 ( .A(n8138), .B(n8139), .ZN(n8143) );
  NAND2_X1 U8042 ( .A1(n8032), .A2(n8147), .ZN(n8039) );
  NAND2_X1 U8043 ( .A1(n8029), .A2(n8031), .ZN(n8147) );
  NAND2_X1 U8044 ( .A1(n8148), .A2(n8149), .ZN(n8031) );
  XNOR2_X1 U8045 ( .A(n8146), .B(n8145), .ZN(n8148) );
  NAND2_X1 U8046 ( .A1(n8027), .A2(n8150), .ZN(n8029) );
  NAND2_X1 U8047 ( .A1(n8024), .A2(n8026), .ZN(n8150) );
  NAND2_X1 U8048 ( .A1(n8151), .A2(n8152), .ZN(n8026) );
  NAND2_X1 U8049 ( .A1(n8153), .A2(n8149), .ZN(n8152) );
  NAND2_X1 U8050 ( .A1(n8154), .A2(n8155), .ZN(n8151) );
  NAND2_X1 U8051 ( .A1(n8021), .A2(n8156), .ZN(n8024) );
  NAND2_X1 U8052 ( .A1(n8019), .A2(n8022), .ZN(n8156) );
  NAND2_X1 U8053 ( .A1(n8157), .A2(n8158), .ZN(n8022) );
  NAND2_X1 U8054 ( .A1(n8159), .A2(n8160), .ZN(n8158) );
  XNOR2_X1 U8055 ( .A(n8155), .B(n8154), .ZN(n8157) );
  NAND2_X1 U8056 ( .A1(n8016), .A2(n8161), .ZN(n8019) );
  NAND2_X1 U8057 ( .A1(n8014), .A2(n8017), .ZN(n8161) );
  NAND2_X1 U8058 ( .A1(n8162), .A2(n8163), .ZN(n8017) );
  NAND2_X1 U8059 ( .A1(n8164), .A2(n8165), .ZN(n8163) );
  XNOR2_X1 U8060 ( .A(n8160), .B(n8159), .ZN(n8162) );
  NAND2_X1 U8061 ( .A1(n8012), .A2(n8166), .ZN(n8014) );
  NAND2_X1 U8062 ( .A1(n8009), .A2(n8011), .ZN(n8166) );
  NAND2_X1 U8063 ( .A1(n8167), .A2(n8168), .ZN(n8011) );
  XOR2_X1 U8064 ( .A(n8165), .B(n8169), .Z(n8167) );
  NAND2_X1 U8065 ( .A1(n8007), .A2(n8170), .ZN(n8009) );
  NAND2_X1 U8066 ( .A1(n8004), .A2(n8006), .ZN(n8170) );
  NAND2_X1 U8067 ( .A1(n8171), .A2(n8172), .ZN(n8006) );
  NAND2_X1 U8068 ( .A1(n8173), .A2(n8168), .ZN(n8172) );
  NAND2_X1 U8069 ( .A1(n8174), .A2(n8175), .ZN(n8171) );
  NAND2_X1 U8070 ( .A1(n8002), .A2(n8176), .ZN(n8004) );
  NAND2_X1 U8071 ( .A1(n8000), .A2(n8001), .ZN(n8176) );
  NAND2_X1 U8072 ( .A1(n8177), .A2(n8178), .ZN(n8001) );
  XNOR2_X1 U8073 ( .A(n8174), .B(n8175), .ZN(n8177) );
  NAND2_X1 U8074 ( .A1(n8179), .A2(n8180), .ZN(n8000) );
  OR2_X1 U8075 ( .A1(n7994), .A2(n7996), .ZN(n8180) );
  AND2_X1 U8076 ( .A1(n8181), .A2(n8182), .ZN(n7996) );
  NOR2_X1 U8077 ( .A1(n8183), .A2(n7991), .ZN(n7994) );
  NOR2_X1 U8078 ( .A1(n8184), .A2(n8185), .ZN(n7991) );
  NOR2_X1 U8079 ( .A1(n7992), .A2(n7989), .ZN(n8183) );
  AND2_X1 U8080 ( .A1(n7986), .A2(n8186), .ZN(n7989) );
  NAND2_X1 U8081 ( .A1(n7975), .A2(n7987), .ZN(n8186) );
  NAND2_X1 U8082 ( .A1(n8187), .A2(n8188), .ZN(n7987) );
  NAND2_X1 U8083 ( .A1(n8189), .A2(n8190), .ZN(n8188) );
  XNOR2_X1 U8084 ( .A(n8191), .B(n8192), .ZN(n8187) );
  AND3_X1 U8085 ( .A1(n7978), .A2(n7974), .A3(n7973), .ZN(n7975) );
  XOR2_X1 U8086 ( .A(n8193), .B(n8194), .Z(n7973) );
  XOR2_X1 U8087 ( .A(n8195), .B(n8196), .Z(n8193) );
  NOR2_X1 U8088 ( .A1(n8197), .A2(n7447), .ZN(n8196) );
  NAND2_X1 U8089 ( .A1(n8198), .A2(n8199), .ZN(n7974) );
  NAND3_X1 U8090 ( .A1(a_0_), .A2(n8200), .A3(b_31_), .ZN(n8199) );
  NAND2_X1 U8091 ( .A1(n7970), .A2(n7968), .ZN(n8200) );
  OR2_X1 U8092 ( .A1(n7968), .A2(n7970), .ZN(n8198) );
  AND2_X1 U8093 ( .A1(n8201), .A2(n8202), .ZN(n7970) );
  NAND3_X1 U8094 ( .A1(a_1_), .A2(n8203), .A3(b_31_), .ZN(n8202) );
  OR2_X1 U8095 ( .A1(n7870), .A2(n7869), .ZN(n8203) );
  NAND2_X1 U8096 ( .A1(n7869), .A2(n7870), .ZN(n8201) );
  NAND2_X1 U8097 ( .A1(n8204), .A2(n8205), .ZN(n7870) );
  NAND3_X1 U8098 ( .A1(a_2_), .A2(n8206), .A3(b_31_), .ZN(n8205) );
  NAND2_X1 U8099 ( .A1(n7863), .A2(n7861), .ZN(n8206) );
  OR2_X1 U8100 ( .A1(n7861), .A2(n7863), .ZN(n8204) );
  AND2_X1 U8101 ( .A1(n8207), .A2(n8208), .ZN(n7863) );
  NAND3_X1 U8102 ( .A1(a_3_), .A2(n8209), .A3(b_31_), .ZN(n8208) );
  OR2_X1 U8103 ( .A1(n7850), .A2(n7849), .ZN(n8209) );
  NAND2_X1 U8104 ( .A1(n7849), .A2(n7850), .ZN(n8207) );
  NAND2_X1 U8105 ( .A1(n8210), .A2(n8211), .ZN(n7850) );
  NAND3_X1 U8106 ( .A1(a_4_), .A2(n8212), .A3(b_31_), .ZN(n8211) );
  OR2_X1 U8107 ( .A1(n7834), .A2(n7833), .ZN(n8212) );
  NAND2_X1 U8108 ( .A1(n7833), .A2(n7834), .ZN(n8210) );
  NAND2_X1 U8109 ( .A1(n8213), .A2(n8214), .ZN(n7834) );
  NAND3_X1 U8110 ( .A1(a_5_), .A2(n8215), .A3(b_31_), .ZN(n8214) );
  OR2_X1 U8111 ( .A1(n7821), .A2(n7820), .ZN(n8215) );
  NAND2_X1 U8112 ( .A1(n7820), .A2(n7821), .ZN(n8213) );
  NAND2_X1 U8113 ( .A1(n8216), .A2(n8217), .ZN(n7821) );
  NAND3_X1 U8114 ( .A1(a_6_), .A2(n8218), .A3(b_31_), .ZN(n8217) );
  OR2_X1 U8115 ( .A1(n7805), .A2(n7804), .ZN(n8218) );
  NAND2_X1 U8116 ( .A1(n7804), .A2(n7805), .ZN(n8216) );
  NAND2_X1 U8117 ( .A1(n8219), .A2(n8220), .ZN(n7805) );
  NAND3_X1 U8118 ( .A1(a_7_), .A2(n8221), .A3(b_31_), .ZN(n8220) );
  OR2_X1 U8119 ( .A1(n7793), .A2(n7791), .ZN(n8221) );
  NAND2_X1 U8120 ( .A1(n7791), .A2(n7793), .ZN(n8219) );
  NAND2_X1 U8121 ( .A1(n8222), .A2(n8223), .ZN(n7793) );
  NAND3_X1 U8122 ( .A1(a_8_), .A2(n8224), .A3(b_31_), .ZN(n8223) );
  NAND2_X1 U8123 ( .A1(n7771), .A2(n7769), .ZN(n8224) );
  OR2_X1 U8124 ( .A1(n7769), .A2(n7771), .ZN(n8222) );
  AND2_X1 U8125 ( .A1(n8225), .A2(n8226), .ZN(n7771) );
  NAND3_X1 U8126 ( .A1(a_9_), .A2(n8227), .A3(b_31_), .ZN(n8226) );
  NAND2_X1 U8127 ( .A1(n7759), .A2(n7757), .ZN(n8227) );
  OR2_X1 U8128 ( .A1(n7757), .A2(n7759), .ZN(n8225) );
  AND2_X1 U8129 ( .A1(n8228), .A2(n8229), .ZN(n7759) );
  NAND3_X1 U8130 ( .A1(a_10_), .A2(n8230), .A3(b_31_), .ZN(n8229) );
  NAND2_X1 U8131 ( .A1(n7742), .A2(n7740), .ZN(n8230) );
  OR2_X1 U8132 ( .A1(n7740), .A2(n7742), .ZN(n8228) );
  AND2_X1 U8133 ( .A1(n8231), .A2(n8232), .ZN(n7742) );
  NAND3_X1 U8134 ( .A1(a_11_), .A2(n8233), .A3(b_31_), .ZN(n8232) );
  OR2_X1 U8135 ( .A1(n7730), .A2(n7728), .ZN(n8233) );
  NAND2_X1 U8136 ( .A1(n7728), .A2(n7730), .ZN(n8231) );
  NAND2_X1 U8137 ( .A1(n8234), .A2(n8235), .ZN(n7730) );
  NAND3_X1 U8138 ( .A1(a_12_), .A2(n8236), .A3(b_31_), .ZN(n8235) );
  NAND2_X1 U8139 ( .A1(n7713), .A2(n7711), .ZN(n8236) );
  OR2_X1 U8140 ( .A1(n7711), .A2(n7713), .ZN(n8234) );
  AND2_X1 U8141 ( .A1(n8237), .A2(n8238), .ZN(n7713) );
  NAND3_X1 U8142 ( .A1(a_13_), .A2(n8239), .A3(b_31_), .ZN(n8238) );
  OR2_X1 U8143 ( .A1(n7700), .A2(n7699), .ZN(n8239) );
  NAND2_X1 U8144 ( .A1(n7699), .A2(n7700), .ZN(n8237) );
  NAND2_X1 U8145 ( .A1(n8240), .A2(n8241), .ZN(n7700) );
  NAND3_X1 U8146 ( .A1(a_14_), .A2(n8242), .A3(b_31_), .ZN(n8241) );
  NAND2_X1 U8147 ( .A1(n7685), .A2(n7683), .ZN(n8242) );
  OR2_X1 U8148 ( .A1(n7683), .A2(n7685), .ZN(n8240) );
  AND2_X1 U8149 ( .A1(n8243), .A2(n8244), .ZN(n7685) );
  NAND3_X1 U8150 ( .A1(a_15_), .A2(n8245), .A3(b_31_), .ZN(n8244) );
  OR2_X1 U8151 ( .A1(n7673), .A2(n7672), .ZN(n8245) );
  NAND2_X1 U8152 ( .A1(n7672), .A2(n7673), .ZN(n8243) );
  NAND2_X1 U8153 ( .A1(n8246), .A2(n8247), .ZN(n7673) );
  NAND3_X1 U8154 ( .A1(a_16_), .A2(n8248), .A3(b_31_), .ZN(n8247) );
  NAND2_X1 U8155 ( .A1(n7656), .A2(n7654), .ZN(n8248) );
  OR2_X1 U8156 ( .A1(n7654), .A2(n7656), .ZN(n8246) );
  AND2_X1 U8157 ( .A1(n8249), .A2(n8250), .ZN(n7656) );
  NAND3_X1 U8158 ( .A1(a_17_), .A2(n8251), .A3(b_31_), .ZN(n8250) );
  OR2_X1 U8159 ( .A1(n7643), .A2(n7642), .ZN(n8251) );
  NAND2_X1 U8160 ( .A1(n7642), .A2(n7643), .ZN(n8249) );
  NAND2_X1 U8161 ( .A1(n8252), .A2(n8253), .ZN(n7643) );
  NAND3_X1 U8162 ( .A1(a_18_), .A2(n8254), .A3(b_31_), .ZN(n8253) );
  NAND2_X1 U8163 ( .A1(n7623), .A2(n7621), .ZN(n8254) );
  OR2_X1 U8164 ( .A1(n7621), .A2(n7623), .ZN(n8252) );
  AND2_X1 U8165 ( .A1(n8255), .A2(n8256), .ZN(n7623) );
  NAND3_X1 U8166 ( .A1(a_19_), .A2(n8257), .A3(b_31_), .ZN(n8256) );
  OR2_X1 U8167 ( .A1(n7611), .A2(n7609), .ZN(n8257) );
  NAND2_X1 U8168 ( .A1(n7609), .A2(n7611), .ZN(n8255) );
  NAND2_X1 U8169 ( .A1(n8258), .A2(n8259), .ZN(n7611) );
  NAND3_X1 U8170 ( .A1(a_20_), .A2(n8260), .A3(b_31_), .ZN(n8259) );
  NAND2_X1 U8171 ( .A1(n7596), .A2(n7594), .ZN(n8260) );
  OR2_X1 U8172 ( .A1(n7594), .A2(n7596), .ZN(n8258) );
  AND2_X1 U8173 ( .A1(n8261), .A2(n8262), .ZN(n7596) );
  NAND3_X1 U8174 ( .A1(a_21_), .A2(n8263), .A3(b_31_), .ZN(n8262) );
  NAND2_X1 U8175 ( .A1(n7584), .A2(n7582), .ZN(n8263) );
  OR2_X1 U8176 ( .A1(n7582), .A2(n7584), .ZN(n8261) );
  AND2_X1 U8177 ( .A1(n8264), .A2(n8265), .ZN(n7584) );
  NAND3_X1 U8178 ( .A1(a_22_), .A2(n8266), .A3(b_31_), .ZN(n8265) );
  NAND2_X1 U8179 ( .A1(n7566), .A2(n7564), .ZN(n8266) );
  OR2_X1 U8180 ( .A1(n7564), .A2(n7566), .ZN(n8264) );
  AND2_X1 U8181 ( .A1(n7554), .A2(n8267), .ZN(n7566) );
  NAND2_X1 U8182 ( .A1(n7553), .A2(n7555), .ZN(n8267) );
  NAND2_X1 U8183 ( .A1(n8268), .A2(n8269), .ZN(n7555) );
  NAND2_X1 U8184 ( .A1(b_31_), .A2(a_23_), .ZN(n8269) );
  INV_X1 U8185 ( .A(n8270), .ZN(n8268) );
  XOR2_X1 U8186 ( .A(n8271), .B(n8272), .Z(n7553) );
  XOR2_X1 U8187 ( .A(n8273), .B(n8274), .Z(n8271) );
  NOR2_X1 U8188 ( .A1(n7954), .A2(n7447), .ZN(n8274) );
  NAND2_X1 U8189 ( .A1(a_23_), .A2(n8270), .ZN(n7554) );
  NAND2_X1 U8190 ( .A1(n8275), .A2(n8276), .ZN(n8270) );
  NAND3_X1 U8191 ( .A1(a_24_), .A2(n8277), .A3(b_31_), .ZN(n8276) );
  OR2_X1 U8192 ( .A1(n7540), .A2(n7537), .ZN(n8277) );
  NAND2_X1 U8193 ( .A1(n7537), .A2(n7540), .ZN(n8275) );
  NAND2_X1 U8194 ( .A1(n7527), .A2(n8278), .ZN(n7540) );
  NAND2_X1 U8195 ( .A1(n7526), .A2(n7528), .ZN(n8278) );
  NAND2_X1 U8196 ( .A1(n8279), .A2(n8280), .ZN(n7528) );
  NAND2_X1 U8197 ( .A1(b_31_), .A2(a_25_), .ZN(n8280) );
  INV_X1 U8198 ( .A(n8281), .ZN(n8279) );
  XNOR2_X1 U8199 ( .A(n8282), .B(n8283), .ZN(n7526) );
  NAND2_X1 U8200 ( .A1(n8284), .A2(n8285), .ZN(n8282) );
  NAND2_X1 U8201 ( .A1(a_25_), .A2(n8281), .ZN(n7527) );
  NAND2_X1 U8202 ( .A1(n8286), .A2(n8287), .ZN(n8281) );
  NAND3_X1 U8203 ( .A1(a_26_), .A2(n8288), .A3(b_31_), .ZN(n8287) );
  OR2_X1 U8204 ( .A1(n7511), .A2(n7510), .ZN(n8288) );
  NAND2_X1 U8205 ( .A1(n7510), .A2(n7511), .ZN(n8286) );
  NAND2_X1 U8206 ( .A1(n7499), .A2(n8289), .ZN(n7511) );
  NAND2_X1 U8207 ( .A1(n7498), .A2(n7500), .ZN(n8289) );
  NAND2_X1 U8208 ( .A1(n8290), .A2(n8291), .ZN(n7500) );
  NAND2_X1 U8209 ( .A1(b_31_), .A2(a_27_), .ZN(n8291) );
  INV_X1 U8210 ( .A(n8292), .ZN(n8290) );
  XNOR2_X1 U8211 ( .A(n8293), .B(n8294), .ZN(n7498) );
  XOR2_X1 U8212 ( .A(n8295), .B(n8296), .Z(n8293) );
  NAND2_X1 U8213 ( .A1(b_30_), .A2(a_28_), .ZN(n8295) );
  NAND2_X1 U8214 ( .A1(a_27_), .A2(n8292), .ZN(n7499) );
  NAND2_X1 U8215 ( .A1(n8297), .A2(n8298), .ZN(n8292) );
  NAND3_X1 U8216 ( .A1(a_28_), .A2(n8299), .A3(b_31_), .ZN(n8298) );
  NAND2_X1 U8217 ( .A1(n7478), .A2(n7476), .ZN(n8299) );
  OR2_X1 U8218 ( .A1(n7476), .A2(n7478), .ZN(n8297) );
  AND2_X1 U8219 ( .A1(n8300), .A2(n8301), .ZN(n7478) );
  NAND3_X1 U8220 ( .A1(a_29_), .A2(n8302), .A3(b_31_), .ZN(n8301) );
  OR2_X1 U8221 ( .A1(n7466), .A2(n7467), .ZN(n8302) );
  NAND2_X1 U8222 ( .A1(n7467), .A2(n7466), .ZN(n8300) );
  NAND2_X1 U8223 ( .A1(n8303), .A2(n8304), .ZN(n7466) );
  NAND2_X1 U8224 ( .A1(b_29_), .A2(n8305), .ZN(n8304) );
  NAND2_X1 U8225 ( .A1(n7441), .A2(n8306), .ZN(n8305) );
  NAND2_X1 U8226 ( .A1(a_31_), .A2(n7447), .ZN(n8306) );
  NAND2_X1 U8227 ( .A1(b_30_), .A2(n8307), .ZN(n8303) );
  NAND2_X1 U8228 ( .A1(n7445), .A2(n8308), .ZN(n8307) );
  NAND2_X1 U8229 ( .A1(a_30_), .A2(n7462), .ZN(n8308) );
  AND3_X1 U8230 ( .A1(b_30_), .A2(n7409), .A3(b_31_), .ZN(n7467) );
  XNOR2_X1 U8231 ( .A(n8309), .B(n8310), .ZN(n7476) );
  XOR2_X1 U8232 ( .A(n8311), .B(n8312), .Z(n8309) );
  XNOR2_X1 U8233 ( .A(n8313), .B(n8314), .ZN(n7510) );
  NAND2_X1 U8234 ( .A1(n8315), .A2(n8316), .ZN(n8313) );
  XOR2_X1 U8235 ( .A(n8317), .B(n8318), .Z(n7537) );
  XOR2_X1 U8236 ( .A(n8319), .B(n8320), .Z(n8317) );
  XNOR2_X1 U8237 ( .A(n8321), .B(n8322), .ZN(n7564) );
  XOR2_X1 U8238 ( .A(n8323), .B(n8324), .Z(n8321) );
  XNOR2_X1 U8239 ( .A(n8325), .B(n8326), .ZN(n7582) );
  XOR2_X1 U8240 ( .A(n8327), .B(n8328), .Z(n8325) );
  NOR2_X1 U8241 ( .A1(n7568), .A2(n7447), .ZN(n8328) );
  XNOR2_X1 U8242 ( .A(n8329), .B(n8330), .ZN(n7594) );
  XOR2_X1 U8243 ( .A(n8331), .B(n8332), .Z(n8329) );
  XNOR2_X1 U8244 ( .A(n8333), .B(n8334), .ZN(n7609) );
  XOR2_X1 U8245 ( .A(n8335), .B(n8336), .Z(n8334) );
  NAND2_X1 U8246 ( .A1(b_30_), .A2(a_20_), .ZN(n8336) );
  XOR2_X1 U8247 ( .A(n8337), .B(n8338), .Z(n7621) );
  XNOR2_X1 U8248 ( .A(n8339), .B(n8340), .ZN(n8338) );
  XNOR2_X1 U8249 ( .A(n8341), .B(n8342), .ZN(n7642) );
  XNOR2_X1 U8250 ( .A(n8343), .B(n8344), .ZN(n8341) );
  NOR2_X1 U8251 ( .A1(n7960), .A2(n7447), .ZN(n8344) );
  XOR2_X1 U8252 ( .A(n8345), .B(n8346), .Z(n7654) );
  XNOR2_X1 U8253 ( .A(n8347), .B(n8348), .ZN(n8346) );
  XNOR2_X1 U8254 ( .A(n8349), .B(n8350), .ZN(n7672) );
  XNOR2_X1 U8255 ( .A(n8351), .B(n8352), .ZN(n8349) );
  NOR2_X1 U8256 ( .A1(n8353), .A2(n7447), .ZN(n8352) );
  XOR2_X1 U8257 ( .A(n8354), .B(n8355), .Z(n7683) );
  XNOR2_X1 U8258 ( .A(n8356), .B(n8357), .ZN(n8355) );
  XNOR2_X1 U8259 ( .A(n8358), .B(n8359), .ZN(n7699) );
  XNOR2_X1 U8260 ( .A(n8360), .B(n8361), .ZN(n8358) );
  NOR2_X1 U8261 ( .A1(n7962), .A2(n7447), .ZN(n8361) );
  XNOR2_X1 U8262 ( .A(n8362), .B(n8363), .ZN(n7711) );
  XOR2_X1 U8263 ( .A(n8364), .B(n8365), .Z(n8362) );
  XNOR2_X1 U8264 ( .A(n8366), .B(n8367), .ZN(n7728) );
  XOR2_X1 U8265 ( .A(n8368), .B(n8369), .Z(n8367) );
  NAND2_X1 U8266 ( .A1(b_30_), .A2(a_12_), .ZN(n8369) );
  XOR2_X1 U8267 ( .A(n8370), .B(n8371), .Z(n7740) );
  XNOR2_X1 U8268 ( .A(n8372), .B(n8373), .ZN(n8371) );
  XNOR2_X1 U8269 ( .A(n8374), .B(n8375), .ZN(n7757) );
  XOR2_X1 U8270 ( .A(n8376), .B(n8377), .Z(n8374) );
  NOR2_X1 U8271 ( .A1(n8378), .A2(n7447), .ZN(n8377) );
  XNOR2_X1 U8272 ( .A(n8379), .B(n8380), .ZN(n7769) );
  XOR2_X1 U8273 ( .A(n8381), .B(n8382), .Z(n8379) );
  XNOR2_X1 U8274 ( .A(n8383), .B(n8384), .ZN(n7791) );
  XOR2_X1 U8275 ( .A(n8385), .B(n8386), .Z(n8384) );
  NAND2_X1 U8276 ( .A1(b_30_), .A2(a_8_), .ZN(n8386) );
  XNOR2_X1 U8277 ( .A(n8387), .B(n8388), .ZN(n7804) );
  XNOR2_X1 U8278 ( .A(n8389), .B(n8390), .ZN(n8388) );
  XNOR2_X1 U8279 ( .A(n8391), .B(n8392), .ZN(n7820) );
  XNOR2_X1 U8280 ( .A(n8393), .B(n8394), .ZN(n8391) );
  NOR2_X1 U8281 ( .A1(n7807), .A2(n7447), .ZN(n8394) );
  XNOR2_X1 U8282 ( .A(n8395), .B(n8396), .ZN(n7833) );
  XNOR2_X1 U8283 ( .A(n8397), .B(n8398), .ZN(n8396) );
  XNOR2_X1 U8284 ( .A(n8399), .B(n8400), .ZN(n7849) );
  XOR2_X1 U8285 ( .A(n8401), .B(n8402), .Z(n8400) );
  NAND2_X1 U8286 ( .A1(b_30_), .A2(a_4_), .ZN(n8402) );
  XOR2_X1 U8287 ( .A(n8403), .B(n8404), .Z(n7861) );
  XNOR2_X1 U8288 ( .A(n8405), .B(n8406), .ZN(n8404) );
  XNOR2_X1 U8289 ( .A(n8407), .B(n8408), .ZN(n7869) );
  XNOR2_X1 U8290 ( .A(n8409), .B(n8410), .ZN(n8407) );
  NOR2_X1 U8291 ( .A1(n7966), .A2(n7447), .ZN(n8410) );
  XOR2_X1 U8292 ( .A(n8411), .B(n8412), .Z(n7968) );
  XOR2_X1 U8293 ( .A(n8413), .B(n8414), .Z(n8412) );
  NAND2_X1 U8294 ( .A1(b_30_), .A2(a_1_), .ZN(n8414) );
  XOR2_X1 U8295 ( .A(n8190), .B(n8189), .Z(n7978) );
  NAND4_X1 U8296 ( .A1(n8189), .A2(n8415), .A3(n8190), .A4(n8185), .ZN(n7986)
         );
  NAND2_X1 U8297 ( .A1(n8416), .A2(n8417), .ZN(n8190) );
  NAND3_X1 U8298 ( .A1(a_0_), .A2(n8418), .A3(b_30_), .ZN(n8417) );
  OR2_X1 U8299 ( .A1(n8195), .A2(n8194), .ZN(n8418) );
  NAND2_X1 U8300 ( .A1(n8194), .A2(n8195), .ZN(n8416) );
  NAND2_X1 U8301 ( .A1(n8419), .A2(n8420), .ZN(n8195) );
  NAND3_X1 U8302 ( .A1(a_1_), .A2(n8421), .A3(b_30_), .ZN(n8420) );
  OR2_X1 U8303 ( .A1(n8411), .A2(n8413), .ZN(n8421) );
  NAND2_X1 U8304 ( .A1(n8411), .A2(n8413), .ZN(n8419) );
  NAND2_X1 U8305 ( .A1(n8422), .A2(n8423), .ZN(n8413) );
  NAND3_X1 U8306 ( .A1(a_2_), .A2(n8424), .A3(b_30_), .ZN(n8423) );
  NAND2_X1 U8307 ( .A1(n8409), .A2(n8408), .ZN(n8424) );
  OR2_X1 U8308 ( .A1(n8408), .A2(n8409), .ZN(n8422) );
  AND2_X1 U8309 ( .A1(n8425), .A2(n8426), .ZN(n8409) );
  NAND2_X1 U8310 ( .A1(n8406), .A2(n8427), .ZN(n8426) );
  OR2_X1 U8311 ( .A1(n8403), .A2(n8405), .ZN(n8427) );
  NOR2_X1 U8312 ( .A1(n7447), .A2(n7852), .ZN(n8406) );
  NAND2_X1 U8313 ( .A1(n8403), .A2(n8405), .ZN(n8425) );
  NAND2_X1 U8314 ( .A1(n8428), .A2(n8429), .ZN(n8405) );
  NAND3_X1 U8315 ( .A1(a_4_), .A2(n8430), .A3(b_30_), .ZN(n8429) );
  OR2_X1 U8316 ( .A1(n8401), .A2(n8399), .ZN(n8430) );
  NAND2_X1 U8317 ( .A1(n8399), .A2(n8401), .ZN(n8428) );
  NAND2_X1 U8318 ( .A1(n8431), .A2(n8432), .ZN(n8401) );
  NAND2_X1 U8319 ( .A1(n8398), .A2(n8433), .ZN(n8432) );
  OR2_X1 U8320 ( .A1(n8397), .A2(n8395), .ZN(n8433) );
  NOR2_X1 U8321 ( .A1(n7447), .A2(n7823), .ZN(n8398) );
  NAND2_X1 U8322 ( .A1(n8395), .A2(n8397), .ZN(n8431) );
  NAND2_X1 U8323 ( .A1(n8434), .A2(n8435), .ZN(n8397) );
  NAND3_X1 U8324 ( .A1(a_6_), .A2(n8436), .A3(b_30_), .ZN(n8435) );
  NAND2_X1 U8325 ( .A1(n8393), .A2(n8392), .ZN(n8436) );
  OR2_X1 U8326 ( .A1(n8392), .A2(n8393), .ZN(n8434) );
  AND2_X1 U8327 ( .A1(n8437), .A2(n8438), .ZN(n8393) );
  NAND2_X1 U8328 ( .A1(n8390), .A2(n8439), .ZN(n8438) );
  OR2_X1 U8329 ( .A1(n8389), .A2(n8387), .ZN(n8439) );
  NOR2_X1 U8330 ( .A1(n7447), .A2(n7787), .ZN(n8390) );
  NAND2_X1 U8331 ( .A1(n8387), .A2(n8389), .ZN(n8437) );
  NAND2_X1 U8332 ( .A1(n8440), .A2(n8441), .ZN(n8389) );
  NAND3_X1 U8333 ( .A1(a_8_), .A2(n8442), .A3(b_30_), .ZN(n8441) );
  OR2_X1 U8334 ( .A1(n8385), .A2(n8383), .ZN(n8442) );
  NAND2_X1 U8335 ( .A1(n8383), .A2(n8385), .ZN(n8440) );
  NAND2_X1 U8336 ( .A1(n8443), .A2(n8444), .ZN(n8385) );
  NAND2_X1 U8337 ( .A1(n8382), .A2(n8445), .ZN(n8444) );
  OR2_X1 U8338 ( .A1(n8380), .A2(n8381), .ZN(n8445) );
  NOR2_X1 U8339 ( .A1(n7447), .A2(n7753), .ZN(n8382) );
  NAND2_X1 U8340 ( .A1(n8380), .A2(n8381), .ZN(n8443) );
  NAND2_X1 U8341 ( .A1(n8446), .A2(n8447), .ZN(n8381) );
  NAND3_X1 U8342 ( .A1(a_10_), .A2(n8448), .A3(b_30_), .ZN(n8447) );
  OR2_X1 U8343 ( .A1(n8375), .A2(n8376), .ZN(n8448) );
  NAND2_X1 U8344 ( .A1(n8375), .A2(n8376), .ZN(n8446) );
  NAND2_X1 U8345 ( .A1(n8449), .A2(n8450), .ZN(n8376) );
  NAND2_X1 U8346 ( .A1(n8373), .A2(n8451), .ZN(n8450) );
  OR2_X1 U8347 ( .A1(n8370), .A2(n8372), .ZN(n8451) );
  NOR2_X1 U8348 ( .A1(n7447), .A2(n7724), .ZN(n8373) );
  NAND2_X1 U8349 ( .A1(n8370), .A2(n8372), .ZN(n8449) );
  NAND2_X1 U8350 ( .A1(n8452), .A2(n8453), .ZN(n8372) );
  NAND3_X1 U8351 ( .A1(a_12_), .A2(n8454), .A3(b_30_), .ZN(n8453) );
  OR2_X1 U8352 ( .A1(n8368), .A2(n8366), .ZN(n8454) );
  NAND2_X1 U8353 ( .A1(n8366), .A2(n8368), .ZN(n8452) );
  NAND2_X1 U8354 ( .A1(n8455), .A2(n8456), .ZN(n8368) );
  NAND2_X1 U8355 ( .A1(n8365), .A2(n8457), .ZN(n8456) );
  OR2_X1 U8356 ( .A1(n8363), .A2(n8364), .ZN(n8457) );
  NOR2_X1 U8357 ( .A1(n7447), .A2(n7702), .ZN(n8365) );
  NAND2_X1 U8358 ( .A1(n8363), .A2(n8364), .ZN(n8455) );
  NAND2_X1 U8359 ( .A1(n8458), .A2(n8459), .ZN(n8364) );
  NAND3_X1 U8360 ( .A1(a_14_), .A2(n8460), .A3(b_30_), .ZN(n8459) );
  NAND2_X1 U8361 ( .A1(n8360), .A2(n8359), .ZN(n8460) );
  OR2_X1 U8362 ( .A1(n8359), .A2(n8360), .ZN(n8458) );
  AND2_X1 U8363 ( .A1(n8461), .A2(n8462), .ZN(n8360) );
  NAND2_X1 U8364 ( .A1(n8357), .A2(n8463), .ZN(n8462) );
  OR2_X1 U8365 ( .A1(n8354), .A2(n8356), .ZN(n8463) );
  NOR2_X1 U8366 ( .A1(n7447), .A2(n7667), .ZN(n8357) );
  NAND2_X1 U8367 ( .A1(n8354), .A2(n8356), .ZN(n8461) );
  NAND2_X1 U8368 ( .A1(n8464), .A2(n8465), .ZN(n8356) );
  NAND3_X1 U8369 ( .A1(a_16_), .A2(n8466), .A3(b_30_), .ZN(n8465) );
  NAND2_X1 U8370 ( .A1(n8351), .A2(n8350), .ZN(n8466) );
  OR2_X1 U8371 ( .A1(n8350), .A2(n8351), .ZN(n8464) );
  AND2_X1 U8372 ( .A1(n8467), .A2(n8468), .ZN(n8351) );
  NAND2_X1 U8373 ( .A1(n8348), .A2(n8469), .ZN(n8468) );
  OR2_X1 U8374 ( .A1(n8345), .A2(n8347), .ZN(n8469) );
  NOR2_X1 U8375 ( .A1(n7447), .A2(n7645), .ZN(n8348) );
  NAND2_X1 U8376 ( .A1(n8345), .A2(n8347), .ZN(n8467) );
  NAND2_X1 U8377 ( .A1(n8470), .A2(n8471), .ZN(n8347) );
  NAND3_X1 U8378 ( .A1(a_18_), .A2(n8472), .A3(b_30_), .ZN(n8471) );
  NAND2_X1 U8379 ( .A1(n8343), .A2(n8342), .ZN(n8472) );
  OR2_X1 U8380 ( .A1(n8342), .A2(n8343), .ZN(n8470) );
  AND2_X1 U8381 ( .A1(n8473), .A2(n8474), .ZN(n8343) );
  NAND2_X1 U8382 ( .A1(n8340), .A2(n8475), .ZN(n8474) );
  OR2_X1 U8383 ( .A1(n8337), .A2(n8339), .ZN(n8475) );
  NOR2_X1 U8384 ( .A1(n7447), .A2(n7958), .ZN(n8340) );
  NAND2_X1 U8385 ( .A1(n8337), .A2(n8339), .ZN(n8473) );
  NAND2_X1 U8386 ( .A1(n8476), .A2(n8477), .ZN(n8339) );
  NAND3_X1 U8387 ( .A1(a_20_), .A2(n8478), .A3(b_30_), .ZN(n8477) );
  OR2_X1 U8388 ( .A1(n8335), .A2(n8333), .ZN(n8478) );
  NAND2_X1 U8389 ( .A1(n8333), .A2(n8335), .ZN(n8476) );
  NAND2_X1 U8390 ( .A1(n8479), .A2(n8480), .ZN(n8335) );
  NAND2_X1 U8391 ( .A1(n8332), .A2(n8481), .ZN(n8480) );
  OR2_X1 U8392 ( .A1(n8330), .A2(n8331), .ZN(n8481) );
  NOR2_X1 U8393 ( .A1(n7447), .A2(n7578), .ZN(n8332) );
  NAND2_X1 U8394 ( .A1(n8330), .A2(n8331), .ZN(n8479) );
  NAND2_X1 U8395 ( .A1(n8482), .A2(n8483), .ZN(n8331) );
  NAND3_X1 U8396 ( .A1(a_22_), .A2(n8484), .A3(b_30_), .ZN(n8483) );
  OR2_X1 U8397 ( .A1(n8326), .A2(n8327), .ZN(n8484) );
  NAND2_X1 U8398 ( .A1(n8326), .A2(n8327), .ZN(n8482) );
  NAND2_X1 U8399 ( .A1(n8485), .A2(n8486), .ZN(n8327) );
  NAND2_X1 U8400 ( .A1(n8324), .A2(n8487), .ZN(n8486) );
  OR2_X1 U8401 ( .A1(n8322), .A2(n8323), .ZN(n8487) );
  NOR2_X1 U8402 ( .A1(n7447), .A2(n7955), .ZN(n8324) );
  NAND2_X1 U8403 ( .A1(n8322), .A2(n8323), .ZN(n8485) );
  NAND2_X1 U8404 ( .A1(n8488), .A2(n8489), .ZN(n8323) );
  NAND3_X1 U8405 ( .A1(a_24_), .A2(n8490), .A3(b_30_), .ZN(n8489) );
  OR2_X1 U8406 ( .A1(n8272), .A2(n8273), .ZN(n8490) );
  NAND2_X1 U8407 ( .A1(n8272), .A2(n8273), .ZN(n8488) );
  NAND2_X1 U8408 ( .A1(n8491), .A2(n8492), .ZN(n8273) );
  NAND2_X1 U8409 ( .A1(n8320), .A2(n8493), .ZN(n8492) );
  OR2_X1 U8410 ( .A1(n8318), .A2(n8319), .ZN(n8493) );
  NOR2_X1 U8411 ( .A1(n7447), .A2(n7952), .ZN(n8320) );
  NAND2_X1 U8412 ( .A1(n8318), .A2(n8319), .ZN(n8491) );
  NAND2_X1 U8413 ( .A1(n8284), .A2(n8494), .ZN(n8319) );
  NAND2_X1 U8414 ( .A1(n8283), .A2(n8285), .ZN(n8494) );
  NAND2_X1 U8415 ( .A1(n8495), .A2(n8496), .ZN(n8285) );
  NAND2_X1 U8416 ( .A1(b_30_), .A2(a_26_), .ZN(n8496) );
  INV_X1 U8417 ( .A(n8497), .ZN(n8495) );
  XNOR2_X1 U8418 ( .A(n8498), .B(n8499), .ZN(n8283) );
  NAND2_X1 U8419 ( .A1(n8500), .A2(n8501), .ZN(n8498) );
  NAND2_X1 U8420 ( .A1(a_26_), .A2(n8497), .ZN(n8284) );
  NAND2_X1 U8421 ( .A1(n8315), .A2(n8502), .ZN(n8497) );
  NAND2_X1 U8422 ( .A1(n8314), .A2(n8316), .ZN(n8502) );
  NAND2_X1 U8423 ( .A1(n8503), .A2(n8504), .ZN(n8316) );
  NAND2_X1 U8424 ( .A1(b_30_), .A2(a_27_), .ZN(n8504) );
  INV_X1 U8425 ( .A(n8505), .ZN(n8503) );
  XNOR2_X1 U8426 ( .A(n8506), .B(n8507), .ZN(n8314) );
  XOR2_X1 U8427 ( .A(n8508), .B(n8509), .Z(n8506) );
  NAND2_X1 U8428 ( .A1(b_29_), .A2(a_28_), .ZN(n8508) );
  NAND2_X1 U8429 ( .A1(a_27_), .A2(n8505), .ZN(n8315) );
  NAND2_X1 U8430 ( .A1(n8510), .A2(n8511), .ZN(n8505) );
  NAND3_X1 U8431 ( .A1(a_28_), .A2(n8512), .A3(b_30_), .ZN(n8511) );
  NAND2_X1 U8432 ( .A1(n8296), .A2(n8294), .ZN(n8512) );
  OR2_X1 U8433 ( .A1(n8294), .A2(n8296), .ZN(n8510) );
  AND2_X1 U8434 ( .A1(n8513), .A2(n8514), .ZN(n8296) );
  NAND2_X1 U8435 ( .A1(n8310), .A2(n8515), .ZN(n8514) );
  OR2_X1 U8436 ( .A1(n8311), .A2(n8312), .ZN(n8515) );
  NOR2_X1 U8437 ( .A1(n7447), .A2(n7460), .ZN(n8310) );
  INV_X1 U8438 ( .A(b_30_), .ZN(n7447) );
  NAND2_X1 U8439 ( .A1(n8312), .A2(n8311), .ZN(n8513) );
  NAND2_X1 U8440 ( .A1(n8516), .A2(n8517), .ZN(n8311) );
  NAND2_X1 U8441 ( .A1(b_28_), .A2(n8518), .ZN(n8517) );
  NAND2_X1 U8442 ( .A1(n7441), .A2(n8519), .ZN(n8518) );
  NAND2_X1 U8443 ( .A1(a_31_), .A2(n7462), .ZN(n8519) );
  NAND2_X1 U8444 ( .A1(b_29_), .A2(n8520), .ZN(n8516) );
  NAND2_X1 U8445 ( .A1(n7445), .A2(n8521), .ZN(n8520) );
  NAND2_X1 U8446 ( .A1(a_30_), .A2(n7949), .ZN(n8521) );
  AND3_X1 U8447 ( .A1(b_29_), .A2(n7409), .A3(b_30_), .ZN(n8312) );
  XNOR2_X1 U8448 ( .A(n8522), .B(n7457), .ZN(n8294) );
  XOR2_X1 U8449 ( .A(n8523), .B(n8524), .Z(n8522) );
  XNOR2_X1 U8450 ( .A(n8525), .B(n8526), .ZN(n8318) );
  NAND2_X1 U8451 ( .A1(n8527), .A2(n8528), .ZN(n8525) );
  XNOR2_X1 U8452 ( .A(n8529), .B(n8530), .ZN(n8272) );
  XNOR2_X1 U8453 ( .A(n8531), .B(n8532), .ZN(n8529) );
  XNOR2_X1 U8454 ( .A(n8533), .B(n8534), .ZN(n8322) );
  XOR2_X1 U8455 ( .A(n8535), .B(n8536), .Z(n8534) );
  NAND2_X1 U8456 ( .A1(b_29_), .A2(a_24_), .ZN(n8536) );
  XNOR2_X1 U8457 ( .A(n8537), .B(n8538), .ZN(n8326) );
  XNOR2_X1 U8458 ( .A(n8539), .B(n8540), .ZN(n8538) );
  XNOR2_X1 U8459 ( .A(n8541), .B(n8542), .ZN(n8330) );
  XOR2_X1 U8460 ( .A(n8543), .B(n8544), .Z(n8542) );
  NAND2_X1 U8461 ( .A1(b_29_), .A2(a_22_), .ZN(n8544) );
  XOR2_X1 U8462 ( .A(n8545), .B(n8546), .Z(n8333) );
  XOR2_X1 U8463 ( .A(n8547), .B(n8548), .Z(n8545) );
  XNOR2_X1 U8464 ( .A(n8549), .B(n8550), .ZN(n8337) );
  XNOR2_X1 U8465 ( .A(n8551), .B(n8552), .ZN(n8549) );
  NOR2_X1 U8466 ( .A1(n7957), .A2(n7462), .ZN(n8552) );
  XOR2_X1 U8467 ( .A(n8553), .B(n8554), .Z(n8342) );
  XNOR2_X1 U8468 ( .A(n8555), .B(n8556), .ZN(n8554) );
  XNOR2_X1 U8469 ( .A(n8557), .B(n8558), .ZN(n8345) );
  XNOR2_X1 U8470 ( .A(n8559), .B(n8560), .ZN(n8557) );
  NOR2_X1 U8471 ( .A1(n7960), .A2(n7462), .ZN(n8560) );
  XNOR2_X1 U8472 ( .A(n8561), .B(n8562), .ZN(n8350) );
  XOR2_X1 U8473 ( .A(n8563), .B(n8564), .Z(n8561) );
  XNOR2_X1 U8474 ( .A(n8565), .B(n8566), .ZN(n8354) );
  XOR2_X1 U8475 ( .A(n8567), .B(n8568), .Z(n8566) );
  NAND2_X1 U8476 ( .A1(b_29_), .A2(a_16_), .ZN(n8568) );
  XOR2_X1 U8477 ( .A(n8569), .B(n8570), .Z(n8359) );
  XNOR2_X1 U8478 ( .A(n8571), .B(n8572), .ZN(n8570) );
  XNOR2_X1 U8479 ( .A(n8573), .B(n8574), .ZN(n8363) );
  XNOR2_X1 U8480 ( .A(n8575), .B(n8576), .ZN(n8573) );
  NOR2_X1 U8481 ( .A1(n7962), .A2(n7462), .ZN(n8576) );
  XNOR2_X1 U8482 ( .A(n8577), .B(n8578), .ZN(n8366) );
  XNOR2_X1 U8483 ( .A(n8579), .B(n8580), .ZN(n8578) );
  XNOR2_X1 U8484 ( .A(n8581), .B(n8582), .ZN(n8370) );
  XNOR2_X1 U8485 ( .A(n8583), .B(n8584), .ZN(n8581) );
  NOR2_X1 U8486 ( .A1(n8585), .A2(n7462), .ZN(n8584) );
  XNOR2_X1 U8487 ( .A(n8586), .B(n8587), .ZN(n8375) );
  XNOR2_X1 U8488 ( .A(n8588), .B(n8589), .ZN(n8587) );
  XNOR2_X1 U8489 ( .A(n8590), .B(n8591), .ZN(n8380) );
  XNOR2_X1 U8490 ( .A(n8592), .B(n8593), .ZN(n8590) );
  NOR2_X1 U8491 ( .A1(n8378), .A2(n7462), .ZN(n8593) );
  XOR2_X1 U8492 ( .A(n8594), .B(n8595), .Z(n8383) );
  XOR2_X1 U8493 ( .A(n8596), .B(n8597), .Z(n8594) );
  XOR2_X1 U8494 ( .A(n8598), .B(n8599), .Z(n8387) );
  XOR2_X1 U8495 ( .A(n8600), .B(n8601), .Z(n8598) );
  NOR2_X1 U8496 ( .A1(n8602), .A2(n7462), .ZN(n8601) );
  XOR2_X1 U8497 ( .A(n8603), .B(n8604), .Z(n8392) );
  XNOR2_X1 U8498 ( .A(n8605), .B(n8606), .ZN(n8604) );
  XOR2_X1 U8499 ( .A(n8607), .B(n8608), .Z(n8395) );
  XOR2_X1 U8500 ( .A(n8609), .B(n8610), .Z(n8607) );
  NOR2_X1 U8501 ( .A1(n7807), .A2(n7462), .ZN(n8610) );
  XOR2_X1 U8502 ( .A(n8611), .B(n8612), .Z(n8399) );
  XOR2_X1 U8503 ( .A(n8613), .B(n8614), .Z(n8611) );
  XNOR2_X1 U8504 ( .A(n8615), .B(n8616), .ZN(n8403) );
  XNOR2_X1 U8505 ( .A(n8617), .B(n8618), .ZN(n8615) );
  NOR2_X1 U8506 ( .A1(n7836), .A2(n7462), .ZN(n8618) );
  XOR2_X1 U8507 ( .A(n8619), .B(n8620), .Z(n8408) );
  XOR2_X1 U8508 ( .A(n8621), .B(n8622), .Z(n8620) );
  NAND2_X1 U8509 ( .A1(b_29_), .A2(a_3_), .ZN(n8622) );
  XNOR2_X1 U8510 ( .A(n8623), .B(n8624), .ZN(n8411) );
  XNOR2_X1 U8511 ( .A(n8625), .B(n8626), .ZN(n8623) );
  XNOR2_X1 U8512 ( .A(n8627), .B(n8628), .ZN(n8194) );
  XNOR2_X1 U8513 ( .A(n8629), .B(n8630), .ZN(n8627) );
  NOR2_X1 U8514 ( .A1(n7872), .A2(n7462), .ZN(n8630) );
  NAND2_X1 U8515 ( .A1(n8191), .A2(n8192), .ZN(n8415) );
  XNOR2_X1 U8516 ( .A(n8631), .B(n8632), .ZN(n8189) );
  NAND2_X1 U8517 ( .A1(n8633), .A2(n8634), .ZN(n8631) );
  AND2_X1 U8518 ( .A1(n8185), .A2(n8184), .ZN(n7992) );
  NAND2_X1 U8519 ( .A1(n8181), .A2(n8635), .ZN(n8184) );
  NAND2_X1 U8520 ( .A1(n8636), .A2(n8637), .ZN(n8635) );
  OR2_X1 U8521 ( .A1(n8192), .A2(n8191), .ZN(n8185) );
  AND2_X1 U8522 ( .A1(n8633), .A2(n8638), .ZN(n8191) );
  NAND2_X1 U8523 ( .A1(n8632), .A2(n8634), .ZN(n8638) );
  NAND2_X1 U8524 ( .A1(n8639), .A2(n8640), .ZN(n8634) );
  NAND2_X1 U8525 ( .A1(b_29_), .A2(a_0_), .ZN(n8640) );
  INV_X1 U8526 ( .A(n8641), .ZN(n8639) );
  XOR2_X1 U8527 ( .A(n8642), .B(n8643), .Z(n8632) );
  XOR2_X1 U8528 ( .A(n8644), .B(n8645), .Z(n8642) );
  NAND2_X1 U8529 ( .A1(a_0_), .A2(n8641), .ZN(n8633) );
  NAND2_X1 U8530 ( .A1(n8646), .A2(n8647), .ZN(n8641) );
  NAND3_X1 U8531 ( .A1(a_1_), .A2(n8648), .A3(b_29_), .ZN(n8647) );
  NAND2_X1 U8532 ( .A1(n8629), .A2(n8628), .ZN(n8648) );
  OR2_X1 U8533 ( .A1(n8628), .A2(n8629), .ZN(n8646) );
  AND2_X1 U8534 ( .A1(n8649), .A2(n8650), .ZN(n8629) );
  NAND2_X1 U8535 ( .A1(n8625), .A2(n8651), .ZN(n8650) );
  NAND2_X1 U8536 ( .A1(n8624), .A2(n8626), .ZN(n8651) );
  NAND2_X1 U8537 ( .A1(n8652), .A2(n8653), .ZN(n8625) );
  NAND3_X1 U8538 ( .A1(a_3_), .A2(n8654), .A3(b_29_), .ZN(n8653) );
  OR2_X1 U8539 ( .A1(n8621), .A2(n8619), .ZN(n8654) );
  NAND2_X1 U8540 ( .A1(n8619), .A2(n8621), .ZN(n8652) );
  NAND2_X1 U8541 ( .A1(n8655), .A2(n8656), .ZN(n8621) );
  NAND3_X1 U8542 ( .A1(a_4_), .A2(n8657), .A3(b_29_), .ZN(n8656) );
  NAND2_X1 U8543 ( .A1(n8617), .A2(n8616), .ZN(n8657) );
  OR2_X1 U8544 ( .A1(n8616), .A2(n8617), .ZN(n8655) );
  AND2_X1 U8545 ( .A1(n8658), .A2(n8659), .ZN(n8617) );
  NAND2_X1 U8546 ( .A1(n8614), .A2(n8660), .ZN(n8659) );
  OR2_X1 U8547 ( .A1(n8613), .A2(n8612), .ZN(n8660) );
  NOR2_X1 U8548 ( .A1(n7462), .A2(n7823), .ZN(n8614) );
  NAND2_X1 U8549 ( .A1(n8612), .A2(n8613), .ZN(n8658) );
  NAND2_X1 U8550 ( .A1(n8661), .A2(n8662), .ZN(n8613) );
  NAND3_X1 U8551 ( .A1(a_6_), .A2(n8663), .A3(b_29_), .ZN(n8662) );
  OR2_X1 U8552 ( .A1(n8609), .A2(n8608), .ZN(n8663) );
  NAND2_X1 U8553 ( .A1(n8608), .A2(n8609), .ZN(n8661) );
  NAND2_X1 U8554 ( .A1(n8664), .A2(n8665), .ZN(n8609) );
  NAND2_X1 U8555 ( .A1(n8606), .A2(n8666), .ZN(n8665) );
  OR2_X1 U8556 ( .A1(n8605), .A2(n8603), .ZN(n8666) );
  NOR2_X1 U8557 ( .A1(n7462), .A2(n7787), .ZN(n8606) );
  NAND2_X1 U8558 ( .A1(n8603), .A2(n8605), .ZN(n8664) );
  NAND2_X1 U8559 ( .A1(n8667), .A2(n8668), .ZN(n8605) );
  NAND3_X1 U8560 ( .A1(a_8_), .A2(n8669), .A3(b_29_), .ZN(n8668) );
  OR2_X1 U8561 ( .A1(n8600), .A2(n8599), .ZN(n8669) );
  NAND2_X1 U8562 ( .A1(n8599), .A2(n8600), .ZN(n8667) );
  NAND2_X1 U8563 ( .A1(n8670), .A2(n8671), .ZN(n8600) );
  NAND2_X1 U8564 ( .A1(n8597), .A2(n8672), .ZN(n8671) );
  OR2_X1 U8565 ( .A1(n8596), .A2(n8595), .ZN(n8672) );
  NOR2_X1 U8566 ( .A1(n7462), .A2(n7753), .ZN(n8597) );
  NAND2_X1 U8567 ( .A1(n8595), .A2(n8596), .ZN(n8670) );
  NAND2_X1 U8568 ( .A1(n8673), .A2(n8674), .ZN(n8596) );
  NAND3_X1 U8569 ( .A1(a_10_), .A2(n8675), .A3(b_29_), .ZN(n8674) );
  NAND2_X1 U8570 ( .A1(n8592), .A2(n8591), .ZN(n8675) );
  OR2_X1 U8571 ( .A1(n8591), .A2(n8592), .ZN(n8673) );
  AND2_X1 U8572 ( .A1(n8676), .A2(n8677), .ZN(n8592) );
  NAND2_X1 U8573 ( .A1(n8589), .A2(n8678), .ZN(n8677) );
  OR2_X1 U8574 ( .A1(n8588), .A2(n8586), .ZN(n8678) );
  NOR2_X1 U8575 ( .A1(n7462), .A2(n7724), .ZN(n8589) );
  NAND2_X1 U8576 ( .A1(n8586), .A2(n8588), .ZN(n8676) );
  NAND2_X1 U8577 ( .A1(n8679), .A2(n8680), .ZN(n8588) );
  NAND3_X1 U8578 ( .A1(a_12_), .A2(n8681), .A3(b_29_), .ZN(n8680) );
  NAND2_X1 U8579 ( .A1(n8583), .A2(n8582), .ZN(n8681) );
  OR2_X1 U8580 ( .A1(n8582), .A2(n8583), .ZN(n8679) );
  AND2_X1 U8581 ( .A1(n8682), .A2(n8683), .ZN(n8583) );
  NAND2_X1 U8582 ( .A1(n8580), .A2(n8684), .ZN(n8683) );
  OR2_X1 U8583 ( .A1(n8579), .A2(n8577), .ZN(n8684) );
  NOR2_X1 U8584 ( .A1(n7462), .A2(n7702), .ZN(n8580) );
  NAND2_X1 U8585 ( .A1(n8577), .A2(n8579), .ZN(n8682) );
  NAND2_X1 U8586 ( .A1(n8685), .A2(n8686), .ZN(n8579) );
  NAND3_X1 U8587 ( .A1(a_14_), .A2(n8687), .A3(b_29_), .ZN(n8686) );
  NAND2_X1 U8588 ( .A1(n8575), .A2(n8574), .ZN(n8687) );
  OR2_X1 U8589 ( .A1(n8574), .A2(n8575), .ZN(n8685) );
  AND2_X1 U8590 ( .A1(n8688), .A2(n8689), .ZN(n8575) );
  NAND2_X1 U8591 ( .A1(n8572), .A2(n8690), .ZN(n8689) );
  OR2_X1 U8592 ( .A1(n8571), .A2(n8569), .ZN(n8690) );
  NOR2_X1 U8593 ( .A1(n7462), .A2(n7667), .ZN(n8572) );
  NAND2_X1 U8594 ( .A1(n8569), .A2(n8571), .ZN(n8688) );
  NAND2_X1 U8595 ( .A1(n8691), .A2(n8692), .ZN(n8571) );
  NAND3_X1 U8596 ( .A1(a_16_), .A2(n8693), .A3(b_29_), .ZN(n8692) );
  OR2_X1 U8597 ( .A1(n8567), .A2(n8565), .ZN(n8693) );
  NAND2_X1 U8598 ( .A1(n8565), .A2(n8567), .ZN(n8691) );
  NAND2_X1 U8599 ( .A1(n8694), .A2(n8695), .ZN(n8567) );
  NAND2_X1 U8600 ( .A1(n8564), .A2(n8696), .ZN(n8695) );
  OR2_X1 U8601 ( .A1(n8563), .A2(n8562), .ZN(n8696) );
  NOR2_X1 U8602 ( .A1(n7462), .A2(n7645), .ZN(n8564) );
  NAND2_X1 U8603 ( .A1(n8562), .A2(n8563), .ZN(n8694) );
  NAND2_X1 U8604 ( .A1(n8697), .A2(n8698), .ZN(n8563) );
  NAND3_X1 U8605 ( .A1(a_18_), .A2(n8699), .A3(b_29_), .ZN(n8698) );
  NAND2_X1 U8606 ( .A1(n8559), .A2(n8558), .ZN(n8699) );
  OR2_X1 U8607 ( .A1(n8558), .A2(n8559), .ZN(n8697) );
  AND2_X1 U8608 ( .A1(n8700), .A2(n8701), .ZN(n8559) );
  NAND2_X1 U8609 ( .A1(n8556), .A2(n8702), .ZN(n8701) );
  OR2_X1 U8610 ( .A1(n8555), .A2(n8553), .ZN(n8702) );
  NOR2_X1 U8611 ( .A1(n7462), .A2(n7958), .ZN(n8556) );
  NAND2_X1 U8612 ( .A1(n8553), .A2(n8555), .ZN(n8700) );
  NAND2_X1 U8613 ( .A1(n8703), .A2(n8704), .ZN(n8555) );
  NAND3_X1 U8614 ( .A1(a_20_), .A2(n8705), .A3(b_29_), .ZN(n8704) );
  NAND2_X1 U8615 ( .A1(n8551), .A2(n8550), .ZN(n8705) );
  OR2_X1 U8616 ( .A1(n8550), .A2(n8551), .ZN(n8703) );
  AND2_X1 U8617 ( .A1(n8706), .A2(n8707), .ZN(n8551) );
  NAND2_X1 U8618 ( .A1(n8548), .A2(n8708), .ZN(n8707) );
  OR2_X1 U8619 ( .A1(n8547), .A2(n8546), .ZN(n8708) );
  NOR2_X1 U8620 ( .A1(n7462), .A2(n7578), .ZN(n8548) );
  NAND2_X1 U8621 ( .A1(n8546), .A2(n8547), .ZN(n8706) );
  NAND2_X1 U8622 ( .A1(n8709), .A2(n8710), .ZN(n8547) );
  NAND3_X1 U8623 ( .A1(a_22_), .A2(n8711), .A3(b_29_), .ZN(n8710) );
  OR2_X1 U8624 ( .A1(n8543), .A2(n8541), .ZN(n8711) );
  NAND2_X1 U8625 ( .A1(n8541), .A2(n8543), .ZN(n8709) );
  NAND2_X1 U8626 ( .A1(n8712), .A2(n8713), .ZN(n8543) );
  NAND2_X1 U8627 ( .A1(n8540), .A2(n8714), .ZN(n8713) );
  OR2_X1 U8628 ( .A1(n8539), .A2(n8537), .ZN(n8714) );
  NOR2_X1 U8629 ( .A1(n7462), .A2(n7955), .ZN(n8540) );
  NAND2_X1 U8630 ( .A1(n8537), .A2(n8539), .ZN(n8712) );
  NAND2_X1 U8631 ( .A1(n8715), .A2(n8716), .ZN(n8539) );
  NAND3_X1 U8632 ( .A1(a_24_), .A2(n8717), .A3(b_29_), .ZN(n8716) );
  OR2_X1 U8633 ( .A1(n8535), .A2(n8533), .ZN(n8717) );
  NAND2_X1 U8634 ( .A1(n8533), .A2(n8535), .ZN(n8715) );
  NAND2_X1 U8635 ( .A1(n8718), .A2(n8719), .ZN(n8535) );
  NAND2_X1 U8636 ( .A1(n8532), .A2(n8720), .ZN(n8719) );
  NAND2_X1 U8637 ( .A1(n8531), .A2(n8530), .ZN(n8720) );
  NOR2_X1 U8638 ( .A1(n7462), .A2(n7952), .ZN(n8532) );
  INV_X1 U8639 ( .A(b_29_), .ZN(n7462) );
  OR2_X1 U8640 ( .A1(n8530), .A2(n8531), .ZN(n8718) );
  AND2_X1 U8641 ( .A1(n8527), .A2(n8721), .ZN(n8531) );
  NAND2_X1 U8642 ( .A1(n8526), .A2(n8528), .ZN(n8721) );
  NAND2_X1 U8643 ( .A1(n8722), .A2(n8723), .ZN(n8528) );
  NAND2_X1 U8644 ( .A1(b_29_), .A2(a_26_), .ZN(n8723) );
  INV_X1 U8645 ( .A(n8724), .ZN(n8722) );
  XNOR2_X1 U8646 ( .A(n8725), .B(n8726), .ZN(n8526) );
  NAND2_X1 U8647 ( .A1(n8727), .A2(n8728), .ZN(n8725) );
  NAND2_X1 U8648 ( .A1(a_26_), .A2(n8724), .ZN(n8527) );
  NAND2_X1 U8649 ( .A1(n8500), .A2(n8729), .ZN(n8724) );
  NAND2_X1 U8650 ( .A1(n8499), .A2(n8501), .ZN(n8729) );
  NAND2_X1 U8651 ( .A1(n8730), .A2(n8731), .ZN(n8501) );
  NAND2_X1 U8652 ( .A1(b_29_), .A2(a_27_), .ZN(n8731) );
  INV_X1 U8653 ( .A(n8732), .ZN(n8730) );
  XOR2_X1 U8654 ( .A(n8733), .B(n8734), .Z(n8499) );
  XOR2_X1 U8655 ( .A(n7473), .B(n8735), .Z(n8733) );
  NAND2_X1 U8656 ( .A1(a_27_), .A2(n8732), .ZN(n8500) );
  NAND2_X1 U8657 ( .A1(n8736), .A2(n8737), .ZN(n8732) );
  NAND3_X1 U8658 ( .A1(a_28_), .A2(n8738), .A3(b_29_), .ZN(n8737) );
  NAND2_X1 U8659 ( .A1(n8509), .A2(n8507), .ZN(n8738) );
  OR2_X1 U8660 ( .A1(n8507), .A2(n8509), .ZN(n8736) );
  AND2_X1 U8661 ( .A1(n8739), .A2(n8740), .ZN(n8509) );
  NAND2_X1 U8662 ( .A1(n7457), .A2(n8741), .ZN(n8740) );
  OR2_X1 U8663 ( .A1(n8523), .A2(n8524), .ZN(n8741) );
  INV_X1 U8664 ( .A(n7942), .ZN(n7457) );
  NAND2_X1 U8665 ( .A1(b_29_), .A2(a_29_), .ZN(n7942) );
  NAND2_X1 U8666 ( .A1(n8524), .A2(n8523), .ZN(n8739) );
  NAND2_X1 U8667 ( .A1(n8742), .A2(n8743), .ZN(n8523) );
  NAND2_X1 U8668 ( .A1(b_27_), .A2(n8744), .ZN(n8743) );
  NAND2_X1 U8669 ( .A1(n7441), .A2(n8745), .ZN(n8744) );
  NAND2_X1 U8670 ( .A1(a_31_), .A2(n7949), .ZN(n8745) );
  NAND2_X1 U8671 ( .A1(b_28_), .A2(n8746), .ZN(n8742) );
  NAND2_X1 U8672 ( .A1(n7445), .A2(n8747), .ZN(n8746) );
  NAND2_X1 U8673 ( .A1(a_30_), .A2(n7494), .ZN(n8747) );
  AND3_X1 U8674 ( .A1(b_28_), .A2(n7409), .A3(b_29_), .ZN(n8524) );
  XNOR2_X1 U8675 ( .A(n8748), .B(n8749), .ZN(n8507) );
  XOR2_X1 U8676 ( .A(n8750), .B(n8751), .Z(n8748) );
  XOR2_X1 U8677 ( .A(n8752), .B(n8753), .Z(n8530) );
  NAND2_X1 U8678 ( .A1(n8754), .A2(n8755), .ZN(n8752) );
  XOR2_X1 U8679 ( .A(n8756), .B(n8757), .Z(n8533) );
  XOR2_X1 U8680 ( .A(n8758), .B(n8759), .Z(n8756) );
  XOR2_X1 U8681 ( .A(n8760), .B(n8761), .Z(n8537) );
  XOR2_X1 U8682 ( .A(n8762), .B(n8763), .Z(n8760) );
  NOR2_X1 U8683 ( .A1(n7954), .A2(n7949), .ZN(n8763) );
  XNOR2_X1 U8684 ( .A(n8764), .B(n8765), .ZN(n8541) );
  XNOR2_X1 U8685 ( .A(n8766), .B(n8767), .ZN(n8765) );
  XNOR2_X1 U8686 ( .A(n8768), .B(n8769), .ZN(n8546) );
  XNOR2_X1 U8687 ( .A(n8770), .B(n8771), .ZN(n8768) );
  NOR2_X1 U8688 ( .A1(n7568), .A2(n7949), .ZN(n8771) );
  XOR2_X1 U8689 ( .A(n8772), .B(n8773), .Z(n8550) );
  XNOR2_X1 U8690 ( .A(n8774), .B(n8775), .ZN(n8773) );
  XNOR2_X1 U8691 ( .A(n8776), .B(n8777), .ZN(n8553) );
  XNOR2_X1 U8692 ( .A(n8778), .B(n8779), .ZN(n8776) );
  NOR2_X1 U8693 ( .A1(n7957), .A2(n7949), .ZN(n8779) );
  XOR2_X1 U8694 ( .A(n8780), .B(n8781), .Z(n8558) );
  XNOR2_X1 U8695 ( .A(n8782), .B(n8783), .ZN(n8781) );
  XNOR2_X1 U8696 ( .A(n8784), .B(n8785), .ZN(n8562) );
  XNOR2_X1 U8697 ( .A(n8786), .B(n8787), .ZN(n8784) );
  NOR2_X1 U8698 ( .A1(n7960), .A2(n7949), .ZN(n8787) );
  XOR2_X1 U8699 ( .A(n8788), .B(n8789), .Z(n8565) );
  XOR2_X1 U8700 ( .A(n8790), .B(n8791), .Z(n8788) );
  XNOR2_X1 U8701 ( .A(n8792), .B(n8793), .ZN(n8569) );
  XOR2_X1 U8702 ( .A(n8794), .B(n8795), .Z(n8793) );
  NAND2_X1 U8703 ( .A1(b_28_), .A2(a_16_), .ZN(n8795) );
  XOR2_X1 U8704 ( .A(n8796), .B(n8797), .Z(n8574) );
  XNOR2_X1 U8705 ( .A(n8798), .B(n8799), .ZN(n8797) );
  XNOR2_X1 U8706 ( .A(n8800), .B(n8801), .ZN(n8577) );
  XNOR2_X1 U8707 ( .A(n8802), .B(n8803), .ZN(n8800) );
  NOR2_X1 U8708 ( .A1(n7962), .A2(n7949), .ZN(n8803) );
  XNOR2_X1 U8709 ( .A(n8804), .B(n8805), .ZN(n8582) );
  XOR2_X1 U8710 ( .A(n8806), .B(n8807), .Z(n8804) );
  XNOR2_X1 U8711 ( .A(n8808), .B(n8809), .ZN(n8586) );
  XOR2_X1 U8712 ( .A(n8810), .B(n8811), .Z(n8809) );
  NAND2_X1 U8713 ( .A1(b_28_), .A2(a_12_), .ZN(n8811) );
  XOR2_X1 U8714 ( .A(n8812), .B(n8813), .Z(n8591) );
  XNOR2_X1 U8715 ( .A(n8814), .B(n8815), .ZN(n8813) );
  XNOR2_X1 U8716 ( .A(n8816), .B(n8817), .ZN(n8595) );
  XOR2_X1 U8717 ( .A(n8818), .B(n8819), .Z(n8816) );
  NAND2_X1 U8718 ( .A1(b_28_), .A2(a_10_), .ZN(n8818) );
  XNOR2_X1 U8719 ( .A(n8820), .B(n8821), .ZN(n8599) );
  XNOR2_X1 U8720 ( .A(n8822), .B(n8823), .ZN(n8820) );
  XNOR2_X1 U8721 ( .A(n8824), .B(n8825), .ZN(n8603) );
  XNOR2_X1 U8722 ( .A(n8826), .B(n8827), .ZN(n8824) );
  NOR2_X1 U8723 ( .A1(n8602), .A2(n7949), .ZN(n8827) );
  XNOR2_X1 U8724 ( .A(n8828), .B(n8829), .ZN(n8608) );
  XNOR2_X1 U8725 ( .A(n8830), .B(n8831), .ZN(n8829) );
  XNOR2_X1 U8726 ( .A(n8832), .B(n8833), .ZN(n8612) );
  XNOR2_X1 U8727 ( .A(n8834), .B(n8835), .ZN(n8832) );
  NOR2_X1 U8728 ( .A1(n7807), .A2(n7949), .ZN(n8835) );
  XOR2_X1 U8729 ( .A(n8836), .B(n8837), .Z(n8616) );
  XNOR2_X1 U8730 ( .A(n8838), .B(n8839), .ZN(n8837) );
  XNOR2_X1 U8731 ( .A(n8840), .B(n8841), .ZN(n8619) );
  XNOR2_X1 U8732 ( .A(n8842), .B(n8843), .ZN(n8840) );
  NOR2_X1 U8733 ( .A1(n7836), .A2(n7949), .ZN(n8843) );
  OR2_X1 U8734 ( .A1(n8626), .A2(n8624), .ZN(n8649) );
  XOR2_X1 U8735 ( .A(n8844), .B(n8845), .Z(n8624) );
  XOR2_X1 U8736 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND2_X1 U8737 ( .A1(b_28_), .A2(a_3_), .ZN(n8847) );
  NAND2_X1 U8738 ( .A1(b_29_), .A2(a_2_), .ZN(n8626) );
  XNOR2_X1 U8739 ( .A(n8848), .B(n8849), .ZN(n8628) );
  XOR2_X1 U8740 ( .A(n8850), .B(n8851), .Z(n8848) );
  XOR2_X1 U8741 ( .A(n8852), .B(n8853), .Z(n8192) );
  XNOR2_X1 U8742 ( .A(n8854), .B(n8855), .ZN(n8852) );
  NOR2_X1 U8743 ( .A1(n8197), .A2(n7949), .ZN(n8855) );
  INV_X1 U8744 ( .A(n7997), .ZN(n8179) );
  NOR2_X1 U8745 ( .A1(n8182), .A2(n8181), .ZN(n7997) );
  OR2_X1 U8746 ( .A1(n8637), .A2(n8636), .ZN(n8181) );
  AND2_X1 U8747 ( .A1(n8856), .A2(n8857), .ZN(n8636) );
  NAND3_X1 U8748 ( .A1(a_0_), .A2(n8858), .A3(b_28_), .ZN(n8857) );
  NAND2_X1 U8749 ( .A1(n8854), .A2(n8853), .ZN(n8858) );
  OR2_X1 U8750 ( .A1(n8853), .A2(n8854), .ZN(n8856) );
  AND2_X1 U8751 ( .A1(n8859), .A2(n8860), .ZN(n8854) );
  NAND2_X1 U8752 ( .A1(n8645), .A2(n8861), .ZN(n8860) );
  OR2_X1 U8753 ( .A1(n8644), .A2(n8643), .ZN(n8861) );
  NOR2_X1 U8754 ( .A1(n7949), .A2(n7872), .ZN(n8645) );
  NAND2_X1 U8755 ( .A1(n8643), .A2(n8644), .ZN(n8859) );
  NAND2_X1 U8756 ( .A1(n8862), .A2(n8863), .ZN(n8644) );
  NAND2_X1 U8757 ( .A1(n8850), .A2(n8864), .ZN(n8863) );
  OR2_X1 U8758 ( .A1(n8849), .A2(n8851), .ZN(n8864) );
  NAND2_X1 U8759 ( .A1(n8865), .A2(n8866), .ZN(n8850) );
  NAND3_X1 U8760 ( .A1(a_3_), .A2(n8867), .A3(b_28_), .ZN(n8866) );
  OR2_X1 U8761 ( .A1(n8846), .A2(n8844), .ZN(n8867) );
  NAND2_X1 U8762 ( .A1(n8844), .A2(n8846), .ZN(n8865) );
  NAND2_X1 U8763 ( .A1(n8868), .A2(n8869), .ZN(n8846) );
  NAND3_X1 U8764 ( .A1(a_4_), .A2(n8870), .A3(b_28_), .ZN(n8869) );
  NAND2_X1 U8765 ( .A1(n8842), .A2(n8841), .ZN(n8870) );
  OR2_X1 U8766 ( .A1(n8841), .A2(n8842), .ZN(n8868) );
  AND2_X1 U8767 ( .A1(n8871), .A2(n8872), .ZN(n8842) );
  NAND2_X1 U8768 ( .A1(n8839), .A2(n8873), .ZN(n8872) );
  OR2_X1 U8769 ( .A1(n8838), .A2(n8836), .ZN(n8873) );
  NOR2_X1 U8770 ( .A1(n7949), .A2(n7823), .ZN(n8839) );
  NAND2_X1 U8771 ( .A1(n8836), .A2(n8838), .ZN(n8871) );
  NAND2_X1 U8772 ( .A1(n8874), .A2(n8875), .ZN(n8838) );
  NAND3_X1 U8773 ( .A1(a_6_), .A2(n8876), .A3(b_28_), .ZN(n8875) );
  NAND2_X1 U8774 ( .A1(n8834), .A2(n8833), .ZN(n8876) );
  OR2_X1 U8775 ( .A1(n8833), .A2(n8834), .ZN(n8874) );
  AND2_X1 U8776 ( .A1(n8877), .A2(n8878), .ZN(n8834) );
  NAND2_X1 U8777 ( .A1(n8831), .A2(n8879), .ZN(n8878) );
  OR2_X1 U8778 ( .A1(n8830), .A2(n8828), .ZN(n8879) );
  NOR2_X1 U8779 ( .A1(n7949), .A2(n7787), .ZN(n8831) );
  NAND2_X1 U8780 ( .A1(n8828), .A2(n8830), .ZN(n8877) );
  NAND2_X1 U8781 ( .A1(n8880), .A2(n8881), .ZN(n8830) );
  NAND3_X1 U8782 ( .A1(a_8_), .A2(n8882), .A3(b_28_), .ZN(n8881) );
  NAND2_X1 U8783 ( .A1(n8826), .A2(n8825), .ZN(n8882) );
  OR2_X1 U8784 ( .A1(n8825), .A2(n8826), .ZN(n8880) );
  AND2_X1 U8785 ( .A1(n8883), .A2(n8884), .ZN(n8826) );
  NAND2_X1 U8786 ( .A1(n8823), .A2(n8885), .ZN(n8884) );
  NAND2_X1 U8787 ( .A1(n8822), .A2(n8821), .ZN(n8885) );
  NOR2_X1 U8788 ( .A1(n7949), .A2(n7753), .ZN(n8823) );
  OR2_X1 U8789 ( .A1(n8821), .A2(n8822), .ZN(n8883) );
  AND2_X1 U8790 ( .A1(n8886), .A2(n8887), .ZN(n8822) );
  NAND3_X1 U8791 ( .A1(a_10_), .A2(n8888), .A3(b_28_), .ZN(n8887) );
  NAND2_X1 U8792 ( .A1(n8819), .A2(n8817), .ZN(n8888) );
  OR2_X1 U8793 ( .A1(n8817), .A2(n8819), .ZN(n8886) );
  AND2_X1 U8794 ( .A1(n8889), .A2(n8890), .ZN(n8819) );
  NAND2_X1 U8795 ( .A1(n8815), .A2(n8891), .ZN(n8890) );
  OR2_X1 U8796 ( .A1(n8814), .A2(n8812), .ZN(n8891) );
  NOR2_X1 U8797 ( .A1(n7949), .A2(n7724), .ZN(n8815) );
  NAND2_X1 U8798 ( .A1(n8812), .A2(n8814), .ZN(n8889) );
  NAND2_X1 U8799 ( .A1(n8892), .A2(n8893), .ZN(n8814) );
  NAND3_X1 U8800 ( .A1(a_12_), .A2(n8894), .A3(b_28_), .ZN(n8893) );
  OR2_X1 U8801 ( .A1(n8810), .A2(n8808), .ZN(n8894) );
  NAND2_X1 U8802 ( .A1(n8808), .A2(n8810), .ZN(n8892) );
  NAND2_X1 U8803 ( .A1(n8895), .A2(n8896), .ZN(n8810) );
  NAND2_X1 U8804 ( .A1(n8807), .A2(n8897), .ZN(n8896) );
  OR2_X1 U8805 ( .A1(n8806), .A2(n8805), .ZN(n8897) );
  NOR2_X1 U8806 ( .A1(n7949), .A2(n7702), .ZN(n8807) );
  NAND2_X1 U8807 ( .A1(n8805), .A2(n8806), .ZN(n8895) );
  NAND2_X1 U8808 ( .A1(n8898), .A2(n8899), .ZN(n8806) );
  NAND3_X1 U8809 ( .A1(a_14_), .A2(n8900), .A3(b_28_), .ZN(n8899) );
  NAND2_X1 U8810 ( .A1(n8802), .A2(n8801), .ZN(n8900) );
  OR2_X1 U8811 ( .A1(n8801), .A2(n8802), .ZN(n8898) );
  AND2_X1 U8812 ( .A1(n8901), .A2(n8902), .ZN(n8802) );
  NAND2_X1 U8813 ( .A1(n8799), .A2(n8903), .ZN(n8902) );
  OR2_X1 U8814 ( .A1(n8798), .A2(n8796), .ZN(n8903) );
  NOR2_X1 U8815 ( .A1(n7949), .A2(n7667), .ZN(n8799) );
  NAND2_X1 U8816 ( .A1(n8796), .A2(n8798), .ZN(n8901) );
  NAND2_X1 U8817 ( .A1(n8904), .A2(n8905), .ZN(n8798) );
  NAND3_X1 U8818 ( .A1(a_16_), .A2(n8906), .A3(b_28_), .ZN(n8905) );
  OR2_X1 U8819 ( .A1(n8794), .A2(n8792), .ZN(n8906) );
  NAND2_X1 U8820 ( .A1(n8792), .A2(n8794), .ZN(n8904) );
  NAND2_X1 U8821 ( .A1(n8907), .A2(n8908), .ZN(n8794) );
  NAND2_X1 U8822 ( .A1(n8791), .A2(n8909), .ZN(n8908) );
  OR2_X1 U8823 ( .A1(n8790), .A2(n8789), .ZN(n8909) );
  NOR2_X1 U8824 ( .A1(n7949), .A2(n7645), .ZN(n8791) );
  NAND2_X1 U8825 ( .A1(n8789), .A2(n8790), .ZN(n8907) );
  NAND2_X1 U8826 ( .A1(n8910), .A2(n8911), .ZN(n8790) );
  NAND3_X1 U8827 ( .A1(a_18_), .A2(n8912), .A3(b_28_), .ZN(n8911) );
  NAND2_X1 U8828 ( .A1(n8786), .A2(n8785), .ZN(n8912) );
  OR2_X1 U8829 ( .A1(n8785), .A2(n8786), .ZN(n8910) );
  AND2_X1 U8830 ( .A1(n8913), .A2(n8914), .ZN(n8786) );
  NAND2_X1 U8831 ( .A1(n8783), .A2(n8915), .ZN(n8914) );
  OR2_X1 U8832 ( .A1(n8782), .A2(n8780), .ZN(n8915) );
  NOR2_X1 U8833 ( .A1(n7949), .A2(n7958), .ZN(n8783) );
  NAND2_X1 U8834 ( .A1(n8780), .A2(n8782), .ZN(n8913) );
  NAND2_X1 U8835 ( .A1(n8916), .A2(n8917), .ZN(n8782) );
  NAND3_X1 U8836 ( .A1(a_20_), .A2(n8918), .A3(b_28_), .ZN(n8917) );
  NAND2_X1 U8837 ( .A1(n8778), .A2(n8777), .ZN(n8918) );
  OR2_X1 U8838 ( .A1(n8777), .A2(n8778), .ZN(n8916) );
  AND2_X1 U8839 ( .A1(n8919), .A2(n8920), .ZN(n8778) );
  NAND2_X1 U8840 ( .A1(n8775), .A2(n8921), .ZN(n8920) );
  OR2_X1 U8841 ( .A1(n8774), .A2(n8772), .ZN(n8921) );
  NOR2_X1 U8842 ( .A1(n7949), .A2(n7578), .ZN(n8775) );
  NAND2_X1 U8843 ( .A1(n8772), .A2(n8774), .ZN(n8919) );
  NAND2_X1 U8844 ( .A1(n8922), .A2(n8923), .ZN(n8774) );
  NAND3_X1 U8845 ( .A1(a_22_), .A2(n8924), .A3(b_28_), .ZN(n8923) );
  NAND2_X1 U8846 ( .A1(n8770), .A2(n8769), .ZN(n8924) );
  OR2_X1 U8847 ( .A1(n8769), .A2(n8770), .ZN(n8922) );
  AND2_X1 U8848 ( .A1(n8925), .A2(n8926), .ZN(n8770) );
  NAND2_X1 U8849 ( .A1(n8767), .A2(n8927), .ZN(n8926) );
  OR2_X1 U8850 ( .A1(n8766), .A2(n8764), .ZN(n8927) );
  NOR2_X1 U8851 ( .A1(n7949), .A2(n7955), .ZN(n8767) );
  NAND2_X1 U8852 ( .A1(n8764), .A2(n8766), .ZN(n8925) );
  NAND2_X1 U8853 ( .A1(n8928), .A2(n8929), .ZN(n8766) );
  NAND3_X1 U8854 ( .A1(a_24_), .A2(n8930), .A3(b_28_), .ZN(n8929) );
  OR2_X1 U8855 ( .A1(n8762), .A2(n8761), .ZN(n8930) );
  NAND2_X1 U8856 ( .A1(n8761), .A2(n8762), .ZN(n8928) );
  NAND2_X1 U8857 ( .A1(n8931), .A2(n8932), .ZN(n8762) );
  NAND2_X1 U8858 ( .A1(n8759), .A2(n8933), .ZN(n8932) );
  OR2_X1 U8859 ( .A1(n8758), .A2(n8757), .ZN(n8933) );
  NOR2_X1 U8860 ( .A1(n7949), .A2(n7952), .ZN(n8759) );
  NAND2_X1 U8861 ( .A1(n8757), .A2(n8758), .ZN(n8931) );
  NAND2_X1 U8862 ( .A1(n8754), .A2(n8934), .ZN(n8758) );
  NAND2_X1 U8863 ( .A1(n8753), .A2(n8755), .ZN(n8934) );
  NAND2_X1 U8864 ( .A1(n8935), .A2(n8936), .ZN(n8755) );
  NAND2_X1 U8865 ( .A1(b_28_), .A2(a_26_), .ZN(n8936) );
  INV_X1 U8866 ( .A(n8937), .ZN(n8935) );
  XOR2_X1 U8867 ( .A(n8938), .B(n8939), .Z(n8753) );
  XOR2_X1 U8868 ( .A(n8940), .B(n7492), .Z(n8938) );
  NAND2_X1 U8869 ( .A1(a_26_), .A2(n8937), .ZN(n8754) );
  NAND2_X1 U8870 ( .A1(n8727), .A2(n8941), .ZN(n8937) );
  NAND2_X1 U8871 ( .A1(n8726), .A2(n8728), .ZN(n8941) );
  NAND2_X1 U8872 ( .A1(n8942), .A2(n8943), .ZN(n8728) );
  NAND2_X1 U8873 ( .A1(b_28_), .A2(a_27_), .ZN(n8943) );
  INV_X1 U8874 ( .A(n8944), .ZN(n8942) );
  XNOR2_X1 U8875 ( .A(n8945), .B(n8946), .ZN(n8726) );
  XOR2_X1 U8876 ( .A(n8947), .B(n8948), .Z(n8945) );
  NAND2_X1 U8877 ( .A1(b_27_), .A2(a_28_), .ZN(n8947) );
  NAND2_X1 U8878 ( .A1(a_27_), .A2(n8944), .ZN(n8727) );
  NAND2_X1 U8879 ( .A1(n8949), .A2(n8950), .ZN(n8944) );
  NAND2_X1 U8880 ( .A1(n8734), .A2(n8951), .ZN(n8950) );
  NAND2_X1 U8881 ( .A1(n8735), .A2(n7473), .ZN(n8951) );
  INV_X1 U8882 ( .A(n8952), .ZN(n8735) );
  XOR2_X1 U8883 ( .A(n8953), .B(n8954), .Z(n8734) );
  XOR2_X1 U8884 ( .A(n8955), .B(n8956), .Z(n8953) );
  NAND2_X1 U8885 ( .A1(n8957), .A2(n8952), .ZN(n8949) );
  NAND2_X1 U8886 ( .A1(n8958), .A2(n8959), .ZN(n8952) );
  NAND2_X1 U8887 ( .A1(n8749), .A2(n8960), .ZN(n8959) );
  OR2_X1 U8888 ( .A1(n8750), .A2(n8751), .ZN(n8960) );
  NOR2_X1 U8889 ( .A1(n7949), .A2(n7460), .ZN(n8749) );
  NAND2_X1 U8890 ( .A1(n8751), .A2(n8750), .ZN(n8958) );
  NAND2_X1 U8891 ( .A1(n8961), .A2(n8962), .ZN(n8750) );
  NAND2_X1 U8892 ( .A1(b_26_), .A2(n8963), .ZN(n8962) );
  NAND2_X1 U8893 ( .A1(n7441), .A2(n8964), .ZN(n8963) );
  NAND2_X1 U8894 ( .A1(a_31_), .A2(n7494), .ZN(n8964) );
  NAND2_X1 U8895 ( .A1(b_27_), .A2(n8965), .ZN(n8961) );
  NAND2_X1 U8896 ( .A1(n7445), .A2(n8966), .ZN(n8965) );
  NAND2_X1 U8897 ( .A1(a_30_), .A2(n7951), .ZN(n8966) );
  AND3_X1 U8898 ( .A1(b_27_), .A2(n7409), .A3(b_28_), .ZN(n8751) );
  INV_X1 U8899 ( .A(n7473), .ZN(n8957) );
  NAND2_X1 U8900 ( .A1(b_28_), .A2(a_28_), .ZN(n7473) );
  XNOR2_X1 U8901 ( .A(n8967), .B(n8968), .ZN(n8757) );
  NAND2_X1 U8902 ( .A1(n8969), .A2(n8970), .ZN(n8967) );
  XNOR2_X1 U8903 ( .A(n8971), .B(n8972), .ZN(n8761) );
  XNOR2_X1 U8904 ( .A(n8973), .B(n8974), .ZN(n8971) );
  XNOR2_X1 U8905 ( .A(n8975), .B(n8976), .ZN(n8764) );
  XOR2_X1 U8906 ( .A(n8977), .B(n8978), .Z(n8976) );
  NAND2_X1 U8907 ( .A1(b_27_), .A2(a_24_), .ZN(n8978) );
  XOR2_X1 U8908 ( .A(n8979), .B(n8980), .Z(n8769) );
  XNOR2_X1 U8909 ( .A(n8981), .B(n8982), .ZN(n8980) );
  XNOR2_X1 U8910 ( .A(n8983), .B(n8984), .ZN(n8772) );
  XOR2_X1 U8911 ( .A(n8985), .B(n8986), .Z(n8984) );
  NAND2_X1 U8912 ( .A1(b_27_), .A2(a_22_), .ZN(n8986) );
  XNOR2_X1 U8913 ( .A(n8987), .B(n8988), .ZN(n8777) );
  XOR2_X1 U8914 ( .A(n8989), .B(n8990), .Z(n8987) );
  XNOR2_X1 U8915 ( .A(n8991), .B(n8992), .ZN(n8780) );
  XNOR2_X1 U8916 ( .A(n8993), .B(n8994), .ZN(n8991) );
  NOR2_X1 U8917 ( .A1(n7957), .A2(n7494), .ZN(n8994) );
  XOR2_X1 U8918 ( .A(n8995), .B(n8996), .Z(n8785) );
  XNOR2_X1 U8919 ( .A(n8997), .B(n8998), .ZN(n8996) );
  XNOR2_X1 U8920 ( .A(n8999), .B(n9000), .ZN(n8789) );
  XNOR2_X1 U8921 ( .A(n9001), .B(n9002), .ZN(n8999) );
  NOR2_X1 U8922 ( .A1(n7960), .A2(n7494), .ZN(n9002) );
  XNOR2_X1 U8923 ( .A(n9003), .B(n9004), .ZN(n8792) );
  XNOR2_X1 U8924 ( .A(n9005), .B(n9006), .ZN(n9004) );
  XNOR2_X1 U8925 ( .A(n9007), .B(n9008), .ZN(n8796) );
  XNOR2_X1 U8926 ( .A(n9009), .B(n9010), .ZN(n9007) );
  NOR2_X1 U8927 ( .A1(n8353), .A2(n7494), .ZN(n9010) );
  XOR2_X1 U8928 ( .A(n9011), .B(n9012), .Z(n8801) );
  XNOR2_X1 U8929 ( .A(n9013), .B(n9014), .ZN(n9012) );
  XNOR2_X1 U8930 ( .A(n9015), .B(n9016), .ZN(n8805) );
  XNOR2_X1 U8931 ( .A(n9017), .B(n9018), .ZN(n9015) );
  NOR2_X1 U8932 ( .A1(n7962), .A2(n7494), .ZN(n9018) );
  XNOR2_X1 U8933 ( .A(n9019), .B(n9020), .ZN(n8808) );
  XNOR2_X1 U8934 ( .A(n9021), .B(n9022), .ZN(n9019) );
  XNOR2_X1 U8935 ( .A(n9023), .B(n9024), .ZN(n8812) );
  XOR2_X1 U8936 ( .A(n9025), .B(n9026), .Z(n9024) );
  NAND2_X1 U8937 ( .A1(b_27_), .A2(a_12_), .ZN(n9026) );
  XOR2_X1 U8938 ( .A(n9027), .B(n9028), .Z(n8817) );
  XNOR2_X1 U8939 ( .A(n9029), .B(n9030), .ZN(n9028) );
  XNOR2_X1 U8940 ( .A(n9031), .B(n9032), .ZN(n8821) );
  XOR2_X1 U8941 ( .A(n9033), .B(n9034), .Z(n9031) );
  NOR2_X1 U8942 ( .A1(n8378), .A2(n7494), .ZN(n9034) );
  XNOR2_X1 U8943 ( .A(n9035), .B(n9036), .ZN(n8825) );
  XOR2_X1 U8944 ( .A(n9037), .B(n9038), .Z(n9035) );
  XOR2_X1 U8945 ( .A(n9039), .B(n9040), .Z(n8828) );
  XOR2_X1 U8946 ( .A(n9041), .B(n9042), .Z(n9039) );
  NOR2_X1 U8947 ( .A1(n8602), .A2(n7494), .ZN(n9042) );
  XOR2_X1 U8948 ( .A(n9043), .B(n9044), .Z(n8833) );
  XOR2_X1 U8949 ( .A(n9045), .B(n9046), .Z(n9044) );
  NAND2_X1 U8950 ( .A1(b_27_), .A2(a_7_), .ZN(n9046) );
  XNOR2_X1 U8951 ( .A(n9047), .B(n9048), .ZN(n8836) );
  XNOR2_X1 U8952 ( .A(n9049), .B(n9050), .ZN(n9047) );
  NOR2_X1 U8953 ( .A1(n7807), .A2(n7494), .ZN(n9050) );
  XOR2_X1 U8954 ( .A(n9051), .B(n9052), .Z(n8841) );
  XNOR2_X1 U8955 ( .A(n9053), .B(n9054), .ZN(n9052) );
  XNOR2_X1 U8956 ( .A(n9055), .B(n9056), .ZN(n8844) );
  XNOR2_X1 U8957 ( .A(n9057), .B(n9058), .ZN(n9055) );
  NOR2_X1 U8958 ( .A1(n7836), .A2(n7494), .ZN(n9058) );
  NAND2_X1 U8959 ( .A1(n8851), .A2(n8849), .ZN(n8862) );
  XNOR2_X1 U8960 ( .A(n9059), .B(n9060), .ZN(n8849) );
  NAND2_X1 U8961 ( .A1(n9061), .A2(n9062), .ZN(n9059) );
  NOR2_X1 U8962 ( .A1(n7949), .A2(n7966), .ZN(n8851) );
  XNOR2_X1 U8963 ( .A(n9063), .B(n9064), .ZN(n8643) );
  NAND2_X1 U8964 ( .A1(n9065), .A2(n9066), .ZN(n9063) );
  XNOR2_X1 U8965 ( .A(n9067), .B(n9068), .ZN(n8853) );
  XOR2_X1 U8966 ( .A(n9069), .B(n9070), .Z(n9067) );
  NOR2_X1 U8967 ( .A1(n7872), .A2(n7494), .ZN(n9070) );
  XNOR2_X1 U8968 ( .A(n9071), .B(n9072), .ZN(n8637) );
  XNOR2_X1 U8969 ( .A(n9073), .B(n9074), .ZN(n9072) );
  NAND2_X1 U8970 ( .A1(n9075), .A2(n8178), .ZN(n8182) );
  INV_X1 U8971 ( .A(n9076), .ZN(n8178) );
  NAND2_X1 U8972 ( .A1(n9077), .A2(n9078), .ZN(n9075) );
  NAND2_X1 U8973 ( .A1(n9076), .A2(n9079), .ZN(n8002) );
  XOR2_X1 U8974 ( .A(n8175), .B(n8174), .Z(n9079) );
  NOR2_X1 U8975 ( .A1(n9078), .A2(n9077), .ZN(n9076) );
  XOR2_X1 U8976 ( .A(n9080), .B(n9081), .Z(n9077) );
  XNOR2_X1 U8977 ( .A(n9082), .B(n9083), .ZN(n9080) );
  NOR2_X1 U8978 ( .A1(n8197), .A2(n7951), .ZN(n9083) );
  NAND2_X1 U8979 ( .A1(n9084), .A2(n9085), .ZN(n9078) );
  NAND2_X1 U8980 ( .A1(n9073), .A2(n9086), .ZN(n9085) );
  OR2_X1 U8981 ( .A1(n9074), .A2(n9071), .ZN(n9086) );
  AND2_X1 U8982 ( .A1(n9087), .A2(n9088), .ZN(n9073) );
  NAND3_X1 U8983 ( .A1(a_1_), .A2(n9089), .A3(b_27_), .ZN(n9088) );
  OR2_X1 U8984 ( .A1(n9069), .A2(n9068), .ZN(n9089) );
  NAND2_X1 U8985 ( .A1(n9068), .A2(n9069), .ZN(n9087) );
  NAND2_X1 U8986 ( .A1(n9065), .A2(n9090), .ZN(n9069) );
  NAND2_X1 U8987 ( .A1(n9064), .A2(n9066), .ZN(n9090) );
  NAND2_X1 U8988 ( .A1(n9091), .A2(n9092), .ZN(n9066) );
  NAND2_X1 U8989 ( .A1(b_27_), .A2(a_2_), .ZN(n9092) );
  INV_X1 U8990 ( .A(n9093), .ZN(n9091) );
  XNOR2_X1 U8991 ( .A(n9094), .B(n9095), .ZN(n9064) );
  XNOR2_X1 U8992 ( .A(n9096), .B(n9097), .ZN(n9094) );
  NOR2_X1 U8993 ( .A1(n7852), .A2(n7951), .ZN(n9097) );
  NAND2_X1 U8994 ( .A1(a_2_), .A2(n9093), .ZN(n9065) );
  NAND2_X1 U8995 ( .A1(n9061), .A2(n9098), .ZN(n9093) );
  NAND2_X1 U8996 ( .A1(n9060), .A2(n9062), .ZN(n9098) );
  NAND2_X1 U8997 ( .A1(n9099), .A2(n9100), .ZN(n9062) );
  NAND2_X1 U8998 ( .A1(b_27_), .A2(a_3_), .ZN(n9100) );
  INV_X1 U8999 ( .A(n9101), .ZN(n9099) );
  XNOR2_X1 U9000 ( .A(n9102), .B(n9103), .ZN(n9060) );
  XNOR2_X1 U9001 ( .A(n9104), .B(n9105), .ZN(n9103) );
  NAND2_X1 U9002 ( .A1(a_3_), .A2(n9101), .ZN(n9061) );
  NAND2_X1 U9003 ( .A1(n9106), .A2(n9107), .ZN(n9101) );
  NAND3_X1 U9004 ( .A1(a_4_), .A2(n9108), .A3(b_27_), .ZN(n9107) );
  NAND2_X1 U9005 ( .A1(n9057), .A2(n9056), .ZN(n9108) );
  OR2_X1 U9006 ( .A1(n9056), .A2(n9057), .ZN(n9106) );
  AND2_X1 U9007 ( .A1(n9109), .A2(n9110), .ZN(n9057) );
  NAND2_X1 U9008 ( .A1(n9054), .A2(n9111), .ZN(n9110) );
  OR2_X1 U9009 ( .A1(n9053), .A2(n9051), .ZN(n9111) );
  NOR2_X1 U9010 ( .A1(n7494), .A2(n7823), .ZN(n9054) );
  NAND2_X1 U9011 ( .A1(n9051), .A2(n9053), .ZN(n9109) );
  NAND2_X1 U9012 ( .A1(n9112), .A2(n9113), .ZN(n9053) );
  NAND3_X1 U9013 ( .A1(a_6_), .A2(n9114), .A3(b_27_), .ZN(n9113) );
  NAND2_X1 U9014 ( .A1(n9049), .A2(n9048), .ZN(n9114) );
  OR2_X1 U9015 ( .A1(n9048), .A2(n9049), .ZN(n9112) );
  AND2_X1 U9016 ( .A1(n9115), .A2(n9116), .ZN(n9049) );
  NAND3_X1 U9017 ( .A1(a_7_), .A2(n9117), .A3(b_27_), .ZN(n9116) );
  OR2_X1 U9018 ( .A1(n9045), .A2(n9043), .ZN(n9117) );
  NAND2_X1 U9019 ( .A1(n9043), .A2(n9045), .ZN(n9115) );
  NAND2_X1 U9020 ( .A1(n9118), .A2(n9119), .ZN(n9045) );
  NAND3_X1 U9021 ( .A1(a_8_), .A2(n9120), .A3(b_27_), .ZN(n9119) );
  OR2_X1 U9022 ( .A1(n9041), .A2(n9040), .ZN(n9120) );
  NAND2_X1 U9023 ( .A1(n9040), .A2(n9041), .ZN(n9118) );
  NAND2_X1 U9024 ( .A1(n9121), .A2(n9122), .ZN(n9041) );
  NAND2_X1 U9025 ( .A1(n9038), .A2(n9123), .ZN(n9122) );
  OR2_X1 U9026 ( .A1(n9037), .A2(n9036), .ZN(n9123) );
  NOR2_X1 U9027 ( .A1(n7494), .A2(n7753), .ZN(n9038) );
  NAND2_X1 U9028 ( .A1(n9036), .A2(n9037), .ZN(n9121) );
  NAND2_X1 U9029 ( .A1(n9124), .A2(n9125), .ZN(n9037) );
  NAND3_X1 U9030 ( .A1(a_10_), .A2(n9126), .A3(b_27_), .ZN(n9125) );
  OR2_X1 U9031 ( .A1(n9033), .A2(n9032), .ZN(n9126) );
  NAND2_X1 U9032 ( .A1(n9032), .A2(n9033), .ZN(n9124) );
  NAND2_X1 U9033 ( .A1(n9127), .A2(n9128), .ZN(n9033) );
  NAND2_X1 U9034 ( .A1(n9030), .A2(n9129), .ZN(n9128) );
  OR2_X1 U9035 ( .A1(n9029), .A2(n9027), .ZN(n9129) );
  NOR2_X1 U9036 ( .A1(n7494), .A2(n7724), .ZN(n9030) );
  NAND2_X1 U9037 ( .A1(n9027), .A2(n9029), .ZN(n9127) );
  NAND2_X1 U9038 ( .A1(n9130), .A2(n9131), .ZN(n9029) );
  NAND3_X1 U9039 ( .A1(a_12_), .A2(n9132), .A3(b_27_), .ZN(n9131) );
  OR2_X1 U9040 ( .A1(n9025), .A2(n9023), .ZN(n9132) );
  NAND2_X1 U9041 ( .A1(n9023), .A2(n9025), .ZN(n9130) );
  NAND2_X1 U9042 ( .A1(n9133), .A2(n9134), .ZN(n9025) );
  NAND2_X1 U9043 ( .A1(n9022), .A2(n9135), .ZN(n9134) );
  NAND2_X1 U9044 ( .A1(n9021), .A2(n9020), .ZN(n9135) );
  NOR2_X1 U9045 ( .A1(n7494), .A2(n7702), .ZN(n9022) );
  OR2_X1 U9046 ( .A1(n9020), .A2(n9021), .ZN(n9133) );
  AND2_X1 U9047 ( .A1(n9136), .A2(n9137), .ZN(n9021) );
  NAND3_X1 U9048 ( .A1(a_14_), .A2(n9138), .A3(b_27_), .ZN(n9137) );
  NAND2_X1 U9049 ( .A1(n9017), .A2(n9016), .ZN(n9138) );
  OR2_X1 U9050 ( .A1(n9016), .A2(n9017), .ZN(n9136) );
  AND2_X1 U9051 ( .A1(n9139), .A2(n9140), .ZN(n9017) );
  NAND2_X1 U9052 ( .A1(n9014), .A2(n9141), .ZN(n9140) );
  OR2_X1 U9053 ( .A1(n9013), .A2(n9011), .ZN(n9141) );
  NOR2_X1 U9054 ( .A1(n7494), .A2(n7667), .ZN(n9014) );
  NAND2_X1 U9055 ( .A1(n9011), .A2(n9013), .ZN(n9139) );
  NAND2_X1 U9056 ( .A1(n9142), .A2(n9143), .ZN(n9013) );
  NAND3_X1 U9057 ( .A1(a_16_), .A2(n9144), .A3(b_27_), .ZN(n9143) );
  NAND2_X1 U9058 ( .A1(n9009), .A2(n9008), .ZN(n9144) );
  OR2_X1 U9059 ( .A1(n9008), .A2(n9009), .ZN(n9142) );
  AND2_X1 U9060 ( .A1(n9145), .A2(n9146), .ZN(n9009) );
  NAND2_X1 U9061 ( .A1(n9006), .A2(n9147), .ZN(n9146) );
  OR2_X1 U9062 ( .A1(n9005), .A2(n9003), .ZN(n9147) );
  NOR2_X1 U9063 ( .A1(n7494), .A2(n7645), .ZN(n9006) );
  NAND2_X1 U9064 ( .A1(n9003), .A2(n9005), .ZN(n9145) );
  NAND2_X1 U9065 ( .A1(n9148), .A2(n9149), .ZN(n9005) );
  NAND3_X1 U9066 ( .A1(a_18_), .A2(n9150), .A3(b_27_), .ZN(n9149) );
  NAND2_X1 U9067 ( .A1(n9001), .A2(n9000), .ZN(n9150) );
  OR2_X1 U9068 ( .A1(n9000), .A2(n9001), .ZN(n9148) );
  AND2_X1 U9069 ( .A1(n9151), .A2(n9152), .ZN(n9001) );
  NAND2_X1 U9070 ( .A1(n8998), .A2(n9153), .ZN(n9152) );
  OR2_X1 U9071 ( .A1(n8997), .A2(n8995), .ZN(n9153) );
  NOR2_X1 U9072 ( .A1(n7494), .A2(n7958), .ZN(n8998) );
  NAND2_X1 U9073 ( .A1(n8995), .A2(n8997), .ZN(n9151) );
  NAND2_X1 U9074 ( .A1(n9154), .A2(n9155), .ZN(n8997) );
  NAND3_X1 U9075 ( .A1(a_20_), .A2(n9156), .A3(b_27_), .ZN(n9155) );
  NAND2_X1 U9076 ( .A1(n8993), .A2(n8992), .ZN(n9156) );
  OR2_X1 U9077 ( .A1(n8992), .A2(n8993), .ZN(n9154) );
  AND2_X1 U9078 ( .A1(n9157), .A2(n9158), .ZN(n8993) );
  NAND2_X1 U9079 ( .A1(n8990), .A2(n9159), .ZN(n9158) );
  OR2_X1 U9080 ( .A1(n8989), .A2(n8988), .ZN(n9159) );
  NOR2_X1 U9081 ( .A1(n7494), .A2(n7578), .ZN(n8990) );
  NAND2_X1 U9082 ( .A1(n8988), .A2(n8989), .ZN(n9157) );
  NAND2_X1 U9083 ( .A1(n9160), .A2(n9161), .ZN(n8989) );
  NAND3_X1 U9084 ( .A1(a_22_), .A2(n9162), .A3(b_27_), .ZN(n9161) );
  OR2_X1 U9085 ( .A1(n8985), .A2(n8983), .ZN(n9162) );
  NAND2_X1 U9086 ( .A1(n8983), .A2(n8985), .ZN(n9160) );
  NAND2_X1 U9087 ( .A1(n9163), .A2(n9164), .ZN(n8985) );
  NAND2_X1 U9088 ( .A1(n8982), .A2(n9165), .ZN(n9164) );
  OR2_X1 U9089 ( .A1(n8981), .A2(n8979), .ZN(n9165) );
  NOR2_X1 U9090 ( .A1(n7494), .A2(n7955), .ZN(n8982) );
  NAND2_X1 U9091 ( .A1(n8979), .A2(n8981), .ZN(n9163) );
  NAND2_X1 U9092 ( .A1(n9166), .A2(n9167), .ZN(n8981) );
  NAND3_X1 U9093 ( .A1(a_24_), .A2(n9168), .A3(b_27_), .ZN(n9167) );
  OR2_X1 U9094 ( .A1(n8977), .A2(n8975), .ZN(n9168) );
  NAND2_X1 U9095 ( .A1(n8975), .A2(n8977), .ZN(n9166) );
  NAND2_X1 U9096 ( .A1(n9169), .A2(n9170), .ZN(n8977) );
  NAND2_X1 U9097 ( .A1(n8974), .A2(n9171), .ZN(n9170) );
  NAND2_X1 U9098 ( .A1(n8973), .A2(n8972), .ZN(n9171) );
  NOR2_X1 U9099 ( .A1(n7494), .A2(n7952), .ZN(n8974) );
  OR2_X1 U9100 ( .A1(n8972), .A2(n8973), .ZN(n9169) );
  AND2_X1 U9101 ( .A1(n8969), .A2(n9172), .ZN(n8973) );
  NAND2_X1 U9102 ( .A1(n8968), .A2(n8970), .ZN(n9172) );
  NAND2_X1 U9103 ( .A1(n9173), .A2(n9174), .ZN(n8970) );
  NAND2_X1 U9104 ( .A1(b_27_), .A2(a_26_), .ZN(n9174) );
  INV_X1 U9105 ( .A(n9175), .ZN(n9173) );
  XNOR2_X1 U9106 ( .A(n9176), .B(n9177), .ZN(n8968) );
  NAND2_X1 U9107 ( .A1(n9178), .A2(n9179), .ZN(n9176) );
  NAND2_X1 U9108 ( .A1(a_26_), .A2(n9175), .ZN(n8969) );
  NAND2_X1 U9109 ( .A1(n9180), .A2(n9181), .ZN(n9175) );
  NAND2_X1 U9110 ( .A1(n8939), .A2(n9182), .ZN(n9181) );
  OR2_X1 U9111 ( .A1(n8940), .A2(n7492), .ZN(n9182) );
  XNOR2_X1 U9112 ( .A(n9183), .B(n9184), .ZN(n8939) );
  XOR2_X1 U9113 ( .A(n9185), .B(n9186), .Z(n9183) );
  NAND2_X1 U9114 ( .A1(b_26_), .A2(a_28_), .ZN(n9185) );
  NAND2_X1 U9115 ( .A1(n7492), .A2(n8940), .ZN(n9180) );
  NAND2_X1 U9116 ( .A1(n9187), .A2(n9188), .ZN(n8940) );
  NAND3_X1 U9117 ( .A1(a_28_), .A2(n9189), .A3(b_27_), .ZN(n9188) );
  NAND2_X1 U9118 ( .A1(n8948), .A2(n8946), .ZN(n9189) );
  OR2_X1 U9119 ( .A1(n8946), .A2(n8948), .ZN(n9187) );
  AND2_X1 U9120 ( .A1(n9190), .A2(n9191), .ZN(n8948) );
  NAND2_X1 U9121 ( .A1(n8954), .A2(n9192), .ZN(n9191) );
  OR2_X1 U9122 ( .A1(n8955), .A2(n8956), .ZN(n9192) );
  NOR2_X1 U9123 ( .A1(n7494), .A2(n7460), .ZN(n8954) );
  INV_X1 U9124 ( .A(b_27_), .ZN(n7494) );
  NAND2_X1 U9125 ( .A1(n8956), .A2(n8955), .ZN(n9190) );
  NAND2_X1 U9126 ( .A1(n9193), .A2(n9194), .ZN(n8955) );
  NAND2_X1 U9127 ( .A1(b_25_), .A2(n9195), .ZN(n9194) );
  NAND2_X1 U9128 ( .A1(n7441), .A2(n9196), .ZN(n9195) );
  NAND2_X1 U9129 ( .A1(a_31_), .A2(n7951), .ZN(n9196) );
  NAND2_X1 U9130 ( .A1(b_26_), .A2(n9197), .ZN(n9193) );
  NAND2_X1 U9131 ( .A1(n7445), .A2(n9198), .ZN(n9197) );
  NAND2_X1 U9132 ( .A1(a_30_), .A2(n7522), .ZN(n9198) );
  AND3_X1 U9133 ( .A1(b_26_), .A2(n7409), .A3(b_27_), .ZN(n8956) );
  XNOR2_X1 U9134 ( .A(n9199), .B(n9200), .ZN(n8946) );
  XOR2_X1 U9135 ( .A(n9201), .B(n9202), .Z(n9199) );
  INV_X1 U9136 ( .A(n7938), .ZN(n7492) );
  NAND2_X1 U9137 ( .A1(b_27_), .A2(a_27_), .ZN(n7938) );
  XNOR2_X1 U9138 ( .A(n9203), .B(n9204), .ZN(n8972) );
  XOR2_X1 U9139 ( .A(n9205), .B(n9206), .Z(n9203) );
  XOR2_X1 U9140 ( .A(n9207), .B(n9208), .Z(n8975) );
  XOR2_X1 U9141 ( .A(n9209), .B(n9210), .Z(n9207) );
  XNOR2_X1 U9142 ( .A(n9211), .B(n9212), .ZN(n8979) );
  XNOR2_X1 U9143 ( .A(n9213), .B(n9214), .ZN(n9211) );
  NOR2_X1 U9144 ( .A1(n7954), .A2(n7951), .ZN(n9214) );
  XNOR2_X1 U9145 ( .A(n9215), .B(n9216), .ZN(n8983) );
  XNOR2_X1 U9146 ( .A(n9217), .B(n9218), .ZN(n9216) );
  XNOR2_X1 U9147 ( .A(n9219), .B(n9220), .ZN(n8988) );
  XOR2_X1 U9148 ( .A(n9221), .B(n9222), .Z(n9220) );
  NAND2_X1 U9149 ( .A1(b_26_), .A2(a_22_), .ZN(n9222) );
  XNOR2_X1 U9150 ( .A(n9223), .B(n9224), .ZN(n8992) );
  XOR2_X1 U9151 ( .A(n9225), .B(n9226), .Z(n9223) );
  XNOR2_X1 U9152 ( .A(n9227), .B(n9228), .ZN(n8995) );
  XNOR2_X1 U9153 ( .A(n9229), .B(n9230), .ZN(n9227) );
  NOR2_X1 U9154 ( .A1(n7957), .A2(n7951), .ZN(n9230) );
  XOR2_X1 U9155 ( .A(n9231), .B(n9232), .Z(n9000) );
  XNOR2_X1 U9156 ( .A(n9233), .B(n9234), .ZN(n9232) );
  XNOR2_X1 U9157 ( .A(n9235), .B(n9236), .ZN(n9003) );
  XNOR2_X1 U9158 ( .A(n9237), .B(n9238), .ZN(n9235) );
  NOR2_X1 U9159 ( .A1(n7960), .A2(n7951), .ZN(n9238) );
  XNOR2_X1 U9160 ( .A(n9239), .B(n9240), .ZN(n9008) );
  XOR2_X1 U9161 ( .A(n9241), .B(n9242), .Z(n9239) );
  XNOR2_X1 U9162 ( .A(n9243), .B(n9244), .ZN(n9011) );
  XOR2_X1 U9163 ( .A(n9245), .B(n9246), .Z(n9244) );
  NAND2_X1 U9164 ( .A1(b_26_), .A2(a_16_), .ZN(n9246) );
  XOR2_X1 U9165 ( .A(n9247), .B(n9248), .Z(n9016) );
  XNOR2_X1 U9166 ( .A(n9249), .B(n9250), .ZN(n9248) );
  XNOR2_X1 U9167 ( .A(n9251), .B(n9252), .ZN(n9020) );
  XOR2_X1 U9168 ( .A(n9253), .B(n9254), .Z(n9251) );
  NOR2_X1 U9169 ( .A1(n7962), .A2(n7951), .ZN(n9254) );
  XOR2_X1 U9170 ( .A(n9255), .B(n9256), .Z(n9023) );
  XOR2_X1 U9171 ( .A(n9257), .B(n9258), .Z(n9255) );
  XNOR2_X1 U9172 ( .A(n9259), .B(n9260), .ZN(n9027) );
  XNOR2_X1 U9173 ( .A(n9261), .B(n9262), .ZN(n9259) );
  NOR2_X1 U9174 ( .A1(n8585), .A2(n7951), .ZN(n9262) );
  XNOR2_X1 U9175 ( .A(n9263), .B(n9264), .ZN(n9032) );
  XNOR2_X1 U9176 ( .A(n9265), .B(n9266), .ZN(n9264) );
  XNOR2_X1 U9177 ( .A(n9267), .B(n9268), .ZN(n9036) );
  XNOR2_X1 U9178 ( .A(n9269), .B(n9270), .ZN(n9267) );
  NOR2_X1 U9179 ( .A1(n8378), .A2(n7951), .ZN(n9270) );
  XNOR2_X1 U9180 ( .A(n9271), .B(n9272), .ZN(n9040) );
  XNOR2_X1 U9181 ( .A(n9273), .B(n9274), .ZN(n9271) );
  XNOR2_X1 U9182 ( .A(n9275), .B(n9276), .ZN(n9043) );
  XOR2_X1 U9183 ( .A(n9277), .B(n9278), .Z(n9276) );
  NAND2_X1 U9184 ( .A1(b_26_), .A2(a_8_), .ZN(n9278) );
  XOR2_X1 U9185 ( .A(n9279), .B(n9280), .Z(n9048) );
  NAND2_X1 U9186 ( .A1(n9281), .A2(n9282), .ZN(n9279) );
  XNOR2_X1 U9187 ( .A(n9283), .B(n9284), .ZN(n9051) );
  XOR2_X1 U9188 ( .A(n9285), .B(n9286), .Z(n9283) );
  NAND2_X1 U9189 ( .A1(b_26_), .A2(a_6_), .ZN(n9285) );
  XOR2_X1 U9190 ( .A(n9287), .B(n9288), .Z(n9056) );
  XOR2_X1 U9191 ( .A(n9289), .B(n9290), .Z(n9288) );
  NAND2_X1 U9192 ( .A1(b_26_), .A2(a_5_), .ZN(n9290) );
  XNOR2_X1 U9193 ( .A(n9291), .B(n9292), .ZN(n9068) );
  XNOR2_X1 U9194 ( .A(n9293), .B(n9294), .ZN(n9292) );
  NAND2_X1 U9195 ( .A1(n9071), .A2(n9074), .ZN(n9084) );
  NAND2_X1 U9196 ( .A1(b_27_), .A2(a_0_), .ZN(n9074) );
  XOR2_X1 U9197 ( .A(n9295), .B(n9296), .Z(n9071) );
  XNOR2_X1 U9198 ( .A(n9297), .B(n9298), .ZN(n9295) );
  NAND4_X1 U9199 ( .A1(n8174), .A2(n8173), .A3(n8175), .A4(n8168), .ZN(n8007)
         );
  INV_X1 U9200 ( .A(n9299), .ZN(n8168) );
  NAND2_X1 U9201 ( .A1(n9300), .A2(n9301), .ZN(n8175) );
  NAND3_X1 U9202 ( .A1(a_0_), .A2(n9302), .A3(b_26_), .ZN(n9301) );
  NAND2_X1 U9203 ( .A1(n9082), .A2(n9081), .ZN(n9302) );
  OR2_X1 U9204 ( .A1(n9081), .A2(n9082), .ZN(n9300) );
  AND2_X1 U9205 ( .A1(n9303), .A2(n9304), .ZN(n9082) );
  NAND2_X1 U9206 ( .A1(n9298), .A2(n9305), .ZN(n9304) );
  NAND2_X1 U9207 ( .A1(n9297), .A2(n9296), .ZN(n9305) );
  NOR2_X1 U9208 ( .A1(n7951), .A2(n7872), .ZN(n9298) );
  OR2_X1 U9209 ( .A1(n9296), .A2(n9297), .ZN(n9303) );
  AND2_X1 U9210 ( .A1(n9306), .A2(n9307), .ZN(n9297) );
  NAND2_X1 U9211 ( .A1(n9294), .A2(n9308), .ZN(n9307) );
  OR2_X1 U9212 ( .A1(n9293), .A2(n9291), .ZN(n9308) );
  NOR2_X1 U9213 ( .A1(n7951), .A2(n7966), .ZN(n9294) );
  NAND2_X1 U9214 ( .A1(n9291), .A2(n9293), .ZN(n9306) );
  NAND2_X1 U9215 ( .A1(n9309), .A2(n9310), .ZN(n9293) );
  NAND3_X1 U9216 ( .A1(a_3_), .A2(n9311), .A3(b_26_), .ZN(n9310) );
  NAND2_X1 U9217 ( .A1(n9096), .A2(n9095), .ZN(n9311) );
  OR2_X1 U9218 ( .A1(n9095), .A2(n9096), .ZN(n9309) );
  AND2_X1 U9219 ( .A1(n9312), .A2(n9313), .ZN(n9096) );
  NAND2_X1 U9220 ( .A1(n9105), .A2(n9314), .ZN(n9313) );
  OR2_X1 U9221 ( .A1(n9104), .A2(n9102), .ZN(n9314) );
  NOR2_X1 U9222 ( .A1(n7951), .A2(n7836), .ZN(n9105) );
  NAND2_X1 U9223 ( .A1(n9102), .A2(n9104), .ZN(n9312) );
  NAND2_X1 U9224 ( .A1(n9315), .A2(n9316), .ZN(n9104) );
  NAND3_X1 U9225 ( .A1(a_5_), .A2(n9317), .A3(b_26_), .ZN(n9316) );
  OR2_X1 U9226 ( .A1(n9289), .A2(n9287), .ZN(n9317) );
  NAND2_X1 U9227 ( .A1(n9287), .A2(n9289), .ZN(n9315) );
  NAND2_X1 U9228 ( .A1(n9318), .A2(n9319), .ZN(n9289) );
  NAND3_X1 U9229 ( .A1(a_6_), .A2(n9320), .A3(b_26_), .ZN(n9319) );
  NAND2_X1 U9230 ( .A1(n9286), .A2(n9284), .ZN(n9320) );
  OR2_X1 U9231 ( .A1(n9284), .A2(n9286), .ZN(n9318) );
  AND2_X1 U9232 ( .A1(n9281), .A2(n9321), .ZN(n9286) );
  NAND2_X1 U9233 ( .A1(n9280), .A2(n9282), .ZN(n9321) );
  NAND2_X1 U9234 ( .A1(n9322), .A2(n9323), .ZN(n9282) );
  NAND2_X1 U9235 ( .A1(b_26_), .A2(a_7_), .ZN(n9323) );
  INV_X1 U9236 ( .A(n9324), .ZN(n9322) );
  XOR2_X1 U9237 ( .A(n9325), .B(n9326), .Z(n9280) );
  XOR2_X1 U9238 ( .A(n9327), .B(n9328), .Z(n9325) );
  NOR2_X1 U9239 ( .A1(n8602), .A2(n7522), .ZN(n9328) );
  NAND2_X1 U9240 ( .A1(a_7_), .A2(n9324), .ZN(n9281) );
  NAND2_X1 U9241 ( .A1(n9329), .A2(n9330), .ZN(n9324) );
  NAND3_X1 U9242 ( .A1(a_8_), .A2(n9331), .A3(b_26_), .ZN(n9330) );
  OR2_X1 U9243 ( .A1(n9277), .A2(n9275), .ZN(n9331) );
  NAND2_X1 U9244 ( .A1(n9275), .A2(n9277), .ZN(n9329) );
  NAND2_X1 U9245 ( .A1(n9332), .A2(n9333), .ZN(n9277) );
  NAND2_X1 U9246 ( .A1(n9274), .A2(n9334), .ZN(n9333) );
  NAND2_X1 U9247 ( .A1(n9273), .A2(n9272), .ZN(n9334) );
  NOR2_X1 U9248 ( .A1(n7951), .A2(n7753), .ZN(n9274) );
  OR2_X1 U9249 ( .A1(n9272), .A2(n9273), .ZN(n9332) );
  AND2_X1 U9250 ( .A1(n9335), .A2(n9336), .ZN(n9273) );
  NAND3_X1 U9251 ( .A1(a_10_), .A2(n9337), .A3(b_26_), .ZN(n9336) );
  NAND2_X1 U9252 ( .A1(n9269), .A2(n9268), .ZN(n9337) );
  OR2_X1 U9253 ( .A1(n9268), .A2(n9269), .ZN(n9335) );
  AND2_X1 U9254 ( .A1(n9338), .A2(n9339), .ZN(n9269) );
  NAND2_X1 U9255 ( .A1(n9266), .A2(n9340), .ZN(n9339) );
  OR2_X1 U9256 ( .A1(n9265), .A2(n9263), .ZN(n9340) );
  NOR2_X1 U9257 ( .A1(n7951), .A2(n7724), .ZN(n9266) );
  NAND2_X1 U9258 ( .A1(n9263), .A2(n9265), .ZN(n9338) );
  NAND2_X1 U9259 ( .A1(n9341), .A2(n9342), .ZN(n9265) );
  NAND3_X1 U9260 ( .A1(a_12_), .A2(n9343), .A3(b_26_), .ZN(n9342) );
  NAND2_X1 U9261 ( .A1(n9261), .A2(n9260), .ZN(n9343) );
  OR2_X1 U9262 ( .A1(n9260), .A2(n9261), .ZN(n9341) );
  AND2_X1 U9263 ( .A1(n9344), .A2(n9345), .ZN(n9261) );
  NAND2_X1 U9264 ( .A1(n9258), .A2(n9346), .ZN(n9345) );
  OR2_X1 U9265 ( .A1(n9257), .A2(n9256), .ZN(n9346) );
  NOR2_X1 U9266 ( .A1(n7951), .A2(n7702), .ZN(n9258) );
  NAND2_X1 U9267 ( .A1(n9256), .A2(n9257), .ZN(n9344) );
  NAND2_X1 U9268 ( .A1(n9347), .A2(n9348), .ZN(n9257) );
  NAND3_X1 U9269 ( .A1(a_14_), .A2(n9349), .A3(b_26_), .ZN(n9348) );
  OR2_X1 U9270 ( .A1(n9253), .A2(n9252), .ZN(n9349) );
  NAND2_X1 U9271 ( .A1(n9252), .A2(n9253), .ZN(n9347) );
  NAND2_X1 U9272 ( .A1(n9350), .A2(n9351), .ZN(n9253) );
  NAND2_X1 U9273 ( .A1(n9250), .A2(n9352), .ZN(n9351) );
  OR2_X1 U9274 ( .A1(n9249), .A2(n9247), .ZN(n9352) );
  NOR2_X1 U9275 ( .A1(n7951), .A2(n7667), .ZN(n9250) );
  NAND2_X1 U9276 ( .A1(n9247), .A2(n9249), .ZN(n9350) );
  NAND2_X1 U9277 ( .A1(n9353), .A2(n9354), .ZN(n9249) );
  NAND3_X1 U9278 ( .A1(a_16_), .A2(n9355), .A3(b_26_), .ZN(n9354) );
  OR2_X1 U9279 ( .A1(n9245), .A2(n9243), .ZN(n9355) );
  NAND2_X1 U9280 ( .A1(n9243), .A2(n9245), .ZN(n9353) );
  NAND2_X1 U9281 ( .A1(n9356), .A2(n9357), .ZN(n9245) );
  NAND2_X1 U9282 ( .A1(n9242), .A2(n9358), .ZN(n9357) );
  OR2_X1 U9283 ( .A1(n9241), .A2(n9240), .ZN(n9358) );
  NOR2_X1 U9284 ( .A1(n7951), .A2(n7645), .ZN(n9242) );
  NAND2_X1 U9285 ( .A1(n9240), .A2(n9241), .ZN(n9356) );
  NAND2_X1 U9286 ( .A1(n9359), .A2(n9360), .ZN(n9241) );
  NAND3_X1 U9287 ( .A1(a_18_), .A2(n9361), .A3(b_26_), .ZN(n9360) );
  NAND2_X1 U9288 ( .A1(n9237), .A2(n9236), .ZN(n9361) );
  OR2_X1 U9289 ( .A1(n9236), .A2(n9237), .ZN(n9359) );
  AND2_X1 U9290 ( .A1(n9362), .A2(n9363), .ZN(n9237) );
  NAND2_X1 U9291 ( .A1(n9234), .A2(n9364), .ZN(n9363) );
  OR2_X1 U9292 ( .A1(n9233), .A2(n9231), .ZN(n9364) );
  NOR2_X1 U9293 ( .A1(n7951), .A2(n7958), .ZN(n9234) );
  NAND2_X1 U9294 ( .A1(n9231), .A2(n9233), .ZN(n9362) );
  NAND2_X1 U9295 ( .A1(n9365), .A2(n9366), .ZN(n9233) );
  NAND3_X1 U9296 ( .A1(a_20_), .A2(n9367), .A3(b_26_), .ZN(n9366) );
  NAND2_X1 U9297 ( .A1(n9229), .A2(n9228), .ZN(n9367) );
  OR2_X1 U9298 ( .A1(n9228), .A2(n9229), .ZN(n9365) );
  AND2_X1 U9299 ( .A1(n9368), .A2(n9369), .ZN(n9229) );
  NAND2_X1 U9300 ( .A1(n9226), .A2(n9370), .ZN(n9369) );
  OR2_X1 U9301 ( .A1(n9225), .A2(n9224), .ZN(n9370) );
  NOR2_X1 U9302 ( .A1(n7951), .A2(n7578), .ZN(n9226) );
  NAND2_X1 U9303 ( .A1(n9224), .A2(n9225), .ZN(n9368) );
  NAND2_X1 U9304 ( .A1(n9371), .A2(n9372), .ZN(n9225) );
  NAND3_X1 U9305 ( .A1(a_22_), .A2(n9373), .A3(b_26_), .ZN(n9372) );
  OR2_X1 U9306 ( .A1(n9221), .A2(n9219), .ZN(n9373) );
  NAND2_X1 U9307 ( .A1(n9219), .A2(n9221), .ZN(n9371) );
  NAND2_X1 U9308 ( .A1(n9374), .A2(n9375), .ZN(n9221) );
  NAND2_X1 U9309 ( .A1(n9218), .A2(n9376), .ZN(n9375) );
  OR2_X1 U9310 ( .A1(n9217), .A2(n9215), .ZN(n9376) );
  NOR2_X1 U9311 ( .A1(n7951), .A2(n7955), .ZN(n9218) );
  NAND2_X1 U9312 ( .A1(n9215), .A2(n9217), .ZN(n9374) );
  NAND2_X1 U9313 ( .A1(n9377), .A2(n9378), .ZN(n9217) );
  NAND3_X1 U9314 ( .A1(a_24_), .A2(n9379), .A3(b_26_), .ZN(n9378) );
  NAND2_X1 U9315 ( .A1(n9213), .A2(n9212), .ZN(n9379) );
  OR2_X1 U9316 ( .A1(n9212), .A2(n9213), .ZN(n9377) );
  AND2_X1 U9317 ( .A1(n9380), .A2(n9381), .ZN(n9213) );
  NAND2_X1 U9318 ( .A1(n9210), .A2(n9382), .ZN(n9381) );
  OR2_X1 U9319 ( .A1(n9209), .A2(n9208), .ZN(n9382) );
  NOR2_X1 U9320 ( .A1(n7951), .A2(n7952), .ZN(n9210) );
  NAND2_X1 U9321 ( .A1(n9208), .A2(n9209), .ZN(n9380) );
  NAND2_X1 U9322 ( .A1(n9383), .A2(n9384), .ZN(n9209) );
  NAND2_X1 U9323 ( .A1(n9204), .A2(n9385), .ZN(n9384) );
  OR2_X1 U9324 ( .A1(n9205), .A2(n9206), .ZN(n9385) );
  XNOR2_X1 U9325 ( .A(n9386), .B(n9387), .ZN(n9204) );
  NAND2_X1 U9326 ( .A1(n9388), .A2(n9389), .ZN(n9386) );
  NAND2_X1 U9327 ( .A1(n9206), .A2(n9205), .ZN(n9383) );
  NAND2_X1 U9328 ( .A1(n9178), .A2(n9390), .ZN(n9205) );
  NAND2_X1 U9329 ( .A1(n9177), .A2(n9179), .ZN(n9390) );
  NAND2_X1 U9330 ( .A1(n9391), .A2(n9392), .ZN(n9179) );
  NAND2_X1 U9331 ( .A1(b_26_), .A2(a_27_), .ZN(n9392) );
  INV_X1 U9332 ( .A(n9393), .ZN(n9391) );
  XNOR2_X1 U9333 ( .A(n9394), .B(n9395), .ZN(n9177) );
  XOR2_X1 U9334 ( .A(n9396), .B(n9397), .Z(n9394) );
  NAND2_X1 U9335 ( .A1(b_25_), .A2(a_28_), .ZN(n9396) );
  NAND2_X1 U9336 ( .A1(a_27_), .A2(n9393), .ZN(n9178) );
  NAND2_X1 U9337 ( .A1(n9398), .A2(n9399), .ZN(n9393) );
  NAND3_X1 U9338 ( .A1(a_28_), .A2(n9400), .A3(b_26_), .ZN(n9399) );
  NAND2_X1 U9339 ( .A1(n9186), .A2(n9184), .ZN(n9400) );
  OR2_X1 U9340 ( .A1(n9184), .A2(n9186), .ZN(n9398) );
  AND2_X1 U9341 ( .A1(n9401), .A2(n9402), .ZN(n9186) );
  NAND2_X1 U9342 ( .A1(n9200), .A2(n9403), .ZN(n9402) );
  OR2_X1 U9343 ( .A1(n9201), .A2(n9202), .ZN(n9403) );
  NOR2_X1 U9344 ( .A1(n7951), .A2(n7460), .ZN(n9200) );
  INV_X1 U9345 ( .A(b_26_), .ZN(n7951) );
  NAND2_X1 U9346 ( .A1(n9202), .A2(n9201), .ZN(n9401) );
  NAND2_X1 U9347 ( .A1(n9404), .A2(n9405), .ZN(n9201) );
  NAND2_X1 U9348 ( .A1(b_24_), .A2(n9406), .ZN(n9405) );
  NAND2_X1 U9349 ( .A1(n7441), .A2(n9407), .ZN(n9406) );
  NAND2_X1 U9350 ( .A1(a_31_), .A2(n7522), .ZN(n9407) );
  NAND2_X1 U9351 ( .A1(b_25_), .A2(n9408), .ZN(n9404) );
  NAND2_X1 U9352 ( .A1(n7445), .A2(n9409), .ZN(n9408) );
  NAND2_X1 U9353 ( .A1(a_30_), .A2(n7953), .ZN(n9409) );
  AND3_X1 U9354 ( .A1(b_25_), .A2(n7409), .A3(b_26_), .ZN(n9202) );
  XNOR2_X1 U9355 ( .A(n9410), .B(n9411), .ZN(n9184) );
  XOR2_X1 U9356 ( .A(n9412), .B(n9413), .Z(n9410) );
  INV_X1 U9357 ( .A(n7507), .ZN(n9206) );
  NAND2_X1 U9358 ( .A1(b_26_), .A2(a_26_), .ZN(n7507) );
  XNOR2_X1 U9359 ( .A(n9414), .B(n9415), .ZN(n9208) );
  NAND2_X1 U9360 ( .A1(n9416), .A2(n9417), .ZN(n9414) );
  XNOR2_X1 U9361 ( .A(n9418), .B(n9419), .ZN(n9212) );
  XOR2_X1 U9362 ( .A(n9420), .B(n7520), .Z(n9418) );
  XNOR2_X1 U9363 ( .A(n9421), .B(n9422), .ZN(n9215) );
  XNOR2_X1 U9364 ( .A(n9423), .B(n9424), .ZN(n9421) );
  NOR2_X1 U9365 ( .A1(n7954), .A2(n7522), .ZN(n9424) );
  XNOR2_X1 U9366 ( .A(n9425), .B(n9426), .ZN(n9219) );
  XNOR2_X1 U9367 ( .A(n9427), .B(n9428), .ZN(n9426) );
  XNOR2_X1 U9368 ( .A(n9429), .B(n9430), .ZN(n9224) );
  XOR2_X1 U9369 ( .A(n9431), .B(n9432), .Z(n9430) );
  NAND2_X1 U9370 ( .A1(b_25_), .A2(a_22_), .ZN(n9432) );
  XOR2_X1 U9371 ( .A(n9433), .B(n9434), .Z(n9228) );
  XNOR2_X1 U9372 ( .A(n9435), .B(n9436), .ZN(n9434) );
  XNOR2_X1 U9373 ( .A(n9437), .B(n9438), .ZN(n9231) );
  XNOR2_X1 U9374 ( .A(n9439), .B(n9440), .ZN(n9437) );
  NOR2_X1 U9375 ( .A1(n7957), .A2(n7522), .ZN(n9440) );
  XOR2_X1 U9376 ( .A(n9441), .B(n9442), .Z(n9236) );
  XNOR2_X1 U9377 ( .A(n9443), .B(n9444), .ZN(n9442) );
  XNOR2_X1 U9378 ( .A(n9445), .B(n9446), .ZN(n9240) );
  XNOR2_X1 U9379 ( .A(n9447), .B(n9448), .ZN(n9445) );
  NOR2_X1 U9380 ( .A1(n7960), .A2(n7522), .ZN(n9448) );
  XOR2_X1 U9381 ( .A(n9449), .B(n9450), .Z(n9243) );
  XOR2_X1 U9382 ( .A(n9451), .B(n9452), .Z(n9449) );
  XNOR2_X1 U9383 ( .A(n9453), .B(n9454), .ZN(n9247) );
  XOR2_X1 U9384 ( .A(n9455), .B(n9456), .Z(n9454) );
  NAND2_X1 U9385 ( .A1(b_25_), .A2(a_16_), .ZN(n9456) );
  XNOR2_X1 U9386 ( .A(n9457), .B(n9458), .ZN(n9252) );
  XNOR2_X1 U9387 ( .A(n9459), .B(n9460), .ZN(n9458) );
  XNOR2_X1 U9388 ( .A(n9461), .B(n9462), .ZN(n9256) );
  XNOR2_X1 U9389 ( .A(n9463), .B(n9464), .ZN(n9461) );
  NOR2_X1 U9390 ( .A1(n7962), .A2(n7522), .ZN(n9464) );
  XNOR2_X1 U9391 ( .A(n9465), .B(n9466), .ZN(n9260) );
  XOR2_X1 U9392 ( .A(n9467), .B(n9468), .Z(n9465) );
  XOR2_X1 U9393 ( .A(n9469), .B(n9470), .Z(n9263) );
  XOR2_X1 U9394 ( .A(n9471), .B(n9472), .Z(n9469) );
  NOR2_X1 U9395 ( .A1(n8585), .A2(n7522), .ZN(n9472) );
  XOR2_X1 U9396 ( .A(n9473), .B(n9474), .Z(n9268) );
  XOR2_X1 U9397 ( .A(n9475), .B(n9476), .Z(n9474) );
  NAND2_X1 U9398 ( .A1(b_25_), .A2(a_11_), .ZN(n9476) );
  XNOR2_X1 U9399 ( .A(n9477), .B(n9478), .ZN(n9272) );
  XOR2_X1 U9400 ( .A(n9479), .B(n9480), .Z(n9477) );
  NOR2_X1 U9401 ( .A1(n8378), .A2(n7522), .ZN(n9480) );
  XOR2_X1 U9402 ( .A(n9481), .B(n9482), .Z(n9275) );
  XOR2_X1 U9403 ( .A(n9483), .B(n9484), .Z(n9481) );
  XNOR2_X1 U9404 ( .A(n9485), .B(n9486), .ZN(n9284) );
  XOR2_X1 U9405 ( .A(n9487), .B(n9488), .Z(n9485) );
  NOR2_X1 U9406 ( .A1(n7787), .A2(n7522), .ZN(n9488) );
  XNOR2_X1 U9407 ( .A(n9489), .B(n9490), .ZN(n9287) );
  XOR2_X1 U9408 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR2_X1 U9409 ( .A(n9493), .B(n9494), .Z(n9102) );
  XOR2_X1 U9410 ( .A(n9495), .B(n9496), .Z(n9493) );
  NOR2_X1 U9411 ( .A1(n7823), .A2(n7522), .ZN(n9496) );
  XOR2_X1 U9412 ( .A(n9497), .B(n9498), .Z(n9095) );
  XOR2_X1 U9413 ( .A(n9499), .B(n9500), .Z(n9498) );
  NAND2_X1 U9414 ( .A1(b_25_), .A2(a_4_), .ZN(n9500) );
  XNOR2_X1 U9415 ( .A(n9501), .B(n9502), .ZN(n9291) );
  XOR2_X1 U9416 ( .A(n9503), .B(n9504), .Z(n9502) );
  NAND2_X1 U9417 ( .A1(b_25_), .A2(a_3_), .ZN(n9504) );
  XOR2_X1 U9418 ( .A(n9505), .B(n9506), .Z(n9296) );
  XOR2_X1 U9419 ( .A(n9507), .B(n9508), .Z(n9506) );
  NAND2_X1 U9420 ( .A1(b_25_), .A2(a_2_), .ZN(n9508) );
  XNOR2_X1 U9421 ( .A(n9509), .B(n9510), .ZN(n9081) );
  XOR2_X1 U9422 ( .A(n9511), .B(n9512), .Z(n9509) );
  NOR2_X1 U9423 ( .A1(n7872), .A2(n7522), .ZN(n9512) );
  NAND2_X1 U9424 ( .A1(n9513), .A2(n9514), .ZN(n8173) );
  XNOR2_X1 U9425 ( .A(n9515), .B(n9516), .ZN(n8174) );
  XNOR2_X1 U9426 ( .A(n9517), .B(n9518), .ZN(n9516) );
  NAND2_X1 U9427 ( .A1(n9519), .A2(n9299), .ZN(n8012) );
  NOR2_X1 U9428 ( .A1(n9514), .A2(n9513), .ZN(n9299) );
  AND2_X1 U9429 ( .A1(n9520), .A2(n9521), .ZN(n9513) );
  NAND2_X1 U9430 ( .A1(n9518), .A2(n9522), .ZN(n9521) );
  OR2_X1 U9431 ( .A1(n9517), .A2(n9515), .ZN(n9522) );
  NOR2_X1 U9432 ( .A1(n7522), .A2(n8197), .ZN(n9518) );
  NAND2_X1 U9433 ( .A1(n9515), .A2(n9517), .ZN(n9520) );
  NAND2_X1 U9434 ( .A1(n9523), .A2(n9524), .ZN(n9517) );
  NAND3_X1 U9435 ( .A1(a_1_), .A2(n9525), .A3(b_25_), .ZN(n9524) );
  OR2_X1 U9436 ( .A1(n9511), .A2(n9510), .ZN(n9525) );
  NAND2_X1 U9437 ( .A1(n9510), .A2(n9511), .ZN(n9523) );
  NAND2_X1 U9438 ( .A1(n9526), .A2(n9527), .ZN(n9511) );
  NAND3_X1 U9439 ( .A1(a_2_), .A2(n9528), .A3(b_25_), .ZN(n9527) );
  OR2_X1 U9440 ( .A1(n9507), .A2(n9505), .ZN(n9528) );
  NAND2_X1 U9441 ( .A1(n9505), .A2(n9507), .ZN(n9526) );
  NAND2_X1 U9442 ( .A1(n9529), .A2(n9530), .ZN(n9507) );
  NAND3_X1 U9443 ( .A1(a_3_), .A2(n9531), .A3(b_25_), .ZN(n9530) );
  OR2_X1 U9444 ( .A1(n9503), .A2(n9501), .ZN(n9531) );
  NAND2_X1 U9445 ( .A1(n9501), .A2(n9503), .ZN(n9529) );
  NAND2_X1 U9446 ( .A1(n9532), .A2(n9533), .ZN(n9503) );
  NAND3_X1 U9447 ( .A1(a_4_), .A2(n9534), .A3(b_25_), .ZN(n9533) );
  OR2_X1 U9448 ( .A1(n9499), .A2(n9497), .ZN(n9534) );
  NAND2_X1 U9449 ( .A1(n9497), .A2(n9499), .ZN(n9532) );
  NAND2_X1 U9450 ( .A1(n9535), .A2(n9536), .ZN(n9499) );
  NAND3_X1 U9451 ( .A1(a_5_), .A2(n9537), .A3(b_25_), .ZN(n9536) );
  OR2_X1 U9452 ( .A1(n9495), .A2(n9494), .ZN(n9537) );
  NAND2_X1 U9453 ( .A1(n9494), .A2(n9495), .ZN(n9535) );
  NAND2_X1 U9454 ( .A1(n9538), .A2(n9539), .ZN(n9495) );
  NAND2_X1 U9455 ( .A1(n9491), .A2(n9540), .ZN(n9539) );
  NAND2_X1 U9456 ( .A1(n9541), .A2(n9492), .ZN(n9540) );
  INV_X1 U9457 ( .A(n9489), .ZN(n9541) );
  NAND2_X1 U9458 ( .A1(n9542), .A2(n9543), .ZN(n9491) );
  NAND3_X1 U9459 ( .A1(a_7_), .A2(n9544), .A3(b_25_), .ZN(n9543) );
  OR2_X1 U9460 ( .A1(n9487), .A2(n9486), .ZN(n9544) );
  NAND2_X1 U9461 ( .A1(n9486), .A2(n9487), .ZN(n9542) );
  NAND2_X1 U9462 ( .A1(n9545), .A2(n9546), .ZN(n9487) );
  NAND3_X1 U9463 ( .A1(a_8_), .A2(n9547), .A3(b_25_), .ZN(n9546) );
  OR2_X1 U9464 ( .A1(n9327), .A2(n9326), .ZN(n9547) );
  NAND2_X1 U9465 ( .A1(n9326), .A2(n9327), .ZN(n9545) );
  NAND2_X1 U9466 ( .A1(n9548), .A2(n9549), .ZN(n9327) );
  NAND2_X1 U9467 ( .A1(n9484), .A2(n9550), .ZN(n9549) );
  OR2_X1 U9468 ( .A1(n9483), .A2(n9482), .ZN(n9550) );
  NOR2_X1 U9469 ( .A1(n7522), .A2(n7753), .ZN(n9484) );
  NAND2_X1 U9470 ( .A1(n9482), .A2(n9483), .ZN(n9548) );
  NAND2_X1 U9471 ( .A1(n9551), .A2(n9552), .ZN(n9483) );
  NAND3_X1 U9472 ( .A1(a_10_), .A2(n9553), .A3(b_25_), .ZN(n9552) );
  OR2_X1 U9473 ( .A1(n9479), .A2(n9478), .ZN(n9553) );
  NAND2_X1 U9474 ( .A1(n9478), .A2(n9479), .ZN(n9551) );
  NAND2_X1 U9475 ( .A1(n9554), .A2(n9555), .ZN(n9479) );
  NAND3_X1 U9476 ( .A1(a_11_), .A2(n9556), .A3(b_25_), .ZN(n9555) );
  OR2_X1 U9477 ( .A1(n9475), .A2(n9473), .ZN(n9556) );
  NAND2_X1 U9478 ( .A1(n9473), .A2(n9475), .ZN(n9554) );
  NAND2_X1 U9479 ( .A1(n9557), .A2(n9558), .ZN(n9475) );
  NAND3_X1 U9480 ( .A1(a_12_), .A2(n9559), .A3(b_25_), .ZN(n9558) );
  OR2_X1 U9481 ( .A1(n9471), .A2(n9470), .ZN(n9559) );
  NAND2_X1 U9482 ( .A1(n9470), .A2(n9471), .ZN(n9557) );
  NAND2_X1 U9483 ( .A1(n9560), .A2(n9561), .ZN(n9471) );
  NAND2_X1 U9484 ( .A1(n9468), .A2(n9562), .ZN(n9561) );
  OR2_X1 U9485 ( .A1(n9467), .A2(n9466), .ZN(n9562) );
  NOR2_X1 U9486 ( .A1(n7522), .A2(n7702), .ZN(n9468) );
  NAND2_X1 U9487 ( .A1(n9466), .A2(n9467), .ZN(n9560) );
  NAND2_X1 U9488 ( .A1(n9563), .A2(n9564), .ZN(n9467) );
  NAND3_X1 U9489 ( .A1(a_14_), .A2(n9565), .A3(b_25_), .ZN(n9564) );
  NAND2_X1 U9490 ( .A1(n9463), .A2(n9462), .ZN(n9565) );
  OR2_X1 U9491 ( .A1(n9462), .A2(n9463), .ZN(n9563) );
  AND2_X1 U9492 ( .A1(n9566), .A2(n9567), .ZN(n9463) );
  NAND2_X1 U9493 ( .A1(n9460), .A2(n9568), .ZN(n9567) );
  OR2_X1 U9494 ( .A1(n9459), .A2(n9457), .ZN(n9568) );
  NOR2_X1 U9495 ( .A1(n7522), .A2(n7667), .ZN(n9460) );
  NAND2_X1 U9496 ( .A1(n9457), .A2(n9459), .ZN(n9566) );
  NAND2_X1 U9497 ( .A1(n9569), .A2(n9570), .ZN(n9459) );
  NAND3_X1 U9498 ( .A1(a_16_), .A2(n9571), .A3(b_25_), .ZN(n9570) );
  OR2_X1 U9499 ( .A1(n9455), .A2(n9453), .ZN(n9571) );
  NAND2_X1 U9500 ( .A1(n9453), .A2(n9455), .ZN(n9569) );
  NAND2_X1 U9501 ( .A1(n9572), .A2(n9573), .ZN(n9455) );
  NAND2_X1 U9502 ( .A1(n9452), .A2(n9574), .ZN(n9573) );
  OR2_X1 U9503 ( .A1(n9451), .A2(n9450), .ZN(n9574) );
  NOR2_X1 U9504 ( .A1(n7522), .A2(n7645), .ZN(n9452) );
  NAND2_X1 U9505 ( .A1(n9450), .A2(n9451), .ZN(n9572) );
  NAND2_X1 U9506 ( .A1(n9575), .A2(n9576), .ZN(n9451) );
  NAND3_X1 U9507 ( .A1(a_18_), .A2(n9577), .A3(b_25_), .ZN(n9576) );
  NAND2_X1 U9508 ( .A1(n9447), .A2(n9446), .ZN(n9577) );
  OR2_X1 U9509 ( .A1(n9446), .A2(n9447), .ZN(n9575) );
  AND2_X1 U9510 ( .A1(n9578), .A2(n9579), .ZN(n9447) );
  NAND2_X1 U9511 ( .A1(n9444), .A2(n9580), .ZN(n9579) );
  OR2_X1 U9512 ( .A1(n9443), .A2(n9441), .ZN(n9580) );
  NOR2_X1 U9513 ( .A1(n7522), .A2(n7958), .ZN(n9444) );
  NAND2_X1 U9514 ( .A1(n9441), .A2(n9443), .ZN(n9578) );
  NAND2_X1 U9515 ( .A1(n9581), .A2(n9582), .ZN(n9443) );
  NAND3_X1 U9516 ( .A1(a_20_), .A2(n9583), .A3(b_25_), .ZN(n9582) );
  NAND2_X1 U9517 ( .A1(n9439), .A2(n9438), .ZN(n9583) );
  OR2_X1 U9518 ( .A1(n9438), .A2(n9439), .ZN(n9581) );
  AND2_X1 U9519 ( .A1(n9584), .A2(n9585), .ZN(n9439) );
  NAND2_X1 U9520 ( .A1(n9436), .A2(n9586), .ZN(n9585) );
  OR2_X1 U9521 ( .A1(n9435), .A2(n9433), .ZN(n9586) );
  NOR2_X1 U9522 ( .A1(n7522), .A2(n7578), .ZN(n9436) );
  NAND2_X1 U9523 ( .A1(n9433), .A2(n9435), .ZN(n9584) );
  NAND2_X1 U9524 ( .A1(n9587), .A2(n9588), .ZN(n9435) );
  NAND3_X1 U9525 ( .A1(a_22_), .A2(n9589), .A3(b_25_), .ZN(n9588) );
  OR2_X1 U9526 ( .A1(n9431), .A2(n9429), .ZN(n9589) );
  NAND2_X1 U9527 ( .A1(n9429), .A2(n9431), .ZN(n9587) );
  NAND2_X1 U9528 ( .A1(n9590), .A2(n9591), .ZN(n9431) );
  NAND2_X1 U9529 ( .A1(n9428), .A2(n9592), .ZN(n9591) );
  OR2_X1 U9530 ( .A1(n9427), .A2(n9425), .ZN(n9592) );
  NOR2_X1 U9531 ( .A1(n7522), .A2(n7955), .ZN(n9428) );
  NAND2_X1 U9532 ( .A1(n9425), .A2(n9427), .ZN(n9590) );
  NAND2_X1 U9533 ( .A1(n9593), .A2(n9594), .ZN(n9427) );
  NAND3_X1 U9534 ( .A1(a_24_), .A2(n9595), .A3(b_25_), .ZN(n9594) );
  NAND2_X1 U9535 ( .A1(n9423), .A2(n9422), .ZN(n9595) );
  OR2_X1 U9536 ( .A1(n9422), .A2(n9423), .ZN(n9593) );
  AND2_X1 U9537 ( .A1(n9596), .A2(n9597), .ZN(n9423) );
  NAND2_X1 U9538 ( .A1(n7520), .A2(n9598), .ZN(n9597) );
  OR2_X1 U9539 ( .A1(n9420), .A2(n9419), .ZN(n9598) );
  INV_X1 U9540 ( .A(n7934), .ZN(n7520) );
  NAND2_X1 U9541 ( .A1(b_25_), .A2(a_25_), .ZN(n7934) );
  NAND2_X1 U9542 ( .A1(n9419), .A2(n9420), .ZN(n9596) );
  NAND2_X1 U9543 ( .A1(n9416), .A2(n9599), .ZN(n9420) );
  NAND2_X1 U9544 ( .A1(n9415), .A2(n9417), .ZN(n9599) );
  NAND2_X1 U9545 ( .A1(n9600), .A2(n9601), .ZN(n9417) );
  NAND2_X1 U9546 ( .A1(b_25_), .A2(a_26_), .ZN(n9601) );
  INV_X1 U9547 ( .A(n9602), .ZN(n9600) );
  XNOR2_X1 U9548 ( .A(n9603), .B(n9604), .ZN(n9415) );
  NAND2_X1 U9549 ( .A1(n9605), .A2(n9606), .ZN(n9603) );
  NAND2_X1 U9550 ( .A1(a_26_), .A2(n9602), .ZN(n9416) );
  NAND2_X1 U9551 ( .A1(n9388), .A2(n9607), .ZN(n9602) );
  NAND2_X1 U9552 ( .A1(n9387), .A2(n9389), .ZN(n9607) );
  NAND2_X1 U9553 ( .A1(n9608), .A2(n9609), .ZN(n9389) );
  NAND2_X1 U9554 ( .A1(b_25_), .A2(a_27_), .ZN(n9609) );
  INV_X1 U9555 ( .A(n9610), .ZN(n9608) );
  XNOR2_X1 U9556 ( .A(n9611), .B(n9612), .ZN(n9387) );
  XOR2_X1 U9557 ( .A(n9613), .B(n9614), .Z(n9611) );
  NAND2_X1 U9558 ( .A1(b_24_), .A2(a_28_), .ZN(n9613) );
  NAND2_X1 U9559 ( .A1(a_27_), .A2(n9610), .ZN(n9388) );
  NAND2_X1 U9560 ( .A1(n9615), .A2(n9616), .ZN(n9610) );
  NAND3_X1 U9561 ( .A1(a_28_), .A2(n9617), .A3(b_25_), .ZN(n9616) );
  NAND2_X1 U9562 ( .A1(n9397), .A2(n9395), .ZN(n9617) );
  OR2_X1 U9563 ( .A1(n9395), .A2(n9397), .ZN(n9615) );
  AND2_X1 U9564 ( .A1(n9618), .A2(n9619), .ZN(n9397) );
  NAND2_X1 U9565 ( .A1(n9411), .A2(n9620), .ZN(n9619) );
  OR2_X1 U9566 ( .A1(n9412), .A2(n9413), .ZN(n9620) );
  NOR2_X1 U9567 ( .A1(n7522), .A2(n7460), .ZN(n9411) );
  INV_X1 U9568 ( .A(b_25_), .ZN(n7522) );
  NAND2_X1 U9569 ( .A1(n9413), .A2(n9412), .ZN(n9618) );
  NAND2_X1 U9570 ( .A1(n9621), .A2(n9622), .ZN(n9412) );
  NAND2_X1 U9571 ( .A1(b_23_), .A2(n9623), .ZN(n9622) );
  NAND2_X1 U9572 ( .A1(n7441), .A2(n9624), .ZN(n9623) );
  NAND2_X1 U9573 ( .A1(a_31_), .A2(n7953), .ZN(n9624) );
  NAND2_X1 U9574 ( .A1(b_24_), .A2(n9625), .ZN(n9621) );
  NAND2_X1 U9575 ( .A1(n7445), .A2(n9626), .ZN(n9625) );
  NAND2_X1 U9576 ( .A1(a_30_), .A2(n7549), .ZN(n9626) );
  AND3_X1 U9577 ( .A1(b_24_), .A2(n7409), .A3(b_25_), .ZN(n9413) );
  XNOR2_X1 U9578 ( .A(n9627), .B(n9628), .ZN(n9395) );
  XOR2_X1 U9579 ( .A(n9629), .B(n9630), .Z(n9627) );
  XNOR2_X1 U9580 ( .A(n9631), .B(n9632), .ZN(n9419) );
  NAND2_X1 U9581 ( .A1(n9633), .A2(n9634), .ZN(n9631) );
  XNOR2_X1 U9582 ( .A(n9635), .B(n9636), .ZN(n9422) );
  XOR2_X1 U9583 ( .A(n9637), .B(n9638), .Z(n9635) );
  XOR2_X1 U9584 ( .A(n9639), .B(n9640), .Z(n9425) );
  XOR2_X1 U9585 ( .A(n9641), .B(n9642), .Z(n9639) );
  XOR2_X1 U9586 ( .A(n9643), .B(n9644), .Z(n9429) );
  XOR2_X1 U9587 ( .A(n9645), .B(n9646), .Z(n9643) );
  XNOR2_X1 U9588 ( .A(n9647), .B(n9648), .ZN(n9433) );
  XOR2_X1 U9589 ( .A(n9649), .B(n9650), .Z(n9648) );
  NAND2_X1 U9590 ( .A1(b_24_), .A2(a_22_), .ZN(n9650) );
  XNOR2_X1 U9591 ( .A(n9651), .B(n9652), .ZN(n9438) );
  XOR2_X1 U9592 ( .A(n9653), .B(n9654), .Z(n9651) );
  XNOR2_X1 U9593 ( .A(n9655), .B(n9656), .ZN(n9441) );
  XNOR2_X1 U9594 ( .A(n9657), .B(n9658), .ZN(n9655) );
  NOR2_X1 U9595 ( .A1(n7957), .A2(n7953), .ZN(n9658) );
  XOR2_X1 U9596 ( .A(n9659), .B(n9660), .Z(n9446) );
  XNOR2_X1 U9597 ( .A(n9661), .B(n9662), .ZN(n9660) );
  XNOR2_X1 U9598 ( .A(n9663), .B(n9664), .ZN(n9450) );
  XNOR2_X1 U9599 ( .A(n9665), .B(n9666), .ZN(n9663) );
  NOR2_X1 U9600 ( .A1(n7960), .A2(n7953), .ZN(n9666) );
  XOR2_X1 U9601 ( .A(n9667), .B(n9668), .Z(n9453) );
  XOR2_X1 U9602 ( .A(n9669), .B(n9670), .Z(n9667) );
  XOR2_X1 U9603 ( .A(n9671), .B(n9672), .Z(n9457) );
  XOR2_X1 U9604 ( .A(n9673), .B(n9674), .Z(n9671) );
  NOR2_X1 U9605 ( .A1(n8353), .A2(n7953), .ZN(n9674) );
  XOR2_X1 U9606 ( .A(n9675), .B(n9676), .Z(n9462) );
  XNOR2_X1 U9607 ( .A(n9677), .B(n9678), .ZN(n9676) );
  XNOR2_X1 U9608 ( .A(n9679), .B(n9680), .ZN(n9466) );
  XOR2_X1 U9609 ( .A(n9681), .B(n9682), .Z(n9679) );
  NAND2_X1 U9610 ( .A1(b_24_), .A2(a_14_), .ZN(n9681) );
  XNOR2_X1 U9611 ( .A(n9683), .B(n9684), .ZN(n9470) );
  XNOR2_X1 U9612 ( .A(n9685), .B(n9686), .ZN(n9683) );
  XNOR2_X1 U9613 ( .A(n9687), .B(n9688), .ZN(n9473) );
  XOR2_X1 U9614 ( .A(n9689), .B(n9690), .Z(n9688) );
  NAND2_X1 U9615 ( .A1(b_24_), .A2(a_12_), .ZN(n9690) );
  XNOR2_X1 U9616 ( .A(n9691), .B(n9692), .ZN(n9478) );
  NAND2_X1 U9617 ( .A1(n9693), .A2(n9694), .ZN(n9691) );
  XNOR2_X1 U9618 ( .A(n9695), .B(n9696), .ZN(n9482) );
  XNOR2_X1 U9619 ( .A(n9697), .B(n9698), .ZN(n9696) );
  NOR2_X1 U9620 ( .A1(n8378), .A2(n7953), .ZN(n9698) );
  XNOR2_X1 U9621 ( .A(n9699), .B(n9700), .ZN(n9326) );
  XNOR2_X1 U9622 ( .A(n9701), .B(n9702), .ZN(n9700) );
  XNOR2_X1 U9623 ( .A(n9703), .B(n9704), .ZN(n9486) );
  XOR2_X1 U9624 ( .A(n9705), .B(n9706), .Z(n9703) );
  NAND2_X1 U9625 ( .A1(b_24_), .A2(a_8_), .ZN(n9705) );
  NAND2_X1 U9626 ( .A1(n9707), .A2(n9489), .ZN(n9538) );
  XNOR2_X1 U9627 ( .A(n9708), .B(n9709), .ZN(n9489) );
  NAND2_X1 U9628 ( .A1(n9710), .A2(n9711), .ZN(n9708) );
  INV_X1 U9629 ( .A(n9492), .ZN(n9707) );
  NAND2_X1 U9630 ( .A1(b_25_), .A2(a_6_), .ZN(n9492) );
  XNOR2_X1 U9631 ( .A(n9712), .B(n9713), .ZN(n9494) );
  XNOR2_X1 U9632 ( .A(n9714), .B(n9715), .ZN(n9712) );
  XNOR2_X1 U9633 ( .A(n9716), .B(n9717), .ZN(n9497) );
  XNOR2_X1 U9634 ( .A(n9718), .B(n9719), .ZN(n9717) );
  XNOR2_X1 U9635 ( .A(n9720), .B(n9721), .ZN(n9501) );
  XOR2_X1 U9636 ( .A(n9722), .B(n9723), .Z(n9720) );
  NAND2_X1 U9637 ( .A1(b_24_), .A2(a_4_), .ZN(n9722) );
  XNOR2_X1 U9638 ( .A(n9724), .B(n9725), .ZN(n9505) );
  NAND2_X1 U9639 ( .A1(n9726), .A2(n9727), .ZN(n9724) );
  XNOR2_X1 U9640 ( .A(n9728), .B(n9729), .ZN(n9510) );
  NAND2_X1 U9641 ( .A1(n9730), .A2(n9731), .ZN(n9728) );
  XNOR2_X1 U9642 ( .A(n9732), .B(n9733), .ZN(n9515) );
  NAND2_X1 U9643 ( .A1(n9734), .A2(n9735), .ZN(n9732) );
  XOR2_X1 U9644 ( .A(n9736), .B(n9737), .Z(n9514) );
  NAND2_X1 U9645 ( .A1(n9738), .A2(n9739), .ZN(n9736) );
  XOR2_X1 U9646 ( .A(n8164), .B(n8165), .Z(n9519) );
  NAND3_X1 U9647 ( .A1(n8164), .A2(n8165), .A3(n9740), .ZN(n8016) );
  XOR2_X1 U9648 ( .A(n8160), .B(n8159), .Z(n9740) );
  NAND2_X1 U9649 ( .A1(n9738), .A2(n9741), .ZN(n8165) );
  NAND2_X1 U9650 ( .A1(n9737), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U9651 ( .A1(n9742), .A2(n9743), .ZN(n9739) );
  NAND2_X1 U9652 ( .A1(b_24_), .A2(a_0_), .ZN(n9743) );
  INV_X1 U9653 ( .A(n9744), .ZN(n9742) );
  XNOR2_X1 U9654 ( .A(n9745), .B(n9746), .ZN(n9737) );
  XOR2_X1 U9655 ( .A(n9747), .B(n9748), .Z(n9746) );
  NAND2_X1 U9656 ( .A1(b_23_), .A2(a_1_), .ZN(n9748) );
  NAND2_X1 U9657 ( .A1(a_0_), .A2(n9744), .ZN(n9738) );
  NAND2_X1 U9658 ( .A1(n9734), .A2(n9749), .ZN(n9744) );
  NAND2_X1 U9659 ( .A1(n9733), .A2(n9735), .ZN(n9749) );
  NAND2_X1 U9660 ( .A1(n9750), .A2(n9751), .ZN(n9735) );
  NAND2_X1 U9661 ( .A1(b_24_), .A2(a_1_), .ZN(n9751) );
  INV_X1 U9662 ( .A(n9752), .ZN(n9750) );
  XNOR2_X1 U9663 ( .A(n9753), .B(n9754), .ZN(n9733) );
  XNOR2_X1 U9664 ( .A(n9755), .B(n9756), .ZN(n9753) );
  NOR2_X1 U9665 ( .A1(n7966), .A2(n7549), .ZN(n9756) );
  NAND2_X1 U9666 ( .A1(a_1_), .A2(n9752), .ZN(n9734) );
  NAND2_X1 U9667 ( .A1(n9730), .A2(n9757), .ZN(n9752) );
  NAND2_X1 U9668 ( .A1(n9729), .A2(n9731), .ZN(n9757) );
  NAND2_X1 U9669 ( .A1(n9758), .A2(n9759), .ZN(n9731) );
  NAND2_X1 U9670 ( .A1(b_24_), .A2(a_2_), .ZN(n9759) );
  INV_X1 U9671 ( .A(n9760), .ZN(n9758) );
  XNOR2_X1 U9672 ( .A(n9761), .B(n9762), .ZN(n9729) );
  XOR2_X1 U9673 ( .A(n9763), .B(n9764), .Z(n9762) );
  NAND2_X1 U9674 ( .A1(b_23_), .A2(a_3_), .ZN(n9764) );
  NAND2_X1 U9675 ( .A1(a_2_), .A2(n9760), .ZN(n9730) );
  NAND2_X1 U9676 ( .A1(n9726), .A2(n9765), .ZN(n9760) );
  NAND2_X1 U9677 ( .A1(n9725), .A2(n9727), .ZN(n9765) );
  NAND2_X1 U9678 ( .A1(n9766), .A2(n9767), .ZN(n9727) );
  NAND2_X1 U9679 ( .A1(b_24_), .A2(a_3_), .ZN(n9767) );
  INV_X1 U9680 ( .A(n9768), .ZN(n9766) );
  XNOR2_X1 U9681 ( .A(n9769), .B(n9770), .ZN(n9725) );
  XOR2_X1 U9682 ( .A(n9771), .B(n9772), .Z(n9770) );
  NAND2_X1 U9683 ( .A1(b_23_), .A2(a_4_), .ZN(n9772) );
  NAND2_X1 U9684 ( .A1(a_3_), .A2(n9768), .ZN(n9726) );
  NAND2_X1 U9685 ( .A1(n9773), .A2(n9774), .ZN(n9768) );
  NAND3_X1 U9686 ( .A1(a_4_), .A2(n9775), .A3(b_24_), .ZN(n9774) );
  NAND2_X1 U9687 ( .A1(n9723), .A2(n9721), .ZN(n9775) );
  OR2_X1 U9688 ( .A1(n9721), .A2(n9723), .ZN(n9773) );
  AND2_X1 U9689 ( .A1(n9776), .A2(n9777), .ZN(n9723) );
  NAND2_X1 U9690 ( .A1(n9719), .A2(n9778), .ZN(n9777) );
  OR2_X1 U9691 ( .A1(n9718), .A2(n9716), .ZN(n9778) );
  NOR2_X1 U9692 ( .A1(n7953), .A2(n7823), .ZN(n9719) );
  NAND2_X1 U9693 ( .A1(n9716), .A2(n9718), .ZN(n9776) );
  NAND2_X1 U9694 ( .A1(n9779), .A2(n9780), .ZN(n9718) );
  NAND2_X1 U9695 ( .A1(n9715), .A2(n9781), .ZN(n9780) );
  NAND2_X1 U9696 ( .A1(n9713), .A2(n9714), .ZN(n9781) );
  NAND2_X1 U9697 ( .A1(n9710), .A2(n9782), .ZN(n9715) );
  NAND2_X1 U9698 ( .A1(n9709), .A2(n9711), .ZN(n9782) );
  NAND2_X1 U9699 ( .A1(n9783), .A2(n9784), .ZN(n9711) );
  NAND2_X1 U9700 ( .A1(b_24_), .A2(a_7_), .ZN(n9784) );
  INV_X1 U9701 ( .A(n9785), .ZN(n9783) );
  XNOR2_X1 U9702 ( .A(n9786), .B(n9787), .ZN(n9709) );
  XNOR2_X1 U9703 ( .A(n9788), .B(n9789), .ZN(n9787) );
  NAND2_X1 U9704 ( .A1(a_7_), .A2(n9785), .ZN(n9710) );
  NAND2_X1 U9705 ( .A1(n9790), .A2(n9791), .ZN(n9785) );
  NAND3_X1 U9706 ( .A1(a_8_), .A2(n9792), .A3(b_24_), .ZN(n9791) );
  NAND2_X1 U9707 ( .A1(n9706), .A2(n9704), .ZN(n9792) );
  OR2_X1 U9708 ( .A1(n9704), .A2(n9706), .ZN(n9790) );
  AND2_X1 U9709 ( .A1(n9793), .A2(n9794), .ZN(n9706) );
  NAND2_X1 U9710 ( .A1(n9702), .A2(n9795), .ZN(n9794) );
  OR2_X1 U9711 ( .A1(n9701), .A2(n9699), .ZN(n9795) );
  NOR2_X1 U9712 ( .A1(n7953), .A2(n7753), .ZN(n9702) );
  NAND2_X1 U9713 ( .A1(n9699), .A2(n9701), .ZN(n9793) );
  NAND2_X1 U9714 ( .A1(n9796), .A2(n9797), .ZN(n9701) );
  NAND3_X1 U9715 ( .A1(a_10_), .A2(n9798), .A3(b_24_), .ZN(n9797) );
  OR2_X1 U9716 ( .A1(n9697), .A2(n9695), .ZN(n9798) );
  NAND2_X1 U9717 ( .A1(n9695), .A2(n9697), .ZN(n9796) );
  NAND2_X1 U9718 ( .A1(n9693), .A2(n9799), .ZN(n9697) );
  NAND2_X1 U9719 ( .A1(n9692), .A2(n9694), .ZN(n9799) );
  NAND2_X1 U9720 ( .A1(n9800), .A2(n9801), .ZN(n9694) );
  NAND2_X1 U9721 ( .A1(b_24_), .A2(a_11_), .ZN(n9801) );
  INV_X1 U9722 ( .A(n9802), .ZN(n9800) );
  XNOR2_X1 U9723 ( .A(n9803), .B(n9804), .ZN(n9692) );
  XNOR2_X1 U9724 ( .A(n9805), .B(n9806), .ZN(n9803) );
  NOR2_X1 U9725 ( .A1(n8585), .A2(n7549), .ZN(n9806) );
  NAND2_X1 U9726 ( .A1(a_11_), .A2(n9802), .ZN(n9693) );
  NAND2_X1 U9727 ( .A1(n9807), .A2(n9808), .ZN(n9802) );
  NAND3_X1 U9728 ( .A1(a_12_), .A2(n9809), .A3(b_24_), .ZN(n9808) );
  OR2_X1 U9729 ( .A1(n9689), .A2(n9687), .ZN(n9809) );
  NAND2_X1 U9730 ( .A1(n9687), .A2(n9689), .ZN(n9807) );
  NAND2_X1 U9731 ( .A1(n9810), .A2(n9811), .ZN(n9689) );
  NAND2_X1 U9732 ( .A1(n9686), .A2(n9812), .ZN(n9811) );
  NAND2_X1 U9733 ( .A1(n9685), .A2(n9684), .ZN(n9812) );
  NOR2_X1 U9734 ( .A1(n7953), .A2(n7702), .ZN(n9686) );
  OR2_X1 U9735 ( .A1(n9684), .A2(n9685), .ZN(n9810) );
  AND2_X1 U9736 ( .A1(n9813), .A2(n9814), .ZN(n9685) );
  NAND3_X1 U9737 ( .A1(a_14_), .A2(n9815), .A3(b_24_), .ZN(n9814) );
  NAND2_X1 U9738 ( .A1(n9682), .A2(n9680), .ZN(n9815) );
  OR2_X1 U9739 ( .A1(n9680), .A2(n9682), .ZN(n9813) );
  AND2_X1 U9740 ( .A1(n9816), .A2(n9817), .ZN(n9682) );
  NAND2_X1 U9741 ( .A1(n9678), .A2(n9818), .ZN(n9817) );
  OR2_X1 U9742 ( .A1(n9677), .A2(n9675), .ZN(n9818) );
  NOR2_X1 U9743 ( .A1(n7953), .A2(n7667), .ZN(n9678) );
  NAND2_X1 U9744 ( .A1(n9675), .A2(n9677), .ZN(n9816) );
  NAND2_X1 U9745 ( .A1(n9819), .A2(n9820), .ZN(n9677) );
  NAND3_X1 U9746 ( .A1(a_16_), .A2(n9821), .A3(b_24_), .ZN(n9820) );
  OR2_X1 U9747 ( .A1(n9673), .A2(n9672), .ZN(n9821) );
  NAND2_X1 U9748 ( .A1(n9672), .A2(n9673), .ZN(n9819) );
  NAND2_X1 U9749 ( .A1(n9822), .A2(n9823), .ZN(n9673) );
  NAND2_X1 U9750 ( .A1(n9670), .A2(n9824), .ZN(n9823) );
  OR2_X1 U9751 ( .A1(n9669), .A2(n9668), .ZN(n9824) );
  NOR2_X1 U9752 ( .A1(n7953), .A2(n7645), .ZN(n9670) );
  NAND2_X1 U9753 ( .A1(n9668), .A2(n9669), .ZN(n9822) );
  NAND2_X1 U9754 ( .A1(n9825), .A2(n9826), .ZN(n9669) );
  NAND3_X1 U9755 ( .A1(a_18_), .A2(n9827), .A3(b_24_), .ZN(n9826) );
  NAND2_X1 U9756 ( .A1(n9665), .A2(n9664), .ZN(n9827) );
  OR2_X1 U9757 ( .A1(n9664), .A2(n9665), .ZN(n9825) );
  AND2_X1 U9758 ( .A1(n9828), .A2(n9829), .ZN(n9665) );
  NAND2_X1 U9759 ( .A1(n9662), .A2(n9830), .ZN(n9829) );
  OR2_X1 U9760 ( .A1(n9661), .A2(n9659), .ZN(n9830) );
  NOR2_X1 U9761 ( .A1(n7953), .A2(n7958), .ZN(n9662) );
  NAND2_X1 U9762 ( .A1(n9659), .A2(n9661), .ZN(n9828) );
  NAND2_X1 U9763 ( .A1(n9831), .A2(n9832), .ZN(n9661) );
  NAND3_X1 U9764 ( .A1(a_20_), .A2(n9833), .A3(b_24_), .ZN(n9832) );
  NAND2_X1 U9765 ( .A1(n9657), .A2(n9656), .ZN(n9833) );
  OR2_X1 U9766 ( .A1(n9656), .A2(n9657), .ZN(n9831) );
  AND2_X1 U9767 ( .A1(n9834), .A2(n9835), .ZN(n9657) );
  NAND2_X1 U9768 ( .A1(n9654), .A2(n9836), .ZN(n9835) );
  OR2_X1 U9769 ( .A1(n9653), .A2(n9652), .ZN(n9836) );
  NOR2_X1 U9770 ( .A1(n7953), .A2(n7578), .ZN(n9654) );
  NAND2_X1 U9771 ( .A1(n9652), .A2(n9653), .ZN(n9834) );
  NAND2_X1 U9772 ( .A1(n9837), .A2(n9838), .ZN(n9653) );
  NAND3_X1 U9773 ( .A1(a_22_), .A2(n9839), .A3(b_24_), .ZN(n9838) );
  OR2_X1 U9774 ( .A1(n9649), .A2(n9647), .ZN(n9839) );
  NAND2_X1 U9775 ( .A1(n9647), .A2(n9649), .ZN(n9837) );
  NAND2_X1 U9776 ( .A1(n9840), .A2(n9841), .ZN(n9649) );
  NAND2_X1 U9777 ( .A1(n9646), .A2(n9842), .ZN(n9841) );
  OR2_X1 U9778 ( .A1(n9645), .A2(n9644), .ZN(n9842) );
  NOR2_X1 U9779 ( .A1(n7953), .A2(n7955), .ZN(n9646) );
  NAND2_X1 U9780 ( .A1(n9644), .A2(n9645), .ZN(n9840) );
  NAND2_X1 U9781 ( .A1(n9843), .A2(n9844), .ZN(n9645) );
  NAND2_X1 U9782 ( .A1(n9640), .A2(n9845), .ZN(n9844) );
  OR2_X1 U9783 ( .A1(n9641), .A2(n9642), .ZN(n9845) );
  XOR2_X1 U9784 ( .A(n9846), .B(n9847), .Z(n9640) );
  XOR2_X1 U9785 ( .A(n9848), .B(n9849), .Z(n9846) );
  NAND2_X1 U9786 ( .A1(n9642), .A2(n9641), .ZN(n9843) );
  NAND2_X1 U9787 ( .A1(n9850), .A2(n9851), .ZN(n9641) );
  NAND2_X1 U9788 ( .A1(n9638), .A2(n9852), .ZN(n9851) );
  OR2_X1 U9789 ( .A1(n9637), .A2(n9636), .ZN(n9852) );
  NOR2_X1 U9790 ( .A1(n7953), .A2(n7952), .ZN(n9638) );
  NAND2_X1 U9791 ( .A1(n9636), .A2(n9637), .ZN(n9850) );
  NAND2_X1 U9792 ( .A1(n9633), .A2(n9853), .ZN(n9637) );
  NAND2_X1 U9793 ( .A1(n9632), .A2(n9634), .ZN(n9853) );
  NAND2_X1 U9794 ( .A1(n9854), .A2(n9855), .ZN(n9634) );
  NAND2_X1 U9795 ( .A1(b_24_), .A2(a_26_), .ZN(n9855) );
  INV_X1 U9796 ( .A(n9856), .ZN(n9854) );
  XNOR2_X1 U9797 ( .A(n9857), .B(n9858), .ZN(n9632) );
  NAND2_X1 U9798 ( .A1(n9859), .A2(n9860), .ZN(n9857) );
  NAND2_X1 U9799 ( .A1(a_26_), .A2(n9856), .ZN(n9633) );
  NAND2_X1 U9800 ( .A1(n9605), .A2(n9861), .ZN(n9856) );
  NAND2_X1 U9801 ( .A1(n9604), .A2(n9606), .ZN(n9861) );
  NAND2_X1 U9802 ( .A1(n9862), .A2(n9863), .ZN(n9606) );
  NAND2_X1 U9803 ( .A1(b_24_), .A2(a_27_), .ZN(n9863) );
  INV_X1 U9804 ( .A(n9864), .ZN(n9862) );
  XNOR2_X1 U9805 ( .A(n9865), .B(n9866), .ZN(n9604) );
  XOR2_X1 U9806 ( .A(n9867), .B(n9868), .Z(n9865) );
  NAND2_X1 U9807 ( .A1(b_23_), .A2(a_28_), .ZN(n9867) );
  NAND2_X1 U9808 ( .A1(a_27_), .A2(n9864), .ZN(n9605) );
  NAND2_X1 U9809 ( .A1(n9869), .A2(n9870), .ZN(n9864) );
  NAND3_X1 U9810 ( .A1(a_28_), .A2(n9871), .A3(b_24_), .ZN(n9870) );
  NAND2_X1 U9811 ( .A1(n9614), .A2(n9612), .ZN(n9871) );
  OR2_X1 U9812 ( .A1(n9612), .A2(n9614), .ZN(n9869) );
  AND2_X1 U9813 ( .A1(n9872), .A2(n9873), .ZN(n9614) );
  NAND2_X1 U9814 ( .A1(n9628), .A2(n9874), .ZN(n9873) );
  OR2_X1 U9815 ( .A1(n9629), .A2(n9630), .ZN(n9874) );
  NOR2_X1 U9816 ( .A1(n7953), .A2(n7460), .ZN(n9628) );
  INV_X1 U9817 ( .A(b_24_), .ZN(n7953) );
  NAND2_X1 U9818 ( .A1(n9630), .A2(n9629), .ZN(n9872) );
  NAND2_X1 U9819 ( .A1(n9875), .A2(n9876), .ZN(n9629) );
  NAND2_X1 U9820 ( .A1(b_22_), .A2(n9877), .ZN(n9876) );
  NAND2_X1 U9821 ( .A1(n7441), .A2(n9878), .ZN(n9877) );
  NAND2_X1 U9822 ( .A1(a_31_), .A2(n7549), .ZN(n9878) );
  NAND2_X1 U9823 ( .A1(b_23_), .A2(n9879), .ZN(n9875) );
  NAND2_X1 U9824 ( .A1(n7445), .A2(n9880), .ZN(n9879) );
  NAND2_X1 U9825 ( .A1(a_30_), .A2(n9881), .ZN(n9880) );
  AND3_X1 U9826 ( .A1(b_23_), .A2(n7409), .A3(b_24_), .ZN(n9630) );
  XNOR2_X1 U9827 ( .A(n9882), .B(n9883), .ZN(n9612) );
  XOR2_X1 U9828 ( .A(n9884), .B(n9885), .Z(n9882) );
  XNOR2_X1 U9829 ( .A(n9886), .B(n9887), .ZN(n9636) );
  NAND2_X1 U9830 ( .A1(n9888), .A2(n9889), .ZN(n9886) );
  INV_X1 U9831 ( .A(n7535), .ZN(n9642) );
  NAND2_X1 U9832 ( .A1(b_24_), .A2(a_24_), .ZN(n7535) );
  XNOR2_X1 U9833 ( .A(n9890), .B(n9891), .ZN(n9644) );
  XNOR2_X1 U9834 ( .A(n9892), .B(n9893), .ZN(n9890) );
  NOR2_X1 U9835 ( .A1(n7954), .A2(n7549), .ZN(n9893) );
  XNOR2_X1 U9836 ( .A(n9894), .B(n9895), .ZN(n9647) );
  XNOR2_X1 U9837 ( .A(n9896), .B(n7547), .ZN(n9895) );
  XNOR2_X1 U9838 ( .A(n9897), .B(n9898), .ZN(n9652) );
  XOR2_X1 U9839 ( .A(n9899), .B(n9900), .Z(n9898) );
  NAND2_X1 U9840 ( .A1(b_23_), .A2(a_22_), .ZN(n9900) );
  XNOR2_X1 U9841 ( .A(n9901), .B(n9902), .ZN(n9656) );
  XOR2_X1 U9842 ( .A(n9903), .B(n9904), .Z(n9901) );
  XNOR2_X1 U9843 ( .A(n9905), .B(n9906), .ZN(n9659) );
  XNOR2_X1 U9844 ( .A(n9907), .B(n9908), .ZN(n9905) );
  NOR2_X1 U9845 ( .A1(n7957), .A2(n7549), .ZN(n9908) );
  XOR2_X1 U9846 ( .A(n9909), .B(n9910), .Z(n9664) );
  XNOR2_X1 U9847 ( .A(n9911), .B(n9912), .ZN(n9910) );
  XNOR2_X1 U9848 ( .A(n9913), .B(n9914), .ZN(n9668) );
  XNOR2_X1 U9849 ( .A(n9915), .B(n9916), .ZN(n9913) );
  NOR2_X1 U9850 ( .A1(n7960), .A2(n7549), .ZN(n9916) );
  XNOR2_X1 U9851 ( .A(n9917), .B(n9918), .ZN(n9672) );
  XNOR2_X1 U9852 ( .A(n9919), .B(n9920), .ZN(n9917) );
  XNOR2_X1 U9853 ( .A(n9921), .B(n9922), .ZN(n9675) );
  XOR2_X1 U9854 ( .A(n9923), .B(n9924), .Z(n9922) );
  NAND2_X1 U9855 ( .A1(b_23_), .A2(a_16_), .ZN(n9924) );
  XOR2_X1 U9856 ( .A(n9925), .B(n9926), .Z(n9680) );
  XOR2_X1 U9857 ( .A(n9927), .B(n9928), .Z(n9926) );
  NAND2_X1 U9858 ( .A1(b_23_), .A2(a_15_), .ZN(n9928) );
  XOR2_X1 U9859 ( .A(n9929), .B(n9930), .Z(n9684) );
  NAND2_X1 U9860 ( .A1(n9931), .A2(n9932), .ZN(n9929) );
  XOR2_X1 U9861 ( .A(n9933), .B(n9934), .Z(n9687) );
  XOR2_X1 U9862 ( .A(n9935), .B(n9936), .Z(n9933) );
  XOR2_X1 U9863 ( .A(n9937), .B(n9938), .Z(n9695) );
  XOR2_X1 U9864 ( .A(n9939), .B(n9940), .Z(n9937) );
  NOR2_X1 U9865 ( .A1(n7724), .A2(n7549), .ZN(n9940) );
  XNOR2_X1 U9866 ( .A(n9941), .B(n9942), .ZN(n9699) );
  NAND2_X1 U9867 ( .A1(n9943), .A2(n9944), .ZN(n9941) );
  XOR2_X1 U9868 ( .A(n9945), .B(n9946), .Z(n9704) );
  XNOR2_X1 U9869 ( .A(n9947), .B(n9948), .ZN(n9946) );
  OR2_X1 U9870 ( .A1(n9714), .A2(n9713), .ZN(n9779) );
  XNOR2_X1 U9871 ( .A(n9949), .B(n9950), .ZN(n9713) );
  XOR2_X1 U9872 ( .A(n9951), .B(n9952), .Z(n9949) );
  NOR2_X1 U9873 ( .A1(n7787), .A2(n7549), .ZN(n9952) );
  NAND2_X1 U9874 ( .A1(b_24_), .A2(a_6_), .ZN(n9714) );
  XNOR2_X1 U9875 ( .A(n9953), .B(n9954), .ZN(n9716) );
  NAND2_X1 U9876 ( .A1(n9955), .A2(n9956), .ZN(n9953) );
  XOR2_X1 U9877 ( .A(n9957), .B(n9958), .Z(n9721) );
  XOR2_X1 U9878 ( .A(n9959), .B(n9960), .Z(n9958) );
  NAND2_X1 U9879 ( .A1(b_23_), .A2(a_5_), .ZN(n9960) );
  INV_X1 U9880 ( .A(n8169), .ZN(n8164) );
  XOR2_X1 U9881 ( .A(n9961), .B(n9962), .Z(n8169) );
  XNOR2_X1 U9882 ( .A(n9963), .B(n9964), .ZN(n9961) );
  NOR2_X1 U9883 ( .A1(n8197), .A2(n7549), .ZN(n9964) );
  NAND3_X1 U9884 ( .A1(n9965), .A2(n8160), .A3(n8159), .ZN(n8021) );
  XNOR2_X1 U9885 ( .A(n9966), .B(n9967), .ZN(n8159) );
  NAND2_X1 U9886 ( .A1(n9968), .A2(n9969), .ZN(n9966) );
  NAND2_X1 U9887 ( .A1(n9970), .A2(n9971), .ZN(n8160) );
  NAND3_X1 U9888 ( .A1(a_0_), .A2(n9972), .A3(b_23_), .ZN(n9971) );
  NAND2_X1 U9889 ( .A1(n9963), .A2(n9962), .ZN(n9972) );
  OR2_X1 U9890 ( .A1(n9962), .A2(n9963), .ZN(n9970) );
  AND2_X1 U9891 ( .A1(n9973), .A2(n9974), .ZN(n9963) );
  NAND3_X1 U9892 ( .A1(a_1_), .A2(n9975), .A3(b_23_), .ZN(n9974) );
  OR2_X1 U9893 ( .A1(n9747), .A2(n9745), .ZN(n9975) );
  NAND2_X1 U9894 ( .A1(n9745), .A2(n9747), .ZN(n9973) );
  NAND2_X1 U9895 ( .A1(n9976), .A2(n9977), .ZN(n9747) );
  NAND3_X1 U9896 ( .A1(a_2_), .A2(n9978), .A3(b_23_), .ZN(n9977) );
  NAND2_X1 U9897 ( .A1(n9755), .A2(n9754), .ZN(n9978) );
  OR2_X1 U9898 ( .A1(n9754), .A2(n9755), .ZN(n9976) );
  AND2_X1 U9899 ( .A1(n9979), .A2(n9980), .ZN(n9755) );
  NAND3_X1 U9900 ( .A1(a_3_), .A2(n9981), .A3(b_23_), .ZN(n9980) );
  OR2_X1 U9901 ( .A1(n9763), .A2(n9761), .ZN(n9981) );
  NAND2_X1 U9902 ( .A1(n9761), .A2(n9763), .ZN(n9979) );
  NAND2_X1 U9903 ( .A1(n9982), .A2(n9983), .ZN(n9763) );
  NAND3_X1 U9904 ( .A1(a_4_), .A2(n9984), .A3(b_23_), .ZN(n9983) );
  OR2_X1 U9905 ( .A1(n9771), .A2(n9769), .ZN(n9984) );
  NAND2_X1 U9906 ( .A1(n9769), .A2(n9771), .ZN(n9982) );
  NAND2_X1 U9907 ( .A1(n9985), .A2(n9986), .ZN(n9771) );
  NAND3_X1 U9908 ( .A1(a_5_), .A2(n9987), .A3(b_23_), .ZN(n9986) );
  OR2_X1 U9909 ( .A1(n9959), .A2(n9957), .ZN(n9987) );
  NAND2_X1 U9910 ( .A1(n9957), .A2(n9959), .ZN(n9985) );
  NAND2_X1 U9911 ( .A1(n9955), .A2(n9988), .ZN(n9959) );
  NAND2_X1 U9912 ( .A1(n9954), .A2(n9956), .ZN(n9988) );
  NAND2_X1 U9913 ( .A1(n9989), .A2(n9990), .ZN(n9956) );
  NAND2_X1 U9914 ( .A1(b_23_), .A2(a_6_), .ZN(n9990) );
  INV_X1 U9915 ( .A(n9991), .ZN(n9989) );
  XNOR2_X1 U9916 ( .A(n9992), .B(n9993), .ZN(n9954) );
  XNOR2_X1 U9917 ( .A(n9994), .B(n9995), .ZN(n9993) );
  NAND2_X1 U9918 ( .A1(a_6_), .A2(n9991), .ZN(n9955) );
  NAND2_X1 U9919 ( .A1(n9996), .A2(n9997), .ZN(n9991) );
  NAND3_X1 U9920 ( .A1(a_7_), .A2(n9998), .A3(b_23_), .ZN(n9997) );
  OR2_X1 U9921 ( .A1(n9951), .A2(n9950), .ZN(n9998) );
  NAND2_X1 U9922 ( .A1(n9950), .A2(n9951), .ZN(n9996) );
  NAND2_X1 U9923 ( .A1(n9999), .A2(n10000), .ZN(n9951) );
  NAND2_X1 U9924 ( .A1(n9789), .A2(n10001), .ZN(n10000) );
  OR2_X1 U9925 ( .A1(n9788), .A2(n9786), .ZN(n10001) );
  NOR2_X1 U9926 ( .A1(n7549), .A2(n8602), .ZN(n9789) );
  NAND2_X1 U9927 ( .A1(n9786), .A2(n9788), .ZN(n9999) );
  NAND2_X1 U9928 ( .A1(n10002), .A2(n10003), .ZN(n9788) );
  NAND2_X1 U9929 ( .A1(n9948), .A2(n10004), .ZN(n10003) );
  OR2_X1 U9930 ( .A1(n9947), .A2(n9945), .ZN(n10004) );
  NOR2_X1 U9931 ( .A1(n7549), .A2(n7753), .ZN(n9948) );
  NAND2_X1 U9932 ( .A1(n9945), .A2(n9947), .ZN(n10002) );
  NAND2_X1 U9933 ( .A1(n9943), .A2(n10005), .ZN(n9947) );
  NAND2_X1 U9934 ( .A1(n9942), .A2(n9944), .ZN(n10005) );
  NAND2_X1 U9935 ( .A1(n10006), .A2(n10007), .ZN(n9944) );
  NAND2_X1 U9936 ( .A1(b_23_), .A2(a_10_), .ZN(n10007) );
  INV_X1 U9937 ( .A(n10008), .ZN(n10006) );
  XNOR2_X1 U9938 ( .A(n10009), .B(n10010), .ZN(n9942) );
  XNOR2_X1 U9939 ( .A(n10011), .B(n10012), .ZN(n10010) );
  NAND2_X1 U9940 ( .A1(a_10_), .A2(n10008), .ZN(n9943) );
  NAND2_X1 U9941 ( .A1(n10013), .A2(n10014), .ZN(n10008) );
  NAND3_X1 U9942 ( .A1(a_11_), .A2(n10015), .A3(b_23_), .ZN(n10014) );
  OR2_X1 U9943 ( .A1(n9939), .A2(n9938), .ZN(n10015) );
  NAND2_X1 U9944 ( .A1(n9938), .A2(n9939), .ZN(n10013) );
  NAND2_X1 U9945 ( .A1(n10016), .A2(n10017), .ZN(n9939) );
  NAND3_X1 U9946 ( .A1(a_12_), .A2(n10018), .A3(b_23_), .ZN(n10017) );
  NAND2_X1 U9947 ( .A1(n9805), .A2(n9804), .ZN(n10018) );
  OR2_X1 U9948 ( .A1(n9804), .A2(n9805), .ZN(n10016) );
  AND2_X1 U9949 ( .A1(n10019), .A2(n10020), .ZN(n9805) );
  NAND2_X1 U9950 ( .A1(n9936), .A2(n10021), .ZN(n10020) );
  OR2_X1 U9951 ( .A1(n9935), .A2(n9934), .ZN(n10021) );
  NOR2_X1 U9952 ( .A1(n7549), .A2(n7702), .ZN(n9936) );
  NAND2_X1 U9953 ( .A1(n9934), .A2(n9935), .ZN(n10019) );
  NAND2_X1 U9954 ( .A1(n9931), .A2(n10022), .ZN(n9935) );
  NAND2_X1 U9955 ( .A1(n9930), .A2(n9932), .ZN(n10022) );
  NAND2_X1 U9956 ( .A1(n10023), .A2(n10024), .ZN(n9932) );
  NAND2_X1 U9957 ( .A1(b_23_), .A2(a_14_), .ZN(n10024) );
  INV_X1 U9958 ( .A(n10025), .ZN(n10023) );
  XOR2_X1 U9959 ( .A(n10026), .B(n10027), .Z(n9930) );
  XOR2_X1 U9960 ( .A(n10028), .B(n10029), .Z(n10026) );
  NAND2_X1 U9961 ( .A1(a_14_), .A2(n10025), .ZN(n9931) );
  NAND2_X1 U9962 ( .A1(n10030), .A2(n10031), .ZN(n10025) );
  NAND3_X1 U9963 ( .A1(a_15_), .A2(n10032), .A3(b_23_), .ZN(n10031) );
  OR2_X1 U9964 ( .A1(n9927), .A2(n9925), .ZN(n10032) );
  NAND2_X1 U9965 ( .A1(n9925), .A2(n9927), .ZN(n10030) );
  NAND2_X1 U9966 ( .A1(n10033), .A2(n10034), .ZN(n9927) );
  NAND3_X1 U9967 ( .A1(a_16_), .A2(n10035), .A3(b_23_), .ZN(n10034) );
  OR2_X1 U9968 ( .A1(n9923), .A2(n9921), .ZN(n10035) );
  NAND2_X1 U9969 ( .A1(n9921), .A2(n9923), .ZN(n10033) );
  NAND2_X1 U9970 ( .A1(n10036), .A2(n10037), .ZN(n9923) );
  NAND2_X1 U9971 ( .A1(n9920), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U9972 ( .A1(n9919), .A2(n9918), .ZN(n10038) );
  NOR2_X1 U9973 ( .A1(n7549), .A2(n7645), .ZN(n9920) );
  OR2_X1 U9974 ( .A1(n9918), .A2(n9919), .ZN(n10036) );
  AND2_X1 U9975 ( .A1(n10039), .A2(n10040), .ZN(n9919) );
  NAND3_X1 U9976 ( .A1(a_18_), .A2(n10041), .A3(b_23_), .ZN(n10040) );
  NAND2_X1 U9977 ( .A1(n9915), .A2(n9914), .ZN(n10041) );
  OR2_X1 U9978 ( .A1(n9914), .A2(n9915), .ZN(n10039) );
  AND2_X1 U9979 ( .A1(n10042), .A2(n10043), .ZN(n9915) );
  NAND2_X1 U9980 ( .A1(n9912), .A2(n10044), .ZN(n10043) );
  OR2_X1 U9981 ( .A1(n9911), .A2(n9909), .ZN(n10044) );
  NOR2_X1 U9982 ( .A1(n7549), .A2(n7958), .ZN(n9912) );
  NAND2_X1 U9983 ( .A1(n9909), .A2(n9911), .ZN(n10042) );
  NAND2_X1 U9984 ( .A1(n10045), .A2(n10046), .ZN(n9911) );
  NAND3_X1 U9985 ( .A1(a_20_), .A2(n10047), .A3(b_23_), .ZN(n10046) );
  NAND2_X1 U9986 ( .A1(n9907), .A2(n9906), .ZN(n10047) );
  OR2_X1 U9987 ( .A1(n9906), .A2(n9907), .ZN(n10045) );
  AND2_X1 U9988 ( .A1(n10048), .A2(n10049), .ZN(n9907) );
  NAND2_X1 U9989 ( .A1(n9904), .A2(n10050), .ZN(n10049) );
  OR2_X1 U9990 ( .A1(n9903), .A2(n9902), .ZN(n10050) );
  NOR2_X1 U9991 ( .A1(n7549), .A2(n7578), .ZN(n9904) );
  NAND2_X1 U9992 ( .A1(n9902), .A2(n9903), .ZN(n10048) );
  NAND2_X1 U9993 ( .A1(n10051), .A2(n10052), .ZN(n9903) );
  NAND3_X1 U9994 ( .A1(a_22_), .A2(n10053), .A3(b_23_), .ZN(n10052) );
  OR2_X1 U9995 ( .A1(n9899), .A2(n9897), .ZN(n10053) );
  NAND2_X1 U9996 ( .A1(n9897), .A2(n9899), .ZN(n10051) );
  NAND2_X1 U9997 ( .A1(n10054), .A2(n10055), .ZN(n9899) );
  NAND2_X1 U9998 ( .A1(n7547), .A2(n10056), .ZN(n10055) );
  OR2_X1 U9999 ( .A1(n9896), .A2(n9894), .ZN(n10056) );
  NOR2_X1 U10000 ( .A1(n7549), .A2(n7955), .ZN(n7547) );
  NAND2_X1 U10001 ( .A1(n9894), .A2(n9896), .ZN(n10054) );
  NAND2_X1 U10002 ( .A1(n10057), .A2(n10058), .ZN(n9896) );
  NAND3_X1 U10003 ( .A1(a_24_), .A2(n10059), .A3(b_23_), .ZN(n10058) );
  NAND2_X1 U10004 ( .A1(n9892), .A2(n9891), .ZN(n10059) );
  OR2_X1 U10005 ( .A1(n9891), .A2(n9892), .ZN(n10057) );
  AND2_X1 U10006 ( .A1(n10060), .A2(n10061), .ZN(n9892) );
  NAND2_X1 U10007 ( .A1(n9849), .A2(n10062), .ZN(n10061) );
  OR2_X1 U10008 ( .A1(n9848), .A2(n9847), .ZN(n10062) );
  NOR2_X1 U10009 ( .A1(n7549), .A2(n7952), .ZN(n9849) );
  NAND2_X1 U10010 ( .A1(n9847), .A2(n9848), .ZN(n10060) );
  NAND2_X1 U10011 ( .A1(n9888), .A2(n10063), .ZN(n9848) );
  NAND2_X1 U10012 ( .A1(n9887), .A2(n9889), .ZN(n10063) );
  NAND2_X1 U10013 ( .A1(n10064), .A2(n10065), .ZN(n9889) );
  NAND2_X1 U10014 ( .A1(b_23_), .A2(a_26_), .ZN(n10065) );
  INV_X1 U10015 ( .A(n10066), .ZN(n10064) );
  XNOR2_X1 U10016 ( .A(n10067), .B(n10068), .ZN(n9887) );
  NAND2_X1 U10017 ( .A1(n10069), .A2(n10070), .ZN(n10067) );
  NAND2_X1 U10018 ( .A1(a_26_), .A2(n10066), .ZN(n9888) );
  NAND2_X1 U10019 ( .A1(n9859), .A2(n10071), .ZN(n10066) );
  NAND2_X1 U10020 ( .A1(n9858), .A2(n9860), .ZN(n10071) );
  NAND2_X1 U10021 ( .A1(n10072), .A2(n10073), .ZN(n9860) );
  NAND2_X1 U10022 ( .A1(b_23_), .A2(a_27_), .ZN(n10073) );
  INV_X1 U10023 ( .A(n10074), .ZN(n10072) );
  XNOR2_X1 U10024 ( .A(n10075), .B(n10076), .ZN(n9858) );
  XOR2_X1 U10025 ( .A(n10077), .B(n10078), .Z(n10075) );
  NAND2_X1 U10026 ( .A1(b_22_), .A2(a_28_), .ZN(n10077) );
  NAND2_X1 U10027 ( .A1(a_27_), .A2(n10074), .ZN(n9859) );
  NAND2_X1 U10028 ( .A1(n10079), .A2(n10080), .ZN(n10074) );
  NAND3_X1 U10029 ( .A1(a_28_), .A2(n10081), .A3(b_23_), .ZN(n10080) );
  NAND2_X1 U10030 ( .A1(n9868), .A2(n9866), .ZN(n10081) );
  OR2_X1 U10031 ( .A1(n9866), .A2(n9868), .ZN(n10079) );
  AND2_X1 U10032 ( .A1(n10082), .A2(n10083), .ZN(n9868) );
  NAND2_X1 U10033 ( .A1(n9883), .A2(n10084), .ZN(n10083) );
  OR2_X1 U10034 ( .A1(n9884), .A2(n9885), .ZN(n10084) );
  NOR2_X1 U10035 ( .A1(n7549), .A2(n7460), .ZN(n9883) );
  INV_X1 U10036 ( .A(b_23_), .ZN(n7549) );
  NAND2_X1 U10037 ( .A1(n9885), .A2(n9884), .ZN(n10082) );
  NAND2_X1 U10038 ( .A1(n10085), .A2(n10086), .ZN(n9884) );
  NAND2_X1 U10039 ( .A1(b_21_), .A2(n10087), .ZN(n10086) );
  NAND2_X1 U10040 ( .A1(n7441), .A2(n10088), .ZN(n10087) );
  NAND2_X1 U10041 ( .A1(a_31_), .A2(n9881), .ZN(n10088) );
  NAND2_X1 U10042 ( .A1(b_22_), .A2(n10089), .ZN(n10085) );
  NAND2_X1 U10043 ( .A1(n7445), .A2(n10090), .ZN(n10089) );
  NAND2_X1 U10044 ( .A1(a_30_), .A2(n7580), .ZN(n10090) );
  AND3_X1 U10045 ( .A1(b_22_), .A2(n7409), .A3(b_23_), .ZN(n9885) );
  XNOR2_X1 U10046 ( .A(n10091), .B(n10092), .ZN(n9866) );
  XOR2_X1 U10047 ( .A(n10093), .B(n10094), .Z(n10091) );
  XNOR2_X1 U10048 ( .A(n10095), .B(n10096), .ZN(n9847) );
  NAND2_X1 U10049 ( .A1(n10097), .A2(n10098), .ZN(n10095) );
  XNOR2_X1 U10050 ( .A(n10099), .B(n10100), .ZN(n9891) );
  XOR2_X1 U10051 ( .A(n10101), .B(n10102), .Z(n10099) );
  XNOR2_X1 U10052 ( .A(n10103), .B(n10104), .ZN(n9894) );
  XNOR2_X1 U10053 ( .A(n10105), .B(n10106), .ZN(n10103) );
  NOR2_X1 U10054 ( .A1(n7954), .A2(n9881), .ZN(n10106) );
  XNOR2_X1 U10055 ( .A(n10107), .B(n10108), .ZN(n9897) );
  XNOR2_X1 U10056 ( .A(n10109), .B(n10110), .ZN(n10108) );
  XNOR2_X1 U10057 ( .A(n10111), .B(n10112), .ZN(n9902) );
  XNOR2_X1 U10058 ( .A(n10113), .B(n7562), .ZN(n10112) );
  XNOR2_X1 U10059 ( .A(n10114), .B(n10115), .ZN(n9906) );
  XOR2_X1 U10060 ( .A(n10116), .B(n10117), .Z(n10114) );
  XNOR2_X1 U10061 ( .A(n10118), .B(n10119), .ZN(n9909) );
  XNOR2_X1 U10062 ( .A(n10120), .B(n10121), .ZN(n10118) );
  NOR2_X1 U10063 ( .A1(n7957), .A2(n9881), .ZN(n10121) );
  XOR2_X1 U10064 ( .A(n10122), .B(n10123), .Z(n9914) );
  XNOR2_X1 U10065 ( .A(n10124), .B(n10125), .ZN(n10123) );
  XNOR2_X1 U10066 ( .A(n10126), .B(n10127), .ZN(n9918) );
  XOR2_X1 U10067 ( .A(n10128), .B(n10129), .Z(n10126) );
  NOR2_X1 U10068 ( .A1(n7960), .A2(n9881), .ZN(n10129) );
  XOR2_X1 U10069 ( .A(n10130), .B(n10131), .Z(n9921) );
  XOR2_X1 U10070 ( .A(n10132), .B(n10133), .Z(n10130) );
  XNOR2_X1 U10071 ( .A(n10134), .B(n10135), .ZN(n9925) );
  XOR2_X1 U10072 ( .A(n10136), .B(n10137), .Z(n10135) );
  NAND2_X1 U10073 ( .A1(b_22_), .A2(a_16_), .ZN(n10137) );
  XNOR2_X1 U10074 ( .A(n10138), .B(n10139), .ZN(n9934) );
  XNOR2_X1 U10075 ( .A(n10140), .B(n10141), .ZN(n10138) );
  NOR2_X1 U10076 ( .A1(n7962), .A2(n9881), .ZN(n10141) );
  XOR2_X1 U10077 ( .A(n10142), .B(n10143), .Z(n9804) );
  XNOR2_X1 U10078 ( .A(n10144), .B(n10145), .ZN(n10143) );
  XNOR2_X1 U10079 ( .A(n10146), .B(n10147), .ZN(n9938) );
  XNOR2_X1 U10080 ( .A(n10148), .B(n10149), .ZN(n10146) );
  NOR2_X1 U10081 ( .A1(n8585), .A2(n9881), .ZN(n10149) );
  XNOR2_X1 U10082 ( .A(n10150), .B(n10151), .ZN(n9945) );
  XNOR2_X1 U10083 ( .A(n10152), .B(n10153), .ZN(n10150) );
  NOR2_X1 U10084 ( .A1(n8378), .A2(n9881), .ZN(n10153) );
  XNOR2_X1 U10085 ( .A(n10154), .B(n10155), .ZN(n9786) );
  XOR2_X1 U10086 ( .A(n10156), .B(n10157), .Z(n10155) );
  NAND2_X1 U10087 ( .A1(b_22_), .A2(a_9_), .ZN(n10157) );
  XNOR2_X1 U10088 ( .A(n10158), .B(n10159), .ZN(n9950) );
  XNOR2_X1 U10089 ( .A(n10160), .B(n10161), .ZN(n10158) );
  XNOR2_X1 U10090 ( .A(n10162), .B(n10163), .ZN(n9957) );
  XNOR2_X1 U10091 ( .A(n10164), .B(n10165), .ZN(n10162) );
  NOR2_X1 U10092 ( .A1(n7807), .A2(n9881), .ZN(n10165) );
  XNOR2_X1 U10093 ( .A(n10166), .B(n10167), .ZN(n9769) );
  XNOR2_X1 U10094 ( .A(n10168), .B(n10169), .ZN(n10167) );
  XOR2_X1 U10095 ( .A(n10170), .B(n10171), .Z(n9761) );
  XOR2_X1 U10096 ( .A(n10172), .B(n10173), .Z(n10170) );
  XNOR2_X1 U10097 ( .A(n10174), .B(n10175), .ZN(n9754) );
  XOR2_X1 U10098 ( .A(n10176), .B(n10177), .Z(n10174) );
  XOR2_X1 U10099 ( .A(n10178), .B(n10179), .Z(n9745) );
  XOR2_X1 U10100 ( .A(n10180), .B(n10181), .Z(n10178) );
  XNOR2_X1 U10101 ( .A(n10182), .B(n10183), .ZN(n9962) );
  XOR2_X1 U10102 ( .A(n10184), .B(n10185), .Z(n10182) );
  NOR2_X1 U10103 ( .A1(n7872), .A2(n9881), .ZN(n10185) );
  XOR2_X1 U10104 ( .A(n8155), .B(n8154), .Z(n9965) );
  NAND4_X1 U10105 ( .A1(n8154), .A2(n8153), .A3(n8155), .A4(n8149), .ZN(n8027)
         );
  INV_X1 U10106 ( .A(n10186), .ZN(n8149) );
  NAND2_X1 U10107 ( .A1(n9968), .A2(n10187), .ZN(n8155) );
  NAND2_X1 U10108 ( .A1(n9967), .A2(n9969), .ZN(n10187) );
  NAND2_X1 U10109 ( .A1(n10188), .A2(n10189), .ZN(n9969) );
  NAND2_X1 U10110 ( .A1(b_22_), .A2(a_0_), .ZN(n10189) );
  INV_X1 U10111 ( .A(n10190), .ZN(n10188) );
  XOR2_X1 U10112 ( .A(n10191), .B(n10192), .Z(n9967) );
  XOR2_X1 U10113 ( .A(n10193), .B(n10194), .Z(n10191) );
  NOR2_X1 U10114 ( .A1(n7872), .A2(n7580), .ZN(n10194) );
  NAND2_X1 U10115 ( .A1(a_0_), .A2(n10190), .ZN(n9968) );
  NAND2_X1 U10116 ( .A1(n10195), .A2(n10196), .ZN(n10190) );
  NAND3_X1 U10117 ( .A1(a_1_), .A2(n10197), .A3(b_22_), .ZN(n10196) );
  OR2_X1 U10118 ( .A1(n10184), .A2(n10183), .ZN(n10197) );
  NAND2_X1 U10119 ( .A1(n10183), .A2(n10184), .ZN(n10195) );
  NAND2_X1 U10120 ( .A1(n10198), .A2(n10199), .ZN(n10184) );
  NAND2_X1 U10121 ( .A1(n10181), .A2(n10200), .ZN(n10199) );
  OR2_X1 U10122 ( .A1(n10180), .A2(n10179), .ZN(n10200) );
  NOR2_X1 U10123 ( .A1(n9881), .A2(n7966), .ZN(n10181) );
  NAND2_X1 U10124 ( .A1(n10179), .A2(n10180), .ZN(n10198) );
  NAND2_X1 U10125 ( .A1(n10201), .A2(n10202), .ZN(n10180) );
  NAND2_X1 U10126 ( .A1(n10177), .A2(n10203), .ZN(n10202) );
  OR2_X1 U10127 ( .A1(n10176), .A2(n10175), .ZN(n10203) );
  NOR2_X1 U10128 ( .A1(n9881), .A2(n7852), .ZN(n10177) );
  NAND2_X1 U10129 ( .A1(n10175), .A2(n10176), .ZN(n10201) );
  NAND2_X1 U10130 ( .A1(n10204), .A2(n10205), .ZN(n10176) );
  NAND2_X1 U10131 ( .A1(n10173), .A2(n10206), .ZN(n10205) );
  OR2_X1 U10132 ( .A1(n10172), .A2(n10171), .ZN(n10206) );
  NOR2_X1 U10133 ( .A1(n9881), .A2(n7836), .ZN(n10173) );
  NAND2_X1 U10134 ( .A1(n10171), .A2(n10172), .ZN(n10204) );
  NAND2_X1 U10135 ( .A1(n10207), .A2(n10208), .ZN(n10172) );
  NAND2_X1 U10136 ( .A1(n10169), .A2(n10209), .ZN(n10208) );
  OR2_X1 U10137 ( .A1(n10168), .A2(n10166), .ZN(n10209) );
  NOR2_X1 U10138 ( .A1(n9881), .A2(n7823), .ZN(n10169) );
  NAND2_X1 U10139 ( .A1(n10166), .A2(n10168), .ZN(n10207) );
  NAND2_X1 U10140 ( .A1(n10210), .A2(n10211), .ZN(n10168) );
  NAND3_X1 U10141 ( .A1(a_6_), .A2(n10212), .A3(b_22_), .ZN(n10211) );
  NAND2_X1 U10142 ( .A1(n10164), .A2(n10163), .ZN(n10212) );
  OR2_X1 U10143 ( .A1(n10163), .A2(n10164), .ZN(n10210) );
  AND2_X1 U10144 ( .A1(n10213), .A2(n10214), .ZN(n10164) );
  NAND2_X1 U10145 ( .A1(n9995), .A2(n10215), .ZN(n10214) );
  OR2_X1 U10146 ( .A1(n9994), .A2(n9992), .ZN(n10215) );
  NOR2_X1 U10147 ( .A1(n9881), .A2(n7787), .ZN(n9995) );
  NAND2_X1 U10148 ( .A1(n9992), .A2(n9994), .ZN(n10213) );
  NAND2_X1 U10149 ( .A1(n10216), .A2(n10217), .ZN(n9994) );
  NAND2_X1 U10150 ( .A1(n10161), .A2(n10218), .ZN(n10217) );
  NAND2_X1 U10151 ( .A1(n10160), .A2(n10159), .ZN(n10218) );
  NOR2_X1 U10152 ( .A1(n9881), .A2(n8602), .ZN(n10161) );
  OR2_X1 U10153 ( .A1(n10159), .A2(n10160), .ZN(n10216) );
  AND2_X1 U10154 ( .A1(n10219), .A2(n10220), .ZN(n10160) );
  NAND3_X1 U10155 ( .A1(a_9_), .A2(n10221), .A3(b_22_), .ZN(n10220) );
  OR2_X1 U10156 ( .A1(n10156), .A2(n10154), .ZN(n10221) );
  NAND2_X1 U10157 ( .A1(n10154), .A2(n10156), .ZN(n10219) );
  NAND2_X1 U10158 ( .A1(n10222), .A2(n10223), .ZN(n10156) );
  NAND3_X1 U10159 ( .A1(a_10_), .A2(n10224), .A3(b_22_), .ZN(n10223) );
  NAND2_X1 U10160 ( .A1(n10152), .A2(n10151), .ZN(n10224) );
  OR2_X1 U10161 ( .A1(n10151), .A2(n10152), .ZN(n10222) );
  AND2_X1 U10162 ( .A1(n10225), .A2(n10226), .ZN(n10152) );
  NAND2_X1 U10163 ( .A1(n10012), .A2(n10227), .ZN(n10226) );
  OR2_X1 U10164 ( .A1(n10011), .A2(n10009), .ZN(n10227) );
  NOR2_X1 U10165 ( .A1(n9881), .A2(n7724), .ZN(n10012) );
  NAND2_X1 U10166 ( .A1(n10009), .A2(n10011), .ZN(n10225) );
  NAND2_X1 U10167 ( .A1(n10228), .A2(n10229), .ZN(n10011) );
  NAND3_X1 U10168 ( .A1(a_12_), .A2(n10230), .A3(b_22_), .ZN(n10229) );
  NAND2_X1 U10169 ( .A1(n10148), .A2(n10147), .ZN(n10230) );
  OR2_X1 U10170 ( .A1(n10147), .A2(n10148), .ZN(n10228) );
  AND2_X1 U10171 ( .A1(n10231), .A2(n10232), .ZN(n10148) );
  NAND2_X1 U10172 ( .A1(n10145), .A2(n10233), .ZN(n10232) );
  OR2_X1 U10173 ( .A1(n10144), .A2(n10142), .ZN(n10233) );
  NOR2_X1 U10174 ( .A1(n9881), .A2(n7702), .ZN(n10145) );
  NAND2_X1 U10175 ( .A1(n10142), .A2(n10144), .ZN(n10231) );
  NAND2_X1 U10176 ( .A1(n10234), .A2(n10235), .ZN(n10144) );
  NAND3_X1 U10177 ( .A1(a_14_), .A2(n10236), .A3(b_22_), .ZN(n10235) );
  NAND2_X1 U10178 ( .A1(n10140), .A2(n10139), .ZN(n10236) );
  OR2_X1 U10179 ( .A1(n10139), .A2(n10140), .ZN(n10234) );
  AND2_X1 U10180 ( .A1(n10237), .A2(n10238), .ZN(n10140) );
  NAND2_X1 U10181 ( .A1(n10029), .A2(n10239), .ZN(n10238) );
  OR2_X1 U10182 ( .A1(n10028), .A2(n10027), .ZN(n10239) );
  NOR2_X1 U10183 ( .A1(n9881), .A2(n7667), .ZN(n10029) );
  NAND2_X1 U10184 ( .A1(n10027), .A2(n10028), .ZN(n10237) );
  NAND2_X1 U10185 ( .A1(n10240), .A2(n10241), .ZN(n10028) );
  NAND3_X1 U10186 ( .A1(a_16_), .A2(n10242), .A3(b_22_), .ZN(n10241) );
  OR2_X1 U10187 ( .A1(n10136), .A2(n10134), .ZN(n10242) );
  NAND2_X1 U10188 ( .A1(n10134), .A2(n10136), .ZN(n10240) );
  NAND2_X1 U10189 ( .A1(n10243), .A2(n10244), .ZN(n10136) );
  NAND2_X1 U10190 ( .A1(n10133), .A2(n10245), .ZN(n10244) );
  OR2_X1 U10191 ( .A1(n10132), .A2(n10131), .ZN(n10245) );
  NOR2_X1 U10192 ( .A1(n9881), .A2(n7645), .ZN(n10133) );
  NAND2_X1 U10193 ( .A1(n10131), .A2(n10132), .ZN(n10243) );
  NAND2_X1 U10194 ( .A1(n10246), .A2(n10247), .ZN(n10132) );
  NAND3_X1 U10195 ( .A1(a_18_), .A2(n10248), .A3(b_22_), .ZN(n10247) );
  OR2_X1 U10196 ( .A1(n10128), .A2(n10127), .ZN(n10248) );
  NAND2_X1 U10197 ( .A1(n10127), .A2(n10128), .ZN(n10246) );
  NAND2_X1 U10198 ( .A1(n10249), .A2(n10250), .ZN(n10128) );
  NAND2_X1 U10199 ( .A1(n10125), .A2(n10251), .ZN(n10250) );
  OR2_X1 U10200 ( .A1(n10124), .A2(n10122), .ZN(n10251) );
  NOR2_X1 U10201 ( .A1(n9881), .A2(n7958), .ZN(n10125) );
  NAND2_X1 U10202 ( .A1(n10122), .A2(n10124), .ZN(n10249) );
  NAND2_X1 U10203 ( .A1(n10252), .A2(n10253), .ZN(n10124) );
  NAND3_X1 U10204 ( .A1(a_20_), .A2(n10254), .A3(b_22_), .ZN(n10253) );
  NAND2_X1 U10205 ( .A1(n10120), .A2(n10119), .ZN(n10254) );
  OR2_X1 U10206 ( .A1(n10119), .A2(n10120), .ZN(n10252) );
  AND2_X1 U10207 ( .A1(n10255), .A2(n10256), .ZN(n10120) );
  NAND2_X1 U10208 ( .A1(n10117), .A2(n10257), .ZN(n10256) );
  OR2_X1 U10209 ( .A1(n10116), .A2(n10115), .ZN(n10257) );
  NOR2_X1 U10210 ( .A1(n9881), .A2(n7578), .ZN(n10117) );
  NAND2_X1 U10211 ( .A1(n10115), .A2(n10116), .ZN(n10255) );
  NAND2_X1 U10212 ( .A1(n10258), .A2(n10259), .ZN(n10116) );
  NAND2_X1 U10213 ( .A1(n10111), .A2(n10260), .ZN(n10259) );
  OR2_X1 U10214 ( .A1(n10113), .A2(n7562), .ZN(n10260) );
  XNOR2_X1 U10215 ( .A(n10261), .B(n10262), .ZN(n10111) );
  XNOR2_X1 U10216 ( .A(n10263), .B(n10264), .ZN(n10262) );
  NAND2_X1 U10217 ( .A1(n7562), .A2(n10113), .ZN(n10258) );
  NAND2_X1 U10218 ( .A1(n10265), .A2(n10266), .ZN(n10113) );
  NAND2_X1 U10219 ( .A1(n10110), .A2(n10267), .ZN(n10266) );
  OR2_X1 U10220 ( .A1(n10109), .A2(n10107), .ZN(n10267) );
  NOR2_X1 U10221 ( .A1(n9881), .A2(n7955), .ZN(n10110) );
  NAND2_X1 U10222 ( .A1(n10107), .A2(n10109), .ZN(n10265) );
  NAND2_X1 U10223 ( .A1(n10268), .A2(n10269), .ZN(n10109) );
  NAND3_X1 U10224 ( .A1(a_24_), .A2(n10270), .A3(b_22_), .ZN(n10269) );
  NAND2_X1 U10225 ( .A1(n10105), .A2(n10104), .ZN(n10270) );
  OR2_X1 U10226 ( .A1(n10104), .A2(n10105), .ZN(n10268) );
  AND2_X1 U10227 ( .A1(n10271), .A2(n10272), .ZN(n10105) );
  NAND2_X1 U10228 ( .A1(n10102), .A2(n10273), .ZN(n10272) );
  OR2_X1 U10229 ( .A1(n10101), .A2(n10100), .ZN(n10273) );
  NOR2_X1 U10230 ( .A1(n9881), .A2(n7952), .ZN(n10102) );
  NAND2_X1 U10231 ( .A1(n10100), .A2(n10101), .ZN(n10271) );
  NAND2_X1 U10232 ( .A1(n10097), .A2(n10274), .ZN(n10101) );
  NAND2_X1 U10233 ( .A1(n10096), .A2(n10098), .ZN(n10274) );
  NAND2_X1 U10234 ( .A1(n10275), .A2(n10276), .ZN(n10098) );
  NAND2_X1 U10235 ( .A1(b_22_), .A2(a_26_), .ZN(n10276) );
  INV_X1 U10236 ( .A(n10277), .ZN(n10275) );
  XNOR2_X1 U10237 ( .A(n10278), .B(n10279), .ZN(n10096) );
  NAND2_X1 U10238 ( .A1(n10280), .A2(n10281), .ZN(n10278) );
  NAND2_X1 U10239 ( .A1(a_26_), .A2(n10277), .ZN(n10097) );
  NAND2_X1 U10240 ( .A1(n10069), .A2(n10282), .ZN(n10277) );
  NAND2_X1 U10241 ( .A1(n10068), .A2(n10070), .ZN(n10282) );
  NAND2_X1 U10242 ( .A1(n10283), .A2(n10284), .ZN(n10070) );
  NAND2_X1 U10243 ( .A1(b_22_), .A2(a_27_), .ZN(n10284) );
  INV_X1 U10244 ( .A(n10285), .ZN(n10283) );
  XNOR2_X1 U10245 ( .A(n10286), .B(n10287), .ZN(n10068) );
  XOR2_X1 U10246 ( .A(n10288), .B(n10289), .Z(n10286) );
  NAND2_X1 U10247 ( .A1(b_21_), .A2(a_28_), .ZN(n10288) );
  NAND2_X1 U10248 ( .A1(a_27_), .A2(n10285), .ZN(n10069) );
  NAND2_X1 U10249 ( .A1(n10290), .A2(n10291), .ZN(n10285) );
  NAND3_X1 U10250 ( .A1(a_28_), .A2(n10292), .A3(b_22_), .ZN(n10291) );
  NAND2_X1 U10251 ( .A1(n10078), .A2(n10076), .ZN(n10292) );
  OR2_X1 U10252 ( .A1(n10076), .A2(n10078), .ZN(n10290) );
  AND2_X1 U10253 ( .A1(n10293), .A2(n10294), .ZN(n10078) );
  NAND2_X1 U10254 ( .A1(n10092), .A2(n10295), .ZN(n10294) );
  OR2_X1 U10255 ( .A1(n10093), .A2(n10094), .ZN(n10295) );
  NOR2_X1 U10256 ( .A1(n9881), .A2(n7460), .ZN(n10092) );
  NAND2_X1 U10257 ( .A1(n10094), .A2(n10093), .ZN(n10293) );
  NAND2_X1 U10258 ( .A1(n10296), .A2(n10297), .ZN(n10093) );
  NAND2_X1 U10259 ( .A1(b_20_), .A2(n10298), .ZN(n10297) );
  NAND2_X1 U10260 ( .A1(n7441), .A2(n10299), .ZN(n10298) );
  NAND2_X1 U10261 ( .A1(a_31_), .A2(n7580), .ZN(n10299) );
  NAND2_X1 U10262 ( .A1(b_21_), .A2(n10300), .ZN(n10296) );
  NAND2_X1 U10263 ( .A1(n7445), .A2(n10301), .ZN(n10300) );
  NAND2_X1 U10264 ( .A1(a_30_), .A2(n7956), .ZN(n10301) );
  AND3_X1 U10265 ( .A1(b_21_), .A2(n7409), .A3(b_22_), .ZN(n10094) );
  XNOR2_X1 U10266 ( .A(n10302), .B(n10303), .ZN(n10076) );
  XOR2_X1 U10267 ( .A(n10304), .B(n10305), .Z(n10302) );
  XNOR2_X1 U10268 ( .A(n10306), .B(n10307), .ZN(n10100) );
  NAND2_X1 U10269 ( .A1(n10308), .A2(n10309), .ZN(n10306) );
  XNOR2_X1 U10270 ( .A(n10310), .B(n10311), .ZN(n10104) );
  XOR2_X1 U10271 ( .A(n10312), .B(n10313), .Z(n10310) );
  XNOR2_X1 U10272 ( .A(n10314), .B(n10315), .ZN(n10107) );
  XNOR2_X1 U10273 ( .A(n10316), .B(n10317), .ZN(n10314) );
  NOR2_X1 U10274 ( .A1(n7954), .A2(n7580), .ZN(n10317) );
  NOR2_X1 U10275 ( .A1(n9881), .A2(n7568), .ZN(n7562) );
  XNOR2_X1 U10276 ( .A(n10318), .B(n10319), .ZN(n10115) );
  XOR2_X1 U10277 ( .A(n10320), .B(n10321), .Z(n10319) );
  NAND2_X1 U10278 ( .A1(b_21_), .A2(a_22_), .ZN(n10321) );
  XNOR2_X1 U10279 ( .A(n10322), .B(n10323), .ZN(n10119) );
  XOR2_X1 U10280 ( .A(n10324), .B(n7575), .Z(n10322) );
  XNOR2_X1 U10281 ( .A(n10325), .B(n10326), .ZN(n10122) );
  XNOR2_X1 U10282 ( .A(n10327), .B(n10328), .ZN(n10325) );
  NOR2_X1 U10283 ( .A1(n7957), .A2(n7580), .ZN(n10328) );
  XNOR2_X1 U10284 ( .A(n10329), .B(n10330), .ZN(n10127) );
  XNOR2_X1 U10285 ( .A(n10331), .B(n10332), .ZN(n10330) );
  XNOR2_X1 U10286 ( .A(n10333), .B(n10334), .ZN(n10131) );
  XNOR2_X1 U10287 ( .A(n10335), .B(n10336), .ZN(n10333) );
  NOR2_X1 U10288 ( .A1(n7960), .A2(n7580), .ZN(n10336) );
  XNOR2_X1 U10289 ( .A(n10337), .B(n10338), .ZN(n10134) );
  XNOR2_X1 U10290 ( .A(n10339), .B(n10340), .ZN(n10338) );
  XNOR2_X1 U10291 ( .A(n10341), .B(n10342), .ZN(n10027) );
  XNOR2_X1 U10292 ( .A(n10343), .B(n10344), .ZN(n10341) );
  NOR2_X1 U10293 ( .A1(n8353), .A2(n7580), .ZN(n10344) );
  XNOR2_X1 U10294 ( .A(n10345), .B(n10346), .ZN(n10139) );
  XOR2_X1 U10295 ( .A(n10347), .B(n10348), .Z(n10345) );
  XNOR2_X1 U10296 ( .A(n10349), .B(n10350), .ZN(n10142) );
  XNOR2_X1 U10297 ( .A(n10351), .B(n10352), .ZN(n10349) );
  NOR2_X1 U10298 ( .A1(n7962), .A2(n7580), .ZN(n10352) );
  XNOR2_X1 U10299 ( .A(n10353), .B(n10354), .ZN(n10147) );
  XOR2_X1 U10300 ( .A(n10355), .B(n10356), .Z(n10353) );
  XNOR2_X1 U10301 ( .A(n10357), .B(n10358), .ZN(n10009) );
  XOR2_X1 U10302 ( .A(n10359), .B(n10360), .Z(n10358) );
  NAND2_X1 U10303 ( .A1(b_21_), .A2(a_12_), .ZN(n10360) );
  XOR2_X1 U10304 ( .A(n10361), .B(n10362), .Z(n10151) );
  XNOR2_X1 U10305 ( .A(n10363), .B(n10364), .ZN(n10362) );
  XOR2_X1 U10306 ( .A(n10365), .B(n10366), .Z(n10154) );
  XOR2_X1 U10307 ( .A(n10367), .B(n10368), .Z(n10365) );
  XNOR2_X1 U10308 ( .A(n10369), .B(n10370), .ZN(n10159) );
  XOR2_X1 U10309 ( .A(n10371), .B(n10372), .Z(n10369) );
  NOR2_X1 U10310 ( .A1(n7753), .A2(n7580), .ZN(n10372) );
  XNOR2_X1 U10311 ( .A(n10373), .B(n10374), .ZN(n9992) );
  XOR2_X1 U10312 ( .A(n10375), .B(n10376), .Z(n10374) );
  NAND2_X1 U10313 ( .A1(b_21_), .A2(a_8_), .ZN(n10376) );
  XOR2_X1 U10314 ( .A(n10377), .B(n10378), .Z(n10163) );
  XOR2_X1 U10315 ( .A(n10379), .B(n10380), .Z(n10378) );
  NAND2_X1 U10316 ( .A1(b_21_), .A2(a_7_), .ZN(n10380) );
  XNOR2_X1 U10317 ( .A(n10381), .B(n10382), .ZN(n10166) );
  XNOR2_X1 U10318 ( .A(n10383), .B(n10384), .ZN(n10381) );
  NOR2_X1 U10319 ( .A1(n7807), .A2(n7580), .ZN(n10384) );
  XNOR2_X1 U10320 ( .A(n10385), .B(n10386), .ZN(n10171) );
  XNOR2_X1 U10321 ( .A(n10387), .B(n10388), .ZN(n10385) );
  NOR2_X1 U10322 ( .A1(n7823), .A2(n7580), .ZN(n10388) );
  XNOR2_X1 U10323 ( .A(n10389), .B(n10390), .ZN(n10175) );
  XOR2_X1 U10324 ( .A(n10391), .B(n10392), .Z(n10390) );
  NAND2_X1 U10325 ( .A1(b_21_), .A2(a_4_), .ZN(n10392) );
  XNOR2_X1 U10326 ( .A(n10393), .B(n10394), .ZN(n10179) );
  XOR2_X1 U10327 ( .A(n10395), .B(n10396), .Z(n10394) );
  NAND2_X1 U10328 ( .A1(b_21_), .A2(a_3_), .ZN(n10396) );
  XNOR2_X1 U10329 ( .A(n10397), .B(n10398), .ZN(n10183) );
  XOR2_X1 U10330 ( .A(n10399), .B(n10400), .Z(n10398) );
  NAND2_X1 U10331 ( .A1(b_21_), .A2(a_2_), .ZN(n10400) );
  NAND2_X1 U10332 ( .A1(n10401), .A2(n10402), .ZN(n8153) );
  XNOR2_X1 U10333 ( .A(n10403), .B(n10404), .ZN(n8154) );
  XNOR2_X1 U10334 ( .A(n10405), .B(n10406), .ZN(n10404) );
  NAND2_X1 U10335 ( .A1(n10407), .A2(n10186), .ZN(n8032) );
  NOR2_X1 U10336 ( .A1(n10402), .A2(n10401), .ZN(n10186) );
  AND2_X1 U10337 ( .A1(n10408), .A2(n10409), .ZN(n10401) );
  NAND2_X1 U10338 ( .A1(n10406), .A2(n10410), .ZN(n10409) );
  OR2_X1 U10339 ( .A1(n10405), .A2(n10403), .ZN(n10410) );
  NOR2_X1 U10340 ( .A1(n7580), .A2(n8197), .ZN(n10406) );
  NAND2_X1 U10341 ( .A1(n10403), .A2(n10405), .ZN(n10408) );
  NAND2_X1 U10342 ( .A1(n10411), .A2(n10412), .ZN(n10405) );
  NAND3_X1 U10343 ( .A1(a_1_), .A2(n10413), .A3(b_21_), .ZN(n10412) );
  OR2_X1 U10344 ( .A1(n10193), .A2(n10192), .ZN(n10413) );
  NAND2_X1 U10345 ( .A1(n10192), .A2(n10193), .ZN(n10411) );
  NAND2_X1 U10346 ( .A1(n10414), .A2(n10415), .ZN(n10193) );
  NAND3_X1 U10347 ( .A1(a_2_), .A2(n10416), .A3(b_21_), .ZN(n10415) );
  OR2_X1 U10348 ( .A1(n10399), .A2(n10397), .ZN(n10416) );
  NAND2_X1 U10349 ( .A1(n10397), .A2(n10399), .ZN(n10414) );
  NAND2_X1 U10350 ( .A1(n10417), .A2(n10418), .ZN(n10399) );
  NAND3_X1 U10351 ( .A1(a_3_), .A2(n10419), .A3(b_21_), .ZN(n10418) );
  OR2_X1 U10352 ( .A1(n10395), .A2(n10393), .ZN(n10419) );
  NAND2_X1 U10353 ( .A1(n10393), .A2(n10395), .ZN(n10417) );
  NAND2_X1 U10354 ( .A1(n10420), .A2(n10421), .ZN(n10395) );
  NAND3_X1 U10355 ( .A1(a_4_), .A2(n10422), .A3(b_21_), .ZN(n10421) );
  OR2_X1 U10356 ( .A1(n10391), .A2(n10389), .ZN(n10422) );
  NAND2_X1 U10357 ( .A1(n10389), .A2(n10391), .ZN(n10420) );
  NAND2_X1 U10358 ( .A1(n10423), .A2(n10424), .ZN(n10391) );
  NAND3_X1 U10359 ( .A1(a_5_), .A2(n10425), .A3(b_21_), .ZN(n10424) );
  NAND2_X1 U10360 ( .A1(n10387), .A2(n10386), .ZN(n10425) );
  OR2_X1 U10361 ( .A1(n10386), .A2(n10387), .ZN(n10423) );
  AND2_X1 U10362 ( .A1(n10426), .A2(n10427), .ZN(n10387) );
  NAND3_X1 U10363 ( .A1(a_6_), .A2(n10428), .A3(b_21_), .ZN(n10427) );
  NAND2_X1 U10364 ( .A1(n10383), .A2(n10382), .ZN(n10428) );
  OR2_X1 U10365 ( .A1(n10382), .A2(n10383), .ZN(n10426) );
  AND2_X1 U10366 ( .A1(n10429), .A2(n10430), .ZN(n10383) );
  NAND3_X1 U10367 ( .A1(a_7_), .A2(n10431), .A3(b_21_), .ZN(n10430) );
  OR2_X1 U10368 ( .A1(n10379), .A2(n10377), .ZN(n10431) );
  NAND2_X1 U10369 ( .A1(n10377), .A2(n10379), .ZN(n10429) );
  NAND2_X1 U10370 ( .A1(n10432), .A2(n10433), .ZN(n10379) );
  NAND3_X1 U10371 ( .A1(a_8_), .A2(n10434), .A3(b_21_), .ZN(n10433) );
  OR2_X1 U10372 ( .A1(n10375), .A2(n10373), .ZN(n10434) );
  NAND2_X1 U10373 ( .A1(n10373), .A2(n10375), .ZN(n10432) );
  NAND2_X1 U10374 ( .A1(n10435), .A2(n10436), .ZN(n10375) );
  NAND3_X1 U10375 ( .A1(a_9_), .A2(n10437), .A3(b_21_), .ZN(n10436) );
  OR2_X1 U10376 ( .A1(n10371), .A2(n10370), .ZN(n10437) );
  NAND2_X1 U10377 ( .A1(n10370), .A2(n10371), .ZN(n10435) );
  NAND2_X1 U10378 ( .A1(n10438), .A2(n10439), .ZN(n10371) );
  NAND2_X1 U10379 ( .A1(n10368), .A2(n10440), .ZN(n10439) );
  OR2_X1 U10380 ( .A1(n10367), .A2(n10366), .ZN(n10440) );
  NOR2_X1 U10381 ( .A1(n7580), .A2(n8378), .ZN(n10368) );
  NAND2_X1 U10382 ( .A1(n10366), .A2(n10367), .ZN(n10438) );
  NAND2_X1 U10383 ( .A1(n10441), .A2(n10442), .ZN(n10367) );
  NAND2_X1 U10384 ( .A1(n10364), .A2(n10443), .ZN(n10442) );
  OR2_X1 U10385 ( .A1(n10363), .A2(n10361), .ZN(n10443) );
  NOR2_X1 U10386 ( .A1(n7580), .A2(n7724), .ZN(n10364) );
  NAND2_X1 U10387 ( .A1(n10361), .A2(n10363), .ZN(n10441) );
  NAND2_X1 U10388 ( .A1(n10444), .A2(n10445), .ZN(n10363) );
  NAND3_X1 U10389 ( .A1(a_12_), .A2(n10446), .A3(b_21_), .ZN(n10445) );
  OR2_X1 U10390 ( .A1(n10359), .A2(n10357), .ZN(n10446) );
  NAND2_X1 U10391 ( .A1(n10357), .A2(n10359), .ZN(n10444) );
  NAND2_X1 U10392 ( .A1(n10447), .A2(n10448), .ZN(n10359) );
  NAND2_X1 U10393 ( .A1(n10356), .A2(n10449), .ZN(n10448) );
  OR2_X1 U10394 ( .A1(n10355), .A2(n10354), .ZN(n10449) );
  NOR2_X1 U10395 ( .A1(n7580), .A2(n7702), .ZN(n10356) );
  NAND2_X1 U10396 ( .A1(n10354), .A2(n10355), .ZN(n10447) );
  NAND2_X1 U10397 ( .A1(n10450), .A2(n10451), .ZN(n10355) );
  NAND3_X1 U10398 ( .A1(a_14_), .A2(n10452), .A3(b_21_), .ZN(n10451) );
  NAND2_X1 U10399 ( .A1(n10351), .A2(n10350), .ZN(n10452) );
  OR2_X1 U10400 ( .A1(n10350), .A2(n10351), .ZN(n10450) );
  AND2_X1 U10401 ( .A1(n10453), .A2(n10454), .ZN(n10351) );
  NAND2_X1 U10402 ( .A1(n10348), .A2(n10455), .ZN(n10454) );
  OR2_X1 U10403 ( .A1(n10347), .A2(n10346), .ZN(n10455) );
  NOR2_X1 U10404 ( .A1(n7580), .A2(n7667), .ZN(n10348) );
  NAND2_X1 U10405 ( .A1(n10346), .A2(n10347), .ZN(n10453) );
  NAND2_X1 U10406 ( .A1(n10456), .A2(n10457), .ZN(n10347) );
  NAND3_X1 U10407 ( .A1(a_16_), .A2(n10458), .A3(b_21_), .ZN(n10457) );
  NAND2_X1 U10408 ( .A1(n10343), .A2(n10342), .ZN(n10458) );
  OR2_X1 U10409 ( .A1(n10342), .A2(n10343), .ZN(n10456) );
  AND2_X1 U10410 ( .A1(n10459), .A2(n10460), .ZN(n10343) );
  NAND2_X1 U10411 ( .A1(n10340), .A2(n10461), .ZN(n10460) );
  OR2_X1 U10412 ( .A1(n10339), .A2(n10337), .ZN(n10461) );
  NOR2_X1 U10413 ( .A1(n7580), .A2(n7645), .ZN(n10340) );
  NAND2_X1 U10414 ( .A1(n10337), .A2(n10339), .ZN(n10459) );
  NAND2_X1 U10415 ( .A1(n10462), .A2(n10463), .ZN(n10339) );
  NAND3_X1 U10416 ( .A1(a_18_), .A2(n10464), .A3(b_21_), .ZN(n10463) );
  NAND2_X1 U10417 ( .A1(n10335), .A2(n10334), .ZN(n10464) );
  OR2_X1 U10418 ( .A1(n10334), .A2(n10335), .ZN(n10462) );
  AND2_X1 U10419 ( .A1(n10465), .A2(n10466), .ZN(n10335) );
  NAND2_X1 U10420 ( .A1(n10332), .A2(n10467), .ZN(n10466) );
  OR2_X1 U10421 ( .A1(n10331), .A2(n10329), .ZN(n10467) );
  NOR2_X1 U10422 ( .A1(n7580), .A2(n7958), .ZN(n10332) );
  NAND2_X1 U10423 ( .A1(n10329), .A2(n10331), .ZN(n10465) );
  NAND2_X1 U10424 ( .A1(n10468), .A2(n10469), .ZN(n10331) );
  NAND3_X1 U10425 ( .A1(a_20_), .A2(n10470), .A3(b_21_), .ZN(n10469) );
  NAND2_X1 U10426 ( .A1(n10327), .A2(n10326), .ZN(n10470) );
  OR2_X1 U10427 ( .A1(n10326), .A2(n10327), .ZN(n10468) );
  AND2_X1 U10428 ( .A1(n10471), .A2(n10472), .ZN(n10327) );
  NAND2_X1 U10429 ( .A1(n7575), .A2(n10473), .ZN(n10472) );
  OR2_X1 U10430 ( .A1(n10324), .A2(n10323), .ZN(n10473) );
  INV_X1 U10431 ( .A(n7927), .ZN(n7575) );
  NAND2_X1 U10432 ( .A1(b_21_), .A2(a_21_), .ZN(n7927) );
  NAND2_X1 U10433 ( .A1(n10323), .A2(n10324), .ZN(n10471) );
  NAND2_X1 U10434 ( .A1(n10474), .A2(n10475), .ZN(n10324) );
  NAND3_X1 U10435 ( .A1(a_22_), .A2(n10476), .A3(b_21_), .ZN(n10475) );
  OR2_X1 U10436 ( .A1(n10320), .A2(n10318), .ZN(n10476) );
  NAND2_X1 U10437 ( .A1(n10318), .A2(n10320), .ZN(n10474) );
  NAND2_X1 U10438 ( .A1(n10477), .A2(n10478), .ZN(n10320) );
  NAND2_X1 U10439 ( .A1(n10264), .A2(n10479), .ZN(n10478) );
  OR2_X1 U10440 ( .A1(n10263), .A2(n10261), .ZN(n10479) );
  NOR2_X1 U10441 ( .A1(n7580), .A2(n7955), .ZN(n10264) );
  NAND2_X1 U10442 ( .A1(n10261), .A2(n10263), .ZN(n10477) );
  NAND2_X1 U10443 ( .A1(n10480), .A2(n10481), .ZN(n10263) );
  NAND3_X1 U10444 ( .A1(a_24_), .A2(n10482), .A3(b_21_), .ZN(n10481) );
  NAND2_X1 U10445 ( .A1(n10316), .A2(n10315), .ZN(n10482) );
  OR2_X1 U10446 ( .A1(n10315), .A2(n10316), .ZN(n10480) );
  AND2_X1 U10447 ( .A1(n10483), .A2(n10484), .ZN(n10316) );
  NAND2_X1 U10448 ( .A1(n10313), .A2(n10485), .ZN(n10484) );
  OR2_X1 U10449 ( .A1(n10312), .A2(n10311), .ZN(n10485) );
  NOR2_X1 U10450 ( .A1(n7580), .A2(n7952), .ZN(n10313) );
  NAND2_X1 U10451 ( .A1(n10311), .A2(n10312), .ZN(n10483) );
  NAND2_X1 U10452 ( .A1(n10308), .A2(n10486), .ZN(n10312) );
  NAND2_X1 U10453 ( .A1(n10307), .A2(n10309), .ZN(n10486) );
  NAND2_X1 U10454 ( .A1(n10487), .A2(n10488), .ZN(n10309) );
  NAND2_X1 U10455 ( .A1(b_21_), .A2(a_26_), .ZN(n10488) );
  INV_X1 U10456 ( .A(n10489), .ZN(n10487) );
  XNOR2_X1 U10457 ( .A(n10490), .B(n10491), .ZN(n10307) );
  NAND2_X1 U10458 ( .A1(n10492), .A2(n10493), .ZN(n10490) );
  NAND2_X1 U10459 ( .A1(a_26_), .A2(n10489), .ZN(n10308) );
  NAND2_X1 U10460 ( .A1(n10280), .A2(n10494), .ZN(n10489) );
  NAND2_X1 U10461 ( .A1(n10279), .A2(n10281), .ZN(n10494) );
  NAND2_X1 U10462 ( .A1(n10495), .A2(n10496), .ZN(n10281) );
  NAND2_X1 U10463 ( .A1(b_21_), .A2(a_27_), .ZN(n10496) );
  INV_X1 U10464 ( .A(n10497), .ZN(n10495) );
  XNOR2_X1 U10465 ( .A(n10498), .B(n10499), .ZN(n10279) );
  XOR2_X1 U10466 ( .A(n10500), .B(n10501), .Z(n10498) );
  NAND2_X1 U10467 ( .A1(b_20_), .A2(a_28_), .ZN(n10500) );
  NAND2_X1 U10468 ( .A1(a_27_), .A2(n10497), .ZN(n10280) );
  NAND2_X1 U10469 ( .A1(n10502), .A2(n10503), .ZN(n10497) );
  NAND3_X1 U10470 ( .A1(a_28_), .A2(n10504), .A3(b_21_), .ZN(n10503) );
  NAND2_X1 U10471 ( .A1(n10289), .A2(n10287), .ZN(n10504) );
  OR2_X1 U10472 ( .A1(n10287), .A2(n10289), .ZN(n10502) );
  AND2_X1 U10473 ( .A1(n10505), .A2(n10506), .ZN(n10289) );
  NAND2_X1 U10474 ( .A1(n10303), .A2(n10507), .ZN(n10506) );
  OR2_X1 U10475 ( .A1(n10304), .A2(n10305), .ZN(n10507) );
  NOR2_X1 U10476 ( .A1(n7580), .A2(n7460), .ZN(n10303) );
  INV_X1 U10477 ( .A(b_21_), .ZN(n7580) );
  NAND2_X1 U10478 ( .A1(n10305), .A2(n10304), .ZN(n10505) );
  NAND2_X1 U10479 ( .A1(n10508), .A2(n10509), .ZN(n10304) );
  NAND2_X1 U10480 ( .A1(b_19_), .A2(n10510), .ZN(n10509) );
  NAND2_X1 U10481 ( .A1(n7441), .A2(n10511), .ZN(n10510) );
  NAND2_X1 U10482 ( .A1(a_31_), .A2(n7956), .ZN(n10511) );
  NAND2_X1 U10483 ( .A1(b_20_), .A2(n10512), .ZN(n10508) );
  NAND2_X1 U10484 ( .A1(n7445), .A2(n10513), .ZN(n10512) );
  NAND2_X1 U10485 ( .A1(a_30_), .A2(n7606), .ZN(n10513) );
  AND3_X1 U10486 ( .A1(b_20_), .A2(n7409), .A3(b_21_), .ZN(n10305) );
  XNOR2_X1 U10487 ( .A(n10514), .B(n10515), .ZN(n10287) );
  XOR2_X1 U10488 ( .A(n10516), .B(n10517), .Z(n10514) );
  XNOR2_X1 U10489 ( .A(n10518), .B(n10519), .ZN(n10311) );
  NAND2_X1 U10490 ( .A1(n10520), .A2(n10521), .ZN(n10518) );
  XNOR2_X1 U10491 ( .A(n10522), .B(n10523), .ZN(n10315) );
  XOR2_X1 U10492 ( .A(n10524), .B(n10525), .Z(n10522) );
  XNOR2_X1 U10493 ( .A(n10526), .B(n10527), .ZN(n10261) );
  XNOR2_X1 U10494 ( .A(n10528), .B(n10529), .ZN(n10526) );
  NOR2_X1 U10495 ( .A1(n7954), .A2(n7956), .ZN(n10529) );
  XNOR2_X1 U10496 ( .A(n10530), .B(n10531), .ZN(n10318) );
  XNOR2_X1 U10497 ( .A(n10532), .B(n10533), .ZN(n10531) );
  XNOR2_X1 U10498 ( .A(n10534), .B(n10535), .ZN(n10323) );
  XOR2_X1 U10499 ( .A(n10536), .B(n10537), .Z(n10535) );
  NAND2_X1 U10500 ( .A1(b_20_), .A2(a_22_), .ZN(n10537) );
  XNOR2_X1 U10501 ( .A(n10538), .B(n10539), .ZN(n10326) );
  XOR2_X1 U10502 ( .A(n10540), .B(n10541), .Z(n10538) );
  XOR2_X1 U10503 ( .A(n10542), .B(n10543), .Z(n10329) );
  XOR2_X1 U10504 ( .A(n10544), .B(n10545), .Z(n10542) );
  XNOR2_X1 U10505 ( .A(n10546), .B(n10547), .ZN(n10334) );
  XOR2_X1 U10506 ( .A(n10548), .B(n10549), .Z(n10546) );
  XNOR2_X1 U10507 ( .A(n10550), .B(n10551), .ZN(n10337) );
  XNOR2_X1 U10508 ( .A(n10552), .B(n10553), .ZN(n10550) );
  NOR2_X1 U10509 ( .A1(n7960), .A2(n7956), .ZN(n10553) );
  XOR2_X1 U10510 ( .A(n10554), .B(n10555), .Z(n10342) );
  XNOR2_X1 U10511 ( .A(n10556), .B(n10557), .ZN(n10555) );
  XNOR2_X1 U10512 ( .A(n10558), .B(n10559), .ZN(n10346) );
  XNOR2_X1 U10513 ( .A(n10560), .B(n10561), .ZN(n10558) );
  NOR2_X1 U10514 ( .A1(n8353), .A2(n7956), .ZN(n10561) );
  XOR2_X1 U10515 ( .A(n10562), .B(n10563), .Z(n10350) );
  XNOR2_X1 U10516 ( .A(n10564), .B(n10565), .ZN(n10563) );
  XNOR2_X1 U10517 ( .A(n10566), .B(n10567), .ZN(n10354) );
  XNOR2_X1 U10518 ( .A(n10568), .B(n10569), .ZN(n10566) );
  NOR2_X1 U10519 ( .A1(n7962), .A2(n7956), .ZN(n10569) );
  XNOR2_X1 U10520 ( .A(n10570), .B(n10571), .ZN(n10357) );
  XNOR2_X1 U10521 ( .A(n10572), .B(n10573), .ZN(n10571) );
  XNOR2_X1 U10522 ( .A(n10574), .B(n10575), .ZN(n10361) );
  XOR2_X1 U10523 ( .A(n10576), .B(n10577), .Z(n10575) );
  NAND2_X1 U10524 ( .A1(b_20_), .A2(a_12_), .ZN(n10577) );
  XNOR2_X1 U10525 ( .A(n10578), .B(n10579), .ZN(n10366) );
  XOR2_X1 U10526 ( .A(n10580), .B(n10581), .Z(n10579) );
  NAND2_X1 U10527 ( .A1(b_20_), .A2(a_11_), .ZN(n10581) );
  XNOR2_X1 U10528 ( .A(n10582), .B(n10583), .ZN(n10370) );
  XNOR2_X1 U10529 ( .A(n10584), .B(n10585), .ZN(n10582) );
  XOR2_X1 U10530 ( .A(n10586), .B(n10587), .Z(n10373) );
  XOR2_X1 U10531 ( .A(n10588), .B(n10589), .Z(n10586) );
  XNOR2_X1 U10532 ( .A(n10590), .B(n10591), .ZN(n10377) );
  XNOR2_X1 U10533 ( .A(n10592), .B(n10593), .ZN(n10590) );
  NOR2_X1 U10534 ( .A1(n8602), .A2(n7956), .ZN(n10593) );
  XOR2_X1 U10535 ( .A(n10594), .B(n10595), .Z(n10382) );
  NAND2_X1 U10536 ( .A1(n10596), .A2(n10597), .ZN(n10594) );
  XNOR2_X1 U10537 ( .A(n10598), .B(n10599), .ZN(n10386) );
  NOR2_X1 U10538 ( .A1(n10600), .A2(n10601), .ZN(n10599) );
  NOR2_X1 U10539 ( .A1(n10602), .A2(n10603), .ZN(n10600) );
  NOR2_X1 U10540 ( .A1(n7807), .A2(n7956), .ZN(n10602) );
  XOR2_X1 U10541 ( .A(n10604), .B(n10605), .Z(n10389) );
  XOR2_X1 U10542 ( .A(n10606), .B(n10607), .Z(n10604) );
  XOR2_X1 U10543 ( .A(n10608), .B(n10609), .Z(n10393) );
  XOR2_X1 U10544 ( .A(n10610), .B(n10611), .Z(n10608) );
  NOR2_X1 U10545 ( .A1(n7836), .A2(n7956), .ZN(n10611) );
  XNOR2_X1 U10546 ( .A(n10612), .B(n10613), .ZN(n10397) );
  NAND2_X1 U10547 ( .A1(n10614), .A2(n10615), .ZN(n10612) );
  XNOR2_X1 U10548 ( .A(n10616), .B(n10617), .ZN(n10192) );
  NAND2_X1 U10549 ( .A1(n10618), .A2(n10619), .ZN(n10616) );
  XNOR2_X1 U10550 ( .A(n10620), .B(n10621), .ZN(n10403) );
  XNOR2_X1 U10551 ( .A(n10622), .B(n10623), .ZN(n10620) );
  XNOR2_X1 U10552 ( .A(n10624), .B(n10625), .ZN(n10402) );
  XOR2_X1 U10553 ( .A(n10626), .B(n10627), .Z(n10624) );
  NOR2_X1 U10554 ( .A1(n8197), .A2(n7956), .ZN(n10627) );
  XOR2_X1 U10555 ( .A(n8146), .B(n8145), .Z(n10407) );
  NAND3_X1 U10556 ( .A1(n8145), .A2(n8146), .A3(n10628), .ZN(n8041) );
  XOR2_X1 U10557 ( .A(n8139), .B(n8138), .Z(n10628) );
  NAND2_X1 U10558 ( .A1(n10629), .A2(n10630), .ZN(n8146) );
  NAND3_X1 U10559 ( .A1(a_0_), .A2(n10631), .A3(b_20_), .ZN(n10630) );
  OR2_X1 U10560 ( .A1(n10626), .A2(n10625), .ZN(n10631) );
  NAND2_X1 U10561 ( .A1(n10625), .A2(n10626), .ZN(n10629) );
  NAND2_X1 U10562 ( .A1(n10632), .A2(n10633), .ZN(n10626) );
  NAND2_X1 U10563 ( .A1(n10623), .A2(n10634), .ZN(n10633) );
  NAND2_X1 U10564 ( .A1(n10622), .A2(n10621), .ZN(n10634) );
  NOR2_X1 U10565 ( .A1(n7956), .A2(n7872), .ZN(n10623) );
  OR2_X1 U10566 ( .A1(n10621), .A2(n10622), .ZN(n10632) );
  AND2_X1 U10567 ( .A1(n10618), .A2(n10635), .ZN(n10622) );
  NAND2_X1 U10568 ( .A1(n10617), .A2(n10619), .ZN(n10635) );
  NAND2_X1 U10569 ( .A1(n10636), .A2(n10637), .ZN(n10619) );
  NAND2_X1 U10570 ( .A1(b_20_), .A2(a_2_), .ZN(n10637) );
  INV_X1 U10571 ( .A(n10638), .ZN(n10636) );
  XNOR2_X1 U10572 ( .A(n10639), .B(n10640), .ZN(n10617) );
  XOR2_X1 U10573 ( .A(n10641), .B(n10642), .Z(n10640) );
  NAND2_X1 U10574 ( .A1(b_19_), .A2(a_3_), .ZN(n10642) );
  NAND2_X1 U10575 ( .A1(a_2_), .A2(n10638), .ZN(n10618) );
  NAND2_X1 U10576 ( .A1(n10614), .A2(n10643), .ZN(n10638) );
  NAND2_X1 U10577 ( .A1(n10613), .A2(n10615), .ZN(n10643) );
  NAND2_X1 U10578 ( .A1(n10644), .A2(n10645), .ZN(n10615) );
  NAND2_X1 U10579 ( .A1(b_20_), .A2(a_3_), .ZN(n10645) );
  INV_X1 U10580 ( .A(n10646), .ZN(n10644) );
  XOR2_X1 U10581 ( .A(n10647), .B(n10648), .Z(n10613) );
  XOR2_X1 U10582 ( .A(n10649), .B(n10650), .Z(n10647) );
  NOR2_X1 U10583 ( .A1(n7836), .A2(n7606), .ZN(n10650) );
  NAND2_X1 U10584 ( .A1(a_3_), .A2(n10646), .ZN(n10614) );
  NAND2_X1 U10585 ( .A1(n10651), .A2(n10652), .ZN(n10646) );
  NAND3_X1 U10586 ( .A1(a_4_), .A2(n10653), .A3(b_20_), .ZN(n10652) );
  OR2_X1 U10587 ( .A1(n10610), .A2(n10609), .ZN(n10653) );
  NAND2_X1 U10588 ( .A1(n10609), .A2(n10610), .ZN(n10651) );
  NAND2_X1 U10589 ( .A1(n10654), .A2(n10655), .ZN(n10610) );
  NAND2_X1 U10590 ( .A1(n10607), .A2(n10656), .ZN(n10655) );
  OR2_X1 U10591 ( .A1(n10606), .A2(n10605), .ZN(n10656) );
  NOR2_X1 U10592 ( .A1(n7956), .A2(n7823), .ZN(n10607) );
  NAND2_X1 U10593 ( .A1(n10605), .A2(n10606), .ZN(n10654) );
  OR2_X1 U10594 ( .A1(n10601), .A2(n10657), .ZN(n10606) );
  AND2_X1 U10595 ( .A1(n10598), .A2(n10658), .ZN(n10657) );
  NAND2_X1 U10596 ( .A1(n10659), .A2(n10660), .ZN(n10658) );
  NAND2_X1 U10597 ( .A1(b_20_), .A2(a_6_), .ZN(n10660) );
  XNOR2_X1 U10598 ( .A(n10661), .B(n10662), .ZN(n10598) );
  XOR2_X1 U10599 ( .A(n10663), .B(n10664), .Z(n10662) );
  NAND2_X1 U10600 ( .A1(b_19_), .A2(a_7_), .ZN(n10664) );
  NOR2_X1 U10601 ( .A1(n7807), .A2(n10659), .ZN(n10601) );
  INV_X1 U10602 ( .A(n10603), .ZN(n10659) );
  NAND2_X1 U10603 ( .A1(n10596), .A2(n10665), .ZN(n10603) );
  NAND2_X1 U10604 ( .A1(n10595), .A2(n10597), .ZN(n10665) );
  NAND2_X1 U10605 ( .A1(n10666), .A2(n10667), .ZN(n10597) );
  NAND2_X1 U10606 ( .A1(b_20_), .A2(a_7_), .ZN(n10667) );
  INV_X1 U10607 ( .A(n10668), .ZN(n10666) );
  XOR2_X1 U10608 ( .A(n10669), .B(n10670), .Z(n10595) );
  XOR2_X1 U10609 ( .A(n10671), .B(n10672), .Z(n10669) );
  NOR2_X1 U10610 ( .A1(n8602), .A2(n7606), .ZN(n10672) );
  NAND2_X1 U10611 ( .A1(a_7_), .A2(n10668), .ZN(n10596) );
  NAND2_X1 U10612 ( .A1(n10673), .A2(n10674), .ZN(n10668) );
  NAND3_X1 U10613 ( .A1(a_8_), .A2(n10675), .A3(b_20_), .ZN(n10674) );
  NAND2_X1 U10614 ( .A1(n10592), .A2(n10591), .ZN(n10675) );
  OR2_X1 U10615 ( .A1(n10591), .A2(n10592), .ZN(n10673) );
  AND2_X1 U10616 ( .A1(n10676), .A2(n10677), .ZN(n10592) );
  NAND2_X1 U10617 ( .A1(n10588), .A2(n10678), .ZN(n10677) );
  OR2_X1 U10618 ( .A1(n10589), .A2(n10587), .ZN(n10678) );
  NOR2_X1 U10619 ( .A1(n7956), .A2(n7753), .ZN(n10588) );
  NAND2_X1 U10620 ( .A1(n10587), .A2(n10589), .ZN(n10676) );
  NAND2_X1 U10621 ( .A1(n10679), .A2(n10680), .ZN(n10589) );
  NAND2_X1 U10622 ( .A1(n10585), .A2(n10681), .ZN(n10680) );
  NAND2_X1 U10623 ( .A1(n10584), .A2(n10583), .ZN(n10681) );
  NOR2_X1 U10624 ( .A1(n7956), .A2(n8378), .ZN(n10585) );
  OR2_X1 U10625 ( .A1(n10583), .A2(n10584), .ZN(n10679) );
  AND2_X1 U10626 ( .A1(n10682), .A2(n10683), .ZN(n10584) );
  NAND3_X1 U10627 ( .A1(a_11_), .A2(n10684), .A3(b_20_), .ZN(n10683) );
  OR2_X1 U10628 ( .A1(n10580), .A2(n10578), .ZN(n10684) );
  NAND2_X1 U10629 ( .A1(n10578), .A2(n10580), .ZN(n10682) );
  NAND2_X1 U10630 ( .A1(n10685), .A2(n10686), .ZN(n10580) );
  NAND3_X1 U10631 ( .A1(a_12_), .A2(n10687), .A3(b_20_), .ZN(n10686) );
  OR2_X1 U10632 ( .A1(n10576), .A2(n10574), .ZN(n10687) );
  NAND2_X1 U10633 ( .A1(n10574), .A2(n10576), .ZN(n10685) );
  NAND2_X1 U10634 ( .A1(n10688), .A2(n10689), .ZN(n10576) );
  NAND2_X1 U10635 ( .A1(n10573), .A2(n10690), .ZN(n10689) );
  OR2_X1 U10636 ( .A1(n10572), .A2(n10570), .ZN(n10690) );
  NOR2_X1 U10637 ( .A1(n7956), .A2(n7702), .ZN(n10573) );
  NAND2_X1 U10638 ( .A1(n10570), .A2(n10572), .ZN(n10688) );
  NAND2_X1 U10639 ( .A1(n10691), .A2(n10692), .ZN(n10572) );
  NAND3_X1 U10640 ( .A1(a_14_), .A2(n10693), .A3(b_20_), .ZN(n10692) );
  NAND2_X1 U10641 ( .A1(n10568), .A2(n10567), .ZN(n10693) );
  OR2_X1 U10642 ( .A1(n10567), .A2(n10568), .ZN(n10691) );
  AND2_X1 U10643 ( .A1(n10694), .A2(n10695), .ZN(n10568) );
  NAND2_X1 U10644 ( .A1(n10565), .A2(n10696), .ZN(n10695) );
  OR2_X1 U10645 ( .A1(n10564), .A2(n10562), .ZN(n10696) );
  NOR2_X1 U10646 ( .A1(n7956), .A2(n7667), .ZN(n10565) );
  NAND2_X1 U10647 ( .A1(n10562), .A2(n10564), .ZN(n10694) );
  NAND2_X1 U10648 ( .A1(n10697), .A2(n10698), .ZN(n10564) );
  NAND3_X1 U10649 ( .A1(a_16_), .A2(n10699), .A3(b_20_), .ZN(n10698) );
  NAND2_X1 U10650 ( .A1(n10560), .A2(n10559), .ZN(n10699) );
  OR2_X1 U10651 ( .A1(n10559), .A2(n10560), .ZN(n10697) );
  AND2_X1 U10652 ( .A1(n10700), .A2(n10701), .ZN(n10560) );
  NAND2_X1 U10653 ( .A1(n10557), .A2(n10702), .ZN(n10701) );
  OR2_X1 U10654 ( .A1(n10556), .A2(n10554), .ZN(n10702) );
  NOR2_X1 U10655 ( .A1(n7956), .A2(n7645), .ZN(n10557) );
  NAND2_X1 U10656 ( .A1(n10554), .A2(n10556), .ZN(n10700) );
  NAND2_X1 U10657 ( .A1(n10703), .A2(n10704), .ZN(n10556) );
  NAND3_X1 U10658 ( .A1(a_18_), .A2(n10705), .A3(b_20_), .ZN(n10704) );
  NAND2_X1 U10659 ( .A1(n10552), .A2(n10551), .ZN(n10705) );
  OR2_X1 U10660 ( .A1(n10551), .A2(n10552), .ZN(n10703) );
  AND2_X1 U10661 ( .A1(n10706), .A2(n10707), .ZN(n10552) );
  NAND2_X1 U10662 ( .A1(n10549), .A2(n10708), .ZN(n10707) );
  OR2_X1 U10663 ( .A1(n10548), .A2(n10547), .ZN(n10708) );
  NOR2_X1 U10664 ( .A1(n7956), .A2(n7958), .ZN(n10549) );
  NAND2_X1 U10665 ( .A1(n10547), .A2(n10548), .ZN(n10706) );
  NAND2_X1 U10666 ( .A1(n10709), .A2(n10710), .ZN(n10548) );
  NAND2_X1 U10667 ( .A1(n10543), .A2(n10711), .ZN(n10710) );
  OR2_X1 U10668 ( .A1(n10544), .A2(n10545), .ZN(n10711) );
  XNOR2_X1 U10669 ( .A(n10712), .B(n10713), .ZN(n10543) );
  XNOR2_X1 U10670 ( .A(n10714), .B(n10715), .ZN(n10712) );
  NAND2_X1 U10671 ( .A1(n10545), .A2(n10544), .ZN(n10709) );
  NAND2_X1 U10672 ( .A1(n10716), .A2(n10717), .ZN(n10544) );
  NAND2_X1 U10673 ( .A1(n10541), .A2(n10718), .ZN(n10717) );
  OR2_X1 U10674 ( .A1(n10540), .A2(n10539), .ZN(n10718) );
  NOR2_X1 U10675 ( .A1(n7956), .A2(n7578), .ZN(n10541) );
  NAND2_X1 U10676 ( .A1(n10539), .A2(n10540), .ZN(n10716) );
  NAND2_X1 U10677 ( .A1(n10719), .A2(n10720), .ZN(n10540) );
  NAND3_X1 U10678 ( .A1(a_22_), .A2(n10721), .A3(b_20_), .ZN(n10720) );
  OR2_X1 U10679 ( .A1(n10536), .A2(n10534), .ZN(n10721) );
  NAND2_X1 U10680 ( .A1(n10534), .A2(n10536), .ZN(n10719) );
  NAND2_X1 U10681 ( .A1(n10722), .A2(n10723), .ZN(n10536) );
  NAND2_X1 U10682 ( .A1(n10533), .A2(n10724), .ZN(n10723) );
  OR2_X1 U10683 ( .A1(n10532), .A2(n10530), .ZN(n10724) );
  NOR2_X1 U10684 ( .A1(n7956), .A2(n7955), .ZN(n10533) );
  NAND2_X1 U10685 ( .A1(n10530), .A2(n10532), .ZN(n10722) );
  NAND2_X1 U10686 ( .A1(n10725), .A2(n10726), .ZN(n10532) );
  NAND3_X1 U10687 ( .A1(a_24_), .A2(n10727), .A3(b_20_), .ZN(n10726) );
  NAND2_X1 U10688 ( .A1(n10528), .A2(n10527), .ZN(n10727) );
  OR2_X1 U10689 ( .A1(n10527), .A2(n10528), .ZN(n10725) );
  AND2_X1 U10690 ( .A1(n10728), .A2(n10729), .ZN(n10528) );
  NAND2_X1 U10691 ( .A1(n10525), .A2(n10730), .ZN(n10729) );
  OR2_X1 U10692 ( .A1(n10524), .A2(n10523), .ZN(n10730) );
  NOR2_X1 U10693 ( .A1(n7956), .A2(n7952), .ZN(n10525) );
  NAND2_X1 U10694 ( .A1(n10523), .A2(n10524), .ZN(n10728) );
  NAND2_X1 U10695 ( .A1(n10520), .A2(n10731), .ZN(n10524) );
  NAND2_X1 U10696 ( .A1(n10519), .A2(n10521), .ZN(n10731) );
  NAND2_X1 U10697 ( .A1(n10732), .A2(n10733), .ZN(n10521) );
  NAND2_X1 U10698 ( .A1(b_20_), .A2(a_26_), .ZN(n10733) );
  INV_X1 U10699 ( .A(n10734), .ZN(n10732) );
  XNOR2_X1 U10700 ( .A(n10735), .B(n10736), .ZN(n10519) );
  NAND2_X1 U10701 ( .A1(n10737), .A2(n10738), .ZN(n10735) );
  NAND2_X1 U10702 ( .A1(a_26_), .A2(n10734), .ZN(n10520) );
  NAND2_X1 U10703 ( .A1(n10492), .A2(n10739), .ZN(n10734) );
  NAND2_X1 U10704 ( .A1(n10491), .A2(n10493), .ZN(n10739) );
  NAND2_X1 U10705 ( .A1(n10740), .A2(n10741), .ZN(n10493) );
  NAND2_X1 U10706 ( .A1(b_20_), .A2(a_27_), .ZN(n10741) );
  INV_X1 U10707 ( .A(n10742), .ZN(n10740) );
  XNOR2_X1 U10708 ( .A(n10743), .B(n10744), .ZN(n10491) );
  XOR2_X1 U10709 ( .A(n10745), .B(n10746), .Z(n10743) );
  NAND2_X1 U10710 ( .A1(b_19_), .A2(a_28_), .ZN(n10745) );
  NAND2_X1 U10711 ( .A1(a_27_), .A2(n10742), .ZN(n10492) );
  NAND2_X1 U10712 ( .A1(n10747), .A2(n10748), .ZN(n10742) );
  NAND3_X1 U10713 ( .A1(a_28_), .A2(n10749), .A3(b_20_), .ZN(n10748) );
  NAND2_X1 U10714 ( .A1(n10501), .A2(n10499), .ZN(n10749) );
  OR2_X1 U10715 ( .A1(n10499), .A2(n10501), .ZN(n10747) );
  AND2_X1 U10716 ( .A1(n10750), .A2(n10751), .ZN(n10501) );
  NAND2_X1 U10717 ( .A1(n10515), .A2(n10752), .ZN(n10751) );
  OR2_X1 U10718 ( .A1(n10516), .A2(n10517), .ZN(n10752) );
  NOR2_X1 U10719 ( .A1(n7956), .A2(n7460), .ZN(n10515) );
  INV_X1 U10720 ( .A(b_20_), .ZN(n7956) );
  NAND2_X1 U10721 ( .A1(n10517), .A2(n10516), .ZN(n10750) );
  NAND2_X1 U10722 ( .A1(n10753), .A2(n10754), .ZN(n10516) );
  NAND2_X1 U10723 ( .A1(b_18_), .A2(n10755), .ZN(n10754) );
  NAND2_X1 U10724 ( .A1(n7441), .A2(n10756), .ZN(n10755) );
  NAND2_X1 U10725 ( .A1(a_31_), .A2(n7606), .ZN(n10756) );
  NAND2_X1 U10726 ( .A1(b_19_), .A2(n10757), .ZN(n10753) );
  NAND2_X1 U10727 ( .A1(n7445), .A2(n10758), .ZN(n10757) );
  NAND2_X1 U10728 ( .A1(a_30_), .A2(n7959), .ZN(n10758) );
  AND3_X1 U10729 ( .A1(b_19_), .A2(n7409), .A3(b_20_), .ZN(n10517) );
  XNOR2_X1 U10730 ( .A(n10759), .B(n10760), .ZN(n10499) );
  XOR2_X1 U10731 ( .A(n10761), .B(n10762), .Z(n10759) );
  XNOR2_X1 U10732 ( .A(n10763), .B(n10764), .ZN(n10523) );
  NAND2_X1 U10733 ( .A1(n10765), .A2(n10766), .ZN(n10763) );
  XNOR2_X1 U10734 ( .A(n10767), .B(n10768), .ZN(n10527) );
  XOR2_X1 U10735 ( .A(n10769), .B(n10770), .Z(n10767) );
  XNOR2_X1 U10736 ( .A(n10771), .B(n10772), .ZN(n10530) );
  XNOR2_X1 U10737 ( .A(n10773), .B(n10774), .ZN(n10771) );
  NOR2_X1 U10738 ( .A1(n7954), .A2(n7606), .ZN(n10774) );
  XNOR2_X1 U10739 ( .A(n10775), .B(n10776), .ZN(n10534) );
  XNOR2_X1 U10740 ( .A(n10777), .B(n10778), .ZN(n10776) );
  XNOR2_X1 U10741 ( .A(n10779), .B(n10780), .ZN(n10539) );
  XOR2_X1 U10742 ( .A(n10781), .B(n10782), .Z(n10780) );
  NAND2_X1 U10743 ( .A1(b_19_), .A2(a_22_), .ZN(n10782) );
  INV_X1 U10744 ( .A(n7592), .ZN(n10545) );
  NAND2_X1 U10745 ( .A1(b_20_), .A2(a_20_), .ZN(n7592) );
  XNOR2_X1 U10746 ( .A(n10783), .B(n10784), .ZN(n10547) );
  XOR2_X1 U10747 ( .A(n10785), .B(n10786), .Z(n10783) );
  NAND2_X1 U10748 ( .A1(b_19_), .A2(a_20_), .ZN(n10785) );
  XNOR2_X1 U10749 ( .A(n10787), .B(n10788), .ZN(n10551) );
  XOR2_X1 U10750 ( .A(n10789), .B(n7604), .Z(n10787) );
  XNOR2_X1 U10751 ( .A(n10790), .B(n10791), .ZN(n10554) );
  XNOR2_X1 U10752 ( .A(n10792), .B(n10793), .ZN(n10790) );
  NOR2_X1 U10753 ( .A1(n7960), .A2(n7606), .ZN(n10793) );
  XNOR2_X1 U10754 ( .A(n10794), .B(n10795), .ZN(n10559) );
  XOR2_X1 U10755 ( .A(n10796), .B(n10797), .Z(n10794) );
  XNOR2_X1 U10756 ( .A(n10798), .B(n10799), .ZN(n10562) );
  XOR2_X1 U10757 ( .A(n10800), .B(n10801), .Z(n10799) );
  NAND2_X1 U10758 ( .A1(b_19_), .A2(a_16_), .ZN(n10801) );
  XOR2_X1 U10759 ( .A(n10802), .B(n10803), .Z(n10567) );
  XNOR2_X1 U10760 ( .A(n10804), .B(n10805), .ZN(n10803) );
  XNOR2_X1 U10761 ( .A(n10806), .B(n10807), .ZN(n10570) );
  XNOR2_X1 U10762 ( .A(n10808), .B(n10809), .ZN(n10806) );
  NOR2_X1 U10763 ( .A1(n7962), .A2(n7606), .ZN(n10809) );
  XOR2_X1 U10764 ( .A(n10810), .B(n10811), .Z(n10574) );
  XOR2_X1 U10765 ( .A(n10812), .B(n10813), .Z(n10810) );
  XOR2_X1 U10766 ( .A(n10814), .B(n10815), .Z(n10578) );
  XOR2_X1 U10767 ( .A(n10816), .B(n10817), .Z(n10814) );
  NOR2_X1 U10768 ( .A1(n8585), .A2(n7606), .ZN(n10817) );
  XOR2_X1 U10769 ( .A(n10818), .B(n10819), .Z(n10583) );
  NAND2_X1 U10770 ( .A1(n10820), .A2(n10821), .ZN(n10818) );
  XNOR2_X1 U10771 ( .A(n10822), .B(n10823), .ZN(n10587) );
  NAND2_X1 U10772 ( .A1(n10824), .A2(n10825), .ZN(n10822) );
  XNOR2_X1 U10773 ( .A(n10826), .B(n10827), .ZN(n10591) );
  XOR2_X1 U10774 ( .A(n10828), .B(n10829), .Z(n10826) );
  NOR2_X1 U10775 ( .A1(n7753), .A2(n7606), .ZN(n10829) );
  XNOR2_X1 U10776 ( .A(n10830), .B(n10831), .ZN(n10605) );
  XNOR2_X1 U10777 ( .A(n10832), .B(n10833), .ZN(n10830) );
  NOR2_X1 U10778 ( .A1(n7807), .A2(n7606), .ZN(n10833) );
  XNOR2_X1 U10779 ( .A(n10834), .B(n10835), .ZN(n10609) );
  XNOR2_X1 U10780 ( .A(n10836), .B(n10837), .ZN(n10834) );
  NOR2_X1 U10781 ( .A1(n7823), .A2(n7606), .ZN(n10837) );
  XOR2_X1 U10782 ( .A(n10838), .B(n10839), .Z(n10621) );
  XOR2_X1 U10783 ( .A(n10840), .B(n10841), .Z(n10839) );
  NAND2_X1 U10784 ( .A1(b_19_), .A2(a_2_), .ZN(n10841) );
  XNOR2_X1 U10785 ( .A(n10842), .B(n10843), .ZN(n10625) );
  XNOR2_X1 U10786 ( .A(n10844), .B(n10845), .ZN(n10842) );
  NOR2_X1 U10787 ( .A1(n7872), .A2(n7606), .ZN(n10845) );
  XNOR2_X1 U10788 ( .A(n10846), .B(n10847), .ZN(n8145) );
  XOR2_X1 U10789 ( .A(n10848), .B(n10849), .Z(n10847) );
  NAND2_X1 U10790 ( .A1(b_19_), .A2(a_0_), .ZN(n10849) );
  NAND3_X1 U10791 ( .A1(n10850), .A2(n8139), .A3(n8138), .ZN(n8046) );
  XOR2_X1 U10792 ( .A(n10851), .B(n10852), .Z(n8138) );
  XOR2_X1 U10793 ( .A(n10853), .B(n10854), .Z(n10851) );
  NOR2_X1 U10794 ( .A1(n8197), .A2(n7959), .ZN(n10854) );
  NAND2_X1 U10795 ( .A1(n10855), .A2(n10856), .ZN(n8139) );
  NAND3_X1 U10796 ( .A1(a_0_), .A2(n10857), .A3(b_19_), .ZN(n10856) );
  OR2_X1 U10797 ( .A1(n10848), .A2(n10846), .ZN(n10857) );
  NAND2_X1 U10798 ( .A1(n10846), .A2(n10848), .ZN(n10855) );
  NAND2_X1 U10799 ( .A1(n10858), .A2(n10859), .ZN(n10848) );
  NAND3_X1 U10800 ( .A1(a_1_), .A2(n10860), .A3(b_19_), .ZN(n10859) );
  NAND2_X1 U10801 ( .A1(n10844), .A2(n10843), .ZN(n10860) );
  OR2_X1 U10802 ( .A1(n10843), .A2(n10844), .ZN(n10858) );
  AND2_X1 U10803 ( .A1(n10861), .A2(n10862), .ZN(n10844) );
  NAND3_X1 U10804 ( .A1(a_2_), .A2(n10863), .A3(b_19_), .ZN(n10862) );
  OR2_X1 U10805 ( .A1(n10840), .A2(n10838), .ZN(n10863) );
  NAND2_X1 U10806 ( .A1(n10838), .A2(n10840), .ZN(n10861) );
  NAND2_X1 U10807 ( .A1(n10864), .A2(n10865), .ZN(n10840) );
  NAND3_X1 U10808 ( .A1(a_3_), .A2(n10866), .A3(b_19_), .ZN(n10865) );
  OR2_X1 U10809 ( .A1(n10641), .A2(n10639), .ZN(n10866) );
  NAND2_X1 U10810 ( .A1(n10639), .A2(n10641), .ZN(n10864) );
  NAND2_X1 U10811 ( .A1(n10867), .A2(n10868), .ZN(n10641) );
  NAND3_X1 U10812 ( .A1(a_4_), .A2(n10869), .A3(b_19_), .ZN(n10868) );
  OR2_X1 U10813 ( .A1(n10649), .A2(n10648), .ZN(n10869) );
  NAND2_X1 U10814 ( .A1(n10648), .A2(n10649), .ZN(n10867) );
  NAND2_X1 U10815 ( .A1(n10870), .A2(n10871), .ZN(n10649) );
  NAND3_X1 U10816 ( .A1(a_5_), .A2(n10872), .A3(b_19_), .ZN(n10871) );
  NAND2_X1 U10817 ( .A1(n10836), .A2(n10835), .ZN(n10872) );
  OR2_X1 U10818 ( .A1(n10835), .A2(n10836), .ZN(n10870) );
  AND2_X1 U10819 ( .A1(n10873), .A2(n10874), .ZN(n10836) );
  NAND3_X1 U10820 ( .A1(a_6_), .A2(n10875), .A3(b_19_), .ZN(n10874) );
  NAND2_X1 U10821 ( .A1(n10832), .A2(n10831), .ZN(n10875) );
  OR2_X1 U10822 ( .A1(n10831), .A2(n10832), .ZN(n10873) );
  AND2_X1 U10823 ( .A1(n10876), .A2(n10877), .ZN(n10832) );
  NAND3_X1 U10824 ( .A1(a_7_), .A2(n10878), .A3(b_19_), .ZN(n10877) );
  OR2_X1 U10825 ( .A1(n10663), .A2(n10661), .ZN(n10878) );
  NAND2_X1 U10826 ( .A1(n10661), .A2(n10663), .ZN(n10876) );
  NAND2_X1 U10827 ( .A1(n10879), .A2(n10880), .ZN(n10663) );
  NAND3_X1 U10828 ( .A1(a_8_), .A2(n10881), .A3(b_19_), .ZN(n10880) );
  OR2_X1 U10829 ( .A1(n10671), .A2(n10670), .ZN(n10881) );
  NAND2_X1 U10830 ( .A1(n10670), .A2(n10671), .ZN(n10879) );
  NAND2_X1 U10831 ( .A1(n10882), .A2(n10883), .ZN(n10671) );
  NAND3_X1 U10832 ( .A1(a_9_), .A2(n10884), .A3(b_19_), .ZN(n10883) );
  OR2_X1 U10833 ( .A1(n10828), .A2(n10827), .ZN(n10884) );
  NAND2_X1 U10834 ( .A1(n10827), .A2(n10828), .ZN(n10882) );
  NAND2_X1 U10835 ( .A1(n10824), .A2(n10885), .ZN(n10828) );
  NAND2_X1 U10836 ( .A1(n10823), .A2(n10825), .ZN(n10885) );
  NAND2_X1 U10837 ( .A1(n10886), .A2(n10887), .ZN(n10825) );
  NAND2_X1 U10838 ( .A1(b_19_), .A2(a_10_), .ZN(n10887) );
  INV_X1 U10839 ( .A(n10888), .ZN(n10886) );
  XNOR2_X1 U10840 ( .A(n10889), .B(n10890), .ZN(n10823) );
  XNOR2_X1 U10841 ( .A(n10891), .B(n10892), .ZN(n10889) );
  NAND2_X1 U10842 ( .A1(a_10_), .A2(n10888), .ZN(n10824) );
  NAND2_X1 U10843 ( .A1(n10820), .A2(n10893), .ZN(n10888) );
  NAND2_X1 U10844 ( .A1(n10819), .A2(n10821), .ZN(n10893) );
  NAND2_X1 U10845 ( .A1(n10894), .A2(n10895), .ZN(n10821) );
  NAND2_X1 U10846 ( .A1(b_19_), .A2(a_11_), .ZN(n10895) );
  INV_X1 U10847 ( .A(n10896), .ZN(n10894) );
  XNOR2_X1 U10848 ( .A(n10897), .B(n10898), .ZN(n10819) );
  XNOR2_X1 U10849 ( .A(n10899), .B(n10900), .ZN(n10898) );
  NAND2_X1 U10850 ( .A1(a_11_), .A2(n10896), .ZN(n10820) );
  NAND2_X1 U10851 ( .A1(n10901), .A2(n10902), .ZN(n10896) );
  NAND3_X1 U10852 ( .A1(a_12_), .A2(n10903), .A3(b_19_), .ZN(n10902) );
  OR2_X1 U10853 ( .A1(n10816), .A2(n10815), .ZN(n10903) );
  NAND2_X1 U10854 ( .A1(n10815), .A2(n10816), .ZN(n10901) );
  NAND2_X1 U10855 ( .A1(n10904), .A2(n10905), .ZN(n10816) );
  NAND2_X1 U10856 ( .A1(n10813), .A2(n10906), .ZN(n10905) );
  OR2_X1 U10857 ( .A1(n10812), .A2(n10811), .ZN(n10906) );
  NOR2_X1 U10858 ( .A1(n7606), .A2(n7702), .ZN(n10813) );
  NAND2_X1 U10859 ( .A1(n10811), .A2(n10812), .ZN(n10904) );
  NAND2_X1 U10860 ( .A1(n10907), .A2(n10908), .ZN(n10812) );
  NAND3_X1 U10861 ( .A1(a_14_), .A2(n10909), .A3(b_19_), .ZN(n10908) );
  NAND2_X1 U10862 ( .A1(n10808), .A2(n10807), .ZN(n10909) );
  OR2_X1 U10863 ( .A1(n10807), .A2(n10808), .ZN(n10907) );
  AND2_X1 U10864 ( .A1(n10910), .A2(n10911), .ZN(n10808) );
  NAND2_X1 U10865 ( .A1(n10805), .A2(n10912), .ZN(n10911) );
  OR2_X1 U10866 ( .A1(n10804), .A2(n10802), .ZN(n10912) );
  NOR2_X1 U10867 ( .A1(n7606), .A2(n7667), .ZN(n10805) );
  NAND2_X1 U10868 ( .A1(n10802), .A2(n10804), .ZN(n10910) );
  NAND2_X1 U10869 ( .A1(n10913), .A2(n10914), .ZN(n10804) );
  NAND3_X1 U10870 ( .A1(a_16_), .A2(n10915), .A3(b_19_), .ZN(n10914) );
  OR2_X1 U10871 ( .A1(n10800), .A2(n10798), .ZN(n10915) );
  NAND2_X1 U10872 ( .A1(n10798), .A2(n10800), .ZN(n10913) );
  NAND2_X1 U10873 ( .A1(n10916), .A2(n10917), .ZN(n10800) );
  NAND2_X1 U10874 ( .A1(n10797), .A2(n10918), .ZN(n10917) );
  OR2_X1 U10875 ( .A1(n10796), .A2(n10795), .ZN(n10918) );
  NOR2_X1 U10876 ( .A1(n7606), .A2(n7645), .ZN(n10797) );
  NAND2_X1 U10877 ( .A1(n10795), .A2(n10796), .ZN(n10916) );
  NAND2_X1 U10878 ( .A1(n10919), .A2(n10920), .ZN(n10796) );
  NAND3_X1 U10879 ( .A1(a_18_), .A2(n10921), .A3(b_19_), .ZN(n10920) );
  NAND2_X1 U10880 ( .A1(n10792), .A2(n10791), .ZN(n10921) );
  OR2_X1 U10881 ( .A1(n10791), .A2(n10792), .ZN(n10919) );
  AND2_X1 U10882 ( .A1(n10922), .A2(n10923), .ZN(n10792) );
  NAND2_X1 U10883 ( .A1(n7604), .A2(n10924), .ZN(n10923) );
  OR2_X1 U10884 ( .A1(n10789), .A2(n10788), .ZN(n10924) );
  INV_X1 U10885 ( .A(n7923), .ZN(n7604) );
  NAND2_X1 U10886 ( .A1(b_19_), .A2(a_19_), .ZN(n7923) );
  NAND2_X1 U10887 ( .A1(n10788), .A2(n10789), .ZN(n10922) );
  NAND2_X1 U10888 ( .A1(n10925), .A2(n10926), .ZN(n10789) );
  NAND3_X1 U10889 ( .A1(a_20_), .A2(n10927), .A3(b_19_), .ZN(n10926) );
  NAND2_X1 U10890 ( .A1(n10786), .A2(n10784), .ZN(n10927) );
  OR2_X1 U10891 ( .A1(n10784), .A2(n10786), .ZN(n10925) );
  AND2_X1 U10892 ( .A1(n10928), .A2(n10929), .ZN(n10786) );
  NAND2_X1 U10893 ( .A1(n10715), .A2(n10930), .ZN(n10929) );
  NAND2_X1 U10894 ( .A1(n10714), .A2(n10713), .ZN(n10930) );
  NOR2_X1 U10895 ( .A1(n7606), .A2(n7578), .ZN(n10715) );
  OR2_X1 U10896 ( .A1(n10713), .A2(n10714), .ZN(n10928) );
  AND2_X1 U10897 ( .A1(n10931), .A2(n10932), .ZN(n10714) );
  NAND3_X1 U10898 ( .A1(a_22_), .A2(n10933), .A3(b_19_), .ZN(n10932) );
  OR2_X1 U10899 ( .A1(n10781), .A2(n10779), .ZN(n10933) );
  NAND2_X1 U10900 ( .A1(n10779), .A2(n10781), .ZN(n10931) );
  NAND2_X1 U10901 ( .A1(n10934), .A2(n10935), .ZN(n10781) );
  NAND2_X1 U10902 ( .A1(n10778), .A2(n10936), .ZN(n10935) );
  OR2_X1 U10903 ( .A1(n10777), .A2(n10775), .ZN(n10936) );
  NOR2_X1 U10904 ( .A1(n7606), .A2(n7955), .ZN(n10778) );
  NAND2_X1 U10905 ( .A1(n10775), .A2(n10777), .ZN(n10934) );
  NAND2_X1 U10906 ( .A1(n10937), .A2(n10938), .ZN(n10777) );
  NAND3_X1 U10907 ( .A1(a_24_), .A2(n10939), .A3(b_19_), .ZN(n10938) );
  NAND2_X1 U10908 ( .A1(n10773), .A2(n10772), .ZN(n10939) );
  OR2_X1 U10909 ( .A1(n10772), .A2(n10773), .ZN(n10937) );
  AND2_X1 U10910 ( .A1(n10940), .A2(n10941), .ZN(n10773) );
  NAND2_X1 U10911 ( .A1(n10770), .A2(n10942), .ZN(n10941) );
  OR2_X1 U10912 ( .A1(n10769), .A2(n10768), .ZN(n10942) );
  NOR2_X1 U10913 ( .A1(n7606), .A2(n7952), .ZN(n10770) );
  NAND2_X1 U10914 ( .A1(n10768), .A2(n10769), .ZN(n10940) );
  NAND2_X1 U10915 ( .A1(n10765), .A2(n10943), .ZN(n10769) );
  NAND2_X1 U10916 ( .A1(n10764), .A2(n10766), .ZN(n10943) );
  NAND2_X1 U10917 ( .A1(n10944), .A2(n10945), .ZN(n10766) );
  NAND2_X1 U10918 ( .A1(b_19_), .A2(a_26_), .ZN(n10945) );
  INV_X1 U10919 ( .A(n10946), .ZN(n10944) );
  XNOR2_X1 U10920 ( .A(n10947), .B(n10948), .ZN(n10764) );
  NAND2_X1 U10921 ( .A1(n10949), .A2(n10950), .ZN(n10947) );
  NAND2_X1 U10922 ( .A1(a_26_), .A2(n10946), .ZN(n10765) );
  NAND2_X1 U10923 ( .A1(n10737), .A2(n10951), .ZN(n10946) );
  NAND2_X1 U10924 ( .A1(n10736), .A2(n10738), .ZN(n10951) );
  NAND2_X1 U10925 ( .A1(n10952), .A2(n10953), .ZN(n10738) );
  NAND2_X1 U10926 ( .A1(b_19_), .A2(a_27_), .ZN(n10953) );
  INV_X1 U10927 ( .A(n10954), .ZN(n10952) );
  XNOR2_X1 U10928 ( .A(n10955), .B(n10956), .ZN(n10736) );
  XOR2_X1 U10929 ( .A(n10957), .B(n10958), .Z(n10955) );
  NAND2_X1 U10930 ( .A1(b_18_), .A2(a_28_), .ZN(n10957) );
  NAND2_X1 U10931 ( .A1(a_27_), .A2(n10954), .ZN(n10737) );
  NAND2_X1 U10932 ( .A1(n10959), .A2(n10960), .ZN(n10954) );
  NAND3_X1 U10933 ( .A1(a_28_), .A2(n10961), .A3(b_19_), .ZN(n10960) );
  NAND2_X1 U10934 ( .A1(n10746), .A2(n10744), .ZN(n10961) );
  OR2_X1 U10935 ( .A1(n10744), .A2(n10746), .ZN(n10959) );
  AND2_X1 U10936 ( .A1(n10962), .A2(n10963), .ZN(n10746) );
  NAND2_X1 U10937 ( .A1(n10760), .A2(n10964), .ZN(n10963) );
  OR2_X1 U10938 ( .A1(n10761), .A2(n10762), .ZN(n10964) );
  NOR2_X1 U10939 ( .A1(n7606), .A2(n7460), .ZN(n10760) );
  INV_X1 U10940 ( .A(b_19_), .ZN(n7606) );
  NAND2_X1 U10941 ( .A1(n10762), .A2(n10761), .ZN(n10962) );
  NAND2_X1 U10942 ( .A1(n10965), .A2(n10966), .ZN(n10761) );
  NAND2_X1 U10943 ( .A1(b_17_), .A2(n10967), .ZN(n10966) );
  NAND2_X1 U10944 ( .A1(n7441), .A2(n10968), .ZN(n10967) );
  NAND2_X1 U10945 ( .A1(a_31_), .A2(n7959), .ZN(n10968) );
  NAND2_X1 U10946 ( .A1(b_18_), .A2(n10969), .ZN(n10965) );
  NAND2_X1 U10947 ( .A1(n7445), .A2(n10970), .ZN(n10969) );
  NAND2_X1 U10948 ( .A1(a_30_), .A2(n7638), .ZN(n10970) );
  AND3_X1 U10949 ( .A1(b_19_), .A2(n7409), .A3(b_18_), .ZN(n10762) );
  XNOR2_X1 U10950 ( .A(n10971), .B(n10972), .ZN(n10744) );
  XOR2_X1 U10951 ( .A(n10973), .B(n10974), .Z(n10971) );
  XNOR2_X1 U10952 ( .A(n10975), .B(n10976), .ZN(n10768) );
  NAND2_X1 U10953 ( .A1(n10977), .A2(n10978), .ZN(n10975) );
  XNOR2_X1 U10954 ( .A(n10979), .B(n10980), .ZN(n10772) );
  XOR2_X1 U10955 ( .A(n10981), .B(n10982), .Z(n10979) );
  XNOR2_X1 U10956 ( .A(n10983), .B(n10984), .ZN(n10775) );
  XNOR2_X1 U10957 ( .A(n10985), .B(n10986), .ZN(n10983) );
  NOR2_X1 U10958 ( .A1(n7954), .A2(n7959), .ZN(n10986) );
  XNOR2_X1 U10959 ( .A(n10987), .B(n10988), .ZN(n10779) );
  XOR2_X1 U10960 ( .A(n10989), .B(n10990), .Z(n10988) );
  NAND2_X1 U10961 ( .A1(b_18_), .A2(a_23_), .ZN(n10990) );
  XOR2_X1 U10962 ( .A(n10991), .B(n10992), .Z(n10713) );
  NAND2_X1 U10963 ( .A1(n10993), .A2(n10994), .ZN(n10991) );
  XNOR2_X1 U10964 ( .A(n10995), .B(n10996), .ZN(n10784) );
  XOR2_X1 U10965 ( .A(n10997), .B(n10998), .Z(n10995) );
  XNOR2_X1 U10966 ( .A(n10999), .B(n11000), .ZN(n10788) );
  XNOR2_X1 U10967 ( .A(n11001), .B(n11002), .ZN(n10999) );
  NOR2_X1 U10968 ( .A1(n7957), .A2(n7959), .ZN(n11002) );
  XOR2_X1 U10969 ( .A(n11003), .B(n11004), .Z(n10791) );
  XNOR2_X1 U10970 ( .A(n11005), .B(n11006), .ZN(n11004) );
  XOR2_X1 U10971 ( .A(n11007), .B(n11008), .Z(n10795) );
  XOR2_X1 U10972 ( .A(n11009), .B(n11010), .Z(n11007) );
  XNOR2_X1 U10973 ( .A(n11011), .B(n11012), .ZN(n10798) );
  XNOR2_X1 U10974 ( .A(n11013), .B(n11014), .ZN(n11012) );
  XNOR2_X1 U10975 ( .A(n11015), .B(n11016), .ZN(n10802) );
  XOR2_X1 U10976 ( .A(n11017), .B(n11018), .Z(n11016) );
  NAND2_X1 U10977 ( .A1(b_18_), .A2(a_16_), .ZN(n11018) );
  XOR2_X1 U10978 ( .A(n11019), .B(n11020), .Z(n10807) );
  XNOR2_X1 U10979 ( .A(n11021), .B(n11022), .ZN(n11020) );
  XNOR2_X1 U10980 ( .A(n11023), .B(n11024), .ZN(n10811) );
  XNOR2_X1 U10981 ( .A(n11025), .B(n11026), .ZN(n11023) );
  NOR2_X1 U10982 ( .A1(n7962), .A2(n7959), .ZN(n11026) );
  XNOR2_X1 U10983 ( .A(n11027), .B(n11028), .ZN(n10815) );
  XNOR2_X1 U10984 ( .A(n11029), .B(n11030), .ZN(n11027) );
  NOR2_X1 U10985 ( .A1(n7702), .A2(n7959), .ZN(n11030) );
  XNOR2_X1 U10986 ( .A(n11031), .B(n11032), .ZN(n10827) );
  XNOR2_X1 U10987 ( .A(n11033), .B(n11034), .ZN(n11031) );
  NOR2_X1 U10988 ( .A1(n8378), .A2(n7959), .ZN(n11034) );
  XNOR2_X1 U10989 ( .A(n11035), .B(n11036), .ZN(n10670) );
  NAND2_X1 U10990 ( .A1(n11037), .A2(n11038), .ZN(n11035) );
  XNOR2_X1 U10991 ( .A(n11039), .B(n11040), .ZN(n10661) );
  NAND2_X1 U10992 ( .A1(n11041), .A2(n11042), .ZN(n11039) );
  XOR2_X1 U10993 ( .A(n11043), .B(n11044), .Z(n10831) );
  NAND2_X1 U10994 ( .A1(n11045), .A2(n11046), .ZN(n11043) );
  XOR2_X1 U10995 ( .A(n11047), .B(n11048), .Z(n10835) );
  NAND2_X1 U10996 ( .A1(n11049), .A2(n11050), .ZN(n11047) );
  XNOR2_X1 U10997 ( .A(n11051), .B(n11052), .ZN(n10648) );
  NAND2_X1 U10998 ( .A1(n11053), .A2(n11054), .ZN(n11051) );
  XNOR2_X1 U10999 ( .A(n11055), .B(n11056), .ZN(n10639) );
  NAND2_X1 U11000 ( .A1(n11057), .A2(n11058), .ZN(n11055) );
  XNOR2_X1 U11001 ( .A(n11059), .B(n11060), .ZN(n10838) );
  NAND2_X1 U11002 ( .A1(n11061), .A2(n11062), .ZN(n11059) );
  XOR2_X1 U11003 ( .A(n11063), .B(n11064), .Z(n10843) );
  NAND2_X1 U11004 ( .A1(n11065), .A2(n11066), .ZN(n11063) );
  XNOR2_X1 U11005 ( .A(n11067), .B(n11068), .ZN(n10846) );
  XNOR2_X1 U11006 ( .A(n11069), .B(n11070), .ZN(n11068) );
  XOR2_X1 U11007 ( .A(n8140), .B(n8141), .Z(n10850) );
  NAND2_X1 U11008 ( .A1(n11071), .A2(n11072), .ZN(n8052) );
  NAND2_X1 U11009 ( .A1(n8141), .A2(n8140), .ZN(n11072) );
  XNOR2_X1 U11010 ( .A(n8131), .B(n8130), .ZN(n11071) );
  NAND3_X1 U11011 ( .A1(n11073), .A2(n8140), .A3(n8141), .ZN(n8051) );
  XNOR2_X1 U11012 ( .A(n11074), .B(n11075), .ZN(n8141) );
  XOR2_X1 U11013 ( .A(n11076), .B(n11077), .Z(n11075) );
  NAND2_X1 U11014 ( .A1(b_17_), .A2(a_0_), .ZN(n11077) );
  NAND2_X1 U11015 ( .A1(n11078), .A2(n11079), .ZN(n8140) );
  NAND3_X1 U11016 ( .A1(a_0_), .A2(n11080), .A3(b_18_), .ZN(n11079) );
  OR2_X1 U11017 ( .A1(n10852), .A2(n10853), .ZN(n11080) );
  NAND2_X1 U11018 ( .A1(n10852), .A2(n10853), .ZN(n11078) );
  NAND2_X1 U11019 ( .A1(n11081), .A2(n11082), .ZN(n10853) );
  NAND2_X1 U11020 ( .A1(n11070), .A2(n11083), .ZN(n11082) );
  OR2_X1 U11021 ( .A1(n11067), .A2(n11069), .ZN(n11083) );
  NOR2_X1 U11022 ( .A1(n7959), .A2(n7872), .ZN(n11070) );
  NAND2_X1 U11023 ( .A1(n11067), .A2(n11069), .ZN(n11081) );
  NAND2_X1 U11024 ( .A1(n11065), .A2(n11084), .ZN(n11069) );
  NAND2_X1 U11025 ( .A1(n11064), .A2(n11066), .ZN(n11084) );
  NAND2_X1 U11026 ( .A1(n11085), .A2(n11086), .ZN(n11066) );
  NAND2_X1 U11027 ( .A1(b_18_), .A2(a_2_), .ZN(n11086) );
  INV_X1 U11028 ( .A(n11087), .ZN(n11085) );
  XNOR2_X1 U11029 ( .A(n11088), .B(n11089), .ZN(n11064) );
  XOR2_X1 U11030 ( .A(n11090), .B(n11091), .Z(n11089) );
  NAND2_X1 U11031 ( .A1(b_17_), .A2(a_3_), .ZN(n11091) );
  NAND2_X1 U11032 ( .A1(a_2_), .A2(n11087), .ZN(n11065) );
  NAND2_X1 U11033 ( .A1(n11061), .A2(n11092), .ZN(n11087) );
  NAND2_X1 U11034 ( .A1(n11060), .A2(n11062), .ZN(n11092) );
  NAND2_X1 U11035 ( .A1(n11093), .A2(n11094), .ZN(n11062) );
  NAND2_X1 U11036 ( .A1(b_18_), .A2(a_3_), .ZN(n11094) );
  INV_X1 U11037 ( .A(n11095), .ZN(n11093) );
  XNOR2_X1 U11038 ( .A(n11096), .B(n11097), .ZN(n11060) );
  XOR2_X1 U11039 ( .A(n11098), .B(n11099), .Z(n11097) );
  NAND2_X1 U11040 ( .A1(b_17_), .A2(a_4_), .ZN(n11099) );
  NAND2_X1 U11041 ( .A1(a_3_), .A2(n11095), .ZN(n11061) );
  NAND2_X1 U11042 ( .A1(n11057), .A2(n11100), .ZN(n11095) );
  NAND2_X1 U11043 ( .A1(n11056), .A2(n11058), .ZN(n11100) );
  NAND2_X1 U11044 ( .A1(n11101), .A2(n11102), .ZN(n11058) );
  NAND2_X1 U11045 ( .A1(b_18_), .A2(a_4_), .ZN(n11102) );
  INV_X1 U11046 ( .A(n11103), .ZN(n11101) );
  XNOR2_X1 U11047 ( .A(n11104), .B(n11105), .ZN(n11056) );
  XOR2_X1 U11048 ( .A(n11106), .B(n11107), .Z(n11105) );
  NAND2_X1 U11049 ( .A1(b_17_), .A2(a_5_), .ZN(n11107) );
  NAND2_X1 U11050 ( .A1(a_4_), .A2(n11103), .ZN(n11057) );
  NAND2_X1 U11051 ( .A1(n11053), .A2(n11108), .ZN(n11103) );
  NAND2_X1 U11052 ( .A1(n11052), .A2(n11054), .ZN(n11108) );
  NAND2_X1 U11053 ( .A1(n11109), .A2(n11110), .ZN(n11054) );
  NAND2_X1 U11054 ( .A1(b_18_), .A2(a_5_), .ZN(n11110) );
  INV_X1 U11055 ( .A(n11111), .ZN(n11109) );
  XNOR2_X1 U11056 ( .A(n11112), .B(n11113), .ZN(n11052) );
  XOR2_X1 U11057 ( .A(n11114), .B(n11115), .Z(n11113) );
  NAND2_X1 U11058 ( .A1(b_17_), .A2(a_6_), .ZN(n11115) );
  NAND2_X1 U11059 ( .A1(a_5_), .A2(n11111), .ZN(n11053) );
  NAND2_X1 U11060 ( .A1(n11049), .A2(n11116), .ZN(n11111) );
  NAND2_X1 U11061 ( .A1(n11048), .A2(n11050), .ZN(n11116) );
  NAND2_X1 U11062 ( .A1(n11117), .A2(n11118), .ZN(n11050) );
  NAND2_X1 U11063 ( .A1(b_18_), .A2(a_6_), .ZN(n11118) );
  INV_X1 U11064 ( .A(n11119), .ZN(n11117) );
  XNOR2_X1 U11065 ( .A(n11120), .B(n11121), .ZN(n11048) );
  XOR2_X1 U11066 ( .A(n11122), .B(n11123), .Z(n11121) );
  NAND2_X1 U11067 ( .A1(b_17_), .A2(a_7_), .ZN(n11123) );
  NAND2_X1 U11068 ( .A1(a_6_), .A2(n11119), .ZN(n11049) );
  NAND2_X1 U11069 ( .A1(n11045), .A2(n11124), .ZN(n11119) );
  NAND2_X1 U11070 ( .A1(n11044), .A2(n11046), .ZN(n11124) );
  NAND2_X1 U11071 ( .A1(n11125), .A2(n11126), .ZN(n11046) );
  NAND2_X1 U11072 ( .A1(b_18_), .A2(a_7_), .ZN(n11126) );
  INV_X1 U11073 ( .A(n11127), .ZN(n11125) );
  XNOR2_X1 U11074 ( .A(n11128), .B(n11129), .ZN(n11044) );
  XOR2_X1 U11075 ( .A(n11130), .B(n11131), .Z(n11129) );
  NAND2_X1 U11076 ( .A1(b_17_), .A2(a_8_), .ZN(n11131) );
  NAND2_X1 U11077 ( .A1(a_7_), .A2(n11127), .ZN(n11045) );
  NAND2_X1 U11078 ( .A1(n11041), .A2(n11132), .ZN(n11127) );
  NAND2_X1 U11079 ( .A1(n11040), .A2(n11042), .ZN(n11132) );
  NAND2_X1 U11080 ( .A1(n11133), .A2(n11134), .ZN(n11042) );
  NAND2_X1 U11081 ( .A1(b_18_), .A2(a_8_), .ZN(n11134) );
  INV_X1 U11082 ( .A(n11135), .ZN(n11133) );
  XNOR2_X1 U11083 ( .A(n11136), .B(n11137), .ZN(n11040) );
  XNOR2_X1 U11084 ( .A(n11138), .B(n11139), .ZN(n11136) );
  NOR2_X1 U11085 ( .A1(n7753), .A2(n7638), .ZN(n11139) );
  NAND2_X1 U11086 ( .A1(a_8_), .A2(n11135), .ZN(n11041) );
  NAND2_X1 U11087 ( .A1(n11037), .A2(n11140), .ZN(n11135) );
  NAND2_X1 U11088 ( .A1(n11036), .A2(n11038), .ZN(n11140) );
  NAND2_X1 U11089 ( .A1(n11141), .A2(n11142), .ZN(n11038) );
  NAND2_X1 U11090 ( .A1(b_18_), .A2(a_9_), .ZN(n11142) );
  INV_X1 U11091 ( .A(n11143), .ZN(n11141) );
  XNOR2_X1 U11092 ( .A(n11144), .B(n11145), .ZN(n11036) );
  XNOR2_X1 U11093 ( .A(n11146), .B(n11147), .ZN(n11144) );
  NOR2_X1 U11094 ( .A1(n8378), .A2(n7638), .ZN(n11147) );
  NAND2_X1 U11095 ( .A1(a_9_), .A2(n11143), .ZN(n11037) );
  NAND2_X1 U11096 ( .A1(n11148), .A2(n11149), .ZN(n11143) );
  NAND3_X1 U11097 ( .A1(a_10_), .A2(n11150), .A3(b_18_), .ZN(n11149) );
  NAND2_X1 U11098 ( .A1(n11033), .A2(n11032), .ZN(n11150) );
  OR2_X1 U11099 ( .A1(n11032), .A2(n11033), .ZN(n11148) );
  AND2_X1 U11100 ( .A1(n11151), .A2(n11152), .ZN(n11033) );
  NAND2_X1 U11101 ( .A1(n10891), .A2(n11153), .ZN(n11152) );
  NAND2_X1 U11102 ( .A1(n10892), .A2(n10890), .ZN(n11153) );
  NOR2_X1 U11103 ( .A1(n7959), .A2(n7724), .ZN(n10891) );
  OR2_X1 U11104 ( .A1(n10890), .A2(n10892), .ZN(n11151) );
  AND2_X1 U11105 ( .A1(n11154), .A2(n11155), .ZN(n10892) );
  NAND2_X1 U11106 ( .A1(n10900), .A2(n11156), .ZN(n11155) );
  OR2_X1 U11107 ( .A1(n10897), .A2(n10899), .ZN(n11156) );
  NOR2_X1 U11108 ( .A1(n7959), .A2(n8585), .ZN(n10900) );
  NAND2_X1 U11109 ( .A1(n10897), .A2(n10899), .ZN(n11154) );
  NAND2_X1 U11110 ( .A1(n11157), .A2(n11158), .ZN(n10899) );
  NAND3_X1 U11111 ( .A1(a_13_), .A2(n11159), .A3(b_18_), .ZN(n11158) );
  NAND2_X1 U11112 ( .A1(n11029), .A2(n11028), .ZN(n11159) );
  OR2_X1 U11113 ( .A1(n11028), .A2(n11029), .ZN(n11157) );
  AND2_X1 U11114 ( .A1(n11160), .A2(n11161), .ZN(n11029) );
  NAND3_X1 U11115 ( .A1(a_14_), .A2(n11162), .A3(b_18_), .ZN(n11161) );
  NAND2_X1 U11116 ( .A1(n11025), .A2(n11024), .ZN(n11162) );
  OR2_X1 U11117 ( .A1(n11024), .A2(n11025), .ZN(n11160) );
  AND2_X1 U11118 ( .A1(n11163), .A2(n11164), .ZN(n11025) );
  NAND2_X1 U11119 ( .A1(n11022), .A2(n11165), .ZN(n11164) );
  OR2_X1 U11120 ( .A1(n11019), .A2(n11021), .ZN(n11165) );
  NOR2_X1 U11121 ( .A1(n7959), .A2(n7667), .ZN(n11022) );
  NAND2_X1 U11122 ( .A1(n11019), .A2(n11021), .ZN(n11163) );
  NAND2_X1 U11123 ( .A1(n11166), .A2(n11167), .ZN(n11021) );
  NAND3_X1 U11124 ( .A1(a_16_), .A2(n11168), .A3(b_18_), .ZN(n11167) );
  OR2_X1 U11125 ( .A1(n11017), .A2(n11015), .ZN(n11168) );
  NAND2_X1 U11126 ( .A1(n11015), .A2(n11017), .ZN(n11166) );
  NAND2_X1 U11127 ( .A1(n11169), .A2(n11170), .ZN(n11017) );
  NAND2_X1 U11128 ( .A1(n11014), .A2(n11171), .ZN(n11170) );
  OR2_X1 U11129 ( .A1(n11011), .A2(n11013), .ZN(n11171) );
  NOR2_X1 U11130 ( .A1(n7959), .A2(n7645), .ZN(n11014) );
  NAND2_X1 U11131 ( .A1(n11011), .A2(n11013), .ZN(n11169) );
  NAND2_X1 U11132 ( .A1(n11172), .A2(n11173), .ZN(n11013) );
  NAND2_X1 U11133 ( .A1(n11008), .A2(n11174), .ZN(n11173) );
  OR2_X1 U11134 ( .A1(n11009), .A2(n11010), .ZN(n11174) );
  XNOR2_X1 U11135 ( .A(n11175), .B(n11176), .ZN(n11008) );
  XNOR2_X1 U11136 ( .A(n11177), .B(n11178), .ZN(n11176) );
  NAND2_X1 U11137 ( .A1(n11010), .A2(n11009), .ZN(n11172) );
  NAND2_X1 U11138 ( .A1(n11179), .A2(n11180), .ZN(n11009) );
  NAND2_X1 U11139 ( .A1(n11006), .A2(n11181), .ZN(n11180) );
  OR2_X1 U11140 ( .A1(n11003), .A2(n11005), .ZN(n11181) );
  NOR2_X1 U11141 ( .A1(n7959), .A2(n7958), .ZN(n11006) );
  NAND2_X1 U11142 ( .A1(n11003), .A2(n11005), .ZN(n11179) );
  NAND2_X1 U11143 ( .A1(n11182), .A2(n11183), .ZN(n11005) );
  NAND3_X1 U11144 ( .A1(a_20_), .A2(n11184), .A3(b_18_), .ZN(n11183) );
  NAND2_X1 U11145 ( .A1(n11001), .A2(n11000), .ZN(n11184) );
  OR2_X1 U11146 ( .A1(n11000), .A2(n11001), .ZN(n11182) );
  AND2_X1 U11147 ( .A1(n11185), .A2(n11186), .ZN(n11001) );
  NAND2_X1 U11148 ( .A1(n10997), .A2(n11187), .ZN(n11186) );
  OR2_X1 U11149 ( .A1(n10996), .A2(n10998), .ZN(n11187) );
  NOR2_X1 U11150 ( .A1(n7959), .A2(n7578), .ZN(n10997) );
  NAND2_X1 U11151 ( .A1(n10996), .A2(n10998), .ZN(n11185) );
  NAND2_X1 U11152 ( .A1(n10993), .A2(n11188), .ZN(n10998) );
  NAND2_X1 U11153 ( .A1(n10992), .A2(n10994), .ZN(n11188) );
  NAND2_X1 U11154 ( .A1(n11189), .A2(n11190), .ZN(n10994) );
  NAND2_X1 U11155 ( .A1(b_18_), .A2(a_22_), .ZN(n11190) );
  INV_X1 U11156 ( .A(n11191), .ZN(n11189) );
  XNOR2_X1 U11157 ( .A(n11192), .B(n11193), .ZN(n10992) );
  XNOR2_X1 U11158 ( .A(n11194), .B(n11195), .ZN(n11193) );
  NAND2_X1 U11159 ( .A1(a_22_), .A2(n11191), .ZN(n10993) );
  NAND2_X1 U11160 ( .A1(n11196), .A2(n11197), .ZN(n11191) );
  NAND3_X1 U11161 ( .A1(a_23_), .A2(n11198), .A3(b_18_), .ZN(n11197) );
  OR2_X1 U11162 ( .A1(n10987), .A2(n10989), .ZN(n11198) );
  NAND2_X1 U11163 ( .A1(n10987), .A2(n10989), .ZN(n11196) );
  NAND2_X1 U11164 ( .A1(n11199), .A2(n11200), .ZN(n10989) );
  NAND3_X1 U11165 ( .A1(a_24_), .A2(n11201), .A3(b_18_), .ZN(n11200) );
  NAND2_X1 U11166 ( .A1(n10985), .A2(n10984), .ZN(n11201) );
  OR2_X1 U11167 ( .A1(n10984), .A2(n10985), .ZN(n11199) );
  AND2_X1 U11168 ( .A1(n11202), .A2(n11203), .ZN(n10985) );
  NAND2_X1 U11169 ( .A1(n10982), .A2(n11204), .ZN(n11203) );
  OR2_X1 U11170 ( .A1(n10980), .A2(n10981), .ZN(n11204) );
  NOR2_X1 U11171 ( .A1(n7959), .A2(n7952), .ZN(n10982) );
  NAND2_X1 U11172 ( .A1(n10980), .A2(n10981), .ZN(n11202) );
  NAND2_X1 U11173 ( .A1(n10977), .A2(n11205), .ZN(n10981) );
  NAND2_X1 U11174 ( .A1(n10976), .A2(n10978), .ZN(n11205) );
  NAND2_X1 U11175 ( .A1(n11206), .A2(n11207), .ZN(n10978) );
  NAND2_X1 U11176 ( .A1(b_18_), .A2(a_26_), .ZN(n11207) );
  INV_X1 U11177 ( .A(n11208), .ZN(n11206) );
  XNOR2_X1 U11178 ( .A(n11209), .B(n11210), .ZN(n10976) );
  NAND2_X1 U11179 ( .A1(n11211), .A2(n11212), .ZN(n11209) );
  NAND2_X1 U11180 ( .A1(a_26_), .A2(n11208), .ZN(n10977) );
  NAND2_X1 U11181 ( .A1(n10949), .A2(n11213), .ZN(n11208) );
  NAND2_X1 U11182 ( .A1(n10948), .A2(n10950), .ZN(n11213) );
  NAND2_X1 U11183 ( .A1(n11214), .A2(n11215), .ZN(n10950) );
  NAND2_X1 U11184 ( .A1(b_18_), .A2(a_27_), .ZN(n11215) );
  INV_X1 U11185 ( .A(n11216), .ZN(n11214) );
  XNOR2_X1 U11186 ( .A(n11217), .B(n11218), .ZN(n10948) );
  XOR2_X1 U11187 ( .A(n11219), .B(n11220), .Z(n11217) );
  NAND2_X1 U11188 ( .A1(b_17_), .A2(a_28_), .ZN(n11219) );
  NAND2_X1 U11189 ( .A1(a_27_), .A2(n11216), .ZN(n10949) );
  NAND2_X1 U11190 ( .A1(n11221), .A2(n11222), .ZN(n11216) );
  NAND3_X1 U11191 ( .A1(a_28_), .A2(n11223), .A3(b_18_), .ZN(n11222) );
  NAND2_X1 U11192 ( .A1(n10958), .A2(n10956), .ZN(n11223) );
  OR2_X1 U11193 ( .A1(n10956), .A2(n10958), .ZN(n11221) );
  AND2_X1 U11194 ( .A1(n11224), .A2(n11225), .ZN(n10958) );
  NAND2_X1 U11195 ( .A1(n10972), .A2(n11226), .ZN(n11225) );
  OR2_X1 U11196 ( .A1(n10973), .A2(n10974), .ZN(n11226) );
  NOR2_X1 U11197 ( .A1(n7959), .A2(n7460), .ZN(n10972) );
  INV_X1 U11198 ( .A(b_18_), .ZN(n7959) );
  NAND2_X1 U11199 ( .A1(n10974), .A2(n10973), .ZN(n11224) );
  NAND2_X1 U11200 ( .A1(n11227), .A2(n11228), .ZN(n10973) );
  NAND2_X1 U11201 ( .A1(b_16_), .A2(n11229), .ZN(n11228) );
  NAND2_X1 U11202 ( .A1(n7441), .A2(n11230), .ZN(n11229) );
  NAND2_X1 U11203 ( .A1(a_31_), .A2(n7638), .ZN(n11230) );
  NAND2_X1 U11204 ( .A1(b_17_), .A2(n11231), .ZN(n11227) );
  NAND2_X1 U11205 ( .A1(n7445), .A2(n11232), .ZN(n11231) );
  NAND2_X1 U11206 ( .A1(a_30_), .A2(n11233), .ZN(n11232) );
  AND3_X1 U11207 ( .A1(b_17_), .A2(n7409), .A3(b_18_), .ZN(n10974) );
  XNOR2_X1 U11208 ( .A(n11234), .B(n11235), .ZN(n10956) );
  XOR2_X1 U11209 ( .A(n11236), .B(n11237), .Z(n11234) );
  XNOR2_X1 U11210 ( .A(n11238), .B(n11239), .ZN(n10980) );
  NAND2_X1 U11211 ( .A1(n11240), .A2(n11241), .ZN(n11238) );
  XNOR2_X1 U11212 ( .A(n11242), .B(n11243), .ZN(n10984) );
  XOR2_X1 U11213 ( .A(n11244), .B(n11245), .Z(n11242) );
  XNOR2_X1 U11214 ( .A(n11246), .B(n11247), .ZN(n10987) );
  XNOR2_X1 U11215 ( .A(n11248), .B(n11249), .ZN(n11246) );
  NOR2_X1 U11216 ( .A1(n7954), .A2(n7638), .ZN(n11249) );
  XNOR2_X1 U11217 ( .A(n11250), .B(n11251), .ZN(n10996) );
  XOR2_X1 U11218 ( .A(n11252), .B(n11253), .Z(n11251) );
  NAND2_X1 U11219 ( .A1(b_17_), .A2(a_22_), .ZN(n11253) );
  XNOR2_X1 U11220 ( .A(n11254), .B(n11255), .ZN(n11000) );
  XOR2_X1 U11221 ( .A(n11256), .B(n11257), .Z(n11254) );
  XNOR2_X1 U11222 ( .A(n11258), .B(n11259), .ZN(n11003) );
  XNOR2_X1 U11223 ( .A(n11260), .B(n11261), .ZN(n11258) );
  NOR2_X1 U11224 ( .A1(n7957), .A2(n7638), .ZN(n11261) );
  INV_X1 U11225 ( .A(n7619), .ZN(n11010) );
  NAND2_X1 U11226 ( .A1(b_18_), .A2(a_18_), .ZN(n7619) );
  XNOR2_X1 U11227 ( .A(n11262), .B(n11263), .ZN(n11011) );
  XNOR2_X1 U11228 ( .A(n11264), .B(n11265), .ZN(n11262) );
  NOR2_X1 U11229 ( .A1(n7960), .A2(n7638), .ZN(n11265) );
  XOR2_X1 U11230 ( .A(n11266), .B(n11267), .Z(n11015) );
  XOR2_X1 U11231 ( .A(n11268), .B(n7636), .Z(n11266) );
  XNOR2_X1 U11232 ( .A(n11269), .B(n11270), .ZN(n11019) );
  XOR2_X1 U11233 ( .A(n11271), .B(n11272), .Z(n11270) );
  NAND2_X1 U11234 ( .A1(b_17_), .A2(a_16_), .ZN(n11272) );
  XOR2_X1 U11235 ( .A(n11273), .B(n11274), .Z(n11024) );
  XNOR2_X1 U11236 ( .A(n11275), .B(n11276), .ZN(n11274) );
  XNOR2_X1 U11237 ( .A(n11277), .B(n11278), .ZN(n11028) );
  XOR2_X1 U11238 ( .A(n11279), .B(n11280), .Z(n11277) );
  XNOR2_X1 U11239 ( .A(n11281), .B(n11282), .ZN(n10897) );
  XNOR2_X1 U11240 ( .A(n11283), .B(n11284), .ZN(n11281) );
  NOR2_X1 U11241 ( .A1(n7702), .A2(n7638), .ZN(n11284) );
  XOR2_X1 U11242 ( .A(n11285), .B(n11286), .Z(n10890) );
  XOR2_X1 U11243 ( .A(n11287), .B(n11288), .Z(n11286) );
  NAND2_X1 U11244 ( .A1(b_17_), .A2(a_12_), .ZN(n11288) );
  XOR2_X1 U11245 ( .A(n11289), .B(n11290), .Z(n11032) );
  XOR2_X1 U11246 ( .A(n11291), .B(n11292), .Z(n11290) );
  NAND2_X1 U11247 ( .A1(b_17_), .A2(a_11_), .ZN(n11292) );
  XNOR2_X1 U11248 ( .A(n11293), .B(n11294), .ZN(n11067) );
  XOR2_X1 U11249 ( .A(n11295), .B(n11296), .Z(n11294) );
  NAND2_X1 U11250 ( .A1(b_17_), .A2(a_2_), .ZN(n11296) );
  XNOR2_X1 U11251 ( .A(n11297), .B(n11298), .ZN(n10852) );
  XOR2_X1 U11252 ( .A(n11299), .B(n11300), .Z(n11298) );
  NAND2_X1 U11253 ( .A1(b_17_), .A2(a_1_), .ZN(n11300) );
  XOR2_X1 U11254 ( .A(n8131), .B(n8130), .Z(n11073) );
  NAND3_X1 U11255 ( .A1(n8130), .A2(n8131), .A3(n11301), .ZN(n8056) );
  XOR2_X1 U11256 ( .A(n8133), .B(n8132), .Z(n11301) );
  NAND2_X1 U11257 ( .A1(n11302), .A2(n11303), .ZN(n8131) );
  NAND3_X1 U11258 ( .A1(a_0_), .A2(n11304), .A3(b_17_), .ZN(n11303) );
  OR2_X1 U11259 ( .A1(n11076), .A2(n11074), .ZN(n11304) );
  NAND2_X1 U11260 ( .A1(n11074), .A2(n11076), .ZN(n11302) );
  NAND2_X1 U11261 ( .A1(n11305), .A2(n11306), .ZN(n11076) );
  NAND3_X1 U11262 ( .A1(a_1_), .A2(n11307), .A3(b_17_), .ZN(n11306) );
  OR2_X1 U11263 ( .A1(n11299), .A2(n11297), .ZN(n11307) );
  NAND2_X1 U11264 ( .A1(n11297), .A2(n11299), .ZN(n11305) );
  NAND2_X1 U11265 ( .A1(n11308), .A2(n11309), .ZN(n11299) );
  NAND3_X1 U11266 ( .A1(a_2_), .A2(n11310), .A3(b_17_), .ZN(n11309) );
  OR2_X1 U11267 ( .A1(n11295), .A2(n11293), .ZN(n11310) );
  NAND2_X1 U11268 ( .A1(n11293), .A2(n11295), .ZN(n11308) );
  NAND2_X1 U11269 ( .A1(n11311), .A2(n11312), .ZN(n11295) );
  NAND3_X1 U11270 ( .A1(a_3_), .A2(n11313), .A3(b_17_), .ZN(n11312) );
  OR2_X1 U11271 ( .A1(n11090), .A2(n11088), .ZN(n11313) );
  NAND2_X1 U11272 ( .A1(n11088), .A2(n11090), .ZN(n11311) );
  NAND2_X1 U11273 ( .A1(n11314), .A2(n11315), .ZN(n11090) );
  NAND3_X1 U11274 ( .A1(a_4_), .A2(n11316), .A3(b_17_), .ZN(n11315) );
  OR2_X1 U11275 ( .A1(n11098), .A2(n11096), .ZN(n11316) );
  NAND2_X1 U11276 ( .A1(n11096), .A2(n11098), .ZN(n11314) );
  NAND2_X1 U11277 ( .A1(n11317), .A2(n11318), .ZN(n11098) );
  NAND3_X1 U11278 ( .A1(a_5_), .A2(n11319), .A3(b_17_), .ZN(n11318) );
  OR2_X1 U11279 ( .A1(n11106), .A2(n11104), .ZN(n11319) );
  NAND2_X1 U11280 ( .A1(n11104), .A2(n11106), .ZN(n11317) );
  NAND2_X1 U11281 ( .A1(n11320), .A2(n11321), .ZN(n11106) );
  NAND3_X1 U11282 ( .A1(a_6_), .A2(n11322), .A3(b_17_), .ZN(n11321) );
  OR2_X1 U11283 ( .A1(n11114), .A2(n11112), .ZN(n11322) );
  NAND2_X1 U11284 ( .A1(n11112), .A2(n11114), .ZN(n11320) );
  NAND2_X1 U11285 ( .A1(n11323), .A2(n11324), .ZN(n11114) );
  NAND3_X1 U11286 ( .A1(a_7_), .A2(n11325), .A3(b_17_), .ZN(n11324) );
  OR2_X1 U11287 ( .A1(n11122), .A2(n11120), .ZN(n11325) );
  NAND2_X1 U11288 ( .A1(n11120), .A2(n11122), .ZN(n11323) );
  NAND2_X1 U11289 ( .A1(n11326), .A2(n11327), .ZN(n11122) );
  NAND3_X1 U11290 ( .A1(a_8_), .A2(n11328), .A3(b_17_), .ZN(n11327) );
  OR2_X1 U11291 ( .A1(n11130), .A2(n11128), .ZN(n11328) );
  NAND2_X1 U11292 ( .A1(n11128), .A2(n11130), .ZN(n11326) );
  NAND2_X1 U11293 ( .A1(n11329), .A2(n11330), .ZN(n11130) );
  NAND3_X1 U11294 ( .A1(a_9_), .A2(n11331), .A3(b_17_), .ZN(n11330) );
  NAND2_X1 U11295 ( .A1(n11138), .A2(n11137), .ZN(n11331) );
  OR2_X1 U11296 ( .A1(n11137), .A2(n11138), .ZN(n11329) );
  AND2_X1 U11297 ( .A1(n11332), .A2(n11333), .ZN(n11138) );
  NAND3_X1 U11298 ( .A1(a_10_), .A2(n11334), .A3(b_17_), .ZN(n11333) );
  NAND2_X1 U11299 ( .A1(n11146), .A2(n11145), .ZN(n11334) );
  OR2_X1 U11300 ( .A1(n11145), .A2(n11146), .ZN(n11332) );
  AND2_X1 U11301 ( .A1(n11335), .A2(n11336), .ZN(n11146) );
  NAND3_X1 U11302 ( .A1(a_11_), .A2(n11337), .A3(b_17_), .ZN(n11336) );
  OR2_X1 U11303 ( .A1(n11291), .A2(n11289), .ZN(n11337) );
  NAND2_X1 U11304 ( .A1(n11289), .A2(n11291), .ZN(n11335) );
  NAND2_X1 U11305 ( .A1(n11338), .A2(n11339), .ZN(n11291) );
  NAND3_X1 U11306 ( .A1(a_12_), .A2(n11340), .A3(b_17_), .ZN(n11339) );
  OR2_X1 U11307 ( .A1(n11287), .A2(n11285), .ZN(n11340) );
  NAND2_X1 U11308 ( .A1(n11285), .A2(n11287), .ZN(n11338) );
  NAND2_X1 U11309 ( .A1(n11341), .A2(n11342), .ZN(n11287) );
  NAND3_X1 U11310 ( .A1(a_13_), .A2(n11343), .A3(b_17_), .ZN(n11342) );
  NAND2_X1 U11311 ( .A1(n11283), .A2(n11282), .ZN(n11343) );
  OR2_X1 U11312 ( .A1(n11282), .A2(n11283), .ZN(n11341) );
  AND2_X1 U11313 ( .A1(n11344), .A2(n11345), .ZN(n11283) );
  NAND2_X1 U11314 ( .A1(n11280), .A2(n11346), .ZN(n11345) );
  OR2_X1 U11315 ( .A1(n11279), .A2(n11278), .ZN(n11346) );
  NOR2_X1 U11316 ( .A1(n7638), .A2(n7962), .ZN(n11280) );
  NAND2_X1 U11317 ( .A1(n11278), .A2(n11279), .ZN(n11344) );
  NAND2_X1 U11318 ( .A1(n11347), .A2(n11348), .ZN(n11279) );
  NAND2_X1 U11319 ( .A1(n11276), .A2(n11349), .ZN(n11348) );
  OR2_X1 U11320 ( .A1(n11275), .A2(n11273), .ZN(n11349) );
  NOR2_X1 U11321 ( .A1(n7638), .A2(n7667), .ZN(n11276) );
  NAND2_X1 U11322 ( .A1(n11273), .A2(n11275), .ZN(n11347) );
  NAND2_X1 U11323 ( .A1(n11350), .A2(n11351), .ZN(n11275) );
  NAND3_X1 U11324 ( .A1(a_16_), .A2(n11352), .A3(b_17_), .ZN(n11351) );
  OR2_X1 U11325 ( .A1(n11271), .A2(n11269), .ZN(n11352) );
  NAND2_X1 U11326 ( .A1(n11269), .A2(n11271), .ZN(n11350) );
  NAND2_X1 U11327 ( .A1(n11353), .A2(n11354), .ZN(n11271) );
  NAND2_X1 U11328 ( .A1(n7636), .A2(n11355), .ZN(n11354) );
  OR2_X1 U11329 ( .A1(n11268), .A2(n11267), .ZN(n11355) );
  INV_X1 U11330 ( .A(n7919), .ZN(n7636) );
  NAND2_X1 U11331 ( .A1(b_17_), .A2(a_17_), .ZN(n7919) );
  NAND2_X1 U11332 ( .A1(n11267), .A2(n11268), .ZN(n11353) );
  NAND2_X1 U11333 ( .A1(n11356), .A2(n11357), .ZN(n11268) );
  NAND3_X1 U11334 ( .A1(a_18_), .A2(n11358), .A3(b_17_), .ZN(n11357) );
  NAND2_X1 U11335 ( .A1(n11264), .A2(n11263), .ZN(n11358) );
  OR2_X1 U11336 ( .A1(n11263), .A2(n11264), .ZN(n11356) );
  AND2_X1 U11337 ( .A1(n11359), .A2(n11360), .ZN(n11264) );
  NAND2_X1 U11338 ( .A1(n11178), .A2(n11361), .ZN(n11360) );
  OR2_X1 U11339 ( .A1(n11177), .A2(n11175), .ZN(n11361) );
  NOR2_X1 U11340 ( .A1(n7638), .A2(n7958), .ZN(n11178) );
  NAND2_X1 U11341 ( .A1(n11175), .A2(n11177), .ZN(n11359) );
  NAND2_X1 U11342 ( .A1(n11362), .A2(n11363), .ZN(n11177) );
  NAND3_X1 U11343 ( .A1(a_20_), .A2(n11364), .A3(b_17_), .ZN(n11363) );
  NAND2_X1 U11344 ( .A1(n11260), .A2(n11259), .ZN(n11364) );
  OR2_X1 U11345 ( .A1(n11259), .A2(n11260), .ZN(n11362) );
  AND2_X1 U11346 ( .A1(n11365), .A2(n11366), .ZN(n11260) );
  NAND2_X1 U11347 ( .A1(n11257), .A2(n11367), .ZN(n11366) );
  OR2_X1 U11348 ( .A1(n11256), .A2(n11255), .ZN(n11367) );
  NOR2_X1 U11349 ( .A1(n7638), .A2(n7578), .ZN(n11257) );
  NAND2_X1 U11350 ( .A1(n11255), .A2(n11256), .ZN(n11365) );
  NAND2_X1 U11351 ( .A1(n11368), .A2(n11369), .ZN(n11256) );
  NAND3_X1 U11352 ( .A1(a_22_), .A2(n11370), .A3(b_17_), .ZN(n11369) );
  OR2_X1 U11353 ( .A1(n11252), .A2(n11250), .ZN(n11370) );
  NAND2_X1 U11354 ( .A1(n11250), .A2(n11252), .ZN(n11368) );
  NAND2_X1 U11355 ( .A1(n11371), .A2(n11372), .ZN(n11252) );
  NAND2_X1 U11356 ( .A1(n11195), .A2(n11373), .ZN(n11372) );
  OR2_X1 U11357 ( .A1(n11194), .A2(n11192), .ZN(n11373) );
  NOR2_X1 U11358 ( .A1(n7638), .A2(n7955), .ZN(n11195) );
  NAND2_X1 U11359 ( .A1(n11192), .A2(n11194), .ZN(n11371) );
  NAND2_X1 U11360 ( .A1(n11374), .A2(n11375), .ZN(n11194) );
  NAND3_X1 U11361 ( .A1(a_24_), .A2(n11376), .A3(b_17_), .ZN(n11375) );
  NAND2_X1 U11362 ( .A1(n11248), .A2(n11247), .ZN(n11376) );
  OR2_X1 U11363 ( .A1(n11247), .A2(n11248), .ZN(n11374) );
  AND2_X1 U11364 ( .A1(n11377), .A2(n11378), .ZN(n11248) );
  NAND2_X1 U11365 ( .A1(n11245), .A2(n11379), .ZN(n11378) );
  OR2_X1 U11366 ( .A1(n11244), .A2(n11243), .ZN(n11379) );
  NOR2_X1 U11367 ( .A1(n7638), .A2(n7952), .ZN(n11245) );
  NAND2_X1 U11368 ( .A1(n11243), .A2(n11244), .ZN(n11377) );
  NAND2_X1 U11369 ( .A1(n11240), .A2(n11380), .ZN(n11244) );
  NAND2_X1 U11370 ( .A1(n11239), .A2(n11241), .ZN(n11380) );
  NAND2_X1 U11371 ( .A1(n11381), .A2(n11382), .ZN(n11241) );
  NAND2_X1 U11372 ( .A1(b_17_), .A2(a_26_), .ZN(n11382) );
  INV_X1 U11373 ( .A(n11383), .ZN(n11381) );
  XNOR2_X1 U11374 ( .A(n11384), .B(n11385), .ZN(n11239) );
  NAND2_X1 U11375 ( .A1(n11386), .A2(n11387), .ZN(n11384) );
  NAND2_X1 U11376 ( .A1(a_26_), .A2(n11383), .ZN(n11240) );
  NAND2_X1 U11377 ( .A1(n11211), .A2(n11388), .ZN(n11383) );
  NAND2_X1 U11378 ( .A1(n11210), .A2(n11212), .ZN(n11388) );
  NAND2_X1 U11379 ( .A1(n11389), .A2(n11390), .ZN(n11212) );
  NAND2_X1 U11380 ( .A1(b_17_), .A2(a_27_), .ZN(n11390) );
  INV_X1 U11381 ( .A(n11391), .ZN(n11389) );
  XNOR2_X1 U11382 ( .A(n11392), .B(n11393), .ZN(n11210) );
  XOR2_X1 U11383 ( .A(n11394), .B(n11395), .Z(n11392) );
  NAND2_X1 U11384 ( .A1(b_16_), .A2(a_28_), .ZN(n11394) );
  NAND2_X1 U11385 ( .A1(a_27_), .A2(n11391), .ZN(n11211) );
  NAND2_X1 U11386 ( .A1(n11396), .A2(n11397), .ZN(n11391) );
  NAND3_X1 U11387 ( .A1(a_28_), .A2(n11398), .A3(b_17_), .ZN(n11397) );
  NAND2_X1 U11388 ( .A1(n11220), .A2(n11218), .ZN(n11398) );
  OR2_X1 U11389 ( .A1(n11218), .A2(n11220), .ZN(n11396) );
  AND2_X1 U11390 ( .A1(n11399), .A2(n11400), .ZN(n11220) );
  NAND2_X1 U11391 ( .A1(n11235), .A2(n11401), .ZN(n11400) );
  OR2_X1 U11392 ( .A1(n11236), .A2(n11237), .ZN(n11401) );
  NOR2_X1 U11393 ( .A1(n7638), .A2(n7460), .ZN(n11235) );
  INV_X1 U11394 ( .A(b_17_), .ZN(n7638) );
  NAND2_X1 U11395 ( .A1(n11237), .A2(n11236), .ZN(n11399) );
  NAND2_X1 U11396 ( .A1(n11402), .A2(n11403), .ZN(n11236) );
  NAND2_X1 U11397 ( .A1(b_15_), .A2(n11404), .ZN(n11403) );
  NAND2_X1 U11398 ( .A1(n7441), .A2(n11405), .ZN(n11404) );
  NAND2_X1 U11399 ( .A1(a_31_), .A2(n11233), .ZN(n11405) );
  NAND2_X1 U11400 ( .A1(b_16_), .A2(n11406), .ZN(n11402) );
  NAND2_X1 U11401 ( .A1(n7445), .A2(n11407), .ZN(n11406) );
  NAND2_X1 U11402 ( .A1(a_30_), .A2(n7669), .ZN(n11407) );
  AND3_X1 U11403 ( .A1(b_17_), .A2(n7409), .A3(b_16_), .ZN(n11237) );
  XNOR2_X1 U11404 ( .A(n11408), .B(n11409), .ZN(n11218) );
  XOR2_X1 U11405 ( .A(n11410), .B(n11411), .Z(n11408) );
  XNOR2_X1 U11406 ( .A(n11412), .B(n11413), .ZN(n11243) );
  NAND2_X1 U11407 ( .A1(n11414), .A2(n11415), .ZN(n11412) );
  XNOR2_X1 U11408 ( .A(n11416), .B(n11417), .ZN(n11247) );
  XOR2_X1 U11409 ( .A(n11418), .B(n11419), .Z(n11416) );
  XNOR2_X1 U11410 ( .A(n11420), .B(n11421), .ZN(n11192) );
  XNOR2_X1 U11411 ( .A(n11422), .B(n11423), .ZN(n11420) );
  NOR2_X1 U11412 ( .A1(n7954), .A2(n11233), .ZN(n11423) );
  XNOR2_X1 U11413 ( .A(n11424), .B(n11425), .ZN(n11250) );
  XNOR2_X1 U11414 ( .A(n11426), .B(n11427), .ZN(n11425) );
  XNOR2_X1 U11415 ( .A(n11428), .B(n11429), .ZN(n11255) );
  XNOR2_X1 U11416 ( .A(n11430), .B(n11431), .ZN(n11428) );
  NOR2_X1 U11417 ( .A1(n7568), .A2(n11233), .ZN(n11431) );
  XNOR2_X1 U11418 ( .A(n11432), .B(n11433), .ZN(n11259) );
  XOR2_X1 U11419 ( .A(n11434), .B(n11435), .Z(n11432) );
  XNOR2_X1 U11420 ( .A(n11436), .B(n11437), .ZN(n11175) );
  XNOR2_X1 U11421 ( .A(n11438), .B(n11439), .ZN(n11436) );
  NOR2_X1 U11422 ( .A1(n7957), .A2(n11233), .ZN(n11439) );
  XOR2_X1 U11423 ( .A(n11440), .B(n11441), .Z(n11263) );
  XNOR2_X1 U11424 ( .A(n11442), .B(n11443), .ZN(n11441) );
  XNOR2_X1 U11425 ( .A(n11444), .B(n11445), .ZN(n11267) );
  XNOR2_X1 U11426 ( .A(n11446), .B(n11447), .ZN(n11444) );
  NOR2_X1 U11427 ( .A1(n7960), .A2(n11233), .ZN(n11447) );
  XOR2_X1 U11428 ( .A(n11448), .B(n11449), .Z(n11269) );
  XOR2_X1 U11429 ( .A(n11450), .B(n11451), .Z(n11448) );
  XNOR2_X1 U11430 ( .A(n11452), .B(n11453), .ZN(n11273) );
  XNOR2_X1 U11431 ( .A(n11454), .B(n7652), .ZN(n11453) );
  XNOR2_X1 U11432 ( .A(n11455), .B(n11456), .ZN(n11278) );
  NAND2_X1 U11433 ( .A1(n11457), .A2(n11458), .ZN(n11455) );
  XNOR2_X1 U11434 ( .A(n11459), .B(n11460), .ZN(n11282) );
  XOR2_X1 U11435 ( .A(n11461), .B(n11462), .Z(n11459) );
  XNOR2_X1 U11436 ( .A(n11463), .B(n11464), .ZN(n11285) );
  XNOR2_X1 U11437 ( .A(n11465), .B(n11466), .ZN(n11463) );
  XNOR2_X1 U11438 ( .A(n11467), .B(n11468), .ZN(n11289) );
  XNOR2_X1 U11439 ( .A(n11469), .B(n11470), .ZN(n11467) );
  XNOR2_X1 U11440 ( .A(n11471), .B(n11472), .ZN(n11145) );
  XOR2_X1 U11441 ( .A(n11473), .B(n11474), .Z(n11471) );
  XNOR2_X1 U11442 ( .A(n11475), .B(n11476), .ZN(n11137) );
  XOR2_X1 U11443 ( .A(n11477), .B(n11478), .Z(n11475) );
  XNOR2_X1 U11444 ( .A(n11479), .B(n11480), .ZN(n11128) );
  XNOR2_X1 U11445 ( .A(n11481), .B(n11482), .ZN(n11480) );
  XNOR2_X1 U11446 ( .A(n11483), .B(n11484), .ZN(n11120) );
  XNOR2_X1 U11447 ( .A(n11485), .B(n11486), .ZN(n11483) );
  NOR2_X1 U11448 ( .A1(n8602), .A2(n11233), .ZN(n11486) );
  XOR2_X1 U11449 ( .A(n11487), .B(n11488), .Z(n11112) );
  XOR2_X1 U11450 ( .A(n11489), .B(n11490), .Z(n11487) );
  XNOR2_X1 U11451 ( .A(n11491), .B(n11492), .ZN(n11104) );
  XOR2_X1 U11452 ( .A(n11493), .B(n11494), .Z(n11492) );
  NAND2_X1 U11453 ( .A1(b_16_), .A2(a_6_), .ZN(n11494) );
  XNOR2_X1 U11454 ( .A(n11495), .B(n11496), .ZN(n11096) );
  NAND2_X1 U11455 ( .A1(n11497), .A2(n11498), .ZN(n11495) );
  XNOR2_X1 U11456 ( .A(n11499), .B(n11500), .ZN(n11088) );
  XNOR2_X1 U11457 ( .A(n11501), .B(n11502), .ZN(n11499) );
  XOR2_X1 U11458 ( .A(n11503), .B(n11504), .Z(n11293) );
  XOR2_X1 U11459 ( .A(n11505), .B(n11506), .Z(n11503) );
  XOR2_X1 U11460 ( .A(n11507), .B(n11508), .Z(n11297) );
  XOR2_X1 U11461 ( .A(n11509), .B(n11510), .Z(n11507) );
  XNOR2_X1 U11462 ( .A(n11511), .B(n11512), .ZN(n11074) );
  XNOR2_X1 U11463 ( .A(n11513), .B(n11514), .ZN(n11511) );
  NOR2_X1 U11464 ( .A1(n7872), .A2(n11233), .ZN(n11514) );
  XNOR2_X1 U11465 ( .A(n11515), .B(n11516), .ZN(n8130) );
  NAND2_X1 U11466 ( .A1(n11517), .A2(n11518), .ZN(n11515) );
  NAND2_X1 U11467 ( .A1(n11519), .A2(n11520), .ZN(n8062) );
  NAND2_X1 U11468 ( .A1(n8133), .A2(n8132), .ZN(n11520) );
  XOR2_X1 U11469 ( .A(n11521), .B(n11522), .Z(n11519) );
  NAND3_X1 U11470 ( .A1(n8133), .A2(n8132), .A3(n11523), .ZN(n8061) );
  XOR2_X1 U11471 ( .A(n11524), .B(n11521), .Z(n11523) );
  NAND2_X1 U11472 ( .A1(n11517), .A2(n11525), .ZN(n8132) );
  NAND2_X1 U11473 ( .A1(n11516), .A2(n11518), .ZN(n11525) );
  NAND2_X1 U11474 ( .A1(n11526), .A2(n11527), .ZN(n11518) );
  NAND2_X1 U11475 ( .A1(b_16_), .A2(a_0_), .ZN(n11527) );
  INV_X1 U11476 ( .A(n11528), .ZN(n11526) );
  XOR2_X1 U11477 ( .A(n11529), .B(n11530), .Z(n11516) );
  XOR2_X1 U11478 ( .A(n11531), .B(n11532), .Z(n11529) );
  NOR2_X1 U11479 ( .A1(n7872), .A2(n7669), .ZN(n11532) );
  NAND2_X1 U11480 ( .A1(a_0_), .A2(n11528), .ZN(n11517) );
  NAND2_X1 U11481 ( .A1(n11533), .A2(n11534), .ZN(n11528) );
  NAND3_X1 U11482 ( .A1(a_1_), .A2(n11535), .A3(b_16_), .ZN(n11534) );
  NAND2_X1 U11483 ( .A1(n11513), .A2(n11512), .ZN(n11535) );
  OR2_X1 U11484 ( .A1(n11512), .A2(n11513), .ZN(n11533) );
  AND2_X1 U11485 ( .A1(n11536), .A2(n11537), .ZN(n11513) );
  NAND2_X1 U11486 ( .A1(n11510), .A2(n11538), .ZN(n11537) );
  OR2_X1 U11487 ( .A1(n11508), .A2(n11509), .ZN(n11538) );
  NOR2_X1 U11488 ( .A1(n11233), .A2(n7966), .ZN(n11510) );
  NAND2_X1 U11489 ( .A1(n11508), .A2(n11509), .ZN(n11536) );
  NAND2_X1 U11490 ( .A1(n11539), .A2(n11540), .ZN(n11509) );
  NAND2_X1 U11491 ( .A1(n11506), .A2(n11541), .ZN(n11540) );
  OR2_X1 U11492 ( .A1(n11504), .A2(n11505), .ZN(n11541) );
  NOR2_X1 U11493 ( .A1(n11233), .A2(n7852), .ZN(n11506) );
  NAND2_X1 U11494 ( .A1(n11504), .A2(n11505), .ZN(n11539) );
  NAND2_X1 U11495 ( .A1(n11542), .A2(n11543), .ZN(n11505) );
  NAND2_X1 U11496 ( .A1(n11502), .A2(n11544), .ZN(n11543) );
  NAND2_X1 U11497 ( .A1(n11501), .A2(n11500), .ZN(n11544) );
  NOR2_X1 U11498 ( .A1(n11233), .A2(n7836), .ZN(n11502) );
  OR2_X1 U11499 ( .A1(n11500), .A2(n11501), .ZN(n11542) );
  AND2_X1 U11500 ( .A1(n11497), .A2(n11545), .ZN(n11501) );
  NAND2_X1 U11501 ( .A1(n11496), .A2(n11498), .ZN(n11545) );
  NAND2_X1 U11502 ( .A1(n11546), .A2(n11547), .ZN(n11498) );
  NAND2_X1 U11503 ( .A1(b_16_), .A2(a_5_), .ZN(n11547) );
  INV_X1 U11504 ( .A(n11548), .ZN(n11546) );
  XOR2_X1 U11505 ( .A(n11549), .B(n11550), .Z(n11496) );
  XOR2_X1 U11506 ( .A(n11551), .B(n11552), .Z(n11549) );
  NOR2_X1 U11507 ( .A1(n7807), .A2(n7669), .ZN(n11552) );
  NAND2_X1 U11508 ( .A1(a_5_), .A2(n11548), .ZN(n11497) );
  NAND2_X1 U11509 ( .A1(n11553), .A2(n11554), .ZN(n11548) );
  NAND3_X1 U11510 ( .A1(a_6_), .A2(n11555), .A3(b_16_), .ZN(n11554) );
  OR2_X1 U11511 ( .A1(n11493), .A2(n11491), .ZN(n11555) );
  NAND2_X1 U11512 ( .A1(n11491), .A2(n11493), .ZN(n11553) );
  NAND2_X1 U11513 ( .A1(n11556), .A2(n11557), .ZN(n11493) );
  NAND2_X1 U11514 ( .A1(n11490), .A2(n11558), .ZN(n11557) );
  OR2_X1 U11515 ( .A1(n11488), .A2(n11489), .ZN(n11558) );
  NOR2_X1 U11516 ( .A1(n11233), .A2(n7787), .ZN(n11490) );
  NAND2_X1 U11517 ( .A1(n11488), .A2(n11489), .ZN(n11556) );
  NAND2_X1 U11518 ( .A1(n11559), .A2(n11560), .ZN(n11489) );
  NAND3_X1 U11519 ( .A1(a_8_), .A2(n11561), .A3(b_16_), .ZN(n11560) );
  NAND2_X1 U11520 ( .A1(n11485), .A2(n11484), .ZN(n11561) );
  OR2_X1 U11521 ( .A1(n11484), .A2(n11485), .ZN(n11559) );
  AND2_X1 U11522 ( .A1(n11562), .A2(n11563), .ZN(n11485) );
  NAND2_X1 U11523 ( .A1(n11482), .A2(n11564), .ZN(n11563) );
  OR2_X1 U11524 ( .A1(n11481), .A2(n11479), .ZN(n11564) );
  NOR2_X1 U11525 ( .A1(n11233), .A2(n7753), .ZN(n11482) );
  NAND2_X1 U11526 ( .A1(n11479), .A2(n11481), .ZN(n11562) );
  NAND2_X1 U11527 ( .A1(n11565), .A2(n11566), .ZN(n11481) );
  NAND2_X1 U11528 ( .A1(n11478), .A2(n11567), .ZN(n11566) );
  OR2_X1 U11529 ( .A1(n11476), .A2(n11477), .ZN(n11567) );
  NOR2_X1 U11530 ( .A1(n11233), .A2(n8378), .ZN(n11478) );
  NAND2_X1 U11531 ( .A1(n11476), .A2(n11477), .ZN(n11565) );
  NAND2_X1 U11532 ( .A1(n11568), .A2(n11569), .ZN(n11477) );
  NAND2_X1 U11533 ( .A1(n11474), .A2(n11570), .ZN(n11569) );
  OR2_X1 U11534 ( .A1(n11472), .A2(n11473), .ZN(n11570) );
  NOR2_X1 U11535 ( .A1(n11233), .A2(n7724), .ZN(n11474) );
  NAND2_X1 U11536 ( .A1(n11472), .A2(n11473), .ZN(n11568) );
  NAND2_X1 U11537 ( .A1(n11571), .A2(n11572), .ZN(n11473) );
  NAND2_X1 U11538 ( .A1(n11470), .A2(n11573), .ZN(n11572) );
  NAND2_X1 U11539 ( .A1(n11469), .A2(n11468), .ZN(n11573) );
  NOR2_X1 U11540 ( .A1(n11233), .A2(n8585), .ZN(n11470) );
  OR2_X1 U11541 ( .A1(n11468), .A2(n11469), .ZN(n11571) );
  AND2_X1 U11542 ( .A1(n11574), .A2(n11575), .ZN(n11469) );
  NAND2_X1 U11543 ( .A1(n11466), .A2(n11576), .ZN(n11575) );
  NAND2_X1 U11544 ( .A1(n11465), .A2(n11464), .ZN(n11576) );
  NOR2_X1 U11545 ( .A1(n11233), .A2(n7702), .ZN(n11466) );
  OR2_X1 U11546 ( .A1(n11464), .A2(n11465), .ZN(n11574) );
  AND2_X1 U11547 ( .A1(n11577), .A2(n11578), .ZN(n11465) );
  NAND2_X1 U11548 ( .A1(n11462), .A2(n11579), .ZN(n11578) );
  OR2_X1 U11549 ( .A1(n11460), .A2(n11461), .ZN(n11579) );
  NOR2_X1 U11550 ( .A1(n11233), .A2(n7962), .ZN(n11462) );
  NAND2_X1 U11551 ( .A1(n11460), .A2(n11461), .ZN(n11577) );
  NAND2_X1 U11552 ( .A1(n11457), .A2(n11580), .ZN(n11461) );
  NAND2_X1 U11553 ( .A1(n11456), .A2(n11458), .ZN(n11580) );
  NAND2_X1 U11554 ( .A1(n11581), .A2(n11582), .ZN(n11458) );
  NAND2_X1 U11555 ( .A1(b_16_), .A2(a_15_), .ZN(n11582) );
  INV_X1 U11556 ( .A(n11583), .ZN(n11581) );
  XNOR2_X1 U11557 ( .A(n11584), .B(n11585), .ZN(n11456) );
  XOR2_X1 U11558 ( .A(n11586), .B(n11587), .Z(n11585) );
  NAND2_X1 U11559 ( .A1(b_15_), .A2(a_16_), .ZN(n11587) );
  NAND2_X1 U11560 ( .A1(a_15_), .A2(n11583), .ZN(n11457) );
  NAND2_X1 U11561 ( .A1(n11588), .A2(n11589), .ZN(n11583) );
  NAND2_X1 U11562 ( .A1(n11452), .A2(n11590), .ZN(n11589) );
  OR2_X1 U11563 ( .A1(n11454), .A2(n7652), .ZN(n11590) );
  XOR2_X1 U11564 ( .A(n11591), .B(n11592), .Z(n11452) );
  XOR2_X1 U11565 ( .A(n11593), .B(n11594), .Z(n11591) );
  NAND2_X1 U11566 ( .A1(n7652), .A2(n11454), .ZN(n11588) );
  NAND2_X1 U11567 ( .A1(n11595), .A2(n11596), .ZN(n11454) );
  NAND2_X1 U11568 ( .A1(n11451), .A2(n11597), .ZN(n11596) );
  OR2_X1 U11569 ( .A1(n11449), .A2(n11450), .ZN(n11597) );
  NOR2_X1 U11570 ( .A1(n11233), .A2(n7645), .ZN(n11451) );
  NAND2_X1 U11571 ( .A1(n11449), .A2(n11450), .ZN(n11595) );
  NAND2_X1 U11572 ( .A1(n11598), .A2(n11599), .ZN(n11450) );
  NAND3_X1 U11573 ( .A1(a_18_), .A2(n11600), .A3(b_16_), .ZN(n11599) );
  NAND2_X1 U11574 ( .A1(n11446), .A2(n11445), .ZN(n11600) );
  OR2_X1 U11575 ( .A1(n11445), .A2(n11446), .ZN(n11598) );
  AND2_X1 U11576 ( .A1(n11601), .A2(n11602), .ZN(n11446) );
  NAND2_X1 U11577 ( .A1(n11443), .A2(n11603), .ZN(n11602) );
  OR2_X1 U11578 ( .A1(n11440), .A2(n11442), .ZN(n11603) );
  NOR2_X1 U11579 ( .A1(n11233), .A2(n7958), .ZN(n11443) );
  NAND2_X1 U11580 ( .A1(n11440), .A2(n11442), .ZN(n11601) );
  NAND2_X1 U11581 ( .A1(n11604), .A2(n11605), .ZN(n11442) );
  NAND3_X1 U11582 ( .A1(a_20_), .A2(n11606), .A3(b_16_), .ZN(n11605) );
  NAND2_X1 U11583 ( .A1(n11438), .A2(n11437), .ZN(n11606) );
  OR2_X1 U11584 ( .A1(n11437), .A2(n11438), .ZN(n11604) );
  AND2_X1 U11585 ( .A1(n11607), .A2(n11608), .ZN(n11438) );
  NAND2_X1 U11586 ( .A1(n11435), .A2(n11609), .ZN(n11608) );
  OR2_X1 U11587 ( .A1(n11433), .A2(n11434), .ZN(n11609) );
  NOR2_X1 U11588 ( .A1(n11233), .A2(n7578), .ZN(n11435) );
  NAND2_X1 U11589 ( .A1(n11433), .A2(n11434), .ZN(n11607) );
  NAND2_X1 U11590 ( .A1(n11610), .A2(n11611), .ZN(n11434) );
  NAND3_X1 U11591 ( .A1(a_22_), .A2(n11612), .A3(b_16_), .ZN(n11611) );
  NAND2_X1 U11592 ( .A1(n11430), .A2(n11429), .ZN(n11612) );
  OR2_X1 U11593 ( .A1(n11429), .A2(n11430), .ZN(n11610) );
  AND2_X1 U11594 ( .A1(n11613), .A2(n11614), .ZN(n11430) );
  NAND2_X1 U11595 ( .A1(n11427), .A2(n11615), .ZN(n11614) );
  OR2_X1 U11596 ( .A1(n11424), .A2(n11426), .ZN(n11615) );
  NOR2_X1 U11597 ( .A1(n11233), .A2(n7955), .ZN(n11427) );
  NAND2_X1 U11598 ( .A1(n11424), .A2(n11426), .ZN(n11613) );
  NAND2_X1 U11599 ( .A1(n11616), .A2(n11617), .ZN(n11426) );
  NAND3_X1 U11600 ( .A1(a_24_), .A2(n11618), .A3(b_16_), .ZN(n11617) );
  NAND2_X1 U11601 ( .A1(n11422), .A2(n11421), .ZN(n11618) );
  OR2_X1 U11602 ( .A1(n11421), .A2(n11422), .ZN(n11616) );
  AND2_X1 U11603 ( .A1(n11619), .A2(n11620), .ZN(n11422) );
  NAND2_X1 U11604 ( .A1(n11419), .A2(n11621), .ZN(n11620) );
  OR2_X1 U11605 ( .A1(n11417), .A2(n11418), .ZN(n11621) );
  NOR2_X1 U11606 ( .A1(n11233), .A2(n7952), .ZN(n11419) );
  NAND2_X1 U11607 ( .A1(n11417), .A2(n11418), .ZN(n11619) );
  NAND2_X1 U11608 ( .A1(n11414), .A2(n11622), .ZN(n11418) );
  NAND2_X1 U11609 ( .A1(n11413), .A2(n11415), .ZN(n11622) );
  NAND2_X1 U11610 ( .A1(n11623), .A2(n11624), .ZN(n11415) );
  NAND2_X1 U11611 ( .A1(b_16_), .A2(a_26_), .ZN(n11624) );
  INV_X1 U11612 ( .A(n11625), .ZN(n11623) );
  XNOR2_X1 U11613 ( .A(n11626), .B(n11627), .ZN(n11413) );
  NAND2_X1 U11614 ( .A1(n11628), .A2(n11629), .ZN(n11626) );
  NAND2_X1 U11615 ( .A1(a_26_), .A2(n11625), .ZN(n11414) );
  NAND2_X1 U11616 ( .A1(n11386), .A2(n11630), .ZN(n11625) );
  NAND2_X1 U11617 ( .A1(n11385), .A2(n11387), .ZN(n11630) );
  NAND2_X1 U11618 ( .A1(n11631), .A2(n11632), .ZN(n11387) );
  NAND2_X1 U11619 ( .A1(b_16_), .A2(a_27_), .ZN(n11632) );
  INV_X1 U11620 ( .A(n11633), .ZN(n11631) );
  XNOR2_X1 U11621 ( .A(n11634), .B(n11635), .ZN(n11385) );
  XOR2_X1 U11622 ( .A(n11636), .B(n11637), .Z(n11634) );
  NAND2_X1 U11623 ( .A1(b_15_), .A2(a_28_), .ZN(n11636) );
  NAND2_X1 U11624 ( .A1(a_27_), .A2(n11633), .ZN(n11386) );
  NAND2_X1 U11625 ( .A1(n11638), .A2(n11639), .ZN(n11633) );
  NAND3_X1 U11626 ( .A1(a_28_), .A2(n11640), .A3(b_16_), .ZN(n11639) );
  NAND2_X1 U11627 ( .A1(n11395), .A2(n11393), .ZN(n11640) );
  OR2_X1 U11628 ( .A1(n11393), .A2(n11395), .ZN(n11638) );
  AND2_X1 U11629 ( .A1(n11641), .A2(n11642), .ZN(n11395) );
  NAND2_X1 U11630 ( .A1(n11409), .A2(n11643), .ZN(n11642) );
  OR2_X1 U11631 ( .A1(n11410), .A2(n11411), .ZN(n11643) );
  NOR2_X1 U11632 ( .A1(n11233), .A2(n7460), .ZN(n11409) );
  NAND2_X1 U11633 ( .A1(n11411), .A2(n11410), .ZN(n11641) );
  NAND2_X1 U11634 ( .A1(n11644), .A2(n11645), .ZN(n11410) );
  NAND2_X1 U11635 ( .A1(b_14_), .A2(n11646), .ZN(n11645) );
  NAND2_X1 U11636 ( .A1(n7441), .A2(n11647), .ZN(n11646) );
  NAND2_X1 U11637 ( .A1(a_31_), .A2(n7669), .ZN(n11647) );
  NAND2_X1 U11638 ( .A1(b_15_), .A2(n11648), .ZN(n11644) );
  NAND2_X1 U11639 ( .A1(n7445), .A2(n11649), .ZN(n11648) );
  NAND2_X1 U11640 ( .A1(a_30_), .A2(n7961), .ZN(n11649) );
  AND3_X1 U11641 ( .A1(b_16_), .A2(n7409), .A3(b_15_), .ZN(n11411) );
  XNOR2_X1 U11642 ( .A(n11650), .B(n11651), .ZN(n11393) );
  XOR2_X1 U11643 ( .A(n11652), .B(n11653), .Z(n11650) );
  XNOR2_X1 U11644 ( .A(n11654), .B(n11655), .ZN(n11417) );
  NAND2_X1 U11645 ( .A1(n11656), .A2(n11657), .ZN(n11654) );
  XNOR2_X1 U11646 ( .A(n11658), .B(n11659), .ZN(n11421) );
  XOR2_X1 U11647 ( .A(n11660), .B(n11661), .Z(n11658) );
  XNOR2_X1 U11648 ( .A(n11662), .B(n11663), .ZN(n11424) );
  XNOR2_X1 U11649 ( .A(n11664), .B(n11665), .ZN(n11662) );
  NOR2_X1 U11650 ( .A1(n7954), .A2(n7669), .ZN(n11665) );
  XOR2_X1 U11651 ( .A(n11666), .B(n11667), .Z(n11429) );
  XNOR2_X1 U11652 ( .A(n11668), .B(n11669), .ZN(n11667) );
  XNOR2_X1 U11653 ( .A(n11670), .B(n11671), .ZN(n11433) );
  XNOR2_X1 U11654 ( .A(n11672), .B(n11673), .ZN(n11670) );
  NOR2_X1 U11655 ( .A1(n7568), .A2(n7669), .ZN(n11673) );
  XNOR2_X1 U11656 ( .A(n11674), .B(n11675), .ZN(n11437) );
  XOR2_X1 U11657 ( .A(n11676), .B(n11677), .Z(n11674) );
  XNOR2_X1 U11658 ( .A(n11678), .B(n11679), .ZN(n11440) );
  XNOR2_X1 U11659 ( .A(n11680), .B(n11681), .ZN(n11678) );
  NOR2_X1 U11660 ( .A1(n7957), .A2(n7669), .ZN(n11681) );
  XOR2_X1 U11661 ( .A(n11682), .B(n11683), .Z(n11445) );
  XNOR2_X1 U11662 ( .A(n11684), .B(n11685), .ZN(n11683) );
  XNOR2_X1 U11663 ( .A(n11686), .B(n11687), .ZN(n11449) );
  XNOR2_X1 U11664 ( .A(n11688), .B(n11689), .ZN(n11686) );
  NOR2_X1 U11665 ( .A1(n7960), .A2(n7669), .ZN(n11689) );
  NOR2_X1 U11666 ( .A1(n11233), .A2(n8353), .ZN(n7652) );
  INV_X1 U11667 ( .A(b_16_), .ZN(n11233) );
  XNOR2_X1 U11668 ( .A(n11690), .B(n11691), .ZN(n11460) );
  XOR2_X1 U11669 ( .A(n7915), .B(n11692), .Z(n11691) );
  XOR2_X1 U11670 ( .A(n11693), .B(n11694), .Z(n11464) );
  NAND2_X1 U11671 ( .A1(n11695), .A2(n11696), .ZN(n11693) );
  XOR2_X1 U11672 ( .A(n11697), .B(n11698), .Z(n11468) );
  XOR2_X1 U11673 ( .A(n11699), .B(n11700), .Z(n11698) );
  NAND2_X1 U11674 ( .A1(b_15_), .A2(a_13_), .ZN(n11700) );
  XNOR2_X1 U11675 ( .A(n11701), .B(n11702), .ZN(n11472) );
  XOR2_X1 U11676 ( .A(n11703), .B(n11704), .Z(n11702) );
  NAND2_X1 U11677 ( .A1(b_15_), .A2(a_12_), .ZN(n11704) );
  XNOR2_X1 U11678 ( .A(n11705), .B(n11706), .ZN(n11476) );
  XNOR2_X1 U11679 ( .A(n11707), .B(n11708), .ZN(n11705) );
  NOR2_X1 U11680 ( .A1(n7724), .A2(n7669), .ZN(n11708) );
  XNOR2_X1 U11681 ( .A(n11709), .B(n11710), .ZN(n11479) );
  XOR2_X1 U11682 ( .A(n11711), .B(n11712), .Z(n11710) );
  NAND2_X1 U11683 ( .A1(b_15_), .A2(a_10_), .ZN(n11712) );
  XOR2_X1 U11684 ( .A(n11713), .B(n11714), .Z(n11484) );
  XOR2_X1 U11685 ( .A(n11715), .B(n11716), .Z(n11714) );
  NAND2_X1 U11686 ( .A1(b_15_), .A2(a_9_), .ZN(n11716) );
  XNOR2_X1 U11687 ( .A(n11717), .B(n11718), .ZN(n11488) );
  XNOR2_X1 U11688 ( .A(n11719), .B(n11720), .ZN(n11717) );
  NOR2_X1 U11689 ( .A1(n8602), .A2(n7669), .ZN(n11720) );
  XOR2_X1 U11690 ( .A(n11721), .B(n11722), .Z(n11491) );
  XOR2_X1 U11691 ( .A(n11723), .B(n11724), .Z(n11721) );
  NOR2_X1 U11692 ( .A1(n7787), .A2(n7669), .ZN(n11724) );
  XNOR2_X1 U11693 ( .A(n11725), .B(n11726), .ZN(n11500) );
  XNOR2_X1 U11694 ( .A(n11727), .B(n11728), .ZN(n11725) );
  NAND2_X1 U11695 ( .A1(b_15_), .A2(a_5_), .ZN(n11727) );
  XNOR2_X1 U11696 ( .A(n11729), .B(n11730), .ZN(n11504) );
  XNOR2_X1 U11697 ( .A(n11731), .B(n11732), .ZN(n11729) );
  NOR2_X1 U11698 ( .A1(n7836), .A2(n7669), .ZN(n11732) );
  XNOR2_X1 U11699 ( .A(n11733), .B(n11734), .ZN(n11508) );
  XOR2_X1 U11700 ( .A(n11735), .B(n11736), .Z(n11734) );
  NAND2_X1 U11701 ( .A1(b_15_), .A2(a_3_), .ZN(n11736) );
  XOR2_X1 U11702 ( .A(n11737), .B(n11738), .Z(n11512) );
  XOR2_X1 U11703 ( .A(n11739), .B(n11740), .Z(n11738) );
  NAND2_X1 U11704 ( .A1(b_15_), .A2(a_2_), .ZN(n11740) );
  XNOR2_X1 U11705 ( .A(n11741), .B(n11742), .ZN(n8133) );
  XOR2_X1 U11706 ( .A(n11743), .B(n11744), .Z(n11742) );
  NAND2_X1 U11707 ( .A1(b_15_), .A2(a_0_), .ZN(n11744) );
  NAND2_X1 U11708 ( .A1(n11745), .A2(n11746), .ZN(n8067) );
  NAND2_X1 U11709 ( .A1(n11524), .A2(n11521), .ZN(n11746) );
  XNOR2_X1 U11710 ( .A(n8123), .B(n8124), .ZN(n11745) );
  NAND3_X1 U11711 ( .A1(n11524), .A2(n11521), .A3(n11747), .ZN(n8066) );
  XOR2_X1 U11712 ( .A(n8124), .B(n8123), .Z(n11747) );
  NAND2_X1 U11713 ( .A1(n11748), .A2(n11749), .ZN(n11521) );
  NAND3_X1 U11714 ( .A1(a_0_), .A2(n11750), .A3(b_15_), .ZN(n11749) );
  OR2_X1 U11715 ( .A1(n11743), .A2(n11741), .ZN(n11750) );
  NAND2_X1 U11716 ( .A1(n11741), .A2(n11743), .ZN(n11748) );
  NAND2_X1 U11717 ( .A1(n11751), .A2(n11752), .ZN(n11743) );
  NAND3_X1 U11718 ( .A1(a_1_), .A2(n11753), .A3(b_15_), .ZN(n11752) );
  OR2_X1 U11719 ( .A1(n11530), .A2(n11531), .ZN(n11753) );
  NAND2_X1 U11720 ( .A1(n11530), .A2(n11531), .ZN(n11751) );
  NAND2_X1 U11721 ( .A1(n11754), .A2(n11755), .ZN(n11531) );
  NAND3_X1 U11722 ( .A1(a_2_), .A2(n11756), .A3(b_15_), .ZN(n11755) );
  OR2_X1 U11723 ( .A1(n11737), .A2(n11739), .ZN(n11756) );
  NAND2_X1 U11724 ( .A1(n11737), .A2(n11739), .ZN(n11754) );
  NAND2_X1 U11725 ( .A1(n11757), .A2(n11758), .ZN(n11739) );
  NAND3_X1 U11726 ( .A1(a_3_), .A2(n11759), .A3(b_15_), .ZN(n11758) );
  OR2_X1 U11727 ( .A1(n11735), .A2(n11733), .ZN(n11759) );
  NAND2_X1 U11728 ( .A1(n11733), .A2(n11735), .ZN(n11757) );
  NAND2_X1 U11729 ( .A1(n11760), .A2(n11761), .ZN(n11735) );
  NAND3_X1 U11730 ( .A1(a_4_), .A2(n11762), .A3(b_15_), .ZN(n11761) );
  NAND2_X1 U11731 ( .A1(n11731), .A2(n11730), .ZN(n11762) );
  OR2_X1 U11732 ( .A1(n11730), .A2(n11731), .ZN(n11760) );
  AND2_X1 U11733 ( .A1(n11763), .A2(n11764), .ZN(n11731) );
  NAND3_X1 U11734 ( .A1(a_5_), .A2(n11765), .A3(b_15_), .ZN(n11764) );
  OR2_X1 U11735 ( .A1(n11726), .A2(n11728), .ZN(n11765) );
  NAND2_X1 U11736 ( .A1(n11726), .A2(n11728), .ZN(n11763) );
  NAND2_X1 U11737 ( .A1(n11766), .A2(n11767), .ZN(n11728) );
  NAND3_X1 U11738 ( .A1(a_6_), .A2(n11768), .A3(b_15_), .ZN(n11767) );
  OR2_X1 U11739 ( .A1(n11550), .A2(n11551), .ZN(n11768) );
  NAND2_X1 U11740 ( .A1(n11550), .A2(n11551), .ZN(n11766) );
  NAND2_X1 U11741 ( .A1(n11769), .A2(n11770), .ZN(n11551) );
  NAND3_X1 U11742 ( .A1(a_7_), .A2(n11771), .A3(b_15_), .ZN(n11770) );
  OR2_X1 U11743 ( .A1(n11722), .A2(n11723), .ZN(n11771) );
  NAND2_X1 U11744 ( .A1(n11722), .A2(n11723), .ZN(n11769) );
  NAND2_X1 U11745 ( .A1(n11772), .A2(n11773), .ZN(n11723) );
  NAND3_X1 U11746 ( .A1(a_8_), .A2(n11774), .A3(b_15_), .ZN(n11773) );
  NAND2_X1 U11747 ( .A1(n11719), .A2(n11718), .ZN(n11774) );
  OR2_X1 U11748 ( .A1(n11718), .A2(n11719), .ZN(n11772) );
  AND2_X1 U11749 ( .A1(n11775), .A2(n11776), .ZN(n11719) );
  NAND3_X1 U11750 ( .A1(a_9_), .A2(n11777), .A3(b_15_), .ZN(n11776) );
  OR2_X1 U11751 ( .A1(n11713), .A2(n11715), .ZN(n11777) );
  NAND2_X1 U11752 ( .A1(n11713), .A2(n11715), .ZN(n11775) );
  NAND2_X1 U11753 ( .A1(n11778), .A2(n11779), .ZN(n11715) );
  NAND3_X1 U11754 ( .A1(a_10_), .A2(n11780), .A3(b_15_), .ZN(n11779) );
  OR2_X1 U11755 ( .A1(n11709), .A2(n11711), .ZN(n11780) );
  NAND2_X1 U11756 ( .A1(n11709), .A2(n11711), .ZN(n11778) );
  NAND2_X1 U11757 ( .A1(n11781), .A2(n11782), .ZN(n11711) );
  NAND3_X1 U11758 ( .A1(a_11_), .A2(n11783), .A3(b_15_), .ZN(n11782) );
  NAND2_X1 U11759 ( .A1(n11707), .A2(n11706), .ZN(n11783) );
  OR2_X1 U11760 ( .A1(n11706), .A2(n11707), .ZN(n11781) );
  AND2_X1 U11761 ( .A1(n11784), .A2(n11785), .ZN(n11707) );
  NAND3_X1 U11762 ( .A1(a_12_), .A2(n11786), .A3(b_15_), .ZN(n11785) );
  OR2_X1 U11763 ( .A1(n11703), .A2(n11701), .ZN(n11786) );
  NAND2_X1 U11764 ( .A1(n11701), .A2(n11703), .ZN(n11784) );
  NAND2_X1 U11765 ( .A1(n11787), .A2(n11788), .ZN(n11703) );
  NAND3_X1 U11766 ( .A1(a_13_), .A2(n11789), .A3(b_15_), .ZN(n11788) );
  OR2_X1 U11767 ( .A1(n11697), .A2(n11699), .ZN(n11789) );
  NAND2_X1 U11768 ( .A1(n11697), .A2(n11699), .ZN(n11787) );
  NAND2_X1 U11769 ( .A1(n11695), .A2(n11790), .ZN(n11699) );
  NAND2_X1 U11770 ( .A1(n11694), .A2(n11696), .ZN(n11790) );
  NAND2_X1 U11771 ( .A1(n11791), .A2(n11792), .ZN(n11696) );
  NAND2_X1 U11772 ( .A1(b_15_), .A2(a_14_), .ZN(n11792) );
  INV_X1 U11773 ( .A(n11793), .ZN(n11791) );
  XOR2_X1 U11774 ( .A(n11794), .B(n11795), .Z(n11694) );
  XOR2_X1 U11775 ( .A(n11796), .B(n11797), .Z(n11794) );
  NAND2_X1 U11776 ( .A1(a_14_), .A2(n11793), .ZN(n11695) );
  NAND2_X1 U11777 ( .A1(n11798), .A2(n11799), .ZN(n11793) );
  NAND2_X1 U11778 ( .A1(n11690), .A2(n11800), .ZN(n11799) );
  OR2_X1 U11779 ( .A1(n11692), .A2(n7664), .ZN(n11800) );
  XNOR2_X1 U11780 ( .A(n11801), .B(n11802), .ZN(n11690) );
  XNOR2_X1 U11781 ( .A(n11803), .B(n11804), .ZN(n11802) );
  NAND2_X1 U11782 ( .A1(n7664), .A2(n11692), .ZN(n11798) );
  NAND2_X1 U11783 ( .A1(n11805), .A2(n11806), .ZN(n11692) );
  NAND3_X1 U11784 ( .A1(a_16_), .A2(n11807), .A3(b_15_), .ZN(n11806) );
  OR2_X1 U11785 ( .A1(n11586), .A2(n11584), .ZN(n11807) );
  NAND2_X1 U11786 ( .A1(n11584), .A2(n11586), .ZN(n11805) );
  NAND2_X1 U11787 ( .A1(n11808), .A2(n11809), .ZN(n11586) );
  NAND2_X1 U11788 ( .A1(n11594), .A2(n11810), .ZN(n11809) );
  OR2_X1 U11789 ( .A1(n11592), .A2(n11593), .ZN(n11810) );
  NOR2_X1 U11790 ( .A1(n7669), .A2(n7645), .ZN(n11594) );
  NAND2_X1 U11791 ( .A1(n11592), .A2(n11593), .ZN(n11808) );
  NAND2_X1 U11792 ( .A1(n11811), .A2(n11812), .ZN(n11593) );
  NAND3_X1 U11793 ( .A1(a_18_), .A2(n11813), .A3(b_15_), .ZN(n11812) );
  NAND2_X1 U11794 ( .A1(n11688), .A2(n11687), .ZN(n11813) );
  OR2_X1 U11795 ( .A1(n11687), .A2(n11688), .ZN(n11811) );
  AND2_X1 U11796 ( .A1(n11814), .A2(n11815), .ZN(n11688) );
  NAND2_X1 U11797 ( .A1(n11685), .A2(n11816), .ZN(n11815) );
  OR2_X1 U11798 ( .A1(n11682), .A2(n11684), .ZN(n11816) );
  NOR2_X1 U11799 ( .A1(n7669), .A2(n7958), .ZN(n11685) );
  NAND2_X1 U11800 ( .A1(n11682), .A2(n11684), .ZN(n11814) );
  NAND2_X1 U11801 ( .A1(n11817), .A2(n11818), .ZN(n11684) );
  NAND3_X1 U11802 ( .A1(a_20_), .A2(n11819), .A3(b_15_), .ZN(n11818) );
  NAND2_X1 U11803 ( .A1(n11680), .A2(n11679), .ZN(n11819) );
  OR2_X1 U11804 ( .A1(n11679), .A2(n11680), .ZN(n11817) );
  AND2_X1 U11805 ( .A1(n11820), .A2(n11821), .ZN(n11680) );
  NAND2_X1 U11806 ( .A1(n11677), .A2(n11822), .ZN(n11821) );
  OR2_X1 U11807 ( .A1(n11675), .A2(n11676), .ZN(n11822) );
  NOR2_X1 U11808 ( .A1(n7669), .A2(n7578), .ZN(n11677) );
  NAND2_X1 U11809 ( .A1(n11675), .A2(n11676), .ZN(n11820) );
  NAND2_X1 U11810 ( .A1(n11823), .A2(n11824), .ZN(n11676) );
  NAND3_X1 U11811 ( .A1(a_22_), .A2(n11825), .A3(b_15_), .ZN(n11824) );
  NAND2_X1 U11812 ( .A1(n11672), .A2(n11671), .ZN(n11825) );
  OR2_X1 U11813 ( .A1(n11671), .A2(n11672), .ZN(n11823) );
  AND2_X1 U11814 ( .A1(n11826), .A2(n11827), .ZN(n11672) );
  NAND2_X1 U11815 ( .A1(n11669), .A2(n11828), .ZN(n11827) );
  OR2_X1 U11816 ( .A1(n11666), .A2(n11668), .ZN(n11828) );
  NOR2_X1 U11817 ( .A1(n7669), .A2(n7955), .ZN(n11669) );
  NAND2_X1 U11818 ( .A1(n11666), .A2(n11668), .ZN(n11826) );
  NAND2_X1 U11819 ( .A1(n11829), .A2(n11830), .ZN(n11668) );
  NAND3_X1 U11820 ( .A1(a_24_), .A2(n11831), .A3(b_15_), .ZN(n11830) );
  NAND2_X1 U11821 ( .A1(n11664), .A2(n11663), .ZN(n11831) );
  OR2_X1 U11822 ( .A1(n11663), .A2(n11664), .ZN(n11829) );
  AND2_X1 U11823 ( .A1(n11832), .A2(n11833), .ZN(n11664) );
  NAND2_X1 U11824 ( .A1(n11661), .A2(n11834), .ZN(n11833) );
  OR2_X1 U11825 ( .A1(n11659), .A2(n11660), .ZN(n11834) );
  NOR2_X1 U11826 ( .A1(n7669), .A2(n7952), .ZN(n11661) );
  NAND2_X1 U11827 ( .A1(n11659), .A2(n11660), .ZN(n11832) );
  NAND2_X1 U11828 ( .A1(n11656), .A2(n11835), .ZN(n11660) );
  NAND2_X1 U11829 ( .A1(n11655), .A2(n11657), .ZN(n11835) );
  NAND2_X1 U11830 ( .A1(n11836), .A2(n11837), .ZN(n11657) );
  NAND2_X1 U11831 ( .A1(b_15_), .A2(a_26_), .ZN(n11837) );
  INV_X1 U11832 ( .A(n11838), .ZN(n11836) );
  XNOR2_X1 U11833 ( .A(n11839), .B(n11840), .ZN(n11655) );
  NAND2_X1 U11834 ( .A1(n11841), .A2(n11842), .ZN(n11839) );
  NAND2_X1 U11835 ( .A1(a_26_), .A2(n11838), .ZN(n11656) );
  NAND2_X1 U11836 ( .A1(n11628), .A2(n11843), .ZN(n11838) );
  NAND2_X1 U11837 ( .A1(n11627), .A2(n11629), .ZN(n11843) );
  NAND2_X1 U11838 ( .A1(n11844), .A2(n11845), .ZN(n11629) );
  NAND2_X1 U11839 ( .A1(b_15_), .A2(a_27_), .ZN(n11845) );
  INV_X1 U11840 ( .A(n11846), .ZN(n11844) );
  XNOR2_X1 U11841 ( .A(n11847), .B(n11848), .ZN(n11627) );
  XOR2_X1 U11842 ( .A(n11849), .B(n11850), .Z(n11847) );
  NAND2_X1 U11843 ( .A1(b_14_), .A2(a_28_), .ZN(n11849) );
  NAND2_X1 U11844 ( .A1(a_27_), .A2(n11846), .ZN(n11628) );
  NAND2_X1 U11845 ( .A1(n11851), .A2(n11852), .ZN(n11846) );
  NAND3_X1 U11846 ( .A1(a_28_), .A2(n11853), .A3(b_15_), .ZN(n11852) );
  NAND2_X1 U11847 ( .A1(n11637), .A2(n11635), .ZN(n11853) );
  OR2_X1 U11848 ( .A1(n11635), .A2(n11637), .ZN(n11851) );
  AND2_X1 U11849 ( .A1(n11854), .A2(n11855), .ZN(n11637) );
  NAND2_X1 U11850 ( .A1(n11651), .A2(n11856), .ZN(n11855) );
  OR2_X1 U11851 ( .A1(n11652), .A2(n11653), .ZN(n11856) );
  NOR2_X1 U11852 ( .A1(n7669), .A2(n7460), .ZN(n11651) );
  INV_X1 U11853 ( .A(b_15_), .ZN(n7669) );
  NAND2_X1 U11854 ( .A1(n11653), .A2(n11652), .ZN(n11854) );
  NAND2_X1 U11855 ( .A1(n11857), .A2(n11858), .ZN(n11652) );
  NAND2_X1 U11856 ( .A1(b_13_), .A2(n11859), .ZN(n11858) );
  NAND2_X1 U11857 ( .A1(n7441), .A2(n11860), .ZN(n11859) );
  NAND2_X1 U11858 ( .A1(a_31_), .A2(n7961), .ZN(n11860) );
  NAND2_X1 U11859 ( .A1(b_14_), .A2(n11861), .ZN(n11857) );
  NAND2_X1 U11860 ( .A1(n7445), .A2(n11862), .ZN(n11861) );
  NAND2_X1 U11861 ( .A1(a_30_), .A2(n7695), .ZN(n11862) );
  AND3_X1 U11862 ( .A1(b_14_), .A2(n7409), .A3(b_15_), .ZN(n11653) );
  XNOR2_X1 U11863 ( .A(n11863), .B(n11864), .ZN(n11635) );
  XOR2_X1 U11864 ( .A(n11865), .B(n11866), .Z(n11863) );
  XNOR2_X1 U11865 ( .A(n11867), .B(n11868), .ZN(n11659) );
  NAND2_X1 U11866 ( .A1(n11869), .A2(n11870), .ZN(n11867) );
  XNOR2_X1 U11867 ( .A(n11871), .B(n11872), .ZN(n11663) );
  XOR2_X1 U11868 ( .A(n11873), .B(n11874), .Z(n11871) );
  XNOR2_X1 U11869 ( .A(n11875), .B(n11876), .ZN(n11666) );
  XNOR2_X1 U11870 ( .A(n11877), .B(n11878), .ZN(n11875) );
  NOR2_X1 U11871 ( .A1(n7954), .A2(n7961), .ZN(n11878) );
  XOR2_X1 U11872 ( .A(n11879), .B(n11880), .Z(n11671) );
  XNOR2_X1 U11873 ( .A(n11881), .B(n11882), .ZN(n11880) );
  XNOR2_X1 U11874 ( .A(n11883), .B(n11884), .ZN(n11675) );
  XOR2_X1 U11875 ( .A(n11885), .B(n11886), .Z(n11884) );
  NAND2_X1 U11876 ( .A1(b_14_), .A2(a_22_), .ZN(n11886) );
  XNOR2_X1 U11877 ( .A(n11887), .B(n11888), .ZN(n11679) );
  XOR2_X1 U11878 ( .A(n11889), .B(n11890), .Z(n11887) );
  XNOR2_X1 U11879 ( .A(n11891), .B(n11892), .ZN(n11682) );
  XNOR2_X1 U11880 ( .A(n11893), .B(n11894), .ZN(n11891) );
  NOR2_X1 U11881 ( .A1(n7957), .A2(n7961), .ZN(n11894) );
  XOR2_X1 U11882 ( .A(n11895), .B(n11896), .Z(n11687) );
  XNOR2_X1 U11883 ( .A(n11897), .B(n11898), .ZN(n11896) );
  XNOR2_X1 U11884 ( .A(n11899), .B(n11900), .ZN(n11592) );
  XNOR2_X1 U11885 ( .A(n11901), .B(n11902), .ZN(n11899) );
  NOR2_X1 U11886 ( .A1(n7960), .A2(n7961), .ZN(n11902) );
  XOR2_X1 U11887 ( .A(n11903), .B(n11904), .Z(n11584) );
  XOR2_X1 U11888 ( .A(n11905), .B(n11906), .Z(n11903) );
  NOR2_X1 U11889 ( .A1(n7645), .A2(n7961), .ZN(n11906) );
  INV_X1 U11890 ( .A(n7915), .ZN(n7664) );
  NAND2_X1 U11891 ( .A1(b_15_), .A2(a_15_), .ZN(n7915) );
  XOR2_X1 U11892 ( .A(n11907), .B(n11908), .Z(n11697) );
  XOR2_X1 U11893 ( .A(n11909), .B(n11910), .Z(n11907) );
  XNOR2_X1 U11894 ( .A(n11911), .B(n11912), .ZN(n11701) );
  NAND2_X1 U11895 ( .A1(n11913), .A2(n11914), .ZN(n11911) );
  XNOR2_X1 U11896 ( .A(n11915), .B(n11916), .ZN(n11706) );
  XOR2_X1 U11897 ( .A(n11917), .B(n11918), .Z(n11915) );
  XNOR2_X1 U11898 ( .A(n11919), .B(n11920), .ZN(n11709) );
  XNOR2_X1 U11899 ( .A(n11921), .B(n11922), .ZN(n11919) );
  NOR2_X1 U11900 ( .A1(n7724), .A2(n7961), .ZN(n11922) );
  XNOR2_X1 U11901 ( .A(n11923), .B(n11924), .ZN(n11713) );
  XNOR2_X1 U11902 ( .A(n11925), .B(n11926), .ZN(n11923) );
  XOR2_X1 U11903 ( .A(n11927), .B(n11928), .Z(n11718) );
  XOR2_X1 U11904 ( .A(n11929), .B(n11930), .Z(n11928) );
  NAND2_X1 U11905 ( .A1(b_14_), .A2(a_9_), .ZN(n11930) );
  XNOR2_X1 U11906 ( .A(n11931), .B(n11932), .ZN(n11722) );
  NAND2_X1 U11907 ( .A1(n11933), .A2(n11934), .ZN(n11931) );
  XNOR2_X1 U11908 ( .A(n11935), .B(n11936), .ZN(n11550) );
  NAND2_X1 U11909 ( .A1(n11937), .A2(n11938), .ZN(n11935) );
  XNOR2_X1 U11910 ( .A(n11939), .B(n11940), .ZN(n11726) );
  NAND2_X1 U11911 ( .A1(n11941), .A2(n11942), .ZN(n11939) );
  XOR2_X1 U11912 ( .A(n11943), .B(n11944), .Z(n11730) );
  NAND2_X1 U11913 ( .A1(n11945), .A2(n11946), .ZN(n11943) );
  XNOR2_X1 U11914 ( .A(n11947), .B(n11948), .ZN(n11733) );
  XNOR2_X1 U11915 ( .A(n11949), .B(n11950), .ZN(n11948) );
  XNOR2_X1 U11916 ( .A(n11951), .B(n11952), .ZN(n11737) );
  XNOR2_X1 U11917 ( .A(n11953), .B(n11954), .ZN(n11952) );
  XNOR2_X1 U11918 ( .A(n11955), .B(n11956), .ZN(n11530) );
  XNOR2_X1 U11919 ( .A(n11957), .B(n11958), .ZN(n11955) );
  NOR2_X1 U11920 ( .A1(n7966), .A2(n7961), .ZN(n11958) );
  XNOR2_X1 U11921 ( .A(n11959), .B(n11960), .ZN(n11741) );
  XNOR2_X1 U11922 ( .A(n11961), .B(n11962), .ZN(n11960) );
  INV_X1 U11923 ( .A(n11522), .ZN(n11524) );
  XOR2_X1 U11924 ( .A(n11963), .B(n11964), .Z(n11522) );
  XOR2_X1 U11925 ( .A(n11965), .B(n11966), .Z(n11964) );
  NAND2_X1 U11926 ( .A1(b_14_), .A2(a_0_), .ZN(n11966) );
  NAND4_X1 U11927 ( .A1(n8123), .A2(n8122), .A3(n8124), .A4(n8118), .ZN(n8071)
         );
  INV_X1 U11928 ( .A(n11967), .ZN(n8118) );
  NAND2_X1 U11929 ( .A1(n11968), .A2(n11969), .ZN(n8124) );
  NAND3_X1 U11930 ( .A1(a_0_), .A2(n11970), .A3(b_14_), .ZN(n11969) );
  OR2_X1 U11931 ( .A1(n11965), .A2(n11963), .ZN(n11970) );
  NAND2_X1 U11932 ( .A1(n11963), .A2(n11965), .ZN(n11968) );
  NAND2_X1 U11933 ( .A1(n11971), .A2(n11972), .ZN(n11965) );
  NAND2_X1 U11934 ( .A1(n11962), .A2(n11973), .ZN(n11972) );
  OR2_X1 U11935 ( .A1(n11961), .A2(n11959), .ZN(n11973) );
  NOR2_X1 U11936 ( .A1(n7961), .A2(n7872), .ZN(n11962) );
  NAND2_X1 U11937 ( .A1(n11959), .A2(n11961), .ZN(n11971) );
  NAND2_X1 U11938 ( .A1(n11974), .A2(n11975), .ZN(n11961) );
  NAND3_X1 U11939 ( .A1(a_2_), .A2(n11976), .A3(b_14_), .ZN(n11975) );
  NAND2_X1 U11940 ( .A1(n11957), .A2(n11956), .ZN(n11976) );
  OR2_X1 U11941 ( .A1(n11956), .A2(n11957), .ZN(n11974) );
  AND2_X1 U11942 ( .A1(n11977), .A2(n11978), .ZN(n11957) );
  NAND2_X1 U11943 ( .A1(n11954), .A2(n11979), .ZN(n11978) );
  OR2_X1 U11944 ( .A1(n11953), .A2(n11951), .ZN(n11979) );
  NOR2_X1 U11945 ( .A1(n7961), .A2(n7852), .ZN(n11954) );
  NAND2_X1 U11946 ( .A1(n11951), .A2(n11953), .ZN(n11977) );
  NAND2_X1 U11947 ( .A1(n11980), .A2(n11981), .ZN(n11953) );
  NAND2_X1 U11948 ( .A1(n11950), .A2(n11982), .ZN(n11981) );
  OR2_X1 U11949 ( .A1(n11949), .A2(n11947), .ZN(n11982) );
  NOR2_X1 U11950 ( .A1(n7961), .A2(n7836), .ZN(n11950) );
  NAND2_X1 U11951 ( .A1(n11947), .A2(n11949), .ZN(n11980) );
  NAND2_X1 U11952 ( .A1(n11945), .A2(n11983), .ZN(n11949) );
  NAND2_X1 U11953 ( .A1(n11944), .A2(n11946), .ZN(n11983) );
  NAND2_X1 U11954 ( .A1(n11984), .A2(n11985), .ZN(n11946) );
  NAND2_X1 U11955 ( .A1(b_14_), .A2(a_5_), .ZN(n11985) );
  INV_X1 U11956 ( .A(n11986), .ZN(n11984) );
  XNOR2_X1 U11957 ( .A(n11987), .B(n11988), .ZN(n11944) );
  XOR2_X1 U11958 ( .A(n11989), .B(n11990), .Z(n11988) );
  NAND2_X1 U11959 ( .A1(b_13_), .A2(a_6_), .ZN(n11990) );
  NAND2_X1 U11960 ( .A1(a_5_), .A2(n11986), .ZN(n11945) );
  NAND2_X1 U11961 ( .A1(n11941), .A2(n11991), .ZN(n11986) );
  NAND2_X1 U11962 ( .A1(n11940), .A2(n11942), .ZN(n11991) );
  NAND2_X1 U11963 ( .A1(n11992), .A2(n11993), .ZN(n11942) );
  NAND2_X1 U11964 ( .A1(b_14_), .A2(a_6_), .ZN(n11993) );
  INV_X1 U11965 ( .A(n11994), .ZN(n11992) );
  XNOR2_X1 U11966 ( .A(n11995), .B(n11996), .ZN(n11940) );
  XOR2_X1 U11967 ( .A(n11997), .B(n11998), .Z(n11996) );
  NAND2_X1 U11968 ( .A1(b_13_), .A2(a_7_), .ZN(n11998) );
  NAND2_X1 U11969 ( .A1(a_6_), .A2(n11994), .ZN(n11941) );
  NAND2_X1 U11970 ( .A1(n11937), .A2(n11999), .ZN(n11994) );
  NAND2_X1 U11971 ( .A1(n11936), .A2(n11938), .ZN(n11999) );
  NAND2_X1 U11972 ( .A1(n12000), .A2(n12001), .ZN(n11938) );
  NAND2_X1 U11973 ( .A1(b_14_), .A2(a_7_), .ZN(n12001) );
  INV_X1 U11974 ( .A(n12002), .ZN(n12000) );
  XNOR2_X1 U11975 ( .A(n12003), .B(n12004), .ZN(n11936) );
  XNOR2_X1 U11976 ( .A(n12005), .B(n12006), .ZN(n12003) );
  NOR2_X1 U11977 ( .A1(n8602), .A2(n7695), .ZN(n12006) );
  NAND2_X1 U11978 ( .A1(a_7_), .A2(n12002), .ZN(n11937) );
  NAND2_X1 U11979 ( .A1(n11933), .A2(n12007), .ZN(n12002) );
  NAND2_X1 U11980 ( .A1(n11932), .A2(n11934), .ZN(n12007) );
  NAND2_X1 U11981 ( .A1(n12008), .A2(n12009), .ZN(n11934) );
  NAND2_X1 U11982 ( .A1(b_14_), .A2(a_8_), .ZN(n12009) );
  INV_X1 U11983 ( .A(n12010), .ZN(n12008) );
  XNOR2_X1 U11984 ( .A(n12011), .B(n12012), .ZN(n11932) );
  XOR2_X1 U11985 ( .A(n12013), .B(n12014), .Z(n12012) );
  NAND2_X1 U11986 ( .A1(b_13_), .A2(a_9_), .ZN(n12014) );
  NAND2_X1 U11987 ( .A1(a_8_), .A2(n12010), .ZN(n11933) );
  NAND2_X1 U11988 ( .A1(n12015), .A2(n12016), .ZN(n12010) );
  NAND3_X1 U11989 ( .A1(a_9_), .A2(n12017), .A3(b_14_), .ZN(n12016) );
  OR2_X1 U11990 ( .A1(n11929), .A2(n11927), .ZN(n12017) );
  NAND2_X1 U11991 ( .A1(n11927), .A2(n11929), .ZN(n12015) );
  NAND2_X1 U11992 ( .A1(n12018), .A2(n12019), .ZN(n11929) );
  NAND2_X1 U11993 ( .A1(n11926), .A2(n12020), .ZN(n12019) );
  NAND2_X1 U11994 ( .A1(n11925), .A2(n11924), .ZN(n12020) );
  NOR2_X1 U11995 ( .A1(n7961), .A2(n8378), .ZN(n11926) );
  OR2_X1 U11996 ( .A1(n11924), .A2(n11925), .ZN(n12018) );
  AND2_X1 U11997 ( .A1(n12021), .A2(n12022), .ZN(n11925) );
  NAND3_X1 U11998 ( .A1(a_11_), .A2(n12023), .A3(b_14_), .ZN(n12022) );
  NAND2_X1 U11999 ( .A1(n11921), .A2(n11920), .ZN(n12023) );
  OR2_X1 U12000 ( .A1(n11920), .A2(n11921), .ZN(n12021) );
  AND2_X1 U12001 ( .A1(n12024), .A2(n12025), .ZN(n11921) );
  NAND2_X1 U12002 ( .A1(n11918), .A2(n12026), .ZN(n12025) );
  OR2_X1 U12003 ( .A1(n11917), .A2(n11916), .ZN(n12026) );
  NOR2_X1 U12004 ( .A1(n7961), .A2(n8585), .ZN(n11918) );
  NAND2_X1 U12005 ( .A1(n11916), .A2(n11917), .ZN(n12024) );
  NAND2_X1 U12006 ( .A1(n11913), .A2(n12027), .ZN(n11917) );
  NAND2_X1 U12007 ( .A1(n11912), .A2(n11914), .ZN(n12027) );
  NAND2_X1 U12008 ( .A1(n12028), .A2(n12029), .ZN(n11914) );
  NAND2_X1 U12009 ( .A1(b_14_), .A2(a_13_), .ZN(n12029) );
  INV_X1 U12010 ( .A(n12030), .ZN(n12028) );
  XOR2_X1 U12011 ( .A(n12031), .B(n12032), .Z(n11912) );
  XOR2_X1 U12012 ( .A(n12033), .B(n12034), .Z(n12031) );
  NOR2_X1 U12013 ( .A1(n7962), .A2(n7695), .ZN(n12034) );
  NAND2_X1 U12014 ( .A1(a_13_), .A2(n12030), .ZN(n11913) );
  NAND2_X1 U12015 ( .A1(n12035), .A2(n12036), .ZN(n12030) );
  NAND2_X1 U12016 ( .A1(n11908), .A2(n12037), .ZN(n12036) );
  OR2_X1 U12017 ( .A1(n11909), .A2(n11910), .ZN(n12037) );
  XNOR2_X1 U12018 ( .A(n12038), .B(n12039), .ZN(n11908) );
  XOR2_X1 U12019 ( .A(n12040), .B(n12041), .Z(n12039) );
  NAND2_X1 U12020 ( .A1(b_13_), .A2(a_15_), .ZN(n12041) );
  NAND2_X1 U12021 ( .A1(n11910), .A2(n11909), .ZN(n12035) );
  NAND2_X1 U12022 ( .A1(n12042), .A2(n12043), .ZN(n11909) );
  NAND2_X1 U12023 ( .A1(n11797), .A2(n12044), .ZN(n12043) );
  OR2_X1 U12024 ( .A1(n11796), .A2(n11795), .ZN(n12044) );
  NOR2_X1 U12025 ( .A1(n7961), .A2(n7667), .ZN(n11797) );
  NAND2_X1 U12026 ( .A1(n11795), .A2(n11796), .ZN(n12042) );
  NAND2_X1 U12027 ( .A1(n12045), .A2(n12046), .ZN(n11796) );
  NAND2_X1 U12028 ( .A1(n11804), .A2(n12047), .ZN(n12046) );
  OR2_X1 U12029 ( .A1(n11803), .A2(n11801), .ZN(n12047) );
  NOR2_X1 U12030 ( .A1(n7961), .A2(n8353), .ZN(n11804) );
  NAND2_X1 U12031 ( .A1(n11801), .A2(n11803), .ZN(n12045) );
  NAND2_X1 U12032 ( .A1(n12048), .A2(n12049), .ZN(n11803) );
  NAND3_X1 U12033 ( .A1(a_17_), .A2(n12050), .A3(b_14_), .ZN(n12049) );
  OR2_X1 U12034 ( .A1(n11905), .A2(n11904), .ZN(n12050) );
  NAND2_X1 U12035 ( .A1(n11904), .A2(n11905), .ZN(n12048) );
  NAND2_X1 U12036 ( .A1(n12051), .A2(n12052), .ZN(n11905) );
  NAND3_X1 U12037 ( .A1(a_18_), .A2(n12053), .A3(b_14_), .ZN(n12052) );
  NAND2_X1 U12038 ( .A1(n11901), .A2(n11900), .ZN(n12053) );
  OR2_X1 U12039 ( .A1(n11900), .A2(n11901), .ZN(n12051) );
  AND2_X1 U12040 ( .A1(n12054), .A2(n12055), .ZN(n11901) );
  NAND2_X1 U12041 ( .A1(n11898), .A2(n12056), .ZN(n12055) );
  OR2_X1 U12042 ( .A1(n11897), .A2(n11895), .ZN(n12056) );
  NOR2_X1 U12043 ( .A1(n7961), .A2(n7958), .ZN(n11898) );
  NAND2_X1 U12044 ( .A1(n11895), .A2(n11897), .ZN(n12054) );
  NAND2_X1 U12045 ( .A1(n12057), .A2(n12058), .ZN(n11897) );
  NAND3_X1 U12046 ( .A1(a_20_), .A2(n12059), .A3(b_14_), .ZN(n12058) );
  NAND2_X1 U12047 ( .A1(n11893), .A2(n11892), .ZN(n12059) );
  OR2_X1 U12048 ( .A1(n11892), .A2(n11893), .ZN(n12057) );
  AND2_X1 U12049 ( .A1(n12060), .A2(n12061), .ZN(n11893) );
  NAND2_X1 U12050 ( .A1(n11890), .A2(n12062), .ZN(n12061) );
  OR2_X1 U12051 ( .A1(n11889), .A2(n11888), .ZN(n12062) );
  NOR2_X1 U12052 ( .A1(n7961), .A2(n7578), .ZN(n11890) );
  NAND2_X1 U12053 ( .A1(n11888), .A2(n11889), .ZN(n12060) );
  NAND2_X1 U12054 ( .A1(n12063), .A2(n12064), .ZN(n11889) );
  NAND3_X1 U12055 ( .A1(a_22_), .A2(n12065), .A3(b_14_), .ZN(n12064) );
  OR2_X1 U12056 ( .A1(n11885), .A2(n11883), .ZN(n12065) );
  NAND2_X1 U12057 ( .A1(n11883), .A2(n11885), .ZN(n12063) );
  NAND2_X1 U12058 ( .A1(n12066), .A2(n12067), .ZN(n11885) );
  NAND2_X1 U12059 ( .A1(n11882), .A2(n12068), .ZN(n12067) );
  OR2_X1 U12060 ( .A1(n11881), .A2(n11879), .ZN(n12068) );
  NOR2_X1 U12061 ( .A1(n7961), .A2(n7955), .ZN(n11882) );
  NAND2_X1 U12062 ( .A1(n11879), .A2(n11881), .ZN(n12066) );
  NAND2_X1 U12063 ( .A1(n12069), .A2(n12070), .ZN(n11881) );
  NAND3_X1 U12064 ( .A1(a_24_), .A2(n12071), .A3(b_14_), .ZN(n12070) );
  NAND2_X1 U12065 ( .A1(n11877), .A2(n11876), .ZN(n12071) );
  OR2_X1 U12066 ( .A1(n11876), .A2(n11877), .ZN(n12069) );
  AND2_X1 U12067 ( .A1(n12072), .A2(n12073), .ZN(n11877) );
  NAND2_X1 U12068 ( .A1(n11874), .A2(n12074), .ZN(n12073) );
  OR2_X1 U12069 ( .A1(n11873), .A2(n11872), .ZN(n12074) );
  NOR2_X1 U12070 ( .A1(n7961), .A2(n7952), .ZN(n11874) );
  NAND2_X1 U12071 ( .A1(n11872), .A2(n11873), .ZN(n12072) );
  NAND2_X1 U12072 ( .A1(n11869), .A2(n12075), .ZN(n11873) );
  NAND2_X1 U12073 ( .A1(n11868), .A2(n11870), .ZN(n12075) );
  NAND2_X1 U12074 ( .A1(n12076), .A2(n12077), .ZN(n11870) );
  NAND2_X1 U12075 ( .A1(b_14_), .A2(a_26_), .ZN(n12077) );
  INV_X1 U12076 ( .A(n12078), .ZN(n12076) );
  XNOR2_X1 U12077 ( .A(n12079), .B(n12080), .ZN(n11868) );
  NAND2_X1 U12078 ( .A1(n12081), .A2(n12082), .ZN(n12079) );
  NAND2_X1 U12079 ( .A1(a_26_), .A2(n12078), .ZN(n11869) );
  NAND2_X1 U12080 ( .A1(n11841), .A2(n12083), .ZN(n12078) );
  NAND2_X1 U12081 ( .A1(n11840), .A2(n11842), .ZN(n12083) );
  NAND2_X1 U12082 ( .A1(n12084), .A2(n12085), .ZN(n11842) );
  NAND2_X1 U12083 ( .A1(b_14_), .A2(a_27_), .ZN(n12085) );
  INV_X1 U12084 ( .A(n12086), .ZN(n12084) );
  XNOR2_X1 U12085 ( .A(n12087), .B(n12088), .ZN(n11840) );
  XOR2_X1 U12086 ( .A(n12089), .B(n12090), .Z(n12087) );
  NAND2_X1 U12087 ( .A1(b_13_), .A2(a_28_), .ZN(n12089) );
  NAND2_X1 U12088 ( .A1(a_27_), .A2(n12086), .ZN(n11841) );
  NAND2_X1 U12089 ( .A1(n12091), .A2(n12092), .ZN(n12086) );
  NAND3_X1 U12090 ( .A1(a_28_), .A2(n12093), .A3(b_14_), .ZN(n12092) );
  NAND2_X1 U12091 ( .A1(n11850), .A2(n11848), .ZN(n12093) );
  OR2_X1 U12092 ( .A1(n11848), .A2(n11850), .ZN(n12091) );
  AND2_X1 U12093 ( .A1(n12094), .A2(n12095), .ZN(n11850) );
  NAND2_X1 U12094 ( .A1(n11864), .A2(n12096), .ZN(n12095) );
  OR2_X1 U12095 ( .A1(n11865), .A2(n11866), .ZN(n12096) );
  NOR2_X1 U12096 ( .A1(n7961), .A2(n7460), .ZN(n11864) );
  INV_X1 U12097 ( .A(b_14_), .ZN(n7961) );
  NAND2_X1 U12098 ( .A1(n11866), .A2(n11865), .ZN(n12094) );
  NAND2_X1 U12099 ( .A1(n12097), .A2(n12098), .ZN(n11865) );
  NAND2_X1 U12100 ( .A1(b_12_), .A2(n12099), .ZN(n12098) );
  NAND2_X1 U12101 ( .A1(n7441), .A2(n12100), .ZN(n12099) );
  NAND2_X1 U12102 ( .A1(a_31_), .A2(n7695), .ZN(n12100) );
  NAND2_X1 U12103 ( .A1(b_13_), .A2(n12101), .ZN(n12097) );
  NAND2_X1 U12104 ( .A1(n7445), .A2(n12102), .ZN(n12101) );
  NAND2_X1 U12105 ( .A1(a_30_), .A2(n12103), .ZN(n12102) );
  AND3_X1 U12106 ( .A1(b_13_), .A2(n7409), .A3(b_14_), .ZN(n11866) );
  XNOR2_X1 U12107 ( .A(n12104), .B(n12105), .ZN(n11848) );
  XOR2_X1 U12108 ( .A(n12106), .B(n12107), .Z(n12104) );
  XNOR2_X1 U12109 ( .A(n12108), .B(n12109), .ZN(n11872) );
  NAND2_X1 U12110 ( .A1(n12110), .A2(n12111), .ZN(n12108) );
  XNOR2_X1 U12111 ( .A(n12112), .B(n12113), .ZN(n11876) );
  XOR2_X1 U12112 ( .A(n12114), .B(n12115), .Z(n12112) );
  XNOR2_X1 U12113 ( .A(n12116), .B(n12117), .ZN(n11879) );
  XNOR2_X1 U12114 ( .A(n12118), .B(n12119), .ZN(n12116) );
  NOR2_X1 U12115 ( .A1(n7954), .A2(n7695), .ZN(n12119) );
  XNOR2_X1 U12116 ( .A(n12120), .B(n12121), .ZN(n11883) );
  XNOR2_X1 U12117 ( .A(n12122), .B(n12123), .ZN(n12121) );
  XNOR2_X1 U12118 ( .A(n12124), .B(n12125), .ZN(n11888) );
  XOR2_X1 U12119 ( .A(n12126), .B(n12127), .Z(n12125) );
  NAND2_X1 U12120 ( .A1(b_13_), .A2(a_22_), .ZN(n12127) );
  XNOR2_X1 U12121 ( .A(n12128), .B(n12129), .ZN(n11892) );
  XOR2_X1 U12122 ( .A(n12130), .B(n12131), .Z(n12128) );
  XNOR2_X1 U12123 ( .A(n12132), .B(n12133), .ZN(n11895) );
  XNOR2_X1 U12124 ( .A(n12134), .B(n12135), .ZN(n12132) );
  NOR2_X1 U12125 ( .A1(n7957), .A2(n7695), .ZN(n12135) );
  XOR2_X1 U12126 ( .A(n12136), .B(n12137), .Z(n11900) );
  XNOR2_X1 U12127 ( .A(n12138), .B(n12139), .ZN(n12137) );
  XNOR2_X1 U12128 ( .A(n12140), .B(n12141), .ZN(n11904) );
  XNOR2_X1 U12129 ( .A(n12142), .B(n12143), .ZN(n12140) );
  XNOR2_X1 U12130 ( .A(n12144), .B(n12145), .ZN(n11801) );
  XOR2_X1 U12131 ( .A(n12146), .B(n12147), .Z(n12144) );
  NAND2_X1 U12132 ( .A1(b_13_), .A2(a_17_), .ZN(n12146) );
  XNOR2_X1 U12133 ( .A(n12148), .B(n12149), .ZN(n11795) );
  XNOR2_X1 U12134 ( .A(n12150), .B(n12151), .ZN(n12148) );
  NOR2_X1 U12135 ( .A1(n8353), .A2(n7695), .ZN(n12151) );
  INV_X1 U12136 ( .A(n7681), .ZN(n11910) );
  NAND2_X1 U12137 ( .A1(b_14_), .A2(a_14_), .ZN(n7681) );
  XOR2_X1 U12138 ( .A(n12152), .B(n12153), .Z(n11916) );
  XOR2_X1 U12139 ( .A(n12154), .B(n7693), .Z(n12152) );
  XNOR2_X1 U12140 ( .A(n12155), .B(n12156), .ZN(n11920) );
  XNOR2_X1 U12141 ( .A(n12157), .B(n12158), .ZN(n12155) );
  NAND2_X1 U12142 ( .A1(b_13_), .A2(a_12_), .ZN(n12157) );
  XNOR2_X1 U12143 ( .A(n12159), .B(n12160), .ZN(n11924) );
  XOR2_X1 U12144 ( .A(n12161), .B(n12162), .Z(n12159) );
  NOR2_X1 U12145 ( .A1(n7724), .A2(n7695), .ZN(n12162) );
  XNOR2_X1 U12146 ( .A(n12163), .B(n12164), .ZN(n11927) );
  XNOR2_X1 U12147 ( .A(n12165), .B(n12166), .ZN(n12163) );
  NOR2_X1 U12148 ( .A1(n8378), .A2(n7695), .ZN(n12166) );
  XNOR2_X1 U12149 ( .A(n12167), .B(n12168), .ZN(n11947) );
  XNOR2_X1 U12150 ( .A(n12169), .B(n12170), .ZN(n12167) );
  NOR2_X1 U12151 ( .A1(n7823), .A2(n7695), .ZN(n12170) );
  XNOR2_X1 U12152 ( .A(n12171), .B(n12172), .ZN(n11951) );
  XOR2_X1 U12153 ( .A(n12173), .B(n12174), .Z(n12172) );
  NAND2_X1 U12154 ( .A1(b_13_), .A2(a_4_), .ZN(n12174) );
  XOR2_X1 U12155 ( .A(n12175), .B(n12176), .Z(n11956) );
  XOR2_X1 U12156 ( .A(n12177), .B(n12178), .Z(n12176) );
  NAND2_X1 U12157 ( .A1(b_13_), .A2(a_3_), .ZN(n12178) );
  XNOR2_X1 U12158 ( .A(n12179), .B(n12180), .ZN(n11959) );
  XNOR2_X1 U12159 ( .A(n12181), .B(n12182), .ZN(n12179) );
  NOR2_X1 U12160 ( .A1(n7966), .A2(n7695), .ZN(n12182) );
  XNOR2_X1 U12161 ( .A(n12183), .B(n12184), .ZN(n11963) );
  XOR2_X1 U12162 ( .A(n12185), .B(n12186), .Z(n12184) );
  NAND2_X1 U12163 ( .A1(b_13_), .A2(a_1_), .ZN(n12186) );
  NAND2_X1 U12164 ( .A1(n12187), .A2(n12188), .ZN(n8122) );
  XNOR2_X1 U12165 ( .A(n12189), .B(n12190), .ZN(n8123) );
  XNOR2_X1 U12166 ( .A(n12191), .B(n12192), .ZN(n12190) );
  NAND2_X1 U12167 ( .A1(n11967), .A2(n12193), .ZN(n8076) );
  XOR2_X1 U12168 ( .A(n8115), .B(n8114), .Z(n12193) );
  NOR2_X1 U12169 ( .A1(n12188), .A2(n12187), .ZN(n11967) );
  AND2_X1 U12170 ( .A1(n12194), .A2(n12195), .ZN(n12187) );
  NAND2_X1 U12171 ( .A1(n12192), .A2(n12196), .ZN(n12195) );
  OR2_X1 U12172 ( .A1(n12191), .A2(n12189), .ZN(n12196) );
  NOR2_X1 U12173 ( .A1(n7695), .A2(n8197), .ZN(n12192) );
  NAND2_X1 U12174 ( .A1(n12189), .A2(n12191), .ZN(n12194) );
  NAND2_X1 U12175 ( .A1(n12197), .A2(n12198), .ZN(n12191) );
  NAND3_X1 U12176 ( .A1(a_1_), .A2(n12199), .A3(b_13_), .ZN(n12198) );
  OR2_X1 U12177 ( .A1(n12185), .A2(n12183), .ZN(n12199) );
  NAND2_X1 U12178 ( .A1(n12183), .A2(n12185), .ZN(n12197) );
  NAND2_X1 U12179 ( .A1(n12200), .A2(n12201), .ZN(n12185) );
  NAND3_X1 U12180 ( .A1(a_2_), .A2(n12202), .A3(b_13_), .ZN(n12201) );
  NAND2_X1 U12181 ( .A1(n12181), .A2(n12180), .ZN(n12202) );
  OR2_X1 U12182 ( .A1(n12180), .A2(n12181), .ZN(n12200) );
  AND2_X1 U12183 ( .A1(n12203), .A2(n12204), .ZN(n12181) );
  NAND3_X1 U12184 ( .A1(a_3_), .A2(n12205), .A3(b_13_), .ZN(n12204) );
  OR2_X1 U12185 ( .A1(n12177), .A2(n12175), .ZN(n12205) );
  NAND2_X1 U12186 ( .A1(n12175), .A2(n12177), .ZN(n12203) );
  NAND2_X1 U12187 ( .A1(n12206), .A2(n12207), .ZN(n12177) );
  NAND3_X1 U12188 ( .A1(a_4_), .A2(n12208), .A3(b_13_), .ZN(n12207) );
  OR2_X1 U12189 ( .A1(n12173), .A2(n12171), .ZN(n12208) );
  NAND2_X1 U12190 ( .A1(n12171), .A2(n12173), .ZN(n12206) );
  NAND2_X1 U12191 ( .A1(n12209), .A2(n12210), .ZN(n12173) );
  NAND3_X1 U12192 ( .A1(a_5_), .A2(n12211), .A3(b_13_), .ZN(n12210) );
  NAND2_X1 U12193 ( .A1(n12169), .A2(n12168), .ZN(n12211) );
  OR2_X1 U12194 ( .A1(n12168), .A2(n12169), .ZN(n12209) );
  AND2_X1 U12195 ( .A1(n12212), .A2(n12213), .ZN(n12169) );
  NAND3_X1 U12196 ( .A1(a_6_), .A2(n12214), .A3(b_13_), .ZN(n12213) );
  OR2_X1 U12197 ( .A1(n11989), .A2(n11987), .ZN(n12214) );
  NAND2_X1 U12198 ( .A1(n11987), .A2(n11989), .ZN(n12212) );
  NAND2_X1 U12199 ( .A1(n12215), .A2(n12216), .ZN(n11989) );
  NAND3_X1 U12200 ( .A1(a_7_), .A2(n12217), .A3(b_13_), .ZN(n12216) );
  OR2_X1 U12201 ( .A1(n11997), .A2(n11995), .ZN(n12217) );
  NAND2_X1 U12202 ( .A1(n11995), .A2(n11997), .ZN(n12215) );
  NAND2_X1 U12203 ( .A1(n12218), .A2(n12219), .ZN(n11997) );
  NAND3_X1 U12204 ( .A1(a_8_), .A2(n12220), .A3(b_13_), .ZN(n12219) );
  NAND2_X1 U12205 ( .A1(n12005), .A2(n12004), .ZN(n12220) );
  OR2_X1 U12206 ( .A1(n12004), .A2(n12005), .ZN(n12218) );
  AND2_X1 U12207 ( .A1(n12221), .A2(n12222), .ZN(n12005) );
  NAND3_X1 U12208 ( .A1(a_9_), .A2(n12223), .A3(b_13_), .ZN(n12222) );
  OR2_X1 U12209 ( .A1(n12013), .A2(n12011), .ZN(n12223) );
  NAND2_X1 U12210 ( .A1(n12011), .A2(n12013), .ZN(n12221) );
  NAND2_X1 U12211 ( .A1(n12224), .A2(n12225), .ZN(n12013) );
  NAND3_X1 U12212 ( .A1(a_10_), .A2(n12226), .A3(b_13_), .ZN(n12225) );
  NAND2_X1 U12213 ( .A1(n12165), .A2(n12164), .ZN(n12226) );
  OR2_X1 U12214 ( .A1(n12164), .A2(n12165), .ZN(n12224) );
  AND2_X1 U12215 ( .A1(n12227), .A2(n12228), .ZN(n12165) );
  NAND3_X1 U12216 ( .A1(a_11_), .A2(n12229), .A3(b_13_), .ZN(n12228) );
  OR2_X1 U12217 ( .A1(n12161), .A2(n12160), .ZN(n12229) );
  NAND2_X1 U12218 ( .A1(n12160), .A2(n12161), .ZN(n12227) );
  NAND2_X1 U12219 ( .A1(n12230), .A2(n12231), .ZN(n12161) );
  NAND3_X1 U12220 ( .A1(a_12_), .A2(n12232), .A3(b_13_), .ZN(n12231) );
  OR2_X1 U12221 ( .A1(n12158), .A2(n12156), .ZN(n12232) );
  NAND2_X1 U12222 ( .A1(n12156), .A2(n12158), .ZN(n12230) );
  NAND2_X1 U12223 ( .A1(n12233), .A2(n12234), .ZN(n12158) );
  NAND2_X1 U12224 ( .A1(n12153), .A2(n12235), .ZN(n12234) );
  OR2_X1 U12225 ( .A1(n12154), .A2(n7693), .ZN(n12235) );
  XNOR2_X1 U12226 ( .A(n12236), .B(n12237), .ZN(n12153) );
  NAND2_X1 U12227 ( .A1(n12238), .A2(n12239), .ZN(n12236) );
  NAND2_X1 U12228 ( .A1(n7693), .A2(n12154), .ZN(n12233) );
  NAND2_X1 U12229 ( .A1(n12240), .A2(n12241), .ZN(n12154) );
  NAND3_X1 U12230 ( .A1(a_14_), .A2(n12242), .A3(b_13_), .ZN(n12241) );
  OR2_X1 U12231 ( .A1(n12033), .A2(n12032), .ZN(n12242) );
  NAND2_X1 U12232 ( .A1(n12032), .A2(n12033), .ZN(n12240) );
  NAND2_X1 U12233 ( .A1(n12243), .A2(n12244), .ZN(n12033) );
  NAND3_X1 U12234 ( .A1(a_15_), .A2(n12245), .A3(b_13_), .ZN(n12244) );
  OR2_X1 U12235 ( .A1(n12040), .A2(n12038), .ZN(n12245) );
  NAND2_X1 U12236 ( .A1(n12038), .A2(n12040), .ZN(n12243) );
  NAND2_X1 U12237 ( .A1(n12246), .A2(n12247), .ZN(n12040) );
  NAND3_X1 U12238 ( .A1(a_16_), .A2(n12248), .A3(b_13_), .ZN(n12247) );
  NAND2_X1 U12239 ( .A1(n12150), .A2(n12149), .ZN(n12248) );
  OR2_X1 U12240 ( .A1(n12149), .A2(n12150), .ZN(n12246) );
  AND2_X1 U12241 ( .A1(n12249), .A2(n12250), .ZN(n12150) );
  NAND3_X1 U12242 ( .A1(a_17_), .A2(n12251), .A3(b_13_), .ZN(n12250) );
  NAND2_X1 U12243 ( .A1(n12147), .A2(n12145), .ZN(n12251) );
  OR2_X1 U12244 ( .A1(n12145), .A2(n12147), .ZN(n12249) );
  AND2_X1 U12245 ( .A1(n12252), .A2(n12253), .ZN(n12147) );
  NAND2_X1 U12246 ( .A1(n12143), .A2(n12254), .ZN(n12253) );
  NAND2_X1 U12247 ( .A1(n12142), .A2(n12141), .ZN(n12254) );
  NOR2_X1 U12248 ( .A1(n7695), .A2(n7960), .ZN(n12143) );
  OR2_X1 U12249 ( .A1(n12141), .A2(n12142), .ZN(n12252) );
  AND2_X1 U12250 ( .A1(n12255), .A2(n12256), .ZN(n12142) );
  NAND2_X1 U12251 ( .A1(n12139), .A2(n12257), .ZN(n12256) );
  OR2_X1 U12252 ( .A1(n12138), .A2(n12136), .ZN(n12257) );
  NOR2_X1 U12253 ( .A1(n7695), .A2(n7958), .ZN(n12139) );
  NAND2_X1 U12254 ( .A1(n12136), .A2(n12138), .ZN(n12255) );
  NAND2_X1 U12255 ( .A1(n12258), .A2(n12259), .ZN(n12138) );
  NAND3_X1 U12256 ( .A1(a_20_), .A2(n12260), .A3(b_13_), .ZN(n12259) );
  NAND2_X1 U12257 ( .A1(n12134), .A2(n12133), .ZN(n12260) );
  OR2_X1 U12258 ( .A1(n12133), .A2(n12134), .ZN(n12258) );
  AND2_X1 U12259 ( .A1(n12261), .A2(n12262), .ZN(n12134) );
  NAND2_X1 U12260 ( .A1(n12131), .A2(n12263), .ZN(n12262) );
  OR2_X1 U12261 ( .A1(n12130), .A2(n12129), .ZN(n12263) );
  NOR2_X1 U12262 ( .A1(n7695), .A2(n7578), .ZN(n12131) );
  NAND2_X1 U12263 ( .A1(n12129), .A2(n12130), .ZN(n12261) );
  NAND2_X1 U12264 ( .A1(n12264), .A2(n12265), .ZN(n12130) );
  NAND3_X1 U12265 ( .A1(a_22_), .A2(n12266), .A3(b_13_), .ZN(n12265) );
  OR2_X1 U12266 ( .A1(n12126), .A2(n12124), .ZN(n12266) );
  NAND2_X1 U12267 ( .A1(n12124), .A2(n12126), .ZN(n12264) );
  NAND2_X1 U12268 ( .A1(n12267), .A2(n12268), .ZN(n12126) );
  NAND2_X1 U12269 ( .A1(n12123), .A2(n12269), .ZN(n12268) );
  OR2_X1 U12270 ( .A1(n12122), .A2(n12120), .ZN(n12269) );
  NOR2_X1 U12271 ( .A1(n7695), .A2(n7955), .ZN(n12123) );
  NAND2_X1 U12272 ( .A1(n12120), .A2(n12122), .ZN(n12267) );
  NAND2_X1 U12273 ( .A1(n12270), .A2(n12271), .ZN(n12122) );
  NAND3_X1 U12274 ( .A1(a_24_), .A2(n12272), .A3(b_13_), .ZN(n12271) );
  NAND2_X1 U12275 ( .A1(n12118), .A2(n12117), .ZN(n12272) );
  OR2_X1 U12276 ( .A1(n12117), .A2(n12118), .ZN(n12270) );
  AND2_X1 U12277 ( .A1(n12273), .A2(n12274), .ZN(n12118) );
  NAND2_X1 U12278 ( .A1(n12115), .A2(n12275), .ZN(n12274) );
  OR2_X1 U12279 ( .A1(n12114), .A2(n12113), .ZN(n12275) );
  NOR2_X1 U12280 ( .A1(n7695), .A2(n7952), .ZN(n12115) );
  NAND2_X1 U12281 ( .A1(n12113), .A2(n12114), .ZN(n12273) );
  NAND2_X1 U12282 ( .A1(n12110), .A2(n12276), .ZN(n12114) );
  NAND2_X1 U12283 ( .A1(n12109), .A2(n12111), .ZN(n12276) );
  NAND2_X1 U12284 ( .A1(n12277), .A2(n12278), .ZN(n12111) );
  NAND2_X1 U12285 ( .A1(b_13_), .A2(a_26_), .ZN(n12278) );
  INV_X1 U12286 ( .A(n12279), .ZN(n12277) );
  XNOR2_X1 U12287 ( .A(n12280), .B(n12281), .ZN(n12109) );
  NAND2_X1 U12288 ( .A1(n12282), .A2(n12283), .ZN(n12280) );
  NAND2_X1 U12289 ( .A1(a_26_), .A2(n12279), .ZN(n12110) );
  NAND2_X1 U12290 ( .A1(n12081), .A2(n12284), .ZN(n12279) );
  NAND2_X1 U12291 ( .A1(n12080), .A2(n12082), .ZN(n12284) );
  NAND2_X1 U12292 ( .A1(n12285), .A2(n12286), .ZN(n12082) );
  NAND2_X1 U12293 ( .A1(b_13_), .A2(a_27_), .ZN(n12286) );
  INV_X1 U12294 ( .A(n12287), .ZN(n12285) );
  XNOR2_X1 U12295 ( .A(n12288), .B(n12289), .ZN(n12080) );
  XOR2_X1 U12296 ( .A(n12290), .B(n12291), .Z(n12288) );
  NAND2_X1 U12297 ( .A1(b_12_), .A2(a_28_), .ZN(n12290) );
  NAND2_X1 U12298 ( .A1(a_27_), .A2(n12287), .ZN(n12081) );
  NAND2_X1 U12299 ( .A1(n12292), .A2(n12293), .ZN(n12287) );
  NAND3_X1 U12300 ( .A1(a_28_), .A2(n12294), .A3(b_13_), .ZN(n12293) );
  NAND2_X1 U12301 ( .A1(n12090), .A2(n12088), .ZN(n12294) );
  OR2_X1 U12302 ( .A1(n12088), .A2(n12090), .ZN(n12292) );
  AND2_X1 U12303 ( .A1(n12295), .A2(n12296), .ZN(n12090) );
  NAND2_X1 U12304 ( .A1(n12105), .A2(n12297), .ZN(n12296) );
  OR2_X1 U12305 ( .A1(n12106), .A2(n12107), .ZN(n12297) );
  NOR2_X1 U12306 ( .A1(n7695), .A2(n7460), .ZN(n12105) );
  INV_X1 U12307 ( .A(b_13_), .ZN(n7695) );
  NAND2_X1 U12308 ( .A1(n12107), .A2(n12106), .ZN(n12295) );
  NAND2_X1 U12309 ( .A1(n12298), .A2(n12299), .ZN(n12106) );
  NAND2_X1 U12310 ( .A1(b_11_), .A2(n12300), .ZN(n12299) );
  NAND2_X1 U12311 ( .A1(n7441), .A2(n12301), .ZN(n12300) );
  NAND2_X1 U12312 ( .A1(a_31_), .A2(n12103), .ZN(n12301) );
  NAND2_X1 U12313 ( .A1(b_12_), .A2(n12302), .ZN(n12298) );
  NAND2_X1 U12314 ( .A1(n7445), .A2(n12303), .ZN(n12302) );
  NAND2_X1 U12315 ( .A1(a_30_), .A2(n7726), .ZN(n12303) );
  AND3_X1 U12316 ( .A1(b_12_), .A2(n7409), .A3(b_13_), .ZN(n12107) );
  XNOR2_X1 U12317 ( .A(n12304), .B(n12305), .ZN(n12088) );
  XOR2_X1 U12318 ( .A(n12306), .B(n12307), .Z(n12304) );
  XNOR2_X1 U12319 ( .A(n12308), .B(n12309), .ZN(n12113) );
  NAND2_X1 U12320 ( .A1(n12310), .A2(n12311), .ZN(n12308) );
  XNOR2_X1 U12321 ( .A(n12312), .B(n12313), .ZN(n12117) );
  XOR2_X1 U12322 ( .A(n12314), .B(n12315), .Z(n12312) );
  XNOR2_X1 U12323 ( .A(n12316), .B(n12317), .ZN(n12120) );
  XNOR2_X1 U12324 ( .A(n12318), .B(n12319), .ZN(n12316) );
  NOR2_X1 U12325 ( .A1(n7954), .A2(n12103), .ZN(n12319) );
  XNOR2_X1 U12326 ( .A(n12320), .B(n12321), .ZN(n12124) );
  XNOR2_X1 U12327 ( .A(n12322), .B(n12323), .ZN(n12321) );
  XNOR2_X1 U12328 ( .A(n12324), .B(n12325), .ZN(n12129) );
  XOR2_X1 U12329 ( .A(n12326), .B(n12327), .Z(n12325) );
  NAND2_X1 U12330 ( .A1(b_12_), .A2(a_22_), .ZN(n12327) );
  XNOR2_X1 U12331 ( .A(n12328), .B(n12329), .ZN(n12133) );
  XOR2_X1 U12332 ( .A(n12330), .B(n12331), .Z(n12328) );
  XNOR2_X1 U12333 ( .A(n12332), .B(n12333), .ZN(n12136) );
  XNOR2_X1 U12334 ( .A(n12334), .B(n12335), .ZN(n12332) );
  NOR2_X1 U12335 ( .A1(n7957), .A2(n12103), .ZN(n12335) );
  XOR2_X1 U12336 ( .A(n12336), .B(n12337), .Z(n12141) );
  NAND2_X1 U12337 ( .A1(n12338), .A2(n12339), .ZN(n12336) );
  XNOR2_X1 U12338 ( .A(n12340), .B(n12341), .ZN(n12145) );
  XOR2_X1 U12339 ( .A(n12342), .B(n12343), .Z(n12340) );
  XNOR2_X1 U12340 ( .A(n12344), .B(n12345), .ZN(n12149) );
  XOR2_X1 U12341 ( .A(n12346), .B(n12347), .Z(n12344) );
  XNOR2_X1 U12342 ( .A(n12348), .B(n12349), .ZN(n12038) );
  XNOR2_X1 U12343 ( .A(n12350), .B(n12351), .ZN(n12348) );
  NOR2_X1 U12344 ( .A1(n8353), .A2(n12103), .ZN(n12351) );
  XNOR2_X1 U12345 ( .A(n12352), .B(n12353), .ZN(n12032) );
  NAND2_X1 U12346 ( .A1(n12354), .A2(n12355), .ZN(n12352) );
  INV_X1 U12347 ( .A(n7911), .ZN(n7693) );
  NAND2_X1 U12348 ( .A1(b_13_), .A2(a_13_), .ZN(n7911) );
  XNOR2_X1 U12349 ( .A(n12356), .B(n12357), .ZN(n12156) );
  XNOR2_X1 U12350 ( .A(n12358), .B(n12359), .ZN(n12357) );
  XNOR2_X1 U12351 ( .A(n12360), .B(n12361), .ZN(n12160) );
  XNOR2_X1 U12352 ( .A(n12362), .B(n7709), .ZN(n12361) );
  XOR2_X1 U12353 ( .A(n12363), .B(n12364), .Z(n12164) );
  NAND2_X1 U12354 ( .A1(n12365), .A2(n12366), .ZN(n12363) );
  XNOR2_X1 U12355 ( .A(n12367), .B(n12368), .ZN(n12011) );
  NAND2_X1 U12356 ( .A1(n12369), .A2(n12370), .ZN(n12367) );
  XOR2_X1 U12357 ( .A(n12371), .B(n12372), .Z(n12004) );
  XNOR2_X1 U12358 ( .A(n12373), .B(n12374), .ZN(n12372) );
  XOR2_X1 U12359 ( .A(n12375), .B(n12376), .Z(n11995) );
  XOR2_X1 U12360 ( .A(n12377), .B(n12378), .Z(n12375) );
  NOR2_X1 U12361 ( .A1(n8602), .A2(n12103), .ZN(n12378) );
  XNOR2_X1 U12362 ( .A(n12379), .B(n12380), .ZN(n11987) );
  NAND2_X1 U12363 ( .A1(n12381), .A2(n12382), .ZN(n12379) );
  XNOR2_X1 U12364 ( .A(n12383), .B(n12384), .ZN(n12168) );
  XOR2_X1 U12365 ( .A(n12385), .B(n12386), .Z(n12383) );
  XNOR2_X1 U12366 ( .A(n12387), .B(n12388), .ZN(n12171) );
  XOR2_X1 U12367 ( .A(n12389), .B(n12390), .Z(n12388) );
  NAND2_X1 U12368 ( .A1(b_12_), .A2(a_5_), .ZN(n12390) );
  XNOR2_X1 U12369 ( .A(n12391), .B(n12392), .ZN(n12175) );
  XNOR2_X1 U12370 ( .A(n12393), .B(n12394), .ZN(n12392) );
  XNOR2_X1 U12371 ( .A(n12395), .B(n12396), .ZN(n12180) );
  XOR2_X1 U12372 ( .A(n12397), .B(n12398), .Z(n12395) );
  NOR2_X1 U12373 ( .A1(n7852), .A2(n12103), .ZN(n12398) );
  XNOR2_X1 U12374 ( .A(n12399), .B(n12400), .ZN(n12183) );
  XNOR2_X1 U12375 ( .A(n12401), .B(n12402), .ZN(n12400) );
  XNOR2_X1 U12376 ( .A(n12403), .B(n12404), .ZN(n12189) );
  XNOR2_X1 U12377 ( .A(n12405), .B(n12406), .ZN(n12403) );
  XOR2_X1 U12378 ( .A(n12407), .B(n12408), .Z(n12188) );
  XOR2_X1 U12379 ( .A(n12409), .B(n12410), .Z(n12408) );
  NAND2_X1 U12380 ( .A1(b_12_), .A2(a_0_), .ZN(n12410) );
  NAND4_X1 U12381 ( .A1(n8114), .A2(n8113), .A3(n8115), .A4(n8107), .ZN(n8081)
         );
  INV_X1 U12382 ( .A(n12411), .ZN(n8107) );
  NAND2_X1 U12383 ( .A1(n12412), .A2(n12413), .ZN(n8115) );
  NAND3_X1 U12384 ( .A1(a_0_), .A2(n12414), .A3(b_12_), .ZN(n12413) );
  OR2_X1 U12385 ( .A1(n12409), .A2(n12407), .ZN(n12414) );
  NAND2_X1 U12386 ( .A1(n12407), .A2(n12409), .ZN(n12412) );
  NAND2_X1 U12387 ( .A1(n12415), .A2(n12416), .ZN(n12409) );
  NAND2_X1 U12388 ( .A1(n12406), .A2(n12417), .ZN(n12416) );
  NAND2_X1 U12389 ( .A1(n12405), .A2(n12404), .ZN(n12417) );
  NOR2_X1 U12390 ( .A1(n12103), .A2(n7872), .ZN(n12406) );
  OR2_X1 U12391 ( .A1(n12404), .A2(n12405), .ZN(n12415) );
  AND2_X1 U12392 ( .A1(n12418), .A2(n12419), .ZN(n12405) );
  NAND2_X1 U12393 ( .A1(n12402), .A2(n12420), .ZN(n12419) );
  OR2_X1 U12394 ( .A1(n12401), .A2(n12399), .ZN(n12420) );
  NOR2_X1 U12395 ( .A1(n12103), .A2(n7966), .ZN(n12402) );
  NAND2_X1 U12396 ( .A1(n12399), .A2(n12401), .ZN(n12418) );
  NAND2_X1 U12397 ( .A1(n12421), .A2(n12422), .ZN(n12401) );
  NAND3_X1 U12398 ( .A1(a_3_), .A2(n12423), .A3(b_12_), .ZN(n12422) );
  OR2_X1 U12399 ( .A1(n12397), .A2(n12396), .ZN(n12423) );
  NAND2_X1 U12400 ( .A1(n12396), .A2(n12397), .ZN(n12421) );
  NAND2_X1 U12401 ( .A1(n12424), .A2(n12425), .ZN(n12397) );
  NAND2_X1 U12402 ( .A1(n12394), .A2(n12426), .ZN(n12425) );
  OR2_X1 U12403 ( .A1(n12393), .A2(n12391), .ZN(n12426) );
  NOR2_X1 U12404 ( .A1(n12103), .A2(n7836), .ZN(n12394) );
  NAND2_X1 U12405 ( .A1(n12391), .A2(n12393), .ZN(n12424) );
  NAND2_X1 U12406 ( .A1(n12427), .A2(n12428), .ZN(n12393) );
  NAND3_X1 U12407 ( .A1(a_5_), .A2(n12429), .A3(b_12_), .ZN(n12428) );
  OR2_X1 U12408 ( .A1(n12389), .A2(n12387), .ZN(n12429) );
  NAND2_X1 U12409 ( .A1(n12387), .A2(n12389), .ZN(n12427) );
  NAND2_X1 U12410 ( .A1(n12430), .A2(n12431), .ZN(n12389) );
  NAND2_X1 U12411 ( .A1(n12385), .A2(n12432), .ZN(n12431) );
  OR2_X1 U12412 ( .A1(n12386), .A2(n12384), .ZN(n12432) );
  NOR2_X1 U12413 ( .A1(n12103), .A2(n7807), .ZN(n12385) );
  NAND2_X1 U12414 ( .A1(n12384), .A2(n12386), .ZN(n12430) );
  NAND2_X1 U12415 ( .A1(n12381), .A2(n12433), .ZN(n12386) );
  NAND2_X1 U12416 ( .A1(n12380), .A2(n12382), .ZN(n12433) );
  NAND2_X1 U12417 ( .A1(n12434), .A2(n12435), .ZN(n12382) );
  NAND2_X1 U12418 ( .A1(b_12_), .A2(a_7_), .ZN(n12435) );
  INV_X1 U12419 ( .A(n12436), .ZN(n12434) );
  XNOR2_X1 U12420 ( .A(n12437), .B(n12438), .ZN(n12380) );
  XOR2_X1 U12421 ( .A(n12439), .B(n12440), .Z(n12438) );
  NAND2_X1 U12422 ( .A1(a_8_), .A2(b_11_), .ZN(n12440) );
  NAND2_X1 U12423 ( .A1(a_7_), .A2(n12436), .ZN(n12381) );
  NAND2_X1 U12424 ( .A1(n12441), .A2(n12442), .ZN(n12436) );
  NAND3_X1 U12425 ( .A1(a_8_), .A2(n12443), .A3(b_12_), .ZN(n12442) );
  OR2_X1 U12426 ( .A1(n12377), .A2(n12376), .ZN(n12443) );
  NAND2_X1 U12427 ( .A1(n12376), .A2(n12377), .ZN(n12441) );
  NAND2_X1 U12428 ( .A1(n12444), .A2(n12445), .ZN(n12377) );
  NAND2_X1 U12429 ( .A1(n12374), .A2(n12446), .ZN(n12445) );
  OR2_X1 U12430 ( .A1(n12373), .A2(n12371), .ZN(n12446) );
  NOR2_X1 U12431 ( .A1(n12103), .A2(n7753), .ZN(n12374) );
  NAND2_X1 U12432 ( .A1(n12371), .A2(n12373), .ZN(n12444) );
  NAND2_X1 U12433 ( .A1(n12369), .A2(n12447), .ZN(n12373) );
  NAND2_X1 U12434 ( .A1(n12368), .A2(n12370), .ZN(n12447) );
  NAND2_X1 U12435 ( .A1(n12448), .A2(n12449), .ZN(n12370) );
  NAND2_X1 U12436 ( .A1(b_12_), .A2(a_10_), .ZN(n12449) );
  INV_X1 U12437 ( .A(n12450), .ZN(n12448) );
  XOR2_X1 U12438 ( .A(n12451), .B(n12452), .Z(n12368) );
  XOR2_X1 U12439 ( .A(n12453), .B(n7721), .Z(n12451) );
  NAND2_X1 U12440 ( .A1(a_10_), .A2(n12450), .ZN(n12369) );
  NAND2_X1 U12441 ( .A1(n12365), .A2(n12454), .ZN(n12450) );
  NAND2_X1 U12442 ( .A1(n12364), .A2(n12366), .ZN(n12454) );
  NAND2_X1 U12443 ( .A1(n12455), .A2(n12456), .ZN(n12366) );
  NAND2_X1 U12444 ( .A1(b_12_), .A2(a_11_), .ZN(n12456) );
  INV_X1 U12445 ( .A(n12457), .ZN(n12455) );
  XOR2_X1 U12446 ( .A(n12458), .B(n12459), .Z(n12364) );
  XOR2_X1 U12447 ( .A(n12460), .B(n12461), .Z(n12458) );
  NOR2_X1 U12448 ( .A1(n7726), .A2(n8585), .ZN(n12461) );
  NAND2_X1 U12449 ( .A1(a_11_), .A2(n12457), .ZN(n12365) );
  NAND2_X1 U12450 ( .A1(n12462), .A2(n12463), .ZN(n12457) );
  NAND2_X1 U12451 ( .A1(n12360), .A2(n12464), .ZN(n12463) );
  OR2_X1 U12452 ( .A1(n12362), .A2(n7709), .ZN(n12464) );
  XNOR2_X1 U12453 ( .A(n12465), .B(n12466), .ZN(n12360) );
  XOR2_X1 U12454 ( .A(n12467), .B(n12468), .Z(n12466) );
  NAND2_X1 U12455 ( .A1(a_13_), .A2(b_11_), .ZN(n12468) );
  NAND2_X1 U12456 ( .A1(n7709), .A2(n12362), .ZN(n12462) );
  NAND2_X1 U12457 ( .A1(n12469), .A2(n12470), .ZN(n12362) );
  NAND2_X1 U12458 ( .A1(n12359), .A2(n12471), .ZN(n12470) );
  OR2_X1 U12459 ( .A1(n12358), .A2(n12356), .ZN(n12471) );
  NOR2_X1 U12460 ( .A1(n12103), .A2(n7702), .ZN(n12359) );
  NAND2_X1 U12461 ( .A1(n12356), .A2(n12358), .ZN(n12469) );
  NAND2_X1 U12462 ( .A1(n12238), .A2(n12472), .ZN(n12358) );
  NAND2_X1 U12463 ( .A1(n12237), .A2(n12239), .ZN(n12472) );
  NAND2_X1 U12464 ( .A1(n12473), .A2(n12474), .ZN(n12239) );
  NAND2_X1 U12465 ( .A1(b_12_), .A2(a_14_), .ZN(n12474) );
  INV_X1 U12466 ( .A(n12475), .ZN(n12473) );
  XNOR2_X1 U12467 ( .A(n12476), .B(n12477), .ZN(n12237) );
  XOR2_X1 U12468 ( .A(n12478), .B(n12479), .Z(n12477) );
  NAND2_X1 U12469 ( .A1(a_15_), .A2(b_11_), .ZN(n12479) );
  NAND2_X1 U12470 ( .A1(a_14_), .A2(n12475), .ZN(n12238) );
  NAND2_X1 U12471 ( .A1(n12354), .A2(n12480), .ZN(n12475) );
  NAND2_X1 U12472 ( .A1(n12353), .A2(n12355), .ZN(n12480) );
  NAND2_X1 U12473 ( .A1(n12481), .A2(n12482), .ZN(n12355) );
  NAND2_X1 U12474 ( .A1(b_12_), .A2(a_15_), .ZN(n12482) );
  INV_X1 U12475 ( .A(n12483), .ZN(n12481) );
  XNOR2_X1 U12476 ( .A(n12484), .B(n12485), .ZN(n12353) );
  XNOR2_X1 U12477 ( .A(n12486), .B(n12487), .ZN(n12484) );
  NOR2_X1 U12478 ( .A1(n7726), .A2(n8353), .ZN(n12487) );
  NAND2_X1 U12479 ( .A1(a_15_), .A2(n12483), .ZN(n12354) );
  NAND2_X1 U12480 ( .A1(n12488), .A2(n12489), .ZN(n12483) );
  NAND3_X1 U12481 ( .A1(a_16_), .A2(n12490), .A3(b_12_), .ZN(n12489) );
  NAND2_X1 U12482 ( .A1(n12350), .A2(n12349), .ZN(n12490) );
  OR2_X1 U12483 ( .A1(n12349), .A2(n12350), .ZN(n12488) );
  AND2_X1 U12484 ( .A1(n12491), .A2(n12492), .ZN(n12350) );
  NAND2_X1 U12485 ( .A1(n12346), .A2(n12493), .ZN(n12492) );
  OR2_X1 U12486 ( .A1(n12347), .A2(n12345), .ZN(n12493) );
  NOR2_X1 U12487 ( .A1(n12103), .A2(n7645), .ZN(n12346) );
  NAND2_X1 U12488 ( .A1(n12345), .A2(n12347), .ZN(n12491) );
  NAND2_X1 U12489 ( .A1(n12494), .A2(n12495), .ZN(n12347) );
  NAND2_X1 U12490 ( .A1(n12342), .A2(n12496), .ZN(n12495) );
  OR2_X1 U12491 ( .A1(n12343), .A2(n12341), .ZN(n12496) );
  NOR2_X1 U12492 ( .A1(n12103), .A2(n7960), .ZN(n12342) );
  NAND2_X1 U12493 ( .A1(n12341), .A2(n12343), .ZN(n12494) );
  NAND2_X1 U12494 ( .A1(n12338), .A2(n12497), .ZN(n12343) );
  NAND2_X1 U12495 ( .A1(n12337), .A2(n12339), .ZN(n12497) );
  NAND2_X1 U12496 ( .A1(n12498), .A2(n12499), .ZN(n12339) );
  NAND2_X1 U12497 ( .A1(b_12_), .A2(a_19_), .ZN(n12499) );
  INV_X1 U12498 ( .A(n12500), .ZN(n12498) );
  XOR2_X1 U12499 ( .A(n12501), .B(n12502), .Z(n12337) );
  XOR2_X1 U12500 ( .A(n12503), .B(n12504), .Z(n12501) );
  NOR2_X1 U12501 ( .A1(n7726), .A2(n7957), .ZN(n12504) );
  NAND2_X1 U12502 ( .A1(a_19_), .A2(n12500), .ZN(n12338) );
  NAND2_X1 U12503 ( .A1(n12505), .A2(n12506), .ZN(n12500) );
  NAND3_X1 U12504 ( .A1(a_20_), .A2(n12507), .A3(b_12_), .ZN(n12506) );
  NAND2_X1 U12505 ( .A1(n12334), .A2(n12333), .ZN(n12507) );
  OR2_X1 U12506 ( .A1(n12333), .A2(n12334), .ZN(n12505) );
  AND2_X1 U12507 ( .A1(n12508), .A2(n12509), .ZN(n12334) );
  NAND2_X1 U12508 ( .A1(n12331), .A2(n12510), .ZN(n12509) );
  OR2_X1 U12509 ( .A1(n12330), .A2(n12329), .ZN(n12510) );
  NOR2_X1 U12510 ( .A1(n12103), .A2(n7578), .ZN(n12331) );
  NAND2_X1 U12511 ( .A1(n12329), .A2(n12330), .ZN(n12508) );
  NAND2_X1 U12512 ( .A1(n12511), .A2(n12512), .ZN(n12330) );
  NAND3_X1 U12513 ( .A1(a_22_), .A2(n12513), .A3(b_12_), .ZN(n12512) );
  OR2_X1 U12514 ( .A1(n12326), .A2(n12324), .ZN(n12513) );
  NAND2_X1 U12515 ( .A1(n12324), .A2(n12326), .ZN(n12511) );
  NAND2_X1 U12516 ( .A1(n12514), .A2(n12515), .ZN(n12326) );
  NAND2_X1 U12517 ( .A1(n12323), .A2(n12516), .ZN(n12515) );
  OR2_X1 U12518 ( .A1(n12322), .A2(n12320), .ZN(n12516) );
  NOR2_X1 U12519 ( .A1(n12103), .A2(n7955), .ZN(n12323) );
  NAND2_X1 U12520 ( .A1(n12320), .A2(n12322), .ZN(n12514) );
  NAND2_X1 U12521 ( .A1(n12517), .A2(n12518), .ZN(n12322) );
  NAND3_X1 U12522 ( .A1(a_24_), .A2(n12519), .A3(b_12_), .ZN(n12518) );
  NAND2_X1 U12523 ( .A1(n12318), .A2(n12317), .ZN(n12519) );
  OR2_X1 U12524 ( .A1(n12317), .A2(n12318), .ZN(n12517) );
  AND2_X1 U12525 ( .A1(n12520), .A2(n12521), .ZN(n12318) );
  NAND2_X1 U12526 ( .A1(n12315), .A2(n12522), .ZN(n12521) );
  OR2_X1 U12527 ( .A1(n12314), .A2(n12313), .ZN(n12522) );
  NOR2_X1 U12528 ( .A1(n12103), .A2(n7952), .ZN(n12315) );
  NAND2_X1 U12529 ( .A1(n12313), .A2(n12314), .ZN(n12520) );
  NAND2_X1 U12530 ( .A1(n12310), .A2(n12523), .ZN(n12314) );
  NAND2_X1 U12531 ( .A1(n12309), .A2(n12311), .ZN(n12523) );
  NAND2_X1 U12532 ( .A1(n12524), .A2(n12525), .ZN(n12311) );
  NAND2_X1 U12533 ( .A1(b_12_), .A2(a_26_), .ZN(n12525) );
  INV_X1 U12534 ( .A(n12526), .ZN(n12524) );
  XNOR2_X1 U12535 ( .A(n12527), .B(n12528), .ZN(n12309) );
  NAND2_X1 U12536 ( .A1(n12529), .A2(n12530), .ZN(n12527) );
  NAND2_X1 U12537 ( .A1(a_26_), .A2(n12526), .ZN(n12310) );
  NAND2_X1 U12538 ( .A1(n12282), .A2(n12531), .ZN(n12526) );
  NAND2_X1 U12539 ( .A1(n12281), .A2(n12283), .ZN(n12531) );
  NAND2_X1 U12540 ( .A1(n12532), .A2(n12533), .ZN(n12283) );
  NAND2_X1 U12541 ( .A1(b_12_), .A2(a_27_), .ZN(n12533) );
  INV_X1 U12542 ( .A(n12534), .ZN(n12532) );
  XNOR2_X1 U12543 ( .A(n12535), .B(n12536), .ZN(n12281) );
  XOR2_X1 U12544 ( .A(n12537), .B(n12538), .Z(n12535) );
  NAND2_X1 U12545 ( .A1(a_28_), .A2(b_11_), .ZN(n12537) );
  NAND2_X1 U12546 ( .A1(a_27_), .A2(n12534), .ZN(n12282) );
  NAND2_X1 U12547 ( .A1(n12539), .A2(n12540), .ZN(n12534) );
  NAND3_X1 U12548 ( .A1(a_28_), .A2(n12541), .A3(b_12_), .ZN(n12540) );
  NAND2_X1 U12549 ( .A1(n12291), .A2(n12289), .ZN(n12541) );
  OR2_X1 U12550 ( .A1(n12289), .A2(n12291), .ZN(n12539) );
  AND2_X1 U12551 ( .A1(n12542), .A2(n12543), .ZN(n12291) );
  NAND2_X1 U12552 ( .A1(n12305), .A2(n12544), .ZN(n12543) );
  OR2_X1 U12553 ( .A1(n12306), .A2(n12307), .ZN(n12544) );
  NOR2_X1 U12554 ( .A1(n12103), .A2(n7460), .ZN(n12305) );
  NAND2_X1 U12555 ( .A1(n12307), .A2(n12306), .ZN(n12542) );
  NAND2_X1 U12556 ( .A1(n12545), .A2(n12546), .ZN(n12306) );
  NAND2_X1 U12557 ( .A1(b_10_), .A2(n12547), .ZN(n12546) );
  NAND2_X1 U12558 ( .A1(n7441), .A2(n12548), .ZN(n12547) );
  NAND2_X1 U12559 ( .A1(a_31_), .A2(n7726), .ZN(n12548) );
  NAND2_X1 U12560 ( .A1(b_11_), .A2(n12549), .ZN(n12545) );
  NAND2_X1 U12561 ( .A1(n7445), .A2(n12550), .ZN(n12549) );
  NAND2_X1 U12562 ( .A1(a_30_), .A2(n12551), .ZN(n12550) );
  AND3_X1 U12563 ( .A1(n7409), .A2(b_11_), .A3(b_12_), .ZN(n12307) );
  XNOR2_X1 U12564 ( .A(n12552), .B(n12553), .ZN(n12289) );
  XOR2_X1 U12565 ( .A(n12554), .B(n12555), .Z(n12552) );
  XNOR2_X1 U12566 ( .A(n12556), .B(n12557), .ZN(n12313) );
  NAND2_X1 U12567 ( .A1(n12558), .A2(n12559), .ZN(n12556) );
  XNOR2_X1 U12568 ( .A(n12560), .B(n12561), .ZN(n12317) );
  XOR2_X1 U12569 ( .A(n12562), .B(n12563), .Z(n12560) );
  XNOR2_X1 U12570 ( .A(n12564), .B(n12565), .ZN(n12320) );
  XNOR2_X1 U12571 ( .A(n12566), .B(n12567), .ZN(n12564) );
  NOR2_X1 U12572 ( .A1(n7726), .A2(n7954), .ZN(n12567) );
  XNOR2_X1 U12573 ( .A(n12568), .B(n12569), .ZN(n12324) );
  XNOR2_X1 U12574 ( .A(n12570), .B(n12571), .ZN(n12569) );
  XNOR2_X1 U12575 ( .A(n12572), .B(n12573), .ZN(n12329) );
  XOR2_X1 U12576 ( .A(n12574), .B(n12575), .Z(n12573) );
  NAND2_X1 U12577 ( .A1(a_22_), .A2(b_11_), .ZN(n12575) );
  XNOR2_X1 U12578 ( .A(n12576), .B(n12577), .ZN(n12333) );
  XOR2_X1 U12579 ( .A(n12578), .B(n12579), .Z(n12576) );
  XNOR2_X1 U12580 ( .A(n12580), .B(n12581), .ZN(n12341) );
  NAND2_X1 U12581 ( .A1(n12582), .A2(n12583), .ZN(n12580) );
  XNOR2_X1 U12582 ( .A(n12584), .B(n12585), .ZN(n12345) );
  NAND2_X1 U12583 ( .A1(n12586), .A2(n12587), .ZN(n12584) );
  XOR2_X1 U12584 ( .A(n12588), .B(n12589), .Z(n12349) );
  XOR2_X1 U12585 ( .A(n12590), .B(n12591), .Z(n12589) );
  NAND2_X1 U12586 ( .A1(a_17_), .A2(b_11_), .ZN(n12591) );
  XOR2_X1 U12587 ( .A(n12592), .B(n12593), .Z(n12356) );
  XOR2_X1 U12588 ( .A(n12594), .B(n12595), .Z(n12592) );
  NOR2_X1 U12589 ( .A1(n7726), .A2(n7962), .ZN(n12595) );
  NOR2_X1 U12590 ( .A1(n12103), .A2(n8585), .ZN(n7709) );
  INV_X1 U12591 ( .A(b_12_), .ZN(n12103) );
  XNOR2_X1 U12592 ( .A(n12596), .B(n12597), .ZN(n12371) );
  XNOR2_X1 U12593 ( .A(n12598), .B(n12599), .ZN(n12596) );
  NOR2_X1 U12594 ( .A1(n7726), .A2(n8378), .ZN(n12599) );
  XNOR2_X1 U12595 ( .A(n12600), .B(n12601), .ZN(n12376) );
  XNOR2_X1 U12596 ( .A(n12602), .B(n12603), .ZN(n12600) );
  NOR2_X1 U12597 ( .A1(n7726), .A2(n7753), .ZN(n12603) );
  XNOR2_X1 U12598 ( .A(n12604), .B(n12605), .ZN(n12384) );
  XNOR2_X1 U12599 ( .A(n12606), .B(n12607), .ZN(n12604) );
  NOR2_X1 U12600 ( .A1(n7726), .A2(n7787), .ZN(n12607) );
  XOR2_X1 U12601 ( .A(n12608), .B(n12609), .Z(n12387) );
  XOR2_X1 U12602 ( .A(n12610), .B(n12611), .Z(n12608) );
  NOR2_X1 U12603 ( .A1(n7726), .A2(n7807), .ZN(n12611) );
  XNOR2_X1 U12604 ( .A(n12612), .B(n12613), .ZN(n12391) );
  XOR2_X1 U12605 ( .A(n12614), .B(n12615), .Z(n12613) );
  NAND2_X1 U12606 ( .A1(a_5_), .A2(b_11_), .ZN(n12615) );
  XNOR2_X1 U12607 ( .A(n12616), .B(n12617), .ZN(n12396) );
  XNOR2_X1 U12608 ( .A(n12618), .B(n12619), .ZN(n12616) );
  NOR2_X1 U12609 ( .A1(n7726), .A2(n7836), .ZN(n12619) );
  XNOR2_X1 U12610 ( .A(n12620), .B(n12621), .ZN(n12399) );
  XOR2_X1 U12611 ( .A(n12622), .B(n12623), .Z(n12621) );
  NAND2_X1 U12612 ( .A1(a_3_), .A2(b_11_), .ZN(n12623) );
  XNOR2_X1 U12613 ( .A(n12624), .B(n12625), .ZN(n12404) );
  XOR2_X1 U12614 ( .A(n12626), .B(n12627), .Z(n12624) );
  NOR2_X1 U12615 ( .A1(n7726), .A2(n7966), .ZN(n12627) );
  XOR2_X1 U12616 ( .A(n12628), .B(n12629), .Z(n12407) );
  XOR2_X1 U12617 ( .A(n12630), .B(n12631), .Z(n12628) );
  NOR2_X1 U12618 ( .A1(n7726), .A2(n7872), .ZN(n12631) );
  NAND2_X1 U12619 ( .A1(n12632), .A2(n12633), .ZN(n8113) );
  XNOR2_X1 U12620 ( .A(n12634), .B(n12635), .ZN(n8114) );
  XNOR2_X1 U12621 ( .A(n12636), .B(n12637), .ZN(n12635) );
  NAND2_X1 U12622 ( .A1(n12411), .A2(n12638), .ZN(n8086) );
  XOR2_X1 U12623 ( .A(n8108), .B(n8109), .Z(n12638) );
  NOR2_X1 U12624 ( .A1(n12633), .A2(n12632), .ZN(n12411) );
  AND2_X1 U12625 ( .A1(n12639), .A2(n12640), .ZN(n12632) );
  NAND2_X1 U12626 ( .A1(n12637), .A2(n12641), .ZN(n12640) );
  OR2_X1 U12627 ( .A1(n12636), .A2(n12634), .ZN(n12641) );
  NOR2_X1 U12628 ( .A1(n7726), .A2(n8197), .ZN(n12637) );
  NAND2_X1 U12629 ( .A1(n12634), .A2(n12636), .ZN(n12639) );
  NAND2_X1 U12630 ( .A1(n12642), .A2(n12643), .ZN(n12636) );
  NAND3_X1 U12631 ( .A1(b_11_), .A2(n12644), .A3(a_1_), .ZN(n12643) );
  OR2_X1 U12632 ( .A1(n12630), .A2(n12629), .ZN(n12644) );
  NAND2_X1 U12633 ( .A1(n12629), .A2(n12630), .ZN(n12642) );
  NAND2_X1 U12634 ( .A1(n12645), .A2(n12646), .ZN(n12630) );
  NAND3_X1 U12635 ( .A1(b_11_), .A2(n12647), .A3(a_2_), .ZN(n12646) );
  OR2_X1 U12636 ( .A1(n12626), .A2(n12625), .ZN(n12647) );
  NAND2_X1 U12637 ( .A1(n12625), .A2(n12626), .ZN(n12645) );
  NAND2_X1 U12638 ( .A1(n12648), .A2(n12649), .ZN(n12626) );
  NAND3_X1 U12639 ( .A1(b_11_), .A2(n12650), .A3(a_3_), .ZN(n12649) );
  OR2_X1 U12640 ( .A1(n12622), .A2(n12620), .ZN(n12650) );
  NAND2_X1 U12641 ( .A1(n12620), .A2(n12622), .ZN(n12648) );
  NAND2_X1 U12642 ( .A1(n12651), .A2(n12652), .ZN(n12622) );
  NAND3_X1 U12643 ( .A1(b_11_), .A2(n12653), .A3(a_4_), .ZN(n12652) );
  NAND2_X1 U12644 ( .A1(n12618), .A2(n12617), .ZN(n12653) );
  OR2_X1 U12645 ( .A1(n12617), .A2(n12618), .ZN(n12651) );
  AND2_X1 U12646 ( .A1(n12654), .A2(n12655), .ZN(n12618) );
  NAND3_X1 U12647 ( .A1(b_11_), .A2(n12656), .A3(a_5_), .ZN(n12655) );
  OR2_X1 U12648 ( .A1(n12614), .A2(n12612), .ZN(n12656) );
  NAND2_X1 U12649 ( .A1(n12612), .A2(n12614), .ZN(n12654) );
  NAND2_X1 U12650 ( .A1(n12657), .A2(n12658), .ZN(n12614) );
  NAND3_X1 U12651 ( .A1(b_11_), .A2(n12659), .A3(a_6_), .ZN(n12658) );
  OR2_X1 U12652 ( .A1(n12610), .A2(n12609), .ZN(n12659) );
  NAND2_X1 U12653 ( .A1(n12609), .A2(n12610), .ZN(n12657) );
  NAND2_X1 U12654 ( .A1(n12660), .A2(n12661), .ZN(n12610) );
  NAND3_X1 U12655 ( .A1(b_11_), .A2(n12662), .A3(a_7_), .ZN(n12661) );
  NAND2_X1 U12656 ( .A1(n12606), .A2(n12605), .ZN(n12662) );
  OR2_X1 U12657 ( .A1(n12605), .A2(n12606), .ZN(n12660) );
  AND2_X1 U12658 ( .A1(n12663), .A2(n12664), .ZN(n12606) );
  NAND3_X1 U12659 ( .A1(b_11_), .A2(n12665), .A3(a_8_), .ZN(n12664) );
  OR2_X1 U12660 ( .A1(n12439), .A2(n12437), .ZN(n12665) );
  NAND2_X1 U12661 ( .A1(n12437), .A2(n12439), .ZN(n12663) );
  NAND2_X1 U12662 ( .A1(n12666), .A2(n12667), .ZN(n12439) );
  NAND3_X1 U12663 ( .A1(b_11_), .A2(n12668), .A3(a_9_), .ZN(n12667) );
  NAND2_X1 U12664 ( .A1(n12602), .A2(n12601), .ZN(n12668) );
  OR2_X1 U12665 ( .A1(n12601), .A2(n12602), .ZN(n12666) );
  AND2_X1 U12666 ( .A1(n12669), .A2(n12670), .ZN(n12602) );
  NAND3_X1 U12667 ( .A1(b_11_), .A2(n12671), .A3(a_10_), .ZN(n12670) );
  NAND2_X1 U12668 ( .A1(n12598), .A2(n12597), .ZN(n12671) );
  OR2_X1 U12669 ( .A1(n12597), .A2(n12598), .ZN(n12669) );
  AND2_X1 U12670 ( .A1(n12672), .A2(n12673), .ZN(n12598) );
  NAND2_X1 U12671 ( .A1(n12452), .A2(n12674), .ZN(n12673) );
  OR2_X1 U12672 ( .A1(n12453), .A2(n7721), .ZN(n12674) );
  XNOR2_X1 U12673 ( .A(n12675), .B(n12676), .ZN(n12452) );
  NAND2_X1 U12674 ( .A1(n12677), .A2(n12678), .ZN(n12675) );
  NAND2_X1 U12675 ( .A1(n7721), .A2(n12453), .ZN(n12672) );
  NAND2_X1 U12676 ( .A1(n12679), .A2(n12680), .ZN(n12453) );
  NAND3_X1 U12677 ( .A1(b_11_), .A2(n12681), .A3(a_12_), .ZN(n12680) );
  OR2_X1 U12678 ( .A1(n12460), .A2(n12459), .ZN(n12681) );
  NAND2_X1 U12679 ( .A1(n12459), .A2(n12460), .ZN(n12679) );
  NAND2_X1 U12680 ( .A1(n12682), .A2(n12683), .ZN(n12460) );
  NAND3_X1 U12681 ( .A1(b_11_), .A2(n12684), .A3(a_13_), .ZN(n12683) );
  OR2_X1 U12682 ( .A1(n12467), .A2(n12465), .ZN(n12684) );
  NAND2_X1 U12683 ( .A1(n12465), .A2(n12467), .ZN(n12682) );
  NAND2_X1 U12684 ( .A1(n12685), .A2(n12686), .ZN(n12467) );
  NAND3_X1 U12685 ( .A1(b_11_), .A2(n12687), .A3(a_14_), .ZN(n12686) );
  OR2_X1 U12686 ( .A1(n12594), .A2(n12593), .ZN(n12687) );
  NAND2_X1 U12687 ( .A1(n12593), .A2(n12594), .ZN(n12685) );
  NAND2_X1 U12688 ( .A1(n12688), .A2(n12689), .ZN(n12594) );
  NAND3_X1 U12689 ( .A1(b_11_), .A2(n12690), .A3(a_15_), .ZN(n12689) );
  OR2_X1 U12690 ( .A1(n12478), .A2(n12476), .ZN(n12690) );
  NAND2_X1 U12691 ( .A1(n12476), .A2(n12478), .ZN(n12688) );
  NAND2_X1 U12692 ( .A1(n12691), .A2(n12692), .ZN(n12478) );
  NAND3_X1 U12693 ( .A1(b_11_), .A2(n12693), .A3(a_16_), .ZN(n12692) );
  NAND2_X1 U12694 ( .A1(n12486), .A2(n12485), .ZN(n12693) );
  OR2_X1 U12695 ( .A1(n12485), .A2(n12486), .ZN(n12691) );
  AND2_X1 U12696 ( .A1(n12694), .A2(n12695), .ZN(n12486) );
  NAND3_X1 U12697 ( .A1(b_11_), .A2(n12696), .A3(a_17_), .ZN(n12695) );
  OR2_X1 U12698 ( .A1(n12590), .A2(n12588), .ZN(n12696) );
  NAND2_X1 U12699 ( .A1(n12588), .A2(n12590), .ZN(n12694) );
  NAND2_X1 U12700 ( .A1(n12586), .A2(n12697), .ZN(n12590) );
  NAND2_X1 U12701 ( .A1(n12585), .A2(n12587), .ZN(n12697) );
  NAND2_X1 U12702 ( .A1(n12698), .A2(n12699), .ZN(n12587) );
  NAND2_X1 U12703 ( .A1(a_18_), .A2(b_11_), .ZN(n12699) );
  INV_X1 U12704 ( .A(n12700), .ZN(n12698) );
  XNOR2_X1 U12705 ( .A(n12701), .B(n12702), .ZN(n12585) );
  XNOR2_X1 U12706 ( .A(n12703), .B(n12704), .ZN(n12702) );
  NAND2_X1 U12707 ( .A1(a_18_), .A2(n12700), .ZN(n12586) );
  NAND2_X1 U12708 ( .A1(n12582), .A2(n12705), .ZN(n12700) );
  NAND2_X1 U12709 ( .A1(n12581), .A2(n12583), .ZN(n12705) );
  NAND2_X1 U12710 ( .A1(n12706), .A2(n12707), .ZN(n12583) );
  NAND2_X1 U12711 ( .A1(a_19_), .A2(b_11_), .ZN(n12707) );
  INV_X1 U12712 ( .A(n12708), .ZN(n12706) );
  XNOR2_X1 U12713 ( .A(n12709), .B(n12710), .ZN(n12581) );
  XNOR2_X1 U12714 ( .A(n12711), .B(n12712), .ZN(n12710) );
  NAND2_X1 U12715 ( .A1(a_19_), .A2(n12708), .ZN(n12582) );
  NAND2_X1 U12716 ( .A1(n12713), .A2(n12714), .ZN(n12708) );
  NAND3_X1 U12717 ( .A1(b_11_), .A2(n12715), .A3(a_20_), .ZN(n12714) );
  OR2_X1 U12718 ( .A1(n12503), .A2(n12502), .ZN(n12715) );
  NAND2_X1 U12719 ( .A1(n12502), .A2(n12503), .ZN(n12713) );
  NAND2_X1 U12720 ( .A1(n12716), .A2(n12717), .ZN(n12503) );
  NAND2_X1 U12721 ( .A1(n12579), .A2(n12718), .ZN(n12717) );
  OR2_X1 U12722 ( .A1(n12578), .A2(n12577), .ZN(n12718) );
  NOR2_X1 U12723 ( .A1(n7578), .A2(n7726), .ZN(n12579) );
  NAND2_X1 U12724 ( .A1(n12577), .A2(n12578), .ZN(n12716) );
  NAND2_X1 U12725 ( .A1(n12719), .A2(n12720), .ZN(n12578) );
  NAND3_X1 U12726 ( .A1(b_11_), .A2(n12721), .A3(a_22_), .ZN(n12720) );
  OR2_X1 U12727 ( .A1(n12574), .A2(n12572), .ZN(n12721) );
  NAND2_X1 U12728 ( .A1(n12572), .A2(n12574), .ZN(n12719) );
  NAND2_X1 U12729 ( .A1(n12722), .A2(n12723), .ZN(n12574) );
  NAND2_X1 U12730 ( .A1(n12571), .A2(n12724), .ZN(n12723) );
  OR2_X1 U12731 ( .A1(n12570), .A2(n12568), .ZN(n12724) );
  NOR2_X1 U12732 ( .A1(n7955), .A2(n7726), .ZN(n12571) );
  NAND2_X1 U12733 ( .A1(n12568), .A2(n12570), .ZN(n12722) );
  NAND2_X1 U12734 ( .A1(n12725), .A2(n12726), .ZN(n12570) );
  NAND3_X1 U12735 ( .A1(b_11_), .A2(n12727), .A3(a_24_), .ZN(n12726) );
  NAND2_X1 U12736 ( .A1(n12566), .A2(n12565), .ZN(n12727) );
  OR2_X1 U12737 ( .A1(n12565), .A2(n12566), .ZN(n12725) );
  AND2_X1 U12738 ( .A1(n12728), .A2(n12729), .ZN(n12566) );
  NAND2_X1 U12739 ( .A1(n12563), .A2(n12730), .ZN(n12729) );
  OR2_X1 U12740 ( .A1(n12562), .A2(n12561), .ZN(n12730) );
  NOR2_X1 U12741 ( .A1(n7952), .A2(n7726), .ZN(n12563) );
  NAND2_X1 U12742 ( .A1(n12561), .A2(n12562), .ZN(n12728) );
  NAND2_X1 U12743 ( .A1(n12558), .A2(n12731), .ZN(n12562) );
  NAND2_X1 U12744 ( .A1(n12557), .A2(n12559), .ZN(n12731) );
  NAND2_X1 U12745 ( .A1(n12732), .A2(n12733), .ZN(n12559) );
  NAND2_X1 U12746 ( .A1(a_26_), .A2(b_11_), .ZN(n12733) );
  INV_X1 U12747 ( .A(n12734), .ZN(n12732) );
  XNOR2_X1 U12748 ( .A(n12735), .B(n12736), .ZN(n12557) );
  NAND2_X1 U12749 ( .A1(n12737), .A2(n12738), .ZN(n12735) );
  NAND2_X1 U12750 ( .A1(a_26_), .A2(n12734), .ZN(n12558) );
  NAND2_X1 U12751 ( .A1(n12529), .A2(n12739), .ZN(n12734) );
  NAND2_X1 U12752 ( .A1(n12528), .A2(n12530), .ZN(n12739) );
  NAND2_X1 U12753 ( .A1(n12740), .A2(n12741), .ZN(n12530) );
  NAND2_X1 U12754 ( .A1(a_27_), .A2(b_11_), .ZN(n12741) );
  INV_X1 U12755 ( .A(n12742), .ZN(n12740) );
  XNOR2_X1 U12756 ( .A(n12743), .B(n12744), .ZN(n12528) );
  XOR2_X1 U12757 ( .A(n12745), .B(n12746), .Z(n12743) );
  NAND2_X1 U12758 ( .A1(a_28_), .A2(b_10_), .ZN(n12745) );
  NAND2_X1 U12759 ( .A1(a_27_), .A2(n12742), .ZN(n12529) );
  NAND2_X1 U12760 ( .A1(n12747), .A2(n12748), .ZN(n12742) );
  NAND3_X1 U12761 ( .A1(b_11_), .A2(n12749), .A3(a_28_), .ZN(n12748) );
  NAND2_X1 U12762 ( .A1(n12538), .A2(n12536), .ZN(n12749) );
  OR2_X1 U12763 ( .A1(n12536), .A2(n12538), .ZN(n12747) );
  AND2_X1 U12764 ( .A1(n12750), .A2(n12751), .ZN(n12538) );
  NAND2_X1 U12765 ( .A1(n12553), .A2(n12752), .ZN(n12751) );
  OR2_X1 U12766 ( .A1(n12554), .A2(n12555), .ZN(n12752) );
  NOR2_X1 U12767 ( .A1(n7460), .A2(n7726), .ZN(n12553) );
  INV_X1 U12768 ( .A(b_11_), .ZN(n7726) );
  NAND2_X1 U12769 ( .A1(n12555), .A2(n12554), .ZN(n12750) );
  NAND2_X1 U12770 ( .A1(n12753), .A2(n12754), .ZN(n12554) );
  NAND2_X1 U12771 ( .A1(b_10_), .A2(n12755), .ZN(n12754) );
  NAND2_X1 U12772 ( .A1(n7445), .A2(n12756), .ZN(n12755) );
  NAND2_X1 U12773 ( .A1(a_30_), .A2(n7755), .ZN(n12756) );
  NAND2_X1 U12774 ( .A1(b_9_), .A2(n12757), .ZN(n12753) );
  NAND2_X1 U12775 ( .A1(n7441), .A2(n12758), .ZN(n12757) );
  NAND2_X1 U12776 ( .A1(a_31_), .A2(n12551), .ZN(n12758) );
  AND3_X1 U12777 ( .A1(n7409), .A2(b_11_), .A3(b_10_), .ZN(n12555) );
  XNOR2_X1 U12778 ( .A(n12759), .B(n12760), .ZN(n12536) );
  XOR2_X1 U12779 ( .A(n12761), .B(n12762), .Z(n12759) );
  XNOR2_X1 U12780 ( .A(n12763), .B(n12764), .ZN(n12561) );
  NAND2_X1 U12781 ( .A1(n12765), .A2(n12766), .ZN(n12763) );
  XNOR2_X1 U12782 ( .A(n12767), .B(n12768), .ZN(n12565) );
  XOR2_X1 U12783 ( .A(n12769), .B(n12770), .Z(n12767) );
  XNOR2_X1 U12784 ( .A(n12771), .B(n12772), .ZN(n12568) );
  XNOR2_X1 U12785 ( .A(n12773), .B(n12774), .ZN(n12771) );
  NOR2_X1 U12786 ( .A1(n12551), .A2(n7954), .ZN(n12774) );
  XNOR2_X1 U12787 ( .A(n12775), .B(n12776), .ZN(n12572) );
  XNOR2_X1 U12788 ( .A(n12777), .B(n12778), .ZN(n12776) );
  XNOR2_X1 U12789 ( .A(n12779), .B(n12780), .ZN(n12577) );
  XNOR2_X1 U12790 ( .A(n12781), .B(n12782), .ZN(n12779) );
  NOR2_X1 U12791 ( .A1(n12551), .A2(n7568), .ZN(n12782) );
  XNOR2_X1 U12792 ( .A(n12783), .B(n12784), .ZN(n12502) );
  XNOR2_X1 U12793 ( .A(n12785), .B(n12786), .ZN(n12783) );
  NOR2_X1 U12794 ( .A1(n7578), .A2(n12551), .ZN(n12786) );
  XNOR2_X1 U12795 ( .A(n12787), .B(n12788), .ZN(n12588) );
  XNOR2_X1 U12796 ( .A(n12789), .B(n12790), .ZN(n12788) );
  XNOR2_X1 U12797 ( .A(n12791), .B(n12792), .ZN(n12485) );
  XOR2_X1 U12798 ( .A(n12793), .B(n12794), .Z(n12791) );
  NOR2_X1 U12799 ( .A1(n12551), .A2(n7645), .ZN(n12794) );
  XNOR2_X1 U12800 ( .A(n12795), .B(n12796), .ZN(n12476) );
  NAND2_X1 U12801 ( .A1(n12797), .A2(n12798), .ZN(n12795) );
  XNOR2_X1 U12802 ( .A(n12799), .B(n12800), .ZN(n12593) );
  NAND2_X1 U12803 ( .A1(n12801), .A2(n12802), .ZN(n12799) );
  XNOR2_X1 U12804 ( .A(n12803), .B(n12804), .ZN(n12465) );
  XNOR2_X1 U12805 ( .A(n12805), .B(n12806), .ZN(n12804) );
  XNOR2_X1 U12806 ( .A(n12807), .B(n12808), .ZN(n12459) );
  XOR2_X1 U12807 ( .A(n12809), .B(n12810), .Z(n12808) );
  NAND2_X1 U12808 ( .A1(a_13_), .A2(b_10_), .ZN(n12810) );
  INV_X1 U12809 ( .A(n7907), .ZN(n7721) );
  NAND2_X1 U12810 ( .A1(a_11_), .A2(b_11_), .ZN(n7907) );
  XOR2_X1 U12811 ( .A(n12811), .B(n12812), .Z(n12597) );
  NAND2_X1 U12812 ( .A1(n12813), .A2(n12814), .ZN(n12811) );
  XOR2_X1 U12813 ( .A(n12815), .B(n12816), .Z(n12601) );
  XNOR2_X1 U12814 ( .A(n7738), .B(n12817), .ZN(n12816) );
  XNOR2_X1 U12815 ( .A(n12818), .B(n12819), .ZN(n12437) );
  NAND2_X1 U12816 ( .A1(n12820), .A2(n12821), .ZN(n12818) );
  XOR2_X1 U12817 ( .A(n12822), .B(n12823), .Z(n12605) );
  NAND2_X1 U12818 ( .A1(n12824), .A2(n12825), .ZN(n12822) );
  XNOR2_X1 U12819 ( .A(n12826), .B(n12827), .ZN(n12609) );
  XNOR2_X1 U12820 ( .A(n12828), .B(n12829), .ZN(n12826) );
  XNOR2_X1 U12821 ( .A(n12830), .B(n12831), .ZN(n12612) );
  XNOR2_X1 U12822 ( .A(n12832), .B(n12833), .ZN(n12831) );
  XNOR2_X1 U12823 ( .A(n12834), .B(n12835), .ZN(n12617) );
  XOR2_X1 U12824 ( .A(n12836), .B(n12837), .Z(n12834) );
  XNOR2_X1 U12825 ( .A(n12838), .B(n12839), .ZN(n12620) );
  XNOR2_X1 U12826 ( .A(n12840), .B(n12841), .ZN(n12839) );
  XNOR2_X1 U12827 ( .A(n12842), .B(n12843), .ZN(n12625) );
  XNOR2_X1 U12828 ( .A(n12844), .B(n12845), .ZN(n12842) );
  XNOR2_X1 U12829 ( .A(n12846), .B(n12847), .ZN(n12629) );
  XNOR2_X1 U12830 ( .A(n12848), .B(n12849), .ZN(n12847) );
  XNOR2_X1 U12831 ( .A(n12850), .B(n12851), .ZN(n12634) );
  XNOR2_X1 U12832 ( .A(n12852), .B(n12853), .ZN(n12850) );
  NOR2_X1 U12833 ( .A1(n12551), .A2(n7872), .ZN(n12853) );
  XNOR2_X1 U12834 ( .A(n12854), .B(n12855), .ZN(n12633) );
  XNOR2_X1 U12835 ( .A(n12856), .B(n12857), .ZN(n12855) );
  NAND2_X1 U12836 ( .A1(b_10_), .A2(a_0_), .ZN(n12857) );
  NAND2_X1 U12837 ( .A1(n12858), .A2(n12859), .ZN(n7415) );
  NAND2_X1 U12838 ( .A1(n12860), .A2(n12861), .ZN(n12859) );
  NAND2_X1 U12839 ( .A1(n8109), .A2(n8108), .ZN(n12858) );
  NAND4_X1 U12840 ( .A1(n8109), .A2(n12860), .A3(n8108), .A4(n12861), .ZN(
        n7414) );
  NAND2_X1 U12841 ( .A1(n12862), .A2(n12863), .ZN(n8108) );
  NAND3_X1 U12842 ( .A1(a_0_), .A2(n12864), .A3(b_10_), .ZN(n12863) );
  NAND2_X1 U12843 ( .A1(n12856), .A2(n12854), .ZN(n12864) );
  OR2_X1 U12844 ( .A1(n12854), .A2(n12856), .ZN(n12862) );
  AND2_X1 U12845 ( .A1(n12865), .A2(n12866), .ZN(n12856) );
  NAND3_X1 U12846 ( .A1(b_10_), .A2(n12867), .A3(a_1_), .ZN(n12866) );
  NAND2_X1 U12847 ( .A1(n12852), .A2(n12851), .ZN(n12867) );
  OR2_X1 U12848 ( .A1(n12851), .A2(n12852), .ZN(n12865) );
  AND2_X1 U12849 ( .A1(n12868), .A2(n12869), .ZN(n12852) );
  NAND2_X1 U12850 ( .A1(n12849), .A2(n12870), .ZN(n12869) );
  OR2_X1 U12851 ( .A1(n12848), .A2(n12846), .ZN(n12870) );
  NOR2_X1 U12852 ( .A1(n7966), .A2(n12551), .ZN(n12849) );
  NAND2_X1 U12853 ( .A1(n12846), .A2(n12848), .ZN(n12868) );
  NAND2_X1 U12854 ( .A1(n12871), .A2(n12872), .ZN(n12848) );
  NAND2_X1 U12855 ( .A1(n12844), .A2(n12873), .ZN(n12872) );
  NAND2_X1 U12856 ( .A1(n12845), .A2(n12843), .ZN(n12873) );
  NOR2_X1 U12857 ( .A1(n7852), .A2(n12551), .ZN(n12844) );
  OR2_X1 U12858 ( .A1(n12843), .A2(n12845), .ZN(n12871) );
  AND2_X1 U12859 ( .A1(n12874), .A2(n12875), .ZN(n12845) );
  NAND2_X1 U12860 ( .A1(n12841), .A2(n12876), .ZN(n12875) );
  OR2_X1 U12861 ( .A1(n12840), .A2(n12838), .ZN(n12876) );
  NOR2_X1 U12862 ( .A1(n7836), .A2(n12551), .ZN(n12841) );
  NAND2_X1 U12863 ( .A1(n12838), .A2(n12840), .ZN(n12874) );
  NAND2_X1 U12864 ( .A1(n12877), .A2(n12878), .ZN(n12840) );
  NAND2_X1 U12865 ( .A1(n12837), .A2(n12879), .ZN(n12878) );
  OR2_X1 U12866 ( .A1(n12835), .A2(n12836), .ZN(n12879) );
  NOR2_X1 U12867 ( .A1(n7823), .A2(n12551), .ZN(n12837) );
  NAND2_X1 U12868 ( .A1(n12835), .A2(n12836), .ZN(n12877) );
  NAND2_X1 U12869 ( .A1(n12880), .A2(n12881), .ZN(n12836) );
  NAND2_X1 U12870 ( .A1(n12833), .A2(n12882), .ZN(n12881) );
  OR2_X1 U12871 ( .A1(n12832), .A2(n12830), .ZN(n12882) );
  NOR2_X1 U12872 ( .A1(n7807), .A2(n12551), .ZN(n12833) );
  NAND2_X1 U12873 ( .A1(n12830), .A2(n12832), .ZN(n12880) );
  NAND2_X1 U12874 ( .A1(n12883), .A2(n12884), .ZN(n12832) );
  NAND2_X1 U12875 ( .A1(n12829), .A2(n12885), .ZN(n12884) );
  NAND2_X1 U12876 ( .A1(n12828), .A2(n12827), .ZN(n12885) );
  NOR2_X1 U12877 ( .A1(n7787), .A2(n12551), .ZN(n12829) );
  OR2_X1 U12878 ( .A1(n12827), .A2(n12828), .ZN(n12883) );
  AND2_X1 U12879 ( .A1(n12824), .A2(n12886), .ZN(n12828) );
  NAND2_X1 U12880 ( .A1(n12823), .A2(n12825), .ZN(n12886) );
  NAND2_X1 U12881 ( .A1(n12887), .A2(n12888), .ZN(n12825) );
  NAND2_X1 U12882 ( .A1(a_8_), .A2(b_10_), .ZN(n12888) );
  INV_X1 U12883 ( .A(n12889), .ZN(n12887) );
  XOR2_X1 U12884 ( .A(n12890), .B(n12891), .Z(n12823) );
  XOR2_X1 U12885 ( .A(n12892), .B(n7750), .Z(n12890) );
  NAND2_X1 U12886 ( .A1(a_8_), .A2(n12889), .ZN(n12824) );
  NAND2_X1 U12887 ( .A1(n12820), .A2(n12893), .ZN(n12889) );
  NAND2_X1 U12888 ( .A1(n12819), .A2(n12821), .ZN(n12893) );
  NAND2_X1 U12889 ( .A1(n12894), .A2(n12895), .ZN(n12821) );
  NAND2_X1 U12890 ( .A1(a_9_), .A2(b_10_), .ZN(n12895) );
  INV_X1 U12891 ( .A(n12896), .ZN(n12894) );
  XNOR2_X1 U12892 ( .A(n12897), .B(n12898), .ZN(n12819) );
  XOR2_X1 U12893 ( .A(n12899), .B(n12900), .Z(n12898) );
  NAND2_X1 U12894 ( .A1(a_10_), .A2(b_9_), .ZN(n12900) );
  NAND2_X1 U12895 ( .A1(a_9_), .A2(n12896), .ZN(n12820) );
  NAND2_X1 U12896 ( .A1(n12901), .A2(n12902), .ZN(n12896) );
  NAND2_X1 U12897 ( .A1(n12815), .A2(n12903), .ZN(n12902) );
  OR2_X1 U12898 ( .A1(n12817), .A2(n7738), .ZN(n12903) );
  XNOR2_X1 U12899 ( .A(n12904), .B(n12905), .ZN(n12815) );
  XNOR2_X1 U12900 ( .A(n12906), .B(n12907), .ZN(n12904) );
  NOR2_X1 U12901 ( .A1(n7724), .A2(n7755), .ZN(n12907) );
  NAND2_X1 U12902 ( .A1(n7738), .A2(n12817), .ZN(n12901) );
  NAND2_X1 U12903 ( .A1(n12813), .A2(n12908), .ZN(n12817) );
  NAND2_X1 U12904 ( .A1(n12812), .A2(n12814), .ZN(n12908) );
  NAND2_X1 U12905 ( .A1(n12909), .A2(n12910), .ZN(n12814) );
  NAND2_X1 U12906 ( .A1(b_10_), .A2(a_11_), .ZN(n12910) );
  INV_X1 U12907 ( .A(n12911), .ZN(n12909) );
  XNOR2_X1 U12908 ( .A(n12912), .B(n12913), .ZN(n12812) );
  XOR2_X1 U12909 ( .A(n12914), .B(n12915), .Z(n12913) );
  NAND2_X1 U12910 ( .A1(a_12_), .A2(b_9_), .ZN(n12915) );
  NAND2_X1 U12911 ( .A1(a_11_), .A2(n12911), .ZN(n12813) );
  NAND2_X1 U12912 ( .A1(n12677), .A2(n12916), .ZN(n12911) );
  NAND2_X1 U12913 ( .A1(n12676), .A2(n12678), .ZN(n12916) );
  NAND2_X1 U12914 ( .A1(n12917), .A2(n12918), .ZN(n12678) );
  NAND2_X1 U12915 ( .A1(a_12_), .A2(b_10_), .ZN(n12918) );
  INV_X1 U12916 ( .A(n12919), .ZN(n12917) );
  XNOR2_X1 U12917 ( .A(n12920), .B(n12921), .ZN(n12676) );
  XOR2_X1 U12918 ( .A(n12922), .B(n12923), .Z(n12921) );
  NAND2_X1 U12919 ( .A1(a_13_), .A2(b_9_), .ZN(n12923) );
  NAND2_X1 U12920 ( .A1(a_12_), .A2(n12919), .ZN(n12677) );
  NAND2_X1 U12921 ( .A1(n12924), .A2(n12925), .ZN(n12919) );
  NAND3_X1 U12922 ( .A1(b_10_), .A2(n12926), .A3(a_13_), .ZN(n12925) );
  OR2_X1 U12923 ( .A1(n12809), .A2(n12807), .ZN(n12926) );
  NAND2_X1 U12924 ( .A1(n12807), .A2(n12809), .ZN(n12924) );
  NAND2_X1 U12925 ( .A1(n12927), .A2(n12928), .ZN(n12809) );
  NAND2_X1 U12926 ( .A1(n12806), .A2(n12929), .ZN(n12928) );
  OR2_X1 U12927 ( .A1(n12805), .A2(n12803), .ZN(n12929) );
  NOR2_X1 U12928 ( .A1(n7962), .A2(n12551), .ZN(n12806) );
  NAND2_X1 U12929 ( .A1(n12803), .A2(n12805), .ZN(n12927) );
  NAND2_X1 U12930 ( .A1(n12801), .A2(n12930), .ZN(n12805) );
  NAND2_X1 U12931 ( .A1(n12800), .A2(n12802), .ZN(n12930) );
  NAND2_X1 U12932 ( .A1(n12931), .A2(n12932), .ZN(n12802) );
  NAND2_X1 U12933 ( .A1(a_15_), .A2(b_10_), .ZN(n12932) );
  INV_X1 U12934 ( .A(n12933), .ZN(n12931) );
  XNOR2_X1 U12935 ( .A(n12934), .B(n12935), .ZN(n12800) );
  XOR2_X1 U12936 ( .A(n12936), .B(n12937), .Z(n12935) );
  NAND2_X1 U12937 ( .A1(a_16_), .A2(b_9_), .ZN(n12937) );
  NAND2_X1 U12938 ( .A1(a_15_), .A2(n12933), .ZN(n12801) );
  NAND2_X1 U12939 ( .A1(n12797), .A2(n12938), .ZN(n12933) );
  NAND2_X1 U12940 ( .A1(n12796), .A2(n12798), .ZN(n12938) );
  NAND2_X1 U12941 ( .A1(n12939), .A2(n12940), .ZN(n12798) );
  NAND2_X1 U12942 ( .A1(a_16_), .A2(b_10_), .ZN(n12940) );
  INV_X1 U12943 ( .A(n12941), .ZN(n12939) );
  XNOR2_X1 U12944 ( .A(n12942), .B(n12943), .ZN(n12796) );
  XNOR2_X1 U12945 ( .A(n12944), .B(n12945), .ZN(n12942) );
  NOR2_X1 U12946 ( .A1(n7755), .A2(n7645), .ZN(n12945) );
  NAND2_X1 U12947 ( .A1(a_16_), .A2(n12941), .ZN(n12797) );
  NAND2_X1 U12948 ( .A1(n12946), .A2(n12947), .ZN(n12941) );
  NAND3_X1 U12949 ( .A1(b_10_), .A2(n12948), .A3(a_17_), .ZN(n12947) );
  OR2_X1 U12950 ( .A1(n12792), .A2(n12793), .ZN(n12948) );
  NAND2_X1 U12951 ( .A1(n12792), .A2(n12793), .ZN(n12946) );
  NAND2_X1 U12952 ( .A1(n12949), .A2(n12950), .ZN(n12793) );
  NAND2_X1 U12953 ( .A1(n12790), .A2(n12951), .ZN(n12950) );
  OR2_X1 U12954 ( .A1(n12789), .A2(n12787), .ZN(n12951) );
  NOR2_X1 U12955 ( .A1(n7960), .A2(n12551), .ZN(n12790) );
  NAND2_X1 U12956 ( .A1(n12787), .A2(n12789), .ZN(n12949) );
  NAND2_X1 U12957 ( .A1(n12952), .A2(n12953), .ZN(n12789) );
  NAND2_X1 U12958 ( .A1(n12704), .A2(n12954), .ZN(n12953) );
  OR2_X1 U12959 ( .A1(n12703), .A2(n12701), .ZN(n12954) );
  NOR2_X1 U12960 ( .A1(n7958), .A2(n12551), .ZN(n12704) );
  NAND2_X1 U12961 ( .A1(n12701), .A2(n12703), .ZN(n12952) );
  NAND2_X1 U12962 ( .A1(n12955), .A2(n12956), .ZN(n12703) );
  NAND2_X1 U12963 ( .A1(n12712), .A2(n12957), .ZN(n12956) );
  OR2_X1 U12964 ( .A1(n12711), .A2(n12709), .ZN(n12957) );
  NOR2_X1 U12965 ( .A1(n7957), .A2(n12551), .ZN(n12712) );
  NAND2_X1 U12966 ( .A1(n12709), .A2(n12711), .ZN(n12955) );
  NAND2_X1 U12967 ( .A1(n12958), .A2(n12959), .ZN(n12711) );
  NAND3_X1 U12968 ( .A1(a_21_), .A2(n12960), .A3(b_10_), .ZN(n12959) );
  NAND2_X1 U12969 ( .A1(n12785), .A2(n12784), .ZN(n12960) );
  OR2_X1 U12970 ( .A1(n12784), .A2(n12785), .ZN(n12958) );
  AND2_X1 U12971 ( .A1(n12961), .A2(n12962), .ZN(n12785) );
  NAND3_X1 U12972 ( .A1(b_10_), .A2(n12963), .A3(a_22_), .ZN(n12962) );
  NAND2_X1 U12973 ( .A1(n12781), .A2(n12780), .ZN(n12963) );
  OR2_X1 U12974 ( .A1(n12780), .A2(n12781), .ZN(n12961) );
  AND2_X1 U12975 ( .A1(n12964), .A2(n12965), .ZN(n12781) );
  NAND2_X1 U12976 ( .A1(n12778), .A2(n12966), .ZN(n12965) );
  OR2_X1 U12977 ( .A1(n12775), .A2(n12777), .ZN(n12966) );
  NOR2_X1 U12978 ( .A1(n12551), .A2(n7955), .ZN(n12778) );
  NAND2_X1 U12979 ( .A1(n12775), .A2(n12777), .ZN(n12964) );
  NAND2_X1 U12980 ( .A1(n12967), .A2(n12968), .ZN(n12777) );
  NAND3_X1 U12981 ( .A1(b_10_), .A2(n12969), .A3(a_24_), .ZN(n12968) );
  NAND2_X1 U12982 ( .A1(n12773), .A2(n12772), .ZN(n12969) );
  OR2_X1 U12983 ( .A1(n12772), .A2(n12773), .ZN(n12967) );
  AND2_X1 U12984 ( .A1(n12970), .A2(n12971), .ZN(n12773) );
  NAND2_X1 U12985 ( .A1(n12770), .A2(n12972), .ZN(n12971) );
  OR2_X1 U12986 ( .A1(n12768), .A2(n12769), .ZN(n12972) );
  NOR2_X1 U12987 ( .A1(n12551), .A2(n7952), .ZN(n12770) );
  NAND2_X1 U12988 ( .A1(n12768), .A2(n12769), .ZN(n12970) );
  NAND2_X1 U12989 ( .A1(n12765), .A2(n12973), .ZN(n12769) );
  NAND2_X1 U12990 ( .A1(n12764), .A2(n12766), .ZN(n12973) );
  NAND2_X1 U12991 ( .A1(n12974), .A2(n12975), .ZN(n12766) );
  NAND2_X1 U12992 ( .A1(a_26_), .A2(b_10_), .ZN(n12975) );
  INV_X1 U12993 ( .A(n12976), .ZN(n12974) );
  XNOR2_X1 U12994 ( .A(n12977), .B(n12978), .ZN(n12764) );
  NAND2_X1 U12995 ( .A1(n12979), .A2(n12980), .ZN(n12977) );
  NAND2_X1 U12996 ( .A1(a_26_), .A2(n12976), .ZN(n12765) );
  NAND2_X1 U12997 ( .A1(n12737), .A2(n12981), .ZN(n12976) );
  NAND2_X1 U12998 ( .A1(n12736), .A2(n12738), .ZN(n12981) );
  NAND2_X1 U12999 ( .A1(n12982), .A2(n12983), .ZN(n12738) );
  NAND2_X1 U13000 ( .A1(a_27_), .A2(b_10_), .ZN(n12983) );
  INV_X1 U13001 ( .A(n12984), .ZN(n12982) );
  XNOR2_X1 U13002 ( .A(n12985), .B(n12986), .ZN(n12736) );
  XOR2_X1 U13003 ( .A(n12987), .B(n12988), .Z(n12985) );
  NAND2_X1 U13004 ( .A1(a_28_), .A2(b_9_), .ZN(n12987) );
  NAND2_X1 U13005 ( .A1(a_27_), .A2(n12984), .ZN(n12737) );
  NAND2_X1 U13006 ( .A1(n12989), .A2(n12990), .ZN(n12984) );
  NAND3_X1 U13007 ( .A1(b_10_), .A2(n12991), .A3(a_28_), .ZN(n12990) );
  NAND2_X1 U13008 ( .A1(n12746), .A2(n12744), .ZN(n12991) );
  OR2_X1 U13009 ( .A1(n12744), .A2(n12746), .ZN(n12989) );
  AND2_X1 U13010 ( .A1(n12992), .A2(n12993), .ZN(n12746) );
  NAND2_X1 U13011 ( .A1(n12760), .A2(n12994), .ZN(n12993) );
  OR2_X1 U13012 ( .A1(n12761), .A2(n12762), .ZN(n12994) );
  NOR2_X1 U13013 ( .A1(n12551), .A2(n7460), .ZN(n12760) );
  NAND2_X1 U13014 ( .A1(n12762), .A2(n12761), .ZN(n12992) );
  NAND2_X1 U13015 ( .A1(n12995), .A2(n12996), .ZN(n12761) );
  NAND2_X1 U13016 ( .A1(b_8_), .A2(n12997), .ZN(n12996) );
  NAND2_X1 U13017 ( .A1(n7441), .A2(n12998), .ZN(n12997) );
  NAND2_X1 U13018 ( .A1(a_31_), .A2(n7755), .ZN(n12998) );
  NAND2_X1 U13019 ( .A1(b_9_), .A2(n12999), .ZN(n12995) );
  NAND2_X1 U13020 ( .A1(n7445), .A2(n13000), .ZN(n12999) );
  NAND2_X1 U13021 ( .A1(a_30_), .A2(n13001), .ZN(n13000) );
  AND3_X1 U13022 ( .A1(b_10_), .A2(n7409), .A3(b_9_), .ZN(n12762) );
  XNOR2_X1 U13023 ( .A(n13002), .B(n13003), .ZN(n12744) );
  XOR2_X1 U13024 ( .A(n13004), .B(n13005), .Z(n13002) );
  XNOR2_X1 U13025 ( .A(n13006), .B(n13007), .ZN(n12768) );
  NAND2_X1 U13026 ( .A1(n13008), .A2(n13009), .ZN(n13006) );
  XNOR2_X1 U13027 ( .A(n13010), .B(n13011), .ZN(n12772) );
  XOR2_X1 U13028 ( .A(n13012), .B(n13013), .Z(n13010) );
  XNOR2_X1 U13029 ( .A(n13014), .B(n13015), .ZN(n12775) );
  XNOR2_X1 U13030 ( .A(n13016), .B(n13017), .ZN(n13014) );
  NOR2_X1 U13031 ( .A1(n7755), .A2(n7954), .ZN(n13017) );
  XOR2_X1 U13032 ( .A(n13018), .B(n13019), .Z(n12780) );
  XNOR2_X1 U13033 ( .A(n13020), .B(n13021), .ZN(n13019) );
  XNOR2_X1 U13034 ( .A(n13022), .B(n13023), .ZN(n12784) );
  XOR2_X1 U13035 ( .A(n13024), .B(n13025), .Z(n13022) );
  XOR2_X1 U13036 ( .A(n13026), .B(n13027), .Z(n12709) );
  XOR2_X1 U13037 ( .A(n13028), .B(n13029), .Z(n13026) );
  NOR2_X1 U13038 ( .A1(n7578), .A2(n7755), .ZN(n13029) );
  XOR2_X1 U13039 ( .A(n13030), .B(n13031), .Z(n12701) );
  XOR2_X1 U13040 ( .A(n13032), .B(n13033), .Z(n13030) );
  NOR2_X1 U13041 ( .A1(n7755), .A2(n7957), .ZN(n13033) );
  XNOR2_X1 U13042 ( .A(n13034), .B(n13035), .ZN(n12787) );
  XOR2_X1 U13043 ( .A(n13036), .B(n13037), .Z(n13035) );
  NAND2_X1 U13044 ( .A1(a_19_), .A2(b_9_), .ZN(n13037) );
  XNOR2_X1 U13045 ( .A(n13038), .B(n13039), .ZN(n12792) );
  XNOR2_X1 U13046 ( .A(n13040), .B(n13041), .ZN(n13038) );
  NOR2_X1 U13047 ( .A1(n7755), .A2(n7960), .ZN(n13041) );
  XOR2_X1 U13048 ( .A(n13042), .B(n13043), .Z(n12803) );
  XOR2_X1 U13049 ( .A(n13044), .B(n13045), .Z(n13042) );
  NOR2_X1 U13050 ( .A1(n7755), .A2(n7667), .ZN(n13045) );
  XNOR2_X1 U13051 ( .A(n13046), .B(n13047), .ZN(n12807) );
  XOR2_X1 U13052 ( .A(n13048), .B(n13049), .Z(n13047) );
  NAND2_X1 U13053 ( .A1(a_14_), .A2(b_9_), .ZN(n13049) );
  NOR2_X1 U13054 ( .A1(n8378), .A2(n12551), .ZN(n7738) );
  INV_X1 U13055 ( .A(b_10_), .ZN(n12551) );
  XNOR2_X1 U13056 ( .A(n13050), .B(n13051), .ZN(n12827) );
  XOR2_X1 U13057 ( .A(n13052), .B(n13053), .Z(n13050) );
  NOR2_X1 U13058 ( .A1(n7755), .A2(n8602), .ZN(n13053) );
  XNOR2_X1 U13059 ( .A(n13054), .B(n13055), .ZN(n12830) );
  XOR2_X1 U13060 ( .A(n13056), .B(n13057), .Z(n13055) );
  NAND2_X1 U13061 ( .A1(a_7_), .A2(b_9_), .ZN(n13057) );
  XNOR2_X1 U13062 ( .A(n13058), .B(n13059), .ZN(n12835) );
  XNOR2_X1 U13063 ( .A(n13060), .B(n13061), .ZN(n13058) );
  NOR2_X1 U13064 ( .A1(n7755), .A2(n7807), .ZN(n13061) );
  XOR2_X1 U13065 ( .A(n13062), .B(n13063), .Z(n12838) );
  XOR2_X1 U13066 ( .A(n13064), .B(n13065), .Z(n13062) );
  NOR2_X1 U13067 ( .A1(n7755), .A2(n7823), .ZN(n13065) );
  XNOR2_X1 U13068 ( .A(n13066), .B(n13067), .ZN(n12843) );
  XOR2_X1 U13069 ( .A(n13068), .B(n13069), .Z(n13066) );
  NOR2_X1 U13070 ( .A1(n7755), .A2(n7836), .ZN(n13069) );
  XOR2_X1 U13071 ( .A(n13070), .B(n13071), .Z(n12846) );
  XOR2_X1 U13072 ( .A(n13072), .B(n13073), .Z(n13070) );
  NOR2_X1 U13073 ( .A1(n7755), .A2(n7852), .ZN(n13073) );
  XNOR2_X1 U13074 ( .A(n13074), .B(n13075), .ZN(n12851) );
  XOR2_X1 U13075 ( .A(n13076), .B(n13077), .Z(n13074) );
  NOR2_X1 U13076 ( .A1(n7755), .A2(n7966), .ZN(n13077) );
  XNOR2_X1 U13077 ( .A(n13078), .B(n13079), .ZN(n12854) );
  XOR2_X1 U13078 ( .A(n13080), .B(n13081), .Z(n13078) );
  NAND2_X1 U13079 ( .A1(n13082), .A2(n13083), .ZN(n12860) );
  XOR2_X1 U13080 ( .A(n13084), .B(n13085), .Z(n8109) );
  XOR2_X1 U13081 ( .A(n13086), .B(n13087), .Z(n13084) );
  NAND2_X1 U13082 ( .A1(n13088), .A2(n12861), .ZN(n7420) );
  INV_X1 U13083 ( .A(n13089), .ZN(n12861) );
  XNOR2_X1 U13084 ( .A(n13090), .B(n13091), .ZN(n13088) );
  NAND2_X1 U13085 ( .A1(n13089), .A2(n13092), .ZN(n7419) );
  XOR2_X1 U13086 ( .A(n13090), .B(n13091), .Z(n13092) );
  NOR2_X1 U13087 ( .A1(n13083), .A2(n13082), .ZN(n13089) );
  AND2_X1 U13088 ( .A1(n13093), .A2(n13094), .ZN(n13082) );
  NAND2_X1 U13089 ( .A1(n13087), .A2(n13095), .ZN(n13094) );
  OR2_X1 U13090 ( .A1(n13085), .A2(n13086), .ZN(n13095) );
  NOR2_X1 U13091 ( .A1(n7755), .A2(n8197), .ZN(n13087) );
  NAND2_X1 U13092 ( .A1(n13085), .A2(n13086), .ZN(n13093) );
  NAND2_X1 U13093 ( .A1(n13096), .A2(n13097), .ZN(n13086) );
  NAND2_X1 U13094 ( .A1(n13081), .A2(n13098), .ZN(n13097) );
  OR2_X1 U13095 ( .A1(n13079), .A2(n13080), .ZN(n13098) );
  NOR2_X1 U13096 ( .A1(n7872), .A2(n7755), .ZN(n13081) );
  NAND2_X1 U13097 ( .A1(n13079), .A2(n13080), .ZN(n13096) );
  NAND2_X1 U13098 ( .A1(n13099), .A2(n13100), .ZN(n13080) );
  NAND3_X1 U13099 ( .A1(b_9_), .A2(n13101), .A3(a_2_), .ZN(n13100) );
  OR2_X1 U13100 ( .A1(n13075), .A2(n13076), .ZN(n13101) );
  NAND2_X1 U13101 ( .A1(n13075), .A2(n13076), .ZN(n13099) );
  NAND2_X1 U13102 ( .A1(n13102), .A2(n13103), .ZN(n13076) );
  NAND3_X1 U13103 ( .A1(b_9_), .A2(n13104), .A3(a_3_), .ZN(n13103) );
  OR2_X1 U13104 ( .A1(n13071), .A2(n13072), .ZN(n13104) );
  NAND2_X1 U13105 ( .A1(n13071), .A2(n13072), .ZN(n13102) );
  NAND2_X1 U13106 ( .A1(n13105), .A2(n13106), .ZN(n13072) );
  NAND3_X1 U13107 ( .A1(b_9_), .A2(n13107), .A3(a_4_), .ZN(n13106) );
  OR2_X1 U13108 ( .A1(n13067), .A2(n13068), .ZN(n13107) );
  NAND2_X1 U13109 ( .A1(n13067), .A2(n13068), .ZN(n13105) );
  NAND2_X1 U13110 ( .A1(n13108), .A2(n13109), .ZN(n13068) );
  NAND3_X1 U13111 ( .A1(b_9_), .A2(n13110), .A3(a_5_), .ZN(n13109) );
  OR2_X1 U13112 ( .A1(n13063), .A2(n13064), .ZN(n13110) );
  NAND2_X1 U13113 ( .A1(n13063), .A2(n13064), .ZN(n13108) );
  NAND2_X1 U13114 ( .A1(n13111), .A2(n13112), .ZN(n13064) );
  NAND3_X1 U13115 ( .A1(b_9_), .A2(n13113), .A3(a_6_), .ZN(n13112) );
  NAND2_X1 U13116 ( .A1(n13060), .A2(n13059), .ZN(n13113) );
  OR2_X1 U13117 ( .A1(n13059), .A2(n13060), .ZN(n13111) );
  AND2_X1 U13118 ( .A1(n13114), .A2(n13115), .ZN(n13060) );
  NAND3_X1 U13119 ( .A1(b_9_), .A2(n13116), .A3(a_7_), .ZN(n13115) );
  OR2_X1 U13120 ( .A1(n13054), .A2(n13056), .ZN(n13116) );
  NAND2_X1 U13121 ( .A1(n13054), .A2(n13056), .ZN(n13114) );
  NAND2_X1 U13122 ( .A1(n13117), .A2(n13118), .ZN(n13056) );
  NAND3_X1 U13123 ( .A1(b_9_), .A2(n13119), .A3(a_8_), .ZN(n13118) );
  OR2_X1 U13124 ( .A1(n13051), .A2(n13052), .ZN(n13119) );
  NAND2_X1 U13125 ( .A1(n13051), .A2(n13052), .ZN(n13117) );
  NAND2_X1 U13126 ( .A1(n13120), .A2(n13121), .ZN(n13052) );
  NAND2_X1 U13127 ( .A1(n12891), .A2(n13122), .ZN(n13121) );
  OR2_X1 U13128 ( .A1(n12892), .A2(n7750), .ZN(n13122) );
  XNOR2_X1 U13129 ( .A(n13123), .B(n13124), .ZN(n12891) );
  XNOR2_X1 U13130 ( .A(n13125), .B(n13126), .ZN(n13124) );
  NAND2_X1 U13131 ( .A1(n7750), .A2(n12892), .ZN(n13120) );
  NAND2_X1 U13132 ( .A1(n13127), .A2(n13128), .ZN(n12892) );
  NAND3_X1 U13133 ( .A1(b_9_), .A2(n13129), .A3(a_10_), .ZN(n13128) );
  OR2_X1 U13134 ( .A1(n12897), .A2(n12899), .ZN(n13129) );
  NAND2_X1 U13135 ( .A1(n12897), .A2(n12899), .ZN(n13127) );
  NAND2_X1 U13136 ( .A1(n13130), .A2(n13131), .ZN(n12899) );
  NAND3_X1 U13137 ( .A1(a_11_), .A2(n13132), .A3(b_9_), .ZN(n13131) );
  NAND2_X1 U13138 ( .A1(n12906), .A2(n12905), .ZN(n13132) );
  OR2_X1 U13139 ( .A1(n12905), .A2(n12906), .ZN(n13130) );
  AND2_X1 U13140 ( .A1(n13133), .A2(n13134), .ZN(n12906) );
  NAND3_X1 U13141 ( .A1(b_9_), .A2(n13135), .A3(a_12_), .ZN(n13134) );
  OR2_X1 U13142 ( .A1(n12912), .A2(n12914), .ZN(n13135) );
  NAND2_X1 U13143 ( .A1(n12912), .A2(n12914), .ZN(n13133) );
  NAND2_X1 U13144 ( .A1(n13136), .A2(n13137), .ZN(n12914) );
  NAND3_X1 U13145 ( .A1(b_9_), .A2(n13138), .A3(a_13_), .ZN(n13137) );
  OR2_X1 U13146 ( .A1(n12922), .A2(n12920), .ZN(n13138) );
  NAND2_X1 U13147 ( .A1(n12920), .A2(n12922), .ZN(n13136) );
  NAND2_X1 U13148 ( .A1(n13139), .A2(n13140), .ZN(n12922) );
  NAND3_X1 U13149 ( .A1(b_9_), .A2(n13141), .A3(a_14_), .ZN(n13140) );
  OR2_X1 U13150 ( .A1(n13046), .A2(n13048), .ZN(n13141) );
  NAND2_X1 U13151 ( .A1(n13046), .A2(n13048), .ZN(n13139) );
  NAND2_X1 U13152 ( .A1(n13142), .A2(n13143), .ZN(n13048) );
  NAND3_X1 U13153 ( .A1(b_9_), .A2(n13144), .A3(a_15_), .ZN(n13143) );
  OR2_X1 U13154 ( .A1(n13043), .A2(n13044), .ZN(n13144) );
  NAND2_X1 U13155 ( .A1(n13043), .A2(n13044), .ZN(n13142) );
  NAND2_X1 U13156 ( .A1(n13145), .A2(n13146), .ZN(n13044) );
  NAND3_X1 U13157 ( .A1(b_9_), .A2(n13147), .A3(a_16_), .ZN(n13146) );
  OR2_X1 U13158 ( .A1(n12936), .A2(n12934), .ZN(n13147) );
  NAND2_X1 U13159 ( .A1(n12934), .A2(n12936), .ZN(n13145) );
  NAND2_X1 U13160 ( .A1(n13148), .A2(n13149), .ZN(n12936) );
  NAND3_X1 U13161 ( .A1(b_9_), .A2(n13150), .A3(a_17_), .ZN(n13149) );
  NAND2_X1 U13162 ( .A1(n12944), .A2(n12943), .ZN(n13150) );
  OR2_X1 U13163 ( .A1(n12943), .A2(n12944), .ZN(n13148) );
  AND2_X1 U13164 ( .A1(n13151), .A2(n13152), .ZN(n12944) );
  NAND3_X1 U13165 ( .A1(b_9_), .A2(n13153), .A3(a_18_), .ZN(n13152) );
  NAND2_X1 U13166 ( .A1(n13040), .A2(n13039), .ZN(n13153) );
  OR2_X1 U13167 ( .A1(n13039), .A2(n13040), .ZN(n13151) );
  AND2_X1 U13168 ( .A1(n13154), .A2(n13155), .ZN(n13040) );
  NAND3_X1 U13169 ( .A1(b_9_), .A2(n13156), .A3(a_19_), .ZN(n13155) );
  OR2_X1 U13170 ( .A1(n13034), .A2(n13036), .ZN(n13156) );
  NAND2_X1 U13171 ( .A1(n13034), .A2(n13036), .ZN(n13154) );
  NAND2_X1 U13172 ( .A1(n13157), .A2(n13158), .ZN(n13036) );
  NAND3_X1 U13173 ( .A1(b_9_), .A2(n13159), .A3(a_20_), .ZN(n13158) );
  OR2_X1 U13174 ( .A1(n13031), .A2(n13032), .ZN(n13159) );
  NAND2_X1 U13175 ( .A1(n13031), .A2(n13032), .ZN(n13157) );
  NAND2_X1 U13176 ( .A1(n13160), .A2(n13161), .ZN(n13032) );
  NAND3_X1 U13177 ( .A1(a_21_), .A2(n13162), .A3(b_9_), .ZN(n13161) );
  OR2_X1 U13178 ( .A1(n13027), .A2(n13028), .ZN(n13162) );
  NAND2_X1 U13179 ( .A1(n13027), .A2(n13028), .ZN(n13160) );
  NAND2_X1 U13180 ( .A1(n13163), .A2(n13164), .ZN(n13028) );
  NAND2_X1 U13181 ( .A1(n13025), .A2(n13165), .ZN(n13164) );
  OR2_X1 U13182 ( .A1(n13023), .A2(n13024), .ZN(n13165) );
  NOR2_X1 U13183 ( .A1(n7568), .A2(n7755), .ZN(n13025) );
  NAND2_X1 U13184 ( .A1(n13023), .A2(n13024), .ZN(n13163) );
  NAND2_X1 U13185 ( .A1(n13166), .A2(n13167), .ZN(n13024) );
  NAND2_X1 U13186 ( .A1(n13021), .A2(n13168), .ZN(n13167) );
  OR2_X1 U13187 ( .A1(n13018), .A2(n13020), .ZN(n13168) );
  NOR2_X1 U13188 ( .A1(n7755), .A2(n7955), .ZN(n13021) );
  NAND2_X1 U13189 ( .A1(n13018), .A2(n13020), .ZN(n13166) );
  NAND2_X1 U13190 ( .A1(n13169), .A2(n13170), .ZN(n13020) );
  NAND3_X1 U13191 ( .A1(b_9_), .A2(n13171), .A3(a_24_), .ZN(n13170) );
  NAND2_X1 U13192 ( .A1(n13016), .A2(n13015), .ZN(n13171) );
  OR2_X1 U13193 ( .A1(n13015), .A2(n13016), .ZN(n13169) );
  AND2_X1 U13194 ( .A1(n13172), .A2(n13173), .ZN(n13016) );
  NAND2_X1 U13195 ( .A1(n13013), .A2(n13174), .ZN(n13173) );
  OR2_X1 U13196 ( .A1(n13011), .A2(n13012), .ZN(n13174) );
  NOR2_X1 U13197 ( .A1(n7755), .A2(n7952), .ZN(n13013) );
  NAND2_X1 U13198 ( .A1(n13011), .A2(n13012), .ZN(n13172) );
  NAND2_X1 U13199 ( .A1(n13008), .A2(n13175), .ZN(n13012) );
  NAND2_X1 U13200 ( .A1(n13007), .A2(n13009), .ZN(n13175) );
  NAND2_X1 U13201 ( .A1(n13176), .A2(n13177), .ZN(n13009) );
  NAND2_X1 U13202 ( .A1(a_26_), .A2(b_9_), .ZN(n13177) );
  INV_X1 U13203 ( .A(n13178), .ZN(n13176) );
  XNOR2_X1 U13204 ( .A(n13179), .B(n13180), .ZN(n13007) );
  NAND2_X1 U13205 ( .A1(n13181), .A2(n13182), .ZN(n13179) );
  NAND2_X1 U13206 ( .A1(a_26_), .A2(n13178), .ZN(n13008) );
  NAND2_X1 U13207 ( .A1(n12979), .A2(n13183), .ZN(n13178) );
  NAND2_X1 U13208 ( .A1(n12978), .A2(n12980), .ZN(n13183) );
  NAND2_X1 U13209 ( .A1(n13184), .A2(n13185), .ZN(n12980) );
  NAND2_X1 U13210 ( .A1(a_27_), .A2(b_9_), .ZN(n13185) );
  INV_X1 U13211 ( .A(n13186), .ZN(n13184) );
  XNOR2_X1 U13212 ( .A(n13187), .B(n13188), .ZN(n12978) );
  XOR2_X1 U13213 ( .A(n13189), .B(n13190), .Z(n13187) );
  NAND2_X1 U13214 ( .A1(a_28_), .A2(b_8_), .ZN(n13189) );
  NAND2_X1 U13215 ( .A1(a_27_), .A2(n13186), .ZN(n12979) );
  NAND2_X1 U13216 ( .A1(n13191), .A2(n13192), .ZN(n13186) );
  NAND3_X1 U13217 ( .A1(b_9_), .A2(n13193), .A3(a_28_), .ZN(n13192) );
  NAND2_X1 U13218 ( .A1(n12988), .A2(n12986), .ZN(n13193) );
  OR2_X1 U13219 ( .A1(n12986), .A2(n12988), .ZN(n13191) );
  AND2_X1 U13220 ( .A1(n13194), .A2(n13195), .ZN(n12988) );
  NAND2_X1 U13221 ( .A1(n13003), .A2(n13196), .ZN(n13195) );
  OR2_X1 U13222 ( .A1(n13004), .A2(n13005), .ZN(n13196) );
  NOR2_X1 U13223 ( .A1(n7755), .A2(n7460), .ZN(n13003) );
  INV_X1 U13224 ( .A(b_9_), .ZN(n7755) );
  NAND2_X1 U13225 ( .A1(n13005), .A2(n13004), .ZN(n13194) );
  NAND2_X1 U13226 ( .A1(n13197), .A2(n13198), .ZN(n13004) );
  NAND2_X1 U13227 ( .A1(b_7_), .A2(n13199), .ZN(n13198) );
  NAND2_X1 U13228 ( .A1(n7441), .A2(n13200), .ZN(n13199) );
  NAND2_X1 U13229 ( .A1(a_31_), .A2(n13001), .ZN(n13200) );
  NAND2_X1 U13230 ( .A1(b_8_), .A2(n13201), .ZN(n13197) );
  NAND2_X1 U13231 ( .A1(n7445), .A2(n13202), .ZN(n13201) );
  NAND2_X1 U13232 ( .A1(a_30_), .A2(n7789), .ZN(n13202) );
  AND3_X1 U13233 ( .A1(b_9_), .A2(n7409), .A3(b_8_), .ZN(n13005) );
  XNOR2_X1 U13234 ( .A(n13203), .B(n13204), .ZN(n12986) );
  XOR2_X1 U13235 ( .A(n13205), .B(n13206), .Z(n13203) );
  XNOR2_X1 U13236 ( .A(n13207), .B(n13208), .ZN(n13011) );
  NAND2_X1 U13237 ( .A1(n13209), .A2(n13210), .ZN(n13207) );
  XNOR2_X1 U13238 ( .A(n13211), .B(n13212), .ZN(n13015) );
  XOR2_X1 U13239 ( .A(n13213), .B(n13214), .Z(n13211) );
  XNOR2_X1 U13240 ( .A(n13215), .B(n13216), .ZN(n13018) );
  XNOR2_X1 U13241 ( .A(n13217), .B(n13218), .ZN(n13215) );
  NOR2_X1 U13242 ( .A1(n13001), .A2(n7954), .ZN(n13218) );
  XNOR2_X1 U13243 ( .A(n13219), .B(n13220), .ZN(n13023) );
  XOR2_X1 U13244 ( .A(n13221), .B(n13222), .Z(n13220) );
  NAND2_X1 U13245 ( .A1(b_8_), .A2(a_23_), .ZN(n13222) );
  XNOR2_X1 U13246 ( .A(n13223), .B(n13224), .ZN(n13027) );
  XNOR2_X1 U13247 ( .A(n13225), .B(n13226), .ZN(n13224) );
  XNOR2_X1 U13248 ( .A(n13227), .B(n13228), .ZN(n13031) );
  XNOR2_X1 U13249 ( .A(n13229), .B(n13230), .ZN(n13227) );
  XNOR2_X1 U13250 ( .A(n13231), .B(n13232), .ZN(n13034) );
  XNOR2_X1 U13251 ( .A(n13233), .B(n13234), .ZN(n13231) );
  XOR2_X1 U13252 ( .A(n13235), .B(n13236), .Z(n13039) );
  XNOR2_X1 U13253 ( .A(n13237), .B(n13238), .ZN(n13236) );
  XOR2_X1 U13254 ( .A(n13239), .B(n13240), .Z(n12943) );
  XOR2_X1 U13255 ( .A(n13241), .B(n13242), .Z(n13240) );
  NAND2_X1 U13256 ( .A1(a_18_), .A2(b_8_), .ZN(n13242) );
  XNOR2_X1 U13257 ( .A(n13243), .B(n13244), .ZN(n12934) );
  NAND2_X1 U13258 ( .A1(n13245), .A2(n13246), .ZN(n13243) );
  XNOR2_X1 U13259 ( .A(n13247), .B(n13248), .ZN(n13043) );
  NAND2_X1 U13260 ( .A1(n13249), .A2(n13250), .ZN(n13247) );
  XNOR2_X1 U13261 ( .A(n13251), .B(n13252), .ZN(n13046) );
  XNOR2_X1 U13262 ( .A(n13253), .B(n13254), .ZN(n13251) );
  XOR2_X1 U13263 ( .A(n13255), .B(n13256), .Z(n12920) );
  XOR2_X1 U13264 ( .A(n13257), .B(n13258), .Z(n13255) );
  NOR2_X1 U13265 ( .A1(n13001), .A2(n7962), .ZN(n13258) );
  XNOR2_X1 U13266 ( .A(n13259), .B(n13260), .ZN(n12912) );
  XNOR2_X1 U13267 ( .A(n13261), .B(n13262), .ZN(n13260) );
  XNOR2_X1 U13268 ( .A(n13263), .B(n13264), .ZN(n12905) );
  XOR2_X1 U13269 ( .A(n13265), .B(n13266), .Z(n13263) );
  XNOR2_X1 U13270 ( .A(n13267), .B(n13268), .ZN(n12897) );
  XNOR2_X1 U13271 ( .A(n13269), .B(n13270), .ZN(n13267) );
  INV_X1 U13272 ( .A(n7903), .ZN(n7750) );
  NAND2_X1 U13273 ( .A1(a_9_), .A2(b_9_), .ZN(n7903) );
  XNOR2_X1 U13274 ( .A(n13271), .B(n13272), .ZN(n13051) );
  XNOR2_X1 U13275 ( .A(n13273), .B(n13274), .ZN(n13271) );
  XOR2_X1 U13276 ( .A(n13275), .B(n13276), .Z(n13054) );
  XNOR2_X1 U13277 ( .A(n13277), .B(n7767), .ZN(n13276) );
  XNOR2_X1 U13278 ( .A(n13278), .B(n13279), .ZN(n13059) );
  XOR2_X1 U13279 ( .A(n13280), .B(n13281), .Z(n13278) );
  XNOR2_X1 U13280 ( .A(n13282), .B(n13283), .ZN(n13063) );
  XNOR2_X1 U13281 ( .A(n13284), .B(n13285), .ZN(n13283) );
  XNOR2_X1 U13282 ( .A(n13286), .B(n13287), .ZN(n13067) );
  XNOR2_X1 U13283 ( .A(n13288), .B(n13289), .ZN(n13286) );
  NOR2_X1 U13284 ( .A1(n13001), .A2(n7823), .ZN(n13289) );
  XNOR2_X1 U13285 ( .A(n13290), .B(n13291), .ZN(n13071) );
  XOR2_X1 U13286 ( .A(n13292), .B(n13293), .Z(n13291) );
  NAND2_X1 U13287 ( .A1(a_4_), .A2(b_8_), .ZN(n13293) );
  XOR2_X1 U13288 ( .A(n13294), .B(n13295), .Z(n13075) );
  XOR2_X1 U13289 ( .A(n13296), .B(n13297), .Z(n13294) );
  NOR2_X1 U13290 ( .A1(n13001), .A2(n7852), .ZN(n13297) );
  XOR2_X1 U13291 ( .A(n13298), .B(n13299), .Z(n13079) );
  XNOR2_X1 U13292 ( .A(n13300), .B(n13301), .ZN(n13299) );
  NAND2_X1 U13293 ( .A1(a_2_), .A2(b_8_), .ZN(n13301) );
  XOR2_X1 U13294 ( .A(n13302), .B(n13303), .Z(n13085) );
  XOR2_X1 U13295 ( .A(n13304), .B(n13305), .Z(n13302) );
  NOR2_X1 U13296 ( .A1(n13001), .A2(n7872), .ZN(n13305) );
  XNOR2_X1 U13297 ( .A(n13306), .B(n13307), .ZN(n13083) );
  XOR2_X1 U13298 ( .A(n13308), .B(n13309), .Z(n13306) );
  NOR2_X1 U13299 ( .A1(n8197), .A2(n13001), .ZN(n13309) );
  NAND2_X1 U13300 ( .A1(n13310), .A2(n13311), .ZN(n7425) );
  NAND2_X1 U13301 ( .A1(n13312), .A2(n13313), .ZN(n13311) );
  NAND2_X1 U13302 ( .A1(n13091), .A2(n13090), .ZN(n13310) );
  NAND4_X1 U13303 ( .A1(n13091), .A2(n13312), .A3(n13090), .A4(n13313), .ZN(
        n7424) );
  NAND2_X1 U13304 ( .A1(n13314), .A2(n13315), .ZN(n13090) );
  NAND3_X1 U13305 ( .A1(a_0_), .A2(n13316), .A3(b_8_), .ZN(n13315) );
  OR2_X1 U13306 ( .A1(n13308), .A2(n13307), .ZN(n13316) );
  NAND2_X1 U13307 ( .A1(n13307), .A2(n13308), .ZN(n13314) );
  NAND2_X1 U13308 ( .A1(n13317), .A2(n13318), .ZN(n13308) );
  NAND3_X1 U13309 ( .A1(b_8_), .A2(n13319), .A3(a_1_), .ZN(n13318) );
  OR2_X1 U13310 ( .A1(n13304), .A2(n13303), .ZN(n13319) );
  NAND2_X1 U13311 ( .A1(n13303), .A2(n13304), .ZN(n13317) );
  NAND2_X1 U13312 ( .A1(n13320), .A2(n13321), .ZN(n13304) );
  NAND3_X1 U13313 ( .A1(b_8_), .A2(n13322), .A3(a_2_), .ZN(n13321) );
  NAND2_X1 U13314 ( .A1(n13300), .A2(n13298), .ZN(n13322) );
  OR2_X1 U13315 ( .A1(n13298), .A2(n13300), .ZN(n13320) );
  AND2_X1 U13316 ( .A1(n13323), .A2(n13324), .ZN(n13300) );
  NAND3_X1 U13317 ( .A1(b_8_), .A2(n13325), .A3(a_3_), .ZN(n13324) );
  OR2_X1 U13318 ( .A1(n13296), .A2(n13295), .ZN(n13325) );
  NAND2_X1 U13319 ( .A1(n13295), .A2(n13296), .ZN(n13323) );
  NAND2_X1 U13320 ( .A1(n13326), .A2(n13327), .ZN(n13296) );
  NAND3_X1 U13321 ( .A1(b_8_), .A2(n13328), .A3(a_4_), .ZN(n13327) );
  OR2_X1 U13322 ( .A1(n13292), .A2(n13290), .ZN(n13328) );
  NAND2_X1 U13323 ( .A1(n13290), .A2(n13292), .ZN(n13326) );
  NAND2_X1 U13324 ( .A1(n13329), .A2(n13330), .ZN(n13292) );
  NAND3_X1 U13325 ( .A1(b_8_), .A2(n13331), .A3(a_5_), .ZN(n13330) );
  NAND2_X1 U13326 ( .A1(n13288), .A2(n13287), .ZN(n13331) );
  OR2_X1 U13327 ( .A1(n13287), .A2(n13288), .ZN(n13329) );
  AND2_X1 U13328 ( .A1(n13332), .A2(n13333), .ZN(n13288) );
  NAND2_X1 U13329 ( .A1(n13285), .A2(n13334), .ZN(n13333) );
  OR2_X1 U13330 ( .A1(n13284), .A2(n13282), .ZN(n13334) );
  NOR2_X1 U13331 ( .A1(n7807), .A2(n13001), .ZN(n13285) );
  NAND2_X1 U13332 ( .A1(n13282), .A2(n13284), .ZN(n13332) );
  NAND2_X1 U13333 ( .A1(n13335), .A2(n13336), .ZN(n13284) );
  NAND2_X1 U13334 ( .A1(n13281), .A2(n13337), .ZN(n13336) );
  NAND2_X1 U13335 ( .A1(n13279), .A2(n13280), .ZN(n13337) );
  NOR2_X1 U13336 ( .A1(n7787), .A2(n13001), .ZN(n13281) );
  OR2_X1 U13337 ( .A1(n13279), .A2(n13280), .ZN(n13335) );
  NAND2_X1 U13338 ( .A1(n13338), .A2(n13339), .ZN(n13280) );
  NAND2_X1 U13339 ( .A1(n13275), .A2(n13340), .ZN(n13339) );
  NAND2_X1 U13340 ( .A1(n7767), .A2(n13277), .ZN(n13340) );
  XNOR2_X1 U13341 ( .A(n13341), .B(n13342), .ZN(n13275) );
  XOR2_X1 U13342 ( .A(n13343), .B(n13344), .Z(n13341) );
  NOR2_X1 U13343 ( .A1(n7789), .A2(n7753), .ZN(n13344) );
  OR2_X1 U13344 ( .A1(n13277), .A2(n7767), .ZN(n13338) );
  NOR2_X1 U13345 ( .A1(n8602), .A2(n13001), .ZN(n7767) );
  NAND2_X1 U13346 ( .A1(n13345), .A2(n13346), .ZN(n13277) );
  NAND2_X1 U13347 ( .A1(n13274), .A2(n13347), .ZN(n13346) );
  NAND2_X1 U13348 ( .A1(n13273), .A2(n13272), .ZN(n13347) );
  NOR2_X1 U13349 ( .A1(n7753), .A2(n13001), .ZN(n13274) );
  OR2_X1 U13350 ( .A1(n13272), .A2(n13273), .ZN(n13345) );
  AND2_X1 U13351 ( .A1(n13348), .A2(n13349), .ZN(n13273) );
  NAND2_X1 U13352 ( .A1(n13126), .A2(n13350), .ZN(n13349) );
  OR2_X1 U13353 ( .A1(n13125), .A2(n13123), .ZN(n13350) );
  NOR2_X1 U13354 ( .A1(n8378), .A2(n13001), .ZN(n13126) );
  NAND2_X1 U13355 ( .A1(n13123), .A2(n13125), .ZN(n13348) );
  NAND2_X1 U13356 ( .A1(n13351), .A2(n13352), .ZN(n13125) );
  NAND2_X1 U13357 ( .A1(n13270), .A2(n13353), .ZN(n13352) );
  NAND2_X1 U13358 ( .A1(n13269), .A2(n13268), .ZN(n13353) );
  NOR2_X1 U13359 ( .A1(n13001), .A2(n7724), .ZN(n13270) );
  OR2_X1 U13360 ( .A1(n13268), .A2(n13269), .ZN(n13351) );
  AND2_X1 U13361 ( .A1(n13354), .A2(n13355), .ZN(n13269) );
  NAND2_X1 U13362 ( .A1(n13266), .A2(n13356), .ZN(n13355) );
  OR2_X1 U13363 ( .A1(n13264), .A2(n13265), .ZN(n13356) );
  NOR2_X1 U13364 ( .A1(n8585), .A2(n13001), .ZN(n13266) );
  NAND2_X1 U13365 ( .A1(n13264), .A2(n13265), .ZN(n13354) );
  NAND2_X1 U13366 ( .A1(n13357), .A2(n13358), .ZN(n13265) );
  NAND2_X1 U13367 ( .A1(n13262), .A2(n13359), .ZN(n13358) );
  OR2_X1 U13368 ( .A1(n13261), .A2(n13259), .ZN(n13359) );
  NOR2_X1 U13369 ( .A1(n7702), .A2(n13001), .ZN(n13262) );
  NAND2_X1 U13370 ( .A1(n13259), .A2(n13261), .ZN(n13357) );
  NAND2_X1 U13371 ( .A1(n13360), .A2(n13361), .ZN(n13261) );
  NAND3_X1 U13372 ( .A1(b_8_), .A2(n13362), .A3(a_14_), .ZN(n13361) );
  OR2_X1 U13373 ( .A1(n13256), .A2(n13257), .ZN(n13362) );
  NAND2_X1 U13374 ( .A1(n13256), .A2(n13257), .ZN(n13360) );
  NAND2_X1 U13375 ( .A1(n13363), .A2(n13364), .ZN(n13257) );
  NAND2_X1 U13376 ( .A1(n13254), .A2(n13365), .ZN(n13364) );
  NAND2_X1 U13377 ( .A1(n13253), .A2(n13252), .ZN(n13365) );
  NOR2_X1 U13378 ( .A1(n7667), .A2(n13001), .ZN(n13254) );
  OR2_X1 U13379 ( .A1(n13252), .A2(n13253), .ZN(n13363) );
  AND2_X1 U13380 ( .A1(n13249), .A2(n13366), .ZN(n13253) );
  NAND2_X1 U13381 ( .A1(n13248), .A2(n13250), .ZN(n13366) );
  NAND2_X1 U13382 ( .A1(n13367), .A2(n13368), .ZN(n13250) );
  NAND2_X1 U13383 ( .A1(a_16_), .A2(b_8_), .ZN(n13368) );
  INV_X1 U13384 ( .A(n13369), .ZN(n13367) );
  XNOR2_X1 U13385 ( .A(n13370), .B(n13371), .ZN(n13248) );
  XNOR2_X1 U13386 ( .A(n13372), .B(n13373), .ZN(n13370) );
  NOR2_X1 U13387 ( .A1(n7789), .A2(n7645), .ZN(n13373) );
  NAND2_X1 U13388 ( .A1(a_16_), .A2(n13369), .ZN(n13249) );
  NAND2_X1 U13389 ( .A1(n13245), .A2(n13374), .ZN(n13369) );
  NAND2_X1 U13390 ( .A1(n13244), .A2(n13246), .ZN(n13374) );
  NAND2_X1 U13391 ( .A1(n13375), .A2(n13376), .ZN(n13246) );
  NAND2_X1 U13392 ( .A1(a_17_), .A2(b_8_), .ZN(n13376) );
  INV_X1 U13393 ( .A(n13377), .ZN(n13375) );
  XNOR2_X1 U13394 ( .A(n13378), .B(n13379), .ZN(n13244) );
  XOR2_X1 U13395 ( .A(n13380), .B(n13381), .Z(n13379) );
  NAND2_X1 U13396 ( .A1(a_18_), .A2(b_7_), .ZN(n13381) );
  NAND2_X1 U13397 ( .A1(a_17_), .A2(n13377), .ZN(n13245) );
  NAND2_X1 U13398 ( .A1(n13382), .A2(n13383), .ZN(n13377) );
  NAND3_X1 U13399 ( .A1(b_8_), .A2(n13384), .A3(a_18_), .ZN(n13383) );
  OR2_X1 U13400 ( .A1(n13239), .A2(n13241), .ZN(n13384) );
  NAND2_X1 U13401 ( .A1(n13239), .A2(n13241), .ZN(n13382) );
  NAND2_X1 U13402 ( .A1(n13385), .A2(n13386), .ZN(n13241) );
  NAND2_X1 U13403 ( .A1(n13238), .A2(n13387), .ZN(n13386) );
  OR2_X1 U13404 ( .A1(n13235), .A2(n13237), .ZN(n13387) );
  NOR2_X1 U13405 ( .A1(n7958), .A2(n13001), .ZN(n13238) );
  NAND2_X1 U13406 ( .A1(n13235), .A2(n13237), .ZN(n13385) );
  NAND2_X1 U13407 ( .A1(n13388), .A2(n13389), .ZN(n13237) );
  NAND2_X1 U13408 ( .A1(n13233), .A2(n13390), .ZN(n13389) );
  NAND2_X1 U13409 ( .A1(n13234), .A2(n13232), .ZN(n13390) );
  NOR2_X1 U13410 ( .A1(n7957), .A2(n13001), .ZN(n13233) );
  OR2_X1 U13411 ( .A1(n13232), .A2(n13234), .ZN(n13388) );
  AND2_X1 U13412 ( .A1(n13391), .A2(n13392), .ZN(n13234) );
  NAND2_X1 U13413 ( .A1(n13230), .A2(n13393), .ZN(n13392) );
  NAND2_X1 U13414 ( .A1(n13229), .A2(n13228), .ZN(n13393) );
  NOR2_X1 U13415 ( .A1(n13001), .A2(n7578), .ZN(n13230) );
  OR2_X1 U13416 ( .A1(n13228), .A2(n13229), .ZN(n13391) );
  AND2_X1 U13417 ( .A1(n13394), .A2(n13395), .ZN(n13229) );
  NAND2_X1 U13418 ( .A1(n13226), .A2(n13396), .ZN(n13395) );
  OR2_X1 U13419 ( .A1(n13225), .A2(n13223), .ZN(n13396) );
  NOR2_X1 U13420 ( .A1(n7568), .A2(n13001), .ZN(n13226) );
  NAND2_X1 U13421 ( .A1(n13223), .A2(n13225), .ZN(n13394) );
  NAND2_X1 U13422 ( .A1(n13397), .A2(n13398), .ZN(n13225) );
  NAND3_X1 U13423 ( .A1(a_23_), .A2(n13399), .A3(b_8_), .ZN(n13398) );
  OR2_X1 U13424 ( .A1(n13221), .A2(n13219), .ZN(n13399) );
  NAND2_X1 U13425 ( .A1(n13219), .A2(n13221), .ZN(n13397) );
  NAND2_X1 U13426 ( .A1(n13400), .A2(n13401), .ZN(n13221) );
  NAND3_X1 U13427 ( .A1(b_8_), .A2(n13402), .A3(a_24_), .ZN(n13401) );
  NAND2_X1 U13428 ( .A1(n13217), .A2(n13216), .ZN(n13402) );
  OR2_X1 U13429 ( .A1(n13216), .A2(n13217), .ZN(n13400) );
  AND2_X1 U13430 ( .A1(n13403), .A2(n13404), .ZN(n13217) );
  NAND2_X1 U13431 ( .A1(n13214), .A2(n13405), .ZN(n13404) );
  OR2_X1 U13432 ( .A1(n13212), .A2(n13213), .ZN(n13405) );
  NOR2_X1 U13433 ( .A1(n13001), .A2(n7952), .ZN(n13214) );
  NAND2_X1 U13434 ( .A1(n13212), .A2(n13213), .ZN(n13403) );
  NAND2_X1 U13435 ( .A1(n13209), .A2(n13406), .ZN(n13213) );
  NAND2_X1 U13436 ( .A1(n13208), .A2(n13210), .ZN(n13406) );
  NAND2_X1 U13437 ( .A1(n13407), .A2(n13408), .ZN(n13210) );
  NAND2_X1 U13438 ( .A1(a_26_), .A2(b_8_), .ZN(n13408) );
  INV_X1 U13439 ( .A(n13409), .ZN(n13407) );
  XNOR2_X1 U13440 ( .A(n13410), .B(n13411), .ZN(n13208) );
  NAND2_X1 U13441 ( .A1(n13412), .A2(n13413), .ZN(n13410) );
  NAND2_X1 U13442 ( .A1(a_26_), .A2(n13409), .ZN(n13209) );
  NAND2_X1 U13443 ( .A1(n13181), .A2(n13414), .ZN(n13409) );
  NAND2_X1 U13444 ( .A1(n13180), .A2(n13182), .ZN(n13414) );
  NAND2_X1 U13445 ( .A1(n13415), .A2(n13416), .ZN(n13182) );
  NAND2_X1 U13446 ( .A1(a_27_), .A2(b_8_), .ZN(n13416) );
  INV_X1 U13447 ( .A(n13417), .ZN(n13415) );
  XNOR2_X1 U13448 ( .A(n13418), .B(n13419), .ZN(n13180) );
  XOR2_X1 U13449 ( .A(n13420), .B(n13421), .Z(n13418) );
  NAND2_X1 U13450 ( .A1(b_7_), .A2(a_28_), .ZN(n13420) );
  NAND2_X1 U13451 ( .A1(a_27_), .A2(n13417), .ZN(n13181) );
  NAND2_X1 U13452 ( .A1(n13422), .A2(n13423), .ZN(n13417) );
  NAND3_X1 U13453 ( .A1(b_8_), .A2(n13424), .A3(a_28_), .ZN(n13423) );
  NAND2_X1 U13454 ( .A1(n13190), .A2(n13188), .ZN(n13424) );
  OR2_X1 U13455 ( .A1(n13188), .A2(n13190), .ZN(n13422) );
  AND2_X1 U13456 ( .A1(n13425), .A2(n13426), .ZN(n13190) );
  NAND2_X1 U13457 ( .A1(n13204), .A2(n13427), .ZN(n13426) );
  OR2_X1 U13458 ( .A1(n13205), .A2(n13206), .ZN(n13427) );
  NOR2_X1 U13459 ( .A1(n13001), .A2(n7460), .ZN(n13204) );
  INV_X1 U13460 ( .A(b_8_), .ZN(n13001) );
  NAND2_X1 U13461 ( .A1(n13206), .A2(n13205), .ZN(n13425) );
  NAND2_X1 U13462 ( .A1(n13428), .A2(n13429), .ZN(n13205) );
  NAND2_X1 U13463 ( .A1(b_6_), .A2(n13430), .ZN(n13429) );
  NAND2_X1 U13464 ( .A1(n7441), .A2(n13431), .ZN(n13430) );
  NAND2_X1 U13465 ( .A1(a_31_), .A2(n7789), .ZN(n13431) );
  NAND2_X1 U13466 ( .A1(b_7_), .A2(n13432), .ZN(n13428) );
  NAND2_X1 U13467 ( .A1(n7445), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U13468 ( .A1(a_30_), .A2(n7963), .ZN(n13433) );
  AND3_X1 U13469 ( .A1(b_8_), .A2(n7409), .A3(b_7_), .ZN(n13206) );
  XNOR2_X1 U13470 ( .A(n13434), .B(n13435), .ZN(n13188) );
  XOR2_X1 U13471 ( .A(n13436), .B(n13437), .Z(n13434) );
  XNOR2_X1 U13472 ( .A(n13438), .B(n13439), .ZN(n13212) );
  NAND2_X1 U13473 ( .A1(n13440), .A2(n13441), .ZN(n13438) );
  XNOR2_X1 U13474 ( .A(n13442), .B(n13443), .ZN(n13216) );
  XOR2_X1 U13475 ( .A(n13444), .B(n13445), .Z(n13442) );
  XOR2_X1 U13476 ( .A(n13446), .B(n13447), .Z(n13219) );
  XOR2_X1 U13477 ( .A(n13448), .B(n13449), .Z(n13446) );
  XOR2_X1 U13478 ( .A(n13450), .B(n13451), .Z(n13223) );
  XOR2_X1 U13479 ( .A(n13452), .B(n13453), .Z(n13450) );
  NOR2_X1 U13480 ( .A1(n7955), .A2(n7789), .ZN(n13453) );
  XOR2_X1 U13481 ( .A(n13454), .B(n13455), .Z(n13228) );
  NAND2_X1 U13482 ( .A1(n13456), .A2(n13457), .ZN(n13454) );
  XNOR2_X1 U13483 ( .A(n13458), .B(n13459), .ZN(n13232) );
  XOR2_X1 U13484 ( .A(n13460), .B(n13461), .Z(n13458) );
  NOR2_X1 U13485 ( .A1(n7578), .A2(n7789), .ZN(n13461) );
  XNOR2_X1 U13486 ( .A(n13462), .B(n13463), .ZN(n13235) );
  XNOR2_X1 U13487 ( .A(n13464), .B(n13465), .ZN(n13462) );
  NOR2_X1 U13488 ( .A1(n7789), .A2(n7957), .ZN(n13465) );
  XNOR2_X1 U13489 ( .A(n13466), .B(n13467), .ZN(n13239) );
  XOR2_X1 U13490 ( .A(n13468), .B(n13469), .Z(n13467) );
  NAND2_X1 U13491 ( .A1(a_19_), .A2(b_7_), .ZN(n13469) );
  XOR2_X1 U13492 ( .A(n13470), .B(n13471), .Z(n13252) );
  XOR2_X1 U13493 ( .A(n13472), .B(n13473), .Z(n13471) );
  NAND2_X1 U13494 ( .A1(a_16_), .A2(b_7_), .ZN(n13473) );
  XNOR2_X1 U13495 ( .A(n13474), .B(n13475), .ZN(n13256) );
  XNOR2_X1 U13496 ( .A(n13476), .B(n13477), .ZN(n13474) );
  NOR2_X1 U13497 ( .A1(n7789), .A2(n7667), .ZN(n13477) );
  XOR2_X1 U13498 ( .A(n13478), .B(n13479), .Z(n13259) );
  XOR2_X1 U13499 ( .A(n13480), .B(n13481), .Z(n13478) );
  NOR2_X1 U13500 ( .A1(n7789), .A2(n7962), .ZN(n13481) );
  XNOR2_X1 U13501 ( .A(n13482), .B(n13483), .ZN(n13264) );
  XOR2_X1 U13502 ( .A(n13484), .B(n13485), .Z(n13483) );
  NAND2_X1 U13503 ( .A1(a_13_), .A2(b_7_), .ZN(n13485) );
  XNOR2_X1 U13504 ( .A(n13486), .B(n13487), .ZN(n13268) );
  XOR2_X1 U13505 ( .A(n13488), .B(n13489), .Z(n13486) );
  NOR2_X1 U13506 ( .A1(n7789), .A2(n8585), .ZN(n13489) );
  XOR2_X1 U13507 ( .A(n13490), .B(n13491), .Z(n13123) );
  XOR2_X1 U13508 ( .A(n13492), .B(n13493), .Z(n13490) );
  NOR2_X1 U13509 ( .A1(n7724), .A2(n7789), .ZN(n13493) );
  XNOR2_X1 U13510 ( .A(n13494), .B(n13495), .ZN(n13272) );
  XOR2_X1 U13511 ( .A(n13496), .B(n13497), .Z(n13494) );
  NOR2_X1 U13512 ( .A1(n7789), .A2(n8378), .ZN(n13497) );
  XNOR2_X1 U13513 ( .A(n13498), .B(n13499), .ZN(n13279) );
  XOR2_X1 U13514 ( .A(n13500), .B(n13501), .Z(n13498) );
  NOR2_X1 U13515 ( .A1(n7789), .A2(n8602), .ZN(n13501) );
  XOR2_X1 U13516 ( .A(n13502), .B(n13503), .Z(n13282) );
  XOR2_X1 U13517 ( .A(n13504), .B(n7784), .Z(n13502) );
  XNOR2_X1 U13518 ( .A(n13505), .B(n13506), .ZN(n13287) );
  XOR2_X1 U13519 ( .A(n13507), .B(n13508), .Z(n13505) );
  NOR2_X1 U13520 ( .A1(n7789), .A2(n7807), .ZN(n13508) );
  XOR2_X1 U13521 ( .A(n13509), .B(n13510), .Z(n13290) );
  XOR2_X1 U13522 ( .A(n13511), .B(n13512), .Z(n13509) );
  NOR2_X1 U13523 ( .A1(n7789), .A2(n7823), .ZN(n13512) );
  XOR2_X1 U13524 ( .A(n13513), .B(n13514), .Z(n13295) );
  XOR2_X1 U13525 ( .A(n13515), .B(n13516), .Z(n13513) );
  NOR2_X1 U13526 ( .A1(n7789), .A2(n7836), .ZN(n13516) );
  XNOR2_X1 U13527 ( .A(n13517), .B(n13518), .ZN(n13298) );
  XOR2_X1 U13528 ( .A(n13519), .B(n13520), .Z(n13517) );
  NOR2_X1 U13529 ( .A1(n7789), .A2(n7852), .ZN(n13520) );
  XOR2_X1 U13530 ( .A(n13521), .B(n13522), .Z(n13303) );
  XOR2_X1 U13531 ( .A(n13523), .B(n13524), .Z(n13521) );
  NOR2_X1 U13532 ( .A1(n7789), .A2(n7966), .ZN(n13524) );
  XOR2_X1 U13533 ( .A(n13525), .B(n13526), .Z(n13307) );
  XOR2_X1 U13534 ( .A(n13527), .B(n13528), .Z(n13525) );
  NAND2_X1 U13535 ( .A1(n13529), .A2(n13530), .ZN(n13312) );
  XOR2_X1 U13536 ( .A(n13531), .B(n13532), .Z(n13091) );
  XOR2_X1 U13537 ( .A(n13533), .B(n13534), .Z(n13531) );
  NAND2_X1 U13538 ( .A1(n13535), .A2(n13313), .ZN(n7430) );
  INV_X1 U13539 ( .A(n13536), .ZN(n13313) );
  XNOR2_X1 U13540 ( .A(n13537), .B(n13538), .ZN(n13535) );
  NAND2_X1 U13541 ( .A1(n13536), .A2(n13539), .ZN(n7429) );
  XOR2_X1 U13542 ( .A(n13537), .B(n13538), .Z(n13539) );
  NOR2_X1 U13543 ( .A1(n13530), .A2(n13529), .ZN(n13536) );
  AND2_X1 U13544 ( .A1(n13540), .A2(n13541), .ZN(n13529) );
  NAND2_X1 U13545 ( .A1(n13534), .A2(n13542), .ZN(n13541) );
  OR2_X1 U13546 ( .A1(n13532), .A2(n13533), .ZN(n13542) );
  NOR2_X1 U13547 ( .A1(n7789), .A2(n8197), .ZN(n13534) );
  NAND2_X1 U13548 ( .A1(n13532), .A2(n13533), .ZN(n13540) );
  NAND2_X1 U13549 ( .A1(n13543), .A2(n13544), .ZN(n13533) );
  NAND2_X1 U13550 ( .A1(n13528), .A2(n13545), .ZN(n13544) );
  OR2_X1 U13551 ( .A1(n13526), .A2(n13527), .ZN(n13545) );
  NOR2_X1 U13552 ( .A1(n7872), .A2(n7789), .ZN(n13528) );
  NAND2_X1 U13553 ( .A1(n13526), .A2(n13527), .ZN(n13543) );
  NAND2_X1 U13554 ( .A1(n13546), .A2(n13547), .ZN(n13527) );
  NAND3_X1 U13555 ( .A1(b_7_), .A2(n13548), .A3(a_2_), .ZN(n13547) );
  OR2_X1 U13556 ( .A1(n13522), .A2(n13523), .ZN(n13548) );
  NAND2_X1 U13557 ( .A1(n13522), .A2(n13523), .ZN(n13546) );
  NAND2_X1 U13558 ( .A1(n13549), .A2(n13550), .ZN(n13523) );
  NAND3_X1 U13559 ( .A1(b_7_), .A2(n13551), .A3(a_3_), .ZN(n13550) );
  OR2_X1 U13560 ( .A1(n13518), .A2(n13519), .ZN(n13551) );
  NAND2_X1 U13561 ( .A1(n13518), .A2(n13519), .ZN(n13549) );
  NAND2_X1 U13562 ( .A1(n13552), .A2(n13553), .ZN(n13519) );
  NAND3_X1 U13563 ( .A1(b_7_), .A2(n13554), .A3(a_4_), .ZN(n13553) );
  OR2_X1 U13564 ( .A1(n13514), .A2(n13515), .ZN(n13554) );
  NAND2_X1 U13565 ( .A1(n13514), .A2(n13515), .ZN(n13552) );
  NAND2_X1 U13566 ( .A1(n13555), .A2(n13556), .ZN(n13515) );
  NAND3_X1 U13567 ( .A1(b_7_), .A2(n13557), .A3(a_5_), .ZN(n13556) );
  OR2_X1 U13568 ( .A1(n13510), .A2(n13511), .ZN(n13557) );
  NAND2_X1 U13569 ( .A1(n13510), .A2(n13511), .ZN(n13555) );
  NAND2_X1 U13570 ( .A1(n13558), .A2(n13559), .ZN(n13511) );
  NAND3_X1 U13571 ( .A1(b_7_), .A2(n13560), .A3(a_6_), .ZN(n13559) );
  OR2_X1 U13572 ( .A1(n13506), .A2(n13507), .ZN(n13560) );
  NAND2_X1 U13573 ( .A1(n13506), .A2(n13507), .ZN(n13558) );
  NAND2_X1 U13574 ( .A1(n13561), .A2(n13562), .ZN(n13507) );
  NAND2_X1 U13575 ( .A1(n13503), .A2(n13563), .ZN(n13562) );
  OR2_X1 U13576 ( .A1(n13504), .A2(n7784), .ZN(n13563) );
  XNOR2_X1 U13577 ( .A(n13564), .B(n13565), .ZN(n13503) );
  XOR2_X1 U13578 ( .A(n13566), .B(n13567), .Z(n13565) );
  NAND2_X1 U13579 ( .A1(a_8_), .A2(b_6_), .ZN(n13567) );
  NAND2_X1 U13580 ( .A1(n7784), .A2(n13504), .ZN(n13561) );
  NAND2_X1 U13581 ( .A1(n13568), .A2(n13569), .ZN(n13504) );
  NAND3_X1 U13582 ( .A1(b_7_), .A2(n13570), .A3(a_8_), .ZN(n13569) );
  OR2_X1 U13583 ( .A1(n13499), .A2(n13500), .ZN(n13570) );
  NAND2_X1 U13584 ( .A1(n13499), .A2(n13500), .ZN(n13568) );
  NAND2_X1 U13585 ( .A1(n13571), .A2(n13572), .ZN(n13500) );
  NAND3_X1 U13586 ( .A1(b_7_), .A2(n13573), .A3(a_9_), .ZN(n13572) );
  OR2_X1 U13587 ( .A1(n13342), .A2(n13343), .ZN(n13573) );
  NAND2_X1 U13588 ( .A1(n13342), .A2(n13343), .ZN(n13571) );
  NAND2_X1 U13589 ( .A1(n13574), .A2(n13575), .ZN(n13343) );
  NAND3_X1 U13590 ( .A1(b_7_), .A2(n13576), .A3(a_10_), .ZN(n13575) );
  OR2_X1 U13591 ( .A1(n13495), .A2(n13496), .ZN(n13576) );
  NAND2_X1 U13592 ( .A1(n13495), .A2(n13496), .ZN(n13574) );
  NAND2_X1 U13593 ( .A1(n13577), .A2(n13578), .ZN(n13496) );
  NAND3_X1 U13594 ( .A1(a_11_), .A2(n13579), .A3(b_7_), .ZN(n13578) );
  OR2_X1 U13595 ( .A1(n13491), .A2(n13492), .ZN(n13579) );
  NAND2_X1 U13596 ( .A1(n13491), .A2(n13492), .ZN(n13577) );
  NAND2_X1 U13597 ( .A1(n13580), .A2(n13581), .ZN(n13492) );
  NAND3_X1 U13598 ( .A1(b_7_), .A2(n13582), .A3(a_12_), .ZN(n13581) );
  OR2_X1 U13599 ( .A1(n13487), .A2(n13488), .ZN(n13582) );
  NAND2_X1 U13600 ( .A1(n13487), .A2(n13488), .ZN(n13580) );
  NAND2_X1 U13601 ( .A1(n13583), .A2(n13584), .ZN(n13488) );
  NAND3_X1 U13602 ( .A1(b_7_), .A2(n13585), .A3(a_13_), .ZN(n13584) );
  OR2_X1 U13603 ( .A1(n13484), .A2(n13482), .ZN(n13585) );
  NAND2_X1 U13604 ( .A1(n13482), .A2(n13484), .ZN(n13583) );
  NAND2_X1 U13605 ( .A1(n13586), .A2(n13587), .ZN(n13484) );
  NAND3_X1 U13606 ( .A1(b_7_), .A2(n13588), .A3(a_14_), .ZN(n13587) );
  OR2_X1 U13607 ( .A1(n13479), .A2(n13480), .ZN(n13588) );
  NAND2_X1 U13608 ( .A1(n13479), .A2(n13480), .ZN(n13586) );
  NAND2_X1 U13609 ( .A1(n13589), .A2(n13590), .ZN(n13480) );
  NAND3_X1 U13610 ( .A1(b_7_), .A2(n13591), .A3(a_15_), .ZN(n13590) );
  NAND2_X1 U13611 ( .A1(n13476), .A2(n13475), .ZN(n13591) );
  OR2_X1 U13612 ( .A1(n13475), .A2(n13476), .ZN(n13589) );
  AND2_X1 U13613 ( .A1(n13592), .A2(n13593), .ZN(n13476) );
  NAND3_X1 U13614 ( .A1(b_7_), .A2(n13594), .A3(a_16_), .ZN(n13593) );
  OR2_X1 U13615 ( .A1(n13470), .A2(n13472), .ZN(n13594) );
  NAND2_X1 U13616 ( .A1(n13470), .A2(n13472), .ZN(n13592) );
  NAND2_X1 U13617 ( .A1(n13595), .A2(n13596), .ZN(n13472) );
  NAND3_X1 U13618 ( .A1(b_7_), .A2(n13597), .A3(a_17_), .ZN(n13596) );
  NAND2_X1 U13619 ( .A1(n13372), .A2(n13371), .ZN(n13597) );
  OR2_X1 U13620 ( .A1(n13371), .A2(n13372), .ZN(n13595) );
  AND2_X1 U13621 ( .A1(n13598), .A2(n13599), .ZN(n13372) );
  NAND3_X1 U13622 ( .A1(b_7_), .A2(n13600), .A3(a_18_), .ZN(n13599) );
  OR2_X1 U13623 ( .A1(n13378), .A2(n13380), .ZN(n13600) );
  NAND2_X1 U13624 ( .A1(n13378), .A2(n13380), .ZN(n13598) );
  NAND2_X1 U13625 ( .A1(n13601), .A2(n13602), .ZN(n13380) );
  NAND3_X1 U13626 ( .A1(b_7_), .A2(n13603), .A3(a_19_), .ZN(n13602) );
  OR2_X1 U13627 ( .A1(n13468), .A2(n13466), .ZN(n13603) );
  NAND2_X1 U13628 ( .A1(n13466), .A2(n13468), .ZN(n13601) );
  NAND2_X1 U13629 ( .A1(n13604), .A2(n13605), .ZN(n13468) );
  NAND3_X1 U13630 ( .A1(b_7_), .A2(n13606), .A3(a_20_), .ZN(n13605) );
  NAND2_X1 U13631 ( .A1(n13464), .A2(n13463), .ZN(n13606) );
  OR2_X1 U13632 ( .A1(n13463), .A2(n13464), .ZN(n13604) );
  AND2_X1 U13633 ( .A1(n13607), .A2(n13608), .ZN(n13464) );
  NAND3_X1 U13634 ( .A1(a_21_), .A2(n13609), .A3(b_7_), .ZN(n13608) );
  OR2_X1 U13635 ( .A1(n13459), .A2(n13460), .ZN(n13609) );
  NAND2_X1 U13636 ( .A1(n13459), .A2(n13460), .ZN(n13607) );
  NAND2_X1 U13637 ( .A1(n13456), .A2(n13610), .ZN(n13460) );
  NAND2_X1 U13638 ( .A1(n13455), .A2(n13457), .ZN(n13610) );
  NAND2_X1 U13639 ( .A1(n13611), .A2(n13612), .ZN(n13457) );
  NAND2_X1 U13640 ( .A1(a_22_), .A2(b_7_), .ZN(n13612) );
  INV_X1 U13641 ( .A(n13613), .ZN(n13611) );
  XOR2_X1 U13642 ( .A(n13614), .B(n13615), .Z(n13455) );
  XOR2_X1 U13643 ( .A(n13616), .B(n13617), .Z(n13614) );
  NOR2_X1 U13644 ( .A1(n7955), .A2(n7963), .ZN(n13617) );
  NAND2_X1 U13645 ( .A1(a_22_), .A2(n13613), .ZN(n13456) );
  NAND2_X1 U13646 ( .A1(n13618), .A2(n13619), .ZN(n13613) );
  NAND3_X1 U13647 ( .A1(a_23_), .A2(n13620), .A3(b_7_), .ZN(n13619) );
  OR2_X1 U13648 ( .A1(n13451), .A2(n13452), .ZN(n13620) );
  NAND2_X1 U13649 ( .A1(n13451), .A2(n13452), .ZN(n13618) );
  NAND2_X1 U13650 ( .A1(n13621), .A2(n13622), .ZN(n13452) );
  NAND2_X1 U13651 ( .A1(n13449), .A2(n13623), .ZN(n13622) );
  OR2_X1 U13652 ( .A1(n13447), .A2(n13448), .ZN(n13623) );
  NOR2_X1 U13653 ( .A1(n7954), .A2(n7789), .ZN(n13449) );
  NAND2_X1 U13654 ( .A1(n13447), .A2(n13448), .ZN(n13621) );
  NAND2_X1 U13655 ( .A1(n13624), .A2(n13625), .ZN(n13448) );
  NAND2_X1 U13656 ( .A1(n13445), .A2(n13626), .ZN(n13625) );
  OR2_X1 U13657 ( .A1(n13443), .A2(n13444), .ZN(n13626) );
  NOR2_X1 U13658 ( .A1(n7789), .A2(n7952), .ZN(n13445) );
  NAND2_X1 U13659 ( .A1(n13443), .A2(n13444), .ZN(n13624) );
  NAND2_X1 U13660 ( .A1(n13440), .A2(n13627), .ZN(n13444) );
  NAND2_X1 U13661 ( .A1(n13439), .A2(n13441), .ZN(n13627) );
  NAND2_X1 U13662 ( .A1(n13628), .A2(n13629), .ZN(n13441) );
  NAND2_X1 U13663 ( .A1(a_26_), .A2(b_7_), .ZN(n13629) );
  INV_X1 U13664 ( .A(n13630), .ZN(n13628) );
  XNOR2_X1 U13665 ( .A(n13631), .B(n13632), .ZN(n13439) );
  NAND2_X1 U13666 ( .A1(n13633), .A2(n13634), .ZN(n13631) );
  NAND2_X1 U13667 ( .A1(a_26_), .A2(n13630), .ZN(n13440) );
  NAND2_X1 U13668 ( .A1(n13412), .A2(n13635), .ZN(n13630) );
  NAND2_X1 U13669 ( .A1(n13411), .A2(n13413), .ZN(n13635) );
  NAND2_X1 U13670 ( .A1(n13636), .A2(n13637), .ZN(n13413) );
  NAND2_X1 U13671 ( .A1(b_7_), .A2(a_27_), .ZN(n13637) );
  INV_X1 U13672 ( .A(n13638), .ZN(n13636) );
  XNOR2_X1 U13673 ( .A(n13639), .B(n13640), .ZN(n13411) );
  XOR2_X1 U13674 ( .A(n13641), .B(n13642), .Z(n13639) );
  NAND2_X1 U13675 ( .A1(b_6_), .A2(a_28_), .ZN(n13641) );
  NAND2_X1 U13676 ( .A1(a_27_), .A2(n13638), .ZN(n13412) );
  NAND2_X1 U13677 ( .A1(n13643), .A2(n13644), .ZN(n13638) );
  NAND3_X1 U13678 ( .A1(a_28_), .A2(n13645), .A3(b_7_), .ZN(n13644) );
  NAND2_X1 U13679 ( .A1(n13421), .A2(n13419), .ZN(n13645) );
  OR2_X1 U13680 ( .A1(n13419), .A2(n13421), .ZN(n13643) );
  AND2_X1 U13681 ( .A1(n13646), .A2(n13647), .ZN(n13421) );
  NAND2_X1 U13682 ( .A1(n13435), .A2(n13648), .ZN(n13647) );
  OR2_X1 U13683 ( .A1(n13436), .A2(n13437), .ZN(n13648) );
  NOR2_X1 U13684 ( .A1(n7789), .A2(n7460), .ZN(n13435) );
  INV_X1 U13685 ( .A(b_7_), .ZN(n7789) );
  NAND2_X1 U13686 ( .A1(n13437), .A2(n13436), .ZN(n13646) );
  NAND2_X1 U13687 ( .A1(n13649), .A2(n13650), .ZN(n13436) );
  NAND2_X1 U13688 ( .A1(b_5_), .A2(n13651), .ZN(n13650) );
  NAND2_X1 U13689 ( .A1(n7441), .A2(n13652), .ZN(n13651) );
  NAND2_X1 U13690 ( .A1(a_31_), .A2(n7963), .ZN(n13652) );
  NAND2_X1 U13691 ( .A1(b_6_), .A2(n13653), .ZN(n13649) );
  NAND2_X1 U13692 ( .A1(n7445), .A2(n13654), .ZN(n13653) );
  NAND2_X1 U13693 ( .A1(a_30_), .A2(n7816), .ZN(n13654) );
  AND3_X1 U13694 ( .A1(b_7_), .A2(n7409), .A3(b_6_), .ZN(n13437) );
  XNOR2_X1 U13695 ( .A(n13655), .B(n13656), .ZN(n13419) );
  XOR2_X1 U13696 ( .A(n13657), .B(n13658), .Z(n13655) );
  XNOR2_X1 U13697 ( .A(n13659), .B(n13660), .ZN(n13443) );
  NAND2_X1 U13698 ( .A1(n13661), .A2(n13662), .ZN(n13659) );
  XNOR2_X1 U13699 ( .A(n13663), .B(n13664), .ZN(n13447) );
  NAND2_X1 U13700 ( .A1(n13665), .A2(n13666), .ZN(n13663) );
  XNOR2_X1 U13701 ( .A(n13667), .B(n13668), .ZN(n13451) );
  XNOR2_X1 U13702 ( .A(n13669), .B(n13670), .ZN(n13668) );
  XNOR2_X1 U13703 ( .A(n13671), .B(n13672), .ZN(n13459) );
  NAND2_X1 U13704 ( .A1(n13673), .A2(n13674), .ZN(n13671) );
  XOR2_X1 U13705 ( .A(n13675), .B(n13676), .Z(n13463) );
  XNOR2_X1 U13706 ( .A(n13677), .B(n13678), .ZN(n13676) );
  XOR2_X1 U13707 ( .A(n13679), .B(n13680), .Z(n13466) );
  XOR2_X1 U13708 ( .A(n13681), .B(n13682), .Z(n13679) );
  NOR2_X1 U13709 ( .A1(n7963), .A2(n7957), .ZN(n13682) );
  XNOR2_X1 U13710 ( .A(n13683), .B(n13684), .ZN(n13378) );
  XNOR2_X1 U13711 ( .A(n13685), .B(n13686), .ZN(n13684) );
  XNOR2_X1 U13712 ( .A(n13687), .B(n13688), .ZN(n13371) );
  XOR2_X1 U13713 ( .A(n13689), .B(n13690), .Z(n13687) );
  XNOR2_X1 U13714 ( .A(n13691), .B(n13692), .ZN(n13470) );
  XNOR2_X1 U13715 ( .A(n13693), .B(n13694), .ZN(n13691) );
  XOR2_X1 U13716 ( .A(n13695), .B(n13696), .Z(n13475) );
  XNOR2_X1 U13717 ( .A(n13697), .B(n13698), .ZN(n13696) );
  XNOR2_X1 U13718 ( .A(n13699), .B(n13700), .ZN(n13479) );
  XNOR2_X1 U13719 ( .A(n13701), .B(n13702), .ZN(n13699) );
  XOR2_X1 U13720 ( .A(n13703), .B(n13704), .Z(n13482) );
  XOR2_X1 U13721 ( .A(n13705), .B(n13706), .Z(n13703) );
  XNOR2_X1 U13722 ( .A(n13707), .B(n13708), .ZN(n13487) );
  XNOR2_X1 U13723 ( .A(n13709), .B(n13710), .ZN(n13707) );
  XNOR2_X1 U13724 ( .A(n13711), .B(n13712), .ZN(n13491) );
  XNOR2_X1 U13725 ( .A(n13713), .B(n13714), .ZN(n13711) );
  XNOR2_X1 U13726 ( .A(n13715), .B(n13716), .ZN(n13495) );
  XNOR2_X1 U13727 ( .A(n13717), .B(n13718), .ZN(n13716) );
  XNOR2_X1 U13728 ( .A(n13719), .B(n13720), .ZN(n13342) );
  XNOR2_X1 U13729 ( .A(n13721), .B(n13722), .ZN(n13719) );
  XNOR2_X1 U13730 ( .A(n13723), .B(n13724), .ZN(n13499) );
  XOR2_X1 U13731 ( .A(n13725), .B(n13726), .Z(n13724) );
  NAND2_X1 U13732 ( .A1(a_9_), .A2(b_6_), .ZN(n13726) );
  INV_X1 U13733 ( .A(n7899), .ZN(n7784) );
  NAND2_X1 U13734 ( .A1(a_7_), .A2(b_7_), .ZN(n7899) );
  XOR2_X1 U13735 ( .A(n13727), .B(n13728), .Z(n13506) );
  XOR2_X1 U13736 ( .A(n13729), .B(n13730), .Z(n13727) );
  NOR2_X1 U13737 ( .A1(n7963), .A2(n7787), .ZN(n13730) );
  XOR2_X1 U13738 ( .A(n13731), .B(n13732), .Z(n13510) );
  XOR2_X1 U13739 ( .A(n13733), .B(n13734), .Z(n13731) );
  XOR2_X1 U13740 ( .A(n13735), .B(n13736), .Z(n13514) );
  XOR2_X1 U13741 ( .A(n13737), .B(n13738), .Z(n13735) );
  NOR2_X1 U13742 ( .A1(n7963), .A2(n7823), .ZN(n13738) );
  XOR2_X1 U13743 ( .A(n13739), .B(n13740), .Z(n13518) );
  XNOR2_X1 U13744 ( .A(n13741), .B(n13742), .ZN(n13740) );
  NAND2_X1 U13745 ( .A1(a_4_), .A2(b_6_), .ZN(n13742) );
  XOR2_X1 U13746 ( .A(n13743), .B(n13744), .Z(n13522) );
  XOR2_X1 U13747 ( .A(n13745), .B(n13746), .Z(n13743) );
  NOR2_X1 U13748 ( .A1(n7963), .A2(n7852), .ZN(n13746) );
  XOR2_X1 U13749 ( .A(n13747), .B(n13748), .Z(n13526) );
  XOR2_X1 U13750 ( .A(n13749), .B(n13750), .Z(n13747) );
  NOR2_X1 U13751 ( .A1(n7963), .A2(n7966), .ZN(n13750) );
  XOR2_X1 U13752 ( .A(n13751), .B(n13752), .Z(n13532) );
  XOR2_X1 U13753 ( .A(n13753), .B(n13754), .Z(n13751) );
  NOR2_X1 U13754 ( .A1(n7963), .A2(n7872), .ZN(n13754) );
  XNOR2_X1 U13755 ( .A(n13755), .B(n13756), .ZN(n13530) );
  XOR2_X1 U13756 ( .A(n13757), .B(n13758), .Z(n13755) );
  NOR2_X1 U13757 ( .A1(n8197), .A2(n7963), .ZN(n13758) );
  NAND2_X1 U13758 ( .A1(n13759), .A2(n13760), .ZN(n7485) );
  NAND2_X1 U13759 ( .A1(n13761), .A2(n13762), .ZN(n13760) );
  NAND2_X1 U13760 ( .A1(n13538), .A2(n13537), .ZN(n13759) );
  NAND4_X1 U13761 ( .A1(n13538), .A2(n13761), .A3(n13537), .A4(n13762), .ZN(
        n7484) );
  NAND2_X1 U13762 ( .A1(n13763), .A2(n13764), .ZN(n13537) );
  NAND3_X1 U13763 ( .A1(a_0_), .A2(n13765), .A3(b_6_), .ZN(n13764) );
  OR2_X1 U13764 ( .A1(n13756), .A2(n13757), .ZN(n13765) );
  NAND2_X1 U13765 ( .A1(n13756), .A2(n13757), .ZN(n13763) );
  NAND2_X1 U13766 ( .A1(n13766), .A2(n13767), .ZN(n13757) );
  NAND3_X1 U13767 ( .A1(b_6_), .A2(n13768), .A3(a_1_), .ZN(n13767) );
  OR2_X1 U13768 ( .A1(n13753), .A2(n13752), .ZN(n13768) );
  NAND2_X1 U13769 ( .A1(n13752), .A2(n13753), .ZN(n13766) );
  NAND2_X1 U13770 ( .A1(n13769), .A2(n13770), .ZN(n13753) );
  NAND3_X1 U13771 ( .A1(b_6_), .A2(n13771), .A3(a_2_), .ZN(n13770) );
  OR2_X1 U13772 ( .A1(n13749), .A2(n13748), .ZN(n13771) );
  NAND2_X1 U13773 ( .A1(n13748), .A2(n13749), .ZN(n13769) );
  NAND2_X1 U13774 ( .A1(n13772), .A2(n13773), .ZN(n13749) );
  NAND3_X1 U13775 ( .A1(b_6_), .A2(n13774), .A3(a_3_), .ZN(n13773) );
  OR2_X1 U13776 ( .A1(n13745), .A2(n13744), .ZN(n13774) );
  NAND2_X1 U13777 ( .A1(n13744), .A2(n13745), .ZN(n13772) );
  NAND2_X1 U13778 ( .A1(n13775), .A2(n13776), .ZN(n13745) );
  NAND3_X1 U13779 ( .A1(b_6_), .A2(n13777), .A3(a_4_), .ZN(n13776) );
  NAND2_X1 U13780 ( .A1(n13741), .A2(n13739), .ZN(n13777) );
  OR2_X1 U13781 ( .A1(n13739), .A2(n13741), .ZN(n13775) );
  AND2_X1 U13782 ( .A1(n13778), .A2(n13779), .ZN(n13741) );
  NAND3_X1 U13783 ( .A1(b_6_), .A2(n13780), .A3(a_5_), .ZN(n13779) );
  OR2_X1 U13784 ( .A1(n13737), .A2(n13736), .ZN(n13780) );
  NAND2_X1 U13785 ( .A1(n13736), .A2(n13737), .ZN(n13778) );
  NAND2_X1 U13786 ( .A1(n13781), .A2(n13782), .ZN(n13737) );
  NAND2_X1 U13787 ( .A1(n13732), .A2(n13783), .ZN(n13782) );
  OR2_X1 U13788 ( .A1(n13733), .A2(n13734), .ZN(n13783) );
  XNOR2_X1 U13789 ( .A(n13784), .B(n13785), .ZN(n13732) );
  XNOR2_X1 U13790 ( .A(n13786), .B(n13787), .ZN(n13784) );
  NOR2_X1 U13791 ( .A1(n7816), .A2(n7787), .ZN(n13787) );
  NAND2_X1 U13792 ( .A1(n13734), .A2(n13733), .ZN(n13781) );
  NAND2_X1 U13793 ( .A1(n13788), .A2(n13789), .ZN(n13733) );
  NAND3_X1 U13794 ( .A1(b_6_), .A2(n13790), .A3(a_7_), .ZN(n13789) );
  OR2_X1 U13795 ( .A1(n13729), .A2(n13728), .ZN(n13790) );
  NAND2_X1 U13796 ( .A1(n13728), .A2(n13729), .ZN(n13788) );
  NAND2_X1 U13797 ( .A1(n13791), .A2(n13792), .ZN(n13729) );
  NAND3_X1 U13798 ( .A1(b_6_), .A2(n13793), .A3(a_8_), .ZN(n13792) );
  OR2_X1 U13799 ( .A1(n13566), .A2(n13564), .ZN(n13793) );
  NAND2_X1 U13800 ( .A1(n13564), .A2(n13566), .ZN(n13791) );
  NAND2_X1 U13801 ( .A1(n13794), .A2(n13795), .ZN(n13566) );
  NAND3_X1 U13802 ( .A1(b_6_), .A2(n13796), .A3(a_9_), .ZN(n13795) );
  OR2_X1 U13803 ( .A1(n13725), .A2(n13723), .ZN(n13796) );
  NAND2_X1 U13804 ( .A1(n13723), .A2(n13725), .ZN(n13794) );
  NAND2_X1 U13805 ( .A1(n13797), .A2(n13798), .ZN(n13725) );
  NAND2_X1 U13806 ( .A1(n13722), .A2(n13799), .ZN(n13798) );
  NAND2_X1 U13807 ( .A1(n13721), .A2(n13720), .ZN(n13799) );
  NOR2_X1 U13808 ( .A1(n8378), .A2(n7963), .ZN(n13722) );
  OR2_X1 U13809 ( .A1(n13720), .A2(n13721), .ZN(n13797) );
  AND2_X1 U13810 ( .A1(n13800), .A2(n13801), .ZN(n13721) );
  NAND2_X1 U13811 ( .A1(n13718), .A2(n13802), .ZN(n13801) );
  OR2_X1 U13812 ( .A1(n13717), .A2(n13715), .ZN(n13802) );
  NOR2_X1 U13813 ( .A1(n7963), .A2(n7724), .ZN(n13718) );
  NAND2_X1 U13814 ( .A1(n13715), .A2(n13717), .ZN(n13800) );
  NAND2_X1 U13815 ( .A1(n13803), .A2(n13804), .ZN(n13717) );
  NAND2_X1 U13816 ( .A1(n13714), .A2(n13805), .ZN(n13804) );
  NAND2_X1 U13817 ( .A1(n13713), .A2(n13712), .ZN(n13805) );
  NOR2_X1 U13818 ( .A1(n8585), .A2(n7963), .ZN(n13714) );
  OR2_X1 U13819 ( .A1(n13712), .A2(n13713), .ZN(n13803) );
  AND2_X1 U13820 ( .A1(n13806), .A2(n13807), .ZN(n13713) );
  NAND2_X1 U13821 ( .A1(n13710), .A2(n13808), .ZN(n13807) );
  NAND2_X1 U13822 ( .A1(n13709), .A2(n13708), .ZN(n13808) );
  NOR2_X1 U13823 ( .A1(n7702), .A2(n7963), .ZN(n13710) );
  OR2_X1 U13824 ( .A1(n13708), .A2(n13709), .ZN(n13806) );
  AND2_X1 U13825 ( .A1(n13809), .A2(n13810), .ZN(n13709) );
  NAND2_X1 U13826 ( .A1(n13706), .A2(n13811), .ZN(n13810) );
  OR2_X1 U13827 ( .A1(n13704), .A2(n13705), .ZN(n13811) );
  NOR2_X1 U13828 ( .A1(n7962), .A2(n7963), .ZN(n13706) );
  NAND2_X1 U13829 ( .A1(n13704), .A2(n13705), .ZN(n13809) );
  NAND2_X1 U13830 ( .A1(n13812), .A2(n13813), .ZN(n13705) );
  NAND2_X1 U13831 ( .A1(n13702), .A2(n13814), .ZN(n13813) );
  NAND2_X1 U13832 ( .A1(n13701), .A2(n13700), .ZN(n13814) );
  NOR2_X1 U13833 ( .A1(n7667), .A2(n7963), .ZN(n13702) );
  OR2_X1 U13834 ( .A1(n13700), .A2(n13701), .ZN(n13812) );
  AND2_X1 U13835 ( .A1(n13815), .A2(n13816), .ZN(n13701) );
  NAND2_X1 U13836 ( .A1(n13698), .A2(n13817), .ZN(n13816) );
  OR2_X1 U13837 ( .A1(n13695), .A2(n13697), .ZN(n13817) );
  NOR2_X1 U13838 ( .A1(n8353), .A2(n7963), .ZN(n13698) );
  NAND2_X1 U13839 ( .A1(n13695), .A2(n13697), .ZN(n13815) );
  NAND2_X1 U13840 ( .A1(n13818), .A2(n13819), .ZN(n13697) );
  NAND2_X1 U13841 ( .A1(n13694), .A2(n13820), .ZN(n13819) );
  NAND2_X1 U13842 ( .A1(n13693), .A2(n13692), .ZN(n13820) );
  NOR2_X1 U13843 ( .A1(n7645), .A2(n7963), .ZN(n13694) );
  OR2_X1 U13844 ( .A1(n13692), .A2(n13693), .ZN(n13818) );
  AND2_X1 U13845 ( .A1(n13821), .A2(n13822), .ZN(n13693) );
  NAND2_X1 U13846 ( .A1(n13690), .A2(n13823), .ZN(n13822) );
  OR2_X1 U13847 ( .A1(n13688), .A2(n13689), .ZN(n13823) );
  NOR2_X1 U13848 ( .A1(n7960), .A2(n7963), .ZN(n13690) );
  NAND2_X1 U13849 ( .A1(n13688), .A2(n13689), .ZN(n13821) );
  NAND2_X1 U13850 ( .A1(n13824), .A2(n13825), .ZN(n13689) );
  NAND2_X1 U13851 ( .A1(n13686), .A2(n13826), .ZN(n13825) );
  OR2_X1 U13852 ( .A1(n13685), .A2(n13683), .ZN(n13826) );
  NOR2_X1 U13853 ( .A1(n7958), .A2(n7963), .ZN(n13686) );
  NAND2_X1 U13854 ( .A1(n13683), .A2(n13685), .ZN(n13824) );
  NAND2_X1 U13855 ( .A1(n13827), .A2(n13828), .ZN(n13685) );
  NAND3_X1 U13856 ( .A1(b_6_), .A2(n13829), .A3(a_20_), .ZN(n13828) );
  OR2_X1 U13857 ( .A1(n13680), .A2(n13681), .ZN(n13829) );
  NAND2_X1 U13858 ( .A1(n13680), .A2(n13681), .ZN(n13827) );
  NAND2_X1 U13859 ( .A1(n13830), .A2(n13831), .ZN(n13681) );
  NAND2_X1 U13860 ( .A1(n13678), .A2(n13832), .ZN(n13831) );
  OR2_X1 U13861 ( .A1(n13675), .A2(n13677), .ZN(n13832) );
  NOR2_X1 U13862 ( .A1(n7963), .A2(n7578), .ZN(n13678) );
  NAND2_X1 U13863 ( .A1(n13675), .A2(n13677), .ZN(n13830) );
  NAND2_X1 U13864 ( .A1(n13673), .A2(n13833), .ZN(n13677) );
  NAND2_X1 U13865 ( .A1(n13672), .A2(n13674), .ZN(n13833) );
  NAND2_X1 U13866 ( .A1(n13834), .A2(n13835), .ZN(n13674) );
  NAND2_X1 U13867 ( .A1(a_22_), .A2(b_6_), .ZN(n13835) );
  INV_X1 U13868 ( .A(n13836), .ZN(n13834) );
  XNOR2_X1 U13869 ( .A(n13837), .B(n13838), .ZN(n13672) );
  XOR2_X1 U13870 ( .A(n13839), .B(n13840), .Z(n13838) );
  NAND2_X1 U13871 ( .A1(b_5_), .A2(a_23_), .ZN(n13840) );
  NAND2_X1 U13872 ( .A1(a_22_), .A2(n13836), .ZN(n13673) );
  NAND2_X1 U13873 ( .A1(n13841), .A2(n13842), .ZN(n13836) );
  NAND3_X1 U13874 ( .A1(a_23_), .A2(n13843), .A3(b_6_), .ZN(n13842) );
  OR2_X1 U13875 ( .A1(n13615), .A2(n13616), .ZN(n13843) );
  NAND2_X1 U13876 ( .A1(n13615), .A2(n13616), .ZN(n13841) );
  NAND2_X1 U13877 ( .A1(n13844), .A2(n13845), .ZN(n13616) );
  NAND2_X1 U13878 ( .A1(n13670), .A2(n13846), .ZN(n13845) );
  OR2_X1 U13879 ( .A1(n13669), .A2(n13667), .ZN(n13846) );
  NOR2_X1 U13880 ( .A1(n7954), .A2(n7963), .ZN(n13670) );
  NAND2_X1 U13881 ( .A1(n13667), .A2(n13669), .ZN(n13844) );
  NAND2_X1 U13882 ( .A1(n13665), .A2(n13847), .ZN(n13669) );
  NAND2_X1 U13883 ( .A1(n13664), .A2(n13666), .ZN(n13847) );
  NAND2_X1 U13884 ( .A1(n13848), .A2(n13849), .ZN(n13666) );
  NAND2_X1 U13885 ( .A1(b_6_), .A2(a_25_), .ZN(n13849) );
  INV_X1 U13886 ( .A(n13850), .ZN(n13848) );
  XNOR2_X1 U13887 ( .A(n13851), .B(n13852), .ZN(n13664) );
  NAND2_X1 U13888 ( .A1(n13853), .A2(n13854), .ZN(n13851) );
  NAND2_X1 U13889 ( .A1(a_25_), .A2(n13850), .ZN(n13665) );
  NAND2_X1 U13890 ( .A1(n13661), .A2(n13855), .ZN(n13850) );
  NAND2_X1 U13891 ( .A1(n13660), .A2(n13662), .ZN(n13855) );
  NAND2_X1 U13892 ( .A1(n13856), .A2(n13857), .ZN(n13662) );
  NAND2_X1 U13893 ( .A1(b_6_), .A2(a_26_), .ZN(n13857) );
  INV_X1 U13894 ( .A(n13858), .ZN(n13856) );
  XNOR2_X1 U13895 ( .A(n13859), .B(n13860), .ZN(n13660) );
  NAND2_X1 U13896 ( .A1(n13861), .A2(n13862), .ZN(n13859) );
  NAND2_X1 U13897 ( .A1(a_26_), .A2(n13858), .ZN(n13661) );
  NAND2_X1 U13898 ( .A1(n13633), .A2(n13863), .ZN(n13858) );
  NAND2_X1 U13899 ( .A1(n13632), .A2(n13634), .ZN(n13863) );
  NAND2_X1 U13900 ( .A1(n13864), .A2(n13865), .ZN(n13634) );
  NAND2_X1 U13901 ( .A1(b_6_), .A2(a_27_), .ZN(n13865) );
  INV_X1 U13902 ( .A(n13866), .ZN(n13864) );
  XNOR2_X1 U13903 ( .A(n13867), .B(n13868), .ZN(n13632) );
  XOR2_X1 U13904 ( .A(n13869), .B(n13870), .Z(n13867) );
  NAND2_X1 U13905 ( .A1(b_5_), .A2(a_28_), .ZN(n13869) );
  NAND2_X1 U13906 ( .A1(a_27_), .A2(n13866), .ZN(n13633) );
  NAND2_X1 U13907 ( .A1(n13871), .A2(n13872), .ZN(n13866) );
  NAND3_X1 U13908 ( .A1(a_28_), .A2(n13873), .A3(b_6_), .ZN(n13872) );
  NAND2_X1 U13909 ( .A1(n13642), .A2(n13640), .ZN(n13873) );
  OR2_X1 U13910 ( .A1(n13640), .A2(n13642), .ZN(n13871) );
  AND2_X1 U13911 ( .A1(n13874), .A2(n13875), .ZN(n13642) );
  NAND2_X1 U13912 ( .A1(n13656), .A2(n13876), .ZN(n13875) );
  OR2_X1 U13913 ( .A1(n13657), .A2(n13658), .ZN(n13876) );
  NOR2_X1 U13914 ( .A1(n7963), .A2(n7460), .ZN(n13656) );
  INV_X1 U13915 ( .A(b_6_), .ZN(n7963) );
  NAND2_X1 U13916 ( .A1(n13658), .A2(n13657), .ZN(n13874) );
  NAND2_X1 U13917 ( .A1(n13877), .A2(n13878), .ZN(n13657) );
  NAND2_X1 U13918 ( .A1(b_4_), .A2(n13879), .ZN(n13878) );
  NAND2_X1 U13919 ( .A1(n7441), .A2(n13880), .ZN(n13879) );
  NAND2_X1 U13920 ( .A1(a_31_), .A2(n7816), .ZN(n13880) );
  NAND2_X1 U13921 ( .A1(b_5_), .A2(n13881), .ZN(n13877) );
  NAND2_X1 U13922 ( .A1(n7445), .A2(n13882), .ZN(n13881) );
  NAND2_X1 U13923 ( .A1(a_30_), .A2(n7964), .ZN(n13882) );
  AND3_X1 U13924 ( .A1(b_6_), .A2(n7409), .A3(b_5_), .ZN(n13658) );
  XNOR2_X1 U13925 ( .A(n13883), .B(n13884), .ZN(n13640) );
  XOR2_X1 U13926 ( .A(n13885), .B(n13886), .Z(n13883) );
  XNOR2_X1 U13927 ( .A(n13887), .B(n13888), .ZN(n13667) );
  NAND2_X1 U13928 ( .A1(n13889), .A2(n13890), .ZN(n13887) );
  XNOR2_X1 U13929 ( .A(n13891), .B(n13892), .ZN(n13615) );
  XOR2_X1 U13930 ( .A(n13893), .B(n13894), .Z(n13892) );
  NAND2_X1 U13931 ( .A1(a_24_), .A2(b_5_), .ZN(n13894) );
  XNOR2_X1 U13932 ( .A(n13895), .B(n13896), .ZN(n13675) );
  XOR2_X1 U13933 ( .A(n13897), .B(n13898), .Z(n13896) );
  NAND2_X1 U13934 ( .A1(a_22_), .A2(b_5_), .ZN(n13898) );
  XNOR2_X1 U13935 ( .A(n13899), .B(n13900), .ZN(n13680) );
  XOR2_X1 U13936 ( .A(n13901), .B(n13902), .Z(n13900) );
  NAND2_X1 U13937 ( .A1(b_5_), .A2(a_21_), .ZN(n13902) );
  XOR2_X1 U13938 ( .A(n13903), .B(n13904), .Z(n13683) );
  XOR2_X1 U13939 ( .A(n13905), .B(n13906), .Z(n13903) );
  NOR2_X1 U13940 ( .A1(n7816), .A2(n7957), .ZN(n13906) );
  XNOR2_X1 U13941 ( .A(n13907), .B(n13908), .ZN(n13688) );
  XOR2_X1 U13942 ( .A(n13909), .B(n13910), .Z(n13908) );
  NAND2_X1 U13943 ( .A1(a_19_), .A2(b_5_), .ZN(n13910) );
  XNOR2_X1 U13944 ( .A(n13911), .B(n13912), .ZN(n13692) );
  XOR2_X1 U13945 ( .A(n13913), .B(n13914), .Z(n13911) );
  NOR2_X1 U13946 ( .A1(n7816), .A2(n7960), .ZN(n13914) );
  XNOR2_X1 U13947 ( .A(n13915), .B(n13916), .ZN(n13695) );
  XNOR2_X1 U13948 ( .A(n13917), .B(n13918), .ZN(n13915) );
  NOR2_X1 U13949 ( .A1(n7816), .A2(n7645), .ZN(n13918) );
  XNOR2_X1 U13950 ( .A(n13919), .B(n13920), .ZN(n13700) );
  XOR2_X1 U13951 ( .A(n13921), .B(n13922), .Z(n13919) );
  NOR2_X1 U13952 ( .A1(n7816), .A2(n8353), .ZN(n13922) );
  XNOR2_X1 U13953 ( .A(n13923), .B(n13924), .ZN(n13704) );
  XNOR2_X1 U13954 ( .A(n13925), .B(n13926), .ZN(n13923) );
  NOR2_X1 U13955 ( .A1(n7816), .A2(n7667), .ZN(n13926) );
  XNOR2_X1 U13956 ( .A(n13927), .B(n13928), .ZN(n13708) );
  XOR2_X1 U13957 ( .A(n13929), .B(n13930), .Z(n13927) );
  NOR2_X1 U13958 ( .A1(n7816), .A2(n7962), .ZN(n13930) );
  XNOR2_X1 U13959 ( .A(n13931), .B(n13932), .ZN(n13712) );
  XOR2_X1 U13960 ( .A(n13933), .B(n13934), .Z(n13931) );
  NOR2_X1 U13961 ( .A1(n7816), .A2(n7702), .ZN(n13934) );
  XOR2_X1 U13962 ( .A(n13935), .B(n13936), .Z(n13715) );
  XOR2_X1 U13963 ( .A(n13937), .B(n13938), .Z(n13935) );
  NOR2_X1 U13964 ( .A1(n7816), .A2(n8585), .ZN(n13938) );
  XNOR2_X1 U13965 ( .A(n13939), .B(n13940), .ZN(n13720) );
  XOR2_X1 U13966 ( .A(n13941), .B(n13942), .Z(n13939) );
  NOR2_X1 U13967 ( .A1(n7724), .A2(n7816), .ZN(n13942) );
  XOR2_X1 U13968 ( .A(n13943), .B(n13944), .Z(n13723) );
  XOR2_X1 U13969 ( .A(n13945), .B(n13946), .Z(n13943) );
  NOR2_X1 U13970 ( .A1(n7816), .A2(n8378), .ZN(n13946) );
  XNOR2_X1 U13971 ( .A(n13947), .B(n13948), .ZN(n13564) );
  XNOR2_X1 U13972 ( .A(n13949), .B(n13950), .ZN(n13947) );
  NOR2_X1 U13973 ( .A1(n7816), .A2(n7753), .ZN(n13950) );
  XOR2_X1 U13974 ( .A(n13951), .B(n13952), .Z(n13728) );
  XOR2_X1 U13975 ( .A(n13953), .B(n13954), .Z(n13951) );
  NOR2_X1 U13976 ( .A1(n7816), .A2(n8602), .ZN(n13954) );
  INV_X1 U13977 ( .A(n7801), .ZN(n13734) );
  NAND2_X1 U13978 ( .A1(a_6_), .A2(b_6_), .ZN(n7801) );
  XOR2_X1 U13979 ( .A(n13955), .B(n13956), .Z(n13736) );
  XOR2_X1 U13980 ( .A(n13957), .B(n13958), .Z(n13955) );
  NOR2_X1 U13981 ( .A1(n7816), .A2(n7807), .ZN(n13958) );
  XNOR2_X1 U13982 ( .A(n13959), .B(n13960), .ZN(n13739) );
  XOR2_X1 U13983 ( .A(n13961), .B(n7814), .Z(n13959) );
  XOR2_X1 U13984 ( .A(n13962), .B(n13963), .Z(n13744) );
  XOR2_X1 U13985 ( .A(n13964), .B(n13965), .Z(n13962) );
  NOR2_X1 U13986 ( .A1(n7816), .A2(n7836), .ZN(n13965) );
  XOR2_X1 U13987 ( .A(n13966), .B(n13967), .Z(n13748) );
  XOR2_X1 U13988 ( .A(n13968), .B(n13969), .Z(n13966) );
  NOR2_X1 U13989 ( .A1(n7816), .A2(n7852), .ZN(n13969) );
  XOR2_X1 U13990 ( .A(n13970), .B(n13971), .Z(n13752) );
  XOR2_X1 U13991 ( .A(n13972), .B(n13973), .Z(n13970) );
  NOR2_X1 U13992 ( .A1(n7816), .A2(n7966), .ZN(n13973) );
  XOR2_X1 U13993 ( .A(n13974), .B(n13975), .Z(n13756) );
  XOR2_X1 U13994 ( .A(n13976), .B(n13977), .Z(n13974) );
  NAND2_X1 U13995 ( .A1(n13978), .A2(n13979), .ZN(n13761) );
  XOR2_X1 U13996 ( .A(n13980), .B(n13981), .Z(n13538) );
  XOR2_X1 U13997 ( .A(n13982), .B(n13983), .Z(n13980) );
  NAND2_X1 U13998 ( .A1(n13984), .A2(n13762), .ZN(n7629) );
  INV_X1 U13999 ( .A(n13985), .ZN(n13762) );
  XNOR2_X1 U14000 ( .A(n13986), .B(n13987), .ZN(n13984) );
  NAND2_X1 U14001 ( .A1(n13985), .A2(n13988), .ZN(n7628) );
  XOR2_X1 U14002 ( .A(n13986), .B(n13987), .Z(n13988) );
  NOR2_X1 U14003 ( .A1(n13979), .A2(n13978), .ZN(n13985) );
  AND2_X1 U14004 ( .A1(n13989), .A2(n13990), .ZN(n13978) );
  NAND2_X1 U14005 ( .A1(n13983), .A2(n13991), .ZN(n13990) );
  OR2_X1 U14006 ( .A1(n13981), .A2(n13982), .ZN(n13991) );
  NOR2_X1 U14007 ( .A1(n7816), .A2(n8197), .ZN(n13983) );
  NAND2_X1 U14008 ( .A1(n13981), .A2(n13982), .ZN(n13989) );
  NAND2_X1 U14009 ( .A1(n13992), .A2(n13993), .ZN(n13982) );
  NAND2_X1 U14010 ( .A1(n13977), .A2(n13994), .ZN(n13993) );
  OR2_X1 U14011 ( .A1(n13976), .A2(n13975), .ZN(n13994) );
  NOR2_X1 U14012 ( .A1(n7872), .A2(n7816), .ZN(n13977) );
  NAND2_X1 U14013 ( .A1(n13975), .A2(n13976), .ZN(n13992) );
  NAND2_X1 U14014 ( .A1(n13995), .A2(n13996), .ZN(n13976) );
  NAND3_X1 U14015 ( .A1(b_5_), .A2(n13997), .A3(a_2_), .ZN(n13996) );
  OR2_X1 U14016 ( .A1(n13971), .A2(n13972), .ZN(n13997) );
  NAND2_X1 U14017 ( .A1(n13971), .A2(n13972), .ZN(n13995) );
  NAND2_X1 U14018 ( .A1(n13998), .A2(n13999), .ZN(n13972) );
  NAND3_X1 U14019 ( .A1(b_5_), .A2(n14000), .A3(a_3_), .ZN(n13999) );
  OR2_X1 U14020 ( .A1(n13967), .A2(n13968), .ZN(n14000) );
  NAND2_X1 U14021 ( .A1(n13967), .A2(n13968), .ZN(n13998) );
  NAND2_X1 U14022 ( .A1(n14001), .A2(n14002), .ZN(n13968) );
  NAND3_X1 U14023 ( .A1(b_5_), .A2(n14003), .A3(a_4_), .ZN(n14002) );
  OR2_X1 U14024 ( .A1(n13963), .A2(n13964), .ZN(n14003) );
  NAND2_X1 U14025 ( .A1(n13963), .A2(n13964), .ZN(n14001) );
  NAND2_X1 U14026 ( .A1(n14004), .A2(n14005), .ZN(n13964) );
  NAND2_X1 U14027 ( .A1(n13960), .A2(n14006), .ZN(n14005) );
  OR2_X1 U14028 ( .A1(n13961), .A2(n7814), .ZN(n14006) );
  XNOR2_X1 U14029 ( .A(n14007), .B(n14008), .ZN(n13960) );
  XNOR2_X1 U14030 ( .A(n14009), .B(n14010), .ZN(n14007) );
  NOR2_X1 U14031 ( .A1(n7964), .A2(n7807), .ZN(n14010) );
  NAND2_X1 U14032 ( .A1(n7814), .A2(n13961), .ZN(n14004) );
  NAND2_X1 U14033 ( .A1(n14011), .A2(n14012), .ZN(n13961) );
  NAND3_X1 U14034 ( .A1(b_5_), .A2(n14013), .A3(a_6_), .ZN(n14012) );
  OR2_X1 U14035 ( .A1(n13956), .A2(n13957), .ZN(n14013) );
  NAND2_X1 U14036 ( .A1(n13956), .A2(n13957), .ZN(n14011) );
  NAND2_X1 U14037 ( .A1(n14014), .A2(n14015), .ZN(n13957) );
  NAND3_X1 U14038 ( .A1(b_5_), .A2(n14016), .A3(a_7_), .ZN(n14015) );
  NAND2_X1 U14039 ( .A1(n13785), .A2(n13786), .ZN(n14016) );
  OR2_X1 U14040 ( .A1(n13785), .A2(n13786), .ZN(n14014) );
  AND2_X1 U14041 ( .A1(n14017), .A2(n14018), .ZN(n13786) );
  NAND3_X1 U14042 ( .A1(b_5_), .A2(n14019), .A3(a_8_), .ZN(n14018) );
  OR2_X1 U14043 ( .A1(n13952), .A2(n13953), .ZN(n14019) );
  NAND2_X1 U14044 ( .A1(n13952), .A2(n13953), .ZN(n14017) );
  NAND2_X1 U14045 ( .A1(n14020), .A2(n14021), .ZN(n13953) );
  NAND3_X1 U14046 ( .A1(b_5_), .A2(n14022), .A3(a_9_), .ZN(n14021) );
  NAND2_X1 U14047 ( .A1(n13948), .A2(n13949), .ZN(n14022) );
  OR2_X1 U14048 ( .A1(n13948), .A2(n13949), .ZN(n14020) );
  AND2_X1 U14049 ( .A1(n14023), .A2(n14024), .ZN(n13949) );
  NAND3_X1 U14050 ( .A1(b_5_), .A2(n14025), .A3(a_10_), .ZN(n14024) );
  OR2_X1 U14051 ( .A1(n13944), .A2(n13945), .ZN(n14025) );
  NAND2_X1 U14052 ( .A1(n13944), .A2(n13945), .ZN(n14023) );
  NAND2_X1 U14053 ( .A1(n14026), .A2(n14027), .ZN(n13945) );
  NAND3_X1 U14054 ( .A1(a_11_), .A2(n14028), .A3(b_5_), .ZN(n14027) );
  OR2_X1 U14055 ( .A1(n13940), .A2(n13941), .ZN(n14028) );
  NAND2_X1 U14056 ( .A1(n13940), .A2(n13941), .ZN(n14026) );
  NAND2_X1 U14057 ( .A1(n14029), .A2(n14030), .ZN(n13941) );
  NAND3_X1 U14058 ( .A1(b_5_), .A2(n14031), .A3(a_12_), .ZN(n14030) );
  OR2_X1 U14059 ( .A1(n13936), .A2(n13937), .ZN(n14031) );
  NAND2_X1 U14060 ( .A1(n13936), .A2(n13937), .ZN(n14029) );
  NAND2_X1 U14061 ( .A1(n14032), .A2(n14033), .ZN(n13937) );
  NAND3_X1 U14062 ( .A1(b_5_), .A2(n14034), .A3(a_13_), .ZN(n14033) );
  OR2_X1 U14063 ( .A1(n13932), .A2(n13933), .ZN(n14034) );
  NAND2_X1 U14064 ( .A1(n13932), .A2(n13933), .ZN(n14032) );
  NAND2_X1 U14065 ( .A1(n14035), .A2(n14036), .ZN(n13933) );
  NAND3_X1 U14066 ( .A1(b_5_), .A2(n14037), .A3(a_14_), .ZN(n14036) );
  OR2_X1 U14067 ( .A1(n13928), .A2(n13929), .ZN(n14037) );
  NAND2_X1 U14068 ( .A1(n13928), .A2(n13929), .ZN(n14035) );
  NAND2_X1 U14069 ( .A1(n14038), .A2(n14039), .ZN(n13929) );
  NAND3_X1 U14070 ( .A1(b_5_), .A2(n14040), .A3(a_15_), .ZN(n14039) );
  NAND2_X1 U14071 ( .A1(n13925), .A2(n13924), .ZN(n14040) );
  OR2_X1 U14072 ( .A1(n13924), .A2(n13925), .ZN(n14038) );
  AND2_X1 U14073 ( .A1(n14041), .A2(n14042), .ZN(n13925) );
  NAND3_X1 U14074 ( .A1(b_5_), .A2(n14043), .A3(a_16_), .ZN(n14042) );
  OR2_X1 U14075 ( .A1(n13920), .A2(n13921), .ZN(n14043) );
  NAND2_X1 U14076 ( .A1(n13920), .A2(n13921), .ZN(n14041) );
  NAND2_X1 U14077 ( .A1(n14044), .A2(n14045), .ZN(n13921) );
  NAND3_X1 U14078 ( .A1(b_5_), .A2(n14046), .A3(a_17_), .ZN(n14045) );
  NAND2_X1 U14079 ( .A1(n13917), .A2(n13916), .ZN(n14046) );
  OR2_X1 U14080 ( .A1(n13916), .A2(n13917), .ZN(n14044) );
  AND2_X1 U14081 ( .A1(n14047), .A2(n14048), .ZN(n13917) );
  NAND3_X1 U14082 ( .A1(b_5_), .A2(n14049), .A3(a_18_), .ZN(n14048) );
  OR2_X1 U14083 ( .A1(n13912), .A2(n13913), .ZN(n14049) );
  NAND2_X1 U14084 ( .A1(n13912), .A2(n13913), .ZN(n14047) );
  NAND2_X1 U14085 ( .A1(n14050), .A2(n14051), .ZN(n13913) );
  NAND3_X1 U14086 ( .A1(b_5_), .A2(n14052), .A3(a_19_), .ZN(n14051) );
  OR2_X1 U14087 ( .A1(n13909), .A2(n13907), .ZN(n14052) );
  NAND2_X1 U14088 ( .A1(n13907), .A2(n13909), .ZN(n14050) );
  NAND2_X1 U14089 ( .A1(n14053), .A2(n14054), .ZN(n13909) );
  NAND3_X1 U14090 ( .A1(b_5_), .A2(n14055), .A3(a_20_), .ZN(n14054) );
  OR2_X1 U14091 ( .A1(n13904), .A2(n13905), .ZN(n14055) );
  NAND2_X1 U14092 ( .A1(n13904), .A2(n13905), .ZN(n14053) );
  NAND2_X1 U14093 ( .A1(n14056), .A2(n14057), .ZN(n13905) );
  NAND3_X1 U14094 ( .A1(a_21_), .A2(n14058), .A3(b_5_), .ZN(n14057) );
  OR2_X1 U14095 ( .A1(n13901), .A2(n13899), .ZN(n14058) );
  NAND2_X1 U14096 ( .A1(n13899), .A2(n13901), .ZN(n14056) );
  NAND2_X1 U14097 ( .A1(n14059), .A2(n14060), .ZN(n13901) );
  NAND3_X1 U14098 ( .A1(b_5_), .A2(n14061), .A3(a_22_), .ZN(n14060) );
  OR2_X1 U14099 ( .A1(n13897), .A2(n13895), .ZN(n14061) );
  NAND2_X1 U14100 ( .A1(n13895), .A2(n13897), .ZN(n14059) );
  NAND2_X1 U14101 ( .A1(n14062), .A2(n14063), .ZN(n13897) );
  NAND3_X1 U14102 ( .A1(a_23_), .A2(n14064), .A3(b_5_), .ZN(n14063) );
  OR2_X1 U14103 ( .A1(n13839), .A2(n13837), .ZN(n14064) );
  NAND2_X1 U14104 ( .A1(n13837), .A2(n13839), .ZN(n14062) );
  NAND2_X1 U14105 ( .A1(n14065), .A2(n14066), .ZN(n13839) );
  NAND3_X1 U14106 ( .A1(b_5_), .A2(n14067), .A3(a_24_), .ZN(n14066) );
  OR2_X1 U14107 ( .A1(n13893), .A2(n13891), .ZN(n14067) );
  NAND2_X1 U14108 ( .A1(n13891), .A2(n13893), .ZN(n14065) );
  NAND2_X1 U14109 ( .A1(n13889), .A2(n14068), .ZN(n13893) );
  NAND2_X1 U14110 ( .A1(n13888), .A2(n13890), .ZN(n14068) );
  NAND2_X1 U14111 ( .A1(n14069), .A2(n14070), .ZN(n13890) );
  NAND2_X1 U14112 ( .A1(b_5_), .A2(a_25_), .ZN(n14070) );
  INV_X1 U14113 ( .A(n14071), .ZN(n14069) );
  XNOR2_X1 U14114 ( .A(n14072), .B(n14073), .ZN(n13888) );
  NAND2_X1 U14115 ( .A1(n14074), .A2(n14075), .ZN(n14072) );
  NAND2_X1 U14116 ( .A1(a_25_), .A2(n14071), .ZN(n13889) );
  NAND2_X1 U14117 ( .A1(n13853), .A2(n14076), .ZN(n14071) );
  NAND2_X1 U14118 ( .A1(n13852), .A2(n13854), .ZN(n14076) );
  NAND2_X1 U14119 ( .A1(n14077), .A2(n14078), .ZN(n13854) );
  NAND2_X1 U14120 ( .A1(b_5_), .A2(a_26_), .ZN(n14078) );
  INV_X1 U14121 ( .A(n14079), .ZN(n14077) );
  XNOR2_X1 U14122 ( .A(n14080), .B(n14081), .ZN(n13852) );
  NAND2_X1 U14123 ( .A1(n14082), .A2(n14083), .ZN(n14080) );
  NAND2_X1 U14124 ( .A1(a_26_), .A2(n14079), .ZN(n13853) );
  NAND2_X1 U14125 ( .A1(n13861), .A2(n14084), .ZN(n14079) );
  NAND2_X1 U14126 ( .A1(n13860), .A2(n13862), .ZN(n14084) );
  NAND2_X1 U14127 ( .A1(n14085), .A2(n14086), .ZN(n13862) );
  NAND2_X1 U14128 ( .A1(b_5_), .A2(a_27_), .ZN(n14086) );
  INV_X1 U14129 ( .A(n14087), .ZN(n14085) );
  XNOR2_X1 U14130 ( .A(n14088), .B(n14089), .ZN(n13860) );
  XOR2_X1 U14131 ( .A(n14090), .B(n14091), .Z(n14088) );
  NAND2_X1 U14132 ( .A1(b_4_), .A2(a_28_), .ZN(n14090) );
  NAND2_X1 U14133 ( .A1(a_27_), .A2(n14087), .ZN(n13861) );
  NAND2_X1 U14134 ( .A1(n14092), .A2(n14093), .ZN(n14087) );
  NAND3_X1 U14135 ( .A1(a_28_), .A2(n14094), .A3(b_5_), .ZN(n14093) );
  NAND2_X1 U14136 ( .A1(n13870), .A2(n13868), .ZN(n14094) );
  OR2_X1 U14137 ( .A1(n13868), .A2(n13870), .ZN(n14092) );
  AND2_X1 U14138 ( .A1(n14095), .A2(n14096), .ZN(n13870) );
  NAND2_X1 U14139 ( .A1(n13884), .A2(n14097), .ZN(n14096) );
  OR2_X1 U14140 ( .A1(n13885), .A2(n13886), .ZN(n14097) );
  NOR2_X1 U14141 ( .A1(n7816), .A2(n7460), .ZN(n13884) );
  INV_X1 U14142 ( .A(b_5_), .ZN(n7816) );
  NAND2_X1 U14143 ( .A1(n13886), .A2(n13885), .ZN(n14095) );
  NAND2_X1 U14144 ( .A1(n14098), .A2(n14099), .ZN(n13885) );
  NAND2_X1 U14145 ( .A1(b_3_), .A2(n14100), .ZN(n14099) );
  NAND2_X1 U14146 ( .A1(n7441), .A2(n14101), .ZN(n14100) );
  NAND2_X1 U14147 ( .A1(a_31_), .A2(n7964), .ZN(n14101) );
  NAND2_X1 U14148 ( .A1(b_4_), .A2(n14102), .ZN(n14098) );
  NAND2_X1 U14149 ( .A1(n7445), .A2(n14103), .ZN(n14102) );
  NAND2_X1 U14150 ( .A1(a_30_), .A2(n7845), .ZN(n14103) );
  AND3_X1 U14151 ( .A1(b_5_), .A2(n7409), .A3(b_4_), .ZN(n13886) );
  XNOR2_X1 U14152 ( .A(n14104), .B(n14105), .ZN(n13868) );
  XOR2_X1 U14153 ( .A(n14106), .B(n14107), .Z(n14104) );
  XOR2_X1 U14154 ( .A(n14108), .B(n14109), .Z(n13891) );
  XOR2_X1 U14155 ( .A(n14110), .B(n14111), .Z(n14108) );
  XOR2_X1 U14156 ( .A(n14112), .B(n14113), .Z(n13837) );
  XOR2_X1 U14157 ( .A(n14114), .B(n14115), .Z(n14112) );
  XOR2_X1 U14158 ( .A(n14116), .B(n14117), .Z(n13895) );
  XOR2_X1 U14159 ( .A(n14118), .B(n14119), .Z(n14116) );
  XNOR2_X1 U14160 ( .A(n14120), .B(n14121), .ZN(n13899) );
  XNOR2_X1 U14161 ( .A(n14122), .B(n14123), .ZN(n14121) );
  XNOR2_X1 U14162 ( .A(n14124), .B(n14125), .ZN(n13904) );
  XNOR2_X1 U14163 ( .A(n14126), .B(n14127), .ZN(n14124) );
  XOR2_X1 U14164 ( .A(n14128), .B(n14129), .Z(n13907) );
  XOR2_X1 U14165 ( .A(n14130), .B(n14131), .Z(n14128) );
  XNOR2_X1 U14166 ( .A(n14132), .B(n14133), .ZN(n13912) );
  XNOR2_X1 U14167 ( .A(n14134), .B(n14135), .ZN(n14132) );
  XNOR2_X1 U14168 ( .A(n14136), .B(n14137), .ZN(n13916) );
  XOR2_X1 U14169 ( .A(n14138), .B(n14139), .Z(n14136) );
  XNOR2_X1 U14170 ( .A(n14140), .B(n14141), .ZN(n13920) );
  XNOR2_X1 U14171 ( .A(n14142), .B(n14143), .ZN(n14140) );
  XNOR2_X1 U14172 ( .A(n14144), .B(n14145), .ZN(n13924) );
  XOR2_X1 U14173 ( .A(n14146), .B(n14147), .Z(n14144) );
  XNOR2_X1 U14174 ( .A(n14148), .B(n14149), .ZN(n13928) );
  XNOR2_X1 U14175 ( .A(n14150), .B(n14151), .ZN(n14148) );
  XNOR2_X1 U14176 ( .A(n14152), .B(n14153), .ZN(n13932) );
  XNOR2_X1 U14177 ( .A(n14154), .B(n14155), .ZN(n14152) );
  XNOR2_X1 U14178 ( .A(n14156), .B(n14157), .ZN(n13936) );
  XNOR2_X1 U14179 ( .A(n14158), .B(n14159), .ZN(n14156) );
  NOR2_X1 U14180 ( .A1(n7964), .A2(n7702), .ZN(n14159) );
  XNOR2_X1 U14181 ( .A(n14160), .B(n14161), .ZN(n13940) );
  XNOR2_X1 U14182 ( .A(n14162), .B(n14163), .ZN(n14160) );
  NOR2_X1 U14183 ( .A1(n7964), .A2(n8585), .ZN(n14163) );
  XOR2_X1 U14184 ( .A(n14164), .B(n14165), .Z(n13944) );
  XNOR2_X1 U14185 ( .A(n14166), .B(n14167), .ZN(n14165) );
  NAND2_X1 U14186 ( .A1(b_4_), .A2(a_11_), .ZN(n14167) );
  XNOR2_X1 U14187 ( .A(n14168), .B(n14169), .ZN(n13948) );
  XNOR2_X1 U14188 ( .A(n14170), .B(n14171), .ZN(n14169) );
  NAND2_X1 U14189 ( .A1(a_10_), .A2(b_4_), .ZN(n14171) );
  XOR2_X1 U14190 ( .A(n14172), .B(n14173), .Z(n13952) );
  XNOR2_X1 U14191 ( .A(n14174), .B(n14175), .ZN(n14173) );
  NAND2_X1 U14192 ( .A1(a_9_), .A2(b_4_), .ZN(n14175) );
  XNOR2_X1 U14193 ( .A(n14176), .B(n14177), .ZN(n13785) );
  XNOR2_X1 U14194 ( .A(n14178), .B(n14179), .ZN(n14177) );
  NAND2_X1 U14195 ( .A1(a_8_), .A2(b_4_), .ZN(n14179) );
  XOR2_X1 U14196 ( .A(n14180), .B(n14181), .Z(n13956) );
  XOR2_X1 U14197 ( .A(n14182), .B(n14183), .Z(n14180) );
  NOR2_X1 U14198 ( .A1(n7964), .A2(n7787), .ZN(n14183) );
  INV_X1 U14199 ( .A(n7895), .ZN(n7814) );
  NAND2_X1 U14200 ( .A1(a_5_), .A2(b_5_), .ZN(n7895) );
  XOR2_X1 U14201 ( .A(n14184), .B(n14185), .Z(n13963) );
  XOR2_X1 U14202 ( .A(n14186), .B(n14187), .Z(n14184) );
  NOR2_X1 U14203 ( .A1(n7964), .A2(n7823), .ZN(n14187) );
  XOR2_X1 U14204 ( .A(n14188), .B(n14189), .Z(n13967) );
  XOR2_X1 U14205 ( .A(n14190), .B(n14191), .Z(n14188) );
  XOR2_X1 U14206 ( .A(n14192), .B(n14193), .Z(n13971) );
  XOR2_X1 U14207 ( .A(n14194), .B(n14195), .Z(n14192) );
  NOR2_X1 U14208 ( .A1(n7964), .A2(n7852), .ZN(n14195) );
  XOR2_X1 U14209 ( .A(n14196), .B(n14197), .Z(n13975) );
  XOR2_X1 U14210 ( .A(n14198), .B(n14199), .Z(n14196) );
  NOR2_X1 U14211 ( .A1(n7964), .A2(n7966), .ZN(n14199) );
  XOR2_X1 U14212 ( .A(n14200), .B(n14201), .Z(n13981) );
  XNOR2_X1 U14213 ( .A(n14202), .B(n14203), .ZN(n14200) );
  NAND2_X1 U14214 ( .A1(a_1_), .A2(b_4_), .ZN(n14202) );
  XNOR2_X1 U14215 ( .A(n14204), .B(n14205), .ZN(n13979) );
  XOR2_X1 U14216 ( .A(n14206), .B(n14207), .Z(n14204) );
  NOR2_X1 U14217 ( .A1(n8197), .A2(n7964), .ZN(n14207) );
  NAND2_X1 U14218 ( .A1(n14208), .A2(n14209), .ZN(n7777) );
  NAND2_X1 U14219 ( .A1(n14210), .A2(n14211), .ZN(n14209) );
  NAND2_X1 U14220 ( .A1(n13987), .A2(n13986), .ZN(n14208) );
  NAND4_X1 U14221 ( .A1(n13987), .A2(n14210), .A3(n13986), .A4(n14211), .ZN(
        n7776) );
  NAND2_X1 U14222 ( .A1(n14212), .A2(n14213), .ZN(n13986) );
  NAND3_X1 U14223 ( .A1(a_0_), .A2(n14214), .A3(b_4_), .ZN(n14213) );
  OR2_X1 U14224 ( .A1(n14206), .A2(n14205), .ZN(n14214) );
  NAND2_X1 U14225 ( .A1(n14205), .A2(n14206), .ZN(n14212) );
  NAND2_X1 U14226 ( .A1(n14215), .A2(n14216), .ZN(n14206) );
  NAND3_X1 U14227 ( .A1(b_4_), .A2(n14217), .A3(a_1_), .ZN(n14216) );
  OR2_X1 U14228 ( .A1(n14203), .A2(n14201), .ZN(n14217) );
  NAND2_X1 U14229 ( .A1(n14201), .A2(n14203), .ZN(n14215) );
  NAND2_X1 U14230 ( .A1(n14218), .A2(n14219), .ZN(n14203) );
  NAND3_X1 U14231 ( .A1(b_4_), .A2(n14220), .A3(a_2_), .ZN(n14219) );
  OR2_X1 U14232 ( .A1(n14197), .A2(n14198), .ZN(n14220) );
  NAND2_X1 U14233 ( .A1(n14197), .A2(n14198), .ZN(n14218) );
  NAND2_X1 U14234 ( .A1(n14221), .A2(n14222), .ZN(n14198) );
  NAND3_X1 U14235 ( .A1(b_4_), .A2(n14223), .A3(a_3_), .ZN(n14222) );
  OR2_X1 U14236 ( .A1(n14194), .A2(n14193), .ZN(n14223) );
  NAND2_X1 U14237 ( .A1(n14193), .A2(n14194), .ZN(n14221) );
  NAND2_X1 U14238 ( .A1(n14224), .A2(n14225), .ZN(n14194) );
  NAND2_X1 U14239 ( .A1(n14189), .A2(n14226), .ZN(n14225) );
  OR2_X1 U14240 ( .A1(n14190), .A2(n14191), .ZN(n14226) );
  XNOR2_X1 U14241 ( .A(n14227), .B(n14228), .ZN(n14189) );
  NAND2_X1 U14242 ( .A1(n14229), .A2(n14230), .ZN(n14227) );
  NAND2_X1 U14243 ( .A1(n14191), .A2(n14190), .ZN(n14224) );
  NAND2_X1 U14244 ( .A1(n14231), .A2(n14232), .ZN(n14190) );
  NAND3_X1 U14245 ( .A1(b_4_), .A2(n14233), .A3(a_5_), .ZN(n14232) );
  OR2_X1 U14246 ( .A1(n14186), .A2(n14185), .ZN(n14233) );
  NAND2_X1 U14247 ( .A1(n14185), .A2(n14186), .ZN(n14231) );
  NAND2_X1 U14248 ( .A1(n14234), .A2(n14235), .ZN(n14186) );
  NAND3_X1 U14249 ( .A1(b_4_), .A2(n14236), .A3(a_6_), .ZN(n14235) );
  NAND2_X1 U14250 ( .A1(n14009), .A2(n14008), .ZN(n14236) );
  OR2_X1 U14251 ( .A1(n14008), .A2(n14009), .ZN(n14234) );
  AND2_X1 U14252 ( .A1(n14237), .A2(n14238), .ZN(n14009) );
  NAND3_X1 U14253 ( .A1(b_4_), .A2(n14239), .A3(a_7_), .ZN(n14238) );
  OR2_X1 U14254 ( .A1(n14182), .A2(n14181), .ZN(n14239) );
  NAND2_X1 U14255 ( .A1(n14181), .A2(n14182), .ZN(n14237) );
  NAND2_X1 U14256 ( .A1(n14240), .A2(n14241), .ZN(n14182) );
  NAND3_X1 U14257 ( .A1(b_4_), .A2(n14242), .A3(a_8_), .ZN(n14241) );
  NAND2_X1 U14258 ( .A1(n14178), .A2(n14176), .ZN(n14242) );
  OR2_X1 U14259 ( .A1(n14176), .A2(n14178), .ZN(n14240) );
  AND2_X1 U14260 ( .A1(n14243), .A2(n14244), .ZN(n14178) );
  NAND3_X1 U14261 ( .A1(b_4_), .A2(n14245), .A3(a_9_), .ZN(n14244) );
  NAND2_X1 U14262 ( .A1(n14174), .A2(n14172), .ZN(n14245) );
  OR2_X1 U14263 ( .A1(n14172), .A2(n14174), .ZN(n14243) );
  AND2_X1 U14264 ( .A1(n14246), .A2(n14247), .ZN(n14174) );
  NAND3_X1 U14265 ( .A1(b_4_), .A2(n14248), .A3(a_10_), .ZN(n14247) );
  NAND2_X1 U14266 ( .A1(n14170), .A2(n14168), .ZN(n14248) );
  OR2_X1 U14267 ( .A1(n14168), .A2(n14170), .ZN(n14246) );
  AND2_X1 U14268 ( .A1(n14249), .A2(n14250), .ZN(n14170) );
  NAND3_X1 U14269 ( .A1(a_11_), .A2(n14251), .A3(b_4_), .ZN(n14250) );
  NAND2_X1 U14270 ( .A1(n14166), .A2(n14164), .ZN(n14251) );
  OR2_X1 U14271 ( .A1(n14164), .A2(n14166), .ZN(n14249) );
  AND2_X1 U14272 ( .A1(n14252), .A2(n14253), .ZN(n14166) );
  NAND3_X1 U14273 ( .A1(b_4_), .A2(n14254), .A3(a_12_), .ZN(n14253) );
  NAND2_X1 U14274 ( .A1(n14162), .A2(n14161), .ZN(n14254) );
  OR2_X1 U14275 ( .A1(n14161), .A2(n14162), .ZN(n14252) );
  AND2_X1 U14276 ( .A1(n14255), .A2(n14256), .ZN(n14162) );
  NAND3_X1 U14277 ( .A1(b_4_), .A2(n14257), .A3(a_13_), .ZN(n14256) );
  NAND2_X1 U14278 ( .A1(n14158), .A2(n14157), .ZN(n14257) );
  OR2_X1 U14279 ( .A1(n14157), .A2(n14158), .ZN(n14255) );
  AND2_X1 U14280 ( .A1(n14258), .A2(n14259), .ZN(n14158) );
  NAND2_X1 U14281 ( .A1(n14155), .A2(n14260), .ZN(n14259) );
  NAND2_X1 U14282 ( .A1(n14154), .A2(n14153), .ZN(n14260) );
  NOR2_X1 U14283 ( .A1(n7962), .A2(n7964), .ZN(n14155) );
  OR2_X1 U14284 ( .A1(n14153), .A2(n14154), .ZN(n14258) );
  AND2_X1 U14285 ( .A1(n14261), .A2(n14262), .ZN(n14154) );
  NAND2_X1 U14286 ( .A1(n14150), .A2(n14263), .ZN(n14262) );
  NAND2_X1 U14287 ( .A1(n14151), .A2(n14149), .ZN(n14263) );
  NOR2_X1 U14288 ( .A1(n7667), .A2(n7964), .ZN(n14150) );
  OR2_X1 U14289 ( .A1(n14149), .A2(n14151), .ZN(n14261) );
  AND2_X1 U14290 ( .A1(n14264), .A2(n14265), .ZN(n14151) );
  NAND2_X1 U14291 ( .A1(n14147), .A2(n14266), .ZN(n14265) );
  OR2_X1 U14292 ( .A1(n14145), .A2(n14146), .ZN(n14266) );
  NOR2_X1 U14293 ( .A1(n8353), .A2(n7964), .ZN(n14147) );
  NAND2_X1 U14294 ( .A1(n14145), .A2(n14146), .ZN(n14264) );
  NAND2_X1 U14295 ( .A1(n14267), .A2(n14268), .ZN(n14146) );
  NAND2_X1 U14296 ( .A1(n14142), .A2(n14269), .ZN(n14268) );
  NAND2_X1 U14297 ( .A1(n14143), .A2(n14141), .ZN(n14269) );
  NOR2_X1 U14298 ( .A1(n7645), .A2(n7964), .ZN(n14142) );
  OR2_X1 U14299 ( .A1(n14141), .A2(n14143), .ZN(n14267) );
  AND2_X1 U14300 ( .A1(n14270), .A2(n14271), .ZN(n14143) );
  NAND2_X1 U14301 ( .A1(n14139), .A2(n14272), .ZN(n14271) );
  OR2_X1 U14302 ( .A1(n14137), .A2(n14138), .ZN(n14272) );
  NOR2_X1 U14303 ( .A1(n7960), .A2(n7964), .ZN(n14139) );
  NAND2_X1 U14304 ( .A1(n14137), .A2(n14138), .ZN(n14270) );
  NAND2_X1 U14305 ( .A1(n14273), .A2(n14274), .ZN(n14138) );
  NAND2_X1 U14306 ( .A1(n14135), .A2(n14275), .ZN(n14274) );
  NAND2_X1 U14307 ( .A1(n14134), .A2(n14133), .ZN(n14275) );
  NOR2_X1 U14308 ( .A1(n7958), .A2(n7964), .ZN(n14135) );
  OR2_X1 U14309 ( .A1(n14133), .A2(n14134), .ZN(n14273) );
  AND2_X1 U14310 ( .A1(n14276), .A2(n14277), .ZN(n14134) );
  NAND2_X1 U14311 ( .A1(n14131), .A2(n14278), .ZN(n14277) );
  OR2_X1 U14312 ( .A1(n14129), .A2(n14130), .ZN(n14278) );
  NOR2_X1 U14313 ( .A1(n7957), .A2(n7964), .ZN(n14131) );
  NAND2_X1 U14314 ( .A1(n14129), .A2(n14130), .ZN(n14276) );
  NAND2_X1 U14315 ( .A1(n14279), .A2(n14280), .ZN(n14130) );
  NAND2_X1 U14316 ( .A1(n14126), .A2(n14281), .ZN(n14280) );
  NAND2_X1 U14317 ( .A1(n14127), .A2(n14125), .ZN(n14281) );
  NOR2_X1 U14318 ( .A1(n7964), .A2(n7578), .ZN(n14126) );
  OR2_X1 U14319 ( .A1(n14125), .A2(n14127), .ZN(n14279) );
  AND2_X1 U14320 ( .A1(n14282), .A2(n14283), .ZN(n14127) );
  NAND2_X1 U14321 ( .A1(n14123), .A2(n14284), .ZN(n14283) );
  OR2_X1 U14322 ( .A1(n14120), .A2(n14122), .ZN(n14284) );
  NOR2_X1 U14323 ( .A1(n7568), .A2(n7964), .ZN(n14123) );
  NAND2_X1 U14324 ( .A1(n14120), .A2(n14122), .ZN(n14282) );
  NAND2_X1 U14325 ( .A1(n14285), .A2(n14286), .ZN(n14122) );
  NAND2_X1 U14326 ( .A1(n14119), .A2(n14287), .ZN(n14286) );
  OR2_X1 U14327 ( .A1(n14117), .A2(n14118), .ZN(n14287) );
  NOR2_X1 U14328 ( .A1(n7964), .A2(n7955), .ZN(n14119) );
  NAND2_X1 U14329 ( .A1(n14117), .A2(n14118), .ZN(n14285) );
  NAND2_X1 U14330 ( .A1(n14288), .A2(n14289), .ZN(n14118) );
  NAND2_X1 U14331 ( .A1(n14115), .A2(n14290), .ZN(n14289) );
  OR2_X1 U14332 ( .A1(n14113), .A2(n14114), .ZN(n14290) );
  NOR2_X1 U14333 ( .A1(n7954), .A2(n7964), .ZN(n14115) );
  NAND2_X1 U14334 ( .A1(n14113), .A2(n14114), .ZN(n14288) );
  NAND2_X1 U14335 ( .A1(n14291), .A2(n14292), .ZN(n14114) );
  NAND2_X1 U14336 ( .A1(n14111), .A2(n14293), .ZN(n14292) );
  OR2_X1 U14337 ( .A1(n14109), .A2(n14110), .ZN(n14293) );
  NOR2_X1 U14338 ( .A1(n7964), .A2(n7952), .ZN(n14111) );
  NAND2_X1 U14339 ( .A1(n14109), .A2(n14110), .ZN(n14291) );
  NAND2_X1 U14340 ( .A1(n14074), .A2(n14294), .ZN(n14110) );
  NAND2_X1 U14341 ( .A1(n14073), .A2(n14075), .ZN(n14294) );
  NAND2_X1 U14342 ( .A1(n14295), .A2(n14296), .ZN(n14075) );
  NAND2_X1 U14343 ( .A1(b_4_), .A2(a_26_), .ZN(n14296) );
  INV_X1 U14344 ( .A(n14297), .ZN(n14295) );
  XNOR2_X1 U14345 ( .A(n14298), .B(n14299), .ZN(n14073) );
  NAND2_X1 U14346 ( .A1(n14300), .A2(n14301), .ZN(n14298) );
  NAND2_X1 U14347 ( .A1(a_26_), .A2(n14297), .ZN(n14074) );
  NAND2_X1 U14348 ( .A1(n14082), .A2(n14302), .ZN(n14297) );
  NAND2_X1 U14349 ( .A1(n14081), .A2(n14083), .ZN(n14302) );
  NAND2_X1 U14350 ( .A1(n14303), .A2(n14304), .ZN(n14083) );
  NAND2_X1 U14351 ( .A1(b_4_), .A2(a_27_), .ZN(n14304) );
  INV_X1 U14352 ( .A(n14305), .ZN(n14303) );
  XNOR2_X1 U14353 ( .A(n14306), .B(n14307), .ZN(n14081) );
  XOR2_X1 U14354 ( .A(n14308), .B(n14309), .Z(n14306) );
  NAND2_X1 U14355 ( .A1(b_3_), .A2(a_28_), .ZN(n14308) );
  NAND2_X1 U14356 ( .A1(a_27_), .A2(n14305), .ZN(n14082) );
  NAND2_X1 U14357 ( .A1(n14310), .A2(n14311), .ZN(n14305) );
  NAND3_X1 U14358 ( .A1(a_28_), .A2(n14312), .A3(b_4_), .ZN(n14311) );
  NAND2_X1 U14359 ( .A1(n14091), .A2(n14089), .ZN(n14312) );
  OR2_X1 U14360 ( .A1(n14089), .A2(n14091), .ZN(n14310) );
  AND2_X1 U14361 ( .A1(n14313), .A2(n14314), .ZN(n14091) );
  NAND2_X1 U14362 ( .A1(n14105), .A2(n14315), .ZN(n14314) );
  OR2_X1 U14363 ( .A1(n14106), .A2(n14107), .ZN(n14315) );
  NOR2_X1 U14364 ( .A1(n7964), .A2(n7460), .ZN(n14105) );
  INV_X1 U14365 ( .A(b_4_), .ZN(n7964) );
  NAND2_X1 U14366 ( .A1(n14107), .A2(n14106), .ZN(n14313) );
  NAND2_X1 U14367 ( .A1(n14316), .A2(n14317), .ZN(n14106) );
  NAND2_X1 U14368 ( .A1(b_2_), .A2(n14318), .ZN(n14317) );
  NAND2_X1 U14369 ( .A1(n7441), .A2(n14319), .ZN(n14318) );
  NAND2_X1 U14370 ( .A1(a_31_), .A2(n7845), .ZN(n14319) );
  NAND2_X1 U14371 ( .A1(b_3_), .A2(n14320), .ZN(n14316) );
  NAND2_X1 U14372 ( .A1(n7445), .A2(n14321), .ZN(n14320) );
  NAND2_X1 U14373 ( .A1(a_30_), .A2(n7965), .ZN(n14321) );
  AND3_X1 U14374 ( .A1(b_4_), .A2(n7409), .A3(b_3_), .ZN(n14107) );
  XNOR2_X1 U14375 ( .A(n14322), .B(n14323), .ZN(n14089) );
  XOR2_X1 U14376 ( .A(n14324), .B(n14325), .Z(n14322) );
  XNOR2_X1 U14377 ( .A(n14326), .B(n14327), .ZN(n14109) );
  NAND2_X1 U14378 ( .A1(n14328), .A2(n14329), .ZN(n14326) );
  XNOR2_X1 U14379 ( .A(n14330), .B(n14331), .ZN(n14113) );
  NAND2_X1 U14380 ( .A1(n14332), .A2(n14333), .ZN(n14330) );
  XNOR2_X1 U14381 ( .A(n14334), .B(n14335), .ZN(n14117) );
  XNOR2_X1 U14382 ( .A(n14336), .B(n14337), .ZN(n14334) );
  NOR2_X1 U14383 ( .A1(n7954), .A2(n7845), .ZN(n14337) );
  XNOR2_X1 U14384 ( .A(n14338), .B(n14339), .ZN(n14120) );
  NAND2_X1 U14385 ( .A1(n14340), .A2(n14341), .ZN(n14338) );
  XNOR2_X1 U14386 ( .A(n14342), .B(n14343), .ZN(n14125) );
  XNOR2_X1 U14387 ( .A(n14344), .B(n14345), .ZN(n14342) );
  NAND2_X1 U14388 ( .A1(a_22_), .A2(b_3_), .ZN(n14344) );
  XNOR2_X1 U14389 ( .A(n14346), .B(n14347), .ZN(n14129) );
  NAND2_X1 U14390 ( .A1(n14348), .A2(n14349), .ZN(n14346) );
  XNOR2_X1 U14391 ( .A(n14350), .B(n14351), .ZN(n14133) );
  XNOR2_X1 U14392 ( .A(n14352), .B(n14353), .ZN(n14350) );
  NAND2_X1 U14393 ( .A1(a_20_), .A2(b_3_), .ZN(n14352) );
  XNOR2_X1 U14394 ( .A(n14354), .B(n14355), .ZN(n14137) );
  NAND2_X1 U14395 ( .A1(n14356), .A2(n14357), .ZN(n14354) );
  XNOR2_X1 U14396 ( .A(n14358), .B(n14359), .ZN(n14141) );
  XNOR2_X1 U14397 ( .A(n14360), .B(n14361), .ZN(n14358) );
  NAND2_X1 U14398 ( .A1(a_18_), .A2(b_3_), .ZN(n14360) );
  XNOR2_X1 U14399 ( .A(n14362), .B(n14363), .ZN(n14145) );
  NAND2_X1 U14400 ( .A1(n14364), .A2(n14365), .ZN(n14362) );
  XNOR2_X1 U14401 ( .A(n14366), .B(n14367), .ZN(n14149) );
  XNOR2_X1 U14402 ( .A(n14368), .B(n14369), .ZN(n14366) );
  NAND2_X1 U14403 ( .A1(a_16_), .A2(b_3_), .ZN(n14368) );
  XOR2_X1 U14404 ( .A(n14370), .B(n14371), .Z(n14153) );
  NAND2_X1 U14405 ( .A1(n14372), .A2(n14373), .ZN(n14370) );
  XNOR2_X1 U14406 ( .A(n14374), .B(n14375), .ZN(n14157) );
  XNOR2_X1 U14407 ( .A(n14376), .B(n14377), .ZN(n14374) );
  NAND2_X1 U14408 ( .A1(a_14_), .A2(b_3_), .ZN(n14376) );
  XOR2_X1 U14409 ( .A(n14378), .B(n14379), .Z(n14161) );
  NAND2_X1 U14410 ( .A1(n14380), .A2(n14381), .ZN(n14378) );
  XNOR2_X1 U14411 ( .A(n14382), .B(n14383), .ZN(n14164) );
  XNOR2_X1 U14412 ( .A(n14384), .B(n14385), .ZN(n14382) );
  NAND2_X1 U14413 ( .A1(a_12_), .A2(b_3_), .ZN(n14384) );
  XOR2_X1 U14414 ( .A(n14386), .B(n14387), .Z(n14168) );
  NAND2_X1 U14415 ( .A1(n14388), .A2(n14389), .ZN(n14386) );
  XNOR2_X1 U14416 ( .A(n14390), .B(n14391), .ZN(n14172) );
  XNOR2_X1 U14417 ( .A(n14392), .B(n14393), .ZN(n14390) );
  NAND2_X1 U14418 ( .A1(a_10_), .A2(b_3_), .ZN(n14392) );
  XOR2_X1 U14419 ( .A(n14394), .B(n14395), .Z(n14176) );
  NAND2_X1 U14420 ( .A1(n14396), .A2(n14397), .ZN(n14394) );
  XOR2_X1 U14421 ( .A(n14398), .B(n14399), .Z(n14181) );
  XNOR2_X1 U14422 ( .A(n14400), .B(n14401), .ZN(n14398) );
  NAND2_X1 U14423 ( .A1(a_8_), .A2(b_3_), .ZN(n14400) );
  XOR2_X1 U14424 ( .A(n14402), .B(n14403), .Z(n14008) );
  NAND2_X1 U14425 ( .A1(n14404), .A2(n14405), .ZN(n14402) );
  XOR2_X1 U14426 ( .A(n14406), .B(n14407), .Z(n14185) );
  XNOR2_X1 U14427 ( .A(n14408), .B(n14409), .ZN(n14406) );
  NAND2_X1 U14428 ( .A1(a_6_), .A2(b_3_), .ZN(n14408) );
  INV_X1 U14429 ( .A(n7830), .ZN(n14191) );
  NAND2_X1 U14430 ( .A1(a_4_), .A2(b_4_), .ZN(n7830) );
  XOR2_X1 U14431 ( .A(n14410), .B(n14411), .Z(n14193) );
  XNOR2_X1 U14432 ( .A(n14412), .B(n14413), .ZN(n14410) );
  NAND2_X1 U14433 ( .A1(a_4_), .A2(b_3_), .ZN(n14412) );
  XOR2_X1 U14434 ( .A(n14414), .B(n14415), .Z(n14197) );
  XOR2_X1 U14435 ( .A(n14416), .B(n7843), .Z(n14414) );
  XOR2_X1 U14436 ( .A(n14417), .B(n14418), .Z(n14201) );
  XNOR2_X1 U14437 ( .A(n14419), .B(n14420), .ZN(n14417) );
  NAND2_X1 U14438 ( .A1(a_2_), .A2(b_3_), .ZN(n14419) );
  XOR2_X1 U14439 ( .A(n14421), .B(n14422), .Z(n14205) );
  XOR2_X1 U14440 ( .A(n14423), .B(n14424), .Z(n14421) );
  NAND2_X1 U14441 ( .A1(n14425), .A2(n14426), .ZN(n14210) );
  XOR2_X1 U14442 ( .A(n14427), .B(n14428), .Z(n13987) );
  XOR2_X1 U14443 ( .A(n14429), .B(n14430), .Z(n14427) );
  NAND2_X1 U14444 ( .A1(n14431), .A2(n14211), .ZN(n7983) );
  INV_X1 U14445 ( .A(n14432), .ZN(n14211) );
  XNOR2_X1 U14446 ( .A(n8094), .B(n8095), .ZN(n14431) );
  NAND2_X1 U14447 ( .A1(n14432), .A2(n14433), .ZN(n7982) );
  XOR2_X1 U14448 ( .A(n8095), .B(n8094), .Z(n14433) );
  NOR2_X1 U14449 ( .A1(n14426), .A2(n14425), .ZN(n14432) );
  AND2_X1 U14450 ( .A1(n14434), .A2(n14435), .ZN(n14425) );
  NAND2_X1 U14451 ( .A1(n14429), .A2(n14436), .ZN(n14435) );
  OR2_X1 U14452 ( .A1(n14428), .A2(n14430), .ZN(n14436) );
  NOR2_X1 U14453 ( .A1(n7845), .A2(n8197), .ZN(n14429) );
  NAND2_X1 U14454 ( .A1(n14428), .A2(n14430), .ZN(n14434) );
  NAND2_X1 U14455 ( .A1(n14437), .A2(n14438), .ZN(n14430) );
  NAND2_X1 U14456 ( .A1(n14424), .A2(n14439), .ZN(n14438) );
  OR2_X1 U14457 ( .A1(n14422), .A2(n14423), .ZN(n14439) );
  NOR2_X1 U14458 ( .A1(n7872), .A2(n7845), .ZN(n14424) );
  NAND2_X1 U14459 ( .A1(n14422), .A2(n14423), .ZN(n14437) );
  NAND2_X1 U14460 ( .A1(n14440), .A2(n14441), .ZN(n14423) );
  NAND3_X1 U14461 ( .A1(b_3_), .A2(n14442), .A3(a_2_), .ZN(n14441) );
  OR2_X1 U14462 ( .A1(n14418), .A2(n14420), .ZN(n14442) );
  NAND2_X1 U14463 ( .A1(n14418), .A2(n14420), .ZN(n14440) );
  NAND2_X1 U14464 ( .A1(n14443), .A2(n14444), .ZN(n14420) );
  NAND2_X1 U14465 ( .A1(n14415), .A2(n14445), .ZN(n14444) );
  OR2_X1 U14466 ( .A1(n14416), .A2(n7843), .ZN(n14445) );
  XNOR2_X1 U14467 ( .A(n14446), .B(n14447), .ZN(n14415) );
  NAND2_X1 U14468 ( .A1(n14448), .A2(n14449), .ZN(n14446) );
  NAND2_X1 U14469 ( .A1(n7843), .A2(n14416), .ZN(n14443) );
  NAND2_X1 U14470 ( .A1(n14450), .A2(n14451), .ZN(n14416) );
  NAND3_X1 U14471 ( .A1(b_3_), .A2(n14452), .A3(a_4_), .ZN(n14451) );
  OR2_X1 U14472 ( .A1(n14411), .A2(n14413), .ZN(n14452) );
  NAND2_X1 U14473 ( .A1(n14411), .A2(n14413), .ZN(n14450) );
  NAND2_X1 U14474 ( .A1(n14229), .A2(n14453), .ZN(n14413) );
  NAND2_X1 U14475 ( .A1(n14228), .A2(n14230), .ZN(n14453) );
  NAND2_X1 U14476 ( .A1(n14454), .A2(n14455), .ZN(n14230) );
  NAND2_X1 U14477 ( .A1(a_5_), .A2(b_3_), .ZN(n14455) );
  INV_X1 U14478 ( .A(n14456), .ZN(n14454) );
  XNOR2_X1 U14479 ( .A(n14457), .B(n14458), .ZN(n14228) );
  NAND2_X1 U14480 ( .A1(n14459), .A2(n14460), .ZN(n14457) );
  NAND2_X1 U14481 ( .A1(a_5_), .A2(n14456), .ZN(n14229) );
  NAND2_X1 U14482 ( .A1(n14461), .A2(n14462), .ZN(n14456) );
  NAND3_X1 U14483 ( .A1(b_3_), .A2(n14463), .A3(a_6_), .ZN(n14462) );
  OR2_X1 U14484 ( .A1(n14407), .A2(n14409), .ZN(n14463) );
  NAND2_X1 U14485 ( .A1(n14407), .A2(n14409), .ZN(n14461) );
  NAND2_X1 U14486 ( .A1(n14404), .A2(n14464), .ZN(n14409) );
  NAND2_X1 U14487 ( .A1(n14403), .A2(n14405), .ZN(n14464) );
  NAND2_X1 U14488 ( .A1(n14465), .A2(n14466), .ZN(n14405) );
  NAND2_X1 U14489 ( .A1(a_7_), .A2(b_3_), .ZN(n14466) );
  INV_X1 U14490 ( .A(n14467), .ZN(n14465) );
  XNOR2_X1 U14491 ( .A(n14468), .B(n14469), .ZN(n14403) );
  NAND2_X1 U14492 ( .A1(n14470), .A2(n14471), .ZN(n14468) );
  NAND2_X1 U14493 ( .A1(a_7_), .A2(n14467), .ZN(n14404) );
  NAND2_X1 U14494 ( .A1(n14472), .A2(n14473), .ZN(n14467) );
  NAND3_X1 U14495 ( .A1(b_3_), .A2(n14474), .A3(a_8_), .ZN(n14473) );
  OR2_X1 U14496 ( .A1(n14399), .A2(n14401), .ZN(n14474) );
  NAND2_X1 U14497 ( .A1(n14399), .A2(n14401), .ZN(n14472) );
  NAND2_X1 U14498 ( .A1(n14396), .A2(n14475), .ZN(n14401) );
  NAND2_X1 U14499 ( .A1(n14395), .A2(n14397), .ZN(n14475) );
  NAND2_X1 U14500 ( .A1(n14476), .A2(n14477), .ZN(n14397) );
  NAND2_X1 U14501 ( .A1(a_9_), .A2(b_3_), .ZN(n14477) );
  INV_X1 U14502 ( .A(n14478), .ZN(n14476) );
  XNOR2_X1 U14503 ( .A(n14479), .B(n14480), .ZN(n14395) );
  NAND2_X1 U14504 ( .A1(n14481), .A2(n14482), .ZN(n14479) );
  NAND2_X1 U14505 ( .A1(a_9_), .A2(n14478), .ZN(n14396) );
  NAND2_X1 U14506 ( .A1(n14483), .A2(n14484), .ZN(n14478) );
  NAND3_X1 U14507 ( .A1(b_3_), .A2(n14485), .A3(a_10_), .ZN(n14484) );
  OR2_X1 U14508 ( .A1(n14391), .A2(n14393), .ZN(n14485) );
  NAND2_X1 U14509 ( .A1(n14391), .A2(n14393), .ZN(n14483) );
  NAND2_X1 U14510 ( .A1(n14388), .A2(n14486), .ZN(n14393) );
  NAND2_X1 U14511 ( .A1(n14387), .A2(n14389), .ZN(n14486) );
  NAND2_X1 U14512 ( .A1(n14487), .A2(n14488), .ZN(n14389) );
  NAND2_X1 U14513 ( .A1(b_3_), .A2(a_11_), .ZN(n14488) );
  INV_X1 U14514 ( .A(n14489), .ZN(n14487) );
  XNOR2_X1 U14515 ( .A(n14490), .B(n14491), .ZN(n14387) );
  NAND2_X1 U14516 ( .A1(n14492), .A2(n14493), .ZN(n14490) );
  NAND2_X1 U14517 ( .A1(a_11_), .A2(n14489), .ZN(n14388) );
  NAND2_X1 U14518 ( .A1(n14494), .A2(n14495), .ZN(n14489) );
  NAND3_X1 U14519 ( .A1(b_3_), .A2(n14496), .A3(a_12_), .ZN(n14495) );
  OR2_X1 U14520 ( .A1(n14383), .A2(n14385), .ZN(n14496) );
  NAND2_X1 U14521 ( .A1(n14383), .A2(n14385), .ZN(n14494) );
  NAND2_X1 U14522 ( .A1(n14380), .A2(n14497), .ZN(n14385) );
  NAND2_X1 U14523 ( .A1(n14379), .A2(n14381), .ZN(n14497) );
  NAND2_X1 U14524 ( .A1(n14498), .A2(n14499), .ZN(n14381) );
  NAND2_X1 U14525 ( .A1(a_13_), .A2(b_3_), .ZN(n14499) );
  INV_X1 U14526 ( .A(n14500), .ZN(n14498) );
  XNOR2_X1 U14527 ( .A(n14501), .B(n14502), .ZN(n14379) );
  NAND2_X1 U14528 ( .A1(n14503), .A2(n14504), .ZN(n14501) );
  NAND2_X1 U14529 ( .A1(a_13_), .A2(n14500), .ZN(n14380) );
  NAND2_X1 U14530 ( .A1(n14505), .A2(n14506), .ZN(n14500) );
  NAND3_X1 U14531 ( .A1(b_3_), .A2(n14507), .A3(a_14_), .ZN(n14506) );
  OR2_X1 U14532 ( .A1(n14375), .A2(n14377), .ZN(n14507) );
  NAND2_X1 U14533 ( .A1(n14375), .A2(n14377), .ZN(n14505) );
  NAND2_X1 U14534 ( .A1(n14372), .A2(n14508), .ZN(n14377) );
  NAND2_X1 U14535 ( .A1(n14371), .A2(n14373), .ZN(n14508) );
  NAND2_X1 U14536 ( .A1(n14509), .A2(n14510), .ZN(n14373) );
  NAND2_X1 U14537 ( .A1(a_15_), .A2(b_3_), .ZN(n14510) );
  INV_X1 U14538 ( .A(n14511), .ZN(n14509) );
  XNOR2_X1 U14539 ( .A(n14512), .B(n14513), .ZN(n14371) );
  NAND2_X1 U14540 ( .A1(n14514), .A2(n14515), .ZN(n14512) );
  NAND2_X1 U14541 ( .A1(a_15_), .A2(n14511), .ZN(n14372) );
  NAND2_X1 U14542 ( .A1(n14516), .A2(n14517), .ZN(n14511) );
  NAND3_X1 U14543 ( .A1(b_3_), .A2(n14518), .A3(a_16_), .ZN(n14517) );
  OR2_X1 U14544 ( .A1(n14367), .A2(n14369), .ZN(n14518) );
  NAND2_X1 U14545 ( .A1(n14367), .A2(n14369), .ZN(n14516) );
  NAND2_X1 U14546 ( .A1(n14364), .A2(n14519), .ZN(n14369) );
  NAND2_X1 U14547 ( .A1(n14363), .A2(n14365), .ZN(n14519) );
  NAND2_X1 U14548 ( .A1(n14520), .A2(n14521), .ZN(n14365) );
  NAND2_X1 U14549 ( .A1(a_17_), .A2(b_3_), .ZN(n14521) );
  INV_X1 U14550 ( .A(n14522), .ZN(n14520) );
  XNOR2_X1 U14551 ( .A(n14523), .B(n14524), .ZN(n14363) );
  XNOR2_X1 U14552 ( .A(n14525), .B(n14526), .ZN(n14524) );
  NAND2_X1 U14553 ( .A1(a_17_), .A2(n14522), .ZN(n14364) );
  NAND2_X1 U14554 ( .A1(n14527), .A2(n14528), .ZN(n14522) );
  NAND3_X1 U14555 ( .A1(b_3_), .A2(n14529), .A3(a_18_), .ZN(n14528) );
  OR2_X1 U14556 ( .A1(n14359), .A2(n14361), .ZN(n14529) );
  NAND2_X1 U14557 ( .A1(n14359), .A2(n14361), .ZN(n14527) );
  NAND2_X1 U14558 ( .A1(n14356), .A2(n14530), .ZN(n14361) );
  NAND2_X1 U14559 ( .A1(n14355), .A2(n14357), .ZN(n14530) );
  NAND2_X1 U14560 ( .A1(n14531), .A2(n14532), .ZN(n14357) );
  NAND2_X1 U14561 ( .A1(a_19_), .A2(b_3_), .ZN(n14532) );
  INV_X1 U14562 ( .A(n14533), .ZN(n14531) );
  XNOR2_X1 U14563 ( .A(n14534), .B(n14535), .ZN(n14355) );
  XNOR2_X1 U14564 ( .A(n14536), .B(n14537), .ZN(n14535) );
  NAND2_X1 U14565 ( .A1(a_19_), .A2(n14533), .ZN(n14356) );
  NAND2_X1 U14566 ( .A1(n14538), .A2(n14539), .ZN(n14533) );
  NAND3_X1 U14567 ( .A1(b_3_), .A2(n14540), .A3(a_20_), .ZN(n14539) );
  OR2_X1 U14568 ( .A1(n14351), .A2(n14353), .ZN(n14540) );
  NAND2_X1 U14569 ( .A1(n14351), .A2(n14353), .ZN(n14538) );
  NAND2_X1 U14570 ( .A1(n14348), .A2(n14541), .ZN(n14353) );
  NAND2_X1 U14571 ( .A1(n14347), .A2(n14349), .ZN(n14541) );
  NAND2_X1 U14572 ( .A1(n14542), .A2(n14543), .ZN(n14349) );
  NAND2_X1 U14573 ( .A1(b_3_), .A2(a_21_), .ZN(n14543) );
  INV_X1 U14574 ( .A(n14544), .ZN(n14542) );
  XNOR2_X1 U14575 ( .A(n14545), .B(n14546), .ZN(n14347) );
  XNOR2_X1 U14576 ( .A(n14547), .B(n14548), .ZN(n14546) );
  NAND2_X1 U14577 ( .A1(a_21_), .A2(n14544), .ZN(n14348) );
  NAND2_X1 U14578 ( .A1(n14549), .A2(n14550), .ZN(n14544) );
  NAND3_X1 U14579 ( .A1(b_3_), .A2(n14551), .A3(a_22_), .ZN(n14550) );
  OR2_X1 U14580 ( .A1(n14343), .A2(n14345), .ZN(n14551) );
  NAND2_X1 U14581 ( .A1(n14343), .A2(n14345), .ZN(n14549) );
  NAND2_X1 U14582 ( .A1(n14340), .A2(n14552), .ZN(n14345) );
  NAND2_X1 U14583 ( .A1(n14339), .A2(n14341), .ZN(n14552) );
  NAND2_X1 U14584 ( .A1(n14553), .A2(n14554), .ZN(n14341) );
  NAND2_X1 U14585 ( .A1(b_3_), .A2(a_23_), .ZN(n14554) );
  INV_X1 U14586 ( .A(n14555), .ZN(n14553) );
  XNOR2_X1 U14587 ( .A(n14556), .B(n14557), .ZN(n14339) );
  XNOR2_X1 U14588 ( .A(n14558), .B(n14559), .ZN(n14557) );
  NAND2_X1 U14589 ( .A1(a_23_), .A2(n14555), .ZN(n14340) );
  NAND2_X1 U14590 ( .A1(n14560), .A2(n14561), .ZN(n14555) );
  NAND3_X1 U14591 ( .A1(a_24_), .A2(n14562), .A3(b_3_), .ZN(n14561) );
  NAND2_X1 U14592 ( .A1(n14336), .A2(n14335), .ZN(n14562) );
  OR2_X1 U14593 ( .A1(n14335), .A2(n14336), .ZN(n14560) );
  AND2_X1 U14594 ( .A1(n14332), .A2(n14563), .ZN(n14336) );
  NAND2_X1 U14595 ( .A1(n14331), .A2(n14333), .ZN(n14563) );
  NAND2_X1 U14596 ( .A1(n14564), .A2(n14565), .ZN(n14333) );
  NAND2_X1 U14597 ( .A1(b_3_), .A2(a_25_), .ZN(n14565) );
  INV_X1 U14598 ( .A(n14566), .ZN(n14564) );
  XNOR2_X1 U14599 ( .A(n14567), .B(n14568), .ZN(n14331) );
  XOR2_X1 U14600 ( .A(n14569), .B(n14570), .Z(n14567) );
  NAND2_X1 U14601 ( .A1(b_2_), .A2(a_26_), .ZN(n14569) );
  NAND2_X1 U14602 ( .A1(a_25_), .A2(n14566), .ZN(n14332) );
  NAND2_X1 U14603 ( .A1(n14328), .A2(n14571), .ZN(n14566) );
  NAND2_X1 U14604 ( .A1(n14327), .A2(n14329), .ZN(n14571) );
  NAND2_X1 U14605 ( .A1(n14572), .A2(n14573), .ZN(n14329) );
  NAND2_X1 U14606 ( .A1(b_3_), .A2(a_26_), .ZN(n14573) );
  INV_X1 U14607 ( .A(n14574), .ZN(n14572) );
  XNOR2_X1 U14608 ( .A(n14575), .B(n14576), .ZN(n14327) );
  XNOR2_X1 U14609 ( .A(n14577), .B(n14578), .ZN(n14576) );
  NAND2_X1 U14610 ( .A1(a_26_), .A2(n14574), .ZN(n14328) );
  NAND2_X1 U14611 ( .A1(n14300), .A2(n14579), .ZN(n14574) );
  NAND2_X1 U14612 ( .A1(n14299), .A2(n14301), .ZN(n14579) );
  NAND2_X1 U14613 ( .A1(n14580), .A2(n14581), .ZN(n14301) );
  NAND2_X1 U14614 ( .A1(b_3_), .A2(a_27_), .ZN(n14581) );
  INV_X1 U14615 ( .A(n14582), .ZN(n14580) );
  XOR2_X1 U14616 ( .A(n14583), .B(n14584), .Z(n14299) );
  XNOR2_X1 U14617 ( .A(n14585), .B(n14586), .ZN(n14583) );
  NAND2_X1 U14618 ( .A1(b_2_), .A2(a_28_), .ZN(n14585) );
  NAND2_X1 U14619 ( .A1(a_27_), .A2(n14582), .ZN(n14300) );
  NAND2_X1 U14620 ( .A1(n14587), .A2(n14588), .ZN(n14582) );
  NAND3_X1 U14621 ( .A1(a_28_), .A2(n14589), .A3(b_3_), .ZN(n14588) );
  NAND2_X1 U14622 ( .A1(n14309), .A2(n14307), .ZN(n14589) );
  OR2_X1 U14623 ( .A1(n14307), .A2(n14309), .ZN(n14587) );
  AND2_X1 U14624 ( .A1(n14590), .A2(n14591), .ZN(n14309) );
  NAND2_X1 U14625 ( .A1(n14323), .A2(n14592), .ZN(n14591) );
  OR2_X1 U14626 ( .A1(n14324), .A2(n14325), .ZN(n14592) );
  NOR2_X1 U14627 ( .A1(n7845), .A2(n7460), .ZN(n14323) );
  INV_X1 U14628 ( .A(b_3_), .ZN(n7845) );
  NAND2_X1 U14629 ( .A1(n14325), .A2(n14324), .ZN(n14590) );
  NAND2_X1 U14630 ( .A1(n14593), .A2(n14594), .ZN(n14324) );
  NAND2_X1 U14631 ( .A1(b_1_), .A2(n14595), .ZN(n14594) );
  NAND2_X1 U14632 ( .A1(n7441), .A2(n14596), .ZN(n14595) );
  NAND2_X1 U14633 ( .A1(a_31_), .A2(n7965), .ZN(n14596) );
  NAND2_X1 U14634 ( .A1(b_2_), .A2(n14597), .ZN(n14593) );
  NAND2_X1 U14635 ( .A1(n7445), .A2(n14598), .ZN(n14597) );
  NAND2_X1 U14636 ( .A1(a_30_), .A2(n14599), .ZN(n14598) );
  AND3_X1 U14637 ( .A1(b_3_), .A2(n7409), .A3(b_2_), .ZN(n14325) );
  XNOR2_X1 U14638 ( .A(n14600), .B(n14601), .ZN(n14307) );
  NOR2_X1 U14639 ( .A1(n7460), .A2(n7965), .ZN(n14601) );
  XOR2_X1 U14640 ( .A(n14602), .B(n14603), .Z(n14600) );
  XOR2_X1 U14641 ( .A(n14604), .B(n14605), .Z(n14335) );
  NAND2_X1 U14642 ( .A1(n14606), .A2(n14607), .ZN(n14604) );
  XNOR2_X1 U14643 ( .A(n14608), .B(n14609), .ZN(n14343) );
  XOR2_X1 U14644 ( .A(n14610), .B(n14611), .Z(n14609) );
  NAND2_X1 U14645 ( .A1(b_2_), .A2(a_23_), .ZN(n14611) );
  XNOR2_X1 U14646 ( .A(n14612), .B(n14613), .ZN(n14351) );
  XOR2_X1 U14647 ( .A(n14614), .B(n14615), .Z(n14612) );
  NAND2_X1 U14648 ( .A1(b_2_), .A2(a_21_), .ZN(n14614) );
  XNOR2_X1 U14649 ( .A(n14616), .B(n14617), .ZN(n14359) );
  XOR2_X1 U14650 ( .A(n14618), .B(n14619), .Z(n14616) );
  NAND2_X1 U14651 ( .A1(a_19_), .A2(b_2_), .ZN(n14618) );
  XNOR2_X1 U14652 ( .A(n14620), .B(n14621), .ZN(n14367) );
  XNOR2_X1 U14653 ( .A(n14622), .B(n14623), .ZN(n14620) );
  XOR2_X1 U14654 ( .A(n14624), .B(n14625), .Z(n14375) );
  XOR2_X1 U14655 ( .A(n14626), .B(n14627), .Z(n14624) );
  XOR2_X1 U14656 ( .A(n14628), .B(n14629), .Z(n14383) );
  XOR2_X1 U14657 ( .A(n14630), .B(n14631), .Z(n14628) );
  XOR2_X1 U14658 ( .A(n14632), .B(n14633), .Z(n14391) );
  XOR2_X1 U14659 ( .A(n14634), .B(n14635), .Z(n14632) );
  XOR2_X1 U14660 ( .A(n14636), .B(n14637), .Z(n14399) );
  XOR2_X1 U14661 ( .A(n14638), .B(n14639), .Z(n14636) );
  XOR2_X1 U14662 ( .A(n14640), .B(n14641), .Z(n14407) );
  XOR2_X1 U14663 ( .A(n14642), .B(n14643), .Z(n14640) );
  XOR2_X1 U14664 ( .A(n14644), .B(n14645), .Z(n14411) );
  XOR2_X1 U14665 ( .A(n14646), .B(n14647), .Z(n14644) );
  INV_X1 U14666 ( .A(n7891), .ZN(n7843) );
  NAND2_X1 U14667 ( .A1(a_3_), .A2(b_3_), .ZN(n7891) );
  XOR2_X1 U14668 ( .A(n14648), .B(n14649), .Z(n14418) );
  XOR2_X1 U14669 ( .A(n14650), .B(n14651), .Z(n14648) );
  XNOR2_X1 U14670 ( .A(n14652), .B(n14653), .ZN(n14422) );
  XOR2_X1 U14671 ( .A(n14654), .B(n7859), .Z(n14653) );
  XOR2_X1 U14672 ( .A(n14655), .B(n14656), .Z(n14428) );
  XOR2_X1 U14673 ( .A(n14657), .B(n14658), .Z(n14655) );
  XOR2_X1 U14674 ( .A(n14659), .B(n14660), .Z(n14426) );
  NAND2_X1 U14675 ( .A1(n14661), .A2(n14662), .ZN(n14659) );
  INV_X1 U14676 ( .A(n8037), .ZN(n8090) );
  NAND4_X1 U14677 ( .A1(n7888), .A2(n8096), .A3(n8094), .A4(n8095), .ZN(n8037)
         );
  NAND2_X1 U14678 ( .A1(n14661), .A2(n14663), .ZN(n8095) );
  NAND2_X1 U14679 ( .A1(n14660), .A2(n14662), .ZN(n14663) );
  NAND2_X1 U14680 ( .A1(n14664), .A2(n14665), .ZN(n14662) );
  NAND2_X1 U14681 ( .A1(b_2_), .A2(a_0_), .ZN(n14665) );
  INV_X1 U14682 ( .A(n14666), .ZN(n14664) );
  XNOR2_X1 U14683 ( .A(n14667), .B(n14668), .ZN(n14660) );
  XNOR2_X1 U14684 ( .A(n7878), .B(n14669), .ZN(n14668) );
  NAND2_X1 U14685 ( .A1(a_0_), .A2(n14666), .ZN(n14661) );
  NAND2_X1 U14686 ( .A1(n14670), .A2(n14671), .ZN(n14666) );
  NAND2_X1 U14687 ( .A1(n14657), .A2(n14672), .ZN(n14671) );
  OR2_X1 U14688 ( .A1(n14658), .A2(n14656), .ZN(n14672) );
  NOR2_X1 U14689 ( .A1(n7872), .A2(n7965), .ZN(n14657) );
  NAND2_X1 U14690 ( .A1(n14656), .A2(n14658), .ZN(n14670) );
  NAND2_X1 U14691 ( .A1(n14673), .A2(n14674), .ZN(n14658) );
  NAND2_X1 U14692 ( .A1(n14652), .A2(n14675), .ZN(n14674) );
  OR2_X1 U14693 ( .A1(n14654), .A2(n14676), .ZN(n14675) );
  XOR2_X1 U14694 ( .A(n14677), .B(n14678), .Z(n14652) );
  XNOR2_X1 U14695 ( .A(n14679), .B(n14680), .ZN(n14678) );
  NAND2_X1 U14696 ( .A1(a_3_), .A2(b_1_), .ZN(n14677) );
  NAND2_X1 U14697 ( .A1(n14676), .A2(n14654), .ZN(n14673) );
  NAND2_X1 U14698 ( .A1(n14681), .A2(n14682), .ZN(n14654) );
  NAND2_X1 U14699 ( .A1(n14650), .A2(n14683), .ZN(n14682) );
  OR2_X1 U14700 ( .A1(n14651), .A2(n14649), .ZN(n14683) );
  NOR2_X1 U14701 ( .A1(n7852), .A2(n7965), .ZN(n14650) );
  NAND2_X1 U14702 ( .A1(n14649), .A2(n14651), .ZN(n14681) );
  NAND2_X1 U14703 ( .A1(n14448), .A2(n14684), .ZN(n14651) );
  NAND2_X1 U14704 ( .A1(n14447), .A2(n14449), .ZN(n14684) );
  NAND2_X1 U14705 ( .A1(n14685), .A2(n14686), .ZN(n14449) );
  NAND2_X1 U14706 ( .A1(a_4_), .A2(b_2_), .ZN(n14686) );
  INV_X1 U14707 ( .A(n14687), .ZN(n14685) );
  XOR2_X1 U14708 ( .A(n14688), .B(n14689), .Z(n14447) );
  XNOR2_X1 U14709 ( .A(n14690), .B(n14691), .ZN(n14689) );
  NAND2_X1 U14710 ( .A1(a_5_), .A2(b_1_), .ZN(n14688) );
  NAND2_X1 U14711 ( .A1(a_4_), .A2(n14687), .ZN(n14448) );
  NAND2_X1 U14712 ( .A1(n14692), .A2(n14693), .ZN(n14687) );
  NAND2_X1 U14713 ( .A1(n14646), .A2(n14694), .ZN(n14693) );
  OR2_X1 U14714 ( .A1(n14647), .A2(n14645), .ZN(n14694) );
  NOR2_X1 U14715 ( .A1(n7823), .A2(n7965), .ZN(n14646) );
  NAND2_X1 U14716 ( .A1(n14645), .A2(n14647), .ZN(n14692) );
  NAND2_X1 U14717 ( .A1(n14459), .A2(n14695), .ZN(n14647) );
  NAND2_X1 U14718 ( .A1(n14458), .A2(n14460), .ZN(n14695) );
  NAND2_X1 U14719 ( .A1(n14696), .A2(n14697), .ZN(n14460) );
  NAND2_X1 U14720 ( .A1(a_6_), .A2(b_2_), .ZN(n14697) );
  INV_X1 U14721 ( .A(n14698), .ZN(n14696) );
  XOR2_X1 U14722 ( .A(n14699), .B(n14700), .Z(n14458) );
  XNOR2_X1 U14723 ( .A(n14701), .B(n14702), .ZN(n14700) );
  NAND2_X1 U14724 ( .A1(a_7_), .A2(b_1_), .ZN(n14699) );
  NAND2_X1 U14725 ( .A1(a_6_), .A2(n14698), .ZN(n14459) );
  NAND2_X1 U14726 ( .A1(n14703), .A2(n14704), .ZN(n14698) );
  NAND2_X1 U14727 ( .A1(n14642), .A2(n14705), .ZN(n14704) );
  OR2_X1 U14728 ( .A1(n14643), .A2(n14641), .ZN(n14705) );
  NOR2_X1 U14729 ( .A1(n7787), .A2(n7965), .ZN(n14642) );
  NAND2_X1 U14730 ( .A1(n14641), .A2(n14643), .ZN(n14703) );
  NAND2_X1 U14731 ( .A1(n14470), .A2(n14706), .ZN(n14643) );
  NAND2_X1 U14732 ( .A1(n14469), .A2(n14471), .ZN(n14706) );
  NAND2_X1 U14733 ( .A1(n14707), .A2(n14708), .ZN(n14471) );
  NAND2_X1 U14734 ( .A1(a_8_), .A2(b_2_), .ZN(n14708) );
  INV_X1 U14735 ( .A(n14709), .ZN(n14707) );
  XOR2_X1 U14736 ( .A(n14710), .B(n14711), .Z(n14469) );
  XNOR2_X1 U14737 ( .A(n14712), .B(n14713), .ZN(n14711) );
  NAND2_X1 U14738 ( .A1(a_9_), .A2(b_1_), .ZN(n14710) );
  NAND2_X1 U14739 ( .A1(a_8_), .A2(n14709), .ZN(n14470) );
  NAND2_X1 U14740 ( .A1(n14714), .A2(n14715), .ZN(n14709) );
  NAND2_X1 U14741 ( .A1(n14638), .A2(n14716), .ZN(n14715) );
  OR2_X1 U14742 ( .A1(n14639), .A2(n14637), .ZN(n14716) );
  NOR2_X1 U14743 ( .A1(n7753), .A2(n7965), .ZN(n14638) );
  NAND2_X1 U14744 ( .A1(n14637), .A2(n14639), .ZN(n14714) );
  NAND2_X1 U14745 ( .A1(n14481), .A2(n14717), .ZN(n14639) );
  NAND2_X1 U14746 ( .A1(n14480), .A2(n14482), .ZN(n14717) );
  NAND2_X1 U14747 ( .A1(n14718), .A2(n14719), .ZN(n14482) );
  NAND2_X1 U14748 ( .A1(a_10_), .A2(b_2_), .ZN(n14719) );
  INV_X1 U14749 ( .A(n14720), .ZN(n14718) );
  XOR2_X1 U14750 ( .A(n14721), .B(n14722), .Z(n14480) );
  XNOR2_X1 U14751 ( .A(n14723), .B(n14724), .ZN(n14722) );
  NAND2_X1 U14752 ( .A1(b_1_), .A2(a_11_), .ZN(n14721) );
  NAND2_X1 U14753 ( .A1(a_10_), .A2(n14720), .ZN(n14481) );
  NAND2_X1 U14754 ( .A1(n14725), .A2(n14726), .ZN(n14720) );
  NAND2_X1 U14755 ( .A1(n14634), .A2(n14727), .ZN(n14726) );
  OR2_X1 U14756 ( .A1(n14635), .A2(n14633), .ZN(n14727) );
  NOR2_X1 U14757 ( .A1(n7965), .A2(n7724), .ZN(n14634) );
  NAND2_X1 U14758 ( .A1(n14633), .A2(n14635), .ZN(n14725) );
  NAND2_X1 U14759 ( .A1(n14492), .A2(n14728), .ZN(n14635) );
  NAND2_X1 U14760 ( .A1(n14491), .A2(n14493), .ZN(n14728) );
  NAND2_X1 U14761 ( .A1(n14729), .A2(n14730), .ZN(n14493) );
  NAND2_X1 U14762 ( .A1(a_12_), .A2(b_2_), .ZN(n14730) );
  INV_X1 U14763 ( .A(n14731), .ZN(n14729) );
  XOR2_X1 U14764 ( .A(n14732), .B(n14733), .Z(n14491) );
  XNOR2_X1 U14765 ( .A(n14734), .B(n14735), .ZN(n14733) );
  NAND2_X1 U14766 ( .A1(a_13_), .A2(b_1_), .ZN(n14732) );
  NAND2_X1 U14767 ( .A1(a_12_), .A2(n14731), .ZN(n14492) );
  NAND2_X1 U14768 ( .A1(n14736), .A2(n14737), .ZN(n14731) );
  NAND2_X1 U14769 ( .A1(n14630), .A2(n14738), .ZN(n14737) );
  OR2_X1 U14770 ( .A1(n14631), .A2(n14629), .ZN(n14738) );
  NOR2_X1 U14771 ( .A1(n7702), .A2(n7965), .ZN(n14630) );
  NAND2_X1 U14772 ( .A1(n14629), .A2(n14631), .ZN(n14736) );
  NAND2_X1 U14773 ( .A1(n14503), .A2(n14739), .ZN(n14631) );
  NAND2_X1 U14774 ( .A1(n14502), .A2(n14504), .ZN(n14739) );
  NAND2_X1 U14775 ( .A1(n14740), .A2(n14741), .ZN(n14504) );
  NAND2_X1 U14776 ( .A1(a_14_), .A2(b_2_), .ZN(n14741) );
  INV_X1 U14777 ( .A(n14742), .ZN(n14740) );
  XOR2_X1 U14778 ( .A(n14743), .B(n14744), .Z(n14502) );
  XNOR2_X1 U14779 ( .A(n14745), .B(n14746), .ZN(n14744) );
  NAND2_X1 U14780 ( .A1(a_15_), .A2(b_1_), .ZN(n14743) );
  NAND2_X1 U14781 ( .A1(a_14_), .A2(n14742), .ZN(n14503) );
  NAND2_X1 U14782 ( .A1(n14747), .A2(n14748), .ZN(n14742) );
  NAND2_X1 U14783 ( .A1(n14626), .A2(n14749), .ZN(n14748) );
  OR2_X1 U14784 ( .A1(n14627), .A2(n14625), .ZN(n14749) );
  NOR2_X1 U14785 ( .A1(n7667), .A2(n7965), .ZN(n14626) );
  NAND2_X1 U14786 ( .A1(n14625), .A2(n14627), .ZN(n14747) );
  NAND2_X1 U14787 ( .A1(n14514), .A2(n14750), .ZN(n14627) );
  NAND2_X1 U14788 ( .A1(n14513), .A2(n14515), .ZN(n14750) );
  NAND2_X1 U14789 ( .A1(n14751), .A2(n14752), .ZN(n14515) );
  NAND2_X1 U14790 ( .A1(a_16_), .A2(b_2_), .ZN(n14752) );
  INV_X1 U14791 ( .A(n14753), .ZN(n14751) );
  XOR2_X1 U14792 ( .A(n14754), .B(n14755), .Z(n14513) );
  XNOR2_X1 U14793 ( .A(n14756), .B(n14757), .ZN(n14755) );
  NAND2_X1 U14794 ( .A1(a_17_), .A2(b_1_), .ZN(n14754) );
  NAND2_X1 U14795 ( .A1(a_16_), .A2(n14753), .ZN(n14514) );
  NAND2_X1 U14796 ( .A1(n14758), .A2(n14759), .ZN(n14753) );
  NAND2_X1 U14797 ( .A1(n14622), .A2(n14760), .ZN(n14759) );
  NAND2_X1 U14798 ( .A1(n14623), .A2(n14621), .ZN(n14760) );
  NOR2_X1 U14799 ( .A1(n7645), .A2(n7965), .ZN(n14622) );
  OR2_X1 U14800 ( .A1(n14621), .A2(n14623), .ZN(n14758) );
  AND2_X1 U14801 ( .A1(n14761), .A2(n14762), .ZN(n14623) );
  NAND2_X1 U14802 ( .A1(n14526), .A2(n14763), .ZN(n14762) );
  OR2_X1 U14803 ( .A1(n14525), .A2(n14523), .ZN(n14763) );
  NOR2_X1 U14804 ( .A1(n7960), .A2(n7965), .ZN(n14526) );
  NAND2_X1 U14805 ( .A1(n14523), .A2(n14525), .ZN(n14761) );
  NAND2_X1 U14806 ( .A1(n14764), .A2(n14765), .ZN(n14525) );
  NAND3_X1 U14807 ( .A1(b_2_), .A2(n14766), .A3(a_19_), .ZN(n14765) );
  NAND2_X1 U14808 ( .A1(n14619), .A2(n14617), .ZN(n14766) );
  OR2_X1 U14809 ( .A1(n14617), .A2(n14619), .ZN(n14764) );
  AND2_X1 U14810 ( .A1(n14767), .A2(n14768), .ZN(n14619) );
  NAND2_X1 U14811 ( .A1(n14537), .A2(n14769), .ZN(n14768) );
  OR2_X1 U14812 ( .A1(n14536), .A2(n14534), .ZN(n14769) );
  NOR2_X1 U14813 ( .A1(n7957), .A2(n7965), .ZN(n14537) );
  NAND2_X1 U14814 ( .A1(n14534), .A2(n14536), .ZN(n14767) );
  NAND2_X1 U14815 ( .A1(n14770), .A2(n14771), .ZN(n14536) );
  NAND3_X1 U14816 ( .A1(a_21_), .A2(n14772), .A3(b_2_), .ZN(n14771) );
  NAND2_X1 U14817 ( .A1(n14615), .A2(n14613), .ZN(n14772) );
  OR2_X1 U14818 ( .A1(n14613), .A2(n14615), .ZN(n14770) );
  AND2_X1 U14819 ( .A1(n14773), .A2(n14774), .ZN(n14615) );
  NAND2_X1 U14820 ( .A1(n14548), .A2(n14775), .ZN(n14774) );
  OR2_X1 U14821 ( .A1(n14547), .A2(n14545), .ZN(n14775) );
  NOR2_X1 U14822 ( .A1(n7568), .A2(n7965), .ZN(n14548) );
  INV_X1 U14823 ( .A(a_22_), .ZN(n7568) );
  NAND2_X1 U14824 ( .A1(n14545), .A2(n14547), .ZN(n14773) );
  NAND2_X1 U14825 ( .A1(n14776), .A2(n14777), .ZN(n14547) );
  NAND3_X1 U14826 ( .A1(a_23_), .A2(n14778), .A3(b_2_), .ZN(n14777) );
  OR2_X1 U14827 ( .A1(n14610), .A2(n14608), .ZN(n14778) );
  NAND2_X1 U14828 ( .A1(n14608), .A2(n14610), .ZN(n14776) );
  NAND2_X1 U14829 ( .A1(n14779), .A2(n14780), .ZN(n14610) );
  NAND2_X1 U14830 ( .A1(n14559), .A2(n14781), .ZN(n14780) );
  OR2_X1 U14831 ( .A1(n14558), .A2(n14556), .ZN(n14781) );
  NOR2_X1 U14832 ( .A1(n7965), .A2(n7954), .ZN(n14559) );
  NAND2_X1 U14833 ( .A1(n14556), .A2(n14558), .ZN(n14779) );
  NAND2_X1 U14834 ( .A1(n14606), .A2(n14782), .ZN(n14558) );
  NAND2_X1 U14835 ( .A1(n14605), .A2(n14607), .ZN(n14782) );
  NAND2_X1 U14836 ( .A1(n14783), .A2(n14784), .ZN(n14607) );
  NAND2_X1 U14837 ( .A1(b_2_), .A2(a_25_), .ZN(n14784) );
  INV_X1 U14838 ( .A(n14785), .ZN(n14783) );
  XOR2_X1 U14839 ( .A(n14786), .B(n14787), .Z(n14605) );
  NOR2_X1 U14840 ( .A1(n7950), .A2(n14788), .ZN(n14787) );
  XOR2_X1 U14841 ( .A(n14789), .B(n14790), .Z(n14786) );
  NAND2_X1 U14842 ( .A1(a_25_), .A2(n14785), .ZN(n14606) );
  NAND2_X1 U14843 ( .A1(n14791), .A2(n14792), .ZN(n14785) );
  NAND3_X1 U14844 ( .A1(a_26_), .A2(n14793), .A3(b_2_), .ZN(n14792) );
  NAND2_X1 U14845 ( .A1(n14570), .A2(n14568), .ZN(n14793) );
  OR2_X1 U14846 ( .A1(n14568), .A2(n14570), .ZN(n14791) );
  AND2_X1 U14847 ( .A1(n14794), .A2(n14795), .ZN(n14570) );
  NAND2_X1 U14848 ( .A1(n14578), .A2(n14796), .ZN(n14795) );
  OR2_X1 U14849 ( .A1(n14577), .A2(n14575), .ZN(n14796) );
  NOR2_X1 U14850 ( .A1(n7965), .A2(n7950), .ZN(n14578) );
  INV_X1 U14851 ( .A(b_2_), .ZN(n7965) );
  NAND2_X1 U14852 ( .A1(n14575), .A2(n14577), .ZN(n14794) );
  NAND2_X1 U14853 ( .A1(n14797), .A2(n14798), .ZN(n14577) );
  NAND3_X1 U14854 ( .A1(a_28_), .A2(n14799), .A3(b_2_), .ZN(n14798) );
  OR2_X1 U14855 ( .A1(n14584), .A2(n14586), .ZN(n14799) );
  NAND2_X1 U14856 ( .A1(n14584), .A2(n14586), .ZN(n14797) );
  NAND2_X1 U14857 ( .A1(n14800), .A2(n14801), .ZN(n14586) );
  NAND3_X1 U14858 ( .A1(a_29_), .A2(n14802), .A3(b_2_), .ZN(n14801) );
  OR2_X1 U14859 ( .A1(n14602), .A2(n14603), .ZN(n14802) );
  NAND2_X1 U14860 ( .A1(n14603), .A2(n14602), .ZN(n14800) );
  NAND2_X1 U14861 ( .A1(n14803), .A2(n14804), .ZN(n14602) );
  NAND2_X1 U14862 ( .A1(b_0_), .A2(n14805), .ZN(n14804) );
  NAND2_X1 U14863 ( .A1(n7441), .A2(n14806), .ZN(n14805) );
  NAND2_X1 U14864 ( .A1(a_31_), .A2(n14599), .ZN(n14806) );
  NAND2_X1 U14865 ( .A1(b_1_), .A2(n14807), .ZN(n14803) );
  NAND2_X1 U14866 ( .A1(n7445), .A2(n14808), .ZN(n14807) );
  NAND2_X1 U14867 ( .A1(a_30_), .A2(n14788), .ZN(n14808) );
  AND3_X1 U14868 ( .A1(b_2_), .A2(n7409), .A3(b_1_), .ZN(n14603) );
  XNOR2_X1 U14869 ( .A(n14809), .B(n14810), .ZN(n14584) );
  NOR2_X1 U14870 ( .A1(n7450), .A2(n14788), .ZN(n14810) );
  XOR2_X1 U14871 ( .A(n14811), .B(n14812), .Z(n14809) );
  XOR2_X1 U14872 ( .A(n14813), .B(n14814), .Z(n14575) );
  XNOR2_X1 U14873 ( .A(n14815), .B(n14816), .ZN(n14814) );
  NAND2_X1 U14874 ( .A1(b_0_), .A2(a_29_), .ZN(n14813) );
  XNOR2_X1 U14875 ( .A(n14817), .B(n14818), .ZN(n14568) );
  XNOR2_X1 U14876 ( .A(n14819), .B(n14820), .ZN(n14818) );
  NAND2_X1 U14877 ( .A1(b_0_), .A2(a_28_), .ZN(n14817) );
  XOR2_X1 U14878 ( .A(n14821), .B(n14822), .Z(n14556) );
  XNOR2_X1 U14879 ( .A(n14823), .B(n14824), .ZN(n14822) );
  NAND2_X1 U14880 ( .A1(b_0_), .A2(a_26_), .ZN(n14821) );
  XOR2_X1 U14881 ( .A(n14825), .B(n14826), .Z(n14608) );
  NOR2_X1 U14882 ( .A1(n7952), .A2(n14788), .ZN(n14826) );
  XOR2_X1 U14883 ( .A(n14827), .B(n14828), .Z(n14825) );
  XOR2_X1 U14884 ( .A(n14829), .B(n14830), .Z(n14545) );
  XNOR2_X1 U14885 ( .A(n14831), .B(n14832), .ZN(n14830) );
  NAND2_X1 U14886 ( .A1(b_0_), .A2(a_24_), .ZN(n14829) );
  XNOR2_X1 U14887 ( .A(n14833), .B(n14834), .ZN(n14613) );
  NOR2_X1 U14888 ( .A1(n7955), .A2(n14788), .ZN(n14834) );
  XOR2_X1 U14889 ( .A(n14835), .B(n14836), .Z(n14833) );
  XOR2_X1 U14890 ( .A(n14837), .B(n14838), .Z(n14534) );
  XNOR2_X1 U14891 ( .A(n14839), .B(n14840), .ZN(n14838) );
  NAND2_X1 U14892 ( .A1(b_0_), .A2(a_22_), .ZN(n14837) );
  XNOR2_X1 U14893 ( .A(n14841), .B(n14842), .ZN(n14617) );
  NOR2_X1 U14894 ( .A1(n7578), .A2(n14788), .ZN(n14842) );
  XOR2_X1 U14895 ( .A(n14843), .B(n14844), .Z(n14841) );
  XOR2_X1 U14896 ( .A(n14845), .B(n14846), .Z(n14523) );
  XNOR2_X1 U14897 ( .A(n14847), .B(n14848), .ZN(n14846) );
  NAND2_X1 U14898 ( .A1(a_20_), .A2(b_0_), .ZN(n14845) );
  XNOR2_X1 U14899 ( .A(n14849), .B(n14850), .ZN(n14621) );
  NOR2_X1 U14900 ( .A1(n14788), .A2(n7958), .ZN(n14850) );
  XOR2_X1 U14901 ( .A(n14851), .B(n14852), .Z(n14849) );
  XOR2_X1 U14902 ( .A(n14853), .B(n14854), .Z(n14625) );
  NOR2_X1 U14903 ( .A1(n14599), .A2(n8353), .ZN(n14854) );
  XOR2_X1 U14904 ( .A(n14855), .B(n14856), .Z(n14853) );
  XOR2_X1 U14905 ( .A(n14857), .B(n14858), .Z(n14629) );
  NOR2_X1 U14906 ( .A1(n14599), .A2(n7962), .ZN(n14858) );
  XOR2_X1 U14907 ( .A(n14859), .B(n14860), .Z(n14857) );
  XOR2_X1 U14908 ( .A(n14861), .B(n14862), .Z(n14633) );
  NOR2_X1 U14909 ( .A1(n14599), .A2(n8585), .ZN(n14862) );
  XOR2_X1 U14910 ( .A(n14863), .B(n14864), .Z(n14861) );
  XOR2_X1 U14911 ( .A(n14865), .B(n14866), .Z(n14637) );
  NOR2_X1 U14912 ( .A1(n14599), .A2(n8378), .ZN(n14866) );
  XOR2_X1 U14913 ( .A(n14867), .B(n14868), .Z(n14865) );
  XOR2_X1 U14914 ( .A(n14869), .B(n14870), .Z(n14641) );
  NOR2_X1 U14915 ( .A1(n14599), .A2(n8602), .ZN(n14870) );
  XOR2_X1 U14916 ( .A(n14871), .B(n14872), .Z(n14869) );
  XOR2_X1 U14917 ( .A(n14873), .B(n14874), .Z(n14645) );
  NOR2_X1 U14918 ( .A1(n14599), .A2(n7807), .ZN(n14874) );
  XOR2_X1 U14919 ( .A(n14875), .B(n14876), .Z(n14873) );
  XOR2_X1 U14920 ( .A(n14877), .B(n14878), .Z(n14649) );
  NOR2_X1 U14921 ( .A1(n14599), .A2(n7836), .ZN(n14878) );
  XOR2_X1 U14922 ( .A(n14879), .B(n14880), .Z(n14877) );
  INV_X1 U14923 ( .A(n7859), .ZN(n14676) );
  NAND2_X1 U14924 ( .A1(a_2_), .A2(b_2_), .ZN(n7859) );
  XOR2_X1 U14925 ( .A(n14881), .B(n14882), .Z(n14656) );
  NOR2_X1 U14926 ( .A1(n14599), .A2(n7966), .ZN(n14882) );
  XOR2_X1 U14927 ( .A(n14883), .B(n14884), .Z(n14881) );
  XOR2_X1 U14928 ( .A(n14885), .B(n14886), .Z(n8094) );
  NOR2_X1 U14929 ( .A1(n14788), .A2(n7872), .ZN(n14886) );
  XOR2_X1 U14930 ( .A(n14887), .B(n14888), .Z(n14885) );
  NOR2_X1 U14931 ( .A1(n14788), .A2(n8197), .ZN(n7888) );
  NOR2_X1 U14932 ( .A1(n8096), .A2(n8197), .ZN(n8089) );
  AND2_X1 U14933 ( .A1(n14889), .A2(n14890), .ZN(n8096) );
  NAND3_X1 U14934 ( .A1(b_0_), .A2(n14891), .A3(a_1_), .ZN(n14890) );
  OR2_X1 U14935 ( .A1(n14888), .A2(n14887), .ZN(n14891) );
  NAND2_X1 U14936 ( .A1(n14887), .A2(n14888), .ZN(n14889) );
  NAND2_X1 U14937 ( .A1(n14892), .A2(n14893), .ZN(n14888) );
  NAND2_X1 U14938 ( .A1(n14667), .A2(n14894), .ZN(n14893) );
  OR2_X1 U14939 ( .A1(n14669), .A2(n7878), .ZN(n14894) );
  NOR2_X1 U14940 ( .A1(n7966), .A2(n14788), .ZN(n14667) );
  INV_X1 U14941 ( .A(a_2_), .ZN(n7966) );
  NAND2_X1 U14942 ( .A1(n7878), .A2(n14669), .ZN(n14892) );
  NAND2_X1 U14943 ( .A1(n14895), .A2(n14896), .ZN(n14669) );
  NAND3_X1 U14944 ( .A1(b_1_), .A2(n14897), .A3(a_2_), .ZN(n14896) );
  OR2_X1 U14945 ( .A1(n14884), .A2(n14883), .ZN(n14897) );
  NAND2_X1 U14946 ( .A1(n14883), .A2(n14884), .ZN(n14895) );
  NAND2_X1 U14947 ( .A1(n14898), .A2(n14899), .ZN(n14884) );
  NAND3_X1 U14948 ( .A1(b_1_), .A2(n14900), .A3(a_3_), .ZN(n14899) );
  OR2_X1 U14949 ( .A1(n14680), .A2(n14679), .ZN(n14900) );
  NAND2_X1 U14950 ( .A1(n14679), .A2(n14680), .ZN(n14898) );
  NAND2_X1 U14951 ( .A1(n14901), .A2(n14902), .ZN(n14680) );
  NAND3_X1 U14952 ( .A1(b_1_), .A2(n14903), .A3(a_4_), .ZN(n14902) );
  OR2_X1 U14953 ( .A1(n14880), .A2(n14879), .ZN(n14903) );
  NAND2_X1 U14954 ( .A1(n14879), .A2(n14880), .ZN(n14901) );
  NAND2_X1 U14955 ( .A1(n14904), .A2(n14905), .ZN(n14880) );
  NAND3_X1 U14956 ( .A1(b_1_), .A2(n14906), .A3(a_5_), .ZN(n14905) );
  OR2_X1 U14957 ( .A1(n14691), .A2(n14690), .ZN(n14906) );
  NAND2_X1 U14958 ( .A1(n14690), .A2(n14691), .ZN(n14904) );
  NAND2_X1 U14959 ( .A1(n14907), .A2(n14908), .ZN(n14691) );
  NAND3_X1 U14960 ( .A1(b_1_), .A2(n14909), .A3(a_6_), .ZN(n14908) );
  OR2_X1 U14961 ( .A1(n14876), .A2(n14875), .ZN(n14909) );
  NAND2_X1 U14962 ( .A1(n14875), .A2(n14876), .ZN(n14907) );
  NAND2_X1 U14963 ( .A1(n14910), .A2(n14911), .ZN(n14876) );
  NAND3_X1 U14964 ( .A1(b_1_), .A2(n14912), .A3(a_7_), .ZN(n14911) );
  OR2_X1 U14965 ( .A1(n14702), .A2(n14701), .ZN(n14912) );
  NAND2_X1 U14966 ( .A1(n14701), .A2(n14702), .ZN(n14910) );
  NAND2_X1 U14967 ( .A1(n14913), .A2(n14914), .ZN(n14702) );
  NAND3_X1 U14968 ( .A1(b_1_), .A2(n14915), .A3(a_8_), .ZN(n14914) );
  OR2_X1 U14969 ( .A1(n14872), .A2(n14871), .ZN(n14915) );
  NAND2_X1 U14970 ( .A1(n14871), .A2(n14872), .ZN(n14913) );
  NAND2_X1 U14971 ( .A1(n14916), .A2(n14917), .ZN(n14872) );
  NAND3_X1 U14972 ( .A1(b_1_), .A2(n14918), .A3(a_9_), .ZN(n14917) );
  OR2_X1 U14973 ( .A1(n14713), .A2(n14712), .ZN(n14918) );
  NAND2_X1 U14974 ( .A1(n14712), .A2(n14713), .ZN(n14916) );
  NAND2_X1 U14975 ( .A1(n14919), .A2(n14920), .ZN(n14713) );
  NAND3_X1 U14976 ( .A1(b_1_), .A2(n14921), .A3(a_10_), .ZN(n14920) );
  OR2_X1 U14977 ( .A1(n14868), .A2(n14867), .ZN(n14921) );
  NAND2_X1 U14978 ( .A1(n14867), .A2(n14868), .ZN(n14919) );
  NAND2_X1 U14979 ( .A1(n14922), .A2(n14923), .ZN(n14868) );
  NAND3_X1 U14980 ( .A1(a_11_), .A2(n14924), .A3(b_1_), .ZN(n14923) );
  OR2_X1 U14981 ( .A1(n14724), .A2(n14723), .ZN(n14924) );
  NAND2_X1 U14982 ( .A1(n14723), .A2(n14724), .ZN(n14922) );
  NAND2_X1 U14983 ( .A1(n14925), .A2(n14926), .ZN(n14724) );
  NAND3_X1 U14984 ( .A1(b_1_), .A2(n14927), .A3(a_12_), .ZN(n14926) );
  OR2_X1 U14985 ( .A1(n14864), .A2(n14863), .ZN(n14927) );
  NAND2_X1 U14986 ( .A1(n14863), .A2(n14864), .ZN(n14925) );
  NAND2_X1 U14987 ( .A1(n14928), .A2(n14929), .ZN(n14864) );
  NAND3_X1 U14988 ( .A1(b_1_), .A2(n14930), .A3(a_13_), .ZN(n14929) );
  OR2_X1 U14989 ( .A1(n14735), .A2(n14734), .ZN(n14930) );
  NAND2_X1 U14990 ( .A1(n14734), .A2(n14735), .ZN(n14928) );
  NAND2_X1 U14991 ( .A1(n14931), .A2(n14932), .ZN(n14735) );
  NAND3_X1 U14992 ( .A1(b_1_), .A2(n14933), .A3(a_14_), .ZN(n14932) );
  OR2_X1 U14993 ( .A1(n14860), .A2(n14859), .ZN(n14933) );
  NAND2_X1 U14994 ( .A1(n14859), .A2(n14860), .ZN(n14931) );
  NAND2_X1 U14995 ( .A1(n14934), .A2(n14935), .ZN(n14860) );
  NAND3_X1 U14996 ( .A1(b_1_), .A2(n14936), .A3(a_15_), .ZN(n14935) );
  OR2_X1 U14997 ( .A1(n14746), .A2(n14745), .ZN(n14936) );
  NAND2_X1 U14998 ( .A1(n14745), .A2(n14746), .ZN(n14934) );
  NAND2_X1 U14999 ( .A1(n14937), .A2(n14938), .ZN(n14746) );
  NAND3_X1 U15000 ( .A1(b_1_), .A2(n14939), .A3(a_16_), .ZN(n14938) );
  OR2_X1 U15001 ( .A1(n14856), .A2(n14855), .ZN(n14939) );
  NAND2_X1 U15002 ( .A1(n14855), .A2(n14856), .ZN(n14937) );
  NAND2_X1 U15003 ( .A1(n14940), .A2(n14941), .ZN(n14856) );
  NAND3_X1 U15004 ( .A1(b_1_), .A2(n14942), .A3(a_17_), .ZN(n14941) );
  OR2_X1 U15005 ( .A1(n14757), .A2(n14756), .ZN(n14942) );
  NAND2_X1 U15006 ( .A1(n14756), .A2(n14757), .ZN(n14940) );
  NAND2_X1 U15007 ( .A1(n14943), .A2(n14944), .ZN(n14757) );
  NAND3_X1 U15008 ( .A1(b_0_), .A2(n14945), .A3(a_19_), .ZN(n14944) );
  OR2_X1 U15009 ( .A1(n14852), .A2(n14851), .ZN(n14945) );
  NAND2_X1 U15010 ( .A1(n14851), .A2(n14852), .ZN(n14943) );
  NAND2_X1 U15011 ( .A1(n14946), .A2(n14947), .ZN(n14852) );
  NAND3_X1 U15012 ( .A1(b_0_), .A2(n14948), .A3(a_20_), .ZN(n14947) );
  OR2_X1 U15013 ( .A1(n14848), .A2(n14847), .ZN(n14948) );
  NAND2_X1 U15014 ( .A1(n14847), .A2(n14848), .ZN(n14946) );
  NAND2_X1 U15015 ( .A1(n14949), .A2(n14950), .ZN(n14848) );
  NAND3_X1 U15016 ( .A1(a_21_), .A2(n14951), .A3(b_0_), .ZN(n14950) );
  NAND2_X1 U15017 ( .A1(n14844), .A2(n14843), .ZN(n14951) );
  INV_X1 U15018 ( .A(n14952), .ZN(n14844) );
  NAND2_X1 U15019 ( .A1(n14953), .A2(n14952), .ZN(n14949) );
  NAND2_X1 U15020 ( .A1(n14954), .A2(n14955), .ZN(n14952) );
  NAND3_X1 U15021 ( .A1(a_22_), .A2(n14956), .A3(b_0_), .ZN(n14955) );
  OR2_X1 U15022 ( .A1(n14840), .A2(n14839), .ZN(n14956) );
  NAND2_X1 U15023 ( .A1(n14839), .A2(n14840), .ZN(n14954) );
  NAND2_X1 U15024 ( .A1(n14957), .A2(n14958), .ZN(n14840) );
  NAND3_X1 U15025 ( .A1(a_23_), .A2(n14959), .A3(b_0_), .ZN(n14958) );
  NAND2_X1 U15026 ( .A1(n14836), .A2(n14835), .ZN(n14959) );
  INV_X1 U15027 ( .A(n14960), .ZN(n14836) );
  NAND2_X1 U15028 ( .A1(n14961), .A2(n14960), .ZN(n14957) );
  NAND2_X1 U15029 ( .A1(n14962), .A2(n14963), .ZN(n14960) );
  NAND3_X1 U15030 ( .A1(a_24_), .A2(n14964), .A3(b_0_), .ZN(n14963) );
  OR2_X1 U15031 ( .A1(n14832), .A2(n14831), .ZN(n14964) );
  NAND2_X1 U15032 ( .A1(n14831), .A2(n14832), .ZN(n14962) );
  NAND2_X1 U15033 ( .A1(n14965), .A2(n14966), .ZN(n14832) );
  NAND3_X1 U15034 ( .A1(a_25_), .A2(n14967), .A3(b_0_), .ZN(n14966) );
  NAND2_X1 U15035 ( .A1(n14828), .A2(n14827), .ZN(n14967) );
  INV_X1 U15036 ( .A(n14968), .ZN(n14828) );
  NAND2_X1 U15037 ( .A1(n14969), .A2(n14968), .ZN(n14965) );
  NAND2_X1 U15038 ( .A1(n14970), .A2(n14971), .ZN(n14968) );
  NAND3_X1 U15039 ( .A1(a_26_), .A2(n14972), .A3(b_0_), .ZN(n14971) );
  OR2_X1 U15040 ( .A1(n14824), .A2(n14823), .ZN(n14972) );
  NAND2_X1 U15041 ( .A1(n14823), .A2(n14824), .ZN(n14970) );
  NAND2_X1 U15042 ( .A1(n14973), .A2(n14974), .ZN(n14824) );
  NAND3_X1 U15043 ( .A1(a_27_), .A2(n14975), .A3(b_0_), .ZN(n14974) );
  NAND2_X1 U15044 ( .A1(n14790), .A2(n14789), .ZN(n14975) );
  INV_X1 U15045 ( .A(n14976), .ZN(n14790) );
  NAND2_X1 U15046 ( .A1(n14977), .A2(n14976), .ZN(n14973) );
  NAND2_X1 U15047 ( .A1(n14978), .A2(n14979), .ZN(n14976) );
  NAND3_X1 U15048 ( .A1(a_28_), .A2(n14980), .A3(b_0_), .ZN(n14979) );
  OR2_X1 U15049 ( .A1(n14820), .A2(n14819), .ZN(n14980) );
  NAND2_X1 U15050 ( .A1(n14819), .A2(n14820), .ZN(n14978) );
  NAND2_X1 U15051 ( .A1(n14981), .A2(n14982), .ZN(n14820) );
  NAND3_X1 U15052 ( .A1(a_29_), .A2(n14983), .A3(b_0_), .ZN(n14982) );
  OR2_X1 U15053 ( .A1(n14816), .A2(n14815), .ZN(n14983) );
  NAND2_X1 U15054 ( .A1(n14815), .A2(n14816), .ZN(n14981) );
  NAND2_X1 U15055 ( .A1(n14812), .A2(n14984), .ZN(n14816) );
  NAND3_X1 U15056 ( .A1(b_0_), .A2(a_30_), .A3(n14811), .ZN(n14984) );
  NOR2_X1 U15057 ( .A1(n14599), .A2(n7460), .ZN(n14811) );
  NAND3_X1 U15058 ( .A1(b_1_), .A2(n7409), .A3(b_0_), .ZN(n14812) );
  INV_X1 U15059 ( .A(a_30_), .ZN(n7450) );
  INV_X1 U15060 ( .A(a_31_), .ZN(n7948) );
  NOR2_X1 U15061 ( .A1(n14599), .A2(n7480), .ZN(n14815) );
  INV_X1 U15062 ( .A(a_28_), .ZN(n7480) );
  NOR2_X1 U15063 ( .A1(n14599), .A2(n7950), .ZN(n14819) );
  INV_X1 U15064 ( .A(a_27_), .ZN(n7950) );
  INV_X1 U15065 ( .A(n14789), .ZN(n14977) );
  NAND2_X1 U15066 ( .A1(b_1_), .A2(a_26_), .ZN(n14789) );
  NOR2_X1 U15067 ( .A1(n14599), .A2(n7952), .ZN(n14823) );
  INV_X1 U15068 ( .A(n14827), .ZN(n14969) );
  NAND2_X1 U15069 ( .A1(b_1_), .A2(a_24_), .ZN(n14827) );
  NOR2_X1 U15070 ( .A1(n14599), .A2(n7955), .ZN(n14831) );
  INV_X1 U15071 ( .A(n14835), .ZN(n14961) );
  NAND2_X1 U15072 ( .A1(b_1_), .A2(a_22_), .ZN(n14835) );
  NOR2_X1 U15073 ( .A1(n14599), .A2(n7578), .ZN(n14839) );
  INV_X1 U15074 ( .A(n14843), .ZN(n14953) );
  NAND2_X1 U15075 ( .A1(a_20_), .A2(b_1_), .ZN(n14843) );
  NOR2_X1 U15076 ( .A1(n7958), .A2(n14599), .ZN(n14847) );
  INV_X1 U15077 ( .A(a_19_), .ZN(n7958) );
  NOR2_X1 U15078 ( .A1(n7960), .A2(n14599), .ZN(n14851) );
  NOR2_X1 U15079 ( .A1(n7960), .A2(n14788), .ZN(n14756) );
  NOR2_X1 U15080 ( .A1(n7645), .A2(n14788), .ZN(n14855) );
  NOR2_X1 U15081 ( .A1(n8353), .A2(n14788), .ZN(n14745) );
  INV_X1 U15082 ( .A(a_16_), .ZN(n8353) );
  NOR2_X1 U15083 ( .A1(n7667), .A2(n14788), .ZN(n14859) );
  INV_X1 U15084 ( .A(a_15_), .ZN(n7667) );
  NOR2_X1 U15085 ( .A1(n7962), .A2(n14788), .ZN(n14734) );
  INV_X1 U15086 ( .A(a_14_), .ZN(n7962) );
  NOR2_X1 U15087 ( .A1(n7702), .A2(n14788), .ZN(n14863) );
  INV_X1 U15088 ( .A(a_13_), .ZN(n7702) );
  NOR2_X1 U15089 ( .A1(n8585), .A2(n14788), .ZN(n14723) );
  INV_X1 U15090 ( .A(a_12_), .ZN(n8585) );
  NOR2_X1 U15091 ( .A1(n14788), .A2(n7724), .ZN(n14867) );
  INV_X1 U15092 ( .A(a_11_), .ZN(n7724) );
  NOR2_X1 U15093 ( .A1(n8378), .A2(n14788), .ZN(n14712) );
  INV_X1 U15094 ( .A(a_10_), .ZN(n8378) );
  NOR2_X1 U15095 ( .A1(n7753), .A2(n14788), .ZN(n14871) );
  INV_X1 U15096 ( .A(a_9_), .ZN(n7753) );
  NOR2_X1 U15097 ( .A1(n8602), .A2(n14788), .ZN(n14701) );
  INV_X1 U15098 ( .A(a_8_), .ZN(n8602) );
  NOR2_X1 U15099 ( .A1(n7787), .A2(n14788), .ZN(n14875) );
  INV_X1 U15100 ( .A(a_7_), .ZN(n7787) );
  NOR2_X1 U15101 ( .A1(n7807), .A2(n14788), .ZN(n14690) );
  INV_X1 U15102 ( .A(a_6_), .ZN(n7807) );
  NOR2_X1 U15103 ( .A1(n7823), .A2(n14788), .ZN(n14879) );
  INV_X1 U15104 ( .A(a_5_), .ZN(n7823) );
  NOR2_X1 U15105 ( .A1(n7836), .A2(n14788), .ZN(n14679) );
  INV_X1 U15106 ( .A(a_4_), .ZN(n7836) );
  NOR2_X1 U15107 ( .A1(n7852), .A2(n14788), .ZN(n14883) );
  INV_X1 U15108 ( .A(a_3_), .ZN(n7852) );
  NOR2_X1 U15109 ( .A1(n7872), .A2(n14599), .ZN(n7878) );
  NOR2_X1 U15110 ( .A1(n14599), .A2(n8197), .ZN(n14887) );
  INV_X1 U15111 ( .A(a_0_), .ZN(n8197) );
  INV_X1 U15112 ( .A(b_1_), .ZN(n14599) );
endmodule

