module add_mul_comp_4_bit ( a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_ );
  input a_0_, a_1_, a_2_, a_3_, b_0_, b_1_, b_2_, b_3_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_;
  wire   n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201;

  NAND2_X1 U110 ( .A1(n102), .A2(n103), .ZN(Result_7_) );
  NAND2_X1 U111 ( .A1(n104), .A2(n105), .ZN(n103) );
  NAND2_X1 U112 ( .A1(n106), .A2(n107), .ZN(n102) );
  NAND2_X1 U113 ( .A1(n108), .A2(n109), .ZN(n107) );
  NAND2_X1 U114 ( .A1(b_3_), .A2(n110), .ZN(n109) );
  NAND2_X1 U115 ( .A1(n111), .A2(n112), .ZN(Result_6_) );
  NAND2_X1 U116 ( .A1(n113), .A2(n105), .ZN(n112) );
  XNOR2_X1 U117 ( .A(n114), .B(n115), .ZN(n113) );
  NAND2_X1 U118 ( .A1(b_2_), .A2(a_3_), .ZN(n115) );
  NAND2_X1 U119 ( .A1(n116), .A2(n106), .ZN(n111) );
  XOR2_X1 U120 ( .A(n104), .B(n117), .Z(n116) );
  XOR2_X1 U121 ( .A(b_2_), .B(a_2_), .Z(n117) );
  NAND2_X1 U122 ( .A1(n118), .A2(n119), .ZN(Result_5_) );
  NAND2_X1 U123 ( .A1(n106), .A2(n120), .ZN(n119) );
  NAND3_X1 U124 ( .A1(n121), .A2(n122), .A3(n123), .ZN(n120) );
  OR2_X1 U125 ( .A1(n124), .A2(n125), .ZN(n123) );
  NAND3_X1 U126 ( .A1(n125), .A2(n126), .A3(b_1_), .ZN(n122) );
  NAND2_X1 U127 ( .A1(n127), .A2(n128), .ZN(n121) );
  XOR2_X1 U128 ( .A(n126), .B(n125), .Z(n127) );
  NAND2_X1 U129 ( .A1(n129), .A2(n105), .ZN(n118) );
  XNOR2_X1 U130 ( .A(n130), .B(n131), .ZN(n129) );
  XNOR2_X1 U131 ( .A(n132), .B(n133), .ZN(n131) );
  NAND2_X1 U132 ( .A1(n134), .A2(n135), .ZN(Result_4_) );
  NAND2_X1 U133 ( .A1(n136), .A2(n105), .ZN(n135) );
  XNOR2_X1 U134 ( .A(n137), .B(n138), .ZN(n136) );
  XOR2_X1 U135 ( .A(n139), .B(n140), .Z(n138) );
  NOR2_X1 U136 ( .A1(n141), .A2(n142), .ZN(n140) );
  NAND2_X1 U137 ( .A1(n143), .A2(n106), .ZN(n134) );
  XOR2_X1 U138 ( .A(n144), .B(n145), .Z(n143) );
  NAND2_X1 U139 ( .A1(n146), .A2(n147), .ZN(n145) );
  NAND2_X1 U140 ( .A1(n125), .A2(n124), .ZN(n147) );
  NOR2_X1 U141 ( .A1(n148), .A2(n149), .ZN(n125) );
  AND2_X1 U142 ( .A1(n104), .A2(n150), .ZN(n148) );
  NAND2_X1 U143 ( .A1(n151), .A2(n152), .ZN(n150) );
  NOR2_X1 U144 ( .A1(n142), .A2(n110), .ZN(n104) );
  NAND2_X1 U145 ( .A1(n126), .A2(n128), .ZN(n146) );
  NOR2_X1 U146 ( .A1(n106), .A2(n153), .ZN(Result_3_) );
  XNOR2_X1 U147 ( .A(n154), .B(n155), .ZN(n153) );
  NOR2_X1 U148 ( .A1(n106), .A2(n156), .ZN(Result_2_) );
  XNOR2_X1 U149 ( .A(n157), .B(n158), .ZN(n156) );
  NOR2_X1 U150 ( .A1(n106), .A2(n159), .ZN(Result_1_) );
  XNOR2_X1 U151 ( .A(n160), .B(n161), .ZN(n159) );
  NOR2_X1 U152 ( .A1(n106), .A2(n162), .ZN(Result_0_) );
  NOR3_X1 U153 ( .A1(n163), .A2(n164), .A3(n165), .ZN(n162) );
  NOR3_X1 U154 ( .A1(n166), .A2(n167), .A3(n168), .ZN(n165) );
  NOR2_X1 U155 ( .A1(n160), .A2(n161), .ZN(n163) );
  NAND2_X1 U156 ( .A1(n157), .A2(n158), .ZN(n161) );
  XOR2_X1 U157 ( .A(n168), .B(n167), .Z(n158) );
  AND2_X1 U158 ( .A1(n155), .A2(n154), .ZN(n157) );
  NAND2_X1 U159 ( .A1(n139), .A2(n169), .ZN(n154) );
  NAND3_X1 U160 ( .A1(a_0_), .A2(n137), .A3(b_3_), .ZN(n169) );
  XNOR2_X1 U161 ( .A(n170), .B(n171), .ZN(n137) );
  XOR2_X1 U162 ( .A(n172), .B(n173), .Z(n170) );
  AND2_X1 U163 ( .A1(n174), .A2(n175), .ZN(n139) );
  NAND2_X1 U164 ( .A1(n133), .A2(n176), .ZN(n175) );
  OR2_X1 U165 ( .A1(n130), .A2(n132), .ZN(n176) );
  AND3_X1 U166 ( .A1(b_2_), .A2(a_3_), .A3(n114), .ZN(n133) );
  NOR2_X1 U167 ( .A1(n142), .A2(n151), .ZN(n114) );
  NAND2_X1 U168 ( .A1(n132), .A2(n130), .ZN(n174) );
  XOR2_X1 U169 ( .A(n149), .B(n177), .Z(n130) );
  NOR2_X1 U170 ( .A1(n142), .A2(n126), .ZN(n132) );
  XNOR2_X1 U171 ( .A(n178), .B(n179), .ZN(n155) );
  XNOR2_X1 U172 ( .A(n180), .B(n181), .ZN(n179) );
  NAND2_X1 U173 ( .A1(a_0_), .A2(b_2_), .ZN(n181) );
  XOR2_X1 U174 ( .A(n182), .B(n183), .Z(n160) );
  NOR2_X1 U175 ( .A1(n167), .A2(n168), .ZN(n183) );
  XOR2_X1 U176 ( .A(n184), .B(n185), .Z(n168) );
  NOR2_X1 U177 ( .A1(n166), .A2(n126), .ZN(n185) );
  OR3_X1 U178 ( .A1(n128), .A2(n186), .A3(n141), .ZN(n184) );
  AND2_X1 U179 ( .A1(n180), .A2(n187), .ZN(n167) );
  NAND2_X1 U180 ( .A1(b_2_), .A2(n178), .ZN(n187) );
  NAND2_X1 U181 ( .A1(n188), .A2(n189), .ZN(n178) );
  NAND2_X1 U182 ( .A1(n190), .A2(a_2_), .ZN(n189) );
  XOR2_X1 U183 ( .A(n124), .B(n186), .Z(n188) );
  NOR2_X1 U184 ( .A1(n151), .A2(n166), .ZN(n186) );
  AND2_X1 U185 ( .A1(n191), .A2(n173), .ZN(n180) );
  NAND2_X1 U186 ( .A1(n177), .A2(n149), .ZN(n173) );
  NOR2_X1 U187 ( .A1(n152), .A2(n151), .ZN(n149) );
  NOR2_X1 U188 ( .A1(n128), .A2(n110), .ZN(n177) );
  NAND2_X1 U189 ( .A1(n172), .A2(n171), .ZN(n191) );
  XOR2_X1 U190 ( .A(n190), .B(n192), .Z(n171) );
  NOR2_X1 U191 ( .A1(n151), .A2(n128), .ZN(n192) );
  NOR2_X1 U192 ( .A1(n110), .A2(n166), .ZN(n190) );
  INV_X1 U193 ( .A(a_3_), .ZN(n110) );
  NOR2_X1 U194 ( .A1(n152), .A2(n126), .ZN(n172) );
  INV_X1 U195 ( .A(b_2_), .ZN(n152) );
  OR2_X1 U196 ( .A1(n166), .A2(n164), .ZN(n182) );
  NOR2_X1 U197 ( .A1(n124), .A2(n166), .ZN(n164) );
  NAND2_X1 U198 ( .A1(b_1_), .A2(a_1_), .ZN(n124) );
  INV_X1 U199 ( .A(n105), .ZN(n106) );
  NAND2_X1 U200 ( .A1(n193), .A2(n194), .ZN(n105) );
  NAND2_X1 U201 ( .A1(n195), .A2(n144), .ZN(n194) );
  NAND2_X1 U202 ( .A1(b_0_), .A2(n141), .ZN(n144) );
  INV_X1 U203 ( .A(a_0_), .ZN(n141) );
  NAND2_X1 U204 ( .A1(n196), .A2(n197), .ZN(n195) );
  NAND2_X1 U205 ( .A1(a_1_), .A2(n128), .ZN(n197) );
  INV_X1 U206 ( .A(b_1_), .ZN(n128) );
  NAND3_X1 U207 ( .A1(n198), .A2(n199), .A3(n200), .ZN(n196) );
  NAND2_X1 U208 ( .A1(b_1_), .A2(n126), .ZN(n200) );
  INV_X1 U209 ( .A(a_1_), .ZN(n126) );
  NAND2_X1 U210 ( .A1(b_2_), .A2(n201), .ZN(n199) );
  OR2_X1 U211 ( .A1(n151), .A2(n108), .ZN(n201) );
  NAND2_X1 U212 ( .A1(n108), .A2(n151), .ZN(n198) );
  INV_X1 U213 ( .A(a_2_), .ZN(n151) );
  NAND2_X1 U214 ( .A1(a_3_), .A2(n142), .ZN(n108) );
  INV_X1 U215 ( .A(b_3_), .ZN(n142) );
  NAND2_X1 U216 ( .A1(a_0_), .A2(n166), .ZN(n193) );
  INV_X1 U217 ( .A(b_0_), .ZN(n166) );
endmodule

