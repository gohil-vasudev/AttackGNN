module add_mul_32_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, 
        a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, 
        a_19_, a_20_, a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, 
        a_29_, a_30_, a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, 
        b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, 
        b_18_, b_19_, b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, 
        b_28_, b_29_, b_30_, b_31_, operation, Result_0_, Result_1_, Result_2_, 
        Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, Result_8_, 
        Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, Result_14_, 
        Result_15_, Result_16_, Result_17_, Result_18_, Result_19_, Result_20_, 
        Result_21_, Result_22_, Result_23_, Result_24_, Result_25_, Result_26_, 
        Result_27_, Result_28_, Result_29_, Result_30_, Result_31_, Result_32_, 
        Result_33_, Result_34_, Result_35_, Result_36_, Result_37_, Result_38_, 
        Result_39_, Result_40_, Result_41_, Result_42_, Result_43_, Result_44_, 
        Result_45_, Result_46_, Result_47_, Result_48_, Result_49_, Result_50_, 
        Result_51_, Result_52_, Result_53_, Result_54_, Result_55_, Result_56_, 
        Result_57_, Result_58_, Result_59_, Result_60_, Result_61_, Result_62_, 
        Result_63_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, a_16_, a_17_, a_18_, a_19_, a_20_,
         a_21_, a_22_, a_23_, a_24_, a_25_, a_26_, a_27_, a_28_, a_29_, a_30_,
         a_31_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_,
         b_10_, b_11_, b_12_, b_13_, b_14_, b_15_, b_16_, b_17_, b_18_, b_19_,
         b_20_, b_21_, b_22_, b_23_, b_24_, b_25_, b_26_, b_27_, b_28_, b_29_,
         b_30_, b_31_, operation;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_,
         Result_32_, Result_33_, Result_34_, Result_35_, Result_36_,
         Result_37_, Result_38_, Result_39_, Result_40_, Result_41_,
         Result_42_, Result_43_, Result_44_, Result_45_, Result_46_,
         Result_47_, Result_48_, Result_49_, Result_50_, Result_51_,
         Result_52_, Result_53_, Result_54_, Result_55_, Result_56_,
         Result_57_, Result_58_, Result_59_, Result_60_, Result_61_,
         Result_62_, Result_63_;
  wire   n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653;

  INV_X2 U7539 ( .A(b_23_), .ZN(n7625) );
  INV_X2 U7540 ( .A(b_28_), .ZN(n8050) );
  INV_X2 U7541 ( .A(b_29_), .ZN(n7527) );
  NAND2_X2 U7542 ( .A1(a_31_), .A2(a_30_), .ZN(n8451) );
  INV_X2 U7543 ( .A(b_21_), .ZN(n7657) );
  INV_X2 U7544 ( .A(b_3_), .ZN(n7946) );
  INV_X2 U7545 ( .A(b_27_), .ZN(n7564) );
  INV_X2 U7546 ( .A(b_25_), .ZN(n7594) );
  INV_X4 U7547 ( .A(b_11_), .ZN(n7818) );
  INV_X4 U7548 ( .A(a_29_), .ZN(n7529) );
  INV_X4 U7549 ( .A(operation), .ZN(n7475) );
  INV_X2 U7550 ( .A(a_31_), .ZN(n8048) );
  INV_X2 U7551 ( .A(b_8_), .ZN(n8058) );
  INV_X2 U7552 ( .A(b_19_), .ZN(n7688) );
  INV_X2 U7553 ( .A(b_30_), .ZN(n7512) );
  INV_X2 U7554 ( .A(a_6_), .ZN(n8061) );
  INV_X2 U7555 ( .A(n7506), .ZN(n8676) );
  INV_X2 U7556 ( .A(n7510), .ZN(n8679) );
  INV_X2 U7557 ( .A(a_13_), .ZN(n7786) );
  INV_X2 U7558 ( .A(b_10_), .ZN(n13001) );
  INV_X2 U7559 ( .A(a_30_), .ZN(n7515) );
  INV_X2 U7560 ( .A(a_17_), .ZN(n7723) );
  INV_X2 U7561 ( .A(a_19_), .ZN(n7687) );
  INV_X2 U7562 ( .A(b_0_), .ZN(n15294) );
  INV_X2 U7563 ( .A(b_4_), .ZN(n8062) );
  INV_X2 U7564 ( .A(a_8_), .ZN(n8059) );
  INV_X2 U7565 ( .A(a_27_), .ZN(n7563) );
  INV_X2 U7566 ( .A(a_23_), .ZN(n7624) );
  INV_X2 U7567 ( .A(a_25_), .ZN(n7593) );
  INV_X2 U7568 ( .A(a_15_), .ZN(n7754) );
  INV_X2 U7569 ( .A(a_7_), .ZN(n7884) );
  INV_X2 U7570 ( .A(a_10_), .ZN(n7837) );
  INV_X2 U7571 ( .A(a_9_), .ZN(n7848) );
  INV_X2 U7572 ( .A(a_3_), .ZN(n7945) );
  INV_X2 U7573 ( .A(a_16_), .ZN(n7743) );
  INV_X2 U7574 ( .A(a_21_), .ZN(n7656) );
  INV_X2 U7575 ( .A(a_0_), .ZN(n8307) );
  INV_X2 U7576 ( .A(a_1_), .ZN(n7973) );
  INV_X2 U7577 ( .A(a_14_), .ZN(n7775) );
  INV_X2 U7578 ( .A(a_12_), .ZN(n7806) );
  INV_X2 U7579 ( .A(a_4_), .ZN(n7934) );
  INV_X2 U7580 ( .A(b_6_), .ZN(n8060) );
  INV_X2 U7581 ( .A(a_5_), .ZN(n7914) );
  INV_X2 U7582 ( .A(b_9_), .ZN(n7849) );
  INV_X2 U7583 ( .A(a_18_), .ZN(n7707) );
  INV_X2 U7584 ( .A(b_1_), .ZN(n15217) );
  INV_X2 U7585 ( .A(a_11_), .ZN(n7817) );
  INV_X2 U7586 ( .A(b_7_), .ZN(n7885) );
  INV_X2 U7587 ( .A(a_20_), .ZN(n7676) );
  INV_X2 U7588 ( .A(b_5_), .ZN(n7915) );
  INV_X2 U7589 ( .A(a_22_), .ZN(n7645) );
  NOR2_X1 U7590 ( .A1(n7475), .A2(n7476), .ZN(Result_9_) );
  XOR2_X1 U7591 ( .A(n7477), .B(n7478), .Z(n7476) );
  NAND2_X1 U7592 ( .A1(n7479), .A2(n7480), .ZN(n7478) );
  NOR2_X1 U7593 ( .A1(n7475), .A2(n7481), .ZN(Result_8_) );
  XOR2_X1 U7594 ( .A(n7482), .B(n7483), .Z(n7481) );
  NAND2_X1 U7595 ( .A1(n7484), .A2(n7485), .ZN(n7483) );
  NOR2_X1 U7596 ( .A1(n7475), .A2(n7486), .ZN(Result_7_) );
  XOR2_X1 U7597 ( .A(n7487), .B(n7488), .Z(n7486) );
  NAND2_X1 U7598 ( .A1(n7489), .A2(n7490), .ZN(n7488) );
  NOR2_X1 U7599 ( .A1(n7475), .A2(n7491), .ZN(Result_6_) );
  XOR2_X1 U7600 ( .A(n7492), .B(n7493), .Z(n7491) );
  NAND2_X1 U7601 ( .A1(n7494), .A2(n7495), .ZN(n7493) );
  NAND2_X1 U7602 ( .A1(n7496), .A2(n7497), .ZN(Result_63_) );
  NAND2_X1 U7603 ( .A1(n7498), .A2(n7475), .ZN(n7497) );
  XOR2_X1 U7604 ( .A(b_31_), .B(a_31_), .Z(n7498) );
  NAND2_X1 U7605 ( .A1(n7499), .A2(operation), .ZN(n7496) );
  NAND2_X1 U7606 ( .A1(n7500), .A2(n7501), .ZN(Result_62_) );
  NAND2_X1 U7607 ( .A1(operation), .A2(n7502), .ZN(n7501) );
  NAND2_X1 U7608 ( .A1(n7503), .A2(n7504), .ZN(n7502) );
  NAND2_X1 U7609 ( .A1(b_30_), .A2(n7505), .ZN(n7504) );
  NAND2_X1 U7610 ( .A1(n7506), .A2(n7507), .ZN(n7505) );
  NAND2_X1 U7611 ( .A1(a_31_), .A2(n7508), .ZN(n7507) );
  NAND2_X1 U7612 ( .A1(b_31_), .A2(n7509), .ZN(n7503) );
  NAND2_X1 U7613 ( .A1(n7510), .A2(n7511), .ZN(n7509) );
  NAND2_X1 U7614 ( .A1(a_30_), .A2(n7512), .ZN(n7511) );
  NAND2_X1 U7615 ( .A1(n7513), .A2(n7475), .ZN(n7500) );
  XNOR2_X1 U7616 ( .A(n7499), .B(n7514), .ZN(n7513) );
  XOR2_X1 U7617 ( .A(n7515), .B(b_30_), .Z(n7514) );
  NAND2_X1 U7618 ( .A1(n7516), .A2(n7517), .ZN(Result_61_) );
  NAND2_X1 U7619 ( .A1(n7518), .A2(n7475), .ZN(n7517) );
  NAND2_X1 U7620 ( .A1(n7519), .A2(n7520), .ZN(n7518) );
  NAND2_X1 U7621 ( .A1(n7521), .A2(n7522), .ZN(n7520) );
  NOR2_X1 U7622 ( .A1(n7523), .A2(n7524), .ZN(n7519) );
  NOR2_X1 U7623 ( .A1(b_29_), .A2(n7525), .ZN(n7524) );
  XOR2_X1 U7624 ( .A(a_29_), .B(n7526), .Z(n7525) );
  NOR2_X1 U7625 ( .A1(n7527), .A2(n7528), .ZN(n7523) );
  NAND2_X1 U7626 ( .A1(n7526), .A2(n7529), .ZN(n7528) );
  INV_X1 U7627 ( .A(n7522), .ZN(n7526) );
  NAND2_X1 U7628 ( .A1(n7530), .A2(operation), .ZN(n7516) );
  XOR2_X1 U7629 ( .A(n7531), .B(n7532), .Z(n7530) );
  XNOR2_X1 U7630 ( .A(n7533), .B(n7534), .ZN(n7532) );
  NAND2_X1 U7631 ( .A1(b_31_), .A2(a_29_), .ZN(n7531) );
  NAND2_X1 U7632 ( .A1(n7535), .A2(n7536), .ZN(Result_60_) );
  NAND2_X1 U7633 ( .A1(n7537), .A2(n7475), .ZN(n7536) );
  XNOR2_X1 U7634 ( .A(n7538), .B(n7539), .ZN(n7537) );
  NAND2_X1 U7635 ( .A1(n7540), .A2(n7541), .ZN(n7538) );
  NAND2_X1 U7636 ( .A1(n7542), .A2(operation), .ZN(n7535) );
  XNOR2_X1 U7637 ( .A(n7543), .B(n7544), .ZN(n7542) );
  XNOR2_X1 U7638 ( .A(n7545), .B(n7546), .ZN(n7544) );
  NOR2_X1 U7639 ( .A1(n7547), .A2(n7508), .ZN(n7546) );
  NOR2_X1 U7640 ( .A1(n7475), .A2(n7548), .ZN(Result_5_) );
  XOR2_X1 U7641 ( .A(n7549), .B(n7550), .Z(n7548) );
  NAND2_X1 U7642 ( .A1(n7551), .A2(n7552), .ZN(n7550) );
  NAND2_X1 U7643 ( .A1(n7553), .A2(n7554), .ZN(Result_59_) );
  NAND2_X1 U7644 ( .A1(n7555), .A2(n7475), .ZN(n7554) );
  NAND2_X1 U7645 ( .A1(n7556), .A2(n7557), .ZN(n7555) );
  NAND2_X1 U7646 ( .A1(n7558), .A2(n7559), .ZN(n7557) );
  NOR2_X1 U7647 ( .A1(n7560), .A2(n7561), .ZN(n7556) );
  NOR2_X1 U7648 ( .A1(b_27_), .A2(n7562), .ZN(n7561) );
  XOR2_X1 U7649 ( .A(n7563), .B(n7559), .Z(n7562) );
  NOR2_X1 U7650 ( .A1(n7564), .A2(n7565), .ZN(n7560) );
  OR2_X1 U7651 ( .A1(n7559), .A2(a_27_), .ZN(n7565) );
  NAND2_X1 U7652 ( .A1(n7566), .A2(operation), .ZN(n7553) );
  XNOR2_X1 U7653 ( .A(n7567), .B(n7568), .ZN(n7566) );
  XNOR2_X1 U7654 ( .A(n7569), .B(n7570), .ZN(n7568) );
  NOR2_X1 U7655 ( .A1(n7563), .A2(n7508), .ZN(n7570) );
  NAND2_X1 U7656 ( .A1(n7571), .A2(n7572), .ZN(Result_58_) );
  NAND2_X1 U7657 ( .A1(n7573), .A2(n7475), .ZN(n7572) );
  XOR2_X1 U7658 ( .A(n7574), .B(n7575), .Z(n7573) );
  AND2_X1 U7659 ( .A1(n7576), .A2(n7577), .ZN(n7575) );
  NAND2_X1 U7660 ( .A1(n7578), .A2(operation), .ZN(n7571) );
  XNOR2_X1 U7661 ( .A(n7579), .B(n7580), .ZN(n7578) );
  NAND2_X1 U7662 ( .A1(n7581), .A2(n7582), .ZN(n7579) );
  NAND2_X1 U7663 ( .A1(n7583), .A2(n7584), .ZN(Result_57_) );
  NAND2_X1 U7664 ( .A1(n7585), .A2(n7475), .ZN(n7584) );
  NAND2_X1 U7665 ( .A1(n7586), .A2(n7587), .ZN(n7585) );
  NAND2_X1 U7666 ( .A1(n7588), .A2(n7589), .ZN(n7587) );
  NOR2_X1 U7667 ( .A1(n7590), .A2(n7591), .ZN(n7586) );
  NOR2_X1 U7668 ( .A1(b_25_), .A2(n7592), .ZN(n7591) );
  XOR2_X1 U7669 ( .A(n7593), .B(n7589), .Z(n7592) );
  NOR2_X1 U7670 ( .A1(n7594), .A2(n7595), .ZN(n7590) );
  OR2_X1 U7671 ( .A1(n7589), .A2(a_25_), .ZN(n7595) );
  NAND2_X1 U7672 ( .A1(n7596), .A2(operation), .ZN(n7583) );
  XNOR2_X1 U7673 ( .A(n7597), .B(n7598), .ZN(n7596) );
  NAND2_X1 U7674 ( .A1(n7599), .A2(n7600), .ZN(n7597) );
  NAND2_X1 U7675 ( .A1(n7601), .A2(n7602), .ZN(Result_56_) );
  NAND2_X1 U7676 ( .A1(n7603), .A2(n7475), .ZN(n7602) );
  XNOR2_X1 U7677 ( .A(n7604), .B(n7605), .ZN(n7603) );
  NOR2_X1 U7678 ( .A1(n7606), .A2(n7607), .ZN(n7605) );
  NAND2_X1 U7679 ( .A1(n7608), .A2(operation), .ZN(n7601) );
  XOR2_X1 U7680 ( .A(n7609), .B(n7610), .Z(n7608) );
  XOR2_X1 U7681 ( .A(n7611), .B(n7612), .Z(n7609) );
  NOR2_X1 U7682 ( .A1(n7613), .A2(n7508), .ZN(n7612) );
  NAND2_X1 U7683 ( .A1(n7614), .A2(n7615), .ZN(Result_55_) );
  NAND2_X1 U7684 ( .A1(n7616), .A2(n7475), .ZN(n7615) );
  NAND2_X1 U7685 ( .A1(n7617), .A2(n7618), .ZN(n7616) );
  NAND2_X1 U7686 ( .A1(n7619), .A2(n7620), .ZN(n7618) );
  NOR2_X1 U7687 ( .A1(n7621), .A2(n7622), .ZN(n7617) );
  NOR2_X1 U7688 ( .A1(b_23_), .A2(n7623), .ZN(n7622) );
  XOR2_X1 U7689 ( .A(n7624), .B(n7620), .Z(n7623) );
  NOR2_X1 U7690 ( .A1(n7625), .A2(n7626), .ZN(n7621) );
  NAND2_X1 U7691 ( .A1(n7627), .A2(n7624), .ZN(n7626) );
  NAND2_X1 U7692 ( .A1(n7628), .A2(operation), .ZN(n7614) );
  XNOR2_X1 U7693 ( .A(n7629), .B(n7630), .ZN(n7628) );
  NAND2_X1 U7694 ( .A1(n7631), .A2(n7632), .ZN(n7629) );
  NAND2_X1 U7695 ( .A1(n7633), .A2(n7634), .ZN(Result_54_) );
  NAND2_X1 U7696 ( .A1(n7635), .A2(n7475), .ZN(n7634) );
  XOR2_X1 U7697 ( .A(n7636), .B(n7637), .Z(n7635) );
  AND2_X1 U7698 ( .A1(n7638), .A2(n7639), .ZN(n7637) );
  NAND2_X1 U7699 ( .A1(n7640), .A2(operation), .ZN(n7633) );
  XOR2_X1 U7700 ( .A(n7641), .B(n7642), .Z(n7640) );
  XOR2_X1 U7701 ( .A(n7643), .B(n7644), .Z(n7641) );
  NOR2_X1 U7702 ( .A1(n7645), .A2(n7508), .ZN(n7644) );
  NAND2_X1 U7703 ( .A1(n7646), .A2(n7647), .ZN(Result_53_) );
  NAND2_X1 U7704 ( .A1(n7648), .A2(n7475), .ZN(n7647) );
  NAND2_X1 U7705 ( .A1(n7649), .A2(n7650), .ZN(n7648) );
  NAND2_X1 U7706 ( .A1(n7651), .A2(n7652), .ZN(n7650) );
  NOR2_X1 U7707 ( .A1(n7653), .A2(n7654), .ZN(n7649) );
  NOR2_X1 U7708 ( .A1(b_21_), .A2(n7655), .ZN(n7654) );
  XOR2_X1 U7709 ( .A(n7656), .B(n7652), .Z(n7655) );
  NOR2_X1 U7710 ( .A1(n7657), .A2(n7658), .ZN(n7653) );
  OR2_X1 U7711 ( .A1(n7652), .A2(a_21_), .ZN(n7658) );
  NAND2_X1 U7712 ( .A1(n7659), .A2(operation), .ZN(n7646) );
  XNOR2_X1 U7713 ( .A(n7660), .B(n7661), .ZN(n7659) );
  NAND2_X1 U7714 ( .A1(n7662), .A2(n7663), .ZN(n7660) );
  NAND2_X1 U7715 ( .A1(n7664), .A2(n7665), .ZN(Result_52_) );
  NAND2_X1 U7716 ( .A1(n7666), .A2(n7475), .ZN(n7665) );
  XOR2_X1 U7717 ( .A(n7667), .B(n7668), .Z(n7666) );
  AND2_X1 U7718 ( .A1(n7669), .A2(n7670), .ZN(n7668) );
  NAND2_X1 U7719 ( .A1(n7671), .A2(operation), .ZN(n7664) );
  XOR2_X1 U7720 ( .A(n7672), .B(n7673), .Z(n7671) );
  XOR2_X1 U7721 ( .A(n7674), .B(n7675), .Z(n7672) );
  NOR2_X1 U7722 ( .A1(n7676), .A2(n7508), .ZN(n7675) );
  NAND2_X1 U7723 ( .A1(n7677), .A2(n7678), .ZN(Result_51_) );
  NAND2_X1 U7724 ( .A1(n7679), .A2(n7475), .ZN(n7678) );
  NAND2_X1 U7725 ( .A1(n7680), .A2(n7681), .ZN(n7679) );
  NAND2_X1 U7726 ( .A1(n7682), .A2(n7683), .ZN(n7681) );
  NOR2_X1 U7727 ( .A1(n7684), .A2(n7685), .ZN(n7680) );
  NOR2_X1 U7728 ( .A1(b_19_), .A2(n7686), .ZN(n7685) );
  XOR2_X1 U7729 ( .A(n7687), .B(n7683), .Z(n7686) );
  NOR2_X1 U7730 ( .A1(n7688), .A2(n7689), .ZN(n7684) );
  OR2_X1 U7731 ( .A1(n7683), .A2(a_19_), .ZN(n7689) );
  NAND2_X1 U7732 ( .A1(n7690), .A2(operation), .ZN(n7677) );
  XNOR2_X1 U7733 ( .A(n7691), .B(n7692), .ZN(n7690) );
  XOR2_X1 U7734 ( .A(n7693), .B(n7694), .Z(n7692) );
  NAND2_X1 U7735 ( .A1(b_31_), .A2(a_19_), .ZN(n7694) );
  NAND2_X1 U7736 ( .A1(n7695), .A2(n7696), .ZN(Result_50_) );
  NAND2_X1 U7737 ( .A1(n7697), .A2(n7475), .ZN(n7696) );
  XOR2_X1 U7738 ( .A(n7698), .B(n7699), .Z(n7697) );
  AND2_X1 U7739 ( .A1(n7700), .A2(n7701), .ZN(n7699) );
  NAND2_X1 U7740 ( .A1(n7702), .A2(operation), .ZN(n7695) );
  XOR2_X1 U7741 ( .A(n7703), .B(n7704), .Z(n7702) );
  XOR2_X1 U7742 ( .A(n7705), .B(n7706), .Z(n7703) );
  NOR2_X1 U7743 ( .A1(n7707), .A2(n7508), .ZN(n7706) );
  NOR2_X1 U7744 ( .A1(n7475), .A2(n7708), .ZN(Result_4_) );
  XOR2_X1 U7745 ( .A(n7709), .B(n7710), .Z(n7708) );
  NAND2_X1 U7746 ( .A1(n7711), .A2(n7712), .ZN(n7710) );
  NAND2_X1 U7747 ( .A1(n7713), .A2(n7714), .ZN(Result_49_) );
  NAND2_X1 U7748 ( .A1(n7715), .A2(n7475), .ZN(n7714) );
  NAND2_X1 U7749 ( .A1(n7716), .A2(n7717), .ZN(n7715) );
  NAND2_X1 U7750 ( .A1(n7718), .A2(n7719), .ZN(n7717) );
  NOR2_X1 U7751 ( .A1(n7720), .A2(n7721), .ZN(n7716) );
  NOR2_X1 U7752 ( .A1(b_17_), .A2(n7722), .ZN(n7721) );
  XOR2_X1 U7753 ( .A(n7723), .B(n7719), .Z(n7722) );
  NOR2_X1 U7754 ( .A1(n7724), .A2(n7725), .ZN(n7720) );
  OR2_X1 U7755 ( .A1(n7719), .A2(a_17_), .ZN(n7725) );
  NAND2_X1 U7756 ( .A1(n7726), .A2(operation), .ZN(n7713) );
  XNOR2_X1 U7757 ( .A(n7727), .B(n7728), .ZN(n7726) );
  XOR2_X1 U7758 ( .A(n7729), .B(n7730), .Z(n7728) );
  NAND2_X1 U7759 ( .A1(b_31_), .A2(a_17_), .ZN(n7730) );
  NAND2_X1 U7760 ( .A1(n7731), .A2(n7732), .ZN(Result_48_) );
  NAND2_X1 U7761 ( .A1(n7733), .A2(n7475), .ZN(n7732) );
  XNOR2_X1 U7762 ( .A(n7734), .B(n7735), .ZN(n7733) );
  NOR2_X1 U7763 ( .A1(n7736), .A2(n7737), .ZN(n7735) );
  NAND2_X1 U7764 ( .A1(n7738), .A2(operation), .ZN(n7731) );
  XOR2_X1 U7765 ( .A(n7739), .B(n7740), .Z(n7738) );
  XOR2_X1 U7766 ( .A(n7741), .B(n7742), .Z(n7739) );
  NOR2_X1 U7767 ( .A1(n7743), .A2(n7508), .ZN(n7742) );
  NAND2_X1 U7768 ( .A1(n7744), .A2(n7745), .ZN(Result_47_) );
  NAND2_X1 U7769 ( .A1(n7746), .A2(n7475), .ZN(n7745) );
  NAND2_X1 U7770 ( .A1(n7747), .A2(n7748), .ZN(n7746) );
  NAND2_X1 U7771 ( .A1(n7749), .A2(n7750), .ZN(n7748) );
  NOR2_X1 U7772 ( .A1(n7751), .A2(n7752), .ZN(n7747) );
  NOR2_X1 U7773 ( .A1(b_15_), .A2(n7753), .ZN(n7752) );
  XOR2_X1 U7774 ( .A(n7754), .B(n7750), .Z(n7753) );
  NOR2_X1 U7775 ( .A1(n7755), .A2(n7756), .ZN(n7751) );
  NAND2_X1 U7776 ( .A1(n7757), .A2(n7754), .ZN(n7756) );
  NAND2_X1 U7777 ( .A1(n7758), .A2(operation), .ZN(n7744) );
  XNOR2_X1 U7778 ( .A(n7759), .B(n7760), .ZN(n7758) );
  XOR2_X1 U7779 ( .A(n7761), .B(n7762), .Z(n7760) );
  NAND2_X1 U7780 ( .A1(b_31_), .A2(a_15_), .ZN(n7762) );
  NAND2_X1 U7781 ( .A1(n7763), .A2(n7764), .ZN(Result_46_) );
  NAND2_X1 U7782 ( .A1(n7765), .A2(n7475), .ZN(n7764) );
  XOR2_X1 U7783 ( .A(n7766), .B(n7767), .Z(n7765) );
  AND2_X1 U7784 ( .A1(n7768), .A2(n7769), .ZN(n7767) );
  NAND2_X1 U7785 ( .A1(n7770), .A2(operation), .ZN(n7763) );
  XOR2_X1 U7786 ( .A(n7771), .B(n7772), .Z(n7770) );
  XOR2_X1 U7787 ( .A(n7773), .B(n7774), .Z(n7771) );
  NOR2_X1 U7788 ( .A1(n7775), .A2(n7508), .ZN(n7774) );
  NAND2_X1 U7789 ( .A1(n7776), .A2(n7777), .ZN(Result_45_) );
  NAND2_X1 U7790 ( .A1(n7778), .A2(n7475), .ZN(n7777) );
  NAND2_X1 U7791 ( .A1(n7779), .A2(n7780), .ZN(n7778) );
  NAND2_X1 U7792 ( .A1(n7781), .A2(n7782), .ZN(n7780) );
  NOR2_X1 U7793 ( .A1(n7783), .A2(n7784), .ZN(n7779) );
  NOR2_X1 U7794 ( .A1(b_13_), .A2(n7785), .ZN(n7784) );
  XOR2_X1 U7795 ( .A(n7786), .B(n7782), .Z(n7785) );
  NOR2_X1 U7796 ( .A1(n7787), .A2(n7788), .ZN(n7783) );
  OR2_X1 U7797 ( .A1(n7782), .A2(a_13_), .ZN(n7788) );
  NAND2_X1 U7798 ( .A1(n7789), .A2(operation), .ZN(n7776) );
  XNOR2_X1 U7799 ( .A(n7790), .B(n7791), .ZN(n7789) );
  XOR2_X1 U7800 ( .A(n7792), .B(n7793), .Z(n7791) );
  NAND2_X1 U7801 ( .A1(b_31_), .A2(a_13_), .ZN(n7793) );
  NAND2_X1 U7802 ( .A1(n7794), .A2(n7795), .ZN(Result_44_) );
  NAND2_X1 U7803 ( .A1(n7796), .A2(n7475), .ZN(n7795) );
  XOR2_X1 U7804 ( .A(n7797), .B(n7798), .Z(n7796) );
  AND2_X1 U7805 ( .A1(n7799), .A2(n7800), .ZN(n7798) );
  NAND2_X1 U7806 ( .A1(n7801), .A2(operation), .ZN(n7794) );
  XOR2_X1 U7807 ( .A(n7802), .B(n7803), .Z(n7801) );
  XOR2_X1 U7808 ( .A(n7804), .B(n7805), .Z(n7802) );
  NOR2_X1 U7809 ( .A1(n7806), .A2(n7508), .ZN(n7805) );
  NAND2_X1 U7810 ( .A1(n7807), .A2(n7808), .ZN(Result_43_) );
  NAND2_X1 U7811 ( .A1(n7809), .A2(n7475), .ZN(n7808) );
  NAND2_X1 U7812 ( .A1(n7810), .A2(n7811), .ZN(n7809) );
  NAND2_X1 U7813 ( .A1(n7812), .A2(n7813), .ZN(n7811) );
  NOR2_X1 U7814 ( .A1(n7814), .A2(n7815), .ZN(n7810) );
  NOR2_X1 U7815 ( .A1(b_11_), .A2(n7816), .ZN(n7815) );
  XOR2_X1 U7816 ( .A(n7817), .B(n7813), .Z(n7816) );
  NOR2_X1 U7817 ( .A1(n7818), .A2(n7819), .ZN(n7814) );
  OR2_X1 U7818 ( .A1(n7813), .A2(a_11_), .ZN(n7819) );
  NAND2_X1 U7819 ( .A1(n7820), .A2(operation), .ZN(n7807) );
  XOR2_X1 U7820 ( .A(n7821), .B(n7822), .Z(n7820) );
  XOR2_X1 U7821 ( .A(n7823), .B(n7824), .Z(n7821) );
  NOR2_X1 U7822 ( .A1(n7817), .A2(n7508), .ZN(n7824) );
  NAND2_X1 U7823 ( .A1(n7825), .A2(n7826), .ZN(Result_42_) );
  NAND2_X1 U7824 ( .A1(n7827), .A2(n7475), .ZN(n7826) );
  XNOR2_X1 U7825 ( .A(n7828), .B(n7829), .ZN(n7827) );
  NOR2_X1 U7826 ( .A1(n7830), .A2(n7831), .ZN(n7829) );
  NAND2_X1 U7827 ( .A1(n7832), .A2(operation), .ZN(n7825) );
  XOR2_X1 U7828 ( .A(n7833), .B(n7834), .Z(n7832) );
  XOR2_X1 U7829 ( .A(n7835), .B(n7836), .Z(n7833) );
  NOR2_X1 U7830 ( .A1(n7837), .A2(n7508), .ZN(n7836) );
  NAND2_X1 U7831 ( .A1(n7838), .A2(n7839), .ZN(Result_41_) );
  NAND2_X1 U7832 ( .A1(n7840), .A2(n7475), .ZN(n7839) );
  NAND2_X1 U7833 ( .A1(n7841), .A2(n7842), .ZN(n7840) );
  NAND2_X1 U7834 ( .A1(n7843), .A2(n7844), .ZN(n7842) );
  NOR2_X1 U7835 ( .A1(n7845), .A2(n7846), .ZN(n7841) );
  NOR2_X1 U7836 ( .A1(b_9_), .A2(n7847), .ZN(n7846) );
  XOR2_X1 U7837 ( .A(n7848), .B(n7844), .Z(n7847) );
  NOR2_X1 U7838 ( .A1(n7849), .A2(n7850), .ZN(n7845) );
  NAND2_X1 U7839 ( .A1(n7851), .A2(n7848), .ZN(n7850) );
  NAND2_X1 U7840 ( .A1(n7852), .A2(operation), .ZN(n7838) );
  XNOR2_X1 U7841 ( .A(n7853), .B(n7854), .ZN(n7852) );
  XOR2_X1 U7842 ( .A(n7855), .B(n7856), .Z(n7854) );
  NAND2_X1 U7843 ( .A1(b_31_), .A2(a_9_), .ZN(n7856) );
  NAND2_X1 U7844 ( .A1(n7857), .A2(n7858), .ZN(Result_40_) );
  NAND2_X1 U7845 ( .A1(n7859), .A2(n7475), .ZN(n7858) );
  XOR2_X1 U7846 ( .A(n7860), .B(n7861), .Z(n7859) );
  AND2_X1 U7847 ( .A1(n7862), .A2(n7863), .ZN(n7861) );
  NAND2_X1 U7848 ( .A1(n7864), .A2(operation), .ZN(n7857) );
  XNOR2_X1 U7849 ( .A(n7865), .B(n7866), .ZN(n7864) );
  XOR2_X1 U7850 ( .A(n7867), .B(n7868), .Z(n7866) );
  NAND2_X1 U7851 ( .A1(b_31_), .A2(a_8_), .ZN(n7868) );
  NOR2_X1 U7852 ( .A1(n7475), .A2(n7869), .ZN(Result_3_) );
  XOR2_X1 U7853 ( .A(n7870), .B(n7871), .Z(n7869) );
  NAND2_X1 U7854 ( .A1(n7872), .A2(n7873), .ZN(n7871) );
  NAND2_X1 U7855 ( .A1(n7874), .A2(n7875), .ZN(Result_39_) );
  NAND2_X1 U7856 ( .A1(n7876), .A2(n7475), .ZN(n7875) );
  NAND2_X1 U7857 ( .A1(n7877), .A2(n7878), .ZN(n7876) );
  NAND2_X1 U7858 ( .A1(n7879), .A2(n7880), .ZN(n7878) );
  NOR2_X1 U7859 ( .A1(n7881), .A2(n7882), .ZN(n7877) );
  NOR2_X1 U7860 ( .A1(b_7_), .A2(n7883), .ZN(n7882) );
  XOR2_X1 U7861 ( .A(n7884), .B(n7880), .Z(n7883) );
  NOR2_X1 U7862 ( .A1(n7885), .A2(n7886), .ZN(n7881) );
  OR2_X1 U7863 ( .A1(n7880), .A2(a_7_), .ZN(n7886) );
  NAND2_X1 U7864 ( .A1(n7887), .A2(operation), .ZN(n7874) );
  XOR2_X1 U7865 ( .A(n7888), .B(n7889), .Z(n7887) );
  XOR2_X1 U7866 ( .A(n7890), .B(n7891), .Z(n7888) );
  NOR2_X1 U7867 ( .A1(n7884), .A2(n7508), .ZN(n7891) );
  NAND2_X1 U7868 ( .A1(n7892), .A2(n7893), .ZN(Result_38_) );
  NAND2_X1 U7869 ( .A1(n7894), .A2(n7475), .ZN(n7893) );
  XOR2_X1 U7870 ( .A(n7895), .B(n7896), .Z(n7894) );
  AND2_X1 U7871 ( .A1(n7897), .A2(n7898), .ZN(n7896) );
  NAND2_X1 U7872 ( .A1(n7899), .A2(operation), .ZN(n7892) );
  XNOR2_X1 U7873 ( .A(n7900), .B(n7901), .ZN(n7899) );
  XOR2_X1 U7874 ( .A(n7902), .B(n7903), .Z(n7901) );
  NAND2_X1 U7875 ( .A1(b_31_), .A2(a_6_), .ZN(n7903) );
  NAND2_X1 U7876 ( .A1(n7904), .A2(n7905), .ZN(Result_37_) );
  NAND2_X1 U7877 ( .A1(n7906), .A2(n7475), .ZN(n7905) );
  NAND2_X1 U7878 ( .A1(n7907), .A2(n7908), .ZN(n7906) );
  NAND2_X1 U7879 ( .A1(n7909), .A2(n7910), .ZN(n7908) );
  NOR2_X1 U7880 ( .A1(n7911), .A2(n7912), .ZN(n7907) );
  NOR2_X1 U7881 ( .A1(b_5_), .A2(n7913), .ZN(n7912) );
  XOR2_X1 U7882 ( .A(n7914), .B(n7910), .Z(n7913) );
  NOR2_X1 U7883 ( .A1(n7915), .A2(n7916), .ZN(n7911) );
  OR2_X1 U7884 ( .A1(n7910), .A2(a_5_), .ZN(n7916) );
  NAND2_X1 U7885 ( .A1(n7917), .A2(operation), .ZN(n7904) );
  XOR2_X1 U7886 ( .A(n7918), .B(n7919), .Z(n7917) );
  XOR2_X1 U7887 ( .A(n7920), .B(n7921), .Z(n7918) );
  NOR2_X1 U7888 ( .A1(n7914), .A2(n7508), .ZN(n7921) );
  NAND2_X1 U7889 ( .A1(n7922), .A2(n7923), .ZN(Result_36_) );
  NAND2_X1 U7890 ( .A1(n7924), .A2(n7475), .ZN(n7923) );
  XOR2_X1 U7891 ( .A(n7925), .B(n7926), .Z(n7924) );
  AND2_X1 U7892 ( .A1(n7927), .A2(n7928), .ZN(n7926) );
  NAND2_X1 U7893 ( .A1(n7929), .A2(operation), .ZN(n7922) );
  XOR2_X1 U7894 ( .A(n7930), .B(n7931), .Z(n7929) );
  XOR2_X1 U7895 ( .A(n7932), .B(n7933), .Z(n7930) );
  NOR2_X1 U7896 ( .A1(n7934), .A2(n7508), .ZN(n7933) );
  NAND2_X1 U7897 ( .A1(n7935), .A2(n7936), .ZN(Result_35_) );
  NAND2_X1 U7898 ( .A1(n7937), .A2(n7475), .ZN(n7936) );
  NAND2_X1 U7899 ( .A1(n7938), .A2(n7939), .ZN(n7937) );
  NAND2_X1 U7900 ( .A1(n7940), .A2(n7941), .ZN(n7939) );
  NOR2_X1 U7901 ( .A1(n7942), .A2(n7943), .ZN(n7938) );
  NOR2_X1 U7902 ( .A1(b_3_), .A2(n7944), .ZN(n7943) );
  XOR2_X1 U7903 ( .A(n7945), .B(n7941), .Z(n7944) );
  NOR2_X1 U7904 ( .A1(n7946), .A2(n7947), .ZN(n7942) );
  OR2_X1 U7905 ( .A1(n7941), .A2(a_3_), .ZN(n7947) );
  NAND2_X1 U7906 ( .A1(n7948), .A2(operation), .ZN(n7935) );
  XNOR2_X1 U7907 ( .A(n7949), .B(n7950), .ZN(n7948) );
  XOR2_X1 U7908 ( .A(n7951), .B(n7952), .Z(n7950) );
  NAND2_X1 U7909 ( .A1(b_31_), .A2(a_3_), .ZN(n7952) );
  NAND2_X1 U7910 ( .A1(n7953), .A2(n7954), .ZN(Result_34_) );
  NAND2_X1 U7911 ( .A1(n7955), .A2(n7475), .ZN(n7954) );
  XOR2_X1 U7912 ( .A(n7956), .B(n7957), .Z(n7955) );
  AND2_X1 U7913 ( .A1(n7958), .A2(n7959), .ZN(n7957) );
  NAND2_X1 U7914 ( .A1(n7960), .A2(operation), .ZN(n7953) );
  XOR2_X1 U7915 ( .A(n7961), .B(n7962), .Z(n7960) );
  XOR2_X1 U7916 ( .A(n7963), .B(n7964), .Z(n7961) );
  NOR2_X1 U7917 ( .A1(n7965), .A2(n7508), .ZN(n7964) );
  NAND2_X1 U7918 ( .A1(n7966), .A2(n7967), .ZN(Result_33_) );
  NAND2_X1 U7919 ( .A1(n7968), .A2(operation), .ZN(n7967) );
  XOR2_X1 U7920 ( .A(n7969), .B(n7970), .Z(n7968) );
  XOR2_X1 U7921 ( .A(n7971), .B(n7972), .Z(n7969) );
  NOR2_X1 U7922 ( .A1(n7973), .A2(n7508), .ZN(n7972) );
  NAND2_X1 U7923 ( .A1(n7974), .A2(n7475), .ZN(n7966) );
  NAND2_X1 U7924 ( .A1(n7975), .A2(n7976), .ZN(n7974) );
  NAND2_X1 U7925 ( .A1(n7977), .A2(n7978), .ZN(n7976) );
  OR2_X1 U7926 ( .A1(n7979), .A2(n7980), .ZN(n7977) );
  NAND2_X1 U7927 ( .A1(n7981), .A2(n7982), .ZN(n7975) );
  INV_X1 U7928 ( .A(n7978), .ZN(n7982) );
  XOR2_X1 U7929 ( .A(b_1_), .B(a_1_), .Z(n7981) );
  NAND2_X1 U7930 ( .A1(n7983), .A2(n7984), .ZN(Result_32_) );
  NAND2_X1 U7931 ( .A1(n7985), .A2(n7475), .ZN(n7984) );
  XOR2_X1 U7932 ( .A(n7986), .B(n7987), .Z(n7985) );
  NOR2_X1 U7933 ( .A1(n7988), .A2(n7989), .ZN(n7987) );
  NOR2_X1 U7934 ( .A1(b_0_), .A2(a_0_), .ZN(n7988) );
  NOR2_X1 U7935 ( .A1(n7980), .A2(n7990), .ZN(n7986) );
  NOR2_X1 U7936 ( .A1(n7979), .A2(n7978), .ZN(n7990) );
  NAND2_X1 U7937 ( .A1(n7959), .A2(n7991), .ZN(n7978) );
  NAND2_X1 U7938 ( .A1(n7958), .A2(n7956), .ZN(n7991) );
  NAND2_X1 U7939 ( .A1(n7992), .A2(n7993), .ZN(n7956) );
  NAND2_X1 U7940 ( .A1(n7994), .A2(n7941), .ZN(n7993) );
  NAND2_X1 U7941 ( .A1(n7928), .A2(n7995), .ZN(n7941) );
  NAND2_X1 U7942 ( .A1(n7927), .A2(n7925), .ZN(n7995) );
  NAND2_X1 U7943 ( .A1(n7996), .A2(n7997), .ZN(n7925) );
  NAND2_X1 U7944 ( .A1(n7998), .A2(n7910), .ZN(n7997) );
  NAND2_X1 U7945 ( .A1(n7898), .A2(n7999), .ZN(n7910) );
  NAND2_X1 U7946 ( .A1(n7897), .A2(n7895), .ZN(n7999) );
  NAND2_X1 U7947 ( .A1(n8000), .A2(n8001), .ZN(n7895) );
  NAND2_X1 U7948 ( .A1(n8002), .A2(n7880), .ZN(n8001) );
  NAND2_X1 U7949 ( .A1(n7863), .A2(n8003), .ZN(n7880) );
  NAND2_X1 U7950 ( .A1(n7862), .A2(n7860), .ZN(n8003) );
  NAND2_X1 U7951 ( .A1(n8004), .A2(n8005), .ZN(n7860) );
  NAND2_X1 U7952 ( .A1(n8006), .A2(n7844), .ZN(n8005) );
  INV_X1 U7953 ( .A(n7851), .ZN(n7844) );
  NOR2_X1 U7954 ( .A1(n7831), .A2(n8007), .ZN(n7851) );
  NOR2_X1 U7955 ( .A1(n7830), .A2(n7828), .ZN(n8007) );
  NOR2_X1 U7956 ( .A1(n7812), .A2(n8008), .ZN(n7828) );
  AND2_X1 U7957 ( .A1(n8009), .A2(n7813), .ZN(n8008) );
  NAND2_X1 U7958 ( .A1(n7800), .A2(n8010), .ZN(n7813) );
  NAND2_X1 U7959 ( .A1(n7799), .A2(n7797), .ZN(n8010) );
  NAND2_X1 U7960 ( .A1(n8011), .A2(n8012), .ZN(n7797) );
  NAND2_X1 U7961 ( .A1(n8013), .A2(n7782), .ZN(n8012) );
  NAND2_X1 U7962 ( .A1(n7769), .A2(n8014), .ZN(n7782) );
  NAND2_X1 U7963 ( .A1(n7768), .A2(n7766), .ZN(n8014) );
  NAND2_X1 U7964 ( .A1(n8015), .A2(n8016), .ZN(n7766) );
  NAND2_X1 U7965 ( .A1(n8017), .A2(n7750), .ZN(n8016) );
  INV_X1 U7966 ( .A(n7757), .ZN(n7750) );
  NOR2_X1 U7967 ( .A1(n7737), .A2(n8018), .ZN(n7757) );
  NOR2_X1 U7968 ( .A1(n7736), .A2(n7734), .ZN(n8018) );
  AND2_X1 U7969 ( .A1(n8019), .A2(n8020), .ZN(n7734) );
  NAND2_X1 U7970 ( .A1(n8021), .A2(n7719), .ZN(n8020) );
  NAND2_X1 U7971 ( .A1(n7701), .A2(n8022), .ZN(n7719) );
  NAND2_X1 U7972 ( .A1(n7700), .A2(n7698), .ZN(n8022) );
  NAND2_X1 U7973 ( .A1(n8023), .A2(n8024), .ZN(n7698) );
  NAND2_X1 U7974 ( .A1(n8025), .A2(n7683), .ZN(n8024) );
  NAND2_X1 U7975 ( .A1(n7670), .A2(n8026), .ZN(n7683) );
  NAND2_X1 U7976 ( .A1(n7669), .A2(n7667), .ZN(n8026) );
  NAND2_X1 U7977 ( .A1(n8027), .A2(n8028), .ZN(n7667) );
  NAND2_X1 U7978 ( .A1(n8029), .A2(n7652), .ZN(n8028) );
  NAND2_X1 U7979 ( .A1(n7639), .A2(n8030), .ZN(n7652) );
  NAND2_X1 U7980 ( .A1(n7638), .A2(n7636), .ZN(n8030) );
  NAND2_X1 U7981 ( .A1(n8031), .A2(n8032), .ZN(n7636) );
  NAND2_X1 U7982 ( .A1(n8033), .A2(n7620), .ZN(n8032) );
  INV_X1 U7983 ( .A(n7627), .ZN(n7620) );
  NOR2_X1 U7984 ( .A1(n7607), .A2(n8034), .ZN(n7627) );
  NOR2_X1 U7985 ( .A1(n7606), .A2(n7604), .ZN(n8034) );
  NOR2_X1 U7986 ( .A1(n7588), .A2(n8035), .ZN(n7604) );
  AND2_X1 U7987 ( .A1(n8036), .A2(n7589), .ZN(n8035) );
  NAND2_X1 U7988 ( .A1(n7577), .A2(n8037), .ZN(n7589) );
  NAND2_X1 U7989 ( .A1(n7576), .A2(n7574), .ZN(n8037) );
  NAND2_X1 U7990 ( .A1(n8038), .A2(n8039), .ZN(n7574) );
  NAND2_X1 U7991 ( .A1(n8040), .A2(n7559), .ZN(n8039) );
  NAND2_X1 U7992 ( .A1(n7540), .A2(n8041), .ZN(n7559) );
  NAND2_X1 U7993 ( .A1(n7541), .A2(n7539), .ZN(n8041) );
  NAND2_X1 U7994 ( .A1(n8042), .A2(n8043), .ZN(n7539) );
  NAND2_X1 U7995 ( .A1(n8044), .A2(n7522), .ZN(n8043) );
  NAND2_X1 U7996 ( .A1(n8045), .A2(n8046), .ZN(n7522) );
  NAND2_X1 U7997 ( .A1(b_30_), .A2(n8047), .ZN(n8046) );
  OR2_X1 U7998 ( .A1(a_30_), .A2(n7499), .ZN(n8047) );
  NOR2_X1 U7999 ( .A1(n7508), .A2(n8048), .ZN(n7499) );
  INV_X1 U8000 ( .A(b_31_), .ZN(n7508) );
  NAND2_X1 U8001 ( .A1(b_31_), .A2(n8049), .ZN(n8045) );
  NAND2_X1 U8002 ( .A1(n7527), .A2(n7529), .ZN(n8044) );
  NAND2_X1 U8003 ( .A1(n8050), .A2(n7547), .ZN(n7541) );
  NAND2_X1 U8004 ( .A1(n7564), .A2(n7563), .ZN(n8040) );
  NAND2_X1 U8005 ( .A1(n8051), .A2(n8052), .ZN(n7576) );
  NAND2_X1 U8006 ( .A1(n7594), .A2(n7593), .ZN(n8036) );
  NOR2_X1 U8007 ( .A1(b_24_), .A2(a_24_), .ZN(n7606) );
  NAND2_X1 U8008 ( .A1(n7625), .A2(n7624), .ZN(n8033) );
  NAND2_X1 U8009 ( .A1(n8053), .A2(n7645), .ZN(n7638) );
  NAND2_X1 U8010 ( .A1(n7657), .A2(n7656), .ZN(n8029) );
  NAND2_X1 U8011 ( .A1(n8054), .A2(n7676), .ZN(n7669) );
  NAND2_X1 U8012 ( .A1(n7688), .A2(n7687), .ZN(n8025) );
  NAND2_X1 U8013 ( .A1(n8055), .A2(n7707), .ZN(n7700) );
  NAND2_X1 U8014 ( .A1(n7724), .A2(n7723), .ZN(n8021) );
  NOR2_X1 U8015 ( .A1(b_16_), .A2(a_16_), .ZN(n7736) );
  NAND2_X1 U8016 ( .A1(n7755), .A2(n7754), .ZN(n8017) );
  NAND2_X1 U8017 ( .A1(n8056), .A2(n7775), .ZN(n7768) );
  NAND2_X1 U8018 ( .A1(n7787), .A2(n7786), .ZN(n8013) );
  NAND2_X1 U8019 ( .A1(n8057), .A2(n7806), .ZN(n7799) );
  NAND2_X1 U8020 ( .A1(n7818), .A2(n7817), .ZN(n8009) );
  NOR2_X1 U8021 ( .A1(b_10_), .A2(a_10_), .ZN(n7830) );
  NAND2_X1 U8022 ( .A1(n7849), .A2(n7848), .ZN(n8006) );
  NAND2_X1 U8023 ( .A1(n8058), .A2(n8059), .ZN(n7862) );
  NAND2_X1 U8024 ( .A1(n7885), .A2(n7884), .ZN(n8002) );
  NAND2_X1 U8025 ( .A1(n8060), .A2(n8061), .ZN(n7897) );
  NAND2_X1 U8026 ( .A1(n7915), .A2(n7914), .ZN(n7998) );
  NAND2_X1 U8027 ( .A1(n8062), .A2(n7934), .ZN(n7927) );
  NAND2_X1 U8028 ( .A1(n7946), .A2(n7945), .ZN(n7994) );
  NAND2_X1 U8029 ( .A1(n8063), .A2(n7965), .ZN(n7958) );
  NOR2_X1 U8030 ( .A1(b_1_), .A2(a_1_), .ZN(n7980) );
  NAND2_X1 U8031 ( .A1(n8064), .A2(operation), .ZN(n7983) );
  XNOR2_X1 U8032 ( .A(n8065), .B(n8066), .ZN(n8064) );
  XOR2_X1 U8033 ( .A(n8067), .B(n8068), .Z(n8066) );
  NAND2_X1 U8034 ( .A1(b_31_), .A2(a_0_), .ZN(n8068) );
  NOR2_X1 U8035 ( .A1(n7475), .A2(n8069), .ZN(Result_31_) );
  XOR2_X1 U8036 ( .A(n8070), .B(n8071), .Z(n8069) );
  NOR2_X1 U8037 ( .A1(n7475), .A2(n8072), .ZN(Result_30_) );
  NAND2_X1 U8038 ( .A1(n8073), .A2(n8074), .ZN(n8072) );
  NAND2_X1 U8039 ( .A1(n8075), .A2(n8076), .ZN(n8073) );
  NAND2_X1 U8040 ( .A1(n8071), .A2(n8077), .ZN(n8076) );
  NOR2_X1 U8041 ( .A1(n7475), .A2(n8078), .ZN(Result_2_) );
  XOR2_X1 U8042 ( .A(n8079), .B(n8080), .Z(n8078) );
  NAND2_X1 U8043 ( .A1(n8081), .A2(n8082), .ZN(n8080) );
  NOR2_X1 U8044 ( .A1(n8083), .A2(n7475), .ZN(Result_29_) );
  XNOR2_X1 U8045 ( .A(n8084), .B(n8085), .ZN(n8083) );
  AND2_X1 U8046 ( .A1(n8086), .A2(n8087), .ZN(n8085) );
  NOR2_X1 U8047 ( .A1(n7475), .A2(n8088), .ZN(Result_28_) );
  XNOR2_X1 U8048 ( .A(n8089), .B(n8090), .ZN(n8088) );
  AND2_X1 U8049 ( .A1(n8091), .A2(n8092), .ZN(n8090) );
  NOR2_X1 U8050 ( .A1(n7475), .A2(n8093), .ZN(Result_27_) );
  XOR2_X1 U8051 ( .A(n8094), .B(n8095), .Z(n8093) );
  NAND2_X1 U8052 ( .A1(n8096), .A2(n8097), .ZN(n8095) );
  NOR2_X1 U8053 ( .A1(n7475), .A2(n8098), .ZN(Result_26_) );
  XOR2_X1 U8054 ( .A(n8099), .B(n8100), .Z(n8098) );
  NAND2_X1 U8055 ( .A1(n8101), .A2(n8102), .ZN(n8100) );
  NOR2_X1 U8056 ( .A1(n7475), .A2(n8103), .ZN(Result_25_) );
  XOR2_X1 U8057 ( .A(n8104), .B(n8105), .Z(n8103) );
  NAND2_X1 U8058 ( .A1(n8106), .A2(n8107), .ZN(n8105) );
  NOR2_X1 U8059 ( .A1(n7475), .A2(n8108), .ZN(Result_24_) );
  XOR2_X1 U8060 ( .A(n8109), .B(n8110), .Z(n8108) );
  NAND2_X1 U8061 ( .A1(n8111), .A2(n8112), .ZN(n8110) );
  NOR2_X1 U8062 ( .A1(n7475), .A2(n8113), .ZN(Result_23_) );
  XOR2_X1 U8063 ( .A(n8114), .B(n8115), .Z(n8113) );
  NAND2_X1 U8064 ( .A1(n8116), .A2(n8117), .ZN(n8115) );
  NOR2_X1 U8065 ( .A1(n7475), .A2(n8118), .ZN(Result_22_) );
  XOR2_X1 U8066 ( .A(n8119), .B(n8120), .Z(n8118) );
  NAND2_X1 U8067 ( .A1(n8121), .A2(n8122), .ZN(n8120) );
  NOR2_X1 U8068 ( .A1(n7475), .A2(n8123), .ZN(Result_21_) );
  XOR2_X1 U8069 ( .A(n8124), .B(n8125), .Z(n8123) );
  NAND2_X1 U8070 ( .A1(n8126), .A2(n8127), .ZN(n8125) );
  NOR2_X1 U8071 ( .A1(n7475), .A2(n8128), .ZN(Result_20_) );
  XOR2_X1 U8072 ( .A(n8129), .B(n8130), .Z(n8128) );
  NAND2_X1 U8073 ( .A1(n8131), .A2(n8132), .ZN(n8130) );
  NOR2_X1 U8074 ( .A1(n7475), .A2(n8133), .ZN(Result_1_) );
  XOR2_X1 U8075 ( .A(n8134), .B(n8135), .Z(n8133) );
  NAND2_X1 U8076 ( .A1(n8136), .A2(n8137), .ZN(n8135) );
  NOR2_X1 U8077 ( .A1(n7475), .A2(n8138), .ZN(Result_19_) );
  XOR2_X1 U8078 ( .A(n8139), .B(n8140), .Z(n8138) );
  NAND2_X1 U8079 ( .A1(n8141), .A2(n8142), .ZN(n8140) );
  NOR2_X1 U8080 ( .A1(n7475), .A2(n8143), .ZN(Result_18_) );
  XOR2_X1 U8081 ( .A(n8144), .B(n8145), .Z(n8143) );
  NAND2_X1 U8082 ( .A1(n8146), .A2(n8147), .ZN(n8145) );
  NOR2_X1 U8083 ( .A1(n7475), .A2(n8148), .ZN(Result_17_) );
  XOR2_X1 U8084 ( .A(n8149), .B(n8150), .Z(n8148) );
  NAND2_X1 U8085 ( .A1(n8151), .A2(n8152), .ZN(n8150) );
  NOR2_X1 U8086 ( .A1(n7475), .A2(n8153), .ZN(Result_16_) );
  XOR2_X1 U8087 ( .A(n8154), .B(n8155), .Z(n8153) );
  NAND2_X1 U8088 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  NOR2_X1 U8089 ( .A1(n7475), .A2(n8158), .ZN(Result_15_) );
  XOR2_X1 U8090 ( .A(n8159), .B(n8160), .Z(n8158) );
  NAND2_X1 U8091 ( .A1(n8161), .A2(n8162), .ZN(n8160) );
  NOR2_X1 U8092 ( .A1(n7475), .A2(n8163), .ZN(Result_14_) );
  XOR2_X1 U8093 ( .A(n8164), .B(n8165), .Z(n8163) );
  NAND2_X1 U8094 ( .A1(n8166), .A2(n8167), .ZN(n8165) );
  NOR2_X1 U8095 ( .A1(n7475), .A2(n8168), .ZN(Result_13_) );
  XOR2_X1 U8096 ( .A(n8169), .B(n8170), .Z(n8168) );
  NAND2_X1 U8097 ( .A1(n8171), .A2(n8172), .ZN(n8170) );
  NOR2_X1 U8098 ( .A1(n7475), .A2(n8173), .ZN(Result_12_) );
  XOR2_X1 U8099 ( .A(n8174), .B(n8175), .Z(n8173) );
  NAND2_X1 U8100 ( .A1(n8176), .A2(n8177), .ZN(n8175) );
  NOR2_X1 U8101 ( .A1(n7475), .A2(n8178), .ZN(Result_11_) );
  XOR2_X1 U8102 ( .A(n8179), .B(n8180), .Z(n8178) );
  NAND2_X1 U8103 ( .A1(n8181), .A2(n8182), .ZN(n8180) );
  NOR2_X1 U8104 ( .A1(n7475), .A2(n8183), .ZN(Result_10_) );
  XOR2_X1 U8105 ( .A(n8184), .B(n8185), .Z(n8183) );
  NAND2_X1 U8106 ( .A1(n8186), .A2(n8187), .ZN(n8185) );
  NOR2_X1 U8107 ( .A1(n8188), .A2(n7475), .ZN(Result_0_) );
  NOR2_X1 U8108 ( .A1(n8189), .A2(n8190), .ZN(n8188) );
  NAND2_X1 U8109 ( .A1(n8191), .A2(n8137), .ZN(n8190) );
  NAND2_X1 U8110 ( .A1(n8192), .A2(n8193), .ZN(n8137) );
  AND2_X1 U8111 ( .A1(n8194), .A2(n8195), .ZN(n8193) );
  AND2_X1 U8112 ( .A1(n8196), .A2(n7989), .ZN(n8192) );
  NAND2_X1 U8113 ( .A1(n8136), .A2(n8134), .ZN(n8191) );
  NAND2_X1 U8114 ( .A1(n8081), .A2(n8197), .ZN(n8134) );
  NAND2_X1 U8115 ( .A1(n8082), .A2(n8079), .ZN(n8197) );
  NAND2_X1 U8116 ( .A1(n7872), .A2(n8198), .ZN(n8079) );
  NAND2_X1 U8117 ( .A1(n7873), .A2(n7870), .ZN(n8198) );
  NAND2_X1 U8118 ( .A1(n7711), .A2(n8199), .ZN(n7870) );
  NAND2_X1 U8119 ( .A1(n7712), .A2(n7709), .ZN(n8199) );
  NAND2_X1 U8120 ( .A1(n7551), .A2(n8200), .ZN(n7709) );
  NAND2_X1 U8121 ( .A1(n7552), .A2(n7549), .ZN(n8200) );
  NAND2_X1 U8122 ( .A1(n7494), .A2(n8201), .ZN(n7549) );
  NAND2_X1 U8123 ( .A1(n7495), .A2(n7492), .ZN(n8201) );
  NAND2_X1 U8124 ( .A1(n7489), .A2(n8202), .ZN(n7492) );
  NAND2_X1 U8125 ( .A1(n7490), .A2(n7487), .ZN(n8202) );
  NAND2_X1 U8126 ( .A1(n7484), .A2(n8203), .ZN(n7487) );
  NAND2_X1 U8127 ( .A1(n7485), .A2(n7482), .ZN(n8203) );
  NAND2_X1 U8128 ( .A1(n7479), .A2(n8204), .ZN(n7482) );
  NAND2_X1 U8129 ( .A1(n7480), .A2(n7477), .ZN(n8204) );
  NAND2_X1 U8130 ( .A1(n8186), .A2(n8205), .ZN(n7477) );
  NAND2_X1 U8131 ( .A1(n8184), .A2(n8187), .ZN(n8205) );
  NAND2_X1 U8132 ( .A1(n8206), .A2(n8207), .ZN(n8187) );
  XOR2_X1 U8133 ( .A(n8208), .B(n8209), .Z(n8206) );
  NAND2_X1 U8134 ( .A1(n8181), .A2(n8210), .ZN(n8184) );
  NAND2_X1 U8135 ( .A1(n8179), .A2(n8182), .ZN(n8210) );
  NAND2_X1 U8136 ( .A1(n8211), .A2(n8212), .ZN(n8182) );
  NAND2_X1 U8137 ( .A1(n8213), .A2(n8207), .ZN(n8212) );
  INV_X1 U8138 ( .A(n8214), .ZN(n8207) );
  NAND2_X1 U8139 ( .A1(n8215), .A2(n8216), .ZN(n8213) );
  OR2_X1 U8140 ( .A1(n8217), .A2(n8218), .ZN(n8211) );
  NAND2_X1 U8141 ( .A1(n8176), .A2(n8219), .ZN(n8179) );
  NAND2_X1 U8142 ( .A1(n8174), .A2(n8177), .ZN(n8219) );
  NAND2_X1 U8143 ( .A1(n8220), .A2(n8221), .ZN(n8177) );
  XOR2_X1 U8144 ( .A(n8222), .B(n8217), .Z(n8220) );
  NAND2_X1 U8145 ( .A1(n8171), .A2(n8223), .ZN(n8174) );
  NAND2_X1 U8146 ( .A1(n8169), .A2(n8172), .ZN(n8223) );
  NAND2_X1 U8147 ( .A1(n8224), .A2(n8225), .ZN(n8172) );
  NAND2_X1 U8148 ( .A1(n8226), .A2(n8221), .ZN(n8225) );
  INV_X1 U8149 ( .A(n8227), .ZN(n8221) );
  NAND2_X1 U8150 ( .A1(n8228), .A2(n8229), .ZN(n8226) );
  NAND2_X1 U8151 ( .A1(n8230), .A2(n8231), .ZN(n8224) );
  NAND2_X1 U8152 ( .A1(n8166), .A2(n8232), .ZN(n8169) );
  NAND2_X1 U8153 ( .A1(n8167), .A2(n8164), .ZN(n8232) );
  NAND2_X1 U8154 ( .A1(n8161), .A2(n8233), .ZN(n8164) );
  NAND2_X1 U8155 ( .A1(n8162), .A2(n8159), .ZN(n8233) );
  NAND2_X1 U8156 ( .A1(n8156), .A2(n8234), .ZN(n8159) );
  NAND2_X1 U8157 ( .A1(n8154), .A2(n8157), .ZN(n8234) );
  NAND2_X1 U8158 ( .A1(n8235), .A2(n8236), .ZN(n8157) );
  NAND2_X1 U8159 ( .A1(n8237), .A2(n8238), .ZN(n8236) );
  XOR2_X1 U8160 ( .A(n8239), .B(n8240), .Z(n8235) );
  NAND2_X1 U8161 ( .A1(n8151), .A2(n8241), .ZN(n8154) );
  NAND2_X1 U8162 ( .A1(n8152), .A2(n8149), .ZN(n8241) );
  NAND2_X1 U8163 ( .A1(n8146), .A2(n8242), .ZN(n8149) );
  NAND2_X1 U8164 ( .A1(n8144), .A2(n8147), .ZN(n8242) );
  NAND2_X1 U8165 ( .A1(n8243), .A2(n8244), .ZN(n8147) );
  NAND2_X1 U8166 ( .A1(n8245), .A2(n8246), .ZN(n8244) );
  XNOR2_X1 U8167 ( .A(n8247), .B(n8248), .ZN(n8243) );
  NAND2_X1 U8168 ( .A1(n8141), .A2(n8249), .ZN(n8144) );
  NAND2_X1 U8169 ( .A1(n8139), .A2(n8142), .ZN(n8249) );
  NAND2_X1 U8170 ( .A1(n8250), .A2(n8251), .ZN(n8142) );
  NAND2_X1 U8171 ( .A1(n8252), .A2(n8253), .ZN(n8251) );
  XOR2_X1 U8172 ( .A(n8246), .B(n8254), .Z(n8250) );
  NAND2_X1 U8173 ( .A1(n8131), .A2(n8255), .ZN(n8139) );
  NAND2_X1 U8174 ( .A1(n8129), .A2(n8132), .ZN(n8255) );
  NAND2_X1 U8175 ( .A1(n8256), .A2(n8257), .ZN(n8132) );
  NAND2_X1 U8176 ( .A1(n8127), .A2(n8258), .ZN(n8129) );
  NAND2_X1 U8177 ( .A1(n8126), .A2(n8124), .ZN(n8258) );
  NAND2_X1 U8178 ( .A1(n8121), .A2(n8259), .ZN(n8124) );
  NAND2_X1 U8179 ( .A1(n8119), .A2(n8122), .ZN(n8259) );
  NAND2_X1 U8180 ( .A1(n8260), .A2(n8261), .ZN(n8122) );
  NAND2_X1 U8181 ( .A1(n8262), .A2(n8263), .ZN(n8261) );
  XNOR2_X1 U8182 ( .A(n8264), .B(n8265), .ZN(n8260) );
  NAND2_X1 U8183 ( .A1(n8116), .A2(n8266), .ZN(n8119) );
  NAND2_X1 U8184 ( .A1(n8114), .A2(n8117), .ZN(n8266) );
  NAND2_X1 U8185 ( .A1(n8267), .A2(n8268), .ZN(n8117) );
  NAND2_X1 U8186 ( .A1(n8269), .A2(n8270), .ZN(n8268) );
  XOR2_X1 U8187 ( .A(n8263), .B(n8271), .Z(n8267) );
  NAND2_X1 U8188 ( .A1(n8111), .A2(n8272), .ZN(n8114) );
  NAND2_X1 U8189 ( .A1(n8109), .A2(n8112), .ZN(n8272) );
  NAND2_X1 U8190 ( .A1(n8273), .A2(n8274), .ZN(n8112) );
  NAND2_X1 U8191 ( .A1(n8107), .A2(n8275), .ZN(n8109) );
  NAND2_X1 U8192 ( .A1(n8106), .A2(n8104), .ZN(n8275) );
  NAND2_X1 U8193 ( .A1(n8101), .A2(n8276), .ZN(n8104) );
  NAND2_X1 U8194 ( .A1(n8099), .A2(n8102), .ZN(n8276) );
  NAND2_X1 U8195 ( .A1(n8277), .A2(n8278), .ZN(n8102) );
  XNOR2_X1 U8196 ( .A(n8279), .B(n8280), .ZN(n8277) );
  NAND2_X1 U8197 ( .A1(n8096), .A2(n8281), .ZN(n8099) );
  NAND2_X1 U8198 ( .A1(n8094), .A2(n8097), .ZN(n8281) );
  NAND2_X1 U8199 ( .A1(n8282), .A2(n8283), .ZN(n8097) );
  NAND2_X1 U8200 ( .A1(n8284), .A2(n8278), .ZN(n8283) );
  INV_X1 U8201 ( .A(n8285), .ZN(n8278) );
  NAND2_X1 U8202 ( .A1(n8286), .A2(n8287), .ZN(n8284) );
  OR2_X1 U8203 ( .A1(n8288), .A2(n8289), .ZN(n8282) );
  NAND2_X1 U8204 ( .A1(n8092), .A2(n8290), .ZN(n8094) );
  NAND2_X1 U8205 ( .A1(n8089), .A2(n8091), .ZN(n8290) );
  NAND2_X1 U8206 ( .A1(n8291), .A2(n8292), .ZN(n8091) );
  NAND2_X1 U8207 ( .A1(n8293), .A2(n8294), .ZN(n8292) );
  XOR2_X1 U8208 ( .A(n8295), .B(n8288), .Z(n8291) );
  NAND2_X1 U8209 ( .A1(n8086), .A2(n8296), .ZN(n8089) );
  NAND2_X1 U8210 ( .A1(n8084), .A2(n8087), .ZN(n8296) );
  NAND2_X1 U8211 ( .A1(n8297), .A2(n8298), .ZN(n8087) );
  NAND2_X1 U8212 ( .A1(n8299), .A2(n8300), .ZN(n8298) );
  XOR2_X1 U8213 ( .A(n8294), .B(n8301), .Z(n8297) );
  INV_X1 U8214 ( .A(n8074), .ZN(n8084) );
  NAND2_X1 U8215 ( .A1(n8302), .A2(n8071), .ZN(n8074) );
  XOR2_X1 U8216 ( .A(n8303), .B(n8304), .Z(n8071) );
  XOR2_X1 U8217 ( .A(n8305), .B(n8306), .Z(n8303) );
  NOR2_X1 U8218 ( .A1(n8307), .A2(n7512), .ZN(n8306) );
  NOR2_X1 U8219 ( .A1(n8070), .A2(n8075), .ZN(n8302) );
  XNOR2_X1 U8220 ( .A(n8300), .B(n8299), .ZN(n8075) );
  INV_X1 U8221 ( .A(n8077), .ZN(n8070) );
  NAND2_X1 U8222 ( .A1(n8308), .A2(n8309), .ZN(n8077) );
  NAND2_X1 U8223 ( .A1(n8310), .A2(b_31_), .ZN(n8309) );
  NOR2_X1 U8224 ( .A1(n8311), .A2(n8307), .ZN(n8310) );
  NOR2_X1 U8225 ( .A1(n8065), .A2(n8067), .ZN(n8311) );
  NAND2_X1 U8226 ( .A1(n8065), .A2(n8067), .ZN(n8308) );
  NAND2_X1 U8227 ( .A1(n8312), .A2(n8313), .ZN(n8067) );
  NAND2_X1 U8228 ( .A1(n8314), .A2(b_31_), .ZN(n8313) );
  NOR2_X1 U8229 ( .A1(n8315), .A2(n7973), .ZN(n8314) );
  NOR2_X1 U8230 ( .A1(n7970), .A2(n7971), .ZN(n8315) );
  NAND2_X1 U8231 ( .A1(n7970), .A2(n7971), .ZN(n8312) );
  NAND2_X1 U8232 ( .A1(n8316), .A2(n8317), .ZN(n7971) );
  NAND2_X1 U8233 ( .A1(n8318), .A2(b_31_), .ZN(n8317) );
  NOR2_X1 U8234 ( .A1(n8319), .A2(n7965), .ZN(n8318) );
  NOR2_X1 U8235 ( .A1(n7962), .A2(n7963), .ZN(n8319) );
  NAND2_X1 U8236 ( .A1(n7962), .A2(n7963), .ZN(n8316) );
  NAND2_X1 U8237 ( .A1(n8320), .A2(n8321), .ZN(n7963) );
  NAND2_X1 U8238 ( .A1(n8322), .A2(b_31_), .ZN(n8321) );
  NOR2_X1 U8239 ( .A1(n8323), .A2(n7945), .ZN(n8322) );
  NOR2_X1 U8240 ( .A1(n7949), .A2(n7951), .ZN(n8323) );
  NAND2_X1 U8241 ( .A1(n7949), .A2(n7951), .ZN(n8320) );
  NAND2_X1 U8242 ( .A1(n8324), .A2(n8325), .ZN(n7951) );
  NAND2_X1 U8243 ( .A1(n8326), .A2(b_31_), .ZN(n8325) );
  NOR2_X1 U8244 ( .A1(n8327), .A2(n7934), .ZN(n8326) );
  NOR2_X1 U8245 ( .A1(n7931), .A2(n7932), .ZN(n8327) );
  NAND2_X1 U8246 ( .A1(n7931), .A2(n7932), .ZN(n8324) );
  NAND2_X1 U8247 ( .A1(n8328), .A2(n8329), .ZN(n7932) );
  NAND2_X1 U8248 ( .A1(n8330), .A2(b_31_), .ZN(n8329) );
  NOR2_X1 U8249 ( .A1(n8331), .A2(n7914), .ZN(n8330) );
  NOR2_X1 U8250 ( .A1(n7919), .A2(n7920), .ZN(n8331) );
  NAND2_X1 U8251 ( .A1(n7919), .A2(n7920), .ZN(n8328) );
  NAND2_X1 U8252 ( .A1(n8332), .A2(n8333), .ZN(n7920) );
  NAND2_X1 U8253 ( .A1(n8334), .A2(b_31_), .ZN(n8333) );
  NOR2_X1 U8254 ( .A1(n8335), .A2(n8061), .ZN(n8334) );
  NOR2_X1 U8255 ( .A1(n7900), .A2(n7902), .ZN(n8335) );
  NAND2_X1 U8256 ( .A1(n7900), .A2(n7902), .ZN(n8332) );
  NAND2_X1 U8257 ( .A1(n8336), .A2(n8337), .ZN(n7902) );
  NAND2_X1 U8258 ( .A1(n8338), .A2(b_31_), .ZN(n8337) );
  NOR2_X1 U8259 ( .A1(n8339), .A2(n7884), .ZN(n8338) );
  NOR2_X1 U8260 ( .A1(n7889), .A2(n7890), .ZN(n8339) );
  NAND2_X1 U8261 ( .A1(n7889), .A2(n7890), .ZN(n8336) );
  NAND2_X1 U8262 ( .A1(n8340), .A2(n8341), .ZN(n7890) );
  NAND2_X1 U8263 ( .A1(n8342), .A2(b_31_), .ZN(n8341) );
  NOR2_X1 U8264 ( .A1(n8343), .A2(n8059), .ZN(n8342) );
  NOR2_X1 U8265 ( .A1(n7865), .A2(n7867), .ZN(n8343) );
  NAND2_X1 U8266 ( .A1(n7865), .A2(n7867), .ZN(n8340) );
  NAND2_X1 U8267 ( .A1(n8344), .A2(n8345), .ZN(n7867) );
  NAND2_X1 U8268 ( .A1(n8346), .A2(b_31_), .ZN(n8345) );
  NOR2_X1 U8269 ( .A1(n8347), .A2(n7848), .ZN(n8346) );
  NOR2_X1 U8270 ( .A1(n7853), .A2(n7855), .ZN(n8347) );
  NAND2_X1 U8271 ( .A1(n7853), .A2(n7855), .ZN(n8344) );
  NAND2_X1 U8272 ( .A1(n8348), .A2(n8349), .ZN(n7855) );
  NAND2_X1 U8273 ( .A1(n8350), .A2(b_31_), .ZN(n8349) );
  NOR2_X1 U8274 ( .A1(n8351), .A2(n7837), .ZN(n8350) );
  NOR2_X1 U8275 ( .A1(n7834), .A2(n7835), .ZN(n8351) );
  NAND2_X1 U8276 ( .A1(n7834), .A2(n7835), .ZN(n8348) );
  NAND2_X1 U8277 ( .A1(n8352), .A2(n8353), .ZN(n7835) );
  NAND2_X1 U8278 ( .A1(n8354), .A2(b_31_), .ZN(n8353) );
  NOR2_X1 U8279 ( .A1(n8355), .A2(n7817), .ZN(n8354) );
  NOR2_X1 U8280 ( .A1(n7822), .A2(n7823), .ZN(n8355) );
  NAND2_X1 U8281 ( .A1(n7822), .A2(n7823), .ZN(n8352) );
  NAND2_X1 U8282 ( .A1(n8356), .A2(n8357), .ZN(n7823) );
  NAND2_X1 U8283 ( .A1(n8358), .A2(b_31_), .ZN(n8357) );
  NOR2_X1 U8284 ( .A1(n8359), .A2(n7806), .ZN(n8358) );
  NOR2_X1 U8285 ( .A1(n7803), .A2(n7804), .ZN(n8359) );
  NAND2_X1 U8286 ( .A1(n7803), .A2(n7804), .ZN(n8356) );
  NAND2_X1 U8287 ( .A1(n8360), .A2(n8361), .ZN(n7804) );
  NAND2_X1 U8288 ( .A1(n8362), .A2(b_31_), .ZN(n8361) );
  NOR2_X1 U8289 ( .A1(n8363), .A2(n7786), .ZN(n8362) );
  NOR2_X1 U8290 ( .A1(n7790), .A2(n7792), .ZN(n8363) );
  NAND2_X1 U8291 ( .A1(n7790), .A2(n7792), .ZN(n8360) );
  NAND2_X1 U8292 ( .A1(n8364), .A2(n8365), .ZN(n7792) );
  NAND2_X1 U8293 ( .A1(n8366), .A2(b_31_), .ZN(n8365) );
  NOR2_X1 U8294 ( .A1(n8367), .A2(n7775), .ZN(n8366) );
  NOR2_X1 U8295 ( .A1(n7772), .A2(n7773), .ZN(n8367) );
  NAND2_X1 U8296 ( .A1(n7772), .A2(n7773), .ZN(n8364) );
  NAND2_X1 U8297 ( .A1(n8368), .A2(n8369), .ZN(n7773) );
  NAND2_X1 U8298 ( .A1(n8370), .A2(b_31_), .ZN(n8369) );
  NOR2_X1 U8299 ( .A1(n8371), .A2(n7754), .ZN(n8370) );
  NOR2_X1 U8300 ( .A1(n7759), .A2(n7761), .ZN(n8371) );
  NAND2_X1 U8301 ( .A1(n7759), .A2(n7761), .ZN(n8368) );
  NAND2_X1 U8302 ( .A1(n8372), .A2(n8373), .ZN(n7761) );
  NAND2_X1 U8303 ( .A1(n8374), .A2(b_31_), .ZN(n8373) );
  NOR2_X1 U8304 ( .A1(n8375), .A2(n7743), .ZN(n8374) );
  NOR2_X1 U8305 ( .A1(n7740), .A2(n7741), .ZN(n8375) );
  NAND2_X1 U8306 ( .A1(n7740), .A2(n7741), .ZN(n8372) );
  NAND2_X1 U8307 ( .A1(n8376), .A2(n8377), .ZN(n7741) );
  NAND2_X1 U8308 ( .A1(n8378), .A2(b_31_), .ZN(n8377) );
  NOR2_X1 U8309 ( .A1(n8379), .A2(n7723), .ZN(n8378) );
  NOR2_X1 U8310 ( .A1(n7727), .A2(n7729), .ZN(n8379) );
  NAND2_X1 U8311 ( .A1(n7727), .A2(n7729), .ZN(n8376) );
  NAND2_X1 U8312 ( .A1(n8380), .A2(n8381), .ZN(n7729) );
  NAND2_X1 U8313 ( .A1(n8382), .A2(b_31_), .ZN(n8381) );
  NOR2_X1 U8314 ( .A1(n8383), .A2(n7707), .ZN(n8382) );
  NOR2_X1 U8315 ( .A1(n7704), .A2(n7705), .ZN(n8383) );
  NAND2_X1 U8316 ( .A1(n7704), .A2(n7705), .ZN(n8380) );
  NAND2_X1 U8317 ( .A1(n8384), .A2(n8385), .ZN(n7705) );
  NAND2_X1 U8318 ( .A1(n8386), .A2(b_31_), .ZN(n8385) );
  NOR2_X1 U8319 ( .A1(n8387), .A2(n7687), .ZN(n8386) );
  NOR2_X1 U8320 ( .A1(n7691), .A2(n7693), .ZN(n8387) );
  NAND2_X1 U8321 ( .A1(n7691), .A2(n7693), .ZN(n8384) );
  NAND2_X1 U8322 ( .A1(n8388), .A2(n8389), .ZN(n7693) );
  NAND2_X1 U8323 ( .A1(n8390), .A2(b_31_), .ZN(n8389) );
  NOR2_X1 U8324 ( .A1(n8391), .A2(n7676), .ZN(n8390) );
  NOR2_X1 U8325 ( .A1(n7673), .A2(n7674), .ZN(n8391) );
  NAND2_X1 U8326 ( .A1(n7673), .A2(n7674), .ZN(n8388) );
  NAND2_X1 U8327 ( .A1(n7662), .A2(n8392), .ZN(n7674) );
  NAND2_X1 U8328 ( .A1(n7661), .A2(n7663), .ZN(n8392) );
  NAND2_X1 U8329 ( .A1(n8393), .A2(n8394), .ZN(n7663) );
  NAND2_X1 U8330 ( .A1(b_31_), .A2(a_21_), .ZN(n8394) );
  INV_X1 U8331 ( .A(n8395), .ZN(n8393) );
  XOR2_X1 U8332 ( .A(n8396), .B(n8397), .Z(n7661) );
  XOR2_X1 U8333 ( .A(n8398), .B(n8399), .Z(n8396) );
  NOR2_X1 U8334 ( .A1(n7645), .A2(n7512), .ZN(n8399) );
  NAND2_X1 U8335 ( .A1(a_21_), .A2(n8395), .ZN(n7662) );
  NAND2_X1 U8336 ( .A1(n8400), .A2(n8401), .ZN(n8395) );
  NAND2_X1 U8337 ( .A1(n8402), .A2(b_31_), .ZN(n8401) );
  NOR2_X1 U8338 ( .A1(n8403), .A2(n7645), .ZN(n8402) );
  NOR2_X1 U8339 ( .A1(n7642), .A2(n7643), .ZN(n8403) );
  NAND2_X1 U8340 ( .A1(n7642), .A2(n7643), .ZN(n8400) );
  NAND2_X1 U8341 ( .A1(n7631), .A2(n8404), .ZN(n7643) );
  NAND2_X1 U8342 ( .A1(n7630), .A2(n7632), .ZN(n8404) );
  NAND2_X1 U8343 ( .A1(n8405), .A2(n8406), .ZN(n7632) );
  NAND2_X1 U8344 ( .A1(b_31_), .A2(a_23_), .ZN(n8406) );
  INV_X1 U8345 ( .A(n8407), .ZN(n8405) );
  XOR2_X1 U8346 ( .A(n8408), .B(n8409), .Z(n7630) );
  XOR2_X1 U8347 ( .A(n8410), .B(n8411), .Z(n8408) );
  NOR2_X1 U8348 ( .A1(n7613), .A2(n7512), .ZN(n8411) );
  NAND2_X1 U8349 ( .A1(a_23_), .A2(n8407), .ZN(n7631) );
  NAND2_X1 U8350 ( .A1(n8412), .A2(n8413), .ZN(n8407) );
  NAND2_X1 U8351 ( .A1(n8414), .A2(b_31_), .ZN(n8413) );
  NOR2_X1 U8352 ( .A1(n8415), .A2(n7613), .ZN(n8414) );
  NOR2_X1 U8353 ( .A1(n7610), .A2(n7611), .ZN(n8415) );
  NAND2_X1 U8354 ( .A1(n7610), .A2(n7611), .ZN(n8412) );
  NAND2_X1 U8355 ( .A1(n7599), .A2(n8416), .ZN(n7611) );
  NAND2_X1 U8356 ( .A1(n7598), .A2(n7600), .ZN(n8416) );
  NAND2_X1 U8357 ( .A1(n8417), .A2(n8418), .ZN(n7600) );
  NAND2_X1 U8358 ( .A1(b_31_), .A2(a_25_), .ZN(n8418) );
  INV_X1 U8359 ( .A(n8419), .ZN(n8417) );
  XNOR2_X1 U8360 ( .A(n8420), .B(n8421), .ZN(n7598) );
  XOR2_X1 U8361 ( .A(n8422), .B(n8423), .Z(n8421) );
  NAND2_X1 U8362 ( .A1(b_30_), .A2(a_26_), .ZN(n8423) );
  NAND2_X1 U8363 ( .A1(a_25_), .A2(n8419), .ZN(n7599) );
  NAND2_X1 U8364 ( .A1(n7581), .A2(n8424), .ZN(n8419) );
  NAND2_X1 U8365 ( .A1(n7580), .A2(n7582), .ZN(n8424) );
  NAND2_X1 U8366 ( .A1(n8425), .A2(n8426), .ZN(n7582) );
  NAND2_X1 U8367 ( .A1(b_31_), .A2(a_26_), .ZN(n8426) );
  INV_X1 U8368 ( .A(n8427), .ZN(n8425) );
  XNOR2_X1 U8369 ( .A(n8428), .B(n8429), .ZN(n7580) );
  XNOR2_X1 U8370 ( .A(n8430), .B(n8431), .ZN(n8429) );
  NAND2_X1 U8371 ( .A1(a_26_), .A2(n8427), .ZN(n7581) );
  NAND2_X1 U8372 ( .A1(n8432), .A2(n8433), .ZN(n8427) );
  NAND2_X1 U8373 ( .A1(n8434), .A2(b_31_), .ZN(n8433) );
  NOR2_X1 U8374 ( .A1(n8435), .A2(n7563), .ZN(n8434) );
  NOR2_X1 U8375 ( .A1(n7567), .A2(n7569), .ZN(n8435) );
  NAND2_X1 U8376 ( .A1(n7567), .A2(n7569), .ZN(n8432) );
  NAND2_X1 U8377 ( .A1(n8436), .A2(n8437), .ZN(n7569) );
  NAND2_X1 U8378 ( .A1(n8438), .A2(b_31_), .ZN(n8437) );
  NOR2_X1 U8379 ( .A1(n8439), .A2(n7547), .ZN(n8438) );
  NOR2_X1 U8380 ( .A1(n7543), .A2(n7545), .ZN(n8439) );
  NAND2_X1 U8381 ( .A1(n7543), .A2(n7545), .ZN(n8436) );
  NAND2_X1 U8382 ( .A1(n8440), .A2(n8441), .ZN(n7545) );
  NAND2_X1 U8383 ( .A1(n8442), .A2(b_31_), .ZN(n8441) );
  NOR2_X1 U8384 ( .A1(n8443), .A2(n7529), .ZN(n8442) );
  NOR2_X1 U8385 ( .A1(n7533), .A2(n7534), .ZN(n8443) );
  NAND2_X1 U8386 ( .A1(n7533), .A2(n7534), .ZN(n8440) );
  NAND2_X1 U8387 ( .A1(n8444), .A2(n8445), .ZN(n7534) );
  NAND2_X1 U8388 ( .A1(b_29_), .A2(n8446), .ZN(n8445) );
  NAND2_X1 U8389 ( .A1(n7506), .A2(n8447), .ZN(n8446) );
  NAND2_X1 U8390 ( .A1(a_31_), .A2(n7512), .ZN(n8447) );
  NAND2_X1 U8391 ( .A1(b_30_), .A2(n8448), .ZN(n8444) );
  NAND2_X1 U8392 ( .A1(n7510), .A2(n8449), .ZN(n8448) );
  NAND2_X1 U8393 ( .A1(a_30_), .A2(n7527), .ZN(n8449) );
  AND2_X1 U8394 ( .A1(n8450), .A2(b_31_), .ZN(n7533) );
  NOR2_X1 U8395 ( .A1(n8451), .A2(n7512), .ZN(n8450) );
  XOR2_X1 U8396 ( .A(n8452), .B(n8453), .Z(n7543) );
  NOR2_X1 U8397 ( .A1(n7529), .A2(n7512), .ZN(n8453) );
  XOR2_X1 U8398 ( .A(n8454), .B(n8455), .Z(n8452) );
  XNOR2_X1 U8399 ( .A(n8456), .B(n8457), .ZN(n7567) );
  NAND2_X1 U8400 ( .A1(n8458), .A2(n8459), .ZN(n8456) );
  XNOR2_X1 U8401 ( .A(n8460), .B(n8461), .ZN(n7610) );
  XNOR2_X1 U8402 ( .A(n8462), .B(n8463), .ZN(n8461) );
  XNOR2_X1 U8403 ( .A(n8464), .B(n8465), .ZN(n7642) );
  XNOR2_X1 U8404 ( .A(n8466), .B(n8467), .ZN(n8465) );
  XNOR2_X1 U8405 ( .A(n8468), .B(n8469), .ZN(n7673) );
  XNOR2_X1 U8406 ( .A(n8470), .B(n8471), .ZN(n8468) );
  XOR2_X1 U8407 ( .A(n8472), .B(n8473), .Z(n7691) );
  XOR2_X1 U8408 ( .A(n8474), .B(n8475), .Z(n8472) );
  NOR2_X1 U8409 ( .A1(n7676), .A2(n7512), .ZN(n8475) );
  XNOR2_X1 U8410 ( .A(n8476), .B(n8477), .ZN(n7704) );
  XNOR2_X1 U8411 ( .A(n8478), .B(n8479), .ZN(n8476) );
  XOR2_X1 U8412 ( .A(n8480), .B(n8481), .Z(n7727) );
  XOR2_X1 U8413 ( .A(n8482), .B(n8483), .Z(n8480) );
  NOR2_X1 U8414 ( .A1(n7707), .A2(n7512), .ZN(n8483) );
  XNOR2_X1 U8415 ( .A(n8484), .B(n8485), .ZN(n7740) );
  XNOR2_X1 U8416 ( .A(n8486), .B(n8487), .ZN(n8484) );
  XNOR2_X1 U8417 ( .A(n8488), .B(n8489), .ZN(n7759) );
  XOR2_X1 U8418 ( .A(n8490), .B(n8491), .Z(n8489) );
  NAND2_X1 U8419 ( .A1(b_30_), .A2(a_16_), .ZN(n8491) );
  XNOR2_X1 U8420 ( .A(n8492), .B(n8493), .ZN(n7772) );
  XNOR2_X1 U8421 ( .A(n8494), .B(n8495), .ZN(n8492) );
  XOR2_X1 U8422 ( .A(n8496), .B(n8497), .Z(n7790) );
  XOR2_X1 U8423 ( .A(n8498), .B(n8499), .Z(n8496) );
  NOR2_X1 U8424 ( .A1(n7775), .A2(n7512), .ZN(n8499) );
  XNOR2_X1 U8425 ( .A(n8500), .B(n8501), .ZN(n7803) );
  XNOR2_X1 U8426 ( .A(n8502), .B(n8503), .ZN(n8500) );
  XOR2_X1 U8427 ( .A(n8504), .B(n8505), .Z(n7822) );
  XOR2_X1 U8428 ( .A(n8506), .B(n8507), .Z(n8504) );
  NOR2_X1 U8429 ( .A1(n7806), .A2(n7512), .ZN(n8507) );
  XNOR2_X1 U8430 ( .A(n8508), .B(n8509), .ZN(n7834) );
  XNOR2_X1 U8431 ( .A(n8510), .B(n8511), .ZN(n8508) );
  XOR2_X1 U8432 ( .A(n8512), .B(n8513), .Z(n7853) );
  XOR2_X1 U8433 ( .A(n8514), .B(n8515), .Z(n8512) );
  NOR2_X1 U8434 ( .A1(n7837), .A2(n7512), .ZN(n8515) );
  XOR2_X1 U8435 ( .A(n8516), .B(n8517), .Z(n7865) );
  XOR2_X1 U8436 ( .A(n8518), .B(n8519), .Z(n8516) );
  XOR2_X1 U8437 ( .A(n8520), .B(n8521), .Z(n7889) );
  XOR2_X1 U8438 ( .A(n8522), .B(n8523), .Z(n8520) );
  NOR2_X1 U8439 ( .A1(n8059), .A2(n7512), .ZN(n8523) );
  XOR2_X1 U8440 ( .A(n8524), .B(n8525), .Z(n7900) );
  XOR2_X1 U8441 ( .A(n8526), .B(n8527), .Z(n8524) );
  XOR2_X1 U8442 ( .A(n8528), .B(n8529), .Z(n7919) );
  XOR2_X1 U8443 ( .A(n8530), .B(n8531), .Z(n8528) );
  NOR2_X1 U8444 ( .A1(n8061), .A2(n7512), .ZN(n8531) );
  XNOR2_X1 U8445 ( .A(n8532), .B(n8533), .ZN(n7931) );
  XNOR2_X1 U8446 ( .A(n8534), .B(n8535), .ZN(n8532) );
  XOR2_X1 U8447 ( .A(n8536), .B(n8537), .Z(n7949) );
  XOR2_X1 U8448 ( .A(n8538), .B(n8539), .Z(n8536) );
  NOR2_X1 U8449 ( .A1(n7934), .A2(n7512), .ZN(n8539) );
  XNOR2_X1 U8450 ( .A(n8540), .B(n8541), .ZN(n7962) );
  XNOR2_X1 U8451 ( .A(n8542), .B(n8543), .ZN(n8540) );
  XOR2_X1 U8452 ( .A(n8544), .B(n8545), .Z(n7970) );
  XOR2_X1 U8453 ( .A(n8546), .B(n8547), .Z(n8544) );
  NOR2_X1 U8454 ( .A1(n7965), .A2(n7512), .ZN(n8547) );
  XNOR2_X1 U8455 ( .A(n8548), .B(n8549), .ZN(n8065) );
  NAND2_X1 U8456 ( .A1(n8550), .A2(n8551), .ZN(n8548) );
  NAND2_X1 U8457 ( .A1(n8552), .A2(n8553), .ZN(n8086) );
  XOR2_X1 U8458 ( .A(n8294), .B(n8293), .Z(n8553) );
  AND2_X1 U8459 ( .A1(n8300), .A2(n8299), .ZN(n8552) );
  XNOR2_X1 U8460 ( .A(n8554), .B(n8555), .ZN(n8299) );
  NAND2_X1 U8461 ( .A1(n8556), .A2(n8557), .ZN(n8554) );
  NAND2_X1 U8462 ( .A1(n8558), .A2(n8559), .ZN(n8300) );
  NAND2_X1 U8463 ( .A1(n8560), .A2(b_30_), .ZN(n8559) );
  NOR2_X1 U8464 ( .A1(n8561), .A2(n8307), .ZN(n8560) );
  NOR2_X1 U8465 ( .A1(n8304), .A2(n8305), .ZN(n8561) );
  NAND2_X1 U8466 ( .A1(n8304), .A2(n8305), .ZN(n8558) );
  NAND2_X1 U8467 ( .A1(n8550), .A2(n8562), .ZN(n8305) );
  NAND2_X1 U8468 ( .A1(n8549), .A2(n8551), .ZN(n8562) );
  NAND2_X1 U8469 ( .A1(n8563), .A2(n8564), .ZN(n8551) );
  NAND2_X1 U8470 ( .A1(b_30_), .A2(a_1_), .ZN(n8564) );
  INV_X1 U8471 ( .A(n8565), .ZN(n8563) );
  XOR2_X1 U8472 ( .A(n8566), .B(n8567), .Z(n8549) );
  XOR2_X1 U8473 ( .A(n8568), .B(n8569), .Z(n8566) );
  NAND2_X1 U8474 ( .A1(a_1_), .A2(n8565), .ZN(n8550) );
  NAND2_X1 U8475 ( .A1(n8570), .A2(n8571), .ZN(n8565) );
  NAND2_X1 U8476 ( .A1(n8572), .A2(b_30_), .ZN(n8571) );
  NOR2_X1 U8477 ( .A1(n8573), .A2(n7965), .ZN(n8572) );
  NOR2_X1 U8478 ( .A1(n8545), .A2(n8546), .ZN(n8573) );
  NAND2_X1 U8479 ( .A1(n8545), .A2(n8546), .ZN(n8570) );
  NAND2_X1 U8480 ( .A1(n8574), .A2(n8575), .ZN(n8546) );
  NAND2_X1 U8481 ( .A1(n8543), .A2(n8576), .ZN(n8575) );
  NAND2_X1 U8482 ( .A1(n8542), .A2(n8541), .ZN(n8576) );
  NOR2_X1 U8483 ( .A1(n7512), .A2(n7945), .ZN(n8543) );
  OR2_X1 U8484 ( .A1(n8541), .A2(n8542), .ZN(n8574) );
  AND2_X1 U8485 ( .A1(n8577), .A2(n8578), .ZN(n8542) );
  NAND2_X1 U8486 ( .A1(n8579), .A2(b_30_), .ZN(n8578) );
  NOR2_X1 U8487 ( .A1(n8580), .A2(n7934), .ZN(n8579) );
  NOR2_X1 U8488 ( .A1(n8538), .A2(n8537), .ZN(n8580) );
  NAND2_X1 U8489 ( .A1(n8537), .A2(n8538), .ZN(n8577) );
  NAND2_X1 U8490 ( .A1(n8581), .A2(n8582), .ZN(n8538) );
  NAND2_X1 U8491 ( .A1(n8535), .A2(n8583), .ZN(n8582) );
  NAND2_X1 U8492 ( .A1(n8534), .A2(n8533), .ZN(n8583) );
  NOR2_X1 U8493 ( .A1(n7512), .A2(n7914), .ZN(n8535) );
  OR2_X1 U8494 ( .A1(n8533), .A2(n8534), .ZN(n8581) );
  AND2_X1 U8495 ( .A1(n8584), .A2(n8585), .ZN(n8534) );
  NAND2_X1 U8496 ( .A1(n8586), .A2(b_30_), .ZN(n8585) );
  NOR2_X1 U8497 ( .A1(n8587), .A2(n8061), .ZN(n8586) );
  NOR2_X1 U8498 ( .A1(n8529), .A2(n8530), .ZN(n8587) );
  NAND2_X1 U8499 ( .A1(n8529), .A2(n8530), .ZN(n8584) );
  NAND2_X1 U8500 ( .A1(n8588), .A2(n8589), .ZN(n8530) );
  NAND2_X1 U8501 ( .A1(n8527), .A2(n8590), .ZN(n8589) );
  OR2_X1 U8502 ( .A1(n8525), .A2(n8526), .ZN(n8590) );
  NOR2_X1 U8503 ( .A1(n7512), .A2(n7884), .ZN(n8527) );
  NAND2_X1 U8504 ( .A1(n8525), .A2(n8526), .ZN(n8588) );
  NAND2_X1 U8505 ( .A1(n8591), .A2(n8592), .ZN(n8526) );
  NAND2_X1 U8506 ( .A1(n8593), .A2(b_30_), .ZN(n8592) );
  NOR2_X1 U8507 ( .A1(n8594), .A2(n8059), .ZN(n8593) );
  NOR2_X1 U8508 ( .A1(n8521), .A2(n8522), .ZN(n8594) );
  NAND2_X1 U8509 ( .A1(n8521), .A2(n8522), .ZN(n8591) );
  NAND2_X1 U8510 ( .A1(n8595), .A2(n8596), .ZN(n8522) );
  NAND2_X1 U8511 ( .A1(n8519), .A2(n8597), .ZN(n8596) );
  OR2_X1 U8512 ( .A1(n8517), .A2(n8518), .ZN(n8597) );
  NOR2_X1 U8513 ( .A1(n7512), .A2(n7848), .ZN(n8519) );
  NAND2_X1 U8514 ( .A1(n8517), .A2(n8518), .ZN(n8595) );
  NAND2_X1 U8515 ( .A1(n8598), .A2(n8599), .ZN(n8518) );
  NAND2_X1 U8516 ( .A1(n8600), .A2(b_30_), .ZN(n8599) );
  NOR2_X1 U8517 ( .A1(n8601), .A2(n7837), .ZN(n8600) );
  NOR2_X1 U8518 ( .A1(n8514), .A2(n8513), .ZN(n8601) );
  NAND2_X1 U8519 ( .A1(n8513), .A2(n8514), .ZN(n8598) );
  NAND2_X1 U8520 ( .A1(n8602), .A2(n8603), .ZN(n8514) );
  NAND2_X1 U8521 ( .A1(n8511), .A2(n8604), .ZN(n8603) );
  NAND2_X1 U8522 ( .A1(n8510), .A2(n8509), .ZN(n8604) );
  NOR2_X1 U8523 ( .A1(n7512), .A2(n7817), .ZN(n8511) );
  OR2_X1 U8524 ( .A1(n8509), .A2(n8510), .ZN(n8602) );
  AND2_X1 U8525 ( .A1(n8605), .A2(n8606), .ZN(n8510) );
  NAND2_X1 U8526 ( .A1(n8607), .A2(b_30_), .ZN(n8606) );
  NOR2_X1 U8527 ( .A1(n8608), .A2(n7806), .ZN(n8607) );
  NOR2_X1 U8528 ( .A1(n8505), .A2(n8506), .ZN(n8608) );
  NAND2_X1 U8529 ( .A1(n8505), .A2(n8506), .ZN(n8605) );
  NAND2_X1 U8530 ( .A1(n8609), .A2(n8610), .ZN(n8506) );
  NAND2_X1 U8531 ( .A1(n8503), .A2(n8611), .ZN(n8610) );
  NAND2_X1 U8532 ( .A1(n8502), .A2(n8501), .ZN(n8611) );
  NOR2_X1 U8533 ( .A1(n7512), .A2(n7786), .ZN(n8503) );
  OR2_X1 U8534 ( .A1(n8501), .A2(n8502), .ZN(n8609) );
  AND2_X1 U8535 ( .A1(n8612), .A2(n8613), .ZN(n8502) );
  NAND2_X1 U8536 ( .A1(n8614), .A2(b_30_), .ZN(n8613) );
  NOR2_X1 U8537 ( .A1(n8615), .A2(n7775), .ZN(n8614) );
  NOR2_X1 U8538 ( .A1(n8498), .A2(n8497), .ZN(n8615) );
  NAND2_X1 U8539 ( .A1(n8497), .A2(n8498), .ZN(n8612) );
  NAND2_X1 U8540 ( .A1(n8616), .A2(n8617), .ZN(n8498) );
  NAND2_X1 U8541 ( .A1(n8494), .A2(n8618), .ZN(n8617) );
  NAND2_X1 U8542 ( .A1(n8495), .A2(n8493), .ZN(n8618) );
  NOR2_X1 U8543 ( .A1(n7512), .A2(n7754), .ZN(n8494) );
  OR2_X1 U8544 ( .A1(n8493), .A2(n8495), .ZN(n8616) );
  AND2_X1 U8545 ( .A1(n8619), .A2(n8620), .ZN(n8495) );
  NAND2_X1 U8546 ( .A1(n8621), .A2(b_30_), .ZN(n8620) );
  NOR2_X1 U8547 ( .A1(n8622), .A2(n7743), .ZN(n8621) );
  NOR2_X1 U8548 ( .A1(n8490), .A2(n8488), .ZN(n8622) );
  NAND2_X1 U8549 ( .A1(n8488), .A2(n8490), .ZN(n8619) );
  NAND2_X1 U8550 ( .A1(n8623), .A2(n8624), .ZN(n8490) );
  NAND2_X1 U8551 ( .A1(n8487), .A2(n8625), .ZN(n8624) );
  NAND2_X1 U8552 ( .A1(n8486), .A2(n8485), .ZN(n8625) );
  NOR2_X1 U8553 ( .A1(n7512), .A2(n7723), .ZN(n8487) );
  OR2_X1 U8554 ( .A1(n8485), .A2(n8486), .ZN(n8623) );
  AND2_X1 U8555 ( .A1(n8626), .A2(n8627), .ZN(n8486) );
  NAND2_X1 U8556 ( .A1(n8628), .A2(b_30_), .ZN(n8627) );
  NOR2_X1 U8557 ( .A1(n8629), .A2(n7707), .ZN(n8628) );
  NOR2_X1 U8558 ( .A1(n8482), .A2(n8481), .ZN(n8629) );
  NAND2_X1 U8559 ( .A1(n8481), .A2(n8482), .ZN(n8626) );
  NAND2_X1 U8560 ( .A1(n8630), .A2(n8631), .ZN(n8482) );
  NAND2_X1 U8561 ( .A1(n8479), .A2(n8632), .ZN(n8631) );
  NAND2_X1 U8562 ( .A1(n8478), .A2(n8477), .ZN(n8632) );
  NOR2_X1 U8563 ( .A1(n7512), .A2(n7687), .ZN(n8479) );
  OR2_X1 U8564 ( .A1(n8477), .A2(n8478), .ZN(n8630) );
  AND2_X1 U8565 ( .A1(n8633), .A2(n8634), .ZN(n8478) );
  NAND2_X1 U8566 ( .A1(n8635), .A2(b_30_), .ZN(n8634) );
  NOR2_X1 U8567 ( .A1(n8636), .A2(n7676), .ZN(n8635) );
  NOR2_X1 U8568 ( .A1(n8474), .A2(n8473), .ZN(n8636) );
  NAND2_X1 U8569 ( .A1(n8473), .A2(n8474), .ZN(n8633) );
  NAND2_X1 U8570 ( .A1(n8637), .A2(n8638), .ZN(n8474) );
  NAND2_X1 U8571 ( .A1(n8471), .A2(n8639), .ZN(n8638) );
  NAND2_X1 U8572 ( .A1(n8470), .A2(n8469), .ZN(n8639) );
  NOR2_X1 U8573 ( .A1(n7512), .A2(n7656), .ZN(n8471) );
  OR2_X1 U8574 ( .A1(n8469), .A2(n8470), .ZN(n8637) );
  AND2_X1 U8575 ( .A1(n8640), .A2(n8641), .ZN(n8470) );
  NAND2_X1 U8576 ( .A1(n8642), .A2(b_30_), .ZN(n8641) );
  NOR2_X1 U8577 ( .A1(n8643), .A2(n7645), .ZN(n8642) );
  NOR2_X1 U8578 ( .A1(n8398), .A2(n8397), .ZN(n8643) );
  NAND2_X1 U8579 ( .A1(n8397), .A2(n8398), .ZN(n8640) );
  NAND2_X1 U8580 ( .A1(n8644), .A2(n8645), .ZN(n8398) );
  NAND2_X1 U8581 ( .A1(n8467), .A2(n8646), .ZN(n8645) );
  OR2_X1 U8582 ( .A1(n8466), .A2(n8464), .ZN(n8646) );
  NOR2_X1 U8583 ( .A1(n7512), .A2(n7624), .ZN(n8467) );
  NAND2_X1 U8584 ( .A1(n8464), .A2(n8466), .ZN(n8644) );
  NAND2_X1 U8585 ( .A1(n8647), .A2(n8648), .ZN(n8466) );
  NAND2_X1 U8586 ( .A1(n8649), .A2(b_30_), .ZN(n8648) );
  NOR2_X1 U8587 ( .A1(n8650), .A2(n7613), .ZN(n8649) );
  NOR2_X1 U8588 ( .A1(n8410), .A2(n8409), .ZN(n8650) );
  NAND2_X1 U8589 ( .A1(n8409), .A2(n8410), .ZN(n8647) );
  NAND2_X1 U8590 ( .A1(n8651), .A2(n8652), .ZN(n8410) );
  NAND2_X1 U8591 ( .A1(n8463), .A2(n8653), .ZN(n8652) );
  OR2_X1 U8592 ( .A1(n8462), .A2(n8460), .ZN(n8653) );
  NOR2_X1 U8593 ( .A1(n7512), .A2(n7593), .ZN(n8463) );
  NAND2_X1 U8594 ( .A1(n8460), .A2(n8462), .ZN(n8651) );
  NAND2_X1 U8595 ( .A1(n8654), .A2(n8655), .ZN(n8462) );
  NAND2_X1 U8596 ( .A1(n8656), .A2(b_30_), .ZN(n8655) );
  NOR2_X1 U8597 ( .A1(n8657), .A2(n8052), .ZN(n8656) );
  NOR2_X1 U8598 ( .A1(n8420), .A2(n8422), .ZN(n8657) );
  NAND2_X1 U8599 ( .A1(n8420), .A2(n8422), .ZN(n8654) );
  NAND2_X1 U8600 ( .A1(n8658), .A2(n8659), .ZN(n8422) );
  NAND2_X1 U8601 ( .A1(n8431), .A2(n8660), .ZN(n8659) );
  OR2_X1 U8602 ( .A1(n8430), .A2(n8428), .ZN(n8660) );
  NOR2_X1 U8603 ( .A1(n7512), .A2(n7563), .ZN(n8431) );
  NAND2_X1 U8604 ( .A1(n8428), .A2(n8430), .ZN(n8658) );
  NAND2_X1 U8605 ( .A1(n8458), .A2(n8661), .ZN(n8430) );
  NAND2_X1 U8606 ( .A1(n8457), .A2(n8459), .ZN(n8661) );
  NAND2_X1 U8607 ( .A1(n8662), .A2(n8663), .ZN(n8459) );
  NAND2_X1 U8608 ( .A1(b_30_), .A2(a_28_), .ZN(n8663) );
  INV_X1 U8609 ( .A(n8664), .ZN(n8662) );
  XOR2_X1 U8610 ( .A(n8665), .B(n8666), .Z(n8457) );
  XOR2_X1 U8611 ( .A(n8042), .B(n8667), .Z(n8665) );
  NAND2_X1 U8612 ( .A1(a_28_), .A2(n8664), .ZN(n8458) );
  NAND2_X1 U8613 ( .A1(n8668), .A2(n8669), .ZN(n8664) );
  NAND2_X1 U8614 ( .A1(n8670), .A2(b_30_), .ZN(n8669) );
  NOR2_X1 U8615 ( .A1(n8671), .A2(n7529), .ZN(n8670) );
  NOR2_X1 U8616 ( .A1(n8454), .A2(n8455), .ZN(n8671) );
  NAND2_X1 U8617 ( .A1(n8454), .A2(n8455), .ZN(n8668) );
  NAND2_X1 U8618 ( .A1(n8672), .A2(n8673), .ZN(n8455) );
  NAND2_X1 U8619 ( .A1(n8674), .A2(b_28_), .ZN(n8673) );
  NOR2_X1 U8620 ( .A1(n8675), .A2(n8048), .ZN(n8674) );
  NOR2_X1 U8621 ( .A1(n8676), .A2(n7527), .ZN(n8675) );
  NAND2_X1 U8622 ( .A1(n8677), .A2(b_29_), .ZN(n8672) );
  NOR2_X1 U8623 ( .A1(n8678), .A2(n7515), .ZN(n8677) );
  NOR2_X1 U8624 ( .A1(n8679), .A2(n8050), .ZN(n8678) );
  AND2_X1 U8625 ( .A1(n8680), .A2(b_30_), .ZN(n8454) );
  NOR2_X1 U8626 ( .A1(n8451), .A2(n7527), .ZN(n8680) );
  XNOR2_X1 U8627 ( .A(n8681), .B(n8682), .ZN(n8428) );
  NAND2_X1 U8628 ( .A1(n8683), .A2(n8684), .ZN(n8681) );
  XNOR2_X1 U8629 ( .A(n8685), .B(n8686), .ZN(n8420) );
  XNOR2_X1 U8630 ( .A(n8687), .B(n8688), .ZN(n8686) );
  XNOR2_X1 U8631 ( .A(n8689), .B(n8690), .ZN(n8460) );
  XOR2_X1 U8632 ( .A(n8691), .B(n8692), .Z(n8690) );
  NAND2_X1 U8633 ( .A1(b_29_), .A2(a_26_), .ZN(n8692) );
  XNOR2_X1 U8634 ( .A(n8693), .B(n8694), .ZN(n8409) );
  XNOR2_X1 U8635 ( .A(n8695), .B(n8696), .ZN(n8694) );
  XNOR2_X1 U8636 ( .A(n8697), .B(n8698), .ZN(n8464) );
  XOR2_X1 U8637 ( .A(n8699), .B(n8700), .Z(n8698) );
  NAND2_X1 U8638 ( .A1(b_29_), .A2(a_24_), .ZN(n8700) );
  XNOR2_X1 U8639 ( .A(n8701), .B(n8702), .ZN(n8397) );
  XNOR2_X1 U8640 ( .A(n8703), .B(n8704), .ZN(n8701) );
  XNOR2_X1 U8641 ( .A(n8705), .B(n8706), .ZN(n8469) );
  XOR2_X1 U8642 ( .A(n8707), .B(n8708), .Z(n8705) );
  NOR2_X1 U8643 ( .A1(n7645), .A2(n7527), .ZN(n8708) );
  XNOR2_X1 U8644 ( .A(n8709), .B(n8710), .ZN(n8473) );
  XNOR2_X1 U8645 ( .A(n8711), .B(n8712), .ZN(n8709) );
  XNOR2_X1 U8646 ( .A(n8713), .B(n8714), .ZN(n8477) );
  XOR2_X1 U8647 ( .A(n8715), .B(n8716), .Z(n8713) );
  NOR2_X1 U8648 ( .A1(n7676), .A2(n7527), .ZN(n8716) );
  XNOR2_X1 U8649 ( .A(n8717), .B(n8718), .ZN(n8481) );
  XNOR2_X1 U8650 ( .A(n8719), .B(n8720), .ZN(n8717) );
  XOR2_X1 U8651 ( .A(n8721), .B(n8722), .Z(n8485) );
  XOR2_X1 U8652 ( .A(n8723), .B(n8724), .Z(n8722) );
  NAND2_X1 U8653 ( .A1(b_29_), .A2(a_18_), .ZN(n8724) );
  XNOR2_X1 U8654 ( .A(n8725), .B(n8726), .ZN(n8488) );
  XNOR2_X1 U8655 ( .A(n8727), .B(n8728), .ZN(n8725) );
  XNOR2_X1 U8656 ( .A(n8729), .B(n8730), .ZN(n8493) );
  XOR2_X1 U8657 ( .A(n8731), .B(n8732), .Z(n8729) );
  NOR2_X1 U8658 ( .A1(n7743), .A2(n7527), .ZN(n8732) );
  XNOR2_X1 U8659 ( .A(n8733), .B(n8734), .ZN(n8497) );
  XNOR2_X1 U8660 ( .A(n8735), .B(n8736), .ZN(n8733) );
  XNOR2_X1 U8661 ( .A(n8737), .B(n8738), .ZN(n8501) );
  XOR2_X1 U8662 ( .A(n8739), .B(n8740), .Z(n8737) );
  NOR2_X1 U8663 ( .A1(n7775), .A2(n7527), .ZN(n8740) );
  XOR2_X1 U8664 ( .A(n8741), .B(n8742), .Z(n8505) );
  XOR2_X1 U8665 ( .A(n8743), .B(n8744), .Z(n8741) );
  XOR2_X1 U8666 ( .A(n8745), .B(n8746), .Z(n8509) );
  XOR2_X1 U8667 ( .A(n8747), .B(n8748), .Z(n8746) );
  NAND2_X1 U8668 ( .A1(b_29_), .A2(a_12_), .ZN(n8748) );
  XNOR2_X1 U8669 ( .A(n8749), .B(n8750), .ZN(n8513) );
  XNOR2_X1 U8670 ( .A(n8751), .B(n8752), .ZN(n8749) );
  XOR2_X1 U8671 ( .A(n8753), .B(n8754), .Z(n8517) );
  XOR2_X1 U8672 ( .A(n8755), .B(n8756), .Z(n8753) );
  NOR2_X1 U8673 ( .A1(n7837), .A2(n7527), .ZN(n8756) );
  XOR2_X1 U8674 ( .A(n8757), .B(n8758), .Z(n8521) );
  XOR2_X1 U8675 ( .A(n8759), .B(n8760), .Z(n8757) );
  XOR2_X1 U8676 ( .A(n8761), .B(n8762), .Z(n8525) );
  XOR2_X1 U8677 ( .A(n8763), .B(n8764), .Z(n8761) );
  NOR2_X1 U8678 ( .A1(n8059), .A2(n7527), .ZN(n8764) );
  XOR2_X1 U8679 ( .A(n8765), .B(n8766), .Z(n8529) );
  XOR2_X1 U8680 ( .A(n8767), .B(n8768), .Z(n8765) );
  XOR2_X1 U8681 ( .A(n8769), .B(n8770), .Z(n8533) );
  XOR2_X1 U8682 ( .A(n8771), .B(n8772), .Z(n8770) );
  NAND2_X1 U8683 ( .A1(b_29_), .A2(a_6_), .ZN(n8772) );
  XNOR2_X1 U8684 ( .A(n8773), .B(n8774), .ZN(n8537) );
  XNOR2_X1 U8685 ( .A(n8775), .B(n8776), .ZN(n8773) );
  XNOR2_X1 U8686 ( .A(n8777), .B(n8778), .ZN(n8541) );
  XOR2_X1 U8687 ( .A(n8779), .B(n8780), .Z(n8777) );
  NOR2_X1 U8688 ( .A1(n7934), .A2(n7527), .ZN(n8780) );
  XOR2_X1 U8689 ( .A(n8781), .B(n8782), .Z(n8545) );
  XOR2_X1 U8690 ( .A(n8783), .B(n8784), .Z(n8781) );
  NOR2_X1 U8691 ( .A1(n7945), .A2(n7527), .ZN(n8784) );
  XNOR2_X1 U8692 ( .A(n8785), .B(n8786), .ZN(n8304) );
  XOR2_X1 U8693 ( .A(n8787), .B(n8788), .Z(n8786) );
  NAND2_X1 U8694 ( .A1(b_29_), .A2(a_1_), .ZN(n8788) );
  NAND2_X1 U8695 ( .A1(n8789), .A2(n8790), .ZN(n8092) );
  XOR2_X1 U8696 ( .A(n8289), .B(n8288), .Z(n8790) );
  AND2_X1 U8697 ( .A1(n8294), .A2(n8293), .ZN(n8789) );
  INV_X1 U8698 ( .A(n8301), .ZN(n8293) );
  XOR2_X1 U8699 ( .A(n8791), .B(n8792), .Z(n8301) );
  XNOR2_X1 U8700 ( .A(n8793), .B(n8794), .ZN(n8792) );
  NAND2_X1 U8701 ( .A1(n8556), .A2(n8795), .ZN(n8294) );
  NAND2_X1 U8702 ( .A1(n8555), .A2(n8557), .ZN(n8795) );
  NAND2_X1 U8703 ( .A1(n8796), .A2(n8797), .ZN(n8557) );
  NAND2_X1 U8704 ( .A1(b_29_), .A2(a_0_), .ZN(n8797) );
  INV_X1 U8705 ( .A(n8798), .ZN(n8796) );
  XOR2_X1 U8706 ( .A(n8799), .B(n8800), .Z(n8555) );
  XOR2_X1 U8707 ( .A(n8801), .B(n8802), .Z(n8799) );
  NAND2_X1 U8708 ( .A1(a_0_), .A2(n8798), .ZN(n8556) );
  NAND2_X1 U8709 ( .A1(n8803), .A2(n8804), .ZN(n8798) );
  NAND2_X1 U8710 ( .A1(n8805), .A2(b_29_), .ZN(n8804) );
  NOR2_X1 U8711 ( .A1(n8806), .A2(n7973), .ZN(n8805) );
  NOR2_X1 U8712 ( .A1(n8785), .A2(n8787), .ZN(n8806) );
  NAND2_X1 U8713 ( .A1(n8785), .A2(n8787), .ZN(n8803) );
  NAND2_X1 U8714 ( .A1(n8807), .A2(n8808), .ZN(n8787) );
  NAND2_X1 U8715 ( .A1(n8568), .A2(n8809), .ZN(n8808) );
  OR2_X1 U8716 ( .A1(n8567), .A2(n8569), .ZN(n8809) );
  NAND2_X1 U8717 ( .A1(n8810), .A2(n8811), .ZN(n8568) );
  NAND2_X1 U8718 ( .A1(n8812), .A2(b_29_), .ZN(n8811) );
  NOR2_X1 U8719 ( .A1(n8813), .A2(n7945), .ZN(n8812) );
  NOR2_X1 U8720 ( .A1(n8782), .A2(n8783), .ZN(n8813) );
  NAND2_X1 U8721 ( .A1(n8782), .A2(n8783), .ZN(n8810) );
  NAND2_X1 U8722 ( .A1(n8814), .A2(n8815), .ZN(n8783) );
  NAND2_X1 U8723 ( .A1(n8816), .A2(b_29_), .ZN(n8815) );
  NOR2_X1 U8724 ( .A1(n8817), .A2(n7934), .ZN(n8816) );
  NOR2_X1 U8725 ( .A1(n8778), .A2(n8779), .ZN(n8817) );
  NAND2_X1 U8726 ( .A1(n8778), .A2(n8779), .ZN(n8814) );
  NAND2_X1 U8727 ( .A1(n8818), .A2(n8819), .ZN(n8779) );
  NAND2_X1 U8728 ( .A1(n8775), .A2(n8820), .ZN(n8819) );
  NAND2_X1 U8729 ( .A1(n8776), .A2(n8774), .ZN(n8820) );
  NOR2_X1 U8730 ( .A1(n7527), .A2(n7914), .ZN(n8775) );
  OR2_X1 U8731 ( .A1(n8774), .A2(n8776), .ZN(n8818) );
  AND2_X1 U8732 ( .A1(n8821), .A2(n8822), .ZN(n8776) );
  NAND2_X1 U8733 ( .A1(n8823), .A2(b_29_), .ZN(n8822) );
  NOR2_X1 U8734 ( .A1(n8824), .A2(n8061), .ZN(n8823) );
  NOR2_X1 U8735 ( .A1(n8769), .A2(n8771), .ZN(n8824) );
  NAND2_X1 U8736 ( .A1(n8769), .A2(n8771), .ZN(n8821) );
  NAND2_X1 U8737 ( .A1(n8825), .A2(n8826), .ZN(n8771) );
  NAND2_X1 U8738 ( .A1(n8768), .A2(n8827), .ZN(n8826) );
  OR2_X1 U8739 ( .A1(n8767), .A2(n8766), .ZN(n8827) );
  NOR2_X1 U8740 ( .A1(n7527), .A2(n7884), .ZN(n8768) );
  NAND2_X1 U8741 ( .A1(n8766), .A2(n8767), .ZN(n8825) );
  NAND2_X1 U8742 ( .A1(n8828), .A2(n8829), .ZN(n8767) );
  NAND2_X1 U8743 ( .A1(n8830), .A2(b_29_), .ZN(n8829) );
  NOR2_X1 U8744 ( .A1(n8831), .A2(n8059), .ZN(n8830) );
  NOR2_X1 U8745 ( .A1(n8762), .A2(n8763), .ZN(n8831) );
  NAND2_X1 U8746 ( .A1(n8762), .A2(n8763), .ZN(n8828) );
  NAND2_X1 U8747 ( .A1(n8832), .A2(n8833), .ZN(n8763) );
  NAND2_X1 U8748 ( .A1(n8760), .A2(n8834), .ZN(n8833) );
  OR2_X1 U8749 ( .A1(n8759), .A2(n8758), .ZN(n8834) );
  NOR2_X1 U8750 ( .A1(n7527), .A2(n7848), .ZN(n8760) );
  NAND2_X1 U8751 ( .A1(n8758), .A2(n8759), .ZN(n8832) );
  NAND2_X1 U8752 ( .A1(n8835), .A2(n8836), .ZN(n8759) );
  NAND2_X1 U8753 ( .A1(n8837), .A2(b_29_), .ZN(n8836) );
  NOR2_X1 U8754 ( .A1(n8838), .A2(n7837), .ZN(n8837) );
  NOR2_X1 U8755 ( .A1(n8754), .A2(n8755), .ZN(n8838) );
  NAND2_X1 U8756 ( .A1(n8754), .A2(n8755), .ZN(n8835) );
  NAND2_X1 U8757 ( .A1(n8839), .A2(n8840), .ZN(n8755) );
  NAND2_X1 U8758 ( .A1(n8751), .A2(n8841), .ZN(n8840) );
  NAND2_X1 U8759 ( .A1(n8752), .A2(n8750), .ZN(n8841) );
  NOR2_X1 U8760 ( .A1(n7527), .A2(n7817), .ZN(n8751) );
  OR2_X1 U8761 ( .A1(n8750), .A2(n8752), .ZN(n8839) );
  AND2_X1 U8762 ( .A1(n8842), .A2(n8843), .ZN(n8752) );
  NAND2_X1 U8763 ( .A1(n8844), .A2(b_29_), .ZN(n8843) );
  NOR2_X1 U8764 ( .A1(n8845), .A2(n7806), .ZN(n8844) );
  NOR2_X1 U8765 ( .A1(n8745), .A2(n8747), .ZN(n8845) );
  NAND2_X1 U8766 ( .A1(n8745), .A2(n8747), .ZN(n8842) );
  NAND2_X1 U8767 ( .A1(n8846), .A2(n8847), .ZN(n8747) );
  NAND2_X1 U8768 ( .A1(n8744), .A2(n8848), .ZN(n8847) );
  OR2_X1 U8769 ( .A1(n8743), .A2(n8742), .ZN(n8848) );
  NOR2_X1 U8770 ( .A1(n7527), .A2(n7786), .ZN(n8744) );
  NAND2_X1 U8771 ( .A1(n8742), .A2(n8743), .ZN(n8846) );
  NAND2_X1 U8772 ( .A1(n8849), .A2(n8850), .ZN(n8743) );
  NAND2_X1 U8773 ( .A1(n8851), .A2(b_29_), .ZN(n8850) );
  NOR2_X1 U8774 ( .A1(n8852), .A2(n7775), .ZN(n8851) );
  NOR2_X1 U8775 ( .A1(n8738), .A2(n8739), .ZN(n8852) );
  NAND2_X1 U8776 ( .A1(n8738), .A2(n8739), .ZN(n8849) );
  NAND2_X1 U8777 ( .A1(n8853), .A2(n8854), .ZN(n8739) );
  NAND2_X1 U8778 ( .A1(n8735), .A2(n8855), .ZN(n8854) );
  NAND2_X1 U8779 ( .A1(n8736), .A2(n8734), .ZN(n8855) );
  NOR2_X1 U8780 ( .A1(n7527), .A2(n7754), .ZN(n8735) );
  OR2_X1 U8781 ( .A1(n8734), .A2(n8736), .ZN(n8853) );
  AND2_X1 U8782 ( .A1(n8856), .A2(n8857), .ZN(n8736) );
  NAND2_X1 U8783 ( .A1(n8858), .A2(b_29_), .ZN(n8857) );
  NOR2_X1 U8784 ( .A1(n8859), .A2(n7743), .ZN(n8858) );
  NOR2_X1 U8785 ( .A1(n8730), .A2(n8731), .ZN(n8859) );
  NAND2_X1 U8786 ( .A1(n8730), .A2(n8731), .ZN(n8856) );
  NAND2_X1 U8787 ( .A1(n8860), .A2(n8861), .ZN(n8731) );
  NAND2_X1 U8788 ( .A1(n8728), .A2(n8862), .ZN(n8861) );
  NAND2_X1 U8789 ( .A1(n8727), .A2(n8726), .ZN(n8862) );
  NOR2_X1 U8790 ( .A1(n7527), .A2(n7723), .ZN(n8728) );
  OR2_X1 U8791 ( .A1(n8726), .A2(n8727), .ZN(n8860) );
  AND2_X1 U8792 ( .A1(n8863), .A2(n8864), .ZN(n8727) );
  NAND2_X1 U8793 ( .A1(n8865), .A2(b_29_), .ZN(n8864) );
  NOR2_X1 U8794 ( .A1(n8866), .A2(n7707), .ZN(n8865) );
  NOR2_X1 U8795 ( .A1(n8721), .A2(n8723), .ZN(n8866) );
  NAND2_X1 U8796 ( .A1(n8721), .A2(n8723), .ZN(n8863) );
  NAND2_X1 U8797 ( .A1(n8867), .A2(n8868), .ZN(n8723) );
  NAND2_X1 U8798 ( .A1(n8720), .A2(n8869), .ZN(n8868) );
  NAND2_X1 U8799 ( .A1(n8719), .A2(n8718), .ZN(n8869) );
  NOR2_X1 U8800 ( .A1(n7527), .A2(n7687), .ZN(n8720) );
  OR2_X1 U8801 ( .A1(n8718), .A2(n8719), .ZN(n8867) );
  AND2_X1 U8802 ( .A1(n8870), .A2(n8871), .ZN(n8719) );
  NAND2_X1 U8803 ( .A1(n8872), .A2(b_29_), .ZN(n8871) );
  NOR2_X1 U8804 ( .A1(n8873), .A2(n7676), .ZN(n8872) );
  NOR2_X1 U8805 ( .A1(n8714), .A2(n8715), .ZN(n8873) );
  NAND2_X1 U8806 ( .A1(n8714), .A2(n8715), .ZN(n8870) );
  NAND2_X1 U8807 ( .A1(n8874), .A2(n8875), .ZN(n8715) );
  NAND2_X1 U8808 ( .A1(n8712), .A2(n8876), .ZN(n8875) );
  NAND2_X1 U8809 ( .A1(n8711), .A2(n8710), .ZN(n8876) );
  NOR2_X1 U8810 ( .A1(n7527), .A2(n7656), .ZN(n8712) );
  OR2_X1 U8811 ( .A1(n8710), .A2(n8711), .ZN(n8874) );
  AND2_X1 U8812 ( .A1(n8877), .A2(n8878), .ZN(n8711) );
  NAND2_X1 U8813 ( .A1(n8879), .A2(b_29_), .ZN(n8878) );
  NOR2_X1 U8814 ( .A1(n8880), .A2(n7645), .ZN(n8879) );
  NOR2_X1 U8815 ( .A1(n8706), .A2(n8707), .ZN(n8880) );
  NAND2_X1 U8816 ( .A1(n8706), .A2(n8707), .ZN(n8877) );
  NAND2_X1 U8817 ( .A1(n8881), .A2(n8882), .ZN(n8707) );
  NAND2_X1 U8818 ( .A1(n8703), .A2(n8883), .ZN(n8882) );
  NAND2_X1 U8819 ( .A1(n8704), .A2(n8702), .ZN(n8883) );
  NOR2_X1 U8820 ( .A1(n7527), .A2(n7624), .ZN(n8703) );
  OR2_X1 U8821 ( .A1(n8702), .A2(n8704), .ZN(n8881) );
  AND2_X1 U8822 ( .A1(n8884), .A2(n8885), .ZN(n8704) );
  NAND2_X1 U8823 ( .A1(n8886), .A2(b_29_), .ZN(n8885) );
  NOR2_X1 U8824 ( .A1(n8887), .A2(n7613), .ZN(n8886) );
  NOR2_X1 U8825 ( .A1(n8697), .A2(n8699), .ZN(n8887) );
  NAND2_X1 U8826 ( .A1(n8697), .A2(n8699), .ZN(n8884) );
  NAND2_X1 U8827 ( .A1(n8888), .A2(n8889), .ZN(n8699) );
  NAND2_X1 U8828 ( .A1(n8696), .A2(n8890), .ZN(n8889) );
  OR2_X1 U8829 ( .A1(n8695), .A2(n8693), .ZN(n8890) );
  NOR2_X1 U8830 ( .A1(n7527), .A2(n7593), .ZN(n8696) );
  NAND2_X1 U8831 ( .A1(n8693), .A2(n8695), .ZN(n8888) );
  NAND2_X1 U8832 ( .A1(n8891), .A2(n8892), .ZN(n8695) );
  NAND2_X1 U8833 ( .A1(n8893), .A2(b_29_), .ZN(n8892) );
  NOR2_X1 U8834 ( .A1(n8894), .A2(n8052), .ZN(n8893) );
  NOR2_X1 U8835 ( .A1(n8689), .A2(n8691), .ZN(n8894) );
  NAND2_X1 U8836 ( .A1(n8689), .A2(n8691), .ZN(n8891) );
  NAND2_X1 U8837 ( .A1(n8895), .A2(n8896), .ZN(n8691) );
  NAND2_X1 U8838 ( .A1(n8688), .A2(n8897), .ZN(n8896) );
  OR2_X1 U8839 ( .A1(n8687), .A2(n8685), .ZN(n8897) );
  NOR2_X1 U8840 ( .A1(n7527), .A2(n7563), .ZN(n8688) );
  NAND2_X1 U8841 ( .A1(n8685), .A2(n8687), .ZN(n8895) );
  NAND2_X1 U8842 ( .A1(n8683), .A2(n8898), .ZN(n8687) );
  NAND2_X1 U8843 ( .A1(n8682), .A2(n8684), .ZN(n8898) );
  NAND2_X1 U8844 ( .A1(n8899), .A2(n8900), .ZN(n8684) );
  NAND2_X1 U8845 ( .A1(b_29_), .A2(a_28_), .ZN(n8900) );
  INV_X1 U8846 ( .A(n8901), .ZN(n8899) );
  XOR2_X1 U8847 ( .A(n8902), .B(n8903), .Z(n8682) );
  NOR2_X1 U8848 ( .A1(n7529), .A2(n8050), .ZN(n8903) );
  XOR2_X1 U8849 ( .A(n8904), .B(n8905), .Z(n8902) );
  NAND2_X1 U8850 ( .A1(a_28_), .A2(n8901), .ZN(n8683) );
  NAND2_X1 U8851 ( .A1(n8906), .A2(n8907), .ZN(n8901) );
  NAND2_X1 U8852 ( .A1(n8666), .A2(n8908), .ZN(n8907) );
  NAND2_X1 U8853 ( .A1(n8667), .A2(n8042), .ZN(n8908) );
  INV_X1 U8854 ( .A(n8909), .ZN(n8667) );
  AND2_X1 U8855 ( .A1(n8910), .A2(b_29_), .ZN(n8666) );
  NOR2_X1 U8856 ( .A1(n8451), .A2(n8050), .ZN(n8910) );
  NAND2_X1 U8857 ( .A1(n7521), .A2(n8909), .ZN(n8906) );
  NAND2_X1 U8858 ( .A1(n8911), .A2(n8912), .ZN(n8909) );
  NAND2_X1 U8859 ( .A1(n8913), .A2(b_27_), .ZN(n8912) );
  NOR2_X1 U8860 ( .A1(n8914), .A2(n8048), .ZN(n8913) );
  NOR2_X1 U8861 ( .A1(n8676), .A2(n8050), .ZN(n8914) );
  NAND2_X1 U8862 ( .A1(n8915), .A2(b_28_), .ZN(n8911) );
  NOR2_X1 U8863 ( .A1(n8916), .A2(n7515), .ZN(n8915) );
  NOR2_X1 U8864 ( .A1(n8679), .A2(n7564), .ZN(n8916) );
  INV_X1 U8865 ( .A(n8042), .ZN(n7521) );
  NAND2_X1 U8866 ( .A1(b_29_), .A2(a_29_), .ZN(n8042) );
  XOR2_X1 U8867 ( .A(n8917), .B(n8918), .Z(n8685) );
  XOR2_X1 U8868 ( .A(n7540), .B(n8919), .Z(n8917) );
  XNOR2_X1 U8869 ( .A(n8920), .B(n8921), .ZN(n8689) );
  XNOR2_X1 U8870 ( .A(n8922), .B(n8923), .ZN(n8920) );
  XOR2_X1 U8871 ( .A(n8924), .B(n8925), .Z(n8693) );
  XNOR2_X1 U8872 ( .A(n8926), .B(n8927), .ZN(n8924) );
  NAND2_X1 U8873 ( .A1(b_28_), .A2(a_26_), .ZN(n8926) );
  XNOR2_X1 U8874 ( .A(n8928), .B(n8929), .ZN(n8697) );
  XNOR2_X1 U8875 ( .A(n8930), .B(n8931), .ZN(n8928) );
  XOR2_X1 U8876 ( .A(n8932), .B(n8933), .Z(n8702) );
  XOR2_X1 U8877 ( .A(n8934), .B(n8935), .Z(n8933) );
  NAND2_X1 U8878 ( .A1(b_28_), .A2(a_24_), .ZN(n8935) );
  XNOR2_X1 U8879 ( .A(n8936), .B(n8937), .ZN(n8706) );
  XNOR2_X1 U8880 ( .A(n8938), .B(n8939), .ZN(n8936) );
  XNOR2_X1 U8881 ( .A(n8940), .B(n8941), .ZN(n8710) );
  XOR2_X1 U8882 ( .A(n8942), .B(n8943), .Z(n8940) );
  NOR2_X1 U8883 ( .A1(n7645), .A2(n8050), .ZN(n8943) );
  XNOR2_X1 U8884 ( .A(n8944), .B(n8945), .ZN(n8714) );
  XNOR2_X1 U8885 ( .A(n8946), .B(n8947), .ZN(n8944) );
  XNOR2_X1 U8886 ( .A(n8948), .B(n8949), .ZN(n8718) );
  XOR2_X1 U8887 ( .A(n8950), .B(n8951), .Z(n8948) );
  NOR2_X1 U8888 ( .A1(n7676), .A2(n8050), .ZN(n8951) );
  XNOR2_X1 U8889 ( .A(n8952), .B(n8953), .ZN(n8721) );
  XNOR2_X1 U8890 ( .A(n8954), .B(n8955), .ZN(n8952) );
  XNOR2_X1 U8891 ( .A(n8956), .B(n8957), .ZN(n8726) );
  XOR2_X1 U8892 ( .A(n8958), .B(n8959), .Z(n8956) );
  NOR2_X1 U8893 ( .A1(n7707), .A2(n8050), .ZN(n8959) );
  XNOR2_X1 U8894 ( .A(n8960), .B(n8961), .ZN(n8730) );
  XNOR2_X1 U8895 ( .A(n8962), .B(n8963), .ZN(n8960) );
  XNOR2_X1 U8896 ( .A(n8964), .B(n8965), .ZN(n8734) );
  XOR2_X1 U8897 ( .A(n8966), .B(n8967), .Z(n8964) );
  NOR2_X1 U8898 ( .A1(n7743), .A2(n8050), .ZN(n8967) );
  XNOR2_X1 U8899 ( .A(n8968), .B(n8969), .ZN(n8738) );
  XNOR2_X1 U8900 ( .A(n8970), .B(n8971), .ZN(n8968) );
  XNOR2_X1 U8901 ( .A(n8972), .B(n8973), .ZN(n8742) );
  XOR2_X1 U8902 ( .A(n8974), .B(n8975), .Z(n8973) );
  NAND2_X1 U8903 ( .A1(b_28_), .A2(a_14_), .ZN(n8975) );
  XNOR2_X1 U8904 ( .A(n8976), .B(n8977), .ZN(n8745) );
  XNOR2_X1 U8905 ( .A(n8978), .B(n8979), .ZN(n8976) );
  XNOR2_X1 U8906 ( .A(n8980), .B(n8981), .ZN(n8750) );
  XOR2_X1 U8907 ( .A(n8982), .B(n8983), .Z(n8980) );
  NOR2_X1 U8908 ( .A1(n7806), .A2(n8050), .ZN(n8983) );
  XOR2_X1 U8909 ( .A(n8984), .B(n8985), .Z(n8754) );
  XOR2_X1 U8910 ( .A(n8986), .B(n8987), .Z(n8984) );
  XNOR2_X1 U8911 ( .A(n8988), .B(n8989), .ZN(n8758) );
  XOR2_X1 U8912 ( .A(n8990), .B(n8991), .Z(n8989) );
  NAND2_X1 U8913 ( .A1(b_28_), .A2(a_10_), .ZN(n8991) );
  XOR2_X1 U8914 ( .A(n8992), .B(n8993), .Z(n8762) );
  XOR2_X1 U8915 ( .A(n8994), .B(n8995), .Z(n8992) );
  XNOR2_X1 U8916 ( .A(n8996), .B(n8997), .ZN(n8766) );
  XOR2_X1 U8917 ( .A(n8998), .B(n8999), .Z(n8997) );
  NAND2_X1 U8918 ( .A1(b_28_), .A2(a_8_), .ZN(n8999) );
  XNOR2_X1 U8919 ( .A(n9000), .B(n9001), .ZN(n8769) );
  XNOR2_X1 U8920 ( .A(n9002), .B(n9003), .ZN(n9000) );
  XNOR2_X1 U8921 ( .A(n9004), .B(n9005), .ZN(n8774) );
  XOR2_X1 U8922 ( .A(n9006), .B(n9007), .Z(n9004) );
  NOR2_X1 U8923 ( .A1(n8061), .A2(n8050), .ZN(n9007) );
  XNOR2_X1 U8924 ( .A(n9008), .B(n9009), .ZN(n8778) );
  XNOR2_X1 U8925 ( .A(n9010), .B(n9011), .ZN(n9009) );
  XNOR2_X1 U8926 ( .A(n9012), .B(n9013), .ZN(n8782) );
  XOR2_X1 U8927 ( .A(n9014), .B(n9015), .Z(n9013) );
  NAND2_X1 U8928 ( .A1(b_28_), .A2(a_4_), .ZN(n9015) );
  NAND2_X1 U8929 ( .A1(n8569), .A2(n8567), .ZN(n8807) );
  XOR2_X1 U8930 ( .A(n9016), .B(n9017), .Z(n8567) );
  XOR2_X1 U8931 ( .A(n9018), .B(n9019), .Z(n9016) );
  NOR2_X1 U8932 ( .A1(n7945), .A2(n8050), .ZN(n9019) );
  NOR2_X1 U8933 ( .A1(n7527), .A2(n7965), .ZN(n8569) );
  XNOR2_X1 U8934 ( .A(n9020), .B(n9021), .ZN(n8785) );
  XNOR2_X1 U8935 ( .A(n9022), .B(n9023), .ZN(n9020) );
  NAND2_X1 U8936 ( .A1(n9024), .A2(n9025), .ZN(n8096) );
  NOR2_X1 U8937 ( .A1(n8285), .A2(n8289), .ZN(n9025) );
  INV_X1 U8938 ( .A(n8295), .ZN(n8289) );
  NAND2_X1 U8939 ( .A1(n9026), .A2(n9027), .ZN(n8295) );
  NAND2_X1 U8940 ( .A1(n8794), .A2(n9028), .ZN(n9027) );
  OR2_X1 U8941 ( .A1(n8793), .A2(n8791), .ZN(n9028) );
  NOR2_X1 U8942 ( .A1(n8050), .A2(n8307), .ZN(n8794) );
  NAND2_X1 U8943 ( .A1(n8791), .A2(n8793), .ZN(n9026) );
  NAND2_X1 U8944 ( .A1(n9029), .A2(n9030), .ZN(n8793) );
  NAND2_X1 U8945 ( .A1(n8802), .A2(n9031), .ZN(n9030) );
  OR2_X1 U8946 ( .A1(n8801), .A2(n8800), .ZN(n9031) );
  NOR2_X1 U8947 ( .A1(n8050), .A2(n7973), .ZN(n8802) );
  NAND2_X1 U8948 ( .A1(n8800), .A2(n8801), .ZN(n9029) );
  NAND2_X1 U8949 ( .A1(n9032), .A2(n9033), .ZN(n8801) );
  NAND2_X1 U8950 ( .A1(n9022), .A2(n9034), .ZN(n9033) );
  NAND2_X1 U8951 ( .A1(n9021), .A2(n9023), .ZN(n9034) );
  NAND2_X1 U8952 ( .A1(n9035), .A2(n9036), .ZN(n9022) );
  NAND2_X1 U8953 ( .A1(n9037), .A2(b_28_), .ZN(n9036) );
  NOR2_X1 U8954 ( .A1(n9038), .A2(n7945), .ZN(n9037) );
  NOR2_X1 U8955 ( .A1(n9017), .A2(n9018), .ZN(n9038) );
  NAND2_X1 U8956 ( .A1(n9017), .A2(n9018), .ZN(n9035) );
  NAND2_X1 U8957 ( .A1(n9039), .A2(n9040), .ZN(n9018) );
  NAND2_X1 U8958 ( .A1(n9041), .A2(b_28_), .ZN(n9040) );
  NOR2_X1 U8959 ( .A1(n9042), .A2(n7934), .ZN(n9041) );
  NOR2_X1 U8960 ( .A1(n9012), .A2(n9014), .ZN(n9042) );
  NAND2_X1 U8961 ( .A1(n9012), .A2(n9014), .ZN(n9039) );
  NAND2_X1 U8962 ( .A1(n9043), .A2(n9044), .ZN(n9014) );
  NAND2_X1 U8963 ( .A1(n9011), .A2(n9045), .ZN(n9044) );
  OR2_X1 U8964 ( .A1(n9010), .A2(n9008), .ZN(n9045) );
  NOR2_X1 U8965 ( .A1(n8050), .A2(n7914), .ZN(n9011) );
  NAND2_X1 U8966 ( .A1(n9008), .A2(n9010), .ZN(n9043) );
  NAND2_X1 U8967 ( .A1(n9046), .A2(n9047), .ZN(n9010) );
  NAND2_X1 U8968 ( .A1(n9048), .A2(b_28_), .ZN(n9047) );
  NOR2_X1 U8969 ( .A1(n9049), .A2(n8061), .ZN(n9048) );
  NOR2_X1 U8970 ( .A1(n9005), .A2(n9006), .ZN(n9049) );
  NAND2_X1 U8971 ( .A1(n9005), .A2(n9006), .ZN(n9046) );
  NAND2_X1 U8972 ( .A1(n9050), .A2(n9051), .ZN(n9006) );
  NAND2_X1 U8973 ( .A1(n9003), .A2(n9052), .ZN(n9051) );
  NAND2_X1 U8974 ( .A1(n9002), .A2(n9001), .ZN(n9052) );
  NOR2_X1 U8975 ( .A1(n8050), .A2(n7884), .ZN(n9003) );
  OR2_X1 U8976 ( .A1(n9001), .A2(n9002), .ZN(n9050) );
  AND2_X1 U8977 ( .A1(n9053), .A2(n9054), .ZN(n9002) );
  NAND2_X1 U8978 ( .A1(n9055), .A2(b_28_), .ZN(n9054) );
  NOR2_X1 U8979 ( .A1(n9056), .A2(n8059), .ZN(n9055) );
  NOR2_X1 U8980 ( .A1(n8996), .A2(n8998), .ZN(n9056) );
  NAND2_X1 U8981 ( .A1(n8996), .A2(n8998), .ZN(n9053) );
  NAND2_X1 U8982 ( .A1(n9057), .A2(n9058), .ZN(n8998) );
  NAND2_X1 U8983 ( .A1(n8995), .A2(n9059), .ZN(n9058) );
  OR2_X1 U8984 ( .A1(n8994), .A2(n8993), .ZN(n9059) );
  NOR2_X1 U8985 ( .A1(n8050), .A2(n7848), .ZN(n8995) );
  NAND2_X1 U8986 ( .A1(n8993), .A2(n8994), .ZN(n9057) );
  NAND2_X1 U8987 ( .A1(n9060), .A2(n9061), .ZN(n8994) );
  NAND2_X1 U8988 ( .A1(n9062), .A2(b_28_), .ZN(n9061) );
  NOR2_X1 U8989 ( .A1(n9063), .A2(n7837), .ZN(n9062) );
  NOR2_X1 U8990 ( .A1(n8988), .A2(n8990), .ZN(n9063) );
  NAND2_X1 U8991 ( .A1(n8988), .A2(n8990), .ZN(n9060) );
  NAND2_X1 U8992 ( .A1(n9064), .A2(n9065), .ZN(n8990) );
  NAND2_X1 U8993 ( .A1(n8987), .A2(n9066), .ZN(n9065) );
  OR2_X1 U8994 ( .A1(n8986), .A2(n8985), .ZN(n9066) );
  NOR2_X1 U8995 ( .A1(n8050), .A2(n7817), .ZN(n8987) );
  NAND2_X1 U8996 ( .A1(n8985), .A2(n8986), .ZN(n9064) );
  NAND2_X1 U8997 ( .A1(n9067), .A2(n9068), .ZN(n8986) );
  NAND2_X1 U8998 ( .A1(n9069), .A2(b_28_), .ZN(n9068) );
  NOR2_X1 U8999 ( .A1(n9070), .A2(n7806), .ZN(n9069) );
  NOR2_X1 U9000 ( .A1(n8981), .A2(n8982), .ZN(n9070) );
  NAND2_X1 U9001 ( .A1(n8981), .A2(n8982), .ZN(n9067) );
  NAND2_X1 U9002 ( .A1(n9071), .A2(n9072), .ZN(n8982) );
  NAND2_X1 U9003 ( .A1(n8979), .A2(n9073), .ZN(n9072) );
  NAND2_X1 U9004 ( .A1(n8978), .A2(n8977), .ZN(n9073) );
  NOR2_X1 U9005 ( .A1(n8050), .A2(n7786), .ZN(n8979) );
  OR2_X1 U9006 ( .A1(n8977), .A2(n8978), .ZN(n9071) );
  AND2_X1 U9007 ( .A1(n9074), .A2(n9075), .ZN(n8978) );
  NAND2_X1 U9008 ( .A1(n9076), .A2(b_28_), .ZN(n9075) );
  NOR2_X1 U9009 ( .A1(n9077), .A2(n7775), .ZN(n9076) );
  NOR2_X1 U9010 ( .A1(n8972), .A2(n8974), .ZN(n9077) );
  NAND2_X1 U9011 ( .A1(n8972), .A2(n8974), .ZN(n9074) );
  NAND2_X1 U9012 ( .A1(n9078), .A2(n9079), .ZN(n8974) );
  NAND2_X1 U9013 ( .A1(n8971), .A2(n9080), .ZN(n9079) );
  NAND2_X1 U9014 ( .A1(n8970), .A2(n8969), .ZN(n9080) );
  NOR2_X1 U9015 ( .A1(n8050), .A2(n7754), .ZN(n8971) );
  OR2_X1 U9016 ( .A1(n8969), .A2(n8970), .ZN(n9078) );
  AND2_X1 U9017 ( .A1(n9081), .A2(n9082), .ZN(n8970) );
  NAND2_X1 U9018 ( .A1(n9083), .A2(b_28_), .ZN(n9082) );
  NOR2_X1 U9019 ( .A1(n9084), .A2(n7743), .ZN(n9083) );
  NOR2_X1 U9020 ( .A1(n8965), .A2(n8966), .ZN(n9084) );
  NAND2_X1 U9021 ( .A1(n8965), .A2(n8966), .ZN(n9081) );
  NAND2_X1 U9022 ( .A1(n9085), .A2(n9086), .ZN(n8966) );
  NAND2_X1 U9023 ( .A1(n8963), .A2(n9087), .ZN(n9086) );
  NAND2_X1 U9024 ( .A1(n8962), .A2(n8961), .ZN(n9087) );
  NOR2_X1 U9025 ( .A1(n8050), .A2(n7723), .ZN(n8963) );
  OR2_X1 U9026 ( .A1(n8961), .A2(n8962), .ZN(n9085) );
  AND2_X1 U9027 ( .A1(n9088), .A2(n9089), .ZN(n8962) );
  NAND2_X1 U9028 ( .A1(n9090), .A2(b_28_), .ZN(n9089) );
  NOR2_X1 U9029 ( .A1(n9091), .A2(n7707), .ZN(n9090) );
  NOR2_X1 U9030 ( .A1(n8957), .A2(n8958), .ZN(n9091) );
  NAND2_X1 U9031 ( .A1(n8957), .A2(n8958), .ZN(n9088) );
  NAND2_X1 U9032 ( .A1(n9092), .A2(n9093), .ZN(n8958) );
  NAND2_X1 U9033 ( .A1(n8955), .A2(n9094), .ZN(n9093) );
  NAND2_X1 U9034 ( .A1(n8954), .A2(n8953), .ZN(n9094) );
  NOR2_X1 U9035 ( .A1(n8050), .A2(n7687), .ZN(n8955) );
  OR2_X1 U9036 ( .A1(n8953), .A2(n8954), .ZN(n9092) );
  AND2_X1 U9037 ( .A1(n9095), .A2(n9096), .ZN(n8954) );
  NAND2_X1 U9038 ( .A1(n9097), .A2(b_28_), .ZN(n9096) );
  NOR2_X1 U9039 ( .A1(n9098), .A2(n7676), .ZN(n9097) );
  NOR2_X1 U9040 ( .A1(n8949), .A2(n8950), .ZN(n9098) );
  NAND2_X1 U9041 ( .A1(n8949), .A2(n8950), .ZN(n9095) );
  NAND2_X1 U9042 ( .A1(n9099), .A2(n9100), .ZN(n8950) );
  NAND2_X1 U9043 ( .A1(n8947), .A2(n9101), .ZN(n9100) );
  NAND2_X1 U9044 ( .A1(n8946), .A2(n8945), .ZN(n9101) );
  NOR2_X1 U9045 ( .A1(n8050), .A2(n7656), .ZN(n8947) );
  OR2_X1 U9046 ( .A1(n8945), .A2(n8946), .ZN(n9099) );
  AND2_X1 U9047 ( .A1(n9102), .A2(n9103), .ZN(n8946) );
  NAND2_X1 U9048 ( .A1(n9104), .A2(b_28_), .ZN(n9103) );
  NOR2_X1 U9049 ( .A1(n9105), .A2(n7645), .ZN(n9104) );
  NOR2_X1 U9050 ( .A1(n8941), .A2(n8942), .ZN(n9105) );
  NAND2_X1 U9051 ( .A1(n8941), .A2(n8942), .ZN(n9102) );
  NAND2_X1 U9052 ( .A1(n9106), .A2(n9107), .ZN(n8942) );
  NAND2_X1 U9053 ( .A1(n8938), .A2(n9108), .ZN(n9107) );
  NAND2_X1 U9054 ( .A1(n8939), .A2(n8937), .ZN(n9108) );
  NOR2_X1 U9055 ( .A1(n8050), .A2(n7624), .ZN(n8938) );
  OR2_X1 U9056 ( .A1(n8937), .A2(n8939), .ZN(n9106) );
  AND2_X1 U9057 ( .A1(n9109), .A2(n9110), .ZN(n8939) );
  NAND2_X1 U9058 ( .A1(n9111), .A2(b_28_), .ZN(n9110) );
  NOR2_X1 U9059 ( .A1(n9112), .A2(n7613), .ZN(n9111) );
  NOR2_X1 U9060 ( .A1(n8932), .A2(n8934), .ZN(n9112) );
  NAND2_X1 U9061 ( .A1(n8932), .A2(n8934), .ZN(n9109) );
  NAND2_X1 U9062 ( .A1(n9113), .A2(n9114), .ZN(n8934) );
  NAND2_X1 U9063 ( .A1(n8931), .A2(n9115), .ZN(n9114) );
  NAND2_X1 U9064 ( .A1(n8930), .A2(n8929), .ZN(n9115) );
  NOR2_X1 U9065 ( .A1(n8050), .A2(n7593), .ZN(n8931) );
  OR2_X1 U9066 ( .A1(n8929), .A2(n8930), .ZN(n9113) );
  AND2_X1 U9067 ( .A1(n9116), .A2(n9117), .ZN(n8930) );
  NAND2_X1 U9068 ( .A1(n9118), .A2(b_28_), .ZN(n9117) );
  NOR2_X1 U9069 ( .A1(n9119), .A2(n8052), .ZN(n9118) );
  NOR2_X1 U9070 ( .A1(n8925), .A2(n8927), .ZN(n9119) );
  NAND2_X1 U9071 ( .A1(n8925), .A2(n8927), .ZN(n9116) );
  NAND2_X1 U9072 ( .A1(n9120), .A2(n9121), .ZN(n8927) );
  NAND2_X1 U9073 ( .A1(n8923), .A2(n9122), .ZN(n9121) );
  NAND2_X1 U9074 ( .A1(n8922), .A2(n8921), .ZN(n9122) );
  NOR2_X1 U9075 ( .A1(n8050), .A2(n7563), .ZN(n8923) );
  OR2_X1 U9076 ( .A1(n8921), .A2(n8922), .ZN(n9120) );
  AND2_X1 U9077 ( .A1(n9123), .A2(n9124), .ZN(n8922) );
  NAND2_X1 U9078 ( .A1(n8918), .A2(n9125), .ZN(n9124) );
  NAND2_X1 U9079 ( .A1(n8919), .A2(n7540), .ZN(n9125) );
  INV_X1 U9080 ( .A(n9126), .ZN(n8919) );
  XOR2_X1 U9081 ( .A(n9127), .B(n9128), .Z(n8918) );
  NOR2_X1 U9082 ( .A1(n7529), .A2(n7564), .ZN(n9128) );
  XOR2_X1 U9083 ( .A(n9129), .B(n9130), .Z(n9127) );
  NAND2_X1 U9084 ( .A1(n9131), .A2(n9126), .ZN(n9123) );
  NAND2_X1 U9085 ( .A1(n9132), .A2(n9133), .ZN(n9126) );
  NAND2_X1 U9086 ( .A1(n9134), .A2(b_28_), .ZN(n9133) );
  NOR2_X1 U9087 ( .A1(n9135), .A2(n7529), .ZN(n9134) );
  NOR2_X1 U9088 ( .A1(n8904), .A2(n8905), .ZN(n9135) );
  NAND2_X1 U9089 ( .A1(n8904), .A2(n8905), .ZN(n9132) );
  NAND2_X1 U9090 ( .A1(n9136), .A2(n9137), .ZN(n8905) );
  NAND2_X1 U9091 ( .A1(n9138), .A2(b_26_), .ZN(n9137) );
  NOR2_X1 U9092 ( .A1(n9139), .A2(n8048), .ZN(n9138) );
  NOR2_X1 U9093 ( .A1(n8676), .A2(n7564), .ZN(n9139) );
  NAND2_X1 U9094 ( .A1(n9140), .A2(b_27_), .ZN(n9136) );
  NOR2_X1 U9095 ( .A1(n9141), .A2(n7515), .ZN(n9140) );
  NOR2_X1 U9096 ( .A1(n8679), .A2(n8051), .ZN(n9141) );
  AND2_X1 U9097 ( .A1(n9142), .A2(b_28_), .ZN(n8904) );
  INV_X1 U9098 ( .A(n7540), .ZN(n9131) );
  NAND2_X1 U9099 ( .A1(b_28_), .A2(a_28_), .ZN(n7540) );
  XOR2_X1 U9100 ( .A(n9143), .B(n9144), .Z(n8921) );
  NAND2_X1 U9101 ( .A1(n9145), .A2(n9146), .ZN(n9143) );
  XNOR2_X1 U9102 ( .A(n9147), .B(n9148), .ZN(n8925) );
  XOR2_X1 U9103 ( .A(n9149), .B(n8038), .Z(n9147) );
  XNOR2_X1 U9104 ( .A(n9150), .B(n9151), .ZN(n8929) );
  XNOR2_X1 U9105 ( .A(n9152), .B(n9153), .ZN(n9150) );
  NAND2_X1 U9106 ( .A1(b_27_), .A2(a_26_), .ZN(n9152) );
  XNOR2_X1 U9107 ( .A(n9154), .B(n9155), .ZN(n8932) );
  XNOR2_X1 U9108 ( .A(n9156), .B(n9157), .ZN(n9154) );
  XOR2_X1 U9109 ( .A(n9158), .B(n9159), .Z(n8937) );
  XOR2_X1 U9110 ( .A(n9160), .B(n9161), .Z(n9159) );
  NAND2_X1 U9111 ( .A1(b_27_), .A2(a_24_), .ZN(n9161) );
  XNOR2_X1 U9112 ( .A(n9162), .B(n9163), .ZN(n8941) );
  XNOR2_X1 U9113 ( .A(n9164), .B(n9165), .ZN(n9162) );
  XNOR2_X1 U9114 ( .A(n9166), .B(n9167), .ZN(n8945) );
  XOR2_X1 U9115 ( .A(n9168), .B(n9169), .Z(n9166) );
  NOR2_X1 U9116 ( .A1(n7645), .A2(n7564), .ZN(n9169) );
  XNOR2_X1 U9117 ( .A(n9170), .B(n9171), .ZN(n8949) );
  XNOR2_X1 U9118 ( .A(n9172), .B(n9173), .ZN(n9171) );
  XNOR2_X1 U9119 ( .A(n9174), .B(n9175), .ZN(n8953) );
  XOR2_X1 U9120 ( .A(n9176), .B(n9177), .Z(n9174) );
  NOR2_X1 U9121 ( .A1(n7676), .A2(n7564), .ZN(n9177) );
  XNOR2_X1 U9122 ( .A(n9178), .B(n9179), .ZN(n8957) );
  XNOR2_X1 U9123 ( .A(n9180), .B(n9181), .ZN(n9178) );
  XNOR2_X1 U9124 ( .A(n9182), .B(n9183), .ZN(n8961) );
  XOR2_X1 U9125 ( .A(n9184), .B(n9185), .Z(n9182) );
  NOR2_X1 U9126 ( .A1(n7707), .A2(n7564), .ZN(n9185) );
  XNOR2_X1 U9127 ( .A(n9186), .B(n9187), .ZN(n8965) );
  XNOR2_X1 U9128 ( .A(n9188), .B(n9189), .ZN(n9186) );
  XOR2_X1 U9129 ( .A(n9190), .B(n9191), .Z(n8969) );
  XOR2_X1 U9130 ( .A(n9192), .B(n9193), .Z(n9191) );
  NAND2_X1 U9131 ( .A1(b_27_), .A2(a_16_), .ZN(n9193) );
  XOR2_X1 U9132 ( .A(n9194), .B(n9195), .Z(n8972) );
  XOR2_X1 U9133 ( .A(n9196), .B(n9197), .Z(n9194) );
  XNOR2_X1 U9134 ( .A(n9198), .B(n9199), .ZN(n8977) );
  XOR2_X1 U9135 ( .A(n9200), .B(n9201), .Z(n9198) );
  NOR2_X1 U9136 ( .A1(n7775), .A2(n7564), .ZN(n9201) );
  XNOR2_X1 U9137 ( .A(n9202), .B(n9203), .ZN(n8981) );
  XNOR2_X1 U9138 ( .A(n9204), .B(n9205), .ZN(n9203) );
  XOR2_X1 U9139 ( .A(n9206), .B(n9207), .Z(n8985) );
  XOR2_X1 U9140 ( .A(n9208), .B(n9209), .Z(n9206) );
  NOR2_X1 U9141 ( .A1(n7806), .A2(n7564), .ZN(n9209) );
  XOR2_X1 U9142 ( .A(n9210), .B(n9211), .Z(n8988) );
  XOR2_X1 U9143 ( .A(n9212), .B(n9213), .Z(n9210) );
  XNOR2_X1 U9144 ( .A(n9214), .B(n9215), .ZN(n8993) );
  XOR2_X1 U9145 ( .A(n9216), .B(n9217), .Z(n9215) );
  NAND2_X1 U9146 ( .A1(b_27_), .A2(a_10_), .ZN(n9217) );
  XOR2_X1 U9147 ( .A(n9218), .B(n9219), .Z(n8996) );
  XOR2_X1 U9148 ( .A(n9220), .B(n9221), .Z(n9218) );
  XNOR2_X1 U9149 ( .A(n9222), .B(n9223), .ZN(n9001) );
  XOR2_X1 U9150 ( .A(n9224), .B(n9225), .Z(n9222) );
  NOR2_X1 U9151 ( .A1(n8059), .A2(n7564), .ZN(n9225) );
  XOR2_X1 U9152 ( .A(n9226), .B(n9227), .Z(n9005) );
  XOR2_X1 U9153 ( .A(n9228), .B(n9229), .Z(n9226) );
  NOR2_X1 U9154 ( .A1(n7884), .A2(n7564), .ZN(n9229) );
  XOR2_X1 U9155 ( .A(n9230), .B(n9231), .Z(n9008) );
  XOR2_X1 U9156 ( .A(n9232), .B(n9233), .Z(n9230) );
  NOR2_X1 U9157 ( .A1(n8061), .A2(n7564), .ZN(n9233) );
  XOR2_X1 U9158 ( .A(n9234), .B(n9235), .Z(n9012) );
  XOR2_X1 U9159 ( .A(n9236), .B(n9237), .Z(n9234) );
  XOR2_X1 U9160 ( .A(n9238), .B(n9239), .Z(n9017) );
  XOR2_X1 U9161 ( .A(n9240), .B(n9241), .Z(n9238) );
  OR2_X1 U9162 ( .A1(n9023), .A2(n9021), .ZN(n9032) );
  XNOR2_X1 U9163 ( .A(n9242), .B(n9243), .ZN(n9021) );
  XOR2_X1 U9164 ( .A(n9244), .B(n9245), .Z(n9242) );
  NOR2_X1 U9165 ( .A1(n7945), .A2(n7564), .ZN(n9245) );
  NAND2_X1 U9166 ( .A1(b_28_), .A2(a_2_), .ZN(n9023) );
  XNOR2_X1 U9167 ( .A(n9246), .B(n9247), .ZN(n8800) );
  NAND2_X1 U9168 ( .A1(n9248), .A2(n9249), .ZN(n9246) );
  XOR2_X1 U9169 ( .A(n9250), .B(n9251), .Z(n8791) );
  XOR2_X1 U9170 ( .A(n9252), .B(n9253), .Z(n9250) );
  NOR2_X1 U9171 ( .A1(n7973), .A2(n7564), .ZN(n9253) );
  NOR2_X1 U9172 ( .A1(n9254), .A2(n8288), .ZN(n9024) );
  XNOR2_X1 U9173 ( .A(n9255), .B(n9256), .ZN(n8288) );
  XNOR2_X1 U9174 ( .A(n9257), .B(n9258), .ZN(n9256) );
  AND2_X1 U9175 ( .A1(n8287), .A2(n8286), .ZN(n9254) );
  NAND2_X1 U9176 ( .A1(n9259), .A2(n8285), .ZN(n8101) );
  NOR2_X1 U9177 ( .A1(n8287), .A2(n8286), .ZN(n8285) );
  XOR2_X1 U9178 ( .A(n9260), .B(n9261), .Z(n8286) );
  XNOR2_X1 U9179 ( .A(n9262), .B(n9263), .ZN(n9261) );
  NAND2_X1 U9180 ( .A1(n9264), .A2(n9265), .ZN(n8287) );
  NAND2_X1 U9181 ( .A1(n9257), .A2(n9266), .ZN(n9265) );
  OR2_X1 U9182 ( .A1(n9258), .A2(n9255), .ZN(n9266) );
  AND2_X1 U9183 ( .A1(n9267), .A2(n9268), .ZN(n9257) );
  NAND2_X1 U9184 ( .A1(n9269), .A2(b_27_), .ZN(n9268) );
  NOR2_X1 U9185 ( .A1(n9270), .A2(n7973), .ZN(n9269) );
  NOR2_X1 U9186 ( .A1(n9251), .A2(n9252), .ZN(n9270) );
  NAND2_X1 U9187 ( .A1(n9251), .A2(n9252), .ZN(n9267) );
  NAND2_X1 U9188 ( .A1(n9248), .A2(n9271), .ZN(n9252) );
  NAND2_X1 U9189 ( .A1(n9247), .A2(n9249), .ZN(n9271) );
  NAND2_X1 U9190 ( .A1(n9272), .A2(n9273), .ZN(n9249) );
  NAND2_X1 U9191 ( .A1(b_27_), .A2(a_2_), .ZN(n9273) );
  INV_X1 U9192 ( .A(n9274), .ZN(n9272) );
  XNOR2_X1 U9193 ( .A(n9275), .B(n9276), .ZN(n9247) );
  XNOR2_X1 U9194 ( .A(n9277), .B(n9278), .ZN(n9276) );
  NAND2_X1 U9195 ( .A1(a_2_), .A2(n9274), .ZN(n9248) );
  NAND2_X1 U9196 ( .A1(n9279), .A2(n9280), .ZN(n9274) );
  NAND2_X1 U9197 ( .A1(n9281), .A2(b_27_), .ZN(n9280) );
  NOR2_X1 U9198 ( .A1(n9282), .A2(n7945), .ZN(n9281) );
  NOR2_X1 U9199 ( .A1(n9243), .A2(n9244), .ZN(n9282) );
  NAND2_X1 U9200 ( .A1(n9243), .A2(n9244), .ZN(n9279) );
  NAND2_X1 U9201 ( .A1(n9283), .A2(n9284), .ZN(n9244) );
  NAND2_X1 U9202 ( .A1(n9241), .A2(n9285), .ZN(n9284) );
  OR2_X1 U9203 ( .A1(n9240), .A2(n9239), .ZN(n9285) );
  NOR2_X1 U9204 ( .A1(n7564), .A2(n7934), .ZN(n9241) );
  NAND2_X1 U9205 ( .A1(n9239), .A2(n9240), .ZN(n9283) );
  NAND2_X1 U9206 ( .A1(n9286), .A2(n9287), .ZN(n9240) );
  NAND2_X1 U9207 ( .A1(n9237), .A2(n9288), .ZN(n9287) );
  OR2_X1 U9208 ( .A1(n9236), .A2(n9235), .ZN(n9288) );
  NOR2_X1 U9209 ( .A1(n7564), .A2(n7914), .ZN(n9237) );
  NAND2_X1 U9210 ( .A1(n9235), .A2(n9236), .ZN(n9286) );
  NAND2_X1 U9211 ( .A1(n9289), .A2(n9290), .ZN(n9236) );
  NAND2_X1 U9212 ( .A1(n9291), .A2(b_27_), .ZN(n9290) );
  NOR2_X1 U9213 ( .A1(n9292), .A2(n8061), .ZN(n9291) );
  NOR2_X1 U9214 ( .A1(n9231), .A2(n9232), .ZN(n9292) );
  NAND2_X1 U9215 ( .A1(n9231), .A2(n9232), .ZN(n9289) );
  NAND2_X1 U9216 ( .A1(n9293), .A2(n9294), .ZN(n9232) );
  NAND2_X1 U9217 ( .A1(n9295), .A2(b_27_), .ZN(n9294) );
  NOR2_X1 U9218 ( .A1(n9296), .A2(n7884), .ZN(n9295) );
  NOR2_X1 U9219 ( .A1(n9227), .A2(n9228), .ZN(n9296) );
  NAND2_X1 U9220 ( .A1(n9227), .A2(n9228), .ZN(n9293) );
  NAND2_X1 U9221 ( .A1(n9297), .A2(n9298), .ZN(n9228) );
  NAND2_X1 U9222 ( .A1(n9299), .A2(b_27_), .ZN(n9298) );
  NOR2_X1 U9223 ( .A1(n9300), .A2(n8059), .ZN(n9299) );
  NOR2_X1 U9224 ( .A1(n9223), .A2(n9224), .ZN(n9300) );
  NAND2_X1 U9225 ( .A1(n9223), .A2(n9224), .ZN(n9297) );
  NAND2_X1 U9226 ( .A1(n9301), .A2(n9302), .ZN(n9224) );
  NAND2_X1 U9227 ( .A1(n9221), .A2(n9303), .ZN(n9302) );
  OR2_X1 U9228 ( .A1(n9220), .A2(n9219), .ZN(n9303) );
  NOR2_X1 U9229 ( .A1(n7564), .A2(n7848), .ZN(n9221) );
  NAND2_X1 U9230 ( .A1(n9219), .A2(n9220), .ZN(n9301) );
  NAND2_X1 U9231 ( .A1(n9304), .A2(n9305), .ZN(n9220) );
  NAND2_X1 U9232 ( .A1(n9306), .A2(b_27_), .ZN(n9305) );
  NOR2_X1 U9233 ( .A1(n9307), .A2(n7837), .ZN(n9306) );
  NOR2_X1 U9234 ( .A1(n9214), .A2(n9216), .ZN(n9307) );
  NAND2_X1 U9235 ( .A1(n9214), .A2(n9216), .ZN(n9304) );
  NAND2_X1 U9236 ( .A1(n9308), .A2(n9309), .ZN(n9216) );
  NAND2_X1 U9237 ( .A1(n9213), .A2(n9310), .ZN(n9309) );
  OR2_X1 U9238 ( .A1(n9212), .A2(n9211), .ZN(n9310) );
  NOR2_X1 U9239 ( .A1(n7564), .A2(n7817), .ZN(n9213) );
  NAND2_X1 U9240 ( .A1(n9211), .A2(n9212), .ZN(n9308) );
  NAND2_X1 U9241 ( .A1(n9311), .A2(n9312), .ZN(n9212) );
  NAND2_X1 U9242 ( .A1(n9313), .A2(b_27_), .ZN(n9312) );
  NOR2_X1 U9243 ( .A1(n9314), .A2(n7806), .ZN(n9313) );
  NOR2_X1 U9244 ( .A1(n9207), .A2(n9208), .ZN(n9314) );
  NAND2_X1 U9245 ( .A1(n9207), .A2(n9208), .ZN(n9311) );
  NAND2_X1 U9246 ( .A1(n9315), .A2(n9316), .ZN(n9208) );
  NAND2_X1 U9247 ( .A1(n9205), .A2(n9317), .ZN(n9316) );
  OR2_X1 U9248 ( .A1(n9204), .A2(n9202), .ZN(n9317) );
  NOR2_X1 U9249 ( .A1(n7564), .A2(n7786), .ZN(n9205) );
  NAND2_X1 U9250 ( .A1(n9202), .A2(n9204), .ZN(n9315) );
  NAND2_X1 U9251 ( .A1(n9318), .A2(n9319), .ZN(n9204) );
  NAND2_X1 U9252 ( .A1(n9320), .A2(b_27_), .ZN(n9319) );
  NOR2_X1 U9253 ( .A1(n9321), .A2(n7775), .ZN(n9320) );
  NOR2_X1 U9254 ( .A1(n9199), .A2(n9200), .ZN(n9321) );
  NAND2_X1 U9255 ( .A1(n9199), .A2(n9200), .ZN(n9318) );
  NAND2_X1 U9256 ( .A1(n9322), .A2(n9323), .ZN(n9200) );
  NAND2_X1 U9257 ( .A1(n9197), .A2(n9324), .ZN(n9323) );
  OR2_X1 U9258 ( .A1(n9196), .A2(n9195), .ZN(n9324) );
  NOR2_X1 U9259 ( .A1(n7564), .A2(n7754), .ZN(n9197) );
  NAND2_X1 U9260 ( .A1(n9195), .A2(n9196), .ZN(n9322) );
  NAND2_X1 U9261 ( .A1(n9325), .A2(n9326), .ZN(n9196) );
  NAND2_X1 U9262 ( .A1(n9327), .A2(b_27_), .ZN(n9326) );
  NOR2_X1 U9263 ( .A1(n9328), .A2(n7743), .ZN(n9327) );
  NOR2_X1 U9264 ( .A1(n9190), .A2(n9192), .ZN(n9328) );
  NAND2_X1 U9265 ( .A1(n9190), .A2(n9192), .ZN(n9325) );
  NAND2_X1 U9266 ( .A1(n9329), .A2(n9330), .ZN(n9192) );
  NAND2_X1 U9267 ( .A1(n9189), .A2(n9331), .ZN(n9330) );
  NAND2_X1 U9268 ( .A1(n9188), .A2(n9187), .ZN(n9331) );
  NOR2_X1 U9269 ( .A1(n7564), .A2(n7723), .ZN(n9189) );
  OR2_X1 U9270 ( .A1(n9187), .A2(n9188), .ZN(n9329) );
  AND2_X1 U9271 ( .A1(n9332), .A2(n9333), .ZN(n9188) );
  NAND2_X1 U9272 ( .A1(n9334), .A2(b_27_), .ZN(n9333) );
  NOR2_X1 U9273 ( .A1(n9335), .A2(n7707), .ZN(n9334) );
  NOR2_X1 U9274 ( .A1(n9183), .A2(n9184), .ZN(n9335) );
  NAND2_X1 U9275 ( .A1(n9183), .A2(n9184), .ZN(n9332) );
  NAND2_X1 U9276 ( .A1(n9336), .A2(n9337), .ZN(n9184) );
  NAND2_X1 U9277 ( .A1(n9181), .A2(n9338), .ZN(n9337) );
  NAND2_X1 U9278 ( .A1(n9180), .A2(n9179), .ZN(n9338) );
  NOR2_X1 U9279 ( .A1(n7564), .A2(n7687), .ZN(n9181) );
  OR2_X1 U9280 ( .A1(n9179), .A2(n9180), .ZN(n9336) );
  AND2_X1 U9281 ( .A1(n9339), .A2(n9340), .ZN(n9180) );
  NAND2_X1 U9282 ( .A1(n9341), .A2(b_27_), .ZN(n9340) );
  NOR2_X1 U9283 ( .A1(n9342), .A2(n7676), .ZN(n9341) );
  NOR2_X1 U9284 ( .A1(n9175), .A2(n9176), .ZN(n9342) );
  NAND2_X1 U9285 ( .A1(n9175), .A2(n9176), .ZN(n9339) );
  NAND2_X1 U9286 ( .A1(n9343), .A2(n9344), .ZN(n9176) );
  NAND2_X1 U9287 ( .A1(n9173), .A2(n9345), .ZN(n9344) );
  OR2_X1 U9288 ( .A1(n9172), .A2(n9170), .ZN(n9345) );
  NOR2_X1 U9289 ( .A1(n7564), .A2(n7656), .ZN(n9173) );
  NAND2_X1 U9290 ( .A1(n9170), .A2(n9172), .ZN(n9343) );
  NAND2_X1 U9291 ( .A1(n9346), .A2(n9347), .ZN(n9172) );
  NAND2_X1 U9292 ( .A1(n9348), .A2(b_27_), .ZN(n9347) );
  NOR2_X1 U9293 ( .A1(n9349), .A2(n7645), .ZN(n9348) );
  NOR2_X1 U9294 ( .A1(n9167), .A2(n9168), .ZN(n9349) );
  NAND2_X1 U9295 ( .A1(n9167), .A2(n9168), .ZN(n9346) );
  NAND2_X1 U9296 ( .A1(n9350), .A2(n9351), .ZN(n9168) );
  NAND2_X1 U9297 ( .A1(n9165), .A2(n9352), .ZN(n9351) );
  NAND2_X1 U9298 ( .A1(n9164), .A2(n9163), .ZN(n9352) );
  NOR2_X1 U9299 ( .A1(n7564), .A2(n7624), .ZN(n9165) );
  OR2_X1 U9300 ( .A1(n9163), .A2(n9164), .ZN(n9350) );
  AND2_X1 U9301 ( .A1(n9353), .A2(n9354), .ZN(n9164) );
  NAND2_X1 U9302 ( .A1(n9355), .A2(b_27_), .ZN(n9354) );
  NOR2_X1 U9303 ( .A1(n9356), .A2(n7613), .ZN(n9355) );
  NOR2_X1 U9304 ( .A1(n9158), .A2(n9160), .ZN(n9356) );
  NAND2_X1 U9305 ( .A1(n9158), .A2(n9160), .ZN(n9353) );
  NAND2_X1 U9306 ( .A1(n9357), .A2(n9358), .ZN(n9160) );
  NAND2_X1 U9307 ( .A1(n9157), .A2(n9359), .ZN(n9358) );
  NAND2_X1 U9308 ( .A1(n9156), .A2(n9155), .ZN(n9359) );
  NOR2_X1 U9309 ( .A1(n7564), .A2(n7593), .ZN(n9157) );
  OR2_X1 U9310 ( .A1(n9155), .A2(n9156), .ZN(n9357) );
  AND2_X1 U9311 ( .A1(n9360), .A2(n9361), .ZN(n9156) );
  NAND2_X1 U9312 ( .A1(n9362), .A2(b_27_), .ZN(n9361) );
  NOR2_X1 U9313 ( .A1(n9363), .A2(n8052), .ZN(n9362) );
  NOR2_X1 U9314 ( .A1(n9151), .A2(n9153), .ZN(n9363) );
  NAND2_X1 U9315 ( .A1(n9151), .A2(n9153), .ZN(n9360) );
  NAND2_X1 U9316 ( .A1(n9364), .A2(n9365), .ZN(n9153) );
  NAND2_X1 U9317 ( .A1(n7558), .A2(n9366), .ZN(n9365) );
  NAND2_X1 U9318 ( .A1(n9149), .A2(n9148), .ZN(n9366) );
  INV_X1 U9319 ( .A(n8038), .ZN(n7558) );
  NAND2_X1 U9320 ( .A1(b_27_), .A2(a_27_), .ZN(n8038) );
  OR2_X1 U9321 ( .A1(n9148), .A2(n9149), .ZN(n9364) );
  AND2_X1 U9322 ( .A1(n9145), .A2(n9367), .ZN(n9149) );
  NAND2_X1 U9323 ( .A1(n9144), .A2(n9146), .ZN(n9367) );
  NAND2_X1 U9324 ( .A1(n9368), .A2(n9369), .ZN(n9146) );
  NAND2_X1 U9325 ( .A1(b_27_), .A2(a_28_), .ZN(n9369) );
  INV_X1 U9326 ( .A(n9370), .ZN(n9368) );
  XOR2_X1 U9327 ( .A(n9371), .B(n9372), .Z(n9144) );
  NOR2_X1 U9328 ( .A1(n7529), .A2(n8051), .ZN(n9372) );
  XOR2_X1 U9329 ( .A(n9373), .B(n9374), .Z(n9371) );
  NAND2_X1 U9330 ( .A1(a_28_), .A2(n9370), .ZN(n9145) );
  NAND2_X1 U9331 ( .A1(n9375), .A2(n9376), .ZN(n9370) );
  NAND2_X1 U9332 ( .A1(n9377), .A2(b_27_), .ZN(n9376) );
  NOR2_X1 U9333 ( .A1(n9378), .A2(n7529), .ZN(n9377) );
  NOR2_X1 U9334 ( .A1(n9129), .A2(n9130), .ZN(n9378) );
  NAND2_X1 U9335 ( .A1(n9129), .A2(n9130), .ZN(n9375) );
  NAND2_X1 U9336 ( .A1(n9379), .A2(n9380), .ZN(n9130) );
  NAND2_X1 U9337 ( .A1(n9381), .A2(b_25_), .ZN(n9380) );
  NOR2_X1 U9338 ( .A1(n9382), .A2(n8048), .ZN(n9381) );
  NOR2_X1 U9339 ( .A1(n8676), .A2(n8051), .ZN(n9382) );
  NAND2_X1 U9340 ( .A1(n9383), .A2(b_26_), .ZN(n9379) );
  NOR2_X1 U9341 ( .A1(n9384), .A2(n7515), .ZN(n9383) );
  NOR2_X1 U9342 ( .A1(n8679), .A2(n7594), .ZN(n9384) );
  AND2_X1 U9343 ( .A1(n9142), .A2(b_26_), .ZN(n9129) );
  NOR2_X1 U9344 ( .A1(n8451), .A2(n7564), .ZN(n9142) );
  XOR2_X1 U9345 ( .A(n9385), .B(n9386), .Z(n9148) );
  NAND2_X1 U9346 ( .A1(n9387), .A2(n9388), .ZN(n9385) );
  XNOR2_X1 U9347 ( .A(n9389), .B(n9390), .ZN(n9151) );
  XNOR2_X1 U9348 ( .A(n9391), .B(n9392), .ZN(n9389) );
  XNOR2_X1 U9349 ( .A(n9393), .B(n9394), .ZN(n9155) );
  XOR2_X1 U9350 ( .A(n7577), .B(n9395), .Z(n9393) );
  XNOR2_X1 U9351 ( .A(n9396), .B(n9397), .ZN(n9158) );
  XNOR2_X1 U9352 ( .A(n9398), .B(n9399), .ZN(n9396) );
  XOR2_X1 U9353 ( .A(n9400), .B(n9401), .Z(n9163) );
  XOR2_X1 U9354 ( .A(n9402), .B(n9403), .Z(n9401) );
  NAND2_X1 U9355 ( .A1(b_26_), .A2(a_24_), .ZN(n9403) );
  XNOR2_X1 U9356 ( .A(n9404), .B(n9405), .ZN(n9167) );
  XNOR2_X1 U9357 ( .A(n9406), .B(n9407), .ZN(n9404) );
  XOR2_X1 U9358 ( .A(n9408), .B(n9409), .Z(n9170) );
  XOR2_X1 U9359 ( .A(n9410), .B(n9411), .Z(n9408) );
  NOR2_X1 U9360 ( .A1(n7645), .A2(n8051), .ZN(n9411) );
  XNOR2_X1 U9361 ( .A(n9412), .B(n9413), .ZN(n9175) );
  XNOR2_X1 U9362 ( .A(n9414), .B(n9415), .ZN(n9413) );
  XNOR2_X1 U9363 ( .A(n9416), .B(n9417), .ZN(n9179) );
  XOR2_X1 U9364 ( .A(n9418), .B(n9419), .Z(n9416) );
  NOR2_X1 U9365 ( .A1(n7676), .A2(n8051), .ZN(n9419) );
  XNOR2_X1 U9366 ( .A(n9420), .B(n9421), .ZN(n9183) );
  XNOR2_X1 U9367 ( .A(n9422), .B(n9423), .ZN(n9420) );
  XOR2_X1 U9368 ( .A(n9424), .B(n9425), .Z(n9187) );
  XOR2_X1 U9369 ( .A(n9426), .B(n9427), .Z(n9425) );
  NAND2_X1 U9370 ( .A1(b_26_), .A2(a_18_), .ZN(n9427) );
  XNOR2_X1 U9371 ( .A(n9428), .B(n9429), .ZN(n9190) );
  XNOR2_X1 U9372 ( .A(n9430), .B(n9431), .ZN(n9428) );
  XOR2_X1 U9373 ( .A(n9432), .B(n9433), .Z(n9195) );
  XOR2_X1 U9374 ( .A(n9434), .B(n9435), .Z(n9432) );
  NOR2_X1 U9375 ( .A1(n7743), .A2(n8051), .ZN(n9435) );
  XNOR2_X1 U9376 ( .A(n9436), .B(n9437), .ZN(n9199) );
  XNOR2_X1 U9377 ( .A(n9438), .B(n9439), .ZN(n9436) );
  XOR2_X1 U9378 ( .A(n9440), .B(n9441), .Z(n9202) );
  XOR2_X1 U9379 ( .A(n9442), .B(n9443), .Z(n9440) );
  NOR2_X1 U9380 ( .A1(n7775), .A2(n8051), .ZN(n9443) );
  XOR2_X1 U9381 ( .A(n9444), .B(n9445), .Z(n9207) );
  XOR2_X1 U9382 ( .A(n9446), .B(n9447), .Z(n9444) );
  XNOR2_X1 U9383 ( .A(n9448), .B(n9449), .ZN(n9211) );
  XOR2_X1 U9384 ( .A(n9450), .B(n9451), .Z(n9449) );
  NAND2_X1 U9385 ( .A1(b_26_), .A2(a_12_), .ZN(n9451) );
  XOR2_X1 U9386 ( .A(n9452), .B(n9453), .Z(n9214) );
  XOR2_X1 U9387 ( .A(n9454), .B(n9455), .Z(n9452) );
  XOR2_X1 U9388 ( .A(n9456), .B(n9457), .Z(n9219) );
  XOR2_X1 U9389 ( .A(n9458), .B(n9459), .Z(n9456) );
  NOR2_X1 U9390 ( .A1(n7837), .A2(n8051), .ZN(n9459) );
  XNOR2_X1 U9391 ( .A(n9460), .B(n9461), .ZN(n9223) );
  XNOR2_X1 U9392 ( .A(n9462), .B(n9463), .ZN(n9460) );
  XOR2_X1 U9393 ( .A(n9464), .B(n9465), .Z(n9227) );
  XOR2_X1 U9394 ( .A(n9466), .B(n9467), .Z(n9464) );
  NOR2_X1 U9395 ( .A1(n8059), .A2(n8051), .ZN(n9467) );
  XNOR2_X1 U9396 ( .A(n9468), .B(n9469), .ZN(n9231) );
  NAND2_X1 U9397 ( .A1(n9470), .A2(n9471), .ZN(n9468) );
  XNOR2_X1 U9398 ( .A(n9472), .B(n9473), .ZN(n9235) );
  NAND2_X1 U9399 ( .A1(n9474), .A2(n9475), .ZN(n9472) );
  XOR2_X1 U9400 ( .A(n9476), .B(n9477), .Z(n9239) );
  XOR2_X1 U9401 ( .A(n9478), .B(n9479), .Z(n9476) );
  NOR2_X1 U9402 ( .A1(n7914), .A2(n8051), .ZN(n9479) );
  XNOR2_X1 U9403 ( .A(n9480), .B(n9481), .ZN(n9243) );
  XNOR2_X1 U9404 ( .A(n9482), .B(n9483), .ZN(n9481) );
  XNOR2_X1 U9405 ( .A(n9484), .B(n9485), .ZN(n9251) );
  NAND2_X1 U9406 ( .A1(n9486), .A2(n9487), .ZN(n9484) );
  NAND2_X1 U9407 ( .A1(n9255), .A2(n9258), .ZN(n9264) );
  NAND2_X1 U9408 ( .A1(b_27_), .A2(a_0_), .ZN(n9258) );
  XNOR2_X1 U9409 ( .A(n9488), .B(n9489), .ZN(n9255) );
  XOR2_X1 U9410 ( .A(n9490), .B(n9491), .Z(n9488) );
  NOR2_X1 U9411 ( .A1(n7973), .A2(n8051), .ZN(n9491) );
  NOR2_X1 U9412 ( .A1(n9492), .A2(n9493), .ZN(n9259) );
  NOR2_X1 U9413 ( .A1(n8279), .A2(n8280), .ZN(n9493) );
  NAND2_X1 U9414 ( .A1(n9494), .A2(n9495), .ZN(n8106) );
  NAND2_X1 U9415 ( .A1(n9496), .A2(n8274), .ZN(n9495) );
  NAND2_X1 U9416 ( .A1(n9497), .A2(n9492), .ZN(n8107) );
  INV_X1 U9417 ( .A(n9494), .ZN(n9492) );
  NAND2_X1 U9418 ( .A1(n8279), .A2(n8280), .ZN(n9494) );
  NAND2_X1 U9419 ( .A1(n9498), .A2(n9499), .ZN(n8280) );
  NAND2_X1 U9420 ( .A1(n9263), .A2(n9500), .ZN(n9499) );
  OR2_X1 U9421 ( .A1(n9262), .A2(n9260), .ZN(n9500) );
  NOR2_X1 U9422 ( .A1(n8051), .A2(n8307), .ZN(n9263) );
  NAND2_X1 U9423 ( .A1(n9260), .A2(n9262), .ZN(n9498) );
  NAND2_X1 U9424 ( .A1(n9501), .A2(n9502), .ZN(n9262) );
  NAND2_X1 U9425 ( .A1(n9503), .A2(b_26_), .ZN(n9502) );
  NOR2_X1 U9426 ( .A1(n9504), .A2(n7973), .ZN(n9503) );
  NOR2_X1 U9427 ( .A1(n9489), .A2(n9490), .ZN(n9504) );
  NAND2_X1 U9428 ( .A1(n9489), .A2(n9490), .ZN(n9501) );
  NAND2_X1 U9429 ( .A1(n9486), .A2(n9505), .ZN(n9490) );
  NAND2_X1 U9430 ( .A1(n9485), .A2(n9487), .ZN(n9505) );
  NAND2_X1 U9431 ( .A1(n9506), .A2(n9507), .ZN(n9487) );
  NAND2_X1 U9432 ( .A1(b_26_), .A2(a_2_), .ZN(n9507) );
  INV_X1 U9433 ( .A(n9508), .ZN(n9506) );
  XOR2_X1 U9434 ( .A(n9509), .B(n9510), .Z(n9485) );
  XOR2_X1 U9435 ( .A(n9511), .B(n9512), .Z(n9509) );
  NOR2_X1 U9436 ( .A1(n7945), .A2(n7594), .ZN(n9512) );
  NAND2_X1 U9437 ( .A1(a_2_), .A2(n9508), .ZN(n9486) );
  NAND2_X1 U9438 ( .A1(n9513), .A2(n9514), .ZN(n9508) );
  NAND2_X1 U9439 ( .A1(n9278), .A2(n9515), .ZN(n9514) );
  OR2_X1 U9440 ( .A1(n9277), .A2(n9275), .ZN(n9515) );
  NOR2_X1 U9441 ( .A1(n8051), .A2(n7945), .ZN(n9278) );
  NAND2_X1 U9442 ( .A1(n9275), .A2(n9277), .ZN(n9513) );
  NAND2_X1 U9443 ( .A1(n9516), .A2(n9517), .ZN(n9277) );
  NAND2_X1 U9444 ( .A1(n9483), .A2(n9518), .ZN(n9517) );
  OR2_X1 U9445 ( .A1(n9482), .A2(n9480), .ZN(n9518) );
  NOR2_X1 U9446 ( .A1(n8051), .A2(n7934), .ZN(n9483) );
  NAND2_X1 U9447 ( .A1(n9480), .A2(n9482), .ZN(n9516) );
  NAND2_X1 U9448 ( .A1(n9519), .A2(n9520), .ZN(n9482) );
  NAND2_X1 U9449 ( .A1(n9521), .A2(b_26_), .ZN(n9520) );
  NOR2_X1 U9450 ( .A1(n9522), .A2(n7914), .ZN(n9521) );
  NOR2_X1 U9451 ( .A1(n9477), .A2(n9478), .ZN(n9522) );
  NAND2_X1 U9452 ( .A1(n9477), .A2(n9478), .ZN(n9519) );
  NAND2_X1 U9453 ( .A1(n9474), .A2(n9523), .ZN(n9478) );
  NAND2_X1 U9454 ( .A1(n9473), .A2(n9475), .ZN(n9523) );
  NAND2_X1 U9455 ( .A1(n9524), .A2(n9525), .ZN(n9475) );
  NAND2_X1 U9456 ( .A1(b_26_), .A2(a_6_), .ZN(n9525) );
  INV_X1 U9457 ( .A(n9526), .ZN(n9524) );
  XNOR2_X1 U9458 ( .A(n9527), .B(n9528), .ZN(n9473) );
  NAND2_X1 U9459 ( .A1(n9529), .A2(n9530), .ZN(n9527) );
  NAND2_X1 U9460 ( .A1(a_6_), .A2(n9526), .ZN(n9474) );
  NAND2_X1 U9461 ( .A1(n9470), .A2(n9531), .ZN(n9526) );
  NAND2_X1 U9462 ( .A1(n9469), .A2(n9471), .ZN(n9531) );
  NAND2_X1 U9463 ( .A1(n9532), .A2(n9533), .ZN(n9471) );
  NAND2_X1 U9464 ( .A1(b_26_), .A2(a_7_), .ZN(n9533) );
  INV_X1 U9465 ( .A(n9534), .ZN(n9532) );
  XNOR2_X1 U9466 ( .A(n9535), .B(n9536), .ZN(n9469) );
  XOR2_X1 U9467 ( .A(n9537), .B(n9538), .Z(n9536) );
  NAND2_X1 U9468 ( .A1(b_25_), .A2(a_8_), .ZN(n9538) );
  NAND2_X1 U9469 ( .A1(a_7_), .A2(n9534), .ZN(n9470) );
  NAND2_X1 U9470 ( .A1(n9539), .A2(n9540), .ZN(n9534) );
  NAND2_X1 U9471 ( .A1(n9541), .A2(b_26_), .ZN(n9540) );
  NOR2_X1 U9472 ( .A1(n9542), .A2(n8059), .ZN(n9541) );
  NOR2_X1 U9473 ( .A1(n9466), .A2(n9465), .ZN(n9542) );
  NAND2_X1 U9474 ( .A1(n9465), .A2(n9466), .ZN(n9539) );
  NAND2_X1 U9475 ( .A1(n9543), .A2(n9544), .ZN(n9466) );
  NAND2_X1 U9476 ( .A1(n9463), .A2(n9545), .ZN(n9544) );
  NAND2_X1 U9477 ( .A1(n9462), .A2(n9461), .ZN(n9545) );
  NOR2_X1 U9478 ( .A1(n8051), .A2(n7848), .ZN(n9463) );
  OR2_X1 U9479 ( .A1(n9461), .A2(n9462), .ZN(n9543) );
  AND2_X1 U9480 ( .A1(n9546), .A2(n9547), .ZN(n9462) );
  NAND2_X1 U9481 ( .A1(n9548), .A2(b_26_), .ZN(n9547) );
  NOR2_X1 U9482 ( .A1(n9549), .A2(n7837), .ZN(n9548) );
  NOR2_X1 U9483 ( .A1(n9457), .A2(n9458), .ZN(n9549) );
  NAND2_X1 U9484 ( .A1(n9457), .A2(n9458), .ZN(n9546) );
  NAND2_X1 U9485 ( .A1(n9550), .A2(n9551), .ZN(n9458) );
  NAND2_X1 U9486 ( .A1(n9455), .A2(n9552), .ZN(n9551) );
  OR2_X1 U9487 ( .A1(n9453), .A2(n9454), .ZN(n9552) );
  NOR2_X1 U9488 ( .A1(n8051), .A2(n7817), .ZN(n9455) );
  NAND2_X1 U9489 ( .A1(n9453), .A2(n9454), .ZN(n9550) );
  NAND2_X1 U9490 ( .A1(n9553), .A2(n9554), .ZN(n9454) );
  NAND2_X1 U9491 ( .A1(n9555), .A2(b_26_), .ZN(n9554) );
  NOR2_X1 U9492 ( .A1(n9556), .A2(n7806), .ZN(n9555) );
  NOR2_X1 U9493 ( .A1(n9448), .A2(n9450), .ZN(n9556) );
  NAND2_X1 U9494 ( .A1(n9448), .A2(n9450), .ZN(n9553) );
  NAND2_X1 U9495 ( .A1(n9557), .A2(n9558), .ZN(n9450) );
  NAND2_X1 U9496 ( .A1(n9447), .A2(n9559), .ZN(n9558) );
  OR2_X1 U9497 ( .A1(n9445), .A2(n9446), .ZN(n9559) );
  NOR2_X1 U9498 ( .A1(n8051), .A2(n7786), .ZN(n9447) );
  NAND2_X1 U9499 ( .A1(n9445), .A2(n9446), .ZN(n9557) );
  NAND2_X1 U9500 ( .A1(n9560), .A2(n9561), .ZN(n9446) );
  NAND2_X1 U9501 ( .A1(n9562), .A2(b_26_), .ZN(n9561) );
  NOR2_X1 U9502 ( .A1(n9563), .A2(n7775), .ZN(n9562) );
  NOR2_X1 U9503 ( .A1(n9442), .A2(n9441), .ZN(n9563) );
  NAND2_X1 U9504 ( .A1(n9441), .A2(n9442), .ZN(n9560) );
  NAND2_X1 U9505 ( .A1(n9564), .A2(n9565), .ZN(n9442) );
  NAND2_X1 U9506 ( .A1(n9439), .A2(n9566), .ZN(n9565) );
  NAND2_X1 U9507 ( .A1(n9438), .A2(n9437), .ZN(n9566) );
  NOR2_X1 U9508 ( .A1(n8051), .A2(n7754), .ZN(n9439) );
  OR2_X1 U9509 ( .A1(n9437), .A2(n9438), .ZN(n9564) );
  AND2_X1 U9510 ( .A1(n9567), .A2(n9568), .ZN(n9438) );
  NAND2_X1 U9511 ( .A1(n9569), .A2(b_26_), .ZN(n9568) );
  NOR2_X1 U9512 ( .A1(n9570), .A2(n7743), .ZN(n9569) );
  NOR2_X1 U9513 ( .A1(n9433), .A2(n9434), .ZN(n9570) );
  NAND2_X1 U9514 ( .A1(n9433), .A2(n9434), .ZN(n9567) );
  NAND2_X1 U9515 ( .A1(n9571), .A2(n9572), .ZN(n9434) );
  NAND2_X1 U9516 ( .A1(n9431), .A2(n9573), .ZN(n9572) );
  NAND2_X1 U9517 ( .A1(n9430), .A2(n9429), .ZN(n9573) );
  NOR2_X1 U9518 ( .A1(n8051), .A2(n7723), .ZN(n9431) );
  OR2_X1 U9519 ( .A1(n9429), .A2(n9430), .ZN(n9571) );
  AND2_X1 U9520 ( .A1(n9574), .A2(n9575), .ZN(n9430) );
  NAND2_X1 U9521 ( .A1(n9576), .A2(b_26_), .ZN(n9575) );
  NOR2_X1 U9522 ( .A1(n9577), .A2(n7707), .ZN(n9576) );
  NOR2_X1 U9523 ( .A1(n9426), .A2(n9424), .ZN(n9577) );
  NAND2_X1 U9524 ( .A1(n9424), .A2(n9426), .ZN(n9574) );
  NAND2_X1 U9525 ( .A1(n9578), .A2(n9579), .ZN(n9426) );
  NAND2_X1 U9526 ( .A1(n9423), .A2(n9580), .ZN(n9579) );
  NAND2_X1 U9527 ( .A1(n9422), .A2(n9421), .ZN(n9580) );
  NOR2_X1 U9528 ( .A1(n8051), .A2(n7687), .ZN(n9423) );
  OR2_X1 U9529 ( .A1(n9421), .A2(n9422), .ZN(n9578) );
  AND2_X1 U9530 ( .A1(n9581), .A2(n9582), .ZN(n9422) );
  NAND2_X1 U9531 ( .A1(n9583), .A2(b_26_), .ZN(n9582) );
  NOR2_X1 U9532 ( .A1(n9584), .A2(n7676), .ZN(n9583) );
  NOR2_X1 U9533 ( .A1(n9418), .A2(n9417), .ZN(n9584) );
  NAND2_X1 U9534 ( .A1(n9417), .A2(n9418), .ZN(n9581) );
  NAND2_X1 U9535 ( .A1(n9585), .A2(n9586), .ZN(n9418) );
  NAND2_X1 U9536 ( .A1(n9415), .A2(n9587), .ZN(n9586) );
  OR2_X1 U9537 ( .A1(n9414), .A2(n9412), .ZN(n9587) );
  NOR2_X1 U9538 ( .A1(n8051), .A2(n7656), .ZN(n9415) );
  NAND2_X1 U9539 ( .A1(n9412), .A2(n9414), .ZN(n9585) );
  NAND2_X1 U9540 ( .A1(n9588), .A2(n9589), .ZN(n9414) );
  NAND2_X1 U9541 ( .A1(n9590), .A2(b_26_), .ZN(n9589) );
  NOR2_X1 U9542 ( .A1(n9591), .A2(n7645), .ZN(n9590) );
  NOR2_X1 U9543 ( .A1(n9410), .A2(n9409), .ZN(n9591) );
  NAND2_X1 U9544 ( .A1(n9409), .A2(n9410), .ZN(n9588) );
  NAND2_X1 U9545 ( .A1(n9592), .A2(n9593), .ZN(n9410) );
  NAND2_X1 U9546 ( .A1(n9406), .A2(n9594), .ZN(n9593) );
  NAND2_X1 U9547 ( .A1(n9407), .A2(n9405), .ZN(n9594) );
  NOR2_X1 U9548 ( .A1(n8051), .A2(n7624), .ZN(n9406) );
  OR2_X1 U9549 ( .A1(n9405), .A2(n9407), .ZN(n9592) );
  AND2_X1 U9550 ( .A1(n9595), .A2(n9596), .ZN(n9407) );
  NAND2_X1 U9551 ( .A1(n9597), .A2(b_26_), .ZN(n9596) );
  NOR2_X1 U9552 ( .A1(n9598), .A2(n7613), .ZN(n9597) );
  NOR2_X1 U9553 ( .A1(n9402), .A2(n9400), .ZN(n9598) );
  NAND2_X1 U9554 ( .A1(n9400), .A2(n9402), .ZN(n9595) );
  NAND2_X1 U9555 ( .A1(n9599), .A2(n9600), .ZN(n9402) );
  NAND2_X1 U9556 ( .A1(n9399), .A2(n9601), .ZN(n9600) );
  NAND2_X1 U9557 ( .A1(n9398), .A2(n9397), .ZN(n9601) );
  NOR2_X1 U9558 ( .A1(n8051), .A2(n7593), .ZN(n9399) );
  OR2_X1 U9559 ( .A1(n9397), .A2(n9398), .ZN(n9599) );
  AND2_X1 U9560 ( .A1(n9602), .A2(n9603), .ZN(n9398) );
  NAND2_X1 U9561 ( .A1(n9394), .A2(n9604), .ZN(n9603) );
  NAND2_X1 U9562 ( .A1(n9395), .A2(n7577), .ZN(n9604) );
  INV_X1 U9563 ( .A(n9605), .ZN(n9395) );
  XNOR2_X1 U9564 ( .A(n9606), .B(n9607), .ZN(n9394) );
  XNOR2_X1 U9565 ( .A(n9608), .B(n9609), .ZN(n9606) );
  NAND2_X1 U9566 ( .A1(n9610), .A2(n9605), .ZN(n9602) );
  NAND2_X1 U9567 ( .A1(n9611), .A2(n9612), .ZN(n9605) );
  NAND2_X1 U9568 ( .A1(n9392), .A2(n9613), .ZN(n9612) );
  NAND2_X1 U9569 ( .A1(n9391), .A2(n9390), .ZN(n9613) );
  NOR2_X1 U9570 ( .A1(n8051), .A2(n7563), .ZN(n9392) );
  INV_X1 U9571 ( .A(b_26_), .ZN(n8051) );
  OR2_X1 U9572 ( .A1(n9390), .A2(n9391), .ZN(n9611) );
  AND2_X1 U9573 ( .A1(n9387), .A2(n9614), .ZN(n9391) );
  NAND2_X1 U9574 ( .A1(n9386), .A2(n9388), .ZN(n9614) );
  NAND2_X1 U9575 ( .A1(n9615), .A2(n9616), .ZN(n9388) );
  NAND2_X1 U9576 ( .A1(b_26_), .A2(a_28_), .ZN(n9616) );
  INV_X1 U9577 ( .A(n9617), .ZN(n9615) );
  XOR2_X1 U9578 ( .A(n9618), .B(n9619), .Z(n9386) );
  NOR2_X1 U9579 ( .A1(n7529), .A2(n7594), .ZN(n9619) );
  XOR2_X1 U9580 ( .A(n9620), .B(n9621), .Z(n9618) );
  NAND2_X1 U9581 ( .A1(a_28_), .A2(n9617), .ZN(n9387) );
  NAND2_X1 U9582 ( .A1(n9622), .A2(n9623), .ZN(n9617) );
  NAND2_X1 U9583 ( .A1(n9624), .A2(b_26_), .ZN(n9623) );
  NOR2_X1 U9584 ( .A1(n9625), .A2(n7529), .ZN(n9624) );
  NOR2_X1 U9585 ( .A1(n9373), .A2(n9374), .ZN(n9625) );
  NAND2_X1 U9586 ( .A1(n9373), .A2(n9374), .ZN(n9622) );
  NAND2_X1 U9587 ( .A1(n9626), .A2(n9627), .ZN(n9374) );
  NAND2_X1 U9588 ( .A1(n9628), .A2(b_24_), .ZN(n9627) );
  NOR2_X1 U9589 ( .A1(n9629), .A2(n8048), .ZN(n9628) );
  NOR2_X1 U9590 ( .A1(n8676), .A2(n7594), .ZN(n9629) );
  NAND2_X1 U9591 ( .A1(n9630), .A2(b_25_), .ZN(n9626) );
  NOR2_X1 U9592 ( .A1(n9631), .A2(n7515), .ZN(n9630) );
  NOR2_X1 U9593 ( .A1(n8679), .A2(n9632), .ZN(n9631) );
  AND2_X1 U9594 ( .A1(n9633), .A2(b_26_), .ZN(n9373) );
  NOR2_X1 U9595 ( .A1(n8451), .A2(n7594), .ZN(n9633) );
  XOR2_X1 U9596 ( .A(n9634), .B(n9635), .Z(n9390) );
  NAND2_X1 U9597 ( .A1(n9636), .A2(n9637), .ZN(n9634) );
  INV_X1 U9598 ( .A(n7577), .ZN(n9610) );
  NAND2_X1 U9599 ( .A1(b_26_), .A2(a_26_), .ZN(n7577) );
  XNOR2_X1 U9600 ( .A(n9638), .B(n9639), .ZN(n9397) );
  XNOR2_X1 U9601 ( .A(n9640), .B(n9641), .ZN(n9638) );
  NAND2_X1 U9602 ( .A1(b_25_), .A2(a_26_), .ZN(n9640) );
  XNOR2_X1 U9603 ( .A(n9642), .B(n9643), .ZN(n9400) );
  XNOR2_X1 U9604 ( .A(n9644), .B(n7588), .ZN(n9642) );
  XOR2_X1 U9605 ( .A(n9645), .B(n9646), .Z(n9405) );
  XOR2_X1 U9606 ( .A(n9647), .B(n9648), .Z(n9646) );
  NAND2_X1 U9607 ( .A1(b_25_), .A2(a_24_), .ZN(n9648) );
  XNOR2_X1 U9608 ( .A(n9649), .B(n9650), .ZN(n9409) );
  XNOR2_X1 U9609 ( .A(n9651), .B(n9652), .ZN(n9650) );
  XOR2_X1 U9610 ( .A(n9653), .B(n9654), .Z(n9412) );
  XOR2_X1 U9611 ( .A(n9655), .B(n9656), .Z(n9653) );
  NOR2_X1 U9612 ( .A1(n7645), .A2(n7594), .ZN(n9656) );
  XNOR2_X1 U9613 ( .A(n9657), .B(n9658), .ZN(n9417) );
  XNOR2_X1 U9614 ( .A(n9659), .B(n9660), .ZN(n9657) );
  XOR2_X1 U9615 ( .A(n9661), .B(n9662), .Z(n9421) );
  XOR2_X1 U9616 ( .A(n9663), .B(n9664), .Z(n9662) );
  NAND2_X1 U9617 ( .A1(b_25_), .A2(a_20_), .ZN(n9664) );
  XNOR2_X1 U9618 ( .A(n9665), .B(n9666), .ZN(n9424) );
  XNOR2_X1 U9619 ( .A(n9667), .B(n9668), .ZN(n9665) );
  XNOR2_X1 U9620 ( .A(n9669), .B(n9670), .ZN(n9429) );
  XOR2_X1 U9621 ( .A(n9671), .B(n9672), .Z(n9669) );
  NOR2_X1 U9622 ( .A1(n7707), .A2(n7594), .ZN(n9672) );
  XOR2_X1 U9623 ( .A(n9673), .B(n9674), .Z(n9433) );
  XOR2_X1 U9624 ( .A(n9675), .B(n9676), .Z(n9673) );
  XNOR2_X1 U9625 ( .A(n9677), .B(n9678), .ZN(n9437) );
  XOR2_X1 U9626 ( .A(n9679), .B(n9680), .Z(n9677) );
  NOR2_X1 U9627 ( .A1(n7743), .A2(n7594), .ZN(n9680) );
  XNOR2_X1 U9628 ( .A(n9681), .B(n9682), .ZN(n9441) );
  XNOR2_X1 U9629 ( .A(n9683), .B(n9684), .ZN(n9681) );
  XNOR2_X1 U9630 ( .A(n9685), .B(n9686), .ZN(n9445) );
  XOR2_X1 U9631 ( .A(n9687), .B(n9688), .Z(n9686) );
  NAND2_X1 U9632 ( .A1(b_25_), .A2(a_14_), .ZN(n9688) );
  XOR2_X1 U9633 ( .A(n9689), .B(n9690), .Z(n9448) );
  XOR2_X1 U9634 ( .A(n9691), .B(n9692), .Z(n9689) );
  XOR2_X1 U9635 ( .A(n9693), .B(n9694), .Z(n9453) );
  XOR2_X1 U9636 ( .A(n9695), .B(n9696), .Z(n9693) );
  NOR2_X1 U9637 ( .A1(n7806), .A2(n7594), .ZN(n9696) );
  XOR2_X1 U9638 ( .A(n9697), .B(n9698), .Z(n9457) );
  XOR2_X1 U9639 ( .A(n9699), .B(n9700), .Z(n9697) );
  NOR2_X1 U9640 ( .A1(n7817), .A2(n7594), .ZN(n9700) );
  XNOR2_X1 U9641 ( .A(n9701), .B(n9702), .ZN(n9461) );
  XOR2_X1 U9642 ( .A(n9703), .B(n9704), .Z(n9701) );
  NOR2_X1 U9643 ( .A1(n7837), .A2(n7594), .ZN(n9704) );
  XNOR2_X1 U9644 ( .A(n9705), .B(n9706), .ZN(n9465) );
  XNOR2_X1 U9645 ( .A(n9707), .B(n9708), .ZN(n9705) );
  XOR2_X1 U9646 ( .A(n9709), .B(n9710), .Z(n9477) );
  XOR2_X1 U9647 ( .A(n9711), .B(n9712), .Z(n9709) );
  XOR2_X1 U9648 ( .A(n9713), .B(n9714), .Z(n9480) );
  XOR2_X1 U9649 ( .A(n9715), .B(n9716), .Z(n9713) );
  NOR2_X1 U9650 ( .A1(n7914), .A2(n7594), .ZN(n9716) );
  XOR2_X1 U9651 ( .A(n9717), .B(n9718), .Z(n9275) );
  XOR2_X1 U9652 ( .A(n9719), .B(n9720), .Z(n9717) );
  NOR2_X1 U9653 ( .A1(n7934), .A2(n7594), .ZN(n9720) );
  XNOR2_X1 U9654 ( .A(n9721), .B(n9722), .ZN(n9489) );
  NAND2_X1 U9655 ( .A1(n9723), .A2(n9724), .ZN(n9721) );
  XOR2_X1 U9656 ( .A(n9725), .B(n9726), .Z(n9260) );
  XOR2_X1 U9657 ( .A(n9727), .B(n9728), .Z(n9725) );
  NOR2_X1 U9658 ( .A1(n7973), .A2(n7594), .ZN(n9728) );
  XNOR2_X1 U9659 ( .A(n9729), .B(n9730), .ZN(n8279) );
  XNOR2_X1 U9660 ( .A(n9731), .B(n9732), .ZN(n9729) );
  AND2_X1 U9661 ( .A1(n8274), .A2(n9496), .ZN(n9497) );
  NAND2_X1 U9662 ( .A1(n9733), .A2(n9734), .ZN(n9496) );
  XOR2_X1 U9663 ( .A(n9735), .B(n9736), .Z(n9734) );
  NOR2_X1 U9664 ( .A1(n9737), .A2(n9738), .ZN(n9733) );
  NOR2_X1 U9665 ( .A1(n9731), .A2(n9730), .ZN(n9738) );
  INV_X1 U9666 ( .A(n9739), .ZN(n9737) );
  OR2_X1 U9667 ( .A1(n8274), .A2(n8273), .ZN(n8111) );
  XNOR2_X1 U9668 ( .A(n8270), .B(n8269), .ZN(n8273) );
  NAND2_X1 U9669 ( .A1(n9740), .A2(n9741), .ZN(n8274) );
  NAND2_X1 U9670 ( .A1(n9742), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U9671 ( .A1(n9732), .A2(n9743), .ZN(n9739) );
  NAND2_X1 U9672 ( .A1(n9731), .A2(n9730), .ZN(n9743) );
  NOR2_X1 U9673 ( .A1(n7594), .A2(n8307), .ZN(n9732) );
  OR2_X1 U9674 ( .A1(n9730), .A2(n9731), .ZN(n9742) );
  AND2_X1 U9675 ( .A1(n9744), .A2(n9745), .ZN(n9731) );
  NAND2_X1 U9676 ( .A1(n9746), .A2(b_25_), .ZN(n9745) );
  NOR2_X1 U9677 ( .A1(n9747), .A2(n7973), .ZN(n9746) );
  NOR2_X1 U9678 ( .A1(n9726), .A2(n9727), .ZN(n9747) );
  NAND2_X1 U9679 ( .A1(n9726), .A2(n9727), .ZN(n9744) );
  NAND2_X1 U9680 ( .A1(n9723), .A2(n9748), .ZN(n9727) );
  NAND2_X1 U9681 ( .A1(n9722), .A2(n9724), .ZN(n9748) );
  NAND2_X1 U9682 ( .A1(n9749), .A2(n9750), .ZN(n9724) );
  NAND2_X1 U9683 ( .A1(b_25_), .A2(a_2_), .ZN(n9750) );
  INV_X1 U9684 ( .A(n9751), .ZN(n9749) );
  XNOR2_X1 U9685 ( .A(n9752), .B(n9753), .ZN(n9722) );
  NAND2_X1 U9686 ( .A1(n9754), .A2(n9755), .ZN(n9752) );
  NAND2_X1 U9687 ( .A1(a_2_), .A2(n9751), .ZN(n9723) );
  NAND2_X1 U9688 ( .A1(n9756), .A2(n9757), .ZN(n9751) );
  NAND2_X1 U9689 ( .A1(n9758), .A2(b_25_), .ZN(n9757) );
  NOR2_X1 U9690 ( .A1(n9759), .A2(n7945), .ZN(n9758) );
  NOR2_X1 U9691 ( .A1(n9510), .A2(n9511), .ZN(n9759) );
  NAND2_X1 U9692 ( .A1(n9510), .A2(n9511), .ZN(n9756) );
  NAND2_X1 U9693 ( .A1(n9760), .A2(n9761), .ZN(n9511) );
  NAND2_X1 U9694 ( .A1(n9762), .A2(b_25_), .ZN(n9761) );
  NOR2_X1 U9695 ( .A1(n9763), .A2(n7934), .ZN(n9762) );
  NOR2_X1 U9696 ( .A1(n9718), .A2(n9719), .ZN(n9763) );
  NAND2_X1 U9697 ( .A1(n9718), .A2(n9719), .ZN(n9760) );
  NAND2_X1 U9698 ( .A1(n9764), .A2(n9765), .ZN(n9719) );
  NAND2_X1 U9699 ( .A1(n9766), .A2(b_25_), .ZN(n9765) );
  NOR2_X1 U9700 ( .A1(n9767), .A2(n7914), .ZN(n9766) );
  NOR2_X1 U9701 ( .A1(n9714), .A2(n9715), .ZN(n9767) );
  NAND2_X1 U9702 ( .A1(n9714), .A2(n9715), .ZN(n9764) );
  NAND2_X1 U9703 ( .A1(n9768), .A2(n9769), .ZN(n9715) );
  NAND2_X1 U9704 ( .A1(n9711), .A2(n9770), .ZN(n9769) );
  OR2_X1 U9705 ( .A1(n9710), .A2(n9712), .ZN(n9770) );
  NAND2_X1 U9706 ( .A1(n9529), .A2(n9771), .ZN(n9711) );
  NAND2_X1 U9707 ( .A1(n9528), .A2(n9530), .ZN(n9771) );
  NAND2_X1 U9708 ( .A1(n9772), .A2(n9773), .ZN(n9530) );
  NAND2_X1 U9709 ( .A1(b_25_), .A2(a_7_), .ZN(n9773) );
  INV_X1 U9710 ( .A(n9774), .ZN(n9772) );
  XNOR2_X1 U9711 ( .A(n9775), .B(n9776), .ZN(n9528) );
  XOR2_X1 U9712 ( .A(n9777), .B(n9778), .Z(n9776) );
  NAND2_X1 U9713 ( .A1(b_24_), .A2(a_8_), .ZN(n9778) );
  NAND2_X1 U9714 ( .A1(a_7_), .A2(n9774), .ZN(n9529) );
  NAND2_X1 U9715 ( .A1(n9779), .A2(n9780), .ZN(n9774) );
  NAND2_X1 U9716 ( .A1(n9781), .A2(b_25_), .ZN(n9780) );
  NOR2_X1 U9717 ( .A1(n9782), .A2(n8059), .ZN(n9781) );
  NOR2_X1 U9718 ( .A1(n9535), .A2(n9537), .ZN(n9782) );
  NAND2_X1 U9719 ( .A1(n9535), .A2(n9537), .ZN(n9779) );
  NAND2_X1 U9720 ( .A1(n9783), .A2(n9784), .ZN(n9537) );
  NAND2_X1 U9721 ( .A1(n9708), .A2(n9785), .ZN(n9784) );
  NAND2_X1 U9722 ( .A1(n9707), .A2(n9706), .ZN(n9785) );
  NOR2_X1 U9723 ( .A1(n7594), .A2(n7848), .ZN(n9708) );
  OR2_X1 U9724 ( .A1(n9706), .A2(n9707), .ZN(n9783) );
  AND2_X1 U9725 ( .A1(n9786), .A2(n9787), .ZN(n9707) );
  NAND2_X1 U9726 ( .A1(n9788), .A2(b_25_), .ZN(n9787) );
  NOR2_X1 U9727 ( .A1(n9789), .A2(n7837), .ZN(n9788) );
  NOR2_X1 U9728 ( .A1(n9702), .A2(n9703), .ZN(n9789) );
  NAND2_X1 U9729 ( .A1(n9702), .A2(n9703), .ZN(n9786) );
  NAND2_X1 U9730 ( .A1(n9790), .A2(n9791), .ZN(n9703) );
  NAND2_X1 U9731 ( .A1(n9792), .A2(b_25_), .ZN(n9791) );
  NOR2_X1 U9732 ( .A1(n9793), .A2(n7817), .ZN(n9792) );
  NOR2_X1 U9733 ( .A1(n9698), .A2(n9699), .ZN(n9793) );
  NAND2_X1 U9734 ( .A1(n9698), .A2(n9699), .ZN(n9790) );
  NAND2_X1 U9735 ( .A1(n9794), .A2(n9795), .ZN(n9699) );
  NAND2_X1 U9736 ( .A1(n9796), .A2(b_25_), .ZN(n9795) );
  NOR2_X1 U9737 ( .A1(n9797), .A2(n7806), .ZN(n9796) );
  NOR2_X1 U9738 ( .A1(n9694), .A2(n9695), .ZN(n9797) );
  NAND2_X1 U9739 ( .A1(n9694), .A2(n9695), .ZN(n9794) );
  NAND2_X1 U9740 ( .A1(n9798), .A2(n9799), .ZN(n9695) );
  NAND2_X1 U9741 ( .A1(n9692), .A2(n9800), .ZN(n9799) );
  OR2_X1 U9742 ( .A1(n9691), .A2(n9690), .ZN(n9800) );
  NOR2_X1 U9743 ( .A1(n7594), .A2(n7786), .ZN(n9692) );
  NAND2_X1 U9744 ( .A1(n9690), .A2(n9691), .ZN(n9798) );
  NAND2_X1 U9745 ( .A1(n9801), .A2(n9802), .ZN(n9691) );
  NAND2_X1 U9746 ( .A1(n9803), .A2(b_25_), .ZN(n9802) );
  NOR2_X1 U9747 ( .A1(n9804), .A2(n7775), .ZN(n9803) );
  NOR2_X1 U9748 ( .A1(n9685), .A2(n9687), .ZN(n9804) );
  NAND2_X1 U9749 ( .A1(n9685), .A2(n9687), .ZN(n9801) );
  NAND2_X1 U9750 ( .A1(n9805), .A2(n9806), .ZN(n9687) );
  NAND2_X1 U9751 ( .A1(n9684), .A2(n9807), .ZN(n9806) );
  NAND2_X1 U9752 ( .A1(n9683), .A2(n9682), .ZN(n9807) );
  NOR2_X1 U9753 ( .A1(n7594), .A2(n7754), .ZN(n9684) );
  OR2_X1 U9754 ( .A1(n9682), .A2(n9683), .ZN(n9805) );
  AND2_X1 U9755 ( .A1(n9808), .A2(n9809), .ZN(n9683) );
  NAND2_X1 U9756 ( .A1(n9810), .A2(b_25_), .ZN(n9809) );
  NOR2_X1 U9757 ( .A1(n9811), .A2(n7743), .ZN(n9810) );
  NOR2_X1 U9758 ( .A1(n9678), .A2(n9679), .ZN(n9811) );
  NAND2_X1 U9759 ( .A1(n9678), .A2(n9679), .ZN(n9808) );
  NAND2_X1 U9760 ( .A1(n9812), .A2(n9813), .ZN(n9679) );
  NAND2_X1 U9761 ( .A1(n9676), .A2(n9814), .ZN(n9813) );
  OR2_X1 U9762 ( .A1(n9675), .A2(n9674), .ZN(n9814) );
  NOR2_X1 U9763 ( .A1(n7594), .A2(n7723), .ZN(n9676) );
  NAND2_X1 U9764 ( .A1(n9674), .A2(n9675), .ZN(n9812) );
  NAND2_X1 U9765 ( .A1(n9815), .A2(n9816), .ZN(n9675) );
  NAND2_X1 U9766 ( .A1(n9817), .A2(b_25_), .ZN(n9816) );
  NOR2_X1 U9767 ( .A1(n9818), .A2(n7707), .ZN(n9817) );
  NOR2_X1 U9768 ( .A1(n9670), .A2(n9671), .ZN(n9818) );
  NAND2_X1 U9769 ( .A1(n9670), .A2(n9671), .ZN(n9815) );
  NAND2_X1 U9770 ( .A1(n9819), .A2(n9820), .ZN(n9671) );
  NAND2_X1 U9771 ( .A1(n9667), .A2(n9821), .ZN(n9820) );
  NAND2_X1 U9772 ( .A1(n9668), .A2(n9666), .ZN(n9821) );
  NOR2_X1 U9773 ( .A1(n7594), .A2(n7687), .ZN(n9667) );
  OR2_X1 U9774 ( .A1(n9666), .A2(n9668), .ZN(n9819) );
  AND2_X1 U9775 ( .A1(n9822), .A2(n9823), .ZN(n9668) );
  NAND2_X1 U9776 ( .A1(n9824), .A2(b_25_), .ZN(n9823) );
  NOR2_X1 U9777 ( .A1(n9825), .A2(n7676), .ZN(n9824) );
  NOR2_X1 U9778 ( .A1(n9661), .A2(n9663), .ZN(n9825) );
  NAND2_X1 U9779 ( .A1(n9661), .A2(n9663), .ZN(n9822) );
  NAND2_X1 U9780 ( .A1(n9826), .A2(n9827), .ZN(n9663) );
  NAND2_X1 U9781 ( .A1(n9660), .A2(n9828), .ZN(n9827) );
  NAND2_X1 U9782 ( .A1(n9659), .A2(n9658), .ZN(n9828) );
  NOR2_X1 U9783 ( .A1(n7594), .A2(n7656), .ZN(n9660) );
  OR2_X1 U9784 ( .A1(n9658), .A2(n9659), .ZN(n9826) );
  AND2_X1 U9785 ( .A1(n9829), .A2(n9830), .ZN(n9659) );
  NAND2_X1 U9786 ( .A1(n9831), .A2(b_25_), .ZN(n9830) );
  NOR2_X1 U9787 ( .A1(n9832), .A2(n7645), .ZN(n9831) );
  NOR2_X1 U9788 ( .A1(n9654), .A2(n9655), .ZN(n9832) );
  NAND2_X1 U9789 ( .A1(n9654), .A2(n9655), .ZN(n9829) );
  NAND2_X1 U9790 ( .A1(n9833), .A2(n9834), .ZN(n9655) );
  NAND2_X1 U9791 ( .A1(n9652), .A2(n9835), .ZN(n9834) );
  OR2_X1 U9792 ( .A1(n9651), .A2(n9649), .ZN(n9835) );
  NOR2_X1 U9793 ( .A1(n7594), .A2(n7624), .ZN(n9652) );
  NAND2_X1 U9794 ( .A1(n9649), .A2(n9651), .ZN(n9833) );
  NAND2_X1 U9795 ( .A1(n9836), .A2(n9837), .ZN(n9651) );
  NAND2_X1 U9796 ( .A1(n9838), .A2(b_25_), .ZN(n9837) );
  NOR2_X1 U9797 ( .A1(n9839), .A2(n7613), .ZN(n9838) );
  NOR2_X1 U9798 ( .A1(n9645), .A2(n9647), .ZN(n9839) );
  NAND2_X1 U9799 ( .A1(n9645), .A2(n9647), .ZN(n9836) );
  NAND2_X1 U9800 ( .A1(n9840), .A2(n9841), .ZN(n9647) );
  NAND2_X1 U9801 ( .A1(n7588), .A2(n9842), .ZN(n9841) );
  NAND2_X1 U9802 ( .A1(n9644), .A2(n9643), .ZN(n9842) );
  NOR2_X1 U9803 ( .A1(n7594), .A2(n7593), .ZN(n7588) );
  OR2_X1 U9804 ( .A1(n9643), .A2(n9644), .ZN(n9840) );
  AND2_X1 U9805 ( .A1(n9843), .A2(n9844), .ZN(n9644) );
  NAND2_X1 U9806 ( .A1(n9845), .A2(b_25_), .ZN(n9844) );
  NOR2_X1 U9807 ( .A1(n9846), .A2(n8052), .ZN(n9845) );
  NOR2_X1 U9808 ( .A1(n9639), .A2(n9641), .ZN(n9846) );
  NAND2_X1 U9809 ( .A1(n9639), .A2(n9641), .ZN(n9843) );
  NAND2_X1 U9810 ( .A1(n9847), .A2(n9848), .ZN(n9641) );
  NAND2_X1 U9811 ( .A1(n9609), .A2(n9849), .ZN(n9848) );
  NAND2_X1 U9812 ( .A1(n9608), .A2(n9607), .ZN(n9849) );
  NOR2_X1 U9813 ( .A1(n7594), .A2(n7563), .ZN(n9609) );
  OR2_X1 U9814 ( .A1(n9607), .A2(n9608), .ZN(n9847) );
  AND2_X1 U9815 ( .A1(n9636), .A2(n9850), .ZN(n9608) );
  NAND2_X1 U9816 ( .A1(n9635), .A2(n9637), .ZN(n9850) );
  NAND2_X1 U9817 ( .A1(n9851), .A2(n9852), .ZN(n9637) );
  NAND2_X1 U9818 ( .A1(b_25_), .A2(a_28_), .ZN(n9852) );
  INV_X1 U9819 ( .A(n9853), .ZN(n9851) );
  XOR2_X1 U9820 ( .A(n9854), .B(n9855), .Z(n9635) );
  NOR2_X1 U9821 ( .A1(n7529), .A2(n9632), .ZN(n9855) );
  XOR2_X1 U9822 ( .A(n9856), .B(n9857), .Z(n9854) );
  NAND2_X1 U9823 ( .A1(a_28_), .A2(n9853), .ZN(n9636) );
  NAND2_X1 U9824 ( .A1(n9858), .A2(n9859), .ZN(n9853) );
  NAND2_X1 U9825 ( .A1(n9860), .A2(b_25_), .ZN(n9859) );
  NOR2_X1 U9826 ( .A1(n9861), .A2(n7529), .ZN(n9860) );
  NOR2_X1 U9827 ( .A1(n9620), .A2(n9621), .ZN(n9861) );
  NAND2_X1 U9828 ( .A1(n9620), .A2(n9621), .ZN(n9858) );
  NAND2_X1 U9829 ( .A1(n9862), .A2(n9863), .ZN(n9621) );
  NAND2_X1 U9830 ( .A1(n9864), .A2(b_23_), .ZN(n9863) );
  NOR2_X1 U9831 ( .A1(n9865), .A2(n8048), .ZN(n9864) );
  NOR2_X1 U9832 ( .A1(n8676), .A2(n9632), .ZN(n9865) );
  NAND2_X1 U9833 ( .A1(n9866), .A2(b_24_), .ZN(n9862) );
  NOR2_X1 U9834 ( .A1(n9867), .A2(n7515), .ZN(n9866) );
  NOR2_X1 U9835 ( .A1(n8679), .A2(n7625), .ZN(n9867) );
  AND2_X1 U9836 ( .A1(n9868), .A2(b_25_), .ZN(n9620) );
  NOR2_X1 U9837 ( .A1(n8451), .A2(n9632), .ZN(n9868) );
  XOR2_X1 U9838 ( .A(n9869), .B(n9870), .Z(n9607) );
  NAND2_X1 U9839 ( .A1(n9871), .A2(n9872), .ZN(n9869) );
  XNOR2_X1 U9840 ( .A(n9873), .B(n9874), .ZN(n9639) );
  XNOR2_X1 U9841 ( .A(n9875), .B(n9876), .ZN(n9873) );
  XNOR2_X1 U9842 ( .A(n9877), .B(n9878), .ZN(n9643) );
  XNOR2_X1 U9843 ( .A(n9879), .B(n9880), .ZN(n9877) );
  NAND2_X1 U9844 ( .A1(b_24_), .A2(a_26_), .ZN(n9879) );
  XNOR2_X1 U9845 ( .A(n9881), .B(n9882), .ZN(n9645) );
  XNOR2_X1 U9846 ( .A(n9883), .B(n9884), .ZN(n9881) );
  XNOR2_X1 U9847 ( .A(n9885), .B(n9886), .ZN(n9649) );
  XNOR2_X1 U9848 ( .A(n9887), .B(n7607), .ZN(n9886) );
  XNOR2_X1 U9849 ( .A(n9888), .B(n9889), .ZN(n9654) );
  XNOR2_X1 U9850 ( .A(n9890), .B(n9891), .ZN(n9888) );
  XOR2_X1 U9851 ( .A(n9892), .B(n9893), .Z(n9658) );
  XOR2_X1 U9852 ( .A(n9894), .B(n9895), .Z(n9893) );
  NAND2_X1 U9853 ( .A1(b_24_), .A2(a_22_), .ZN(n9895) );
  XNOR2_X1 U9854 ( .A(n9896), .B(n9897), .ZN(n9661) );
  XNOR2_X1 U9855 ( .A(n9898), .B(n9899), .ZN(n9896) );
  XNOR2_X1 U9856 ( .A(n9900), .B(n9901), .ZN(n9666) );
  XOR2_X1 U9857 ( .A(n9902), .B(n9903), .Z(n9900) );
  NOR2_X1 U9858 ( .A1(n7676), .A2(n9632), .ZN(n9903) );
  XNOR2_X1 U9859 ( .A(n9904), .B(n9905), .ZN(n9670) );
  XNOR2_X1 U9860 ( .A(n9906), .B(n9907), .ZN(n9904) );
  XOR2_X1 U9861 ( .A(n9908), .B(n9909), .Z(n9674) );
  XOR2_X1 U9862 ( .A(n9910), .B(n9911), .Z(n9908) );
  NOR2_X1 U9863 ( .A1(n7707), .A2(n9632), .ZN(n9911) );
  XNOR2_X1 U9864 ( .A(n9912), .B(n9913), .ZN(n9678) );
  XNOR2_X1 U9865 ( .A(n9914), .B(n9915), .ZN(n9912) );
  XOR2_X1 U9866 ( .A(n9916), .B(n9917), .Z(n9682) );
  XOR2_X1 U9867 ( .A(n9918), .B(n9919), .Z(n9917) );
  NAND2_X1 U9868 ( .A1(b_24_), .A2(a_16_), .ZN(n9919) );
  XOR2_X1 U9869 ( .A(n9920), .B(n9921), .Z(n9685) );
  XOR2_X1 U9870 ( .A(n9922), .B(n9923), .Z(n9920) );
  XOR2_X1 U9871 ( .A(n9924), .B(n9925), .Z(n9690) );
  XOR2_X1 U9872 ( .A(n9926), .B(n9927), .Z(n9924) );
  NOR2_X1 U9873 ( .A1(n7775), .A2(n9632), .ZN(n9927) );
  XOR2_X1 U9874 ( .A(n9928), .B(n9929), .Z(n9694) );
  XOR2_X1 U9875 ( .A(n9930), .B(n9931), .Z(n9928) );
  XOR2_X1 U9876 ( .A(n9932), .B(n9933), .Z(n9698) );
  XOR2_X1 U9877 ( .A(n9934), .B(n9935), .Z(n9932) );
  NOR2_X1 U9878 ( .A1(n7806), .A2(n9632), .ZN(n9935) );
  XNOR2_X1 U9879 ( .A(n9936), .B(n9937), .ZN(n9702) );
  NAND2_X1 U9880 ( .A1(n9938), .A2(n9939), .ZN(n9936) );
  XOR2_X1 U9881 ( .A(n9940), .B(n9941), .Z(n9706) );
  NAND2_X1 U9882 ( .A1(n9942), .A2(n9943), .ZN(n9940) );
  XNOR2_X1 U9883 ( .A(n9944), .B(n9945), .ZN(n9535) );
  XNOR2_X1 U9884 ( .A(n9946), .B(n9947), .ZN(n9945) );
  NAND2_X1 U9885 ( .A1(n9712), .A2(n9710), .ZN(n9768) );
  XNOR2_X1 U9886 ( .A(n9948), .B(n9949), .ZN(n9710) );
  NAND2_X1 U9887 ( .A1(n9950), .A2(n9951), .ZN(n9948) );
  NOR2_X1 U9888 ( .A1(n7594), .A2(n8061), .ZN(n9712) );
  XNOR2_X1 U9889 ( .A(n9952), .B(n9953), .ZN(n9714) );
  XNOR2_X1 U9890 ( .A(n9954), .B(n9955), .ZN(n9952) );
  XNOR2_X1 U9891 ( .A(n9956), .B(n9957), .ZN(n9718) );
  XNOR2_X1 U9892 ( .A(n9958), .B(n9959), .ZN(n9957) );
  XOR2_X1 U9893 ( .A(n9960), .B(n9961), .Z(n9510) );
  XOR2_X1 U9894 ( .A(n9962), .B(n9963), .Z(n9960) );
  NOR2_X1 U9895 ( .A1(n7934), .A2(n9632), .ZN(n9963) );
  XNOR2_X1 U9896 ( .A(n9964), .B(n9965), .ZN(n9726) );
  NAND2_X1 U9897 ( .A1(n9966), .A2(n9967), .ZN(n9964) );
  XOR2_X1 U9898 ( .A(n9968), .B(n9969), .Z(n9730) );
  XNOR2_X1 U9899 ( .A(n9970), .B(n9971), .ZN(n9968) );
  XNOR2_X1 U9900 ( .A(n9736), .B(n9735), .ZN(n9740) );
  XNOR2_X1 U9901 ( .A(n9972), .B(n9973), .ZN(n9736) );
  NOR2_X1 U9902 ( .A1(n8307), .A2(n9632), .ZN(n9973) );
  NAND2_X1 U9903 ( .A1(n9974), .A2(n9975), .ZN(n8116) );
  XOR2_X1 U9904 ( .A(n8263), .B(n8262), .Z(n9975) );
  INV_X1 U9905 ( .A(n8271), .ZN(n8262) );
  AND2_X1 U9906 ( .A1(n8270), .A2(n8269), .ZN(n9974) );
  XOR2_X1 U9907 ( .A(n9976), .B(n9977), .Z(n8269) );
  XOR2_X1 U9908 ( .A(n9978), .B(n9979), .Z(n9976) );
  NOR2_X1 U9909 ( .A1(n8307), .A2(n7625), .ZN(n9979) );
  NAND2_X1 U9910 ( .A1(n9980), .A2(n9981), .ZN(n8270) );
  NAND2_X1 U9911 ( .A1(n9982), .A2(b_24_), .ZN(n9981) );
  NOR2_X1 U9912 ( .A1(n9983), .A2(n8307), .ZN(n9982) );
  NOR2_X1 U9913 ( .A1(n9735), .A2(n9972), .ZN(n9983) );
  NAND2_X1 U9914 ( .A1(n9735), .A2(n9972), .ZN(n9980) );
  NAND2_X1 U9915 ( .A1(n9984), .A2(n9985), .ZN(n9972) );
  NAND2_X1 U9916 ( .A1(n9970), .A2(n9986), .ZN(n9985) );
  NAND2_X1 U9917 ( .A1(n9969), .A2(n9971), .ZN(n9986) );
  NAND2_X1 U9918 ( .A1(n9966), .A2(n9987), .ZN(n9970) );
  NAND2_X1 U9919 ( .A1(n9965), .A2(n9967), .ZN(n9987) );
  NAND2_X1 U9920 ( .A1(n9988), .A2(n9989), .ZN(n9967) );
  NAND2_X1 U9921 ( .A1(b_24_), .A2(a_2_), .ZN(n9989) );
  INV_X1 U9922 ( .A(n9990), .ZN(n9988) );
  XOR2_X1 U9923 ( .A(n9991), .B(n9992), .Z(n9965) );
  XOR2_X1 U9924 ( .A(n9993), .B(n9994), .Z(n9991) );
  NOR2_X1 U9925 ( .A1(n7945), .A2(n7625), .ZN(n9994) );
  NAND2_X1 U9926 ( .A1(a_2_), .A2(n9990), .ZN(n9966) );
  NAND2_X1 U9927 ( .A1(n9754), .A2(n9995), .ZN(n9990) );
  NAND2_X1 U9928 ( .A1(n9753), .A2(n9755), .ZN(n9995) );
  NAND2_X1 U9929 ( .A1(n9996), .A2(n9997), .ZN(n9755) );
  NAND2_X1 U9930 ( .A1(b_24_), .A2(a_3_), .ZN(n9997) );
  INV_X1 U9931 ( .A(n9998), .ZN(n9996) );
  XOR2_X1 U9932 ( .A(n9999), .B(n10000), .Z(n9753) );
  XOR2_X1 U9933 ( .A(n10001), .B(n10002), .Z(n9999) );
  NOR2_X1 U9934 ( .A1(n7934), .A2(n7625), .ZN(n10002) );
  NAND2_X1 U9935 ( .A1(a_3_), .A2(n9998), .ZN(n9754) );
  NAND2_X1 U9936 ( .A1(n10003), .A2(n10004), .ZN(n9998) );
  NAND2_X1 U9937 ( .A1(n10005), .A2(b_24_), .ZN(n10004) );
  NOR2_X1 U9938 ( .A1(n10006), .A2(n7934), .ZN(n10005) );
  NOR2_X1 U9939 ( .A1(n9961), .A2(n9962), .ZN(n10006) );
  NAND2_X1 U9940 ( .A1(n9961), .A2(n9962), .ZN(n10003) );
  NAND2_X1 U9941 ( .A1(n10007), .A2(n10008), .ZN(n9962) );
  NAND2_X1 U9942 ( .A1(n9959), .A2(n10009), .ZN(n10008) );
  OR2_X1 U9943 ( .A1(n9958), .A2(n9956), .ZN(n10009) );
  NOR2_X1 U9944 ( .A1(n9632), .A2(n7914), .ZN(n9959) );
  NAND2_X1 U9945 ( .A1(n9956), .A2(n9958), .ZN(n10007) );
  NAND2_X1 U9946 ( .A1(n10010), .A2(n10011), .ZN(n9958) );
  NAND2_X1 U9947 ( .A1(n9954), .A2(n10012), .ZN(n10011) );
  NAND2_X1 U9948 ( .A1(n9953), .A2(n9955), .ZN(n10012) );
  NAND2_X1 U9949 ( .A1(n9950), .A2(n10013), .ZN(n9954) );
  NAND2_X1 U9950 ( .A1(n9949), .A2(n9951), .ZN(n10013) );
  NAND2_X1 U9951 ( .A1(n10014), .A2(n10015), .ZN(n9951) );
  NAND2_X1 U9952 ( .A1(b_24_), .A2(a_7_), .ZN(n10015) );
  INV_X1 U9953 ( .A(n10016), .ZN(n10014) );
  XNOR2_X1 U9954 ( .A(n10017), .B(n10018), .ZN(n9949) );
  XNOR2_X1 U9955 ( .A(n10019), .B(n10020), .ZN(n10017) );
  NAND2_X1 U9956 ( .A1(a_7_), .A2(n10016), .ZN(n9950) );
  NAND2_X1 U9957 ( .A1(n10021), .A2(n10022), .ZN(n10016) );
  NAND2_X1 U9958 ( .A1(n10023), .A2(b_24_), .ZN(n10022) );
  NOR2_X1 U9959 ( .A1(n10024), .A2(n8059), .ZN(n10023) );
  NOR2_X1 U9960 ( .A1(n9775), .A2(n9777), .ZN(n10024) );
  NAND2_X1 U9961 ( .A1(n9775), .A2(n9777), .ZN(n10021) );
  NAND2_X1 U9962 ( .A1(n10025), .A2(n10026), .ZN(n9777) );
  NAND2_X1 U9963 ( .A1(n9947), .A2(n10027), .ZN(n10026) );
  OR2_X1 U9964 ( .A1(n9946), .A2(n9944), .ZN(n10027) );
  NOR2_X1 U9965 ( .A1(n9632), .A2(n7848), .ZN(n9947) );
  NAND2_X1 U9966 ( .A1(n9944), .A2(n9946), .ZN(n10025) );
  NAND2_X1 U9967 ( .A1(n9942), .A2(n10028), .ZN(n9946) );
  NAND2_X1 U9968 ( .A1(n9941), .A2(n9943), .ZN(n10028) );
  NAND2_X1 U9969 ( .A1(n10029), .A2(n10030), .ZN(n9943) );
  NAND2_X1 U9970 ( .A1(b_24_), .A2(a_10_), .ZN(n10030) );
  INV_X1 U9971 ( .A(n10031), .ZN(n10029) );
  XOR2_X1 U9972 ( .A(n10032), .B(n10033), .Z(n9941) );
  XOR2_X1 U9973 ( .A(n10034), .B(n10035), .Z(n10032) );
  NOR2_X1 U9974 ( .A1(n7817), .A2(n7625), .ZN(n10035) );
  NAND2_X1 U9975 ( .A1(a_10_), .A2(n10031), .ZN(n9942) );
  NAND2_X1 U9976 ( .A1(n9938), .A2(n10036), .ZN(n10031) );
  NAND2_X1 U9977 ( .A1(n9937), .A2(n9939), .ZN(n10036) );
  NAND2_X1 U9978 ( .A1(n10037), .A2(n10038), .ZN(n9939) );
  NAND2_X1 U9979 ( .A1(b_24_), .A2(a_11_), .ZN(n10038) );
  INV_X1 U9980 ( .A(n10039), .ZN(n10037) );
  XNOR2_X1 U9981 ( .A(n10040), .B(n10041), .ZN(n9937) );
  XNOR2_X1 U9982 ( .A(n10042), .B(n10043), .ZN(n10041) );
  NOR2_X1 U9983 ( .A1(n7806), .A2(n7625), .ZN(n10043) );
  NAND2_X1 U9984 ( .A1(a_11_), .A2(n10039), .ZN(n9938) );
  NAND2_X1 U9985 ( .A1(n10044), .A2(n10045), .ZN(n10039) );
  NAND2_X1 U9986 ( .A1(n10046), .A2(b_24_), .ZN(n10045) );
  NOR2_X1 U9987 ( .A1(n10047), .A2(n7806), .ZN(n10046) );
  NOR2_X1 U9988 ( .A1(n9933), .A2(n9934), .ZN(n10047) );
  NAND2_X1 U9989 ( .A1(n9933), .A2(n9934), .ZN(n10044) );
  NAND2_X1 U9990 ( .A1(n10048), .A2(n10049), .ZN(n9934) );
  NAND2_X1 U9991 ( .A1(n9931), .A2(n10050), .ZN(n10049) );
  OR2_X1 U9992 ( .A1(n9930), .A2(n9929), .ZN(n10050) );
  NOR2_X1 U9993 ( .A1(n9632), .A2(n7786), .ZN(n9931) );
  NAND2_X1 U9994 ( .A1(n9929), .A2(n9930), .ZN(n10048) );
  NAND2_X1 U9995 ( .A1(n10051), .A2(n10052), .ZN(n9930) );
  NAND2_X1 U9996 ( .A1(n10053), .A2(b_24_), .ZN(n10052) );
  NOR2_X1 U9997 ( .A1(n10054), .A2(n7775), .ZN(n10053) );
  NOR2_X1 U9998 ( .A1(n9925), .A2(n9926), .ZN(n10054) );
  NAND2_X1 U9999 ( .A1(n9925), .A2(n9926), .ZN(n10051) );
  NAND2_X1 U10000 ( .A1(n10055), .A2(n10056), .ZN(n9926) );
  NAND2_X1 U10001 ( .A1(n9923), .A2(n10057), .ZN(n10056) );
  OR2_X1 U10002 ( .A1(n9922), .A2(n9921), .ZN(n10057) );
  NOR2_X1 U10003 ( .A1(n9632), .A2(n7754), .ZN(n9923) );
  NAND2_X1 U10004 ( .A1(n9921), .A2(n9922), .ZN(n10055) );
  NAND2_X1 U10005 ( .A1(n10058), .A2(n10059), .ZN(n9922) );
  NAND2_X1 U10006 ( .A1(n10060), .A2(b_24_), .ZN(n10059) );
  NOR2_X1 U10007 ( .A1(n10061), .A2(n7743), .ZN(n10060) );
  NOR2_X1 U10008 ( .A1(n9916), .A2(n9918), .ZN(n10061) );
  NAND2_X1 U10009 ( .A1(n9916), .A2(n9918), .ZN(n10058) );
  NAND2_X1 U10010 ( .A1(n10062), .A2(n10063), .ZN(n9918) );
  NAND2_X1 U10011 ( .A1(n9915), .A2(n10064), .ZN(n10063) );
  NAND2_X1 U10012 ( .A1(n9914), .A2(n9913), .ZN(n10064) );
  NOR2_X1 U10013 ( .A1(n9632), .A2(n7723), .ZN(n9915) );
  OR2_X1 U10014 ( .A1(n9913), .A2(n9914), .ZN(n10062) );
  AND2_X1 U10015 ( .A1(n10065), .A2(n10066), .ZN(n9914) );
  NAND2_X1 U10016 ( .A1(n10067), .A2(b_24_), .ZN(n10066) );
  NOR2_X1 U10017 ( .A1(n10068), .A2(n7707), .ZN(n10067) );
  NOR2_X1 U10018 ( .A1(n9909), .A2(n9910), .ZN(n10068) );
  NAND2_X1 U10019 ( .A1(n9909), .A2(n9910), .ZN(n10065) );
  NAND2_X1 U10020 ( .A1(n10069), .A2(n10070), .ZN(n9910) );
  NAND2_X1 U10021 ( .A1(n9907), .A2(n10071), .ZN(n10070) );
  NAND2_X1 U10022 ( .A1(n9906), .A2(n9905), .ZN(n10071) );
  NOR2_X1 U10023 ( .A1(n9632), .A2(n7687), .ZN(n9907) );
  OR2_X1 U10024 ( .A1(n9905), .A2(n9906), .ZN(n10069) );
  AND2_X1 U10025 ( .A1(n10072), .A2(n10073), .ZN(n9906) );
  NAND2_X1 U10026 ( .A1(n10074), .A2(b_24_), .ZN(n10073) );
  NOR2_X1 U10027 ( .A1(n10075), .A2(n7676), .ZN(n10074) );
  NOR2_X1 U10028 ( .A1(n9901), .A2(n9902), .ZN(n10075) );
  NAND2_X1 U10029 ( .A1(n9901), .A2(n9902), .ZN(n10072) );
  NAND2_X1 U10030 ( .A1(n10076), .A2(n10077), .ZN(n9902) );
  NAND2_X1 U10031 ( .A1(n9899), .A2(n10078), .ZN(n10077) );
  NAND2_X1 U10032 ( .A1(n9898), .A2(n9897), .ZN(n10078) );
  NOR2_X1 U10033 ( .A1(n9632), .A2(n7656), .ZN(n9899) );
  OR2_X1 U10034 ( .A1(n9897), .A2(n9898), .ZN(n10076) );
  AND2_X1 U10035 ( .A1(n10079), .A2(n10080), .ZN(n9898) );
  NAND2_X1 U10036 ( .A1(n10081), .A2(b_24_), .ZN(n10080) );
  NOR2_X1 U10037 ( .A1(n10082), .A2(n7645), .ZN(n10081) );
  NOR2_X1 U10038 ( .A1(n9892), .A2(n9894), .ZN(n10082) );
  NAND2_X1 U10039 ( .A1(n9892), .A2(n9894), .ZN(n10079) );
  NAND2_X1 U10040 ( .A1(n10083), .A2(n10084), .ZN(n9894) );
  NAND2_X1 U10041 ( .A1(n9891), .A2(n10085), .ZN(n10084) );
  NAND2_X1 U10042 ( .A1(n9890), .A2(n9889), .ZN(n10085) );
  NOR2_X1 U10043 ( .A1(n9632), .A2(n7624), .ZN(n9891) );
  OR2_X1 U10044 ( .A1(n9889), .A2(n9890), .ZN(n10083) );
  AND2_X1 U10045 ( .A1(n10086), .A2(n10087), .ZN(n9890) );
  NAND2_X1 U10046 ( .A1(n9885), .A2(n10088), .ZN(n10087) );
  OR2_X1 U10047 ( .A1(n9887), .A2(n7607), .ZN(n10088) );
  XNOR2_X1 U10048 ( .A(n10089), .B(n10090), .ZN(n9885) );
  XNOR2_X1 U10049 ( .A(n10091), .B(n10092), .ZN(n10089) );
  NAND2_X1 U10050 ( .A1(n7607), .A2(n9887), .ZN(n10086) );
  NAND2_X1 U10051 ( .A1(n10093), .A2(n10094), .ZN(n9887) );
  NAND2_X1 U10052 ( .A1(n9884), .A2(n10095), .ZN(n10094) );
  NAND2_X1 U10053 ( .A1(n9883), .A2(n9882), .ZN(n10095) );
  NOR2_X1 U10054 ( .A1(n9632), .A2(n7593), .ZN(n9884) );
  OR2_X1 U10055 ( .A1(n9882), .A2(n9883), .ZN(n10093) );
  AND2_X1 U10056 ( .A1(n10096), .A2(n10097), .ZN(n9883) );
  NAND2_X1 U10057 ( .A1(n10098), .A2(b_24_), .ZN(n10097) );
  NOR2_X1 U10058 ( .A1(n10099), .A2(n8052), .ZN(n10098) );
  NOR2_X1 U10059 ( .A1(n9878), .A2(n9880), .ZN(n10099) );
  NAND2_X1 U10060 ( .A1(n9878), .A2(n9880), .ZN(n10096) );
  NAND2_X1 U10061 ( .A1(n10100), .A2(n10101), .ZN(n9880) );
  NAND2_X1 U10062 ( .A1(n9876), .A2(n10102), .ZN(n10101) );
  NAND2_X1 U10063 ( .A1(n9875), .A2(n9874), .ZN(n10102) );
  NOR2_X1 U10064 ( .A1(n9632), .A2(n7563), .ZN(n9876) );
  OR2_X1 U10065 ( .A1(n9874), .A2(n9875), .ZN(n10100) );
  AND2_X1 U10066 ( .A1(n9871), .A2(n10103), .ZN(n9875) );
  NAND2_X1 U10067 ( .A1(n9870), .A2(n9872), .ZN(n10103) );
  NAND2_X1 U10068 ( .A1(n10104), .A2(n10105), .ZN(n9872) );
  NAND2_X1 U10069 ( .A1(b_24_), .A2(a_28_), .ZN(n10105) );
  INV_X1 U10070 ( .A(n10106), .ZN(n10104) );
  XOR2_X1 U10071 ( .A(n10107), .B(n10108), .Z(n9870) );
  NOR2_X1 U10072 ( .A1(n7529), .A2(n7625), .ZN(n10108) );
  XOR2_X1 U10073 ( .A(n10109), .B(n10110), .Z(n10107) );
  NAND2_X1 U10074 ( .A1(a_28_), .A2(n10106), .ZN(n9871) );
  NAND2_X1 U10075 ( .A1(n10111), .A2(n10112), .ZN(n10106) );
  NAND2_X1 U10076 ( .A1(n10113), .A2(b_24_), .ZN(n10112) );
  NOR2_X1 U10077 ( .A1(n10114), .A2(n7529), .ZN(n10113) );
  NOR2_X1 U10078 ( .A1(n9856), .A2(n9857), .ZN(n10114) );
  NAND2_X1 U10079 ( .A1(n9856), .A2(n9857), .ZN(n10111) );
  NAND2_X1 U10080 ( .A1(n10115), .A2(n10116), .ZN(n9857) );
  NAND2_X1 U10081 ( .A1(n10117), .A2(b_22_), .ZN(n10116) );
  NOR2_X1 U10082 ( .A1(n10118), .A2(n8048), .ZN(n10117) );
  NOR2_X1 U10083 ( .A1(n8676), .A2(n7625), .ZN(n10118) );
  NAND2_X1 U10084 ( .A1(n10119), .A2(b_23_), .ZN(n10115) );
  NOR2_X1 U10085 ( .A1(n10120), .A2(n7515), .ZN(n10119) );
  NOR2_X1 U10086 ( .A1(n8679), .A2(n8053), .ZN(n10120) );
  AND2_X1 U10087 ( .A1(n10121), .A2(b_24_), .ZN(n9856) );
  XOR2_X1 U10088 ( .A(n10122), .B(n10123), .Z(n9874) );
  NAND2_X1 U10089 ( .A1(n10124), .A2(n10125), .ZN(n10122) );
  XNOR2_X1 U10090 ( .A(n10126), .B(n10127), .ZN(n9878) );
  XNOR2_X1 U10091 ( .A(n10128), .B(n10129), .ZN(n10126) );
  XNOR2_X1 U10092 ( .A(n10130), .B(n10131), .ZN(n9882) );
  XNOR2_X1 U10093 ( .A(n10132), .B(n10133), .ZN(n10130) );
  NAND2_X1 U10094 ( .A1(b_23_), .A2(a_26_), .ZN(n10132) );
  NOR2_X1 U10095 ( .A1(n9632), .A2(n7613), .ZN(n7607) );
  INV_X1 U10096 ( .A(b_24_), .ZN(n9632) );
  XOR2_X1 U10097 ( .A(n10134), .B(n10135), .Z(n9889) );
  XOR2_X1 U10098 ( .A(n10136), .B(n10137), .Z(n10135) );
  NAND2_X1 U10099 ( .A1(b_23_), .A2(a_24_), .ZN(n10137) );
  XNOR2_X1 U10100 ( .A(n10138), .B(n10139), .ZN(n9892) );
  XOR2_X1 U10101 ( .A(n10140), .B(n8031), .Z(n10138) );
  XNOR2_X1 U10102 ( .A(n10141), .B(n10142), .ZN(n9897) );
  XOR2_X1 U10103 ( .A(n10143), .B(n10144), .Z(n10141) );
  NOR2_X1 U10104 ( .A1(n7645), .A2(n7625), .ZN(n10144) );
  XNOR2_X1 U10105 ( .A(n10145), .B(n10146), .ZN(n9901) );
  XNOR2_X1 U10106 ( .A(n10147), .B(n10148), .ZN(n10146) );
  XNOR2_X1 U10107 ( .A(n10149), .B(n10150), .ZN(n9905) );
  XOR2_X1 U10108 ( .A(n10151), .B(n10152), .Z(n10149) );
  NOR2_X1 U10109 ( .A1(n7676), .A2(n7625), .ZN(n10152) );
  XOR2_X1 U10110 ( .A(n10153), .B(n10154), .Z(n9909) );
  XOR2_X1 U10111 ( .A(n10155), .B(n10156), .Z(n10153) );
  XOR2_X1 U10112 ( .A(n10157), .B(n10158), .Z(n9913) );
  XOR2_X1 U10113 ( .A(n10159), .B(n10160), .Z(n10158) );
  NAND2_X1 U10114 ( .A1(b_23_), .A2(a_18_), .ZN(n10160) );
  XNOR2_X1 U10115 ( .A(n10161), .B(n10162), .ZN(n9916) );
  XNOR2_X1 U10116 ( .A(n10163), .B(n10164), .ZN(n10161) );
  XOR2_X1 U10117 ( .A(n10165), .B(n10166), .Z(n9921) );
  XOR2_X1 U10118 ( .A(n10167), .B(n10168), .Z(n10165) );
  NOR2_X1 U10119 ( .A1(n7743), .A2(n7625), .ZN(n10168) );
  XNOR2_X1 U10120 ( .A(n10169), .B(n10170), .ZN(n9925) );
  XOR2_X1 U10121 ( .A(n10171), .B(n10172), .Z(n10170) );
  NAND2_X1 U10122 ( .A1(b_23_), .A2(a_15_), .ZN(n10172) );
  XOR2_X1 U10123 ( .A(n10173), .B(n10174), .Z(n9929) );
  XOR2_X1 U10124 ( .A(n10175), .B(n10176), .Z(n10173) );
  NOR2_X1 U10125 ( .A1(n7775), .A2(n7625), .ZN(n10176) );
  XOR2_X1 U10126 ( .A(n10177), .B(n10178), .Z(n9933) );
  XOR2_X1 U10127 ( .A(n10179), .B(n10180), .Z(n10177) );
  XOR2_X1 U10128 ( .A(n10181), .B(n10182), .Z(n9944) );
  XOR2_X1 U10129 ( .A(n10183), .B(n10184), .Z(n10181) );
  NOR2_X1 U10130 ( .A1(n7837), .A2(n7625), .ZN(n10184) );
  XOR2_X1 U10131 ( .A(n10185), .B(n10186), .Z(n9775) );
  XOR2_X1 U10132 ( .A(n10187), .B(n10188), .Z(n10185) );
  OR2_X1 U10133 ( .A1(n9955), .A2(n9953), .ZN(n10010) );
  XNOR2_X1 U10134 ( .A(n10189), .B(n10190), .ZN(n9953) );
  XOR2_X1 U10135 ( .A(n10191), .B(n10192), .Z(n10189) );
  NOR2_X1 U10136 ( .A1(n7884), .A2(n7625), .ZN(n10192) );
  NAND2_X1 U10137 ( .A1(b_24_), .A2(a_6_), .ZN(n9955) );
  XNOR2_X1 U10138 ( .A(n10193), .B(n10194), .ZN(n9956) );
  NAND2_X1 U10139 ( .A1(n10195), .A2(n10196), .ZN(n10193) );
  XOR2_X1 U10140 ( .A(n10197), .B(n10198), .Z(n9961) );
  XOR2_X1 U10141 ( .A(n10199), .B(n10200), .Z(n10197) );
  NOR2_X1 U10142 ( .A1(n7914), .A2(n7625), .ZN(n10200) );
  OR2_X1 U10143 ( .A1(n9971), .A2(n9969), .ZN(n9984) );
  XOR2_X1 U10144 ( .A(n10201), .B(n10202), .Z(n9969) );
  XOR2_X1 U10145 ( .A(n10203), .B(n10204), .Z(n10202) );
  NAND2_X1 U10146 ( .A1(b_23_), .A2(a_2_), .ZN(n10204) );
  NAND2_X1 U10147 ( .A1(b_24_), .A2(a_1_), .ZN(n9971) );
  XNOR2_X1 U10148 ( .A(n10205), .B(n10206), .ZN(n9735) );
  XOR2_X1 U10149 ( .A(n10207), .B(n10208), .Z(n10206) );
  NAND2_X1 U10150 ( .A1(b_23_), .A2(a_1_), .ZN(n10208) );
  NAND2_X1 U10151 ( .A1(n10209), .A2(n10210), .ZN(n8121) );
  AND2_X1 U10152 ( .A1(n10211), .A2(n8263), .ZN(n10210) );
  NAND2_X1 U10153 ( .A1(n10212), .A2(n10213), .ZN(n8263) );
  NAND2_X1 U10154 ( .A1(n10214), .A2(b_23_), .ZN(n10213) );
  NOR2_X1 U10155 ( .A1(n10215), .A2(n8307), .ZN(n10214) );
  NOR2_X1 U10156 ( .A1(n9977), .A2(n9978), .ZN(n10215) );
  NAND2_X1 U10157 ( .A1(n9977), .A2(n9978), .ZN(n10212) );
  NAND2_X1 U10158 ( .A1(n10216), .A2(n10217), .ZN(n9978) );
  NAND2_X1 U10159 ( .A1(n10218), .A2(b_23_), .ZN(n10217) );
  NOR2_X1 U10160 ( .A1(n10219), .A2(n7973), .ZN(n10218) );
  NOR2_X1 U10161 ( .A1(n10205), .A2(n10207), .ZN(n10219) );
  NAND2_X1 U10162 ( .A1(n10205), .A2(n10207), .ZN(n10216) );
  NAND2_X1 U10163 ( .A1(n10220), .A2(n10221), .ZN(n10207) );
  NAND2_X1 U10164 ( .A1(n10222), .A2(b_23_), .ZN(n10221) );
  NOR2_X1 U10165 ( .A1(n10223), .A2(n7965), .ZN(n10222) );
  NOR2_X1 U10166 ( .A1(n10201), .A2(n10203), .ZN(n10223) );
  NAND2_X1 U10167 ( .A1(n10201), .A2(n10203), .ZN(n10220) );
  NAND2_X1 U10168 ( .A1(n10224), .A2(n10225), .ZN(n10203) );
  NAND2_X1 U10169 ( .A1(n10226), .A2(b_23_), .ZN(n10225) );
  NOR2_X1 U10170 ( .A1(n10227), .A2(n7945), .ZN(n10226) );
  NOR2_X1 U10171 ( .A1(n9992), .A2(n9993), .ZN(n10227) );
  NAND2_X1 U10172 ( .A1(n9992), .A2(n9993), .ZN(n10224) );
  NAND2_X1 U10173 ( .A1(n10228), .A2(n10229), .ZN(n9993) );
  NAND2_X1 U10174 ( .A1(n10230), .A2(b_23_), .ZN(n10229) );
  NOR2_X1 U10175 ( .A1(n10231), .A2(n7934), .ZN(n10230) );
  NOR2_X1 U10176 ( .A1(n10000), .A2(n10001), .ZN(n10231) );
  NAND2_X1 U10177 ( .A1(n10000), .A2(n10001), .ZN(n10228) );
  NAND2_X1 U10178 ( .A1(n10232), .A2(n10233), .ZN(n10001) );
  NAND2_X1 U10179 ( .A1(n10234), .A2(b_23_), .ZN(n10233) );
  NOR2_X1 U10180 ( .A1(n10235), .A2(n7914), .ZN(n10234) );
  NOR2_X1 U10181 ( .A1(n10198), .A2(n10199), .ZN(n10235) );
  NAND2_X1 U10182 ( .A1(n10198), .A2(n10199), .ZN(n10232) );
  NAND2_X1 U10183 ( .A1(n10195), .A2(n10236), .ZN(n10199) );
  NAND2_X1 U10184 ( .A1(n10194), .A2(n10196), .ZN(n10236) );
  NAND2_X1 U10185 ( .A1(n10237), .A2(n10238), .ZN(n10196) );
  NAND2_X1 U10186 ( .A1(b_23_), .A2(a_6_), .ZN(n10238) );
  INV_X1 U10187 ( .A(n10239), .ZN(n10237) );
  XOR2_X1 U10188 ( .A(n10240), .B(n10241), .Z(n10194) );
  XOR2_X1 U10189 ( .A(n10242), .B(n10243), .Z(n10240) );
  NAND2_X1 U10190 ( .A1(a_6_), .A2(n10239), .ZN(n10195) );
  NAND2_X1 U10191 ( .A1(n10244), .A2(n10245), .ZN(n10239) );
  NAND2_X1 U10192 ( .A1(n10246), .A2(b_23_), .ZN(n10245) );
  NOR2_X1 U10193 ( .A1(n10247), .A2(n7884), .ZN(n10246) );
  NOR2_X1 U10194 ( .A1(n10190), .A2(n10191), .ZN(n10247) );
  NAND2_X1 U10195 ( .A1(n10190), .A2(n10191), .ZN(n10244) );
  NAND2_X1 U10196 ( .A1(n10248), .A2(n10249), .ZN(n10191) );
  NAND2_X1 U10197 ( .A1(n10020), .A2(n10250), .ZN(n10249) );
  NAND2_X1 U10198 ( .A1(n10019), .A2(n10018), .ZN(n10250) );
  NOR2_X1 U10199 ( .A1(n7625), .A2(n8059), .ZN(n10020) );
  OR2_X1 U10200 ( .A1(n10018), .A2(n10019), .ZN(n10248) );
  AND2_X1 U10201 ( .A1(n10251), .A2(n10252), .ZN(n10019) );
  NAND2_X1 U10202 ( .A1(n10188), .A2(n10253), .ZN(n10252) );
  OR2_X1 U10203 ( .A1(n10187), .A2(n10186), .ZN(n10253) );
  NOR2_X1 U10204 ( .A1(n7625), .A2(n7848), .ZN(n10188) );
  NAND2_X1 U10205 ( .A1(n10186), .A2(n10187), .ZN(n10251) );
  NAND2_X1 U10206 ( .A1(n10254), .A2(n10255), .ZN(n10187) );
  NAND2_X1 U10207 ( .A1(n10256), .A2(b_23_), .ZN(n10255) );
  NOR2_X1 U10208 ( .A1(n10257), .A2(n7837), .ZN(n10256) );
  NOR2_X1 U10209 ( .A1(n10182), .A2(n10183), .ZN(n10257) );
  NAND2_X1 U10210 ( .A1(n10182), .A2(n10183), .ZN(n10254) );
  NAND2_X1 U10211 ( .A1(n10258), .A2(n10259), .ZN(n10183) );
  NAND2_X1 U10212 ( .A1(n10260), .A2(b_23_), .ZN(n10259) );
  NOR2_X1 U10213 ( .A1(n10261), .A2(n7817), .ZN(n10260) );
  NOR2_X1 U10214 ( .A1(n10033), .A2(n10034), .ZN(n10261) );
  NAND2_X1 U10215 ( .A1(n10033), .A2(n10034), .ZN(n10258) );
  NAND2_X1 U10216 ( .A1(n10262), .A2(n10263), .ZN(n10034) );
  NAND2_X1 U10217 ( .A1(n10264), .A2(b_23_), .ZN(n10263) );
  NOR2_X1 U10218 ( .A1(n10265), .A2(n7806), .ZN(n10264) );
  NOR2_X1 U10219 ( .A1(n10040), .A2(n10042), .ZN(n10265) );
  NAND2_X1 U10220 ( .A1(n10040), .A2(n10042), .ZN(n10262) );
  NAND2_X1 U10221 ( .A1(n10266), .A2(n10267), .ZN(n10042) );
  NAND2_X1 U10222 ( .A1(n10180), .A2(n10268), .ZN(n10267) );
  OR2_X1 U10223 ( .A1(n10179), .A2(n10178), .ZN(n10268) );
  NOR2_X1 U10224 ( .A1(n7625), .A2(n7786), .ZN(n10180) );
  NAND2_X1 U10225 ( .A1(n10178), .A2(n10179), .ZN(n10266) );
  NAND2_X1 U10226 ( .A1(n10269), .A2(n10270), .ZN(n10179) );
  NAND2_X1 U10227 ( .A1(n10271), .A2(b_23_), .ZN(n10270) );
  NOR2_X1 U10228 ( .A1(n10272), .A2(n7775), .ZN(n10271) );
  NOR2_X1 U10229 ( .A1(n10174), .A2(n10175), .ZN(n10272) );
  NAND2_X1 U10230 ( .A1(n10174), .A2(n10175), .ZN(n10269) );
  NAND2_X1 U10231 ( .A1(n10273), .A2(n10274), .ZN(n10175) );
  NAND2_X1 U10232 ( .A1(n10275), .A2(b_23_), .ZN(n10274) );
  NOR2_X1 U10233 ( .A1(n10276), .A2(n7754), .ZN(n10275) );
  NOR2_X1 U10234 ( .A1(n10169), .A2(n10171), .ZN(n10276) );
  NAND2_X1 U10235 ( .A1(n10169), .A2(n10171), .ZN(n10273) );
  NAND2_X1 U10236 ( .A1(n10277), .A2(n10278), .ZN(n10171) );
  NAND2_X1 U10237 ( .A1(n10279), .A2(b_23_), .ZN(n10278) );
  NOR2_X1 U10238 ( .A1(n10280), .A2(n7743), .ZN(n10279) );
  NOR2_X1 U10239 ( .A1(n10166), .A2(n10167), .ZN(n10280) );
  NAND2_X1 U10240 ( .A1(n10166), .A2(n10167), .ZN(n10277) );
  NAND2_X1 U10241 ( .A1(n10281), .A2(n10282), .ZN(n10167) );
  NAND2_X1 U10242 ( .A1(n10164), .A2(n10283), .ZN(n10282) );
  NAND2_X1 U10243 ( .A1(n10163), .A2(n10162), .ZN(n10283) );
  NOR2_X1 U10244 ( .A1(n7625), .A2(n7723), .ZN(n10164) );
  OR2_X1 U10245 ( .A1(n10162), .A2(n10163), .ZN(n10281) );
  AND2_X1 U10246 ( .A1(n10284), .A2(n10285), .ZN(n10163) );
  NAND2_X1 U10247 ( .A1(n10286), .A2(b_23_), .ZN(n10285) );
  NOR2_X1 U10248 ( .A1(n10287), .A2(n7707), .ZN(n10286) );
  NOR2_X1 U10249 ( .A1(n10157), .A2(n10159), .ZN(n10287) );
  NAND2_X1 U10250 ( .A1(n10157), .A2(n10159), .ZN(n10284) );
  NAND2_X1 U10251 ( .A1(n10288), .A2(n10289), .ZN(n10159) );
  NAND2_X1 U10252 ( .A1(n10156), .A2(n10290), .ZN(n10289) );
  OR2_X1 U10253 ( .A1(n10155), .A2(n10154), .ZN(n10290) );
  NOR2_X1 U10254 ( .A1(n7625), .A2(n7687), .ZN(n10156) );
  NAND2_X1 U10255 ( .A1(n10154), .A2(n10155), .ZN(n10288) );
  NAND2_X1 U10256 ( .A1(n10291), .A2(n10292), .ZN(n10155) );
  NAND2_X1 U10257 ( .A1(n10293), .A2(b_23_), .ZN(n10292) );
  NOR2_X1 U10258 ( .A1(n10294), .A2(n7676), .ZN(n10293) );
  NOR2_X1 U10259 ( .A1(n10150), .A2(n10151), .ZN(n10294) );
  NAND2_X1 U10260 ( .A1(n10150), .A2(n10151), .ZN(n10291) );
  NAND2_X1 U10261 ( .A1(n10295), .A2(n10296), .ZN(n10151) );
  NAND2_X1 U10262 ( .A1(n10148), .A2(n10297), .ZN(n10296) );
  OR2_X1 U10263 ( .A1(n10147), .A2(n10145), .ZN(n10297) );
  NOR2_X1 U10264 ( .A1(n7625), .A2(n7656), .ZN(n10148) );
  NAND2_X1 U10265 ( .A1(n10145), .A2(n10147), .ZN(n10295) );
  NAND2_X1 U10266 ( .A1(n10298), .A2(n10299), .ZN(n10147) );
  NAND2_X1 U10267 ( .A1(n10300), .A2(b_23_), .ZN(n10299) );
  NOR2_X1 U10268 ( .A1(n10301), .A2(n7645), .ZN(n10300) );
  NOR2_X1 U10269 ( .A1(n10142), .A2(n10143), .ZN(n10301) );
  NAND2_X1 U10270 ( .A1(n10142), .A2(n10143), .ZN(n10298) );
  NAND2_X1 U10271 ( .A1(n10302), .A2(n10303), .ZN(n10143) );
  NAND2_X1 U10272 ( .A1(n7619), .A2(n10304), .ZN(n10303) );
  NAND2_X1 U10273 ( .A1(n10140), .A2(n10139), .ZN(n10304) );
  INV_X1 U10274 ( .A(n8031), .ZN(n7619) );
  NAND2_X1 U10275 ( .A1(b_23_), .A2(a_23_), .ZN(n8031) );
  OR2_X1 U10276 ( .A1(n10139), .A2(n10140), .ZN(n10302) );
  AND2_X1 U10277 ( .A1(n10305), .A2(n10306), .ZN(n10140) );
  NAND2_X1 U10278 ( .A1(n10307), .A2(b_23_), .ZN(n10306) );
  NOR2_X1 U10279 ( .A1(n10308), .A2(n7613), .ZN(n10307) );
  NOR2_X1 U10280 ( .A1(n10134), .A2(n10136), .ZN(n10308) );
  NAND2_X1 U10281 ( .A1(n10134), .A2(n10136), .ZN(n10305) );
  NAND2_X1 U10282 ( .A1(n10309), .A2(n10310), .ZN(n10136) );
  NAND2_X1 U10283 ( .A1(n10092), .A2(n10311), .ZN(n10310) );
  NAND2_X1 U10284 ( .A1(n10091), .A2(n10090), .ZN(n10311) );
  NOR2_X1 U10285 ( .A1(n7625), .A2(n7593), .ZN(n10092) );
  OR2_X1 U10286 ( .A1(n10090), .A2(n10091), .ZN(n10309) );
  AND2_X1 U10287 ( .A1(n10312), .A2(n10313), .ZN(n10091) );
  NAND2_X1 U10288 ( .A1(n10314), .A2(b_23_), .ZN(n10313) );
  NOR2_X1 U10289 ( .A1(n10315), .A2(n8052), .ZN(n10314) );
  NOR2_X1 U10290 ( .A1(n10131), .A2(n10133), .ZN(n10315) );
  NAND2_X1 U10291 ( .A1(n10131), .A2(n10133), .ZN(n10312) );
  NAND2_X1 U10292 ( .A1(n10316), .A2(n10317), .ZN(n10133) );
  NAND2_X1 U10293 ( .A1(n10129), .A2(n10318), .ZN(n10317) );
  NAND2_X1 U10294 ( .A1(n10128), .A2(n10127), .ZN(n10318) );
  NOR2_X1 U10295 ( .A1(n7625), .A2(n7563), .ZN(n10129) );
  OR2_X1 U10296 ( .A1(n10127), .A2(n10128), .ZN(n10316) );
  AND2_X1 U10297 ( .A1(n10124), .A2(n10319), .ZN(n10128) );
  NAND2_X1 U10298 ( .A1(n10123), .A2(n10125), .ZN(n10319) );
  NAND2_X1 U10299 ( .A1(n10320), .A2(n10321), .ZN(n10125) );
  NAND2_X1 U10300 ( .A1(b_23_), .A2(a_28_), .ZN(n10321) );
  INV_X1 U10301 ( .A(n10322), .ZN(n10320) );
  XOR2_X1 U10302 ( .A(n10323), .B(n10324), .Z(n10123) );
  NOR2_X1 U10303 ( .A1(n7529), .A2(n8053), .ZN(n10324) );
  XOR2_X1 U10304 ( .A(n10325), .B(n10326), .Z(n10323) );
  NAND2_X1 U10305 ( .A1(a_28_), .A2(n10322), .ZN(n10124) );
  NAND2_X1 U10306 ( .A1(n10327), .A2(n10328), .ZN(n10322) );
  NAND2_X1 U10307 ( .A1(n10329), .A2(b_23_), .ZN(n10328) );
  NOR2_X1 U10308 ( .A1(n10330), .A2(n7529), .ZN(n10329) );
  NOR2_X1 U10309 ( .A1(n10109), .A2(n10110), .ZN(n10330) );
  NAND2_X1 U10310 ( .A1(n10109), .A2(n10110), .ZN(n10327) );
  NAND2_X1 U10311 ( .A1(n10331), .A2(n10332), .ZN(n10110) );
  NAND2_X1 U10312 ( .A1(n10333), .A2(b_21_), .ZN(n10332) );
  NOR2_X1 U10313 ( .A1(n10334), .A2(n8048), .ZN(n10333) );
  NOR2_X1 U10314 ( .A1(n8676), .A2(n8053), .ZN(n10334) );
  NAND2_X1 U10315 ( .A1(n10335), .A2(b_22_), .ZN(n10331) );
  NOR2_X1 U10316 ( .A1(n10336), .A2(n7515), .ZN(n10335) );
  NOR2_X1 U10317 ( .A1(n8679), .A2(n7657), .ZN(n10336) );
  AND2_X1 U10318 ( .A1(n10121), .A2(b_22_), .ZN(n10109) );
  NOR2_X1 U10319 ( .A1(n8451), .A2(n7625), .ZN(n10121) );
  XOR2_X1 U10320 ( .A(n10337), .B(n10338), .Z(n10127) );
  NAND2_X1 U10321 ( .A1(n10339), .A2(n10340), .ZN(n10337) );
  XNOR2_X1 U10322 ( .A(n10341), .B(n10342), .ZN(n10131) );
  XNOR2_X1 U10323 ( .A(n10343), .B(n10344), .ZN(n10341) );
  XNOR2_X1 U10324 ( .A(n10345), .B(n10346), .ZN(n10090) );
  XNOR2_X1 U10325 ( .A(n10347), .B(n10348), .ZN(n10345) );
  NAND2_X1 U10326 ( .A1(b_22_), .A2(a_26_), .ZN(n10347) );
  XNOR2_X1 U10327 ( .A(n10349), .B(n10350), .ZN(n10134) );
  XNOR2_X1 U10328 ( .A(n10351), .B(n10352), .ZN(n10350) );
  XOR2_X1 U10329 ( .A(n10353), .B(n10354), .Z(n10139) );
  XOR2_X1 U10330 ( .A(n10355), .B(n10356), .Z(n10354) );
  NAND2_X1 U10331 ( .A1(b_22_), .A2(a_24_), .ZN(n10356) );
  XNOR2_X1 U10332 ( .A(n10357), .B(n10358), .ZN(n10142) );
  XNOR2_X1 U10333 ( .A(n10359), .B(n10360), .ZN(n10357) );
  XOR2_X1 U10334 ( .A(n10361), .B(n10362), .Z(n10145) );
  XOR2_X1 U10335 ( .A(n10363), .B(n10364), .Z(n10361) );
  XNOR2_X1 U10336 ( .A(n10365), .B(n10366), .ZN(n10150) );
  XNOR2_X1 U10337 ( .A(n10367), .B(n10368), .ZN(n10366) );
  XNOR2_X1 U10338 ( .A(n10369), .B(n10370), .ZN(n10154) );
  XOR2_X1 U10339 ( .A(n10371), .B(n10372), .Z(n10370) );
  NAND2_X1 U10340 ( .A1(b_22_), .A2(a_20_), .ZN(n10372) );
  XNOR2_X1 U10341 ( .A(n10373), .B(n10374), .ZN(n10157) );
  XNOR2_X1 U10342 ( .A(n10375), .B(n10376), .ZN(n10373) );
  XNOR2_X1 U10343 ( .A(n10377), .B(n10378), .ZN(n10162) );
  XOR2_X1 U10344 ( .A(n10379), .B(n10380), .Z(n10377) );
  NOR2_X1 U10345 ( .A1(n7707), .A2(n8053), .ZN(n10380) );
  XOR2_X1 U10346 ( .A(n10381), .B(n10382), .Z(n10166) );
  XOR2_X1 U10347 ( .A(n10383), .B(n10384), .Z(n10381) );
  XOR2_X1 U10348 ( .A(n10385), .B(n10386), .Z(n10169) );
  XOR2_X1 U10349 ( .A(n10387), .B(n10388), .Z(n10385) );
  NOR2_X1 U10350 ( .A1(n7743), .A2(n8053), .ZN(n10388) );
  XOR2_X1 U10351 ( .A(n10389), .B(n10390), .Z(n10174) );
  XOR2_X1 U10352 ( .A(n10391), .B(n10392), .Z(n10389) );
  XNOR2_X1 U10353 ( .A(n10393), .B(n10394), .ZN(n10178) );
  XOR2_X1 U10354 ( .A(n10395), .B(n10396), .Z(n10394) );
  NAND2_X1 U10355 ( .A1(b_22_), .A2(a_14_), .ZN(n10396) );
  XOR2_X1 U10356 ( .A(n10397), .B(n10398), .Z(n10040) );
  XOR2_X1 U10357 ( .A(n10399), .B(n10400), .Z(n10397) );
  XOR2_X1 U10358 ( .A(n10401), .B(n10402), .Z(n10033) );
  XOR2_X1 U10359 ( .A(n10403), .B(n10404), .Z(n10401) );
  NOR2_X1 U10360 ( .A1(n7806), .A2(n8053), .ZN(n10404) );
  XOR2_X1 U10361 ( .A(n10405), .B(n10406), .Z(n10182) );
  XOR2_X1 U10362 ( .A(n10407), .B(n10408), .Z(n10405) );
  XOR2_X1 U10363 ( .A(n10409), .B(n10410), .Z(n10186) );
  XOR2_X1 U10364 ( .A(n10411), .B(n10412), .Z(n10409) );
  NOR2_X1 U10365 ( .A1(n7837), .A2(n8053), .ZN(n10412) );
  XNOR2_X1 U10366 ( .A(n10413), .B(n10414), .ZN(n10018) );
  XOR2_X1 U10367 ( .A(n10415), .B(n10416), .Z(n10413) );
  NOR2_X1 U10368 ( .A1(n7848), .A2(n8053), .ZN(n10416) );
  XNOR2_X1 U10369 ( .A(n10417), .B(n10418), .ZN(n10190) );
  XNOR2_X1 U10370 ( .A(n10419), .B(n10420), .ZN(n10417) );
  XOR2_X1 U10371 ( .A(n10421), .B(n10422), .Z(n10198) );
  XOR2_X1 U10372 ( .A(n10423), .B(n10424), .Z(n10421) );
  XNOR2_X1 U10373 ( .A(n10425), .B(n10426), .ZN(n10000) );
  XOR2_X1 U10374 ( .A(n10427), .B(n10428), .Z(n10426) );
  NAND2_X1 U10375 ( .A1(b_22_), .A2(a_5_), .ZN(n10428) );
  XNOR2_X1 U10376 ( .A(n10429), .B(n10430), .ZN(n9992) );
  NAND2_X1 U10377 ( .A1(n10431), .A2(n10432), .ZN(n10429) );
  XNOR2_X1 U10378 ( .A(n10433), .B(n10434), .ZN(n10201) );
  XNOR2_X1 U10379 ( .A(n10435), .B(n10436), .ZN(n10433) );
  XOR2_X1 U10380 ( .A(n10437), .B(n10438), .Z(n10205) );
  XOR2_X1 U10381 ( .A(n10439), .B(n10440), .Z(n10437) );
  XNOR2_X1 U10382 ( .A(n10441), .B(n10442), .ZN(n9977) );
  XOR2_X1 U10383 ( .A(n10443), .B(n10444), .Z(n10442) );
  NAND2_X1 U10384 ( .A1(b_22_), .A2(a_1_), .ZN(n10444) );
  NOR2_X1 U10385 ( .A1(n10445), .A2(n8271), .ZN(n10209) );
  XOR2_X1 U10386 ( .A(n10446), .B(n10447), .Z(n8271) );
  XNOR2_X1 U10387 ( .A(n10448), .B(n10449), .ZN(n10447) );
  NOR2_X1 U10388 ( .A1(n8264), .A2(n8265), .ZN(n10445) );
  NAND2_X1 U10389 ( .A1(n10450), .A2(n10211), .ZN(n8126) );
  OR2_X1 U10390 ( .A1(n10211), .A2(n10450), .ZN(n8127) );
  NAND2_X1 U10391 ( .A1(n8257), .A2(n10451), .ZN(n10450) );
  NAND2_X1 U10392 ( .A1(n10452), .A2(n10453), .ZN(n10451) );
  INV_X1 U10393 ( .A(n10454), .ZN(n10453) );
  XOR2_X1 U10394 ( .A(n10455), .B(n10456), .Z(n10452) );
  NAND2_X1 U10395 ( .A1(n8264), .A2(n8265), .ZN(n10211) );
  NAND2_X1 U10396 ( .A1(n10457), .A2(n10458), .ZN(n8265) );
  NAND2_X1 U10397 ( .A1(n10449), .A2(n10459), .ZN(n10458) );
  OR2_X1 U10398 ( .A1(n10448), .A2(n10446), .ZN(n10459) );
  NOR2_X1 U10399 ( .A1(n8053), .A2(n8307), .ZN(n10449) );
  NAND2_X1 U10400 ( .A1(n10446), .A2(n10448), .ZN(n10457) );
  NAND2_X1 U10401 ( .A1(n10460), .A2(n10461), .ZN(n10448) );
  NAND2_X1 U10402 ( .A1(n10462), .A2(b_22_), .ZN(n10461) );
  NOR2_X1 U10403 ( .A1(n10463), .A2(n7973), .ZN(n10462) );
  NOR2_X1 U10404 ( .A1(n10443), .A2(n10441), .ZN(n10463) );
  NAND2_X1 U10405 ( .A1(n10441), .A2(n10443), .ZN(n10460) );
  NAND2_X1 U10406 ( .A1(n10464), .A2(n10465), .ZN(n10443) );
  NAND2_X1 U10407 ( .A1(n10440), .A2(n10466), .ZN(n10465) );
  OR2_X1 U10408 ( .A1(n10438), .A2(n10439), .ZN(n10466) );
  NOR2_X1 U10409 ( .A1(n8053), .A2(n7965), .ZN(n10440) );
  NAND2_X1 U10410 ( .A1(n10438), .A2(n10439), .ZN(n10464) );
  NAND2_X1 U10411 ( .A1(n10467), .A2(n10468), .ZN(n10439) );
  NAND2_X1 U10412 ( .A1(n10436), .A2(n10469), .ZN(n10468) );
  NAND2_X1 U10413 ( .A1(n10435), .A2(n10434), .ZN(n10469) );
  NOR2_X1 U10414 ( .A1(n8053), .A2(n7945), .ZN(n10436) );
  OR2_X1 U10415 ( .A1(n10434), .A2(n10435), .ZN(n10467) );
  AND2_X1 U10416 ( .A1(n10431), .A2(n10470), .ZN(n10435) );
  NAND2_X1 U10417 ( .A1(n10430), .A2(n10432), .ZN(n10470) );
  NAND2_X1 U10418 ( .A1(n10471), .A2(n10472), .ZN(n10432) );
  NAND2_X1 U10419 ( .A1(b_22_), .A2(a_4_), .ZN(n10472) );
  INV_X1 U10420 ( .A(n10473), .ZN(n10471) );
  XOR2_X1 U10421 ( .A(n10474), .B(n10475), .Z(n10430) );
  XOR2_X1 U10422 ( .A(n10476), .B(n10477), .Z(n10474) );
  NOR2_X1 U10423 ( .A1(n7914), .A2(n7657), .ZN(n10477) );
  NAND2_X1 U10424 ( .A1(a_4_), .A2(n10473), .ZN(n10431) );
  NAND2_X1 U10425 ( .A1(n10478), .A2(n10479), .ZN(n10473) );
  NAND2_X1 U10426 ( .A1(n10480), .A2(b_22_), .ZN(n10479) );
  NOR2_X1 U10427 ( .A1(n10481), .A2(n7914), .ZN(n10480) );
  NOR2_X1 U10428 ( .A1(n10425), .A2(n10427), .ZN(n10481) );
  NAND2_X1 U10429 ( .A1(n10425), .A2(n10427), .ZN(n10478) );
  NAND2_X1 U10430 ( .A1(n10482), .A2(n10483), .ZN(n10427) );
  NAND2_X1 U10431 ( .A1(n10424), .A2(n10484), .ZN(n10483) );
  OR2_X1 U10432 ( .A1(n10422), .A2(n10423), .ZN(n10484) );
  NOR2_X1 U10433 ( .A1(n8053), .A2(n8061), .ZN(n10424) );
  NAND2_X1 U10434 ( .A1(n10422), .A2(n10423), .ZN(n10482) );
  NAND2_X1 U10435 ( .A1(n10485), .A2(n10486), .ZN(n10423) );
  NAND2_X1 U10436 ( .A1(n10243), .A2(n10487), .ZN(n10486) );
  OR2_X1 U10437 ( .A1(n10241), .A2(n10242), .ZN(n10487) );
  NOR2_X1 U10438 ( .A1(n8053), .A2(n7884), .ZN(n10243) );
  NAND2_X1 U10439 ( .A1(n10241), .A2(n10242), .ZN(n10485) );
  NAND2_X1 U10440 ( .A1(n10488), .A2(n10489), .ZN(n10242) );
  NAND2_X1 U10441 ( .A1(n10420), .A2(n10490), .ZN(n10489) );
  NAND2_X1 U10442 ( .A1(n10419), .A2(n10418), .ZN(n10490) );
  NOR2_X1 U10443 ( .A1(n8053), .A2(n8059), .ZN(n10420) );
  OR2_X1 U10444 ( .A1(n10418), .A2(n10419), .ZN(n10488) );
  AND2_X1 U10445 ( .A1(n10491), .A2(n10492), .ZN(n10419) );
  NAND2_X1 U10446 ( .A1(n10493), .A2(b_22_), .ZN(n10492) );
  NOR2_X1 U10447 ( .A1(n10494), .A2(n7848), .ZN(n10493) );
  NOR2_X1 U10448 ( .A1(n10415), .A2(n10414), .ZN(n10494) );
  NAND2_X1 U10449 ( .A1(n10414), .A2(n10415), .ZN(n10491) );
  NAND2_X1 U10450 ( .A1(n10495), .A2(n10496), .ZN(n10415) );
  NAND2_X1 U10451 ( .A1(n10497), .A2(b_22_), .ZN(n10496) );
  NOR2_X1 U10452 ( .A1(n10498), .A2(n7837), .ZN(n10497) );
  NOR2_X1 U10453 ( .A1(n10410), .A2(n10411), .ZN(n10498) );
  NAND2_X1 U10454 ( .A1(n10410), .A2(n10411), .ZN(n10495) );
  NAND2_X1 U10455 ( .A1(n10499), .A2(n10500), .ZN(n10411) );
  NAND2_X1 U10456 ( .A1(n10408), .A2(n10501), .ZN(n10500) );
  OR2_X1 U10457 ( .A1(n10406), .A2(n10407), .ZN(n10501) );
  NOR2_X1 U10458 ( .A1(n8053), .A2(n7817), .ZN(n10408) );
  NAND2_X1 U10459 ( .A1(n10406), .A2(n10407), .ZN(n10499) );
  NAND2_X1 U10460 ( .A1(n10502), .A2(n10503), .ZN(n10407) );
  NAND2_X1 U10461 ( .A1(n10504), .A2(b_22_), .ZN(n10503) );
  NOR2_X1 U10462 ( .A1(n10505), .A2(n7806), .ZN(n10504) );
  NOR2_X1 U10463 ( .A1(n10402), .A2(n10403), .ZN(n10505) );
  NAND2_X1 U10464 ( .A1(n10402), .A2(n10403), .ZN(n10502) );
  NAND2_X1 U10465 ( .A1(n10506), .A2(n10507), .ZN(n10403) );
  NAND2_X1 U10466 ( .A1(n10400), .A2(n10508), .ZN(n10507) );
  OR2_X1 U10467 ( .A1(n10398), .A2(n10399), .ZN(n10508) );
  NOR2_X1 U10468 ( .A1(n8053), .A2(n7786), .ZN(n10400) );
  NAND2_X1 U10469 ( .A1(n10398), .A2(n10399), .ZN(n10506) );
  NAND2_X1 U10470 ( .A1(n10509), .A2(n10510), .ZN(n10399) );
  NAND2_X1 U10471 ( .A1(n10511), .A2(b_22_), .ZN(n10510) );
  NOR2_X1 U10472 ( .A1(n10512), .A2(n7775), .ZN(n10511) );
  NOR2_X1 U10473 ( .A1(n10393), .A2(n10395), .ZN(n10512) );
  NAND2_X1 U10474 ( .A1(n10393), .A2(n10395), .ZN(n10509) );
  NAND2_X1 U10475 ( .A1(n10513), .A2(n10514), .ZN(n10395) );
  NAND2_X1 U10476 ( .A1(n10392), .A2(n10515), .ZN(n10514) );
  OR2_X1 U10477 ( .A1(n10390), .A2(n10391), .ZN(n10515) );
  NOR2_X1 U10478 ( .A1(n8053), .A2(n7754), .ZN(n10392) );
  NAND2_X1 U10479 ( .A1(n10390), .A2(n10391), .ZN(n10513) );
  NAND2_X1 U10480 ( .A1(n10516), .A2(n10517), .ZN(n10391) );
  NAND2_X1 U10481 ( .A1(n10518), .A2(b_22_), .ZN(n10517) );
  NOR2_X1 U10482 ( .A1(n10519), .A2(n7743), .ZN(n10518) );
  NOR2_X1 U10483 ( .A1(n10386), .A2(n10387), .ZN(n10519) );
  NAND2_X1 U10484 ( .A1(n10386), .A2(n10387), .ZN(n10516) );
  NAND2_X1 U10485 ( .A1(n10520), .A2(n10521), .ZN(n10387) );
  NAND2_X1 U10486 ( .A1(n10383), .A2(n10522), .ZN(n10521) );
  OR2_X1 U10487 ( .A1(n10382), .A2(n10384), .ZN(n10522) );
  NOR2_X1 U10488 ( .A1(n8053), .A2(n7723), .ZN(n10383) );
  NAND2_X1 U10489 ( .A1(n10382), .A2(n10384), .ZN(n10520) );
  NAND2_X1 U10490 ( .A1(n10523), .A2(n10524), .ZN(n10384) );
  NAND2_X1 U10491 ( .A1(n10525), .A2(b_22_), .ZN(n10524) );
  NOR2_X1 U10492 ( .A1(n10526), .A2(n7707), .ZN(n10525) );
  NOR2_X1 U10493 ( .A1(n10379), .A2(n10378), .ZN(n10526) );
  NAND2_X1 U10494 ( .A1(n10378), .A2(n10379), .ZN(n10523) );
  NAND2_X1 U10495 ( .A1(n10527), .A2(n10528), .ZN(n10379) );
  NAND2_X1 U10496 ( .A1(n10376), .A2(n10529), .ZN(n10528) );
  NAND2_X1 U10497 ( .A1(n10375), .A2(n10374), .ZN(n10529) );
  NOR2_X1 U10498 ( .A1(n8053), .A2(n7687), .ZN(n10376) );
  OR2_X1 U10499 ( .A1(n10374), .A2(n10375), .ZN(n10527) );
  AND2_X1 U10500 ( .A1(n10530), .A2(n10531), .ZN(n10375) );
  NAND2_X1 U10501 ( .A1(n10532), .A2(b_22_), .ZN(n10531) );
  NOR2_X1 U10502 ( .A1(n10533), .A2(n7676), .ZN(n10532) );
  NOR2_X1 U10503 ( .A1(n10369), .A2(n10371), .ZN(n10533) );
  NAND2_X1 U10504 ( .A1(n10369), .A2(n10371), .ZN(n10530) );
  NAND2_X1 U10505 ( .A1(n10534), .A2(n10535), .ZN(n10371) );
  NAND2_X1 U10506 ( .A1(n10368), .A2(n10536), .ZN(n10535) );
  OR2_X1 U10507 ( .A1(n10367), .A2(n10365), .ZN(n10536) );
  NOR2_X1 U10508 ( .A1(n8053), .A2(n7656), .ZN(n10368) );
  NAND2_X1 U10509 ( .A1(n10365), .A2(n10367), .ZN(n10534) );
  NAND2_X1 U10510 ( .A1(n10537), .A2(n10538), .ZN(n10367) );
  NAND2_X1 U10511 ( .A1(n10362), .A2(n10539), .ZN(n10538) );
  OR2_X1 U10512 ( .A1(n10363), .A2(n10364), .ZN(n10539) );
  XNOR2_X1 U10513 ( .A(n10540), .B(n10541), .ZN(n10362) );
  XNOR2_X1 U10514 ( .A(n10542), .B(n10543), .ZN(n10541) );
  NAND2_X1 U10515 ( .A1(n10364), .A2(n10363), .ZN(n10537) );
  NAND2_X1 U10516 ( .A1(n10544), .A2(n10545), .ZN(n10363) );
  NAND2_X1 U10517 ( .A1(n10359), .A2(n10546), .ZN(n10545) );
  NAND2_X1 U10518 ( .A1(n10360), .A2(n10358), .ZN(n10546) );
  NOR2_X1 U10519 ( .A1(n8053), .A2(n7624), .ZN(n10359) );
  OR2_X1 U10520 ( .A1(n10358), .A2(n10360), .ZN(n10544) );
  AND2_X1 U10521 ( .A1(n10547), .A2(n10548), .ZN(n10360) );
  NAND2_X1 U10522 ( .A1(n10549), .A2(b_22_), .ZN(n10548) );
  NOR2_X1 U10523 ( .A1(n10550), .A2(n7613), .ZN(n10549) );
  NOR2_X1 U10524 ( .A1(n10355), .A2(n10353), .ZN(n10550) );
  NAND2_X1 U10525 ( .A1(n10353), .A2(n10355), .ZN(n10547) );
  NAND2_X1 U10526 ( .A1(n10551), .A2(n10552), .ZN(n10355) );
  NAND2_X1 U10527 ( .A1(n10352), .A2(n10553), .ZN(n10552) );
  OR2_X1 U10528 ( .A1(n10351), .A2(n10349), .ZN(n10553) );
  NOR2_X1 U10529 ( .A1(n8053), .A2(n7593), .ZN(n10352) );
  NAND2_X1 U10530 ( .A1(n10349), .A2(n10351), .ZN(n10551) );
  NAND2_X1 U10531 ( .A1(n10554), .A2(n10555), .ZN(n10351) );
  NAND2_X1 U10532 ( .A1(n10556), .A2(b_22_), .ZN(n10555) );
  NOR2_X1 U10533 ( .A1(n10557), .A2(n8052), .ZN(n10556) );
  NOR2_X1 U10534 ( .A1(n10348), .A2(n10346), .ZN(n10557) );
  NAND2_X1 U10535 ( .A1(n10346), .A2(n10348), .ZN(n10554) );
  NAND2_X1 U10536 ( .A1(n10558), .A2(n10559), .ZN(n10348) );
  NAND2_X1 U10537 ( .A1(n10344), .A2(n10560), .ZN(n10559) );
  NAND2_X1 U10538 ( .A1(n10343), .A2(n10342), .ZN(n10560) );
  NOR2_X1 U10539 ( .A1(n8053), .A2(n7563), .ZN(n10344) );
  INV_X1 U10540 ( .A(b_22_), .ZN(n8053) );
  OR2_X1 U10541 ( .A1(n10342), .A2(n10343), .ZN(n10558) );
  AND2_X1 U10542 ( .A1(n10339), .A2(n10561), .ZN(n10343) );
  NAND2_X1 U10543 ( .A1(n10338), .A2(n10340), .ZN(n10561) );
  NAND2_X1 U10544 ( .A1(n10562), .A2(n10563), .ZN(n10340) );
  NAND2_X1 U10545 ( .A1(b_22_), .A2(a_28_), .ZN(n10563) );
  INV_X1 U10546 ( .A(n10564), .ZN(n10562) );
  XOR2_X1 U10547 ( .A(n10565), .B(n10566), .Z(n10338) );
  NOR2_X1 U10548 ( .A1(n7529), .A2(n7657), .ZN(n10566) );
  XOR2_X1 U10549 ( .A(n10567), .B(n10568), .Z(n10565) );
  NAND2_X1 U10550 ( .A1(a_28_), .A2(n10564), .ZN(n10339) );
  NAND2_X1 U10551 ( .A1(n10569), .A2(n10570), .ZN(n10564) );
  NAND2_X1 U10552 ( .A1(n10571), .A2(b_22_), .ZN(n10570) );
  NOR2_X1 U10553 ( .A1(n10572), .A2(n7529), .ZN(n10571) );
  NOR2_X1 U10554 ( .A1(n10325), .A2(n10326), .ZN(n10572) );
  NAND2_X1 U10555 ( .A1(n10325), .A2(n10326), .ZN(n10569) );
  NAND2_X1 U10556 ( .A1(n10573), .A2(n10574), .ZN(n10326) );
  NAND2_X1 U10557 ( .A1(n10575), .A2(b_20_), .ZN(n10574) );
  NOR2_X1 U10558 ( .A1(n10576), .A2(n8048), .ZN(n10575) );
  NOR2_X1 U10559 ( .A1(n8676), .A2(n7657), .ZN(n10576) );
  NAND2_X1 U10560 ( .A1(n10577), .A2(b_21_), .ZN(n10573) );
  NOR2_X1 U10561 ( .A1(n10578), .A2(n7515), .ZN(n10577) );
  NOR2_X1 U10562 ( .A1(n8679), .A2(n8054), .ZN(n10578) );
  AND2_X1 U10563 ( .A1(n10579), .A2(b_22_), .ZN(n10325) );
  NOR2_X1 U10564 ( .A1(n8451), .A2(n7657), .ZN(n10579) );
  XOR2_X1 U10565 ( .A(n10580), .B(n10581), .Z(n10342) );
  NAND2_X1 U10566 ( .A1(n10582), .A2(n10583), .ZN(n10580) );
  XNOR2_X1 U10567 ( .A(n10584), .B(n10585), .ZN(n10346) );
  XNOR2_X1 U10568 ( .A(n10586), .B(n10587), .ZN(n10584) );
  XOR2_X1 U10569 ( .A(n10588), .B(n10589), .Z(n10349) );
  XNOR2_X1 U10570 ( .A(n10590), .B(n10591), .ZN(n10588) );
  NAND2_X1 U10571 ( .A1(b_21_), .A2(a_26_), .ZN(n10590) );
  XNOR2_X1 U10572 ( .A(n10592), .B(n10593), .ZN(n10353) );
  XNOR2_X1 U10573 ( .A(n10594), .B(n10595), .ZN(n10592) );
  XOR2_X1 U10574 ( .A(n10596), .B(n10597), .Z(n10358) );
  XOR2_X1 U10575 ( .A(n10598), .B(n10599), .Z(n10597) );
  NAND2_X1 U10576 ( .A1(b_21_), .A2(a_24_), .ZN(n10599) );
  INV_X1 U10577 ( .A(n7639), .ZN(n10364) );
  NAND2_X1 U10578 ( .A1(b_22_), .A2(a_22_), .ZN(n7639) );
  XOR2_X1 U10579 ( .A(n10600), .B(n10601), .Z(n10365) );
  XOR2_X1 U10580 ( .A(n10602), .B(n10603), .Z(n10600) );
  NOR2_X1 U10581 ( .A1(n7645), .A2(n7657), .ZN(n10603) );
  XOR2_X1 U10582 ( .A(n10604), .B(n10605), .Z(n10369) );
  XOR2_X1 U10583 ( .A(n10606), .B(n7651), .Z(n10604) );
  XNOR2_X1 U10584 ( .A(n10607), .B(n10608), .ZN(n10374) );
  XOR2_X1 U10585 ( .A(n10609), .B(n10610), .Z(n10607) );
  NOR2_X1 U10586 ( .A1(n7676), .A2(n7657), .ZN(n10610) );
  XNOR2_X1 U10587 ( .A(n10611), .B(n10612), .ZN(n10378) );
  XNOR2_X1 U10588 ( .A(n10613), .B(n10614), .ZN(n10611) );
  XOR2_X1 U10589 ( .A(n10615), .B(n10616), .Z(n10382) );
  XOR2_X1 U10590 ( .A(n10617), .B(n10618), .Z(n10615) );
  NOR2_X1 U10591 ( .A1(n7707), .A2(n7657), .ZN(n10618) );
  XOR2_X1 U10592 ( .A(n10619), .B(n10620), .Z(n10386) );
  XOR2_X1 U10593 ( .A(n10621), .B(n10622), .Z(n10619) );
  XOR2_X1 U10594 ( .A(n10623), .B(n10624), .Z(n10390) );
  XOR2_X1 U10595 ( .A(n10625), .B(n10626), .Z(n10623) );
  NOR2_X1 U10596 ( .A1(n7743), .A2(n7657), .ZN(n10626) );
  XOR2_X1 U10597 ( .A(n10627), .B(n10628), .Z(n10393) );
  XOR2_X1 U10598 ( .A(n10629), .B(n10630), .Z(n10627) );
  XOR2_X1 U10599 ( .A(n10631), .B(n10632), .Z(n10398) );
  XOR2_X1 U10600 ( .A(n10633), .B(n10634), .Z(n10631) );
  NOR2_X1 U10601 ( .A1(n7775), .A2(n7657), .ZN(n10634) );
  XOR2_X1 U10602 ( .A(n10635), .B(n10636), .Z(n10402) );
  XOR2_X1 U10603 ( .A(n10637), .B(n10638), .Z(n10635) );
  XOR2_X1 U10604 ( .A(n10639), .B(n10640), .Z(n10406) );
  XOR2_X1 U10605 ( .A(n10641), .B(n10642), .Z(n10639) );
  NOR2_X1 U10606 ( .A1(n7806), .A2(n7657), .ZN(n10642) );
  XOR2_X1 U10607 ( .A(n10643), .B(n10644), .Z(n10410) );
  XOR2_X1 U10608 ( .A(n10645), .B(n10646), .Z(n10643) );
  XNOR2_X1 U10609 ( .A(n10647), .B(n10648), .ZN(n10414) );
  XNOR2_X1 U10610 ( .A(n10649), .B(n10650), .ZN(n10647) );
  XOR2_X1 U10611 ( .A(n10651), .B(n10652), .Z(n10418) );
  XOR2_X1 U10612 ( .A(n10653), .B(n10654), .Z(n10652) );
  NAND2_X1 U10613 ( .A1(b_21_), .A2(a_9_), .ZN(n10654) );
  XOR2_X1 U10614 ( .A(n10655), .B(n10656), .Z(n10241) );
  XNOR2_X1 U10615 ( .A(n10657), .B(n10658), .ZN(n10655) );
  NAND2_X1 U10616 ( .A1(b_21_), .A2(a_8_), .ZN(n10657) );
  XOR2_X1 U10617 ( .A(n10659), .B(n10660), .Z(n10422) );
  XOR2_X1 U10618 ( .A(n10661), .B(n10662), .Z(n10659) );
  NOR2_X1 U10619 ( .A1(n7884), .A2(n7657), .ZN(n10662) );
  XOR2_X1 U10620 ( .A(n10663), .B(n10664), .Z(n10425) );
  XOR2_X1 U10621 ( .A(n10665), .B(n10666), .Z(n10663) );
  NOR2_X1 U10622 ( .A1(n8061), .A2(n7657), .ZN(n10666) );
  XOR2_X1 U10623 ( .A(n10667), .B(n10668), .Z(n10434) );
  XOR2_X1 U10624 ( .A(n10669), .B(n10670), .Z(n10668) );
  NAND2_X1 U10625 ( .A1(b_21_), .A2(a_4_), .ZN(n10670) );
  XNOR2_X1 U10626 ( .A(n10671), .B(n10672), .ZN(n10438) );
  XOR2_X1 U10627 ( .A(n10673), .B(n10674), .Z(n10672) );
  NAND2_X1 U10628 ( .A1(b_21_), .A2(a_3_), .ZN(n10674) );
  XOR2_X1 U10629 ( .A(n10675), .B(n10676), .Z(n10441) );
  XOR2_X1 U10630 ( .A(n10677), .B(n10678), .Z(n10675) );
  NOR2_X1 U10631 ( .A1(n7965), .A2(n7657), .ZN(n10678) );
  XOR2_X1 U10632 ( .A(n10679), .B(n10680), .Z(n10446) );
  XOR2_X1 U10633 ( .A(n10681), .B(n10682), .Z(n10679) );
  NOR2_X1 U10634 ( .A1(n7973), .A2(n7657), .ZN(n10682) );
  XNOR2_X1 U10635 ( .A(n10683), .B(n10684), .ZN(n8264) );
  XNOR2_X1 U10636 ( .A(n10685), .B(n10686), .ZN(n10684) );
  OR2_X1 U10637 ( .A1(n8257), .A2(n8256), .ZN(n8131) );
  XNOR2_X1 U10638 ( .A(n8253), .B(n8252), .ZN(n8256) );
  NAND2_X1 U10639 ( .A1(n10687), .A2(n10454), .ZN(n8257) );
  NAND2_X1 U10640 ( .A1(n10688), .A2(n10689), .ZN(n10454) );
  NAND2_X1 U10641 ( .A1(n10686), .A2(n10690), .ZN(n10689) );
  OR2_X1 U10642 ( .A1(n10685), .A2(n10683), .ZN(n10690) );
  NOR2_X1 U10643 ( .A1(n7657), .A2(n8307), .ZN(n10686) );
  NAND2_X1 U10644 ( .A1(n10683), .A2(n10685), .ZN(n10688) );
  NAND2_X1 U10645 ( .A1(n10691), .A2(n10692), .ZN(n10685) );
  NAND2_X1 U10646 ( .A1(n10693), .A2(b_21_), .ZN(n10692) );
  NOR2_X1 U10647 ( .A1(n10694), .A2(n7973), .ZN(n10693) );
  NOR2_X1 U10648 ( .A1(n10680), .A2(n10681), .ZN(n10694) );
  NAND2_X1 U10649 ( .A1(n10680), .A2(n10681), .ZN(n10691) );
  NAND2_X1 U10650 ( .A1(n10695), .A2(n10696), .ZN(n10681) );
  NAND2_X1 U10651 ( .A1(n10697), .A2(b_21_), .ZN(n10696) );
  NOR2_X1 U10652 ( .A1(n10698), .A2(n7965), .ZN(n10697) );
  NOR2_X1 U10653 ( .A1(n10676), .A2(n10677), .ZN(n10698) );
  NAND2_X1 U10654 ( .A1(n10676), .A2(n10677), .ZN(n10695) );
  NAND2_X1 U10655 ( .A1(n10699), .A2(n10700), .ZN(n10677) );
  NAND2_X1 U10656 ( .A1(n10701), .A2(b_21_), .ZN(n10700) );
  NOR2_X1 U10657 ( .A1(n10702), .A2(n7945), .ZN(n10701) );
  NOR2_X1 U10658 ( .A1(n10671), .A2(n10673), .ZN(n10702) );
  NAND2_X1 U10659 ( .A1(n10671), .A2(n10673), .ZN(n10699) );
  NAND2_X1 U10660 ( .A1(n10703), .A2(n10704), .ZN(n10673) );
  NAND2_X1 U10661 ( .A1(n10705), .A2(b_21_), .ZN(n10704) );
  NOR2_X1 U10662 ( .A1(n10706), .A2(n7934), .ZN(n10705) );
  NOR2_X1 U10663 ( .A1(n10667), .A2(n10669), .ZN(n10706) );
  NAND2_X1 U10664 ( .A1(n10667), .A2(n10669), .ZN(n10703) );
  NAND2_X1 U10665 ( .A1(n10707), .A2(n10708), .ZN(n10669) );
  NAND2_X1 U10666 ( .A1(n10709), .A2(b_21_), .ZN(n10708) );
  NOR2_X1 U10667 ( .A1(n10710), .A2(n7914), .ZN(n10709) );
  NOR2_X1 U10668 ( .A1(n10475), .A2(n10476), .ZN(n10710) );
  NAND2_X1 U10669 ( .A1(n10475), .A2(n10476), .ZN(n10707) );
  NAND2_X1 U10670 ( .A1(n10711), .A2(n10712), .ZN(n10476) );
  NAND2_X1 U10671 ( .A1(n10713), .A2(b_21_), .ZN(n10712) );
  NOR2_X1 U10672 ( .A1(n10714), .A2(n8061), .ZN(n10713) );
  NOR2_X1 U10673 ( .A1(n10664), .A2(n10665), .ZN(n10714) );
  NAND2_X1 U10674 ( .A1(n10664), .A2(n10665), .ZN(n10711) );
  NAND2_X1 U10675 ( .A1(n10715), .A2(n10716), .ZN(n10665) );
  NAND2_X1 U10676 ( .A1(n10717), .A2(b_21_), .ZN(n10716) );
  NOR2_X1 U10677 ( .A1(n10718), .A2(n7884), .ZN(n10717) );
  NOR2_X1 U10678 ( .A1(n10660), .A2(n10661), .ZN(n10718) );
  NAND2_X1 U10679 ( .A1(n10660), .A2(n10661), .ZN(n10715) );
  NAND2_X1 U10680 ( .A1(n10719), .A2(n10720), .ZN(n10661) );
  NAND2_X1 U10681 ( .A1(n10721), .A2(b_21_), .ZN(n10720) );
  NOR2_X1 U10682 ( .A1(n10722), .A2(n8059), .ZN(n10721) );
  NOR2_X1 U10683 ( .A1(n10656), .A2(n10658), .ZN(n10722) );
  NAND2_X1 U10684 ( .A1(n10656), .A2(n10658), .ZN(n10719) );
  NAND2_X1 U10685 ( .A1(n10723), .A2(n10724), .ZN(n10658) );
  NAND2_X1 U10686 ( .A1(n10725), .A2(b_21_), .ZN(n10724) );
  NOR2_X1 U10687 ( .A1(n10726), .A2(n7848), .ZN(n10725) );
  NOR2_X1 U10688 ( .A1(n10651), .A2(n10653), .ZN(n10726) );
  NAND2_X1 U10689 ( .A1(n10651), .A2(n10653), .ZN(n10723) );
  NAND2_X1 U10690 ( .A1(n10727), .A2(n10728), .ZN(n10653) );
  NAND2_X1 U10691 ( .A1(n10650), .A2(n10729), .ZN(n10728) );
  NAND2_X1 U10692 ( .A1(n10649), .A2(n10648), .ZN(n10729) );
  NOR2_X1 U10693 ( .A1(n7657), .A2(n7837), .ZN(n10650) );
  OR2_X1 U10694 ( .A1(n10648), .A2(n10649), .ZN(n10727) );
  AND2_X1 U10695 ( .A1(n10730), .A2(n10731), .ZN(n10649) );
  NAND2_X1 U10696 ( .A1(n10646), .A2(n10732), .ZN(n10731) );
  OR2_X1 U10697 ( .A1(n10645), .A2(n10644), .ZN(n10732) );
  NOR2_X1 U10698 ( .A1(n7657), .A2(n7817), .ZN(n10646) );
  NAND2_X1 U10699 ( .A1(n10644), .A2(n10645), .ZN(n10730) );
  NAND2_X1 U10700 ( .A1(n10733), .A2(n10734), .ZN(n10645) );
  NAND2_X1 U10701 ( .A1(n10735), .A2(b_21_), .ZN(n10734) );
  NOR2_X1 U10702 ( .A1(n10736), .A2(n7806), .ZN(n10735) );
  NOR2_X1 U10703 ( .A1(n10640), .A2(n10641), .ZN(n10736) );
  NAND2_X1 U10704 ( .A1(n10640), .A2(n10641), .ZN(n10733) );
  NAND2_X1 U10705 ( .A1(n10737), .A2(n10738), .ZN(n10641) );
  NAND2_X1 U10706 ( .A1(n10638), .A2(n10739), .ZN(n10738) );
  OR2_X1 U10707 ( .A1(n10637), .A2(n10636), .ZN(n10739) );
  NOR2_X1 U10708 ( .A1(n7657), .A2(n7786), .ZN(n10638) );
  NAND2_X1 U10709 ( .A1(n10636), .A2(n10637), .ZN(n10737) );
  NAND2_X1 U10710 ( .A1(n10740), .A2(n10741), .ZN(n10637) );
  NAND2_X1 U10711 ( .A1(n10742), .A2(b_21_), .ZN(n10741) );
  NOR2_X1 U10712 ( .A1(n10743), .A2(n7775), .ZN(n10742) );
  NOR2_X1 U10713 ( .A1(n10632), .A2(n10633), .ZN(n10743) );
  NAND2_X1 U10714 ( .A1(n10632), .A2(n10633), .ZN(n10740) );
  NAND2_X1 U10715 ( .A1(n10744), .A2(n10745), .ZN(n10633) );
  NAND2_X1 U10716 ( .A1(n10630), .A2(n10746), .ZN(n10745) );
  OR2_X1 U10717 ( .A1(n10629), .A2(n10628), .ZN(n10746) );
  NOR2_X1 U10718 ( .A1(n7657), .A2(n7754), .ZN(n10630) );
  NAND2_X1 U10719 ( .A1(n10628), .A2(n10629), .ZN(n10744) );
  NAND2_X1 U10720 ( .A1(n10747), .A2(n10748), .ZN(n10629) );
  NAND2_X1 U10721 ( .A1(n10749), .A2(b_21_), .ZN(n10748) );
  NOR2_X1 U10722 ( .A1(n10750), .A2(n7743), .ZN(n10749) );
  NOR2_X1 U10723 ( .A1(n10624), .A2(n10625), .ZN(n10750) );
  NAND2_X1 U10724 ( .A1(n10624), .A2(n10625), .ZN(n10747) );
  NAND2_X1 U10725 ( .A1(n10751), .A2(n10752), .ZN(n10625) );
  NAND2_X1 U10726 ( .A1(n10622), .A2(n10753), .ZN(n10752) );
  OR2_X1 U10727 ( .A1(n10621), .A2(n10620), .ZN(n10753) );
  NOR2_X1 U10728 ( .A1(n7657), .A2(n7723), .ZN(n10622) );
  NAND2_X1 U10729 ( .A1(n10620), .A2(n10621), .ZN(n10751) );
  NAND2_X1 U10730 ( .A1(n10754), .A2(n10755), .ZN(n10621) );
  NAND2_X1 U10731 ( .A1(n10756), .A2(b_21_), .ZN(n10755) );
  NOR2_X1 U10732 ( .A1(n10757), .A2(n7707), .ZN(n10756) );
  NOR2_X1 U10733 ( .A1(n10616), .A2(n10617), .ZN(n10757) );
  NAND2_X1 U10734 ( .A1(n10616), .A2(n10617), .ZN(n10754) );
  NAND2_X1 U10735 ( .A1(n10758), .A2(n10759), .ZN(n10617) );
  NAND2_X1 U10736 ( .A1(n10614), .A2(n10760), .ZN(n10759) );
  NAND2_X1 U10737 ( .A1(n10613), .A2(n10612), .ZN(n10760) );
  NOR2_X1 U10738 ( .A1(n7657), .A2(n7687), .ZN(n10614) );
  OR2_X1 U10739 ( .A1(n10612), .A2(n10613), .ZN(n10758) );
  AND2_X1 U10740 ( .A1(n10761), .A2(n10762), .ZN(n10613) );
  NAND2_X1 U10741 ( .A1(n10763), .A2(b_21_), .ZN(n10762) );
  NOR2_X1 U10742 ( .A1(n10764), .A2(n7676), .ZN(n10763) );
  NOR2_X1 U10743 ( .A1(n10608), .A2(n10609), .ZN(n10764) );
  NAND2_X1 U10744 ( .A1(n10608), .A2(n10609), .ZN(n10761) );
  NAND2_X1 U10745 ( .A1(n10765), .A2(n10766), .ZN(n10609) );
  NAND2_X1 U10746 ( .A1(n7651), .A2(n10767), .ZN(n10766) );
  OR2_X1 U10747 ( .A1(n10606), .A2(n10605), .ZN(n10767) );
  INV_X1 U10748 ( .A(n8027), .ZN(n7651) );
  NAND2_X1 U10749 ( .A1(b_21_), .A2(a_21_), .ZN(n8027) );
  NAND2_X1 U10750 ( .A1(n10605), .A2(n10606), .ZN(n10765) );
  NAND2_X1 U10751 ( .A1(n10768), .A2(n10769), .ZN(n10606) );
  NAND2_X1 U10752 ( .A1(n10770), .A2(b_21_), .ZN(n10769) );
  NOR2_X1 U10753 ( .A1(n10771), .A2(n7645), .ZN(n10770) );
  NOR2_X1 U10754 ( .A1(n10601), .A2(n10602), .ZN(n10771) );
  NAND2_X1 U10755 ( .A1(n10601), .A2(n10602), .ZN(n10768) );
  NAND2_X1 U10756 ( .A1(n10772), .A2(n10773), .ZN(n10602) );
  NAND2_X1 U10757 ( .A1(n10543), .A2(n10774), .ZN(n10773) );
  OR2_X1 U10758 ( .A1(n10542), .A2(n10540), .ZN(n10774) );
  NOR2_X1 U10759 ( .A1(n7657), .A2(n7624), .ZN(n10543) );
  NAND2_X1 U10760 ( .A1(n10540), .A2(n10542), .ZN(n10772) );
  NAND2_X1 U10761 ( .A1(n10775), .A2(n10776), .ZN(n10542) );
  NAND2_X1 U10762 ( .A1(n10777), .A2(b_21_), .ZN(n10776) );
  NOR2_X1 U10763 ( .A1(n10778), .A2(n7613), .ZN(n10777) );
  NOR2_X1 U10764 ( .A1(n10596), .A2(n10598), .ZN(n10778) );
  NAND2_X1 U10765 ( .A1(n10596), .A2(n10598), .ZN(n10775) );
  NAND2_X1 U10766 ( .A1(n10779), .A2(n10780), .ZN(n10598) );
  NAND2_X1 U10767 ( .A1(n10595), .A2(n10781), .ZN(n10780) );
  NAND2_X1 U10768 ( .A1(n10594), .A2(n10593), .ZN(n10781) );
  NOR2_X1 U10769 ( .A1(n7657), .A2(n7593), .ZN(n10595) );
  OR2_X1 U10770 ( .A1(n10593), .A2(n10594), .ZN(n10779) );
  AND2_X1 U10771 ( .A1(n10782), .A2(n10783), .ZN(n10594) );
  NAND2_X1 U10772 ( .A1(n10784), .A2(b_21_), .ZN(n10783) );
  NOR2_X1 U10773 ( .A1(n10785), .A2(n8052), .ZN(n10784) );
  NOR2_X1 U10774 ( .A1(n10589), .A2(n10591), .ZN(n10785) );
  NAND2_X1 U10775 ( .A1(n10589), .A2(n10591), .ZN(n10782) );
  NAND2_X1 U10776 ( .A1(n10786), .A2(n10787), .ZN(n10591) );
  NAND2_X1 U10777 ( .A1(n10587), .A2(n10788), .ZN(n10787) );
  NAND2_X1 U10778 ( .A1(n10586), .A2(n10585), .ZN(n10788) );
  NOR2_X1 U10779 ( .A1(n7657), .A2(n7563), .ZN(n10587) );
  OR2_X1 U10780 ( .A1(n10585), .A2(n10586), .ZN(n10786) );
  AND2_X1 U10781 ( .A1(n10582), .A2(n10789), .ZN(n10586) );
  NAND2_X1 U10782 ( .A1(n10581), .A2(n10583), .ZN(n10789) );
  NAND2_X1 U10783 ( .A1(n10790), .A2(n10791), .ZN(n10583) );
  NAND2_X1 U10784 ( .A1(b_21_), .A2(a_28_), .ZN(n10791) );
  INV_X1 U10785 ( .A(n10792), .ZN(n10790) );
  XOR2_X1 U10786 ( .A(n10793), .B(n10794), .Z(n10581) );
  NOR2_X1 U10787 ( .A1(n7529), .A2(n8054), .ZN(n10794) );
  XOR2_X1 U10788 ( .A(n10795), .B(n10796), .Z(n10793) );
  NAND2_X1 U10789 ( .A1(a_28_), .A2(n10792), .ZN(n10582) );
  NAND2_X1 U10790 ( .A1(n10797), .A2(n10798), .ZN(n10792) );
  NAND2_X1 U10791 ( .A1(n10799), .A2(b_21_), .ZN(n10798) );
  NOR2_X1 U10792 ( .A1(n10800), .A2(n7529), .ZN(n10799) );
  NOR2_X1 U10793 ( .A1(n10567), .A2(n10568), .ZN(n10800) );
  NAND2_X1 U10794 ( .A1(n10567), .A2(n10568), .ZN(n10797) );
  NAND2_X1 U10795 ( .A1(n10801), .A2(n10802), .ZN(n10568) );
  NAND2_X1 U10796 ( .A1(n10803), .A2(b_19_), .ZN(n10802) );
  NOR2_X1 U10797 ( .A1(n10804), .A2(n8048), .ZN(n10803) );
  NOR2_X1 U10798 ( .A1(n8676), .A2(n8054), .ZN(n10804) );
  NAND2_X1 U10799 ( .A1(n10805), .A2(b_20_), .ZN(n10801) );
  NOR2_X1 U10800 ( .A1(n10806), .A2(n7515), .ZN(n10805) );
  NOR2_X1 U10801 ( .A1(n8679), .A2(n7688), .ZN(n10806) );
  AND2_X1 U10802 ( .A1(n10807), .A2(b_21_), .ZN(n10567) );
  NOR2_X1 U10803 ( .A1(n8451), .A2(n8054), .ZN(n10807) );
  XOR2_X1 U10804 ( .A(n10808), .B(n10809), .Z(n10585) );
  NAND2_X1 U10805 ( .A1(n10810), .A2(n10811), .ZN(n10808) );
  XNOR2_X1 U10806 ( .A(n10812), .B(n10813), .ZN(n10589) );
  XNOR2_X1 U10807 ( .A(n10814), .B(n10815), .ZN(n10812) );
  XNOR2_X1 U10808 ( .A(n10816), .B(n10817), .ZN(n10593) );
  XNOR2_X1 U10809 ( .A(n10818), .B(n10819), .ZN(n10816) );
  NAND2_X1 U10810 ( .A1(b_20_), .A2(a_26_), .ZN(n10818) );
  XNOR2_X1 U10811 ( .A(n10820), .B(n10821), .ZN(n10596) );
  XNOR2_X1 U10812 ( .A(n10822), .B(n10823), .ZN(n10820) );
  XNOR2_X1 U10813 ( .A(n10824), .B(n10825), .ZN(n10540) );
  XOR2_X1 U10814 ( .A(n10826), .B(n10827), .Z(n10825) );
  NAND2_X1 U10815 ( .A1(b_20_), .A2(a_24_), .ZN(n10827) );
  XNOR2_X1 U10816 ( .A(n10828), .B(n10829), .ZN(n10601) );
  XNOR2_X1 U10817 ( .A(n10830), .B(n10831), .ZN(n10828) );
  XOR2_X1 U10818 ( .A(n10832), .B(n10833), .Z(n10605) );
  XOR2_X1 U10819 ( .A(n10834), .B(n10835), .Z(n10832) );
  NOR2_X1 U10820 ( .A1(n7645), .A2(n8054), .ZN(n10835) );
  XNOR2_X1 U10821 ( .A(n10836), .B(n10837), .ZN(n10608) );
  XNOR2_X1 U10822 ( .A(n10838), .B(n10839), .ZN(n10836) );
  XNOR2_X1 U10823 ( .A(n10840), .B(n10841), .ZN(n10612) );
  XOR2_X1 U10824 ( .A(n10842), .B(n10843), .Z(n10840) );
  XOR2_X1 U10825 ( .A(n10844), .B(n10845), .Z(n10616) );
  XOR2_X1 U10826 ( .A(n10846), .B(n10847), .Z(n10844) );
  XOR2_X1 U10827 ( .A(n10848), .B(n10849), .Z(n10620) );
  XOR2_X1 U10828 ( .A(n10850), .B(n10851), .Z(n10848) );
  NOR2_X1 U10829 ( .A1(n7707), .A2(n8054), .ZN(n10851) );
  XNOR2_X1 U10830 ( .A(n10852), .B(n10853), .ZN(n10624) );
  XNOR2_X1 U10831 ( .A(n10854), .B(n10855), .ZN(n10853) );
  XOR2_X1 U10832 ( .A(n10856), .B(n10857), .Z(n10628) );
  XOR2_X1 U10833 ( .A(n10858), .B(n10859), .Z(n10856) );
  NOR2_X1 U10834 ( .A1(n7743), .A2(n8054), .ZN(n10859) );
  XOR2_X1 U10835 ( .A(n10860), .B(n10861), .Z(n10632) );
  XOR2_X1 U10836 ( .A(n10862), .B(n10863), .Z(n10860) );
  XOR2_X1 U10837 ( .A(n10864), .B(n10865), .Z(n10636) );
  XOR2_X1 U10838 ( .A(n10866), .B(n10867), .Z(n10864) );
  NOR2_X1 U10839 ( .A1(n7775), .A2(n8054), .ZN(n10867) );
  XOR2_X1 U10840 ( .A(n10868), .B(n10869), .Z(n10640) );
  XOR2_X1 U10841 ( .A(n10870), .B(n10871), .Z(n10868) );
  XOR2_X1 U10842 ( .A(n10872), .B(n10873), .Z(n10644) );
  XOR2_X1 U10843 ( .A(n10874), .B(n10875), .Z(n10872) );
  NOR2_X1 U10844 ( .A1(n7806), .A2(n8054), .ZN(n10875) );
  XNOR2_X1 U10845 ( .A(n10876), .B(n10877), .ZN(n10648) );
  XOR2_X1 U10846 ( .A(n10878), .B(n10879), .Z(n10876) );
  NOR2_X1 U10847 ( .A1(n7817), .A2(n8054), .ZN(n10879) );
  XNOR2_X1 U10848 ( .A(n10880), .B(n10881), .ZN(n10651) );
  XNOR2_X1 U10849 ( .A(n10882), .B(n10883), .ZN(n10880) );
  XOR2_X1 U10850 ( .A(n10884), .B(n10885), .Z(n10656) );
  XOR2_X1 U10851 ( .A(n10886), .B(n10887), .Z(n10884) );
  XNOR2_X1 U10852 ( .A(n10888), .B(n10889), .ZN(n10660) );
  XNOR2_X1 U10853 ( .A(n10890), .B(n10891), .ZN(n10889) );
  XNOR2_X1 U10854 ( .A(n10892), .B(n10893), .ZN(n10664) );
  XOR2_X1 U10855 ( .A(n10894), .B(n10895), .Z(n10893) );
  NAND2_X1 U10856 ( .A1(b_20_), .A2(a_7_), .ZN(n10895) );
  XNOR2_X1 U10857 ( .A(n10896), .B(n10897), .ZN(n10475) );
  NAND2_X1 U10858 ( .A1(n10898), .A2(n10899), .ZN(n10896) );
  XNOR2_X1 U10859 ( .A(n10900), .B(n10901), .ZN(n10667) );
  NAND2_X1 U10860 ( .A1(n10902), .A2(n10903), .ZN(n10900) );
  XOR2_X1 U10861 ( .A(n10904), .B(n10905), .Z(n10671) );
  XOR2_X1 U10862 ( .A(n10906), .B(n10907), .Z(n10904) );
  XNOR2_X1 U10863 ( .A(n10908), .B(n10909), .ZN(n10676) );
  XOR2_X1 U10864 ( .A(n10910), .B(n10911), .Z(n10909) );
  NAND2_X1 U10865 ( .A1(b_20_), .A2(a_3_), .ZN(n10911) );
  XNOR2_X1 U10866 ( .A(n10912), .B(n10913), .ZN(n10680) );
  NAND2_X1 U10867 ( .A1(n10914), .A2(n10915), .ZN(n10912) );
  XNOR2_X1 U10868 ( .A(n10916), .B(n10917), .ZN(n10683) );
  XNOR2_X1 U10869 ( .A(n10918), .B(n10919), .ZN(n10916) );
  XOR2_X1 U10870 ( .A(n10920), .B(n10455), .Z(n10687) );
  XNOR2_X1 U10871 ( .A(n10921), .B(n10922), .ZN(n10455) );
  NOR2_X1 U10872 ( .A1(n8307), .A2(n8054), .ZN(n10922) );
  INV_X1 U10873 ( .A(n10456), .ZN(n10920) );
  NAND2_X1 U10874 ( .A1(n10923), .A2(n10924), .ZN(n8141) );
  XOR2_X1 U10875 ( .A(n8246), .B(n8245), .Z(n10924) );
  AND2_X1 U10876 ( .A1(n8253), .A2(n8252), .ZN(n10923) );
  XOR2_X1 U10877 ( .A(n10925), .B(n10926), .Z(n8252) );
  XOR2_X1 U10878 ( .A(n10927), .B(n10928), .Z(n10925) );
  NOR2_X1 U10879 ( .A1(n8307), .A2(n7688), .ZN(n10928) );
  NAND2_X1 U10880 ( .A1(n10929), .A2(n10930), .ZN(n8253) );
  NAND2_X1 U10881 ( .A1(n10931), .A2(b_20_), .ZN(n10930) );
  NOR2_X1 U10882 ( .A1(n10932), .A2(n8307), .ZN(n10931) );
  NOR2_X1 U10883 ( .A1(n10456), .A2(n10921), .ZN(n10932) );
  NAND2_X1 U10884 ( .A1(n10456), .A2(n10921), .ZN(n10929) );
  NAND2_X1 U10885 ( .A1(n10933), .A2(n10934), .ZN(n10921) );
  NAND2_X1 U10886 ( .A1(n10919), .A2(n10935), .ZN(n10934) );
  NAND2_X1 U10887 ( .A1(n10918), .A2(n10917), .ZN(n10935) );
  NOR2_X1 U10888 ( .A1(n8054), .A2(n7973), .ZN(n10919) );
  OR2_X1 U10889 ( .A1(n10917), .A2(n10918), .ZN(n10933) );
  AND2_X1 U10890 ( .A1(n10914), .A2(n10936), .ZN(n10918) );
  NAND2_X1 U10891 ( .A1(n10913), .A2(n10915), .ZN(n10936) );
  NAND2_X1 U10892 ( .A1(n10937), .A2(n10938), .ZN(n10915) );
  NAND2_X1 U10893 ( .A1(b_20_), .A2(a_2_), .ZN(n10938) );
  INV_X1 U10894 ( .A(n10939), .ZN(n10937) );
  XOR2_X1 U10895 ( .A(n10940), .B(n10941), .Z(n10913) );
  XOR2_X1 U10896 ( .A(n10942), .B(n10943), .Z(n10940) );
  NOR2_X1 U10897 ( .A1(n7945), .A2(n7688), .ZN(n10943) );
  NAND2_X1 U10898 ( .A1(a_2_), .A2(n10939), .ZN(n10914) );
  NAND2_X1 U10899 ( .A1(n10944), .A2(n10945), .ZN(n10939) );
  NAND2_X1 U10900 ( .A1(n10946), .A2(b_20_), .ZN(n10945) );
  NOR2_X1 U10901 ( .A1(n10947), .A2(n7945), .ZN(n10946) );
  NOR2_X1 U10902 ( .A1(n10908), .A2(n10910), .ZN(n10947) );
  NAND2_X1 U10903 ( .A1(n10908), .A2(n10910), .ZN(n10944) );
  NAND2_X1 U10904 ( .A1(n10948), .A2(n10949), .ZN(n10910) );
  NAND2_X1 U10905 ( .A1(n10907), .A2(n10950), .ZN(n10949) );
  OR2_X1 U10906 ( .A1(n10906), .A2(n10905), .ZN(n10950) );
  NOR2_X1 U10907 ( .A1(n8054), .A2(n7934), .ZN(n10907) );
  NAND2_X1 U10908 ( .A1(n10905), .A2(n10906), .ZN(n10948) );
  NAND2_X1 U10909 ( .A1(n10902), .A2(n10951), .ZN(n10906) );
  NAND2_X1 U10910 ( .A1(n10901), .A2(n10903), .ZN(n10951) );
  NAND2_X1 U10911 ( .A1(n10952), .A2(n10953), .ZN(n10903) );
  NAND2_X1 U10912 ( .A1(b_20_), .A2(a_5_), .ZN(n10953) );
  INV_X1 U10913 ( .A(n10954), .ZN(n10952) );
  XOR2_X1 U10914 ( .A(n10955), .B(n10956), .Z(n10901) );
  XOR2_X1 U10915 ( .A(n10957), .B(n10958), .Z(n10955) );
  NOR2_X1 U10916 ( .A1(n8061), .A2(n7688), .ZN(n10958) );
  NAND2_X1 U10917 ( .A1(a_5_), .A2(n10954), .ZN(n10902) );
  NAND2_X1 U10918 ( .A1(n10898), .A2(n10959), .ZN(n10954) );
  NAND2_X1 U10919 ( .A1(n10897), .A2(n10899), .ZN(n10959) );
  NAND2_X1 U10920 ( .A1(n10960), .A2(n10961), .ZN(n10899) );
  NAND2_X1 U10921 ( .A1(b_20_), .A2(a_6_), .ZN(n10961) );
  INV_X1 U10922 ( .A(n10962), .ZN(n10960) );
  XOR2_X1 U10923 ( .A(n10963), .B(n10964), .Z(n10897) );
  XOR2_X1 U10924 ( .A(n10965), .B(n10966), .Z(n10963) );
  NOR2_X1 U10925 ( .A1(n7884), .A2(n7688), .ZN(n10966) );
  NAND2_X1 U10926 ( .A1(a_6_), .A2(n10962), .ZN(n10898) );
  NAND2_X1 U10927 ( .A1(n10967), .A2(n10968), .ZN(n10962) );
  NAND2_X1 U10928 ( .A1(n10969), .A2(b_20_), .ZN(n10968) );
  NOR2_X1 U10929 ( .A1(n10970), .A2(n7884), .ZN(n10969) );
  NOR2_X1 U10930 ( .A1(n10892), .A2(n10894), .ZN(n10970) );
  NAND2_X1 U10931 ( .A1(n10892), .A2(n10894), .ZN(n10967) );
  NAND2_X1 U10932 ( .A1(n10971), .A2(n10972), .ZN(n10894) );
  NAND2_X1 U10933 ( .A1(n10891), .A2(n10973), .ZN(n10972) );
  OR2_X1 U10934 ( .A1(n10890), .A2(n10888), .ZN(n10973) );
  NOR2_X1 U10935 ( .A1(n8054), .A2(n8059), .ZN(n10891) );
  NAND2_X1 U10936 ( .A1(n10888), .A2(n10890), .ZN(n10971) );
  NAND2_X1 U10937 ( .A1(n10974), .A2(n10975), .ZN(n10890) );
  NAND2_X1 U10938 ( .A1(n10887), .A2(n10976), .ZN(n10975) );
  OR2_X1 U10939 ( .A1(n10886), .A2(n10885), .ZN(n10976) );
  NOR2_X1 U10940 ( .A1(n8054), .A2(n7848), .ZN(n10887) );
  NAND2_X1 U10941 ( .A1(n10885), .A2(n10886), .ZN(n10974) );
  NAND2_X1 U10942 ( .A1(n10977), .A2(n10978), .ZN(n10886) );
  NAND2_X1 U10943 ( .A1(n10883), .A2(n10979), .ZN(n10978) );
  NAND2_X1 U10944 ( .A1(n10882), .A2(n10881), .ZN(n10979) );
  NOR2_X1 U10945 ( .A1(n8054), .A2(n7837), .ZN(n10883) );
  OR2_X1 U10946 ( .A1(n10881), .A2(n10882), .ZN(n10977) );
  AND2_X1 U10947 ( .A1(n10980), .A2(n10981), .ZN(n10882) );
  NAND2_X1 U10948 ( .A1(n10982), .A2(b_20_), .ZN(n10981) );
  NOR2_X1 U10949 ( .A1(n10983), .A2(n7817), .ZN(n10982) );
  NOR2_X1 U10950 ( .A1(n10877), .A2(n10878), .ZN(n10983) );
  NAND2_X1 U10951 ( .A1(n10877), .A2(n10878), .ZN(n10980) );
  NAND2_X1 U10952 ( .A1(n10984), .A2(n10985), .ZN(n10878) );
  NAND2_X1 U10953 ( .A1(n10986), .A2(b_20_), .ZN(n10985) );
  NOR2_X1 U10954 ( .A1(n10987), .A2(n7806), .ZN(n10986) );
  NOR2_X1 U10955 ( .A1(n10873), .A2(n10874), .ZN(n10987) );
  NAND2_X1 U10956 ( .A1(n10873), .A2(n10874), .ZN(n10984) );
  NAND2_X1 U10957 ( .A1(n10988), .A2(n10989), .ZN(n10874) );
  NAND2_X1 U10958 ( .A1(n10871), .A2(n10990), .ZN(n10989) );
  OR2_X1 U10959 ( .A1(n10870), .A2(n10869), .ZN(n10990) );
  NOR2_X1 U10960 ( .A1(n8054), .A2(n7786), .ZN(n10871) );
  NAND2_X1 U10961 ( .A1(n10869), .A2(n10870), .ZN(n10988) );
  NAND2_X1 U10962 ( .A1(n10991), .A2(n10992), .ZN(n10870) );
  NAND2_X1 U10963 ( .A1(n10993), .A2(b_20_), .ZN(n10992) );
  NOR2_X1 U10964 ( .A1(n10994), .A2(n7775), .ZN(n10993) );
  NOR2_X1 U10965 ( .A1(n10865), .A2(n10866), .ZN(n10994) );
  NAND2_X1 U10966 ( .A1(n10865), .A2(n10866), .ZN(n10991) );
  NAND2_X1 U10967 ( .A1(n10995), .A2(n10996), .ZN(n10866) );
  NAND2_X1 U10968 ( .A1(n10863), .A2(n10997), .ZN(n10996) );
  OR2_X1 U10969 ( .A1(n10862), .A2(n10861), .ZN(n10997) );
  NOR2_X1 U10970 ( .A1(n8054), .A2(n7754), .ZN(n10863) );
  NAND2_X1 U10971 ( .A1(n10861), .A2(n10862), .ZN(n10995) );
  NAND2_X1 U10972 ( .A1(n10998), .A2(n10999), .ZN(n10862) );
  NAND2_X1 U10973 ( .A1(n11000), .A2(b_20_), .ZN(n10999) );
  NOR2_X1 U10974 ( .A1(n11001), .A2(n7743), .ZN(n11000) );
  NOR2_X1 U10975 ( .A1(n10857), .A2(n10858), .ZN(n11001) );
  NAND2_X1 U10976 ( .A1(n10857), .A2(n10858), .ZN(n10998) );
  NAND2_X1 U10977 ( .A1(n11002), .A2(n11003), .ZN(n10858) );
  NAND2_X1 U10978 ( .A1(n10855), .A2(n11004), .ZN(n11003) );
  OR2_X1 U10979 ( .A1(n10854), .A2(n10852), .ZN(n11004) );
  NOR2_X1 U10980 ( .A1(n8054), .A2(n7723), .ZN(n10855) );
  NAND2_X1 U10981 ( .A1(n10852), .A2(n10854), .ZN(n11002) );
  NAND2_X1 U10982 ( .A1(n11005), .A2(n11006), .ZN(n10854) );
  NAND2_X1 U10983 ( .A1(n11007), .A2(b_20_), .ZN(n11006) );
  NOR2_X1 U10984 ( .A1(n11008), .A2(n7707), .ZN(n11007) );
  NOR2_X1 U10985 ( .A1(n10849), .A2(n10850), .ZN(n11008) );
  NAND2_X1 U10986 ( .A1(n10849), .A2(n10850), .ZN(n11005) );
  NAND2_X1 U10987 ( .A1(n11009), .A2(n11010), .ZN(n10850) );
  NAND2_X1 U10988 ( .A1(n10847), .A2(n11011), .ZN(n11010) );
  OR2_X1 U10989 ( .A1(n10846), .A2(n10845), .ZN(n11011) );
  NOR2_X1 U10990 ( .A1(n8054), .A2(n7687), .ZN(n10847) );
  NAND2_X1 U10991 ( .A1(n10845), .A2(n10846), .ZN(n11009) );
  NAND2_X1 U10992 ( .A1(n11012), .A2(n11013), .ZN(n10846) );
  NAND2_X1 U10993 ( .A1(n10841), .A2(n11014), .ZN(n11013) );
  OR2_X1 U10994 ( .A1(n10842), .A2(n10843), .ZN(n11014) );
  XNOR2_X1 U10995 ( .A(n11015), .B(n11016), .ZN(n10841) );
  XNOR2_X1 U10996 ( .A(n11017), .B(n11018), .ZN(n11015) );
  NAND2_X1 U10997 ( .A1(n10843), .A2(n10842), .ZN(n11012) );
  NAND2_X1 U10998 ( .A1(n11019), .A2(n11020), .ZN(n10842) );
  NAND2_X1 U10999 ( .A1(n10839), .A2(n11021), .ZN(n11020) );
  NAND2_X1 U11000 ( .A1(n10838), .A2(n10837), .ZN(n11021) );
  NOR2_X1 U11001 ( .A1(n8054), .A2(n7656), .ZN(n10839) );
  OR2_X1 U11002 ( .A1(n10837), .A2(n10838), .ZN(n11019) );
  AND2_X1 U11003 ( .A1(n11022), .A2(n11023), .ZN(n10838) );
  NAND2_X1 U11004 ( .A1(n11024), .A2(b_20_), .ZN(n11023) );
  NOR2_X1 U11005 ( .A1(n11025), .A2(n7645), .ZN(n11024) );
  NOR2_X1 U11006 ( .A1(n10833), .A2(n10834), .ZN(n11025) );
  NAND2_X1 U11007 ( .A1(n10833), .A2(n10834), .ZN(n11022) );
  NAND2_X1 U11008 ( .A1(n11026), .A2(n11027), .ZN(n10834) );
  NAND2_X1 U11009 ( .A1(n10830), .A2(n11028), .ZN(n11027) );
  NAND2_X1 U11010 ( .A1(n10831), .A2(n10829), .ZN(n11028) );
  NOR2_X1 U11011 ( .A1(n8054), .A2(n7624), .ZN(n10830) );
  OR2_X1 U11012 ( .A1(n10829), .A2(n10831), .ZN(n11026) );
  AND2_X1 U11013 ( .A1(n11029), .A2(n11030), .ZN(n10831) );
  NAND2_X1 U11014 ( .A1(n11031), .A2(b_20_), .ZN(n11030) );
  NOR2_X1 U11015 ( .A1(n11032), .A2(n7613), .ZN(n11031) );
  NOR2_X1 U11016 ( .A1(n10824), .A2(n10826), .ZN(n11032) );
  NAND2_X1 U11017 ( .A1(n10824), .A2(n10826), .ZN(n11029) );
  NAND2_X1 U11018 ( .A1(n11033), .A2(n11034), .ZN(n10826) );
  NAND2_X1 U11019 ( .A1(n10823), .A2(n11035), .ZN(n11034) );
  NAND2_X1 U11020 ( .A1(n10822), .A2(n10821), .ZN(n11035) );
  NOR2_X1 U11021 ( .A1(n8054), .A2(n7593), .ZN(n10823) );
  OR2_X1 U11022 ( .A1(n10821), .A2(n10822), .ZN(n11033) );
  AND2_X1 U11023 ( .A1(n11036), .A2(n11037), .ZN(n10822) );
  NAND2_X1 U11024 ( .A1(n11038), .A2(b_20_), .ZN(n11037) );
  NOR2_X1 U11025 ( .A1(n11039), .A2(n8052), .ZN(n11038) );
  NOR2_X1 U11026 ( .A1(n10817), .A2(n10819), .ZN(n11039) );
  NAND2_X1 U11027 ( .A1(n10817), .A2(n10819), .ZN(n11036) );
  NAND2_X1 U11028 ( .A1(n11040), .A2(n11041), .ZN(n10819) );
  NAND2_X1 U11029 ( .A1(n10815), .A2(n11042), .ZN(n11041) );
  NAND2_X1 U11030 ( .A1(n10814), .A2(n10813), .ZN(n11042) );
  NOR2_X1 U11031 ( .A1(n8054), .A2(n7563), .ZN(n10815) );
  INV_X1 U11032 ( .A(b_20_), .ZN(n8054) );
  OR2_X1 U11033 ( .A1(n10813), .A2(n10814), .ZN(n11040) );
  AND2_X1 U11034 ( .A1(n10810), .A2(n11043), .ZN(n10814) );
  NAND2_X1 U11035 ( .A1(n10809), .A2(n10811), .ZN(n11043) );
  NAND2_X1 U11036 ( .A1(n11044), .A2(n11045), .ZN(n10811) );
  NAND2_X1 U11037 ( .A1(b_20_), .A2(a_28_), .ZN(n11045) );
  INV_X1 U11038 ( .A(n11046), .ZN(n11044) );
  XOR2_X1 U11039 ( .A(n11047), .B(n11048), .Z(n10809) );
  NOR2_X1 U11040 ( .A1(n7529), .A2(n7688), .ZN(n11048) );
  XOR2_X1 U11041 ( .A(n11049), .B(n11050), .Z(n11047) );
  NAND2_X1 U11042 ( .A1(a_28_), .A2(n11046), .ZN(n10810) );
  NAND2_X1 U11043 ( .A1(n11051), .A2(n11052), .ZN(n11046) );
  NAND2_X1 U11044 ( .A1(n11053), .A2(b_20_), .ZN(n11052) );
  NOR2_X1 U11045 ( .A1(n11054), .A2(n7529), .ZN(n11053) );
  NOR2_X1 U11046 ( .A1(n10795), .A2(n10796), .ZN(n11054) );
  NAND2_X1 U11047 ( .A1(n10795), .A2(n10796), .ZN(n11051) );
  NAND2_X1 U11048 ( .A1(n11055), .A2(n11056), .ZN(n10796) );
  NAND2_X1 U11049 ( .A1(n11057), .A2(b_18_), .ZN(n11056) );
  NOR2_X1 U11050 ( .A1(n11058), .A2(n8048), .ZN(n11057) );
  NOR2_X1 U11051 ( .A1(n8676), .A2(n7688), .ZN(n11058) );
  NAND2_X1 U11052 ( .A1(n11059), .A2(b_19_), .ZN(n11055) );
  NOR2_X1 U11053 ( .A1(n11060), .A2(n7515), .ZN(n11059) );
  NOR2_X1 U11054 ( .A1(n8679), .A2(n8055), .ZN(n11060) );
  AND2_X1 U11055 ( .A1(n11061), .A2(b_20_), .ZN(n10795) );
  XOR2_X1 U11056 ( .A(n11062), .B(n11063), .Z(n10813) );
  NAND2_X1 U11057 ( .A1(n11064), .A2(n11065), .ZN(n11062) );
  XNOR2_X1 U11058 ( .A(n11066), .B(n11067), .ZN(n10817) );
  XNOR2_X1 U11059 ( .A(n11068), .B(n11069), .ZN(n11066) );
  XNOR2_X1 U11060 ( .A(n11070), .B(n11071), .ZN(n10821) );
  XNOR2_X1 U11061 ( .A(n11072), .B(n11073), .ZN(n11070) );
  NAND2_X1 U11062 ( .A1(b_19_), .A2(a_26_), .ZN(n11072) );
  XNOR2_X1 U11063 ( .A(n11074), .B(n11075), .ZN(n10824) );
  XNOR2_X1 U11064 ( .A(n11076), .B(n11077), .ZN(n11074) );
  XOR2_X1 U11065 ( .A(n11078), .B(n11079), .Z(n10829) );
  XOR2_X1 U11066 ( .A(n11080), .B(n11081), .Z(n11079) );
  NAND2_X1 U11067 ( .A1(b_19_), .A2(a_24_), .ZN(n11081) );
  XOR2_X1 U11068 ( .A(n11082), .B(n11083), .Z(n10833) );
  XOR2_X1 U11069 ( .A(n11084), .B(n11085), .Z(n11082) );
  XNOR2_X1 U11070 ( .A(n11086), .B(n11087), .ZN(n10837) );
  XOR2_X1 U11071 ( .A(n11088), .B(n11089), .Z(n11086) );
  NOR2_X1 U11072 ( .A1(n7645), .A2(n7688), .ZN(n11089) );
  INV_X1 U11073 ( .A(n7670), .ZN(n10843) );
  NAND2_X1 U11074 ( .A1(b_20_), .A2(a_20_), .ZN(n7670) );
  XOR2_X1 U11075 ( .A(n11090), .B(n11091), .Z(n10845) );
  XOR2_X1 U11076 ( .A(n11092), .B(n11093), .Z(n11090) );
  NOR2_X1 U11077 ( .A1(n7676), .A2(n7688), .ZN(n11093) );
  XNOR2_X1 U11078 ( .A(n11094), .B(n11095), .ZN(n10849) );
  XOR2_X1 U11079 ( .A(n11096), .B(n8023), .Z(n11095) );
  XOR2_X1 U11080 ( .A(n11097), .B(n11098), .Z(n10852) );
  XOR2_X1 U11081 ( .A(n11099), .B(n11100), .Z(n11097) );
  NOR2_X1 U11082 ( .A1(n7707), .A2(n7688), .ZN(n11100) );
  XOR2_X1 U11083 ( .A(n11101), .B(n11102), .Z(n10857) );
  XOR2_X1 U11084 ( .A(n11103), .B(n11104), .Z(n11101) );
  XOR2_X1 U11085 ( .A(n11105), .B(n11106), .Z(n10861) );
  XOR2_X1 U11086 ( .A(n11107), .B(n11108), .Z(n11105) );
  NOR2_X1 U11087 ( .A1(n7743), .A2(n7688), .ZN(n11108) );
  XOR2_X1 U11088 ( .A(n11109), .B(n11110), .Z(n10865) );
  XOR2_X1 U11089 ( .A(n11111), .B(n11112), .Z(n11109) );
  XNOR2_X1 U11090 ( .A(n11113), .B(n11114), .ZN(n10869) );
  XOR2_X1 U11091 ( .A(n11115), .B(n11116), .Z(n11114) );
  NAND2_X1 U11092 ( .A1(b_19_), .A2(a_14_), .ZN(n11116) );
  XOR2_X1 U11093 ( .A(n11117), .B(n11118), .Z(n10873) );
  XOR2_X1 U11094 ( .A(n11119), .B(n11120), .Z(n11117) );
  XNOR2_X1 U11095 ( .A(n11121), .B(n11122), .ZN(n10877) );
  XNOR2_X1 U11096 ( .A(n11123), .B(n11124), .ZN(n11121) );
  XOR2_X1 U11097 ( .A(n11125), .B(n11126), .Z(n10881) );
  XOR2_X1 U11098 ( .A(n11127), .B(n11128), .Z(n11126) );
  NAND2_X1 U11099 ( .A1(b_19_), .A2(a_11_), .ZN(n11128) );
  XOR2_X1 U11100 ( .A(n11129), .B(n11130), .Z(n10885) );
  XOR2_X1 U11101 ( .A(n11131), .B(n11132), .Z(n11129) );
  NOR2_X1 U11102 ( .A1(n7837), .A2(n7688), .ZN(n11132) );
  XOR2_X1 U11103 ( .A(n11133), .B(n11134), .Z(n10888) );
  XOR2_X1 U11104 ( .A(n11135), .B(n11136), .Z(n11133) );
  NOR2_X1 U11105 ( .A1(n7848), .A2(n7688), .ZN(n11136) );
  XOR2_X1 U11106 ( .A(n11137), .B(n11138), .Z(n10892) );
  XOR2_X1 U11107 ( .A(n11139), .B(n11140), .Z(n11137) );
  NOR2_X1 U11108 ( .A1(n8059), .A2(n7688), .ZN(n11140) );
  XOR2_X1 U11109 ( .A(n11141), .B(n11142), .Z(n10905) );
  XOR2_X1 U11110 ( .A(n11143), .B(n11144), .Z(n11141) );
  NOR2_X1 U11111 ( .A1(n7914), .A2(n7688), .ZN(n11144) );
  XOR2_X1 U11112 ( .A(n11145), .B(n11146), .Z(n10908) );
  XOR2_X1 U11113 ( .A(n11147), .B(n11148), .Z(n11145) );
  NOR2_X1 U11114 ( .A1(n7934), .A2(n7688), .ZN(n11148) );
  XOR2_X1 U11115 ( .A(n11149), .B(n11150), .Z(n10917) );
  NAND2_X1 U11116 ( .A1(n11151), .A2(n11152), .ZN(n11149) );
  XOR2_X1 U11117 ( .A(n11153), .B(n11154), .Z(n10456) );
  XOR2_X1 U11118 ( .A(n11155), .B(n11156), .Z(n11153) );
  NOR2_X1 U11119 ( .A1(n7973), .A2(n7688), .ZN(n11156) );
  NAND2_X1 U11120 ( .A1(n11157), .A2(n11158), .ZN(n8146) );
  XOR2_X1 U11121 ( .A(n8247), .B(n8248), .Z(n11158) );
  AND2_X1 U11122 ( .A1(n8246), .A2(n8245), .ZN(n11157) );
  INV_X1 U11123 ( .A(n8254), .ZN(n8245) );
  XOR2_X1 U11124 ( .A(n11159), .B(n11160), .Z(n8254) );
  XOR2_X1 U11125 ( .A(n11161), .B(n11162), .Z(n11160) );
  NAND2_X1 U11126 ( .A1(b_18_), .A2(a_0_), .ZN(n11162) );
  NAND2_X1 U11127 ( .A1(n11163), .A2(n11164), .ZN(n8246) );
  NAND2_X1 U11128 ( .A1(n11165), .A2(b_19_), .ZN(n11164) );
  NOR2_X1 U11129 ( .A1(n11166), .A2(n8307), .ZN(n11165) );
  NOR2_X1 U11130 ( .A1(n10926), .A2(n10927), .ZN(n11166) );
  NAND2_X1 U11131 ( .A1(n10926), .A2(n10927), .ZN(n11163) );
  NAND2_X1 U11132 ( .A1(n11167), .A2(n11168), .ZN(n10927) );
  NAND2_X1 U11133 ( .A1(n11169), .A2(b_19_), .ZN(n11168) );
  NOR2_X1 U11134 ( .A1(n11170), .A2(n7973), .ZN(n11169) );
  NOR2_X1 U11135 ( .A1(n11154), .A2(n11155), .ZN(n11170) );
  NAND2_X1 U11136 ( .A1(n11154), .A2(n11155), .ZN(n11167) );
  NAND2_X1 U11137 ( .A1(n11151), .A2(n11171), .ZN(n11155) );
  NAND2_X1 U11138 ( .A1(n11150), .A2(n11152), .ZN(n11171) );
  NAND2_X1 U11139 ( .A1(n11172), .A2(n11173), .ZN(n11152) );
  NAND2_X1 U11140 ( .A1(b_19_), .A2(a_2_), .ZN(n11173) );
  INV_X1 U11141 ( .A(n11174), .ZN(n11172) );
  XNOR2_X1 U11142 ( .A(n11175), .B(n11176), .ZN(n11150) );
  NAND2_X1 U11143 ( .A1(n11177), .A2(n11178), .ZN(n11175) );
  NAND2_X1 U11144 ( .A1(a_2_), .A2(n11174), .ZN(n11151) );
  NAND2_X1 U11145 ( .A1(n11179), .A2(n11180), .ZN(n11174) );
  NAND2_X1 U11146 ( .A1(n11181), .A2(b_19_), .ZN(n11180) );
  NOR2_X1 U11147 ( .A1(n11182), .A2(n7945), .ZN(n11181) );
  NOR2_X1 U11148 ( .A1(n10941), .A2(n10942), .ZN(n11182) );
  NAND2_X1 U11149 ( .A1(n10941), .A2(n10942), .ZN(n11179) );
  NAND2_X1 U11150 ( .A1(n11183), .A2(n11184), .ZN(n10942) );
  NAND2_X1 U11151 ( .A1(n11185), .A2(b_19_), .ZN(n11184) );
  NOR2_X1 U11152 ( .A1(n11186), .A2(n7934), .ZN(n11185) );
  NOR2_X1 U11153 ( .A1(n11146), .A2(n11147), .ZN(n11186) );
  NAND2_X1 U11154 ( .A1(n11146), .A2(n11147), .ZN(n11183) );
  NAND2_X1 U11155 ( .A1(n11187), .A2(n11188), .ZN(n11147) );
  NAND2_X1 U11156 ( .A1(n11189), .A2(b_19_), .ZN(n11188) );
  NOR2_X1 U11157 ( .A1(n11190), .A2(n7914), .ZN(n11189) );
  NOR2_X1 U11158 ( .A1(n11142), .A2(n11143), .ZN(n11190) );
  NAND2_X1 U11159 ( .A1(n11142), .A2(n11143), .ZN(n11187) );
  NAND2_X1 U11160 ( .A1(n11191), .A2(n11192), .ZN(n11143) );
  NAND2_X1 U11161 ( .A1(n11193), .A2(b_19_), .ZN(n11192) );
  NOR2_X1 U11162 ( .A1(n11194), .A2(n8061), .ZN(n11193) );
  NOR2_X1 U11163 ( .A1(n10956), .A2(n10957), .ZN(n11194) );
  NAND2_X1 U11164 ( .A1(n10956), .A2(n10957), .ZN(n11191) );
  NAND2_X1 U11165 ( .A1(n11195), .A2(n11196), .ZN(n10957) );
  NAND2_X1 U11166 ( .A1(n11197), .A2(b_19_), .ZN(n11196) );
  NOR2_X1 U11167 ( .A1(n11198), .A2(n7884), .ZN(n11197) );
  NOR2_X1 U11168 ( .A1(n10964), .A2(n10965), .ZN(n11198) );
  NAND2_X1 U11169 ( .A1(n10964), .A2(n10965), .ZN(n11195) );
  NAND2_X1 U11170 ( .A1(n11199), .A2(n11200), .ZN(n10965) );
  NAND2_X1 U11171 ( .A1(n11201), .A2(b_19_), .ZN(n11200) );
  NOR2_X1 U11172 ( .A1(n11202), .A2(n8059), .ZN(n11201) );
  NOR2_X1 U11173 ( .A1(n11138), .A2(n11139), .ZN(n11202) );
  NAND2_X1 U11174 ( .A1(n11138), .A2(n11139), .ZN(n11199) );
  NAND2_X1 U11175 ( .A1(n11203), .A2(n11204), .ZN(n11139) );
  NAND2_X1 U11176 ( .A1(n11205), .A2(b_19_), .ZN(n11204) );
  NOR2_X1 U11177 ( .A1(n11206), .A2(n7848), .ZN(n11205) );
  NOR2_X1 U11178 ( .A1(n11134), .A2(n11135), .ZN(n11206) );
  NAND2_X1 U11179 ( .A1(n11134), .A2(n11135), .ZN(n11203) );
  NAND2_X1 U11180 ( .A1(n11207), .A2(n11208), .ZN(n11135) );
  NAND2_X1 U11181 ( .A1(n11209), .A2(b_19_), .ZN(n11208) );
  NOR2_X1 U11182 ( .A1(n11210), .A2(n7837), .ZN(n11209) );
  NOR2_X1 U11183 ( .A1(n11130), .A2(n11131), .ZN(n11210) );
  NAND2_X1 U11184 ( .A1(n11130), .A2(n11131), .ZN(n11207) );
  NAND2_X1 U11185 ( .A1(n11211), .A2(n11212), .ZN(n11131) );
  NAND2_X1 U11186 ( .A1(n11213), .A2(b_19_), .ZN(n11212) );
  NOR2_X1 U11187 ( .A1(n11214), .A2(n7817), .ZN(n11213) );
  NOR2_X1 U11188 ( .A1(n11125), .A2(n11127), .ZN(n11214) );
  NAND2_X1 U11189 ( .A1(n11125), .A2(n11127), .ZN(n11211) );
  NAND2_X1 U11190 ( .A1(n11215), .A2(n11216), .ZN(n11127) );
  NAND2_X1 U11191 ( .A1(n11124), .A2(n11217), .ZN(n11216) );
  NAND2_X1 U11192 ( .A1(n11123), .A2(n11122), .ZN(n11217) );
  NOR2_X1 U11193 ( .A1(n7688), .A2(n7806), .ZN(n11124) );
  OR2_X1 U11194 ( .A1(n11122), .A2(n11123), .ZN(n11215) );
  AND2_X1 U11195 ( .A1(n11218), .A2(n11219), .ZN(n11123) );
  NAND2_X1 U11196 ( .A1(n11120), .A2(n11220), .ZN(n11219) );
  OR2_X1 U11197 ( .A1(n11119), .A2(n11118), .ZN(n11220) );
  NOR2_X1 U11198 ( .A1(n7688), .A2(n7786), .ZN(n11120) );
  NAND2_X1 U11199 ( .A1(n11118), .A2(n11119), .ZN(n11218) );
  NAND2_X1 U11200 ( .A1(n11221), .A2(n11222), .ZN(n11119) );
  NAND2_X1 U11201 ( .A1(n11223), .A2(b_19_), .ZN(n11222) );
  NOR2_X1 U11202 ( .A1(n11224), .A2(n7775), .ZN(n11223) );
  NOR2_X1 U11203 ( .A1(n11113), .A2(n11115), .ZN(n11224) );
  NAND2_X1 U11204 ( .A1(n11113), .A2(n11115), .ZN(n11221) );
  NAND2_X1 U11205 ( .A1(n11225), .A2(n11226), .ZN(n11115) );
  NAND2_X1 U11206 ( .A1(n11112), .A2(n11227), .ZN(n11226) );
  OR2_X1 U11207 ( .A1(n11111), .A2(n11110), .ZN(n11227) );
  NOR2_X1 U11208 ( .A1(n7688), .A2(n7754), .ZN(n11112) );
  NAND2_X1 U11209 ( .A1(n11110), .A2(n11111), .ZN(n11225) );
  NAND2_X1 U11210 ( .A1(n11228), .A2(n11229), .ZN(n11111) );
  NAND2_X1 U11211 ( .A1(n11230), .A2(b_19_), .ZN(n11229) );
  NOR2_X1 U11212 ( .A1(n11231), .A2(n7743), .ZN(n11230) );
  NOR2_X1 U11213 ( .A1(n11106), .A2(n11107), .ZN(n11231) );
  NAND2_X1 U11214 ( .A1(n11106), .A2(n11107), .ZN(n11228) );
  NAND2_X1 U11215 ( .A1(n11232), .A2(n11233), .ZN(n11107) );
  NAND2_X1 U11216 ( .A1(n11104), .A2(n11234), .ZN(n11233) );
  OR2_X1 U11217 ( .A1(n11103), .A2(n11102), .ZN(n11234) );
  NOR2_X1 U11218 ( .A1(n7688), .A2(n7723), .ZN(n11104) );
  NAND2_X1 U11219 ( .A1(n11102), .A2(n11103), .ZN(n11232) );
  NAND2_X1 U11220 ( .A1(n11235), .A2(n11236), .ZN(n11103) );
  NAND2_X1 U11221 ( .A1(n11237), .A2(b_19_), .ZN(n11236) );
  NOR2_X1 U11222 ( .A1(n11238), .A2(n7707), .ZN(n11237) );
  NOR2_X1 U11223 ( .A1(n11098), .A2(n11099), .ZN(n11238) );
  NAND2_X1 U11224 ( .A1(n11098), .A2(n11099), .ZN(n11235) );
  NAND2_X1 U11225 ( .A1(n11239), .A2(n11240), .ZN(n11099) );
  NAND2_X1 U11226 ( .A1(n7682), .A2(n11241), .ZN(n11240) );
  OR2_X1 U11227 ( .A1(n11096), .A2(n11094), .ZN(n11241) );
  INV_X1 U11228 ( .A(n8023), .ZN(n7682) );
  NAND2_X1 U11229 ( .A1(b_19_), .A2(a_19_), .ZN(n8023) );
  NAND2_X1 U11230 ( .A1(n11094), .A2(n11096), .ZN(n11239) );
  NAND2_X1 U11231 ( .A1(n11242), .A2(n11243), .ZN(n11096) );
  NAND2_X1 U11232 ( .A1(n11244), .A2(b_19_), .ZN(n11243) );
  NOR2_X1 U11233 ( .A1(n11245), .A2(n7676), .ZN(n11244) );
  NOR2_X1 U11234 ( .A1(n11091), .A2(n11092), .ZN(n11245) );
  NAND2_X1 U11235 ( .A1(n11091), .A2(n11092), .ZN(n11242) );
  NAND2_X1 U11236 ( .A1(n11246), .A2(n11247), .ZN(n11092) );
  NAND2_X1 U11237 ( .A1(n11018), .A2(n11248), .ZN(n11247) );
  NAND2_X1 U11238 ( .A1(n11017), .A2(n11016), .ZN(n11248) );
  NOR2_X1 U11239 ( .A1(n7688), .A2(n7656), .ZN(n11018) );
  OR2_X1 U11240 ( .A1(n11016), .A2(n11017), .ZN(n11246) );
  AND2_X1 U11241 ( .A1(n11249), .A2(n11250), .ZN(n11017) );
  NAND2_X1 U11242 ( .A1(n11251), .A2(b_19_), .ZN(n11250) );
  NOR2_X1 U11243 ( .A1(n11252), .A2(n7645), .ZN(n11251) );
  NOR2_X1 U11244 ( .A1(n11087), .A2(n11088), .ZN(n11252) );
  NAND2_X1 U11245 ( .A1(n11087), .A2(n11088), .ZN(n11249) );
  NAND2_X1 U11246 ( .A1(n11253), .A2(n11254), .ZN(n11088) );
  NAND2_X1 U11247 ( .A1(n11085), .A2(n11255), .ZN(n11254) );
  OR2_X1 U11248 ( .A1(n11084), .A2(n11083), .ZN(n11255) );
  NOR2_X1 U11249 ( .A1(n7688), .A2(n7624), .ZN(n11085) );
  NAND2_X1 U11250 ( .A1(n11083), .A2(n11084), .ZN(n11253) );
  NAND2_X1 U11251 ( .A1(n11256), .A2(n11257), .ZN(n11084) );
  NAND2_X1 U11252 ( .A1(n11258), .A2(b_19_), .ZN(n11257) );
  NOR2_X1 U11253 ( .A1(n11259), .A2(n7613), .ZN(n11258) );
  NOR2_X1 U11254 ( .A1(n11078), .A2(n11080), .ZN(n11259) );
  NAND2_X1 U11255 ( .A1(n11078), .A2(n11080), .ZN(n11256) );
  NAND2_X1 U11256 ( .A1(n11260), .A2(n11261), .ZN(n11080) );
  NAND2_X1 U11257 ( .A1(n11077), .A2(n11262), .ZN(n11261) );
  NAND2_X1 U11258 ( .A1(n11076), .A2(n11075), .ZN(n11262) );
  NOR2_X1 U11259 ( .A1(n7688), .A2(n7593), .ZN(n11077) );
  OR2_X1 U11260 ( .A1(n11075), .A2(n11076), .ZN(n11260) );
  AND2_X1 U11261 ( .A1(n11263), .A2(n11264), .ZN(n11076) );
  NAND2_X1 U11262 ( .A1(n11265), .A2(b_19_), .ZN(n11264) );
  NOR2_X1 U11263 ( .A1(n11266), .A2(n8052), .ZN(n11265) );
  NOR2_X1 U11264 ( .A1(n11071), .A2(n11073), .ZN(n11266) );
  NAND2_X1 U11265 ( .A1(n11071), .A2(n11073), .ZN(n11263) );
  NAND2_X1 U11266 ( .A1(n11267), .A2(n11268), .ZN(n11073) );
  NAND2_X1 U11267 ( .A1(n11069), .A2(n11269), .ZN(n11268) );
  NAND2_X1 U11268 ( .A1(n11068), .A2(n11067), .ZN(n11269) );
  NOR2_X1 U11269 ( .A1(n7688), .A2(n7563), .ZN(n11069) );
  OR2_X1 U11270 ( .A1(n11067), .A2(n11068), .ZN(n11267) );
  AND2_X1 U11271 ( .A1(n11064), .A2(n11270), .ZN(n11068) );
  NAND2_X1 U11272 ( .A1(n11063), .A2(n11065), .ZN(n11270) );
  NAND2_X1 U11273 ( .A1(n11271), .A2(n11272), .ZN(n11065) );
  NAND2_X1 U11274 ( .A1(b_19_), .A2(a_28_), .ZN(n11272) );
  INV_X1 U11275 ( .A(n11273), .ZN(n11271) );
  XOR2_X1 U11276 ( .A(n11274), .B(n11275), .Z(n11063) );
  NOR2_X1 U11277 ( .A1(n7529), .A2(n8055), .ZN(n11275) );
  XOR2_X1 U11278 ( .A(n11276), .B(n11277), .Z(n11274) );
  NAND2_X1 U11279 ( .A1(a_28_), .A2(n11273), .ZN(n11064) );
  NAND2_X1 U11280 ( .A1(n11278), .A2(n11279), .ZN(n11273) );
  NAND2_X1 U11281 ( .A1(n11280), .A2(b_19_), .ZN(n11279) );
  NOR2_X1 U11282 ( .A1(n11281), .A2(n7529), .ZN(n11280) );
  NOR2_X1 U11283 ( .A1(n11049), .A2(n11050), .ZN(n11281) );
  NAND2_X1 U11284 ( .A1(n11049), .A2(n11050), .ZN(n11278) );
  NAND2_X1 U11285 ( .A1(n11282), .A2(n11283), .ZN(n11050) );
  NAND2_X1 U11286 ( .A1(n11284), .A2(b_17_), .ZN(n11283) );
  NOR2_X1 U11287 ( .A1(n11285), .A2(n8048), .ZN(n11284) );
  NOR2_X1 U11288 ( .A1(n8676), .A2(n8055), .ZN(n11285) );
  NAND2_X1 U11289 ( .A1(n11286), .A2(b_18_), .ZN(n11282) );
  NOR2_X1 U11290 ( .A1(n11287), .A2(n7515), .ZN(n11286) );
  NOR2_X1 U11291 ( .A1(n8679), .A2(n7724), .ZN(n11287) );
  AND2_X1 U11292 ( .A1(n11061), .A2(b_18_), .ZN(n11049) );
  NOR2_X1 U11293 ( .A1(n8451), .A2(n7688), .ZN(n11061) );
  XOR2_X1 U11294 ( .A(n11288), .B(n11289), .Z(n11067) );
  NAND2_X1 U11295 ( .A1(n11290), .A2(n11291), .ZN(n11288) );
  XNOR2_X1 U11296 ( .A(n11292), .B(n11293), .ZN(n11071) );
  XNOR2_X1 U11297 ( .A(n11294), .B(n11295), .ZN(n11292) );
  XNOR2_X1 U11298 ( .A(n11296), .B(n11297), .ZN(n11075) );
  XNOR2_X1 U11299 ( .A(n11298), .B(n11299), .ZN(n11296) );
  NAND2_X1 U11300 ( .A1(b_18_), .A2(a_26_), .ZN(n11298) );
  XNOR2_X1 U11301 ( .A(n11300), .B(n11301), .ZN(n11078) );
  XOR2_X1 U11302 ( .A(n11302), .B(n11303), .Z(n11301) );
  NAND2_X1 U11303 ( .A1(b_18_), .A2(a_25_), .ZN(n11303) );
  XNOR2_X1 U11304 ( .A(n11304), .B(n11305), .ZN(n11083) );
  NAND2_X1 U11305 ( .A1(n11306), .A2(n11307), .ZN(n11304) );
  XNOR2_X1 U11306 ( .A(n11308), .B(n11309), .ZN(n11087) );
  XNOR2_X1 U11307 ( .A(n11310), .B(n11311), .ZN(n11308) );
  XOR2_X1 U11308 ( .A(n11312), .B(n11313), .Z(n11016) );
  XOR2_X1 U11309 ( .A(n11314), .B(n11315), .Z(n11313) );
  NAND2_X1 U11310 ( .A1(b_18_), .A2(a_22_), .ZN(n11315) );
  XOR2_X1 U11311 ( .A(n11316), .B(n11317), .Z(n11091) );
  XOR2_X1 U11312 ( .A(n11318), .B(n11319), .Z(n11316) );
  XOR2_X1 U11313 ( .A(n11320), .B(n11321), .Z(n11094) );
  XOR2_X1 U11314 ( .A(n11322), .B(n11323), .Z(n11320) );
  NOR2_X1 U11315 ( .A1(n7676), .A2(n8055), .ZN(n11323) );
  XOR2_X1 U11316 ( .A(n11324), .B(n11325), .Z(n11098) );
  XOR2_X1 U11317 ( .A(n11326), .B(n11327), .Z(n11324) );
  XOR2_X1 U11318 ( .A(n11328), .B(n11329), .Z(n11102) );
  XOR2_X1 U11319 ( .A(n11330), .B(n11331), .Z(n11328) );
  XOR2_X1 U11320 ( .A(n11332), .B(n11333), .Z(n11106) );
  XOR2_X1 U11321 ( .A(n11334), .B(n11335), .Z(n11332) );
  XNOR2_X1 U11322 ( .A(n11336), .B(n11337), .ZN(n11110) );
  XOR2_X1 U11323 ( .A(n11338), .B(n11339), .Z(n11337) );
  NAND2_X1 U11324 ( .A1(b_18_), .A2(a_16_), .ZN(n11339) );
  XOR2_X1 U11325 ( .A(n11340), .B(n11341), .Z(n11113) );
  XOR2_X1 U11326 ( .A(n11342), .B(n11343), .Z(n11340) );
  XNOR2_X1 U11327 ( .A(n11344), .B(n11345), .ZN(n11118) );
  XOR2_X1 U11328 ( .A(n11346), .B(n11347), .Z(n11345) );
  NAND2_X1 U11329 ( .A1(b_18_), .A2(a_14_), .ZN(n11347) );
  XNOR2_X1 U11330 ( .A(n11348), .B(n11349), .ZN(n11122) );
  XOR2_X1 U11331 ( .A(n11350), .B(n11351), .Z(n11348) );
  NOR2_X1 U11332 ( .A1(n7786), .A2(n8055), .ZN(n11351) );
  XNOR2_X1 U11333 ( .A(n11352), .B(n11353), .ZN(n11125) );
  XNOR2_X1 U11334 ( .A(n11354), .B(n11355), .ZN(n11352) );
  XOR2_X1 U11335 ( .A(n11356), .B(n11357), .Z(n11130) );
  XOR2_X1 U11336 ( .A(n11358), .B(n11359), .Z(n11356) );
  XOR2_X1 U11337 ( .A(n11360), .B(n11361), .Z(n11134) );
  XOR2_X1 U11338 ( .A(n11362), .B(n11363), .Z(n11360) );
  XOR2_X1 U11339 ( .A(n11364), .B(n11365), .Z(n11138) );
  XOR2_X1 U11340 ( .A(n11366), .B(n11367), .Z(n11364) );
  NOR2_X1 U11341 ( .A1(n7848), .A2(n8055), .ZN(n11367) );
  XNOR2_X1 U11342 ( .A(n11368), .B(n11369), .ZN(n10964) );
  NAND2_X1 U11343 ( .A1(n11370), .A2(n11371), .ZN(n11368) );
  XNOR2_X1 U11344 ( .A(n11372), .B(n11373), .ZN(n10956) );
  NAND2_X1 U11345 ( .A1(n11374), .A2(n11375), .ZN(n11372) );
  XOR2_X1 U11346 ( .A(n11376), .B(n11377), .Z(n11142) );
  XOR2_X1 U11347 ( .A(n11378), .B(n11379), .Z(n11376) );
  XOR2_X1 U11348 ( .A(n11380), .B(n11381), .Z(n11146) );
  XOR2_X1 U11349 ( .A(n11382), .B(n11383), .Z(n11380) );
  NOR2_X1 U11350 ( .A1(n7914), .A2(n8055), .ZN(n11383) );
  XNOR2_X1 U11351 ( .A(n11384), .B(n11385), .ZN(n10941) );
  NAND2_X1 U11352 ( .A1(n11386), .A2(n11387), .ZN(n11384) );
  XNOR2_X1 U11353 ( .A(n11388), .B(n11389), .ZN(n11154) );
  NAND2_X1 U11354 ( .A1(n11390), .A2(n11391), .ZN(n11388) );
  XNOR2_X1 U11355 ( .A(n11392), .B(n11393), .ZN(n10926) );
  XNOR2_X1 U11356 ( .A(n11394), .B(n11395), .ZN(n11393) );
  NAND2_X1 U11357 ( .A1(n11396), .A2(n11397), .ZN(n8152) );
  NAND2_X1 U11358 ( .A1(n8248), .A2(n8247), .ZN(n11397) );
  XOR2_X1 U11359 ( .A(n8238), .B(n11398), .Z(n11396) );
  NAND2_X1 U11360 ( .A1(n11399), .A2(n11400), .ZN(n8151) );
  XOR2_X1 U11361 ( .A(n8238), .B(n8237), .Z(n11400) );
  AND2_X1 U11362 ( .A1(n8247), .A2(n8248), .ZN(n11399) );
  XNOR2_X1 U11363 ( .A(n11401), .B(n11402), .ZN(n8248) );
  XOR2_X1 U11364 ( .A(n11403), .B(n11404), .Z(n11402) );
  NAND2_X1 U11365 ( .A1(b_17_), .A2(a_0_), .ZN(n11404) );
  NAND2_X1 U11366 ( .A1(n11405), .A2(n11406), .ZN(n8247) );
  NAND2_X1 U11367 ( .A1(n11407), .A2(b_18_), .ZN(n11406) );
  NOR2_X1 U11368 ( .A1(n11408), .A2(n8307), .ZN(n11407) );
  NOR2_X1 U11369 ( .A1(n11159), .A2(n11161), .ZN(n11408) );
  NAND2_X1 U11370 ( .A1(n11159), .A2(n11161), .ZN(n11405) );
  NAND2_X1 U11371 ( .A1(n11409), .A2(n11410), .ZN(n11161) );
  NAND2_X1 U11372 ( .A1(n11395), .A2(n11411), .ZN(n11410) );
  OR2_X1 U11373 ( .A1(n11392), .A2(n11394), .ZN(n11411) );
  NOR2_X1 U11374 ( .A1(n8055), .A2(n7973), .ZN(n11395) );
  NAND2_X1 U11375 ( .A1(n11392), .A2(n11394), .ZN(n11409) );
  NAND2_X1 U11376 ( .A1(n11390), .A2(n11412), .ZN(n11394) );
  NAND2_X1 U11377 ( .A1(n11389), .A2(n11391), .ZN(n11412) );
  NAND2_X1 U11378 ( .A1(n11413), .A2(n11414), .ZN(n11391) );
  NAND2_X1 U11379 ( .A1(b_18_), .A2(a_2_), .ZN(n11414) );
  INV_X1 U11380 ( .A(n11415), .ZN(n11413) );
  XOR2_X1 U11381 ( .A(n11416), .B(n11417), .Z(n11389) );
  XOR2_X1 U11382 ( .A(n11418), .B(n11419), .Z(n11416) );
  NOR2_X1 U11383 ( .A1(n7945), .A2(n7724), .ZN(n11419) );
  NAND2_X1 U11384 ( .A1(a_2_), .A2(n11415), .ZN(n11390) );
  NAND2_X1 U11385 ( .A1(n11177), .A2(n11420), .ZN(n11415) );
  NAND2_X1 U11386 ( .A1(n11176), .A2(n11178), .ZN(n11420) );
  NAND2_X1 U11387 ( .A1(n11421), .A2(n11422), .ZN(n11178) );
  NAND2_X1 U11388 ( .A1(b_18_), .A2(a_3_), .ZN(n11422) );
  INV_X1 U11389 ( .A(n11423), .ZN(n11421) );
  XOR2_X1 U11390 ( .A(n11424), .B(n11425), .Z(n11176) );
  XOR2_X1 U11391 ( .A(n11426), .B(n11427), .Z(n11424) );
  NOR2_X1 U11392 ( .A1(n7934), .A2(n7724), .ZN(n11427) );
  NAND2_X1 U11393 ( .A1(a_3_), .A2(n11423), .ZN(n11177) );
  NAND2_X1 U11394 ( .A1(n11386), .A2(n11428), .ZN(n11423) );
  NAND2_X1 U11395 ( .A1(n11385), .A2(n11387), .ZN(n11428) );
  NAND2_X1 U11396 ( .A1(n11429), .A2(n11430), .ZN(n11387) );
  NAND2_X1 U11397 ( .A1(b_18_), .A2(a_4_), .ZN(n11430) );
  INV_X1 U11398 ( .A(n11431), .ZN(n11429) );
  XOR2_X1 U11399 ( .A(n11432), .B(n11433), .Z(n11385) );
  XOR2_X1 U11400 ( .A(n11434), .B(n11435), .Z(n11432) );
  NOR2_X1 U11401 ( .A1(n7914), .A2(n7724), .ZN(n11435) );
  NAND2_X1 U11402 ( .A1(a_4_), .A2(n11431), .ZN(n11386) );
  NAND2_X1 U11403 ( .A1(n11436), .A2(n11437), .ZN(n11431) );
  NAND2_X1 U11404 ( .A1(n11438), .A2(b_18_), .ZN(n11437) );
  NOR2_X1 U11405 ( .A1(n11439), .A2(n7914), .ZN(n11438) );
  NOR2_X1 U11406 ( .A1(n11382), .A2(n11381), .ZN(n11439) );
  NAND2_X1 U11407 ( .A1(n11381), .A2(n11382), .ZN(n11436) );
  NAND2_X1 U11408 ( .A1(n11440), .A2(n11441), .ZN(n11382) );
  NAND2_X1 U11409 ( .A1(n11379), .A2(n11442), .ZN(n11441) );
  OR2_X1 U11410 ( .A1(n11377), .A2(n11378), .ZN(n11442) );
  NOR2_X1 U11411 ( .A1(n8055), .A2(n8061), .ZN(n11379) );
  NAND2_X1 U11412 ( .A1(n11377), .A2(n11378), .ZN(n11440) );
  NAND2_X1 U11413 ( .A1(n11374), .A2(n11443), .ZN(n11378) );
  NAND2_X1 U11414 ( .A1(n11373), .A2(n11375), .ZN(n11443) );
  NAND2_X1 U11415 ( .A1(n11444), .A2(n11445), .ZN(n11375) );
  NAND2_X1 U11416 ( .A1(b_18_), .A2(a_7_), .ZN(n11445) );
  INV_X1 U11417 ( .A(n11446), .ZN(n11444) );
  XNOR2_X1 U11418 ( .A(n11447), .B(n11448), .ZN(n11373) );
  XOR2_X1 U11419 ( .A(n11449), .B(n11450), .Z(n11448) );
  NAND2_X1 U11420 ( .A1(b_17_), .A2(a_8_), .ZN(n11450) );
  NAND2_X1 U11421 ( .A1(a_7_), .A2(n11446), .ZN(n11374) );
  NAND2_X1 U11422 ( .A1(n11370), .A2(n11451), .ZN(n11446) );
  NAND2_X1 U11423 ( .A1(n11369), .A2(n11371), .ZN(n11451) );
  NAND2_X1 U11424 ( .A1(n11452), .A2(n11453), .ZN(n11371) );
  NAND2_X1 U11425 ( .A1(b_18_), .A2(a_8_), .ZN(n11453) );
  INV_X1 U11426 ( .A(n11454), .ZN(n11452) );
  XOR2_X1 U11427 ( .A(n11455), .B(n11456), .Z(n11369) );
  XOR2_X1 U11428 ( .A(n11457), .B(n11458), .Z(n11455) );
  NOR2_X1 U11429 ( .A1(n7848), .A2(n7724), .ZN(n11458) );
  NAND2_X1 U11430 ( .A1(a_8_), .A2(n11454), .ZN(n11370) );
  NAND2_X1 U11431 ( .A1(n11459), .A2(n11460), .ZN(n11454) );
  NAND2_X1 U11432 ( .A1(n11461), .A2(b_18_), .ZN(n11460) );
  NOR2_X1 U11433 ( .A1(n11462), .A2(n7848), .ZN(n11461) );
  NOR2_X1 U11434 ( .A1(n11365), .A2(n11366), .ZN(n11462) );
  NAND2_X1 U11435 ( .A1(n11365), .A2(n11366), .ZN(n11459) );
  NAND2_X1 U11436 ( .A1(n11463), .A2(n11464), .ZN(n11366) );
  NAND2_X1 U11437 ( .A1(n11363), .A2(n11465), .ZN(n11464) );
  OR2_X1 U11438 ( .A1(n11361), .A2(n11362), .ZN(n11465) );
  NOR2_X1 U11439 ( .A1(n8055), .A2(n7837), .ZN(n11363) );
  NAND2_X1 U11440 ( .A1(n11361), .A2(n11362), .ZN(n11463) );
  NAND2_X1 U11441 ( .A1(n11466), .A2(n11467), .ZN(n11362) );
  NAND2_X1 U11442 ( .A1(n11359), .A2(n11468), .ZN(n11467) );
  OR2_X1 U11443 ( .A1(n11357), .A2(n11358), .ZN(n11468) );
  NOR2_X1 U11444 ( .A1(n8055), .A2(n7817), .ZN(n11359) );
  NAND2_X1 U11445 ( .A1(n11357), .A2(n11358), .ZN(n11466) );
  NAND2_X1 U11446 ( .A1(n11469), .A2(n11470), .ZN(n11358) );
  NAND2_X1 U11447 ( .A1(n11355), .A2(n11471), .ZN(n11470) );
  NAND2_X1 U11448 ( .A1(n11354), .A2(n11353), .ZN(n11471) );
  NOR2_X1 U11449 ( .A1(n8055), .A2(n7806), .ZN(n11355) );
  OR2_X1 U11450 ( .A1(n11353), .A2(n11354), .ZN(n11469) );
  AND2_X1 U11451 ( .A1(n11472), .A2(n11473), .ZN(n11354) );
  NAND2_X1 U11452 ( .A1(n11474), .A2(b_18_), .ZN(n11473) );
  NOR2_X1 U11453 ( .A1(n11475), .A2(n7786), .ZN(n11474) );
  NOR2_X1 U11454 ( .A1(n11350), .A2(n11349), .ZN(n11475) );
  NAND2_X1 U11455 ( .A1(n11349), .A2(n11350), .ZN(n11472) );
  NAND2_X1 U11456 ( .A1(n11476), .A2(n11477), .ZN(n11350) );
  NAND2_X1 U11457 ( .A1(n11478), .A2(b_18_), .ZN(n11477) );
  NOR2_X1 U11458 ( .A1(n11479), .A2(n7775), .ZN(n11478) );
  NOR2_X1 U11459 ( .A1(n11344), .A2(n11346), .ZN(n11479) );
  NAND2_X1 U11460 ( .A1(n11344), .A2(n11346), .ZN(n11476) );
  NAND2_X1 U11461 ( .A1(n11480), .A2(n11481), .ZN(n11346) );
  NAND2_X1 U11462 ( .A1(n11343), .A2(n11482), .ZN(n11481) );
  OR2_X1 U11463 ( .A1(n11341), .A2(n11342), .ZN(n11482) );
  NOR2_X1 U11464 ( .A1(n8055), .A2(n7754), .ZN(n11343) );
  NAND2_X1 U11465 ( .A1(n11341), .A2(n11342), .ZN(n11480) );
  NAND2_X1 U11466 ( .A1(n11483), .A2(n11484), .ZN(n11342) );
  NAND2_X1 U11467 ( .A1(n11485), .A2(b_18_), .ZN(n11484) );
  NOR2_X1 U11468 ( .A1(n11486), .A2(n7743), .ZN(n11485) );
  NOR2_X1 U11469 ( .A1(n11336), .A2(n11338), .ZN(n11486) );
  NAND2_X1 U11470 ( .A1(n11336), .A2(n11338), .ZN(n11483) );
  NAND2_X1 U11471 ( .A1(n11487), .A2(n11488), .ZN(n11338) );
  NAND2_X1 U11472 ( .A1(n11335), .A2(n11489), .ZN(n11488) );
  OR2_X1 U11473 ( .A1(n11333), .A2(n11334), .ZN(n11489) );
  NOR2_X1 U11474 ( .A1(n8055), .A2(n7723), .ZN(n11335) );
  NAND2_X1 U11475 ( .A1(n11333), .A2(n11334), .ZN(n11487) );
  NAND2_X1 U11476 ( .A1(n11490), .A2(n11491), .ZN(n11334) );
  NAND2_X1 U11477 ( .A1(n11329), .A2(n11492), .ZN(n11491) );
  OR2_X1 U11478 ( .A1(n11330), .A2(n11331), .ZN(n11492) );
  XOR2_X1 U11479 ( .A(n11493), .B(n11494), .Z(n11329) );
  XOR2_X1 U11480 ( .A(n11495), .B(n11496), .Z(n11493) );
  NAND2_X1 U11481 ( .A1(n11331), .A2(n11330), .ZN(n11490) );
  NAND2_X1 U11482 ( .A1(n11497), .A2(n11498), .ZN(n11330) );
  NAND2_X1 U11483 ( .A1(n11327), .A2(n11499), .ZN(n11498) );
  OR2_X1 U11484 ( .A1(n11325), .A2(n11326), .ZN(n11499) );
  NOR2_X1 U11485 ( .A1(n8055), .A2(n7687), .ZN(n11327) );
  NAND2_X1 U11486 ( .A1(n11325), .A2(n11326), .ZN(n11497) );
  NAND2_X1 U11487 ( .A1(n11500), .A2(n11501), .ZN(n11326) );
  NAND2_X1 U11488 ( .A1(n11502), .A2(b_18_), .ZN(n11501) );
  NOR2_X1 U11489 ( .A1(n11503), .A2(n7676), .ZN(n11502) );
  NOR2_X1 U11490 ( .A1(n11321), .A2(n11322), .ZN(n11503) );
  NAND2_X1 U11491 ( .A1(n11321), .A2(n11322), .ZN(n11500) );
  NAND2_X1 U11492 ( .A1(n11504), .A2(n11505), .ZN(n11322) );
  NAND2_X1 U11493 ( .A1(n11318), .A2(n11506), .ZN(n11505) );
  OR2_X1 U11494 ( .A1(n11317), .A2(n11319), .ZN(n11506) );
  NOR2_X1 U11495 ( .A1(n8055), .A2(n7656), .ZN(n11318) );
  NAND2_X1 U11496 ( .A1(n11317), .A2(n11319), .ZN(n11504) );
  NAND2_X1 U11497 ( .A1(n11507), .A2(n11508), .ZN(n11319) );
  NAND2_X1 U11498 ( .A1(n11509), .A2(b_18_), .ZN(n11508) );
  NOR2_X1 U11499 ( .A1(n11510), .A2(n7645), .ZN(n11509) );
  NOR2_X1 U11500 ( .A1(n11314), .A2(n11312), .ZN(n11510) );
  NAND2_X1 U11501 ( .A1(n11312), .A2(n11314), .ZN(n11507) );
  NAND2_X1 U11502 ( .A1(n11511), .A2(n11512), .ZN(n11314) );
  NAND2_X1 U11503 ( .A1(n11311), .A2(n11513), .ZN(n11512) );
  NAND2_X1 U11504 ( .A1(n11310), .A2(n11309), .ZN(n11513) );
  NOR2_X1 U11505 ( .A1(n8055), .A2(n7624), .ZN(n11311) );
  OR2_X1 U11506 ( .A1(n11309), .A2(n11310), .ZN(n11511) );
  AND2_X1 U11507 ( .A1(n11306), .A2(n11514), .ZN(n11310) );
  NAND2_X1 U11508 ( .A1(n11305), .A2(n11307), .ZN(n11514) );
  NAND2_X1 U11509 ( .A1(n11515), .A2(n11516), .ZN(n11307) );
  NAND2_X1 U11510 ( .A1(b_18_), .A2(a_24_), .ZN(n11516) );
  INV_X1 U11511 ( .A(n11517), .ZN(n11515) );
  XNOR2_X1 U11512 ( .A(n11518), .B(n11519), .ZN(n11305) );
  XNOR2_X1 U11513 ( .A(n11520), .B(n11521), .ZN(n11518) );
  NAND2_X1 U11514 ( .A1(a_24_), .A2(n11517), .ZN(n11306) );
  NAND2_X1 U11515 ( .A1(n11522), .A2(n11523), .ZN(n11517) );
  NAND2_X1 U11516 ( .A1(n11524), .A2(b_18_), .ZN(n11523) );
  NOR2_X1 U11517 ( .A1(n11525), .A2(n7593), .ZN(n11524) );
  NOR2_X1 U11518 ( .A1(n11300), .A2(n11302), .ZN(n11525) );
  NAND2_X1 U11519 ( .A1(n11300), .A2(n11302), .ZN(n11522) );
  NAND2_X1 U11520 ( .A1(n11526), .A2(n11527), .ZN(n11302) );
  NAND2_X1 U11521 ( .A1(n11528), .A2(b_18_), .ZN(n11527) );
  NOR2_X1 U11522 ( .A1(n11529), .A2(n8052), .ZN(n11528) );
  NOR2_X1 U11523 ( .A1(n11299), .A2(n11297), .ZN(n11529) );
  NAND2_X1 U11524 ( .A1(n11297), .A2(n11299), .ZN(n11526) );
  NAND2_X1 U11525 ( .A1(n11530), .A2(n11531), .ZN(n11299) );
  NAND2_X1 U11526 ( .A1(n11295), .A2(n11532), .ZN(n11531) );
  NAND2_X1 U11527 ( .A1(n11294), .A2(n11293), .ZN(n11532) );
  NOR2_X1 U11528 ( .A1(n8055), .A2(n7563), .ZN(n11295) );
  INV_X1 U11529 ( .A(b_18_), .ZN(n8055) );
  OR2_X1 U11530 ( .A1(n11293), .A2(n11294), .ZN(n11530) );
  AND2_X1 U11531 ( .A1(n11290), .A2(n11533), .ZN(n11294) );
  NAND2_X1 U11532 ( .A1(n11289), .A2(n11291), .ZN(n11533) );
  NAND2_X1 U11533 ( .A1(n11534), .A2(n11535), .ZN(n11291) );
  NAND2_X1 U11534 ( .A1(b_18_), .A2(a_28_), .ZN(n11535) );
  INV_X1 U11535 ( .A(n11536), .ZN(n11534) );
  XOR2_X1 U11536 ( .A(n11537), .B(n11538), .Z(n11289) );
  NOR2_X1 U11537 ( .A1(n7529), .A2(n7724), .ZN(n11538) );
  XOR2_X1 U11538 ( .A(n11539), .B(n11540), .Z(n11537) );
  NAND2_X1 U11539 ( .A1(a_28_), .A2(n11536), .ZN(n11290) );
  NAND2_X1 U11540 ( .A1(n11541), .A2(n11542), .ZN(n11536) );
  NAND2_X1 U11541 ( .A1(n11543), .A2(b_18_), .ZN(n11542) );
  NOR2_X1 U11542 ( .A1(n11544), .A2(n7529), .ZN(n11543) );
  NOR2_X1 U11543 ( .A1(n11276), .A2(n11277), .ZN(n11544) );
  NAND2_X1 U11544 ( .A1(n11276), .A2(n11277), .ZN(n11541) );
  NAND2_X1 U11545 ( .A1(n11545), .A2(n11546), .ZN(n11277) );
  NAND2_X1 U11546 ( .A1(n11547), .A2(b_16_), .ZN(n11546) );
  NOR2_X1 U11547 ( .A1(n11548), .A2(n8048), .ZN(n11547) );
  NOR2_X1 U11548 ( .A1(n8676), .A2(n7724), .ZN(n11548) );
  NAND2_X1 U11549 ( .A1(n11549), .A2(b_17_), .ZN(n11545) );
  NOR2_X1 U11550 ( .A1(n11550), .A2(n7515), .ZN(n11549) );
  NOR2_X1 U11551 ( .A1(n8679), .A2(n11551), .ZN(n11550) );
  AND2_X1 U11552 ( .A1(n11552), .A2(b_18_), .ZN(n11276) );
  XOR2_X1 U11553 ( .A(n11553), .B(n11554), .Z(n11293) );
  NAND2_X1 U11554 ( .A1(n11555), .A2(n11556), .ZN(n11553) );
  XNOR2_X1 U11555 ( .A(n11557), .B(n11558), .ZN(n11297) );
  XNOR2_X1 U11556 ( .A(n11559), .B(n11560), .ZN(n11557) );
  XOR2_X1 U11557 ( .A(n11561), .B(n11562), .Z(n11300) );
  XNOR2_X1 U11558 ( .A(n11563), .B(n11564), .ZN(n11561) );
  NAND2_X1 U11559 ( .A1(b_17_), .A2(a_26_), .ZN(n11563) );
  XOR2_X1 U11560 ( .A(n11565), .B(n11566), .Z(n11309) );
  XOR2_X1 U11561 ( .A(n11567), .B(n11568), .Z(n11566) );
  NAND2_X1 U11562 ( .A1(b_17_), .A2(a_24_), .ZN(n11568) );
  XNOR2_X1 U11563 ( .A(n11569), .B(n11570), .ZN(n11312) );
  XNOR2_X1 U11564 ( .A(n11571), .B(n11572), .ZN(n11569) );
  XOR2_X1 U11565 ( .A(n11573), .B(n11574), .Z(n11317) );
  XOR2_X1 U11566 ( .A(n11575), .B(n11576), .Z(n11573) );
  NOR2_X1 U11567 ( .A1(n7645), .A2(n7724), .ZN(n11576) );
  XOR2_X1 U11568 ( .A(n11577), .B(n11578), .Z(n11321) );
  XOR2_X1 U11569 ( .A(n11579), .B(n11580), .Z(n11577) );
  XOR2_X1 U11570 ( .A(n11581), .B(n11582), .Z(n11325) );
  XOR2_X1 U11571 ( .A(n11583), .B(n11584), .Z(n11581) );
  NOR2_X1 U11572 ( .A1(n7676), .A2(n7724), .ZN(n11584) );
  INV_X1 U11573 ( .A(n7701), .ZN(n11331) );
  NAND2_X1 U11574 ( .A1(b_18_), .A2(a_18_), .ZN(n7701) );
  XOR2_X1 U11575 ( .A(n11585), .B(n11586), .Z(n11333) );
  XOR2_X1 U11576 ( .A(n11587), .B(n11588), .Z(n11585) );
  NOR2_X1 U11577 ( .A1(n7707), .A2(n7724), .ZN(n11588) );
  XOR2_X1 U11578 ( .A(n11589), .B(n11590), .Z(n11336) );
  XOR2_X1 U11579 ( .A(n11591), .B(n7718), .Z(n11589) );
  XNOR2_X1 U11580 ( .A(n11592), .B(n11593), .ZN(n11341) );
  XOR2_X1 U11581 ( .A(n11594), .B(n11595), .Z(n11593) );
  NAND2_X1 U11582 ( .A1(b_17_), .A2(a_16_), .ZN(n11595) );
  XOR2_X1 U11583 ( .A(n11596), .B(n11597), .Z(n11344) );
  XOR2_X1 U11584 ( .A(n11598), .B(n11599), .Z(n11596) );
  XNOR2_X1 U11585 ( .A(n11600), .B(n11601), .ZN(n11349) );
  XNOR2_X1 U11586 ( .A(n11602), .B(n11603), .ZN(n11600) );
  XOR2_X1 U11587 ( .A(n11604), .B(n11605), .Z(n11353) );
  XOR2_X1 U11588 ( .A(n11606), .B(n11607), .Z(n11605) );
  NAND2_X1 U11589 ( .A1(b_17_), .A2(a_13_), .ZN(n11607) );
  XNOR2_X1 U11590 ( .A(n11608), .B(n11609), .ZN(n11357) );
  NAND2_X1 U11591 ( .A1(n11610), .A2(n11611), .ZN(n11608) );
  XOR2_X1 U11592 ( .A(n11612), .B(n11613), .Z(n11361) );
  XOR2_X1 U11593 ( .A(n11614), .B(n11615), .Z(n11612) );
  NOR2_X1 U11594 ( .A1(n7817), .A2(n7724), .ZN(n11615) );
  XOR2_X1 U11595 ( .A(n11616), .B(n11617), .Z(n11365) );
  XOR2_X1 U11596 ( .A(n11618), .B(n11619), .Z(n11616) );
  NOR2_X1 U11597 ( .A1(n7837), .A2(n7724), .ZN(n11619) );
  XNOR2_X1 U11598 ( .A(n11620), .B(n11621), .ZN(n11377) );
  XOR2_X1 U11599 ( .A(n11622), .B(n11623), .Z(n11621) );
  NAND2_X1 U11600 ( .A1(b_17_), .A2(a_7_), .ZN(n11623) );
  XNOR2_X1 U11601 ( .A(n11624), .B(n11625), .ZN(n11381) );
  XOR2_X1 U11602 ( .A(n11626), .B(n11627), .Z(n11625) );
  NAND2_X1 U11603 ( .A1(b_17_), .A2(a_6_), .ZN(n11627) );
  XOR2_X1 U11604 ( .A(n11628), .B(n11629), .Z(n11392) );
  XOR2_X1 U11605 ( .A(n11630), .B(n11631), .Z(n11628) );
  NOR2_X1 U11606 ( .A1(n7965), .A2(n7724), .ZN(n11631) );
  XOR2_X1 U11607 ( .A(n11632), .B(n11633), .Z(n11159) );
  XOR2_X1 U11608 ( .A(n11634), .B(n11635), .Z(n11632) );
  NOR2_X1 U11609 ( .A1(n7973), .A2(n7724), .ZN(n11635) );
  NAND2_X1 U11610 ( .A1(n11636), .A2(n11637), .ZN(n8156) );
  XOR2_X1 U11611 ( .A(n8240), .B(n11638), .Z(n11637) );
  AND2_X1 U11612 ( .A1(n8238), .A2(n8237), .ZN(n11636) );
  INV_X1 U11613 ( .A(n11398), .ZN(n8237) );
  XOR2_X1 U11614 ( .A(n11639), .B(n11640), .Z(n11398) );
  XNOR2_X1 U11615 ( .A(n11641), .B(n11642), .ZN(n11639) );
  NAND2_X1 U11616 ( .A1(n11643), .A2(n11644), .ZN(n8238) );
  NAND2_X1 U11617 ( .A1(n11645), .A2(b_17_), .ZN(n11644) );
  NOR2_X1 U11618 ( .A1(n11646), .A2(n8307), .ZN(n11645) );
  NOR2_X1 U11619 ( .A1(n11401), .A2(n11403), .ZN(n11646) );
  NAND2_X1 U11620 ( .A1(n11401), .A2(n11403), .ZN(n11643) );
  NAND2_X1 U11621 ( .A1(n11647), .A2(n11648), .ZN(n11403) );
  NAND2_X1 U11622 ( .A1(n11649), .A2(b_17_), .ZN(n11648) );
  NOR2_X1 U11623 ( .A1(n11650), .A2(n7973), .ZN(n11649) );
  NOR2_X1 U11624 ( .A1(n11633), .A2(n11634), .ZN(n11650) );
  NAND2_X1 U11625 ( .A1(n11633), .A2(n11634), .ZN(n11647) );
  NAND2_X1 U11626 ( .A1(n11651), .A2(n11652), .ZN(n11634) );
  NAND2_X1 U11627 ( .A1(n11653), .A2(b_17_), .ZN(n11652) );
  NOR2_X1 U11628 ( .A1(n11654), .A2(n7965), .ZN(n11653) );
  NOR2_X1 U11629 ( .A1(n11629), .A2(n11630), .ZN(n11654) );
  NAND2_X1 U11630 ( .A1(n11629), .A2(n11630), .ZN(n11651) );
  NAND2_X1 U11631 ( .A1(n11655), .A2(n11656), .ZN(n11630) );
  NAND2_X1 U11632 ( .A1(n11657), .A2(b_17_), .ZN(n11656) );
  NOR2_X1 U11633 ( .A1(n11658), .A2(n7945), .ZN(n11657) );
  NOR2_X1 U11634 ( .A1(n11417), .A2(n11418), .ZN(n11658) );
  NAND2_X1 U11635 ( .A1(n11417), .A2(n11418), .ZN(n11655) );
  NAND2_X1 U11636 ( .A1(n11659), .A2(n11660), .ZN(n11418) );
  NAND2_X1 U11637 ( .A1(n11661), .A2(b_17_), .ZN(n11660) );
  NOR2_X1 U11638 ( .A1(n11662), .A2(n7934), .ZN(n11661) );
  NOR2_X1 U11639 ( .A1(n11425), .A2(n11426), .ZN(n11662) );
  NAND2_X1 U11640 ( .A1(n11425), .A2(n11426), .ZN(n11659) );
  NAND2_X1 U11641 ( .A1(n11663), .A2(n11664), .ZN(n11426) );
  NAND2_X1 U11642 ( .A1(n11665), .A2(b_17_), .ZN(n11664) );
  NOR2_X1 U11643 ( .A1(n11666), .A2(n7914), .ZN(n11665) );
  NOR2_X1 U11644 ( .A1(n11433), .A2(n11434), .ZN(n11666) );
  NAND2_X1 U11645 ( .A1(n11433), .A2(n11434), .ZN(n11663) );
  NAND2_X1 U11646 ( .A1(n11667), .A2(n11668), .ZN(n11434) );
  NAND2_X1 U11647 ( .A1(n11669), .A2(b_17_), .ZN(n11668) );
  NOR2_X1 U11648 ( .A1(n11670), .A2(n8061), .ZN(n11669) );
  NOR2_X1 U11649 ( .A1(n11624), .A2(n11626), .ZN(n11670) );
  NAND2_X1 U11650 ( .A1(n11624), .A2(n11626), .ZN(n11667) );
  NAND2_X1 U11651 ( .A1(n11671), .A2(n11672), .ZN(n11626) );
  NAND2_X1 U11652 ( .A1(n11673), .A2(b_17_), .ZN(n11672) );
  NOR2_X1 U11653 ( .A1(n11674), .A2(n7884), .ZN(n11673) );
  NOR2_X1 U11654 ( .A1(n11620), .A2(n11622), .ZN(n11674) );
  NAND2_X1 U11655 ( .A1(n11620), .A2(n11622), .ZN(n11671) );
  NAND2_X1 U11656 ( .A1(n11675), .A2(n11676), .ZN(n11622) );
  NAND2_X1 U11657 ( .A1(n11677), .A2(b_17_), .ZN(n11676) );
  NOR2_X1 U11658 ( .A1(n11678), .A2(n8059), .ZN(n11677) );
  NOR2_X1 U11659 ( .A1(n11447), .A2(n11449), .ZN(n11678) );
  NAND2_X1 U11660 ( .A1(n11447), .A2(n11449), .ZN(n11675) );
  NAND2_X1 U11661 ( .A1(n11679), .A2(n11680), .ZN(n11449) );
  NAND2_X1 U11662 ( .A1(n11681), .A2(b_17_), .ZN(n11680) );
  NOR2_X1 U11663 ( .A1(n11682), .A2(n7848), .ZN(n11681) );
  NOR2_X1 U11664 ( .A1(n11456), .A2(n11457), .ZN(n11682) );
  NAND2_X1 U11665 ( .A1(n11456), .A2(n11457), .ZN(n11679) );
  NAND2_X1 U11666 ( .A1(n11683), .A2(n11684), .ZN(n11457) );
  NAND2_X1 U11667 ( .A1(n11685), .A2(b_17_), .ZN(n11684) );
  NOR2_X1 U11668 ( .A1(n11686), .A2(n7837), .ZN(n11685) );
  NOR2_X1 U11669 ( .A1(n11617), .A2(n11618), .ZN(n11686) );
  NAND2_X1 U11670 ( .A1(n11617), .A2(n11618), .ZN(n11683) );
  NAND2_X1 U11671 ( .A1(n11687), .A2(n11688), .ZN(n11618) );
  NAND2_X1 U11672 ( .A1(n11689), .A2(b_17_), .ZN(n11688) );
  NOR2_X1 U11673 ( .A1(n11690), .A2(n7817), .ZN(n11689) );
  NOR2_X1 U11674 ( .A1(n11613), .A2(n11614), .ZN(n11690) );
  NAND2_X1 U11675 ( .A1(n11613), .A2(n11614), .ZN(n11687) );
  NAND2_X1 U11676 ( .A1(n11610), .A2(n11691), .ZN(n11614) );
  NAND2_X1 U11677 ( .A1(n11609), .A2(n11611), .ZN(n11691) );
  NAND2_X1 U11678 ( .A1(n11692), .A2(n11693), .ZN(n11611) );
  NAND2_X1 U11679 ( .A1(b_17_), .A2(a_12_), .ZN(n11693) );
  INV_X1 U11680 ( .A(n11694), .ZN(n11692) );
  XNOR2_X1 U11681 ( .A(n11695), .B(n11696), .ZN(n11609) );
  XNOR2_X1 U11682 ( .A(n11697), .B(n11698), .ZN(n11695) );
  NAND2_X1 U11683 ( .A1(a_12_), .A2(n11694), .ZN(n11610) );
  NAND2_X1 U11684 ( .A1(n11699), .A2(n11700), .ZN(n11694) );
  NAND2_X1 U11685 ( .A1(n11701), .A2(b_17_), .ZN(n11700) );
  NOR2_X1 U11686 ( .A1(n11702), .A2(n7786), .ZN(n11701) );
  NOR2_X1 U11687 ( .A1(n11604), .A2(n11606), .ZN(n11702) );
  NAND2_X1 U11688 ( .A1(n11604), .A2(n11606), .ZN(n11699) );
  NAND2_X1 U11689 ( .A1(n11703), .A2(n11704), .ZN(n11606) );
  NAND2_X1 U11690 ( .A1(n11603), .A2(n11705), .ZN(n11704) );
  NAND2_X1 U11691 ( .A1(n11602), .A2(n11601), .ZN(n11705) );
  NOR2_X1 U11692 ( .A1(n7724), .A2(n7775), .ZN(n11603) );
  OR2_X1 U11693 ( .A1(n11601), .A2(n11602), .ZN(n11703) );
  AND2_X1 U11694 ( .A1(n11706), .A2(n11707), .ZN(n11602) );
  NAND2_X1 U11695 ( .A1(n11599), .A2(n11708), .ZN(n11707) );
  OR2_X1 U11696 ( .A1(n11598), .A2(n11597), .ZN(n11708) );
  NOR2_X1 U11697 ( .A1(n7724), .A2(n7754), .ZN(n11599) );
  NAND2_X1 U11698 ( .A1(n11597), .A2(n11598), .ZN(n11706) );
  NAND2_X1 U11699 ( .A1(n11709), .A2(n11710), .ZN(n11598) );
  NAND2_X1 U11700 ( .A1(n11711), .A2(b_17_), .ZN(n11710) );
  NOR2_X1 U11701 ( .A1(n11712), .A2(n7743), .ZN(n11711) );
  NOR2_X1 U11702 ( .A1(n11592), .A2(n11594), .ZN(n11712) );
  NAND2_X1 U11703 ( .A1(n11592), .A2(n11594), .ZN(n11709) );
  NAND2_X1 U11704 ( .A1(n11713), .A2(n11714), .ZN(n11594) );
  NAND2_X1 U11705 ( .A1(n7718), .A2(n11715), .ZN(n11714) );
  OR2_X1 U11706 ( .A1(n11591), .A2(n11590), .ZN(n11715) );
  INV_X1 U11707 ( .A(n8019), .ZN(n7718) );
  NAND2_X1 U11708 ( .A1(b_17_), .A2(a_17_), .ZN(n8019) );
  NAND2_X1 U11709 ( .A1(n11590), .A2(n11591), .ZN(n11713) );
  NAND2_X1 U11710 ( .A1(n11716), .A2(n11717), .ZN(n11591) );
  NAND2_X1 U11711 ( .A1(n11718), .A2(b_17_), .ZN(n11717) );
  NOR2_X1 U11712 ( .A1(n11719), .A2(n7707), .ZN(n11718) );
  NOR2_X1 U11713 ( .A1(n11586), .A2(n11587), .ZN(n11719) );
  NAND2_X1 U11714 ( .A1(n11586), .A2(n11587), .ZN(n11716) );
  NAND2_X1 U11715 ( .A1(n11720), .A2(n11721), .ZN(n11587) );
  NAND2_X1 U11716 ( .A1(n11496), .A2(n11722), .ZN(n11721) );
  OR2_X1 U11717 ( .A1(n11495), .A2(n11494), .ZN(n11722) );
  NOR2_X1 U11718 ( .A1(n7724), .A2(n7687), .ZN(n11496) );
  NAND2_X1 U11719 ( .A1(n11494), .A2(n11495), .ZN(n11720) );
  NAND2_X1 U11720 ( .A1(n11723), .A2(n11724), .ZN(n11495) );
  NAND2_X1 U11721 ( .A1(n11725), .A2(b_17_), .ZN(n11724) );
  NOR2_X1 U11722 ( .A1(n11726), .A2(n7676), .ZN(n11725) );
  NOR2_X1 U11723 ( .A1(n11582), .A2(n11583), .ZN(n11726) );
  NAND2_X1 U11724 ( .A1(n11582), .A2(n11583), .ZN(n11723) );
  NAND2_X1 U11725 ( .A1(n11727), .A2(n11728), .ZN(n11583) );
  NAND2_X1 U11726 ( .A1(n11580), .A2(n11729), .ZN(n11728) );
  OR2_X1 U11727 ( .A1(n11579), .A2(n11578), .ZN(n11729) );
  NOR2_X1 U11728 ( .A1(n7724), .A2(n7656), .ZN(n11580) );
  NAND2_X1 U11729 ( .A1(n11578), .A2(n11579), .ZN(n11727) );
  NAND2_X1 U11730 ( .A1(n11730), .A2(n11731), .ZN(n11579) );
  NAND2_X1 U11731 ( .A1(n11732), .A2(b_17_), .ZN(n11731) );
  NOR2_X1 U11732 ( .A1(n11733), .A2(n7645), .ZN(n11732) );
  NOR2_X1 U11733 ( .A1(n11574), .A2(n11575), .ZN(n11733) );
  NAND2_X1 U11734 ( .A1(n11574), .A2(n11575), .ZN(n11730) );
  NAND2_X1 U11735 ( .A1(n11734), .A2(n11735), .ZN(n11575) );
  NAND2_X1 U11736 ( .A1(n11572), .A2(n11736), .ZN(n11735) );
  NAND2_X1 U11737 ( .A1(n11571), .A2(n11570), .ZN(n11736) );
  NOR2_X1 U11738 ( .A1(n7724), .A2(n7624), .ZN(n11572) );
  OR2_X1 U11739 ( .A1(n11570), .A2(n11571), .ZN(n11734) );
  AND2_X1 U11740 ( .A1(n11737), .A2(n11738), .ZN(n11571) );
  NAND2_X1 U11741 ( .A1(n11739), .A2(b_17_), .ZN(n11738) );
  NOR2_X1 U11742 ( .A1(n11740), .A2(n7613), .ZN(n11739) );
  NOR2_X1 U11743 ( .A1(n11565), .A2(n11567), .ZN(n11740) );
  NAND2_X1 U11744 ( .A1(n11565), .A2(n11567), .ZN(n11737) );
  NAND2_X1 U11745 ( .A1(n11741), .A2(n11742), .ZN(n11567) );
  NAND2_X1 U11746 ( .A1(n11521), .A2(n11743), .ZN(n11742) );
  NAND2_X1 U11747 ( .A1(n11520), .A2(n11519), .ZN(n11743) );
  NOR2_X1 U11748 ( .A1(n7724), .A2(n7593), .ZN(n11521) );
  OR2_X1 U11749 ( .A1(n11519), .A2(n11520), .ZN(n11741) );
  AND2_X1 U11750 ( .A1(n11744), .A2(n11745), .ZN(n11520) );
  NAND2_X1 U11751 ( .A1(n11746), .A2(b_17_), .ZN(n11745) );
  NOR2_X1 U11752 ( .A1(n11747), .A2(n8052), .ZN(n11746) );
  NOR2_X1 U11753 ( .A1(n11562), .A2(n11564), .ZN(n11747) );
  NAND2_X1 U11754 ( .A1(n11562), .A2(n11564), .ZN(n11744) );
  NAND2_X1 U11755 ( .A1(n11748), .A2(n11749), .ZN(n11564) );
  NAND2_X1 U11756 ( .A1(n11560), .A2(n11750), .ZN(n11749) );
  NAND2_X1 U11757 ( .A1(n11559), .A2(n11558), .ZN(n11750) );
  NOR2_X1 U11758 ( .A1(n7724), .A2(n7563), .ZN(n11560) );
  OR2_X1 U11759 ( .A1(n11558), .A2(n11559), .ZN(n11748) );
  AND2_X1 U11760 ( .A1(n11555), .A2(n11751), .ZN(n11559) );
  NAND2_X1 U11761 ( .A1(n11554), .A2(n11556), .ZN(n11751) );
  NAND2_X1 U11762 ( .A1(n11752), .A2(n11753), .ZN(n11556) );
  NAND2_X1 U11763 ( .A1(b_17_), .A2(a_28_), .ZN(n11753) );
  INV_X1 U11764 ( .A(n11754), .ZN(n11752) );
  XOR2_X1 U11765 ( .A(n11755), .B(n11756), .Z(n11554) );
  NOR2_X1 U11766 ( .A1(n7529), .A2(n11551), .ZN(n11756) );
  XOR2_X1 U11767 ( .A(n11757), .B(n11758), .Z(n11755) );
  NAND2_X1 U11768 ( .A1(a_28_), .A2(n11754), .ZN(n11555) );
  NAND2_X1 U11769 ( .A1(n11759), .A2(n11760), .ZN(n11754) );
  NAND2_X1 U11770 ( .A1(n11761), .A2(b_17_), .ZN(n11760) );
  NOR2_X1 U11771 ( .A1(n11762), .A2(n7529), .ZN(n11761) );
  NOR2_X1 U11772 ( .A1(n11539), .A2(n11540), .ZN(n11762) );
  NAND2_X1 U11773 ( .A1(n11539), .A2(n11540), .ZN(n11759) );
  NAND2_X1 U11774 ( .A1(n11763), .A2(n11764), .ZN(n11540) );
  NAND2_X1 U11775 ( .A1(n11765), .A2(b_15_), .ZN(n11764) );
  NOR2_X1 U11776 ( .A1(n11766), .A2(n8048), .ZN(n11765) );
  NOR2_X1 U11777 ( .A1(n8676), .A2(n11551), .ZN(n11766) );
  NAND2_X1 U11778 ( .A1(n11767), .A2(b_16_), .ZN(n11763) );
  NOR2_X1 U11779 ( .A1(n11768), .A2(n7515), .ZN(n11767) );
  NOR2_X1 U11780 ( .A1(n8679), .A2(n7755), .ZN(n11768) );
  AND2_X1 U11781 ( .A1(n11552), .A2(b_16_), .ZN(n11539) );
  NOR2_X1 U11782 ( .A1(n8451), .A2(n7724), .ZN(n11552) );
  INV_X1 U11783 ( .A(b_17_), .ZN(n7724) );
  XOR2_X1 U11784 ( .A(n11769), .B(n11770), .Z(n11558) );
  NAND2_X1 U11785 ( .A1(n11771), .A2(n11772), .ZN(n11769) );
  XNOR2_X1 U11786 ( .A(n11773), .B(n11774), .ZN(n11562) );
  XNOR2_X1 U11787 ( .A(n11775), .B(n11776), .ZN(n11773) );
  XNOR2_X1 U11788 ( .A(n11777), .B(n11778), .ZN(n11519) );
  XNOR2_X1 U11789 ( .A(n11779), .B(n11780), .ZN(n11777) );
  NAND2_X1 U11790 ( .A1(b_16_), .A2(a_26_), .ZN(n11779) );
  XNOR2_X1 U11791 ( .A(n11781), .B(n11782), .ZN(n11565) );
  XNOR2_X1 U11792 ( .A(n11783), .B(n11784), .ZN(n11782) );
  XOR2_X1 U11793 ( .A(n11785), .B(n11786), .Z(n11570) );
  XOR2_X1 U11794 ( .A(n11787), .B(n11788), .Z(n11786) );
  NAND2_X1 U11795 ( .A1(b_16_), .A2(a_24_), .ZN(n11788) );
  XOR2_X1 U11796 ( .A(n11789), .B(n11790), .Z(n11574) );
  XOR2_X1 U11797 ( .A(n11791), .B(n11792), .Z(n11789) );
  XOR2_X1 U11798 ( .A(n11793), .B(n11794), .Z(n11578) );
  XOR2_X1 U11799 ( .A(n11795), .B(n11796), .Z(n11793) );
  NOR2_X1 U11800 ( .A1(n7645), .A2(n11551), .ZN(n11796) );
  XOR2_X1 U11801 ( .A(n11797), .B(n11798), .Z(n11582) );
  XOR2_X1 U11802 ( .A(n11799), .B(n11800), .Z(n11797) );
  XNOR2_X1 U11803 ( .A(n11801), .B(n11802), .ZN(n11494) );
  XOR2_X1 U11804 ( .A(n11803), .B(n11804), .Z(n11802) );
  NAND2_X1 U11805 ( .A1(b_16_), .A2(a_20_), .ZN(n11804) );
  XOR2_X1 U11806 ( .A(n11805), .B(n11806), .Z(n11586) );
  XOR2_X1 U11807 ( .A(n11807), .B(n11808), .Z(n11805) );
  XNOR2_X1 U11808 ( .A(n11809), .B(n11810), .ZN(n11590) );
  XOR2_X1 U11809 ( .A(n11811), .B(n11812), .Z(n11810) );
  NAND2_X1 U11810 ( .A1(b_16_), .A2(a_18_), .ZN(n11812) );
  XOR2_X1 U11811 ( .A(n11813), .B(n11814), .Z(n11592) );
  XOR2_X1 U11812 ( .A(n11815), .B(n11816), .Z(n11813) );
  XNOR2_X1 U11813 ( .A(n11817), .B(n11818), .ZN(n11597) );
  XNOR2_X1 U11814 ( .A(n11819), .B(n7737), .ZN(n11818) );
  XNOR2_X1 U11815 ( .A(n11820), .B(n11821), .ZN(n11601) );
  XOR2_X1 U11816 ( .A(n11822), .B(n11823), .Z(n11820) );
  NOR2_X1 U11817 ( .A1(n7754), .A2(n11551), .ZN(n11823) );
  XNOR2_X1 U11818 ( .A(n11824), .B(n11825), .ZN(n11604) );
  XNOR2_X1 U11819 ( .A(n11826), .B(n11827), .ZN(n11824) );
  XNOR2_X1 U11820 ( .A(n11828), .B(n11829), .ZN(n11613) );
  XNOR2_X1 U11821 ( .A(n11830), .B(n11831), .ZN(n11829) );
  XNOR2_X1 U11822 ( .A(n11832), .B(n11833), .ZN(n11617) );
  XNOR2_X1 U11823 ( .A(n11834), .B(n11835), .ZN(n11832) );
  XNOR2_X1 U11824 ( .A(n11836), .B(n11837), .ZN(n11456) );
  XOR2_X1 U11825 ( .A(n11838), .B(n11839), .Z(n11837) );
  NAND2_X1 U11826 ( .A1(b_16_), .A2(a_10_), .ZN(n11839) );
  XNOR2_X1 U11827 ( .A(n11840), .B(n11841), .ZN(n11447) );
  NAND2_X1 U11828 ( .A1(n11842), .A2(n11843), .ZN(n11840) );
  XNOR2_X1 U11829 ( .A(n11844), .B(n11845), .ZN(n11620) );
  XNOR2_X1 U11830 ( .A(n11846), .B(n11847), .ZN(n11845) );
  XOR2_X1 U11831 ( .A(n11848), .B(n11849), .Z(n11624) );
  XOR2_X1 U11832 ( .A(n11850), .B(n11851), .Z(n11848) );
  XNOR2_X1 U11833 ( .A(n11852), .B(n11853), .ZN(n11433) );
  XNOR2_X1 U11834 ( .A(n11854), .B(n11855), .ZN(n11852) );
  XNOR2_X1 U11835 ( .A(n11856), .B(n11857), .ZN(n11425) );
  XOR2_X1 U11836 ( .A(n11858), .B(n11859), .Z(n11857) );
  NAND2_X1 U11837 ( .A1(b_16_), .A2(a_5_), .ZN(n11859) );
  XOR2_X1 U11838 ( .A(n11860), .B(n11861), .Z(n11417) );
  XOR2_X1 U11839 ( .A(n11862), .B(n11863), .Z(n11860) );
  XOR2_X1 U11840 ( .A(n11864), .B(n11865), .Z(n11629) );
  XOR2_X1 U11841 ( .A(n11866), .B(n11867), .Z(n11864) );
  XNOR2_X1 U11842 ( .A(n11868), .B(n11869), .ZN(n11633) );
  XNOR2_X1 U11843 ( .A(n11870), .B(n11871), .ZN(n11868) );
  XOR2_X1 U11844 ( .A(n11872), .B(n11873), .Z(n11401) );
  XOR2_X1 U11845 ( .A(n11874), .B(n11875), .Z(n11872) );
  NAND2_X1 U11846 ( .A1(n11876), .A2(n11877), .ZN(n8162) );
  NAND2_X1 U11847 ( .A1(n11878), .A2(n8239), .ZN(n11877) );
  INV_X1 U11848 ( .A(n8240), .ZN(n11878) );
  XOR2_X1 U11849 ( .A(n11879), .B(n11880), .Z(n11876) );
  NAND2_X1 U11850 ( .A1(n11881), .A2(n11882), .ZN(n8161) );
  XOR2_X1 U11851 ( .A(n11879), .B(n11883), .Z(n11882) );
  NOR2_X1 U11852 ( .A1(n11638), .A2(n8240), .ZN(n11881) );
  XNOR2_X1 U11853 ( .A(n11884), .B(n11885), .ZN(n8240) );
  XOR2_X1 U11854 ( .A(n11886), .B(n11887), .Z(n11884) );
  NOR2_X1 U11855 ( .A1(n8307), .A2(n7755), .ZN(n11887) );
  INV_X1 U11856 ( .A(n8239), .ZN(n11638) );
  NAND2_X1 U11857 ( .A1(n11888), .A2(n11889), .ZN(n8239) );
  NAND2_X1 U11858 ( .A1(n11642), .A2(n11890), .ZN(n11889) );
  NAND2_X1 U11859 ( .A1(n11641), .A2(n11640), .ZN(n11890) );
  NOR2_X1 U11860 ( .A1(n11551), .A2(n8307), .ZN(n11642) );
  OR2_X1 U11861 ( .A1(n11640), .A2(n11641), .ZN(n11888) );
  AND2_X1 U11862 ( .A1(n11891), .A2(n11892), .ZN(n11641) );
  NAND2_X1 U11863 ( .A1(n11874), .A2(n11893), .ZN(n11892) );
  OR2_X1 U11864 ( .A1(n11873), .A2(n11875), .ZN(n11893) );
  NOR2_X1 U11865 ( .A1(n11551), .A2(n7973), .ZN(n11874) );
  NAND2_X1 U11866 ( .A1(n11873), .A2(n11875), .ZN(n11891) );
  NAND2_X1 U11867 ( .A1(n11894), .A2(n11895), .ZN(n11875) );
  NAND2_X1 U11868 ( .A1(n11871), .A2(n11896), .ZN(n11895) );
  NAND2_X1 U11869 ( .A1(n11870), .A2(n11869), .ZN(n11896) );
  NOR2_X1 U11870 ( .A1(n11551), .A2(n7965), .ZN(n11871) );
  OR2_X1 U11871 ( .A1(n11869), .A2(n11870), .ZN(n11894) );
  AND2_X1 U11872 ( .A1(n11897), .A2(n11898), .ZN(n11870) );
  NAND2_X1 U11873 ( .A1(n11867), .A2(n11899), .ZN(n11898) );
  OR2_X1 U11874 ( .A1(n11865), .A2(n11866), .ZN(n11899) );
  NOR2_X1 U11875 ( .A1(n11551), .A2(n7945), .ZN(n11867) );
  NAND2_X1 U11876 ( .A1(n11865), .A2(n11866), .ZN(n11897) );
  NAND2_X1 U11877 ( .A1(n11900), .A2(n11901), .ZN(n11866) );
  NAND2_X1 U11878 ( .A1(n11863), .A2(n11902), .ZN(n11901) );
  OR2_X1 U11879 ( .A1(n11861), .A2(n11862), .ZN(n11902) );
  NOR2_X1 U11880 ( .A1(n11551), .A2(n7934), .ZN(n11863) );
  NAND2_X1 U11881 ( .A1(n11861), .A2(n11862), .ZN(n11900) );
  NAND2_X1 U11882 ( .A1(n11903), .A2(n11904), .ZN(n11862) );
  NAND2_X1 U11883 ( .A1(n11905), .A2(b_16_), .ZN(n11904) );
  NOR2_X1 U11884 ( .A1(n11906), .A2(n7914), .ZN(n11905) );
  NOR2_X1 U11885 ( .A1(n11856), .A2(n11858), .ZN(n11906) );
  NAND2_X1 U11886 ( .A1(n11856), .A2(n11858), .ZN(n11903) );
  NAND2_X1 U11887 ( .A1(n11907), .A2(n11908), .ZN(n11858) );
  NAND2_X1 U11888 ( .A1(n11855), .A2(n11909), .ZN(n11908) );
  NAND2_X1 U11889 ( .A1(n11854), .A2(n11853), .ZN(n11909) );
  NOR2_X1 U11890 ( .A1(n11551), .A2(n8061), .ZN(n11855) );
  OR2_X1 U11891 ( .A1(n11853), .A2(n11854), .ZN(n11907) );
  AND2_X1 U11892 ( .A1(n11910), .A2(n11911), .ZN(n11854) );
  NAND2_X1 U11893 ( .A1(n11851), .A2(n11912), .ZN(n11911) );
  OR2_X1 U11894 ( .A1(n11849), .A2(n11850), .ZN(n11912) );
  NOR2_X1 U11895 ( .A1(n11551), .A2(n7884), .ZN(n11851) );
  NAND2_X1 U11896 ( .A1(n11849), .A2(n11850), .ZN(n11910) );
  NAND2_X1 U11897 ( .A1(n11913), .A2(n11914), .ZN(n11850) );
  NAND2_X1 U11898 ( .A1(n11847), .A2(n11915), .ZN(n11914) );
  OR2_X1 U11899 ( .A1(n11844), .A2(n11846), .ZN(n11915) );
  NOR2_X1 U11900 ( .A1(n11551), .A2(n8059), .ZN(n11847) );
  NAND2_X1 U11901 ( .A1(n11844), .A2(n11846), .ZN(n11913) );
  NAND2_X1 U11902 ( .A1(n11842), .A2(n11916), .ZN(n11846) );
  NAND2_X1 U11903 ( .A1(n11841), .A2(n11843), .ZN(n11916) );
  NAND2_X1 U11904 ( .A1(n11917), .A2(n11918), .ZN(n11843) );
  NAND2_X1 U11905 ( .A1(b_16_), .A2(a_9_), .ZN(n11918) );
  INV_X1 U11906 ( .A(n11919), .ZN(n11917) );
  XNOR2_X1 U11907 ( .A(n11920), .B(n11921), .ZN(n11841) );
  XOR2_X1 U11908 ( .A(n11922), .B(n11923), .Z(n11921) );
  NAND2_X1 U11909 ( .A1(b_15_), .A2(a_10_), .ZN(n11923) );
  NAND2_X1 U11910 ( .A1(a_9_), .A2(n11919), .ZN(n11842) );
  NAND2_X1 U11911 ( .A1(n11924), .A2(n11925), .ZN(n11919) );
  NAND2_X1 U11912 ( .A1(n11926), .A2(b_16_), .ZN(n11925) );
  NOR2_X1 U11913 ( .A1(n11927), .A2(n7837), .ZN(n11926) );
  NOR2_X1 U11914 ( .A1(n11836), .A2(n11838), .ZN(n11927) );
  NAND2_X1 U11915 ( .A1(n11836), .A2(n11838), .ZN(n11924) );
  NAND2_X1 U11916 ( .A1(n11928), .A2(n11929), .ZN(n11838) );
  NAND2_X1 U11917 ( .A1(n11835), .A2(n11930), .ZN(n11929) );
  NAND2_X1 U11918 ( .A1(n11834), .A2(n11833), .ZN(n11930) );
  NOR2_X1 U11919 ( .A1(n11551), .A2(n7817), .ZN(n11835) );
  OR2_X1 U11920 ( .A1(n11833), .A2(n11834), .ZN(n11928) );
  AND2_X1 U11921 ( .A1(n11931), .A2(n11932), .ZN(n11834) );
  NAND2_X1 U11922 ( .A1(n11831), .A2(n11933), .ZN(n11932) );
  OR2_X1 U11923 ( .A1(n11828), .A2(n11830), .ZN(n11933) );
  NOR2_X1 U11924 ( .A1(n11551), .A2(n7806), .ZN(n11831) );
  NAND2_X1 U11925 ( .A1(n11828), .A2(n11830), .ZN(n11931) );
  NAND2_X1 U11926 ( .A1(n11934), .A2(n11935), .ZN(n11830) );
  NAND2_X1 U11927 ( .A1(n11698), .A2(n11936), .ZN(n11935) );
  NAND2_X1 U11928 ( .A1(n11697), .A2(n11696), .ZN(n11936) );
  NOR2_X1 U11929 ( .A1(n11551), .A2(n7786), .ZN(n11698) );
  OR2_X1 U11930 ( .A1(n11696), .A2(n11697), .ZN(n11934) );
  AND2_X1 U11931 ( .A1(n11937), .A2(n11938), .ZN(n11697) );
  NAND2_X1 U11932 ( .A1(n11827), .A2(n11939), .ZN(n11938) );
  NAND2_X1 U11933 ( .A1(n11826), .A2(n11825), .ZN(n11939) );
  NOR2_X1 U11934 ( .A1(n11551), .A2(n7775), .ZN(n11827) );
  OR2_X1 U11935 ( .A1(n11825), .A2(n11826), .ZN(n11937) );
  AND2_X1 U11936 ( .A1(n11940), .A2(n11941), .ZN(n11826) );
  NAND2_X1 U11937 ( .A1(n11942), .A2(b_16_), .ZN(n11941) );
  NOR2_X1 U11938 ( .A1(n11943), .A2(n7754), .ZN(n11942) );
  NOR2_X1 U11939 ( .A1(n11822), .A2(n11821), .ZN(n11943) );
  NAND2_X1 U11940 ( .A1(n11821), .A2(n11822), .ZN(n11940) );
  NAND2_X1 U11941 ( .A1(n11944), .A2(n11945), .ZN(n11822) );
  NAND2_X1 U11942 ( .A1(n11817), .A2(n11946), .ZN(n11945) );
  OR2_X1 U11943 ( .A1(n11819), .A2(n7737), .ZN(n11946) );
  XOR2_X1 U11944 ( .A(n11947), .B(n11948), .Z(n11817) );
  XOR2_X1 U11945 ( .A(n11949), .B(n11950), .Z(n11947) );
  NAND2_X1 U11946 ( .A1(n7737), .A2(n11819), .ZN(n11944) );
  NAND2_X1 U11947 ( .A1(n11951), .A2(n11952), .ZN(n11819) );
  NAND2_X1 U11948 ( .A1(n11816), .A2(n11953), .ZN(n11952) );
  OR2_X1 U11949 ( .A1(n11814), .A2(n11815), .ZN(n11953) );
  NOR2_X1 U11950 ( .A1(n11551), .A2(n7723), .ZN(n11816) );
  NAND2_X1 U11951 ( .A1(n11814), .A2(n11815), .ZN(n11951) );
  NAND2_X1 U11952 ( .A1(n11954), .A2(n11955), .ZN(n11815) );
  NAND2_X1 U11953 ( .A1(n11956), .A2(b_16_), .ZN(n11955) );
  NOR2_X1 U11954 ( .A1(n11957), .A2(n7707), .ZN(n11956) );
  NOR2_X1 U11955 ( .A1(n11809), .A2(n11811), .ZN(n11957) );
  NAND2_X1 U11956 ( .A1(n11809), .A2(n11811), .ZN(n11954) );
  NAND2_X1 U11957 ( .A1(n11958), .A2(n11959), .ZN(n11811) );
  NAND2_X1 U11958 ( .A1(n11808), .A2(n11960), .ZN(n11959) );
  OR2_X1 U11959 ( .A1(n11806), .A2(n11807), .ZN(n11960) );
  NOR2_X1 U11960 ( .A1(n11551), .A2(n7687), .ZN(n11808) );
  NAND2_X1 U11961 ( .A1(n11806), .A2(n11807), .ZN(n11958) );
  NAND2_X1 U11962 ( .A1(n11961), .A2(n11962), .ZN(n11807) );
  NAND2_X1 U11963 ( .A1(n11963), .A2(b_16_), .ZN(n11962) );
  NOR2_X1 U11964 ( .A1(n11964), .A2(n7676), .ZN(n11963) );
  NOR2_X1 U11965 ( .A1(n11801), .A2(n11803), .ZN(n11964) );
  NAND2_X1 U11966 ( .A1(n11801), .A2(n11803), .ZN(n11961) );
  NAND2_X1 U11967 ( .A1(n11965), .A2(n11966), .ZN(n11803) );
  NAND2_X1 U11968 ( .A1(n11800), .A2(n11967), .ZN(n11966) );
  OR2_X1 U11969 ( .A1(n11798), .A2(n11799), .ZN(n11967) );
  NOR2_X1 U11970 ( .A1(n11551), .A2(n7656), .ZN(n11800) );
  NAND2_X1 U11971 ( .A1(n11798), .A2(n11799), .ZN(n11965) );
  NAND2_X1 U11972 ( .A1(n11968), .A2(n11969), .ZN(n11799) );
  NAND2_X1 U11973 ( .A1(n11970), .A2(b_16_), .ZN(n11969) );
  NOR2_X1 U11974 ( .A1(n11971), .A2(n7645), .ZN(n11970) );
  NOR2_X1 U11975 ( .A1(n11794), .A2(n11795), .ZN(n11971) );
  NAND2_X1 U11976 ( .A1(n11794), .A2(n11795), .ZN(n11968) );
  NAND2_X1 U11977 ( .A1(n11972), .A2(n11973), .ZN(n11795) );
  NAND2_X1 U11978 ( .A1(n11792), .A2(n11974), .ZN(n11973) );
  OR2_X1 U11979 ( .A1(n11790), .A2(n11791), .ZN(n11974) );
  NOR2_X1 U11980 ( .A1(n11551), .A2(n7624), .ZN(n11792) );
  NAND2_X1 U11981 ( .A1(n11790), .A2(n11791), .ZN(n11972) );
  NAND2_X1 U11982 ( .A1(n11975), .A2(n11976), .ZN(n11791) );
  NAND2_X1 U11983 ( .A1(n11977), .A2(b_16_), .ZN(n11976) );
  NOR2_X1 U11984 ( .A1(n11978), .A2(n7613), .ZN(n11977) );
  NOR2_X1 U11985 ( .A1(n11787), .A2(n11785), .ZN(n11978) );
  NAND2_X1 U11986 ( .A1(n11785), .A2(n11787), .ZN(n11975) );
  NAND2_X1 U11987 ( .A1(n11979), .A2(n11980), .ZN(n11787) );
  NAND2_X1 U11988 ( .A1(n11784), .A2(n11981), .ZN(n11980) );
  OR2_X1 U11989 ( .A1(n11783), .A2(n11781), .ZN(n11981) );
  NOR2_X1 U11990 ( .A1(n11551), .A2(n7593), .ZN(n11784) );
  NAND2_X1 U11991 ( .A1(n11781), .A2(n11783), .ZN(n11979) );
  NAND2_X1 U11992 ( .A1(n11982), .A2(n11983), .ZN(n11783) );
  NAND2_X1 U11993 ( .A1(n11984), .A2(b_16_), .ZN(n11983) );
  NOR2_X1 U11994 ( .A1(n11985), .A2(n8052), .ZN(n11984) );
  NOR2_X1 U11995 ( .A1(n11780), .A2(n11778), .ZN(n11985) );
  NAND2_X1 U11996 ( .A1(n11778), .A2(n11780), .ZN(n11982) );
  NAND2_X1 U11997 ( .A1(n11986), .A2(n11987), .ZN(n11780) );
  NAND2_X1 U11998 ( .A1(n11776), .A2(n11988), .ZN(n11987) );
  NAND2_X1 U11999 ( .A1(n11775), .A2(n11774), .ZN(n11988) );
  NOR2_X1 U12000 ( .A1(n11551), .A2(n7563), .ZN(n11776) );
  OR2_X1 U12001 ( .A1(n11774), .A2(n11775), .ZN(n11986) );
  AND2_X1 U12002 ( .A1(n11771), .A2(n11989), .ZN(n11775) );
  NAND2_X1 U12003 ( .A1(n11770), .A2(n11772), .ZN(n11989) );
  NAND2_X1 U12004 ( .A1(n11990), .A2(n11991), .ZN(n11772) );
  NAND2_X1 U12005 ( .A1(b_16_), .A2(a_28_), .ZN(n11991) );
  INV_X1 U12006 ( .A(n11992), .ZN(n11990) );
  XOR2_X1 U12007 ( .A(n11993), .B(n11994), .Z(n11770) );
  NOR2_X1 U12008 ( .A1(n7529), .A2(n7755), .ZN(n11994) );
  XOR2_X1 U12009 ( .A(n11995), .B(n11996), .Z(n11993) );
  NAND2_X1 U12010 ( .A1(a_28_), .A2(n11992), .ZN(n11771) );
  NAND2_X1 U12011 ( .A1(n11997), .A2(n11998), .ZN(n11992) );
  NAND2_X1 U12012 ( .A1(n11999), .A2(b_16_), .ZN(n11998) );
  NOR2_X1 U12013 ( .A1(n12000), .A2(n7529), .ZN(n11999) );
  NOR2_X1 U12014 ( .A1(n11757), .A2(n11758), .ZN(n12000) );
  NAND2_X1 U12015 ( .A1(n11757), .A2(n11758), .ZN(n11997) );
  NAND2_X1 U12016 ( .A1(n12001), .A2(n12002), .ZN(n11758) );
  NAND2_X1 U12017 ( .A1(n12003), .A2(b_14_), .ZN(n12002) );
  NOR2_X1 U12018 ( .A1(n12004), .A2(n8048), .ZN(n12003) );
  NOR2_X1 U12019 ( .A1(n8676), .A2(n7755), .ZN(n12004) );
  NAND2_X1 U12020 ( .A1(n12005), .A2(b_15_), .ZN(n12001) );
  NOR2_X1 U12021 ( .A1(n12006), .A2(n7515), .ZN(n12005) );
  NOR2_X1 U12022 ( .A1(n8679), .A2(n8056), .ZN(n12006) );
  AND2_X1 U12023 ( .A1(n12007), .A2(b_15_), .ZN(n11757) );
  NOR2_X1 U12024 ( .A1(n8451), .A2(n11551), .ZN(n12007) );
  XOR2_X1 U12025 ( .A(n12008), .B(n12009), .Z(n11774) );
  NAND2_X1 U12026 ( .A1(n12010), .A2(n12011), .ZN(n12008) );
  XNOR2_X1 U12027 ( .A(n12012), .B(n12013), .ZN(n11778) );
  XNOR2_X1 U12028 ( .A(n12014), .B(n12015), .ZN(n12012) );
  XOR2_X1 U12029 ( .A(n12016), .B(n12017), .Z(n11781) );
  XNOR2_X1 U12030 ( .A(n12018), .B(n12019), .ZN(n12016) );
  NAND2_X1 U12031 ( .A1(b_15_), .A2(a_26_), .ZN(n12018) );
  XNOR2_X1 U12032 ( .A(n12020), .B(n12021), .ZN(n11785) );
  XOR2_X1 U12033 ( .A(n12022), .B(n12023), .Z(n12021) );
  NAND2_X1 U12034 ( .A1(b_15_), .A2(a_25_), .ZN(n12023) );
  XNOR2_X1 U12035 ( .A(n12024), .B(n12025), .ZN(n11790) );
  NAND2_X1 U12036 ( .A1(n12026), .A2(n12027), .ZN(n12024) );
  XOR2_X1 U12037 ( .A(n12028), .B(n12029), .Z(n11794) );
  XOR2_X1 U12038 ( .A(n12030), .B(n12031), .Z(n12028) );
  XOR2_X1 U12039 ( .A(n12032), .B(n12033), .Z(n11798) );
  XOR2_X1 U12040 ( .A(n12034), .B(n12035), .Z(n12032) );
  NOR2_X1 U12041 ( .A1(n7645), .A2(n7755), .ZN(n12035) );
  XOR2_X1 U12042 ( .A(n12036), .B(n12037), .Z(n11801) );
  XOR2_X1 U12043 ( .A(n12038), .B(n12039), .Z(n12036) );
  XNOR2_X1 U12044 ( .A(n12040), .B(n12041), .ZN(n11806) );
  XOR2_X1 U12045 ( .A(n12042), .B(n12043), .Z(n12041) );
  NAND2_X1 U12046 ( .A1(b_15_), .A2(a_20_), .ZN(n12043) );
  XOR2_X1 U12047 ( .A(n12044), .B(n12045), .Z(n11809) );
  XOR2_X1 U12048 ( .A(n12046), .B(n12047), .Z(n12044) );
  XNOR2_X1 U12049 ( .A(n12048), .B(n12049), .ZN(n11814) );
  XOR2_X1 U12050 ( .A(n12050), .B(n12051), .Z(n12049) );
  NAND2_X1 U12051 ( .A1(b_15_), .A2(a_18_), .ZN(n12051) );
  NOR2_X1 U12052 ( .A1(n11551), .A2(n7743), .ZN(n7737) );
  INV_X1 U12053 ( .A(b_16_), .ZN(n11551) );
  XNOR2_X1 U12054 ( .A(n12052), .B(n12053), .ZN(n11821) );
  XNOR2_X1 U12055 ( .A(n12054), .B(n12055), .ZN(n12053) );
  XOR2_X1 U12056 ( .A(n12056), .B(n12057), .Z(n11825) );
  XOR2_X1 U12057 ( .A(n12058), .B(n8015), .Z(n12057) );
  XNOR2_X1 U12058 ( .A(n12059), .B(n12060), .ZN(n11696) );
  XNOR2_X1 U12059 ( .A(n12061), .B(n12062), .ZN(n12059) );
  NAND2_X1 U12060 ( .A1(b_15_), .A2(a_14_), .ZN(n12061) );
  XOR2_X1 U12061 ( .A(n12063), .B(n12064), .Z(n11828) );
  XNOR2_X1 U12062 ( .A(n12065), .B(n12066), .ZN(n12063) );
  NAND2_X1 U12063 ( .A1(b_15_), .A2(a_13_), .ZN(n12065) );
  XNOR2_X1 U12064 ( .A(n12067), .B(n12068), .ZN(n11833) );
  XOR2_X1 U12065 ( .A(n12069), .B(n12070), .Z(n12067) );
  NOR2_X1 U12066 ( .A1(n7806), .A2(n7755), .ZN(n12070) );
  XOR2_X1 U12067 ( .A(n12071), .B(n12072), .Z(n11836) );
  XOR2_X1 U12068 ( .A(n12073), .B(n12074), .Z(n12071) );
  NOR2_X1 U12069 ( .A1(n7817), .A2(n7755), .ZN(n12074) );
  XNOR2_X1 U12070 ( .A(n12075), .B(n12076), .ZN(n11844) );
  XOR2_X1 U12071 ( .A(n12077), .B(n12078), .Z(n12076) );
  NAND2_X1 U12072 ( .A1(b_15_), .A2(a_9_), .ZN(n12078) );
  XOR2_X1 U12073 ( .A(n12079), .B(n12080), .Z(n11849) );
  XOR2_X1 U12074 ( .A(n12081), .B(n12082), .Z(n12079) );
  NOR2_X1 U12075 ( .A1(n8059), .A2(n7755), .ZN(n12082) );
  XNOR2_X1 U12076 ( .A(n12083), .B(n12084), .ZN(n11853) );
  XOR2_X1 U12077 ( .A(n12085), .B(n12086), .Z(n12083) );
  NOR2_X1 U12078 ( .A1(n7884), .A2(n7755), .ZN(n12086) );
  XOR2_X1 U12079 ( .A(n12087), .B(n12088), .Z(n11856) );
  XOR2_X1 U12080 ( .A(n12089), .B(n12090), .Z(n12087) );
  NOR2_X1 U12081 ( .A1(n8061), .A2(n7755), .ZN(n12090) );
  XOR2_X1 U12082 ( .A(n12091), .B(n12092), .Z(n11861) );
  XOR2_X1 U12083 ( .A(n12093), .B(n12094), .Z(n12091) );
  NOR2_X1 U12084 ( .A1(n7914), .A2(n7755), .ZN(n12094) );
  XOR2_X1 U12085 ( .A(n12095), .B(n12096), .Z(n11865) );
  XOR2_X1 U12086 ( .A(n12097), .B(n12098), .Z(n12095) );
  NOR2_X1 U12087 ( .A1(n7934), .A2(n7755), .ZN(n12098) );
  XOR2_X1 U12088 ( .A(n12099), .B(n12100), .Z(n11869) );
  NAND2_X1 U12089 ( .A1(n12101), .A2(n12102), .ZN(n12099) );
  XNOR2_X1 U12090 ( .A(n12103), .B(n12104), .ZN(n11873) );
  NAND2_X1 U12091 ( .A1(n12105), .A2(n12106), .ZN(n12103) );
  XNOR2_X1 U12092 ( .A(n12107), .B(n12108), .ZN(n11640) );
  XOR2_X1 U12093 ( .A(n12109), .B(n12110), .Z(n12107) );
  NOR2_X1 U12094 ( .A1(n7973), .A2(n7755), .ZN(n12110) );
  NAND2_X1 U12095 ( .A1(n12111), .A2(n12112), .ZN(n8167) );
  NAND2_X1 U12096 ( .A1(n11883), .A2(n11879), .ZN(n12112) );
  XOR2_X1 U12097 ( .A(n12113), .B(n8230), .Z(n12111) );
  NAND2_X1 U12098 ( .A1(n12114), .A2(n12115), .ZN(n8166) );
  XOR2_X1 U12099 ( .A(n8231), .B(n8230), .Z(n12115) );
  INV_X1 U12100 ( .A(n12116), .ZN(n8230) );
  AND2_X1 U12101 ( .A1(n11879), .A2(n11883), .ZN(n12114) );
  INV_X1 U12102 ( .A(n11880), .ZN(n11883) );
  XOR2_X1 U12103 ( .A(n12117), .B(n12118), .Z(n11880) );
  NAND2_X1 U12104 ( .A1(n12119), .A2(n12120), .ZN(n12117) );
  NAND2_X1 U12105 ( .A1(n12121), .A2(n12122), .ZN(n11879) );
  NAND2_X1 U12106 ( .A1(n12123), .A2(b_15_), .ZN(n12122) );
  NOR2_X1 U12107 ( .A1(n12124), .A2(n8307), .ZN(n12123) );
  NOR2_X1 U12108 ( .A1(n11885), .A2(n11886), .ZN(n12124) );
  NAND2_X1 U12109 ( .A1(n11885), .A2(n11886), .ZN(n12121) );
  NAND2_X1 U12110 ( .A1(n12125), .A2(n12126), .ZN(n11886) );
  NAND2_X1 U12111 ( .A1(n12127), .A2(b_15_), .ZN(n12126) );
  NOR2_X1 U12112 ( .A1(n12128), .A2(n7973), .ZN(n12127) );
  NOR2_X1 U12113 ( .A1(n12109), .A2(n12108), .ZN(n12128) );
  NAND2_X1 U12114 ( .A1(n12108), .A2(n12109), .ZN(n12125) );
  NAND2_X1 U12115 ( .A1(n12105), .A2(n12129), .ZN(n12109) );
  NAND2_X1 U12116 ( .A1(n12104), .A2(n12106), .ZN(n12129) );
  NAND2_X1 U12117 ( .A1(n12130), .A2(n12131), .ZN(n12106) );
  NAND2_X1 U12118 ( .A1(b_15_), .A2(a_2_), .ZN(n12131) );
  INV_X1 U12119 ( .A(n12132), .ZN(n12130) );
  XNOR2_X1 U12120 ( .A(n12133), .B(n12134), .ZN(n12104) );
  XNOR2_X1 U12121 ( .A(n12135), .B(n12136), .ZN(n12133) );
  NAND2_X1 U12122 ( .A1(a_2_), .A2(n12132), .ZN(n12105) );
  NAND2_X1 U12123 ( .A1(n12101), .A2(n12137), .ZN(n12132) );
  NAND2_X1 U12124 ( .A1(n12100), .A2(n12102), .ZN(n12137) );
  NAND2_X1 U12125 ( .A1(n12138), .A2(n12139), .ZN(n12102) );
  NAND2_X1 U12126 ( .A1(b_15_), .A2(a_3_), .ZN(n12139) );
  INV_X1 U12127 ( .A(n12140), .ZN(n12138) );
  XOR2_X1 U12128 ( .A(n12141), .B(n12142), .Z(n12100) );
  NOR2_X1 U12129 ( .A1(n12143), .A2(n12144), .ZN(n12142) );
  NOR2_X1 U12130 ( .A1(n12145), .A2(n12146), .ZN(n12143) );
  NOR2_X1 U12131 ( .A1(n7934), .A2(n8056), .ZN(n12145) );
  NAND2_X1 U12132 ( .A1(a_3_), .A2(n12140), .ZN(n12101) );
  NAND2_X1 U12133 ( .A1(n12147), .A2(n12148), .ZN(n12140) );
  NAND2_X1 U12134 ( .A1(n12149), .A2(b_15_), .ZN(n12148) );
  NOR2_X1 U12135 ( .A1(n12150), .A2(n7934), .ZN(n12149) );
  NOR2_X1 U12136 ( .A1(n12096), .A2(n12097), .ZN(n12150) );
  NAND2_X1 U12137 ( .A1(n12096), .A2(n12097), .ZN(n12147) );
  NAND2_X1 U12138 ( .A1(n12151), .A2(n12152), .ZN(n12097) );
  NAND2_X1 U12139 ( .A1(n12153), .A2(b_15_), .ZN(n12152) );
  NOR2_X1 U12140 ( .A1(n12154), .A2(n7914), .ZN(n12153) );
  NOR2_X1 U12141 ( .A1(n12092), .A2(n12093), .ZN(n12154) );
  NAND2_X1 U12142 ( .A1(n12092), .A2(n12093), .ZN(n12151) );
  NAND2_X1 U12143 ( .A1(n12155), .A2(n12156), .ZN(n12093) );
  NAND2_X1 U12144 ( .A1(n12157), .A2(b_15_), .ZN(n12156) );
  NOR2_X1 U12145 ( .A1(n12158), .A2(n8061), .ZN(n12157) );
  NOR2_X1 U12146 ( .A1(n12089), .A2(n12088), .ZN(n12158) );
  NAND2_X1 U12147 ( .A1(n12088), .A2(n12089), .ZN(n12155) );
  NAND2_X1 U12148 ( .A1(n12159), .A2(n12160), .ZN(n12089) );
  NAND2_X1 U12149 ( .A1(n12161), .A2(b_15_), .ZN(n12160) );
  NOR2_X1 U12150 ( .A1(n12162), .A2(n7884), .ZN(n12161) );
  NOR2_X1 U12151 ( .A1(n12085), .A2(n12084), .ZN(n12162) );
  NAND2_X1 U12152 ( .A1(n12084), .A2(n12085), .ZN(n12159) );
  NAND2_X1 U12153 ( .A1(n12163), .A2(n12164), .ZN(n12085) );
  NAND2_X1 U12154 ( .A1(n12165), .A2(b_15_), .ZN(n12164) );
  NOR2_X1 U12155 ( .A1(n12166), .A2(n8059), .ZN(n12165) );
  NOR2_X1 U12156 ( .A1(n12080), .A2(n12081), .ZN(n12166) );
  NAND2_X1 U12157 ( .A1(n12080), .A2(n12081), .ZN(n12163) );
  NAND2_X1 U12158 ( .A1(n12167), .A2(n12168), .ZN(n12081) );
  NAND2_X1 U12159 ( .A1(n12169), .A2(b_15_), .ZN(n12168) );
  NOR2_X1 U12160 ( .A1(n12170), .A2(n7848), .ZN(n12169) );
  NOR2_X1 U12161 ( .A1(n12075), .A2(n12077), .ZN(n12170) );
  NAND2_X1 U12162 ( .A1(n12075), .A2(n12077), .ZN(n12167) );
  NAND2_X1 U12163 ( .A1(n12171), .A2(n12172), .ZN(n12077) );
  NAND2_X1 U12164 ( .A1(n12173), .A2(b_15_), .ZN(n12172) );
  NOR2_X1 U12165 ( .A1(n12174), .A2(n7837), .ZN(n12173) );
  NOR2_X1 U12166 ( .A1(n11920), .A2(n11922), .ZN(n12174) );
  NAND2_X1 U12167 ( .A1(n11920), .A2(n11922), .ZN(n12171) );
  NAND2_X1 U12168 ( .A1(n12175), .A2(n12176), .ZN(n11922) );
  NAND2_X1 U12169 ( .A1(n12177), .A2(b_15_), .ZN(n12176) );
  NOR2_X1 U12170 ( .A1(n12178), .A2(n7817), .ZN(n12177) );
  NOR2_X1 U12171 ( .A1(n12073), .A2(n12072), .ZN(n12178) );
  NAND2_X1 U12172 ( .A1(n12072), .A2(n12073), .ZN(n12175) );
  NAND2_X1 U12173 ( .A1(n12179), .A2(n12180), .ZN(n12073) );
  NAND2_X1 U12174 ( .A1(n12181), .A2(b_15_), .ZN(n12180) );
  NOR2_X1 U12175 ( .A1(n12182), .A2(n7806), .ZN(n12181) );
  NOR2_X1 U12176 ( .A1(n12069), .A2(n12068), .ZN(n12182) );
  NAND2_X1 U12177 ( .A1(n12068), .A2(n12069), .ZN(n12179) );
  NAND2_X1 U12178 ( .A1(n12183), .A2(n12184), .ZN(n12069) );
  NAND2_X1 U12179 ( .A1(n12185), .A2(b_15_), .ZN(n12184) );
  NOR2_X1 U12180 ( .A1(n12186), .A2(n7786), .ZN(n12185) );
  NOR2_X1 U12181 ( .A1(n12064), .A2(n12066), .ZN(n12186) );
  NAND2_X1 U12182 ( .A1(n12064), .A2(n12066), .ZN(n12183) );
  NAND2_X1 U12183 ( .A1(n12187), .A2(n12188), .ZN(n12066) );
  NAND2_X1 U12184 ( .A1(n12189), .A2(b_15_), .ZN(n12188) );
  NOR2_X1 U12185 ( .A1(n12190), .A2(n7775), .ZN(n12189) );
  NOR2_X1 U12186 ( .A1(n12062), .A2(n12060), .ZN(n12190) );
  NAND2_X1 U12187 ( .A1(n12060), .A2(n12062), .ZN(n12187) );
  NAND2_X1 U12188 ( .A1(n12191), .A2(n12192), .ZN(n12062) );
  NAND2_X1 U12189 ( .A1(n12056), .A2(n12193), .ZN(n12192) );
  OR2_X1 U12190 ( .A1(n12058), .A2(n7749), .ZN(n12193) );
  XNOR2_X1 U12191 ( .A(n12194), .B(n12195), .ZN(n12056) );
  XNOR2_X1 U12192 ( .A(n12196), .B(n12197), .ZN(n12194) );
  NAND2_X1 U12193 ( .A1(n7749), .A2(n12058), .ZN(n12191) );
  NAND2_X1 U12194 ( .A1(n12198), .A2(n12199), .ZN(n12058) );
  NAND2_X1 U12195 ( .A1(n12055), .A2(n12200), .ZN(n12199) );
  OR2_X1 U12196 ( .A1(n12054), .A2(n12052), .ZN(n12200) );
  NOR2_X1 U12197 ( .A1(n7755), .A2(n7743), .ZN(n12055) );
  NAND2_X1 U12198 ( .A1(n12052), .A2(n12054), .ZN(n12198) );
  NAND2_X1 U12199 ( .A1(n12201), .A2(n12202), .ZN(n12054) );
  NAND2_X1 U12200 ( .A1(n11950), .A2(n12203), .ZN(n12202) );
  OR2_X1 U12201 ( .A1(n11948), .A2(n11949), .ZN(n12203) );
  NOR2_X1 U12202 ( .A1(n7755), .A2(n7723), .ZN(n11950) );
  NAND2_X1 U12203 ( .A1(n11948), .A2(n11949), .ZN(n12201) );
  NAND2_X1 U12204 ( .A1(n12204), .A2(n12205), .ZN(n11949) );
  NAND2_X1 U12205 ( .A1(n12206), .A2(b_15_), .ZN(n12205) );
  NOR2_X1 U12206 ( .A1(n12207), .A2(n7707), .ZN(n12206) );
  NOR2_X1 U12207 ( .A1(n12048), .A2(n12050), .ZN(n12207) );
  NAND2_X1 U12208 ( .A1(n12048), .A2(n12050), .ZN(n12204) );
  NAND2_X1 U12209 ( .A1(n12208), .A2(n12209), .ZN(n12050) );
  NAND2_X1 U12210 ( .A1(n12047), .A2(n12210), .ZN(n12209) );
  OR2_X1 U12211 ( .A1(n12045), .A2(n12046), .ZN(n12210) );
  NOR2_X1 U12212 ( .A1(n7755), .A2(n7687), .ZN(n12047) );
  NAND2_X1 U12213 ( .A1(n12045), .A2(n12046), .ZN(n12208) );
  NAND2_X1 U12214 ( .A1(n12211), .A2(n12212), .ZN(n12046) );
  NAND2_X1 U12215 ( .A1(n12213), .A2(b_15_), .ZN(n12212) );
  NOR2_X1 U12216 ( .A1(n12214), .A2(n7676), .ZN(n12213) );
  NOR2_X1 U12217 ( .A1(n12040), .A2(n12042), .ZN(n12214) );
  NAND2_X1 U12218 ( .A1(n12040), .A2(n12042), .ZN(n12211) );
  NAND2_X1 U12219 ( .A1(n12215), .A2(n12216), .ZN(n12042) );
  NAND2_X1 U12220 ( .A1(n12039), .A2(n12217), .ZN(n12216) );
  OR2_X1 U12221 ( .A1(n12037), .A2(n12038), .ZN(n12217) );
  NOR2_X1 U12222 ( .A1(n7755), .A2(n7656), .ZN(n12039) );
  NAND2_X1 U12223 ( .A1(n12037), .A2(n12038), .ZN(n12215) );
  NAND2_X1 U12224 ( .A1(n12218), .A2(n12219), .ZN(n12038) );
  NAND2_X1 U12225 ( .A1(n12220), .A2(b_15_), .ZN(n12219) );
  NOR2_X1 U12226 ( .A1(n12221), .A2(n7645), .ZN(n12220) );
  NOR2_X1 U12227 ( .A1(n12033), .A2(n12034), .ZN(n12221) );
  NAND2_X1 U12228 ( .A1(n12033), .A2(n12034), .ZN(n12218) );
  NAND2_X1 U12229 ( .A1(n12222), .A2(n12223), .ZN(n12034) );
  NAND2_X1 U12230 ( .A1(n12031), .A2(n12224), .ZN(n12223) );
  OR2_X1 U12231 ( .A1(n12029), .A2(n12030), .ZN(n12224) );
  NOR2_X1 U12232 ( .A1(n7755), .A2(n7624), .ZN(n12031) );
  NAND2_X1 U12233 ( .A1(n12029), .A2(n12030), .ZN(n12222) );
  NAND2_X1 U12234 ( .A1(n12026), .A2(n12225), .ZN(n12030) );
  NAND2_X1 U12235 ( .A1(n12025), .A2(n12027), .ZN(n12225) );
  NAND2_X1 U12236 ( .A1(n12226), .A2(n12227), .ZN(n12027) );
  NAND2_X1 U12237 ( .A1(b_15_), .A2(a_24_), .ZN(n12227) );
  INV_X1 U12238 ( .A(n12228), .ZN(n12226) );
  XOR2_X1 U12239 ( .A(n12229), .B(n12230), .Z(n12025) );
  XOR2_X1 U12240 ( .A(n12231), .B(n12232), .Z(n12229) );
  NOR2_X1 U12241 ( .A1(n7593), .A2(n8056), .ZN(n12232) );
  NAND2_X1 U12242 ( .A1(a_24_), .A2(n12228), .ZN(n12026) );
  NAND2_X1 U12243 ( .A1(n12233), .A2(n12234), .ZN(n12228) );
  NAND2_X1 U12244 ( .A1(n12235), .A2(b_15_), .ZN(n12234) );
  NOR2_X1 U12245 ( .A1(n12236), .A2(n7593), .ZN(n12235) );
  NOR2_X1 U12246 ( .A1(n12020), .A2(n12022), .ZN(n12236) );
  NAND2_X1 U12247 ( .A1(n12020), .A2(n12022), .ZN(n12233) );
  NAND2_X1 U12248 ( .A1(n12237), .A2(n12238), .ZN(n12022) );
  NAND2_X1 U12249 ( .A1(n12239), .A2(b_15_), .ZN(n12238) );
  NOR2_X1 U12250 ( .A1(n12240), .A2(n8052), .ZN(n12239) );
  NOR2_X1 U12251 ( .A1(n12019), .A2(n12017), .ZN(n12240) );
  NAND2_X1 U12252 ( .A1(n12017), .A2(n12019), .ZN(n12237) );
  NAND2_X1 U12253 ( .A1(n12241), .A2(n12242), .ZN(n12019) );
  NAND2_X1 U12254 ( .A1(n12015), .A2(n12243), .ZN(n12242) );
  NAND2_X1 U12255 ( .A1(n12014), .A2(n12013), .ZN(n12243) );
  NOR2_X1 U12256 ( .A1(n7755), .A2(n7563), .ZN(n12015) );
  INV_X1 U12257 ( .A(b_15_), .ZN(n7755) );
  OR2_X1 U12258 ( .A1(n12013), .A2(n12014), .ZN(n12241) );
  AND2_X1 U12259 ( .A1(n12010), .A2(n12244), .ZN(n12014) );
  NAND2_X1 U12260 ( .A1(n12009), .A2(n12011), .ZN(n12244) );
  NAND2_X1 U12261 ( .A1(n12245), .A2(n12246), .ZN(n12011) );
  NAND2_X1 U12262 ( .A1(b_15_), .A2(a_28_), .ZN(n12246) );
  INV_X1 U12263 ( .A(n12247), .ZN(n12245) );
  XOR2_X1 U12264 ( .A(n12248), .B(n12249), .Z(n12009) );
  NOR2_X1 U12265 ( .A1(n7529), .A2(n8056), .ZN(n12249) );
  XOR2_X1 U12266 ( .A(n12250), .B(n12251), .Z(n12248) );
  NAND2_X1 U12267 ( .A1(a_28_), .A2(n12247), .ZN(n12010) );
  NAND2_X1 U12268 ( .A1(n12252), .A2(n12253), .ZN(n12247) );
  NAND2_X1 U12269 ( .A1(n12254), .A2(b_15_), .ZN(n12253) );
  NOR2_X1 U12270 ( .A1(n12255), .A2(n7529), .ZN(n12254) );
  NOR2_X1 U12271 ( .A1(n11995), .A2(n11996), .ZN(n12255) );
  NAND2_X1 U12272 ( .A1(n11995), .A2(n11996), .ZN(n12252) );
  NAND2_X1 U12273 ( .A1(n12256), .A2(n12257), .ZN(n11996) );
  NAND2_X1 U12274 ( .A1(n12258), .A2(b_13_), .ZN(n12257) );
  NOR2_X1 U12275 ( .A1(n12259), .A2(n8048), .ZN(n12258) );
  NOR2_X1 U12276 ( .A1(n8676), .A2(n8056), .ZN(n12259) );
  NAND2_X1 U12277 ( .A1(n12260), .A2(b_14_), .ZN(n12256) );
  NOR2_X1 U12278 ( .A1(n12261), .A2(n7515), .ZN(n12260) );
  NOR2_X1 U12279 ( .A1(n8679), .A2(n7787), .ZN(n12261) );
  AND2_X1 U12280 ( .A1(n12262), .A2(b_15_), .ZN(n11995) );
  NOR2_X1 U12281 ( .A1(n8451), .A2(n8056), .ZN(n12262) );
  XOR2_X1 U12282 ( .A(n12263), .B(n12264), .Z(n12013) );
  NAND2_X1 U12283 ( .A1(n12265), .A2(n12266), .ZN(n12263) );
  XNOR2_X1 U12284 ( .A(n12267), .B(n12268), .ZN(n12017) );
  XNOR2_X1 U12285 ( .A(n12269), .B(n12270), .ZN(n12267) );
  XOR2_X1 U12286 ( .A(n12271), .B(n12272), .Z(n12020) );
  XNOR2_X1 U12287 ( .A(n12273), .B(n12274), .ZN(n12271) );
  NAND2_X1 U12288 ( .A1(b_14_), .A2(a_26_), .ZN(n12273) );
  XNOR2_X1 U12289 ( .A(n12275), .B(n12276), .ZN(n12029) );
  NAND2_X1 U12290 ( .A1(n12277), .A2(n12278), .ZN(n12275) );
  XOR2_X1 U12291 ( .A(n12279), .B(n12280), .Z(n12033) );
  XOR2_X1 U12292 ( .A(n12281), .B(n12282), .Z(n12279) );
  XOR2_X1 U12293 ( .A(n12283), .B(n12284), .Z(n12037) );
  XOR2_X1 U12294 ( .A(n12285), .B(n12286), .Z(n12283) );
  NOR2_X1 U12295 ( .A1(n7645), .A2(n8056), .ZN(n12286) );
  XOR2_X1 U12296 ( .A(n12287), .B(n12288), .Z(n12040) );
  XOR2_X1 U12297 ( .A(n12289), .B(n12290), .Z(n12287) );
  XNOR2_X1 U12298 ( .A(n12291), .B(n12292), .ZN(n12045) );
  XOR2_X1 U12299 ( .A(n12293), .B(n12294), .Z(n12292) );
  NAND2_X1 U12300 ( .A1(b_14_), .A2(a_20_), .ZN(n12294) );
  XOR2_X1 U12301 ( .A(n12295), .B(n12296), .Z(n12048) );
  XOR2_X1 U12302 ( .A(n12297), .B(n12298), .Z(n12295) );
  XOR2_X1 U12303 ( .A(n12299), .B(n12300), .Z(n11948) );
  XOR2_X1 U12304 ( .A(n12301), .B(n12302), .Z(n12299) );
  NOR2_X1 U12305 ( .A1(n7707), .A2(n8056), .ZN(n12302) );
  XOR2_X1 U12306 ( .A(n12303), .B(n12304), .Z(n12052) );
  XOR2_X1 U12307 ( .A(n12305), .B(n12306), .Z(n12303) );
  NOR2_X1 U12308 ( .A1(n7723), .A2(n8056), .ZN(n12306) );
  INV_X1 U12309 ( .A(n8015), .ZN(n7749) );
  NAND2_X1 U12310 ( .A1(b_15_), .A2(a_15_), .ZN(n8015) );
  XNOR2_X1 U12311 ( .A(n12307), .B(n12308), .ZN(n12060) );
  XNOR2_X1 U12312 ( .A(n12309), .B(n12310), .ZN(n12307) );
  XNOR2_X1 U12313 ( .A(n12311), .B(n12312), .ZN(n12064) );
  XOR2_X1 U12314 ( .A(n12313), .B(n12314), .Z(n12311) );
  XOR2_X1 U12315 ( .A(n12315), .B(n12316), .Z(n12068) );
  XNOR2_X1 U12316 ( .A(n12317), .B(n12318), .ZN(n12316) );
  NAND2_X1 U12317 ( .A1(b_14_), .A2(a_13_), .ZN(n12318) );
  XNOR2_X1 U12318 ( .A(n12319), .B(n12320), .ZN(n12072) );
  NAND2_X1 U12319 ( .A1(n12321), .A2(n12322), .ZN(n12319) );
  XNOR2_X1 U12320 ( .A(n12323), .B(n12324), .ZN(n11920) );
  NAND2_X1 U12321 ( .A1(n12325), .A2(n12326), .ZN(n12323) );
  XNOR2_X1 U12322 ( .A(n12327), .B(n12328), .ZN(n12075) );
  NAND2_X1 U12323 ( .A1(n12329), .A2(n12330), .ZN(n12327) );
  XNOR2_X1 U12324 ( .A(n12331), .B(n12332), .ZN(n12080) );
  NAND2_X1 U12325 ( .A1(n12333), .A2(n12334), .ZN(n12331) );
  XNOR2_X1 U12326 ( .A(n12335), .B(n12336), .ZN(n12084) );
  NAND2_X1 U12327 ( .A1(n12337), .A2(n12338), .ZN(n12335) );
  XNOR2_X1 U12328 ( .A(n12339), .B(n12340), .ZN(n12088) );
  NAND2_X1 U12329 ( .A1(n12341), .A2(n12342), .ZN(n12339) );
  XNOR2_X1 U12330 ( .A(n12343), .B(n12344), .ZN(n12092) );
  NAND2_X1 U12331 ( .A1(n12345), .A2(n12346), .ZN(n12343) );
  XNOR2_X1 U12332 ( .A(n12347), .B(n12348), .ZN(n12096) );
  NAND2_X1 U12333 ( .A1(n12349), .A2(n12350), .ZN(n12347) );
  XOR2_X1 U12334 ( .A(n12351), .B(n12352), .Z(n12108) );
  XOR2_X1 U12335 ( .A(n12353), .B(n12354), .Z(n12351) );
  NOR2_X1 U12336 ( .A1(n7965), .A2(n8056), .ZN(n12354) );
  XNOR2_X1 U12337 ( .A(n12355), .B(n12356), .ZN(n11885) );
  NAND2_X1 U12338 ( .A1(n12357), .A2(n12358), .ZN(n12355) );
  NAND2_X1 U12339 ( .A1(n12359), .A2(n12360), .ZN(n8171) );
  NOR2_X1 U12340 ( .A1(n8227), .A2(n12113), .ZN(n12360) );
  INV_X1 U12341 ( .A(n8231), .ZN(n12113) );
  NAND2_X1 U12342 ( .A1(n12119), .A2(n12361), .ZN(n8231) );
  NAND2_X1 U12343 ( .A1(n12118), .A2(n12120), .ZN(n12361) );
  NAND2_X1 U12344 ( .A1(n12362), .A2(n12363), .ZN(n12120) );
  NAND2_X1 U12345 ( .A1(b_14_), .A2(a_0_), .ZN(n12363) );
  INV_X1 U12346 ( .A(n12364), .ZN(n12362) );
  XOR2_X1 U12347 ( .A(n12365), .B(n12366), .Z(n12118) );
  XOR2_X1 U12348 ( .A(n12367), .B(n12368), .Z(n12365) );
  NOR2_X1 U12349 ( .A1(n7973), .A2(n7787), .ZN(n12368) );
  NAND2_X1 U12350 ( .A1(a_0_), .A2(n12364), .ZN(n12119) );
  NAND2_X1 U12351 ( .A1(n12357), .A2(n12369), .ZN(n12364) );
  NAND2_X1 U12352 ( .A1(n12356), .A2(n12358), .ZN(n12369) );
  NAND2_X1 U12353 ( .A1(n12370), .A2(n12371), .ZN(n12358) );
  NAND2_X1 U12354 ( .A1(b_14_), .A2(a_1_), .ZN(n12371) );
  INV_X1 U12355 ( .A(n12372), .ZN(n12370) );
  XNOR2_X1 U12356 ( .A(n12373), .B(n12374), .ZN(n12356) );
  XOR2_X1 U12357 ( .A(n12375), .B(n12376), .Z(n12374) );
  NAND2_X1 U12358 ( .A1(b_13_), .A2(a_2_), .ZN(n12376) );
  NAND2_X1 U12359 ( .A1(a_1_), .A2(n12372), .ZN(n12357) );
  NAND2_X1 U12360 ( .A1(n12377), .A2(n12378), .ZN(n12372) );
  NAND2_X1 U12361 ( .A1(n12379), .A2(b_14_), .ZN(n12378) );
  NOR2_X1 U12362 ( .A1(n12380), .A2(n7965), .ZN(n12379) );
  NOR2_X1 U12363 ( .A1(n12352), .A2(n12353), .ZN(n12380) );
  NAND2_X1 U12364 ( .A1(n12352), .A2(n12353), .ZN(n12377) );
  NAND2_X1 U12365 ( .A1(n12381), .A2(n12382), .ZN(n12353) );
  NAND2_X1 U12366 ( .A1(n12136), .A2(n12383), .ZN(n12382) );
  NAND2_X1 U12367 ( .A1(n12135), .A2(n12134), .ZN(n12383) );
  NOR2_X1 U12368 ( .A1(n8056), .A2(n7945), .ZN(n12136) );
  OR2_X1 U12369 ( .A1(n12134), .A2(n12135), .ZN(n12381) );
  NOR2_X1 U12370 ( .A1(n12144), .A2(n12384), .ZN(n12135) );
  AND2_X1 U12371 ( .A1(n12141), .A2(n12385), .ZN(n12384) );
  NAND2_X1 U12372 ( .A1(n12386), .A2(n12387), .ZN(n12385) );
  NAND2_X1 U12373 ( .A1(b_14_), .A2(a_4_), .ZN(n12387) );
  XOR2_X1 U12374 ( .A(n12388), .B(n12389), .Z(n12141) );
  XOR2_X1 U12375 ( .A(n12390), .B(n12391), .Z(n12388) );
  NOR2_X1 U12376 ( .A1(n7914), .A2(n7787), .ZN(n12391) );
  NOR2_X1 U12377 ( .A1(n7934), .A2(n12386), .ZN(n12144) );
  INV_X1 U12378 ( .A(n12146), .ZN(n12386) );
  NAND2_X1 U12379 ( .A1(n12349), .A2(n12392), .ZN(n12146) );
  NAND2_X1 U12380 ( .A1(n12348), .A2(n12350), .ZN(n12392) );
  NAND2_X1 U12381 ( .A1(n12393), .A2(n12394), .ZN(n12350) );
  NAND2_X1 U12382 ( .A1(b_14_), .A2(a_5_), .ZN(n12394) );
  INV_X1 U12383 ( .A(n12395), .ZN(n12393) );
  XNOR2_X1 U12384 ( .A(n12396), .B(n12397), .ZN(n12348) );
  XOR2_X1 U12385 ( .A(n12398), .B(n12399), .Z(n12397) );
  NAND2_X1 U12386 ( .A1(b_13_), .A2(a_6_), .ZN(n12399) );
  NAND2_X1 U12387 ( .A1(a_5_), .A2(n12395), .ZN(n12349) );
  NAND2_X1 U12388 ( .A1(n12345), .A2(n12400), .ZN(n12395) );
  NAND2_X1 U12389 ( .A1(n12344), .A2(n12346), .ZN(n12400) );
  NAND2_X1 U12390 ( .A1(n12401), .A2(n12402), .ZN(n12346) );
  NAND2_X1 U12391 ( .A1(b_14_), .A2(a_6_), .ZN(n12402) );
  INV_X1 U12392 ( .A(n12403), .ZN(n12401) );
  XNOR2_X1 U12393 ( .A(n12404), .B(n12405), .ZN(n12344) );
  XOR2_X1 U12394 ( .A(n12406), .B(n12407), .Z(n12405) );
  NAND2_X1 U12395 ( .A1(b_13_), .A2(a_7_), .ZN(n12407) );
  NAND2_X1 U12396 ( .A1(a_6_), .A2(n12403), .ZN(n12345) );
  NAND2_X1 U12397 ( .A1(n12341), .A2(n12408), .ZN(n12403) );
  NAND2_X1 U12398 ( .A1(n12340), .A2(n12342), .ZN(n12408) );
  NAND2_X1 U12399 ( .A1(n12409), .A2(n12410), .ZN(n12342) );
  NAND2_X1 U12400 ( .A1(b_14_), .A2(a_7_), .ZN(n12410) );
  INV_X1 U12401 ( .A(n12411), .ZN(n12409) );
  XNOR2_X1 U12402 ( .A(n12412), .B(n12413), .ZN(n12340) );
  XOR2_X1 U12403 ( .A(n12414), .B(n12415), .Z(n12413) );
  NAND2_X1 U12404 ( .A1(b_13_), .A2(a_8_), .ZN(n12415) );
  NAND2_X1 U12405 ( .A1(a_7_), .A2(n12411), .ZN(n12341) );
  NAND2_X1 U12406 ( .A1(n12337), .A2(n12416), .ZN(n12411) );
  NAND2_X1 U12407 ( .A1(n12336), .A2(n12338), .ZN(n12416) );
  NAND2_X1 U12408 ( .A1(n12417), .A2(n12418), .ZN(n12338) );
  NAND2_X1 U12409 ( .A1(b_14_), .A2(a_8_), .ZN(n12418) );
  INV_X1 U12410 ( .A(n12419), .ZN(n12417) );
  XNOR2_X1 U12411 ( .A(n12420), .B(n12421), .ZN(n12336) );
  XOR2_X1 U12412 ( .A(n12422), .B(n12423), .Z(n12421) );
  NAND2_X1 U12413 ( .A1(b_13_), .A2(a_9_), .ZN(n12423) );
  NAND2_X1 U12414 ( .A1(a_8_), .A2(n12419), .ZN(n12337) );
  NAND2_X1 U12415 ( .A1(n12333), .A2(n12424), .ZN(n12419) );
  NAND2_X1 U12416 ( .A1(n12332), .A2(n12334), .ZN(n12424) );
  NAND2_X1 U12417 ( .A1(n12425), .A2(n12426), .ZN(n12334) );
  NAND2_X1 U12418 ( .A1(b_14_), .A2(a_9_), .ZN(n12426) );
  INV_X1 U12419 ( .A(n12427), .ZN(n12425) );
  XNOR2_X1 U12420 ( .A(n12428), .B(n12429), .ZN(n12332) );
  XOR2_X1 U12421 ( .A(n12430), .B(n12431), .Z(n12429) );
  NAND2_X1 U12422 ( .A1(b_13_), .A2(a_10_), .ZN(n12431) );
  NAND2_X1 U12423 ( .A1(a_9_), .A2(n12427), .ZN(n12333) );
  NAND2_X1 U12424 ( .A1(n12329), .A2(n12432), .ZN(n12427) );
  NAND2_X1 U12425 ( .A1(n12328), .A2(n12330), .ZN(n12432) );
  NAND2_X1 U12426 ( .A1(n12433), .A2(n12434), .ZN(n12330) );
  NAND2_X1 U12427 ( .A1(b_14_), .A2(a_10_), .ZN(n12434) );
  INV_X1 U12428 ( .A(n12435), .ZN(n12433) );
  XNOR2_X1 U12429 ( .A(n12436), .B(n12437), .ZN(n12328) );
  XOR2_X1 U12430 ( .A(n12438), .B(n12439), .Z(n12437) );
  NAND2_X1 U12431 ( .A1(b_13_), .A2(a_11_), .ZN(n12439) );
  NAND2_X1 U12432 ( .A1(a_10_), .A2(n12435), .ZN(n12329) );
  NAND2_X1 U12433 ( .A1(n12325), .A2(n12440), .ZN(n12435) );
  NAND2_X1 U12434 ( .A1(n12324), .A2(n12326), .ZN(n12440) );
  NAND2_X1 U12435 ( .A1(n12441), .A2(n12442), .ZN(n12326) );
  NAND2_X1 U12436 ( .A1(b_14_), .A2(a_11_), .ZN(n12442) );
  INV_X1 U12437 ( .A(n12443), .ZN(n12441) );
  XOR2_X1 U12438 ( .A(n12444), .B(n12445), .Z(n12324) );
  XOR2_X1 U12439 ( .A(n12446), .B(n12447), .Z(n12444) );
  NOR2_X1 U12440 ( .A1(n7806), .A2(n7787), .ZN(n12447) );
  NAND2_X1 U12441 ( .A1(a_11_), .A2(n12443), .ZN(n12325) );
  NAND2_X1 U12442 ( .A1(n12321), .A2(n12448), .ZN(n12443) );
  NAND2_X1 U12443 ( .A1(n12320), .A2(n12322), .ZN(n12448) );
  NAND2_X1 U12444 ( .A1(n12449), .A2(n12450), .ZN(n12322) );
  NAND2_X1 U12445 ( .A1(b_14_), .A2(a_12_), .ZN(n12450) );
  INV_X1 U12446 ( .A(n12451), .ZN(n12449) );
  XOR2_X1 U12447 ( .A(n12452), .B(n12453), .Z(n12320) );
  XOR2_X1 U12448 ( .A(n12454), .B(n7781), .Z(n12452) );
  NAND2_X1 U12449 ( .A1(a_12_), .A2(n12451), .ZN(n12321) );
  NAND2_X1 U12450 ( .A1(n12455), .A2(n12456), .ZN(n12451) );
  NAND2_X1 U12451 ( .A1(n12457), .A2(b_14_), .ZN(n12456) );
  NOR2_X1 U12452 ( .A1(n12458), .A2(n7786), .ZN(n12457) );
  NOR2_X1 U12453 ( .A1(n12317), .A2(n12315), .ZN(n12458) );
  NAND2_X1 U12454 ( .A1(n12317), .A2(n12315), .ZN(n12455) );
  XOR2_X1 U12455 ( .A(n12459), .B(n12460), .Z(n12315) );
  XOR2_X1 U12456 ( .A(n12461), .B(n12462), .Z(n12459) );
  NOR2_X1 U12457 ( .A1(n7775), .A2(n7787), .ZN(n12462) );
  AND2_X1 U12458 ( .A1(n12463), .A2(n12464), .ZN(n12317) );
  NAND2_X1 U12459 ( .A1(n12312), .A2(n12465), .ZN(n12464) );
  NAND2_X1 U12460 ( .A1(n12314), .A2(n12313), .ZN(n12465) );
  XNOR2_X1 U12461 ( .A(n12466), .B(n12467), .ZN(n12312) );
  XOR2_X1 U12462 ( .A(n12468), .B(n12469), .Z(n12466) );
  NOR2_X1 U12463 ( .A1(n7754), .A2(n7787), .ZN(n12469) );
  OR2_X1 U12464 ( .A1(n12313), .A2(n12314), .ZN(n12463) );
  INV_X1 U12465 ( .A(n7769), .ZN(n12314) );
  NAND2_X1 U12466 ( .A1(b_14_), .A2(a_14_), .ZN(n7769) );
  NAND2_X1 U12467 ( .A1(n12470), .A2(n12471), .ZN(n12313) );
  NAND2_X1 U12468 ( .A1(n12310), .A2(n12472), .ZN(n12471) );
  NAND2_X1 U12469 ( .A1(n12309), .A2(n12308), .ZN(n12472) );
  NOR2_X1 U12470 ( .A1(n8056), .A2(n7754), .ZN(n12310) );
  OR2_X1 U12471 ( .A1(n12308), .A2(n12309), .ZN(n12470) );
  AND2_X1 U12472 ( .A1(n12473), .A2(n12474), .ZN(n12309) );
  NAND2_X1 U12473 ( .A1(n12197), .A2(n12475), .ZN(n12474) );
  NAND2_X1 U12474 ( .A1(n12196), .A2(n12195), .ZN(n12475) );
  NOR2_X1 U12475 ( .A1(n8056), .A2(n7743), .ZN(n12197) );
  OR2_X1 U12476 ( .A1(n12195), .A2(n12196), .ZN(n12473) );
  AND2_X1 U12477 ( .A1(n12476), .A2(n12477), .ZN(n12196) );
  NAND2_X1 U12478 ( .A1(n12478), .A2(b_14_), .ZN(n12477) );
  NOR2_X1 U12479 ( .A1(n12479), .A2(n7723), .ZN(n12478) );
  NOR2_X1 U12480 ( .A1(n12304), .A2(n12305), .ZN(n12479) );
  NAND2_X1 U12481 ( .A1(n12304), .A2(n12305), .ZN(n12476) );
  NAND2_X1 U12482 ( .A1(n12480), .A2(n12481), .ZN(n12305) );
  NAND2_X1 U12483 ( .A1(n12482), .A2(b_14_), .ZN(n12481) );
  NOR2_X1 U12484 ( .A1(n12483), .A2(n7707), .ZN(n12482) );
  NOR2_X1 U12485 ( .A1(n12300), .A2(n12301), .ZN(n12483) );
  NAND2_X1 U12486 ( .A1(n12300), .A2(n12301), .ZN(n12480) );
  NAND2_X1 U12487 ( .A1(n12484), .A2(n12485), .ZN(n12301) );
  NAND2_X1 U12488 ( .A1(n12298), .A2(n12486), .ZN(n12485) );
  OR2_X1 U12489 ( .A1(n12297), .A2(n12296), .ZN(n12486) );
  NOR2_X1 U12490 ( .A1(n8056), .A2(n7687), .ZN(n12298) );
  NAND2_X1 U12491 ( .A1(n12296), .A2(n12297), .ZN(n12484) );
  NAND2_X1 U12492 ( .A1(n12487), .A2(n12488), .ZN(n12297) );
  NAND2_X1 U12493 ( .A1(n12489), .A2(b_14_), .ZN(n12488) );
  NOR2_X1 U12494 ( .A1(n12490), .A2(n7676), .ZN(n12489) );
  NOR2_X1 U12495 ( .A1(n12291), .A2(n12293), .ZN(n12490) );
  NAND2_X1 U12496 ( .A1(n12291), .A2(n12293), .ZN(n12487) );
  NAND2_X1 U12497 ( .A1(n12491), .A2(n12492), .ZN(n12293) );
  NAND2_X1 U12498 ( .A1(n12290), .A2(n12493), .ZN(n12492) );
  OR2_X1 U12499 ( .A1(n12289), .A2(n12288), .ZN(n12493) );
  NOR2_X1 U12500 ( .A1(n8056), .A2(n7656), .ZN(n12290) );
  NAND2_X1 U12501 ( .A1(n12288), .A2(n12289), .ZN(n12491) );
  NAND2_X1 U12502 ( .A1(n12494), .A2(n12495), .ZN(n12289) );
  NAND2_X1 U12503 ( .A1(n12496), .A2(b_14_), .ZN(n12495) );
  NOR2_X1 U12504 ( .A1(n12497), .A2(n7645), .ZN(n12496) );
  NOR2_X1 U12505 ( .A1(n12284), .A2(n12285), .ZN(n12497) );
  NAND2_X1 U12506 ( .A1(n12284), .A2(n12285), .ZN(n12494) );
  NAND2_X1 U12507 ( .A1(n12498), .A2(n12499), .ZN(n12285) );
  NAND2_X1 U12508 ( .A1(n12282), .A2(n12500), .ZN(n12499) );
  OR2_X1 U12509 ( .A1(n12281), .A2(n12280), .ZN(n12500) );
  NOR2_X1 U12510 ( .A1(n8056), .A2(n7624), .ZN(n12282) );
  NAND2_X1 U12511 ( .A1(n12280), .A2(n12281), .ZN(n12498) );
  NAND2_X1 U12512 ( .A1(n12277), .A2(n12501), .ZN(n12281) );
  NAND2_X1 U12513 ( .A1(n12276), .A2(n12278), .ZN(n12501) );
  NAND2_X1 U12514 ( .A1(n12502), .A2(n12503), .ZN(n12278) );
  NAND2_X1 U12515 ( .A1(b_14_), .A2(a_24_), .ZN(n12503) );
  INV_X1 U12516 ( .A(n12504), .ZN(n12502) );
  XOR2_X1 U12517 ( .A(n12505), .B(n12506), .Z(n12276) );
  XOR2_X1 U12518 ( .A(n12507), .B(n12508), .Z(n12505) );
  NOR2_X1 U12519 ( .A1(n7593), .A2(n7787), .ZN(n12508) );
  NAND2_X1 U12520 ( .A1(a_24_), .A2(n12504), .ZN(n12277) );
  NAND2_X1 U12521 ( .A1(n12509), .A2(n12510), .ZN(n12504) );
  NAND2_X1 U12522 ( .A1(n12511), .A2(b_14_), .ZN(n12510) );
  NOR2_X1 U12523 ( .A1(n12512), .A2(n7593), .ZN(n12511) );
  NOR2_X1 U12524 ( .A1(n12230), .A2(n12231), .ZN(n12512) );
  NAND2_X1 U12525 ( .A1(n12230), .A2(n12231), .ZN(n12509) );
  NAND2_X1 U12526 ( .A1(n12513), .A2(n12514), .ZN(n12231) );
  NAND2_X1 U12527 ( .A1(n12515), .A2(b_14_), .ZN(n12514) );
  NOR2_X1 U12528 ( .A1(n12516), .A2(n8052), .ZN(n12515) );
  NOR2_X1 U12529 ( .A1(n12272), .A2(n12274), .ZN(n12516) );
  NAND2_X1 U12530 ( .A1(n12272), .A2(n12274), .ZN(n12513) );
  NAND2_X1 U12531 ( .A1(n12517), .A2(n12518), .ZN(n12274) );
  NAND2_X1 U12532 ( .A1(n12270), .A2(n12519), .ZN(n12518) );
  NAND2_X1 U12533 ( .A1(n12269), .A2(n12268), .ZN(n12519) );
  NOR2_X1 U12534 ( .A1(n8056), .A2(n7563), .ZN(n12270) );
  INV_X1 U12535 ( .A(b_14_), .ZN(n8056) );
  OR2_X1 U12536 ( .A1(n12268), .A2(n12269), .ZN(n12517) );
  AND2_X1 U12537 ( .A1(n12265), .A2(n12520), .ZN(n12269) );
  NAND2_X1 U12538 ( .A1(n12264), .A2(n12266), .ZN(n12520) );
  NAND2_X1 U12539 ( .A1(n12521), .A2(n12522), .ZN(n12266) );
  NAND2_X1 U12540 ( .A1(b_14_), .A2(a_28_), .ZN(n12522) );
  INV_X1 U12541 ( .A(n12523), .ZN(n12521) );
  XOR2_X1 U12542 ( .A(n12524), .B(n12525), .Z(n12264) );
  NOR2_X1 U12543 ( .A1(n7529), .A2(n7787), .ZN(n12525) );
  XOR2_X1 U12544 ( .A(n12526), .B(n12527), .Z(n12524) );
  NAND2_X1 U12545 ( .A1(a_28_), .A2(n12523), .ZN(n12265) );
  NAND2_X1 U12546 ( .A1(n12528), .A2(n12529), .ZN(n12523) );
  NAND2_X1 U12547 ( .A1(n12530), .A2(b_14_), .ZN(n12529) );
  NOR2_X1 U12548 ( .A1(n12531), .A2(n7529), .ZN(n12530) );
  NOR2_X1 U12549 ( .A1(n12250), .A2(n12251), .ZN(n12531) );
  NAND2_X1 U12550 ( .A1(n12250), .A2(n12251), .ZN(n12528) );
  NAND2_X1 U12551 ( .A1(n12532), .A2(n12533), .ZN(n12251) );
  NAND2_X1 U12552 ( .A1(n12534), .A2(b_12_), .ZN(n12533) );
  NOR2_X1 U12553 ( .A1(n12535), .A2(n8048), .ZN(n12534) );
  NOR2_X1 U12554 ( .A1(n8676), .A2(n7787), .ZN(n12535) );
  NAND2_X1 U12555 ( .A1(n12536), .A2(b_13_), .ZN(n12532) );
  NOR2_X1 U12556 ( .A1(n12537), .A2(n7515), .ZN(n12536) );
  NOR2_X1 U12557 ( .A1(n8679), .A2(n8057), .ZN(n12537) );
  AND2_X1 U12558 ( .A1(n12538), .A2(b_14_), .ZN(n12250) );
  NOR2_X1 U12559 ( .A1(n8451), .A2(n7787), .ZN(n12538) );
  XOR2_X1 U12560 ( .A(n12539), .B(n12540), .Z(n12268) );
  NAND2_X1 U12561 ( .A1(n12541), .A2(n12542), .ZN(n12539) );
  XNOR2_X1 U12562 ( .A(n12543), .B(n12544), .ZN(n12272) );
  XNOR2_X1 U12563 ( .A(n12545), .B(n12546), .ZN(n12543) );
  XOR2_X1 U12564 ( .A(n12547), .B(n12548), .Z(n12230) );
  XNOR2_X1 U12565 ( .A(n12549), .B(n12550), .ZN(n12547) );
  NAND2_X1 U12566 ( .A1(b_13_), .A2(a_26_), .ZN(n12549) );
  XNOR2_X1 U12567 ( .A(n12551), .B(n12552), .ZN(n12280) );
  NAND2_X1 U12568 ( .A1(n12553), .A2(n12554), .ZN(n12551) );
  XOR2_X1 U12569 ( .A(n12555), .B(n12556), .Z(n12284) );
  XOR2_X1 U12570 ( .A(n12557), .B(n12558), .Z(n12555) );
  XOR2_X1 U12571 ( .A(n12559), .B(n12560), .Z(n12288) );
  XOR2_X1 U12572 ( .A(n12561), .B(n12562), .Z(n12559) );
  NOR2_X1 U12573 ( .A1(n7645), .A2(n7787), .ZN(n12562) );
  XOR2_X1 U12574 ( .A(n12563), .B(n12564), .Z(n12291) );
  XOR2_X1 U12575 ( .A(n12565), .B(n12566), .Z(n12563) );
  XNOR2_X1 U12576 ( .A(n12567), .B(n12568), .ZN(n12296) );
  XOR2_X1 U12577 ( .A(n12569), .B(n12570), .Z(n12568) );
  NAND2_X1 U12578 ( .A1(b_13_), .A2(a_20_), .ZN(n12570) );
  XOR2_X1 U12579 ( .A(n12571), .B(n12572), .Z(n12300) );
  XOR2_X1 U12580 ( .A(n12573), .B(n12574), .Z(n12571) );
  XNOR2_X1 U12581 ( .A(n12575), .B(n12576), .ZN(n12304) );
  XNOR2_X1 U12582 ( .A(n12577), .B(n12578), .ZN(n12575) );
  XOR2_X1 U12583 ( .A(n12579), .B(n12580), .Z(n12195) );
  XOR2_X1 U12584 ( .A(n12581), .B(n12582), .Z(n12580) );
  NAND2_X1 U12585 ( .A1(b_13_), .A2(a_17_), .ZN(n12582) );
  XOR2_X1 U12586 ( .A(n12583), .B(n12584), .Z(n12308) );
  NAND2_X1 U12587 ( .A1(n12585), .A2(n12586), .ZN(n12583) );
  XOR2_X1 U12588 ( .A(n12587), .B(n12588), .Z(n12134) );
  XOR2_X1 U12589 ( .A(n12589), .B(n12590), .Z(n12588) );
  NAND2_X1 U12590 ( .A1(b_13_), .A2(a_4_), .ZN(n12590) );
  XNOR2_X1 U12591 ( .A(n12591), .B(n12592), .ZN(n12352) );
  XOR2_X1 U12592 ( .A(n12593), .B(n12594), .Z(n12592) );
  NAND2_X1 U12593 ( .A1(b_13_), .A2(a_3_), .ZN(n12594) );
  NOR2_X1 U12594 ( .A1(n12595), .A2(n12116), .ZN(n12359) );
  XOR2_X1 U12595 ( .A(n12596), .B(n12597), .Z(n12116) );
  XNOR2_X1 U12596 ( .A(n12598), .B(n12599), .ZN(n12597) );
  AND2_X1 U12597 ( .A1(n8229), .A2(n8228), .ZN(n12595) );
  NAND2_X1 U12598 ( .A1(n12600), .A2(n8227), .ZN(n8176) );
  NOR2_X1 U12599 ( .A1(n8229), .A2(n8228), .ZN(n8227) );
  AND2_X1 U12600 ( .A1(n12601), .A2(n12602), .ZN(n8228) );
  NAND2_X1 U12601 ( .A1(n12599), .A2(n12603), .ZN(n12602) );
  OR2_X1 U12602 ( .A1(n12598), .A2(n12596), .ZN(n12603) );
  NOR2_X1 U12603 ( .A1(n7787), .A2(n8307), .ZN(n12599) );
  NAND2_X1 U12604 ( .A1(n12596), .A2(n12598), .ZN(n12601) );
  NAND2_X1 U12605 ( .A1(n12604), .A2(n12605), .ZN(n12598) );
  NAND2_X1 U12606 ( .A1(n12606), .A2(b_13_), .ZN(n12605) );
  NOR2_X1 U12607 ( .A1(n12607), .A2(n7973), .ZN(n12606) );
  NOR2_X1 U12608 ( .A1(n12366), .A2(n12367), .ZN(n12607) );
  NAND2_X1 U12609 ( .A1(n12366), .A2(n12367), .ZN(n12604) );
  NAND2_X1 U12610 ( .A1(n12608), .A2(n12609), .ZN(n12367) );
  NAND2_X1 U12611 ( .A1(n12610), .A2(b_13_), .ZN(n12609) );
  NOR2_X1 U12612 ( .A1(n12611), .A2(n7965), .ZN(n12610) );
  NOR2_X1 U12613 ( .A1(n12373), .A2(n12375), .ZN(n12611) );
  NAND2_X1 U12614 ( .A1(n12373), .A2(n12375), .ZN(n12608) );
  NAND2_X1 U12615 ( .A1(n12612), .A2(n12613), .ZN(n12375) );
  NAND2_X1 U12616 ( .A1(n12614), .A2(b_13_), .ZN(n12613) );
  NOR2_X1 U12617 ( .A1(n12615), .A2(n7945), .ZN(n12614) );
  NOR2_X1 U12618 ( .A1(n12591), .A2(n12593), .ZN(n12615) );
  NAND2_X1 U12619 ( .A1(n12591), .A2(n12593), .ZN(n12612) );
  NAND2_X1 U12620 ( .A1(n12616), .A2(n12617), .ZN(n12593) );
  NAND2_X1 U12621 ( .A1(n12618), .A2(b_13_), .ZN(n12617) );
  NOR2_X1 U12622 ( .A1(n12619), .A2(n7934), .ZN(n12618) );
  NOR2_X1 U12623 ( .A1(n12587), .A2(n12589), .ZN(n12619) );
  NAND2_X1 U12624 ( .A1(n12587), .A2(n12589), .ZN(n12616) );
  NAND2_X1 U12625 ( .A1(n12620), .A2(n12621), .ZN(n12589) );
  NAND2_X1 U12626 ( .A1(n12622), .A2(b_13_), .ZN(n12621) );
  NOR2_X1 U12627 ( .A1(n12623), .A2(n7914), .ZN(n12622) );
  NOR2_X1 U12628 ( .A1(n12389), .A2(n12390), .ZN(n12623) );
  NAND2_X1 U12629 ( .A1(n12389), .A2(n12390), .ZN(n12620) );
  NAND2_X1 U12630 ( .A1(n12624), .A2(n12625), .ZN(n12390) );
  NAND2_X1 U12631 ( .A1(n12626), .A2(b_13_), .ZN(n12625) );
  NOR2_X1 U12632 ( .A1(n12627), .A2(n8061), .ZN(n12626) );
  NOR2_X1 U12633 ( .A1(n12396), .A2(n12398), .ZN(n12627) );
  NAND2_X1 U12634 ( .A1(n12396), .A2(n12398), .ZN(n12624) );
  NAND2_X1 U12635 ( .A1(n12628), .A2(n12629), .ZN(n12398) );
  NAND2_X1 U12636 ( .A1(n12630), .A2(b_13_), .ZN(n12629) );
  NOR2_X1 U12637 ( .A1(n12631), .A2(n7884), .ZN(n12630) );
  NOR2_X1 U12638 ( .A1(n12404), .A2(n12406), .ZN(n12631) );
  NAND2_X1 U12639 ( .A1(n12404), .A2(n12406), .ZN(n12628) );
  NAND2_X1 U12640 ( .A1(n12632), .A2(n12633), .ZN(n12406) );
  NAND2_X1 U12641 ( .A1(n12634), .A2(b_13_), .ZN(n12633) );
  NOR2_X1 U12642 ( .A1(n12635), .A2(n8059), .ZN(n12634) );
  NOR2_X1 U12643 ( .A1(n12412), .A2(n12414), .ZN(n12635) );
  NAND2_X1 U12644 ( .A1(n12412), .A2(n12414), .ZN(n12632) );
  NAND2_X1 U12645 ( .A1(n12636), .A2(n12637), .ZN(n12414) );
  NAND2_X1 U12646 ( .A1(n12638), .A2(b_13_), .ZN(n12637) );
  NOR2_X1 U12647 ( .A1(n12639), .A2(n7848), .ZN(n12638) );
  NOR2_X1 U12648 ( .A1(n12420), .A2(n12422), .ZN(n12639) );
  NAND2_X1 U12649 ( .A1(n12420), .A2(n12422), .ZN(n12636) );
  NAND2_X1 U12650 ( .A1(n12640), .A2(n12641), .ZN(n12422) );
  NAND2_X1 U12651 ( .A1(n12642), .A2(b_13_), .ZN(n12641) );
  NOR2_X1 U12652 ( .A1(n12643), .A2(n7837), .ZN(n12642) );
  NOR2_X1 U12653 ( .A1(n12428), .A2(n12430), .ZN(n12643) );
  NAND2_X1 U12654 ( .A1(n12428), .A2(n12430), .ZN(n12640) );
  NAND2_X1 U12655 ( .A1(n12644), .A2(n12645), .ZN(n12430) );
  NAND2_X1 U12656 ( .A1(n12646), .A2(b_13_), .ZN(n12645) );
  NOR2_X1 U12657 ( .A1(n12647), .A2(n7817), .ZN(n12646) );
  NOR2_X1 U12658 ( .A1(n12436), .A2(n12438), .ZN(n12647) );
  NAND2_X1 U12659 ( .A1(n12436), .A2(n12438), .ZN(n12644) );
  NAND2_X1 U12660 ( .A1(n12648), .A2(n12649), .ZN(n12438) );
  NAND2_X1 U12661 ( .A1(n12650), .A2(b_13_), .ZN(n12649) );
  NOR2_X1 U12662 ( .A1(n12651), .A2(n7806), .ZN(n12650) );
  NOR2_X1 U12663 ( .A1(n12445), .A2(n12446), .ZN(n12651) );
  NAND2_X1 U12664 ( .A1(n12445), .A2(n12446), .ZN(n12648) );
  NAND2_X1 U12665 ( .A1(n12652), .A2(n12653), .ZN(n12446) );
  NAND2_X1 U12666 ( .A1(n12453), .A2(n12654), .ZN(n12653) );
  OR2_X1 U12667 ( .A1(n12454), .A2(n7781), .ZN(n12654) );
  XNOR2_X1 U12668 ( .A(n12655), .B(n12656), .ZN(n12453) );
  NAND2_X1 U12669 ( .A1(n12657), .A2(n12658), .ZN(n12655) );
  NAND2_X1 U12670 ( .A1(n7781), .A2(n12454), .ZN(n12652) );
  NAND2_X1 U12671 ( .A1(n12659), .A2(n12660), .ZN(n12454) );
  NAND2_X1 U12672 ( .A1(n12661), .A2(b_13_), .ZN(n12660) );
  NOR2_X1 U12673 ( .A1(n12662), .A2(n7775), .ZN(n12661) );
  NOR2_X1 U12674 ( .A1(n12460), .A2(n12461), .ZN(n12662) );
  NAND2_X1 U12675 ( .A1(n12460), .A2(n12461), .ZN(n12659) );
  NAND2_X1 U12676 ( .A1(n12663), .A2(n12664), .ZN(n12461) );
  NAND2_X1 U12677 ( .A1(n12665), .A2(b_13_), .ZN(n12664) );
  NOR2_X1 U12678 ( .A1(n12666), .A2(n7754), .ZN(n12665) );
  NOR2_X1 U12679 ( .A1(n12467), .A2(n12468), .ZN(n12666) );
  NAND2_X1 U12680 ( .A1(n12467), .A2(n12468), .ZN(n12663) );
  NAND2_X1 U12681 ( .A1(n12585), .A2(n12667), .ZN(n12468) );
  NAND2_X1 U12682 ( .A1(n12584), .A2(n12586), .ZN(n12667) );
  NAND2_X1 U12683 ( .A1(n12668), .A2(n12669), .ZN(n12586) );
  NAND2_X1 U12684 ( .A1(b_13_), .A2(a_16_), .ZN(n12669) );
  INV_X1 U12685 ( .A(n12670), .ZN(n12668) );
  XNOR2_X1 U12686 ( .A(n12671), .B(n12672), .ZN(n12584) );
  XNOR2_X1 U12687 ( .A(n12673), .B(n12674), .ZN(n12672) );
  NAND2_X1 U12688 ( .A1(a_16_), .A2(n12670), .ZN(n12585) );
  NAND2_X1 U12689 ( .A1(n12675), .A2(n12676), .ZN(n12670) );
  NAND2_X1 U12690 ( .A1(n12677), .A2(b_13_), .ZN(n12676) );
  NOR2_X1 U12691 ( .A1(n12678), .A2(n7723), .ZN(n12677) );
  NOR2_X1 U12692 ( .A1(n12579), .A2(n12581), .ZN(n12678) );
  NAND2_X1 U12693 ( .A1(n12579), .A2(n12581), .ZN(n12675) );
  NAND2_X1 U12694 ( .A1(n12679), .A2(n12680), .ZN(n12581) );
  NAND2_X1 U12695 ( .A1(n12578), .A2(n12681), .ZN(n12680) );
  NAND2_X1 U12696 ( .A1(n12577), .A2(n12576), .ZN(n12681) );
  NOR2_X1 U12697 ( .A1(n7787), .A2(n7707), .ZN(n12578) );
  OR2_X1 U12698 ( .A1(n12576), .A2(n12577), .ZN(n12679) );
  AND2_X1 U12699 ( .A1(n12682), .A2(n12683), .ZN(n12577) );
  NAND2_X1 U12700 ( .A1(n12574), .A2(n12684), .ZN(n12683) );
  OR2_X1 U12701 ( .A1(n12573), .A2(n12572), .ZN(n12684) );
  NOR2_X1 U12702 ( .A1(n7787), .A2(n7687), .ZN(n12574) );
  NAND2_X1 U12703 ( .A1(n12572), .A2(n12573), .ZN(n12682) );
  NAND2_X1 U12704 ( .A1(n12685), .A2(n12686), .ZN(n12573) );
  NAND2_X1 U12705 ( .A1(n12687), .A2(b_13_), .ZN(n12686) );
  NOR2_X1 U12706 ( .A1(n12688), .A2(n7676), .ZN(n12687) );
  NOR2_X1 U12707 ( .A1(n12567), .A2(n12569), .ZN(n12688) );
  NAND2_X1 U12708 ( .A1(n12567), .A2(n12569), .ZN(n12685) );
  NAND2_X1 U12709 ( .A1(n12689), .A2(n12690), .ZN(n12569) );
  NAND2_X1 U12710 ( .A1(n12566), .A2(n12691), .ZN(n12690) );
  OR2_X1 U12711 ( .A1(n12565), .A2(n12564), .ZN(n12691) );
  NOR2_X1 U12712 ( .A1(n7787), .A2(n7656), .ZN(n12566) );
  NAND2_X1 U12713 ( .A1(n12564), .A2(n12565), .ZN(n12689) );
  NAND2_X1 U12714 ( .A1(n12692), .A2(n12693), .ZN(n12565) );
  NAND2_X1 U12715 ( .A1(n12694), .A2(b_13_), .ZN(n12693) );
  NOR2_X1 U12716 ( .A1(n12695), .A2(n7645), .ZN(n12694) );
  NOR2_X1 U12717 ( .A1(n12560), .A2(n12561), .ZN(n12695) );
  NAND2_X1 U12718 ( .A1(n12560), .A2(n12561), .ZN(n12692) );
  NAND2_X1 U12719 ( .A1(n12696), .A2(n12697), .ZN(n12561) );
  NAND2_X1 U12720 ( .A1(n12558), .A2(n12698), .ZN(n12697) );
  OR2_X1 U12721 ( .A1(n12557), .A2(n12556), .ZN(n12698) );
  NOR2_X1 U12722 ( .A1(n7787), .A2(n7624), .ZN(n12558) );
  NAND2_X1 U12723 ( .A1(n12556), .A2(n12557), .ZN(n12696) );
  NAND2_X1 U12724 ( .A1(n12553), .A2(n12699), .ZN(n12557) );
  NAND2_X1 U12725 ( .A1(n12552), .A2(n12554), .ZN(n12699) );
  NAND2_X1 U12726 ( .A1(n12700), .A2(n12701), .ZN(n12554) );
  NAND2_X1 U12727 ( .A1(b_13_), .A2(a_24_), .ZN(n12701) );
  INV_X1 U12728 ( .A(n12702), .ZN(n12700) );
  XOR2_X1 U12729 ( .A(n12703), .B(n12704), .Z(n12552) );
  XOR2_X1 U12730 ( .A(n12705), .B(n12706), .Z(n12703) );
  NOR2_X1 U12731 ( .A1(n7593), .A2(n8057), .ZN(n12706) );
  NAND2_X1 U12732 ( .A1(a_24_), .A2(n12702), .ZN(n12553) );
  NAND2_X1 U12733 ( .A1(n12707), .A2(n12708), .ZN(n12702) );
  NAND2_X1 U12734 ( .A1(n12709), .A2(b_13_), .ZN(n12708) );
  NOR2_X1 U12735 ( .A1(n12710), .A2(n7593), .ZN(n12709) );
  NOR2_X1 U12736 ( .A1(n12506), .A2(n12507), .ZN(n12710) );
  NAND2_X1 U12737 ( .A1(n12506), .A2(n12507), .ZN(n12707) );
  NAND2_X1 U12738 ( .A1(n12711), .A2(n12712), .ZN(n12507) );
  NAND2_X1 U12739 ( .A1(n12713), .A2(b_13_), .ZN(n12712) );
  NOR2_X1 U12740 ( .A1(n12714), .A2(n8052), .ZN(n12713) );
  NOR2_X1 U12741 ( .A1(n12548), .A2(n12550), .ZN(n12714) );
  NAND2_X1 U12742 ( .A1(n12548), .A2(n12550), .ZN(n12711) );
  NAND2_X1 U12743 ( .A1(n12715), .A2(n12716), .ZN(n12550) );
  NAND2_X1 U12744 ( .A1(n12546), .A2(n12717), .ZN(n12716) );
  NAND2_X1 U12745 ( .A1(n12545), .A2(n12544), .ZN(n12717) );
  NOR2_X1 U12746 ( .A1(n7787), .A2(n7563), .ZN(n12546) );
  INV_X1 U12747 ( .A(b_13_), .ZN(n7787) );
  OR2_X1 U12748 ( .A1(n12544), .A2(n12545), .ZN(n12715) );
  AND2_X1 U12749 ( .A1(n12541), .A2(n12718), .ZN(n12545) );
  NAND2_X1 U12750 ( .A1(n12540), .A2(n12542), .ZN(n12718) );
  NAND2_X1 U12751 ( .A1(n12719), .A2(n12720), .ZN(n12542) );
  NAND2_X1 U12752 ( .A1(b_13_), .A2(a_28_), .ZN(n12720) );
  INV_X1 U12753 ( .A(n12721), .ZN(n12719) );
  XOR2_X1 U12754 ( .A(n12722), .B(n12723), .Z(n12540) );
  NOR2_X1 U12755 ( .A1(n7529), .A2(n8057), .ZN(n12723) );
  XOR2_X1 U12756 ( .A(n12724), .B(n12725), .Z(n12722) );
  NAND2_X1 U12757 ( .A1(a_28_), .A2(n12721), .ZN(n12541) );
  NAND2_X1 U12758 ( .A1(n12726), .A2(n12727), .ZN(n12721) );
  NAND2_X1 U12759 ( .A1(n12728), .A2(b_13_), .ZN(n12727) );
  NOR2_X1 U12760 ( .A1(n12729), .A2(n7529), .ZN(n12728) );
  NOR2_X1 U12761 ( .A1(n12526), .A2(n12527), .ZN(n12729) );
  NAND2_X1 U12762 ( .A1(n12526), .A2(n12527), .ZN(n12726) );
  NAND2_X1 U12763 ( .A1(n12730), .A2(n12731), .ZN(n12527) );
  NAND2_X1 U12764 ( .A1(n12732), .A2(a_31_), .ZN(n12731) );
  NOR2_X1 U12765 ( .A1(n12733), .A2(n7818), .ZN(n12732) );
  NOR2_X1 U12766 ( .A1(n8676), .A2(n8057), .ZN(n12733) );
  NAND2_X1 U12767 ( .A1(n12734), .A2(b_12_), .ZN(n12730) );
  NOR2_X1 U12768 ( .A1(n12735), .A2(n7515), .ZN(n12734) );
  NOR2_X1 U12769 ( .A1(n8679), .A2(n7818), .ZN(n12735) );
  AND2_X1 U12770 ( .A1(n12736), .A2(b_13_), .ZN(n12526) );
  NOR2_X1 U12771 ( .A1(n8451), .A2(n8057), .ZN(n12736) );
  XOR2_X1 U12772 ( .A(n12737), .B(n12738), .Z(n12544) );
  NAND2_X1 U12773 ( .A1(n12739), .A2(n12740), .ZN(n12737) );
  XNOR2_X1 U12774 ( .A(n12741), .B(n12742), .ZN(n12548) );
  XNOR2_X1 U12775 ( .A(n12743), .B(n12744), .ZN(n12741) );
  XOR2_X1 U12776 ( .A(n12745), .B(n12746), .Z(n12506) );
  XNOR2_X1 U12777 ( .A(n12747), .B(n12748), .ZN(n12745) );
  NAND2_X1 U12778 ( .A1(b_12_), .A2(a_26_), .ZN(n12747) );
  XNOR2_X1 U12779 ( .A(n12749), .B(n12750), .ZN(n12556) );
  NAND2_X1 U12780 ( .A1(n12751), .A2(n12752), .ZN(n12749) );
  XOR2_X1 U12781 ( .A(n12753), .B(n12754), .Z(n12560) );
  XOR2_X1 U12782 ( .A(n12755), .B(n12756), .Z(n12753) );
  XOR2_X1 U12783 ( .A(n12757), .B(n12758), .Z(n12564) );
  XOR2_X1 U12784 ( .A(n12759), .B(n12760), .Z(n12757) );
  NOR2_X1 U12785 ( .A1(n7645), .A2(n8057), .ZN(n12760) );
  XOR2_X1 U12786 ( .A(n12761), .B(n12762), .Z(n12567) );
  XOR2_X1 U12787 ( .A(n12763), .B(n12764), .Z(n12761) );
  XNOR2_X1 U12788 ( .A(n12765), .B(n12766), .ZN(n12572) );
  XOR2_X1 U12789 ( .A(n12767), .B(n12768), .Z(n12766) );
  NAND2_X1 U12790 ( .A1(b_12_), .A2(a_20_), .ZN(n12768) );
  XNOR2_X1 U12791 ( .A(n12769), .B(n12770), .ZN(n12576) );
  XOR2_X1 U12792 ( .A(n12771), .B(n12772), .Z(n12769) );
  NOR2_X1 U12793 ( .A1(n7687), .A2(n8057), .ZN(n12772) );
  XNOR2_X1 U12794 ( .A(n12773), .B(n12774), .ZN(n12579) );
  XNOR2_X1 U12795 ( .A(n12775), .B(n12776), .ZN(n12773) );
  XNOR2_X1 U12796 ( .A(n12777), .B(n12778), .ZN(n12467) );
  XNOR2_X1 U12797 ( .A(n12779), .B(n12780), .ZN(n12778) );
  XNOR2_X1 U12798 ( .A(n12781), .B(n12782), .ZN(n12460) );
  XOR2_X1 U12799 ( .A(n12783), .B(n12784), .Z(n12782) );
  NAND2_X1 U12800 ( .A1(b_12_), .A2(a_15_), .ZN(n12784) );
  INV_X1 U12801 ( .A(n8011), .ZN(n7781) );
  NAND2_X1 U12802 ( .A1(b_13_), .A2(a_13_), .ZN(n8011) );
  XNOR2_X1 U12803 ( .A(n12785), .B(n12786), .ZN(n12445) );
  NAND2_X1 U12804 ( .A1(n12787), .A2(n12788), .ZN(n12785) );
  XOR2_X1 U12805 ( .A(n12789), .B(n12790), .Z(n12436) );
  XOR2_X1 U12806 ( .A(n12791), .B(n12792), .Z(n12789) );
  XNOR2_X1 U12807 ( .A(n12793), .B(n12794), .ZN(n12428) );
  NAND2_X1 U12808 ( .A1(n12795), .A2(n12796), .ZN(n12793) );
  XNOR2_X1 U12809 ( .A(n12797), .B(n12798), .ZN(n12420) );
  NAND2_X1 U12810 ( .A1(n12799), .A2(n12800), .ZN(n12797) );
  XNOR2_X1 U12811 ( .A(n12801), .B(n12802), .ZN(n12412) );
  NAND2_X1 U12812 ( .A1(n12803), .A2(n12804), .ZN(n12801) );
  XNOR2_X1 U12813 ( .A(n12805), .B(n12806), .ZN(n12404) );
  XNOR2_X1 U12814 ( .A(n12807), .B(n12808), .ZN(n12805) );
  XOR2_X1 U12815 ( .A(n12809), .B(n12810), .Z(n12396) );
  XOR2_X1 U12816 ( .A(n12811), .B(n12812), .Z(n12809) );
  NOR2_X1 U12817 ( .A1(n7884), .A2(n8057), .ZN(n12812) );
  XNOR2_X1 U12818 ( .A(n12813), .B(n12814), .ZN(n12389) );
  NAND2_X1 U12819 ( .A1(n12815), .A2(n12816), .ZN(n12813) );
  XNOR2_X1 U12820 ( .A(n12817), .B(n12818), .ZN(n12587) );
  NAND2_X1 U12821 ( .A1(n12819), .A2(n12820), .ZN(n12817) );
  XOR2_X1 U12822 ( .A(n12821), .B(n12822), .Z(n12591) );
  NOR2_X1 U12823 ( .A1(n12823), .A2(n12824), .ZN(n12822) );
  NOR2_X1 U12824 ( .A1(n12825), .A2(n12826), .ZN(n12823) );
  NOR2_X1 U12825 ( .A1(n7934), .A2(n8057), .ZN(n12825) );
  XOR2_X1 U12826 ( .A(n12827), .B(n12828), .Z(n12373) );
  XOR2_X1 U12827 ( .A(n12829), .B(n12830), .Z(n12828) );
  XNOR2_X1 U12828 ( .A(n12831), .B(n12832), .ZN(n12366) );
  XNOR2_X1 U12829 ( .A(n12833), .B(n12834), .ZN(n12832) );
  XNOR2_X1 U12830 ( .A(n12835), .B(n12836), .ZN(n12596) );
  XNOR2_X1 U12831 ( .A(n12837), .B(n12838), .ZN(n12836) );
  XOR2_X1 U12832 ( .A(n12839), .B(n12840), .Z(n8229) );
  XOR2_X1 U12833 ( .A(n12841), .B(n12842), .Z(n12840) );
  NAND2_X1 U12834 ( .A1(b_12_), .A2(a_0_), .ZN(n12842) );
  XOR2_X1 U12835 ( .A(n8217), .B(n8218), .Z(n12600) );
  NAND2_X1 U12836 ( .A1(n12843), .A2(n12844), .ZN(n8181) );
  NOR2_X1 U12837 ( .A1(n8214), .A2(n8218), .ZN(n12844) );
  INV_X1 U12838 ( .A(n8222), .ZN(n8218) );
  NAND2_X1 U12839 ( .A1(n12845), .A2(n12846), .ZN(n8222) );
  NAND2_X1 U12840 ( .A1(n12847), .A2(b_12_), .ZN(n12846) );
  NOR2_X1 U12841 ( .A1(n12848), .A2(n8307), .ZN(n12847) );
  NOR2_X1 U12842 ( .A1(n12839), .A2(n12841), .ZN(n12848) );
  NAND2_X1 U12843 ( .A1(n12839), .A2(n12841), .ZN(n12845) );
  NAND2_X1 U12844 ( .A1(n12849), .A2(n12850), .ZN(n12841) );
  NAND2_X1 U12845 ( .A1(n12838), .A2(n12851), .ZN(n12850) );
  OR2_X1 U12846 ( .A1(n12837), .A2(n12835), .ZN(n12851) );
  NOR2_X1 U12847 ( .A1(n8057), .A2(n7973), .ZN(n12838) );
  NAND2_X1 U12848 ( .A1(n12835), .A2(n12837), .ZN(n12849) );
  NAND2_X1 U12849 ( .A1(n12852), .A2(n12853), .ZN(n12837) );
  NAND2_X1 U12850 ( .A1(n12834), .A2(n12854), .ZN(n12853) );
  OR2_X1 U12851 ( .A1(n12833), .A2(n12831), .ZN(n12854) );
  NOR2_X1 U12852 ( .A1(n8057), .A2(n7965), .ZN(n12834) );
  NAND2_X1 U12853 ( .A1(n12831), .A2(n12833), .ZN(n12852) );
  NAND2_X1 U12854 ( .A1(n12855), .A2(n12856), .ZN(n12833) );
  NAND2_X1 U12855 ( .A1(n12830), .A2(n12857), .ZN(n12856) );
  NAND2_X1 U12856 ( .A1(n12829), .A2(n12827), .ZN(n12857) );
  NOR2_X1 U12857 ( .A1(n8057), .A2(n7945), .ZN(n12830) );
  OR2_X1 U12858 ( .A1(n12827), .A2(n12829), .ZN(n12855) );
  NOR2_X1 U12859 ( .A1(n12824), .A2(n12858), .ZN(n12829) );
  AND2_X1 U12860 ( .A1(n12821), .A2(n12859), .ZN(n12858) );
  NAND2_X1 U12861 ( .A1(n12860), .A2(n12861), .ZN(n12859) );
  NAND2_X1 U12862 ( .A1(b_12_), .A2(a_4_), .ZN(n12861) );
  XOR2_X1 U12863 ( .A(n12862), .B(n12863), .Z(n12821) );
  XOR2_X1 U12864 ( .A(n12864), .B(n12865), .Z(n12862) );
  NOR2_X1 U12865 ( .A1(n7818), .A2(n7914), .ZN(n12865) );
  NOR2_X1 U12866 ( .A1(n7934), .A2(n12860), .ZN(n12824) );
  INV_X1 U12867 ( .A(n12826), .ZN(n12860) );
  NAND2_X1 U12868 ( .A1(n12819), .A2(n12866), .ZN(n12826) );
  NAND2_X1 U12869 ( .A1(n12818), .A2(n12820), .ZN(n12866) );
  NAND2_X1 U12870 ( .A1(n12867), .A2(n12868), .ZN(n12820) );
  NAND2_X1 U12871 ( .A1(b_12_), .A2(a_5_), .ZN(n12868) );
  INV_X1 U12872 ( .A(n12869), .ZN(n12867) );
  XOR2_X1 U12873 ( .A(n12870), .B(n12871), .Z(n12818) );
  XOR2_X1 U12874 ( .A(n12872), .B(n12873), .Z(n12870) );
  NOR2_X1 U12875 ( .A1(n7818), .A2(n8061), .ZN(n12873) );
  NAND2_X1 U12876 ( .A1(a_5_), .A2(n12869), .ZN(n12819) );
  NAND2_X1 U12877 ( .A1(n12815), .A2(n12874), .ZN(n12869) );
  NAND2_X1 U12878 ( .A1(n12814), .A2(n12816), .ZN(n12874) );
  NAND2_X1 U12879 ( .A1(n12875), .A2(n12876), .ZN(n12816) );
  NAND2_X1 U12880 ( .A1(b_12_), .A2(a_6_), .ZN(n12876) );
  INV_X1 U12881 ( .A(n12877), .ZN(n12875) );
  XOR2_X1 U12882 ( .A(n12878), .B(n12879), .Z(n12814) );
  XOR2_X1 U12883 ( .A(n12880), .B(n12881), .Z(n12878) );
  NOR2_X1 U12884 ( .A1(n7818), .A2(n7884), .ZN(n12881) );
  NAND2_X1 U12885 ( .A1(a_6_), .A2(n12877), .ZN(n12815) );
  NAND2_X1 U12886 ( .A1(n12882), .A2(n12883), .ZN(n12877) );
  NAND2_X1 U12887 ( .A1(n12884), .A2(b_12_), .ZN(n12883) );
  NOR2_X1 U12888 ( .A1(n12885), .A2(n7884), .ZN(n12884) );
  NOR2_X1 U12889 ( .A1(n12810), .A2(n12811), .ZN(n12885) );
  NAND2_X1 U12890 ( .A1(n12810), .A2(n12811), .ZN(n12882) );
  NAND2_X1 U12891 ( .A1(n12886), .A2(n12887), .ZN(n12811) );
  NAND2_X1 U12892 ( .A1(n12808), .A2(n12888), .ZN(n12887) );
  NAND2_X1 U12893 ( .A1(n12807), .A2(n12806), .ZN(n12888) );
  NOR2_X1 U12894 ( .A1(n8057), .A2(n8059), .ZN(n12808) );
  OR2_X1 U12895 ( .A1(n12806), .A2(n12807), .ZN(n12886) );
  AND2_X1 U12896 ( .A1(n12803), .A2(n12889), .ZN(n12807) );
  NAND2_X1 U12897 ( .A1(n12802), .A2(n12804), .ZN(n12889) );
  NAND2_X1 U12898 ( .A1(n12890), .A2(n12891), .ZN(n12804) );
  NAND2_X1 U12899 ( .A1(b_12_), .A2(a_9_), .ZN(n12891) );
  INV_X1 U12900 ( .A(n12892), .ZN(n12890) );
  XOR2_X1 U12901 ( .A(n12893), .B(n12894), .Z(n12802) );
  XNOR2_X1 U12902 ( .A(n12895), .B(n12896), .ZN(n12893) );
  NAND2_X1 U12903 ( .A1(a_10_), .A2(b_11_), .ZN(n12895) );
  NAND2_X1 U12904 ( .A1(a_9_), .A2(n12892), .ZN(n12803) );
  NAND2_X1 U12905 ( .A1(n12799), .A2(n12897), .ZN(n12892) );
  NAND2_X1 U12906 ( .A1(n12798), .A2(n12800), .ZN(n12897) );
  NAND2_X1 U12907 ( .A1(n12898), .A2(n12899), .ZN(n12800) );
  NAND2_X1 U12908 ( .A1(b_12_), .A2(a_10_), .ZN(n12899) );
  INV_X1 U12909 ( .A(n12900), .ZN(n12898) );
  XNOR2_X1 U12910 ( .A(n12901), .B(n12902), .ZN(n12798) );
  XNOR2_X1 U12911 ( .A(n7812), .B(n12903), .ZN(n12902) );
  NAND2_X1 U12912 ( .A1(a_10_), .A2(n12900), .ZN(n12799) );
  NAND2_X1 U12913 ( .A1(n12795), .A2(n12904), .ZN(n12900) );
  NAND2_X1 U12914 ( .A1(n12794), .A2(n12796), .ZN(n12904) );
  NAND2_X1 U12915 ( .A1(n12905), .A2(n12906), .ZN(n12796) );
  NAND2_X1 U12916 ( .A1(b_12_), .A2(a_11_), .ZN(n12906) );
  INV_X1 U12917 ( .A(n12907), .ZN(n12905) );
  XNOR2_X1 U12918 ( .A(n12908), .B(n12909), .ZN(n12794) );
  XOR2_X1 U12919 ( .A(n12910), .B(n12911), .Z(n12909) );
  NAND2_X1 U12920 ( .A1(a_12_), .A2(b_11_), .ZN(n12911) );
  NAND2_X1 U12921 ( .A1(a_11_), .A2(n12907), .ZN(n12795) );
  NAND2_X1 U12922 ( .A1(n12912), .A2(n12913), .ZN(n12907) );
  NAND2_X1 U12923 ( .A1(n12790), .A2(n12914), .ZN(n12913) );
  OR2_X1 U12924 ( .A1(n12791), .A2(n12792), .ZN(n12914) );
  XOR2_X1 U12925 ( .A(n12915), .B(n12916), .Z(n12790) );
  XOR2_X1 U12926 ( .A(n12917), .B(n12918), .Z(n12915) );
  NOR2_X1 U12927 ( .A1(n7818), .A2(n7786), .ZN(n12918) );
  NAND2_X1 U12928 ( .A1(n12792), .A2(n12791), .ZN(n12912) );
  NAND2_X1 U12929 ( .A1(n12787), .A2(n12919), .ZN(n12791) );
  NAND2_X1 U12930 ( .A1(n12786), .A2(n12788), .ZN(n12919) );
  NAND2_X1 U12931 ( .A1(n12920), .A2(n12921), .ZN(n12788) );
  NAND2_X1 U12932 ( .A1(b_12_), .A2(a_13_), .ZN(n12921) );
  INV_X1 U12933 ( .A(n12922), .ZN(n12920) );
  XOR2_X1 U12934 ( .A(n12923), .B(n12924), .Z(n12786) );
  XOR2_X1 U12935 ( .A(n12925), .B(n12926), .Z(n12923) );
  NOR2_X1 U12936 ( .A1(n7818), .A2(n7775), .ZN(n12926) );
  NAND2_X1 U12937 ( .A1(a_13_), .A2(n12922), .ZN(n12787) );
  NAND2_X1 U12938 ( .A1(n12657), .A2(n12927), .ZN(n12922) );
  NAND2_X1 U12939 ( .A1(n12656), .A2(n12658), .ZN(n12927) );
  NAND2_X1 U12940 ( .A1(n12928), .A2(n12929), .ZN(n12658) );
  NAND2_X1 U12941 ( .A1(b_12_), .A2(a_14_), .ZN(n12929) );
  INV_X1 U12942 ( .A(n12930), .ZN(n12928) );
  XOR2_X1 U12943 ( .A(n12931), .B(n12932), .Z(n12656) );
  XOR2_X1 U12944 ( .A(n12933), .B(n12934), .Z(n12931) );
  NOR2_X1 U12945 ( .A1(n7818), .A2(n7754), .ZN(n12934) );
  NAND2_X1 U12946 ( .A1(a_14_), .A2(n12930), .ZN(n12657) );
  NAND2_X1 U12947 ( .A1(n12935), .A2(n12936), .ZN(n12930) );
  NAND2_X1 U12948 ( .A1(n12937), .A2(b_12_), .ZN(n12936) );
  NOR2_X1 U12949 ( .A1(n12938), .A2(n7754), .ZN(n12937) );
  NOR2_X1 U12950 ( .A1(n12781), .A2(n12783), .ZN(n12938) );
  NAND2_X1 U12951 ( .A1(n12781), .A2(n12783), .ZN(n12935) );
  NAND2_X1 U12952 ( .A1(n12939), .A2(n12940), .ZN(n12783) );
  NAND2_X1 U12953 ( .A1(n12780), .A2(n12941), .ZN(n12940) );
  OR2_X1 U12954 ( .A1(n12779), .A2(n12777), .ZN(n12941) );
  NOR2_X1 U12955 ( .A1(n8057), .A2(n7743), .ZN(n12780) );
  NAND2_X1 U12956 ( .A1(n12777), .A2(n12779), .ZN(n12939) );
  NAND2_X1 U12957 ( .A1(n12942), .A2(n12943), .ZN(n12779) );
  NAND2_X1 U12958 ( .A1(n12674), .A2(n12944), .ZN(n12943) );
  OR2_X1 U12959 ( .A1(n12673), .A2(n12671), .ZN(n12944) );
  NOR2_X1 U12960 ( .A1(n8057), .A2(n7723), .ZN(n12674) );
  NAND2_X1 U12961 ( .A1(n12671), .A2(n12673), .ZN(n12942) );
  NAND2_X1 U12962 ( .A1(n12945), .A2(n12946), .ZN(n12673) );
  NAND2_X1 U12963 ( .A1(n12776), .A2(n12947), .ZN(n12946) );
  NAND2_X1 U12964 ( .A1(n12775), .A2(n12774), .ZN(n12947) );
  NOR2_X1 U12965 ( .A1(n8057), .A2(n7707), .ZN(n12776) );
  OR2_X1 U12966 ( .A1(n12774), .A2(n12775), .ZN(n12945) );
  AND2_X1 U12967 ( .A1(n12948), .A2(n12949), .ZN(n12775) );
  NAND2_X1 U12968 ( .A1(n12950), .A2(b_12_), .ZN(n12949) );
  NOR2_X1 U12969 ( .A1(n12951), .A2(n7687), .ZN(n12950) );
  NOR2_X1 U12970 ( .A1(n12770), .A2(n12771), .ZN(n12951) );
  NAND2_X1 U12971 ( .A1(n12770), .A2(n12771), .ZN(n12948) );
  NAND2_X1 U12972 ( .A1(n12952), .A2(n12953), .ZN(n12771) );
  NAND2_X1 U12973 ( .A1(n12954), .A2(b_12_), .ZN(n12953) );
  NOR2_X1 U12974 ( .A1(n12955), .A2(n7676), .ZN(n12954) );
  NOR2_X1 U12975 ( .A1(n12765), .A2(n12767), .ZN(n12955) );
  NAND2_X1 U12976 ( .A1(n12765), .A2(n12767), .ZN(n12952) );
  NAND2_X1 U12977 ( .A1(n12956), .A2(n12957), .ZN(n12767) );
  NAND2_X1 U12978 ( .A1(n12764), .A2(n12958), .ZN(n12957) );
  OR2_X1 U12979 ( .A1(n12763), .A2(n12762), .ZN(n12958) );
  NOR2_X1 U12980 ( .A1(n8057), .A2(n7656), .ZN(n12764) );
  NAND2_X1 U12981 ( .A1(n12762), .A2(n12763), .ZN(n12956) );
  NAND2_X1 U12982 ( .A1(n12959), .A2(n12960), .ZN(n12763) );
  NAND2_X1 U12983 ( .A1(n12961), .A2(b_12_), .ZN(n12960) );
  NOR2_X1 U12984 ( .A1(n12962), .A2(n7645), .ZN(n12961) );
  NOR2_X1 U12985 ( .A1(n12758), .A2(n12759), .ZN(n12962) );
  NAND2_X1 U12986 ( .A1(n12758), .A2(n12759), .ZN(n12959) );
  NAND2_X1 U12987 ( .A1(n12963), .A2(n12964), .ZN(n12759) );
  NAND2_X1 U12988 ( .A1(n12756), .A2(n12965), .ZN(n12964) );
  OR2_X1 U12989 ( .A1(n12755), .A2(n12754), .ZN(n12965) );
  NOR2_X1 U12990 ( .A1(n8057), .A2(n7624), .ZN(n12756) );
  NAND2_X1 U12991 ( .A1(n12754), .A2(n12755), .ZN(n12963) );
  NAND2_X1 U12992 ( .A1(n12751), .A2(n12966), .ZN(n12755) );
  NAND2_X1 U12993 ( .A1(n12750), .A2(n12752), .ZN(n12966) );
  NAND2_X1 U12994 ( .A1(n12967), .A2(n12968), .ZN(n12752) );
  NAND2_X1 U12995 ( .A1(b_12_), .A2(a_24_), .ZN(n12968) );
  INV_X1 U12996 ( .A(n12969), .ZN(n12967) );
  XOR2_X1 U12997 ( .A(n12970), .B(n12971), .Z(n12750) );
  XOR2_X1 U12998 ( .A(n12972), .B(n12973), .Z(n12970) );
  NOR2_X1 U12999 ( .A1(n7818), .A2(n7593), .ZN(n12973) );
  NAND2_X1 U13000 ( .A1(a_24_), .A2(n12969), .ZN(n12751) );
  NAND2_X1 U13001 ( .A1(n12974), .A2(n12975), .ZN(n12969) );
  NAND2_X1 U13002 ( .A1(n12976), .A2(b_12_), .ZN(n12975) );
  NOR2_X1 U13003 ( .A1(n12977), .A2(n7593), .ZN(n12976) );
  NOR2_X1 U13004 ( .A1(n12704), .A2(n12705), .ZN(n12977) );
  NAND2_X1 U13005 ( .A1(n12704), .A2(n12705), .ZN(n12974) );
  NAND2_X1 U13006 ( .A1(n12978), .A2(n12979), .ZN(n12705) );
  NAND2_X1 U13007 ( .A1(n12980), .A2(b_12_), .ZN(n12979) );
  NOR2_X1 U13008 ( .A1(n12981), .A2(n8052), .ZN(n12980) );
  NOR2_X1 U13009 ( .A1(n12746), .A2(n12748), .ZN(n12981) );
  NAND2_X1 U13010 ( .A1(n12746), .A2(n12748), .ZN(n12978) );
  NAND2_X1 U13011 ( .A1(n12982), .A2(n12983), .ZN(n12748) );
  NAND2_X1 U13012 ( .A1(n12744), .A2(n12984), .ZN(n12983) );
  NAND2_X1 U13013 ( .A1(n12743), .A2(n12742), .ZN(n12984) );
  NOR2_X1 U13014 ( .A1(n8057), .A2(n7563), .ZN(n12744) );
  INV_X1 U13015 ( .A(b_12_), .ZN(n8057) );
  OR2_X1 U13016 ( .A1(n12742), .A2(n12743), .ZN(n12982) );
  AND2_X1 U13017 ( .A1(n12739), .A2(n12985), .ZN(n12743) );
  NAND2_X1 U13018 ( .A1(n12738), .A2(n12740), .ZN(n12985) );
  NAND2_X1 U13019 ( .A1(n12986), .A2(n12987), .ZN(n12740) );
  NAND2_X1 U13020 ( .A1(b_12_), .A2(a_28_), .ZN(n12987) );
  INV_X1 U13021 ( .A(n12988), .ZN(n12986) );
  XOR2_X1 U13022 ( .A(n12989), .B(n12990), .Z(n12738) );
  NOR2_X1 U13023 ( .A1(n7818), .A2(n7529), .ZN(n12990) );
  XOR2_X1 U13024 ( .A(n12991), .B(n12992), .Z(n12989) );
  NAND2_X1 U13025 ( .A1(a_28_), .A2(n12988), .ZN(n12739) );
  NAND2_X1 U13026 ( .A1(n12993), .A2(n12994), .ZN(n12988) );
  NAND2_X1 U13027 ( .A1(n12995), .A2(b_12_), .ZN(n12994) );
  NOR2_X1 U13028 ( .A1(n12996), .A2(n7529), .ZN(n12995) );
  NOR2_X1 U13029 ( .A1(n12724), .A2(n12725), .ZN(n12996) );
  NAND2_X1 U13030 ( .A1(n12724), .A2(n12725), .ZN(n12993) );
  NAND2_X1 U13031 ( .A1(n12997), .A2(n12998), .ZN(n12725) );
  NAND2_X1 U13032 ( .A1(n12999), .A2(a_31_), .ZN(n12998) );
  NOR2_X1 U13033 ( .A1(n13000), .A2(n13001), .ZN(n12999) );
  NOR2_X1 U13034 ( .A1(n8676), .A2(n7818), .ZN(n13000) );
  NAND2_X1 U13035 ( .A1(n13002), .A2(a_30_), .ZN(n12997) );
  NOR2_X1 U13036 ( .A1(n13003), .A2(n7818), .ZN(n13002) );
  NOR2_X1 U13037 ( .A1(n8679), .A2(n13001), .ZN(n13003) );
  AND2_X1 U13038 ( .A1(n13004), .A2(b_12_), .ZN(n12724) );
  NOR2_X1 U13039 ( .A1(n7818), .A2(n8451), .ZN(n13004) );
  XOR2_X1 U13040 ( .A(n13005), .B(n13006), .Z(n12742) );
  NAND2_X1 U13041 ( .A1(n13007), .A2(n13008), .ZN(n13005) );
  XNOR2_X1 U13042 ( .A(n13009), .B(n13010), .ZN(n12746) );
  XNOR2_X1 U13043 ( .A(n13011), .B(n13012), .ZN(n13009) );
  XOR2_X1 U13044 ( .A(n13013), .B(n13014), .Z(n12704) );
  XNOR2_X1 U13045 ( .A(n13015), .B(n13016), .ZN(n13013) );
  NAND2_X1 U13046 ( .A1(a_26_), .A2(b_11_), .ZN(n13015) );
  XNOR2_X1 U13047 ( .A(n13017), .B(n13018), .ZN(n12754) );
  NAND2_X1 U13048 ( .A1(n13019), .A2(n13020), .ZN(n13017) );
  XOR2_X1 U13049 ( .A(n13021), .B(n13022), .Z(n12758) );
  XOR2_X1 U13050 ( .A(n13023), .B(n13024), .Z(n13021) );
  XOR2_X1 U13051 ( .A(n13025), .B(n13026), .Z(n12762) );
  XOR2_X1 U13052 ( .A(n13027), .B(n13028), .Z(n13025) );
  NOR2_X1 U13053 ( .A1(n7818), .A2(n7645), .ZN(n13028) );
  XOR2_X1 U13054 ( .A(n13029), .B(n13030), .Z(n12765) );
  XOR2_X1 U13055 ( .A(n13031), .B(n13032), .Z(n13029) );
  XNOR2_X1 U13056 ( .A(n13033), .B(n13034), .ZN(n12770) );
  XNOR2_X1 U13057 ( .A(n13035), .B(n13036), .ZN(n13034) );
  XOR2_X1 U13058 ( .A(n13037), .B(n13038), .Z(n12774) );
  XOR2_X1 U13059 ( .A(n13039), .B(n13040), .Z(n13038) );
  NAND2_X1 U13060 ( .A1(a_19_), .A2(b_11_), .ZN(n13040) );
  XNOR2_X1 U13061 ( .A(n13041), .B(n13042), .ZN(n12671) );
  XOR2_X1 U13062 ( .A(n13043), .B(n13044), .Z(n13042) );
  NAND2_X1 U13063 ( .A1(a_18_), .A2(b_11_), .ZN(n13044) );
  XOR2_X1 U13064 ( .A(n13045), .B(n13046), .Z(n12777) );
  XOR2_X1 U13065 ( .A(n13047), .B(n13048), .Z(n13045) );
  NOR2_X1 U13066 ( .A1(n7818), .A2(n7723), .ZN(n13048) );
  XOR2_X1 U13067 ( .A(n13049), .B(n13050), .Z(n12781) );
  XOR2_X1 U13068 ( .A(n13051), .B(n13052), .Z(n13049) );
  NOR2_X1 U13069 ( .A1(n7818), .A2(n7743), .ZN(n13052) );
  INV_X1 U13070 ( .A(n7800), .ZN(n12792) );
  NAND2_X1 U13071 ( .A1(b_12_), .A2(a_12_), .ZN(n7800) );
  XOR2_X1 U13072 ( .A(n13053), .B(n13054), .Z(n12806) );
  XOR2_X1 U13073 ( .A(n13055), .B(n13056), .Z(n13054) );
  NAND2_X1 U13074 ( .A1(a_9_), .A2(b_11_), .ZN(n13056) );
  XOR2_X1 U13075 ( .A(n13057), .B(n13058), .Z(n12810) );
  XOR2_X1 U13076 ( .A(n13059), .B(n13060), .Z(n13057) );
  NOR2_X1 U13077 ( .A1(n7818), .A2(n8059), .ZN(n13060) );
  XNOR2_X1 U13078 ( .A(n13061), .B(n13062), .ZN(n12827) );
  XOR2_X1 U13079 ( .A(n13063), .B(n13064), .Z(n13061) );
  NOR2_X1 U13080 ( .A1(n7818), .A2(n7934), .ZN(n13064) );
  XOR2_X1 U13081 ( .A(n13065), .B(n13066), .Z(n12831) );
  XOR2_X1 U13082 ( .A(n13067), .B(n13068), .Z(n13065) );
  NOR2_X1 U13083 ( .A1(n7818), .A2(n7945), .ZN(n13068) );
  XOR2_X1 U13084 ( .A(n13069), .B(n13070), .Z(n12835) );
  XOR2_X1 U13085 ( .A(n13071), .B(n13072), .Z(n13069) );
  NOR2_X1 U13086 ( .A1(n7818), .A2(n7965), .ZN(n13072) );
  XOR2_X1 U13087 ( .A(n13073), .B(n13074), .Z(n12839) );
  XOR2_X1 U13088 ( .A(n13075), .B(n13076), .Z(n13073) );
  NOR2_X1 U13089 ( .A1(n7818), .A2(n7973), .ZN(n13076) );
  NOR2_X1 U13090 ( .A1(n13077), .A2(n8217), .ZN(n12843) );
  XOR2_X1 U13091 ( .A(n13078), .B(n13079), .Z(n8217) );
  XNOR2_X1 U13092 ( .A(n13080), .B(n13081), .ZN(n13078) );
  AND2_X1 U13093 ( .A1(n8216), .A2(n8215), .ZN(n13077) );
  NAND2_X1 U13094 ( .A1(n13082), .A2(n8214), .ZN(n8186) );
  NOR2_X1 U13095 ( .A1(n8216), .A2(n8215), .ZN(n8214) );
  AND2_X1 U13096 ( .A1(n13083), .A2(n13084), .ZN(n8215) );
  NAND2_X1 U13097 ( .A1(n13081), .A2(n13085), .ZN(n13084) );
  NAND2_X1 U13098 ( .A1(n13080), .A2(n13079), .ZN(n13085) );
  NOR2_X1 U13099 ( .A1(n7818), .A2(n8307), .ZN(n13081) );
  OR2_X1 U13100 ( .A1(n13079), .A2(n13080), .ZN(n13083) );
  AND2_X1 U13101 ( .A1(n13086), .A2(n13087), .ZN(n13080) );
  NAND2_X1 U13102 ( .A1(n13088), .A2(a_1_), .ZN(n13087) );
  NOR2_X1 U13103 ( .A1(n13089), .A2(n7818), .ZN(n13088) );
  NOR2_X1 U13104 ( .A1(n13074), .A2(n13075), .ZN(n13089) );
  NAND2_X1 U13105 ( .A1(n13074), .A2(n13075), .ZN(n13086) );
  NAND2_X1 U13106 ( .A1(n13090), .A2(n13091), .ZN(n13075) );
  NAND2_X1 U13107 ( .A1(n13092), .A2(a_2_), .ZN(n13091) );
  NOR2_X1 U13108 ( .A1(n13093), .A2(n7818), .ZN(n13092) );
  NOR2_X1 U13109 ( .A1(n13070), .A2(n13071), .ZN(n13093) );
  NAND2_X1 U13110 ( .A1(n13070), .A2(n13071), .ZN(n13090) );
  NAND2_X1 U13111 ( .A1(n13094), .A2(n13095), .ZN(n13071) );
  NAND2_X1 U13112 ( .A1(n13096), .A2(a_3_), .ZN(n13095) );
  NOR2_X1 U13113 ( .A1(n13097), .A2(n7818), .ZN(n13096) );
  NOR2_X1 U13114 ( .A1(n13066), .A2(n13067), .ZN(n13097) );
  NAND2_X1 U13115 ( .A1(n13066), .A2(n13067), .ZN(n13094) );
  NAND2_X1 U13116 ( .A1(n13098), .A2(n13099), .ZN(n13067) );
  NAND2_X1 U13117 ( .A1(n13100), .A2(a_4_), .ZN(n13099) );
  NOR2_X1 U13118 ( .A1(n13101), .A2(n7818), .ZN(n13100) );
  NOR2_X1 U13119 ( .A1(n13062), .A2(n13063), .ZN(n13101) );
  NAND2_X1 U13120 ( .A1(n13062), .A2(n13063), .ZN(n13098) );
  NAND2_X1 U13121 ( .A1(n13102), .A2(n13103), .ZN(n13063) );
  NAND2_X1 U13122 ( .A1(n13104), .A2(a_5_), .ZN(n13103) );
  NOR2_X1 U13123 ( .A1(n13105), .A2(n7818), .ZN(n13104) );
  NOR2_X1 U13124 ( .A1(n12863), .A2(n12864), .ZN(n13105) );
  NAND2_X1 U13125 ( .A1(n12863), .A2(n12864), .ZN(n13102) );
  NAND2_X1 U13126 ( .A1(n13106), .A2(n13107), .ZN(n12864) );
  NAND2_X1 U13127 ( .A1(n13108), .A2(a_6_), .ZN(n13107) );
  NOR2_X1 U13128 ( .A1(n13109), .A2(n7818), .ZN(n13108) );
  NOR2_X1 U13129 ( .A1(n12871), .A2(n12872), .ZN(n13109) );
  NAND2_X1 U13130 ( .A1(n12871), .A2(n12872), .ZN(n13106) );
  NAND2_X1 U13131 ( .A1(n13110), .A2(n13111), .ZN(n12872) );
  NAND2_X1 U13132 ( .A1(n13112), .A2(a_7_), .ZN(n13111) );
  NOR2_X1 U13133 ( .A1(n13113), .A2(n7818), .ZN(n13112) );
  NOR2_X1 U13134 ( .A1(n12879), .A2(n12880), .ZN(n13113) );
  NAND2_X1 U13135 ( .A1(n12879), .A2(n12880), .ZN(n13110) );
  NAND2_X1 U13136 ( .A1(n13114), .A2(n13115), .ZN(n12880) );
  NAND2_X1 U13137 ( .A1(n13116), .A2(a_8_), .ZN(n13115) );
  NOR2_X1 U13138 ( .A1(n13117), .A2(n7818), .ZN(n13116) );
  NOR2_X1 U13139 ( .A1(n13058), .A2(n13059), .ZN(n13117) );
  NAND2_X1 U13140 ( .A1(n13058), .A2(n13059), .ZN(n13114) );
  NAND2_X1 U13141 ( .A1(n13118), .A2(n13119), .ZN(n13059) );
  NAND2_X1 U13142 ( .A1(n13120), .A2(a_9_), .ZN(n13119) );
  NOR2_X1 U13143 ( .A1(n13121), .A2(n7818), .ZN(n13120) );
  NOR2_X1 U13144 ( .A1(n13053), .A2(n13055), .ZN(n13121) );
  NAND2_X1 U13145 ( .A1(n13053), .A2(n13055), .ZN(n13118) );
  NAND2_X1 U13146 ( .A1(n13122), .A2(n13123), .ZN(n13055) );
  NAND2_X1 U13147 ( .A1(n13124), .A2(a_10_), .ZN(n13123) );
  NOR2_X1 U13148 ( .A1(n13125), .A2(n7818), .ZN(n13124) );
  NOR2_X1 U13149 ( .A1(n12894), .A2(n12896), .ZN(n13125) );
  NAND2_X1 U13150 ( .A1(n12894), .A2(n12896), .ZN(n13122) );
  NAND2_X1 U13151 ( .A1(n13126), .A2(n13127), .ZN(n12896) );
  NAND2_X1 U13152 ( .A1(n12901), .A2(n13128), .ZN(n13127) );
  OR2_X1 U13153 ( .A1(n12903), .A2(n7812), .ZN(n13128) );
  XNOR2_X1 U13154 ( .A(n13129), .B(n13130), .ZN(n12901) );
  NAND2_X1 U13155 ( .A1(n13131), .A2(n13132), .ZN(n13129) );
  NAND2_X1 U13156 ( .A1(n7812), .A2(n12903), .ZN(n13126) );
  NAND2_X1 U13157 ( .A1(n13133), .A2(n13134), .ZN(n12903) );
  NAND2_X1 U13158 ( .A1(n13135), .A2(a_12_), .ZN(n13134) );
  NOR2_X1 U13159 ( .A1(n13136), .A2(n7818), .ZN(n13135) );
  NOR2_X1 U13160 ( .A1(n12908), .A2(n12910), .ZN(n13136) );
  NAND2_X1 U13161 ( .A1(n12908), .A2(n12910), .ZN(n13133) );
  NAND2_X1 U13162 ( .A1(n13137), .A2(n13138), .ZN(n12910) );
  NAND2_X1 U13163 ( .A1(n13139), .A2(a_13_), .ZN(n13138) );
  NOR2_X1 U13164 ( .A1(n13140), .A2(n7818), .ZN(n13139) );
  NOR2_X1 U13165 ( .A1(n12916), .A2(n12917), .ZN(n13140) );
  NAND2_X1 U13166 ( .A1(n12916), .A2(n12917), .ZN(n13137) );
  NAND2_X1 U13167 ( .A1(n13141), .A2(n13142), .ZN(n12917) );
  NAND2_X1 U13168 ( .A1(n13143), .A2(a_14_), .ZN(n13142) );
  NOR2_X1 U13169 ( .A1(n13144), .A2(n7818), .ZN(n13143) );
  NOR2_X1 U13170 ( .A1(n12924), .A2(n12925), .ZN(n13144) );
  NAND2_X1 U13171 ( .A1(n12924), .A2(n12925), .ZN(n13141) );
  NAND2_X1 U13172 ( .A1(n13145), .A2(n13146), .ZN(n12925) );
  NAND2_X1 U13173 ( .A1(n13147), .A2(a_15_), .ZN(n13146) );
  NOR2_X1 U13174 ( .A1(n13148), .A2(n7818), .ZN(n13147) );
  NOR2_X1 U13175 ( .A1(n12932), .A2(n12933), .ZN(n13148) );
  NAND2_X1 U13176 ( .A1(n12932), .A2(n12933), .ZN(n13145) );
  NAND2_X1 U13177 ( .A1(n13149), .A2(n13150), .ZN(n12933) );
  NAND2_X1 U13178 ( .A1(n13151), .A2(a_16_), .ZN(n13150) );
  NOR2_X1 U13179 ( .A1(n13152), .A2(n7818), .ZN(n13151) );
  NOR2_X1 U13180 ( .A1(n13050), .A2(n13051), .ZN(n13152) );
  NAND2_X1 U13181 ( .A1(n13050), .A2(n13051), .ZN(n13149) );
  NAND2_X1 U13182 ( .A1(n13153), .A2(n13154), .ZN(n13051) );
  NAND2_X1 U13183 ( .A1(n13155), .A2(a_17_), .ZN(n13154) );
  NOR2_X1 U13184 ( .A1(n13156), .A2(n7818), .ZN(n13155) );
  NOR2_X1 U13185 ( .A1(n13046), .A2(n13047), .ZN(n13156) );
  NAND2_X1 U13186 ( .A1(n13046), .A2(n13047), .ZN(n13153) );
  NAND2_X1 U13187 ( .A1(n13157), .A2(n13158), .ZN(n13047) );
  NAND2_X1 U13188 ( .A1(n13159), .A2(a_18_), .ZN(n13158) );
  NOR2_X1 U13189 ( .A1(n13160), .A2(n7818), .ZN(n13159) );
  NOR2_X1 U13190 ( .A1(n13041), .A2(n13043), .ZN(n13160) );
  NAND2_X1 U13191 ( .A1(n13041), .A2(n13043), .ZN(n13157) );
  NAND2_X1 U13192 ( .A1(n13161), .A2(n13162), .ZN(n13043) );
  NAND2_X1 U13193 ( .A1(n13163), .A2(a_19_), .ZN(n13162) );
  NOR2_X1 U13194 ( .A1(n13164), .A2(n7818), .ZN(n13163) );
  NOR2_X1 U13195 ( .A1(n13037), .A2(n13039), .ZN(n13164) );
  NAND2_X1 U13196 ( .A1(n13037), .A2(n13039), .ZN(n13161) );
  NAND2_X1 U13197 ( .A1(n13165), .A2(n13166), .ZN(n13039) );
  NAND2_X1 U13198 ( .A1(n13036), .A2(n13167), .ZN(n13166) );
  OR2_X1 U13199 ( .A1(n13035), .A2(n13033), .ZN(n13167) );
  NOR2_X1 U13200 ( .A1(n7676), .A2(n7818), .ZN(n13036) );
  NAND2_X1 U13201 ( .A1(n13033), .A2(n13035), .ZN(n13165) );
  NAND2_X1 U13202 ( .A1(n13168), .A2(n13169), .ZN(n13035) );
  NAND2_X1 U13203 ( .A1(n13032), .A2(n13170), .ZN(n13169) );
  OR2_X1 U13204 ( .A1(n13031), .A2(n13030), .ZN(n13170) );
  NOR2_X1 U13205 ( .A1(n7656), .A2(n7818), .ZN(n13032) );
  NAND2_X1 U13206 ( .A1(n13030), .A2(n13031), .ZN(n13168) );
  NAND2_X1 U13207 ( .A1(n13171), .A2(n13172), .ZN(n13031) );
  NAND2_X1 U13208 ( .A1(n13173), .A2(a_22_), .ZN(n13172) );
  NOR2_X1 U13209 ( .A1(n13174), .A2(n7818), .ZN(n13173) );
  NOR2_X1 U13210 ( .A1(n13026), .A2(n13027), .ZN(n13174) );
  NAND2_X1 U13211 ( .A1(n13026), .A2(n13027), .ZN(n13171) );
  NAND2_X1 U13212 ( .A1(n13175), .A2(n13176), .ZN(n13027) );
  NAND2_X1 U13213 ( .A1(n13024), .A2(n13177), .ZN(n13176) );
  OR2_X1 U13214 ( .A1(n13023), .A2(n13022), .ZN(n13177) );
  NOR2_X1 U13215 ( .A1(n7624), .A2(n7818), .ZN(n13024) );
  NAND2_X1 U13216 ( .A1(n13022), .A2(n13023), .ZN(n13175) );
  NAND2_X1 U13217 ( .A1(n13019), .A2(n13178), .ZN(n13023) );
  NAND2_X1 U13218 ( .A1(n13018), .A2(n13020), .ZN(n13178) );
  NAND2_X1 U13219 ( .A1(n13179), .A2(n13180), .ZN(n13020) );
  NAND2_X1 U13220 ( .A1(a_24_), .A2(b_11_), .ZN(n13180) );
  INV_X1 U13221 ( .A(n13181), .ZN(n13179) );
  XNOR2_X1 U13222 ( .A(n13182), .B(n13183), .ZN(n13018) );
  XOR2_X1 U13223 ( .A(n13184), .B(n13185), .Z(n13183) );
  NAND2_X1 U13224 ( .A1(a_25_), .A2(b_10_), .ZN(n13185) );
  NAND2_X1 U13225 ( .A1(a_24_), .A2(n13181), .ZN(n13019) );
  NAND2_X1 U13226 ( .A1(n13186), .A2(n13187), .ZN(n13181) );
  NAND2_X1 U13227 ( .A1(n13188), .A2(a_25_), .ZN(n13187) );
  NOR2_X1 U13228 ( .A1(n13189), .A2(n7818), .ZN(n13188) );
  NOR2_X1 U13229 ( .A1(n12971), .A2(n12972), .ZN(n13189) );
  NAND2_X1 U13230 ( .A1(n12971), .A2(n12972), .ZN(n13186) );
  NAND2_X1 U13231 ( .A1(n13190), .A2(n13191), .ZN(n12972) );
  NAND2_X1 U13232 ( .A1(n13192), .A2(a_26_), .ZN(n13191) );
  NOR2_X1 U13233 ( .A1(n13193), .A2(n7818), .ZN(n13192) );
  NOR2_X1 U13234 ( .A1(n13014), .A2(n13016), .ZN(n13193) );
  NAND2_X1 U13235 ( .A1(n13014), .A2(n13016), .ZN(n13190) );
  NAND2_X1 U13236 ( .A1(n13194), .A2(n13195), .ZN(n13016) );
  NAND2_X1 U13237 ( .A1(n13012), .A2(n13196), .ZN(n13195) );
  NAND2_X1 U13238 ( .A1(n13011), .A2(n13010), .ZN(n13196) );
  NOR2_X1 U13239 ( .A1(n7563), .A2(n7818), .ZN(n13012) );
  OR2_X1 U13240 ( .A1(n13010), .A2(n13011), .ZN(n13194) );
  AND2_X1 U13241 ( .A1(n13007), .A2(n13197), .ZN(n13011) );
  NAND2_X1 U13242 ( .A1(n13006), .A2(n13008), .ZN(n13197) );
  NAND2_X1 U13243 ( .A1(n13198), .A2(n13199), .ZN(n13008) );
  NAND2_X1 U13244 ( .A1(a_28_), .A2(b_11_), .ZN(n13199) );
  INV_X1 U13245 ( .A(n13200), .ZN(n13198) );
  XOR2_X1 U13246 ( .A(n13201), .B(n13202), .Z(n13006) );
  NOR2_X1 U13247 ( .A1(n13001), .A2(n7529), .ZN(n13202) );
  XOR2_X1 U13248 ( .A(n13203), .B(n13204), .Z(n13201) );
  NAND2_X1 U13249 ( .A1(a_28_), .A2(n13200), .ZN(n13007) );
  NAND2_X1 U13250 ( .A1(n13205), .A2(n13206), .ZN(n13200) );
  NAND2_X1 U13251 ( .A1(n13207), .A2(a_29_), .ZN(n13206) );
  NOR2_X1 U13252 ( .A1(n13208), .A2(n7818), .ZN(n13207) );
  NOR2_X1 U13253 ( .A1(n12991), .A2(n12992), .ZN(n13208) );
  NAND2_X1 U13254 ( .A1(n12991), .A2(n12992), .ZN(n13205) );
  NAND2_X1 U13255 ( .A1(n13209), .A2(n13210), .ZN(n12992) );
  NAND2_X1 U13256 ( .A1(n13211), .A2(b_10_), .ZN(n13210) );
  NOR2_X1 U13257 ( .A1(n13212), .A2(n7515), .ZN(n13211) );
  NOR2_X1 U13258 ( .A1(n8679), .A2(n7849), .ZN(n13212) );
  NAND2_X1 U13259 ( .A1(n13213), .A2(a_31_), .ZN(n13209) );
  NOR2_X1 U13260 ( .A1(n13214), .A2(n7849), .ZN(n13213) );
  NOR2_X1 U13261 ( .A1(n8676), .A2(n13001), .ZN(n13214) );
  AND2_X1 U13262 ( .A1(n13215), .A2(n8049), .ZN(n12991) );
  NOR2_X1 U13263 ( .A1(n7818), .A2(n13001), .ZN(n13215) );
  XOR2_X1 U13264 ( .A(n13216), .B(n13217), .Z(n13010) );
  NAND2_X1 U13265 ( .A1(n13218), .A2(n13219), .ZN(n13216) );
  XNOR2_X1 U13266 ( .A(n13220), .B(n13221), .ZN(n13014) );
  XNOR2_X1 U13267 ( .A(n13222), .B(n13223), .ZN(n13220) );
  XOR2_X1 U13268 ( .A(n13224), .B(n13225), .Z(n12971) );
  XNOR2_X1 U13269 ( .A(n13226), .B(n13227), .ZN(n13224) );
  NAND2_X1 U13270 ( .A1(a_26_), .A2(b_10_), .ZN(n13226) );
  XNOR2_X1 U13271 ( .A(n13228), .B(n13229), .ZN(n13022) );
  NAND2_X1 U13272 ( .A1(n13230), .A2(n13231), .ZN(n13228) );
  XOR2_X1 U13273 ( .A(n13232), .B(n13233), .Z(n13026) );
  XOR2_X1 U13274 ( .A(n13234), .B(n13235), .Z(n13232) );
  XOR2_X1 U13275 ( .A(n13236), .B(n13237), .Z(n13030) );
  XOR2_X1 U13276 ( .A(n13238), .B(n13239), .Z(n13236) );
  NOR2_X1 U13277 ( .A1(n13001), .A2(n7645), .ZN(n13239) );
  XOR2_X1 U13278 ( .A(n13240), .B(n13241), .Z(n13033) );
  XOR2_X1 U13279 ( .A(n13242), .B(n13243), .Z(n13240) );
  NOR2_X1 U13280 ( .A1(n7656), .A2(n13001), .ZN(n13243) );
  XNOR2_X1 U13281 ( .A(n13244), .B(n13245), .ZN(n13037) );
  XNOR2_X1 U13282 ( .A(n13246), .B(n13247), .ZN(n13244) );
  XOR2_X1 U13283 ( .A(n13248), .B(n13249), .Z(n13041) );
  XOR2_X1 U13284 ( .A(n13250), .B(n13251), .Z(n13248) );
  XOR2_X1 U13285 ( .A(n13252), .B(n13253), .Z(n13046) );
  XOR2_X1 U13286 ( .A(n13254), .B(n13255), .Z(n13252) );
  XOR2_X1 U13287 ( .A(n13256), .B(n13257), .Z(n13050) );
  XOR2_X1 U13288 ( .A(n13258), .B(n13259), .Z(n13256) );
  XNOR2_X1 U13289 ( .A(n13260), .B(n13261), .ZN(n12932) );
  XOR2_X1 U13290 ( .A(n13262), .B(n13263), .Z(n13261) );
  NAND2_X1 U13291 ( .A1(a_16_), .A2(b_10_), .ZN(n13263) );
  XNOR2_X1 U13292 ( .A(n13264), .B(n13265), .ZN(n12924) );
  NAND2_X1 U13293 ( .A1(n13266), .A2(n13267), .ZN(n13264) );
  XNOR2_X1 U13294 ( .A(n13268), .B(n13269), .ZN(n12916) );
  NAND2_X1 U13295 ( .A1(n13270), .A2(n13271), .ZN(n13268) );
  XNOR2_X1 U13296 ( .A(n13272), .B(n13273), .ZN(n12908) );
  NAND2_X1 U13297 ( .A1(n13274), .A2(n13275), .ZN(n13272) );
  NOR2_X1 U13298 ( .A1(n7817), .A2(n7818), .ZN(n7812) );
  XNOR2_X1 U13299 ( .A(n13276), .B(n13277), .ZN(n12894) );
  NAND2_X1 U13300 ( .A1(n13278), .A2(n13279), .ZN(n13276) );
  XNOR2_X1 U13301 ( .A(n13280), .B(n13281), .ZN(n13053) );
  XNOR2_X1 U13302 ( .A(n13282), .B(n7831), .ZN(n13281) );
  XOR2_X1 U13303 ( .A(n13283), .B(n13284), .Z(n13058) );
  NOR2_X1 U13304 ( .A1(n13285), .A2(n13286), .ZN(n13284) );
  NOR2_X1 U13305 ( .A1(n13287), .A2(n13288), .ZN(n13285) );
  NOR2_X1 U13306 ( .A1(n13001), .A2(n7848), .ZN(n13287) );
  XOR2_X1 U13307 ( .A(n13289), .B(n13290), .Z(n12879) );
  XOR2_X1 U13308 ( .A(n13291), .B(n13292), .Z(n13289) );
  XOR2_X1 U13309 ( .A(n13293), .B(n13294), .Z(n12871) );
  XOR2_X1 U13310 ( .A(n13295), .B(n13296), .Z(n13293) );
  XOR2_X1 U13311 ( .A(n13297), .B(n13298), .Z(n12863) );
  XOR2_X1 U13312 ( .A(n13299), .B(n13300), .Z(n13297) );
  XNOR2_X1 U13313 ( .A(n13301), .B(n13302), .ZN(n13062) );
  XNOR2_X1 U13314 ( .A(n13303), .B(n13304), .ZN(n13301) );
  XNOR2_X1 U13315 ( .A(n13305), .B(n13306), .ZN(n13066) );
  XNOR2_X1 U13316 ( .A(n13307), .B(n13308), .ZN(n13306) );
  XNOR2_X1 U13317 ( .A(n13309), .B(n13310), .ZN(n13070) );
  XNOR2_X1 U13318 ( .A(n13311), .B(n13312), .ZN(n13310) );
  XOR2_X1 U13319 ( .A(n13313), .B(n13314), .Z(n13074) );
  XOR2_X1 U13320 ( .A(n13315), .B(n13316), .Z(n13313) );
  XNOR2_X1 U13321 ( .A(n13317), .B(n13318), .ZN(n13079) );
  XOR2_X1 U13322 ( .A(n13319), .B(n13320), .Z(n13317) );
  NOR2_X1 U13323 ( .A1(n13001), .A2(n7973), .ZN(n13320) );
  XOR2_X1 U13324 ( .A(n13321), .B(n13322), .Z(n8216) );
  XNOR2_X1 U13325 ( .A(n13323), .B(n13324), .ZN(n13322) );
  XOR2_X1 U13326 ( .A(n8209), .B(n13325), .Z(n13082) );
  NAND2_X1 U13327 ( .A1(n13326), .A2(n13327), .ZN(n7480) );
  NAND2_X1 U13328 ( .A1(n13328), .A2(n13329), .ZN(n13327) );
  OR2_X1 U13329 ( .A1(n13330), .A2(n13331), .ZN(n13328) );
  OR2_X1 U13330 ( .A1(n8209), .A2(n13325), .ZN(n13326) );
  NAND2_X1 U13331 ( .A1(n13332), .A2(n13333), .ZN(n7479) );
  NOR2_X1 U13332 ( .A1(n13334), .A2(n13325), .ZN(n13333) );
  INV_X1 U13333 ( .A(n8208), .ZN(n13325) );
  NAND2_X1 U13334 ( .A1(n13335), .A2(n13336), .ZN(n8208) );
  NAND2_X1 U13335 ( .A1(n13324), .A2(n13337), .ZN(n13336) );
  OR2_X1 U13336 ( .A1(n13321), .A2(n13323), .ZN(n13337) );
  NOR2_X1 U13337 ( .A1(n13001), .A2(n8307), .ZN(n13324) );
  NAND2_X1 U13338 ( .A1(n13321), .A2(n13323), .ZN(n13335) );
  NAND2_X1 U13339 ( .A1(n13338), .A2(n13339), .ZN(n13323) );
  NAND2_X1 U13340 ( .A1(n13340), .A2(a_1_), .ZN(n13339) );
  NOR2_X1 U13341 ( .A1(n13341), .A2(n13001), .ZN(n13340) );
  NOR2_X1 U13342 ( .A1(n13319), .A2(n13318), .ZN(n13341) );
  NAND2_X1 U13343 ( .A1(n13318), .A2(n13319), .ZN(n13338) );
  NAND2_X1 U13344 ( .A1(n13342), .A2(n13343), .ZN(n13319) );
  NAND2_X1 U13345 ( .A1(n13316), .A2(n13344), .ZN(n13343) );
  OR2_X1 U13346 ( .A1(n13314), .A2(n13315), .ZN(n13344) );
  NOR2_X1 U13347 ( .A1(n7965), .A2(n13001), .ZN(n13316) );
  NAND2_X1 U13348 ( .A1(n13314), .A2(n13315), .ZN(n13342) );
  NAND2_X1 U13349 ( .A1(n13345), .A2(n13346), .ZN(n13315) );
  NAND2_X1 U13350 ( .A1(n13312), .A2(n13347), .ZN(n13346) );
  OR2_X1 U13351 ( .A1(n13309), .A2(n13311), .ZN(n13347) );
  NOR2_X1 U13352 ( .A1(n7945), .A2(n13001), .ZN(n13312) );
  NAND2_X1 U13353 ( .A1(n13309), .A2(n13311), .ZN(n13345) );
  NAND2_X1 U13354 ( .A1(n13348), .A2(n13349), .ZN(n13311) );
  NAND2_X1 U13355 ( .A1(n13308), .A2(n13350), .ZN(n13349) );
  OR2_X1 U13356 ( .A1(n13305), .A2(n13307), .ZN(n13350) );
  NOR2_X1 U13357 ( .A1(n7934), .A2(n13001), .ZN(n13308) );
  NAND2_X1 U13358 ( .A1(n13305), .A2(n13307), .ZN(n13348) );
  NAND2_X1 U13359 ( .A1(n13351), .A2(n13352), .ZN(n13307) );
  NAND2_X1 U13360 ( .A1(n13304), .A2(n13353), .ZN(n13352) );
  NAND2_X1 U13361 ( .A1(n13303), .A2(n13302), .ZN(n13353) );
  NOR2_X1 U13362 ( .A1(n7914), .A2(n13001), .ZN(n13304) );
  OR2_X1 U13363 ( .A1(n13302), .A2(n13303), .ZN(n13351) );
  AND2_X1 U13364 ( .A1(n13354), .A2(n13355), .ZN(n13303) );
  NAND2_X1 U13365 ( .A1(n13299), .A2(n13356), .ZN(n13355) );
  OR2_X1 U13366 ( .A1(n13298), .A2(n13300), .ZN(n13356) );
  NOR2_X1 U13367 ( .A1(n8061), .A2(n13001), .ZN(n13299) );
  NAND2_X1 U13368 ( .A1(n13298), .A2(n13300), .ZN(n13354) );
  NAND2_X1 U13369 ( .A1(n13357), .A2(n13358), .ZN(n13300) );
  NAND2_X1 U13370 ( .A1(n13296), .A2(n13359), .ZN(n13358) );
  OR2_X1 U13371 ( .A1(n13294), .A2(n13295), .ZN(n13359) );
  NOR2_X1 U13372 ( .A1(n7884), .A2(n13001), .ZN(n13296) );
  NAND2_X1 U13373 ( .A1(n13294), .A2(n13295), .ZN(n13357) );
  NAND2_X1 U13374 ( .A1(n13360), .A2(n13361), .ZN(n13295) );
  NAND2_X1 U13375 ( .A1(n13292), .A2(n13362), .ZN(n13361) );
  OR2_X1 U13376 ( .A1(n13290), .A2(n13291), .ZN(n13362) );
  NOR2_X1 U13377 ( .A1(n8059), .A2(n13001), .ZN(n13292) );
  NAND2_X1 U13378 ( .A1(n13290), .A2(n13291), .ZN(n13360) );
  OR2_X1 U13379 ( .A1(n13286), .A2(n13363), .ZN(n13291) );
  AND2_X1 U13380 ( .A1(n13283), .A2(n13364), .ZN(n13363) );
  NAND2_X1 U13381 ( .A1(n13365), .A2(n13366), .ZN(n13364) );
  NAND2_X1 U13382 ( .A1(a_9_), .A2(b_10_), .ZN(n13366) );
  XOR2_X1 U13383 ( .A(n13367), .B(n13368), .Z(n13283) );
  XOR2_X1 U13384 ( .A(n13369), .B(n13370), .Z(n13367) );
  NOR2_X1 U13385 ( .A1(n7849), .A2(n7837), .ZN(n13370) );
  NOR2_X1 U13386 ( .A1(n7848), .A2(n13365), .ZN(n13286) );
  INV_X1 U13387 ( .A(n13288), .ZN(n13365) );
  NAND2_X1 U13388 ( .A1(n13371), .A2(n13372), .ZN(n13288) );
  NAND2_X1 U13389 ( .A1(n13280), .A2(n13373), .ZN(n13372) );
  OR2_X1 U13390 ( .A1(n13282), .A2(n7831), .ZN(n13373) );
  XOR2_X1 U13391 ( .A(n13374), .B(n13375), .Z(n13280) );
  XOR2_X1 U13392 ( .A(n13376), .B(n13377), .Z(n13374) );
  NOR2_X1 U13393 ( .A1(n7817), .A2(n7849), .ZN(n13377) );
  NAND2_X1 U13394 ( .A1(n7831), .A2(n13282), .ZN(n13371) );
  NAND2_X1 U13395 ( .A1(n13278), .A2(n13378), .ZN(n13282) );
  NAND2_X1 U13396 ( .A1(n13277), .A2(n13279), .ZN(n13378) );
  NAND2_X1 U13397 ( .A1(n13379), .A2(n13380), .ZN(n13279) );
  NAND2_X1 U13398 ( .A1(b_10_), .A2(a_11_), .ZN(n13380) );
  INV_X1 U13399 ( .A(n13381), .ZN(n13379) );
  XNOR2_X1 U13400 ( .A(n13382), .B(n13383), .ZN(n13277) );
  XOR2_X1 U13401 ( .A(n13384), .B(n13385), .Z(n13383) );
  NAND2_X1 U13402 ( .A1(a_12_), .A2(b_9_), .ZN(n13385) );
  NAND2_X1 U13403 ( .A1(a_11_), .A2(n13381), .ZN(n13278) );
  NAND2_X1 U13404 ( .A1(n13131), .A2(n13386), .ZN(n13381) );
  NAND2_X1 U13405 ( .A1(n13130), .A2(n13132), .ZN(n13386) );
  NAND2_X1 U13406 ( .A1(n13387), .A2(n13388), .ZN(n13132) );
  NAND2_X1 U13407 ( .A1(a_12_), .A2(b_10_), .ZN(n13388) );
  INV_X1 U13408 ( .A(n13389), .ZN(n13387) );
  XNOR2_X1 U13409 ( .A(n13390), .B(n13391), .ZN(n13130) );
  XOR2_X1 U13410 ( .A(n13392), .B(n13393), .Z(n13391) );
  NAND2_X1 U13411 ( .A1(a_13_), .A2(b_9_), .ZN(n13393) );
  NAND2_X1 U13412 ( .A1(a_12_), .A2(n13389), .ZN(n13131) );
  NAND2_X1 U13413 ( .A1(n13274), .A2(n13394), .ZN(n13389) );
  NAND2_X1 U13414 ( .A1(n13273), .A2(n13275), .ZN(n13394) );
  NAND2_X1 U13415 ( .A1(n13395), .A2(n13396), .ZN(n13275) );
  NAND2_X1 U13416 ( .A1(a_13_), .A2(b_10_), .ZN(n13396) );
  INV_X1 U13417 ( .A(n13397), .ZN(n13395) );
  XNOR2_X1 U13418 ( .A(n13398), .B(n13399), .ZN(n13273) );
  XOR2_X1 U13419 ( .A(n13400), .B(n13401), .Z(n13399) );
  NAND2_X1 U13420 ( .A1(a_14_), .A2(b_9_), .ZN(n13401) );
  NAND2_X1 U13421 ( .A1(a_13_), .A2(n13397), .ZN(n13274) );
  NAND2_X1 U13422 ( .A1(n13270), .A2(n13402), .ZN(n13397) );
  NAND2_X1 U13423 ( .A1(n13269), .A2(n13271), .ZN(n13402) );
  NAND2_X1 U13424 ( .A1(n13403), .A2(n13404), .ZN(n13271) );
  NAND2_X1 U13425 ( .A1(a_14_), .A2(b_10_), .ZN(n13404) );
  INV_X1 U13426 ( .A(n13405), .ZN(n13403) );
  XNOR2_X1 U13427 ( .A(n13406), .B(n13407), .ZN(n13269) );
  XOR2_X1 U13428 ( .A(n13408), .B(n13409), .Z(n13407) );
  NAND2_X1 U13429 ( .A1(a_15_), .A2(b_9_), .ZN(n13409) );
  NAND2_X1 U13430 ( .A1(a_14_), .A2(n13405), .ZN(n13270) );
  NAND2_X1 U13431 ( .A1(n13266), .A2(n13410), .ZN(n13405) );
  NAND2_X1 U13432 ( .A1(n13265), .A2(n13267), .ZN(n13410) );
  NAND2_X1 U13433 ( .A1(n13411), .A2(n13412), .ZN(n13267) );
  NAND2_X1 U13434 ( .A1(a_15_), .A2(b_10_), .ZN(n13412) );
  INV_X1 U13435 ( .A(n13413), .ZN(n13411) );
  XNOR2_X1 U13436 ( .A(n13414), .B(n13415), .ZN(n13265) );
  XOR2_X1 U13437 ( .A(n13416), .B(n13417), .Z(n13415) );
  NAND2_X1 U13438 ( .A1(a_16_), .A2(b_9_), .ZN(n13417) );
  NAND2_X1 U13439 ( .A1(a_15_), .A2(n13413), .ZN(n13266) );
  NAND2_X1 U13440 ( .A1(n13418), .A2(n13419), .ZN(n13413) );
  NAND2_X1 U13441 ( .A1(n13420), .A2(a_16_), .ZN(n13419) );
  NOR2_X1 U13442 ( .A1(n13421), .A2(n13001), .ZN(n13420) );
  NOR2_X1 U13443 ( .A1(n13260), .A2(n13262), .ZN(n13421) );
  NAND2_X1 U13444 ( .A1(n13260), .A2(n13262), .ZN(n13418) );
  NAND2_X1 U13445 ( .A1(n13422), .A2(n13423), .ZN(n13262) );
  NAND2_X1 U13446 ( .A1(n13259), .A2(n13424), .ZN(n13423) );
  OR2_X1 U13447 ( .A1(n13257), .A2(n13258), .ZN(n13424) );
  NOR2_X1 U13448 ( .A1(n7723), .A2(n13001), .ZN(n13259) );
  NAND2_X1 U13449 ( .A1(n13257), .A2(n13258), .ZN(n13422) );
  NAND2_X1 U13450 ( .A1(n13425), .A2(n13426), .ZN(n13258) );
  NAND2_X1 U13451 ( .A1(n13255), .A2(n13427), .ZN(n13426) );
  OR2_X1 U13452 ( .A1(n13253), .A2(n13254), .ZN(n13427) );
  NOR2_X1 U13453 ( .A1(n7707), .A2(n13001), .ZN(n13255) );
  NAND2_X1 U13454 ( .A1(n13253), .A2(n13254), .ZN(n13425) );
  NAND2_X1 U13455 ( .A1(n13428), .A2(n13429), .ZN(n13254) );
  NAND2_X1 U13456 ( .A1(n13251), .A2(n13430), .ZN(n13429) );
  OR2_X1 U13457 ( .A1(n13249), .A2(n13250), .ZN(n13430) );
  NOR2_X1 U13458 ( .A1(n7687), .A2(n13001), .ZN(n13251) );
  NAND2_X1 U13459 ( .A1(n13249), .A2(n13250), .ZN(n13428) );
  NAND2_X1 U13460 ( .A1(n13431), .A2(n13432), .ZN(n13250) );
  NAND2_X1 U13461 ( .A1(n13246), .A2(n13433), .ZN(n13432) );
  NAND2_X1 U13462 ( .A1(n13247), .A2(n13245), .ZN(n13433) );
  NOR2_X1 U13463 ( .A1(n13001), .A2(n7676), .ZN(n13246) );
  OR2_X1 U13464 ( .A1(n13245), .A2(n13247), .ZN(n13431) );
  AND2_X1 U13465 ( .A1(n13434), .A2(n13435), .ZN(n13247) );
  NAND2_X1 U13466 ( .A1(n13436), .A2(b_10_), .ZN(n13435) );
  NOR2_X1 U13467 ( .A1(n13437), .A2(n7656), .ZN(n13436) );
  NOR2_X1 U13468 ( .A1(n13242), .A2(n13241), .ZN(n13437) );
  NAND2_X1 U13469 ( .A1(n13241), .A2(n13242), .ZN(n13434) );
  NAND2_X1 U13470 ( .A1(n13438), .A2(n13439), .ZN(n13242) );
  NAND2_X1 U13471 ( .A1(n13440), .A2(a_22_), .ZN(n13439) );
  NOR2_X1 U13472 ( .A1(n13441), .A2(n13001), .ZN(n13440) );
  NOR2_X1 U13473 ( .A1(n13237), .A2(n13238), .ZN(n13441) );
  NAND2_X1 U13474 ( .A1(n13237), .A2(n13238), .ZN(n13438) );
  NAND2_X1 U13475 ( .A1(n13442), .A2(n13443), .ZN(n13238) );
  NAND2_X1 U13476 ( .A1(n13235), .A2(n13444), .ZN(n13443) );
  OR2_X1 U13477 ( .A1(n13233), .A2(n13234), .ZN(n13444) );
  NOR2_X1 U13478 ( .A1(n13001), .A2(n7624), .ZN(n13235) );
  NAND2_X1 U13479 ( .A1(n13233), .A2(n13234), .ZN(n13442) );
  NAND2_X1 U13480 ( .A1(n13230), .A2(n13445), .ZN(n13234) );
  NAND2_X1 U13481 ( .A1(n13229), .A2(n13231), .ZN(n13445) );
  NAND2_X1 U13482 ( .A1(n13446), .A2(n13447), .ZN(n13231) );
  NAND2_X1 U13483 ( .A1(a_24_), .A2(b_10_), .ZN(n13447) );
  INV_X1 U13484 ( .A(n13448), .ZN(n13446) );
  XNOR2_X1 U13485 ( .A(n13449), .B(n13450), .ZN(n13229) );
  XOR2_X1 U13486 ( .A(n13451), .B(n13452), .Z(n13450) );
  NAND2_X1 U13487 ( .A1(a_25_), .A2(b_9_), .ZN(n13452) );
  NAND2_X1 U13488 ( .A1(a_24_), .A2(n13448), .ZN(n13230) );
  NAND2_X1 U13489 ( .A1(n13453), .A2(n13454), .ZN(n13448) );
  NAND2_X1 U13490 ( .A1(n13455), .A2(a_25_), .ZN(n13454) );
  NOR2_X1 U13491 ( .A1(n13456), .A2(n13001), .ZN(n13455) );
  NOR2_X1 U13492 ( .A1(n13182), .A2(n13184), .ZN(n13456) );
  NAND2_X1 U13493 ( .A1(n13182), .A2(n13184), .ZN(n13453) );
  NAND2_X1 U13494 ( .A1(n13457), .A2(n13458), .ZN(n13184) );
  NAND2_X1 U13495 ( .A1(n13459), .A2(a_26_), .ZN(n13458) );
  NOR2_X1 U13496 ( .A1(n13460), .A2(n13001), .ZN(n13459) );
  NOR2_X1 U13497 ( .A1(n13227), .A2(n13225), .ZN(n13460) );
  NAND2_X1 U13498 ( .A1(n13225), .A2(n13227), .ZN(n13457) );
  NAND2_X1 U13499 ( .A1(n13461), .A2(n13462), .ZN(n13227) );
  NAND2_X1 U13500 ( .A1(n13223), .A2(n13463), .ZN(n13462) );
  NAND2_X1 U13501 ( .A1(n13222), .A2(n13221), .ZN(n13463) );
  NOR2_X1 U13502 ( .A1(n13001), .A2(n7563), .ZN(n13223) );
  OR2_X1 U13503 ( .A1(n13221), .A2(n13222), .ZN(n13461) );
  AND2_X1 U13504 ( .A1(n13218), .A2(n13464), .ZN(n13222) );
  NAND2_X1 U13505 ( .A1(n13217), .A2(n13219), .ZN(n13464) );
  NAND2_X1 U13506 ( .A1(n13465), .A2(n13466), .ZN(n13219) );
  NAND2_X1 U13507 ( .A1(a_28_), .A2(b_10_), .ZN(n13466) );
  INV_X1 U13508 ( .A(n13467), .ZN(n13465) );
  XOR2_X1 U13509 ( .A(n13468), .B(n13469), .Z(n13217) );
  NOR2_X1 U13510 ( .A1(n7849), .A2(n7529), .ZN(n13469) );
  XOR2_X1 U13511 ( .A(n13470), .B(n13471), .Z(n13468) );
  NAND2_X1 U13512 ( .A1(a_28_), .A2(n13467), .ZN(n13218) );
  NAND2_X1 U13513 ( .A1(n13472), .A2(n13473), .ZN(n13467) );
  NAND2_X1 U13514 ( .A1(n13474), .A2(a_29_), .ZN(n13473) );
  NOR2_X1 U13515 ( .A1(n13475), .A2(n13001), .ZN(n13474) );
  NOR2_X1 U13516 ( .A1(n13203), .A2(n13204), .ZN(n13475) );
  NAND2_X1 U13517 ( .A1(n13203), .A2(n13204), .ZN(n13472) );
  NAND2_X1 U13518 ( .A1(n13476), .A2(n13477), .ZN(n13204) );
  NAND2_X1 U13519 ( .A1(n13478), .A2(b_8_), .ZN(n13477) );
  NOR2_X1 U13520 ( .A1(n13479), .A2(n8048), .ZN(n13478) );
  NOR2_X1 U13521 ( .A1(n8676), .A2(n7849), .ZN(n13479) );
  NAND2_X1 U13522 ( .A1(n13480), .A2(b_9_), .ZN(n13476) );
  NOR2_X1 U13523 ( .A1(n13481), .A2(n7515), .ZN(n13480) );
  NOR2_X1 U13524 ( .A1(n8679), .A2(n8058), .ZN(n13481) );
  AND2_X1 U13525 ( .A1(n13482), .A2(n8049), .ZN(n13203) );
  INV_X1 U13526 ( .A(n8451), .ZN(n8049) );
  NOR2_X1 U13527 ( .A1(n7849), .A2(n13001), .ZN(n13482) );
  XOR2_X1 U13528 ( .A(n13483), .B(n13484), .Z(n13221) );
  NAND2_X1 U13529 ( .A1(n13485), .A2(n13486), .ZN(n13483) );
  XNOR2_X1 U13530 ( .A(n13487), .B(n13488), .ZN(n13225) );
  XNOR2_X1 U13531 ( .A(n13489), .B(n13490), .ZN(n13487) );
  XOR2_X1 U13532 ( .A(n13491), .B(n13492), .Z(n13182) );
  XNOR2_X1 U13533 ( .A(n13493), .B(n13494), .ZN(n13491) );
  NAND2_X1 U13534 ( .A1(a_26_), .A2(b_9_), .ZN(n13493) );
  XNOR2_X1 U13535 ( .A(n13495), .B(n13496), .ZN(n13233) );
  NAND2_X1 U13536 ( .A1(n13497), .A2(n13498), .ZN(n13495) );
  XOR2_X1 U13537 ( .A(n13499), .B(n13500), .Z(n13237) );
  XOR2_X1 U13538 ( .A(n13501), .B(n13502), .Z(n13499) );
  XNOR2_X1 U13539 ( .A(n13503), .B(n13504), .ZN(n13241) );
  XNOR2_X1 U13540 ( .A(n13505), .B(n13506), .ZN(n13503) );
  XNOR2_X1 U13541 ( .A(n13507), .B(n13508), .ZN(n13245) );
  XOR2_X1 U13542 ( .A(n13509), .B(n13510), .Z(n13507) );
  NOR2_X1 U13543 ( .A1(n7656), .A2(n7849), .ZN(n13510) );
  XNOR2_X1 U13544 ( .A(n13511), .B(n13512), .ZN(n13249) );
  NAND2_X1 U13545 ( .A1(n13513), .A2(n13514), .ZN(n13511) );
  XNOR2_X1 U13546 ( .A(n13515), .B(n13516), .ZN(n13253) );
  NAND2_X1 U13547 ( .A1(n13517), .A2(n13518), .ZN(n13515) );
  XNOR2_X1 U13548 ( .A(n13519), .B(n13520), .ZN(n13257) );
  XOR2_X1 U13549 ( .A(n13521), .B(n13522), .Z(n13520) );
  NAND2_X1 U13550 ( .A1(a_18_), .A2(b_9_), .ZN(n13522) );
  XOR2_X1 U13551 ( .A(n13523), .B(n13524), .Z(n13260) );
  XOR2_X1 U13552 ( .A(n13525), .B(n13526), .Z(n13523) );
  NOR2_X1 U13553 ( .A1(n7849), .A2(n7723), .ZN(n13526) );
  NOR2_X1 U13554 ( .A1(n7837), .A2(n13001), .ZN(n7831) );
  XOR2_X1 U13555 ( .A(n13527), .B(n13528), .Z(n13290) );
  XOR2_X1 U13556 ( .A(n13529), .B(n7843), .Z(n13527) );
  XOR2_X1 U13557 ( .A(n13530), .B(n13531), .Z(n13294) );
  XNOR2_X1 U13558 ( .A(n13532), .B(n13533), .ZN(n13530) );
  NAND2_X1 U13559 ( .A1(a_8_), .A2(b_9_), .ZN(n13532) );
  XOR2_X1 U13560 ( .A(n13534), .B(n13535), .Z(n13298) );
  XNOR2_X1 U13561 ( .A(n13536), .B(n13537), .ZN(n13534) );
  NAND2_X1 U13562 ( .A1(a_7_), .A2(b_9_), .ZN(n13536) );
  XNOR2_X1 U13563 ( .A(n13538), .B(n13539), .ZN(n13302) );
  XOR2_X1 U13564 ( .A(n13540), .B(n13541), .Z(n13538) );
  NOR2_X1 U13565 ( .A1(n7849), .A2(n8061), .ZN(n13541) );
  XOR2_X1 U13566 ( .A(n13542), .B(n13543), .Z(n13305) );
  XOR2_X1 U13567 ( .A(n13544), .B(n13545), .Z(n13542) );
  NOR2_X1 U13568 ( .A1(n7849), .A2(n7914), .ZN(n13545) );
  XOR2_X1 U13569 ( .A(n13546), .B(n13547), .Z(n13309) );
  XOR2_X1 U13570 ( .A(n13548), .B(n13549), .Z(n13546) );
  NOR2_X1 U13571 ( .A1(n7849), .A2(n7934), .ZN(n13549) );
  XOR2_X1 U13572 ( .A(n13550), .B(n13551), .Z(n13314) );
  XOR2_X1 U13573 ( .A(n13552), .B(n13553), .Z(n13550) );
  NOR2_X1 U13574 ( .A1(n7849), .A2(n7945), .ZN(n13553) );
  XNOR2_X1 U13575 ( .A(n13554), .B(n13555), .ZN(n13318) );
  XOR2_X1 U13576 ( .A(n13556), .B(n13557), .Z(n13555) );
  NAND2_X1 U13577 ( .A1(a_2_), .A2(b_9_), .ZN(n13557) );
  XNOR2_X1 U13578 ( .A(n13558), .B(n13559), .ZN(n13321) );
  XOR2_X1 U13579 ( .A(n13560), .B(n13561), .Z(n13559) );
  NAND2_X1 U13580 ( .A1(a_1_), .A2(b_9_), .ZN(n13561) );
  NOR2_X1 U13581 ( .A1(n13562), .A2(n8209), .ZN(n13332) );
  XNOR2_X1 U13582 ( .A(n13563), .B(n13564), .ZN(n8209) );
  XOR2_X1 U13583 ( .A(n13565), .B(n13566), .Z(n13563) );
  NOR2_X1 U13584 ( .A1(n13331), .A2(n13330), .ZN(n13562) );
  NAND2_X1 U13585 ( .A1(n13567), .A2(n13329), .ZN(n7485) );
  XOR2_X1 U13586 ( .A(n13568), .B(n13569), .Z(n13567) );
  NAND2_X1 U13587 ( .A1(n13570), .A2(n13334), .ZN(n7484) );
  INV_X1 U13588 ( .A(n13329), .ZN(n13334) );
  NAND2_X1 U13589 ( .A1(n13331), .A2(n13330), .ZN(n13329) );
  NAND2_X1 U13590 ( .A1(n13571), .A2(n13572), .ZN(n13330) );
  NAND2_X1 U13591 ( .A1(n13566), .A2(n13573), .ZN(n13572) );
  OR2_X1 U13592 ( .A1(n13565), .A2(n13564), .ZN(n13573) );
  NOR2_X1 U13593 ( .A1(n7849), .A2(n8307), .ZN(n13566) );
  NAND2_X1 U13594 ( .A1(n13564), .A2(n13565), .ZN(n13571) );
  NAND2_X1 U13595 ( .A1(n13574), .A2(n13575), .ZN(n13565) );
  NAND2_X1 U13596 ( .A1(n13576), .A2(a_1_), .ZN(n13575) );
  NOR2_X1 U13597 ( .A1(n13577), .A2(n7849), .ZN(n13576) );
  NOR2_X1 U13598 ( .A1(n13558), .A2(n13560), .ZN(n13577) );
  NAND2_X1 U13599 ( .A1(n13558), .A2(n13560), .ZN(n13574) );
  NAND2_X1 U13600 ( .A1(n13578), .A2(n13579), .ZN(n13560) );
  NAND2_X1 U13601 ( .A1(n13580), .A2(a_2_), .ZN(n13579) );
  NOR2_X1 U13602 ( .A1(n13581), .A2(n7849), .ZN(n13580) );
  NOR2_X1 U13603 ( .A1(n13554), .A2(n13556), .ZN(n13581) );
  NAND2_X1 U13604 ( .A1(n13554), .A2(n13556), .ZN(n13578) );
  NAND2_X1 U13605 ( .A1(n13582), .A2(n13583), .ZN(n13556) );
  NAND2_X1 U13606 ( .A1(n13584), .A2(a_3_), .ZN(n13583) );
  NOR2_X1 U13607 ( .A1(n13585), .A2(n7849), .ZN(n13584) );
  NOR2_X1 U13608 ( .A1(n13551), .A2(n13552), .ZN(n13585) );
  NAND2_X1 U13609 ( .A1(n13551), .A2(n13552), .ZN(n13582) );
  NAND2_X1 U13610 ( .A1(n13586), .A2(n13587), .ZN(n13552) );
  NAND2_X1 U13611 ( .A1(n13588), .A2(a_4_), .ZN(n13587) );
  NOR2_X1 U13612 ( .A1(n13589), .A2(n7849), .ZN(n13588) );
  NOR2_X1 U13613 ( .A1(n13547), .A2(n13548), .ZN(n13589) );
  NAND2_X1 U13614 ( .A1(n13547), .A2(n13548), .ZN(n13586) );
  NAND2_X1 U13615 ( .A1(n13590), .A2(n13591), .ZN(n13548) );
  NAND2_X1 U13616 ( .A1(n13592), .A2(a_5_), .ZN(n13591) );
  NOR2_X1 U13617 ( .A1(n13593), .A2(n7849), .ZN(n13592) );
  NOR2_X1 U13618 ( .A1(n13543), .A2(n13544), .ZN(n13593) );
  NAND2_X1 U13619 ( .A1(n13543), .A2(n13544), .ZN(n13590) );
  NAND2_X1 U13620 ( .A1(n13594), .A2(n13595), .ZN(n13544) );
  NAND2_X1 U13621 ( .A1(n13596), .A2(a_6_), .ZN(n13595) );
  NOR2_X1 U13622 ( .A1(n13597), .A2(n7849), .ZN(n13596) );
  NOR2_X1 U13623 ( .A1(n13540), .A2(n13539), .ZN(n13597) );
  NAND2_X1 U13624 ( .A1(n13539), .A2(n13540), .ZN(n13594) );
  NAND2_X1 U13625 ( .A1(n13598), .A2(n13599), .ZN(n13540) );
  NAND2_X1 U13626 ( .A1(n13600), .A2(a_7_), .ZN(n13599) );
  NOR2_X1 U13627 ( .A1(n13601), .A2(n7849), .ZN(n13600) );
  NOR2_X1 U13628 ( .A1(n13535), .A2(n13537), .ZN(n13601) );
  NAND2_X1 U13629 ( .A1(n13535), .A2(n13537), .ZN(n13598) );
  NAND2_X1 U13630 ( .A1(n13602), .A2(n13603), .ZN(n13537) );
  NAND2_X1 U13631 ( .A1(n13604), .A2(a_8_), .ZN(n13603) );
  NOR2_X1 U13632 ( .A1(n13605), .A2(n7849), .ZN(n13604) );
  NOR2_X1 U13633 ( .A1(n13531), .A2(n13533), .ZN(n13605) );
  NAND2_X1 U13634 ( .A1(n13531), .A2(n13533), .ZN(n13602) );
  NAND2_X1 U13635 ( .A1(n13606), .A2(n13607), .ZN(n13533) );
  NAND2_X1 U13636 ( .A1(n13528), .A2(n13608), .ZN(n13607) );
  OR2_X1 U13637 ( .A1(n13529), .A2(n7843), .ZN(n13608) );
  XNOR2_X1 U13638 ( .A(n13609), .B(n13610), .ZN(n13528) );
  XNOR2_X1 U13639 ( .A(n13611), .B(n13612), .ZN(n13610) );
  NAND2_X1 U13640 ( .A1(n7843), .A2(n13529), .ZN(n13606) );
  NAND2_X1 U13641 ( .A1(n13613), .A2(n13614), .ZN(n13529) );
  NAND2_X1 U13642 ( .A1(n13615), .A2(a_10_), .ZN(n13614) );
  NOR2_X1 U13643 ( .A1(n13616), .A2(n7849), .ZN(n13615) );
  NOR2_X1 U13644 ( .A1(n13368), .A2(n13369), .ZN(n13616) );
  NAND2_X1 U13645 ( .A1(n13368), .A2(n13369), .ZN(n13613) );
  NAND2_X1 U13646 ( .A1(n13617), .A2(n13618), .ZN(n13369) );
  NAND2_X1 U13647 ( .A1(n13619), .A2(b_9_), .ZN(n13618) );
  NOR2_X1 U13648 ( .A1(n13620), .A2(n7817), .ZN(n13619) );
  NOR2_X1 U13649 ( .A1(n13376), .A2(n13375), .ZN(n13620) );
  NAND2_X1 U13650 ( .A1(n13375), .A2(n13376), .ZN(n13617) );
  NAND2_X1 U13651 ( .A1(n13621), .A2(n13622), .ZN(n13376) );
  NAND2_X1 U13652 ( .A1(n13623), .A2(a_12_), .ZN(n13622) );
  NOR2_X1 U13653 ( .A1(n13624), .A2(n7849), .ZN(n13623) );
  NOR2_X1 U13654 ( .A1(n13382), .A2(n13384), .ZN(n13624) );
  NAND2_X1 U13655 ( .A1(n13382), .A2(n13384), .ZN(n13621) );
  NAND2_X1 U13656 ( .A1(n13625), .A2(n13626), .ZN(n13384) );
  NAND2_X1 U13657 ( .A1(n13627), .A2(a_13_), .ZN(n13626) );
  NOR2_X1 U13658 ( .A1(n13628), .A2(n7849), .ZN(n13627) );
  NOR2_X1 U13659 ( .A1(n13390), .A2(n13392), .ZN(n13628) );
  NAND2_X1 U13660 ( .A1(n13390), .A2(n13392), .ZN(n13625) );
  NAND2_X1 U13661 ( .A1(n13629), .A2(n13630), .ZN(n13392) );
  NAND2_X1 U13662 ( .A1(n13631), .A2(a_14_), .ZN(n13630) );
  NOR2_X1 U13663 ( .A1(n13632), .A2(n7849), .ZN(n13631) );
  NOR2_X1 U13664 ( .A1(n13400), .A2(n13398), .ZN(n13632) );
  NAND2_X1 U13665 ( .A1(n13398), .A2(n13400), .ZN(n13629) );
  NAND2_X1 U13666 ( .A1(n13633), .A2(n13634), .ZN(n13400) );
  NAND2_X1 U13667 ( .A1(n13635), .A2(a_15_), .ZN(n13634) );
  NOR2_X1 U13668 ( .A1(n13636), .A2(n7849), .ZN(n13635) );
  NOR2_X1 U13669 ( .A1(n13406), .A2(n13408), .ZN(n13636) );
  NAND2_X1 U13670 ( .A1(n13406), .A2(n13408), .ZN(n13633) );
  NAND2_X1 U13671 ( .A1(n13637), .A2(n13638), .ZN(n13408) );
  NAND2_X1 U13672 ( .A1(n13639), .A2(a_16_), .ZN(n13638) );
  NOR2_X1 U13673 ( .A1(n13640), .A2(n7849), .ZN(n13639) );
  NOR2_X1 U13674 ( .A1(n13416), .A2(n13414), .ZN(n13640) );
  NAND2_X1 U13675 ( .A1(n13414), .A2(n13416), .ZN(n13637) );
  NAND2_X1 U13676 ( .A1(n13641), .A2(n13642), .ZN(n13416) );
  NAND2_X1 U13677 ( .A1(n13643), .A2(a_17_), .ZN(n13642) );
  NOR2_X1 U13678 ( .A1(n13644), .A2(n7849), .ZN(n13643) );
  NOR2_X1 U13679 ( .A1(n13525), .A2(n13524), .ZN(n13644) );
  NAND2_X1 U13680 ( .A1(n13524), .A2(n13525), .ZN(n13641) );
  NAND2_X1 U13681 ( .A1(n13645), .A2(n13646), .ZN(n13525) );
  NAND2_X1 U13682 ( .A1(n13647), .A2(a_18_), .ZN(n13646) );
  NOR2_X1 U13683 ( .A1(n13648), .A2(n7849), .ZN(n13647) );
  NOR2_X1 U13684 ( .A1(n13519), .A2(n13521), .ZN(n13648) );
  NAND2_X1 U13685 ( .A1(n13519), .A2(n13521), .ZN(n13645) );
  NAND2_X1 U13686 ( .A1(n13517), .A2(n13649), .ZN(n13521) );
  NAND2_X1 U13687 ( .A1(n13516), .A2(n13518), .ZN(n13649) );
  NAND2_X1 U13688 ( .A1(n13650), .A2(n13651), .ZN(n13518) );
  NAND2_X1 U13689 ( .A1(a_19_), .A2(b_9_), .ZN(n13651) );
  INV_X1 U13690 ( .A(n13652), .ZN(n13650) );
  XNOR2_X1 U13691 ( .A(n13653), .B(n13654), .ZN(n13516) );
  NAND2_X1 U13692 ( .A1(n13655), .A2(n13656), .ZN(n13653) );
  NAND2_X1 U13693 ( .A1(a_19_), .A2(n13652), .ZN(n13517) );
  NAND2_X1 U13694 ( .A1(n13513), .A2(n13657), .ZN(n13652) );
  NAND2_X1 U13695 ( .A1(n13512), .A2(n13514), .ZN(n13657) );
  NAND2_X1 U13696 ( .A1(n13658), .A2(n13659), .ZN(n13514) );
  NAND2_X1 U13697 ( .A1(b_9_), .A2(a_20_), .ZN(n13659) );
  INV_X1 U13698 ( .A(n13660), .ZN(n13658) );
  XOR2_X1 U13699 ( .A(n13661), .B(n13662), .Z(n13512) );
  XNOR2_X1 U13700 ( .A(n13663), .B(n13664), .ZN(n13661) );
  NAND2_X1 U13701 ( .A1(b_8_), .A2(a_21_), .ZN(n13663) );
  NAND2_X1 U13702 ( .A1(a_20_), .A2(n13660), .ZN(n13513) );
  NAND2_X1 U13703 ( .A1(n13665), .A2(n13666), .ZN(n13660) );
  NAND2_X1 U13704 ( .A1(n13667), .A2(b_9_), .ZN(n13666) );
  NOR2_X1 U13705 ( .A1(n13668), .A2(n7656), .ZN(n13667) );
  NOR2_X1 U13706 ( .A1(n13509), .A2(n13508), .ZN(n13668) );
  NAND2_X1 U13707 ( .A1(n13508), .A2(n13509), .ZN(n13665) );
  NAND2_X1 U13708 ( .A1(n13669), .A2(n13670), .ZN(n13509) );
  NAND2_X1 U13709 ( .A1(n13506), .A2(n13671), .ZN(n13670) );
  NAND2_X1 U13710 ( .A1(n13505), .A2(n13504), .ZN(n13671) );
  NOR2_X1 U13711 ( .A1(n7645), .A2(n7849), .ZN(n13506) );
  OR2_X1 U13712 ( .A1(n13504), .A2(n13505), .ZN(n13669) );
  AND2_X1 U13713 ( .A1(n13672), .A2(n13673), .ZN(n13505) );
  NAND2_X1 U13714 ( .A1(n13502), .A2(n13674), .ZN(n13673) );
  OR2_X1 U13715 ( .A1(n13500), .A2(n13501), .ZN(n13674) );
  NOR2_X1 U13716 ( .A1(n7849), .A2(n7624), .ZN(n13502) );
  NAND2_X1 U13717 ( .A1(n13500), .A2(n13501), .ZN(n13672) );
  NAND2_X1 U13718 ( .A1(n13497), .A2(n13675), .ZN(n13501) );
  NAND2_X1 U13719 ( .A1(n13496), .A2(n13498), .ZN(n13675) );
  NAND2_X1 U13720 ( .A1(n13676), .A2(n13677), .ZN(n13498) );
  NAND2_X1 U13721 ( .A1(a_24_), .A2(b_9_), .ZN(n13677) );
  INV_X1 U13722 ( .A(n13678), .ZN(n13676) );
  XNOR2_X1 U13723 ( .A(n13679), .B(n13680), .ZN(n13496) );
  XOR2_X1 U13724 ( .A(n13681), .B(n13682), .Z(n13680) );
  NAND2_X1 U13725 ( .A1(a_25_), .A2(b_8_), .ZN(n13682) );
  NAND2_X1 U13726 ( .A1(a_24_), .A2(n13678), .ZN(n13497) );
  NAND2_X1 U13727 ( .A1(n13683), .A2(n13684), .ZN(n13678) );
  NAND2_X1 U13728 ( .A1(n13685), .A2(a_25_), .ZN(n13684) );
  NOR2_X1 U13729 ( .A1(n13686), .A2(n7849), .ZN(n13685) );
  NOR2_X1 U13730 ( .A1(n13449), .A2(n13451), .ZN(n13686) );
  NAND2_X1 U13731 ( .A1(n13449), .A2(n13451), .ZN(n13683) );
  NAND2_X1 U13732 ( .A1(n13687), .A2(n13688), .ZN(n13451) );
  NAND2_X1 U13733 ( .A1(n13689), .A2(a_26_), .ZN(n13688) );
  NOR2_X1 U13734 ( .A1(n13690), .A2(n7849), .ZN(n13689) );
  NOR2_X1 U13735 ( .A1(n13494), .A2(n13492), .ZN(n13690) );
  NAND2_X1 U13736 ( .A1(n13492), .A2(n13494), .ZN(n13687) );
  NAND2_X1 U13737 ( .A1(n13691), .A2(n13692), .ZN(n13494) );
  NAND2_X1 U13738 ( .A1(n13490), .A2(n13693), .ZN(n13692) );
  NAND2_X1 U13739 ( .A1(n13489), .A2(n13488), .ZN(n13693) );
  NOR2_X1 U13740 ( .A1(n7849), .A2(n7563), .ZN(n13490) );
  OR2_X1 U13741 ( .A1(n13488), .A2(n13489), .ZN(n13691) );
  AND2_X1 U13742 ( .A1(n13485), .A2(n13694), .ZN(n13489) );
  NAND2_X1 U13743 ( .A1(n13484), .A2(n13486), .ZN(n13694) );
  NAND2_X1 U13744 ( .A1(n13695), .A2(n13696), .ZN(n13486) );
  NAND2_X1 U13745 ( .A1(a_28_), .A2(b_9_), .ZN(n13696) );
  INV_X1 U13746 ( .A(n13697), .ZN(n13695) );
  XOR2_X1 U13747 ( .A(n13698), .B(n13699), .Z(n13484) );
  NOR2_X1 U13748 ( .A1(n7529), .A2(n8058), .ZN(n13699) );
  XOR2_X1 U13749 ( .A(n13700), .B(n13701), .Z(n13698) );
  NAND2_X1 U13750 ( .A1(a_28_), .A2(n13697), .ZN(n13485) );
  NAND2_X1 U13751 ( .A1(n13702), .A2(n13703), .ZN(n13697) );
  NAND2_X1 U13752 ( .A1(n13704), .A2(a_29_), .ZN(n13703) );
  NOR2_X1 U13753 ( .A1(n13705), .A2(n7849), .ZN(n13704) );
  NOR2_X1 U13754 ( .A1(n13470), .A2(n13471), .ZN(n13705) );
  NAND2_X1 U13755 ( .A1(n13470), .A2(n13471), .ZN(n13702) );
  NAND2_X1 U13756 ( .A1(n13706), .A2(n13707), .ZN(n13471) );
  NAND2_X1 U13757 ( .A1(n13708), .A2(b_7_), .ZN(n13707) );
  NOR2_X1 U13758 ( .A1(n13709), .A2(n8048), .ZN(n13708) );
  NOR2_X1 U13759 ( .A1(n8676), .A2(n8058), .ZN(n13709) );
  NAND2_X1 U13760 ( .A1(n13710), .A2(b_8_), .ZN(n13706) );
  NOR2_X1 U13761 ( .A1(n13711), .A2(n7515), .ZN(n13710) );
  NOR2_X1 U13762 ( .A1(n8679), .A2(n7885), .ZN(n13711) );
  AND2_X1 U13763 ( .A1(n13712), .A2(b_8_), .ZN(n13470) );
  NOR2_X1 U13764 ( .A1(n7849), .A2(n8451), .ZN(n13712) );
  XOR2_X1 U13765 ( .A(n13713), .B(n13714), .Z(n13488) );
  NAND2_X1 U13766 ( .A1(n13715), .A2(n13716), .ZN(n13713) );
  XNOR2_X1 U13767 ( .A(n13717), .B(n13718), .ZN(n13492) );
  XNOR2_X1 U13768 ( .A(n13719), .B(n13720), .ZN(n13717) );
  XOR2_X1 U13769 ( .A(n13721), .B(n13722), .Z(n13449) );
  XNOR2_X1 U13770 ( .A(n13723), .B(n13724), .ZN(n13721) );
  NAND2_X1 U13771 ( .A1(a_26_), .A2(b_8_), .ZN(n13723) );
  XNOR2_X1 U13772 ( .A(n13725), .B(n13726), .ZN(n13500) );
  NAND2_X1 U13773 ( .A1(n13727), .A2(n13728), .ZN(n13725) );
  XOR2_X1 U13774 ( .A(n13729), .B(n13730), .Z(n13504) );
  NAND2_X1 U13775 ( .A1(n13731), .A2(n13732), .ZN(n13729) );
  XNOR2_X1 U13776 ( .A(n13733), .B(n13734), .ZN(n13508) );
  XNOR2_X1 U13777 ( .A(n13735), .B(n13736), .ZN(n13734) );
  XNOR2_X1 U13778 ( .A(n13737), .B(n13738), .ZN(n13519) );
  XNOR2_X1 U13779 ( .A(n13739), .B(n13740), .ZN(n13738) );
  XOR2_X1 U13780 ( .A(n13741), .B(n13742), .Z(n13524) );
  XOR2_X1 U13781 ( .A(n13743), .B(n13744), .Z(n13741) );
  NOR2_X1 U13782 ( .A1(n8058), .A2(n7707), .ZN(n13744) );
  XNOR2_X1 U13783 ( .A(n13745), .B(n13746), .ZN(n13414) );
  NAND2_X1 U13784 ( .A1(n13747), .A2(n13748), .ZN(n13745) );
  XNOR2_X1 U13785 ( .A(n13749), .B(n13750), .ZN(n13406) );
  NAND2_X1 U13786 ( .A1(n13751), .A2(n13752), .ZN(n13749) );
  XNOR2_X1 U13787 ( .A(n13753), .B(n13754), .ZN(n13398) );
  NAND2_X1 U13788 ( .A1(n13755), .A2(n13756), .ZN(n13753) );
  XNOR2_X1 U13789 ( .A(n13757), .B(n13758), .ZN(n13390) );
  NAND2_X1 U13790 ( .A1(n13759), .A2(n13760), .ZN(n13757) );
  XNOR2_X1 U13791 ( .A(n13761), .B(n13762), .ZN(n13382) );
  XNOR2_X1 U13792 ( .A(n13763), .B(n13764), .ZN(n13762) );
  XNOR2_X1 U13793 ( .A(n13765), .B(n13766), .ZN(n13375) );
  XNOR2_X1 U13794 ( .A(n13767), .B(n13768), .ZN(n13765) );
  XNOR2_X1 U13795 ( .A(n13769), .B(n13770), .ZN(n13368) );
  XNOR2_X1 U13796 ( .A(n13771), .B(n13772), .ZN(n13770) );
  INV_X1 U13797 ( .A(n8004), .ZN(n7843) );
  NAND2_X1 U13798 ( .A1(a_9_), .A2(b_9_), .ZN(n8004) );
  XNOR2_X1 U13799 ( .A(n13773), .B(n13774), .ZN(n13531) );
  XNOR2_X1 U13800 ( .A(n13775), .B(n13776), .ZN(n13774) );
  XNOR2_X1 U13801 ( .A(n13777), .B(n13778), .ZN(n13535) );
  XOR2_X1 U13802 ( .A(n13779), .B(n13780), .Z(n13777) );
  XNOR2_X1 U13803 ( .A(n13781), .B(n13782), .ZN(n13539) );
  XNOR2_X1 U13804 ( .A(n13783), .B(n13784), .ZN(n13782) );
  XNOR2_X1 U13805 ( .A(n13785), .B(n13786), .ZN(n13543) );
  XNOR2_X1 U13806 ( .A(n13787), .B(n13788), .ZN(n13786) );
  XOR2_X1 U13807 ( .A(n13789), .B(n13790), .Z(n13547) );
  XOR2_X1 U13808 ( .A(n13791), .B(n13792), .Z(n13789) );
  NOR2_X1 U13809 ( .A1(n8058), .A2(n7914), .ZN(n13792) );
  XNOR2_X1 U13810 ( .A(n13793), .B(n13794), .ZN(n13551) );
  XOR2_X1 U13811 ( .A(n13795), .B(n13796), .Z(n13794) );
  NAND2_X1 U13812 ( .A1(a_4_), .A2(b_8_), .ZN(n13796) );
  XNOR2_X1 U13813 ( .A(n13797), .B(n13798), .ZN(n13554) );
  XOR2_X1 U13814 ( .A(n13799), .B(n13800), .Z(n13798) );
  NAND2_X1 U13815 ( .A1(a_3_), .A2(b_8_), .ZN(n13800) );
  XOR2_X1 U13816 ( .A(n13801), .B(n13802), .Z(n13558) );
  XOR2_X1 U13817 ( .A(n13803), .B(n13804), .Z(n13801) );
  NOR2_X1 U13818 ( .A1(n8058), .A2(n7965), .ZN(n13804) );
  XOR2_X1 U13819 ( .A(n13805), .B(n13806), .Z(n13564) );
  XOR2_X1 U13820 ( .A(n13807), .B(n13808), .Z(n13805) );
  NOR2_X1 U13821 ( .A1(n8058), .A2(n7973), .ZN(n13808) );
  XOR2_X1 U13822 ( .A(n13809), .B(n13810), .Z(n13331) );
  XOR2_X1 U13823 ( .A(n13811), .B(n13812), .Z(n13809) );
  XOR2_X1 U13824 ( .A(n13813), .B(n13569), .Z(n13570) );
  NAND2_X1 U13825 ( .A1(n13814), .A2(n13815), .ZN(n7490) );
  NAND2_X1 U13826 ( .A1(n13816), .A2(n13817), .ZN(n13815) );
  OR2_X1 U13827 ( .A1(n13818), .A2(n13819), .ZN(n13816) );
  NAND2_X1 U13828 ( .A1(n13569), .A2(n13813), .ZN(n13814) );
  INV_X1 U13829 ( .A(n13820), .ZN(n13569) );
  NAND2_X1 U13830 ( .A1(n13821), .A2(n13822), .ZN(n7489) );
  NOR2_X1 U13831 ( .A1(n13823), .A2(n13568), .ZN(n13822) );
  INV_X1 U13832 ( .A(n13813), .ZN(n13568) );
  NAND2_X1 U13833 ( .A1(n13824), .A2(n13825), .ZN(n13813) );
  NAND2_X1 U13834 ( .A1(n13812), .A2(n13826), .ZN(n13825) );
  OR2_X1 U13835 ( .A1(n13810), .A2(n13811), .ZN(n13826) );
  NOR2_X1 U13836 ( .A1(n8058), .A2(n8307), .ZN(n13812) );
  NAND2_X1 U13837 ( .A1(n13810), .A2(n13811), .ZN(n13824) );
  NAND2_X1 U13838 ( .A1(n13827), .A2(n13828), .ZN(n13811) );
  NAND2_X1 U13839 ( .A1(n13829), .A2(a_1_), .ZN(n13828) );
  NOR2_X1 U13840 ( .A1(n13830), .A2(n8058), .ZN(n13829) );
  NOR2_X1 U13841 ( .A1(n13807), .A2(n13806), .ZN(n13830) );
  NAND2_X1 U13842 ( .A1(n13806), .A2(n13807), .ZN(n13827) );
  NAND2_X1 U13843 ( .A1(n13831), .A2(n13832), .ZN(n13807) );
  NAND2_X1 U13844 ( .A1(n13833), .A2(a_2_), .ZN(n13832) );
  NOR2_X1 U13845 ( .A1(n13834), .A2(n8058), .ZN(n13833) );
  NOR2_X1 U13846 ( .A1(n13803), .A2(n13802), .ZN(n13834) );
  NAND2_X1 U13847 ( .A1(n13802), .A2(n13803), .ZN(n13831) );
  NAND2_X1 U13848 ( .A1(n13835), .A2(n13836), .ZN(n13803) );
  NAND2_X1 U13849 ( .A1(n13837), .A2(a_3_), .ZN(n13836) );
  NOR2_X1 U13850 ( .A1(n13838), .A2(n8058), .ZN(n13837) );
  NOR2_X1 U13851 ( .A1(n13799), .A2(n13797), .ZN(n13838) );
  NAND2_X1 U13852 ( .A1(n13797), .A2(n13799), .ZN(n13835) );
  NAND2_X1 U13853 ( .A1(n13839), .A2(n13840), .ZN(n13799) );
  NAND2_X1 U13854 ( .A1(n13841), .A2(a_4_), .ZN(n13840) );
  NOR2_X1 U13855 ( .A1(n13842), .A2(n8058), .ZN(n13841) );
  NOR2_X1 U13856 ( .A1(n13795), .A2(n13793), .ZN(n13842) );
  NAND2_X1 U13857 ( .A1(n13793), .A2(n13795), .ZN(n13839) );
  NAND2_X1 U13858 ( .A1(n13843), .A2(n13844), .ZN(n13795) );
  NAND2_X1 U13859 ( .A1(n13845), .A2(a_5_), .ZN(n13844) );
  NOR2_X1 U13860 ( .A1(n13846), .A2(n8058), .ZN(n13845) );
  NOR2_X1 U13861 ( .A1(n13791), .A2(n13790), .ZN(n13846) );
  NAND2_X1 U13862 ( .A1(n13790), .A2(n13791), .ZN(n13843) );
  NAND2_X1 U13863 ( .A1(n13847), .A2(n13848), .ZN(n13791) );
  NAND2_X1 U13864 ( .A1(n13788), .A2(n13849), .ZN(n13848) );
  OR2_X1 U13865 ( .A1(n13785), .A2(n13787), .ZN(n13849) );
  NOR2_X1 U13866 ( .A1(n8061), .A2(n8058), .ZN(n13788) );
  NAND2_X1 U13867 ( .A1(n13785), .A2(n13787), .ZN(n13847) );
  NAND2_X1 U13868 ( .A1(n13850), .A2(n13851), .ZN(n13787) );
  NAND2_X1 U13869 ( .A1(n13784), .A2(n13852), .ZN(n13851) );
  NAND2_X1 U13870 ( .A1(n13781), .A2(n13783), .ZN(n13852) );
  NOR2_X1 U13871 ( .A1(n7884), .A2(n8058), .ZN(n13784) );
  OR2_X1 U13872 ( .A1(n13783), .A2(n13781), .ZN(n13850) );
  XNOR2_X1 U13873 ( .A(n13853), .B(n13854), .ZN(n13781) );
  XOR2_X1 U13874 ( .A(n13855), .B(n13856), .Z(n13853) );
  NOR2_X1 U13875 ( .A1(n7885), .A2(n8059), .ZN(n13856) );
  NAND2_X1 U13876 ( .A1(n13857), .A2(n13858), .ZN(n13783) );
  NAND2_X1 U13877 ( .A1(n13778), .A2(n13859), .ZN(n13858) );
  NAND2_X1 U13878 ( .A1(n13780), .A2(n13779), .ZN(n13859) );
  XNOR2_X1 U13879 ( .A(n13860), .B(n13861), .ZN(n13778) );
  XOR2_X1 U13880 ( .A(n13862), .B(n13863), .Z(n13860) );
  NOR2_X1 U13881 ( .A1(n7885), .A2(n7848), .ZN(n13863) );
  OR2_X1 U13882 ( .A1(n13779), .A2(n13780), .ZN(n13857) );
  INV_X1 U13883 ( .A(n7863), .ZN(n13780) );
  NAND2_X1 U13884 ( .A1(a_8_), .A2(b_8_), .ZN(n7863) );
  NAND2_X1 U13885 ( .A1(n13864), .A2(n13865), .ZN(n13779) );
  NAND2_X1 U13886 ( .A1(n13776), .A2(n13866), .ZN(n13865) );
  OR2_X1 U13887 ( .A1(n13773), .A2(n13775), .ZN(n13866) );
  NOR2_X1 U13888 ( .A1(n7848), .A2(n8058), .ZN(n13776) );
  NAND2_X1 U13889 ( .A1(n13773), .A2(n13775), .ZN(n13864) );
  NAND2_X1 U13890 ( .A1(n13867), .A2(n13868), .ZN(n13775) );
  NAND2_X1 U13891 ( .A1(n13612), .A2(n13869), .ZN(n13868) );
  OR2_X1 U13892 ( .A1(n13609), .A2(n13611), .ZN(n13869) );
  NOR2_X1 U13893 ( .A1(n7837), .A2(n8058), .ZN(n13612) );
  NAND2_X1 U13894 ( .A1(n13609), .A2(n13611), .ZN(n13867) );
  NAND2_X1 U13895 ( .A1(n13870), .A2(n13871), .ZN(n13611) );
  NAND2_X1 U13896 ( .A1(n13772), .A2(n13872), .ZN(n13871) );
  OR2_X1 U13897 ( .A1(n13769), .A2(n13771), .ZN(n13872) );
  NOR2_X1 U13898 ( .A1(n8058), .A2(n7817), .ZN(n13772) );
  NAND2_X1 U13899 ( .A1(n13769), .A2(n13771), .ZN(n13870) );
  NAND2_X1 U13900 ( .A1(n13873), .A2(n13874), .ZN(n13771) );
  NAND2_X1 U13901 ( .A1(n13768), .A2(n13875), .ZN(n13874) );
  NAND2_X1 U13902 ( .A1(n13767), .A2(n13766), .ZN(n13875) );
  NOR2_X1 U13903 ( .A1(n7806), .A2(n8058), .ZN(n13768) );
  OR2_X1 U13904 ( .A1(n13766), .A2(n13767), .ZN(n13873) );
  AND2_X1 U13905 ( .A1(n13876), .A2(n13877), .ZN(n13767) );
  NAND2_X1 U13906 ( .A1(n13764), .A2(n13878), .ZN(n13877) );
  OR2_X1 U13907 ( .A1(n13761), .A2(n13763), .ZN(n13878) );
  NOR2_X1 U13908 ( .A1(n7786), .A2(n8058), .ZN(n13764) );
  NAND2_X1 U13909 ( .A1(n13761), .A2(n13763), .ZN(n13876) );
  NAND2_X1 U13910 ( .A1(n13759), .A2(n13879), .ZN(n13763) );
  NAND2_X1 U13911 ( .A1(n13758), .A2(n13760), .ZN(n13879) );
  NAND2_X1 U13912 ( .A1(n13880), .A2(n13881), .ZN(n13760) );
  NAND2_X1 U13913 ( .A1(a_14_), .A2(b_8_), .ZN(n13881) );
  INV_X1 U13914 ( .A(n13882), .ZN(n13880) );
  XOR2_X1 U13915 ( .A(n13883), .B(n13884), .Z(n13758) );
  XOR2_X1 U13916 ( .A(n13885), .B(n13886), .Z(n13883) );
  NOR2_X1 U13917 ( .A1(n7885), .A2(n7754), .ZN(n13886) );
  NAND2_X1 U13918 ( .A1(a_14_), .A2(n13882), .ZN(n13759) );
  NAND2_X1 U13919 ( .A1(n13755), .A2(n13887), .ZN(n13882) );
  NAND2_X1 U13920 ( .A1(n13754), .A2(n13756), .ZN(n13887) );
  NAND2_X1 U13921 ( .A1(n13888), .A2(n13889), .ZN(n13756) );
  NAND2_X1 U13922 ( .A1(a_15_), .A2(b_8_), .ZN(n13889) );
  INV_X1 U13923 ( .A(n13890), .ZN(n13888) );
  XNOR2_X1 U13924 ( .A(n13891), .B(n13892), .ZN(n13754) );
  XOR2_X1 U13925 ( .A(n13893), .B(n13894), .Z(n13892) );
  NAND2_X1 U13926 ( .A1(a_16_), .A2(b_7_), .ZN(n13894) );
  NAND2_X1 U13927 ( .A1(a_15_), .A2(n13890), .ZN(n13755) );
  NAND2_X1 U13928 ( .A1(n13751), .A2(n13895), .ZN(n13890) );
  NAND2_X1 U13929 ( .A1(n13750), .A2(n13752), .ZN(n13895) );
  NAND2_X1 U13930 ( .A1(n13896), .A2(n13897), .ZN(n13752) );
  NAND2_X1 U13931 ( .A1(a_16_), .A2(b_8_), .ZN(n13897) );
  INV_X1 U13932 ( .A(n13898), .ZN(n13896) );
  XNOR2_X1 U13933 ( .A(n13899), .B(n13900), .ZN(n13750) );
  XOR2_X1 U13934 ( .A(n13901), .B(n13902), .Z(n13900) );
  NAND2_X1 U13935 ( .A1(a_17_), .A2(b_7_), .ZN(n13902) );
  NAND2_X1 U13936 ( .A1(a_16_), .A2(n13898), .ZN(n13751) );
  NAND2_X1 U13937 ( .A1(n13747), .A2(n13903), .ZN(n13898) );
  NAND2_X1 U13938 ( .A1(n13746), .A2(n13748), .ZN(n13903) );
  NAND2_X1 U13939 ( .A1(n13904), .A2(n13905), .ZN(n13748) );
  NAND2_X1 U13940 ( .A1(a_17_), .A2(b_8_), .ZN(n13905) );
  INV_X1 U13941 ( .A(n13906), .ZN(n13904) );
  XOR2_X1 U13942 ( .A(n13907), .B(n13908), .Z(n13746) );
  XNOR2_X1 U13943 ( .A(n13909), .B(n13910), .ZN(n13907) );
  NAND2_X1 U13944 ( .A1(a_18_), .A2(b_7_), .ZN(n13909) );
  NAND2_X1 U13945 ( .A1(a_17_), .A2(n13906), .ZN(n13747) );
  NAND2_X1 U13946 ( .A1(n13911), .A2(n13912), .ZN(n13906) );
  NAND2_X1 U13947 ( .A1(n13913), .A2(a_18_), .ZN(n13912) );
  NOR2_X1 U13948 ( .A1(n13914), .A2(n8058), .ZN(n13913) );
  NOR2_X1 U13949 ( .A1(n13742), .A2(n13743), .ZN(n13914) );
  NAND2_X1 U13950 ( .A1(n13742), .A2(n13743), .ZN(n13911) );
  NAND2_X1 U13951 ( .A1(n13915), .A2(n13916), .ZN(n13743) );
  NAND2_X1 U13952 ( .A1(n13740), .A2(n13917), .ZN(n13916) );
  OR2_X1 U13953 ( .A1(n13737), .A2(n13739), .ZN(n13917) );
  NOR2_X1 U13954 ( .A1(n7687), .A2(n8058), .ZN(n13740) );
  NAND2_X1 U13955 ( .A1(n13737), .A2(n13739), .ZN(n13915) );
  NAND2_X1 U13956 ( .A1(n13655), .A2(n13918), .ZN(n13739) );
  NAND2_X1 U13957 ( .A1(n13654), .A2(n13656), .ZN(n13918) );
  NAND2_X1 U13958 ( .A1(n13919), .A2(n13920), .ZN(n13656) );
  NAND2_X1 U13959 ( .A1(b_8_), .A2(a_20_), .ZN(n13920) );
  INV_X1 U13960 ( .A(n13921), .ZN(n13919) );
  XOR2_X1 U13961 ( .A(n13922), .B(n13923), .Z(n13654) );
  XNOR2_X1 U13962 ( .A(n13924), .B(n13925), .ZN(n13922) );
  NAND2_X1 U13963 ( .A1(b_7_), .A2(a_21_), .ZN(n13924) );
  NAND2_X1 U13964 ( .A1(a_20_), .A2(n13921), .ZN(n13655) );
  NAND2_X1 U13965 ( .A1(n13926), .A2(n13927), .ZN(n13921) );
  NAND2_X1 U13966 ( .A1(n13928), .A2(b_8_), .ZN(n13927) );
  NOR2_X1 U13967 ( .A1(n13929), .A2(n7656), .ZN(n13928) );
  NOR2_X1 U13968 ( .A1(n13662), .A2(n13664), .ZN(n13929) );
  NAND2_X1 U13969 ( .A1(n13662), .A2(n13664), .ZN(n13926) );
  NAND2_X1 U13970 ( .A1(n13930), .A2(n13931), .ZN(n13664) );
  NAND2_X1 U13971 ( .A1(n13736), .A2(n13932), .ZN(n13931) );
  OR2_X1 U13972 ( .A1(n13735), .A2(n13733), .ZN(n13932) );
  NOR2_X1 U13973 ( .A1(n7645), .A2(n8058), .ZN(n13736) );
  NAND2_X1 U13974 ( .A1(n13733), .A2(n13735), .ZN(n13930) );
  NAND2_X1 U13975 ( .A1(n13731), .A2(n13933), .ZN(n13735) );
  NAND2_X1 U13976 ( .A1(n13730), .A2(n13732), .ZN(n13933) );
  NAND2_X1 U13977 ( .A1(n13934), .A2(n13935), .ZN(n13732) );
  NAND2_X1 U13978 ( .A1(b_8_), .A2(a_23_), .ZN(n13935) );
  INV_X1 U13979 ( .A(n13936), .ZN(n13934) );
  XNOR2_X1 U13980 ( .A(n13937), .B(n13938), .ZN(n13730) );
  NAND2_X1 U13981 ( .A1(n13939), .A2(n13940), .ZN(n13937) );
  NAND2_X1 U13982 ( .A1(a_23_), .A2(n13936), .ZN(n13731) );
  NAND2_X1 U13983 ( .A1(n13727), .A2(n13941), .ZN(n13936) );
  NAND2_X1 U13984 ( .A1(n13726), .A2(n13728), .ZN(n13941) );
  NAND2_X1 U13985 ( .A1(n13942), .A2(n13943), .ZN(n13728) );
  NAND2_X1 U13986 ( .A1(a_24_), .A2(b_8_), .ZN(n13943) );
  INV_X1 U13987 ( .A(n13944), .ZN(n13942) );
  XOR2_X1 U13988 ( .A(n13945), .B(n13946), .Z(n13726) );
  XOR2_X1 U13989 ( .A(n13947), .B(n13948), .Z(n13945) );
  NOR2_X1 U13990 ( .A1(n7885), .A2(n7593), .ZN(n13948) );
  NAND2_X1 U13991 ( .A1(a_24_), .A2(n13944), .ZN(n13727) );
  NAND2_X1 U13992 ( .A1(n13949), .A2(n13950), .ZN(n13944) );
  NAND2_X1 U13993 ( .A1(n13951), .A2(a_25_), .ZN(n13950) );
  NOR2_X1 U13994 ( .A1(n13952), .A2(n8058), .ZN(n13951) );
  NOR2_X1 U13995 ( .A1(n13679), .A2(n13681), .ZN(n13952) );
  NAND2_X1 U13996 ( .A1(n13679), .A2(n13681), .ZN(n13949) );
  NAND2_X1 U13997 ( .A1(n13953), .A2(n13954), .ZN(n13681) );
  NAND2_X1 U13998 ( .A1(n13955), .A2(a_26_), .ZN(n13954) );
  NOR2_X1 U13999 ( .A1(n13956), .A2(n8058), .ZN(n13955) );
  NOR2_X1 U14000 ( .A1(n13724), .A2(n13722), .ZN(n13956) );
  NAND2_X1 U14001 ( .A1(n13722), .A2(n13724), .ZN(n13953) );
  NAND2_X1 U14002 ( .A1(n13957), .A2(n13958), .ZN(n13724) );
  NAND2_X1 U14003 ( .A1(n13720), .A2(n13959), .ZN(n13958) );
  NAND2_X1 U14004 ( .A1(n13719), .A2(n13718), .ZN(n13959) );
  NOR2_X1 U14005 ( .A1(n8058), .A2(n7563), .ZN(n13720) );
  OR2_X1 U14006 ( .A1(n13718), .A2(n13719), .ZN(n13957) );
  AND2_X1 U14007 ( .A1(n13715), .A2(n13960), .ZN(n13719) );
  NAND2_X1 U14008 ( .A1(n13714), .A2(n13716), .ZN(n13960) );
  NAND2_X1 U14009 ( .A1(n13961), .A2(n13962), .ZN(n13716) );
  NAND2_X1 U14010 ( .A1(b_8_), .A2(a_28_), .ZN(n13962) );
  INV_X1 U14011 ( .A(n13963), .ZN(n13961) );
  XOR2_X1 U14012 ( .A(n13964), .B(n13965), .Z(n13714) );
  NOR2_X1 U14013 ( .A1(n7529), .A2(n7885), .ZN(n13965) );
  XOR2_X1 U14014 ( .A(n13966), .B(n13967), .Z(n13964) );
  NAND2_X1 U14015 ( .A1(a_28_), .A2(n13963), .ZN(n13715) );
  NAND2_X1 U14016 ( .A1(n13968), .A2(n13969), .ZN(n13963) );
  NAND2_X1 U14017 ( .A1(n13970), .A2(b_8_), .ZN(n13969) );
  NOR2_X1 U14018 ( .A1(n13971), .A2(n7529), .ZN(n13970) );
  NOR2_X1 U14019 ( .A1(n13700), .A2(n13701), .ZN(n13971) );
  NAND2_X1 U14020 ( .A1(n13700), .A2(n13701), .ZN(n13968) );
  NAND2_X1 U14021 ( .A1(n13972), .A2(n13973), .ZN(n13701) );
  NAND2_X1 U14022 ( .A1(n13974), .A2(b_6_), .ZN(n13973) );
  NOR2_X1 U14023 ( .A1(n13975), .A2(n8048), .ZN(n13974) );
  NOR2_X1 U14024 ( .A1(n8676), .A2(n7885), .ZN(n13975) );
  NAND2_X1 U14025 ( .A1(n13976), .A2(b_7_), .ZN(n13972) );
  NOR2_X1 U14026 ( .A1(n13977), .A2(n7515), .ZN(n13976) );
  NOR2_X1 U14027 ( .A1(n8679), .A2(n8060), .ZN(n13977) );
  AND2_X1 U14028 ( .A1(n13978), .A2(b_7_), .ZN(n13700) );
  NOR2_X1 U14029 ( .A1(n8451), .A2(n8058), .ZN(n13978) );
  XOR2_X1 U14030 ( .A(n13979), .B(n13980), .Z(n13718) );
  NAND2_X1 U14031 ( .A1(n13981), .A2(n13982), .ZN(n13979) );
  XNOR2_X1 U14032 ( .A(n13983), .B(n13984), .ZN(n13722) );
  XNOR2_X1 U14033 ( .A(n13985), .B(n13986), .ZN(n13983) );
  XOR2_X1 U14034 ( .A(n13987), .B(n13988), .Z(n13679) );
  XNOR2_X1 U14035 ( .A(n13989), .B(n13990), .ZN(n13987) );
  NAND2_X1 U14036 ( .A1(a_26_), .A2(b_7_), .ZN(n13989) );
  XNOR2_X1 U14037 ( .A(n13991), .B(n13992), .ZN(n13733) );
  NAND2_X1 U14038 ( .A1(n13993), .A2(n13994), .ZN(n13991) );
  XNOR2_X1 U14039 ( .A(n13995), .B(n13996), .ZN(n13662) );
  XOR2_X1 U14040 ( .A(n13997), .B(n13998), .Z(n13996) );
  NAND2_X1 U14041 ( .A1(a_22_), .A2(b_7_), .ZN(n13998) );
  XOR2_X1 U14042 ( .A(n13999), .B(n14000), .Z(n13737) );
  XOR2_X1 U14043 ( .A(n14001), .B(n14002), .Z(n13999) );
  NOR2_X1 U14044 ( .A1(n7676), .A2(n7885), .ZN(n14002) );
  XNOR2_X1 U14045 ( .A(n14003), .B(n14004), .ZN(n13742) );
  XOR2_X1 U14046 ( .A(n14005), .B(n14006), .Z(n14004) );
  NAND2_X1 U14047 ( .A1(a_19_), .A2(b_7_), .ZN(n14006) );
  XOR2_X1 U14048 ( .A(n14007), .B(n14008), .Z(n13761) );
  XOR2_X1 U14049 ( .A(n14009), .B(n14010), .Z(n14007) );
  NOR2_X1 U14050 ( .A1(n7885), .A2(n7775), .ZN(n14010) );
  XNOR2_X1 U14051 ( .A(n14011), .B(n14012), .ZN(n13766) );
  XOR2_X1 U14052 ( .A(n14013), .B(n14014), .Z(n14011) );
  NOR2_X1 U14053 ( .A1(n7885), .A2(n7786), .ZN(n14014) );
  XOR2_X1 U14054 ( .A(n14015), .B(n14016), .Z(n13769) );
  XOR2_X1 U14055 ( .A(n14017), .B(n14018), .Z(n14015) );
  NOR2_X1 U14056 ( .A1(n7885), .A2(n7806), .ZN(n14018) );
  XOR2_X1 U14057 ( .A(n14019), .B(n14020), .Z(n13609) );
  XOR2_X1 U14058 ( .A(n14021), .B(n14022), .Z(n14019) );
  NOR2_X1 U14059 ( .A1(n7817), .A2(n7885), .ZN(n14022) );
  XOR2_X1 U14060 ( .A(n14023), .B(n14024), .Z(n13773) );
  XOR2_X1 U14061 ( .A(n14025), .B(n14026), .Z(n14023) );
  NOR2_X1 U14062 ( .A1(n7885), .A2(n7837), .ZN(n14026) );
  XOR2_X1 U14063 ( .A(n14027), .B(n14028), .Z(n13785) );
  XOR2_X1 U14064 ( .A(n14029), .B(n7879), .Z(n14027) );
  XOR2_X1 U14065 ( .A(n14030), .B(n14031), .Z(n13790) );
  XNOR2_X1 U14066 ( .A(n14032), .B(n14033), .ZN(n14030) );
  NAND2_X1 U14067 ( .A1(a_6_), .A2(b_7_), .ZN(n14032) );
  XOR2_X1 U14068 ( .A(n14034), .B(n14035), .Z(n13793) );
  XNOR2_X1 U14069 ( .A(n14036), .B(n14037), .ZN(n14034) );
  NAND2_X1 U14070 ( .A1(a_5_), .A2(b_7_), .ZN(n14036) );
  XOR2_X1 U14071 ( .A(n14038), .B(n14039), .Z(n13797) );
  XOR2_X1 U14072 ( .A(n14040), .B(n14041), .Z(n14038) );
  NOR2_X1 U14073 ( .A1(n7885), .A2(n7934), .ZN(n14041) );
  XOR2_X1 U14074 ( .A(n14042), .B(n14043), .Z(n13802) );
  XOR2_X1 U14075 ( .A(n14044), .B(n14045), .Z(n14042) );
  NOR2_X1 U14076 ( .A1(n7885), .A2(n7945), .ZN(n14045) );
  XOR2_X1 U14077 ( .A(n14046), .B(n14047), .Z(n13806) );
  XOR2_X1 U14078 ( .A(n14048), .B(n14049), .Z(n14046) );
  NOR2_X1 U14079 ( .A1(n7885), .A2(n7965), .ZN(n14049) );
  XOR2_X1 U14080 ( .A(n14050), .B(n14051), .Z(n13810) );
  XOR2_X1 U14081 ( .A(n14052), .B(n14053), .Z(n14050) );
  NOR2_X1 U14082 ( .A1(n7885), .A2(n7973), .ZN(n14053) );
  NOR2_X1 U14083 ( .A1(n14054), .A2(n13820), .ZN(n13821) );
  XNOR2_X1 U14084 ( .A(n14055), .B(n14056), .ZN(n13820) );
  XOR2_X1 U14085 ( .A(n14057), .B(n14058), .Z(n14056) );
  NOR2_X1 U14086 ( .A1(n13819), .A2(n13818), .ZN(n14054) );
  NAND2_X1 U14087 ( .A1(n14059), .A2(n13817), .ZN(n7495) );
  XOR2_X1 U14088 ( .A(n14060), .B(n14061), .Z(n14059) );
  NAND2_X1 U14089 ( .A1(n14062), .A2(n13823), .ZN(n7494) );
  INV_X1 U14090 ( .A(n13817), .ZN(n13823) );
  NAND2_X1 U14091 ( .A1(n13819), .A2(n13818), .ZN(n13817) );
  NAND2_X1 U14092 ( .A1(n14063), .A2(n14064), .ZN(n13818) );
  NAND2_X1 U14093 ( .A1(n14058), .A2(n14065), .ZN(n14064) );
  NAND2_X1 U14094 ( .A1(n14057), .A2(n14055), .ZN(n14065) );
  NOR2_X1 U14095 ( .A1(n7885), .A2(n8307), .ZN(n14058) );
  OR2_X1 U14096 ( .A1(n14055), .A2(n14057), .ZN(n14063) );
  AND2_X1 U14097 ( .A1(n14066), .A2(n14067), .ZN(n14057) );
  NAND2_X1 U14098 ( .A1(n14068), .A2(a_1_), .ZN(n14067) );
  NOR2_X1 U14099 ( .A1(n14069), .A2(n7885), .ZN(n14068) );
  NOR2_X1 U14100 ( .A1(n14051), .A2(n14052), .ZN(n14069) );
  NAND2_X1 U14101 ( .A1(n14051), .A2(n14052), .ZN(n14066) );
  NAND2_X1 U14102 ( .A1(n14070), .A2(n14071), .ZN(n14052) );
  NAND2_X1 U14103 ( .A1(n14072), .A2(a_2_), .ZN(n14071) );
  NOR2_X1 U14104 ( .A1(n14073), .A2(n7885), .ZN(n14072) );
  NOR2_X1 U14105 ( .A1(n14047), .A2(n14048), .ZN(n14073) );
  NAND2_X1 U14106 ( .A1(n14047), .A2(n14048), .ZN(n14070) );
  NAND2_X1 U14107 ( .A1(n14074), .A2(n14075), .ZN(n14048) );
  NAND2_X1 U14108 ( .A1(n14076), .A2(a_3_), .ZN(n14075) );
  NOR2_X1 U14109 ( .A1(n14077), .A2(n7885), .ZN(n14076) );
  NOR2_X1 U14110 ( .A1(n14043), .A2(n14044), .ZN(n14077) );
  NAND2_X1 U14111 ( .A1(n14043), .A2(n14044), .ZN(n14074) );
  NAND2_X1 U14112 ( .A1(n14078), .A2(n14079), .ZN(n14044) );
  NAND2_X1 U14113 ( .A1(n14080), .A2(a_4_), .ZN(n14079) );
  NOR2_X1 U14114 ( .A1(n14081), .A2(n7885), .ZN(n14080) );
  NOR2_X1 U14115 ( .A1(n14039), .A2(n14040), .ZN(n14081) );
  NAND2_X1 U14116 ( .A1(n14039), .A2(n14040), .ZN(n14078) );
  NAND2_X1 U14117 ( .A1(n14082), .A2(n14083), .ZN(n14040) );
  NAND2_X1 U14118 ( .A1(n14084), .A2(a_5_), .ZN(n14083) );
  NOR2_X1 U14119 ( .A1(n14085), .A2(n7885), .ZN(n14084) );
  NOR2_X1 U14120 ( .A1(n14035), .A2(n14037), .ZN(n14085) );
  NAND2_X1 U14121 ( .A1(n14035), .A2(n14037), .ZN(n14082) );
  NAND2_X1 U14122 ( .A1(n14086), .A2(n14087), .ZN(n14037) );
  NAND2_X1 U14123 ( .A1(n14088), .A2(a_6_), .ZN(n14087) );
  NOR2_X1 U14124 ( .A1(n14089), .A2(n7885), .ZN(n14088) );
  NOR2_X1 U14125 ( .A1(n14031), .A2(n14033), .ZN(n14089) );
  NAND2_X1 U14126 ( .A1(n14031), .A2(n14033), .ZN(n14086) );
  NAND2_X1 U14127 ( .A1(n14090), .A2(n14091), .ZN(n14033) );
  NAND2_X1 U14128 ( .A1(n14028), .A2(n14092), .ZN(n14091) );
  OR2_X1 U14129 ( .A1(n14029), .A2(n7879), .ZN(n14092) );
  XOR2_X1 U14130 ( .A(n14093), .B(n14094), .Z(n14028) );
  XOR2_X1 U14131 ( .A(n14095), .B(n14096), .Z(n14093) );
  NOR2_X1 U14132 ( .A1(n8060), .A2(n8059), .ZN(n14096) );
  NAND2_X1 U14133 ( .A1(n7879), .A2(n14029), .ZN(n14090) );
  NAND2_X1 U14134 ( .A1(n14097), .A2(n14098), .ZN(n14029) );
  NAND2_X1 U14135 ( .A1(n14099), .A2(a_8_), .ZN(n14098) );
  NOR2_X1 U14136 ( .A1(n14100), .A2(n7885), .ZN(n14099) );
  NOR2_X1 U14137 ( .A1(n13854), .A2(n13855), .ZN(n14100) );
  NAND2_X1 U14138 ( .A1(n13854), .A2(n13855), .ZN(n14097) );
  NAND2_X1 U14139 ( .A1(n14101), .A2(n14102), .ZN(n13855) );
  NAND2_X1 U14140 ( .A1(n14103), .A2(a_9_), .ZN(n14102) );
  NOR2_X1 U14141 ( .A1(n14104), .A2(n7885), .ZN(n14103) );
  NOR2_X1 U14142 ( .A1(n13861), .A2(n13862), .ZN(n14104) );
  NAND2_X1 U14143 ( .A1(n13861), .A2(n13862), .ZN(n14101) );
  NAND2_X1 U14144 ( .A1(n14105), .A2(n14106), .ZN(n13862) );
  NAND2_X1 U14145 ( .A1(n14107), .A2(a_10_), .ZN(n14106) );
  NOR2_X1 U14146 ( .A1(n14108), .A2(n7885), .ZN(n14107) );
  NOR2_X1 U14147 ( .A1(n14024), .A2(n14025), .ZN(n14108) );
  NAND2_X1 U14148 ( .A1(n14024), .A2(n14025), .ZN(n14105) );
  NAND2_X1 U14149 ( .A1(n14109), .A2(n14110), .ZN(n14025) );
  NAND2_X1 U14150 ( .A1(n14111), .A2(b_7_), .ZN(n14110) );
  NOR2_X1 U14151 ( .A1(n14112), .A2(n7817), .ZN(n14111) );
  NOR2_X1 U14152 ( .A1(n14020), .A2(n14021), .ZN(n14112) );
  NAND2_X1 U14153 ( .A1(n14020), .A2(n14021), .ZN(n14109) );
  NAND2_X1 U14154 ( .A1(n14113), .A2(n14114), .ZN(n14021) );
  NAND2_X1 U14155 ( .A1(n14115), .A2(a_12_), .ZN(n14114) );
  NOR2_X1 U14156 ( .A1(n14116), .A2(n7885), .ZN(n14115) );
  NOR2_X1 U14157 ( .A1(n14016), .A2(n14017), .ZN(n14116) );
  NAND2_X1 U14158 ( .A1(n14016), .A2(n14017), .ZN(n14113) );
  NAND2_X1 U14159 ( .A1(n14117), .A2(n14118), .ZN(n14017) );
  NAND2_X1 U14160 ( .A1(n14119), .A2(a_13_), .ZN(n14118) );
  NOR2_X1 U14161 ( .A1(n14120), .A2(n7885), .ZN(n14119) );
  NOR2_X1 U14162 ( .A1(n14013), .A2(n14012), .ZN(n14120) );
  NAND2_X1 U14163 ( .A1(n14012), .A2(n14013), .ZN(n14117) );
  NAND2_X1 U14164 ( .A1(n14121), .A2(n14122), .ZN(n14013) );
  NAND2_X1 U14165 ( .A1(n14123), .A2(a_14_), .ZN(n14122) );
  NOR2_X1 U14166 ( .A1(n14124), .A2(n7885), .ZN(n14123) );
  NOR2_X1 U14167 ( .A1(n14008), .A2(n14009), .ZN(n14124) );
  NAND2_X1 U14168 ( .A1(n14008), .A2(n14009), .ZN(n14121) );
  NAND2_X1 U14169 ( .A1(n14125), .A2(n14126), .ZN(n14009) );
  NAND2_X1 U14170 ( .A1(n14127), .A2(a_15_), .ZN(n14126) );
  NOR2_X1 U14171 ( .A1(n14128), .A2(n7885), .ZN(n14127) );
  NOR2_X1 U14172 ( .A1(n13885), .A2(n13884), .ZN(n14128) );
  NAND2_X1 U14173 ( .A1(n13884), .A2(n13885), .ZN(n14125) );
  NAND2_X1 U14174 ( .A1(n14129), .A2(n14130), .ZN(n13885) );
  NAND2_X1 U14175 ( .A1(n14131), .A2(a_16_), .ZN(n14130) );
  NOR2_X1 U14176 ( .A1(n14132), .A2(n7885), .ZN(n14131) );
  NOR2_X1 U14177 ( .A1(n13891), .A2(n13893), .ZN(n14132) );
  NAND2_X1 U14178 ( .A1(n13891), .A2(n13893), .ZN(n14129) );
  NAND2_X1 U14179 ( .A1(n14133), .A2(n14134), .ZN(n13893) );
  NAND2_X1 U14180 ( .A1(n14135), .A2(a_17_), .ZN(n14134) );
  NOR2_X1 U14181 ( .A1(n14136), .A2(n7885), .ZN(n14135) );
  NOR2_X1 U14182 ( .A1(n13901), .A2(n13899), .ZN(n14136) );
  NAND2_X1 U14183 ( .A1(n13899), .A2(n13901), .ZN(n14133) );
  NAND2_X1 U14184 ( .A1(n14137), .A2(n14138), .ZN(n13901) );
  NAND2_X1 U14185 ( .A1(n14139), .A2(a_18_), .ZN(n14138) );
  NOR2_X1 U14186 ( .A1(n14140), .A2(n7885), .ZN(n14139) );
  NOR2_X1 U14187 ( .A1(n13908), .A2(n13910), .ZN(n14140) );
  NAND2_X1 U14188 ( .A1(n13908), .A2(n13910), .ZN(n14137) );
  NAND2_X1 U14189 ( .A1(n14141), .A2(n14142), .ZN(n13910) );
  NAND2_X1 U14190 ( .A1(n14143), .A2(a_19_), .ZN(n14142) );
  NOR2_X1 U14191 ( .A1(n14144), .A2(n7885), .ZN(n14143) );
  NOR2_X1 U14192 ( .A1(n14005), .A2(n14003), .ZN(n14144) );
  NAND2_X1 U14193 ( .A1(n14003), .A2(n14005), .ZN(n14141) );
  NAND2_X1 U14194 ( .A1(n14145), .A2(n14146), .ZN(n14005) );
  NAND2_X1 U14195 ( .A1(n14147), .A2(b_7_), .ZN(n14146) );
  NOR2_X1 U14196 ( .A1(n14148), .A2(n7676), .ZN(n14147) );
  NOR2_X1 U14197 ( .A1(n14000), .A2(n14001), .ZN(n14148) );
  NAND2_X1 U14198 ( .A1(n14000), .A2(n14001), .ZN(n14145) );
  NAND2_X1 U14199 ( .A1(n14149), .A2(n14150), .ZN(n14001) );
  NAND2_X1 U14200 ( .A1(n14151), .A2(b_7_), .ZN(n14150) );
  NOR2_X1 U14201 ( .A1(n14152), .A2(n7656), .ZN(n14151) );
  NOR2_X1 U14202 ( .A1(n13923), .A2(n13925), .ZN(n14152) );
  NAND2_X1 U14203 ( .A1(n13923), .A2(n13925), .ZN(n14149) );
  NAND2_X1 U14204 ( .A1(n14153), .A2(n14154), .ZN(n13925) );
  NAND2_X1 U14205 ( .A1(n14155), .A2(a_22_), .ZN(n14154) );
  NOR2_X1 U14206 ( .A1(n14156), .A2(n7885), .ZN(n14155) );
  NOR2_X1 U14207 ( .A1(n13997), .A2(n13995), .ZN(n14156) );
  NAND2_X1 U14208 ( .A1(n13995), .A2(n13997), .ZN(n14153) );
  NAND2_X1 U14209 ( .A1(n13993), .A2(n14157), .ZN(n13997) );
  NAND2_X1 U14210 ( .A1(n13992), .A2(n13994), .ZN(n14157) );
  NAND2_X1 U14211 ( .A1(n14158), .A2(n14159), .ZN(n13994) );
  NAND2_X1 U14212 ( .A1(b_7_), .A2(a_23_), .ZN(n14159) );
  INV_X1 U14213 ( .A(n14160), .ZN(n14158) );
  XNOR2_X1 U14214 ( .A(n14161), .B(n14162), .ZN(n13992) );
  NAND2_X1 U14215 ( .A1(n14163), .A2(n14164), .ZN(n14161) );
  NAND2_X1 U14216 ( .A1(a_23_), .A2(n14160), .ZN(n13993) );
  NAND2_X1 U14217 ( .A1(n13939), .A2(n14165), .ZN(n14160) );
  NAND2_X1 U14218 ( .A1(n13938), .A2(n13940), .ZN(n14165) );
  NAND2_X1 U14219 ( .A1(n14166), .A2(n14167), .ZN(n13940) );
  NAND2_X1 U14220 ( .A1(a_24_), .A2(b_7_), .ZN(n14167) );
  INV_X1 U14221 ( .A(n14168), .ZN(n14166) );
  XNOR2_X1 U14222 ( .A(n14169), .B(n14170), .ZN(n13938) );
  XOR2_X1 U14223 ( .A(n14171), .B(n14172), .Z(n14170) );
  NAND2_X1 U14224 ( .A1(a_25_), .A2(b_6_), .ZN(n14172) );
  NAND2_X1 U14225 ( .A1(a_24_), .A2(n14168), .ZN(n13939) );
  NAND2_X1 U14226 ( .A1(n14173), .A2(n14174), .ZN(n14168) );
  NAND2_X1 U14227 ( .A1(n14175), .A2(a_25_), .ZN(n14174) );
  NOR2_X1 U14228 ( .A1(n14176), .A2(n7885), .ZN(n14175) );
  NOR2_X1 U14229 ( .A1(n13946), .A2(n13947), .ZN(n14176) );
  NAND2_X1 U14230 ( .A1(n13946), .A2(n13947), .ZN(n14173) );
  NAND2_X1 U14231 ( .A1(n14177), .A2(n14178), .ZN(n13947) );
  NAND2_X1 U14232 ( .A1(n14179), .A2(a_26_), .ZN(n14178) );
  NOR2_X1 U14233 ( .A1(n14180), .A2(n7885), .ZN(n14179) );
  NOR2_X1 U14234 ( .A1(n13990), .A2(n13988), .ZN(n14180) );
  NAND2_X1 U14235 ( .A1(n13988), .A2(n13990), .ZN(n14177) );
  NAND2_X1 U14236 ( .A1(n14181), .A2(n14182), .ZN(n13990) );
  NAND2_X1 U14237 ( .A1(n13986), .A2(n14183), .ZN(n14182) );
  NAND2_X1 U14238 ( .A1(n13985), .A2(n13984), .ZN(n14183) );
  NOR2_X1 U14239 ( .A1(n7885), .A2(n7563), .ZN(n13986) );
  OR2_X1 U14240 ( .A1(n13984), .A2(n13985), .ZN(n14181) );
  AND2_X1 U14241 ( .A1(n13981), .A2(n14184), .ZN(n13985) );
  NAND2_X1 U14242 ( .A1(n13980), .A2(n13982), .ZN(n14184) );
  NAND2_X1 U14243 ( .A1(n14185), .A2(n14186), .ZN(n13982) );
  NAND2_X1 U14244 ( .A1(b_7_), .A2(a_28_), .ZN(n14186) );
  INV_X1 U14245 ( .A(n14187), .ZN(n14185) );
  XOR2_X1 U14246 ( .A(n14188), .B(n14189), .Z(n13980) );
  NOR2_X1 U14247 ( .A1(n7529), .A2(n8060), .ZN(n14189) );
  XOR2_X1 U14248 ( .A(n14190), .B(n14191), .Z(n14188) );
  NAND2_X1 U14249 ( .A1(a_28_), .A2(n14187), .ZN(n13981) );
  NAND2_X1 U14250 ( .A1(n14192), .A2(n14193), .ZN(n14187) );
  NAND2_X1 U14251 ( .A1(n14194), .A2(b_7_), .ZN(n14193) );
  NOR2_X1 U14252 ( .A1(n14195), .A2(n7529), .ZN(n14194) );
  NOR2_X1 U14253 ( .A1(n13966), .A2(n13967), .ZN(n14195) );
  NAND2_X1 U14254 ( .A1(n13966), .A2(n13967), .ZN(n14192) );
  NAND2_X1 U14255 ( .A1(n14196), .A2(n14197), .ZN(n13967) );
  NAND2_X1 U14256 ( .A1(n14198), .A2(b_5_), .ZN(n14197) );
  NOR2_X1 U14257 ( .A1(n14199), .A2(n8048), .ZN(n14198) );
  NOR2_X1 U14258 ( .A1(n8676), .A2(n8060), .ZN(n14199) );
  NAND2_X1 U14259 ( .A1(n14200), .A2(b_6_), .ZN(n14196) );
  NOR2_X1 U14260 ( .A1(n14201), .A2(n7515), .ZN(n14200) );
  NOR2_X1 U14261 ( .A1(n8679), .A2(n7915), .ZN(n14201) );
  AND2_X1 U14262 ( .A1(n14202), .A2(b_6_), .ZN(n13966) );
  NOR2_X1 U14263 ( .A1(n8451), .A2(n7885), .ZN(n14202) );
  XOR2_X1 U14264 ( .A(n14203), .B(n14204), .Z(n13984) );
  NAND2_X1 U14265 ( .A1(n14205), .A2(n14206), .ZN(n14203) );
  XNOR2_X1 U14266 ( .A(n14207), .B(n14208), .ZN(n13988) );
  XNOR2_X1 U14267 ( .A(n14209), .B(n14210), .ZN(n14207) );
  XOR2_X1 U14268 ( .A(n14211), .B(n14212), .Z(n13946) );
  XNOR2_X1 U14269 ( .A(n14213), .B(n14214), .ZN(n14211) );
  NAND2_X1 U14270 ( .A1(a_26_), .A2(b_6_), .ZN(n14213) );
  XNOR2_X1 U14271 ( .A(n14215), .B(n14216), .ZN(n13995) );
  XNOR2_X1 U14272 ( .A(n14217), .B(n14218), .ZN(n14215) );
  XOR2_X1 U14273 ( .A(n14219), .B(n14220), .Z(n13923) );
  XOR2_X1 U14274 ( .A(n14221), .B(n14222), .Z(n14219) );
  NOR2_X1 U14275 ( .A1(n8060), .A2(n7645), .ZN(n14222) );
  XNOR2_X1 U14276 ( .A(n14223), .B(n14224), .ZN(n14000) );
  XNOR2_X1 U14277 ( .A(n14225), .B(n14226), .ZN(n14224) );
  XOR2_X1 U14278 ( .A(n14227), .B(n14228), .Z(n14003) );
  XOR2_X1 U14279 ( .A(n14229), .B(n14230), .Z(n14227) );
  NOR2_X1 U14280 ( .A1(n7676), .A2(n8060), .ZN(n14230) );
  XNOR2_X1 U14281 ( .A(n14231), .B(n14232), .ZN(n13908) );
  XNOR2_X1 U14282 ( .A(n14233), .B(n14234), .ZN(n14232) );
  XNOR2_X1 U14283 ( .A(n14235), .B(n14236), .ZN(n13899) );
  XNOR2_X1 U14284 ( .A(n14237), .B(n14238), .ZN(n14235) );
  XNOR2_X1 U14285 ( .A(n14239), .B(n14240), .ZN(n13891) );
  XNOR2_X1 U14286 ( .A(n14241), .B(n14242), .ZN(n14240) );
  XNOR2_X1 U14287 ( .A(n14243), .B(n14244), .ZN(n13884) );
  XNOR2_X1 U14288 ( .A(n14245), .B(n14246), .ZN(n14244) );
  XNOR2_X1 U14289 ( .A(n14247), .B(n14248), .ZN(n14008) );
  XNOR2_X1 U14290 ( .A(n14249), .B(n14250), .ZN(n14248) );
  XNOR2_X1 U14291 ( .A(n14251), .B(n14252), .ZN(n14012) );
  XNOR2_X1 U14292 ( .A(n14253), .B(n14254), .ZN(n14252) );
  XNOR2_X1 U14293 ( .A(n14255), .B(n14256), .ZN(n14016) );
  XNOR2_X1 U14294 ( .A(n14257), .B(n14258), .ZN(n14256) );
  XNOR2_X1 U14295 ( .A(n14259), .B(n14260), .ZN(n14020) );
  XNOR2_X1 U14296 ( .A(n14261), .B(n14262), .ZN(n14260) );
  XOR2_X1 U14297 ( .A(n14263), .B(n14264), .Z(n14024) );
  XOR2_X1 U14298 ( .A(n14265), .B(n14266), .Z(n14263) );
  XOR2_X1 U14299 ( .A(n14267), .B(n14268), .Z(n13861) );
  XOR2_X1 U14300 ( .A(n14269), .B(n14270), .Z(n14267) );
  XOR2_X1 U14301 ( .A(n14271), .B(n14272), .Z(n13854) );
  XOR2_X1 U14302 ( .A(n14273), .B(n14274), .Z(n14271) );
  NOR2_X1 U14303 ( .A1(n8060), .A2(n7848), .ZN(n14274) );
  INV_X1 U14304 ( .A(n8000), .ZN(n7879) );
  NAND2_X1 U14305 ( .A1(a_7_), .A2(b_7_), .ZN(n8000) );
  XOR2_X1 U14306 ( .A(n14275), .B(n14276), .Z(n14031) );
  XOR2_X1 U14307 ( .A(n14277), .B(n14278), .Z(n14275) );
  NOR2_X1 U14308 ( .A1(n8060), .A2(n7884), .ZN(n14278) );
  XOR2_X1 U14309 ( .A(n14279), .B(n14280), .Z(n14035) );
  XOR2_X1 U14310 ( .A(n14281), .B(n14282), .Z(n14279) );
  XOR2_X1 U14311 ( .A(n14283), .B(n14284), .Z(n14039) );
  XOR2_X1 U14312 ( .A(n14285), .B(n14286), .Z(n14283) );
  NOR2_X1 U14313 ( .A1(n8060), .A2(n7914), .ZN(n14286) );
  XOR2_X1 U14314 ( .A(n14287), .B(n14288), .Z(n14043) );
  XOR2_X1 U14315 ( .A(n14289), .B(n14290), .Z(n14287) );
  NOR2_X1 U14316 ( .A1(n8060), .A2(n7934), .ZN(n14290) );
  XOR2_X1 U14317 ( .A(n14291), .B(n14292), .Z(n14047) );
  XOR2_X1 U14318 ( .A(n14293), .B(n14294), .Z(n14291) );
  NOR2_X1 U14319 ( .A1(n8060), .A2(n7945), .ZN(n14294) );
  XNOR2_X1 U14320 ( .A(n14295), .B(n14296), .ZN(n14051) );
  XOR2_X1 U14321 ( .A(n14297), .B(n14298), .Z(n14296) );
  NAND2_X1 U14322 ( .A1(a_2_), .A2(b_6_), .ZN(n14298) );
  XOR2_X1 U14323 ( .A(n14299), .B(n14300), .Z(n14055) );
  XOR2_X1 U14324 ( .A(n14301), .B(n14302), .Z(n14300) );
  NAND2_X1 U14325 ( .A1(a_1_), .A2(b_6_), .ZN(n14302) );
  XOR2_X1 U14326 ( .A(n14303), .B(n14304), .Z(n13819) );
  XOR2_X1 U14327 ( .A(n14305), .B(n14306), .Z(n14303) );
  XOR2_X1 U14328 ( .A(n14061), .B(n14307), .Z(n14062) );
  NAND2_X1 U14329 ( .A1(n14308), .A2(n14309), .ZN(n7552) );
  NAND2_X1 U14330 ( .A1(n14310), .A2(n14311), .ZN(n14309) );
  NAND2_X1 U14331 ( .A1(n14312), .A2(n14313), .ZN(n14310) );
  OR2_X1 U14332 ( .A1(n14061), .A2(n14307), .ZN(n14308) );
  NAND2_X1 U14333 ( .A1(n14314), .A2(n14315), .ZN(n7551) );
  NOR2_X1 U14334 ( .A1(n14316), .A2(n14307), .ZN(n14315) );
  INV_X1 U14335 ( .A(n14060), .ZN(n14307) );
  NAND2_X1 U14336 ( .A1(n14317), .A2(n14318), .ZN(n14060) );
  NAND2_X1 U14337 ( .A1(n14306), .A2(n14319), .ZN(n14318) );
  OR2_X1 U14338 ( .A1(n14304), .A2(n14305), .ZN(n14319) );
  NOR2_X1 U14339 ( .A1(n8060), .A2(n8307), .ZN(n14306) );
  NAND2_X1 U14340 ( .A1(n14304), .A2(n14305), .ZN(n14317) );
  NAND2_X1 U14341 ( .A1(n14320), .A2(n14321), .ZN(n14305) );
  NAND2_X1 U14342 ( .A1(n14322), .A2(a_1_), .ZN(n14321) );
  NOR2_X1 U14343 ( .A1(n14323), .A2(n8060), .ZN(n14322) );
  NOR2_X1 U14344 ( .A1(n14301), .A2(n14299), .ZN(n14323) );
  NAND2_X1 U14345 ( .A1(n14299), .A2(n14301), .ZN(n14320) );
  NAND2_X1 U14346 ( .A1(n14324), .A2(n14325), .ZN(n14301) );
  NAND2_X1 U14347 ( .A1(n14326), .A2(a_2_), .ZN(n14325) );
  NOR2_X1 U14348 ( .A1(n14327), .A2(n8060), .ZN(n14326) );
  NOR2_X1 U14349 ( .A1(n14297), .A2(n14295), .ZN(n14327) );
  NAND2_X1 U14350 ( .A1(n14295), .A2(n14297), .ZN(n14324) );
  NAND2_X1 U14351 ( .A1(n14328), .A2(n14329), .ZN(n14297) );
  NAND2_X1 U14352 ( .A1(n14330), .A2(a_3_), .ZN(n14329) );
  NOR2_X1 U14353 ( .A1(n14331), .A2(n8060), .ZN(n14330) );
  NOR2_X1 U14354 ( .A1(n14293), .A2(n14292), .ZN(n14331) );
  NAND2_X1 U14355 ( .A1(n14292), .A2(n14293), .ZN(n14328) );
  NAND2_X1 U14356 ( .A1(n14332), .A2(n14333), .ZN(n14293) );
  NAND2_X1 U14357 ( .A1(n14334), .A2(a_4_), .ZN(n14333) );
  NOR2_X1 U14358 ( .A1(n14335), .A2(n8060), .ZN(n14334) );
  NOR2_X1 U14359 ( .A1(n14289), .A2(n14288), .ZN(n14335) );
  NAND2_X1 U14360 ( .A1(n14288), .A2(n14289), .ZN(n14332) );
  NAND2_X1 U14361 ( .A1(n14336), .A2(n14337), .ZN(n14289) );
  NAND2_X1 U14362 ( .A1(n14338), .A2(a_5_), .ZN(n14337) );
  NOR2_X1 U14363 ( .A1(n14339), .A2(n8060), .ZN(n14338) );
  NOR2_X1 U14364 ( .A1(n14285), .A2(n14284), .ZN(n14339) );
  NAND2_X1 U14365 ( .A1(n14284), .A2(n14285), .ZN(n14336) );
  NAND2_X1 U14366 ( .A1(n14340), .A2(n14341), .ZN(n14285) );
  NAND2_X1 U14367 ( .A1(n14280), .A2(n14342), .ZN(n14341) );
  OR2_X1 U14368 ( .A1(n14281), .A2(n14282), .ZN(n14342) );
  XOR2_X1 U14369 ( .A(n14343), .B(n14344), .Z(n14280) );
  XOR2_X1 U14370 ( .A(n14345), .B(n14346), .Z(n14343) );
  NOR2_X1 U14371 ( .A1(n7915), .A2(n7884), .ZN(n14346) );
  NAND2_X1 U14372 ( .A1(n14282), .A2(n14281), .ZN(n14340) );
  NAND2_X1 U14373 ( .A1(n14347), .A2(n14348), .ZN(n14281) );
  NAND2_X1 U14374 ( .A1(n14349), .A2(a_7_), .ZN(n14348) );
  NOR2_X1 U14375 ( .A1(n14350), .A2(n8060), .ZN(n14349) );
  NOR2_X1 U14376 ( .A1(n14277), .A2(n14276), .ZN(n14350) );
  NAND2_X1 U14377 ( .A1(n14276), .A2(n14277), .ZN(n14347) );
  NAND2_X1 U14378 ( .A1(n14351), .A2(n14352), .ZN(n14277) );
  NAND2_X1 U14379 ( .A1(n14353), .A2(a_8_), .ZN(n14352) );
  NOR2_X1 U14380 ( .A1(n14354), .A2(n8060), .ZN(n14353) );
  NOR2_X1 U14381 ( .A1(n14095), .A2(n14094), .ZN(n14354) );
  NAND2_X1 U14382 ( .A1(n14094), .A2(n14095), .ZN(n14351) );
  NAND2_X1 U14383 ( .A1(n14355), .A2(n14356), .ZN(n14095) );
  NAND2_X1 U14384 ( .A1(n14357), .A2(a_9_), .ZN(n14356) );
  NOR2_X1 U14385 ( .A1(n14358), .A2(n8060), .ZN(n14357) );
  NOR2_X1 U14386 ( .A1(n14273), .A2(n14272), .ZN(n14358) );
  NAND2_X1 U14387 ( .A1(n14272), .A2(n14273), .ZN(n14355) );
  NAND2_X1 U14388 ( .A1(n14359), .A2(n14360), .ZN(n14273) );
  NAND2_X1 U14389 ( .A1(n14270), .A2(n14361), .ZN(n14360) );
  OR2_X1 U14390 ( .A1(n14268), .A2(n14269), .ZN(n14361) );
  NOR2_X1 U14391 ( .A1(n7837), .A2(n8060), .ZN(n14270) );
  NAND2_X1 U14392 ( .A1(n14268), .A2(n14269), .ZN(n14359) );
  NAND2_X1 U14393 ( .A1(n14362), .A2(n14363), .ZN(n14269) );
  NAND2_X1 U14394 ( .A1(n14266), .A2(n14364), .ZN(n14363) );
  OR2_X1 U14395 ( .A1(n14264), .A2(n14265), .ZN(n14364) );
  NOR2_X1 U14396 ( .A1(n8060), .A2(n7817), .ZN(n14266) );
  NAND2_X1 U14397 ( .A1(n14264), .A2(n14265), .ZN(n14362) );
  NAND2_X1 U14398 ( .A1(n14365), .A2(n14366), .ZN(n14265) );
  NAND2_X1 U14399 ( .A1(n14262), .A2(n14367), .ZN(n14366) );
  OR2_X1 U14400 ( .A1(n14259), .A2(n14261), .ZN(n14367) );
  NOR2_X1 U14401 ( .A1(n7806), .A2(n8060), .ZN(n14262) );
  NAND2_X1 U14402 ( .A1(n14259), .A2(n14261), .ZN(n14365) );
  NAND2_X1 U14403 ( .A1(n14368), .A2(n14369), .ZN(n14261) );
  NAND2_X1 U14404 ( .A1(n14258), .A2(n14370), .ZN(n14369) );
  OR2_X1 U14405 ( .A1(n14255), .A2(n14257), .ZN(n14370) );
  NOR2_X1 U14406 ( .A1(n7786), .A2(n8060), .ZN(n14258) );
  NAND2_X1 U14407 ( .A1(n14255), .A2(n14257), .ZN(n14368) );
  NAND2_X1 U14408 ( .A1(n14371), .A2(n14372), .ZN(n14257) );
  NAND2_X1 U14409 ( .A1(n14254), .A2(n14373), .ZN(n14372) );
  OR2_X1 U14410 ( .A1(n14253), .A2(n14251), .ZN(n14373) );
  NOR2_X1 U14411 ( .A1(n7775), .A2(n8060), .ZN(n14254) );
  NAND2_X1 U14412 ( .A1(n14251), .A2(n14253), .ZN(n14371) );
  NAND2_X1 U14413 ( .A1(n14374), .A2(n14375), .ZN(n14253) );
  NAND2_X1 U14414 ( .A1(n14250), .A2(n14376), .ZN(n14375) );
  OR2_X1 U14415 ( .A1(n14247), .A2(n14249), .ZN(n14376) );
  NOR2_X1 U14416 ( .A1(n7754), .A2(n8060), .ZN(n14250) );
  NAND2_X1 U14417 ( .A1(n14247), .A2(n14249), .ZN(n14374) );
  NAND2_X1 U14418 ( .A1(n14377), .A2(n14378), .ZN(n14249) );
  NAND2_X1 U14419 ( .A1(n14246), .A2(n14379), .ZN(n14378) );
  OR2_X1 U14420 ( .A1(n14245), .A2(n14243), .ZN(n14379) );
  NOR2_X1 U14421 ( .A1(n7743), .A2(n8060), .ZN(n14246) );
  NAND2_X1 U14422 ( .A1(n14243), .A2(n14245), .ZN(n14377) );
  NAND2_X1 U14423 ( .A1(n14380), .A2(n14381), .ZN(n14245) );
  NAND2_X1 U14424 ( .A1(n14242), .A2(n14382), .ZN(n14381) );
  OR2_X1 U14425 ( .A1(n14239), .A2(n14241), .ZN(n14382) );
  NOR2_X1 U14426 ( .A1(n7723), .A2(n8060), .ZN(n14242) );
  NAND2_X1 U14427 ( .A1(n14239), .A2(n14241), .ZN(n14380) );
  NAND2_X1 U14428 ( .A1(n14383), .A2(n14384), .ZN(n14241) );
  NAND2_X1 U14429 ( .A1(n14238), .A2(n14385), .ZN(n14384) );
  NAND2_X1 U14430 ( .A1(n14237), .A2(n14236), .ZN(n14385) );
  NOR2_X1 U14431 ( .A1(n7707), .A2(n8060), .ZN(n14238) );
  OR2_X1 U14432 ( .A1(n14236), .A2(n14237), .ZN(n14383) );
  AND2_X1 U14433 ( .A1(n14386), .A2(n14387), .ZN(n14237) );
  NAND2_X1 U14434 ( .A1(n14234), .A2(n14388), .ZN(n14387) );
  OR2_X1 U14435 ( .A1(n14231), .A2(n14233), .ZN(n14388) );
  NOR2_X1 U14436 ( .A1(n7687), .A2(n8060), .ZN(n14234) );
  NAND2_X1 U14437 ( .A1(n14231), .A2(n14233), .ZN(n14386) );
  NAND2_X1 U14438 ( .A1(n14389), .A2(n14390), .ZN(n14233) );
  NAND2_X1 U14439 ( .A1(n14391), .A2(b_6_), .ZN(n14390) );
  NOR2_X1 U14440 ( .A1(n14392), .A2(n7676), .ZN(n14391) );
  NOR2_X1 U14441 ( .A1(n14228), .A2(n14229), .ZN(n14392) );
  NAND2_X1 U14442 ( .A1(n14228), .A2(n14229), .ZN(n14389) );
  NAND2_X1 U14443 ( .A1(n14393), .A2(n14394), .ZN(n14229) );
  NAND2_X1 U14444 ( .A1(n14226), .A2(n14395), .ZN(n14394) );
  OR2_X1 U14445 ( .A1(n14223), .A2(n14225), .ZN(n14395) );
  NOR2_X1 U14446 ( .A1(n8060), .A2(n7656), .ZN(n14226) );
  NAND2_X1 U14447 ( .A1(n14223), .A2(n14225), .ZN(n14393) );
  NAND2_X1 U14448 ( .A1(n14396), .A2(n14397), .ZN(n14225) );
  NAND2_X1 U14449 ( .A1(n14398), .A2(a_22_), .ZN(n14397) );
  NOR2_X1 U14450 ( .A1(n14399), .A2(n8060), .ZN(n14398) );
  NOR2_X1 U14451 ( .A1(n14221), .A2(n14220), .ZN(n14399) );
  NAND2_X1 U14452 ( .A1(n14220), .A2(n14221), .ZN(n14396) );
  NAND2_X1 U14453 ( .A1(n14400), .A2(n14401), .ZN(n14221) );
  NAND2_X1 U14454 ( .A1(n14218), .A2(n14402), .ZN(n14401) );
  NAND2_X1 U14455 ( .A1(n14217), .A2(n14216), .ZN(n14402) );
  NOR2_X1 U14456 ( .A1(n8060), .A2(n7624), .ZN(n14218) );
  OR2_X1 U14457 ( .A1(n14216), .A2(n14217), .ZN(n14400) );
  AND2_X1 U14458 ( .A1(n14163), .A2(n14403), .ZN(n14217) );
  NAND2_X1 U14459 ( .A1(n14162), .A2(n14164), .ZN(n14403) );
  NAND2_X1 U14460 ( .A1(n14404), .A2(n14405), .ZN(n14164) );
  NAND2_X1 U14461 ( .A1(a_24_), .A2(b_6_), .ZN(n14405) );
  INV_X1 U14462 ( .A(n14406), .ZN(n14404) );
  XOR2_X1 U14463 ( .A(n14407), .B(n14408), .Z(n14162) );
  XOR2_X1 U14464 ( .A(n14409), .B(n14410), .Z(n14407) );
  NOR2_X1 U14465 ( .A1(n7915), .A2(n7593), .ZN(n14410) );
  NAND2_X1 U14466 ( .A1(a_24_), .A2(n14406), .ZN(n14163) );
  NAND2_X1 U14467 ( .A1(n14411), .A2(n14412), .ZN(n14406) );
  NAND2_X1 U14468 ( .A1(n14413), .A2(a_25_), .ZN(n14412) );
  NOR2_X1 U14469 ( .A1(n14414), .A2(n8060), .ZN(n14413) );
  NOR2_X1 U14470 ( .A1(n14171), .A2(n14169), .ZN(n14414) );
  NAND2_X1 U14471 ( .A1(n14169), .A2(n14171), .ZN(n14411) );
  NAND2_X1 U14472 ( .A1(n14415), .A2(n14416), .ZN(n14171) );
  NAND2_X1 U14473 ( .A1(n14417), .A2(a_26_), .ZN(n14416) );
  NOR2_X1 U14474 ( .A1(n14418), .A2(n8060), .ZN(n14417) );
  NOR2_X1 U14475 ( .A1(n14214), .A2(n14212), .ZN(n14418) );
  NAND2_X1 U14476 ( .A1(n14212), .A2(n14214), .ZN(n14415) );
  NAND2_X1 U14477 ( .A1(n14419), .A2(n14420), .ZN(n14214) );
  NAND2_X1 U14478 ( .A1(n14210), .A2(n14421), .ZN(n14420) );
  NAND2_X1 U14479 ( .A1(n14209), .A2(n14208), .ZN(n14421) );
  NOR2_X1 U14480 ( .A1(n8060), .A2(n7563), .ZN(n14210) );
  OR2_X1 U14481 ( .A1(n14208), .A2(n14209), .ZN(n14419) );
  AND2_X1 U14482 ( .A1(n14205), .A2(n14422), .ZN(n14209) );
  NAND2_X1 U14483 ( .A1(n14204), .A2(n14206), .ZN(n14422) );
  NAND2_X1 U14484 ( .A1(n14423), .A2(n14424), .ZN(n14206) );
  NAND2_X1 U14485 ( .A1(b_6_), .A2(a_28_), .ZN(n14424) );
  INV_X1 U14486 ( .A(n14425), .ZN(n14423) );
  XOR2_X1 U14487 ( .A(n14426), .B(n14427), .Z(n14204) );
  NOR2_X1 U14488 ( .A1(n7529), .A2(n7915), .ZN(n14427) );
  XOR2_X1 U14489 ( .A(n14428), .B(n14429), .Z(n14426) );
  NAND2_X1 U14490 ( .A1(a_28_), .A2(n14425), .ZN(n14205) );
  NAND2_X1 U14491 ( .A1(n14430), .A2(n14431), .ZN(n14425) );
  NAND2_X1 U14492 ( .A1(n14432), .A2(b_6_), .ZN(n14431) );
  NOR2_X1 U14493 ( .A1(n14433), .A2(n7529), .ZN(n14432) );
  NOR2_X1 U14494 ( .A1(n14190), .A2(n14191), .ZN(n14433) );
  NAND2_X1 U14495 ( .A1(n14190), .A2(n14191), .ZN(n14430) );
  NAND2_X1 U14496 ( .A1(n14434), .A2(n14435), .ZN(n14191) );
  NAND2_X1 U14497 ( .A1(n14436), .A2(b_4_), .ZN(n14435) );
  NOR2_X1 U14498 ( .A1(n14437), .A2(n8048), .ZN(n14436) );
  NOR2_X1 U14499 ( .A1(n8676), .A2(n7915), .ZN(n14437) );
  NAND2_X1 U14500 ( .A1(n14438), .A2(b_5_), .ZN(n14434) );
  NOR2_X1 U14501 ( .A1(n14439), .A2(n7515), .ZN(n14438) );
  NOR2_X1 U14502 ( .A1(n8679), .A2(n8062), .ZN(n14439) );
  AND2_X1 U14503 ( .A1(n14440), .A2(b_5_), .ZN(n14190) );
  NOR2_X1 U14504 ( .A1(n8451), .A2(n8060), .ZN(n14440) );
  XOR2_X1 U14505 ( .A(n14441), .B(n14442), .Z(n14208) );
  NAND2_X1 U14506 ( .A1(n14443), .A2(n14444), .ZN(n14441) );
  XNOR2_X1 U14507 ( .A(n14445), .B(n14446), .ZN(n14212) );
  XNOR2_X1 U14508 ( .A(n14447), .B(n14448), .ZN(n14445) );
  XNOR2_X1 U14509 ( .A(n14449), .B(n14450), .ZN(n14169) );
  XNOR2_X1 U14510 ( .A(n14451), .B(n14452), .ZN(n14449) );
  XOR2_X1 U14511 ( .A(n14453), .B(n14454), .Z(n14216) );
  NAND2_X1 U14512 ( .A1(n14455), .A2(n14456), .ZN(n14453) );
  XOR2_X1 U14513 ( .A(n14457), .B(n14458), .Z(n14220) );
  XOR2_X1 U14514 ( .A(n14459), .B(n14460), .Z(n14457) );
  NOR2_X1 U14515 ( .A1(n7624), .A2(n7915), .ZN(n14460) );
  XNOR2_X1 U14516 ( .A(n14461), .B(n14462), .ZN(n14223) );
  XOR2_X1 U14517 ( .A(n14463), .B(n14464), .Z(n14462) );
  NAND2_X1 U14518 ( .A1(a_22_), .A2(b_5_), .ZN(n14464) );
  XNOR2_X1 U14519 ( .A(n14465), .B(n14466), .ZN(n14228) );
  XOR2_X1 U14520 ( .A(n14467), .B(n14468), .Z(n14466) );
  NAND2_X1 U14521 ( .A1(b_5_), .A2(a_21_), .ZN(n14468) );
  XOR2_X1 U14522 ( .A(n14469), .B(n14470), .Z(n14231) );
  XOR2_X1 U14523 ( .A(n14471), .B(n14472), .Z(n14469) );
  NOR2_X1 U14524 ( .A1(n7676), .A2(n7915), .ZN(n14472) );
  XNOR2_X1 U14525 ( .A(n14473), .B(n14474), .ZN(n14236) );
  XOR2_X1 U14526 ( .A(n14475), .B(n14476), .Z(n14473) );
  NOR2_X1 U14527 ( .A1(n7915), .A2(n7687), .ZN(n14476) );
  XOR2_X1 U14528 ( .A(n14477), .B(n14478), .Z(n14239) );
  XOR2_X1 U14529 ( .A(n14479), .B(n14480), .Z(n14477) );
  NOR2_X1 U14530 ( .A1(n7915), .A2(n7707), .ZN(n14480) );
  XOR2_X1 U14531 ( .A(n14481), .B(n14482), .Z(n14243) );
  XOR2_X1 U14532 ( .A(n14483), .B(n14484), .Z(n14481) );
  NOR2_X1 U14533 ( .A1(n7915), .A2(n7723), .ZN(n14484) );
  XOR2_X1 U14534 ( .A(n14485), .B(n14486), .Z(n14247) );
  XOR2_X1 U14535 ( .A(n14487), .B(n14488), .Z(n14485) );
  NOR2_X1 U14536 ( .A1(n7915), .A2(n7743), .ZN(n14488) );
  XOR2_X1 U14537 ( .A(n14489), .B(n14490), .Z(n14251) );
  XOR2_X1 U14538 ( .A(n14491), .B(n14492), .Z(n14489) );
  NOR2_X1 U14539 ( .A1(n7915), .A2(n7754), .ZN(n14492) );
  XOR2_X1 U14540 ( .A(n14493), .B(n14494), .Z(n14255) );
  XOR2_X1 U14541 ( .A(n14495), .B(n14496), .Z(n14493) );
  NOR2_X1 U14542 ( .A1(n7915), .A2(n7775), .ZN(n14496) );
  XOR2_X1 U14543 ( .A(n14497), .B(n14498), .Z(n14259) );
  XOR2_X1 U14544 ( .A(n14499), .B(n14500), .Z(n14497) );
  NOR2_X1 U14545 ( .A1(n7915), .A2(n7786), .ZN(n14500) );
  XOR2_X1 U14546 ( .A(n14501), .B(n14502), .Z(n14264) );
  XOR2_X1 U14547 ( .A(n14503), .B(n14504), .Z(n14501) );
  NOR2_X1 U14548 ( .A1(n7915), .A2(n7806), .ZN(n14504) );
  XOR2_X1 U14549 ( .A(n14505), .B(n14506), .Z(n14268) );
  XOR2_X1 U14550 ( .A(n14507), .B(n14508), .Z(n14505) );
  NOR2_X1 U14551 ( .A1(n7817), .A2(n7915), .ZN(n14508) );
  XOR2_X1 U14552 ( .A(n14509), .B(n14510), .Z(n14272) );
  XOR2_X1 U14553 ( .A(n14511), .B(n14512), .Z(n14509) );
  NOR2_X1 U14554 ( .A1(n7915), .A2(n7837), .ZN(n14512) );
  XOR2_X1 U14555 ( .A(n14513), .B(n14514), .Z(n14094) );
  XOR2_X1 U14556 ( .A(n14515), .B(n14516), .Z(n14513) );
  NOR2_X1 U14557 ( .A1(n7915), .A2(n7848), .ZN(n14516) );
  XOR2_X1 U14558 ( .A(n14517), .B(n14518), .Z(n14276) );
  XOR2_X1 U14559 ( .A(n14519), .B(n14520), .Z(n14517) );
  NOR2_X1 U14560 ( .A1(n7915), .A2(n8059), .ZN(n14520) );
  INV_X1 U14561 ( .A(n7898), .ZN(n14282) );
  NAND2_X1 U14562 ( .A1(a_6_), .A2(b_6_), .ZN(n7898) );
  XOR2_X1 U14563 ( .A(n14521), .B(n14522), .Z(n14284) );
  XOR2_X1 U14564 ( .A(n14523), .B(n14524), .Z(n14521) );
  NOR2_X1 U14565 ( .A1(n7915), .A2(n8061), .ZN(n14524) );
  XOR2_X1 U14566 ( .A(n14525), .B(n14526), .Z(n14288) );
  XOR2_X1 U14567 ( .A(n14527), .B(n7909), .Z(n14525) );
  XOR2_X1 U14568 ( .A(n14528), .B(n14529), .Z(n14292) );
  XNOR2_X1 U14569 ( .A(n14530), .B(n14531), .ZN(n14528) );
  NAND2_X1 U14570 ( .A1(a_4_), .A2(b_5_), .ZN(n14530) );
  XOR2_X1 U14571 ( .A(n14532), .B(n14533), .Z(n14295) );
  XNOR2_X1 U14572 ( .A(n14534), .B(n14535), .ZN(n14532) );
  NAND2_X1 U14573 ( .A1(a_3_), .A2(b_5_), .ZN(n14534) );
  XOR2_X1 U14574 ( .A(n14536), .B(n14537), .Z(n14299) );
  XOR2_X1 U14575 ( .A(n14538), .B(n14539), .Z(n14536) );
  NOR2_X1 U14576 ( .A1(n7915), .A2(n7965), .ZN(n14539) );
  XOR2_X1 U14577 ( .A(n14540), .B(n14541), .Z(n14304) );
  XOR2_X1 U14578 ( .A(n14542), .B(n14543), .Z(n14540) );
  NOR2_X1 U14579 ( .A1(n7915), .A2(n7973), .ZN(n14543) );
  NOR2_X1 U14580 ( .A1(n14544), .A2(n14061), .ZN(n14314) );
  XNOR2_X1 U14581 ( .A(n14545), .B(n14546), .ZN(n14061) );
  XOR2_X1 U14582 ( .A(n14547), .B(n14548), .Z(n14545) );
  AND2_X1 U14583 ( .A1(n14313), .A2(n14312), .ZN(n14544) );
  NAND2_X1 U14584 ( .A1(n14549), .A2(n14311), .ZN(n7712) );
  INV_X1 U14585 ( .A(n14316), .ZN(n14311) );
  XOR2_X1 U14586 ( .A(n14550), .B(n14551), .Z(n14549) );
  NAND2_X1 U14587 ( .A1(n14316), .A2(n14552), .ZN(n7711) );
  XOR2_X1 U14588 ( .A(n14550), .B(n14553), .Z(n14552) );
  NOR2_X1 U14589 ( .A1(n14313), .A2(n14312), .ZN(n14316) );
  AND2_X1 U14590 ( .A1(n14554), .A2(n14555), .ZN(n14312) );
  NAND2_X1 U14591 ( .A1(n14548), .A2(n14556), .ZN(n14555) );
  OR2_X1 U14592 ( .A1(n14547), .A2(n14546), .ZN(n14556) );
  NOR2_X1 U14593 ( .A1(n7915), .A2(n8307), .ZN(n14548) );
  NAND2_X1 U14594 ( .A1(n14546), .A2(n14547), .ZN(n14554) );
  NAND2_X1 U14595 ( .A1(n14557), .A2(n14558), .ZN(n14547) );
  NAND2_X1 U14596 ( .A1(n14559), .A2(a_1_), .ZN(n14558) );
  NOR2_X1 U14597 ( .A1(n14560), .A2(n7915), .ZN(n14559) );
  NOR2_X1 U14598 ( .A1(n14541), .A2(n14542), .ZN(n14560) );
  NAND2_X1 U14599 ( .A1(n14541), .A2(n14542), .ZN(n14557) );
  NAND2_X1 U14600 ( .A1(n14561), .A2(n14562), .ZN(n14542) );
  NAND2_X1 U14601 ( .A1(n14563), .A2(a_2_), .ZN(n14562) );
  NOR2_X1 U14602 ( .A1(n14564), .A2(n7915), .ZN(n14563) );
  NOR2_X1 U14603 ( .A1(n14537), .A2(n14538), .ZN(n14564) );
  NAND2_X1 U14604 ( .A1(n14537), .A2(n14538), .ZN(n14561) );
  NAND2_X1 U14605 ( .A1(n14565), .A2(n14566), .ZN(n14538) );
  NAND2_X1 U14606 ( .A1(n14567), .A2(a_3_), .ZN(n14566) );
  NOR2_X1 U14607 ( .A1(n14568), .A2(n7915), .ZN(n14567) );
  NOR2_X1 U14608 ( .A1(n14533), .A2(n14535), .ZN(n14568) );
  NAND2_X1 U14609 ( .A1(n14533), .A2(n14535), .ZN(n14565) );
  NAND2_X1 U14610 ( .A1(n14569), .A2(n14570), .ZN(n14535) );
  NAND2_X1 U14611 ( .A1(n14571), .A2(a_4_), .ZN(n14570) );
  NOR2_X1 U14612 ( .A1(n14572), .A2(n7915), .ZN(n14571) );
  NOR2_X1 U14613 ( .A1(n14529), .A2(n14531), .ZN(n14572) );
  NAND2_X1 U14614 ( .A1(n14529), .A2(n14531), .ZN(n14569) );
  NAND2_X1 U14615 ( .A1(n14573), .A2(n14574), .ZN(n14531) );
  NAND2_X1 U14616 ( .A1(n14526), .A2(n14575), .ZN(n14574) );
  OR2_X1 U14617 ( .A1(n14527), .A2(n7909), .ZN(n14575) );
  XNOR2_X1 U14618 ( .A(n14576), .B(n14577), .ZN(n14526) );
  XOR2_X1 U14619 ( .A(n14578), .B(n14579), .Z(n14577) );
  NAND2_X1 U14620 ( .A1(a_6_), .A2(b_4_), .ZN(n14579) );
  NAND2_X1 U14621 ( .A1(n7909), .A2(n14527), .ZN(n14573) );
  NAND2_X1 U14622 ( .A1(n14580), .A2(n14581), .ZN(n14527) );
  NAND2_X1 U14623 ( .A1(n14582), .A2(a_6_), .ZN(n14581) );
  NOR2_X1 U14624 ( .A1(n14583), .A2(n7915), .ZN(n14582) );
  NOR2_X1 U14625 ( .A1(n14522), .A2(n14523), .ZN(n14583) );
  NAND2_X1 U14626 ( .A1(n14522), .A2(n14523), .ZN(n14580) );
  NAND2_X1 U14627 ( .A1(n14584), .A2(n14585), .ZN(n14523) );
  NAND2_X1 U14628 ( .A1(n14586), .A2(a_7_), .ZN(n14585) );
  NOR2_X1 U14629 ( .A1(n14587), .A2(n7915), .ZN(n14586) );
  NOR2_X1 U14630 ( .A1(n14344), .A2(n14345), .ZN(n14587) );
  NAND2_X1 U14631 ( .A1(n14344), .A2(n14345), .ZN(n14584) );
  NAND2_X1 U14632 ( .A1(n14588), .A2(n14589), .ZN(n14345) );
  NAND2_X1 U14633 ( .A1(n14590), .A2(a_8_), .ZN(n14589) );
  NOR2_X1 U14634 ( .A1(n14591), .A2(n7915), .ZN(n14590) );
  NOR2_X1 U14635 ( .A1(n14518), .A2(n14519), .ZN(n14591) );
  NAND2_X1 U14636 ( .A1(n14518), .A2(n14519), .ZN(n14588) );
  NAND2_X1 U14637 ( .A1(n14592), .A2(n14593), .ZN(n14519) );
  NAND2_X1 U14638 ( .A1(n14594), .A2(a_9_), .ZN(n14593) );
  NOR2_X1 U14639 ( .A1(n14595), .A2(n7915), .ZN(n14594) );
  NOR2_X1 U14640 ( .A1(n14514), .A2(n14515), .ZN(n14595) );
  NAND2_X1 U14641 ( .A1(n14514), .A2(n14515), .ZN(n14592) );
  NAND2_X1 U14642 ( .A1(n14596), .A2(n14597), .ZN(n14515) );
  NAND2_X1 U14643 ( .A1(n14598), .A2(a_10_), .ZN(n14597) );
  NOR2_X1 U14644 ( .A1(n14599), .A2(n7915), .ZN(n14598) );
  NOR2_X1 U14645 ( .A1(n14510), .A2(n14511), .ZN(n14599) );
  NAND2_X1 U14646 ( .A1(n14510), .A2(n14511), .ZN(n14596) );
  NAND2_X1 U14647 ( .A1(n14600), .A2(n14601), .ZN(n14511) );
  NAND2_X1 U14648 ( .A1(n14602), .A2(b_5_), .ZN(n14601) );
  NOR2_X1 U14649 ( .A1(n14603), .A2(n7817), .ZN(n14602) );
  NOR2_X1 U14650 ( .A1(n14506), .A2(n14507), .ZN(n14603) );
  NAND2_X1 U14651 ( .A1(n14506), .A2(n14507), .ZN(n14600) );
  NAND2_X1 U14652 ( .A1(n14604), .A2(n14605), .ZN(n14507) );
  NAND2_X1 U14653 ( .A1(n14606), .A2(a_12_), .ZN(n14605) );
  NOR2_X1 U14654 ( .A1(n14607), .A2(n7915), .ZN(n14606) );
  NOR2_X1 U14655 ( .A1(n14502), .A2(n14503), .ZN(n14607) );
  NAND2_X1 U14656 ( .A1(n14502), .A2(n14503), .ZN(n14604) );
  NAND2_X1 U14657 ( .A1(n14608), .A2(n14609), .ZN(n14503) );
  NAND2_X1 U14658 ( .A1(n14610), .A2(a_13_), .ZN(n14609) );
  NOR2_X1 U14659 ( .A1(n14611), .A2(n7915), .ZN(n14610) );
  NOR2_X1 U14660 ( .A1(n14498), .A2(n14499), .ZN(n14611) );
  NAND2_X1 U14661 ( .A1(n14498), .A2(n14499), .ZN(n14608) );
  NAND2_X1 U14662 ( .A1(n14612), .A2(n14613), .ZN(n14499) );
  NAND2_X1 U14663 ( .A1(n14614), .A2(a_14_), .ZN(n14613) );
  NOR2_X1 U14664 ( .A1(n14615), .A2(n7915), .ZN(n14614) );
  NOR2_X1 U14665 ( .A1(n14494), .A2(n14495), .ZN(n14615) );
  NAND2_X1 U14666 ( .A1(n14494), .A2(n14495), .ZN(n14612) );
  NAND2_X1 U14667 ( .A1(n14616), .A2(n14617), .ZN(n14495) );
  NAND2_X1 U14668 ( .A1(n14618), .A2(a_15_), .ZN(n14617) );
  NOR2_X1 U14669 ( .A1(n14619), .A2(n7915), .ZN(n14618) );
  NOR2_X1 U14670 ( .A1(n14491), .A2(n14490), .ZN(n14619) );
  NAND2_X1 U14671 ( .A1(n14490), .A2(n14491), .ZN(n14616) );
  NAND2_X1 U14672 ( .A1(n14620), .A2(n14621), .ZN(n14491) );
  NAND2_X1 U14673 ( .A1(n14622), .A2(a_16_), .ZN(n14621) );
  NOR2_X1 U14674 ( .A1(n14623), .A2(n7915), .ZN(n14622) );
  NOR2_X1 U14675 ( .A1(n14486), .A2(n14487), .ZN(n14623) );
  NAND2_X1 U14676 ( .A1(n14486), .A2(n14487), .ZN(n14620) );
  NAND2_X1 U14677 ( .A1(n14624), .A2(n14625), .ZN(n14487) );
  NAND2_X1 U14678 ( .A1(n14626), .A2(a_17_), .ZN(n14625) );
  NOR2_X1 U14679 ( .A1(n14627), .A2(n7915), .ZN(n14626) );
  NOR2_X1 U14680 ( .A1(n14483), .A2(n14482), .ZN(n14627) );
  NAND2_X1 U14681 ( .A1(n14482), .A2(n14483), .ZN(n14624) );
  NAND2_X1 U14682 ( .A1(n14628), .A2(n14629), .ZN(n14483) );
  NAND2_X1 U14683 ( .A1(n14630), .A2(a_18_), .ZN(n14629) );
  NOR2_X1 U14684 ( .A1(n14631), .A2(n7915), .ZN(n14630) );
  NOR2_X1 U14685 ( .A1(n14478), .A2(n14479), .ZN(n14631) );
  NAND2_X1 U14686 ( .A1(n14478), .A2(n14479), .ZN(n14628) );
  NAND2_X1 U14687 ( .A1(n14632), .A2(n14633), .ZN(n14479) );
  NAND2_X1 U14688 ( .A1(n14634), .A2(a_19_), .ZN(n14633) );
  NOR2_X1 U14689 ( .A1(n14635), .A2(n7915), .ZN(n14634) );
  NOR2_X1 U14690 ( .A1(n14475), .A2(n14474), .ZN(n14635) );
  NAND2_X1 U14691 ( .A1(n14474), .A2(n14475), .ZN(n14632) );
  NAND2_X1 U14692 ( .A1(n14636), .A2(n14637), .ZN(n14475) );
  NAND2_X1 U14693 ( .A1(n14638), .A2(b_5_), .ZN(n14637) );
  NOR2_X1 U14694 ( .A1(n14639), .A2(n7676), .ZN(n14638) );
  NOR2_X1 U14695 ( .A1(n14470), .A2(n14471), .ZN(n14639) );
  NAND2_X1 U14696 ( .A1(n14470), .A2(n14471), .ZN(n14636) );
  NAND2_X1 U14697 ( .A1(n14640), .A2(n14641), .ZN(n14471) );
  NAND2_X1 U14698 ( .A1(n14642), .A2(b_5_), .ZN(n14641) );
  NOR2_X1 U14699 ( .A1(n14643), .A2(n7656), .ZN(n14642) );
  NOR2_X1 U14700 ( .A1(n14467), .A2(n14465), .ZN(n14643) );
  NAND2_X1 U14701 ( .A1(n14465), .A2(n14467), .ZN(n14640) );
  NAND2_X1 U14702 ( .A1(n14644), .A2(n14645), .ZN(n14467) );
  NAND2_X1 U14703 ( .A1(n14646), .A2(a_22_), .ZN(n14645) );
  NOR2_X1 U14704 ( .A1(n14647), .A2(n7915), .ZN(n14646) );
  NOR2_X1 U14705 ( .A1(n14461), .A2(n14463), .ZN(n14647) );
  NAND2_X1 U14706 ( .A1(n14461), .A2(n14463), .ZN(n14644) );
  NAND2_X1 U14707 ( .A1(n14648), .A2(n14649), .ZN(n14463) );
  NAND2_X1 U14708 ( .A1(n14650), .A2(b_5_), .ZN(n14649) );
  NOR2_X1 U14709 ( .A1(n14651), .A2(n7624), .ZN(n14650) );
  NOR2_X1 U14710 ( .A1(n14458), .A2(n14459), .ZN(n14651) );
  NAND2_X1 U14711 ( .A1(n14458), .A2(n14459), .ZN(n14648) );
  NAND2_X1 U14712 ( .A1(n14455), .A2(n14652), .ZN(n14459) );
  NAND2_X1 U14713 ( .A1(n14454), .A2(n14456), .ZN(n14652) );
  NAND2_X1 U14714 ( .A1(n14653), .A2(n14654), .ZN(n14456) );
  NAND2_X1 U14715 ( .A1(a_24_), .A2(b_5_), .ZN(n14654) );
  INV_X1 U14716 ( .A(n14655), .ZN(n14653) );
  XOR2_X1 U14717 ( .A(n14656), .B(n14657), .Z(n14454) );
  XOR2_X1 U14718 ( .A(n14658), .B(n14659), .Z(n14656) );
  NOR2_X1 U14719 ( .A1(n7593), .A2(n8062), .ZN(n14659) );
  NAND2_X1 U14720 ( .A1(a_24_), .A2(n14655), .ZN(n14455) );
  NAND2_X1 U14721 ( .A1(n14660), .A2(n14661), .ZN(n14655) );
  NAND2_X1 U14722 ( .A1(n14662), .A2(a_25_), .ZN(n14661) );
  NOR2_X1 U14723 ( .A1(n14663), .A2(n7915), .ZN(n14662) );
  NOR2_X1 U14724 ( .A1(n14409), .A2(n14408), .ZN(n14663) );
  NAND2_X1 U14725 ( .A1(n14408), .A2(n14409), .ZN(n14660) );
  NAND2_X1 U14726 ( .A1(n14664), .A2(n14665), .ZN(n14409) );
  NAND2_X1 U14727 ( .A1(n14451), .A2(n14666), .ZN(n14665) );
  NAND2_X1 U14728 ( .A1(n14452), .A2(n14450), .ZN(n14666) );
  NOR2_X1 U14729 ( .A1(n7915), .A2(n8052), .ZN(n14451) );
  OR2_X1 U14730 ( .A1(n14450), .A2(n14452), .ZN(n14664) );
  AND2_X1 U14731 ( .A1(n14667), .A2(n14668), .ZN(n14452) );
  NAND2_X1 U14732 ( .A1(n14448), .A2(n14669), .ZN(n14668) );
  NAND2_X1 U14733 ( .A1(n14447), .A2(n14446), .ZN(n14669) );
  NOR2_X1 U14734 ( .A1(n7915), .A2(n7563), .ZN(n14448) );
  OR2_X1 U14735 ( .A1(n14446), .A2(n14447), .ZN(n14667) );
  AND2_X1 U14736 ( .A1(n14443), .A2(n14670), .ZN(n14447) );
  NAND2_X1 U14737 ( .A1(n14442), .A2(n14444), .ZN(n14670) );
  NAND2_X1 U14738 ( .A1(n14671), .A2(n14672), .ZN(n14444) );
  NAND2_X1 U14739 ( .A1(b_5_), .A2(a_28_), .ZN(n14672) );
  INV_X1 U14740 ( .A(n14673), .ZN(n14671) );
  XOR2_X1 U14741 ( .A(n14674), .B(n14675), .Z(n14442) );
  NOR2_X1 U14742 ( .A1(n7529), .A2(n8062), .ZN(n14675) );
  XOR2_X1 U14743 ( .A(n14676), .B(n14677), .Z(n14674) );
  NAND2_X1 U14744 ( .A1(a_28_), .A2(n14673), .ZN(n14443) );
  NAND2_X1 U14745 ( .A1(n14678), .A2(n14679), .ZN(n14673) );
  NAND2_X1 U14746 ( .A1(n14680), .A2(b_5_), .ZN(n14679) );
  NOR2_X1 U14747 ( .A1(n14681), .A2(n7529), .ZN(n14680) );
  NOR2_X1 U14748 ( .A1(n14428), .A2(n14429), .ZN(n14681) );
  NAND2_X1 U14749 ( .A1(n14428), .A2(n14429), .ZN(n14678) );
  NAND2_X1 U14750 ( .A1(n14682), .A2(n14683), .ZN(n14429) );
  NAND2_X1 U14751 ( .A1(n14684), .A2(b_3_), .ZN(n14683) );
  NOR2_X1 U14752 ( .A1(n14685), .A2(n8048), .ZN(n14684) );
  NOR2_X1 U14753 ( .A1(n8676), .A2(n8062), .ZN(n14685) );
  NAND2_X1 U14754 ( .A1(n14686), .A2(b_4_), .ZN(n14682) );
  NOR2_X1 U14755 ( .A1(n14687), .A2(n7515), .ZN(n14686) );
  NOR2_X1 U14756 ( .A1(n8679), .A2(n7946), .ZN(n14687) );
  AND2_X1 U14757 ( .A1(n14688), .A2(b_4_), .ZN(n14428) );
  NOR2_X1 U14758 ( .A1(n8451), .A2(n7915), .ZN(n14688) );
  XOR2_X1 U14759 ( .A(n14689), .B(n14690), .Z(n14446) );
  NAND2_X1 U14760 ( .A1(n14691), .A2(n14692), .ZN(n14689) );
  XOR2_X1 U14761 ( .A(n14693), .B(n14694), .Z(n14450) );
  XOR2_X1 U14762 ( .A(n14695), .B(n14696), .Z(n14694) );
  NAND2_X1 U14763 ( .A1(b_4_), .A2(a_27_), .ZN(n14696) );
  XNOR2_X1 U14764 ( .A(n14697), .B(n14698), .ZN(n14408) );
  XNOR2_X1 U14765 ( .A(n14699), .B(n14700), .ZN(n14697) );
  XNOR2_X1 U14766 ( .A(n14701), .B(n14702), .ZN(n14458) );
  XNOR2_X1 U14767 ( .A(n14703), .B(n14704), .ZN(n14702) );
  XOR2_X1 U14768 ( .A(n14705), .B(n14706), .Z(n14461) );
  XOR2_X1 U14769 ( .A(n14707), .B(n14708), .Z(n14705) );
  XNOR2_X1 U14770 ( .A(n14709), .B(n14710), .ZN(n14465) );
  XNOR2_X1 U14771 ( .A(n14711), .B(n14712), .ZN(n14709) );
  XNOR2_X1 U14772 ( .A(n14713), .B(n14714), .ZN(n14470) );
  XNOR2_X1 U14773 ( .A(n14715), .B(n14716), .ZN(n14714) );
  XNOR2_X1 U14774 ( .A(n14717), .B(n14718), .ZN(n14474) );
  XNOR2_X1 U14775 ( .A(n14719), .B(n14720), .ZN(n14717) );
  XNOR2_X1 U14776 ( .A(n14721), .B(n14722), .ZN(n14478) );
  XNOR2_X1 U14777 ( .A(n14723), .B(n14724), .ZN(n14722) );
  XNOR2_X1 U14778 ( .A(n14725), .B(n14726), .ZN(n14482) );
  XNOR2_X1 U14779 ( .A(n14727), .B(n14728), .ZN(n14725) );
  XNOR2_X1 U14780 ( .A(n14729), .B(n14730), .ZN(n14486) );
  XNOR2_X1 U14781 ( .A(n14731), .B(n14732), .ZN(n14730) );
  XNOR2_X1 U14782 ( .A(n14733), .B(n14734), .ZN(n14490) );
  XNOR2_X1 U14783 ( .A(n14735), .B(n14736), .ZN(n14733) );
  XNOR2_X1 U14784 ( .A(n14737), .B(n14738), .ZN(n14494) );
  XNOR2_X1 U14785 ( .A(n14739), .B(n14740), .ZN(n14738) );
  XOR2_X1 U14786 ( .A(n14741), .B(n14742), .Z(n14498) );
  XOR2_X1 U14787 ( .A(n14743), .B(n14744), .Z(n14741) );
  XNOR2_X1 U14788 ( .A(n14745), .B(n14746), .ZN(n14502) );
  XOR2_X1 U14789 ( .A(n14747), .B(n14748), .Z(n14746) );
  NAND2_X1 U14790 ( .A1(a_13_), .A2(b_4_), .ZN(n14748) );
  XNOR2_X1 U14791 ( .A(n14749), .B(n14750), .ZN(n14506) );
  XOR2_X1 U14792 ( .A(n14751), .B(n14752), .Z(n14750) );
  NAND2_X1 U14793 ( .A1(a_12_), .A2(b_4_), .ZN(n14752) );
  XNOR2_X1 U14794 ( .A(n14753), .B(n14754), .ZN(n14510) );
  XOR2_X1 U14795 ( .A(n14755), .B(n14756), .Z(n14754) );
  NAND2_X1 U14796 ( .A1(b_4_), .A2(a_11_), .ZN(n14756) );
  XNOR2_X1 U14797 ( .A(n14757), .B(n14758), .ZN(n14514) );
  XOR2_X1 U14798 ( .A(n14759), .B(n14760), .Z(n14758) );
  NAND2_X1 U14799 ( .A1(a_10_), .A2(b_4_), .ZN(n14760) );
  XNOR2_X1 U14800 ( .A(n14761), .B(n14762), .ZN(n14518) );
  XOR2_X1 U14801 ( .A(n14763), .B(n14764), .Z(n14762) );
  NAND2_X1 U14802 ( .A1(a_9_), .A2(b_4_), .ZN(n14764) );
  XNOR2_X1 U14803 ( .A(n14765), .B(n14766), .ZN(n14344) );
  XOR2_X1 U14804 ( .A(n14767), .B(n14768), .Z(n14766) );
  NAND2_X1 U14805 ( .A1(a_8_), .A2(b_4_), .ZN(n14768) );
  XNOR2_X1 U14806 ( .A(n14769), .B(n14770), .ZN(n14522) );
  XOR2_X1 U14807 ( .A(n14771), .B(n14772), .Z(n14770) );
  NAND2_X1 U14808 ( .A1(a_7_), .A2(b_4_), .ZN(n14772) );
  INV_X1 U14809 ( .A(n7996), .ZN(n7909) );
  NAND2_X1 U14810 ( .A1(a_5_), .A2(b_5_), .ZN(n7996) );
  XNOR2_X1 U14811 ( .A(n14773), .B(n14774), .ZN(n14529) );
  XOR2_X1 U14812 ( .A(n14775), .B(n14776), .Z(n14774) );
  NAND2_X1 U14813 ( .A1(a_5_), .A2(b_4_), .ZN(n14776) );
  XOR2_X1 U14814 ( .A(n14777), .B(n14778), .Z(n14533) );
  XOR2_X1 U14815 ( .A(n14779), .B(n14780), .Z(n14777) );
  XOR2_X1 U14816 ( .A(n14781), .B(n14782), .Z(n14537) );
  XNOR2_X1 U14817 ( .A(n14783), .B(n14784), .ZN(n14781) );
  NAND2_X1 U14818 ( .A1(a_3_), .A2(b_4_), .ZN(n14783) );
  XOR2_X1 U14819 ( .A(n14785), .B(n14786), .Z(n14541) );
  XOR2_X1 U14820 ( .A(n14787), .B(n14788), .Z(n14785) );
  NOR2_X1 U14821 ( .A1(n8062), .A2(n7965), .ZN(n14788) );
  XOR2_X1 U14822 ( .A(n14789), .B(n14790), .Z(n14546) );
  XOR2_X1 U14823 ( .A(n14791), .B(n14792), .Z(n14789) );
  NOR2_X1 U14824 ( .A1(n8062), .A2(n7973), .ZN(n14792) );
  XNOR2_X1 U14825 ( .A(n14793), .B(n14794), .ZN(n14313) );
  XOR2_X1 U14826 ( .A(n14795), .B(n14796), .Z(n14793) );
  NOR2_X1 U14827 ( .A1(n8307), .A2(n8062), .ZN(n14796) );
  NAND2_X1 U14828 ( .A1(n14797), .A2(n14798), .ZN(n7873) );
  NAND2_X1 U14829 ( .A1(n14799), .A2(n14800), .ZN(n14798) );
  OR2_X1 U14830 ( .A1(n14801), .A2(n14802), .ZN(n14799) );
  NAND2_X1 U14831 ( .A1(n14553), .A2(n14550), .ZN(n14797) );
  NAND2_X1 U14832 ( .A1(n14803), .A2(n14804), .ZN(n7872) );
  AND2_X1 U14833 ( .A1(n14800), .A2(n14550), .ZN(n14804) );
  NAND2_X1 U14834 ( .A1(n14805), .A2(n14806), .ZN(n14550) );
  NAND2_X1 U14835 ( .A1(n14807), .A2(b_4_), .ZN(n14806) );
  NOR2_X1 U14836 ( .A1(n14808), .A2(n8307), .ZN(n14807) );
  NOR2_X1 U14837 ( .A1(n14794), .A2(n14795), .ZN(n14808) );
  NAND2_X1 U14838 ( .A1(n14794), .A2(n14795), .ZN(n14805) );
  NAND2_X1 U14839 ( .A1(n14809), .A2(n14810), .ZN(n14795) );
  NAND2_X1 U14840 ( .A1(n14811), .A2(a_1_), .ZN(n14810) );
  NOR2_X1 U14841 ( .A1(n14812), .A2(n8062), .ZN(n14811) );
  NOR2_X1 U14842 ( .A1(n14791), .A2(n14790), .ZN(n14812) );
  NAND2_X1 U14843 ( .A1(n14790), .A2(n14791), .ZN(n14809) );
  NAND2_X1 U14844 ( .A1(n14813), .A2(n14814), .ZN(n14791) );
  NAND2_X1 U14845 ( .A1(n14815), .A2(a_2_), .ZN(n14814) );
  NOR2_X1 U14846 ( .A1(n14816), .A2(n8062), .ZN(n14815) );
  NOR2_X1 U14847 ( .A1(n14787), .A2(n14786), .ZN(n14816) );
  NAND2_X1 U14848 ( .A1(n14786), .A2(n14787), .ZN(n14813) );
  NAND2_X1 U14849 ( .A1(n14817), .A2(n14818), .ZN(n14787) );
  NAND2_X1 U14850 ( .A1(n14819), .A2(a_3_), .ZN(n14818) );
  NOR2_X1 U14851 ( .A1(n14820), .A2(n8062), .ZN(n14819) );
  NOR2_X1 U14852 ( .A1(n14784), .A2(n14782), .ZN(n14820) );
  NAND2_X1 U14853 ( .A1(n14782), .A2(n14784), .ZN(n14817) );
  NAND2_X1 U14854 ( .A1(n14821), .A2(n14822), .ZN(n14784) );
  NAND2_X1 U14855 ( .A1(n14778), .A2(n14823), .ZN(n14822) );
  OR2_X1 U14856 ( .A1(n14779), .A2(n14780), .ZN(n14823) );
  XOR2_X1 U14857 ( .A(n14824), .B(n14825), .Z(n14778) );
  XOR2_X1 U14858 ( .A(n14826), .B(n14827), .Z(n14824) );
  NOR2_X1 U14859 ( .A1(n7946), .A2(n7914), .ZN(n14827) );
  NAND2_X1 U14860 ( .A1(n14780), .A2(n14779), .ZN(n14821) );
  NAND2_X1 U14861 ( .A1(n14828), .A2(n14829), .ZN(n14779) );
  NAND2_X1 U14862 ( .A1(n14830), .A2(a_5_), .ZN(n14829) );
  NOR2_X1 U14863 ( .A1(n14831), .A2(n8062), .ZN(n14830) );
  NOR2_X1 U14864 ( .A1(n14775), .A2(n14773), .ZN(n14831) );
  NAND2_X1 U14865 ( .A1(n14773), .A2(n14775), .ZN(n14828) );
  NAND2_X1 U14866 ( .A1(n14832), .A2(n14833), .ZN(n14775) );
  NAND2_X1 U14867 ( .A1(n14834), .A2(a_6_), .ZN(n14833) );
  NOR2_X1 U14868 ( .A1(n14835), .A2(n8062), .ZN(n14834) );
  NOR2_X1 U14869 ( .A1(n14578), .A2(n14576), .ZN(n14835) );
  NAND2_X1 U14870 ( .A1(n14576), .A2(n14578), .ZN(n14832) );
  NAND2_X1 U14871 ( .A1(n14836), .A2(n14837), .ZN(n14578) );
  NAND2_X1 U14872 ( .A1(n14838), .A2(a_7_), .ZN(n14837) );
  NOR2_X1 U14873 ( .A1(n14839), .A2(n8062), .ZN(n14838) );
  NOR2_X1 U14874 ( .A1(n14771), .A2(n14769), .ZN(n14839) );
  NAND2_X1 U14875 ( .A1(n14769), .A2(n14771), .ZN(n14836) );
  NAND2_X1 U14876 ( .A1(n14840), .A2(n14841), .ZN(n14771) );
  NAND2_X1 U14877 ( .A1(n14842), .A2(a_8_), .ZN(n14841) );
  NOR2_X1 U14878 ( .A1(n14843), .A2(n8062), .ZN(n14842) );
  NOR2_X1 U14879 ( .A1(n14767), .A2(n14765), .ZN(n14843) );
  NAND2_X1 U14880 ( .A1(n14765), .A2(n14767), .ZN(n14840) );
  NAND2_X1 U14881 ( .A1(n14844), .A2(n14845), .ZN(n14767) );
  NAND2_X1 U14882 ( .A1(n14846), .A2(a_9_), .ZN(n14845) );
  NOR2_X1 U14883 ( .A1(n14847), .A2(n8062), .ZN(n14846) );
  NOR2_X1 U14884 ( .A1(n14763), .A2(n14761), .ZN(n14847) );
  NAND2_X1 U14885 ( .A1(n14761), .A2(n14763), .ZN(n14844) );
  NAND2_X1 U14886 ( .A1(n14848), .A2(n14849), .ZN(n14763) );
  NAND2_X1 U14887 ( .A1(n14850), .A2(a_10_), .ZN(n14849) );
  NOR2_X1 U14888 ( .A1(n14851), .A2(n8062), .ZN(n14850) );
  NOR2_X1 U14889 ( .A1(n14759), .A2(n14757), .ZN(n14851) );
  NAND2_X1 U14890 ( .A1(n14757), .A2(n14759), .ZN(n14848) );
  NAND2_X1 U14891 ( .A1(n14852), .A2(n14853), .ZN(n14759) );
  NAND2_X1 U14892 ( .A1(n14854), .A2(b_4_), .ZN(n14853) );
  NOR2_X1 U14893 ( .A1(n14855), .A2(n7817), .ZN(n14854) );
  NOR2_X1 U14894 ( .A1(n14755), .A2(n14753), .ZN(n14855) );
  NAND2_X1 U14895 ( .A1(n14753), .A2(n14755), .ZN(n14852) );
  NAND2_X1 U14896 ( .A1(n14856), .A2(n14857), .ZN(n14755) );
  NAND2_X1 U14897 ( .A1(n14858), .A2(a_12_), .ZN(n14857) );
  NOR2_X1 U14898 ( .A1(n14859), .A2(n8062), .ZN(n14858) );
  NOR2_X1 U14899 ( .A1(n14751), .A2(n14749), .ZN(n14859) );
  NAND2_X1 U14900 ( .A1(n14749), .A2(n14751), .ZN(n14856) );
  NAND2_X1 U14901 ( .A1(n14860), .A2(n14861), .ZN(n14751) );
  NAND2_X1 U14902 ( .A1(n14862), .A2(a_13_), .ZN(n14861) );
  NOR2_X1 U14903 ( .A1(n14863), .A2(n8062), .ZN(n14862) );
  NOR2_X1 U14904 ( .A1(n14747), .A2(n14745), .ZN(n14863) );
  NAND2_X1 U14905 ( .A1(n14745), .A2(n14747), .ZN(n14860) );
  NAND2_X1 U14906 ( .A1(n14864), .A2(n14865), .ZN(n14747) );
  NAND2_X1 U14907 ( .A1(n14744), .A2(n14866), .ZN(n14865) );
  OR2_X1 U14908 ( .A1(n14742), .A2(n14743), .ZN(n14866) );
  NOR2_X1 U14909 ( .A1(n7775), .A2(n8062), .ZN(n14744) );
  NAND2_X1 U14910 ( .A1(n14742), .A2(n14743), .ZN(n14864) );
  NAND2_X1 U14911 ( .A1(n14867), .A2(n14868), .ZN(n14743) );
  NAND2_X1 U14912 ( .A1(n14740), .A2(n14869), .ZN(n14868) );
  OR2_X1 U14913 ( .A1(n14737), .A2(n14739), .ZN(n14869) );
  NOR2_X1 U14914 ( .A1(n7754), .A2(n8062), .ZN(n14740) );
  NAND2_X1 U14915 ( .A1(n14737), .A2(n14739), .ZN(n14867) );
  NAND2_X1 U14916 ( .A1(n14870), .A2(n14871), .ZN(n14739) );
  NAND2_X1 U14917 ( .A1(n14736), .A2(n14872), .ZN(n14871) );
  NAND2_X1 U14918 ( .A1(n14735), .A2(n14734), .ZN(n14872) );
  NOR2_X1 U14919 ( .A1(n7743), .A2(n8062), .ZN(n14736) );
  OR2_X1 U14920 ( .A1(n14734), .A2(n14735), .ZN(n14870) );
  AND2_X1 U14921 ( .A1(n14873), .A2(n14874), .ZN(n14735) );
  NAND2_X1 U14922 ( .A1(n14732), .A2(n14875), .ZN(n14874) );
  OR2_X1 U14923 ( .A1(n14729), .A2(n14731), .ZN(n14875) );
  NOR2_X1 U14924 ( .A1(n7723), .A2(n8062), .ZN(n14732) );
  NAND2_X1 U14925 ( .A1(n14729), .A2(n14731), .ZN(n14873) );
  NAND2_X1 U14926 ( .A1(n14876), .A2(n14877), .ZN(n14731) );
  NAND2_X1 U14927 ( .A1(n14728), .A2(n14878), .ZN(n14877) );
  NAND2_X1 U14928 ( .A1(n14727), .A2(n14726), .ZN(n14878) );
  NOR2_X1 U14929 ( .A1(n7707), .A2(n8062), .ZN(n14728) );
  OR2_X1 U14930 ( .A1(n14726), .A2(n14727), .ZN(n14876) );
  AND2_X1 U14931 ( .A1(n14879), .A2(n14880), .ZN(n14727) );
  NAND2_X1 U14932 ( .A1(n14724), .A2(n14881), .ZN(n14880) );
  OR2_X1 U14933 ( .A1(n14721), .A2(n14723), .ZN(n14881) );
  NOR2_X1 U14934 ( .A1(n7687), .A2(n8062), .ZN(n14724) );
  NAND2_X1 U14935 ( .A1(n14721), .A2(n14723), .ZN(n14879) );
  NAND2_X1 U14936 ( .A1(n14882), .A2(n14883), .ZN(n14723) );
  NAND2_X1 U14937 ( .A1(n14720), .A2(n14884), .ZN(n14883) );
  NAND2_X1 U14938 ( .A1(n14719), .A2(n14718), .ZN(n14884) );
  NOR2_X1 U14939 ( .A1(n8062), .A2(n7676), .ZN(n14720) );
  OR2_X1 U14940 ( .A1(n14718), .A2(n14719), .ZN(n14882) );
  AND2_X1 U14941 ( .A1(n14885), .A2(n14886), .ZN(n14719) );
  NAND2_X1 U14942 ( .A1(n14716), .A2(n14887), .ZN(n14886) );
  OR2_X1 U14943 ( .A1(n14713), .A2(n14715), .ZN(n14887) );
  NOR2_X1 U14944 ( .A1(n8062), .A2(n7656), .ZN(n14716) );
  NAND2_X1 U14945 ( .A1(n14713), .A2(n14715), .ZN(n14885) );
  NAND2_X1 U14946 ( .A1(n14888), .A2(n14889), .ZN(n14715) );
  NAND2_X1 U14947 ( .A1(n14712), .A2(n14890), .ZN(n14889) );
  NAND2_X1 U14948 ( .A1(n14711), .A2(n14710), .ZN(n14890) );
  NOR2_X1 U14949 ( .A1(n7645), .A2(n8062), .ZN(n14712) );
  OR2_X1 U14950 ( .A1(n14710), .A2(n14711), .ZN(n14888) );
  AND2_X1 U14951 ( .A1(n14891), .A2(n14892), .ZN(n14711) );
  NAND2_X1 U14952 ( .A1(n14707), .A2(n14893), .ZN(n14892) );
  OR2_X1 U14953 ( .A1(n14706), .A2(n14708), .ZN(n14893) );
  NOR2_X1 U14954 ( .A1(n8062), .A2(n7624), .ZN(n14707) );
  NAND2_X1 U14955 ( .A1(n14706), .A2(n14708), .ZN(n14891) );
  NAND2_X1 U14956 ( .A1(n14894), .A2(n14895), .ZN(n14708) );
  NAND2_X1 U14957 ( .A1(n14704), .A2(n14896), .ZN(n14895) );
  OR2_X1 U14958 ( .A1(n14701), .A2(n14703), .ZN(n14896) );
  NOR2_X1 U14959 ( .A1(n8062), .A2(n7613), .ZN(n14704) );
  NAND2_X1 U14960 ( .A1(n14701), .A2(n14703), .ZN(n14894) );
  NAND2_X1 U14961 ( .A1(n14897), .A2(n14898), .ZN(n14703) );
  NAND2_X1 U14962 ( .A1(n14899), .A2(b_4_), .ZN(n14898) );
  NOR2_X1 U14963 ( .A1(n14900), .A2(n7593), .ZN(n14899) );
  NOR2_X1 U14964 ( .A1(n14658), .A2(n14657), .ZN(n14900) );
  NAND2_X1 U14965 ( .A1(n14657), .A2(n14658), .ZN(n14897) );
  NAND2_X1 U14966 ( .A1(n14901), .A2(n14902), .ZN(n14658) );
  NAND2_X1 U14967 ( .A1(n14699), .A2(n14903), .ZN(n14902) );
  NAND2_X1 U14968 ( .A1(n14700), .A2(n14698), .ZN(n14903) );
  NOR2_X1 U14969 ( .A1(n8062), .A2(n8052), .ZN(n14699) );
  OR2_X1 U14970 ( .A1(n14698), .A2(n14700), .ZN(n14901) );
  AND2_X1 U14971 ( .A1(n14904), .A2(n14905), .ZN(n14700) );
  NAND2_X1 U14972 ( .A1(n14906), .A2(b_4_), .ZN(n14905) );
  NOR2_X1 U14973 ( .A1(n14907), .A2(n7563), .ZN(n14906) );
  NOR2_X1 U14974 ( .A1(n14695), .A2(n14693), .ZN(n14907) );
  NAND2_X1 U14975 ( .A1(n14693), .A2(n14695), .ZN(n14904) );
  NAND2_X1 U14976 ( .A1(n14691), .A2(n14908), .ZN(n14695) );
  NAND2_X1 U14977 ( .A1(n14690), .A2(n14692), .ZN(n14908) );
  NAND2_X1 U14978 ( .A1(n14909), .A2(n14910), .ZN(n14692) );
  NAND2_X1 U14979 ( .A1(b_4_), .A2(a_28_), .ZN(n14910) );
  INV_X1 U14980 ( .A(n14911), .ZN(n14909) );
  XOR2_X1 U14981 ( .A(n14912), .B(n14913), .Z(n14690) );
  NOR2_X1 U14982 ( .A1(n7529), .A2(n7946), .ZN(n14913) );
  XOR2_X1 U14983 ( .A(n14914), .B(n14915), .Z(n14912) );
  NAND2_X1 U14984 ( .A1(a_28_), .A2(n14911), .ZN(n14691) );
  NAND2_X1 U14985 ( .A1(n14916), .A2(n14917), .ZN(n14911) );
  NAND2_X1 U14986 ( .A1(n14918), .A2(b_4_), .ZN(n14917) );
  NOR2_X1 U14987 ( .A1(n14919), .A2(n7529), .ZN(n14918) );
  NOR2_X1 U14988 ( .A1(n14676), .A2(n14677), .ZN(n14919) );
  NAND2_X1 U14989 ( .A1(n14676), .A2(n14677), .ZN(n14916) );
  NAND2_X1 U14990 ( .A1(n14920), .A2(n14921), .ZN(n14677) );
  NAND2_X1 U14991 ( .A1(n14922), .A2(b_2_), .ZN(n14921) );
  NOR2_X1 U14992 ( .A1(n14923), .A2(n8048), .ZN(n14922) );
  NOR2_X1 U14993 ( .A1(n8676), .A2(n7946), .ZN(n14923) );
  NAND2_X1 U14994 ( .A1(n14924), .A2(b_3_), .ZN(n14920) );
  NOR2_X1 U14995 ( .A1(n14925), .A2(n7515), .ZN(n14924) );
  NOR2_X1 U14996 ( .A1(n8679), .A2(n8063), .ZN(n14925) );
  AND2_X1 U14997 ( .A1(n14926), .A2(b_3_), .ZN(n14676) );
  NOR2_X1 U14998 ( .A1(n8451), .A2(n8062), .ZN(n14926) );
  XNOR2_X1 U14999 ( .A(n14927), .B(n14928), .ZN(n14693) );
  XNOR2_X1 U15000 ( .A(n14929), .B(n14930), .ZN(n14927) );
  XOR2_X1 U15001 ( .A(n14931), .B(n14932), .Z(n14698) );
  XOR2_X1 U15002 ( .A(n14933), .B(n14934), .Z(n14932) );
  NAND2_X1 U15003 ( .A1(b_3_), .A2(a_27_), .ZN(n14934) );
  XNOR2_X1 U15004 ( .A(n14935), .B(n14936), .ZN(n14657) );
  XOR2_X1 U15005 ( .A(n14937), .B(n14938), .Z(n14936) );
  NAND2_X1 U15006 ( .A1(b_3_), .A2(a_26_), .ZN(n14938) );
  XNOR2_X1 U15007 ( .A(n14939), .B(n14940), .ZN(n14701) );
  XOR2_X1 U15008 ( .A(n14941), .B(n14942), .Z(n14940) );
  NAND2_X1 U15009 ( .A1(b_3_), .A2(a_25_), .ZN(n14942) );
  XNOR2_X1 U15010 ( .A(n14943), .B(n14944), .ZN(n14706) );
  NAND2_X1 U15011 ( .A1(n14945), .A2(n14946), .ZN(n14943) );
  XNOR2_X1 U15012 ( .A(n14947), .B(n14948), .ZN(n14710) );
  XOR2_X1 U15013 ( .A(n14949), .B(n14950), .Z(n14947) );
  NOR2_X1 U15014 ( .A1(n7624), .A2(n7946), .ZN(n14950) );
  XNOR2_X1 U15015 ( .A(n14951), .B(n14952), .ZN(n14713) );
  NAND2_X1 U15016 ( .A1(n14953), .A2(n14954), .ZN(n14951) );
  XNOR2_X1 U15017 ( .A(n14955), .B(n14956), .ZN(n14718) );
  XOR2_X1 U15018 ( .A(n14957), .B(n14958), .Z(n14955) );
  NOR2_X1 U15019 ( .A1(n7656), .A2(n7946), .ZN(n14958) );
  XNOR2_X1 U15020 ( .A(n14959), .B(n14960), .ZN(n14721) );
  NAND2_X1 U15021 ( .A1(n14961), .A2(n14962), .ZN(n14959) );
  XNOR2_X1 U15022 ( .A(n14963), .B(n14964), .ZN(n14726) );
  XOR2_X1 U15023 ( .A(n14965), .B(n14966), .Z(n14963) );
  NOR2_X1 U15024 ( .A1(n7946), .A2(n7687), .ZN(n14966) );
  XNOR2_X1 U15025 ( .A(n14967), .B(n14968), .ZN(n14729) );
  NAND2_X1 U15026 ( .A1(n14969), .A2(n14970), .ZN(n14967) );
  XNOR2_X1 U15027 ( .A(n14971), .B(n14972), .ZN(n14734) );
  XOR2_X1 U15028 ( .A(n14973), .B(n14974), .Z(n14971) );
  NOR2_X1 U15029 ( .A1(n7946), .A2(n7723), .ZN(n14974) );
  XNOR2_X1 U15030 ( .A(n14975), .B(n14976), .ZN(n14737) );
  NAND2_X1 U15031 ( .A1(n14977), .A2(n14978), .ZN(n14975) );
  XOR2_X1 U15032 ( .A(n14979), .B(n14980), .Z(n14742) );
  XOR2_X1 U15033 ( .A(n14981), .B(n14982), .Z(n14979) );
  NOR2_X1 U15034 ( .A1(n7946), .A2(n7754), .ZN(n14982) );
  XNOR2_X1 U15035 ( .A(n14983), .B(n14984), .ZN(n14745) );
  NAND2_X1 U15036 ( .A1(n14985), .A2(n14986), .ZN(n14983) );
  XOR2_X1 U15037 ( .A(n14987), .B(n14988), .Z(n14749) );
  XOR2_X1 U15038 ( .A(n14989), .B(n14990), .Z(n14987) );
  NOR2_X1 U15039 ( .A1(n7946), .A2(n7786), .ZN(n14990) );
  XNOR2_X1 U15040 ( .A(n14991), .B(n14992), .ZN(n14753) );
  NAND2_X1 U15041 ( .A1(n14993), .A2(n14994), .ZN(n14991) );
  XOR2_X1 U15042 ( .A(n14995), .B(n14996), .Z(n14757) );
  XOR2_X1 U15043 ( .A(n14997), .B(n14998), .Z(n14995) );
  NOR2_X1 U15044 ( .A1(n7817), .A2(n7946), .ZN(n14998) );
  XNOR2_X1 U15045 ( .A(n14999), .B(n15000), .ZN(n14761) );
  NAND2_X1 U15046 ( .A1(n15001), .A2(n15002), .ZN(n14999) );
  XOR2_X1 U15047 ( .A(n15003), .B(n15004), .Z(n14765) );
  XOR2_X1 U15048 ( .A(n15005), .B(n15006), .Z(n15003) );
  NOR2_X1 U15049 ( .A1(n7946), .A2(n7848), .ZN(n15006) );
  XNOR2_X1 U15050 ( .A(n15007), .B(n15008), .ZN(n14769) );
  NAND2_X1 U15051 ( .A1(n15009), .A2(n15010), .ZN(n15007) );
  XOR2_X1 U15052 ( .A(n15011), .B(n15012), .Z(n14576) );
  XOR2_X1 U15053 ( .A(n15013), .B(n15014), .Z(n15011) );
  NOR2_X1 U15054 ( .A1(n7946), .A2(n7884), .ZN(n15014) );
  XNOR2_X1 U15055 ( .A(n15015), .B(n15016), .ZN(n14773) );
  NAND2_X1 U15056 ( .A1(n15017), .A2(n15018), .ZN(n15015) );
  INV_X1 U15057 ( .A(n7928), .ZN(n14780) );
  NAND2_X1 U15058 ( .A1(a_4_), .A2(b_4_), .ZN(n7928) );
  XNOR2_X1 U15059 ( .A(n15019), .B(n15020), .ZN(n14782) );
  NAND2_X1 U15060 ( .A1(n15021), .A2(n15022), .ZN(n15019) );
  XOR2_X1 U15061 ( .A(n15023), .B(n15024), .Z(n14786) );
  XOR2_X1 U15062 ( .A(n15025), .B(n7940), .Z(n15023) );
  XNOR2_X1 U15063 ( .A(n15026), .B(n15027), .ZN(n14790) );
  NAND2_X1 U15064 ( .A1(n15028), .A2(n15029), .ZN(n15026) );
  XOR2_X1 U15065 ( .A(n15030), .B(n15031), .Z(n14794) );
  XOR2_X1 U15066 ( .A(n15032), .B(n15033), .Z(n15030) );
  NOR2_X1 U15067 ( .A1(n7946), .A2(n7973), .ZN(n15033) );
  NOR2_X1 U15068 ( .A1(n15034), .A2(n14551), .ZN(n14803) );
  INV_X1 U15069 ( .A(n14553), .ZN(n14551) );
  XOR2_X1 U15070 ( .A(n15035), .B(n15036), .Z(n14553) );
  XOR2_X1 U15071 ( .A(n15037), .B(n15038), .Z(n15035) );
  NOR2_X1 U15072 ( .A1(n14802), .A2(n14801), .ZN(n15034) );
  NAND2_X1 U15073 ( .A1(n15039), .A2(n14800), .ZN(n8082) );
  XNOR2_X1 U15074 ( .A(n8194), .B(n8195), .ZN(n15039) );
  NAND2_X1 U15075 ( .A1(n15040), .A2(n15041), .ZN(n8081) );
  XOR2_X1 U15076 ( .A(n8194), .B(n8195), .Z(n15041) );
  INV_X1 U15077 ( .A(n14800), .ZN(n15040) );
  NAND2_X1 U15078 ( .A1(n14802), .A2(n14801), .ZN(n14800) );
  NAND2_X1 U15079 ( .A1(n15042), .A2(n15043), .ZN(n14801) );
  NAND2_X1 U15080 ( .A1(n15038), .A2(n15044), .ZN(n15043) );
  OR2_X1 U15081 ( .A1(n15036), .A2(n15037), .ZN(n15044) );
  NOR2_X1 U15082 ( .A1(n7946), .A2(n8307), .ZN(n15038) );
  NAND2_X1 U15083 ( .A1(n15036), .A2(n15037), .ZN(n15042) );
  NAND2_X1 U15084 ( .A1(n15045), .A2(n15046), .ZN(n15037) );
  NAND2_X1 U15085 ( .A1(n15047), .A2(a_1_), .ZN(n15046) );
  NOR2_X1 U15086 ( .A1(n15048), .A2(n7946), .ZN(n15047) );
  NOR2_X1 U15087 ( .A1(n15032), .A2(n15031), .ZN(n15048) );
  NAND2_X1 U15088 ( .A1(n15031), .A2(n15032), .ZN(n15045) );
  NAND2_X1 U15089 ( .A1(n15028), .A2(n15049), .ZN(n15032) );
  NAND2_X1 U15090 ( .A1(n15027), .A2(n15029), .ZN(n15049) );
  NAND2_X1 U15091 ( .A1(n15050), .A2(n15051), .ZN(n15029) );
  NAND2_X1 U15092 ( .A1(a_2_), .A2(b_3_), .ZN(n15051) );
  INV_X1 U15093 ( .A(n15052), .ZN(n15050) );
  XNOR2_X1 U15094 ( .A(n15053), .B(n15054), .ZN(n15027) );
  XNOR2_X1 U15095 ( .A(n15055), .B(n15056), .ZN(n15053) );
  NAND2_X1 U15096 ( .A1(a_2_), .A2(n15052), .ZN(n15028) );
  NAND2_X1 U15097 ( .A1(n15057), .A2(n15058), .ZN(n15052) );
  NAND2_X1 U15098 ( .A1(n15024), .A2(n15059), .ZN(n15058) );
  OR2_X1 U15099 ( .A1(n15025), .A2(n7940), .ZN(n15059) );
  XNOR2_X1 U15100 ( .A(n15060), .B(n15061), .ZN(n15024) );
  NAND2_X1 U15101 ( .A1(n15062), .A2(n15063), .ZN(n15060) );
  NAND2_X1 U15102 ( .A1(n7940), .A2(n15025), .ZN(n15057) );
  NAND2_X1 U15103 ( .A1(n15021), .A2(n15064), .ZN(n15025) );
  NAND2_X1 U15104 ( .A1(n15020), .A2(n15022), .ZN(n15064) );
  NAND2_X1 U15105 ( .A1(n15065), .A2(n15066), .ZN(n15022) );
  NAND2_X1 U15106 ( .A1(a_4_), .A2(b_3_), .ZN(n15066) );
  INV_X1 U15107 ( .A(n15067), .ZN(n15065) );
  XNOR2_X1 U15108 ( .A(n15068), .B(n15069), .ZN(n15020) );
  XNOR2_X1 U15109 ( .A(n15070), .B(n15071), .ZN(n15068) );
  NAND2_X1 U15110 ( .A1(a_4_), .A2(n15067), .ZN(n15021) );
  NAND2_X1 U15111 ( .A1(n15072), .A2(n15073), .ZN(n15067) );
  NAND2_X1 U15112 ( .A1(n15074), .A2(a_5_), .ZN(n15073) );
  NOR2_X1 U15113 ( .A1(n15075), .A2(n7946), .ZN(n15074) );
  NOR2_X1 U15114 ( .A1(n14825), .A2(n14826), .ZN(n15075) );
  NAND2_X1 U15115 ( .A1(n14825), .A2(n14826), .ZN(n15072) );
  NAND2_X1 U15116 ( .A1(n15017), .A2(n15076), .ZN(n14826) );
  NAND2_X1 U15117 ( .A1(n15016), .A2(n15018), .ZN(n15076) );
  NAND2_X1 U15118 ( .A1(n15077), .A2(n15078), .ZN(n15018) );
  NAND2_X1 U15119 ( .A1(a_6_), .A2(b_3_), .ZN(n15078) );
  INV_X1 U15120 ( .A(n15079), .ZN(n15077) );
  XNOR2_X1 U15121 ( .A(n15080), .B(n15081), .ZN(n15016) );
  XNOR2_X1 U15122 ( .A(n15082), .B(n15083), .ZN(n15080) );
  NAND2_X1 U15123 ( .A1(a_6_), .A2(n15079), .ZN(n15017) );
  NAND2_X1 U15124 ( .A1(n15084), .A2(n15085), .ZN(n15079) );
  NAND2_X1 U15125 ( .A1(n15086), .A2(a_7_), .ZN(n15085) );
  NOR2_X1 U15126 ( .A1(n15087), .A2(n7946), .ZN(n15086) );
  NOR2_X1 U15127 ( .A1(n15012), .A2(n15013), .ZN(n15087) );
  NAND2_X1 U15128 ( .A1(n15012), .A2(n15013), .ZN(n15084) );
  NAND2_X1 U15129 ( .A1(n15009), .A2(n15088), .ZN(n15013) );
  NAND2_X1 U15130 ( .A1(n15008), .A2(n15010), .ZN(n15088) );
  NAND2_X1 U15131 ( .A1(n15089), .A2(n15090), .ZN(n15010) );
  NAND2_X1 U15132 ( .A1(a_8_), .A2(b_3_), .ZN(n15090) );
  INV_X1 U15133 ( .A(n15091), .ZN(n15089) );
  XNOR2_X1 U15134 ( .A(n15092), .B(n15093), .ZN(n15008) );
  XNOR2_X1 U15135 ( .A(n15094), .B(n15095), .ZN(n15092) );
  NAND2_X1 U15136 ( .A1(a_8_), .A2(n15091), .ZN(n15009) );
  NAND2_X1 U15137 ( .A1(n15096), .A2(n15097), .ZN(n15091) );
  NAND2_X1 U15138 ( .A1(n15098), .A2(a_9_), .ZN(n15097) );
  NOR2_X1 U15139 ( .A1(n15099), .A2(n7946), .ZN(n15098) );
  NOR2_X1 U15140 ( .A1(n15004), .A2(n15005), .ZN(n15099) );
  NAND2_X1 U15141 ( .A1(n15004), .A2(n15005), .ZN(n15096) );
  NAND2_X1 U15142 ( .A1(n15001), .A2(n15100), .ZN(n15005) );
  NAND2_X1 U15143 ( .A1(n15000), .A2(n15002), .ZN(n15100) );
  NAND2_X1 U15144 ( .A1(n15101), .A2(n15102), .ZN(n15002) );
  NAND2_X1 U15145 ( .A1(a_10_), .A2(b_3_), .ZN(n15102) );
  INV_X1 U15146 ( .A(n15103), .ZN(n15101) );
  XNOR2_X1 U15147 ( .A(n15104), .B(n15105), .ZN(n15000) );
  XNOR2_X1 U15148 ( .A(n15106), .B(n15107), .ZN(n15104) );
  NAND2_X1 U15149 ( .A1(a_10_), .A2(n15103), .ZN(n15001) );
  NAND2_X1 U15150 ( .A1(n15108), .A2(n15109), .ZN(n15103) );
  NAND2_X1 U15151 ( .A1(n15110), .A2(b_3_), .ZN(n15109) );
  NOR2_X1 U15152 ( .A1(n15111), .A2(n7817), .ZN(n15110) );
  NOR2_X1 U15153 ( .A1(n14996), .A2(n14997), .ZN(n15111) );
  NAND2_X1 U15154 ( .A1(n14996), .A2(n14997), .ZN(n15108) );
  NAND2_X1 U15155 ( .A1(n14993), .A2(n15112), .ZN(n14997) );
  NAND2_X1 U15156 ( .A1(n14992), .A2(n14994), .ZN(n15112) );
  NAND2_X1 U15157 ( .A1(n15113), .A2(n15114), .ZN(n14994) );
  NAND2_X1 U15158 ( .A1(a_12_), .A2(b_3_), .ZN(n15114) );
  INV_X1 U15159 ( .A(n15115), .ZN(n15113) );
  XNOR2_X1 U15160 ( .A(n15116), .B(n15117), .ZN(n14992) );
  XNOR2_X1 U15161 ( .A(n15118), .B(n15119), .ZN(n15116) );
  NAND2_X1 U15162 ( .A1(a_12_), .A2(n15115), .ZN(n14993) );
  NAND2_X1 U15163 ( .A1(n15120), .A2(n15121), .ZN(n15115) );
  NAND2_X1 U15164 ( .A1(n15122), .A2(a_13_), .ZN(n15121) );
  NOR2_X1 U15165 ( .A1(n15123), .A2(n7946), .ZN(n15122) );
  NOR2_X1 U15166 ( .A1(n14988), .A2(n14989), .ZN(n15123) );
  NAND2_X1 U15167 ( .A1(n14988), .A2(n14989), .ZN(n15120) );
  NAND2_X1 U15168 ( .A1(n14985), .A2(n15124), .ZN(n14989) );
  NAND2_X1 U15169 ( .A1(n14984), .A2(n14986), .ZN(n15124) );
  NAND2_X1 U15170 ( .A1(n15125), .A2(n15126), .ZN(n14986) );
  NAND2_X1 U15171 ( .A1(a_14_), .A2(b_3_), .ZN(n15126) );
  INV_X1 U15172 ( .A(n15127), .ZN(n15125) );
  XNOR2_X1 U15173 ( .A(n15128), .B(n15129), .ZN(n14984) );
  XNOR2_X1 U15174 ( .A(n15130), .B(n15131), .ZN(n15128) );
  NAND2_X1 U15175 ( .A1(a_14_), .A2(n15127), .ZN(n14985) );
  NAND2_X1 U15176 ( .A1(n15132), .A2(n15133), .ZN(n15127) );
  NAND2_X1 U15177 ( .A1(n15134), .A2(a_15_), .ZN(n15133) );
  NOR2_X1 U15178 ( .A1(n15135), .A2(n7946), .ZN(n15134) );
  NOR2_X1 U15179 ( .A1(n14980), .A2(n14981), .ZN(n15135) );
  NAND2_X1 U15180 ( .A1(n14980), .A2(n14981), .ZN(n15132) );
  NAND2_X1 U15181 ( .A1(n14977), .A2(n15136), .ZN(n14981) );
  NAND2_X1 U15182 ( .A1(n14976), .A2(n14978), .ZN(n15136) );
  NAND2_X1 U15183 ( .A1(n15137), .A2(n15138), .ZN(n14978) );
  NAND2_X1 U15184 ( .A1(a_16_), .A2(b_3_), .ZN(n15138) );
  INV_X1 U15185 ( .A(n15139), .ZN(n15137) );
  XOR2_X1 U15186 ( .A(n15140), .B(n15141), .Z(n14976) );
  XNOR2_X1 U15187 ( .A(n15142), .B(n15143), .ZN(n15140) );
  NAND2_X1 U15188 ( .A1(a_17_), .A2(b_2_), .ZN(n15142) );
  NAND2_X1 U15189 ( .A1(a_16_), .A2(n15139), .ZN(n14977) );
  NAND2_X1 U15190 ( .A1(n15144), .A2(n15145), .ZN(n15139) );
  NAND2_X1 U15191 ( .A1(n15146), .A2(a_17_), .ZN(n15145) );
  NOR2_X1 U15192 ( .A1(n15147), .A2(n7946), .ZN(n15146) );
  NOR2_X1 U15193 ( .A1(n14973), .A2(n14972), .ZN(n15147) );
  NAND2_X1 U15194 ( .A1(n14972), .A2(n14973), .ZN(n15144) );
  NAND2_X1 U15195 ( .A1(n14969), .A2(n15148), .ZN(n14973) );
  NAND2_X1 U15196 ( .A1(n14968), .A2(n14970), .ZN(n15148) );
  NAND2_X1 U15197 ( .A1(n15149), .A2(n15150), .ZN(n14970) );
  NAND2_X1 U15198 ( .A1(a_18_), .A2(b_3_), .ZN(n15150) );
  INV_X1 U15199 ( .A(n15151), .ZN(n15149) );
  XOR2_X1 U15200 ( .A(n15152), .B(n15153), .Z(n14968) );
  XOR2_X1 U15201 ( .A(n15154), .B(n15155), .Z(n15152) );
  NOR2_X1 U15202 ( .A1(n8063), .A2(n7687), .ZN(n15155) );
  NAND2_X1 U15203 ( .A1(a_18_), .A2(n15151), .ZN(n14969) );
  NAND2_X1 U15204 ( .A1(n15156), .A2(n15157), .ZN(n15151) );
  NAND2_X1 U15205 ( .A1(n15158), .A2(a_19_), .ZN(n15157) );
  NOR2_X1 U15206 ( .A1(n15159), .A2(n7946), .ZN(n15158) );
  NOR2_X1 U15207 ( .A1(n14965), .A2(n14964), .ZN(n15159) );
  NAND2_X1 U15208 ( .A1(n14964), .A2(n14965), .ZN(n15156) );
  NAND2_X1 U15209 ( .A1(n14961), .A2(n15160), .ZN(n14965) );
  NAND2_X1 U15210 ( .A1(n14960), .A2(n14962), .ZN(n15160) );
  NAND2_X1 U15211 ( .A1(n15161), .A2(n15162), .ZN(n14962) );
  NAND2_X1 U15212 ( .A1(b_3_), .A2(a_20_), .ZN(n15162) );
  INV_X1 U15213 ( .A(n15163), .ZN(n15161) );
  XOR2_X1 U15214 ( .A(n15164), .B(n15165), .Z(n14960) );
  XNOR2_X1 U15215 ( .A(n15166), .B(n15167), .ZN(n15164) );
  NAND2_X1 U15216 ( .A1(b_2_), .A2(a_21_), .ZN(n15166) );
  NAND2_X1 U15217 ( .A1(a_20_), .A2(n15163), .ZN(n14961) );
  NAND2_X1 U15218 ( .A1(n15168), .A2(n15169), .ZN(n15163) );
  NAND2_X1 U15219 ( .A1(n15170), .A2(b_3_), .ZN(n15169) );
  NOR2_X1 U15220 ( .A1(n15171), .A2(n7656), .ZN(n15170) );
  NOR2_X1 U15221 ( .A1(n14957), .A2(n14956), .ZN(n15171) );
  NAND2_X1 U15222 ( .A1(n14956), .A2(n14957), .ZN(n15168) );
  NAND2_X1 U15223 ( .A1(n14953), .A2(n15172), .ZN(n14957) );
  NAND2_X1 U15224 ( .A1(n14952), .A2(n14954), .ZN(n15172) );
  NAND2_X1 U15225 ( .A1(n15173), .A2(n15174), .ZN(n14954) );
  NAND2_X1 U15226 ( .A1(a_22_), .A2(b_3_), .ZN(n15174) );
  INV_X1 U15227 ( .A(n15175), .ZN(n15173) );
  XNOR2_X1 U15228 ( .A(n15176), .B(n15177), .ZN(n14952) );
  XOR2_X1 U15229 ( .A(n15178), .B(n15179), .Z(n15177) );
  NAND2_X1 U15230 ( .A1(b_2_), .A2(a_23_), .ZN(n15179) );
  NAND2_X1 U15231 ( .A1(a_22_), .A2(n15175), .ZN(n14953) );
  NAND2_X1 U15232 ( .A1(n15180), .A2(n15181), .ZN(n15175) );
  NAND2_X1 U15233 ( .A1(n15182), .A2(b_3_), .ZN(n15181) );
  NOR2_X1 U15234 ( .A1(n15183), .A2(n7624), .ZN(n15182) );
  NOR2_X1 U15235 ( .A1(n14949), .A2(n14948), .ZN(n15183) );
  NAND2_X1 U15236 ( .A1(n14948), .A2(n14949), .ZN(n15180) );
  NAND2_X1 U15237 ( .A1(n14945), .A2(n15184), .ZN(n14949) );
  NAND2_X1 U15238 ( .A1(n14944), .A2(n14946), .ZN(n15184) );
  NAND2_X1 U15239 ( .A1(n15185), .A2(n15186), .ZN(n14946) );
  NAND2_X1 U15240 ( .A1(b_3_), .A2(a_24_), .ZN(n15186) );
  INV_X1 U15241 ( .A(n15187), .ZN(n15185) );
  XNOR2_X1 U15242 ( .A(n15188), .B(n15189), .ZN(n14944) );
  XNOR2_X1 U15243 ( .A(n15190), .B(n15191), .ZN(n15189) );
  NAND2_X1 U15244 ( .A1(a_24_), .A2(n15187), .ZN(n14945) );
  NAND2_X1 U15245 ( .A1(n15192), .A2(n15193), .ZN(n15187) );
  NAND2_X1 U15246 ( .A1(n15194), .A2(b_3_), .ZN(n15193) );
  NOR2_X1 U15247 ( .A1(n15195), .A2(n7593), .ZN(n15194) );
  NOR2_X1 U15248 ( .A1(n14939), .A2(n14941), .ZN(n15195) );
  NAND2_X1 U15249 ( .A1(n14939), .A2(n14941), .ZN(n15192) );
  NAND2_X1 U15250 ( .A1(n15196), .A2(n15197), .ZN(n14941) );
  NAND2_X1 U15251 ( .A1(n15198), .A2(b_3_), .ZN(n15197) );
  NOR2_X1 U15252 ( .A1(n15199), .A2(n8052), .ZN(n15198) );
  NOR2_X1 U15253 ( .A1(n14935), .A2(n14937), .ZN(n15199) );
  NAND2_X1 U15254 ( .A1(n14935), .A2(n14937), .ZN(n15196) );
  NAND2_X1 U15255 ( .A1(n15200), .A2(n15201), .ZN(n14937) );
  NAND2_X1 U15256 ( .A1(n15202), .A2(b_3_), .ZN(n15201) );
  NOR2_X1 U15257 ( .A1(n15203), .A2(n7563), .ZN(n15202) );
  NOR2_X1 U15258 ( .A1(n14933), .A2(n14931), .ZN(n15203) );
  NAND2_X1 U15259 ( .A1(n14931), .A2(n14933), .ZN(n15200) );
  NAND2_X1 U15260 ( .A1(n15204), .A2(n15205), .ZN(n14933) );
  NAND2_X1 U15261 ( .A1(n14929), .A2(n15206), .ZN(n15205) );
  NAND2_X1 U15262 ( .A1(n14930), .A2(n14928), .ZN(n15206) );
  NOR2_X1 U15263 ( .A1(n7946), .A2(n7547), .ZN(n14929) );
  OR2_X1 U15264 ( .A1(n14928), .A2(n14930), .ZN(n15204) );
  AND2_X1 U15265 ( .A1(n15207), .A2(n15208), .ZN(n14930) );
  NAND2_X1 U15266 ( .A1(n15209), .A2(b_3_), .ZN(n15208) );
  NOR2_X1 U15267 ( .A1(n15210), .A2(n7529), .ZN(n15209) );
  NOR2_X1 U15268 ( .A1(n14914), .A2(n14915), .ZN(n15210) );
  NAND2_X1 U15269 ( .A1(n14914), .A2(n14915), .ZN(n15207) );
  NAND2_X1 U15270 ( .A1(n15211), .A2(n15212), .ZN(n14915) );
  NAND2_X1 U15271 ( .A1(n15213), .A2(b_1_), .ZN(n15212) );
  NOR2_X1 U15272 ( .A1(n15214), .A2(n8048), .ZN(n15213) );
  NOR2_X1 U15273 ( .A1(n8676), .A2(n8063), .ZN(n15214) );
  NAND2_X1 U15274 ( .A1(n15215), .A2(b_2_), .ZN(n15211) );
  NOR2_X1 U15275 ( .A1(n15216), .A2(n7515), .ZN(n15215) );
  NOR2_X1 U15276 ( .A1(n8679), .A2(n15217), .ZN(n15216) );
  AND2_X1 U15277 ( .A1(n15218), .A2(b_2_), .ZN(n14914) );
  NOR2_X1 U15278 ( .A1(n8451), .A2(n7946), .ZN(n15218) );
  XNOR2_X1 U15279 ( .A(n15219), .B(n15220), .ZN(n14928) );
  NOR2_X1 U15280 ( .A1(n7529), .A2(n8063), .ZN(n15220) );
  XOR2_X1 U15281 ( .A(n15221), .B(n15222), .Z(n15219) );
  XNOR2_X1 U15282 ( .A(n15223), .B(n15224), .ZN(n14931) );
  NAND2_X1 U15283 ( .A1(n15225), .A2(n15226), .ZN(n15223) );
  XNOR2_X1 U15284 ( .A(n15227), .B(n15228), .ZN(n14935) );
  NAND2_X1 U15285 ( .A1(n15229), .A2(n15230), .ZN(n15227) );
  XNOR2_X1 U15286 ( .A(n15231), .B(n15232), .ZN(n14939) );
  NAND2_X1 U15287 ( .A1(n15233), .A2(n15234), .ZN(n15231) );
  XNOR2_X1 U15288 ( .A(n15235), .B(n15236), .ZN(n14948) );
  XNOR2_X1 U15289 ( .A(n15237), .B(n15238), .ZN(n15236) );
  XNOR2_X1 U15290 ( .A(n15239), .B(n15240), .ZN(n14956) );
  XNOR2_X1 U15291 ( .A(n15241), .B(n15242), .ZN(n15239) );
  XNOR2_X1 U15292 ( .A(n15243), .B(n15244), .ZN(n14964) );
  XNOR2_X1 U15293 ( .A(n15245), .B(n15246), .ZN(n15243) );
  XNOR2_X1 U15294 ( .A(n15247), .B(n15248), .ZN(n14972) );
  XNOR2_X1 U15295 ( .A(n15249), .B(n15250), .ZN(n15247) );
  XNOR2_X1 U15296 ( .A(n15251), .B(n15252), .ZN(n14980) );
  NAND2_X1 U15297 ( .A1(n15253), .A2(n15254), .ZN(n15251) );
  XNOR2_X1 U15298 ( .A(n15255), .B(n15256), .ZN(n14988) );
  NAND2_X1 U15299 ( .A1(n15257), .A2(n15258), .ZN(n15255) );
  XNOR2_X1 U15300 ( .A(n15259), .B(n15260), .ZN(n14996) );
  NAND2_X1 U15301 ( .A1(n15261), .A2(n15262), .ZN(n15259) );
  XNOR2_X1 U15302 ( .A(n15263), .B(n15264), .ZN(n15004) );
  NAND2_X1 U15303 ( .A1(n15265), .A2(n15266), .ZN(n15263) );
  XNOR2_X1 U15304 ( .A(n15267), .B(n15268), .ZN(n15012) );
  NAND2_X1 U15305 ( .A1(n15269), .A2(n15270), .ZN(n15267) );
  XNOR2_X1 U15306 ( .A(n15271), .B(n15272), .ZN(n14825) );
  NAND2_X1 U15307 ( .A1(n15273), .A2(n15274), .ZN(n15271) );
  INV_X1 U15308 ( .A(n7992), .ZN(n7940) );
  NAND2_X1 U15309 ( .A1(a_3_), .A2(b_3_), .ZN(n7992) );
  XOR2_X1 U15310 ( .A(n15275), .B(n15276), .Z(n15031) );
  XOR2_X1 U15311 ( .A(n7959), .B(n15277), .Z(n15275) );
  XOR2_X1 U15312 ( .A(n15278), .B(n15279), .Z(n15036) );
  XOR2_X1 U15313 ( .A(n15280), .B(n15281), .Z(n15278) );
  XNOR2_X1 U15314 ( .A(n15282), .B(n15283), .ZN(n14802) );
  NAND2_X1 U15315 ( .A1(n15284), .A2(n15285), .ZN(n15282) );
  NAND2_X1 U15316 ( .A1(n15286), .A2(n15287), .ZN(n8136) );
  NAND2_X1 U15317 ( .A1(n8195), .A2(n8194), .ZN(n15287) );
  NAND2_X1 U15318 ( .A1(n15284), .A2(n15288), .ZN(n8194) );
  NAND2_X1 U15319 ( .A1(n15283), .A2(n15285), .ZN(n15288) );
  NAND2_X1 U15320 ( .A1(n15289), .A2(n15290), .ZN(n15285) );
  NAND2_X1 U15321 ( .A1(b_2_), .A2(a_0_), .ZN(n15290) );
  INV_X1 U15322 ( .A(n15291), .ZN(n15289) );
  XOR2_X1 U15323 ( .A(n15292), .B(n15293), .Z(n15283) );
  NOR2_X1 U15324 ( .A1(n15294), .A2(n7965), .ZN(n15293) );
  XOR2_X1 U15325 ( .A(n15295), .B(n7979), .Z(n15292) );
  NAND2_X1 U15326 ( .A1(a_0_), .A2(n15291), .ZN(n15284) );
  NAND2_X1 U15327 ( .A1(n15296), .A2(n15297), .ZN(n15291) );
  NAND2_X1 U15328 ( .A1(n15281), .A2(n15298), .ZN(n15297) );
  OR2_X1 U15329 ( .A1(n15280), .A2(n15279), .ZN(n15298) );
  NOR2_X1 U15330 ( .A1(n7973), .A2(n8063), .ZN(n15281) );
  NAND2_X1 U15331 ( .A1(n15279), .A2(n15280), .ZN(n15296) );
  NAND2_X1 U15332 ( .A1(n15299), .A2(n15300), .ZN(n15280) );
  NAND2_X1 U15333 ( .A1(n15276), .A2(n15301), .ZN(n15300) );
  NAND2_X1 U15334 ( .A1(n15277), .A2(n7959), .ZN(n15301) );
  XOR2_X1 U15335 ( .A(n15302), .B(n15303), .Z(n15276) );
  NOR2_X1 U15336 ( .A1(n15217), .A2(n7945), .ZN(n15303) );
  XOR2_X1 U15337 ( .A(n15304), .B(n15305), .Z(n15302) );
  OR2_X1 U15338 ( .A1(n7959), .A2(n15277), .ZN(n15299) );
  AND2_X1 U15339 ( .A1(n15306), .A2(n15307), .ZN(n15277) );
  NAND2_X1 U15340 ( .A1(n15056), .A2(n15308), .ZN(n15307) );
  NAND2_X1 U15341 ( .A1(n15055), .A2(n15054), .ZN(n15308) );
  NOR2_X1 U15342 ( .A1(n7945), .A2(n8063), .ZN(n15056) );
  OR2_X1 U15343 ( .A1(n15054), .A2(n15055), .ZN(n15306) );
  AND2_X1 U15344 ( .A1(n15062), .A2(n15309), .ZN(n15055) );
  NAND2_X1 U15345 ( .A1(n15061), .A2(n15063), .ZN(n15309) );
  NAND2_X1 U15346 ( .A1(n15310), .A2(n15311), .ZN(n15063) );
  NAND2_X1 U15347 ( .A1(a_4_), .A2(b_2_), .ZN(n15311) );
  INV_X1 U15348 ( .A(n15312), .ZN(n15310) );
  XOR2_X1 U15349 ( .A(n15313), .B(n15314), .Z(n15061) );
  NOR2_X1 U15350 ( .A1(n15217), .A2(n7914), .ZN(n15314) );
  XOR2_X1 U15351 ( .A(n15315), .B(n15316), .Z(n15313) );
  NAND2_X1 U15352 ( .A1(a_4_), .A2(n15312), .ZN(n15062) );
  NAND2_X1 U15353 ( .A1(n15317), .A2(n15318), .ZN(n15312) );
  NAND2_X1 U15354 ( .A1(n15071), .A2(n15319), .ZN(n15318) );
  NAND2_X1 U15355 ( .A1(n15070), .A2(n15069), .ZN(n15319) );
  NOR2_X1 U15356 ( .A1(n7914), .A2(n8063), .ZN(n15071) );
  OR2_X1 U15357 ( .A1(n15069), .A2(n15070), .ZN(n15317) );
  AND2_X1 U15358 ( .A1(n15273), .A2(n15320), .ZN(n15070) );
  NAND2_X1 U15359 ( .A1(n15272), .A2(n15274), .ZN(n15320) );
  NAND2_X1 U15360 ( .A1(n15321), .A2(n15322), .ZN(n15274) );
  NAND2_X1 U15361 ( .A1(a_6_), .A2(b_2_), .ZN(n15322) );
  INV_X1 U15362 ( .A(n15323), .ZN(n15321) );
  XOR2_X1 U15363 ( .A(n15324), .B(n15325), .Z(n15272) );
  NOR2_X1 U15364 ( .A1(n15217), .A2(n7884), .ZN(n15325) );
  XOR2_X1 U15365 ( .A(n15326), .B(n15327), .Z(n15324) );
  NAND2_X1 U15366 ( .A1(a_6_), .A2(n15323), .ZN(n15273) );
  NAND2_X1 U15367 ( .A1(n15328), .A2(n15329), .ZN(n15323) );
  NAND2_X1 U15368 ( .A1(n15083), .A2(n15330), .ZN(n15329) );
  NAND2_X1 U15369 ( .A1(n15082), .A2(n15081), .ZN(n15330) );
  NOR2_X1 U15370 ( .A1(n7884), .A2(n8063), .ZN(n15083) );
  OR2_X1 U15371 ( .A1(n15081), .A2(n15082), .ZN(n15328) );
  AND2_X1 U15372 ( .A1(n15269), .A2(n15331), .ZN(n15082) );
  NAND2_X1 U15373 ( .A1(n15268), .A2(n15270), .ZN(n15331) );
  NAND2_X1 U15374 ( .A1(n15332), .A2(n15333), .ZN(n15270) );
  NAND2_X1 U15375 ( .A1(a_8_), .A2(b_2_), .ZN(n15333) );
  INV_X1 U15376 ( .A(n15334), .ZN(n15332) );
  XOR2_X1 U15377 ( .A(n15335), .B(n15336), .Z(n15268) );
  NOR2_X1 U15378 ( .A1(n15217), .A2(n7848), .ZN(n15336) );
  XOR2_X1 U15379 ( .A(n15337), .B(n15338), .Z(n15335) );
  NAND2_X1 U15380 ( .A1(a_8_), .A2(n15334), .ZN(n15269) );
  NAND2_X1 U15381 ( .A1(n15339), .A2(n15340), .ZN(n15334) );
  NAND2_X1 U15382 ( .A1(n15095), .A2(n15341), .ZN(n15340) );
  NAND2_X1 U15383 ( .A1(n15094), .A2(n15093), .ZN(n15341) );
  NOR2_X1 U15384 ( .A1(n7848), .A2(n8063), .ZN(n15095) );
  OR2_X1 U15385 ( .A1(n15093), .A2(n15094), .ZN(n15339) );
  AND2_X1 U15386 ( .A1(n15265), .A2(n15342), .ZN(n15094) );
  NAND2_X1 U15387 ( .A1(n15264), .A2(n15266), .ZN(n15342) );
  NAND2_X1 U15388 ( .A1(n15343), .A2(n15344), .ZN(n15266) );
  NAND2_X1 U15389 ( .A1(a_10_), .A2(b_2_), .ZN(n15344) );
  INV_X1 U15390 ( .A(n15345), .ZN(n15343) );
  XOR2_X1 U15391 ( .A(n15346), .B(n15347), .Z(n15264) );
  NOR2_X1 U15392 ( .A1(n7817), .A2(n15217), .ZN(n15347) );
  XOR2_X1 U15393 ( .A(n15348), .B(n15349), .Z(n15346) );
  NAND2_X1 U15394 ( .A1(a_10_), .A2(n15345), .ZN(n15265) );
  NAND2_X1 U15395 ( .A1(n15350), .A2(n15351), .ZN(n15345) );
  NAND2_X1 U15396 ( .A1(n15107), .A2(n15352), .ZN(n15351) );
  NAND2_X1 U15397 ( .A1(n15106), .A2(n15105), .ZN(n15352) );
  NOR2_X1 U15398 ( .A1(n8063), .A2(n7817), .ZN(n15107) );
  OR2_X1 U15399 ( .A1(n15105), .A2(n15106), .ZN(n15350) );
  AND2_X1 U15400 ( .A1(n15261), .A2(n15353), .ZN(n15106) );
  NAND2_X1 U15401 ( .A1(n15260), .A2(n15262), .ZN(n15353) );
  NAND2_X1 U15402 ( .A1(n15354), .A2(n15355), .ZN(n15262) );
  NAND2_X1 U15403 ( .A1(a_12_), .A2(b_2_), .ZN(n15355) );
  INV_X1 U15404 ( .A(n15356), .ZN(n15354) );
  XOR2_X1 U15405 ( .A(n15357), .B(n15358), .Z(n15260) );
  NOR2_X1 U15406 ( .A1(n15217), .A2(n7786), .ZN(n15358) );
  XOR2_X1 U15407 ( .A(n15359), .B(n15360), .Z(n15357) );
  NAND2_X1 U15408 ( .A1(a_12_), .A2(n15356), .ZN(n15261) );
  NAND2_X1 U15409 ( .A1(n15361), .A2(n15362), .ZN(n15356) );
  NAND2_X1 U15410 ( .A1(n15119), .A2(n15363), .ZN(n15362) );
  NAND2_X1 U15411 ( .A1(n15118), .A2(n15117), .ZN(n15363) );
  NOR2_X1 U15412 ( .A1(n7786), .A2(n8063), .ZN(n15119) );
  OR2_X1 U15413 ( .A1(n15117), .A2(n15118), .ZN(n15361) );
  AND2_X1 U15414 ( .A1(n15257), .A2(n15364), .ZN(n15118) );
  NAND2_X1 U15415 ( .A1(n15256), .A2(n15258), .ZN(n15364) );
  NAND2_X1 U15416 ( .A1(n15365), .A2(n15366), .ZN(n15258) );
  NAND2_X1 U15417 ( .A1(a_14_), .A2(b_2_), .ZN(n15366) );
  INV_X1 U15418 ( .A(n15367), .ZN(n15365) );
  XOR2_X1 U15419 ( .A(n15368), .B(n15369), .Z(n15256) );
  NOR2_X1 U15420 ( .A1(n15217), .A2(n7754), .ZN(n15369) );
  XOR2_X1 U15421 ( .A(n15370), .B(n15371), .Z(n15368) );
  NAND2_X1 U15422 ( .A1(a_14_), .A2(n15367), .ZN(n15257) );
  NAND2_X1 U15423 ( .A1(n15372), .A2(n15373), .ZN(n15367) );
  NAND2_X1 U15424 ( .A1(n15131), .A2(n15374), .ZN(n15373) );
  NAND2_X1 U15425 ( .A1(n15130), .A2(n15129), .ZN(n15374) );
  NOR2_X1 U15426 ( .A1(n7754), .A2(n8063), .ZN(n15131) );
  OR2_X1 U15427 ( .A1(n15129), .A2(n15130), .ZN(n15372) );
  AND2_X1 U15428 ( .A1(n15253), .A2(n15375), .ZN(n15130) );
  NAND2_X1 U15429 ( .A1(n15252), .A2(n15254), .ZN(n15375) );
  NAND2_X1 U15430 ( .A1(n15376), .A2(n15377), .ZN(n15254) );
  NAND2_X1 U15431 ( .A1(a_16_), .A2(b_2_), .ZN(n15377) );
  INV_X1 U15432 ( .A(n15378), .ZN(n15376) );
  XOR2_X1 U15433 ( .A(n15379), .B(n15380), .Z(n15252) );
  NOR2_X1 U15434 ( .A1(n15217), .A2(n7723), .ZN(n15380) );
  XOR2_X1 U15435 ( .A(n15381), .B(n15382), .Z(n15379) );
  NAND2_X1 U15436 ( .A1(a_16_), .A2(n15378), .ZN(n15253) );
  NAND2_X1 U15437 ( .A1(n15383), .A2(n15384), .ZN(n15378) );
  NAND2_X1 U15438 ( .A1(n15385), .A2(a_17_), .ZN(n15384) );
  NOR2_X1 U15439 ( .A1(n15386), .A2(n8063), .ZN(n15385) );
  NOR2_X1 U15440 ( .A1(n15141), .A2(n15143), .ZN(n15386) );
  NAND2_X1 U15441 ( .A1(n15141), .A2(n15143), .ZN(n15383) );
  NAND2_X1 U15442 ( .A1(n15387), .A2(n15388), .ZN(n15143) );
  NAND2_X1 U15443 ( .A1(n15250), .A2(n15389), .ZN(n15388) );
  NAND2_X1 U15444 ( .A1(n15249), .A2(n15248), .ZN(n15389) );
  NOR2_X1 U15445 ( .A1(n7707), .A2(n8063), .ZN(n15250) );
  OR2_X1 U15446 ( .A1(n15248), .A2(n15249), .ZN(n15387) );
  AND2_X1 U15447 ( .A1(n15390), .A2(n15391), .ZN(n15249) );
  NAND2_X1 U15448 ( .A1(n15392), .A2(a_19_), .ZN(n15391) );
  NOR2_X1 U15449 ( .A1(n15393), .A2(n8063), .ZN(n15392) );
  NOR2_X1 U15450 ( .A1(n15153), .A2(n15154), .ZN(n15393) );
  NAND2_X1 U15451 ( .A1(n15153), .A2(n15154), .ZN(n15390) );
  NAND2_X1 U15452 ( .A1(n15394), .A2(n15395), .ZN(n15154) );
  NAND2_X1 U15453 ( .A1(n15246), .A2(n15396), .ZN(n15395) );
  NAND2_X1 U15454 ( .A1(n15245), .A2(n15244), .ZN(n15396) );
  NOR2_X1 U15455 ( .A1(n8063), .A2(n7676), .ZN(n15246) );
  OR2_X1 U15456 ( .A1(n15244), .A2(n15245), .ZN(n15394) );
  AND2_X1 U15457 ( .A1(n15397), .A2(n15398), .ZN(n15245) );
  NAND2_X1 U15458 ( .A1(n15399), .A2(b_2_), .ZN(n15398) );
  NOR2_X1 U15459 ( .A1(n15400), .A2(n7656), .ZN(n15399) );
  NOR2_X1 U15460 ( .A1(n15165), .A2(n15167), .ZN(n15400) );
  NAND2_X1 U15461 ( .A1(n15165), .A2(n15167), .ZN(n15397) );
  NAND2_X1 U15462 ( .A1(n15401), .A2(n15402), .ZN(n15167) );
  NAND2_X1 U15463 ( .A1(n15242), .A2(n15403), .ZN(n15402) );
  NAND2_X1 U15464 ( .A1(n15241), .A2(n15240), .ZN(n15403) );
  NOR2_X1 U15465 ( .A1(n7645), .A2(n8063), .ZN(n15242) );
  OR2_X1 U15466 ( .A1(n15240), .A2(n15241), .ZN(n15401) );
  AND2_X1 U15467 ( .A1(n15404), .A2(n15405), .ZN(n15241) );
  NAND2_X1 U15468 ( .A1(n15406), .A2(b_2_), .ZN(n15405) );
  NOR2_X1 U15469 ( .A1(n15407), .A2(n7624), .ZN(n15406) );
  NOR2_X1 U15470 ( .A1(n15176), .A2(n15178), .ZN(n15407) );
  NAND2_X1 U15471 ( .A1(n15176), .A2(n15178), .ZN(n15404) );
  NAND2_X1 U15472 ( .A1(n15408), .A2(n15409), .ZN(n15178) );
  NAND2_X1 U15473 ( .A1(n15238), .A2(n15410), .ZN(n15409) );
  OR2_X1 U15474 ( .A1(n15237), .A2(n15235), .ZN(n15410) );
  NOR2_X1 U15475 ( .A1(n8063), .A2(n7613), .ZN(n15238) );
  NAND2_X1 U15476 ( .A1(n15235), .A2(n15237), .ZN(n15408) );
  NAND2_X1 U15477 ( .A1(n15411), .A2(n15412), .ZN(n15237) );
  NAND2_X1 U15478 ( .A1(n15191), .A2(n15413), .ZN(n15412) );
  OR2_X1 U15479 ( .A1(n15190), .A2(n15188), .ZN(n15413) );
  NOR2_X1 U15480 ( .A1(n8063), .A2(n7593), .ZN(n15191) );
  NAND2_X1 U15481 ( .A1(n15188), .A2(n15190), .ZN(n15411) );
  NAND2_X1 U15482 ( .A1(n15233), .A2(n15414), .ZN(n15190) );
  NAND2_X1 U15483 ( .A1(n15232), .A2(n15234), .ZN(n15414) );
  NAND2_X1 U15484 ( .A1(n15415), .A2(n15416), .ZN(n15234) );
  NAND2_X1 U15485 ( .A1(b_2_), .A2(a_26_), .ZN(n15416) );
  INV_X1 U15486 ( .A(n15417), .ZN(n15415) );
  XOR2_X1 U15487 ( .A(n15418), .B(n15419), .Z(n15232) );
  NOR2_X1 U15488 ( .A1(n7547), .A2(n15294), .ZN(n15419) );
  XOR2_X1 U15489 ( .A(n15420), .B(n15421), .Z(n15418) );
  NAND2_X1 U15490 ( .A1(a_26_), .A2(n15417), .ZN(n15233) );
  NAND2_X1 U15491 ( .A1(n15229), .A2(n15422), .ZN(n15417) );
  NAND2_X1 U15492 ( .A1(n15228), .A2(n15230), .ZN(n15422) );
  NAND2_X1 U15493 ( .A1(n15423), .A2(n15424), .ZN(n15230) );
  NAND2_X1 U15494 ( .A1(b_2_), .A2(a_27_), .ZN(n15424) );
  INV_X1 U15495 ( .A(n15425), .ZN(n15423) );
  XOR2_X1 U15496 ( .A(n15426), .B(n15427), .Z(n15228) );
  XNOR2_X1 U15497 ( .A(n15428), .B(n15429), .ZN(n15427) );
  NAND2_X1 U15498 ( .A1(b_0_), .A2(a_29_), .ZN(n15426) );
  NAND2_X1 U15499 ( .A1(a_27_), .A2(n15425), .ZN(n15229) );
  NAND2_X1 U15500 ( .A1(n15225), .A2(n15430), .ZN(n15425) );
  NAND2_X1 U15501 ( .A1(n15224), .A2(n15226), .ZN(n15430) );
  NAND2_X1 U15502 ( .A1(n15431), .A2(n15432), .ZN(n15226) );
  NAND2_X1 U15503 ( .A1(b_2_), .A2(a_28_), .ZN(n15432) );
  INV_X1 U15504 ( .A(n15433), .ZN(n15431) );
  XNOR2_X1 U15505 ( .A(n15434), .B(n15435), .ZN(n15224) );
  XNOR2_X1 U15506 ( .A(n15436), .B(n15437), .ZN(n15435) );
  NAND2_X1 U15507 ( .A1(b_0_), .A2(a_30_), .ZN(n15434) );
  NAND2_X1 U15508 ( .A1(a_28_), .A2(n15433), .ZN(n15225) );
  NAND2_X1 U15509 ( .A1(n15438), .A2(n15439), .ZN(n15433) );
  NAND2_X1 U15510 ( .A1(n15440), .A2(b_2_), .ZN(n15439) );
  NOR2_X1 U15511 ( .A1(n15441), .A2(n7529), .ZN(n15440) );
  NOR2_X1 U15512 ( .A1(n15221), .A2(n15222), .ZN(n15441) );
  NAND2_X1 U15513 ( .A1(n15221), .A2(n15222), .ZN(n15438) );
  NAND2_X1 U15514 ( .A1(n15442), .A2(n15443), .ZN(n15222) );
  NAND2_X1 U15515 ( .A1(n15444), .A2(b_0_), .ZN(n15443) );
  NOR2_X1 U15516 ( .A1(n15445), .A2(n8048), .ZN(n15444) );
  NOR2_X1 U15517 ( .A1(n8676), .A2(n15217), .ZN(n15445) );
  NAND2_X1 U15518 ( .A1(a_31_), .A2(n7515), .ZN(n7506) );
  NAND2_X1 U15519 ( .A1(n15446), .A2(b_1_), .ZN(n15442) );
  NOR2_X1 U15520 ( .A1(n15447), .A2(n7515), .ZN(n15446) );
  NOR2_X1 U15521 ( .A1(n8679), .A2(n15294), .ZN(n15447) );
  NAND2_X1 U15522 ( .A1(a_30_), .A2(n8048), .ZN(n7510) );
  AND2_X1 U15523 ( .A1(n15448), .A2(b_1_), .ZN(n15221) );
  NOR2_X1 U15524 ( .A1(n8451), .A2(n8063), .ZN(n15448) );
  INV_X1 U15525 ( .A(b_2_), .ZN(n8063) );
  XOR2_X1 U15526 ( .A(n15449), .B(n15450), .Z(n15188) );
  NOR2_X1 U15527 ( .A1(n15451), .A2(n15452), .ZN(n15450) );
  INV_X1 U15528 ( .A(n15453), .ZN(n15452) );
  NOR2_X1 U15529 ( .A1(n15454), .A2(n15455), .ZN(n15451) );
  XOR2_X1 U15530 ( .A(n15456), .B(n15457), .Z(n15235) );
  NOR2_X1 U15531 ( .A1(n8052), .A2(n15294), .ZN(n15457) );
  XOR2_X1 U15532 ( .A(n15458), .B(n15459), .Z(n15456) );
  XOR2_X1 U15533 ( .A(n15460), .B(n15461), .Z(n15176) );
  NOR2_X1 U15534 ( .A1(n15462), .A2(n15463), .ZN(n15461) );
  INV_X1 U15535 ( .A(n15464), .ZN(n15463) );
  NOR2_X1 U15536 ( .A1(n15465), .A2(n15466), .ZN(n15462) );
  XNOR2_X1 U15537 ( .A(n15467), .B(n15468), .ZN(n15240) );
  NOR2_X1 U15538 ( .A1(n7613), .A2(n15294), .ZN(n15468) );
  XOR2_X1 U15539 ( .A(n15469), .B(n15470), .Z(n15467) );
  XOR2_X1 U15540 ( .A(n15471), .B(n15472), .Z(n15165) );
  NOR2_X1 U15541 ( .A1(n15473), .A2(n15474), .ZN(n15472) );
  INV_X1 U15542 ( .A(n15475), .ZN(n15474) );
  NOR2_X1 U15543 ( .A1(n15476), .A2(n15477), .ZN(n15473) );
  XNOR2_X1 U15544 ( .A(n15478), .B(n15479), .ZN(n15244) );
  NOR2_X1 U15545 ( .A1(n7645), .A2(n15294), .ZN(n15479) );
  XOR2_X1 U15546 ( .A(n15480), .B(n15481), .Z(n15478) );
  XOR2_X1 U15547 ( .A(n15482), .B(n15483), .Z(n15153) );
  NOR2_X1 U15548 ( .A1(n15484), .A2(n15485), .ZN(n15483) );
  INV_X1 U15549 ( .A(n15486), .ZN(n15485) );
  NOR2_X1 U15550 ( .A1(n15487), .A2(n15488), .ZN(n15484) );
  XNOR2_X1 U15551 ( .A(n15489), .B(n15490), .ZN(n15248) );
  NOR2_X1 U15552 ( .A1(n7676), .A2(n15294), .ZN(n15490) );
  XOR2_X1 U15553 ( .A(n15491), .B(n15492), .Z(n15489) );
  XOR2_X1 U15554 ( .A(n15493), .B(n15494), .Z(n15141) );
  NOR2_X1 U15555 ( .A1(n15495), .A2(n15496), .ZN(n15494) );
  INV_X1 U15556 ( .A(n15497), .ZN(n15496) );
  NOR2_X1 U15557 ( .A1(n15498), .A2(n15499), .ZN(n15495) );
  XNOR2_X1 U15558 ( .A(n15500), .B(n15501), .ZN(n15129) );
  NOR2_X1 U15559 ( .A1(n15502), .A2(n15503), .ZN(n15501) );
  INV_X1 U15560 ( .A(n15504), .ZN(n15503) );
  NOR2_X1 U15561 ( .A1(n15505), .A2(n15506), .ZN(n15502) );
  XNOR2_X1 U15562 ( .A(n15507), .B(n15508), .ZN(n15117) );
  NOR2_X1 U15563 ( .A1(n15509), .A2(n15510), .ZN(n15508) );
  INV_X1 U15564 ( .A(n15511), .ZN(n15510) );
  NOR2_X1 U15565 ( .A1(n15512), .A2(n15513), .ZN(n15509) );
  XNOR2_X1 U15566 ( .A(n15514), .B(n15515), .ZN(n15105) );
  NOR2_X1 U15567 ( .A1(n15516), .A2(n15517), .ZN(n15515) );
  INV_X1 U15568 ( .A(n15518), .ZN(n15517) );
  NOR2_X1 U15569 ( .A1(n15519), .A2(n15520), .ZN(n15516) );
  XNOR2_X1 U15570 ( .A(n15521), .B(n15522), .ZN(n15093) );
  NOR2_X1 U15571 ( .A1(n15523), .A2(n15524), .ZN(n15522) );
  INV_X1 U15572 ( .A(n15525), .ZN(n15524) );
  NOR2_X1 U15573 ( .A1(n15526), .A2(n15527), .ZN(n15523) );
  XNOR2_X1 U15574 ( .A(n15528), .B(n15529), .ZN(n15081) );
  NOR2_X1 U15575 ( .A1(n15530), .A2(n15531), .ZN(n15529) );
  INV_X1 U15576 ( .A(n15532), .ZN(n15531) );
  NOR2_X1 U15577 ( .A1(n15533), .A2(n15534), .ZN(n15530) );
  XNOR2_X1 U15578 ( .A(n15535), .B(n15536), .ZN(n15069) );
  NOR2_X1 U15579 ( .A1(n15537), .A2(n15538), .ZN(n15536) );
  INV_X1 U15580 ( .A(n15539), .ZN(n15538) );
  NOR2_X1 U15581 ( .A1(n15540), .A2(n15541), .ZN(n15537) );
  XNOR2_X1 U15582 ( .A(n15542), .B(n15543), .ZN(n15054) );
  NOR2_X1 U15583 ( .A1(n15544), .A2(n15545), .ZN(n15543) );
  INV_X1 U15584 ( .A(n15546), .ZN(n15545) );
  NOR2_X1 U15585 ( .A1(n15547), .A2(n15548), .ZN(n15544) );
  NAND2_X1 U15586 ( .A1(a_2_), .A2(b_2_), .ZN(n7959) );
  XOR2_X1 U15587 ( .A(n15549), .B(n15550), .Z(n15279) );
  NOR2_X1 U15588 ( .A1(n15551), .A2(n15552), .ZN(n15550) );
  INV_X1 U15589 ( .A(n15553), .ZN(n15552) );
  NOR2_X1 U15590 ( .A1(n15554), .A2(n15555), .ZN(n15551) );
  XOR2_X1 U15591 ( .A(n15556), .B(n15557), .Z(n8195) );
  NOR2_X1 U15592 ( .A1(n15558), .A2(n15559), .ZN(n15557) );
  INV_X1 U15593 ( .A(n15560), .ZN(n15559) );
  NOR2_X1 U15594 ( .A1(n15561), .A2(n15562), .ZN(n15558) );
  XOR2_X1 U15595 ( .A(n7989), .B(n8196), .Z(n15286) );
  NOR2_X1 U15596 ( .A1(n15294), .A2(n8307), .ZN(n7989) );
  NOR2_X1 U15597 ( .A1(n8196), .A2(n8307), .ZN(n8189) );
  AND2_X1 U15598 ( .A1(n15560), .A2(n15563), .ZN(n8196) );
  NAND2_X1 U15599 ( .A1(n15564), .A2(n15556), .ZN(n15563) );
  NAND2_X1 U15600 ( .A1(n15565), .A2(n15566), .ZN(n15556) );
  NAND2_X1 U15601 ( .A1(n15567), .A2(a_2_), .ZN(n15566) );
  NOR2_X1 U15602 ( .A1(n15568), .A2(n15294), .ZN(n15567) );
  NOR2_X1 U15603 ( .A1(n7979), .A2(n15295), .ZN(n15568) );
  NAND2_X1 U15604 ( .A1(n7979), .A2(n15295), .ZN(n15565) );
  NAND2_X1 U15605 ( .A1(n15553), .A2(n15569), .ZN(n15295) );
  NAND2_X1 U15606 ( .A1(n15570), .A2(n15549), .ZN(n15569) );
  NAND2_X1 U15607 ( .A1(n15571), .A2(n15572), .ZN(n15549) );
  NAND2_X1 U15608 ( .A1(n15573), .A2(a_3_), .ZN(n15572) );
  NOR2_X1 U15609 ( .A1(n15574), .A2(n15217), .ZN(n15573) );
  NOR2_X1 U15610 ( .A1(n15305), .A2(n15304), .ZN(n15574) );
  NAND2_X1 U15611 ( .A1(n15305), .A2(n15304), .ZN(n15571) );
  NAND2_X1 U15612 ( .A1(n15546), .A2(n15575), .ZN(n15304) );
  NAND2_X1 U15613 ( .A1(n15576), .A2(n15542), .ZN(n15575) );
  NAND2_X1 U15614 ( .A1(n15577), .A2(n15578), .ZN(n15542) );
  NAND2_X1 U15615 ( .A1(n15579), .A2(a_5_), .ZN(n15578) );
  NOR2_X1 U15616 ( .A1(n15580), .A2(n15217), .ZN(n15579) );
  NOR2_X1 U15617 ( .A1(n15316), .A2(n15315), .ZN(n15580) );
  NAND2_X1 U15618 ( .A1(n15316), .A2(n15315), .ZN(n15577) );
  NAND2_X1 U15619 ( .A1(n15539), .A2(n15581), .ZN(n15315) );
  NAND2_X1 U15620 ( .A1(n15582), .A2(n15535), .ZN(n15581) );
  NAND2_X1 U15621 ( .A1(n15583), .A2(n15584), .ZN(n15535) );
  NAND2_X1 U15622 ( .A1(n15585), .A2(a_7_), .ZN(n15584) );
  NOR2_X1 U15623 ( .A1(n15586), .A2(n15217), .ZN(n15585) );
  NOR2_X1 U15624 ( .A1(n15327), .A2(n15326), .ZN(n15586) );
  NAND2_X1 U15625 ( .A1(n15327), .A2(n15326), .ZN(n15583) );
  NAND2_X1 U15626 ( .A1(n15532), .A2(n15587), .ZN(n15326) );
  NAND2_X1 U15627 ( .A1(n15588), .A2(n15528), .ZN(n15587) );
  NAND2_X1 U15628 ( .A1(n15589), .A2(n15590), .ZN(n15528) );
  NAND2_X1 U15629 ( .A1(n15591), .A2(a_9_), .ZN(n15590) );
  NOR2_X1 U15630 ( .A1(n15592), .A2(n15217), .ZN(n15591) );
  NOR2_X1 U15631 ( .A1(n15338), .A2(n15337), .ZN(n15592) );
  NAND2_X1 U15632 ( .A1(n15338), .A2(n15337), .ZN(n15589) );
  NAND2_X1 U15633 ( .A1(n15525), .A2(n15593), .ZN(n15337) );
  NAND2_X1 U15634 ( .A1(n15594), .A2(n15521), .ZN(n15593) );
  NAND2_X1 U15635 ( .A1(n15595), .A2(n15596), .ZN(n15521) );
  NAND2_X1 U15636 ( .A1(n15597), .A2(b_1_), .ZN(n15596) );
  NOR2_X1 U15637 ( .A1(n15598), .A2(n7817), .ZN(n15597) );
  NOR2_X1 U15638 ( .A1(n15349), .A2(n15348), .ZN(n15598) );
  NAND2_X1 U15639 ( .A1(n15349), .A2(n15348), .ZN(n15595) );
  NAND2_X1 U15640 ( .A1(n15518), .A2(n15599), .ZN(n15348) );
  NAND2_X1 U15641 ( .A1(n15600), .A2(n15514), .ZN(n15599) );
  NAND2_X1 U15642 ( .A1(n15601), .A2(n15602), .ZN(n15514) );
  NAND2_X1 U15643 ( .A1(n15603), .A2(a_13_), .ZN(n15602) );
  NOR2_X1 U15644 ( .A1(n15604), .A2(n15217), .ZN(n15603) );
  NOR2_X1 U15645 ( .A1(n15360), .A2(n15359), .ZN(n15604) );
  NAND2_X1 U15646 ( .A1(n15360), .A2(n15359), .ZN(n15601) );
  NAND2_X1 U15647 ( .A1(n15511), .A2(n15605), .ZN(n15359) );
  NAND2_X1 U15648 ( .A1(n15606), .A2(n15507), .ZN(n15605) );
  NAND2_X1 U15649 ( .A1(n15607), .A2(n15608), .ZN(n15507) );
  NAND2_X1 U15650 ( .A1(n15609), .A2(a_15_), .ZN(n15608) );
  NOR2_X1 U15651 ( .A1(n15610), .A2(n15217), .ZN(n15609) );
  NOR2_X1 U15652 ( .A1(n15371), .A2(n15370), .ZN(n15610) );
  NAND2_X1 U15653 ( .A1(n15371), .A2(n15370), .ZN(n15607) );
  NAND2_X1 U15654 ( .A1(n15504), .A2(n15611), .ZN(n15370) );
  NAND2_X1 U15655 ( .A1(n15612), .A2(n15500), .ZN(n15611) );
  NAND2_X1 U15656 ( .A1(n15613), .A2(n15614), .ZN(n15500) );
  NAND2_X1 U15657 ( .A1(n15615), .A2(a_17_), .ZN(n15614) );
  NOR2_X1 U15658 ( .A1(n15616), .A2(n15217), .ZN(n15615) );
  NOR2_X1 U15659 ( .A1(n15382), .A2(n15381), .ZN(n15616) );
  NAND2_X1 U15660 ( .A1(n15382), .A2(n15381), .ZN(n15613) );
  NAND2_X1 U15661 ( .A1(n15497), .A2(n15617), .ZN(n15381) );
  NAND2_X1 U15662 ( .A1(n15618), .A2(n15493), .ZN(n15617) );
  NAND2_X1 U15663 ( .A1(n15619), .A2(n15620), .ZN(n15493) );
  NAND2_X1 U15664 ( .A1(n15621), .A2(b_0_), .ZN(n15620) );
  NOR2_X1 U15665 ( .A1(n15622), .A2(n7676), .ZN(n15621) );
  NOR2_X1 U15666 ( .A1(n15492), .A2(n15491), .ZN(n15622) );
  NAND2_X1 U15667 ( .A1(n15492), .A2(n15491), .ZN(n15619) );
  NAND2_X1 U15668 ( .A1(n15486), .A2(n15623), .ZN(n15491) );
  NAND2_X1 U15669 ( .A1(n15624), .A2(n15482), .ZN(n15623) );
  NAND2_X1 U15670 ( .A1(n15625), .A2(n15626), .ZN(n15482) );
  NAND2_X1 U15671 ( .A1(n15627), .A2(b_0_), .ZN(n15626) );
  NOR2_X1 U15672 ( .A1(n15628), .A2(n7645), .ZN(n15627) );
  NOR2_X1 U15673 ( .A1(n15481), .A2(n15480), .ZN(n15628) );
  NAND2_X1 U15674 ( .A1(n15481), .A2(n15480), .ZN(n15625) );
  NAND2_X1 U15675 ( .A1(n15475), .A2(n15629), .ZN(n15480) );
  NAND2_X1 U15676 ( .A1(n15630), .A2(n15471), .ZN(n15629) );
  NAND2_X1 U15677 ( .A1(n15631), .A2(n15632), .ZN(n15471) );
  NAND2_X1 U15678 ( .A1(n15633), .A2(b_0_), .ZN(n15632) );
  NOR2_X1 U15679 ( .A1(n15634), .A2(n7613), .ZN(n15633) );
  NOR2_X1 U15680 ( .A1(n15470), .A2(n15469), .ZN(n15634) );
  NAND2_X1 U15681 ( .A1(n15470), .A2(n15469), .ZN(n15631) );
  NAND2_X1 U15682 ( .A1(n15464), .A2(n15635), .ZN(n15469) );
  NAND2_X1 U15683 ( .A1(n15636), .A2(n15460), .ZN(n15635) );
  NAND2_X1 U15684 ( .A1(n15637), .A2(n15638), .ZN(n15460) );
  NAND2_X1 U15685 ( .A1(n15639), .A2(b_0_), .ZN(n15638) );
  NOR2_X1 U15686 ( .A1(n15640), .A2(n8052), .ZN(n15639) );
  NOR2_X1 U15687 ( .A1(n15459), .A2(n15458), .ZN(n15640) );
  NAND2_X1 U15688 ( .A1(n15459), .A2(n15458), .ZN(n15637) );
  NAND2_X1 U15689 ( .A1(n15453), .A2(n15641), .ZN(n15458) );
  NAND2_X1 U15690 ( .A1(n15642), .A2(n15449), .ZN(n15641) );
  NAND2_X1 U15691 ( .A1(n15643), .A2(n15644), .ZN(n15449) );
  NAND2_X1 U15692 ( .A1(n15645), .A2(b_0_), .ZN(n15644) );
  NOR2_X1 U15693 ( .A1(n15646), .A2(n7547), .ZN(n15645) );
  NOR2_X1 U15694 ( .A1(n15421), .A2(n15420), .ZN(n15646) );
  NAND2_X1 U15695 ( .A1(n15421), .A2(n15420), .ZN(n15643) );
  NAND2_X1 U15696 ( .A1(n15647), .A2(n15648), .ZN(n15420) );
  NAND2_X1 U15697 ( .A1(n15649), .A2(b_0_), .ZN(n15648) );
  NOR2_X1 U15698 ( .A1(n15650), .A2(n7529), .ZN(n15649) );
  NOR2_X1 U15699 ( .A1(n15428), .A2(n15429), .ZN(n15650) );
  NAND2_X1 U15700 ( .A1(n15428), .A2(n15429), .ZN(n15647) );
  NAND2_X1 U15701 ( .A1(n15437), .A2(n15651), .ZN(n15429) );
  NAND2_X1 U15702 ( .A1(n15652), .A2(n15436), .ZN(n15651) );
  NOR2_X1 U15703 ( .A1(n15217), .A2(n7529), .ZN(n15436) );
  NOR2_X1 U15704 ( .A1(n7515), .A2(n15294), .ZN(n15652) );
  NAND2_X1 U15705 ( .A1(n15653), .A2(b_0_), .ZN(n15437) );
  NOR2_X1 U15706 ( .A1(n8451), .A2(n15217), .ZN(n15653) );
  NOR2_X1 U15707 ( .A1(n15217), .A2(n7547), .ZN(n15428) );
  INV_X1 U15708 ( .A(a_28_), .ZN(n7547) );
  NOR2_X1 U15709 ( .A1(n15217), .A2(n7563), .ZN(n15421) );
  OR2_X1 U15710 ( .A1(n15454), .A2(a_27_), .ZN(n15642) );
  NAND2_X1 U15711 ( .A1(n15455), .A2(n15454), .ZN(n15453) );
  NOR2_X1 U15712 ( .A1(n15217), .A2(n8052), .ZN(n15454) );
  INV_X1 U15713 ( .A(a_26_), .ZN(n8052) );
  NOR2_X1 U15714 ( .A1(n7563), .A2(n15294), .ZN(n15455) );
  NOR2_X1 U15715 ( .A1(n15217), .A2(n7593), .ZN(n15459) );
  OR2_X1 U15716 ( .A1(n15465), .A2(a_25_), .ZN(n15636) );
  NAND2_X1 U15717 ( .A1(n15466), .A2(n15465), .ZN(n15464) );
  NOR2_X1 U15718 ( .A1(n15217), .A2(n7613), .ZN(n15465) );
  INV_X1 U15719 ( .A(a_24_), .ZN(n7613) );
  NOR2_X1 U15720 ( .A1(n7593), .A2(n15294), .ZN(n15466) );
  NOR2_X1 U15721 ( .A1(n15217), .A2(n7624), .ZN(n15470) );
  OR2_X1 U15722 ( .A1(n15476), .A2(a_23_), .ZN(n15630) );
  NAND2_X1 U15723 ( .A1(n15477), .A2(n15476), .ZN(n15475) );
  NOR2_X1 U15724 ( .A1(n15217), .A2(n7645), .ZN(n15476) );
  NOR2_X1 U15725 ( .A1(n7624), .A2(n15294), .ZN(n15477) );
  NOR2_X1 U15726 ( .A1(n15217), .A2(n7656), .ZN(n15481) );
  OR2_X1 U15727 ( .A1(n15487), .A2(a_21_), .ZN(n15624) );
  NAND2_X1 U15728 ( .A1(n15488), .A2(n15487), .ZN(n15486) );
  NOR2_X1 U15729 ( .A1(n15217), .A2(n7676), .ZN(n15487) );
  NOR2_X1 U15730 ( .A1(n7656), .A2(n15294), .ZN(n15488) );
  NOR2_X1 U15731 ( .A1(n7687), .A2(n15217), .ZN(n15492) );
  OR2_X1 U15732 ( .A1(n15498), .A2(a_19_), .ZN(n15618) );
  NAND2_X1 U15733 ( .A1(n15499), .A2(n15498), .ZN(n15497) );
  NOR2_X1 U15734 ( .A1(n7707), .A2(n15217), .ZN(n15498) );
  NOR2_X1 U15735 ( .A1(n15294), .A2(n7687), .ZN(n15499) );
  NOR2_X1 U15736 ( .A1(n7707), .A2(n15294), .ZN(n15382) );
  OR2_X1 U15737 ( .A1(n15505), .A2(a_16_), .ZN(n15612) );
  NAND2_X1 U15738 ( .A1(n15506), .A2(n15505), .ZN(n15504) );
  NOR2_X1 U15739 ( .A1(n7723), .A2(n15294), .ZN(n15505) );
  NOR2_X1 U15740 ( .A1(n15217), .A2(n7743), .ZN(n15506) );
  NOR2_X1 U15741 ( .A1(n7743), .A2(n15294), .ZN(n15371) );
  OR2_X1 U15742 ( .A1(n15512), .A2(a_14_), .ZN(n15606) );
  NAND2_X1 U15743 ( .A1(n15513), .A2(n15512), .ZN(n15511) );
  NOR2_X1 U15744 ( .A1(n7754), .A2(n15294), .ZN(n15512) );
  NOR2_X1 U15745 ( .A1(n15217), .A2(n7775), .ZN(n15513) );
  NOR2_X1 U15746 ( .A1(n7775), .A2(n15294), .ZN(n15360) );
  OR2_X1 U15747 ( .A1(n15519), .A2(a_12_), .ZN(n15600) );
  NAND2_X1 U15748 ( .A1(n15520), .A2(n15519), .ZN(n15518) );
  NOR2_X1 U15749 ( .A1(n7786), .A2(n15294), .ZN(n15519) );
  NOR2_X1 U15750 ( .A1(n15217), .A2(n7806), .ZN(n15520) );
  NOR2_X1 U15751 ( .A1(n7806), .A2(n15294), .ZN(n15349) );
  OR2_X1 U15752 ( .A1(n15526), .A2(a_10_), .ZN(n15594) );
  NAND2_X1 U15753 ( .A1(n15527), .A2(n15526), .ZN(n15525) );
  NOR2_X1 U15754 ( .A1(n15294), .A2(n7817), .ZN(n15526) );
  NOR2_X1 U15755 ( .A1(n15217), .A2(n7837), .ZN(n15527) );
  NOR2_X1 U15756 ( .A1(n7837), .A2(n15294), .ZN(n15338) );
  OR2_X1 U15757 ( .A1(n15533), .A2(a_8_), .ZN(n15588) );
  NAND2_X1 U15758 ( .A1(n15534), .A2(n15533), .ZN(n15532) );
  NOR2_X1 U15759 ( .A1(n7848), .A2(n15294), .ZN(n15533) );
  NOR2_X1 U15760 ( .A1(n15217), .A2(n8059), .ZN(n15534) );
  NOR2_X1 U15761 ( .A1(n8059), .A2(n15294), .ZN(n15327) );
  OR2_X1 U15762 ( .A1(n15540), .A2(a_6_), .ZN(n15582) );
  NAND2_X1 U15763 ( .A1(n15541), .A2(n15540), .ZN(n15539) );
  NOR2_X1 U15764 ( .A1(n7884), .A2(n15294), .ZN(n15540) );
  NOR2_X1 U15765 ( .A1(n15217), .A2(n8061), .ZN(n15541) );
  NOR2_X1 U15766 ( .A1(n8061), .A2(n15294), .ZN(n15316) );
  OR2_X1 U15767 ( .A1(n15547), .A2(a_4_), .ZN(n15576) );
  NAND2_X1 U15768 ( .A1(n15548), .A2(n15547), .ZN(n15546) );
  NOR2_X1 U15769 ( .A1(n7914), .A2(n15294), .ZN(n15547) );
  NOR2_X1 U15770 ( .A1(n15217), .A2(n7934), .ZN(n15548) );
  NOR2_X1 U15771 ( .A1(n7934), .A2(n15294), .ZN(n15305) );
  OR2_X1 U15772 ( .A1(n15554), .A2(a_2_), .ZN(n15570) );
  NAND2_X1 U15773 ( .A1(n15555), .A2(n15554), .ZN(n15553) );
  NOR2_X1 U15774 ( .A1(n7945), .A2(n15294), .ZN(n15554) );
  NOR2_X1 U15775 ( .A1(n15217), .A2(n7965), .ZN(n15555) );
  INV_X1 U15776 ( .A(a_2_), .ZN(n7965) );
  NOR2_X1 U15777 ( .A1(n7973), .A2(n15217), .ZN(n7979) );
  OR2_X1 U15778 ( .A1(n15561), .A2(a_0_), .ZN(n15564) );
  NAND2_X1 U15779 ( .A1(n15562), .A2(n15561), .ZN(n15560) );
  NOR2_X1 U15780 ( .A1(n7973), .A2(n15294), .ZN(n15561) );
  NOR2_X1 U15781 ( .A1(n8307), .A2(n15217), .ZN(n15562) );
endmodule

