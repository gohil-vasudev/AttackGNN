module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137;
output N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n236_, new_n976_, new_n238_, new_n479_, new_n1009_, new_n1105_, new_n955_, new_n608_, new_n847_, new_n250_, new_n501_, new_n288_, new_n1157_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n885_, new_n439_, new_n827_, new_n283_, new_n223_, new_n390_, new_n743_, new_n366_, new_n779_, new_n241_, new_n1025_, new_n566_, new_n186_, new_n339_, new_n365_, new_n641_, new_n197_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n456_, new_n691_, new_n1024_, new_n1125_, new_n170_, new_n246_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n266_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n173_, new_n220_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n214_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n188_, new_n695_, new_n240_, new_n660_, new_n413_, new_n1060_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n211_, new_n552_, new_n678_, new_n342_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n1132_, new_n500_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n317_, new_n344_, new_n287_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n234_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n292_, new_n1167_, new_n215_, new_n626_, new_n152_, new_n959_, new_n990_, new_n774_, new_n157_, new_n716_, new_n153_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n257_, new_n1162_, new_n481_, new_n212_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n272_, new_n282_, new_n1059_, new_n201_, new_n634_, new_n192_, new_n414_, new_n1101_, new_n635_, new_n315_, new_n685_, new_n326_, new_n554_, new_n648_, new_n1050_, new_n164_, new_n230_, new_n983_, new_n281_, new_n430_, new_n822_, new_n482_, new_n844_, new_n1151_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n248_, new_n350_, new_n655_, new_n759_, new_n630_, new_n1054_, new_n167_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n297_, new_n361_, new_n565_, new_n764_, new_n906_, new_n150_, new_n683_, new_n183_, new_n511_, new_n463_, new_n303_, new_n510_, new_n966_, new_n351_, new_n1184_, new_n517_, new_n325_, new_n609_, new_n180_, new_n1031_, new_n961_, new_n530_, new_n890_, new_n318_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n321_, new_n715_, new_n811_, new_n443_, new_n324_, new_n1086_, new_n956_, new_n158_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n262_, new_n970_, new_n995_, new_n1035_, new_n271_, new_n674_, new_n274_, new_n991_, new_n1044_, new_n218_, new_n497_, new_n816_, new_n1170_, new_n845_, new_n768_, new_n773_, new_n305_, new_n420_, new_n568_, new_n876_, new_n899_, new_n1051_, new_n1053_, new_n423_, new_n205_, new_n492_, new_n496_, new_n498_, new_n141_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n1182_, new_n206_, new_n887_, new_n254_, new_n429_, new_n355_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n256_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n1028_, new_n1168_, new_n508_, new_n714_, new_n194_, new_n483_, new_n1004_, new_n1152_, new_n394_, new_n299_, new_n1007_, new_n142_, new_n935_, new_n139_, new_n882_, new_n657_, new_n929_, new_n652_, new_n314_, new_n582_, new_n986_, new_n1020_, new_n363_, new_n1159_, new_n1113_, new_n165_, new_n441_, new_n785_, new_n477_, new_n664_, new_n216_, new_n600_, new_n280_, new_n917_, new_n1041_, new_n426_, new_n1036_, new_n235_, new_n1133_, new_n398_, new_n301_, new_n1177_, new_n169_, new_n646_, new_n395_, new_n538_, new_n383_, new_n343_, new_n210_, new_n458_, new_n541_, new_n447_, new_n854_, new_n1026_, new_n207_, new_n267_, new_n1106_, new_n473_, new_n140_, new_n1147_, new_n790_, new_n1081_, new_n187_, new_n311_, new_n587_, new_n465_, new_n739_, new_n783_, new_n263_, new_n334_, new_n331_, new_n835_, new_n341_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n244_, new_n172_, new_n488_, new_n524_, new_n277_, new_n705_, new_n848_, new_n874_, new_n943_, new_n402_, new_n663_, new_n579_, new_n286_, new_n335_, new_n347_, new_n659_, new_n700_, new_n921_, new_n346_, new_n396_, new_n198_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n208_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n179_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n233_, new_n469_, new_n391_, new_n178_, new_n437_, new_n1085_, new_n1154_, new_n295_, new_n359_, new_n794_, new_n628_, new_n166_, new_n162_, new_n409_, new_n745_, new_n1090_, new_n457_, new_n161_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n333_, new_n1128_, new_n1002_, new_n290_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n276_, new_n688_, new_n155_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n1096_, new_n454_, new_n202_, new_n1034_, new_n296_, new_n661_, new_n308_, new_n1000_, new_n633_, new_n797_, new_n232_, new_n784_, new_n258_, new_n724_, new_n1070_, new_n176_, new_n156_, new_n306_, new_n494_, new_n860_, new_n291_, new_n261_, new_n672_, new_n309_, new_n616_, new_n529_, new_n323_, new_n884_, new_n914_, new_n259_, new_n362_, new_n938_, new_n1160_, new_n809_, new_n1142_, new_n654_, new_n1166_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n227_, new_n1104_, new_n690_, new_n416_, new_n222_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n328_, new_n460_, new_n1136_, new_n693_, new_n1175_, new_n505_, new_n619_, new_n471_, new_n967_, new_n268_, new_n374_, new_n577_, new_n1135_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n138_, new_n749_, new_n861_, new_n1091_, new_n310_, new_n144_, new_n1095_, new_n275_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n177_, new_n1118_, new_n493_, new_n547_, new_n907_, new_n264_, new_n665_, new_n800_, new_n379_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n273_, new_n1178_, new_n224_, new_n586_, new_n963_, new_n270_, new_n570_, new_n598_, new_n993_, new_n1063_, new_n824_, new_n143_, new_n520_, new_n145_, new_n253_, new_n717_, new_n403_, new_n475_, new_n868_, new_n237_, new_n825_, new_n858_, new_n149_, new_n557_, new_n260_, new_n251_, new_n189_, new_n300_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n1144_, new_n1137_, new_n182_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n151_, new_n513_, new_n592_, new_n726_, new_n1123_, new_n558_, new_n219_, new_n231_, new_n313_, new_n382_, new_n239_, new_n583_, new_n617_, new_n718_, new_n1080_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n199_, new_n146_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n546_, new_n612_, new_n919_, new_n1015_, new_n302_, new_n191_, new_n755_, new_n225_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n221_, new_n243_, new_n450_, new_n345_, new_n1179_, new_n298_, new_n184_, new_n499_, new_n154_, new_n255_, new_n533_, new_n1130_, new_n1148_, new_n795_, new_n1146_, new_n459_, new_n569_, new_n555_, new_n174_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n340_, new_n147_, new_n285_, new_n502_, new_n692_, new_n613_, new_n209_, new_n337_, new_n446_, new_n623_, new_n203_, new_n316_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n332_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n163_, new_n997_, new_n519_, new_n563_, new_n148_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n1076_, new_n252_, new_n585_, new_n751_, new_n160_, new_n312_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n242_, new_n503_, new_n527_, new_n772_, new_n852_, new_n307_, new_n190_, new_n597_, new_n978_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n213_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n265_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n278_, new_n304_, new_n523_, new_n638_, new_n857_, new_n909_, new_n1052_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n217_, new_n269_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n327_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n196_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n319_, new_n1008_, new_n640_, new_n684_, new_n338_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n336_, new_n377_, new_n247_, new_n539_, new_n905_, new_n803_, new_n330_, new_n727_, new_n375_, new_n962_, new_n294_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n195_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1153_, new_n357_, new_n320_, new_n780_, new_n984_, new_n1183_, new_n245_, new_n643_, new_n474_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n193_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n159_, new_n843_, new_n322_, new_n228_, new_n545_, new_n611_, new_n703_, new_n289_, new_n698_, new_n1165_, new_n425_, new_n175_, new_n226_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n185_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n171_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n200_, new_n947_, new_n994_, new_n982_, new_n422_, new_n581_, new_n329_, new_n249_, new_n284_, new_n293_, new_n686_, new_n934_, new_n551_, new_n168_, new_n279_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n229_, new_n536_, new_n889_, new_n464_, new_n204_, new_n1089_, new_n181_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g0000 ( new_n138_, keyIn_0_38 );
not g0001 ( new_n139_, keyIn_0_30 );
not g0002 ( new_n140_, keyIn_0_26 );
not g0003 ( new_n141_, N65 );
not g0004 ( new_n142_, N69 );
and g0005 ( new_n143_, new_n141_, new_n142_ );
and g0006 ( new_n144_, N65, N69 );
or g0007 ( new_n145_, new_n143_, new_n144_ );
not g0008 ( new_n146_, N77 );
and g0009 ( new_n147_, new_n146_, N73 );
not g0010 ( new_n148_, N73 );
and g0011 ( new_n149_, new_n148_, N77 );
or g0012 ( new_n150_, new_n147_, new_n149_ );
and g0013 ( new_n151_, new_n150_, keyIn_0_5 );
not g0014 ( new_n152_, keyIn_0_5 );
or g0015 ( new_n153_, new_n148_, N77 );
or g0016 ( new_n154_, new_n146_, N73 );
and g0017 ( new_n155_, new_n153_, new_n154_ );
and g0018 ( new_n156_, new_n155_, new_n152_ );
or g0019 ( new_n157_, new_n151_, new_n156_ );
or g0020 ( new_n158_, new_n157_, new_n145_ );
not g0021 ( new_n159_, new_n145_ );
or g0022 ( new_n160_, new_n155_, new_n152_ );
or g0023 ( new_n161_, new_n150_, keyIn_0_5 );
and g0024 ( new_n162_, new_n161_, new_n160_ );
or g0025 ( new_n163_, new_n162_, new_n159_ );
and g0026 ( new_n164_, new_n158_, new_n163_ );
or g0027 ( new_n165_, new_n164_, keyIn_0_10 );
not g0028 ( new_n166_, keyIn_0_10 );
and g0029 ( new_n167_, new_n162_, new_n159_ );
and g0030 ( new_n168_, new_n157_, new_n145_ );
or g0031 ( new_n169_, new_n168_, new_n167_ );
or g0032 ( new_n170_, new_n169_, new_n166_ );
and g0033 ( new_n171_, new_n170_, new_n165_ );
not g0034 ( new_n172_, keyIn_0_11 );
not g0035 ( new_n173_, N81 );
not g0036 ( new_n174_, N85 );
and g0037 ( new_n175_, new_n173_, new_n174_ );
and g0038 ( new_n176_, N81, N85 );
or g0039 ( new_n177_, new_n175_, new_n176_ );
not g0040 ( new_n178_, N89 );
not g0041 ( new_n179_, N93 );
and g0042 ( new_n180_, new_n178_, new_n179_ );
and g0043 ( new_n181_, N89, N93 );
or g0044 ( new_n182_, new_n180_, new_n181_ );
and g0045 ( new_n183_, new_n177_, new_n182_ );
not g0046 ( new_n184_, new_n183_ );
or g0047 ( new_n185_, new_n177_, new_n182_ );
and g0048 ( new_n186_, new_n184_, new_n185_ );
or g0049 ( new_n187_, new_n186_, new_n172_ );
and g0050 ( new_n188_, new_n186_, new_n172_ );
not g0051 ( new_n189_, new_n188_ );
and g0052 ( new_n190_, new_n189_, new_n187_ );
or g0053 ( new_n191_, new_n171_, new_n190_ );
and g0054 ( new_n192_, new_n169_, new_n166_ );
and g0055 ( new_n193_, new_n164_, keyIn_0_10 );
or g0056 ( new_n194_, new_n192_, new_n193_ );
not g0057 ( new_n195_, new_n190_ );
or g0058 ( new_n196_, new_n194_, new_n195_ );
and g0059 ( new_n197_, new_n196_, new_n191_ );
or g0060 ( new_n198_, new_n197_, new_n140_ );
and g0061 ( new_n199_, new_n194_, new_n195_ );
and g0062 ( new_n200_, new_n171_, new_n190_ );
or g0063 ( new_n201_, new_n199_, new_n200_ );
or g0064 ( new_n202_, new_n201_, keyIn_0_26 );
and g0065 ( new_n203_, new_n202_, new_n198_ );
and g0066 ( new_n204_, N129, N137 );
not g0067 ( new_n205_, new_n204_ );
or g0068 ( new_n206_, new_n203_, new_n205_ );
and g0069 ( new_n207_, new_n201_, keyIn_0_26 );
and g0070 ( new_n208_, new_n197_, new_n140_ );
or g0071 ( new_n209_, new_n207_, new_n208_ );
or g0072 ( new_n210_, new_n209_, new_n204_ );
and g0073 ( new_n211_, new_n210_, new_n206_ );
or g0074 ( new_n212_, new_n211_, new_n139_ );
and g0075 ( new_n213_, new_n209_, new_n204_ );
and g0076 ( new_n214_, new_n203_, new_n205_ );
or g0077 ( new_n215_, new_n213_, new_n214_ );
or g0078 ( new_n216_, new_n215_, keyIn_0_30 );
and g0079 ( new_n217_, new_n216_, new_n212_ );
not g0080 ( new_n218_, N1 );
not g0081 ( new_n219_, N17 );
and g0082 ( new_n220_, new_n218_, new_n219_ );
and g0083 ( new_n221_, N1, N17 );
or g0084 ( new_n222_, new_n220_, new_n221_ );
not g0085 ( new_n223_, N33 );
not g0086 ( new_n224_, N49 );
and g0087 ( new_n225_, new_n223_, new_n224_ );
and g0088 ( new_n226_, N33, N49 );
or g0089 ( new_n227_, new_n225_, new_n226_ );
and g0090 ( new_n228_, new_n222_, new_n227_ );
not g0091 ( new_n229_, new_n228_ );
or g0092 ( new_n230_, new_n222_, new_n227_ );
and g0093 ( new_n231_, new_n229_, new_n230_ );
not g0094 ( new_n232_, new_n231_ );
and g0095 ( new_n233_, new_n232_, keyIn_0_14 );
not g0096 ( new_n234_, new_n233_ );
or g0097 ( new_n235_, new_n232_, keyIn_0_14 );
and g0098 ( new_n236_, new_n234_, new_n235_ );
or g0099 ( new_n237_, new_n217_, new_n236_ );
and g0100 ( new_n238_, new_n215_, keyIn_0_30 );
and g0101 ( new_n239_, new_n211_, new_n139_ );
or g0102 ( new_n240_, new_n238_, new_n239_ );
not g0103 ( new_n241_, new_n236_ );
or g0104 ( new_n242_, new_n240_, new_n241_ );
and g0105 ( new_n243_, new_n242_, new_n237_ );
and g0106 ( new_n244_, new_n243_, new_n138_ );
and g0107 ( new_n245_, new_n240_, new_n241_ );
and g0108 ( new_n246_, new_n217_, new_n236_ );
or g0109 ( new_n247_, new_n245_, new_n246_ );
and g0110 ( new_n248_, new_n247_, keyIn_0_38 );
or g0111 ( new_n249_, new_n248_, new_n244_ );
not g0112 ( new_n250_, keyIn_0_56 );
not g0113 ( new_n251_, keyIn_0_54 );
not g0114 ( new_n252_, keyIn_0_48 );
not g0115 ( new_n253_, keyIn_0_33 );
not g0116 ( new_n254_, keyIn_0_29 );
not g0117 ( new_n255_, keyIn_0_13 );
not g0118 ( new_n256_, N117 );
and g0119 ( new_n257_, new_n256_, N113 );
not g0120 ( new_n258_, N113 );
and g0121 ( new_n259_, new_n258_, N117 );
or g0122 ( new_n260_, new_n257_, new_n259_ );
not g0123 ( new_n261_, N121 );
not g0124 ( new_n262_, N125 );
and g0125 ( new_n263_, new_n261_, new_n262_ );
and g0126 ( new_n264_, N121, N125 );
or g0127 ( new_n265_, new_n263_, new_n264_ );
and g0128 ( new_n266_, new_n260_, new_n265_ );
not g0129 ( new_n267_, new_n266_ );
or g0130 ( new_n268_, new_n260_, new_n265_ );
and g0131 ( new_n269_, new_n267_, new_n268_ );
and g0132 ( new_n270_, new_n269_, new_n255_ );
not g0133 ( new_n271_, new_n270_ );
or g0134 ( new_n272_, new_n269_, new_n255_ );
and g0135 ( new_n273_, new_n271_, new_n272_ );
and g0136 ( new_n274_, new_n273_, new_n190_ );
not g0137 ( new_n275_, new_n273_ );
and g0138 ( new_n276_, new_n275_, new_n195_ );
or g0139 ( new_n277_, new_n276_, new_n274_ );
not g0140 ( new_n278_, new_n277_ );
and g0141 ( new_n279_, new_n278_, new_n254_ );
and g0142 ( new_n280_, new_n277_, keyIn_0_29 );
or g0143 ( new_n281_, new_n279_, new_n280_ );
and g0144 ( new_n282_, N132, N137 );
and g0145 ( new_n283_, new_n281_, new_n282_ );
not g0146 ( new_n284_, new_n283_ );
or g0147 ( new_n285_, new_n281_, new_n282_ );
and g0148 ( new_n286_, new_n284_, new_n285_ );
or g0149 ( new_n287_, new_n286_, new_n253_ );
and g0150 ( new_n288_, new_n286_, new_n253_ );
not g0151 ( new_n289_, new_n288_ );
and g0152 ( new_n290_, new_n289_, new_n287_ );
not g0153 ( new_n291_, N29 );
and g0154 ( new_n292_, new_n291_, N13 );
not g0155 ( new_n293_, N13 );
and g0156 ( new_n294_, new_n293_, N29 );
or g0157 ( new_n295_, new_n292_, new_n294_ );
not g0158 ( new_n296_, N45 );
not g0159 ( new_n297_, N61 );
and g0160 ( new_n298_, new_n296_, new_n297_ );
and g0161 ( new_n299_, N45, N61 );
or g0162 ( new_n300_, new_n298_, new_n299_ );
and g0163 ( new_n301_, new_n295_, new_n300_ );
not g0164 ( new_n302_, new_n301_ );
or g0165 ( new_n303_, new_n295_, new_n300_ );
and g0166 ( new_n304_, new_n302_, new_n303_ );
not g0167 ( new_n305_, new_n304_ );
and g0168 ( new_n306_, new_n305_, keyIn_0_17 );
not g0169 ( new_n307_, new_n306_ );
or g0170 ( new_n308_, new_n305_, keyIn_0_17 );
and g0171 ( new_n309_, new_n307_, new_n308_ );
or g0172 ( new_n310_, new_n290_, new_n309_ );
not g0173 ( new_n311_, new_n285_ );
or g0174 ( new_n312_, new_n311_, new_n283_ );
and g0175 ( new_n313_, new_n312_, keyIn_0_33 );
or g0176 ( new_n314_, new_n313_, new_n288_ );
not g0177 ( new_n315_, new_n309_ );
or g0178 ( new_n316_, new_n314_, new_n315_ );
and g0179 ( new_n317_, new_n310_, new_n316_ );
or g0180 ( new_n318_, new_n317_, keyIn_0_41 );
not g0181 ( new_n319_, keyIn_0_41 );
and g0182 ( new_n320_, new_n314_, new_n315_ );
and g0183 ( new_n321_, new_n290_, new_n309_ );
or g0184 ( new_n322_, new_n321_, new_n320_ );
or g0185 ( new_n323_, new_n322_, new_n319_ );
and g0186 ( new_n324_, new_n323_, new_n318_ );
not g0187 ( new_n325_, keyIn_0_32 );
not g0188 ( new_n326_, keyIn_0_28 );
not g0189 ( new_n327_, N101 );
and g0190 ( new_n328_, new_n327_, N97 );
not g0191 ( new_n329_, N97 );
and g0192 ( new_n330_, new_n329_, N101 );
or g0193 ( new_n331_, new_n328_, new_n330_ );
not g0194 ( new_n332_, N105 );
not g0195 ( new_n333_, N109 );
and g0196 ( new_n334_, new_n332_, new_n333_ );
and g0197 ( new_n335_, N105, N109 );
or g0198 ( new_n336_, new_n334_, new_n335_ );
and g0199 ( new_n337_, new_n331_, new_n336_ );
not g0200 ( new_n338_, new_n337_ );
or g0201 ( new_n339_, new_n331_, new_n336_ );
and g0202 ( new_n340_, new_n338_, new_n339_ );
not g0203 ( new_n341_, new_n340_ );
and g0204 ( new_n342_, new_n341_, keyIn_0_12 );
not g0205 ( new_n343_, new_n342_ );
or g0206 ( new_n344_, new_n341_, keyIn_0_12 );
and g0207 ( new_n345_, new_n343_, new_n344_ );
or g0208 ( new_n346_, new_n171_, new_n345_ );
not g0209 ( new_n347_, new_n345_ );
or g0210 ( new_n348_, new_n194_, new_n347_ );
and g0211 ( new_n349_, new_n348_, new_n346_ );
or g0212 ( new_n350_, new_n349_, new_n326_ );
and g0213 ( new_n351_, new_n194_, new_n347_ );
and g0214 ( new_n352_, new_n171_, new_n345_ );
or g0215 ( new_n353_, new_n351_, new_n352_ );
or g0216 ( new_n354_, new_n353_, keyIn_0_28 );
and g0217 ( new_n355_, new_n354_, new_n350_ );
and g0218 ( new_n356_, N131, N137 );
not g0219 ( new_n357_, new_n356_ );
or g0220 ( new_n358_, new_n355_, new_n357_ );
and g0221 ( new_n359_, new_n353_, keyIn_0_28 );
and g0222 ( new_n360_, new_n349_, new_n326_ );
or g0223 ( new_n361_, new_n359_, new_n360_ );
or g0224 ( new_n362_, new_n361_, new_n356_ );
and g0225 ( new_n363_, new_n362_, new_n358_ );
or g0226 ( new_n364_, new_n363_, new_n325_ );
and g0227 ( new_n365_, new_n361_, new_n356_ );
and g0228 ( new_n366_, new_n355_, new_n357_ );
or g0229 ( new_n367_, new_n365_, new_n366_ );
or g0230 ( new_n368_, new_n367_, keyIn_0_32 );
and g0231 ( new_n369_, new_n368_, new_n364_ );
not g0232 ( new_n370_, N9 );
not g0233 ( new_n371_, N25 );
and g0234 ( new_n372_, new_n370_, new_n371_ );
and g0235 ( new_n373_, N9, N25 );
or g0236 ( new_n374_, new_n372_, new_n373_ );
not g0237 ( new_n375_, N41 );
not g0238 ( new_n376_, N57 );
and g0239 ( new_n377_, new_n375_, new_n376_ );
and g0240 ( new_n378_, N41, N57 );
or g0241 ( new_n379_, new_n377_, new_n378_ );
and g0242 ( new_n380_, new_n374_, new_n379_ );
not g0243 ( new_n381_, new_n380_ );
or g0244 ( new_n382_, new_n374_, new_n379_ );
and g0245 ( new_n383_, new_n381_, new_n382_ );
not g0246 ( new_n384_, new_n383_ );
and g0247 ( new_n385_, new_n384_, keyIn_0_16 );
not g0248 ( new_n386_, new_n385_ );
or g0249 ( new_n387_, new_n384_, keyIn_0_16 );
and g0250 ( new_n388_, new_n386_, new_n387_ );
or g0251 ( new_n389_, new_n369_, new_n388_ );
and g0252 ( new_n390_, new_n367_, keyIn_0_32 );
and g0253 ( new_n391_, new_n363_, new_n325_ );
or g0254 ( new_n392_, new_n390_, new_n391_ );
not g0255 ( new_n393_, new_n388_ );
or g0256 ( new_n394_, new_n392_, new_n393_ );
and g0257 ( new_n395_, new_n394_, new_n389_ );
and g0258 ( new_n396_, new_n395_, keyIn_0_40 );
not g0259 ( new_n397_, keyIn_0_40 );
and g0260 ( new_n398_, new_n392_, new_n393_ );
and g0261 ( new_n399_, new_n369_, new_n388_ );
or g0262 ( new_n400_, new_n398_, new_n399_ );
and g0263 ( new_n401_, new_n400_, new_n397_ );
or g0264 ( new_n402_, new_n401_, new_n396_ );
and g0265 ( new_n403_, new_n249_, new_n402_ );
not g0266 ( new_n404_, keyIn_0_31 );
and g0267 ( new_n405_, new_n345_, new_n273_ );
and g0268 ( new_n406_, new_n347_, new_n275_ );
or g0269 ( new_n407_, new_n406_, new_n405_ );
or g0270 ( new_n408_, new_n407_, keyIn_0_27 );
and g0271 ( new_n409_, new_n407_, keyIn_0_27 );
not g0272 ( new_n410_, new_n409_ );
and g0273 ( new_n411_, new_n410_, new_n408_ );
and g0274 ( new_n412_, N130, N137 );
not g0275 ( new_n413_, new_n412_ );
or g0276 ( new_n414_, new_n411_, new_n413_ );
not g0277 ( new_n415_, keyIn_0_27 );
not g0278 ( new_n416_, new_n407_ );
and g0279 ( new_n417_, new_n416_, new_n415_ );
or g0280 ( new_n418_, new_n417_, new_n409_ );
or g0281 ( new_n419_, new_n418_, new_n412_ );
and g0282 ( new_n420_, new_n419_, new_n414_ );
or g0283 ( new_n421_, new_n420_, new_n404_ );
and g0284 ( new_n422_, new_n418_, new_n412_ );
and g0285 ( new_n423_, new_n411_, new_n413_ );
or g0286 ( new_n424_, new_n422_, new_n423_ );
or g0287 ( new_n425_, new_n424_, keyIn_0_31 );
and g0288 ( new_n426_, new_n425_, new_n421_ );
not g0289 ( new_n427_, N37 );
not g0290 ( new_n428_, N53 );
and g0291 ( new_n429_, new_n427_, new_n428_ );
and g0292 ( new_n430_, N37, N53 );
or g0293 ( new_n431_, new_n429_, new_n430_ );
not g0294 ( new_n432_, new_n431_ );
not g0295 ( new_n433_, N5 );
not g0296 ( new_n434_, N21 );
and g0297 ( new_n435_, new_n433_, new_n434_ );
and g0298 ( new_n436_, N5, N21 );
or g0299 ( new_n437_, new_n435_, new_n436_ );
and g0300 ( new_n438_, new_n432_, new_n437_ );
not g0301 ( new_n439_, new_n438_ );
or g0302 ( new_n440_, new_n432_, new_n437_ );
and g0303 ( new_n441_, new_n439_, new_n440_ );
not g0304 ( new_n442_, new_n441_ );
and g0305 ( new_n443_, new_n442_, keyIn_0_15 );
not g0306 ( new_n444_, new_n443_ );
or g0307 ( new_n445_, new_n442_, keyIn_0_15 );
and g0308 ( new_n446_, new_n444_, new_n445_ );
or g0309 ( new_n447_, new_n426_, new_n446_ );
and g0310 ( new_n448_, new_n424_, keyIn_0_31 );
and g0311 ( new_n449_, new_n420_, new_n404_ );
or g0312 ( new_n450_, new_n448_, new_n449_ );
not g0313 ( new_n451_, new_n446_ );
or g0314 ( new_n452_, new_n450_, new_n451_ );
and g0315 ( new_n453_, new_n452_, new_n447_ );
and g0316 ( new_n454_, new_n453_, keyIn_0_39 );
not g0317 ( new_n455_, keyIn_0_39 );
and g0318 ( new_n456_, new_n450_, new_n451_ );
and g0319 ( new_n457_, new_n426_, new_n446_ );
or g0320 ( new_n458_, new_n456_, new_n457_ );
and g0321 ( new_n459_, new_n458_, new_n455_ );
or g0322 ( new_n460_, new_n459_, new_n454_ );
and g0323 ( new_n461_, new_n403_, new_n460_ );
and g0324 ( new_n462_, new_n461_, new_n324_ );
and g0325 ( new_n463_, new_n462_, new_n252_ );
not g0326 ( new_n464_, new_n463_ );
or g0327 ( new_n465_, new_n462_, new_n252_ );
and g0328 ( new_n466_, new_n464_, new_n465_ );
not g0329 ( new_n467_, new_n244_ );
or g0330 ( new_n468_, new_n243_, new_n138_ );
and g0331 ( new_n469_, new_n467_, new_n468_ );
or g0332 ( new_n470_, new_n400_, new_n397_ );
or g0333 ( new_n471_, new_n395_, keyIn_0_40 );
and g0334 ( new_n472_, new_n470_, new_n471_ );
or g0335 ( new_n473_, new_n469_, new_n472_ );
or g0336 ( new_n474_, new_n324_, new_n460_ );
or g0337 ( new_n475_, new_n473_, new_n474_ );
or g0338 ( new_n476_, new_n475_, keyIn_0_46 );
not g0339 ( new_n477_, keyIn_0_46 );
and g0340 ( new_n478_, new_n322_, new_n319_ );
and g0341 ( new_n479_, new_n317_, keyIn_0_41 );
or g0342 ( new_n480_, new_n478_, new_n479_ );
not g0343 ( new_n481_, new_n460_ );
and g0344 ( new_n482_, new_n481_, new_n480_ );
and g0345 ( new_n483_, new_n482_, new_n403_ );
or g0346 ( new_n484_, new_n483_, new_n477_ );
and g0347 ( new_n485_, new_n476_, new_n484_ );
and g0348 ( new_n486_, new_n472_, new_n324_ );
and g0349 ( new_n487_, new_n486_, new_n249_ );
and g0350 ( new_n488_, new_n481_, keyIn_0_47 );
and g0351 ( new_n489_, new_n487_, new_n488_ );
not g0352 ( new_n490_, new_n489_ );
and g0353 ( new_n491_, new_n481_, new_n249_ );
and g0354 ( new_n492_, new_n491_, new_n486_ );
or g0355 ( new_n493_, new_n492_, keyIn_0_47 );
and g0356 ( new_n494_, new_n490_, new_n493_ );
or g0357 ( new_n495_, new_n485_, new_n494_ );
or g0358 ( new_n496_, new_n249_, new_n460_ );
or g0359 ( new_n497_, new_n496_, new_n472_ );
or g0360 ( new_n498_, new_n497_, new_n480_ );
and g0361 ( new_n499_, new_n498_, keyIn_0_49 );
not g0362 ( new_n500_, keyIn_0_49 );
and g0363 ( new_n501_, new_n481_, new_n469_ );
and g0364 ( new_n502_, new_n501_, new_n402_ );
and g0365 ( new_n503_, new_n502_, new_n324_ );
and g0366 ( new_n504_, new_n503_, new_n500_ );
or g0367 ( new_n505_, new_n499_, new_n504_ );
or g0368 ( new_n506_, new_n495_, new_n505_ );
or g0369 ( new_n507_, new_n506_, new_n466_ );
or g0370 ( new_n508_, new_n507_, new_n251_ );
not g0371 ( new_n509_, new_n466_ );
and g0372 ( new_n510_, new_n483_, new_n477_ );
and g0373 ( new_n511_, new_n475_, keyIn_0_46 );
or g0374 ( new_n512_, new_n511_, new_n510_ );
not g0375 ( new_n513_, keyIn_0_47 );
or g0376 ( new_n514_, new_n402_, new_n480_ );
or g0377 ( new_n515_, new_n469_, new_n460_ );
or g0378 ( new_n516_, new_n515_, new_n514_ );
and g0379 ( new_n517_, new_n516_, new_n513_ );
or g0380 ( new_n518_, new_n517_, new_n489_ );
and g0381 ( new_n519_, new_n512_, new_n518_ );
or g0382 ( new_n520_, new_n503_, new_n500_ );
not g0383 ( new_n521_, new_n504_ );
and g0384 ( new_n522_, new_n521_, new_n520_ );
and g0385 ( new_n523_, new_n522_, new_n519_ );
and g0386 ( new_n524_, new_n523_, new_n509_ );
or g0387 ( new_n525_, new_n524_, keyIn_0_54 );
and g0388 ( new_n526_, new_n508_, new_n525_ );
not g0389 ( new_n527_, keyIn_0_44 );
not g0390 ( new_n528_, keyIn_0_36 );
not g0391 ( new_n529_, keyIn_0_24 );
and g0392 ( new_n530_, new_n223_, new_n427_ );
and g0393 ( new_n531_, N33, N37 );
or g0394 ( new_n532_, new_n530_, new_n531_ );
and g0395 ( new_n533_, new_n532_, keyIn_0_1 );
not g0396 ( new_n534_, new_n531_ );
not g0397 ( new_n535_, keyIn_0_1 );
or g0398 ( new_n536_, N33, N37 );
and g0399 ( new_n537_, new_n536_, new_n535_ );
and g0400 ( new_n538_, new_n537_, new_n534_ );
or g0401 ( new_n539_, new_n533_, new_n538_ );
and g0402 ( new_n540_, new_n375_, new_n296_ );
and g0403 ( new_n541_, N41, N45 );
or g0404 ( new_n542_, new_n540_, new_n541_ );
and g0405 ( new_n543_, new_n542_, keyIn_0_2 );
not g0406 ( new_n544_, keyIn_0_2 );
or g0407 ( new_n545_, N41, N45 );
not g0408 ( new_n546_, new_n541_ );
and g0409 ( new_n547_, new_n546_, new_n545_ );
and g0410 ( new_n548_, new_n547_, new_n544_ );
or g0411 ( new_n549_, new_n543_, new_n548_ );
or g0412 ( new_n550_, new_n549_, new_n539_ );
and g0413 ( new_n551_, new_n534_, new_n536_ );
or g0414 ( new_n552_, new_n551_, new_n535_ );
not g0415 ( new_n553_, new_n538_ );
and g0416 ( new_n554_, new_n553_, new_n552_ );
or g0417 ( new_n555_, new_n547_, new_n544_ );
or g0418 ( new_n556_, new_n542_, keyIn_0_2 );
and g0419 ( new_n557_, new_n556_, new_n555_ );
or g0420 ( new_n558_, new_n557_, new_n554_ );
and g0421 ( new_n559_, new_n550_, new_n558_ );
and g0422 ( new_n560_, new_n559_, keyIn_0_8 );
not g0423 ( new_n561_, keyIn_0_8 );
and g0424 ( new_n562_, new_n557_, new_n554_ );
and g0425 ( new_n563_, new_n549_, new_n539_ );
or g0426 ( new_n564_, new_n563_, new_n562_ );
and g0427 ( new_n565_, new_n564_, new_n561_ );
or g0428 ( new_n566_, new_n560_, new_n565_ );
and g0429 ( new_n567_, new_n218_, new_n433_ );
and g0430 ( new_n568_, N1, N5 );
or g0431 ( new_n569_, new_n567_, new_n568_ );
and g0432 ( new_n570_, new_n370_, new_n293_ );
and g0433 ( new_n571_, N9, N13 );
or g0434 ( new_n572_, new_n570_, new_n571_ );
and g0435 ( new_n573_, new_n569_, new_n572_ );
not g0436 ( new_n574_, new_n573_ );
or g0437 ( new_n575_, new_n569_, new_n572_ );
and g0438 ( new_n576_, new_n574_, new_n575_ );
not g0439 ( new_n577_, new_n576_ );
and g0440 ( new_n578_, new_n577_, keyIn_0_6 );
not g0441 ( new_n579_, new_n578_ );
or g0442 ( new_n580_, new_n577_, keyIn_0_6 );
and g0443 ( new_n581_, new_n579_, new_n580_ );
not g0444 ( new_n582_, new_n581_ );
and g0445 ( new_n583_, new_n566_, new_n582_ );
or g0446 ( new_n584_, new_n564_, new_n561_ );
or g0447 ( new_n585_, new_n559_, keyIn_0_8 );
and g0448 ( new_n586_, new_n584_, new_n585_ );
and g0449 ( new_n587_, new_n586_, new_n581_ );
or g0450 ( new_n588_, new_n583_, new_n587_ );
and g0451 ( new_n589_, new_n588_, new_n529_ );
or g0452 ( new_n590_, new_n586_, new_n581_ );
or g0453 ( new_n591_, new_n566_, new_n582_ );
and g0454 ( new_n592_, new_n591_, new_n590_ );
and g0455 ( new_n593_, new_n592_, keyIn_0_24 );
or g0456 ( new_n594_, new_n589_, new_n593_ );
and g0457 ( new_n595_, N135, N137 );
or g0458 ( new_n596_, new_n594_, new_n595_ );
or g0459 ( new_n597_, new_n592_, keyIn_0_24 );
or g0460 ( new_n598_, new_n588_, new_n529_ );
and g0461 ( new_n599_, new_n598_, new_n597_ );
not g0462 ( new_n600_, new_n595_ );
or g0463 ( new_n601_, new_n599_, new_n600_ );
and g0464 ( new_n602_, new_n596_, new_n601_ );
and g0465 ( new_n603_, new_n602_, new_n528_ );
and g0466 ( new_n604_, new_n599_, new_n600_ );
and g0467 ( new_n605_, new_n594_, new_n595_ );
or g0468 ( new_n606_, new_n605_, new_n604_ );
and g0469 ( new_n607_, new_n606_, keyIn_0_36 );
or g0470 ( new_n608_, new_n607_, new_n603_ );
and g0471 ( new_n609_, new_n178_, N73 );
and g0472 ( new_n610_, new_n148_, N89 );
or g0473 ( new_n611_, new_n609_, new_n610_ );
and g0474 ( new_n612_, new_n332_, new_n261_ );
and g0475 ( new_n613_, N105, N121 );
or g0476 ( new_n614_, new_n612_, new_n613_ );
and g0477 ( new_n615_, new_n611_, new_n614_ );
not g0478 ( new_n616_, new_n615_ );
or g0479 ( new_n617_, new_n611_, new_n614_ );
and g0480 ( new_n618_, new_n616_, new_n617_ );
not g0481 ( new_n619_, new_n618_ );
and g0482 ( new_n620_, new_n619_, keyIn_0_20 );
not g0483 ( new_n621_, new_n620_ );
or g0484 ( new_n622_, new_n619_, keyIn_0_20 );
and g0485 ( new_n623_, new_n621_, new_n622_ );
not g0486 ( new_n624_, new_n623_ );
and g0487 ( new_n625_, new_n608_, new_n624_ );
or g0488 ( new_n626_, new_n606_, keyIn_0_36 );
or g0489 ( new_n627_, new_n602_, new_n528_ );
and g0490 ( new_n628_, new_n626_, new_n627_ );
and g0491 ( new_n629_, new_n628_, new_n623_ );
or g0492 ( new_n630_, new_n625_, new_n629_ );
and g0493 ( new_n631_, new_n630_, new_n527_ );
or g0494 ( new_n632_, new_n628_, new_n623_ );
or g0495 ( new_n633_, new_n608_, new_n624_ );
and g0496 ( new_n634_, new_n633_, new_n632_ );
and g0497 ( new_n635_, new_n634_, keyIn_0_44 );
or g0498 ( new_n636_, new_n631_, new_n635_ );
not g0499 ( new_n637_, keyIn_0_45 );
not g0500 ( new_n638_, keyIn_0_37 );
not g0501 ( new_n639_, keyIn_0_25 );
not g0502 ( new_n640_, keyIn_0_3 );
or g0503 ( new_n641_, N49, N53 );
and g0504 ( new_n642_, N49, N53 );
not g0505 ( new_n643_, new_n642_ );
and g0506 ( new_n644_, new_n643_, new_n641_ );
or g0507 ( new_n645_, new_n644_, new_n640_ );
and g0508 ( new_n646_, new_n641_, new_n640_ );
and g0509 ( new_n647_, new_n646_, new_n643_ );
not g0510 ( new_n648_, new_n647_ );
and g0511 ( new_n649_, new_n648_, new_n645_ );
not g0512 ( new_n650_, keyIn_0_4 );
or g0513 ( new_n651_, N57, N61 );
and g0514 ( new_n652_, N57, N61 );
not g0515 ( new_n653_, new_n652_ );
and g0516 ( new_n654_, new_n653_, new_n651_ );
or g0517 ( new_n655_, new_n654_, new_n650_ );
and g0518 ( new_n656_, new_n376_, new_n297_ );
or g0519 ( new_n657_, new_n656_, new_n652_ );
or g0520 ( new_n658_, new_n657_, keyIn_0_4 );
and g0521 ( new_n659_, new_n658_, new_n655_ );
and g0522 ( new_n660_, new_n659_, new_n649_ );
and g0523 ( new_n661_, new_n224_, new_n428_ );
or g0524 ( new_n662_, new_n661_, new_n642_ );
and g0525 ( new_n663_, new_n662_, keyIn_0_3 );
or g0526 ( new_n664_, new_n663_, new_n647_ );
and g0527 ( new_n665_, new_n657_, keyIn_0_4 );
and g0528 ( new_n666_, new_n654_, new_n650_ );
or g0529 ( new_n667_, new_n665_, new_n666_ );
and g0530 ( new_n668_, new_n667_, new_n664_ );
or g0531 ( new_n669_, new_n668_, new_n660_ );
and g0532 ( new_n670_, new_n669_, keyIn_0_9 );
not g0533 ( new_n671_, keyIn_0_9 );
or g0534 ( new_n672_, new_n667_, new_n664_ );
or g0535 ( new_n673_, new_n659_, new_n649_ );
and g0536 ( new_n674_, new_n672_, new_n673_ );
and g0537 ( new_n675_, new_n674_, new_n671_ );
or g0538 ( new_n676_, new_n670_, new_n675_ );
and g0539 ( new_n677_, new_n371_, new_n291_ );
and g0540 ( new_n678_, N25, N29 );
or g0541 ( new_n679_, new_n677_, new_n678_ );
not g0542 ( new_n680_, new_n679_ );
not g0543 ( new_n681_, keyIn_0_0 );
or g0544 ( new_n682_, new_n219_, N21 );
or g0545 ( new_n683_, new_n434_, N17 );
and g0546 ( new_n684_, new_n682_, new_n683_ );
or g0547 ( new_n685_, new_n684_, new_n681_ );
and g0548 ( new_n686_, new_n434_, N17 );
and g0549 ( new_n687_, new_n219_, N21 );
or g0550 ( new_n688_, new_n686_, new_n687_ );
or g0551 ( new_n689_, new_n688_, keyIn_0_0 );
and g0552 ( new_n690_, new_n689_, new_n685_ );
and g0553 ( new_n691_, new_n690_, new_n680_ );
and g0554 ( new_n692_, new_n688_, keyIn_0_0 );
and g0555 ( new_n693_, new_n684_, new_n681_ );
or g0556 ( new_n694_, new_n692_, new_n693_ );
and g0557 ( new_n695_, new_n694_, new_n679_ );
or g0558 ( new_n696_, new_n695_, new_n691_ );
and g0559 ( new_n697_, new_n696_, keyIn_0_7 );
not g0560 ( new_n698_, keyIn_0_7 );
or g0561 ( new_n699_, new_n694_, new_n679_ );
or g0562 ( new_n700_, new_n690_, new_n680_ );
and g0563 ( new_n701_, new_n699_, new_n700_ );
and g0564 ( new_n702_, new_n701_, new_n698_ );
or g0565 ( new_n703_, new_n697_, new_n702_ );
and g0566 ( new_n704_, new_n676_, new_n703_ );
or g0567 ( new_n705_, new_n674_, new_n671_ );
or g0568 ( new_n706_, new_n669_, keyIn_0_9 );
and g0569 ( new_n707_, new_n705_, new_n706_ );
or g0570 ( new_n708_, new_n701_, new_n698_ );
or g0571 ( new_n709_, new_n696_, keyIn_0_7 );
and g0572 ( new_n710_, new_n709_, new_n708_ );
and g0573 ( new_n711_, new_n710_, new_n707_ );
or g0574 ( new_n712_, new_n704_, new_n711_ );
and g0575 ( new_n713_, new_n712_, new_n639_ );
or g0576 ( new_n714_, new_n710_, new_n707_ );
or g0577 ( new_n715_, new_n676_, new_n703_ );
and g0578 ( new_n716_, new_n715_, new_n714_ );
and g0579 ( new_n717_, new_n716_, keyIn_0_25 );
or g0580 ( new_n718_, new_n717_, new_n713_ );
and g0581 ( new_n719_, N136, N137 );
or g0582 ( new_n720_, new_n718_, new_n719_ );
or g0583 ( new_n721_, new_n716_, keyIn_0_25 );
or g0584 ( new_n722_, new_n712_, new_n639_ );
and g0585 ( new_n723_, new_n721_, new_n722_ );
not g0586 ( new_n724_, new_n719_ );
or g0587 ( new_n725_, new_n723_, new_n724_ );
and g0588 ( new_n726_, new_n720_, new_n725_ );
and g0589 ( new_n727_, new_n726_, new_n638_ );
and g0590 ( new_n728_, new_n723_, new_n724_ );
and g0591 ( new_n729_, new_n718_, new_n719_ );
or g0592 ( new_n730_, new_n729_, new_n728_ );
and g0593 ( new_n731_, new_n730_, keyIn_0_37 );
or g0594 ( new_n732_, new_n731_, new_n727_ );
not g0595 ( new_n733_, keyIn_0_21 );
and g0596 ( new_n734_, new_n179_, N77 );
and g0597 ( new_n735_, new_n146_, N93 );
or g0598 ( new_n736_, new_n734_, new_n735_ );
and g0599 ( new_n737_, new_n333_, new_n262_ );
and g0600 ( new_n738_, N109, N125 );
or g0601 ( new_n739_, new_n737_, new_n738_ );
and g0602 ( new_n740_, new_n736_, new_n739_ );
not g0603 ( new_n741_, new_n740_ );
or g0604 ( new_n742_, new_n736_, new_n739_ );
and g0605 ( new_n743_, new_n741_, new_n742_ );
not g0606 ( new_n744_, new_n743_ );
and g0607 ( new_n745_, new_n744_, new_n733_ );
and g0608 ( new_n746_, new_n743_, keyIn_0_21 );
or g0609 ( new_n747_, new_n745_, new_n746_ );
and g0610 ( new_n748_, new_n732_, new_n747_ );
or g0611 ( new_n749_, new_n730_, keyIn_0_37 );
or g0612 ( new_n750_, new_n726_, new_n638_ );
and g0613 ( new_n751_, new_n749_, new_n750_ );
not g0614 ( new_n752_, new_n747_ );
and g0615 ( new_n753_, new_n751_, new_n752_ );
or g0616 ( new_n754_, new_n748_, new_n753_ );
and g0617 ( new_n755_, new_n754_, new_n637_ );
or g0618 ( new_n756_, new_n751_, new_n752_ );
or g0619 ( new_n757_, new_n732_, new_n747_ );
and g0620 ( new_n758_, new_n757_, new_n756_ );
and g0621 ( new_n759_, new_n758_, keyIn_0_45 );
or g0622 ( new_n760_, new_n755_, new_n759_ );
and g0623 ( new_n761_, new_n760_, new_n636_ );
or g0624 ( new_n762_, new_n566_, new_n676_ );
or g0625 ( new_n763_, new_n586_, new_n707_ );
and g0626 ( new_n764_, new_n762_, new_n763_ );
and g0627 ( new_n765_, new_n764_, keyIn_0_23 );
not g0628 ( new_n766_, keyIn_0_23 );
and g0629 ( new_n767_, new_n586_, new_n707_ );
and g0630 ( new_n768_, new_n566_, new_n676_ );
or g0631 ( new_n769_, new_n768_, new_n767_ );
and g0632 ( new_n770_, new_n769_, new_n766_ );
or g0633 ( new_n771_, new_n765_, new_n770_ );
and g0634 ( new_n772_, N134, N137 );
and g0635 ( new_n773_, new_n771_, new_n772_ );
or g0636 ( new_n774_, new_n769_, new_n766_ );
or g0637 ( new_n775_, new_n764_, keyIn_0_23 );
and g0638 ( new_n776_, new_n775_, new_n774_ );
not g0639 ( new_n777_, new_n772_ );
and g0640 ( new_n778_, new_n776_, new_n777_ );
or g0641 ( new_n779_, new_n773_, new_n778_ );
and g0642 ( new_n780_, new_n779_, keyIn_0_35 );
not g0643 ( new_n781_, keyIn_0_35 );
or g0644 ( new_n782_, new_n776_, new_n777_ );
or g0645 ( new_n783_, new_n771_, new_n772_ );
and g0646 ( new_n784_, new_n783_, new_n782_ );
and g0647 ( new_n785_, new_n784_, new_n781_ );
or g0648 ( new_n786_, new_n780_, new_n785_ );
and g0649 ( new_n787_, new_n142_, new_n174_ );
and g0650 ( new_n788_, N69, N85 );
or g0651 ( new_n789_, new_n787_, new_n788_ );
and g0652 ( new_n790_, new_n327_, new_n256_ );
and g0653 ( new_n791_, N101, N117 );
or g0654 ( new_n792_, new_n790_, new_n791_ );
and g0655 ( new_n793_, new_n789_, new_n792_ );
not g0656 ( new_n794_, new_n793_ );
or g0657 ( new_n795_, new_n789_, new_n792_ );
and g0658 ( new_n796_, new_n794_, new_n795_ );
not g0659 ( new_n797_, new_n796_ );
and g0660 ( new_n798_, new_n797_, keyIn_0_19 );
not g0661 ( new_n799_, new_n798_ );
or g0662 ( new_n800_, new_n797_, keyIn_0_19 );
and g0663 ( new_n801_, new_n799_, new_n800_ );
not g0664 ( new_n802_, new_n801_ );
and g0665 ( new_n803_, new_n786_, new_n802_ );
or g0666 ( new_n804_, new_n784_, new_n781_ );
or g0667 ( new_n805_, new_n779_, keyIn_0_35 );
and g0668 ( new_n806_, new_n805_, new_n804_ );
and g0669 ( new_n807_, new_n806_, new_n801_ );
or g0670 ( new_n808_, new_n803_, new_n807_ );
and g0671 ( new_n809_, new_n808_, keyIn_0_43 );
not g0672 ( new_n810_, keyIn_0_43 );
or g0673 ( new_n811_, new_n806_, new_n801_ );
or g0674 ( new_n812_, new_n786_, new_n802_ );
and g0675 ( new_n813_, new_n812_, new_n811_ );
and g0676 ( new_n814_, new_n813_, new_n810_ );
or g0677 ( new_n815_, new_n809_, new_n814_ );
not g0678 ( new_n816_, keyIn_0_42 );
not g0679 ( new_n817_, keyIn_0_22 );
and g0680 ( new_n818_, new_n703_, new_n582_ );
and g0681 ( new_n819_, new_n710_, new_n581_ );
or g0682 ( new_n820_, new_n818_, new_n819_ );
and g0683 ( new_n821_, new_n820_, new_n817_ );
or g0684 ( new_n822_, new_n710_, new_n581_ );
or g0685 ( new_n823_, new_n703_, new_n582_ );
and g0686 ( new_n824_, new_n823_, new_n822_ );
and g0687 ( new_n825_, new_n824_, keyIn_0_22 );
or g0688 ( new_n826_, new_n821_, new_n825_ );
and g0689 ( new_n827_, N133, N137 );
and g0690 ( new_n828_, new_n826_, new_n827_ );
or g0691 ( new_n829_, new_n824_, keyIn_0_22 );
or g0692 ( new_n830_, new_n820_, new_n817_ );
and g0693 ( new_n831_, new_n830_, new_n829_ );
not g0694 ( new_n832_, new_n827_ );
and g0695 ( new_n833_, new_n831_, new_n832_ );
or g0696 ( new_n834_, new_n828_, new_n833_ );
and g0697 ( new_n835_, new_n834_, keyIn_0_34 );
not g0698 ( new_n836_, keyIn_0_34 );
or g0699 ( new_n837_, new_n831_, new_n832_ );
or g0700 ( new_n838_, new_n826_, new_n827_ );
and g0701 ( new_n839_, new_n838_, new_n837_ );
and g0702 ( new_n840_, new_n839_, new_n836_ );
or g0703 ( new_n841_, new_n835_, new_n840_ );
and g0704 ( new_n842_, new_n141_, new_n173_ );
and g0705 ( new_n843_, N65, N81 );
or g0706 ( new_n844_, new_n842_, new_n843_ );
and g0707 ( new_n845_, new_n329_, new_n258_ );
and g0708 ( new_n846_, N97, N113 );
or g0709 ( new_n847_, new_n845_, new_n846_ );
and g0710 ( new_n848_, new_n844_, new_n847_ );
not g0711 ( new_n849_, new_n848_ );
or g0712 ( new_n850_, new_n844_, new_n847_ );
and g0713 ( new_n851_, new_n849_, new_n850_ );
not g0714 ( new_n852_, new_n851_ );
and g0715 ( new_n853_, new_n852_, keyIn_0_18 );
not g0716 ( new_n854_, new_n853_ );
or g0717 ( new_n855_, new_n852_, keyIn_0_18 );
and g0718 ( new_n856_, new_n854_, new_n855_ );
not g0719 ( new_n857_, new_n856_ );
and g0720 ( new_n858_, new_n841_, new_n857_ );
or g0721 ( new_n859_, new_n839_, new_n836_ );
or g0722 ( new_n860_, new_n834_, keyIn_0_34 );
and g0723 ( new_n861_, new_n860_, new_n859_ );
and g0724 ( new_n862_, new_n861_, new_n856_ );
or g0725 ( new_n863_, new_n858_, new_n862_ );
and g0726 ( new_n864_, new_n863_, new_n816_ );
or g0727 ( new_n865_, new_n861_, new_n856_ );
or g0728 ( new_n866_, new_n841_, new_n857_ );
and g0729 ( new_n867_, new_n866_, new_n865_ );
and g0730 ( new_n868_, new_n867_, keyIn_0_42 );
or g0731 ( new_n869_, new_n864_, new_n868_ );
and g0732 ( new_n870_, new_n815_, new_n869_ );
and g0733 ( new_n871_, new_n761_, new_n870_ );
not g0734 ( new_n872_, new_n871_ );
or g0735 ( new_n873_, new_n526_, new_n872_ );
or g0736 ( new_n874_, new_n873_, new_n250_ );
and g0737 ( new_n875_, new_n524_, keyIn_0_54 );
and g0738 ( new_n876_, new_n507_, new_n251_ );
or g0739 ( new_n877_, new_n876_, new_n875_ );
and g0740 ( new_n878_, new_n877_, new_n871_ );
or g0741 ( new_n879_, new_n878_, keyIn_0_56 );
and g0742 ( new_n880_, new_n874_, new_n879_ );
or g0743 ( new_n881_, new_n880_, new_n249_ );
and g0744 ( new_n882_, new_n881_, N1 );
and g0745 ( new_n883_, new_n878_, keyIn_0_56 );
and g0746 ( new_n884_, new_n873_, new_n250_ );
or g0747 ( new_n885_, new_n884_, new_n883_ );
and g0748 ( new_n886_, new_n885_, new_n469_ );
and g0749 ( new_n887_, new_n886_, new_n218_ );
or g0750 ( N724, new_n882_, new_n887_ );
or g0751 ( new_n889_, new_n880_, new_n481_ );
and g0752 ( new_n890_, new_n889_, N5 );
and g0753 ( new_n891_, new_n885_, new_n460_ );
and g0754 ( new_n892_, new_n891_, new_n433_ );
or g0755 ( N725, new_n890_, new_n892_ );
or g0756 ( new_n894_, new_n880_, new_n402_ );
and g0757 ( new_n895_, new_n894_, N9 );
and g0758 ( new_n896_, new_n885_, new_n472_ );
and g0759 ( new_n897_, new_n896_, new_n370_ );
or g0760 ( N726, new_n895_, new_n897_ );
or g0761 ( new_n899_, new_n880_, new_n324_ );
and g0762 ( new_n900_, new_n899_, N13 );
and g0763 ( new_n901_, new_n885_, new_n480_ );
and g0764 ( new_n902_, new_n901_, new_n293_ );
or g0765 ( N727, new_n900_, new_n902_ );
not g0766 ( new_n904_, keyIn_0_57 );
or g0767 ( new_n905_, new_n758_, keyIn_0_45 );
or g0768 ( new_n906_, new_n754_, new_n637_ );
and g0769 ( new_n907_, new_n906_, new_n905_ );
or g0770 ( new_n908_, new_n634_, keyIn_0_44 );
not g0771 ( new_n909_, new_n635_ );
and g0772 ( new_n910_, new_n909_, new_n908_ );
and g0773 ( new_n911_, new_n870_, new_n910_ );
and g0774 ( new_n912_, new_n911_, new_n907_ );
not g0775 ( new_n913_, new_n912_ );
or g0776 ( new_n914_, new_n526_, new_n913_ );
or g0777 ( new_n915_, new_n914_, new_n904_ );
and g0778 ( new_n916_, new_n877_, new_n912_ );
or g0779 ( new_n917_, new_n916_, keyIn_0_57 );
and g0780 ( new_n918_, new_n915_, new_n917_ );
or g0781 ( new_n919_, new_n918_, new_n249_ );
and g0782 ( new_n920_, new_n919_, N17 );
and g0783 ( new_n921_, new_n916_, keyIn_0_57 );
and g0784 ( new_n922_, new_n914_, new_n904_ );
or g0785 ( new_n923_, new_n922_, new_n921_ );
and g0786 ( new_n924_, new_n923_, new_n469_ );
and g0787 ( new_n925_, new_n924_, new_n219_ );
or g0788 ( N728, new_n920_, new_n925_ );
or g0789 ( new_n927_, new_n918_, new_n481_ );
and g0790 ( new_n928_, new_n927_, N21 );
and g0791 ( new_n929_, new_n923_, new_n460_ );
and g0792 ( new_n930_, new_n929_, new_n434_ );
or g0793 ( N729, new_n928_, new_n930_ );
or g0794 ( new_n932_, new_n918_, new_n402_ );
and g0795 ( new_n933_, new_n932_, N25 );
and g0796 ( new_n934_, new_n923_, new_n472_ );
and g0797 ( new_n935_, new_n934_, new_n371_ );
or g0798 ( N730, new_n933_, new_n935_ );
or g0799 ( new_n937_, new_n918_, new_n324_ );
and g0800 ( new_n938_, new_n937_, N29 );
and g0801 ( new_n939_, new_n923_, new_n480_ );
and g0802 ( new_n940_, new_n939_, new_n291_ );
or g0803 ( N731, new_n938_, new_n940_ );
not g0804 ( new_n942_, keyIn_0_58 );
or g0805 ( new_n943_, new_n813_, new_n810_ );
or g0806 ( new_n944_, new_n808_, keyIn_0_43 );
and g0807 ( new_n945_, new_n944_, new_n943_ );
or g0808 ( new_n946_, new_n867_, keyIn_0_42 );
not g0809 ( new_n947_, new_n868_ );
and g0810 ( new_n948_, new_n947_, new_n946_ );
and g0811 ( new_n949_, new_n948_, new_n945_ );
and g0812 ( new_n950_, new_n949_, new_n761_ );
not g0813 ( new_n951_, new_n950_ );
or g0814 ( new_n952_, new_n526_, new_n951_ );
or g0815 ( new_n953_, new_n952_, new_n942_ );
and g0816 ( new_n954_, new_n877_, new_n950_ );
or g0817 ( new_n955_, new_n954_, keyIn_0_58 );
and g0818 ( new_n956_, new_n953_, new_n955_ );
or g0819 ( new_n957_, new_n956_, new_n249_ );
and g0820 ( new_n958_, new_n957_, N33 );
and g0821 ( new_n959_, new_n954_, keyIn_0_58 );
and g0822 ( new_n960_, new_n952_, new_n942_ );
or g0823 ( new_n961_, new_n960_, new_n959_ );
and g0824 ( new_n962_, new_n961_, new_n469_ );
and g0825 ( new_n963_, new_n962_, new_n223_ );
or g0826 ( N732, new_n958_, new_n963_ );
or g0827 ( new_n965_, new_n956_, new_n481_ );
and g0828 ( new_n966_, new_n965_, N37 );
and g0829 ( new_n967_, new_n961_, new_n460_ );
and g0830 ( new_n968_, new_n967_, new_n427_ );
or g0831 ( N733, new_n966_, new_n968_ );
or g0832 ( new_n970_, new_n956_, new_n402_ );
and g0833 ( new_n971_, new_n970_, N41 );
and g0834 ( new_n972_, new_n961_, new_n472_ );
and g0835 ( new_n973_, new_n972_, new_n375_ );
or g0836 ( N734, new_n971_, new_n973_ );
or g0837 ( new_n975_, new_n956_, new_n324_ );
and g0838 ( new_n976_, new_n975_, N45 );
and g0839 ( new_n977_, new_n961_, new_n480_ );
and g0840 ( new_n978_, new_n977_, new_n296_ );
or g0841 ( N735, new_n976_, new_n978_ );
not g0842 ( new_n980_, keyIn_0_59 );
and g0843 ( new_n981_, new_n910_, new_n907_ );
and g0844 ( new_n982_, new_n981_, new_n949_ );
not g0845 ( new_n983_, new_n982_ );
or g0846 ( new_n984_, new_n526_, new_n983_ );
or g0847 ( new_n985_, new_n984_, new_n980_ );
and g0848 ( new_n986_, new_n877_, new_n982_ );
or g0849 ( new_n987_, new_n986_, keyIn_0_59 );
and g0850 ( new_n988_, new_n985_, new_n987_ );
or g0851 ( new_n989_, new_n988_, new_n249_ );
and g0852 ( new_n990_, new_n989_, N49 );
and g0853 ( new_n991_, new_n986_, keyIn_0_59 );
and g0854 ( new_n992_, new_n984_, new_n980_ );
or g0855 ( new_n993_, new_n992_, new_n991_ );
and g0856 ( new_n994_, new_n993_, new_n469_ );
and g0857 ( new_n995_, new_n994_, new_n224_ );
or g0858 ( N736, new_n990_, new_n995_ );
or g0859 ( new_n997_, new_n988_, new_n481_ );
and g0860 ( new_n998_, new_n997_, N53 );
and g0861 ( new_n999_, new_n993_, new_n460_ );
and g0862 ( new_n1000_, new_n999_, new_n428_ );
or g0863 ( N737, new_n998_, new_n1000_ );
or g0864 ( new_n1002_, new_n988_, new_n402_ );
and g0865 ( new_n1003_, new_n1002_, N57 );
and g0866 ( new_n1004_, new_n993_, new_n472_ );
and g0867 ( new_n1005_, new_n1004_, new_n376_ );
or g0868 ( N738, new_n1003_, new_n1005_ );
or g0869 ( new_n1007_, new_n988_, new_n324_ );
and g0870 ( new_n1008_, new_n1007_, N61 );
and g0871 ( new_n1009_, new_n993_, new_n480_ );
and g0872 ( new_n1010_, new_n1009_, new_n297_ );
or g0873 ( N739, new_n1008_, new_n1010_ );
not g0874 ( new_n1012_, keyIn_0_60 );
not g0875 ( new_n1013_, keyIn_0_55 );
not g0876 ( new_n1014_, keyIn_0_53 );
and g0877 ( new_n1015_, new_n911_, new_n760_ );
and g0878 ( new_n1016_, new_n1015_, new_n1014_ );
not g0879 ( new_n1017_, new_n1016_ );
or g0880 ( new_n1018_, new_n1015_, new_n1014_ );
and g0881 ( new_n1019_, new_n1017_, new_n1018_ );
not g0882 ( new_n1020_, keyIn_0_51 );
and g0883 ( new_n1021_, new_n948_, new_n815_ );
and g0884 ( new_n1022_, new_n1021_, new_n761_ );
and g0885 ( new_n1023_, new_n1022_, new_n1020_ );
not g0886 ( new_n1024_, new_n1023_ );
or g0887 ( new_n1025_, new_n1022_, new_n1020_ );
and g0888 ( new_n1026_, new_n1024_, new_n1025_ );
not g0889 ( new_n1027_, keyIn_0_52 );
or g0890 ( new_n1028_, new_n815_, new_n869_ );
or g0891 ( new_n1029_, new_n907_, new_n636_ );
or g0892 ( new_n1030_, new_n1029_, new_n1028_ );
or g0893 ( new_n1031_, new_n1030_, new_n1027_ );
and g0894 ( new_n1032_, new_n910_, new_n760_ );
and g0895 ( new_n1033_, new_n1032_, new_n949_ );
or g0896 ( new_n1034_, new_n1033_, keyIn_0_52 );
and g0897 ( new_n1035_, new_n1031_, new_n1034_ );
not g0898 ( new_n1036_, keyIn_0_50 );
or g0899 ( new_n1037_, new_n760_, new_n636_ );
or g0900 ( new_n1038_, new_n945_, new_n869_ );
or g0901 ( new_n1039_, new_n1037_, new_n1038_ );
or g0902 ( new_n1040_, new_n1039_, new_n1036_ );
and g0903 ( new_n1041_, new_n981_, new_n1021_ );
or g0904 ( new_n1042_, new_n1041_, keyIn_0_50 );
and g0905 ( new_n1043_, new_n1040_, new_n1042_ );
or g0906 ( new_n1044_, new_n1035_, new_n1043_ );
or g0907 ( new_n1045_, new_n1044_, new_n1026_ );
or g0908 ( new_n1046_, new_n1045_, new_n1019_ );
and g0909 ( new_n1047_, new_n1046_, new_n1013_ );
not g0910 ( new_n1048_, new_n1019_ );
not g0911 ( new_n1049_, new_n1026_ );
and g0912 ( new_n1050_, new_n1033_, keyIn_0_52 );
and g0913 ( new_n1051_, new_n1030_, new_n1027_ );
or g0914 ( new_n1052_, new_n1051_, new_n1050_ );
and g0915 ( new_n1053_, new_n1041_, keyIn_0_50 );
and g0916 ( new_n1054_, new_n1039_, new_n1036_ );
or g0917 ( new_n1055_, new_n1054_, new_n1053_ );
and g0918 ( new_n1056_, new_n1052_, new_n1055_ );
and g0919 ( new_n1057_, new_n1056_, new_n1049_ );
and g0920 ( new_n1058_, new_n1057_, new_n1048_ );
and g0921 ( new_n1059_, new_n1058_, keyIn_0_55 );
or g0922 ( new_n1060_, new_n1047_, new_n1059_ );
and g0923 ( new_n1061_, new_n501_, new_n486_ );
and g0924 ( new_n1062_, new_n1060_, new_n1061_ );
or g0925 ( new_n1063_, new_n1062_, new_n1012_ );
or g0926 ( new_n1064_, new_n1058_, keyIn_0_55 );
not g0927 ( new_n1065_, new_n1059_ );
and g0928 ( new_n1066_, new_n1065_, new_n1064_ );
not g0929 ( new_n1067_, new_n1061_ );
or g0930 ( new_n1068_, new_n1066_, new_n1067_ );
or g0931 ( new_n1069_, new_n1068_, keyIn_0_60 );
and g0932 ( new_n1070_, new_n1069_, new_n1063_ );
or g0933 ( new_n1071_, new_n1070_, new_n948_ );
and g0934 ( new_n1072_, new_n1071_, N65 );
and g0935 ( new_n1073_, new_n1068_, keyIn_0_60 );
and g0936 ( new_n1074_, new_n1062_, new_n1012_ );
or g0937 ( new_n1075_, new_n1073_, new_n1074_ );
and g0938 ( new_n1076_, new_n1075_, new_n869_ );
and g0939 ( new_n1077_, new_n1076_, new_n141_ );
or g0940 ( N740, new_n1072_, new_n1077_ );
or g0941 ( new_n1079_, new_n1070_, new_n815_ );
and g0942 ( new_n1080_, new_n1079_, N69 );
and g0943 ( new_n1081_, new_n1075_, new_n945_ );
and g0944 ( new_n1082_, new_n1081_, new_n142_ );
or g0945 ( N741, new_n1080_, new_n1082_ );
or g0946 ( new_n1084_, new_n1070_, new_n910_ );
and g0947 ( new_n1085_, new_n1084_, N73 );
and g0948 ( new_n1086_, new_n1075_, new_n636_ );
and g0949 ( new_n1087_, new_n1086_, new_n148_ );
or g0950 ( N742, new_n1085_, new_n1087_ );
or g0951 ( new_n1089_, new_n1070_, new_n760_ );
and g0952 ( new_n1090_, new_n1089_, N77 );
and g0953 ( new_n1091_, new_n1075_, new_n907_ );
and g0954 ( new_n1092_, new_n1091_, new_n146_ );
or g0955 ( N743, new_n1090_, new_n1092_ );
not g0956 ( new_n1094_, keyIn_0_61 );
and g0957 ( new_n1095_, new_n502_, new_n480_ );
and g0958 ( new_n1096_, new_n1060_, new_n1095_ );
or g0959 ( new_n1097_, new_n1096_, new_n1094_ );
not g0960 ( new_n1098_, new_n1095_ );
or g0961 ( new_n1099_, new_n1066_, new_n1098_ );
or g0962 ( new_n1100_, new_n1099_, keyIn_0_61 );
and g0963 ( new_n1101_, new_n1100_, new_n1097_ );
or g0964 ( new_n1102_, new_n1101_, new_n948_ );
and g0965 ( new_n1103_, new_n1102_, N81 );
and g0966 ( new_n1104_, new_n1099_, keyIn_0_61 );
and g0967 ( new_n1105_, new_n1096_, new_n1094_ );
or g0968 ( new_n1106_, new_n1104_, new_n1105_ );
and g0969 ( new_n1107_, new_n1106_, new_n869_ );
and g0970 ( new_n1108_, new_n1107_, new_n173_ );
or g0971 ( N744, new_n1103_, new_n1108_ );
or g0972 ( new_n1110_, new_n1101_, new_n815_ );
and g0973 ( new_n1111_, new_n1110_, N85 );
and g0974 ( new_n1112_, new_n1106_, new_n945_ );
and g0975 ( new_n1113_, new_n1112_, new_n174_ );
or g0976 ( N745, new_n1111_, new_n1113_ );
or g0977 ( new_n1115_, new_n1101_, new_n910_ );
and g0978 ( new_n1116_, new_n1115_, N89 );
and g0979 ( new_n1117_, new_n1106_, new_n636_ );
and g0980 ( new_n1118_, new_n1117_, new_n178_ );
or g0981 ( N746, new_n1116_, new_n1118_ );
or g0982 ( new_n1120_, new_n1101_, new_n760_ );
and g0983 ( new_n1121_, new_n1120_, N93 );
and g0984 ( new_n1122_, new_n1106_, new_n907_ );
and g0985 ( new_n1123_, new_n1122_, new_n179_ );
or g0986 ( N747, new_n1121_, new_n1123_ );
not g0987 ( new_n1125_, keyIn_0_62 );
and g0988 ( new_n1126_, new_n487_, new_n460_ );
and g0989 ( new_n1127_, new_n1060_, new_n1126_ );
or g0990 ( new_n1128_, new_n1127_, new_n1125_ );
not g0991 ( new_n1129_, new_n1126_ );
or g0992 ( new_n1130_, new_n1066_, new_n1129_ );
or g0993 ( new_n1131_, new_n1130_, keyIn_0_62 );
and g0994 ( new_n1132_, new_n1131_, new_n1128_ );
or g0995 ( new_n1133_, new_n1132_, new_n948_ );
and g0996 ( new_n1134_, new_n1133_, N97 );
and g0997 ( new_n1135_, new_n1130_, keyIn_0_62 );
and g0998 ( new_n1136_, new_n1127_, new_n1125_ );
or g0999 ( new_n1137_, new_n1135_, new_n1136_ );
and g1000 ( new_n1138_, new_n1137_, new_n869_ );
and g1001 ( new_n1139_, new_n1138_, new_n329_ );
or g1002 ( N748, new_n1134_, new_n1139_ );
or g1003 ( new_n1141_, new_n1132_, new_n815_ );
and g1004 ( new_n1142_, new_n1141_, N101 );
and g1005 ( new_n1143_, new_n1137_, new_n945_ );
and g1006 ( new_n1144_, new_n1143_, new_n327_ );
or g1007 ( N749, new_n1142_, new_n1144_ );
or g1008 ( new_n1146_, new_n1132_, new_n910_ );
and g1009 ( new_n1147_, new_n1146_, N105 );
and g1010 ( new_n1148_, new_n1137_, new_n636_ );
and g1011 ( new_n1149_, new_n1148_, new_n332_ );
or g1012 ( N750, new_n1147_, new_n1149_ );
or g1013 ( new_n1151_, new_n1132_, new_n760_ );
and g1014 ( new_n1152_, new_n1151_, N109 );
and g1015 ( new_n1153_, new_n1137_, new_n907_ );
and g1016 ( new_n1154_, new_n1153_, new_n333_ );
or g1017 ( N751, new_n1152_, new_n1154_ );
not g1018 ( new_n1156_, keyIn_0_63 );
and g1019 ( new_n1157_, new_n461_, new_n480_ );
and g1020 ( new_n1158_, new_n1060_, new_n1157_ );
or g1021 ( new_n1159_, new_n1158_, new_n1156_ );
not g1022 ( new_n1160_, new_n1157_ );
or g1023 ( new_n1161_, new_n1066_, new_n1160_ );
or g1024 ( new_n1162_, new_n1161_, keyIn_0_63 );
and g1025 ( new_n1163_, new_n1162_, new_n1159_ );
or g1026 ( new_n1164_, new_n1163_, new_n948_ );
and g1027 ( new_n1165_, new_n1164_, N113 );
and g1028 ( new_n1166_, new_n1161_, keyIn_0_63 );
and g1029 ( new_n1167_, new_n1158_, new_n1156_ );
or g1030 ( new_n1168_, new_n1166_, new_n1167_ );
and g1031 ( new_n1169_, new_n1168_, new_n869_ );
and g1032 ( new_n1170_, new_n1169_, new_n258_ );
or g1033 ( N752, new_n1165_, new_n1170_ );
or g1034 ( new_n1172_, new_n1163_, new_n815_ );
and g1035 ( new_n1173_, new_n1172_, N117 );
and g1036 ( new_n1174_, new_n1168_, new_n945_ );
and g1037 ( new_n1175_, new_n1174_, new_n256_ );
or g1038 ( N753, new_n1173_, new_n1175_ );
or g1039 ( new_n1177_, new_n1163_, new_n910_ );
and g1040 ( new_n1178_, new_n1177_, N121 );
and g1041 ( new_n1179_, new_n1168_, new_n636_ );
and g1042 ( new_n1180_, new_n1179_, new_n261_ );
or g1043 ( N754, new_n1178_, new_n1180_ );
or g1044 ( new_n1182_, new_n1163_, new_n760_ );
and g1045 ( new_n1183_, new_n1182_, N125 );
and g1046 ( new_n1184_, new_n1168_, new_n907_ );
and g1047 ( new_n1185_, new_n1184_, new_n262_ );
or g1048 ( N755, new_n1183_, new_n1185_ );
endmodule