module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n479_, new_n1105_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n798_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1025_, new_n566_, new_n641_, new_n365_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n840_, new_n735_, new_n1045_, new_n500_, new_n898_, new_n786_, new_n799_, new_n946_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n626_, new_n959_, new_n990_, new_n774_, new_n716_, new_n701_, new_n792_, new_n1058_, new_n953_, new_n481_, new_n1073_, new_n1110_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n350_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n1083_, new_n385_, new_n1049_, new_n829_, new_n988_, new_n478_, new_n694_, new_n461_, new_n710_, new_n971_, new_n565_, new_n764_, new_n906_, new_n683_, new_n511_, new_n463_, new_n510_, new_n966_, new_n351_, new_n517_, new_n609_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1006_, new_n622_, new_n629_, new_n702_, new_n833_, new_n883_, new_n1005_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n650_, new_n708_, new_n750_, new_n887_, new_n429_, new_n926_, new_n353_, new_n432_, new_n734_, new_n912_, new_n925_, new_n1062_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n778_, new_n452_, new_n381_, new_n920_, new_n656_, new_n820_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n394_, new_n1007_, new_n935_, new_n882_, new_n657_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1020_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n398_, new_n646_, new_n395_, new_n538_, new_n383_, new_n854_, new_n541_, new_n458_, new_n1026_, new_n447_, new_n1106_, new_n473_, new_n790_, new_n1081_, new_n587_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n874_, new_n402_, new_n663_, new_n579_, new_n659_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n528_, new_n952_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n399_, new_n596_, new_n870_, new_n945_, new_n805_, new_n559_, new_n948_, new_n762_, new_n1055_, new_n838_, new_n923_, new_n469_, new_n391_, new_n437_, new_n1085_, new_n359_, new_n794_, new_n628_, new_n409_, new_n1090_, new_n457_, new_n553_, new_n1084_, new_n1061_, new_n668_, new_n1002_, new_n834_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n688_, new_n384_, new_n900_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n371_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1000_, new_n633_, new_n797_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n362_, new_n809_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n693_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n376_, new_n380_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n998_, new_n1056_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n562_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n379_, new_n1012_, new_n719_, new_n869_, new_n963_, new_n586_, new_n570_, new_n598_, new_n893_, new_n993_, new_n1063_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n825_, new_n858_, new_n557_, new_n936_, new_n411_, new_n507_, new_n673_, new_n741_, new_n806_, new_n605_, new_n1016_, new_n1074_, new_n748_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n558_, new_n382_, new_n583_, new_n617_, new_n1080_, new_n718_, new_n522_, new_n588_, new_n781_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n546_, new_n919_, new_n1015_, new_n755_, new_n1040_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n499_, new_n533_, new_n1088_, new_n795_, new_n459_, new_n569_, new_n555_, new_n977_, new_n782_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n751_, new_n535_, new_n1038_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n597_, new_n1093_, new_n1092_, new_n408_, new_n470_, new_n1072_, new_n769_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n989_, new_n1112_, new_n711_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n973_, new_n412_, new_n607_, new_n904_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1008_, new_n640_, new_n684_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n905_, new_n539_, new_n803_, new_n727_, new_n962_, new_n760_, new_n627_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n780_, new_n984_, new_n643_, new_n474_, new_n467_, new_n1013_, new_n404_, new_n1077_, new_n490_, new_n560_, new_n1100_, new_n865_, new_n1027_, new_n877_, new_n348_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n425_, new_n896_, new_n802_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n709_, new_n373_, new_n866_, new_n540_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n521_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n647_, new_n889_, new_n536_, new_n464_, new_n1089_, new_n573_, new_n765_, new_n405_, new_n1103_;

and g000 ( N388, N29, N42, N75 );
and g001 ( N389, N29, N36, N80 );
nand g002 ( new_n345_, N29, N36, N42 );
not g003 ( N390, new_n345_ );
and g004 ( N391, N85, N86 );
not g005 ( new_n348_, N1 );
not g006 ( new_n349_, N8 );
not g007 ( new_n350_, N13 );
not g008 ( new_n351_, N17 );
nor g009 ( N418, new_n348_, new_n349_, new_n350_, new_n351_ );
nand g010 ( new_n353_, N1, N13, N17, N26 );
nor g011 ( new_n354_, N390, new_n353_ );
xor g012 ( N419, new_n354_, keyIn_0_8 );
nand g013 ( N420, N59, N75, N80 );
nand g014 ( N421, N36, N59, N80 );
nand g015 ( N422, N36, N42, N59 );
not g016 ( new_n359_, N90 );
nor g017 ( new_n360_, N87, N88 );
nor g018 ( N423, new_n360_, new_n359_ );
nor g019 ( new_n362_, new_n353_, new_n345_ );
xor g020 ( N446, new_n362_, keyIn_0_25 );
not g021 ( new_n364_, keyIn_0_0 );
nand g022 ( new_n365_, N1, N26, N51 );
nand g023 ( new_n366_, new_n365_, new_n364_ );
nand g024 ( new_n367_, keyIn_0_0, N1, N26, N51 );
nand g025 ( N447, new_n366_, new_n367_ );
not g026 ( new_n369_, N55 );
nor g027 ( new_n370_, new_n348_, new_n349_, new_n350_, new_n369_ );
nand g028 ( new_n371_, new_n370_, N29, N68 );
xnor g029 ( N448, new_n371_, keyIn_0_12 );
and g030 ( new_n373_, N59, N68 );
nand g031 ( new_n374_, new_n370_, N74, new_n373_ );
xnor g032 ( N449, new_n374_, keyIn_0_13 );
not g033 ( new_n376_, N89 );
nor g034 ( N450, new_n360_, new_n376_ );
xor g035 ( new_n378_, N111, N116 );
xnor g036 ( new_n379_, new_n378_, keyIn_0_17 );
xor g037 ( new_n380_, new_n379_, keyIn_0_31 );
xnor g038 ( new_n381_, N121, N126 );
xnor g039 ( new_n382_, new_n381_, keyIn_0_18 );
xor g040 ( new_n383_, new_n382_, keyIn_0_32 );
nand g041 ( new_n384_, new_n380_, new_n383_ );
xor g042 ( new_n385_, new_n384_, keyIn_0_43 );
nand g043 ( new_n386_, new_n379_, new_n382_ );
xor g044 ( new_n387_, new_n386_, keyIn_0_33 );
nand g045 ( new_n388_, new_n385_, new_n387_ );
xor g046 ( new_n389_, new_n388_, keyIn_0_53 );
nor g047 ( new_n390_, new_n389_, N135 );
xor g048 ( new_n391_, new_n390_, keyIn_0_73 );
nand g049 ( new_n392_, new_n389_, N135 );
xnor g050 ( new_n393_, new_n392_, keyIn_0_72 );
nand g051 ( new_n394_, new_n391_, new_n393_ );
xor g052 ( new_n395_, new_n394_, keyIn_0_95 );
xor g053 ( new_n396_, N101, N106 );
xnor g054 ( new_n397_, new_n396_, keyIn_0_16 );
xor g055 ( new_n398_, new_n397_, keyIn_0_29 );
xnor g056 ( new_n399_, N91, N96 );
xnor g057 ( new_n400_, new_n399_, keyIn_0_15 );
xor g058 ( new_n401_, new_n400_, keyIn_0_28 );
nand g059 ( new_n402_, new_n398_, new_n401_ );
nand g060 ( new_n403_, new_n402_, keyIn_0_42 );
or g061 ( new_n404_, new_n402_, keyIn_0_42 );
nand g062 ( new_n405_, new_n397_, new_n400_ );
xnor g063 ( new_n406_, new_n405_, keyIn_0_30 );
nand g064 ( new_n407_, new_n404_, new_n403_, new_n406_ );
xnor g065 ( new_n408_, new_n407_, keyIn_0_52 );
nor g066 ( new_n409_, new_n408_, N130 );
xor g067 ( new_n410_, new_n409_, keyIn_0_71 );
nand g068 ( new_n411_, new_n408_, N130 );
xor g069 ( new_n412_, new_n411_, keyIn_0_70 );
nand g070 ( new_n413_, new_n410_, new_n412_ );
xnor g071 ( new_n414_, new_n413_, keyIn_0_94 );
nor g072 ( new_n415_, new_n395_, new_n414_ );
xor g073 ( new_n416_, new_n415_, keyIn_0_116 );
nand g074 ( new_n417_, new_n395_, new_n414_ );
xor g075 ( new_n418_, new_n417_, keyIn_0_106 );
nand g076 ( new_n419_, new_n416_, new_n418_ );
xnor g077 ( N767, new_n419_, keyIn_0_139 );
xor g078 ( new_n421_, N159, N165 );
xnor g079 ( new_n422_, new_n421_, keyIn_0_21 );
xor g080 ( new_n423_, new_n422_, keyIn_0_35 );
xnor g081 ( new_n424_, N171, N177 );
xnor g082 ( new_n425_, new_n424_, keyIn_0_22 );
xor g083 ( new_n426_, new_n425_, keyIn_0_36 );
nand g084 ( new_n427_, new_n423_, new_n426_ );
xnor g085 ( new_n428_, new_n427_, keyIn_0_49 );
nand g086 ( new_n429_, new_n422_, new_n425_ );
xor g087 ( new_n430_, new_n429_, keyIn_0_37 );
nand g088 ( new_n431_, new_n428_, new_n430_ );
xnor g089 ( new_n432_, new_n431_, keyIn_0_68 );
nor g090 ( new_n433_, new_n432_, N130 );
xor g091 ( new_n434_, new_n433_, keyIn_0_91 );
nand g092 ( new_n435_, new_n432_, N130 );
xnor g093 ( new_n436_, new_n435_, keyIn_0_90 );
nand g094 ( new_n437_, new_n434_, new_n436_ );
xnor g095 ( new_n438_, new_n437_, keyIn_0_104 );
not g096 ( new_n439_, N207 );
xnor g097 ( new_n440_, N183, N189 );
xor g098 ( new_n441_, new_n440_, keyIn_0_23 );
not g099 ( new_n442_, new_n441_ );
or g100 ( new_n443_, new_n442_, keyIn_0_38 );
xnor g101 ( new_n444_, N195, N201 );
xor g102 ( new_n445_, new_n444_, keyIn_0_24 );
not g103 ( new_n446_, new_n445_ );
or g104 ( new_n447_, new_n446_, keyIn_0_39 );
nand g105 ( new_n448_, new_n446_, keyIn_0_39 );
nand g106 ( new_n449_, new_n442_, keyIn_0_38 );
nand g107 ( new_n450_, new_n443_, new_n447_, new_n448_, new_n449_ );
nand g108 ( new_n451_, new_n450_, keyIn_0_50 );
or g109 ( new_n452_, new_n450_, keyIn_0_50 );
nand g110 ( new_n453_, new_n441_, new_n445_ );
xnor g111 ( new_n454_, new_n453_, keyIn_0_40 );
nand g112 ( new_n455_, new_n452_, new_n451_, new_n454_ );
xor g113 ( new_n456_, new_n455_, keyIn_0_69 );
nor g114 ( new_n457_, new_n456_, new_n439_ );
xor g115 ( new_n458_, new_n457_, keyIn_0_92 );
nand g116 ( new_n459_, new_n456_, new_n439_ );
xor g117 ( new_n460_, new_n459_, keyIn_0_93 );
nand g118 ( new_n461_, new_n458_, new_n460_ );
xor g119 ( new_n462_, new_n461_, keyIn_0_105 );
nor g120 ( new_n463_, new_n462_, new_n438_ );
xor g121 ( new_n464_, new_n463_, keyIn_0_117 );
nand g122 ( new_n465_, new_n462_, new_n438_ );
xnor g123 ( new_n466_, new_n465_, keyIn_0_115 );
nand g124 ( new_n467_, new_n464_, new_n466_ );
xnor g125 ( N768, new_n467_, keyIn_0_140 );
not g126 ( new_n469_, keyIn_0_210 );
not g127 ( new_n470_, keyIn_0_137 );
not g128 ( new_n471_, keyIn_0_114 );
not g129 ( new_n472_, keyIn_0_63 );
not g130 ( new_n473_, keyIn_0_48 );
not g131 ( new_n474_, keyIn_0_26 );
nand g132 ( new_n475_, N447, keyIn_0_9 );
not g133 ( new_n476_, keyIn_0_9 );
nand g134 ( new_n477_, new_n366_, new_n476_, new_n367_ );
nand g135 ( new_n478_, new_n475_, new_n477_ );
nand g136 ( new_n479_, new_n478_, new_n474_ );
nand g137 ( new_n480_, new_n475_, keyIn_0_26, new_n477_ );
nand g138 ( new_n481_, N59, N156 );
xnor g139 ( new_n482_, new_n481_, keyIn_0_5 );
and g140 ( new_n483_, new_n482_, N17 );
nand g141 ( new_n484_, new_n479_, new_n473_, new_n480_, new_n483_ );
nand g142 ( new_n485_, new_n479_, new_n480_, new_n483_ );
nand g143 ( new_n486_, new_n485_, keyIn_0_48 );
nand g144 ( new_n487_, new_n486_, new_n484_ );
nand g145 ( new_n488_, new_n487_, new_n472_, N1 );
nand g146 ( new_n489_, new_n487_, N1 );
nand g147 ( new_n490_, new_n489_, keyIn_0_63 );
nand g148 ( new_n491_, new_n490_, N153, new_n488_ );
xnor g149 ( new_n492_, new_n491_, keyIn_0_88 );
not g150 ( new_n493_, keyIn_0_89 );
not g151 ( new_n494_, keyIn_0_47 );
not g152 ( new_n495_, new_n481_ );
not g153 ( new_n496_, keyIn_0_7 );
nand g154 ( new_n497_, N17, N42 );
nand g155 ( new_n498_, new_n497_, new_n496_ );
nand g156 ( new_n499_, keyIn_0_7, N17, N42 );
nand g157 ( new_n500_, new_n498_, new_n499_ );
not g158 ( new_n501_, N42 );
nand g159 ( new_n502_, new_n351_, new_n501_, keyIn_0_6 );
not g160 ( new_n503_, keyIn_0_6 );
nand g161 ( new_n504_, new_n351_, new_n501_ );
nand g162 ( new_n505_, new_n504_, new_n503_ );
nand g163 ( new_n506_, new_n500_, new_n505_, keyIn_0_20, new_n502_ );
not g164 ( new_n507_, keyIn_0_20 );
nand g165 ( new_n508_, new_n500_, new_n502_, new_n505_ );
nand g166 ( new_n509_, new_n508_, new_n507_ );
and g167 ( new_n510_, new_n509_, new_n495_, new_n506_ );
nand g168 ( new_n511_, new_n510_, new_n494_, new_n479_, new_n480_ );
and g169 ( new_n512_, new_n509_, new_n495_ );
nand g170 ( new_n513_, new_n512_, new_n479_, new_n480_, new_n506_ );
nand g171 ( new_n514_, new_n513_, keyIn_0_47 );
not g172 ( new_n515_, keyIn_0_3 );
nand g173 ( new_n516_, N42, N59, N75 );
xnor g174 ( new_n517_, new_n516_, new_n515_ );
nand g175 ( new_n518_, new_n517_, keyIn_0_14 );
not g176 ( new_n519_, keyIn_0_14 );
xnor g177 ( new_n520_, new_n516_, keyIn_0_3 );
nand g178 ( new_n521_, new_n520_, new_n519_ );
nand g179 ( new_n522_, new_n518_, new_n521_ );
nor g180 ( new_n523_, new_n348_, new_n349_ );
xnor g181 ( new_n524_, keyIn_0_1, keyIn_0_10 );
nand g182 ( new_n525_, new_n524_, N17, N51, new_n523_ );
nand g183 ( new_n526_, new_n523_, N17, N51 );
not g184 ( new_n527_, new_n524_ );
nand g185 ( new_n528_, new_n527_, new_n526_ );
nand g186 ( new_n529_, new_n528_, new_n525_ );
nand g187 ( new_n530_, new_n522_, new_n529_ );
nand g188 ( new_n531_, new_n530_, keyIn_0_34 );
not g189 ( new_n532_, keyIn_0_34 );
nand g190 ( new_n533_, new_n522_, new_n532_, new_n529_ );
nand g191 ( new_n534_, new_n531_, new_n533_ );
nand g192 ( new_n535_, new_n514_, new_n534_, new_n511_, keyIn_0_54 );
not g193 ( new_n536_, keyIn_0_54 );
nand g194 ( new_n537_, new_n514_, new_n511_, new_n534_ );
nand g195 ( new_n538_, new_n537_, new_n536_ );
nand g196 ( new_n539_, new_n538_, new_n535_ );
nand g197 ( new_n540_, new_n539_, N126 );
nand g198 ( new_n541_, new_n540_, new_n493_ );
nand g199 ( new_n542_, new_n539_, keyIn_0_89, N126 );
nand g200 ( new_n543_, new_n541_, new_n542_ );
nand g201 ( new_n544_, new_n543_, new_n492_, keyIn_0_103 );
not g202 ( new_n545_, keyIn_0_103 );
nand g203 ( new_n546_, new_n543_, new_n492_ );
nand g204 ( new_n547_, new_n546_, new_n545_ );
not g205 ( new_n548_, keyIn_0_46 );
and g206 ( new_n549_, new_n479_, new_n480_ );
nand g207 ( new_n550_, N29, N75, N80 );
xor g208 ( new_n551_, new_n550_, keyIn_0_2 );
nand g209 ( new_n552_, new_n549_, new_n551_ );
nor g210 ( new_n553_, new_n552_, new_n369_ );
or g211 ( new_n554_, new_n553_, new_n548_ );
nand g212 ( new_n555_, new_n553_, new_n548_ );
xor g213 ( new_n556_, keyIn_0_4, N268 );
xor g214 ( new_n557_, new_n556_, keyIn_0_19 );
nand g215 ( new_n558_, new_n554_, new_n555_, new_n557_ );
xnor g216 ( new_n559_, new_n558_, keyIn_0_67 );
nand g217 ( new_n560_, new_n547_, new_n544_, new_n559_ );
nand g218 ( new_n561_, new_n560_, new_n471_ );
nand g219 ( new_n562_, new_n547_, keyIn_0_114, new_n544_, new_n559_ );
nand g220 ( new_n563_, new_n561_, new_n562_ );
nand g221 ( new_n564_, new_n563_, new_n470_, N201 );
nand g222 ( new_n565_, new_n563_, N201 );
nand g223 ( new_n566_, new_n565_, keyIn_0_137 );
nand g224 ( new_n567_, new_n566_, new_n564_ );
not g225 ( new_n568_, keyIn_0_138 );
not g226 ( new_n569_, N201 );
nand g227 ( new_n570_, new_n561_, new_n569_, new_n562_ );
nand g228 ( new_n571_, new_n570_, new_n568_ );
nand g229 ( new_n572_, new_n561_, keyIn_0_138, new_n569_, new_n562_ );
nand g230 ( new_n573_, new_n571_, new_n572_ );
nand g231 ( new_n574_, new_n567_, new_n573_ );
xor g232 ( new_n575_, new_n574_, keyIn_0_163 );
nor g233 ( new_n576_, new_n575_, N261 );
xor g234 ( new_n577_, new_n576_, keyIn_0_184 );
nand g235 ( new_n578_, new_n575_, N261 );
xor g236 ( new_n579_, new_n578_, keyIn_0_185 );
and g237 ( new_n580_, new_n577_, new_n579_ );
or g238 ( new_n581_, new_n580_, keyIn_0_202 );
nand g239 ( new_n582_, new_n580_, keyIn_0_202 );
nand g240 ( new_n583_, new_n581_, N219, new_n582_ );
nand g241 ( new_n584_, new_n583_, new_n469_ );
or g242 ( new_n585_, new_n583_, new_n469_ );
nand g243 ( new_n586_, N121, N210 );
nand g244 ( new_n587_, new_n585_, new_n584_, new_n586_ );
nand g245 ( new_n588_, new_n587_, keyIn_0_216 );
or g246 ( new_n589_, new_n587_, keyIn_0_216 );
nand g247 ( new_n590_, new_n575_, N228 );
not g248 ( new_n591_, keyIn_0_162 );
xnor g249 ( new_n592_, new_n567_, new_n591_ );
nand g250 ( new_n593_, new_n592_, N237 );
and g251 ( new_n594_, new_n590_, new_n593_ );
and g252 ( new_n595_, new_n594_, keyIn_0_203 );
nor g253 ( new_n596_, new_n594_, keyIn_0_203 );
nand g254 ( new_n597_, new_n563_, N246 );
nand g255 ( new_n598_, N255, N267 );
and g256 ( new_n599_, new_n597_, new_n598_ );
nand g257 ( new_n600_, new_n599_, keyIn_0_164 );
or g258 ( new_n601_, new_n599_, keyIn_0_164 );
nand g259 ( new_n602_, new_n370_, N42, N72, new_n373_ );
xor g260 ( new_n603_, new_n602_, keyIn_0_11 );
nand g261 ( new_n604_, new_n603_, N73 );
xor g262 ( new_n605_, new_n604_, keyIn_0_27 );
xnor g263 ( new_n606_, new_n605_, keyIn_0_41 );
xor g264 ( new_n607_, new_n606_, keyIn_0_51 );
nand g265 ( new_n608_, new_n607_, N201 );
nand g266 ( new_n609_, new_n601_, new_n600_, new_n608_ );
nor g267 ( new_n610_, new_n595_, new_n596_, new_n609_ );
nand g268 ( new_n611_, new_n589_, new_n588_, new_n610_ );
xnor g269 ( N850, new_n611_, keyIn_0_222 );
not g270 ( new_n613_, keyIn_0_196 );
not g271 ( new_n614_, N189 );
not g272 ( new_n615_, keyIn_0_112 );
not g273 ( new_n616_, keyIn_0_101 );
not g274 ( new_n617_, keyIn_0_84 );
nand g275 ( new_n618_, new_n490_, new_n617_, N146, new_n488_ );
nand g276 ( new_n619_, new_n490_, N146, new_n488_ );
nand g277 ( new_n620_, new_n619_, keyIn_0_84 );
nand g278 ( new_n621_, new_n620_, new_n618_ );
not g279 ( new_n622_, keyIn_0_85 );
nand g280 ( new_n623_, new_n539_, N116 );
nand g281 ( new_n624_, new_n623_, new_n622_ );
nand g282 ( new_n625_, new_n539_, keyIn_0_85, N116 );
nand g283 ( new_n626_, new_n624_, new_n625_ );
nand g284 ( new_n627_, new_n626_, new_n616_, new_n621_ );
nand g285 ( new_n628_, new_n626_, new_n621_ );
nand g286 ( new_n629_, new_n628_, keyIn_0_101 );
xnor g287 ( new_n630_, new_n558_, keyIn_0_65 );
nand g288 ( new_n631_, new_n629_, new_n615_, new_n627_, new_n630_ );
nand g289 ( new_n632_, new_n629_, new_n627_, new_n630_ );
nand g290 ( new_n633_, new_n632_, keyIn_0_112 );
nand g291 ( new_n634_, new_n633_, new_n631_ );
nand g292 ( new_n635_, new_n634_, new_n614_ );
xnor g293 ( new_n636_, new_n635_, keyIn_0_134 );
not g294 ( new_n637_, N195 );
not g295 ( new_n638_, keyIn_0_113 );
not g296 ( new_n639_, keyIn_0_86 );
nand g297 ( new_n640_, new_n490_, N149, new_n488_ );
xnor g298 ( new_n641_, new_n640_, new_n639_ );
not g299 ( new_n642_, keyIn_0_87 );
nand g300 ( new_n643_, new_n539_, N121 );
nand g301 ( new_n644_, new_n643_, new_n642_ );
nand g302 ( new_n645_, new_n539_, keyIn_0_87, N121 );
nand g303 ( new_n646_, new_n644_, new_n645_ );
nand g304 ( new_n647_, new_n646_, new_n641_, keyIn_0_102 );
not g305 ( new_n648_, keyIn_0_102 );
nand g306 ( new_n649_, new_n646_, new_n641_ );
nand g307 ( new_n650_, new_n649_, new_n648_ );
xnor g308 ( new_n651_, new_n558_, keyIn_0_66 );
nand g309 ( new_n652_, new_n650_, new_n638_, new_n647_, new_n651_ );
nand g310 ( new_n653_, new_n650_, new_n647_, new_n651_ );
nand g311 ( new_n654_, new_n653_, keyIn_0_113 );
nand g312 ( new_n655_, new_n654_, new_n652_ );
nand g313 ( new_n656_, new_n655_, new_n637_ );
xnor g314 ( new_n657_, new_n656_, keyIn_0_136 );
nand g315 ( new_n658_, new_n592_, new_n636_, new_n657_ );
nand g316 ( new_n659_, new_n658_, keyIn_0_188 );
not g317 ( new_n660_, keyIn_0_177 );
not g318 ( new_n661_, keyIn_0_156 );
not g319 ( new_n662_, keyIn_0_133 );
nand g320 ( new_n663_, new_n633_, new_n662_, N189, new_n631_ );
nand g321 ( new_n664_, new_n633_, N189, new_n631_ );
nand g322 ( new_n665_, new_n664_, keyIn_0_133 );
nand g323 ( new_n666_, new_n665_, new_n663_ );
nand g324 ( new_n667_, new_n666_, new_n661_ );
nand g325 ( new_n668_, new_n665_, keyIn_0_156, new_n663_ );
nand g326 ( new_n669_, new_n667_, new_n668_ );
xnor g327 ( new_n670_, new_n669_, new_n660_ );
not g328 ( new_n671_, keyIn_0_167 );
and g329 ( new_n672_, new_n573_, N261 );
nand g330 ( new_n673_, new_n672_, new_n657_, new_n636_, new_n671_ );
nand g331 ( new_n674_, new_n672_, new_n636_, new_n657_ );
nand g332 ( new_n675_, new_n674_, keyIn_0_167 );
and g333 ( new_n676_, new_n670_, new_n673_, new_n675_ );
not g334 ( new_n677_, keyIn_0_188 );
nand g335 ( new_n678_, new_n592_, new_n677_, new_n636_, new_n657_ );
not g336 ( new_n679_, keyIn_0_187 );
not g337 ( new_n680_, keyIn_0_159 );
not g338 ( new_n681_, keyIn_0_135 );
nand g339 ( new_n682_, new_n654_, new_n681_, N195, new_n652_ );
nand g340 ( new_n683_, new_n654_, N195, new_n652_ );
nand g341 ( new_n684_, new_n683_, keyIn_0_135 );
nand g342 ( new_n685_, new_n684_, new_n682_ );
nand g343 ( new_n686_, new_n685_, new_n680_ );
nand g344 ( new_n687_, new_n684_, keyIn_0_159, new_n682_ );
nand g345 ( new_n688_, new_n686_, new_n687_ );
nand g346 ( new_n689_, new_n688_, new_n636_ );
nand g347 ( new_n690_, new_n689_, new_n679_ );
nand g348 ( new_n691_, new_n688_, keyIn_0_187, new_n636_ );
nand g349 ( new_n692_, new_n690_, new_n691_ );
nand g350 ( new_n693_, new_n676_, new_n659_, new_n678_, new_n692_ );
nand g351 ( new_n694_, new_n693_, new_n613_ );
and g352 ( new_n695_, new_n692_, keyIn_0_196, new_n678_ );
nand g353 ( new_n696_, new_n695_, new_n659_, new_n676_ );
nand g354 ( new_n697_, new_n694_, new_n696_ );
nand g355 ( new_n698_, new_n539_, N111 );
xor g356 ( new_n699_, new_n698_, keyIn_0_83 );
nand g357 ( new_n700_, new_n490_, N143, new_n488_ );
xor g358 ( new_n701_, new_n700_, keyIn_0_82 );
nand g359 ( new_n702_, new_n699_, new_n701_ );
xor g360 ( new_n703_, new_n702_, keyIn_0_100 );
xnor g361 ( new_n704_, new_n558_, keyIn_0_64 );
nand g362 ( new_n705_, new_n703_, new_n704_ );
xnor g363 ( new_n706_, new_n705_, keyIn_0_111 );
nor g364 ( new_n707_, new_n706_, N183 );
xnor g365 ( new_n708_, new_n707_, keyIn_0_131 );
nand g366 ( new_n709_, new_n706_, N183 );
xnor g367 ( new_n710_, new_n709_, keyIn_0_130 );
nand g368 ( new_n711_, new_n708_, new_n710_ );
xnor g369 ( new_n712_, new_n711_, keyIn_0_154 );
nor g370 ( new_n713_, new_n697_, new_n712_ );
xnor g371 ( new_n714_, new_n713_, keyIn_0_205 );
nand g372 ( new_n715_, new_n697_, new_n712_ );
xnor g373 ( new_n716_, new_n715_, keyIn_0_204 );
nand g374 ( new_n717_, new_n714_, new_n716_ );
xnor g375 ( new_n718_, new_n717_, keyIn_0_213 );
and g376 ( new_n719_, new_n718_, N219 );
nand g377 ( new_n720_, new_n719_, keyIn_0_219 );
or g378 ( new_n721_, new_n719_, keyIn_0_219 );
nand g379 ( new_n722_, N106, N210 );
nand g380 ( new_n723_, new_n721_, new_n720_, new_n722_ );
or g381 ( new_n724_, new_n723_, keyIn_0_230 );
nand g382 ( new_n725_, new_n723_, keyIn_0_230 );
not g383 ( new_n726_, keyIn_0_197 );
not g384 ( new_n727_, new_n712_ );
and g385 ( new_n728_, new_n727_, N228 );
nand g386 ( new_n729_, new_n728_, keyIn_0_175 );
or g387 ( new_n730_, new_n728_, keyIn_0_175 );
xor g388 ( new_n731_, new_n710_, keyIn_0_153 );
nand g389 ( new_n732_, new_n731_, N237 );
xnor g390 ( new_n733_, new_n732_, keyIn_0_176 );
nand g391 ( new_n734_, new_n730_, new_n733_, new_n729_ );
nor g392 ( new_n735_, new_n734_, new_n726_ );
and g393 ( new_n736_, new_n734_, new_n726_ );
and g394 ( new_n737_, new_n706_, N246 );
nand g395 ( new_n738_, new_n737_, keyIn_0_132 );
or g396 ( new_n739_, new_n737_, keyIn_0_132 );
nand g397 ( new_n740_, new_n607_, N183 );
nand g398 ( new_n741_, new_n739_, new_n738_, new_n740_ );
xnor g399 ( new_n742_, new_n741_, keyIn_0_155 );
nor g400 ( new_n743_, new_n736_, new_n735_, new_n742_ );
nand g401 ( new_n744_, new_n724_, new_n725_, new_n743_ );
xor g402 ( N863, new_n744_, keyIn_0_240 );
xor g403 ( new_n746_, new_n688_, keyIn_0_180 );
nand g404 ( new_n747_, new_n672_, new_n657_ );
xor g405 ( new_n748_, new_n747_, keyIn_0_166 );
nand g406 ( new_n749_, new_n592_, new_n657_ );
xor g407 ( new_n750_, new_n749_, keyIn_0_186 );
nand g408 ( new_n751_, new_n750_, new_n746_, new_n748_ );
xor g409 ( new_n752_, new_n751_, keyIn_0_198 );
nand g410 ( new_n753_, new_n636_, new_n663_, new_n665_ );
xnor g411 ( new_n754_, new_n753_, keyIn_0_157 );
nor g412 ( new_n755_, new_n752_, new_n754_ );
xnor g413 ( new_n756_, new_n755_, keyIn_0_206 );
nand g414 ( new_n757_, new_n752_, new_n754_ );
xnor g415 ( new_n758_, new_n757_, keyIn_0_207 );
nand g416 ( new_n759_, new_n756_, new_n758_ );
xor g417 ( new_n760_, new_n759_, keyIn_0_214 );
and g418 ( new_n761_, new_n760_, N219 );
nand g419 ( new_n762_, new_n761_, keyIn_0_220 );
or g420 ( new_n763_, new_n761_, keyIn_0_220 );
nand g421 ( new_n764_, N111, N210 );
nand g422 ( new_n765_, new_n763_, new_n762_, new_n764_ );
nand g423 ( new_n766_, new_n765_, keyIn_0_231 );
or g424 ( new_n767_, new_n765_, keyIn_0_231 );
nand g425 ( new_n768_, new_n754_, N228 );
xor g426 ( new_n769_, new_n768_, keyIn_0_178 );
nand g427 ( new_n770_, new_n669_, N237 );
xor g428 ( new_n771_, new_n770_, keyIn_0_179 );
and g429 ( new_n772_, new_n769_, new_n771_ );
and g430 ( new_n773_, new_n772_, keyIn_0_199 );
nor g431 ( new_n774_, new_n772_, keyIn_0_199 );
nand g432 ( new_n775_, new_n633_, N246, new_n631_ );
nand g433 ( new_n776_, N255, N259 );
nand g434 ( new_n777_, new_n775_, new_n776_ );
nor g435 ( new_n778_, new_n777_, keyIn_0_158 );
and g436 ( new_n779_, new_n777_, keyIn_0_158 );
and g437 ( new_n780_, new_n607_, N189 );
or g438 ( new_n781_, new_n779_, new_n778_, new_n780_ );
nor g439 ( new_n782_, new_n773_, new_n774_, new_n781_ );
nand g440 ( new_n783_, new_n767_, new_n766_, new_n782_ );
xor g441 ( N864, new_n783_, keyIn_0_241 );
xnor g442 ( new_n785_, new_n592_, keyIn_0_183 );
xor g443 ( new_n786_, new_n672_, keyIn_0_165 );
nand g444 ( new_n787_, new_n785_, new_n786_ );
xnor g445 ( new_n788_, new_n787_, keyIn_0_200 );
nand g446 ( new_n789_, new_n657_, new_n685_ );
xor g447 ( new_n790_, new_n789_, keyIn_0_160 );
not g448 ( new_n791_, new_n790_ );
nand g449 ( new_n792_, new_n788_, new_n791_ );
xor g450 ( new_n793_, new_n792_, keyIn_0_208 );
nor g451 ( new_n794_, new_n788_, new_n791_ );
xnor g452 ( new_n795_, new_n794_, keyIn_0_209 );
and g453 ( new_n796_, new_n793_, new_n795_ );
or g454 ( new_n797_, new_n796_, keyIn_0_215 );
nand g455 ( new_n798_, new_n796_, keyIn_0_215 );
nand g456 ( new_n799_, new_n797_, N219, new_n798_ );
nand g457 ( new_n800_, new_n799_, keyIn_0_221 );
or g458 ( new_n801_, new_n799_, keyIn_0_221 );
nand g459 ( new_n802_, N116, N210 );
nand g460 ( new_n803_, new_n801_, new_n800_, new_n802_ );
xnor g461 ( new_n804_, new_n803_, keyIn_0_232 );
nand g462 ( new_n805_, new_n790_, N228 );
xor g463 ( new_n806_, new_n805_, keyIn_0_181 );
nand g464 ( new_n807_, new_n688_, N237 );
xor g465 ( new_n808_, new_n807_, keyIn_0_182 );
and g466 ( new_n809_, new_n806_, new_n808_ );
nand g467 ( new_n810_, new_n809_, keyIn_0_201 );
nor g468 ( new_n811_, new_n809_, keyIn_0_201 );
nand g469 ( new_n812_, new_n654_, N246, new_n652_ );
nand g470 ( new_n813_, N255, N260 );
nand g471 ( new_n814_, new_n812_, new_n813_ );
xnor g472 ( new_n815_, new_n814_, keyIn_0_161 );
and g473 ( new_n816_, new_n607_, N195 );
nor g474 ( new_n817_, new_n811_, new_n815_, new_n816_ );
nand g475 ( new_n818_, new_n804_, new_n810_, new_n817_ );
xor g476 ( N865, new_n818_, keyIn_0_242 );
not g477 ( new_n820_, keyIn_0_226 );
not g478 ( new_n821_, keyIn_0_99 );
nand g479 ( new_n822_, new_n539_, N106 );
nand g480 ( new_n823_, new_n822_, keyIn_0_80 );
or g481 ( new_n824_, new_n822_, keyIn_0_80 );
nand g482 ( new_n825_, N138, N152 );
nand g483 ( new_n826_, new_n824_, new_n823_, new_n825_ );
nand g484 ( new_n827_, new_n826_, new_n821_ );
nor g485 ( new_n828_, new_n552_, new_n351_ );
not g486 ( new_n829_, new_n828_ );
or g487 ( new_n830_, new_n829_, keyIn_0_45 );
nand g488 ( new_n831_, new_n829_, keyIn_0_45 );
nand g489 ( new_n832_, new_n830_, new_n556_, new_n831_ );
xor g490 ( new_n833_, new_n832_, keyIn_0_62 );
nand g491 ( new_n834_, new_n549_, N55, new_n482_ );
xor g492 ( new_n835_, new_n834_, keyIn_0_44 );
nand g493 ( new_n836_, new_n835_, N153 );
xnor g494 ( new_n837_, new_n836_, keyIn_0_61 );
nand g495 ( new_n838_, new_n833_, new_n837_ );
xnor g496 ( new_n839_, new_n838_, keyIn_0_81 );
or g497 ( new_n840_, new_n826_, new_n821_ );
nand g498 ( new_n841_, new_n839_, new_n827_, new_n840_ );
xnor g499 ( new_n842_, new_n841_, keyIn_0_110 );
nor g500 ( new_n843_, new_n842_, N177 );
xnor g501 ( new_n844_, new_n843_, keyIn_0_128 );
not g502 ( new_n845_, keyIn_0_212 );
nand g503 ( new_n846_, new_n669_, new_n660_ );
nand g504 ( new_n847_, new_n667_, keyIn_0_177, new_n668_ );
nand g505 ( new_n848_, new_n846_, new_n847_ );
and g506 ( new_n849_, new_n848_, new_n675_, new_n673_ );
nand g507 ( new_n850_, new_n849_, new_n659_, new_n678_, new_n692_ );
nand g508 ( new_n851_, new_n850_, new_n613_ );
nand g509 ( new_n852_, new_n695_, new_n659_, new_n849_ );
nand g510 ( new_n853_, new_n851_, new_n708_, new_n852_ );
nand g511 ( new_n854_, new_n853_, keyIn_0_211 );
not g512 ( new_n855_, keyIn_0_211 );
nand g513 ( new_n856_, new_n694_, new_n855_, new_n696_, new_n708_ );
nand g514 ( new_n857_, new_n854_, new_n856_ );
xor g515 ( new_n858_, new_n731_, keyIn_0_174 );
nand g516 ( new_n859_, new_n857_, new_n858_ );
nand g517 ( new_n860_, new_n859_, new_n845_ );
nand g518 ( new_n861_, new_n857_, keyIn_0_212, new_n858_ );
nand g519 ( new_n862_, new_n539_, N101 );
nand g520 ( new_n863_, new_n862_, keyIn_0_78 );
or g521 ( new_n864_, new_n862_, keyIn_0_78 );
nand g522 ( new_n865_, N17, N138 );
nand g523 ( new_n866_, new_n864_, new_n863_, new_n865_ );
xnor g524 ( new_n867_, new_n866_, keyIn_0_98 );
xor g525 ( new_n868_, new_n832_, keyIn_0_60 );
nand g526 ( new_n869_, new_n835_, N149 );
xnor g527 ( new_n870_, new_n869_, keyIn_0_59 );
nand g528 ( new_n871_, new_n868_, new_n870_ );
xor g529 ( new_n872_, new_n871_, keyIn_0_79 );
nand g530 ( new_n873_, new_n872_, new_n867_ );
xor g531 ( new_n874_, new_n873_, keyIn_0_109 );
nor g532 ( new_n875_, new_n874_, N171 );
xnor g533 ( new_n876_, new_n875_, keyIn_0_125 );
xor g534 ( new_n877_, new_n832_, keyIn_0_58 );
nand g535 ( new_n878_, new_n835_, N146 );
xor g536 ( new_n879_, new_n878_, keyIn_0_57 );
nand g537 ( new_n880_, new_n877_, new_n879_ );
xor g538 ( new_n881_, new_n880_, keyIn_0_77 );
nand g539 ( new_n882_, new_n539_, N96 );
nand g540 ( new_n883_, new_n882_, keyIn_0_76 );
or g541 ( new_n884_, new_n882_, keyIn_0_76 );
nand g542 ( new_n885_, N51, N138 );
nand g543 ( new_n886_, new_n884_, new_n883_, new_n885_ );
xor g544 ( new_n887_, new_n886_, keyIn_0_97 );
nand g545 ( new_n888_, new_n881_, new_n887_ );
xnor g546 ( new_n889_, new_n888_, keyIn_0_108 );
nor g547 ( new_n890_, new_n889_, N165 );
xor g548 ( new_n891_, new_n890_, keyIn_0_122 );
and g549 ( new_n892_, new_n876_, new_n891_ );
nand g550 ( new_n893_, new_n860_, new_n844_, new_n861_, new_n892_ );
nand g551 ( new_n894_, new_n893_, keyIn_0_225 );
not g552 ( new_n895_, keyIn_0_225 );
and g553 ( new_n896_, new_n860_, new_n861_ );
nand g554 ( new_n897_, new_n896_, new_n895_, new_n844_, new_n892_ );
nand g555 ( new_n898_, new_n842_, N177 );
xor g556 ( new_n899_, new_n898_, keyIn_0_127 );
xor g557 ( new_n900_, new_n899_, keyIn_0_150 );
and g558 ( new_n901_, new_n900_, new_n876_ );
nand g559 ( new_n902_, new_n901_, new_n891_ );
xnor g560 ( new_n903_, new_n902_, keyIn_0_191 );
nand g561 ( new_n904_, new_n874_, N171 );
xor g562 ( new_n905_, new_n904_, keyIn_0_124 );
xnor g563 ( new_n906_, new_n905_, keyIn_0_147 );
and g564 ( new_n907_, new_n906_, new_n891_ );
nand g565 ( new_n908_, new_n907_, keyIn_0_190 );
or g566 ( new_n909_, new_n907_, keyIn_0_190 );
nand g567 ( new_n910_, new_n889_, N165 );
xnor g568 ( new_n911_, new_n910_, keyIn_0_121 );
xor g569 ( new_n912_, new_n911_, keyIn_0_144 );
xor g570 ( new_n913_, new_n912_, keyIn_0_168 );
and g571 ( new_n914_, new_n903_, new_n908_, new_n909_, new_n913_ );
nand g572 ( new_n915_, new_n897_, new_n894_, new_n914_ );
nand g573 ( new_n916_, new_n915_, new_n820_ );
nand g574 ( new_n917_, new_n897_, keyIn_0_226, new_n894_, new_n914_ );
nand g575 ( new_n918_, new_n916_, new_n917_ );
nand g576 ( new_n919_, new_n539_, N91 );
nand g577 ( new_n920_, new_n919_, keyIn_0_74 );
or g578 ( new_n921_, new_n919_, keyIn_0_74 );
nand g579 ( new_n922_, N8, N138 );
nand g580 ( new_n923_, new_n921_, new_n920_, new_n922_ );
nand g581 ( new_n924_, new_n923_, keyIn_0_96 );
nand g582 ( new_n925_, new_n832_, keyIn_0_56 );
nand g583 ( new_n926_, new_n835_, N143 );
xor g584 ( new_n927_, new_n926_, keyIn_0_55 );
or g585 ( new_n928_, new_n832_, keyIn_0_56 );
nand g586 ( new_n929_, new_n927_, new_n925_, new_n928_ );
xor g587 ( new_n930_, new_n929_, keyIn_0_75 );
or g588 ( new_n931_, new_n923_, keyIn_0_96 );
nand g589 ( new_n932_, new_n930_, new_n924_, new_n931_ );
xnor g590 ( new_n933_, new_n932_, keyIn_0_107 );
nor g591 ( new_n934_, new_n933_, N159 );
xnor g592 ( new_n935_, new_n934_, keyIn_0_119 );
nand g593 ( new_n936_, new_n918_, new_n935_ );
or g594 ( new_n937_, new_n936_, keyIn_0_243 );
nand g595 ( new_n938_, new_n936_, keyIn_0_243 );
nand g596 ( new_n939_, new_n933_, N159 );
xnor g597 ( new_n940_, new_n939_, keyIn_0_118 );
xor g598 ( new_n941_, new_n940_, keyIn_0_141 );
nand g599 ( new_n942_, new_n937_, new_n938_, new_n941_ );
xor g600 ( N866, new_n942_, keyIn_0_248 );
not g601 ( new_n944_, keyIn_0_239 );
nand g602 ( new_n945_, new_n899_, new_n844_ );
xnor g603 ( new_n946_, new_n945_, keyIn_0_151 );
nand g604 ( new_n947_, new_n896_, new_n946_ );
xnor g605 ( new_n948_, new_n947_, keyIn_0_218 );
nor g606 ( new_n949_, new_n896_, new_n946_ );
xor g607 ( new_n950_, new_n949_, keyIn_0_217 );
nand g608 ( new_n951_, new_n950_, new_n948_ );
or g609 ( new_n952_, new_n951_, keyIn_0_229 );
nand g610 ( new_n953_, new_n951_, keyIn_0_229 );
nand g611 ( new_n954_, new_n952_, N219, new_n953_ );
nand g612 ( new_n955_, new_n954_, new_n944_ );
or g613 ( new_n956_, new_n954_, new_n944_ );
nand g614 ( new_n957_, N101, N210 );
nand g615 ( new_n958_, new_n956_, new_n955_, new_n957_ );
nand g616 ( new_n959_, new_n958_, keyIn_0_247 );
or g617 ( new_n960_, new_n958_, keyIn_0_247 );
nand g618 ( new_n961_, new_n946_, keyIn_0_172, N228 );
not g619 ( new_n962_, keyIn_0_172 );
nand g620 ( new_n963_, new_n946_, N228 );
nand g621 ( new_n964_, new_n963_, new_n962_ );
nand g622 ( new_n965_, new_n900_, N237 );
xor g623 ( new_n966_, new_n965_, keyIn_0_173 );
nand g624 ( new_n967_, new_n966_, new_n961_, new_n964_ );
nor g625 ( new_n968_, new_n967_, keyIn_0_195 );
and g626 ( new_n969_, new_n967_, keyIn_0_195 );
nand g627 ( new_n970_, new_n842_, N246 );
or g628 ( new_n971_, new_n970_, keyIn_0_129 );
nand g629 ( new_n972_, new_n970_, keyIn_0_129 );
nand g630 ( new_n973_, new_n607_, N177 );
nand g631 ( new_n974_, new_n971_, new_n972_, new_n973_ );
xor g632 ( new_n975_, new_n974_, keyIn_0_152 );
nor g633 ( new_n976_, new_n969_, new_n968_, new_n975_ );
nand g634 ( new_n977_, new_n960_, new_n959_, new_n976_ );
xnor g635 ( N874, new_n977_, keyIn_0_249 );
not g636 ( new_n979_, keyIn_0_253 );
not g637 ( new_n980_, keyIn_0_244 );
nand g638 ( new_n981_, new_n935_, new_n940_ );
xnor g639 ( new_n982_, new_n981_, keyIn_0_142 );
not g640 ( new_n983_, new_n982_ );
nand g641 ( new_n984_, new_n918_, new_n983_ );
xnor g642 ( new_n985_, new_n984_, keyIn_0_234 );
nand g643 ( new_n986_, new_n916_, new_n917_, new_n982_ );
xnor g644 ( new_n987_, new_n986_, keyIn_0_233 );
nand g645 ( new_n988_, new_n985_, new_n987_ );
nand g646 ( new_n989_, new_n988_, new_n980_ );
nand g647 ( new_n990_, new_n985_, keyIn_0_244, new_n987_ );
nand g648 ( new_n991_, new_n989_, N219, new_n990_ );
not g649 ( new_n992_, N210 );
or g650 ( new_n993_, new_n557_, new_n992_ );
nand g651 ( new_n994_, new_n991_, new_n993_ );
nand g652 ( new_n995_, new_n994_, keyIn_0_250 );
not g653 ( new_n996_, keyIn_0_250 );
nand g654 ( new_n997_, new_n991_, new_n996_, new_n993_ );
nand g655 ( new_n998_, new_n995_, new_n997_ );
nand g656 ( new_n999_, new_n983_, N228 );
not g657 ( new_n1000_, new_n941_ );
nand g658 ( new_n1001_, new_n1000_, N237 );
nand g659 ( new_n1002_, new_n999_, new_n1001_ );
nor g660 ( new_n1003_, new_n1002_, keyIn_0_192 );
and g661 ( new_n1004_, new_n1002_, keyIn_0_192 );
nand g662 ( new_n1005_, new_n933_, N246 );
xor g663 ( new_n1006_, new_n1005_, keyIn_0_120 );
nand g664 ( new_n1007_, new_n607_, N159 );
nand g665 ( new_n1008_, new_n1006_, new_n1007_ );
xnor g666 ( new_n1009_, new_n1008_, keyIn_0_143 );
nor g667 ( new_n1010_, new_n1004_, new_n1003_, new_n1009_ );
nand g668 ( new_n1011_, new_n998_, new_n979_, new_n1010_ );
nand g669 ( new_n1012_, new_n998_, new_n1010_ );
nand g670 ( new_n1013_, new_n1012_, keyIn_0_253 );
nand g671 ( N878, new_n1013_, new_n1011_ );
not g672 ( new_n1015_, keyIn_0_251 );
nand g673 ( new_n1016_, new_n891_, new_n911_ );
xnor g674 ( new_n1017_, new_n1016_, keyIn_0_145 );
not g675 ( new_n1018_, new_n1017_ );
not g676 ( new_n1019_, keyIn_0_227 );
not g677 ( new_n1020_, keyIn_0_224 );
nand g678 ( new_n1021_, new_n860_, new_n844_, new_n861_, new_n876_ );
nand g679 ( new_n1022_, new_n1021_, new_n1020_ );
nand g680 ( new_n1023_, new_n896_, keyIn_0_224, new_n844_, new_n876_ );
nand g681 ( new_n1024_, new_n1023_, new_n1022_ );
and g682 ( new_n1025_, new_n901_, keyIn_0_189 );
nor g683 ( new_n1026_, new_n901_, keyIn_0_189 );
xor g684 ( new_n1027_, new_n906_, keyIn_0_169 );
nor g685 ( new_n1028_, new_n1027_, new_n1025_, new_n1026_ );
nand g686 ( new_n1029_, new_n1024_, new_n1019_, new_n1028_ );
nand g687 ( new_n1030_, new_n1024_, new_n1028_ );
nand g688 ( new_n1031_, new_n1030_, keyIn_0_227 );
nand g689 ( new_n1032_, new_n1031_, new_n1029_ );
nand g690 ( new_n1033_, new_n1032_, keyIn_0_236, new_n1018_ );
not g691 ( new_n1034_, keyIn_0_236 );
nand g692 ( new_n1035_, new_n1032_, new_n1018_ );
nand g693 ( new_n1036_, new_n1035_, new_n1034_ );
nand g694 ( new_n1037_, new_n1036_, new_n1033_ );
nand g695 ( new_n1038_, new_n1031_, new_n1017_, new_n1029_ );
xnor g696 ( new_n1039_, new_n1038_, keyIn_0_235 );
nand g697 ( new_n1040_, new_n1037_, new_n1039_ );
nand g698 ( new_n1041_, new_n1040_, keyIn_0_245 );
not g699 ( new_n1042_, keyIn_0_245 );
nand g700 ( new_n1043_, new_n1037_, new_n1039_, new_n1042_ );
nand g701 ( new_n1044_, new_n1041_, N219, new_n1043_ );
nand g702 ( new_n1045_, N91, N210 );
nand g703 ( new_n1046_, new_n1044_, new_n1045_ );
nand g704 ( new_n1047_, new_n1046_, new_n1015_ );
nand g705 ( new_n1048_, new_n1044_, keyIn_0_251, new_n1045_ );
nand g706 ( new_n1049_, new_n1047_, new_n1048_ );
nand g707 ( new_n1050_, new_n1018_, N228 );
nand g708 ( new_n1051_, new_n912_, N237 );
nand g709 ( new_n1052_, new_n1050_, new_n1051_ );
nor g710 ( new_n1053_, new_n1052_, keyIn_0_193 );
and g711 ( new_n1054_, new_n1052_, keyIn_0_193 );
nand g712 ( new_n1055_, new_n889_, N246 );
xnor g713 ( new_n1056_, new_n1055_, keyIn_0_123 );
nand g714 ( new_n1057_, new_n607_, N165 );
nand g715 ( new_n1058_, new_n1056_, new_n1057_ );
xor g716 ( new_n1059_, new_n1058_, keyIn_0_146 );
nor g717 ( new_n1060_, new_n1054_, new_n1053_, new_n1059_ );
nand g718 ( new_n1061_, new_n1049_, keyIn_0_254, new_n1060_ );
not g719 ( new_n1062_, keyIn_0_254 );
nand g720 ( new_n1063_, new_n1049_, new_n1060_ );
nand g721 ( new_n1064_, new_n1063_, new_n1062_ );
nand g722 ( N879, new_n1064_, new_n1061_ );
not g723 ( new_n1066_, keyIn_0_255 );
not g724 ( new_n1067_, keyIn_0_246 );
not g725 ( new_n1068_, keyIn_0_238 );
nand g726 ( new_n1069_, new_n896_, new_n844_ );
nand g727 ( new_n1070_, new_n1069_, keyIn_0_223 );
or g728 ( new_n1071_, new_n1069_, keyIn_0_223 );
xor g729 ( new_n1072_, new_n900_, keyIn_0_171 );
nand g730 ( new_n1073_, new_n1071_, new_n1070_, new_n1072_ );
nand g731 ( new_n1074_, new_n1073_, keyIn_0_228 );
not g732 ( new_n1075_, keyIn_0_228 );
nand g733 ( new_n1076_, new_n1071_, new_n1075_, new_n1070_, new_n1072_ );
nand g734 ( new_n1077_, new_n1074_, new_n1076_ );
nand g735 ( new_n1078_, new_n905_, new_n876_ );
xor g736 ( new_n1079_, new_n1078_, keyIn_0_148 );
not g737 ( new_n1080_, new_n1079_ );
nand g738 ( new_n1081_, new_n1077_, new_n1080_ );
nand g739 ( new_n1082_, new_n1081_, new_n1068_ );
nand g740 ( new_n1083_, new_n1077_, keyIn_0_238, new_n1080_ );
nand g741 ( new_n1084_, new_n1082_, new_n1083_ );
nand g742 ( new_n1085_, new_n1074_, new_n1076_, new_n1079_ );
xnor g743 ( new_n1086_, new_n1085_, keyIn_0_237 );
nand g744 ( new_n1087_, new_n1084_, new_n1086_, new_n1067_ );
nand g745 ( new_n1088_, new_n1084_, new_n1086_ );
nand g746 ( new_n1089_, new_n1088_, keyIn_0_246 );
nand g747 ( new_n1090_, new_n1089_, N219, new_n1087_ );
nand g748 ( new_n1091_, N96, N210 );
nand g749 ( new_n1092_, new_n1090_, keyIn_0_252, new_n1091_ );
not g750 ( new_n1093_, keyIn_0_252 );
nand g751 ( new_n1094_, new_n1090_, new_n1091_ );
nand g752 ( new_n1095_, new_n1094_, new_n1093_ );
and g753 ( new_n1096_, new_n906_, N237 );
or g754 ( new_n1097_, new_n1096_, keyIn_0_170 );
nand g755 ( new_n1098_, new_n1080_, N228 );
nand g756 ( new_n1099_, new_n1096_, keyIn_0_170 );
nand g757 ( new_n1100_, new_n1098_, new_n1097_, new_n1099_ );
nor g758 ( new_n1101_, new_n1100_, keyIn_0_194 );
and g759 ( new_n1102_, new_n1100_, keyIn_0_194 );
and g760 ( new_n1103_, new_n874_, N246 );
nand g761 ( new_n1104_, new_n1103_, keyIn_0_126 );
or g762 ( new_n1105_, new_n1103_, keyIn_0_126 );
nand g763 ( new_n1106_, new_n607_, N171 );
nand g764 ( new_n1107_, new_n1105_, new_n1104_, new_n1106_ );
xnor g765 ( new_n1108_, new_n1107_, keyIn_0_149 );
nor g766 ( new_n1109_, new_n1102_, new_n1101_, new_n1108_ );
nand g767 ( new_n1110_, new_n1095_, new_n1066_, new_n1092_, new_n1109_ );
nand g768 ( new_n1111_, new_n1095_, new_n1092_, new_n1109_ );
nand g769 ( new_n1112_, new_n1111_, keyIn_0_255 );
nand g770 ( N880, new_n1112_, new_n1110_ );
endmodule