module add_mul_comp_16_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        a_8_, a_9_, a_10_, a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, 
        b_3_, b_4_, b_5_, b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, 
        b_14_, b_15_, Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, 
        Result_5_, Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, 
        Result_11_, Result_12_, Result_13_, Result_14_, Result_15_, Result_16_, 
        Result_17_, Result_18_, Result_19_, Result_20_, Result_21_, Result_22_, 
        Result_23_, Result_24_, Result_25_, Result_26_, Result_27_, Result_28_, 
        Result_29_, Result_30_, Result_31_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, a_8_, a_9_, a_10_,
         a_11_, a_12_, a_13_, a_14_, a_15_, b_0_, b_1_, b_2_, b_3_, b_4_, b_5_,
         b_6_, b_7_, b_8_, b_9_, b_10_, b_11_, b_12_, b_13_, b_14_, b_15_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_, Result_16_,
         Result_17_, Result_18_, Result_19_, Result_20_, Result_21_,
         Result_22_, Result_23_, Result_24_, Result_25_, Result_26_,
         Result_27_, Result_28_, Result_29_, Result_30_, Result_31_;
  wire   n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
         n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
         n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
         n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
         n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
         n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
         n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
         n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896;

  NOR2_X2 U1949 ( .A1(n3792), .A2(n1973), .ZN(n2215) );
  INV_X2 U1950 ( .A(n1957), .ZN(n1917) );
  NOR2_X1 U1951 ( .A1(n1917), .A2(n1918), .ZN(Result_9_) );
  XOR2_X1 U1952 ( .A(n1919), .B(n1920), .Z(n1918) );
  NAND2_X1 U1953 ( .A1(n1921), .A2(n1922), .ZN(n1920) );
  NOR2_X1 U1954 ( .A1(n1917), .A2(n1923), .ZN(Result_8_) );
  XOR2_X1 U1955 ( .A(n1924), .B(n1925), .Z(n1923) );
  NAND2_X1 U1956 ( .A1(n1926), .A2(n1927), .ZN(n1925) );
  NOR2_X1 U1957 ( .A1(n1917), .A2(n1928), .ZN(Result_7_) );
  XOR2_X1 U1958 ( .A(n1929), .B(n1930), .Z(n1928) );
  NAND2_X1 U1959 ( .A1(n1931), .A2(n1932), .ZN(n1930) );
  NOR2_X1 U1960 ( .A1(n1917), .A2(n1933), .ZN(Result_6_) );
  XOR2_X1 U1961 ( .A(n1934), .B(n1935), .Z(n1933) );
  NAND2_X1 U1962 ( .A1(n1936), .A2(n1937), .ZN(n1935) );
  NOR2_X1 U1963 ( .A1(n1917), .A2(n1938), .ZN(Result_5_) );
  XOR2_X1 U1964 ( .A(n1939), .B(n1940), .Z(n1938) );
  NAND2_X1 U1965 ( .A1(n1941), .A2(n1942), .ZN(n1940) );
  NOR2_X1 U1966 ( .A1(n1917), .A2(n1943), .ZN(Result_4_) );
  XOR2_X1 U1967 ( .A(n1944), .B(n1945), .Z(n1943) );
  NAND2_X1 U1968 ( .A1(n1946), .A2(n1947), .ZN(n1945) );
  NOR2_X1 U1969 ( .A1(n1917), .A2(n1948), .ZN(Result_3_) );
  XOR2_X1 U1970 ( .A(n1949), .B(n1950), .Z(n1948) );
  NAND2_X1 U1971 ( .A1(n1951), .A2(n1952), .ZN(n1950) );
  NAND2_X1 U1972 ( .A1(n1953), .A2(n1954), .ZN(Result_31_) );
  NAND3_X1 U1973 ( .A1(n1917), .A2(a_15_), .A3(n1955), .ZN(n1954) );
  NAND2_X1 U1974 ( .A1(n1956), .A2(b_15_), .ZN(n1953) );
  XNOR2_X1 U1975 ( .A(a_15_), .B(n1957), .ZN(n1956) );
  NAND2_X1 U1976 ( .A1(n1958), .A2(n1959), .ZN(Result_30_) );
  NAND2_X1 U1977 ( .A1(n1960), .A2(n1957), .ZN(n1959) );
  NAND2_X1 U1978 ( .A1(n1961), .A2(n1962), .ZN(n1960) );
  NAND2_X1 U1979 ( .A1(b_14_), .A2(n1963), .ZN(n1962) );
  NAND2_X1 U1980 ( .A1(n1964), .A2(n1965), .ZN(n1963) );
  NAND2_X1 U1981 ( .A1(b_15_), .A2(n1966), .ZN(n1961) );
  NAND2_X1 U1982 ( .A1(n1967), .A2(n1968), .ZN(n1966) );
  NAND2_X1 U1983 ( .A1(a_14_), .A2(n1969), .ZN(n1968) );
  NAND2_X1 U1984 ( .A1(n1970), .A2(n1917), .ZN(n1958) );
  XOR2_X1 U1985 ( .A(n1971), .B(n1972), .Z(n1970) );
  XNOR2_X1 U1986 ( .A(n1969), .B(a_14_), .ZN(n1972) );
  NOR2_X1 U1987 ( .A1(n1955), .A2(n1973), .ZN(n1971) );
  NOR2_X1 U1988 ( .A1(n1917), .A2(n1974), .ZN(Result_2_) );
  XOR2_X1 U1989 ( .A(n1975), .B(n1976), .Z(n1974) );
  NAND2_X1 U1990 ( .A1(n1977), .A2(n1978), .ZN(n1976) );
  NAND2_X1 U1991 ( .A1(n1979), .A2(n1980), .ZN(Result_29_) );
  NAND2_X1 U1992 ( .A1(n1917), .A2(n1981), .ZN(n1980) );
  NAND3_X1 U1993 ( .A1(n1982), .A2(n1983), .A3(n1984), .ZN(n1981) );
  NAND2_X1 U1994 ( .A1(n1985), .A2(n1986), .ZN(n1984) );
  NAND3_X1 U1995 ( .A1(n1987), .A2(n1988), .A3(b_13_), .ZN(n1983) );
  NAND2_X1 U1996 ( .A1(n1989), .A2(n1990), .ZN(n1982) );
  XNOR2_X1 U1997 ( .A(a_13_), .B(n1987), .ZN(n1989) );
  INV_X1 U1998 ( .A(n1986), .ZN(n1987) );
  NAND2_X1 U1999 ( .A1(n1991), .A2(n1957), .ZN(n1979) );
  XOR2_X1 U2000 ( .A(n1992), .B(n1993), .Z(n1991) );
  NOR2_X1 U2001 ( .A1(n1955), .A2(n1988), .ZN(n1993) );
  XOR2_X1 U2002 ( .A(n1994), .B(n1995), .Z(n1992) );
  NAND2_X1 U2003 ( .A1(n1996), .A2(n1997), .ZN(Result_28_) );
  NAND2_X1 U2004 ( .A1(n1998), .A2(n1957), .ZN(n1997) );
  XOR2_X1 U2005 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR2_X1 U2006 ( .A(n2001), .B(n2002), .Z(n2000) );
  NOR2_X1 U2007 ( .A1(n1955), .A2(n2003), .ZN(n2002) );
  NAND2_X1 U2008 ( .A1(n2004), .A2(n1917), .ZN(n1996) );
  XOR2_X1 U2009 ( .A(n2005), .B(n2006), .Z(n2004) );
  AND2_X1 U2010 ( .A1(n2007), .A2(n2008), .ZN(n2006) );
  NAND2_X1 U2011 ( .A1(n2009), .A2(n2010), .ZN(Result_27_) );
  NAND2_X1 U2012 ( .A1(n1917), .A2(n2011), .ZN(n2010) );
  NAND3_X1 U2013 ( .A1(n2012), .A2(n2013), .A3(n2014), .ZN(n2011) );
  NAND2_X1 U2014 ( .A1(n2015), .A2(n2016), .ZN(n2014) );
  OR3_X1 U2015 ( .A1(n2016), .A2(a_11_), .A3(n2017), .ZN(n2013) );
  NAND2_X1 U2016 ( .A1(n2018), .A2(n2017), .ZN(n2012) );
  XNOR2_X1 U2017 ( .A(n2016), .B(n2019), .ZN(n2018) );
  NAND2_X1 U2018 ( .A1(n2020), .A2(n1957), .ZN(n2009) );
  XNOR2_X1 U2019 ( .A(n2021), .B(n2022), .ZN(n2020) );
  NAND2_X1 U2020 ( .A1(n2023), .A2(n2024), .ZN(n2021) );
  NAND2_X1 U2021 ( .A1(n2025), .A2(n2026), .ZN(Result_26_) );
  NAND2_X1 U2022 ( .A1(n2027), .A2(n1957), .ZN(n2026) );
  XNOR2_X1 U2023 ( .A(n2028), .B(n2029), .ZN(n2027) );
  XOR2_X1 U2024 ( .A(n2030), .B(n2031), .Z(n2029) );
  NAND2_X1 U2025 ( .A1(a_10_), .A2(b_15_), .ZN(n2031) );
  NAND2_X1 U2026 ( .A1(n2032), .A2(n1917), .ZN(n2025) );
  XNOR2_X1 U2027 ( .A(n2033), .B(n2034), .ZN(n2032) );
  NOR2_X1 U2028 ( .A1(n2035), .A2(n2036), .ZN(n2034) );
  NAND2_X1 U2029 ( .A1(n2037), .A2(n2038), .ZN(Result_25_) );
  NAND2_X1 U2030 ( .A1(n1917), .A2(n2039), .ZN(n2038) );
  NAND3_X1 U2031 ( .A1(n2040), .A2(n2041), .A3(n2042), .ZN(n2039) );
  NAND2_X1 U2032 ( .A1(n2043), .A2(n2044), .ZN(n2042) );
  NAND3_X1 U2033 ( .A1(n2045), .A2(n2046), .A3(b_9_), .ZN(n2041) );
  NAND2_X1 U2034 ( .A1(n2047), .A2(n2048), .ZN(n2040) );
  XNOR2_X1 U2035 ( .A(n2045), .B(a_9_), .ZN(n2047) );
  NAND2_X1 U2036 ( .A1(n2049), .A2(n1957), .ZN(n2037) );
  XNOR2_X1 U2037 ( .A(n2050), .B(n2051), .ZN(n2049) );
  XOR2_X1 U2038 ( .A(n2052), .B(n2053), .Z(n2051) );
  NAND2_X1 U2039 ( .A1(a_9_), .A2(b_15_), .ZN(n2053) );
  NAND2_X1 U2040 ( .A1(n2054), .A2(n2055), .ZN(Result_24_) );
  NAND2_X1 U2041 ( .A1(n2056), .A2(n1957), .ZN(n2055) );
  XOR2_X1 U2042 ( .A(n2057), .B(n2058), .Z(n2056) );
  XNOR2_X1 U2043 ( .A(n2059), .B(n2060), .ZN(n2058) );
  NAND2_X1 U2044 ( .A1(a_8_), .A2(b_15_), .ZN(n2060) );
  NAND2_X1 U2045 ( .A1(n2061), .A2(n1917), .ZN(n2054) );
  XOR2_X1 U2046 ( .A(n2062), .B(n2063), .Z(n2061) );
  AND2_X1 U2047 ( .A1(n2064), .A2(n2065), .ZN(n2063) );
  NAND2_X1 U2048 ( .A1(n2066), .A2(n2067), .ZN(Result_23_) );
  NAND2_X1 U2049 ( .A1(n1917), .A2(n2068), .ZN(n2067) );
  NAND3_X1 U2050 ( .A1(n2069), .A2(n2070), .A3(n2071), .ZN(n2068) );
  NAND2_X1 U2051 ( .A1(n2072), .A2(n2073), .ZN(n2071) );
  OR3_X1 U2052 ( .A1(n2073), .A2(a_7_), .A3(n2074), .ZN(n2070) );
  NAND2_X1 U2053 ( .A1(n2075), .A2(n2074), .ZN(n2069) );
  XNOR2_X1 U2054 ( .A(n2073), .B(n2076), .ZN(n2075) );
  NAND2_X1 U2055 ( .A1(n2077), .A2(n1957), .ZN(n2066) );
  XNOR2_X1 U2056 ( .A(n2078), .B(n2079), .ZN(n2077) );
  NAND2_X1 U2057 ( .A1(n2080), .A2(n2081), .ZN(n2078) );
  NAND2_X1 U2058 ( .A1(n2082), .A2(n2083), .ZN(Result_22_) );
  NAND2_X1 U2059 ( .A1(n2084), .A2(n1957), .ZN(n2083) );
  XOR2_X1 U2060 ( .A(n2085), .B(n2086), .Z(n2084) );
  XOR2_X1 U2061 ( .A(n2087), .B(n2088), .Z(n2086) );
  NOR2_X1 U2062 ( .A1(n1955), .A2(n2089), .ZN(n2088) );
  NAND2_X1 U2063 ( .A1(n2090), .A2(n1917), .ZN(n2082) );
  XNOR2_X1 U2064 ( .A(n2091), .B(n2092), .ZN(n2090) );
  NOR2_X1 U2065 ( .A1(n2093), .A2(n2094), .ZN(n2092) );
  NAND2_X1 U2066 ( .A1(n2095), .A2(n2096), .ZN(Result_21_) );
  NAND2_X1 U2067 ( .A1(n1917), .A2(n2097), .ZN(n2096) );
  NAND3_X1 U2068 ( .A1(n2098), .A2(n2099), .A3(n2100), .ZN(n2097) );
  NAND2_X1 U2069 ( .A1(n2101), .A2(n2102), .ZN(n2100) );
  NAND3_X1 U2070 ( .A1(n2103), .A2(n2104), .A3(b_5_), .ZN(n2099) );
  NAND2_X1 U2071 ( .A1(n2105), .A2(n2106), .ZN(n2098) );
  XNOR2_X1 U2072 ( .A(n2103), .B(a_5_), .ZN(n2105) );
  NAND2_X1 U2073 ( .A1(n2107), .A2(n1957), .ZN(n2095) );
  XNOR2_X1 U2074 ( .A(n2108), .B(n2109), .ZN(n2107) );
  NAND2_X1 U2075 ( .A1(n2110), .A2(n2111), .ZN(n2108) );
  NAND2_X1 U2076 ( .A1(n2112), .A2(n2113), .ZN(Result_20_) );
  NAND2_X1 U2077 ( .A1(n2114), .A2(n1957), .ZN(n2113) );
  XOR2_X1 U2078 ( .A(n2115), .B(n2116), .Z(n2114) );
  XOR2_X1 U2079 ( .A(n2117), .B(n2118), .Z(n2116) );
  NOR2_X1 U2080 ( .A1(n1955), .A2(n2119), .ZN(n2118) );
  NAND2_X1 U2081 ( .A1(n2120), .A2(n1917), .ZN(n2112) );
  XNOR2_X1 U2082 ( .A(n2121), .B(n2122), .ZN(n2120) );
  NOR2_X1 U2083 ( .A1(n2123), .A2(n2124), .ZN(n2122) );
  NOR2_X1 U2084 ( .A1(n1917), .A2(n2125), .ZN(Result_1_) );
  XOR2_X1 U2085 ( .A(n2126), .B(n2127), .Z(n2125) );
  NAND2_X1 U2086 ( .A1(n2128), .A2(n2129), .ZN(n2127) );
  NAND2_X1 U2087 ( .A1(n2130), .A2(n2131), .ZN(Result_19_) );
  NAND2_X1 U2088 ( .A1(n1917), .A2(n2132), .ZN(n2131) );
  NAND3_X1 U2089 ( .A1(n2133), .A2(n2134), .A3(n2135), .ZN(n2132) );
  NAND2_X1 U2090 ( .A1(n2136), .A2(n2137), .ZN(n2135) );
  NAND3_X1 U2091 ( .A1(n2138), .A2(n2139), .A3(b_3_), .ZN(n2134) );
  NAND2_X1 U2092 ( .A1(n2140), .A2(n2141), .ZN(n2133) );
  XNOR2_X1 U2093 ( .A(n2138), .B(a_3_), .ZN(n2140) );
  NAND2_X1 U2094 ( .A1(n2142), .A2(n1957), .ZN(n2130) );
  XNOR2_X1 U2095 ( .A(n2143), .B(n2144), .ZN(n2142) );
  XOR2_X1 U2096 ( .A(n2145), .B(n2146), .Z(n2144) );
  NAND2_X1 U2097 ( .A1(a_3_), .A2(b_15_), .ZN(n2146) );
  NAND2_X1 U2098 ( .A1(n2147), .A2(n2148), .ZN(Result_18_) );
  NAND2_X1 U2099 ( .A1(n2149), .A2(n1957), .ZN(n2148) );
  XOR2_X1 U2100 ( .A(n2150), .B(n2151), .Z(n2149) );
  XNOR2_X1 U2101 ( .A(n2152), .B(n2153), .ZN(n2151) );
  NAND2_X1 U2102 ( .A1(a_2_), .A2(b_15_), .ZN(n2153) );
  NAND2_X1 U2103 ( .A1(n2154), .A2(n1917), .ZN(n2147) );
  XOR2_X1 U2104 ( .A(n2155), .B(n2156), .Z(n2154) );
  AND2_X1 U2105 ( .A1(n2157), .A2(n2158), .ZN(n2156) );
  NAND2_X1 U2106 ( .A1(n2159), .A2(n2160), .ZN(Result_17_) );
  NAND2_X1 U2107 ( .A1(n2161), .A2(n1957), .ZN(n2160) );
  XOR2_X1 U2108 ( .A(n2162), .B(n2163), .Z(n2161) );
  XNOR2_X1 U2109 ( .A(n2164), .B(n2165), .ZN(n2163) );
  NAND2_X1 U2110 ( .A1(b_15_), .A2(a_1_), .ZN(n2165) );
  NAND2_X1 U2111 ( .A1(n2166), .A2(n1917), .ZN(n2159) );
  NAND2_X1 U2112 ( .A1(n2167), .A2(n2168), .ZN(n2166) );
  NAND2_X1 U2113 ( .A1(n2169), .A2(n2170), .ZN(n2168) );
  OR2_X1 U2114 ( .A1(n2171), .A2(n2172), .ZN(n2169) );
  NAND2_X1 U2115 ( .A1(n2173), .A2(n2174), .ZN(n2167) );
  INV_X1 U2116 ( .A(n2170), .ZN(n2174) );
  XNOR2_X1 U2117 ( .A(n2175), .B(a_1_), .ZN(n2173) );
  NAND2_X1 U2118 ( .A1(n2176), .A2(n2177), .ZN(Result_16_) );
  NAND2_X1 U2119 ( .A1(n2178), .A2(n1957), .ZN(n2177) );
  XOR2_X1 U2120 ( .A(n2179), .B(n2180), .Z(n2178) );
  XNOR2_X1 U2121 ( .A(n2181), .B(n2182), .ZN(n2180) );
  NAND2_X1 U2122 ( .A1(a_0_), .A2(b_15_), .ZN(n2182) );
  NAND2_X1 U2123 ( .A1(n2183), .A2(n1917), .ZN(n2176) );
  XNOR2_X1 U2124 ( .A(n2184), .B(n2185), .ZN(n2183) );
  NOR2_X1 U2125 ( .A1(n2172), .A2(n2186), .ZN(n2184) );
  NOR2_X1 U2126 ( .A1(n2171), .A2(n2170), .ZN(n2186) );
  NAND2_X1 U2127 ( .A1(n2158), .A2(n2187), .ZN(n2170) );
  NAND2_X1 U2128 ( .A1(n2157), .A2(n2155), .ZN(n2187) );
  NAND2_X1 U2129 ( .A1(n2188), .A2(n2189), .ZN(n2155) );
  NAND2_X1 U2130 ( .A1(n2190), .A2(n2137), .ZN(n2189) );
  INV_X1 U2131 ( .A(n2138), .ZN(n2137) );
  NOR2_X1 U2132 ( .A1(n2124), .A2(n2191), .ZN(n2138) );
  NOR2_X1 U2133 ( .A1(n2123), .A2(n2121), .ZN(n2191) );
  AND2_X1 U2134 ( .A1(n2192), .A2(n2193), .ZN(n2121) );
  NAND2_X1 U2135 ( .A1(n2194), .A2(n2102), .ZN(n2193) );
  INV_X1 U2136 ( .A(n2103), .ZN(n2102) );
  NOR2_X1 U2137 ( .A1(n2094), .A2(n2195), .ZN(n2103) );
  NOR2_X1 U2138 ( .A1(n2093), .A2(n2091), .ZN(n2195) );
  AND2_X1 U2139 ( .A1(n2196), .A2(n2197), .ZN(n2091) );
  NAND2_X1 U2140 ( .A1(n2198), .A2(n2073), .ZN(n2197) );
  NAND2_X1 U2141 ( .A1(n2065), .A2(n2199), .ZN(n2073) );
  NAND2_X1 U2142 ( .A1(n2064), .A2(n2062), .ZN(n2199) );
  NAND2_X1 U2143 ( .A1(n2200), .A2(n2201), .ZN(n2062) );
  NAND2_X1 U2144 ( .A1(n2202), .A2(n2044), .ZN(n2201) );
  INV_X1 U2145 ( .A(n2045), .ZN(n2044) );
  NOR2_X1 U2146 ( .A1(n2036), .A2(n2203), .ZN(n2045) );
  NOR2_X1 U2147 ( .A1(n2035), .A2(n2033), .ZN(n2203) );
  AND2_X1 U2148 ( .A1(n2204), .A2(n2205), .ZN(n2033) );
  NAND2_X1 U2149 ( .A1(n2206), .A2(n2016), .ZN(n2205) );
  NAND2_X1 U2150 ( .A1(n2008), .A2(n2207), .ZN(n2016) );
  NAND2_X1 U2151 ( .A1(n2007), .A2(n2005), .ZN(n2207) );
  NAND2_X1 U2152 ( .A1(n2208), .A2(n2209), .ZN(n2005) );
  NAND2_X1 U2153 ( .A1(n2210), .A2(n1986), .ZN(n2209) );
  NAND3_X1 U2154 ( .A1(n2211), .A2(n2212), .A3(n2213), .ZN(n1986) );
  NAND2_X1 U2155 ( .A1(a_14_), .A2(b_14_), .ZN(n2213) );
  NAND2_X1 U2156 ( .A1(n2214), .A2(a_15_), .ZN(n2212) );
  NAND2_X1 U2157 ( .A1(n2215), .A2(b_15_), .ZN(n2211) );
  NAND2_X1 U2158 ( .A1(n1990), .A2(n1988), .ZN(n2210) );
  NAND2_X1 U2159 ( .A1(n2216), .A2(n2003), .ZN(n2007) );
  NAND2_X1 U2160 ( .A1(n2017), .A2(n2019), .ZN(n2206) );
  NOR2_X1 U2161 ( .A1(b_10_), .A2(a_10_), .ZN(n2035) );
  NAND2_X1 U2162 ( .A1(n2048), .A2(n2046), .ZN(n2202) );
  NAND2_X1 U2163 ( .A1(n2217), .A2(n2218), .ZN(n2064) );
  NAND2_X1 U2164 ( .A1(n2074), .A2(n2076), .ZN(n2198) );
  NOR2_X1 U2165 ( .A1(b_6_), .A2(a_6_), .ZN(n2093) );
  NAND2_X1 U2166 ( .A1(n2106), .A2(n2104), .ZN(n2194) );
  NOR2_X1 U2167 ( .A1(b_4_), .A2(a_4_), .ZN(n2123) );
  NAND2_X1 U2168 ( .A1(n2141), .A2(n2139), .ZN(n2190) );
  NAND2_X1 U2169 ( .A1(n2219), .A2(n2220), .ZN(n2157) );
  NOR2_X1 U2170 ( .A1(b_1_), .A2(a_1_), .ZN(n2172) );
  NOR2_X1 U2171 ( .A1(n1917), .A2(n2221), .ZN(Result_15_) );
  XNOR2_X1 U2172 ( .A(n2222), .B(n2223), .ZN(n2221) );
  NOR3_X1 U2173 ( .A1(n2224), .A2(n2225), .A3(n1917), .ZN(Result_14_) );
  NOR2_X1 U2174 ( .A1(n2226), .A2(n2227), .ZN(n2224) );
  AND2_X1 U2175 ( .A1(n2223), .A2(n2222), .ZN(n2226) );
  NOR2_X1 U2176 ( .A1(n1917), .A2(n2228), .ZN(Result_13_) );
  XOR2_X1 U2177 ( .A(n2229), .B(n2225), .Z(n2228) );
  NAND2_X1 U2178 ( .A1(n2230), .A2(n2231), .ZN(n2229) );
  NAND2_X1 U2179 ( .A1(n2232), .A2(n2233), .ZN(n2230) );
  NAND2_X1 U2180 ( .A1(n2234), .A2(n2235), .ZN(n2233) );
  NOR2_X1 U2181 ( .A1(n1917), .A2(n2236), .ZN(Result_12_) );
  XNOR2_X1 U2182 ( .A(n2237), .B(n2238), .ZN(n2236) );
  NOR2_X1 U2183 ( .A1(n1917), .A2(n2239), .ZN(Result_11_) );
  XOR2_X1 U2184 ( .A(n2240), .B(n2241), .Z(n2239) );
  NAND2_X1 U2185 ( .A1(n2242), .A2(n2243), .ZN(n2240) );
  NAND2_X1 U2186 ( .A1(n2244), .A2(n2245), .ZN(n2242) );
  NOR2_X1 U2187 ( .A1(n1917), .A2(n2246), .ZN(Result_10_) );
  XOR2_X1 U2188 ( .A(n2247), .B(n2248), .Z(n2246) );
  NAND2_X1 U2189 ( .A1(n2249), .A2(n2250), .ZN(n2248) );
  NOR2_X1 U2190 ( .A1(n1917), .A2(n2251), .ZN(Result_0_) );
  AND3_X1 U2191 ( .A1(n2252), .A2(n2253), .A3(n2129), .ZN(n2251) );
  NAND4_X1 U2192 ( .A1(b_0_), .A2(n2253), .A3(n2254), .A4(n2255), .ZN(n2129)
         );
  NAND2_X1 U2193 ( .A1(n2126), .A2(n2128), .ZN(n2252) );
  NAND2_X1 U2194 ( .A1(n2256), .A2(n2257), .ZN(n2128) );
  NAND2_X1 U2195 ( .A1(b_0_), .A2(n2253), .ZN(n2257) );
  NAND2_X1 U2196 ( .A1(n2258), .A2(n2259), .ZN(n2253) );
  NAND2_X1 U2197 ( .A1(n2254), .A2(n2255), .ZN(n2256) );
  NAND2_X1 U2198 ( .A1(n1977), .A2(n2260), .ZN(n2126) );
  NAND2_X1 U2199 ( .A1(n1978), .A2(n1975), .ZN(n2260) );
  NAND2_X1 U2200 ( .A1(n1951), .A2(n2261), .ZN(n1975) );
  NAND2_X1 U2201 ( .A1(n1952), .A2(n1949), .ZN(n2261) );
  NAND2_X1 U2202 ( .A1(n1946), .A2(n2262), .ZN(n1949) );
  NAND2_X1 U2203 ( .A1(n1947), .A2(n1944), .ZN(n2262) );
  NAND2_X1 U2204 ( .A1(n1941), .A2(n2263), .ZN(n1944) );
  NAND2_X1 U2205 ( .A1(n1942), .A2(n1939), .ZN(n2263) );
  NAND2_X1 U2206 ( .A1(n1936), .A2(n2264), .ZN(n1939) );
  NAND2_X1 U2207 ( .A1(n1937), .A2(n1934), .ZN(n2264) );
  NAND2_X1 U2208 ( .A1(n1931), .A2(n2265), .ZN(n1934) );
  NAND2_X1 U2209 ( .A1(n1932), .A2(n1929), .ZN(n2265) );
  NAND2_X1 U2210 ( .A1(n1926), .A2(n2266), .ZN(n1929) );
  NAND2_X1 U2211 ( .A1(n1927), .A2(n1924), .ZN(n2266) );
  NAND2_X1 U2212 ( .A1(n1921), .A2(n2267), .ZN(n1924) );
  NAND2_X1 U2213 ( .A1(n1922), .A2(n1919), .ZN(n2267) );
  NAND2_X1 U2214 ( .A1(n2268), .A2(n2249), .ZN(n1919) );
  NAND2_X1 U2215 ( .A1(n2269), .A2(n2270), .ZN(n2249) );
  NAND2_X1 U2216 ( .A1(n2247), .A2(n2250), .ZN(n2268) );
  OR2_X1 U2217 ( .A1(n2270), .A2(n2269), .ZN(n2250) );
  XOR2_X1 U2218 ( .A(n2271), .B(n2272), .Z(n2270) );
  NAND2_X1 U2219 ( .A1(n2273), .A2(n2243), .ZN(n2247) );
  OR2_X1 U2220 ( .A1(n2244), .A2(n2245), .ZN(n2243) );
  NAND2_X1 U2221 ( .A1(n2274), .A2(n2275), .ZN(n2245) );
  INV_X1 U2222 ( .A(n2276), .ZN(n2244) );
  NAND2_X1 U2223 ( .A1(n2241), .A2(n2276), .ZN(n2273) );
  NOR2_X1 U2224 ( .A1(n2269), .A2(n2277), .ZN(n2276) );
  AND2_X1 U2225 ( .A1(n2278), .A2(n2279), .ZN(n2277) );
  NOR2_X1 U2226 ( .A1(n2279), .A2(n2278), .ZN(n2269) );
  XOR2_X1 U2227 ( .A(n2280), .B(n2281), .Z(n2278) );
  NAND2_X1 U2228 ( .A1(n2282), .A2(n2283), .ZN(n2280) );
  NAND2_X1 U2229 ( .A1(n2284), .A2(n2285), .ZN(n2279) );
  NAND2_X1 U2230 ( .A1(n2286), .A2(n2287), .ZN(n2285) );
  NAND2_X1 U2231 ( .A1(n2288), .A2(n2289), .ZN(n2287) );
  OR2_X1 U2232 ( .A1(n2289), .A2(n2288), .ZN(n2284) );
  AND2_X1 U2233 ( .A1(n2237), .A2(n2238), .ZN(n2241) );
  NAND3_X1 U2234 ( .A1(n2290), .A2(n2231), .A3(n2291), .ZN(n2238) );
  NAND2_X1 U2235 ( .A1(n2225), .A2(n2292), .ZN(n2291) );
  AND3_X1 U2236 ( .A1(n2222), .A2(n2223), .A3(n2227), .ZN(n2225) );
  XOR2_X1 U2237 ( .A(n2235), .B(n2234), .Z(n2227) );
  NAND2_X1 U2238 ( .A1(n2293), .A2(n2294), .ZN(n2223) );
  NAND3_X1 U2239 ( .A1(b_15_), .A2(n2295), .A3(a_0_), .ZN(n2294) );
  NAND2_X1 U2240 ( .A1(n2181), .A2(n2179), .ZN(n2295) );
  OR2_X1 U2241 ( .A1(n2179), .A2(n2181), .ZN(n2293) );
  AND2_X1 U2242 ( .A1(n2296), .A2(n2297), .ZN(n2181) );
  NAND3_X1 U2243 ( .A1(a_1_), .A2(n2298), .A3(b_15_), .ZN(n2297) );
  NAND2_X1 U2244 ( .A1(n2164), .A2(n2162), .ZN(n2298) );
  OR2_X1 U2245 ( .A1(n2162), .A2(n2164), .ZN(n2296) );
  AND2_X1 U2246 ( .A1(n2299), .A2(n2300), .ZN(n2164) );
  NAND3_X1 U2247 ( .A1(b_15_), .A2(n2301), .A3(a_2_), .ZN(n2300) );
  NAND2_X1 U2248 ( .A1(n2152), .A2(n2150), .ZN(n2301) );
  OR2_X1 U2249 ( .A1(n2150), .A2(n2152), .ZN(n2299) );
  AND2_X1 U2250 ( .A1(n2302), .A2(n2303), .ZN(n2152) );
  NAND3_X1 U2251 ( .A1(b_15_), .A2(n2304), .A3(a_3_), .ZN(n2303) );
  OR2_X1 U2252 ( .A1(n2145), .A2(n2143), .ZN(n2304) );
  NAND2_X1 U2253 ( .A1(n2143), .A2(n2145), .ZN(n2302) );
  NAND2_X1 U2254 ( .A1(n2305), .A2(n2306), .ZN(n2145) );
  NAND3_X1 U2255 ( .A1(b_15_), .A2(n2307), .A3(a_4_), .ZN(n2306) );
  OR2_X1 U2256 ( .A1(n2117), .A2(n2115), .ZN(n2307) );
  NAND2_X1 U2257 ( .A1(n2115), .A2(n2117), .ZN(n2305) );
  NAND2_X1 U2258 ( .A1(n2110), .A2(n2308), .ZN(n2117) );
  NAND2_X1 U2259 ( .A1(n2109), .A2(n2111), .ZN(n2308) );
  NAND2_X1 U2260 ( .A1(n2309), .A2(n2310), .ZN(n2111) );
  NAND2_X1 U2261 ( .A1(a_5_), .A2(b_15_), .ZN(n2310) );
  INV_X1 U2262 ( .A(n2311), .ZN(n2309) );
  XOR2_X1 U2263 ( .A(n2312), .B(n2313), .Z(n2109) );
  XOR2_X1 U2264 ( .A(n2314), .B(n2315), .Z(n2312) );
  NOR2_X1 U2265 ( .A1(n1969), .A2(n2089), .ZN(n2315) );
  NAND2_X1 U2266 ( .A1(a_5_), .A2(n2311), .ZN(n2110) );
  NAND2_X1 U2267 ( .A1(n2316), .A2(n2317), .ZN(n2311) );
  NAND3_X1 U2268 ( .A1(b_15_), .A2(n2318), .A3(a_6_), .ZN(n2317) );
  NAND2_X1 U2269 ( .A1(n2087), .A2(n2085), .ZN(n2318) );
  OR2_X1 U2270 ( .A1(n2085), .A2(n2087), .ZN(n2316) );
  AND2_X1 U2271 ( .A1(n2080), .A2(n2319), .ZN(n2087) );
  NAND2_X1 U2272 ( .A1(n2079), .A2(n2081), .ZN(n2319) );
  NAND2_X1 U2273 ( .A1(n2320), .A2(n2321), .ZN(n2081) );
  NAND2_X1 U2274 ( .A1(a_7_), .A2(b_15_), .ZN(n2321) );
  INV_X1 U2275 ( .A(n2322), .ZN(n2320) );
  XOR2_X1 U2276 ( .A(n2323), .B(n2324), .Z(n2079) );
  XNOR2_X1 U2277 ( .A(n2325), .B(n2326), .ZN(n2323) );
  NAND2_X1 U2278 ( .A1(a_8_), .A2(b_14_), .ZN(n2325) );
  NAND2_X1 U2279 ( .A1(a_7_), .A2(n2322), .ZN(n2080) );
  NAND2_X1 U2280 ( .A1(n2327), .A2(n2328), .ZN(n2322) );
  NAND3_X1 U2281 ( .A1(b_15_), .A2(n2329), .A3(a_8_), .ZN(n2328) );
  NAND2_X1 U2282 ( .A1(n2059), .A2(n2057), .ZN(n2329) );
  OR2_X1 U2283 ( .A1(n2057), .A2(n2059), .ZN(n2327) );
  AND2_X1 U2284 ( .A1(n2330), .A2(n2331), .ZN(n2059) );
  NAND3_X1 U2285 ( .A1(b_15_), .A2(n2332), .A3(a_9_), .ZN(n2331) );
  OR2_X1 U2286 ( .A1(n2052), .A2(n2050), .ZN(n2332) );
  NAND2_X1 U2287 ( .A1(n2050), .A2(n2052), .ZN(n2330) );
  NAND2_X1 U2288 ( .A1(n2333), .A2(n2334), .ZN(n2052) );
  NAND3_X1 U2289 ( .A1(b_15_), .A2(n2335), .A3(a_10_), .ZN(n2334) );
  OR2_X1 U2290 ( .A1(n2030), .A2(n2028), .ZN(n2335) );
  NAND2_X1 U2291 ( .A1(n2028), .A2(n2030), .ZN(n2333) );
  NAND2_X1 U2292 ( .A1(n2023), .A2(n2336), .ZN(n2030) );
  NAND2_X1 U2293 ( .A1(n2022), .A2(n2024), .ZN(n2336) );
  NAND2_X1 U2294 ( .A1(n2337), .A2(n2338), .ZN(n2024) );
  NAND2_X1 U2295 ( .A1(a_11_), .A2(b_15_), .ZN(n2338) );
  INV_X1 U2296 ( .A(n2339), .ZN(n2337) );
  XNOR2_X1 U2297 ( .A(n2340), .B(n2341), .ZN(n2022) );
  XOR2_X1 U2298 ( .A(n2342), .B(n2343), .Z(n2340) );
  NAND2_X1 U2299 ( .A1(a_12_), .A2(b_14_), .ZN(n2342) );
  NAND2_X1 U2300 ( .A1(a_11_), .A2(n2339), .ZN(n2023) );
  NAND2_X1 U2301 ( .A1(n2344), .A2(n2345), .ZN(n2339) );
  NAND3_X1 U2302 ( .A1(b_15_), .A2(n2346), .A3(a_12_), .ZN(n2345) );
  NAND2_X1 U2303 ( .A1(n2001), .A2(n1999), .ZN(n2346) );
  OR2_X1 U2304 ( .A1(n1999), .A2(n2001), .ZN(n2344) );
  AND2_X1 U2305 ( .A1(n2347), .A2(n2348), .ZN(n2001) );
  NAND3_X1 U2306 ( .A1(b_15_), .A2(n2349), .A3(a_13_), .ZN(n2348) );
  OR2_X1 U2307 ( .A1(n1994), .A2(n1995), .ZN(n2349) );
  NAND2_X1 U2308 ( .A1(n1995), .A2(n1994), .ZN(n2347) );
  NAND2_X1 U2309 ( .A1(n2350), .A2(n2351), .ZN(n1994) );
  NAND2_X1 U2310 ( .A1(b_13_), .A2(n2352), .ZN(n2351) );
  NAND2_X1 U2311 ( .A1(n1964), .A2(n2353), .ZN(n2352) );
  NAND2_X1 U2312 ( .A1(a_15_), .A2(n1969), .ZN(n2353) );
  NAND2_X1 U2313 ( .A1(b_14_), .A2(n2354), .ZN(n2350) );
  NAND2_X1 U2314 ( .A1(n1967), .A2(n2355), .ZN(n2354) );
  NAND2_X1 U2315 ( .A1(a_14_), .A2(n1990), .ZN(n2355) );
  AND2_X1 U2316 ( .A1(n2214), .A2(n2215), .ZN(n1995) );
  XNOR2_X1 U2317 ( .A(n2356), .B(n2357), .ZN(n1999) );
  XOR2_X1 U2318 ( .A(n2358), .B(n2359), .Z(n2356) );
  XNOR2_X1 U2319 ( .A(n2360), .B(n2361), .ZN(n2028) );
  NAND2_X1 U2320 ( .A1(n2362), .A2(n2363), .ZN(n2360) );
  XNOR2_X1 U2321 ( .A(n2364), .B(n2365), .ZN(n2050) );
  NAND2_X1 U2322 ( .A1(n2366), .A2(n2367), .ZN(n2364) );
  XNOR2_X1 U2323 ( .A(n2368), .B(n2369), .ZN(n2057) );
  XOR2_X1 U2324 ( .A(n2370), .B(n2371), .Z(n2368) );
  XOR2_X1 U2325 ( .A(n2372), .B(n2373), .Z(n2085) );
  XNOR2_X1 U2326 ( .A(n2374), .B(n2375), .ZN(n2373) );
  XOR2_X1 U2327 ( .A(n2376), .B(n2377), .Z(n2115) );
  XOR2_X1 U2328 ( .A(n2378), .B(n2379), .Z(n2376) );
  XNOR2_X1 U2329 ( .A(n2380), .B(n2381), .ZN(n2143) );
  XNOR2_X1 U2330 ( .A(n2382), .B(n2383), .ZN(n2380) );
  NOR2_X1 U2331 ( .A1(n1969), .A2(n2119), .ZN(n2383) );
  XOR2_X1 U2332 ( .A(n2384), .B(n2385), .Z(n2150) );
  XNOR2_X1 U2333 ( .A(n2386), .B(n2387), .ZN(n2385) );
  XOR2_X1 U2334 ( .A(n2388), .B(n2389), .Z(n2162) );
  XOR2_X1 U2335 ( .A(n2390), .B(n2391), .Z(n2389) );
  NAND2_X1 U2336 ( .A1(a_2_), .A2(b_14_), .ZN(n2391) );
  XNOR2_X1 U2337 ( .A(n2392), .B(n2393), .ZN(n2179) );
  XOR2_X1 U2338 ( .A(n2394), .B(n2395), .Z(n2392) );
  NOR2_X1 U2339 ( .A1(n2396), .A2(n1969), .ZN(n2395) );
  XNOR2_X1 U2340 ( .A(n2397), .B(n2398), .ZN(n2222) );
  XNOR2_X1 U2341 ( .A(n2399), .B(n2400), .ZN(n2398) );
  NAND3_X1 U2342 ( .A1(n2234), .A2(n2235), .A3(n2292), .ZN(n2231) );
  INV_X1 U2343 ( .A(n2232), .ZN(n2292) );
  NAND2_X1 U2344 ( .A1(n2290), .A2(n2401), .ZN(n2232) );
  NAND2_X1 U2345 ( .A1(n2402), .A2(n2403), .ZN(n2401) );
  NAND2_X1 U2346 ( .A1(n2404), .A2(n2405), .ZN(n2235) );
  NAND2_X1 U2347 ( .A1(n2400), .A2(n2406), .ZN(n2405) );
  OR2_X1 U2348 ( .A1(n2399), .A2(n2397), .ZN(n2406) );
  NOR2_X1 U2349 ( .A1(n2407), .A2(n1969), .ZN(n2400) );
  NAND2_X1 U2350 ( .A1(n2397), .A2(n2399), .ZN(n2404) );
  NAND2_X1 U2351 ( .A1(n2408), .A2(n2409), .ZN(n2399) );
  NAND3_X1 U2352 ( .A1(a_1_), .A2(n2410), .A3(b_14_), .ZN(n2409) );
  OR2_X1 U2353 ( .A1(n2394), .A2(n2393), .ZN(n2410) );
  NAND2_X1 U2354 ( .A1(n2393), .A2(n2394), .ZN(n2408) );
  NAND2_X1 U2355 ( .A1(n2411), .A2(n2412), .ZN(n2394) );
  NAND3_X1 U2356 ( .A1(b_14_), .A2(n2413), .A3(a_2_), .ZN(n2412) );
  OR2_X1 U2357 ( .A1(n2390), .A2(n2388), .ZN(n2413) );
  NAND2_X1 U2358 ( .A1(n2388), .A2(n2390), .ZN(n2411) );
  NAND2_X1 U2359 ( .A1(n2414), .A2(n2415), .ZN(n2390) );
  NAND2_X1 U2360 ( .A1(n2387), .A2(n2416), .ZN(n2415) );
  OR2_X1 U2361 ( .A1(n2386), .A2(n2384), .ZN(n2416) );
  NOR2_X1 U2362 ( .A1(n2139), .A2(n1969), .ZN(n2387) );
  NAND2_X1 U2363 ( .A1(n2384), .A2(n2386), .ZN(n2414) );
  NAND2_X1 U2364 ( .A1(n2417), .A2(n2418), .ZN(n2386) );
  NAND3_X1 U2365 ( .A1(b_14_), .A2(n2419), .A3(a_4_), .ZN(n2418) );
  NAND2_X1 U2366 ( .A1(n2382), .A2(n2381), .ZN(n2419) );
  OR2_X1 U2367 ( .A1(n2381), .A2(n2382), .ZN(n2417) );
  AND2_X1 U2368 ( .A1(n2420), .A2(n2421), .ZN(n2382) );
  NAND2_X1 U2369 ( .A1(n2379), .A2(n2422), .ZN(n2421) );
  OR2_X1 U2370 ( .A1(n2378), .A2(n2377), .ZN(n2422) );
  NOR2_X1 U2371 ( .A1(n2104), .A2(n1969), .ZN(n2379) );
  NAND2_X1 U2372 ( .A1(n2377), .A2(n2378), .ZN(n2420) );
  NAND2_X1 U2373 ( .A1(n2423), .A2(n2424), .ZN(n2378) );
  NAND3_X1 U2374 ( .A1(b_14_), .A2(n2425), .A3(a_6_), .ZN(n2424) );
  OR2_X1 U2375 ( .A1(n2314), .A2(n2313), .ZN(n2425) );
  NAND2_X1 U2376 ( .A1(n2313), .A2(n2314), .ZN(n2423) );
  NAND2_X1 U2377 ( .A1(n2426), .A2(n2427), .ZN(n2314) );
  NAND2_X1 U2378 ( .A1(n2375), .A2(n2428), .ZN(n2427) );
  OR2_X1 U2379 ( .A1(n2374), .A2(n2372), .ZN(n2428) );
  NOR2_X1 U2380 ( .A1(n2076), .A2(n1969), .ZN(n2375) );
  NAND2_X1 U2381 ( .A1(n2372), .A2(n2374), .ZN(n2426) );
  NAND2_X1 U2382 ( .A1(n2429), .A2(n2430), .ZN(n2374) );
  NAND3_X1 U2383 ( .A1(b_14_), .A2(n2431), .A3(a_8_), .ZN(n2430) );
  OR2_X1 U2384 ( .A1(n2326), .A2(n2324), .ZN(n2431) );
  NAND2_X1 U2385 ( .A1(n2324), .A2(n2326), .ZN(n2429) );
  NAND2_X1 U2386 ( .A1(n2432), .A2(n2433), .ZN(n2326) );
  NAND2_X1 U2387 ( .A1(n2371), .A2(n2434), .ZN(n2433) );
  OR2_X1 U2388 ( .A1(n2370), .A2(n2369), .ZN(n2434) );
  NOR2_X1 U2389 ( .A1(n2046), .A2(n1969), .ZN(n2371) );
  NAND2_X1 U2390 ( .A1(n2369), .A2(n2370), .ZN(n2432) );
  NAND2_X1 U2391 ( .A1(n2366), .A2(n2435), .ZN(n2370) );
  NAND2_X1 U2392 ( .A1(n2365), .A2(n2367), .ZN(n2435) );
  NAND2_X1 U2393 ( .A1(n2436), .A2(n2437), .ZN(n2367) );
  NAND2_X1 U2394 ( .A1(a_10_), .A2(b_14_), .ZN(n2437) );
  INV_X1 U2395 ( .A(n2438), .ZN(n2436) );
  XNOR2_X1 U2396 ( .A(n2439), .B(n2440), .ZN(n2365) );
  NAND2_X1 U2397 ( .A1(n2441), .A2(n2442), .ZN(n2439) );
  NAND2_X1 U2398 ( .A1(a_10_), .A2(n2438), .ZN(n2366) );
  NAND2_X1 U2399 ( .A1(n2362), .A2(n2443), .ZN(n2438) );
  NAND2_X1 U2400 ( .A1(n2361), .A2(n2363), .ZN(n2443) );
  NAND2_X1 U2401 ( .A1(n2444), .A2(n2445), .ZN(n2363) );
  NAND2_X1 U2402 ( .A1(a_11_), .A2(b_14_), .ZN(n2445) );
  INV_X1 U2403 ( .A(n2446), .ZN(n2444) );
  XNOR2_X1 U2404 ( .A(n2447), .B(n2448), .ZN(n2361) );
  XOR2_X1 U2405 ( .A(n2449), .B(n2450), .Z(n2447) );
  NAND2_X1 U2406 ( .A1(a_12_), .A2(b_13_), .ZN(n2449) );
  NAND2_X1 U2407 ( .A1(a_11_), .A2(n2446), .ZN(n2362) );
  NAND2_X1 U2408 ( .A1(n2451), .A2(n2452), .ZN(n2446) );
  NAND3_X1 U2409 ( .A1(b_14_), .A2(n2453), .A3(a_12_), .ZN(n2452) );
  NAND2_X1 U2410 ( .A1(n2343), .A2(n2341), .ZN(n2453) );
  OR2_X1 U2411 ( .A1(n2341), .A2(n2343), .ZN(n2451) );
  AND2_X1 U2412 ( .A1(n2454), .A2(n2455), .ZN(n2343) );
  NAND2_X1 U2413 ( .A1(n2357), .A2(n2456), .ZN(n2455) );
  OR2_X1 U2414 ( .A1(n2358), .A2(n2359), .ZN(n2456) );
  NOR2_X1 U2415 ( .A1(n1988), .A2(n1969), .ZN(n2357) );
  NAND2_X1 U2416 ( .A1(n2359), .A2(n2358), .ZN(n2454) );
  NAND2_X1 U2417 ( .A1(n2457), .A2(n2458), .ZN(n2358) );
  NAND2_X1 U2418 ( .A1(b_12_), .A2(n2459), .ZN(n2458) );
  NAND2_X1 U2419 ( .A1(n1964), .A2(n2460), .ZN(n2459) );
  NAND2_X1 U2420 ( .A1(a_15_), .A2(n1990), .ZN(n2460) );
  NAND2_X1 U2421 ( .A1(b_13_), .A2(n2461), .ZN(n2457) );
  NAND2_X1 U2422 ( .A1(n1967), .A2(n2462), .ZN(n2461) );
  NAND2_X1 U2423 ( .A1(a_14_), .A2(n2216), .ZN(n2462) );
  AND3_X1 U2424 ( .A1(b_13_), .A2(b_14_), .A3(n2215), .ZN(n2359) );
  XOR2_X1 U2425 ( .A(n2463), .B(n2208), .Z(n2341) );
  INV_X1 U2426 ( .A(n1985), .ZN(n2208) );
  XOR2_X1 U2427 ( .A(n2464), .B(n2465), .Z(n2463) );
  XNOR2_X1 U2428 ( .A(n2466), .B(n2467), .ZN(n2369) );
  NAND2_X1 U2429 ( .A1(n2468), .A2(n2469), .ZN(n2466) );
  XNOR2_X1 U2430 ( .A(n2470), .B(n2471), .ZN(n2324) );
  XNOR2_X1 U2431 ( .A(n2472), .B(n2473), .ZN(n2470) );
  XNOR2_X1 U2432 ( .A(n2474), .B(n2475), .ZN(n2372) );
  XOR2_X1 U2433 ( .A(n2476), .B(n2477), .Z(n2475) );
  NAND2_X1 U2434 ( .A1(a_8_), .A2(b_13_), .ZN(n2477) );
  XNOR2_X1 U2435 ( .A(n2478), .B(n2479), .ZN(n2313) );
  XNOR2_X1 U2436 ( .A(n2480), .B(n2481), .ZN(n2479) );
  XNOR2_X1 U2437 ( .A(n2482), .B(n2483), .ZN(n2377) );
  XOR2_X1 U2438 ( .A(n2484), .B(n2485), .Z(n2483) );
  NAND2_X1 U2439 ( .A1(a_6_), .A2(b_13_), .ZN(n2485) );
  XNOR2_X1 U2440 ( .A(n2486), .B(n2487), .ZN(n2381) );
  XOR2_X1 U2441 ( .A(n2488), .B(n2489), .Z(n2486) );
  XNOR2_X1 U2442 ( .A(n2490), .B(n2491), .ZN(n2384) );
  XNOR2_X1 U2443 ( .A(n2492), .B(n2493), .ZN(n2490) );
  NOR2_X1 U2444 ( .A1(n1990), .A2(n2119), .ZN(n2493) );
  XNOR2_X1 U2445 ( .A(n2494), .B(n2495), .ZN(n2388) );
  XNOR2_X1 U2446 ( .A(n2496), .B(n2497), .ZN(n2495) );
  XNOR2_X1 U2447 ( .A(n2498), .B(n2499), .ZN(n2393) );
  XNOR2_X1 U2448 ( .A(n2500), .B(n2501), .ZN(n2498) );
  XNOR2_X1 U2449 ( .A(n2502), .B(n2503), .ZN(n2397) );
  XNOR2_X1 U2450 ( .A(n2504), .B(n2505), .ZN(n2502) );
  NOR2_X1 U2451 ( .A1(n2396), .A2(n1990), .ZN(n2505) );
  XOR2_X1 U2452 ( .A(n2506), .B(n2507), .Z(n2234) );
  XNOR2_X1 U2453 ( .A(n2508), .B(n2509), .ZN(n2507) );
  OR2_X1 U2454 ( .A1(n2403), .A2(n2402), .ZN(n2290) );
  XOR2_X1 U2455 ( .A(n2510), .B(n2511), .Z(n2402) );
  XNOR2_X1 U2456 ( .A(n2512), .B(n2513), .ZN(n2510) );
  NOR2_X1 U2457 ( .A1(n2216), .A2(n2407), .ZN(n2513) );
  NAND2_X1 U2458 ( .A1(n2514), .A2(n2515), .ZN(n2403) );
  NAND2_X1 U2459 ( .A1(n2506), .A2(n2516), .ZN(n2515) );
  NAND2_X1 U2460 ( .A1(n2509), .A2(n2508), .ZN(n2516) );
  XNOR2_X1 U2461 ( .A(n2517), .B(n2518), .ZN(n2506) );
  XOR2_X1 U2462 ( .A(n2519), .B(n2520), .Z(n2517) );
  OR2_X1 U2463 ( .A1(n2508), .A2(n2509), .ZN(n2514) );
  NOR2_X1 U2464 ( .A1(n2407), .A2(n1990), .ZN(n2509) );
  NAND2_X1 U2465 ( .A1(n2521), .A2(n2522), .ZN(n2508) );
  NAND3_X1 U2466 ( .A1(a_1_), .A2(n2523), .A3(b_13_), .ZN(n2522) );
  NAND2_X1 U2467 ( .A1(n2504), .A2(n2503), .ZN(n2523) );
  OR2_X1 U2468 ( .A1(n2503), .A2(n2504), .ZN(n2521) );
  AND2_X1 U2469 ( .A1(n2524), .A2(n2525), .ZN(n2504) );
  NAND2_X1 U2470 ( .A1(n2501), .A2(n2526), .ZN(n2525) );
  NAND2_X1 U2471 ( .A1(n2500), .A2(n2499), .ZN(n2526) );
  NOR2_X1 U2472 ( .A1(n2220), .A2(n1990), .ZN(n2501) );
  OR2_X1 U2473 ( .A1(n2499), .A2(n2500), .ZN(n2524) );
  AND2_X1 U2474 ( .A1(n2527), .A2(n2528), .ZN(n2500) );
  NAND2_X1 U2475 ( .A1(n2497), .A2(n2529), .ZN(n2528) );
  OR2_X1 U2476 ( .A1(n2496), .A2(n2494), .ZN(n2529) );
  NOR2_X1 U2477 ( .A1(n2139), .A2(n1990), .ZN(n2497) );
  NAND2_X1 U2478 ( .A1(n2494), .A2(n2496), .ZN(n2527) );
  NAND2_X1 U2479 ( .A1(n2530), .A2(n2531), .ZN(n2496) );
  NAND3_X1 U2480 ( .A1(b_13_), .A2(n2532), .A3(a_4_), .ZN(n2531) );
  NAND2_X1 U2481 ( .A1(n2492), .A2(n2491), .ZN(n2532) );
  OR2_X1 U2482 ( .A1(n2491), .A2(n2492), .ZN(n2530) );
  AND2_X1 U2483 ( .A1(n2533), .A2(n2534), .ZN(n2492) );
  NAND2_X1 U2484 ( .A1(n2489), .A2(n2535), .ZN(n2534) );
  OR2_X1 U2485 ( .A1(n2487), .A2(n2488), .ZN(n2535) );
  NOR2_X1 U2486 ( .A1(n2104), .A2(n1990), .ZN(n2489) );
  NAND2_X1 U2487 ( .A1(n2487), .A2(n2488), .ZN(n2533) );
  NAND2_X1 U2488 ( .A1(n2536), .A2(n2537), .ZN(n2488) );
  NAND3_X1 U2489 ( .A1(b_13_), .A2(n2538), .A3(a_6_), .ZN(n2537) );
  OR2_X1 U2490 ( .A1(n2484), .A2(n2482), .ZN(n2538) );
  NAND2_X1 U2491 ( .A1(n2482), .A2(n2484), .ZN(n2536) );
  NAND2_X1 U2492 ( .A1(n2539), .A2(n2540), .ZN(n2484) );
  NAND2_X1 U2493 ( .A1(n2481), .A2(n2541), .ZN(n2540) );
  OR2_X1 U2494 ( .A1(n2480), .A2(n2478), .ZN(n2541) );
  NOR2_X1 U2495 ( .A1(n2076), .A2(n1990), .ZN(n2481) );
  NAND2_X1 U2496 ( .A1(n2478), .A2(n2480), .ZN(n2539) );
  NAND2_X1 U2497 ( .A1(n2542), .A2(n2543), .ZN(n2480) );
  NAND3_X1 U2498 ( .A1(b_13_), .A2(n2544), .A3(a_8_), .ZN(n2543) );
  OR2_X1 U2499 ( .A1(n2476), .A2(n2474), .ZN(n2544) );
  NAND2_X1 U2500 ( .A1(n2474), .A2(n2476), .ZN(n2542) );
  NAND2_X1 U2501 ( .A1(n2545), .A2(n2546), .ZN(n2476) );
  NAND2_X1 U2502 ( .A1(n2473), .A2(n2547), .ZN(n2546) );
  NAND2_X1 U2503 ( .A1(n2472), .A2(n2471), .ZN(n2547) );
  NOR2_X1 U2504 ( .A1(n2046), .A2(n1990), .ZN(n2473) );
  OR2_X1 U2505 ( .A1(n2471), .A2(n2472), .ZN(n2545) );
  AND2_X1 U2506 ( .A1(n2468), .A2(n2548), .ZN(n2472) );
  NAND2_X1 U2507 ( .A1(n2467), .A2(n2469), .ZN(n2548) );
  NAND2_X1 U2508 ( .A1(n2549), .A2(n2550), .ZN(n2469) );
  NAND2_X1 U2509 ( .A1(a_10_), .A2(b_13_), .ZN(n2550) );
  INV_X1 U2510 ( .A(n2551), .ZN(n2549) );
  XNOR2_X1 U2511 ( .A(n2552), .B(n2553), .ZN(n2467) );
  NAND2_X1 U2512 ( .A1(n2554), .A2(n2555), .ZN(n2552) );
  NAND2_X1 U2513 ( .A1(a_10_), .A2(n2551), .ZN(n2468) );
  NAND2_X1 U2514 ( .A1(n2441), .A2(n2556), .ZN(n2551) );
  NAND2_X1 U2515 ( .A1(n2440), .A2(n2442), .ZN(n2556) );
  NAND2_X1 U2516 ( .A1(n2557), .A2(n2558), .ZN(n2442) );
  NAND2_X1 U2517 ( .A1(a_11_), .A2(b_13_), .ZN(n2558) );
  INV_X1 U2518 ( .A(n2559), .ZN(n2557) );
  XOR2_X1 U2519 ( .A(n2560), .B(n2561), .Z(n2440) );
  XNOR2_X1 U2520 ( .A(n2562), .B(n2563), .ZN(n2560) );
  NAND2_X1 U2521 ( .A1(a_11_), .A2(n2559), .ZN(n2441) );
  NAND2_X1 U2522 ( .A1(n2564), .A2(n2565), .ZN(n2559) );
  NAND3_X1 U2523 ( .A1(b_13_), .A2(n2566), .A3(a_12_), .ZN(n2565) );
  NAND2_X1 U2524 ( .A1(n2450), .A2(n2448), .ZN(n2566) );
  OR2_X1 U2525 ( .A1(n2448), .A2(n2450), .ZN(n2564) );
  AND2_X1 U2526 ( .A1(n2567), .A2(n2568), .ZN(n2450) );
  NAND2_X1 U2527 ( .A1(n1985), .A2(n2569), .ZN(n2568) );
  OR2_X1 U2528 ( .A1(n2464), .A2(n2465), .ZN(n2569) );
  NOR2_X1 U2529 ( .A1(n1988), .A2(n1990), .ZN(n1985) );
  NAND2_X1 U2530 ( .A1(n2465), .A2(n2464), .ZN(n2567) );
  NAND2_X1 U2531 ( .A1(n2570), .A2(n2571), .ZN(n2464) );
  NAND2_X1 U2532 ( .A1(b_11_), .A2(n2572), .ZN(n2571) );
  NAND2_X1 U2533 ( .A1(n1964), .A2(n2573), .ZN(n2572) );
  NAND2_X1 U2534 ( .A1(a_15_), .A2(n2216), .ZN(n2573) );
  NAND2_X1 U2535 ( .A1(b_12_), .A2(n2574), .ZN(n2570) );
  NAND2_X1 U2536 ( .A1(n1967), .A2(n2575), .ZN(n2574) );
  NAND2_X1 U2537 ( .A1(a_14_), .A2(n2017), .ZN(n2575) );
  AND3_X1 U2538 ( .A1(b_12_), .A2(b_13_), .A3(n2215), .ZN(n2465) );
  XNOR2_X1 U2539 ( .A(n2576), .B(n2577), .ZN(n2448) );
  XOR2_X1 U2540 ( .A(n2578), .B(n2579), .Z(n2576) );
  XNOR2_X1 U2541 ( .A(n2580), .B(n2581), .ZN(n2471) );
  NOR2_X1 U2542 ( .A1(n2582), .A2(n2583), .ZN(n2581) );
  NOR2_X1 U2543 ( .A1(n2584), .A2(n2585), .ZN(n2582) );
  NOR2_X1 U2544 ( .A1(n2216), .A2(n2586), .ZN(n2584) );
  XOR2_X1 U2545 ( .A(n2587), .B(n2588), .Z(n2474) );
  XOR2_X1 U2546 ( .A(n2589), .B(n2590), .Z(n2587) );
  XOR2_X1 U2547 ( .A(n2591), .B(n2592), .Z(n2478) );
  XOR2_X1 U2548 ( .A(n2593), .B(n2594), .Z(n2591) );
  NOR2_X1 U2549 ( .A1(n2216), .A2(n2218), .ZN(n2594) );
  XNOR2_X1 U2550 ( .A(n2595), .B(n2596), .ZN(n2482) );
  XNOR2_X1 U2551 ( .A(n2597), .B(n2598), .ZN(n2596) );
  XNOR2_X1 U2552 ( .A(n2599), .B(n2600), .ZN(n2487) );
  XNOR2_X1 U2553 ( .A(n2601), .B(n2602), .ZN(n2599) );
  NOR2_X1 U2554 ( .A1(n2216), .A2(n2089), .ZN(n2602) );
  XNOR2_X1 U2555 ( .A(n2603), .B(n2604), .ZN(n2491) );
  XOR2_X1 U2556 ( .A(n2605), .B(n2606), .Z(n2603) );
  XOR2_X1 U2557 ( .A(n2607), .B(n2608), .Z(n2494) );
  XOR2_X1 U2558 ( .A(n2609), .B(n2610), .Z(n2607) );
  NOR2_X1 U2559 ( .A1(n2216), .A2(n2119), .ZN(n2610) );
  XOR2_X1 U2560 ( .A(n2611), .B(n2612), .Z(n2499) );
  XOR2_X1 U2561 ( .A(n2613), .B(n2614), .Z(n2612) );
  NAND2_X1 U2562 ( .A1(a_3_), .A2(b_12_), .ZN(n2614) );
  XNOR2_X1 U2563 ( .A(n2615), .B(n2616), .ZN(n2503) );
  XOR2_X1 U2564 ( .A(n2617), .B(n2618), .Z(n2615) );
  XOR2_X1 U2565 ( .A(n2275), .B(n2274), .Z(n2237) );
  XOR2_X1 U2566 ( .A(n2286), .B(n2619), .Z(n2274) );
  XNOR2_X1 U2567 ( .A(n2289), .B(n2288), .ZN(n2619) );
  NOR2_X1 U2568 ( .A1(n2407), .A2(n2017), .ZN(n2288) );
  NAND2_X1 U2569 ( .A1(n2620), .A2(n2621), .ZN(n2289) );
  NAND3_X1 U2570 ( .A1(a_1_), .A2(n2622), .A3(b_11_), .ZN(n2621) );
  OR2_X1 U2571 ( .A1(n2623), .A2(n2624), .ZN(n2622) );
  NAND2_X1 U2572 ( .A1(n2624), .A2(n2623), .ZN(n2620) );
  XOR2_X1 U2573 ( .A(n2625), .B(n2626), .Z(n2286) );
  XNOR2_X1 U2574 ( .A(n2627), .B(n2628), .ZN(n2626) );
  NAND2_X1 U2575 ( .A1(n2629), .A2(n2630), .ZN(n2275) );
  NAND3_X1 U2576 ( .A1(b_12_), .A2(n2631), .A3(a_0_), .ZN(n2630) );
  NAND2_X1 U2577 ( .A1(n2512), .A2(n2511), .ZN(n2631) );
  OR2_X1 U2578 ( .A1(n2511), .A2(n2512), .ZN(n2629) );
  AND2_X1 U2579 ( .A1(n2632), .A2(n2633), .ZN(n2512) );
  NAND2_X1 U2580 ( .A1(n2520), .A2(n2634), .ZN(n2633) );
  OR2_X1 U2581 ( .A1(n2519), .A2(n2518), .ZN(n2634) );
  NOR2_X1 U2582 ( .A1(n2216), .A2(n2396), .ZN(n2520) );
  NAND2_X1 U2583 ( .A1(n2518), .A2(n2519), .ZN(n2632) );
  NAND2_X1 U2584 ( .A1(n2635), .A2(n2636), .ZN(n2519) );
  NAND2_X1 U2585 ( .A1(n2618), .A2(n2637), .ZN(n2636) );
  OR2_X1 U2586 ( .A1(n2617), .A2(n2616), .ZN(n2637) );
  NOR2_X1 U2587 ( .A1(n2220), .A2(n2216), .ZN(n2618) );
  NAND2_X1 U2588 ( .A1(n2616), .A2(n2617), .ZN(n2635) );
  NAND2_X1 U2589 ( .A1(n2638), .A2(n2639), .ZN(n2617) );
  NAND3_X1 U2590 ( .A1(b_12_), .A2(n2640), .A3(a_3_), .ZN(n2639) );
  OR2_X1 U2591 ( .A1(n2613), .A2(n2611), .ZN(n2640) );
  NAND2_X1 U2592 ( .A1(n2611), .A2(n2613), .ZN(n2638) );
  NAND2_X1 U2593 ( .A1(n2641), .A2(n2642), .ZN(n2613) );
  NAND3_X1 U2594 ( .A1(b_12_), .A2(n2643), .A3(a_4_), .ZN(n2642) );
  OR2_X1 U2595 ( .A1(n2609), .A2(n2608), .ZN(n2643) );
  NAND2_X1 U2596 ( .A1(n2608), .A2(n2609), .ZN(n2641) );
  NAND2_X1 U2597 ( .A1(n2644), .A2(n2645), .ZN(n2609) );
  NAND2_X1 U2598 ( .A1(n2606), .A2(n2646), .ZN(n2645) );
  OR2_X1 U2599 ( .A1(n2605), .A2(n2604), .ZN(n2646) );
  NOR2_X1 U2600 ( .A1(n2104), .A2(n2216), .ZN(n2606) );
  NAND2_X1 U2601 ( .A1(n2604), .A2(n2605), .ZN(n2644) );
  NAND2_X1 U2602 ( .A1(n2647), .A2(n2648), .ZN(n2605) );
  NAND3_X1 U2603 ( .A1(b_12_), .A2(n2649), .A3(a_6_), .ZN(n2648) );
  NAND2_X1 U2604 ( .A1(n2601), .A2(n2600), .ZN(n2649) );
  OR2_X1 U2605 ( .A1(n2600), .A2(n2601), .ZN(n2647) );
  AND2_X1 U2606 ( .A1(n2650), .A2(n2651), .ZN(n2601) );
  NAND2_X1 U2607 ( .A1(n2598), .A2(n2652), .ZN(n2651) );
  OR2_X1 U2608 ( .A1(n2597), .A2(n2595), .ZN(n2652) );
  NOR2_X1 U2609 ( .A1(n2076), .A2(n2216), .ZN(n2598) );
  NAND2_X1 U2610 ( .A1(n2595), .A2(n2597), .ZN(n2650) );
  NAND2_X1 U2611 ( .A1(n2653), .A2(n2654), .ZN(n2597) );
  NAND3_X1 U2612 ( .A1(b_12_), .A2(n2655), .A3(a_8_), .ZN(n2654) );
  OR2_X1 U2613 ( .A1(n2593), .A2(n2592), .ZN(n2655) );
  NAND2_X1 U2614 ( .A1(n2592), .A2(n2593), .ZN(n2653) );
  NAND2_X1 U2615 ( .A1(n2656), .A2(n2657), .ZN(n2593) );
  NAND2_X1 U2616 ( .A1(n2590), .A2(n2658), .ZN(n2657) );
  OR2_X1 U2617 ( .A1(n2589), .A2(n2588), .ZN(n2658) );
  NOR2_X1 U2618 ( .A1(n2046), .A2(n2216), .ZN(n2590) );
  NAND2_X1 U2619 ( .A1(n2588), .A2(n2589), .ZN(n2656) );
  OR2_X1 U2620 ( .A1(n2583), .A2(n2659), .ZN(n2589) );
  AND2_X1 U2621 ( .A1(n2580), .A2(n2660), .ZN(n2659) );
  NAND2_X1 U2622 ( .A1(n2661), .A2(n2662), .ZN(n2660) );
  NAND2_X1 U2623 ( .A1(a_10_), .A2(b_12_), .ZN(n2662) );
  XOR2_X1 U2624 ( .A(n2663), .B(n2664), .Z(n2580) );
  XNOR2_X1 U2625 ( .A(n2665), .B(n2204), .ZN(n2663) );
  INV_X1 U2626 ( .A(n2015), .ZN(n2204) );
  NOR2_X1 U2627 ( .A1(n2586), .A2(n2661), .ZN(n2583) );
  INV_X1 U2628 ( .A(n2585), .ZN(n2661) );
  NAND2_X1 U2629 ( .A1(n2554), .A2(n2666), .ZN(n2585) );
  NAND2_X1 U2630 ( .A1(n2553), .A2(n2555), .ZN(n2666) );
  NAND2_X1 U2631 ( .A1(n2667), .A2(n2668), .ZN(n2555) );
  NAND2_X1 U2632 ( .A1(a_11_), .A2(b_12_), .ZN(n2668) );
  INV_X1 U2633 ( .A(n2669), .ZN(n2667) );
  XNOR2_X1 U2634 ( .A(n2670), .B(n2671), .ZN(n2553) );
  XOR2_X1 U2635 ( .A(n2672), .B(n2673), .Z(n2670) );
  NAND2_X1 U2636 ( .A1(b_11_), .A2(a_12_), .ZN(n2672) );
  NAND2_X1 U2637 ( .A1(a_11_), .A2(n2669), .ZN(n2554) );
  NAND2_X1 U2638 ( .A1(n2674), .A2(n2675), .ZN(n2669) );
  NAND2_X1 U2639 ( .A1(n2561), .A2(n2676), .ZN(n2675) );
  NAND2_X1 U2640 ( .A1(n2563), .A2(n2008), .ZN(n2676) );
  INV_X1 U2641 ( .A(n2562), .ZN(n2008) );
  INV_X1 U2642 ( .A(n2677), .ZN(n2563) );
  XOR2_X1 U2643 ( .A(n2678), .B(n2679), .Z(n2561) );
  XOR2_X1 U2644 ( .A(n2680), .B(n2681), .Z(n2678) );
  NAND2_X1 U2645 ( .A1(n2562), .A2(n2677), .ZN(n2674) );
  NAND2_X1 U2646 ( .A1(n2682), .A2(n2683), .ZN(n2677) );
  NAND2_X1 U2647 ( .A1(n2577), .A2(n2684), .ZN(n2683) );
  OR2_X1 U2648 ( .A1(n2578), .A2(n2579), .ZN(n2684) );
  NOR2_X1 U2649 ( .A1(n2216), .A2(n1988), .ZN(n2577) );
  NAND2_X1 U2650 ( .A1(n2579), .A2(n2578), .ZN(n2682) );
  NAND2_X1 U2651 ( .A1(n2685), .A2(n2686), .ZN(n2578) );
  NAND2_X1 U2652 ( .A1(b_10_), .A2(n2687), .ZN(n2686) );
  NAND2_X1 U2653 ( .A1(n1964), .A2(n2688), .ZN(n2687) );
  NAND2_X1 U2654 ( .A1(a_15_), .A2(n2017), .ZN(n2688) );
  NAND2_X1 U2655 ( .A1(b_11_), .A2(n2689), .ZN(n2685) );
  NAND2_X1 U2656 ( .A1(n1967), .A2(n2690), .ZN(n2689) );
  NAND2_X1 U2657 ( .A1(a_14_), .A2(n2691), .ZN(n2690) );
  AND3_X1 U2658 ( .A1(b_12_), .A2(b_11_), .A3(n2215), .ZN(n2579) );
  NOR2_X1 U2659 ( .A1(n2216), .A2(n2003), .ZN(n2562) );
  XNOR2_X1 U2660 ( .A(n2692), .B(n2693), .ZN(n2588) );
  NAND2_X1 U2661 ( .A1(n2694), .A2(n2695), .ZN(n2692) );
  XNOR2_X1 U2662 ( .A(n2696), .B(n2697), .ZN(n2592) );
  XNOR2_X1 U2663 ( .A(n2698), .B(n2699), .ZN(n2696) );
  XNOR2_X1 U2664 ( .A(n2700), .B(n2701), .ZN(n2595) );
  XNOR2_X1 U2665 ( .A(n2702), .B(n2703), .ZN(n2700) );
  NOR2_X1 U2666 ( .A1(n2017), .A2(n2218), .ZN(n2703) );
  XOR2_X1 U2667 ( .A(n2704), .B(n2705), .Z(n2600) );
  XNOR2_X1 U2668 ( .A(n2706), .B(n2707), .ZN(n2705) );
  XNOR2_X1 U2669 ( .A(n2708), .B(n2709), .ZN(n2604) );
  XOR2_X1 U2670 ( .A(n2710), .B(n2711), .Z(n2709) );
  NAND2_X1 U2671 ( .A1(a_6_), .A2(b_11_), .ZN(n2711) );
  XNOR2_X1 U2672 ( .A(n2712), .B(n2713), .ZN(n2608) );
  XNOR2_X1 U2673 ( .A(n2714), .B(n2715), .ZN(n2712) );
  XNOR2_X1 U2674 ( .A(n2716), .B(n2717), .ZN(n2611) );
  XNOR2_X1 U2675 ( .A(n2718), .B(n2719), .ZN(n2716) );
  XNOR2_X1 U2676 ( .A(n2720), .B(n2721), .ZN(n2616) );
  XOR2_X1 U2677 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND2_X1 U2678 ( .A1(a_3_), .A2(b_11_), .ZN(n2723) );
  XNOR2_X1 U2679 ( .A(n2724), .B(n2725), .ZN(n2518) );
  XOR2_X1 U2680 ( .A(n2726), .B(n2727), .Z(n2725) );
  NAND2_X1 U2681 ( .A1(a_2_), .A2(b_11_), .ZN(n2727) );
  XOR2_X1 U2682 ( .A(n2624), .B(n2728), .Z(n2511) );
  XOR2_X1 U2683 ( .A(n2623), .B(n2729), .Z(n2728) );
  NAND2_X1 U2684 ( .A1(b_11_), .A2(a_1_), .ZN(n2729) );
  NAND2_X1 U2685 ( .A1(n2730), .A2(n2731), .ZN(n2623) );
  NAND3_X1 U2686 ( .A1(b_11_), .A2(n2732), .A3(a_2_), .ZN(n2731) );
  OR2_X1 U2687 ( .A1(n2726), .A2(n2724), .ZN(n2732) );
  NAND2_X1 U2688 ( .A1(n2724), .A2(n2726), .ZN(n2730) );
  NAND2_X1 U2689 ( .A1(n2733), .A2(n2734), .ZN(n2726) );
  NAND3_X1 U2690 ( .A1(b_11_), .A2(n2735), .A3(a_3_), .ZN(n2734) );
  OR2_X1 U2691 ( .A1(n2722), .A2(n2720), .ZN(n2735) );
  NAND2_X1 U2692 ( .A1(n2720), .A2(n2722), .ZN(n2733) );
  NAND2_X1 U2693 ( .A1(n2736), .A2(n2737), .ZN(n2722) );
  NAND2_X1 U2694 ( .A1(n2719), .A2(n2738), .ZN(n2737) );
  NAND2_X1 U2695 ( .A1(n2718), .A2(n2717), .ZN(n2738) );
  NOR2_X1 U2696 ( .A1(n2119), .A2(n2017), .ZN(n2719) );
  OR2_X1 U2697 ( .A1(n2717), .A2(n2718), .ZN(n2736) );
  AND2_X1 U2698 ( .A1(n2739), .A2(n2740), .ZN(n2718) );
  NAND2_X1 U2699 ( .A1(n2715), .A2(n2741), .ZN(n2740) );
  NAND2_X1 U2700 ( .A1(n2714), .A2(n2713), .ZN(n2741) );
  NOR2_X1 U2701 ( .A1(n2104), .A2(n2017), .ZN(n2715) );
  OR2_X1 U2702 ( .A1(n2713), .A2(n2714), .ZN(n2739) );
  AND2_X1 U2703 ( .A1(n2742), .A2(n2743), .ZN(n2714) );
  NAND3_X1 U2704 ( .A1(b_11_), .A2(n2744), .A3(a_6_), .ZN(n2743) );
  OR2_X1 U2705 ( .A1(n2710), .A2(n2708), .ZN(n2744) );
  NAND2_X1 U2706 ( .A1(n2708), .A2(n2710), .ZN(n2742) );
  NAND2_X1 U2707 ( .A1(n2745), .A2(n2746), .ZN(n2710) );
  NAND2_X1 U2708 ( .A1(n2707), .A2(n2747), .ZN(n2746) );
  OR2_X1 U2709 ( .A1(n2706), .A2(n2704), .ZN(n2747) );
  NOR2_X1 U2710 ( .A1(n2076), .A2(n2017), .ZN(n2707) );
  NAND2_X1 U2711 ( .A1(n2704), .A2(n2706), .ZN(n2745) );
  NAND2_X1 U2712 ( .A1(n2748), .A2(n2749), .ZN(n2706) );
  NAND3_X1 U2713 ( .A1(b_11_), .A2(n2750), .A3(a_8_), .ZN(n2749) );
  NAND2_X1 U2714 ( .A1(n2702), .A2(n2701), .ZN(n2750) );
  OR2_X1 U2715 ( .A1(n2701), .A2(n2702), .ZN(n2748) );
  AND2_X1 U2716 ( .A1(n2751), .A2(n2752), .ZN(n2702) );
  NAND2_X1 U2717 ( .A1(n2699), .A2(n2753), .ZN(n2752) );
  NAND2_X1 U2718 ( .A1(n2698), .A2(n2697), .ZN(n2753) );
  NOR2_X1 U2719 ( .A1(n2046), .A2(n2017), .ZN(n2699) );
  OR2_X1 U2720 ( .A1(n2697), .A2(n2698), .ZN(n2751) );
  AND2_X1 U2721 ( .A1(n2694), .A2(n2754), .ZN(n2698) );
  NAND2_X1 U2722 ( .A1(n2693), .A2(n2695), .ZN(n2754) );
  NAND2_X1 U2723 ( .A1(n2755), .A2(n2756), .ZN(n2695) );
  NAND2_X1 U2724 ( .A1(a_10_), .A2(b_11_), .ZN(n2756) );
  INV_X1 U2725 ( .A(n2757), .ZN(n2755) );
  XNOR2_X1 U2726 ( .A(n2758), .B(n2759), .ZN(n2693) );
  NAND2_X1 U2727 ( .A1(n2760), .A2(n2761), .ZN(n2758) );
  NAND2_X1 U2728 ( .A1(a_10_), .A2(n2757), .ZN(n2694) );
  NAND2_X1 U2729 ( .A1(n2762), .A2(n2763), .ZN(n2757) );
  NAND2_X1 U2730 ( .A1(n2664), .A2(n2764), .ZN(n2763) );
  OR2_X1 U2731 ( .A1(n2665), .A2(n2015), .ZN(n2764) );
  XNOR2_X1 U2732 ( .A(n2765), .B(n2766), .ZN(n2664) );
  XOR2_X1 U2733 ( .A(n2767), .B(n2768), .Z(n2765) );
  NAND2_X1 U2734 ( .A1(b_10_), .A2(a_12_), .ZN(n2767) );
  NAND2_X1 U2735 ( .A1(n2015), .A2(n2665), .ZN(n2762) );
  NAND2_X1 U2736 ( .A1(n2769), .A2(n2770), .ZN(n2665) );
  NAND3_X1 U2737 ( .A1(a_12_), .A2(n2771), .A3(b_11_), .ZN(n2770) );
  NAND2_X1 U2738 ( .A1(n2673), .A2(n2671), .ZN(n2771) );
  OR2_X1 U2739 ( .A1(n2671), .A2(n2673), .ZN(n2769) );
  AND2_X1 U2740 ( .A1(n2772), .A2(n2773), .ZN(n2673) );
  NAND2_X1 U2741 ( .A1(n2679), .A2(n2774), .ZN(n2773) );
  OR2_X1 U2742 ( .A1(n2680), .A2(n2681), .ZN(n2774) );
  NOR2_X1 U2743 ( .A1(n2017), .A2(n1988), .ZN(n2679) );
  NAND2_X1 U2744 ( .A1(n2681), .A2(n2680), .ZN(n2772) );
  NAND2_X1 U2745 ( .A1(n2775), .A2(n2776), .ZN(n2680) );
  NAND2_X1 U2746 ( .A1(b_10_), .A2(n2777), .ZN(n2776) );
  NAND2_X1 U2747 ( .A1(n1967), .A2(n2778), .ZN(n2777) );
  NAND2_X1 U2748 ( .A1(a_14_), .A2(n2048), .ZN(n2778) );
  NAND2_X1 U2749 ( .A1(b_9_), .A2(n2779), .ZN(n2775) );
  NAND2_X1 U2750 ( .A1(n1964), .A2(n2780), .ZN(n2779) );
  NAND2_X1 U2751 ( .A1(a_15_), .A2(n2691), .ZN(n2780) );
  AND3_X1 U2752 ( .A1(b_10_), .A2(b_11_), .A3(n2215), .ZN(n2681) );
  XNOR2_X1 U2753 ( .A(n2781), .B(n2782), .ZN(n2671) );
  XOR2_X1 U2754 ( .A(n2783), .B(n2784), .Z(n2781) );
  NOR2_X1 U2755 ( .A1(n2019), .A2(n2017), .ZN(n2015) );
  XOR2_X1 U2756 ( .A(n2785), .B(n2786), .Z(n2697) );
  XNOR2_X1 U2757 ( .A(n2036), .B(n2787), .ZN(n2786) );
  XNOR2_X1 U2758 ( .A(n2788), .B(n2789), .ZN(n2701) );
  XOR2_X1 U2759 ( .A(n2790), .B(n2791), .Z(n2788) );
  XNOR2_X1 U2760 ( .A(n2792), .B(n2793), .ZN(n2704) );
  XNOR2_X1 U2761 ( .A(n2794), .B(n2795), .ZN(n2792) );
  NOR2_X1 U2762 ( .A1(n2691), .A2(n2218), .ZN(n2795) );
  XNOR2_X1 U2763 ( .A(n2796), .B(n2797), .ZN(n2708) );
  XNOR2_X1 U2764 ( .A(n2798), .B(n2799), .ZN(n2797) );
  XOR2_X1 U2765 ( .A(n2800), .B(n2801), .Z(n2713) );
  XOR2_X1 U2766 ( .A(n2802), .B(n2803), .Z(n2801) );
  NAND2_X1 U2767 ( .A1(a_6_), .A2(b_10_), .ZN(n2803) );
  XNOR2_X1 U2768 ( .A(n2804), .B(n2805), .ZN(n2717) );
  XOR2_X1 U2769 ( .A(n2806), .B(n2807), .Z(n2804) );
  NOR2_X1 U2770 ( .A1(n2691), .A2(n2104), .ZN(n2807) );
  XNOR2_X1 U2771 ( .A(n2808), .B(n2809), .ZN(n2720) );
  XNOR2_X1 U2772 ( .A(n2810), .B(n2811), .ZN(n2809) );
  XOR2_X1 U2773 ( .A(n2812), .B(n2813), .Z(n2724) );
  XOR2_X1 U2774 ( .A(n2814), .B(n2815), .Z(n2812) );
  XOR2_X1 U2775 ( .A(n2816), .B(n2817), .Z(n2624) );
  XOR2_X1 U2776 ( .A(n2818), .B(n2819), .Z(n2816) );
  NOR2_X1 U2777 ( .A1(n2691), .A2(n2220), .ZN(n2819) );
  NAND2_X1 U2778 ( .A1(n2820), .A2(n2821), .ZN(n1922) );
  NAND2_X1 U2779 ( .A1(n2271), .A2(n2272), .ZN(n2821) );
  XNOR2_X1 U2780 ( .A(n2822), .B(n2823), .ZN(n2820) );
  NAND3_X1 U2781 ( .A1(n2271), .A2(n2272), .A3(n2824), .ZN(n1921) );
  XNOR2_X1 U2782 ( .A(n2822), .B(n2825), .ZN(n2824) );
  INV_X1 U2783 ( .A(n2823), .ZN(n2825) );
  NAND2_X1 U2784 ( .A1(n2282), .A2(n2826), .ZN(n2272) );
  NAND2_X1 U2785 ( .A1(n2281), .A2(n2283), .ZN(n2826) );
  NAND2_X1 U2786 ( .A1(n2827), .A2(n2828), .ZN(n2283) );
  NAND2_X1 U2787 ( .A1(a_0_), .A2(b_10_), .ZN(n2828) );
  INV_X1 U2788 ( .A(n2829), .ZN(n2827) );
  XNOR2_X1 U2789 ( .A(n2830), .B(n2831), .ZN(n2281) );
  XOR2_X1 U2790 ( .A(n2832), .B(n2833), .Z(n2831) );
  NAND2_X1 U2791 ( .A1(b_9_), .A2(a_1_), .ZN(n2833) );
  NAND2_X1 U2792 ( .A1(a_0_), .A2(n2829), .ZN(n2282) );
  NAND2_X1 U2793 ( .A1(n2834), .A2(n2835), .ZN(n2829) );
  NAND2_X1 U2794 ( .A1(n2628), .A2(n2836), .ZN(n2835) );
  OR2_X1 U2795 ( .A1(n2625), .A2(n2627), .ZN(n2836) );
  NOR2_X1 U2796 ( .A1(n2691), .A2(n2396), .ZN(n2628) );
  NAND2_X1 U2797 ( .A1(n2625), .A2(n2627), .ZN(n2834) );
  NAND2_X1 U2798 ( .A1(n2837), .A2(n2838), .ZN(n2627) );
  NAND3_X1 U2799 ( .A1(b_10_), .A2(n2839), .A3(a_2_), .ZN(n2838) );
  OR2_X1 U2800 ( .A1(n2818), .A2(n2817), .ZN(n2839) );
  NAND2_X1 U2801 ( .A1(n2817), .A2(n2818), .ZN(n2837) );
  NAND2_X1 U2802 ( .A1(n2840), .A2(n2841), .ZN(n2818) );
  NAND2_X1 U2803 ( .A1(n2815), .A2(n2842), .ZN(n2841) );
  OR2_X1 U2804 ( .A1(n2813), .A2(n2814), .ZN(n2842) );
  NOR2_X1 U2805 ( .A1(n2139), .A2(n2691), .ZN(n2815) );
  NAND2_X1 U2806 ( .A1(n2813), .A2(n2814), .ZN(n2840) );
  NAND2_X1 U2807 ( .A1(n2843), .A2(n2844), .ZN(n2814) );
  NAND2_X1 U2808 ( .A1(n2811), .A2(n2845), .ZN(n2844) );
  OR2_X1 U2809 ( .A1(n2808), .A2(n2810), .ZN(n2845) );
  NOR2_X1 U2810 ( .A1(n2119), .A2(n2691), .ZN(n2811) );
  NAND2_X1 U2811 ( .A1(n2808), .A2(n2810), .ZN(n2843) );
  NAND2_X1 U2812 ( .A1(n2846), .A2(n2847), .ZN(n2810) );
  NAND3_X1 U2813 ( .A1(b_10_), .A2(n2848), .A3(a_5_), .ZN(n2847) );
  OR2_X1 U2814 ( .A1(n2805), .A2(n2806), .ZN(n2848) );
  NAND2_X1 U2815 ( .A1(n2805), .A2(n2806), .ZN(n2846) );
  NAND2_X1 U2816 ( .A1(n2849), .A2(n2850), .ZN(n2806) );
  NAND3_X1 U2817 ( .A1(b_10_), .A2(n2851), .A3(a_6_), .ZN(n2850) );
  OR2_X1 U2818 ( .A1(n2800), .A2(n2802), .ZN(n2851) );
  NAND2_X1 U2819 ( .A1(n2800), .A2(n2802), .ZN(n2849) );
  NAND2_X1 U2820 ( .A1(n2852), .A2(n2853), .ZN(n2802) );
  NAND2_X1 U2821 ( .A1(n2799), .A2(n2854), .ZN(n2853) );
  OR2_X1 U2822 ( .A1(n2796), .A2(n2798), .ZN(n2854) );
  NOR2_X1 U2823 ( .A1(n2076), .A2(n2691), .ZN(n2799) );
  NAND2_X1 U2824 ( .A1(n2796), .A2(n2798), .ZN(n2852) );
  NAND2_X1 U2825 ( .A1(n2855), .A2(n2856), .ZN(n2798) );
  NAND3_X1 U2826 ( .A1(b_10_), .A2(n2857), .A3(a_8_), .ZN(n2856) );
  NAND2_X1 U2827 ( .A1(n2794), .A2(n2793), .ZN(n2857) );
  OR2_X1 U2828 ( .A1(n2793), .A2(n2794), .ZN(n2855) );
  AND2_X1 U2829 ( .A1(n2858), .A2(n2859), .ZN(n2794) );
  NAND2_X1 U2830 ( .A1(n2791), .A2(n2860), .ZN(n2859) );
  OR2_X1 U2831 ( .A1(n2789), .A2(n2790), .ZN(n2860) );
  NOR2_X1 U2832 ( .A1(n2046), .A2(n2691), .ZN(n2791) );
  NAND2_X1 U2833 ( .A1(n2789), .A2(n2790), .ZN(n2858) );
  NAND2_X1 U2834 ( .A1(n2861), .A2(n2862), .ZN(n2790) );
  NAND2_X1 U2835 ( .A1(n2785), .A2(n2863), .ZN(n2862) );
  OR2_X1 U2836 ( .A1(n2787), .A2(n2036), .ZN(n2863) );
  XNOR2_X1 U2837 ( .A(n2864), .B(n2865), .ZN(n2785) );
  NAND2_X1 U2838 ( .A1(n2866), .A2(n2867), .ZN(n2864) );
  NAND2_X1 U2839 ( .A1(n2036), .A2(n2787), .ZN(n2861) );
  NAND2_X1 U2840 ( .A1(n2760), .A2(n2868), .ZN(n2787) );
  NAND2_X1 U2841 ( .A1(n2759), .A2(n2761), .ZN(n2868) );
  NAND2_X1 U2842 ( .A1(n2869), .A2(n2870), .ZN(n2761) );
  NAND2_X1 U2843 ( .A1(b_10_), .A2(a_11_), .ZN(n2870) );
  INV_X1 U2844 ( .A(n2871), .ZN(n2869) );
  XNOR2_X1 U2845 ( .A(n2872), .B(n2873), .ZN(n2759) );
  XOR2_X1 U2846 ( .A(n2874), .B(n2875), .Z(n2872) );
  NAND2_X1 U2847 ( .A1(b_9_), .A2(a_12_), .ZN(n2874) );
  NAND2_X1 U2848 ( .A1(a_11_), .A2(n2871), .ZN(n2760) );
  NAND2_X1 U2849 ( .A1(n2876), .A2(n2877), .ZN(n2871) );
  NAND3_X1 U2850 ( .A1(a_12_), .A2(n2878), .A3(b_10_), .ZN(n2877) );
  NAND2_X1 U2851 ( .A1(n2768), .A2(n2766), .ZN(n2878) );
  OR2_X1 U2852 ( .A1(n2766), .A2(n2768), .ZN(n2876) );
  AND2_X1 U2853 ( .A1(n2879), .A2(n2880), .ZN(n2768) );
  NAND2_X1 U2854 ( .A1(n2782), .A2(n2881), .ZN(n2880) );
  OR2_X1 U2855 ( .A1(n2783), .A2(n2784), .ZN(n2881) );
  NOR2_X1 U2856 ( .A1(n2691), .A2(n1988), .ZN(n2782) );
  NAND2_X1 U2857 ( .A1(n2784), .A2(n2783), .ZN(n2879) );
  NAND2_X1 U2858 ( .A1(n2882), .A2(n2883), .ZN(n2783) );
  NAND2_X1 U2859 ( .A1(b_8_), .A2(n2884), .ZN(n2883) );
  NAND2_X1 U2860 ( .A1(n1964), .A2(n2885), .ZN(n2884) );
  NAND2_X1 U2861 ( .A1(a_15_), .A2(n2048), .ZN(n2885) );
  NAND2_X1 U2862 ( .A1(b_9_), .A2(n2886), .ZN(n2882) );
  NAND2_X1 U2863 ( .A1(n1967), .A2(n2887), .ZN(n2886) );
  NAND2_X1 U2864 ( .A1(a_14_), .A2(n2217), .ZN(n2887) );
  AND3_X1 U2865 ( .A1(b_9_), .A2(b_10_), .A3(n2215), .ZN(n2784) );
  XNOR2_X1 U2866 ( .A(n2888), .B(n2889), .ZN(n2766) );
  XOR2_X1 U2867 ( .A(n2890), .B(n2891), .Z(n2888) );
  NOR2_X1 U2868 ( .A1(n2691), .A2(n2586), .ZN(n2036) );
  XNOR2_X1 U2869 ( .A(n2892), .B(n2893), .ZN(n2789) );
  NAND2_X1 U2870 ( .A1(n2894), .A2(n2895), .ZN(n2892) );
  XNOR2_X1 U2871 ( .A(n2896), .B(n2897), .ZN(n2793) );
  XNOR2_X1 U2872 ( .A(n2898), .B(n2200), .ZN(n2896) );
  INV_X1 U2873 ( .A(n2043), .ZN(n2200) );
  XNOR2_X1 U2874 ( .A(n2899), .B(n2900), .ZN(n2796) );
  XNOR2_X1 U2875 ( .A(n2901), .B(n2902), .ZN(n2899) );
  NOR2_X1 U2876 ( .A1(n2048), .A2(n2218), .ZN(n2902) );
  XNOR2_X1 U2877 ( .A(n2903), .B(n2904), .ZN(n2800) );
  XNOR2_X1 U2878 ( .A(n2905), .B(n2906), .ZN(n2904) );
  XNOR2_X1 U2879 ( .A(n2907), .B(n2908), .ZN(n2805) );
  XNOR2_X1 U2880 ( .A(n2909), .B(n2910), .ZN(n2908) );
  XNOR2_X1 U2881 ( .A(n2911), .B(n2912), .ZN(n2808) );
  XOR2_X1 U2882 ( .A(n2913), .B(n2914), .Z(n2912) );
  NAND2_X1 U2883 ( .A1(a_5_), .A2(b_9_), .ZN(n2914) );
  XNOR2_X1 U2884 ( .A(n2915), .B(n2916), .ZN(n2813) );
  NAND2_X1 U2885 ( .A1(n2917), .A2(n2918), .ZN(n2915) );
  XOR2_X1 U2886 ( .A(n2919), .B(n2920), .Z(n2817) );
  XNOR2_X1 U2887 ( .A(n2921), .B(n2922), .ZN(n2919) );
  NAND2_X1 U2888 ( .A1(a_3_), .A2(b_9_), .ZN(n2921) );
  XOR2_X1 U2889 ( .A(n2923), .B(n2924), .Z(n2625) );
  XNOR2_X1 U2890 ( .A(n2925), .B(n2926), .ZN(n2924) );
  NAND2_X1 U2891 ( .A1(a_2_), .A2(b_9_), .ZN(n2926) );
  XOR2_X1 U2892 ( .A(n2927), .B(n2928), .Z(n2271) );
  XOR2_X1 U2893 ( .A(n2929), .B(n2930), .Z(n2927) );
  NOR2_X1 U2894 ( .A1(n2048), .A2(n2407), .ZN(n2930) );
  NAND2_X1 U2895 ( .A1(n2931), .A2(n2932), .ZN(n1927) );
  NAND2_X1 U2896 ( .A1(n2823), .A2(n2822), .ZN(n2932) );
  XNOR2_X1 U2897 ( .A(n2933), .B(n2934), .ZN(n2931) );
  NAND3_X1 U2898 ( .A1(n2823), .A2(n2822), .A3(n2935), .ZN(n1926) );
  XOR2_X1 U2899 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND2_X1 U2900 ( .A1(n2936), .A2(n2937), .ZN(n2822) );
  NAND3_X1 U2901 ( .A1(b_9_), .A2(n2938), .A3(a_0_), .ZN(n2937) );
  OR2_X1 U2902 ( .A1(n2928), .A2(n2929), .ZN(n2938) );
  NAND2_X1 U2903 ( .A1(n2928), .A2(n2929), .ZN(n2936) );
  NAND2_X1 U2904 ( .A1(n2939), .A2(n2940), .ZN(n2929) );
  NAND3_X1 U2905 ( .A1(a_1_), .A2(n2941), .A3(b_9_), .ZN(n2940) );
  OR2_X1 U2906 ( .A1(n2830), .A2(n2832), .ZN(n2941) );
  NAND2_X1 U2907 ( .A1(n2830), .A2(n2832), .ZN(n2939) );
  NAND2_X1 U2908 ( .A1(n2942), .A2(n2943), .ZN(n2832) );
  NAND3_X1 U2909 ( .A1(b_9_), .A2(n2944), .A3(a_2_), .ZN(n2943) );
  NAND2_X1 U2910 ( .A1(n2925), .A2(n2923), .ZN(n2944) );
  OR2_X1 U2911 ( .A1(n2923), .A2(n2925), .ZN(n2942) );
  AND2_X1 U2912 ( .A1(n2945), .A2(n2946), .ZN(n2925) );
  NAND3_X1 U2913 ( .A1(b_9_), .A2(n2947), .A3(a_3_), .ZN(n2946) );
  OR2_X1 U2914 ( .A1(n2920), .A2(n2922), .ZN(n2947) );
  NAND2_X1 U2915 ( .A1(n2920), .A2(n2922), .ZN(n2945) );
  NAND2_X1 U2916 ( .A1(n2917), .A2(n2948), .ZN(n2922) );
  NAND2_X1 U2917 ( .A1(n2916), .A2(n2918), .ZN(n2948) );
  NAND2_X1 U2918 ( .A1(n2949), .A2(n2950), .ZN(n2918) );
  NAND2_X1 U2919 ( .A1(a_4_), .A2(b_9_), .ZN(n2950) );
  INV_X1 U2920 ( .A(n2951), .ZN(n2949) );
  XNOR2_X1 U2921 ( .A(n2952), .B(n2953), .ZN(n2916) );
  XNOR2_X1 U2922 ( .A(n2954), .B(n2955), .ZN(n2952) );
  NOR2_X1 U2923 ( .A1(n2217), .A2(n2104), .ZN(n2955) );
  NAND2_X1 U2924 ( .A1(a_4_), .A2(n2951), .ZN(n2917) );
  NAND2_X1 U2925 ( .A1(n2956), .A2(n2957), .ZN(n2951) );
  NAND3_X1 U2926 ( .A1(b_9_), .A2(n2958), .A3(a_5_), .ZN(n2957) );
  OR2_X1 U2927 ( .A1(n2913), .A2(n2911), .ZN(n2958) );
  NAND2_X1 U2928 ( .A1(n2911), .A2(n2913), .ZN(n2956) );
  NAND2_X1 U2929 ( .A1(n2959), .A2(n2960), .ZN(n2913) );
  NAND2_X1 U2930 ( .A1(n2910), .A2(n2961), .ZN(n2960) );
  OR2_X1 U2931 ( .A1(n2909), .A2(n2907), .ZN(n2961) );
  NOR2_X1 U2932 ( .A1(n2089), .A2(n2048), .ZN(n2910) );
  NAND2_X1 U2933 ( .A1(n2907), .A2(n2909), .ZN(n2959) );
  NAND2_X1 U2934 ( .A1(n2962), .A2(n2963), .ZN(n2909) );
  NAND2_X1 U2935 ( .A1(n2906), .A2(n2964), .ZN(n2963) );
  OR2_X1 U2936 ( .A1(n2905), .A2(n2903), .ZN(n2964) );
  NOR2_X1 U2937 ( .A1(n2076), .A2(n2048), .ZN(n2906) );
  NAND2_X1 U2938 ( .A1(n2903), .A2(n2905), .ZN(n2962) );
  NAND2_X1 U2939 ( .A1(n2965), .A2(n2966), .ZN(n2905) );
  NAND3_X1 U2940 ( .A1(b_9_), .A2(n2967), .A3(a_8_), .ZN(n2966) );
  NAND2_X1 U2941 ( .A1(n2901), .A2(n2900), .ZN(n2967) );
  OR2_X1 U2942 ( .A1(n2900), .A2(n2901), .ZN(n2965) );
  AND2_X1 U2943 ( .A1(n2968), .A2(n2969), .ZN(n2901) );
  NAND2_X1 U2944 ( .A1(n2043), .A2(n2970), .ZN(n2969) );
  OR2_X1 U2945 ( .A1(n2897), .A2(n2898), .ZN(n2970) );
  NOR2_X1 U2946 ( .A1(n2046), .A2(n2048), .ZN(n2043) );
  NAND2_X1 U2947 ( .A1(n2897), .A2(n2898), .ZN(n2968) );
  NAND2_X1 U2948 ( .A1(n2894), .A2(n2971), .ZN(n2898) );
  NAND2_X1 U2949 ( .A1(n2893), .A2(n2895), .ZN(n2971) );
  NAND2_X1 U2950 ( .A1(n2972), .A2(n2973), .ZN(n2895) );
  NAND2_X1 U2951 ( .A1(b_9_), .A2(a_10_), .ZN(n2973) );
  INV_X1 U2952 ( .A(n2974), .ZN(n2972) );
  XNOR2_X1 U2953 ( .A(n2975), .B(n2976), .ZN(n2893) );
  NAND2_X1 U2954 ( .A1(n2977), .A2(n2978), .ZN(n2975) );
  NAND2_X1 U2955 ( .A1(a_10_), .A2(n2974), .ZN(n2894) );
  NAND2_X1 U2956 ( .A1(n2866), .A2(n2979), .ZN(n2974) );
  NAND2_X1 U2957 ( .A1(n2865), .A2(n2867), .ZN(n2979) );
  NAND2_X1 U2958 ( .A1(n2980), .A2(n2981), .ZN(n2867) );
  NAND2_X1 U2959 ( .A1(b_9_), .A2(a_11_), .ZN(n2981) );
  INV_X1 U2960 ( .A(n2982), .ZN(n2980) );
  XNOR2_X1 U2961 ( .A(n2983), .B(n2984), .ZN(n2865) );
  XOR2_X1 U2962 ( .A(n2985), .B(n2986), .Z(n2983) );
  NAND2_X1 U2963 ( .A1(b_8_), .A2(a_12_), .ZN(n2985) );
  NAND2_X1 U2964 ( .A1(a_11_), .A2(n2982), .ZN(n2866) );
  NAND2_X1 U2965 ( .A1(n2987), .A2(n2988), .ZN(n2982) );
  NAND3_X1 U2966 ( .A1(a_12_), .A2(n2989), .A3(b_9_), .ZN(n2988) );
  NAND2_X1 U2967 ( .A1(n2875), .A2(n2873), .ZN(n2989) );
  OR2_X1 U2968 ( .A1(n2873), .A2(n2875), .ZN(n2987) );
  AND2_X1 U2969 ( .A1(n2990), .A2(n2991), .ZN(n2875) );
  NAND2_X1 U2970 ( .A1(n2889), .A2(n2992), .ZN(n2991) );
  OR2_X1 U2971 ( .A1(n2890), .A2(n2891), .ZN(n2992) );
  NOR2_X1 U2972 ( .A1(n2048), .A2(n1988), .ZN(n2889) );
  NAND2_X1 U2973 ( .A1(n2891), .A2(n2890), .ZN(n2990) );
  NAND2_X1 U2974 ( .A1(n2993), .A2(n2994), .ZN(n2890) );
  NAND2_X1 U2975 ( .A1(b_7_), .A2(n2995), .ZN(n2994) );
  NAND2_X1 U2976 ( .A1(n1964), .A2(n2996), .ZN(n2995) );
  NAND2_X1 U2977 ( .A1(a_15_), .A2(n2217), .ZN(n2996) );
  NAND2_X1 U2978 ( .A1(b_8_), .A2(n2997), .ZN(n2993) );
  NAND2_X1 U2979 ( .A1(n1967), .A2(n2998), .ZN(n2997) );
  NAND2_X1 U2980 ( .A1(a_14_), .A2(n2074), .ZN(n2998) );
  AND3_X1 U2981 ( .A1(b_8_), .A2(b_9_), .A3(n2215), .ZN(n2891) );
  XNOR2_X1 U2982 ( .A(n2999), .B(n3000), .ZN(n2873) );
  XOR2_X1 U2983 ( .A(n3001), .B(n3002), .Z(n2999) );
  XNOR2_X1 U2984 ( .A(n3003), .B(n3004), .ZN(n2897) );
  NAND2_X1 U2985 ( .A1(n3005), .A2(n3006), .ZN(n3003) );
  XNOR2_X1 U2986 ( .A(n3007), .B(n3008), .ZN(n2900) );
  XOR2_X1 U2987 ( .A(n3009), .B(n3010), .Z(n3007) );
  XOR2_X1 U2988 ( .A(n3011), .B(n3012), .Z(n2903) );
  XNOR2_X1 U2989 ( .A(n3013), .B(n2065), .ZN(n3011) );
  INV_X1 U2990 ( .A(n3014), .ZN(n2065) );
  XOR2_X1 U2991 ( .A(n3015), .B(n3016), .Z(n2907) );
  XOR2_X1 U2992 ( .A(n3017), .B(n3018), .Z(n3015) );
  NOR2_X1 U2993 ( .A1(n2217), .A2(n2076), .ZN(n3018) );
  XNOR2_X1 U2994 ( .A(n3019), .B(n3020), .ZN(n2911) );
  XOR2_X1 U2995 ( .A(n3021), .B(n3022), .Z(n3020) );
  NAND2_X1 U2996 ( .A1(a_6_), .A2(b_8_), .ZN(n3022) );
  XOR2_X1 U2997 ( .A(n3023), .B(n3024), .Z(n2920) );
  XNOR2_X1 U2998 ( .A(n3025), .B(n3026), .ZN(n3024) );
  NAND2_X1 U2999 ( .A1(a_4_), .A2(b_8_), .ZN(n3026) );
  XNOR2_X1 U3000 ( .A(n3027), .B(n3028), .ZN(n2923) );
  XOR2_X1 U3001 ( .A(n3029), .B(n3030), .Z(n3027) );
  NOR2_X1 U3002 ( .A1(n2217), .A2(n2139), .ZN(n3030) );
  XOR2_X1 U3003 ( .A(n3031), .B(n3032), .Z(n2830) );
  XOR2_X1 U3004 ( .A(n3033), .B(n3034), .Z(n3032) );
  XNOR2_X1 U3005 ( .A(n3035), .B(n3036), .ZN(n2928) );
  NAND2_X1 U3006 ( .A1(n3037), .A2(n3038), .ZN(n3035) );
  XNOR2_X1 U3007 ( .A(n3039), .B(n3040), .ZN(n2823) );
  NAND2_X1 U3008 ( .A1(n3041), .A2(n3042), .ZN(n3039) );
  NAND2_X1 U3009 ( .A1(n3043), .A2(n3044), .ZN(n1932) );
  NAND2_X1 U3010 ( .A1(n2933), .A2(n2934), .ZN(n3044) );
  XNOR2_X1 U3011 ( .A(n3045), .B(n3046), .ZN(n3043) );
  NAND3_X1 U3012 ( .A1(n3047), .A2(n2934), .A3(n2933), .ZN(n1931) );
  XNOR2_X1 U3013 ( .A(n3048), .B(n3049), .ZN(n2933) );
  XOR2_X1 U3014 ( .A(n3050), .B(n3051), .Z(n3049) );
  NAND2_X1 U3015 ( .A1(a_0_), .A2(b_7_), .ZN(n3051) );
  NAND2_X1 U3016 ( .A1(n3041), .A2(n3052), .ZN(n2934) );
  NAND2_X1 U3017 ( .A1(n3040), .A2(n3042), .ZN(n3052) );
  NAND2_X1 U3018 ( .A1(n3053), .A2(n3054), .ZN(n3042) );
  NAND2_X1 U3019 ( .A1(a_0_), .A2(b_8_), .ZN(n3054) );
  INV_X1 U3020 ( .A(n3055), .ZN(n3053) );
  XNOR2_X1 U3021 ( .A(n3056), .B(n3057), .ZN(n3040) );
  XOR2_X1 U3022 ( .A(n3058), .B(n3059), .Z(n3056) );
  NAND2_X1 U3023 ( .A1(b_7_), .A2(a_1_), .ZN(n3058) );
  NAND2_X1 U3024 ( .A1(a_0_), .A2(n3055), .ZN(n3041) );
  NAND2_X1 U3025 ( .A1(n3037), .A2(n3060), .ZN(n3055) );
  NAND2_X1 U3026 ( .A1(n3036), .A2(n3038), .ZN(n3060) );
  NAND2_X1 U3027 ( .A1(n3061), .A2(n3062), .ZN(n3038) );
  NAND2_X1 U3028 ( .A1(b_8_), .A2(a_1_), .ZN(n3062) );
  INV_X1 U3029 ( .A(n3063), .ZN(n3061) );
  XNOR2_X1 U3030 ( .A(n3064), .B(n3065), .ZN(n3036) );
  XNOR2_X1 U3031 ( .A(n3066), .B(n3067), .ZN(n3064) );
  NAND2_X1 U3032 ( .A1(a_1_), .A2(n3063), .ZN(n3037) );
  NAND2_X1 U3033 ( .A1(n3068), .A2(n3069), .ZN(n3063) );
  NAND2_X1 U3034 ( .A1(n3034), .A2(n3070), .ZN(n3069) );
  NAND2_X1 U3035 ( .A1(n3033), .A2(n3031), .ZN(n3070) );
  NOR2_X1 U3036 ( .A1(n2220), .A2(n2217), .ZN(n3034) );
  OR2_X1 U3037 ( .A1(n3031), .A2(n3033), .ZN(n3068) );
  AND2_X1 U3038 ( .A1(n3071), .A2(n3072), .ZN(n3033) );
  NAND3_X1 U3039 ( .A1(b_8_), .A2(n3073), .A3(a_3_), .ZN(n3072) );
  OR2_X1 U3040 ( .A1(n3028), .A2(n3029), .ZN(n3073) );
  NAND2_X1 U3041 ( .A1(n3028), .A2(n3029), .ZN(n3071) );
  NAND2_X1 U3042 ( .A1(n3074), .A2(n3075), .ZN(n3029) );
  NAND3_X1 U3043 ( .A1(b_8_), .A2(n3076), .A3(a_4_), .ZN(n3075) );
  NAND2_X1 U3044 ( .A1(n3025), .A2(n3023), .ZN(n3076) );
  OR2_X1 U3045 ( .A1(n3023), .A2(n3025), .ZN(n3074) );
  AND2_X1 U3046 ( .A1(n3077), .A2(n3078), .ZN(n3025) );
  NAND3_X1 U3047 ( .A1(b_8_), .A2(n3079), .A3(a_5_), .ZN(n3078) );
  NAND2_X1 U3048 ( .A1(n2954), .A2(n2953), .ZN(n3079) );
  OR2_X1 U3049 ( .A1(n2953), .A2(n2954), .ZN(n3077) );
  AND2_X1 U3050 ( .A1(n3080), .A2(n3081), .ZN(n2954) );
  NAND3_X1 U3051 ( .A1(b_8_), .A2(n3082), .A3(a_6_), .ZN(n3081) );
  OR2_X1 U3052 ( .A1(n3019), .A2(n3021), .ZN(n3082) );
  NAND2_X1 U3053 ( .A1(n3019), .A2(n3021), .ZN(n3080) );
  NAND2_X1 U3054 ( .A1(n3083), .A2(n3084), .ZN(n3021) );
  NAND3_X1 U3055 ( .A1(b_8_), .A2(n3085), .A3(a_7_), .ZN(n3084) );
  OR2_X1 U3056 ( .A1(n3016), .A2(n3017), .ZN(n3085) );
  NAND2_X1 U3057 ( .A1(n3016), .A2(n3017), .ZN(n3083) );
  NAND2_X1 U3058 ( .A1(n3086), .A2(n3087), .ZN(n3017) );
  NAND2_X1 U3059 ( .A1(n3012), .A2(n3088), .ZN(n3087) );
  OR2_X1 U3060 ( .A1(n3013), .A2(n3014), .ZN(n3088) );
  XNOR2_X1 U3061 ( .A(n3089), .B(n3090), .ZN(n3012) );
  XNOR2_X1 U3062 ( .A(n3091), .B(n3092), .ZN(n3089) );
  NAND2_X1 U3063 ( .A1(n3014), .A2(n3013), .ZN(n3086) );
  NAND2_X1 U3064 ( .A1(n3093), .A2(n3094), .ZN(n3013) );
  NAND2_X1 U3065 ( .A1(n3010), .A2(n3095), .ZN(n3094) );
  OR2_X1 U3066 ( .A1(n3008), .A2(n3009), .ZN(n3095) );
  NOR2_X1 U3067 ( .A1(n2217), .A2(n2046), .ZN(n3010) );
  NAND2_X1 U3068 ( .A1(n3008), .A2(n3009), .ZN(n3093) );
  NAND2_X1 U3069 ( .A1(n3005), .A2(n3096), .ZN(n3009) );
  NAND2_X1 U3070 ( .A1(n3004), .A2(n3006), .ZN(n3096) );
  NAND2_X1 U3071 ( .A1(n3097), .A2(n3098), .ZN(n3006) );
  NAND2_X1 U3072 ( .A1(b_8_), .A2(a_10_), .ZN(n3098) );
  INV_X1 U3073 ( .A(n3099), .ZN(n3097) );
  XNOR2_X1 U3074 ( .A(n3100), .B(n3101), .ZN(n3004) );
  NAND2_X1 U3075 ( .A1(n3102), .A2(n3103), .ZN(n3100) );
  NAND2_X1 U3076 ( .A1(a_10_), .A2(n3099), .ZN(n3005) );
  NAND2_X1 U3077 ( .A1(n2977), .A2(n3104), .ZN(n3099) );
  NAND2_X1 U3078 ( .A1(n2976), .A2(n2978), .ZN(n3104) );
  NAND2_X1 U3079 ( .A1(n3105), .A2(n3106), .ZN(n2978) );
  NAND2_X1 U3080 ( .A1(b_8_), .A2(a_11_), .ZN(n3106) );
  INV_X1 U3081 ( .A(n3107), .ZN(n3105) );
  XNOR2_X1 U3082 ( .A(n3108), .B(n3109), .ZN(n2976) );
  XOR2_X1 U3083 ( .A(n3110), .B(n3111), .Z(n3108) );
  NAND2_X1 U3084 ( .A1(b_7_), .A2(a_12_), .ZN(n3110) );
  NAND2_X1 U3085 ( .A1(a_11_), .A2(n3107), .ZN(n2977) );
  NAND2_X1 U3086 ( .A1(n3112), .A2(n3113), .ZN(n3107) );
  NAND3_X1 U3087 ( .A1(a_12_), .A2(n3114), .A3(b_8_), .ZN(n3113) );
  NAND2_X1 U3088 ( .A1(n2986), .A2(n2984), .ZN(n3114) );
  OR2_X1 U3089 ( .A1(n2984), .A2(n2986), .ZN(n3112) );
  AND2_X1 U3090 ( .A1(n3115), .A2(n3116), .ZN(n2986) );
  NAND2_X1 U3091 ( .A1(n3000), .A2(n3117), .ZN(n3116) );
  OR2_X1 U3092 ( .A1(n3001), .A2(n3002), .ZN(n3117) );
  NOR2_X1 U3093 ( .A1(n2217), .A2(n1988), .ZN(n3000) );
  NAND2_X1 U3094 ( .A1(n3002), .A2(n3001), .ZN(n3115) );
  NAND2_X1 U3095 ( .A1(n3118), .A2(n3119), .ZN(n3001) );
  NAND2_X1 U3096 ( .A1(b_6_), .A2(n3120), .ZN(n3119) );
  NAND2_X1 U3097 ( .A1(n1964), .A2(n3121), .ZN(n3120) );
  NAND2_X1 U3098 ( .A1(a_15_), .A2(n2074), .ZN(n3121) );
  NAND2_X1 U3099 ( .A1(b_7_), .A2(n3122), .ZN(n3118) );
  NAND2_X1 U3100 ( .A1(n1967), .A2(n3123), .ZN(n3122) );
  NAND2_X1 U3101 ( .A1(a_14_), .A2(n3124), .ZN(n3123) );
  AND3_X1 U3102 ( .A1(b_8_), .A2(b_7_), .A3(n2215), .ZN(n3002) );
  XNOR2_X1 U3103 ( .A(n3125), .B(n3126), .ZN(n2984) );
  XOR2_X1 U3104 ( .A(n3127), .B(n3128), .Z(n3125) );
  XNOR2_X1 U3105 ( .A(n3129), .B(n3130), .ZN(n3008) );
  NAND2_X1 U3106 ( .A1(n3131), .A2(n3132), .ZN(n3129) );
  NOR2_X1 U3107 ( .A1(n2217), .A2(n2218), .ZN(n3014) );
  XNOR2_X1 U3108 ( .A(n3133), .B(n3134), .ZN(n3016) );
  XNOR2_X1 U3109 ( .A(n3135), .B(n3136), .ZN(n3133) );
  XOR2_X1 U3110 ( .A(n3137), .B(n3138), .Z(n3019) );
  XNOR2_X1 U3111 ( .A(n3139), .B(n2196), .ZN(n3137) );
  INV_X1 U3112 ( .A(n2072), .ZN(n2196) );
  XOR2_X1 U3113 ( .A(n3140), .B(n3141), .Z(n2953) );
  XOR2_X1 U3114 ( .A(n3142), .B(n3143), .Z(n3141) );
  NAND2_X1 U3115 ( .A1(a_6_), .A2(b_7_), .ZN(n3143) );
  XOR2_X1 U3116 ( .A(n3144), .B(n3145), .Z(n3023) );
  XOR2_X1 U3117 ( .A(n3146), .B(n3147), .Z(n3145) );
  NAND2_X1 U3118 ( .A1(a_5_), .A2(b_7_), .ZN(n3147) );
  XOR2_X1 U3119 ( .A(n3148), .B(n3149), .Z(n3028) );
  XOR2_X1 U3120 ( .A(n3150), .B(n3151), .Z(n3148) );
  NOR2_X1 U3121 ( .A1(n2074), .A2(n2119), .ZN(n3151) );
  XOR2_X1 U3122 ( .A(n3152), .B(n3153), .Z(n3031) );
  XOR2_X1 U3123 ( .A(n3154), .B(n3155), .Z(n3153) );
  NAND2_X1 U3124 ( .A1(a_3_), .A2(b_7_), .ZN(n3155) );
  XOR2_X1 U3125 ( .A(n3046), .B(n3045), .Z(n3047) );
  NAND2_X1 U3126 ( .A1(n3156), .A2(n3157), .ZN(n1937) );
  NAND2_X1 U3127 ( .A1(n3045), .A2(n3046), .ZN(n3157) );
  XNOR2_X1 U3128 ( .A(n3158), .B(n3159), .ZN(n3156) );
  NAND3_X1 U3129 ( .A1(n3160), .A2(n3046), .A3(n3045), .ZN(n1936) );
  XNOR2_X1 U3130 ( .A(n3161), .B(n3162), .ZN(n3045) );
  XOR2_X1 U3131 ( .A(n3163), .B(n3164), .Z(n3162) );
  NAND2_X1 U3132 ( .A1(a_0_), .A2(b_6_), .ZN(n3164) );
  NAND2_X1 U3133 ( .A1(n3165), .A2(n3166), .ZN(n3046) );
  NAND3_X1 U3134 ( .A1(b_7_), .A2(n3167), .A3(a_0_), .ZN(n3166) );
  OR2_X1 U3135 ( .A1(n3048), .A2(n3050), .ZN(n3167) );
  NAND2_X1 U3136 ( .A1(n3048), .A2(n3050), .ZN(n3165) );
  NAND2_X1 U3137 ( .A1(n3168), .A2(n3169), .ZN(n3050) );
  NAND3_X1 U3138 ( .A1(a_1_), .A2(n3170), .A3(b_7_), .ZN(n3169) );
  NAND2_X1 U3139 ( .A1(n3059), .A2(n3057), .ZN(n3170) );
  OR2_X1 U3140 ( .A1(n3057), .A2(n3059), .ZN(n3168) );
  AND2_X1 U3141 ( .A1(n3171), .A2(n3172), .ZN(n3059) );
  NAND2_X1 U3142 ( .A1(n3067), .A2(n3173), .ZN(n3172) );
  NAND2_X1 U3143 ( .A1(n3066), .A2(n3065), .ZN(n3173) );
  NOR2_X1 U3144 ( .A1(n2220), .A2(n2074), .ZN(n3067) );
  OR2_X1 U3145 ( .A1(n3065), .A2(n3066), .ZN(n3171) );
  AND2_X1 U3146 ( .A1(n3174), .A2(n3175), .ZN(n3066) );
  NAND3_X1 U3147 ( .A1(b_7_), .A2(n3176), .A3(a_3_), .ZN(n3175) );
  OR2_X1 U3148 ( .A1(n3152), .A2(n3154), .ZN(n3176) );
  NAND2_X1 U3149 ( .A1(n3152), .A2(n3154), .ZN(n3174) );
  NAND2_X1 U3150 ( .A1(n3177), .A2(n3178), .ZN(n3154) );
  NAND3_X1 U3151 ( .A1(b_7_), .A2(n3179), .A3(a_4_), .ZN(n3178) );
  OR2_X1 U3152 ( .A1(n3150), .A2(n3149), .ZN(n3179) );
  NAND2_X1 U3153 ( .A1(n3149), .A2(n3150), .ZN(n3177) );
  NAND2_X1 U3154 ( .A1(n3180), .A2(n3181), .ZN(n3150) );
  NAND3_X1 U3155 ( .A1(b_7_), .A2(n3182), .A3(a_5_), .ZN(n3181) );
  OR2_X1 U3156 ( .A1(n3144), .A2(n3146), .ZN(n3182) );
  NAND2_X1 U3157 ( .A1(n3144), .A2(n3146), .ZN(n3180) );
  NAND2_X1 U3158 ( .A1(n3183), .A2(n3184), .ZN(n3146) );
  NAND3_X1 U3159 ( .A1(b_7_), .A2(n3185), .A3(a_6_), .ZN(n3184) );
  OR2_X1 U3160 ( .A1(n3140), .A2(n3142), .ZN(n3185) );
  NAND2_X1 U3161 ( .A1(n3140), .A2(n3142), .ZN(n3183) );
  NAND2_X1 U3162 ( .A1(n3186), .A2(n3187), .ZN(n3142) );
  NAND2_X1 U3163 ( .A1(n3138), .A2(n3188), .ZN(n3187) );
  OR2_X1 U3164 ( .A1(n3139), .A2(n2072), .ZN(n3188) );
  XNOR2_X1 U3165 ( .A(n3189), .B(n3190), .ZN(n3138) );
  XOR2_X1 U3166 ( .A(n3191), .B(n3192), .Z(n3190) );
  NAND2_X1 U3167 ( .A1(b_6_), .A2(a_8_), .ZN(n3192) );
  NAND2_X1 U3168 ( .A1(n2072), .A2(n3139), .ZN(n3186) );
  NAND2_X1 U3169 ( .A1(n3193), .A2(n3194), .ZN(n3139) );
  NAND2_X1 U3170 ( .A1(n3136), .A2(n3195), .ZN(n3194) );
  NAND2_X1 U3171 ( .A1(n3135), .A2(n3134), .ZN(n3195) );
  NOR2_X1 U3172 ( .A1(n2074), .A2(n2218), .ZN(n3136) );
  OR2_X1 U3173 ( .A1(n3134), .A2(n3135), .ZN(n3193) );
  AND2_X1 U3174 ( .A1(n3196), .A2(n3197), .ZN(n3135) );
  NAND2_X1 U3175 ( .A1(n3092), .A2(n3198), .ZN(n3197) );
  NAND2_X1 U3176 ( .A1(n3091), .A2(n3090), .ZN(n3198) );
  NOR2_X1 U3177 ( .A1(n2074), .A2(n2046), .ZN(n3092) );
  OR2_X1 U3178 ( .A1(n3090), .A2(n3091), .ZN(n3196) );
  AND2_X1 U3179 ( .A1(n3131), .A2(n3199), .ZN(n3091) );
  NAND2_X1 U3180 ( .A1(n3130), .A2(n3132), .ZN(n3199) );
  NAND2_X1 U3181 ( .A1(n3200), .A2(n3201), .ZN(n3132) );
  NAND2_X1 U3182 ( .A1(b_7_), .A2(a_10_), .ZN(n3201) );
  INV_X1 U3183 ( .A(n3202), .ZN(n3200) );
  XNOR2_X1 U3184 ( .A(n3203), .B(n3204), .ZN(n3130) );
  NAND2_X1 U3185 ( .A1(n3205), .A2(n3206), .ZN(n3203) );
  NAND2_X1 U3186 ( .A1(a_10_), .A2(n3202), .ZN(n3131) );
  NAND2_X1 U3187 ( .A1(n3102), .A2(n3207), .ZN(n3202) );
  NAND2_X1 U3188 ( .A1(n3101), .A2(n3103), .ZN(n3207) );
  NAND2_X1 U3189 ( .A1(n3208), .A2(n3209), .ZN(n3103) );
  NAND2_X1 U3190 ( .A1(b_7_), .A2(a_11_), .ZN(n3209) );
  INV_X1 U3191 ( .A(n3210), .ZN(n3208) );
  XNOR2_X1 U3192 ( .A(n3211), .B(n3212), .ZN(n3101) );
  XOR2_X1 U3193 ( .A(n3213), .B(n3214), .Z(n3211) );
  NAND2_X1 U3194 ( .A1(b_6_), .A2(a_12_), .ZN(n3213) );
  NAND2_X1 U3195 ( .A1(a_11_), .A2(n3210), .ZN(n3102) );
  NAND2_X1 U3196 ( .A1(n3215), .A2(n3216), .ZN(n3210) );
  NAND3_X1 U3197 ( .A1(a_12_), .A2(n3217), .A3(b_7_), .ZN(n3216) );
  NAND2_X1 U3198 ( .A1(n3111), .A2(n3109), .ZN(n3217) );
  OR2_X1 U3199 ( .A1(n3109), .A2(n3111), .ZN(n3215) );
  AND2_X1 U3200 ( .A1(n3218), .A2(n3219), .ZN(n3111) );
  NAND2_X1 U3201 ( .A1(n3126), .A2(n3220), .ZN(n3219) );
  OR2_X1 U3202 ( .A1(n3127), .A2(n3128), .ZN(n3220) );
  NOR2_X1 U3203 ( .A1(n2074), .A2(n1988), .ZN(n3126) );
  NAND2_X1 U3204 ( .A1(n3128), .A2(n3127), .ZN(n3218) );
  NAND2_X1 U3205 ( .A1(n3221), .A2(n3222), .ZN(n3127) );
  NAND2_X1 U3206 ( .A1(b_5_), .A2(n3223), .ZN(n3222) );
  NAND2_X1 U3207 ( .A1(n1964), .A2(n3224), .ZN(n3223) );
  NAND2_X1 U3208 ( .A1(a_15_), .A2(n3124), .ZN(n3224) );
  NAND2_X1 U3209 ( .A1(b_6_), .A2(n3225), .ZN(n3221) );
  NAND2_X1 U3210 ( .A1(n1967), .A2(n3226), .ZN(n3225) );
  NAND2_X1 U3211 ( .A1(a_14_), .A2(n2106), .ZN(n3226) );
  AND3_X1 U3212 ( .A1(b_6_), .A2(b_7_), .A3(n2215), .ZN(n3128) );
  XNOR2_X1 U3213 ( .A(n3227), .B(n3228), .ZN(n3109) );
  XOR2_X1 U3214 ( .A(n3229), .B(n3230), .Z(n3227) );
  XOR2_X1 U3215 ( .A(n3231), .B(n3232), .Z(n3090) );
  NAND2_X1 U3216 ( .A1(n3233), .A2(n3234), .ZN(n3231) );
  XOR2_X1 U3217 ( .A(n3235), .B(n3236), .Z(n3134) );
  NAND2_X1 U3218 ( .A1(n3237), .A2(n3238), .ZN(n3235) );
  NOR2_X1 U3219 ( .A1(n2076), .A2(n2074), .ZN(n2072) );
  XOR2_X1 U3220 ( .A(n3239), .B(n3240), .Z(n3140) );
  XOR2_X1 U3221 ( .A(n3241), .B(n3242), .Z(n3239) );
  NOR2_X1 U3222 ( .A1(n2076), .A2(n3124), .ZN(n3242) );
  XOR2_X1 U3223 ( .A(n3243), .B(n3244), .Z(n3144) );
  XNOR2_X1 U3224 ( .A(n2094), .B(n3245), .ZN(n3244) );
  XOR2_X1 U3225 ( .A(n3246), .B(n3247), .Z(n3149) );
  NOR2_X1 U3226 ( .A1(n3248), .A2(n3249), .ZN(n3247) );
  NOR2_X1 U3227 ( .A1(n3250), .A2(n3251), .ZN(n3248) );
  NOR2_X1 U3228 ( .A1(n3124), .A2(n2104), .ZN(n3251) );
  INV_X1 U3229 ( .A(n3252), .ZN(n3250) );
  XOR2_X1 U3230 ( .A(n3253), .B(n3254), .Z(n3152) );
  XOR2_X1 U3231 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR2_X1 U3232 ( .A(n3257), .B(n3258), .Z(n3065) );
  NAND2_X1 U3233 ( .A1(n3259), .A2(n3260), .ZN(n3257) );
  XNOR2_X1 U3234 ( .A(n3261), .B(n3262), .ZN(n3057) );
  XNOR2_X1 U3235 ( .A(n3263), .B(n3264), .ZN(n3261) );
  NAND2_X1 U3236 ( .A1(a_2_), .A2(b_6_), .ZN(n3263) );
  XOR2_X1 U3237 ( .A(n3265), .B(n3266), .Z(n3048) );
  XOR2_X1 U3238 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR2_X1 U3239 ( .A(n3158), .B(n3159), .Z(n3160) );
  NAND2_X1 U3240 ( .A1(n3269), .A2(n3270), .ZN(n1942) );
  NAND2_X1 U3241 ( .A1(n3159), .A2(n3158), .ZN(n3270) );
  XNOR2_X1 U3242 ( .A(n3271), .B(n3272), .ZN(n3269) );
  NAND3_X1 U3243 ( .A1(n3159), .A2(n3158), .A3(n3273), .ZN(n1941) );
  XNOR2_X1 U3244 ( .A(n3271), .B(n3274), .ZN(n3273) );
  INV_X1 U3245 ( .A(n3272), .ZN(n3274) );
  NAND2_X1 U3246 ( .A1(n3275), .A2(n3276), .ZN(n3158) );
  NAND3_X1 U3247 ( .A1(b_6_), .A2(n3277), .A3(a_0_), .ZN(n3276) );
  OR2_X1 U3248 ( .A1(n3161), .A2(n3163), .ZN(n3277) );
  NAND2_X1 U3249 ( .A1(n3161), .A2(n3163), .ZN(n3275) );
  NAND2_X1 U3250 ( .A1(n3278), .A2(n3279), .ZN(n3163) );
  NAND2_X1 U3251 ( .A1(n3268), .A2(n3280), .ZN(n3279) );
  NAND2_X1 U3252 ( .A1(n3267), .A2(n3265), .ZN(n3280) );
  NOR2_X1 U3253 ( .A1(n3124), .A2(n2396), .ZN(n3268) );
  OR2_X1 U3254 ( .A1(n3265), .A2(n3267), .ZN(n3278) );
  AND2_X1 U3255 ( .A1(n3281), .A2(n3282), .ZN(n3267) );
  NAND3_X1 U3256 ( .A1(b_6_), .A2(n3283), .A3(a_2_), .ZN(n3282) );
  OR2_X1 U3257 ( .A1(n3262), .A2(n3264), .ZN(n3283) );
  NAND2_X1 U3258 ( .A1(n3262), .A2(n3264), .ZN(n3281) );
  NAND2_X1 U3259 ( .A1(n3259), .A2(n3284), .ZN(n3264) );
  NAND2_X1 U3260 ( .A1(n3258), .A2(n3260), .ZN(n3284) );
  NAND2_X1 U3261 ( .A1(n3285), .A2(n3286), .ZN(n3260) );
  NAND2_X1 U3262 ( .A1(a_3_), .A2(b_6_), .ZN(n3286) );
  INV_X1 U3263 ( .A(n3287), .ZN(n3285) );
  XNOR2_X1 U3264 ( .A(n3288), .B(n3289), .ZN(n3258) );
  XNOR2_X1 U3265 ( .A(n3290), .B(n3291), .ZN(n3288) );
  NOR2_X1 U3266 ( .A1(n2106), .A2(n2119), .ZN(n3291) );
  NAND2_X1 U3267 ( .A1(a_3_), .A2(n3287), .ZN(n3259) );
  NAND2_X1 U3268 ( .A1(n3292), .A2(n3293), .ZN(n3287) );
  NAND2_X1 U3269 ( .A1(n3256), .A2(n3294), .ZN(n3293) );
  NAND2_X1 U3270 ( .A1(n3255), .A2(n3253), .ZN(n3294) );
  NOR2_X1 U3271 ( .A1(n2119), .A2(n3124), .ZN(n3256) );
  OR2_X1 U3272 ( .A1(n3253), .A2(n3255), .ZN(n3292) );
  NOR2_X1 U3273 ( .A1(n3249), .A2(n3295), .ZN(n3255) );
  AND2_X1 U3274 ( .A1(n3246), .A2(n3296), .ZN(n3295) );
  NAND2_X1 U3275 ( .A1(n3252), .A2(n3297), .ZN(n3296) );
  NAND2_X1 U3276 ( .A1(a_5_), .A2(b_6_), .ZN(n3297) );
  XNOR2_X1 U3277 ( .A(n3298), .B(n3299), .ZN(n3246) );
  XOR2_X1 U3278 ( .A(n3300), .B(n3301), .Z(n3299) );
  NAND2_X1 U3279 ( .A1(b_5_), .A2(a_6_), .ZN(n3301) );
  NOR2_X1 U3280 ( .A1(n3252), .A2(n2104), .ZN(n3249) );
  NAND2_X1 U3281 ( .A1(n3302), .A2(n3303), .ZN(n3252) );
  NAND2_X1 U3282 ( .A1(n3243), .A2(n3304), .ZN(n3303) );
  NAND2_X1 U3283 ( .A1(n2094), .A2(n3245), .ZN(n3304) );
  XNOR2_X1 U3284 ( .A(n3305), .B(n3306), .ZN(n3243) );
  XOR2_X1 U3285 ( .A(n3307), .B(n3308), .Z(n3305) );
  NOR2_X1 U3286 ( .A1(n2076), .A2(n2106), .ZN(n3308) );
  OR2_X1 U3287 ( .A1(n3245), .A2(n2094), .ZN(n3302) );
  NOR2_X1 U3288 ( .A1(n3124), .A2(n2089), .ZN(n2094) );
  NAND2_X1 U3289 ( .A1(n3309), .A2(n3310), .ZN(n3245) );
  NAND3_X1 U3290 ( .A1(a_7_), .A2(n3311), .A3(b_6_), .ZN(n3310) );
  OR2_X1 U3291 ( .A1(n3241), .A2(n3240), .ZN(n3311) );
  NAND2_X1 U3292 ( .A1(n3240), .A2(n3241), .ZN(n3309) );
  NAND2_X1 U3293 ( .A1(n3312), .A2(n3313), .ZN(n3241) );
  NAND3_X1 U3294 ( .A1(a_8_), .A2(n3314), .A3(b_6_), .ZN(n3313) );
  OR2_X1 U3295 ( .A1(n3189), .A2(n3191), .ZN(n3314) );
  NAND2_X1 U3296 ( .A1(n3189), .A2(n3191), .ZN(n3312) );
  NAND2_X1 U3297 ( .A1(n3237), .A2(n3315), .ZN(n3191) );
  NAND2_X1 U3298 ( .A1(n3236), .A2(n3238), .ZN(n3315) );
  NAND2_X1 U3299 ( .A1(n3316), .A2(n3317), .ZN(n3238) );
  NAND2_X1 U3300 ( .A1(b_6_), .A2(a_9_), .ZN(n3317) );
  INV_X1 U3301 ( .A(n3318), .ZN(n3316) );
  XNOR2_X1 U3302 ( .A(n3319), .B(n3320), .ZN(n3236) );
  XNOR2_X1 U3303 ( .A(n3321), .B(n3322), .ZN(n3320) );
  NAND2_X1 U3304 ( .A1(a_9_), .A2(n3318), .ZN(n3237) );
  NAND2_X1 U3305 ( .A1(n3233), .A2(n3323), .ZN(n3318) );
  NAND2_X1 U3306 ( .A1(n3232), .A2(n3234), .ZN(n3323) );
  NAND2_X1 U3307 ( .A1(n3324), .A2(n3325), .ZN(n3234) );
  NAND2_X1 U3308 ( .A1(b_6_), .A2(a_10_), .ZN(n3325) );
  INV_X1 U3309 ( .A(n3326), .ZN(n3324) );
  XNOR2_X1 U3310 ( .A(n3327), .B(n3328), .ZN(n3232) );
  XNOR2_X1 U3311 ( .A(n3329), .B(n3330), .ZN(n3327) );
  NAND2_X1 U3312 ( .A1(a_10_), .A2(n3326), .ZN(n3233) );
  NAND2_X1 U3313 ( .A1(n3205), .A2(n3331), .ZN(n3326) );
  NAND2_X1 U3314 ( .A1(n3204), .A2(n3206), .ZN(n3331) );
  NAND2_X1 U3315 ( .A1(n3332), .A2(n3333), .ZN(n3206) );
  NAND2_X1 U3316 ( .A1(b_6_), .A2(a_11_), .ZN(n3333) );
  INV_X1 U3317 ( .A(n3334), .ZN(n3332) );
  XNOR2_X1 U3318 ( .A(n3335), .B(n3336), .ZN(n3204) );
  XOR2_X1 U3319 ( .A(n3337), .B(n3338), .Z(n3335) );
  NAND2_X1 U3320 ( .A1(b_5_), .A2(a_12_), .ZN(n3337) );
  NAND2_X1 U3321 ( .A1(a_11_), .A2(n3334), .ZN(n3205) );
  NAND2_X1 U3322 ( .A1(n3339), .A2(n3340), .ZN(n3334) );
  NAND3_X1 U3323 ( .A1(a_12_), .A2(n3341), .A3(b_6_), .ZN(n3340) );
  NAND2_X1 U3324 ( .A1(n3214), .A2(n3212), .ZN(n3341) );
  OR2_X1 U3325 ( .A1(n3212), .A2(n3214), .ZN(n3339) );
  AND2_X1 U3326 ( .A1(n3342), .A2(n3343), .ZN(n3214) );
  NAND2_X1 U3327 ( .A1(n3228), .A2(n3344), .ZN(n3343) );
  OR2_X1 U3328 ( .A1(n3229), .A2(n3230), .ZN(n3344) );
  NOR2_X1 U3329 ( .A1(n3124), .A2(n1988), .ZN(n3228) );
  NAND2_X1 U3330 ( .A1(n3230), .A2(n3229), .ZN(n3342) );
  NAND2_X1 U3331 ( .A1(n3345), .A2(n3346), .ZN(n3229) );
  NAND2_X1 U3332 ( .A1(b_4_), .A2(n3347), .ZN(n3346) );
  NAND2_X1 U3333 ( .A1(n1964), .A2(n3348), .ZN(n3347) );
  NAND2_X1 U3334 ( .A1(a_15_), .A2(n2106), .ZN(n3348) );
  NAND2_X1 U3335 ( .A1(b_5_), .A2(n3349), .ZN(n3345) );
  NAND2_X1 U3336 ( .A1(n1967), .A2(n3350), .ZN(n3349) );
  NAND2_X1 U3337 ( .A1(a_14_), .A2(n3351), .ZN(n3350) );
  AND3_X1 U3338 ( .A1(b_6_), .A2(b_5_), .A3(n2215), .ZN(n3230) );
  XNOR2_X1 U3339 ( .A(n3352), .B(n3353), .ZN(n3212) );
  XOR2_X1 U3340 ( .A(n3354), .B(n3355), .Z(n3352) );
  XNOR2_X1 U3341 ( .A(n3356), .B(n3357), .ZN(n3189) );
  NAND2_X1 U3342 ( .A1(n3358), .A2(n3359), .ZN(n3356) );
  XOR2_X1 U3343 ( .A(n3360), .B(n3361), .Z(n3240) );
  XNOR2_X1 U3344 ( .A(n3362), .B(n3363), .ZN(n3360) );
  NAND2_X1 U3345 ( .A1(b_5_), .A2(a_8_), .ZN(n3362) );
  XNOR2_X1 U3346 ( .A(n3364), .B(n3365), .ZN(n3253) );
  XNOR2_X1 U3347 ( .A(n3366), .B(n2192), .ZN(n3364) );
  INV_X1 U3348 ( .A(n2101), .ZN(n2192) );
  XOR2_X1 U3349 ( .A(n3367), .B(n3368), .Z(n3262) );
  XOR2_X1 U3350 ( .A(n3369), .B(n3370), .Z(n3367) );
  NOR2_X1 U3351 ( .A1(n2106), .A2(n2139), .ZN(n3370) );
  XNOR2_X1 U3352 ( .A(n3371), .B(n3372), .ZN(n3265) );
  XOR2_X1 U3353 ( .A(n3373), .B(n3374), .Z(n3371) );
  NOR2_X1 U3354 ( .A1(n2106), .A2(n2220), .ZN(n3374) );
  XOR2_X1 U3355 ( .A(n3375), .B(n3376), .Z(n3161) );
  XNOR2_X1 U3356 ( .A(n3377), .B(n3378), .ZN(n3376) );
  NAND2_X1 U3357 ( .A1(b_5_), .A2(a_1_), .ZN(n3378) );
  XOR2_X1 U3358 ( .A(n3379), .B(n3380), .Z(n3159) );
  XOR2_X1 U3359 ( .A(n3381), .B(n3382), .Z(n3379) );
  NOR2_X1 U3360 ( .A1(n2106), .A2(n2407), .ZN(n3382) );
  NAND2_X1 U3361 ( .A1(n3383), .A2(n3384), .ZN(n1947) );
  NAND2_X1 U3362 ( .A1(n3272), .A2(n3271), .ZN(n3384) );
  XNOR2_X1 U3363 ( .A(n3385), .B(n3386), .ZN(n3383) );
  NAND3_X1 U3364 ( .A1(n3272), .A2(n3271), .A3(n3387), .ZN(n1946) );
  XOR2_X1 U3365 ( .A(n3385), .B(n3386), .Z(n3387) );
  NAND2_X1 U3366 ( .A1(n3388), .A2(n3389), .ZN(n3271) );
  NAND3_X1 U3367 ( .A1(b_5_), .A2(n3390), .A3(a_0_), .ZN(n3389) );
  OR2_X1 U3368 ( .A1(n3380), .A2(n3381), .ZN(n3390) );
  NAND2_X1 U3369 ( .A1(n3380), .A2(n3381), .ZN(n3388) );
  NAND2_X1 U3370 ( .A1(n3391), .A2(n3392), .ZN(n3381) );
  NAND3_X1 U3371 ( .A1(a_1_), .A2(n3393), .A3(b_5_), .ZN(n3392) );
  NAND2_X1 U3372 ( .A1(n3377), .A2(n3375), .ZN(n3393) );
  OR2_X1 U3373 ( .A1(n3375), .A2(n3377), .ZN(n3391) );
  AND2_X1 U3374 ( .A1(n3394), .A2(n3395), .ZN(n3377) );
  NAND3_X1 U3375 ( .A1(b_5_), .A2(n3396), .A3(a_2_), .ZN(n3395) );
  OR2_X1 U3376 ( .A1(n3372), .A2(n3373), .ZN(n3396) );
  NAND2_X1 U3377 ( .A1(n3372), .A2(n3373), .ZN(n3394) );
  NAND2_X1 U3378 ( .A1(n3397), .A2(n3398), .ZN(n3373) );
  NAND3_X1 U3379 ( .A1(b_5_), .A2(n3399), .A3(a_3_), .ZN(n3398) );
  OR2_X1 U3380 ( .A1(n3369), .A2(n3368), .ZN(n3399) );
  NAND2_X1 U3381 ( .A1(n3368), .A2(n3369), .ZN(n3397) );
  NAND2_X1 U3382 ( .A1(n3400), .A2(n3401), .ZN(n3369) );
  NAND3_X1 U3383 ( .A1(b_5_), .A2(n3402), .A3(a_4_), .ZN(n3401) );
  NAND2_X1 U3384 ( .A1(n3289), .A2(n3290), .ZN(n3402) );
  OR2_X1 U3385 ( .A1(n3289), .A2(n3290), .ZN(n3400) );
  AND2_X1 U3386 ( .A1(n3403), .A2(n3404), .ZN(n3290) );
  NAND2_X1 U3387 ( .A1(n3365), .A2(n3405), .ZN(n3404) );
  OR2_X1 U3388 ( .A1(n3366), .A2(n2101), .ZN(n3405) );
  XNOR2_X1 U3389 ( .A(n3406), .B(n3407), .ZN(n3365) );
  XOR2_X1 U3390 ( .A(n3408), .B(n3409), .Z(n3407) );
  NAND2_X1 U3391 ( .A1(b_4_), .A2(a_6_), .ZN(n3409) );
  NAND2_X1 U3392 ( .A1(n2101), .A2(n3366), .ZN(n3403) );
  NAND2_X1 U3393 ( .A1(n3410), .A2(n3411), .ZN(n3366) );
  NAND3_X1 U3394 ( .A1(a_6_), .A2(n3412), .A3(b_5_), .ZN(n3411) );
  OR2_X1 U3395 ( .A1(n3298), .A2(n3300), .ZN(n3412) );
  NAND2_X1 U3396 ( .A1(n3298), .A2(n3300), .ZN(n3410) );
  NAND2_X1 U3397 ( .A1(n3413), .A2(n3414), .ZN(n3300) );
  NAND3_X1 U3398 ( .A1(a_7_), .A2(n3415), .A3(b_5_), .ZN(n3414) );
  OR2_X1 U3399 ( .A1(n3306), .A2(n3307), .ZN(n3415) );
  NAND2_X1 U3400 ( .A1(n3306), .A2(n3307), .ZN(n3413) );
  NAND2_X1 U3401 ( .A1(n3416), .A2(n3417), .ZN(n3307) );
  NAND3_X1 U3402 ( .A1(a_8_), .A2(n3418), .A3(b_5_), .ZN(n3417) );
  OR2_X1 U3403 ( .A1(n3361), .A2(n3363), .ZN(n3418) );
  NAND2_X1 U3404 ( .A1(n3361), .A2(n3363), .ZN(n3416) );
  NAND2_X1 U3405 ( .A1(n3358), .A2(n3419), .ZN(n3363) );
  NAND2_X1 U3406 ( .A1(n3357), .A2(n3359), .ZN(n3419) );
  NAND2_X1 U3407 ( .A1(n3420), .A2(n3421), .ZN(n3359) );
  NAND2_X1 U3408 ( .A1(b_5_), .A2(a_9_), .ZN(n3421) );
  INV_X1 U3409 ( .A(n3422), .ZN(n3420) );
  XNOR2_X1 U3410 ( .A(n3423), .B(n3424), .ZN(n3357) );
  XNOR2_X1 U3411 ( .A(n3425), .B(n3426), .ZN(n3424) );
  NAND2_X1 U3412 ( .A1(a_9_), .A2(n3422), .ZN(n3358) );
  NAND2_X1 U3413 ( .A1(n3427), .A2(n3428), .ZN(n3422) );
  NAND2_X1 U3414 ( .A1(n3322), .A2(n3429), .ZN(n3428) );
  OR2_X1 U3415 ( .A1(n3319), .A2(n3321), .ZN(n3429) );
  NOR2_X1 U3416 ( .A1(n2106), .A2(n2586), .ZN(n3322) );
  NAND2_X1 U3417 ( .A1(n3319), .A2(n3321), .ZN(n3427) );
  NAND2_X1 U3418 ( .A1(n3430), .A2(n3431), .ZN(n3321) );
  NAND2_X1 U3419 ( .A1(n3330), .A2(n3432), .ZN(n3431) );
  NAND2_X1 U3420 ( .A1(n3328), .A2(n3329), .ZN(n3432) );
  NOR2_X1 U3421 ( .A1(n2106), .A2(n2019), .ZN(n3330) );
  OR2_X1 U3422 ( .A1(n3328), .A2(n3329), .ZN(n3430) );
  AND2_X1 U3423 ( .A1(n3433), .A2(n3434), .ZN(n3329) );
  NAND3_X1 U3424 ( .A1(a_12_), .A2(n3435), .A3(b_5_), .ZN(n3434) );
  NAND2_X1 U3425 ( .A1(n3338), .A2(n3336), .ZN(n3435) );
  OR2_X1 U3426 ( .A1(n3336), .A2(n3338), .ZN(n3433) );
  AND2_X1 U3427 ( .A1(n3436), .A2(n3437), .ZN(n3338) );
  NAND2_X1 U3428 ( .A1(n3353), .A2(n3438), .ZN(n3437) );
  OR2_X1 U3429 ( .A1(n3354), .A2(n3355), .ZN(n3438) );
  NOR2_X1 U3430 ( .A1(n2106), .A2(n1988), .ZN(n3353) );
  NAND2_X1 U3431 ( .A1(n3355), .A2(n3354), .ZN(n3436) );
  NAND2_X1 U3432 ( .A1(n3439), .A2(n3440), .ZN(n3354) );
  NAND2_X1 U3433 ( .A1(b_3_), .A2(n3441), .ZN(n3440) );
  NAND2_X1 U3434 ( .A1(n1964), .A2(n3442), .ZN(n3441) );
  NAND2_X1 U3435 ( .A1(a_15_), .A2(n3351), .ZN(n3442) );
  NAND2_X1 U3436 ( .A1(b_4_), .A2(n3443), .ZN(n3439) );
  NAND2_X1 U3437 ( .A1(n1967), .A2(n3444), .ZN(n3443) );
  NAND2_X1 U3438 ( .A1(a_14_), .A2(n2141), .ZN(n3444) );
  AND3_X1 U3439 ( .A1(b_4_), .A2(b_5_), .A3(n2215), .ZN(n3355) );
  XNOR2_X1 U3440 ( .A(n3445), .B(n3446), .ZN(n3336) );
  XOR2_X1 U3441 ( .A(n3447), .B(n3448), .Z(n3445) );
  XNOR2_X1 U3442 ( .A(n3449), .B(n3450), .ZN(n3328) );
  XNOR2_X1 U3443 ( .A(n3451), .B(n3452), .ZN(n3449) );
  NAND2_X1 U3444 ( .A1(b_4_), .A2(a_12_), .ZN(n3451) );
  XNOR2_X1 U3445 ( .A(n3453), .B(n3454), .ZN(n3319) );
  NAND2_X1 U3446 ( .A1(n3455), .A2(n3456), .ZN(n3453) );
  XNOR2_X1 U3447 ( .A(n3457), .B(n3458), .ZN(n3361) );
  NAND2_X1 U3448 ( .A1(n3459), .A2(n3460), .ZN(n3457) );
  XOR2_X1 U3449 ( .A(n3461), .B(n3462), .Z(n3306) );
  XOR2_X1 U3450 ( .A(n3463), .B(n3464), .Z(n3461) );
  NOR2_X1 U3451 ( .A1(n2218), .A2(n3351), .ZN(n3464) );
  XOR2_X1 U3452 ( .A(n3465), .B(n3466), .Z(n3298) );
  XNOR2_X1 U3453 ( .A(n3467), .B(n3468), .ZN(n3466) );
  NAND2_X1 U3454 ( .A1(b_4_), .A2(a_7_), .ZN(n3468) );
  NOR2_X1 U3455 ( .A1(n2104), .A2(n2106), .ZN(n2101) );
  XNOR2_X1 U3456 ( .A(n3469), .B(n3470), .ZN(n3289) );
  XOR2_X1 U3457 ( .A(n3471), .B(n3472), .Z(n3469) );
  NOR2_X1 U3458 ( .A1(n2104), .A2(n3351), .ZN(n3472) );
  XNOR2_X1 U3459 ( .A(n3473), .B(n3474), .ZN(n3368) );
  XNOR2_X1 U3460 ( .A(n2124), .B(n3475), .ZN(n3474) );
  XOR2_X1 U3461 ( .A(n3476), .B(n3477), .Z(n3372) );
  XNOR2_X1 U3462 ( .A(n3478), .B(n3479), .ZN(n3476) );
  NAND2_X1 U3463 ( .A1(a_3_), .A2(b_4_), .ZN(n3478) );
  XOR2_X1 U3464 ( .A(n3480), .B(n3481), .Z(n3375) );
  XOR2_X1 U3465 ( .A(n3482), .B(n3483), .Z(n3481) );
  NAND2_X1 U3466 ( .A1(a_2_), .A2(b_4_), .ZN(n3483) );
  XOR2_X1 U3467 ( .A(n3484), .B(n3485), .Z(n3380) );
  XOR2_X1 U3468 ( .A(n3486), .B(n3487), .Z(n3484) );
  XOR2_X1 U3469 ( .A(n3488), .B(n3489), .Z(n3272) );
  XOR2_X1 U3470 ( .A(n3490), .B(n3491), .Z(n3488) );
  NOR2_X1 U3471 ( .A1(n3351), .A2(n2407), .ZN(n3491) );
  NAND2_X1 U3472 ( .A1(n3492), .A2(n3493), .ZN(n1952) );
  NAND2_X1 U3473 ( .A1(n3386), .A2(n3385), .ZN(n3493) );
  XNOR2_X1 U3474 ( .A(n3494), .B(n3495), .ZN(n3492) );
  NAND3_X1 U3475 ( .A1(n3386), .A2(n3385), .A3(n3496), .ZN(n1951) );
  XOR2_X1 U3476 ( .A(n3494), .B(n3495), .Z(n3496) );
  NAND2_X1 U3477 ( .A1(n3497), .A2(n3498), .ZN(n3385) );
  NAND3_X1 U3478 ( .A1(b_4_), .A2(n3499), .A3(a_0_), .ZN(n3498) );
  OR2_X1 U3479 ( .A1(n3490), .A2(n3489), .ZN(n3499) );
  NAND2_X1 U3480 ( .A1(n3489), .A2(n3490), .ZN(n3497) );
  NAND2_X1 U3481 ( .A1(n3500), .A2(n3501), .ZN(n3490) );
  NAND2_X1 U3482 ( .A1(n3487), .A2(n3502), .ZN(n3501) );
  OR2_X1 U3483 ( .A1(n3486), .A2(n3485), .ZN(n3502) );
  NOR2_X1 U3484 ( .A1(n3351), .A2(n2396), .ZN(n3487) );
  NAND2_X1 U3485 ( .A1(n3485), .A2(n3486), .ZN(n3500) );
  NAND2_X1 U3486 ( .A1(n3503), .A2(n3504), .ZN(n3486) );
  NAND3_X1 U3487 ( .A1(b_4_), .A2(n3505), .A3(a_2_), .ZN(n3504) );
  OR2_X1 U3488 ( .A1(n3480), .A2(n3482), .ZN(n3505) );
  NAND2_X1 U3489 ( .A1(n3480), .A2(n3482), .ZN(n3503) );
  NAND2_X1 U3490 ( .A1(n3506), .A2(n3507), .ZN(n3482) );
  NAND3_X1 U3491 ( .A1(b_4_), .A2(n3508), .A3(a_3_), .ZN(n3507) );
  OR2_X1 U3492 ( .A1(n3479), .A2(n3477), .ZN(n3508) );
  NAND2_X1 U3493 ( .A1(n3477), .A2(n3479), .ZN(n3506) );
  NAND2_X1 U3494 ( .A1(n3509), .A2(n3510), .ZN(n3479) );
  NAND2_X1 U3495 ( .A1(n3473), .A2(n3511), .ZN(n3510) );
  OR2_X1 U3496 ( .A1(n3475), .A2(n2124), .ZN(n3511) );
  XOR2_X1 U3497 ( .A(n3512), .B(n3513), .Z(n3473) );
  XOR2_X1 U3498 ( .A(n3514), .B(n3515), .Z(n3512) );
  NOR2_X1 U3499 ( .A1(n2104), .A2(n2141), .ZN(n3515) );
  NAND2_X1 U3500 ( .A1(n2124), .A2(n3475), .ZN(n3509) );
  NAND2_X1 U3501 ( .A1(n3516), .A2(n3517), .ZN(n3475) );
  NAND3_X1 U3502 ( .A1(a_5_), .A2(n3518), .A3(b_4_), .ZN(n3517) );
  OR2_X1 U3503 ( .A1(n3471), .A2(n3470), .ZN(n3518) );
  NAND2_X1 U3504 ( .A1(n3470), .A2(n3471), .ZN(n3516) );
  NAND2_X1 U3505 ( .A1(n3519), .A2(n3520), .ZN(n3471) );
  NAND3_X1 U3506 ( .A1(a_6_), .A2(n3521), .A3(b_4_), .ZN(n3520) );
  OR2_X1 U3507 ( .A1(n3408), .A2(n3406), .ZN(n3521) );
  NAND2_X1 U3508 ( .A1(n3406), .A2(n3408), .ZN(n3519) );
  NAND2_X1 U3509 ( .A1(n3522), .A2(n3523), .ZN(n3408) );
  NAND3_X1 U3510 ( .A1(a_7_), .A2(n3524), .A3(b_4_), .ZN(n3523) );
  NAND2_X1 U3511 ( .A1(n3467), .A2(n3465), .ZN(n3524) );
  OR2_X1 U3512 ( .A1(n3465), .A2(n3467), .ZN(n3522) );
  AND2_X1 U3513 ( .A1(n3525), .A2(n3526), .ZN(n3467) );
  NAND3_X1 U3514 ( .A1(a_8_), .A2(n3527), .A3(b_4_), .ZN(n3526) );
  OR2_X1 U3515 ( .A1(n3463), .A2(n3462), .ZN(n3527) );
  NAND2_X1 U3516 ( .A1(n3462), .A2(n3463), .ZN(n3525) );
  NAND2_X1 U3517 ( .A1(n3459), .A2(n3528), .ZN(n3463) );
  NAND2_X1 U3518 ( .A1(n3458), .A2(n3460), .ZN(n3528) );
  NAND2_X1 U3519 ( .A1(n3529), .A2(n3530), .ZN(n3460) );
  NAND2_X1 U3520 ( .A1(b_4_), .A2(a_9_), .ZN(n3530) );
  INV_X1 U3521 ( .A(n3531), .ZN(n3529) );
  XNOR2_X1 U3522 ( .A(n3532), .B(n3533), .ZN(n3458) );
  NAND2_X1 U3523 ( .A1(n3534), .A2(n3535), .ZN(n3532) );
  NAND2_X1 U3524 ( .A1(a_9_), .A2(n3531), .ZN(n3459) );
  NAND2_X1 U3525 ( .A1(n3536), .A2(n3537), .ZN(n3531) );
  NAND2_X1 U3526 ( .A1(n3426), .A2(n3538), .ZN(n3537) );
  OR2_X1 U3527 ( .A1(n3425), .A2(n3423), .ZN(n3538) );
  NOR2_X1 U3528 ( .A1(n3351), .A2(n2586), .ZN(n3426) );
  NAND2_X1 U3529 ( .A1(n3423), .A2(n3425), .ZN(n3536) );
  NAND2_X1 U3530 ( .A1(n3455), .A2(n3539), .ZN(n3425) );
  NAND2_X1 U3531 ( .A1(n3454), .A2(n3456), .ZN(n3539) );
  NAND2_X1 U3532 ( .A1(n3540), .A2(n3541), .ZN(n3456) );
  NAND2_X1 U3533 ( .A1(b_4_), .A2(a_11_), .ZN(n3541) );
  INV_X1 U3534 ( .A(n3542), .ZN(n3540) );
  XNOR2_X1 U3535 ( .A(n3543), .B(n3544), .ZN(n3454) );
  XNOR2_X1 U3536 ( .A(n3545), .B(n3546), .ZN(n3543) );
  NAND2_X1 U3537 ( .A1(a_11_), .A2(n3542), .ZN(n3455) );
  NAND2_X1 U3538 ( .A1(n3547), .A2(n3548), .ZN(n3542) );
  NAND3_X1 U3539 ( .A1(a_12_), .A2(n3549), .A3(b_4_), .ZN(n3548) );
  OR2_X1 U3540 ( .A1(n3452), .A2(n3450), .ZN(n3549) );
  NAND2_X1 U3541 ( .A1(n3450), .A2(n3452), .ZN(n3547) );
  NAND2_X1 U3542 ( .A1(n3550), .A2(n3551), .ZN(n3452) );
  NAND2_X1 U3543 ( .A1(n3446), .A2(n3552), .ZN(n3551) );
  OR2_X1 U3544 ( .A1(n3447), .A2(n3448), .ZN(n3552) );
  NOR2_X1 U3545 ( .A1(n3351), .A2(n1988), .ZN(n3446) );
  NAND2_X1 U3546 ( .A1(n3448), .A2(n3447), .ZN(n3550) );
  NAND2_X1 U3547 ( .A1(n3553), .A2(n3554), .ZN(n3447) );
  NAND2_X1 U3548 ( .A1(b_2_), .A2(n3555), .ZN(n3554) );
  NAND2_X1 U3549 ( .A1(n1964), .A2(n3556), .ZN(n3555) );
  NAND2_X1 U3550 ( .A1(a_15_), .A2(n2141), .ZN(n3556) );
  NAND2_X1 U3551 ( .A1(b_3_), .A2(n3557), .ZN(n3553) );
  NAND2_X1 U3552 ( .A1(n1967), .A2(n3558), .ZN(n3557) );
  NAND2_X1 U3553 ( .A1(a_14_), .A2(n2219), .ZN(n3558) );
  AND3_X1 U3554 ( .A1(b_4_), .A2(b_3_), .A3(n2215), .ZN(n3448) );
  XOR2_X1 U3555 ( .A(n3559), .B(n3560), .Z(n3450) );
  NOR2_X1 U3556 ( .A1(n1988), .A2(n2141), .ZN(n3560) );
  XOR2_X1 U3557 ( .A(n3561), .B(n3562), .Z(n3559) );
  XNOR2_X1 U3558 ( .A(n3563), .B(n3564), .ZN(n3423) );
  NAND2_X1 U3559 ( .A1(n3565), .A2(n3566), .ZN(n3563) );
  XNOR2_X1 U3560 ( .A(n3567), .B(n3568), .ZN(n3462) );
  NAND2_X1 U3561 ( .A1(n3569), .A2(n3570), .ZN(n3567) );
  XNOR2_X1 U3562 ( .A(n3571), .B(n3572), .ZN(n3465) );
  XOR2_X1 U3563 ( .A(n3573), .B(n3574), .Z(n3571) );
  NOR2_X1 U3564 ( .A1(n2218), .A2(n2141), .ZN(n3574) );
  XNOR2_X1 U3565 ( .A(n3575), .B(n3576), .ZN(n3406) );
  NAND2_X1 U3566 ( .A1(n3577), .A2(n3578), .ZN(n3575) );
  XOR2_X1 U3567 ( .A(n3579), .B(n3580), .Z(n3470) );
  XOR2_X1 U3568 ( .A(n3581), .B(n3582), .Z(n3579) );
  NOR2_X1 U3569 ( .A1(n2089), .A2(n2141), .ZN(n3582) );
  NOR2_X1 U3570 ( .A1(n3351), .A2(n2119), .ZN(n2124) );
  XNOR2_X1 U3571 ( .A(n3583), .B(n3584), .ZN(n3477) );
  XNOR2_X1 U3572 ( .A(n3585), .B(n3586), .ZN(n3583) );
  NOR2_X1 U3573 ( .A1(n2119), .A2(n2141), .ZN(n3586) );
  XOR2_X1 U3574 ( .A(n3587), .B(n3588), .Z(n3480) );
  XNOR2_X1 U3575 ( .A(n3589), .B(n2188), .ZN(n3587) );
  INV_X1 U3576 ( .A(n2136), .ZN(n2188) );
  XOR2_X1 U3577 ( .A(n3590), .B(n3591), .Z(n3485) );
  XOR2_X1 U3578 ( .A(n3592), .B(n3593), .Z(n3590) );
  NOR2_X1 U3579 ( .A1(n2141), .A2(n2220), .ZN(n3593) );
  XOR2_X1 U3580 ( .A(n3594), .B(n3595), .Z(n3489) );
  XOR2_X1 U3581 ( .A(n3596), .B(n3597), .Z(n3594) );
  XOR2_X1 U3582 ( .A(n3598), .B(n3599), .Z(n3386) );
  XOR2_X1 U3583 ( .A(n3600), .B(n3601), .Z(n3598) );
  NOR2_X1 U3584 ( .A1(n2141), .A2(n2407), .ZN(n3601) );
  NAND2_X1 U3585 ( .A1(n3602), .A2(n3603), .ZN(n1978) );
  NAND2_X1 U3586 ( .A1(n3495), .A2(n3494), .ZN(n3603) );
  XNOR2_X1 U3587 ( .A(n2255), .B(n2254), .ZN(n3602) );
  NAND3_X1 U3588 ( .A1(n3495), .A2(n3494), .A3(n3604), .ZN(n1977) );
  XOR2_X1 U3589 ( .A(n2255), .B(n2254), .Z(n3604) );
  NAND3_X1 U3590 ( .A1(n3605), .A2(n3606), .A3(n3607), .ZN(n2254) );
  XNOR2_X1 U3591 ( .A(n2258), .B(n2259), .ZN(n3607) );
  NOR2_X1 U3592 ( .A1(n2396), .A2(n3608), .ZN(n2259) );
  NOR2_X1 U3593 ( .A1(n2407), .A2(n2175), .ZN(n2258) );
  NAND3_X1 U3594 ( .A1(a_2_), .A2(b_0_), .A3(n2171), .ZN(n3606) );
  NAND2_X1 U3595 ( .A1(n3609), .A2(n3610), .ZN(n2255) );
  NAND2_X1 U3596 ( .A1(n3611), .A2(b_2_), .ZN(n3610) );
  NAND2_X1 U3597 ( .A1(n3612), .A2(n3613), .ZN(n3494) );
  NAND3_X1 U3598 ( .A1(b_3_), .A2(n3614), .A3(a_0_), .ZN(n3613) );
  OR2_X1 U3599 ( .A1(n3599), .A2(n3600), .ZN(n3614) );
  NAND2_X1 U3600 ( .A1(n3599), .A2(n3600), .ZN(n3612) );
  NAND2_X1 U3601 ( .A1(n3615), .A2(n3616), .ZN(n3600) );
  NAND2_X1 U3602 ( .A1(n3597), .A2(n3617), .ZN(n3616) );
  OR2_X1 U3603 ( .A1(n3595), .A2(n3596), .ZN(n3617) );
  NOR2_X1 U3604 ( .A1(n2141), .A2(n2396), .ZN(n3597) );
  NAND2_X1 U3605 ( .A1(n3595), .A2(n3596), .ZN(n3615) );
  NAND2_X1 U3606 ( .A1(n3618), .A2(n3619), .ZN(n3596) );
  NAND3_X1 U3607 ( .A1(b_3_), .A2(n3620), .A3(a_2_), .ZN(n3619) );
  OR2_X1 U3608 ( .A1(n3591), .A2(n3592), .ZN(n3620) );
  NAND2_X1 U3609 ( .A1(n3591), .A2(n3592), .ZN(n3618) );
  NAND2_X1 U3610 ( .A1(n3621), .A2(n3622), .ZN(n3592) );
  NAND2_X1 U3611 ( .A1(n3588), .A2(n3623), .ZN(n3622) );
  OR2_X1 U3612 ( .A1(n3589), .A2(n2136), .ZN(n3623) );
  XNOR2_X1 U3613 ( .A(n3624), .B(n3625), .ZN(n3588) );
  NAND2_X1 U3614 ( .A1(n3626), .A2(n3627), .ZN(n3624) );
  NAND2_X1 U3615 ( .A1(n2136), .A2(n3589), .ZN(n3621) );
  NAND2_X1 U3616 ( .A1(n3628), .A2(n3629), .ZN(n3589) );
  NAND3_X1 U3617 ( .A1(a_4_), .A2(n3630), .A3(b_3_), .ZN(n3629) );
  NAND2_X1 U3618 ( .A1(n3584), .A2(n3585), .ZN(n3630) );
  OR2_X1 U3619 ( .A1(n3584), .A2(n3585), .ZN(n3628) );
  AND2_X1 U3620 ( .A1(n3631), .A2(n3632), .ZN(n3585) );
  NAND3_X1 U3621 ( .A1(a_5_), .A2(n3633), .A3(b_3_), .ZN(n3632) );
  OR2_X1 U3622 ( .A1(n3514), .A2(n3513), .ZN(n3633) );
  NAND2_X1 U3623 ( .A1(n3513), .A2(n3514), .ZN(n3631) );
  NAND2_X1 U3624 ( .A1(n3634), .A2(n3635), .ZN(n3514) );
  NAND3_X1 U3625 ( .A1(a_6_), .A2(n3636), .A3(b_3_), .ZN(n3635) );
  OR2_X1 U3626 ( .A1(n3580), .A2(n3581), .ZN(n3636) );
  NAND2_X1 U3627 ( .A1(n3580), .A2(n3581), .ZN(n3634) );
  NAND2_X1 U3628 ( .A1(n3577), .A2(n3637), .ZN(n3581) );
  NAND2_X1 U3629 ( .A1(n3576), .A2(n3578), .ZN(n3637) );
  NAND2_X1 U3630 ( .A1(n3638), .A2(n3639), .ZN(n3578) );
  NAND2_X1 U3631 ( .A1(b_3_), .A2(a_7_), .ZN(n3639) );
  INV_X1 U3632 ( .A(n3640), .ZN(n3638) );
  XNOR2_X1 U3633 ( .A(n3641), .B(n3642), .ZN(n3576) );
  NAND2_X1 U3634 ( .A1(n3643), .A2(n3644), .ZN(n3641) );
  NAND2_X1 U3635 ( .A1(a_7_), .A2(n3640), .ZN(n3577) );
  NAND2_X1 U3636 ( .A1(n3645), .A2(n3646), .ZN(n3640) );
  NAND3_X1 U3637 ( .A1(a_8_), .A2(n3647), .A3(b_3_), .ZN(n3646) );
  OR2_X1 U3638 ( .A1(n3572), .A2(n3573), .ZN(n3647) );
  NAND2_X1 U3639 ( .A1(n3572), .A2(n3573), .ZN(n3645) );
  NAND2_X1 U3640 ( .A1(n3569), .A2(n3648), .ZN(n3573) );
  NAND2_X1 U3641 ( .A1(n3568), .A2(n3570), .ZN(n3648) );
  NAND2_X1 U3642 ( .A1(n3649), .A2(n3650), .ZN(n3570) );
  NAND2_X1 U3643 ( .A1(b_3_), .A2(a_9_), .ZN(n3650) );
  INV_X1 U3644 ( .A(n3651), .ZN(n3649) );
  XNOR2_X1 U3645 ( .A(n3652), .B(n3653), .ZN(n3568) );
  NAND2_X1 U3646 ( .A1(n3654), .A2(n3655), .ZN(n3652) );
  NAND2_X1 U3647 ( .A1(a_9_), .A2(n3651), .ZN(n3569) );
  NAND2_X1 U3648 ( .A1(n3534), .A2(n3656), .ZN(n3651) );
  NAND2_X1 U3649 ( .A1(n3533), .A2(n3535), .ZN(n3656) );
  NAND2_X1 U3650 ( .A1(n3657), .A2(n3658), .ZN(n3535) );
  NAND2_X1 U3651 ( .A1(b_3_), .A2(a_10_), .ZN(n3658) );
  INV_X1 U3652 ( .A(n3659), .ZN(n3657) );
  XNOR2_X1 U3653 ( .A(n3660), .B(n3661), .ZN(n3533) );
  XNOR2_X1 U3654 ( .A(n3662), .B(n3663), .ZN(n3661) );
  NAND2_X1 U3655 ( .A1(a_10_), .A2(n3659), .ZN(n3534) );
  NAND2_X1 U3656 ( .A1(n3565), .A2(n3664), .ZN(n3659) );
  NAND2_X1 U3657 ( .A1(n3564), .A2(n3566), .ZN(n3664) );
  NAND2_X1 U3658 ( .A1(n3665), .A2(n3666), .ZN(n3566) );
  NAND2_X1 U3659 ( .A1(b_3_), .A2(a_11_), .ZN(n3666) );
  INV_X1 U3660 ( .A(n3667), .ZN(n3665) );
  XNOR2_X1 U3661 ( .A(n3668), .B(n3669), .ZN(n3564) );
  XNOR2_X1 U3662 ( .A(n3670), .B(n3671), .ZN(n3668) );
  NOR2_X1 U3663 ( .A1(n2003), .A2(n2219), .ZN(n3671) );
  NAND2_X1 U3664 ( .A1(a_11_), .A2(n3667), .ZN(n3565) );
  NAND2_X1 U3665 ( .A1(n3672), .A2(n3673), .ZN(n3667) );
  NAND2_X1 U3666 ( .A1(n3545), .A2(n3674), .ZN(n3673) );
  NAND2_X1 U3667 ( .A1(n3546), .A2(n3544), .ZN(n3674) );
  NOR2_X1 U3668 ( .A1(n2141), .A2(n2003), .ZN(n3545) );
  OR2_X1 U3669 ( .A1(n3544), .A2(n3546), .ZN(n3672) );
  AND2_X1 U3670 ( .A1(n3675), .A2(n3676), .ZN(n3546) );
  NAND3_X1 U3671 ( .A1(a_13_), .A2(n3677), .A3(b_3_), .ZN(n3676) );
  OR2_X1 U3672 ( .A1(n3561), .A2(n3562), .ZN(n3677) );
  NAND2_X1 U3673 ( .A1(n3562), .A2(n3561), .ZN(n3675) );
  NAND2_X1 U3674 ( .A1(n3678), .A2(n3679), .ZN(n3561) );
  NAND2_X1 U3675 ( .A1(b_1_), .A2(n3680), .ZN(n3679) );
  NAND2_X1 U3676 ( .A1(n1964), .A2(n3681), .ZN(n3680) );
  NAND2_X1 U3677 ( .A1(a_15_), .A2(n2219), .ZN(n3681) );
  NAND2_X1 U3678 ( .A1(b_2_), .A2(n3682), .ZN(n3678) );
  NAND2_X1 U3679 ( .A1(n1967), .A2(n3683), .ZN(n3682) );
  NAND2_X1 U3680 ( .A1(a_14_), .A2(n2175), .ZN(n3683) );
  AND3_X1 U3681 ( .A1(b_2_), .A2(b_3_), .A3(n2215), .ZN(n3562) );
  XNOR2_X1 U3682 ( .A(n3684), .B(n3685), .ZN(n3544) );
  NOR2_X1 U3683 ( .A1(n1988), .A2(n2219), .ZN(n3685) );
  XOR2_X1 U3684 ( .A(n3686), .B(n3687), .Z(n3684) );
  XOR2_X1 U3685 ( .A(n3688), .B(n3689), .Z(n3572) );
  XOR2_X1 U3686 ( .A(n3690), .B(n3691), .Z(n3688) );
  XOR2_X1 U3687 ( .A(n3692), .B(n3693), .Z(n3580) );
  XOR2_X1 U3688 ( .A(n3694), .B(n3695), .Z(n3692) );
  XNOR2_X1 U3689 ( .A(n3696), .B(n3697), .ZN(n3513) );
  NAND2_X1 U3690 ( .A1(n3698), .A2(n3699), .ZN(n3696) );
  XNOR2_X1 U3691 ( .A(n3700), .B(n3701), .ZN(n3584) );
  XOR2_X1 U3692 ( .A(n3702), .B(n3703), .Z(n3700) );
  NOR2_X1 U3693 ( .A1(n2139), .A2(n2141), .ZN(n2136) );
  XOR2_X1 U3694 ( .A(n3704), .B(n3705), .Z(n3591) );
  XOR2_X1 U3695 ( .A(n3706), .B(n3707), .Z(n3704) );
  XOR2_X1 U3696 ( .A(n3708), .B(n3709), .Z(n3595) );
  XOR2_X1 U3697 ( .A(n2158), .B(n3710), .Z(n3708) );
  XOR2_X1 U3698 ( .A(n3711), .B(n3712), .Z(n3599) );
  XOR2_X1 U3699 ( .A(n3713), .B(n3714), .Z(n3711) );
  XOR2_X1 U3700 ( .A(n3715), .B(n3611), .Z(n3495) );
  XNOR2_X1 U3701 ( .A(n3716), .B(n3717), .ZN(n3611) );
  NOR2_X1 U3702 ( .A1(n3608), .A2(n2220), .ZN(n3717) );
  NAND2_X1 U3703 ( .A1(n3605), .A2(n2171), .ZN(n3716) );
  NOR2_X1 U3704 ( .A1(n2175), .A2(n2396), .ZN(n2171) );
  AND2_X1 U3705 ( .A1(n3718), .A2(n3719), .ZN(n3605) );
  NAND2_X1 U3706 ( .A1(n3720), .A2(n3721), .ZN(n3719) );
  OR2_X1 U3707 ( .A1(n3722), .A2(n3723), .ZN(n3721) );
  NAND2_X1 U3708 ( .A1(n3723), .A2(n3722), .ZN(n3718) );
  XOR2_X1 U3709 ( .A(n3724), .B(n3609), .Z(n3715) );
  AND2_X1 U3710 ( .A1(n3725), .A2(n3726), .ZN(n3609) );
  NAND2_X1 U3711 ( .A1(n3714), .A2(n3727), .ZN(n3726) );
  OR2_X1 U3712 ( .A1(n3713), .A2(n3712), .ZN(n3727) );
  NOR2_X1 U3713 ( .A1(n2219), .A2(n2396), .ZN(n3714) );
  NAND2_X1 U3714 ( .A1(n3712), .A2(n3713), .ZN(n3725) );
  NAND2_X1 U3715 ( .A1(n3728), .A2(n3729), .ZN(n3713) );
  NAND2_X1 U3716 ( .A1(n3709), .A2(n3730), .ZN(n3729) );
  NAND2_X1 U3717 ( .A1(n3710), .A2(n2158), .ZN(n3730) );
  XOR2_X1 U3718 ( .A(n3731), .B(n3732), .Z(n3709) );
  NOR2_X1 U3719 ( .A1(n2139), .A2(n2175), .ZN(n3732) );
  XOR2_X1 U3720 ( .A(n3733), .B(n3734), .Z(n3731) );
  OR2_X1 U3721 ( .A1(n2158), .A2(n3710), .ZN(n3728) );
  AND2_X1 U3722 ( .A1(n3735), .A2(n3736), .ZN(n3710) );
  NAND2_X1 U3723 ( .A1(n3707), .A2(n3737), .ZN(n3736) );
  OR2_X1 U3724 ( .A1(n3706), .A2(n3705), .ZN(n3737) );
  NOR2_X1 U3725 ( .A1(n2219), .A2(n2139), .ZN(n3707) );
  NAND2_X1 U3726 ( .A1(n3705), .A2(n3706), .ZN(n3735) );
  NAND2_X1 U3727 ( .A1(n3626), .A2(n3738), .ZN(n3706) );
  NAND2_X1 U3728 ( .A1(n3625), .A2(n3627), .ZN(n3738) );
  NAND2_X1 U3729 ( .A1(n3739), .A2(n3740), .ZN(n3627) );
  NAND2_X1 U3730 ( .A1(b_2_), .A2(a_4_), .ZN(n3740) );
  INV_X1 U3731 ( .A(n3741), .ZN(n3739) );
  XOR2_X1 U3732 ( .A(n3742), .B(n3743), .Z(n3625) );
  NOR2_X1 U3733 ( .A1(n2104), .A2(n2175), .ZN(n3743) );
  XOR2_X1 U3734 ( .A(n3744), .B(n3745), .Z(n3742) );
  NAND2_X1 U3735 ( .A1(a_4_), .A2(n3741), .ZN(n3626) );
  NAND2_X1 U3736 ( .A1(n3746), .A2(n3747), .ZN(n3741) );
  NAND2_X1 U3737 ( .A1(n3703), .A2(n3748), .ZN(n3747) );
  OR2_X1 U3738 ( .A1(n3702), .A2(n3701), .ZN(n3748) );
  NOR2_X1 U3739 ( .A1(n2219), .A2(n2104), .ZN(n3703) );
  NAND2_X1 U3740 ( .A1(n3701), .A2(n3702), .ZN(n3746) );
  NAND2_X1 U3741 ( .A1(n3698), .A2(n3749), .ZN(n3702) );
  NAND2_X1 U3742 ( .A1(n3697), .A2(n3699), .ZN(n3749) );
  NAND2_X1 U3743 ( .A1(n3750), .A2(n3751), .ZN(n3699) );
  NAND2_X1 U3744 ( .A1(b_2_), .A2(a_6_), .ZN(n3751) );
  INV_X1 U3745 ( .A(n3752), .ZN(n3750) );
  XOR2_X1 U3746 ( .A(n3753), .B(n3754), .Z(n3697) );
  NOR2_X1 U3747 ( .A1(n2076), .A2(n2175), .ZN(n3754) );
  XOR2_X1 U3748 ( .A(n3755), .B(n3756), .Z(n3753) );
  NAND2_X1 U3749 ( .A1(a_6_), .A2(n3752), .ZN(n3698) );
  NAND2_X1 U3750 ( .A1(n3757), .A2(n3758), .ZN(n3752) );
  NAND2_X1 U3751 ( .A1(n3695), .A2(n3759), .ZN(n3758) );
  OR2_X1 U3752 ( .A1(n3694), .A2(n3693), .ZN(n3759) );
  NOR2_X1 U3753 ( .A1(n2219), .A2(n2076), .ZN(n3695) );
  NAND2_X1 U3754 ( .A1(n3693), .A2(n3694), .ZN(n3757) );
  NAND2_X1 U3755 ( .A1(n3643), .A2(n3760), .ZN(n3694) );
  NAND2_X1 U3756 ( .A1(n3642), .A2(n3644), .ZN(n3760) );
  NAND2_X1 U3757 ( .A1(n3761), .A2(n3762), .ZN(n3644) );
  NAND2_X1 U3758 ( .A1(b_2_), .A2(a_8_), .ZN(n3762) );
  INV_X1 U3759 ( .A(n3763), .ZN(n3761) );
  XOR2_X1 U3760 ( .A(n3764), .B(n3765), .Z(n3642) );
  NOR2_X1 U3761 ( .A1(n2046), .A2(n2175), .ZN(n3765) );
  XOR2_X1 U3762 ( .A(n3766), .B(n3767), .Z(n3764) );
  NAND2_X1 U3763 ( .A1(a_8_), .A2(n3763), .ZN(n3643) );
  NAND2_X1 U3764 ( .A1(n3768), .A2(n3769), .ZN(n3763) );
  NAND2_X1 U3765 ( .A1(n3691), .A2(n3770), .ZN(n3769) );
  OR2_X1 U3766 ( .A1(n3690), .A2(n3689), .ZN(n3770) );
  NOR2_X1 U3767 ( .A1(n2219), .A2(n2046), .ZN(n3691) );
  NAND2_X1 U3768 ( .A1(n3689), .A2(n3690), .ZN(n3768) );
  NAND2_X1 U3769 ( .A1(n3654), .A2(n3771), .ZN(n3690) );
  NAND2_X1 U3770 ( .A1(n3653), .A2(n3655), .ZN(n3771) );
  NAND2_X1 U3771 ( .A1(n3772), .A2(n3773), .ZN(n3655) );
  NAND2_X1 U3772 ( .A1(b_2_), .A2(a_10_), .ZN(n3773) );
  INV_X1 U3773 ( .A(n3774), .ZN(n3772) );
  XOR2_X1 U3774 ( .A(n3775), .B(n3776), .Z(n3653) );
  NOR2_X1 U3775 ( .A1(n2019), .A2(n2175), .ZN(n3776) );
  XOR2_X1 U3776 ( .A(n3777), .B(n3778), .Z(n3775) );
  NAND2_X1 U3777 ( .A1(a_10_), .A2(n3774), .ZN(n3654) );
  NAND2_X1 U3778 ( .A1(n3779), .A2(n3780), .ZN(n3774) );
  NAND2_X1 U3779 ( .A1(n3663), .A2(n3781), .ZN(n3780) );
  OR2_X1 U3780 ( .A1(n3662), .A2(n3660), .ZN(n3781) );
  NOR2_X1 U3781 ( .A1(n2219), .A2(n2019), .ZN(n3663) );
  NAND2_X1 U3782 ( .A1(n3660), .A2(n3662), .ZN(n3779) );
  NAND2_X1 U3783 ( .A1(n3782), .A2(n3783), .ZN(n3662) );
  NAND3_X1 U3784 ( .A1(a_12_), .A2(n3784), .A3(b_2_), .ZN(n3783) );
  NAND2_X1 U3785 ( .A1(n3669), .A2(n3670), .ZN(n3784) );
  OR2_X1 U3786 ( .A1(n3669), .A2(n3670), .ZN(n3782) );
  AND2_X1 U3787 ( .A1(n3785), .A2(n3786), .ZN(n3670) );
  NAND3_X1 U3788 ( .A1(a_13_), .A2(n3787), .A3(b_2_), .ZN(n3786) );
  OR2_X1 U3789 ( .A1(n3686), .A2(n3687), .ZN(n3787) );
  NAND2_X1 U3790 ( .A1(n3687), .A2(n3686), .ZN(n3785) );
  NAND2_X1 U3791 ( .A1(n3788), .A2(n3789), .ZN(n3686) );
  NAND2_X1 U3792 ( .A1(b_0_), .A2(n3790), .ZN(n3789) );
  NAND2_X1 U3793 ( .A1(n3791), .A2(n1964), .ZN(n3790) );
  NAND2_X1 U3794 ( .A1(a_15_), .A2(n3792), .ZN(n1964) );
  NAND2_X1 U3795 ( .A1(a_15_), .A2(n2175), .ZN(n3791) );
  NAND2_X1 U3796 ( .A1(b_1_), .A2(n3793), .ZN(n3788) );
  NAND2_X1 U3797 ( .A1(n3794), .A2(n1967), .ZN(n3793) );
  NAND2_X1 U3798 ( .A1(a_14_), .A2(n1973), .ZN(n1967) );
  NAND2_X1 U3799 ( .A1(a_14_), .A2(n3608), .ZN(n3794) );
  AND3_X1 U3800 ( .A1(b_2_), .A2(b_1_), .A3(n2215), .ZN(n3687) );
  XOR2_X1 U3801 ( .A(n3795), .B(n3796), .Z(n3669) );
  XNOR2_X1 U3802 ( .A(n3797), .B(n3798), .ZN(n3796) );
  NAND2_X1 U3803 ( .A1(a_14_), .A2(b_0_), .ZN(n3795) );
  XNOR2_X1 U3804 ( .A(n3799), .B(n3800), .ZN(n3660) );
  NAND2_X1 U3805 ( .A1(n3801), .A2(n3802), .ZN(n3799) );
  NAND2_X1 U3806 ( .A1(n3803), .A2(n3804), .ZN(n3802) );
  NAND2_X1 U3807 ( .A1(b_1_), .A2(a_12_), .ZN(n3803) );
  XOR2_X1 U3808 ( .A(n3805), .B(n3806), .Z(n3689) );
  XNOR2_X1 U3809 ( .A(n3807), .B(n3808), .ZN(n3806) );
  NAND2_X1 U3810 ( .A1(b_1_), .A2(a_10_), .ZN(n3805) );
  XOR2_X1 U3811 ( .A(n3809), .B(n3810), .Z(n3693) );
  XNOR2_X1 U3812 ( .A(n3811), .B(n3812), .ZN(n3810) );
  NAND2_X1 U3813 ( .A1(b_1_), .A2(a_8_), .ZN(n3809) );
  XOR2_X1 U3814 ( .A(n3813), .B(n3814), .Z(n3701) );
  XNOR2_X1 U3815 ( .A(n3815), .B(n3816), .ZN(n3814) );
  NAND2_X1 U3816 ( .A1(b_1_), .A2(a_6_), .ZN(n3813) );
  XOR2_X1 U3817 ( .A(n3817), .B(n3818), .Z(n3705) );
  XNOR2_X1 U3818 ( .A(n3819), .B(n3820), .ZN(n3818) );
  NAND2_X1 U3819 ( .A1(b_1_), .A2(a_4_), .ZN(n3817) );
  NAND2_X1 U3820 ( .A1(b_2_), .A2(a_2_), .ZN(n2158) );
  XNOR2_X1 U3821 ( .A(n3720), .B(n3821), .ZN(n3712) );
  XNOR2_X1 U3822 ( .A(n3723), .B(n3722), .ZN(n3821) );
  NAND2_X1 U3823 ( .A1(n3822), .A2(n3823), .ZN(n3722) );
  NAND3_X1 U3824 ( .A1(a_3_), .A2(n3824), .A3(b_1_), .ZN(n3823) );
  OR2_X1 U3825 ( .A1(n3734), .A2(n3733), .ZN(n3824) );
  NAND2_X1 U3826 ( .A1(n3733), .A2(n3734), .ZN(n3822) );
  NAND2_X1 U3827 ( .A1(n3825), .A2(n3826), .ZN(n3734) );
  NAND3_X1 U3828 ( .A1(a_4_), .A2(n3827), .A3(b_1_), .ZN(n3826) );
  OR2_X1 U3829 ( .A1(n3820), .A2(n3819), .ZN(n3827) );
  NAND2_X1 U3830 ( .A1(n3819), .A2(n3820), .ZN(n3825) );
  NAND2_X1 U3831 ( .A1(n3828), .A2(n3829), .ZN(n3820) );
  NAND3_X1 U3832 ( .A1(a_5_), .A2(n3830), .A3(b_1_), .ZN(n3829) );
  OR2_X1 U3833 ( .A1(n3745), .A2(n3744), .ZN(n3830) );
  NAND2_X1 U3834 ( .A1(n3744), .A2(n3745), .ZN(n3828) );
  NAND2_X1 U3835 ( .A1(n3831), .A2(n3832), .ZN(n3745) );
  NAND3_X1 U3836 ( .A1(a_6_), .A2(n3833), .A3(b_1_), .ZN(n3832) );
  OR2_X1 U3837 ( .A1(n3816), .A2(n3815), .ZN(n3833) );
  NAND2_X1 U3838 ( .A1(n3815), .A2(n3816), .ZN(n3831) );
  NAND2_X1 U3839 ( .A1(n3834), .A2(n3835), .ZN(n3816) );
  NAND3_X1 U3840 ( .A1(a_7_), .A2(n3836), .A3(b_1_), .ZN(n3835) );
  OR2_X1 U3841 ( .A1(n3756), .A2(n3755), .ZN(n3836) );
  NAND2_X1 U3842 ( .A1(n3755), .A2(n3756), .ZN(n3834) );
  NAND2_X1 U3843 ( .A1(n3837), .A2(n3838), .ZN(n3756) );
  NAND3_X1 U3844 ( .A1(a_8_), .A2(n3839), .A3(b_1_), .ZN(n3838) );
  OR2_X1 U3845 ( .A1(n3812), .A2(n3811), .ZN(n3839) );
  NAND2_X1 U3846 ( .A1(n3811), .A2(n3812), .ZN(n3837) );
  NAND2_X1 U3847 ( .A1(n3840), .A2(n3841), .ZN(n3812) );
  NAND3_X1 U3848 ( .A1(a_9_), .A2(n3842), .A3(b_1_), .ZN(n3841) );
  OR2_X1 U3849 ( .A1(n3767), .A2(n3766), .ZN(n3842) );
  NAND2_X1 U3850 ( .A1(n3766), .A2(n3767), .ZN(n3840) );
  NAND2_X1 U3851 ( .A1(n3843), .A2(n3844), .ZN(n3767) );
  NAND3_X1 U3852 ( .A1(a_10_), .A2(n3845), .A3(b_1_), .ZN(n3844) );
  OR2_X1 U3853 ( .A1(n3808), .A2(n3807), .ZN(n3845) );
  NAND2_X1 U3854 ( .A1(n3807), .A2(n3808), .ZN(n3843) );
  NAND2_X1 U3855 ( .A1(n3846), .A2(n3847), .ZN(n3808) );
  NAND3_X1 U3856 ( .A1(a_11_), .A2(n3848), .A3(b_1_), .ZN(n3847) );
  OR2_X1 U3857 ( .A1(n3778), .A2(n3777), .ZN(n3848) );
  NAND2_X1 U3858 ( .A1(n3777), .A2(n3778), .ZN(n3846) );
  NAND2_X1 U3859 ( .A1(n3801), .A2(n3849), .ZN(n3778) );
  NAND2_X1 U3860 ( .A1(n3850), .A2(n3800), .ZN(n3849) );
  NAND2_X1 U3861 ( .A1(n3798), .A2(n3851), .ZN(n3800) );
  NAND3_X1 U3862 ( .A1(a_14_), .A2(b_0_), .A3(n3797), .ZN(n3851) );
  NOR2_X1 U3863 ( .A1(n2175), .A2(n1988), .ZN(n3797) );
  NAND3_X1 U3864 ( .A1(b_1_), .A2(b_0_), .A3(n2215), .ZN(n3798) );
  NAND2_X1 U3865 ( .A1(n3804), .A2(n2003), .ZN(n3850) );
  OR3_X1 U3866 ( .A1(n2175), .A2(n2003), .A3(n3804), .ZN(n3801) );
  NAND2_X1 U3867 ( .A1(a_13_), .A2(b_0_), .ZN(n3804) );
  NOR2_X1 U3868 ( .A1(n2003), .A2(n3608), .ZN(n3777) );
  NOR2_X1 U3869 ( .A1(n2019), .A2(n3608), .ZN(n3807) );
  NOR2_X1 U3870 ( .A1(n2586), .A2(n3608), .ZN(n3766) );
  NOR2_X1 U3871 ( .A1(n2046), .A2(n3608), .ZN(n3811) );
  NOR2_X1 U3872 ( .A1(n2218), .A2(n3608), .ZN(n3755) );
  NOR2_X1 U3873 ( .A1(n2076), .A2(n3608), .ZN(n3815) );
  NOR2_X1 U3874 ( .A1(n2089), .A2(n3608), .ZN(n3744) );
  NOR2_X1 U3875 ( .A1(n2104), .A2(n3608), .ZN(n3819) );
  NOR2_X1 U3876 ( .A1(n2119), .A2(n3608), .ZN(n3733) );
  NOR2_X1 U3877 ( .A1(n2139), .A2(n3608), .ZN(n3723) );
  NOR2_X1 U3878 ( .A1(n2175), .A2(n2220), .ZN(n3720) );
  NAND2_X1 U3879 ( .A1(a_0_), .A2(b_2_), .ZN(n3724) );
  NAND2_X1 U3880 ( .A1(n3852), .A2(n3853), .ZN(n1957) );
  NAND2_X1 U3881 ( .A1(n3854), .A2(n2185), .ZN(n3853) );
  NAND2_X1 U3882 ( .A1(b_0_), .A2(n2407), .ZN(n2185) );
  INV_X1 U3883 ( .A(a_0_), .ZN(n2407) );
  NAND2_X1 U3884 ( .A1(n3855), .A2(n3856), .ZN(n3854) );
  NAND2_X1 U3885 ( .A1(a_1_), .A2(n2175), .ZN(n3856) );
  INV_X1 U3886 ( .A(b_1_), .ZN(n2175) );
  NAND3_X1 U3887 ( .A1(n3857), .A2(n3858), .A3(n3859), .ZN(n3855) );
  NAND2_X1 U3888 ( .A1(b_2_), .A2(n2220), .ZN(n3859) );
  INV_X1 U3889 ( .A(a_2_), .ZN(n2220) );
  NAND3_X1 U3890 ( .A1(n3860), .A2(n3861), .A3(n3862), .ZN(n3858) );
  NAND2_X1 U3891 ( .A1(a_3_), .A2(n2141), .ZN(n3862) );
  INV_X1 U3892 ( .A(b_3_), .ZN(n2141) );
  NAND3_X1 U3893 ( .A1(n3863), .A2(n3864), .A3(n3865), .ZN(n3861) );
  NAND2_X1 U3894 ( .A1(b_4_), .A2(n2119), .ZN(n3865) );
  INV_X1 U3895 ( .A(a_4_), .ZN(n2119) );
  NAND3_X1 U3896 ( .A1(n3866), .A2(n3867), .A3(n3868), .ZN(n3864) );
  NAND2_X1 U3897 ( .A1(a_5_), .A2(n2106), .ZN(n3868) );
  INV_X1 U3898 ( .A(b_5_), .ZN(n2106) );
  NAND3_X1 U3899 ( .A1(n3869), .A2(n3870), .A3(n3871), .ZN(n3867) );
  NAND2_X1 U3900 ( .A1(b_6_), .A2(n2089), .ZN(n3871) );
  INV_X1 U3901 ( .A(a_6_), .ZN(n2089) );
  NAND3_X1 U3902 ( .A1(n3872), .A2(n3873), .A3(n3874), .ZN(n3870) );
  NAND2_X1 U3903 ( .A1(a_7_), .A2(n2074), .ZN(n3874) );
  INV_X1 U3904 ( .A(b_7_), .ZN(n2074) );
  NAND3_X1 U3905 ( .A1(n3875), .A2(n3876), .A3(n3877), .ZN(n3873) );
  NAND2_X1 U3906 ( .A1(b_8_), .A2(n2218), .ZN(n3877) );
  INV_X1 U3907 ( .A(a_8_), .ZN(n2218) );
  NAND3_X1 U3908 ( .A1(n3878), .A2(n3879), .A3(n3880), .ZN(n3876) );
  NAND2_X1 U3909 ( .A1(a_9_), .A2(n2048), .ZN(n3880) );
  INV_X1 U3910 ( .A(b_9_), .ZN(n2048) );
  NAND3_X1 U3911 ( .A1(n3881), .A2(n3882), .A3(n3883), .ZN(n3879) );
  NAND2_X1 U3912 ( .A1(b_9_), .A2(n2046), .ZN(n3883) );
  INV_X1 U3913 ( .A(a_9_), .ZN(n2046) );
  NAND3_X1 U3914 ( .A1(n3884), .A2(n3885), .A3(n3886), .ZN(n3882) );
  NAND2_X1 U3915 ( .A1(a_11_), .A2(n2017), .ZN(n3886) );
  INV_X1 U3916 ( .A(b_11_), .ZN(n2017) );
  NAND3_X1 U3917 ( .A1(n3887), .A2(n3888), .A3(n3889), .ZN(n3885) );
  NAND2_X1 U3918 ( .A1(b_12_), .A2(n2003), .ZN(n3889) );
  INV_X1 U3919 ( .A(a_12_), .ZN(n2003) );
  NAND3_X1 U3920 ( .A1(n3890), .A2(n3891), .A3(n3892), .ZN(n3888) );
  NAND2_X1 U3921 ( .A1(a_13_), .A2(n1990), .ZN(n3892) );
  INV_X1 U3922 ( .A(b_13_), .ZN(n1990) );
  NAND4_X1 U3923 ( .A1(n3893), .A2(n3894), .A3(n3895), .A4(n3896), .ZN(n3891)
         );
  INV_X1 U3924 ( .A(n2214), .ZN(n3896) );
  NOR2_X1 U3925 ( .A1(n1955), .A2(n1969), .ZN(n2214) );
  NAND2_X1 U3926 ( .A1(n1965), .A2(n3792), .ZN(n3895) );
  NAND2_X1 U3927 ( .A1(a_15_), .A2(n1955), .ZN(n1965) );
  INV_X1 U3928 ( .A(b_15_), .ZN(n1955) );
  OR2_X1 U3929 ( .A1(n1969), .A2(n2215), .ZN(n3894) );
  INV_X1 U3930 ( .A(a_15_), .ZN(n1973) );
  INV_X1 U3931 ( .A(a_14_), .ZN(n3792) );
  INV_X1 U3932 ( .A(b_14_), .ZN(n1969) );
  NAND2_X1 U3933 ( .A1(b_13_), .A2(n1988), .ZN(n3893) );
  INV_X1 U3934 ( .A(a_13_), .ZN(n1988) );
  NAND2_X1 U3935 ( .A1(a_12_), .A2(n2216), .ZN(n3890) );
  INV_X1 U3936 ( .A(b_12_), .ZN(n2216) );
  NAND2_X1 U3937 ( .A1(b_11_), .A2(n2019), .ZN(n3887) );
  INV_X1 U3938 ( .A(a_11_), .ZN(n2019) );
  NAND2_X1 U3939 ( .A1(a_10_), .A2(n2691), .ZN(n3884) );
  INV_X1 U3940 ( .A(b_10_), .ZN(n2691) );
  NAND2_X1 U3941 ( .A1(b_10_), .A2(n2586), .ZN(n3881) );
  INV_X1 U3942 ( .A(a_10_), .ZN(n2586) );
  NAND2_X1 U3943 ( .A1(a_8_), .A2(n2217), .ZN(n3878) );
  INV_X1 U3944 ( .A(b_8_), .ZN(n2217) );
  NAND2_X1 U3945 ( .A1(b_7_), .A2(n2076), .ZN(n3875) );
  INV_X1 U3946 ( .A(a_7_), .ZN(n2076) );
  NAND2_X1 U3947 ( .A1(a_6_), .A2(n3124), .ZN(n3872) );
  INV_X1 U3948 ( .A(b_6_), .ZN(n3124) );
  NAND2_X1 U3949 ( .A1(b_5_), .A2(n2104), .ZN(n3869) );
  INV_X1 U3950 ( .A(a_5_), .ZN(n2104) );
  NAND2_X1 U3951 ( .A1(a_4_), .A2(n3351), .ZN(n3866) );
  INV_X1 U3952 ( .A(b_4_), .ZN(n3351) );
  NAND2_X1 U3953 ( .A1(b_3_), .A2(n2139), .ZN(n3863) );
  INV_X1 U3954 ( .A(a_3_), .ZN(n2139) );
  NAND2_X1 U3955 ( .A1(a_2_), .A2(n2219), .ZN(n3860) );
  INV_X1 U3956 ( .A(b_2_), .ZN(n2219) );
  NAND2_X1 U3957 ( .A1(b_1_), .A2(n2396), .ZN(n3857) );
  INV_X1 U3958 ( .A(a_1_), .ZN(n2396) );
  NAND2_X1 U3959 ( .A1(a_0_), .A2(n3608), .ZN(n3852) );
  INV_X1 U3960 ( .A(b_0_), .ZN(n3608) );
endmodule

