module add_mul_comp_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, Result_0_, Result_1_, 
        Result_2_, Result_3_, Result_4_, Result_5_, Result_6_, Result_7_, 
        Result_8_, Result_9_, Result_10_, Result_11_, Result_12_, Result_13_, 
        Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992;

  OR2_X1 U505 ( .A1(n489), .A2(n490), .ZN(Result_9_) );
  AND2_X1 U506 ( .A1(n491), .A2(n492), .ZN(n490) );
  XNOR2_X1 U507 ( .A(n493), .B(n494), .ZN(n491) );
  XOR2_X1 U508 ( .A(n495), .B(n496), .Z(n494) );
  AND2_X1 U509 ( .A1(n497), .A2(n498), .ZN(n489) );
  XNOR2_X1 U510 ( .A(n499), .B(n500), .ZN(n497) );
  AND2_X1 U511 ( .A1(n501), .A2(n502), .ZN(n500) );
  INV_X1 U512 ( .A(n503), .ZN(n501) );
  OR2_X1 U513 ( .A1(n504), .A2(n505), .ZN(Result_8_) );
  AND2_X1 U514 ( .A1(n506), .A2(n492), .ZN(n505) );
  XNOR2_X1 U515 ( .A(n507), .B(n508), .ZN(n506) );
  XOR2_X1 U516 ( .A(n509), .B(n510), .Z(n508) );
  AND2_X1 U517 ( .A1(n511), .A2(n498), .ZN(n504) );
  XOR2_X1 U518 ( .A(n512), .B(n513), .Z(n511) );
  AND2_X1 U519 ( .A1(n514), .A2(n515), .ZN(n512) );
  OR2_X1 U520 ( .A1(n499), .A2(n516), .ZN(n515) );
  AND2_X1 U521 ( .A1(n517), .A2(n518), .ZN(n499) );
  INV_X1 U522 ( .A(n519), .ZN(n517) );
  AND2_X1 U523 ( .A1(n520), .A2(n521), .ZN(n519) );
  OR2_X1 U524 ( .A1(b_1_), .A2(a_1_), .ZN(n514) );
  AND2_X1 U525 ( .A1(n492), .A2(n522), .ZN(Result_7_) );
  XOR2_X1 U526 ( .A(n523), .B(n524), .Z(n522) );
  AND2_X1 U527 ( .A1(n525), .A2(n492), .ZN(Result_6_) );
  AND2_X1 U528 ( .A1(n526), .A2(n527), .ZN(n525) );
  OR2_X1 U529 ( .A1(n528), .A2(n529), .ZN(n526) );
  XOR2_X1 U530 ( .A(n530), .B(n531), .Z(n529) );
  INV_X1 U531 ( .A(n532), .ZN(n528) );
  AND2_X1 U532 ( .A1(n492), .A2(n533), .ZN(Result_5_) );
  XOR2_X1 U533 ( .A(n534), .B(n535), .Z(n533) );
  OR2_X1 U534 ( .A1(n536), .A2(n537), .ZN(n534) );
  AND2_X1 U535 ( .A1(n538), .A2(n492), .ZN(Result_4_) );
  XOR2_X1 U536 ( .A(n539), .B(n540), .Z(n538) );
  AND2_X1 U537 ( .A1(n492), .A2(n541), .ZN(Result_3_) );
  XOR2_X1 U538 ( .A(n542), .B(n543), .Z(n541) );
  AND2_X1 U539 ( .A1(n544), .A2(n545), .ZN(n543) );
  OR2_X1 U540 ( .A1(n546), .A2(n547), .ZN(n545) );
  INV_X1 U541 ( .A(n548), .ZN(n544) );
  AND2_X1 U542 ( .A1(n549), .A2(n492), .ZN(Result_2_) );
  XOR2_X1 U543 ( .A(n550), .B(n551), .Z(n549) );
  AND2_X1 U544 ( .A1(n492), .A2(n552), .ZN(Result_1_) );
  XOR2_X1 U545 ( .A(n553), .B(n554), .Z(n552) );
  AND2_X1 U546 ( .A1(n555), .A2(n556), .ZN(n554) );
  OR2_X1 U547 ( .A1(n557), .A2(n558), .ZN(n556) );
  INV_X1 U548 ( .A(n559), .ZN(n555) );
  OR2_X1 U549 ( .A1(n560), .A2(n561), .ZN(Result_15_) );
  AND2_X1 U550 ( .A1(n562), .A2(n498), .ZN(n561) );
  OR2_X1 U551 ( .A1(n563), .A2(n564), .ZN(n562) );
  AND2_X1 U552 ( .A1(b_7_), .A2(n565), .ZN(n563) );
  AND2_X1 U553 ( .A1(n566), .A2(n492), .ZN(n560) );
  OR2_X1 U554 ( .A1(n567), .A2(n568), .ZN(Result_14_) );
  AND2_X1 U555 ( .A1(n569), .A2(n492), .ZN(n568) );
  XNOR2_X1 U556 ( .A(n570), .B(n571), .ZN(n569) );
  AND2_X1 U557 ( .A1(b_7_), .A2(a_6_), .ZN(n571) );
  AND2_X1 U558 ( .A1(n572), .A2(n498), .ZN(n567) );
  XOR2_X1 U559 ( .A(n566), .B(n573), .Z(n572) );
  XNOR2_X1 U560 ( .A(n574), .B(a_6_), .ZN(n573) );
  OR2_X1 U561 ( .A1(n575), .A2(n576), .ZN(Result_13_) );
  AND2_X1 U562 ( .A1(n577), .A2(n492), .ZN(n576) );
  XOR2_X1 U563 ( .A(n578), .B(n579), .Z(n577) );
  XNOR2_X1 U564 ( .A(n580), .B(n581), .ZN(n579) );
  AND2_X1 U565 ( .A1(n582), .A2(n498), .ZN(n575) );
  OR2_X1 U566 ( .A1(n583), .A2(n584), .ZN(n582) );
  OR2_X1 U567 ( .A1(n585), .A2(n586), .ZN(n584) );
  AND2_X1 U568 ( .A1(n587), .A2(n588), .ZN(n586) );
  INV_X1 U569 ( .A(n589), .ZN(n585) );
  OR2_X1 U570 ( .A1(n590), .A2(n588), .ZN(n589) );
  AND2_X1 U571 ( .A1(n591), .A2(n592), .ZN(n583) );
  XNOR2_X1 U572 ( .A(n588), .B(a_5_), .ZN(n591) );
  OR2_X1 U573 ( .A1(n593), .A2(n594), .ZN(Result_12_) );
  AND2_X1 U574 ( .A1(n595), .A2(n492), .ZN(n594) );
  XNOR2_X1 U575 ( .A(n596), .B(n597), .ZN(n595) );
  XOR2_X1 U576 ( .A(n598), .B(n599), .Z(n597) );
  AND2_X1 U577 ( .A1(n600), .A2(n498), .ZN(n593) );
  XNOR2_X1 U578 ( .A(n601), .B(n602), .ZN(n600) );
  AND2_X1 U579 ( .A1(n603), .A2(n604), .ZN(n602) );
  OR2_X1 U580 ( .A1(n605), .A2(n606), .ZN(Result_11_) );
  AND2_X1 U581 ( .A1(n607), .A2(n492), .ZN(n606) );
  XNOR2_X1 U582 ( .A(n608), .B(n609), .ZN(n607) );
  XOR2_X1 U583 ( .A(n610), .B(n611), .Z(n609) );
  AND2_X1 U584 ( .A1(n612), .A2(n498), .ZN(n605) );
  OR2_X1 U585 ( .A1(n613), .A2(n614), .ZN(n612) );
  OR2_X1 U586 ( .A1(n615), .A2(n616), .ZN(n614) );
  AND2_X1 U587 ( .A1(n617), .A2(n618), .ZN(n616) );
  AND2_X1 U588 ( .A1(n619), .A2(n620), .ZN(n615) );
  AND2_X1 U589 ( .A1(n621), .A2(n622), .ZN(n613) );
  XNOR2_X1 U590 ( .A(n623), .B(n617), .ZN(n621) );
  OR2_X1 U591 ( .A1(n624), .A2(n625), .ZN(Result_10_) );
  AND2_X1 U592 ( .A1(n626), .A2(n492), .ZN(n625) );
  XNOR2_X1 U593 ( .A(n627), .B(n628), .ZN(n626) );
  XOR2_X1 U594 ( .A(n629), .B(n630), .Z(n628) );
  AND2_X1 U595 ( .A1(n631), .A2(n498), .ZN(n624) );
  XNOR2_X1 U596 ( .A(n520), .B(n632), .ZN(n631) );
  AND2_X1 U597 ( .A1(n521), .A2(n518), .ZN(n632) );
  OR2_X1 U598 ( .A1(a_2_), .A2(b_2_), .ZN(n518) );
  OR2_X1 U599 ( .A1(n633), .A2(n634), .ZN(n520) );
  AND2_X1 U600 ( .A1(n623), .A2(n622), .ZN(n634) );
  AND2_X1 U601 ( .A1(n620), .A2(n635), .ZN(n633) );
  INV_X1 U602 ( .A(n617), .ZN(n620) );
  AND2_X1 U603 ( .A1(n636), .A2(n604), .ZN(n617) );
  OR2_X1 U604 ( .A1(a_4_), .A2(b_4_), .ZN(n604) );
  INV_X1 U605 ( .A(n637), .ZN(n636) );
  AND2_X1 U606 ( .A1(n601), .A2(n603), .ZN(n637) );
  OR2_X1 U607 ( .A1(n638), .A2(n639), .ZN(n601) );
  AND2_X1 U608 ( .A1(n640), .A2(n592), .ZN(n639) );
  AND2_X1 U609 ( .A1(n588), .A2(n590), .ZN(n638) );
  AND2_X1 U610 ( .A1(n641), .A2(n642), .ZN(n588) );
  OR2_X1 U611 ( .A1(n643), .A2(n570), .ZN(n642) );
  INV_X1 U612 ( .A(n644), .ZN(n641) );
  AND2_X1 U613 ( .A1(a_6_), .A2(n645), .ZN(n644) );
  OR2_X1 U614 ( .A1(n566), .A2(b_6_), .ZN(n645) );
  AND2_X1 U615 ( .A1(a_7_), .A2(b_7_), .ZN(n566) );
  AND2_X1 U616 ( .A1(n492), .A2(n646), .ZN(Result_0_) );
  OR2_X1 U617 ( .A1(n647), .A2(n648), .ZN(n646) );
  OR2_X1 U618 ( .A1(n559), .A2(n649), .ZN(n648) );
  AND2_X1 U619 ( .A1(n650), .A2(b_0_), .ZN(n649) );
  INV_X1 U620 ( .A(n651), .ZN(n650) );
  AND2_X1 U621 ( .A1(n557), .A2(n558), .ZN(n559) );
  AND2_X1 U622 ( .A1(n652), .A2(n653), .ZN(n558) );
  AND2_X1 U623 ( .A1(n553), .A2(n557), .ZN(n647) );
  AND2_X1 U624 ( .A1(n651), .A2(b_0_), .ZN(n557) );
  AND2_X1 U625 ( .A1(n550), .A2(n551), .ZN(n553) );
  XOR2_X1 U626 ( .A(n653), .B(n652), .Z(n551) );
  OR2_X1 U627 ( .A1(n654), .A2(n655), .ZN(n652) );
  OR2_X1 U628 ( .A1(n656), .A2(n657), .ZN(n655) );
  INV_X1 U629 ( .A(n658), .ZN(n657) );
  XNOR2_X1 U630 ( .A(n651), .B(n659), .ZN(n654) );
  AND2_X1 U631 ( .A1(b_0_), .A2(a_1_), .ZN(n659) );
  OR2_X1 U632 ( .A1(n660), .A2(n661), .ZN(n651) );
  OR2_X1 U633 ( .A1(n662), .A2(n663), .ZN(n653) );
  AND2_X1 U634 ( .A1(n664), .A2(n665), .ZN(n663) );
  OR2_X1 U635 ( .A1(n666), .A2(n667), .ZN(n550) );
  OR2_X1 U636 ( .A1(n668), .A2(n548), .ZN(n666) );
  AND2_X1 U637 ( .A1(n546), .A2(n547), .ZN(n548) );
  AND2_X1 U638 ( .A1(n669), .A2(n670), .ZN(n547) );
  INV_X1 U639 ( .A(n671), .ZN(n669) );
  AND2_X1 U640 ( .A1(n542), .A2(n546), .ZN(n668) );
  INV_X1 U641 ( .A(n672), .ZN(n546) );
  OR2_X1 U642 ( .A1(n673), .A2(n667), .ZN(n672) );
  INV_X1 U643 ( .A(n674), .ZN(n667) );
  OR2_X1 U644 ( .A1(n675), .A2(n676), .ZN(n674) );
  AND2_X1 U645 ( .A1(n675), .A2(n676), .ZN(n673) );
  OR2_X1 U646 ( .A1(n677), .A2(n678), .ZN(n676) );
  AND2_X1 U647 ( .A1(n679), .A2(n680), .ZN(n678) );
  AND2_X1 U648 ( .A1(n681), .A2(n682), .ZN(n677) );
  OR2_X1 U649 ( .A1(n680), .A2(n679), .ZN(n682) );
  XNOR2_X1 U650 ( .A(n665), .B(n683), .ZN(n675) );
  XOR2_X1 U651 ( .A(n662), .B(n664), .Z(n683) );
  AND2_X1 U652 ( .A1(b_2_), .A2(a_0_), .ZN(n664) );
  INV_X1 U653 ( .A(n684), .ZN(n662) );
  OR2_X1 U654 ( .A1(n685), .A2(n686), .ZN(n684) );
  AND2_X1 U655 ( .A1(n687), .A2(n688), .ZN(n686) );
  AND2_X1 U656 ( .A1(n689), .A2(n690), .ZN(n685) );
  OR2_X1 U657 ( .A1(n688), .A2(n687), .ZN(n690) );
  XOR2_X1 U658 ( .A(n691), .B(n658), .Z(n665) );
  OR2_X1 U659 ( .A1(n692), .A2(n693), .ZN(n658) );
  AND2_X1 U660 ( .A1(n694), .A2(n695), .ZN(n693) );
  AND2_X1 U661 ( .A1(n696), .A2(n697), .ZN(n692) );
  OR2_X1 U662 ( .A1(n695), .A2(n694), .ZN(n696) );
  OR2_X1 U663 ( .A1(n698), .A2(n656), .ZN(n691) );
  AND2_X1 U664 ( .A1(n516), .A2(n699), .ZN(n656) );
  AND2_X1 U665 ( .A1(a_2_), .A2(b_0_), .ZN(n699) );
  AND2_X1 U666 ( .A1(n700), .A2(n701), .ZN(n698) );
  INV_X1 U667 ( .A(n516), .ZN(n701) );
  AND2_X1 U668 ( .A1(b_1_), .A2(a_1_), .ZN(n516) );
  OR2_X1 U669 ( .A1(n702), .A2(n703), .ZN(n700) );
  AND2_X1 U670 ( .A1(n539), .A2(n540), .ZN(n542) );
  XNOR2_X1 U671 ( .A(n670), .B(n671), .ZN(n540) );
  OR2_X1 U672 ( .A1(n704), .A2(n705), .ZN(n671) );
  AND2_X1 U673 ( .A1(n706), .A2(n707), .ZN(n705) );
  AND2_X1 U674 ( .A1(n708), .A2(n709), .ZN(n704) );
  OR2_X1 U675 ( .A1(n707), .A2(n706), .ZN(n709) );
  XOR2_X1 U676 ( .A(n710), .B(n681), .Z(n670) );
  XOR2_X1 U677 ( .A(n689), .B(n711), .Z(n681) );
  XOR2_X1 U678 ( .A(n688), .B(n687), .Z(n711) );
  OR2_X1 U679 ( .A1(n712), .A2(n713), .ZN(n687) );
  OR2_X1 U680 ( .A1(n714), .A2(n715), .ZN(n688) );
  AND2_X1 U681 ( .A1(n716), .A2(n521), .ZN(n715) );
  AND2_X1 U682 ( .A1(n717), .A2(n718), .ZN(n714) );
  OR2_X1 U683 ( .A1(n521), .A2(n716), .ZN(n718) );
  XOR2_X1 U684 ( .A(n694), .B(n719), .Z(n689) );
  XOR2_X1 U685 ( .A(n695), .B(n697), .Z(n719) );
  OR2_X1 U686 ( .A1(n623), .A2(n703), .ZN(n697) );
  OR2_X1 U687 ( .A1(n720), .A2(n721), .ZN(n695) );
  AND2_X1 U688 ( .A1(n722), .A2(n723), .ZN(n721) );
  AND2_X1 U689 ( .A1(n724), .A2(n725), .ZN(n720) );
  OR2_X1 U690 ( .A1(n723), .A2(n722), .ZN(n724) );
  OR2_X1 U691 ( .A1(n660), .A2(n702), .ZN(n694) );
  XNOR2_X1 U692 ( .A(n680), .B(n679), .ZN(n710) );
  OR2_X1 U693 ( .A1(n726), .A2(n727), .ZN(n679) );
  AND2_X1 U694 ( .A1(n728), .A2(n729), .ZN(n727) );
  AND2_X1 U695 ( .A1(n730), .A2(n731), .ZN(n726) );
  OR2_X1 U696 ( .A1(n729), .A2(n728), .ZN(n731) );
  OR2_X1 U697 ( .A1(n622), .A2(n661), .ZN(n680) );
  OR2_X1 U698 ( .A1(n732), .A2(n733), .ZN(n539) );
  INV_X1 U699 ( .A(n734), .ZN(n733) );
  OR2_X1 U700 ( .A1(n735), .A2(n736), .ZN(n732) );
  AND2_X1 U701 ( .A1(n536), .A2(n535), .ZN(n736) );
  AND2_X1 U702 ( .A1(n537), .A2(n535), .ZN(n735) );
  AND2_X1 U703 ( .A1(n737), .A2(n734), .ZN(n535) );
  OR2_X1 U704 ( .A1(n738), .A2(n739), .ZN(n734) );
  INV_X1 U705 ( .A(n740), .ZN(n737) );
  AND2_X1 U706 ( .A1(n738), .A2(n739), .ZN(n740) );
  OR2_X1 U707 ( .A1(n741), .A2(n742), .ZN(n739) );
  AND2_X1 U708 ( .A1(n743), .A2(n744), .ZN(n742) );
  AND2_X1 U709 ( .A1(n745), .A2(n746), .ZN(n741) );
  OR2_X1 U710 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U711 ( .A(n708), .B(n747), .Z(n738) );
  XOR2_X1 U712 ( .A(n707), .B(n706), .Z(n747) );
  OR2_X1 U713 ( .A1(n748), .A2(n661), .ZN(n706) );
  OR2_X1 U714 ( .A1(n749), .A2(n750), .ZN(n707) );
  AND2_X1 U715 ( .A1(n751), .A2(n752), .ZN(n750) );
  AND2_X1 U716 ( .A1(n753), .A2(n754), .ZN(n749) );
  OR2_X1 U717 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U718 ( .A(n755), .B(n730), .ZN(n708) );
  XNOR2_X1 U719 ( .A(n756), .B(n717), .ZN(n730) );
  XOR2_X1 U720 ( .A(n722), .B(n757), .Z(n717) );
  XOR2_X1 U721 ( .A(n723), .B(n725), .Z(n757) );
  OR2_X1 U722 ( .A1(n660), .A2(n623), .ZN(n725) );
  OR2_X1 U723 ( .A1(n758), .A2(n759), .ZN(n723) );
  AND2_X1 U724 ( .A1(n760), .A2(n761), .ZN(n759) );
  AND2_X1 U725 ( .A1(n762), .A2(n763), .ZN(n758) );
  OR2_X1 U726 ( .A1(n761), .A2(n760), .ZN(n763) );
  OR2_X1 U727 ( .A1(n764), .A2(n703), .ZN(n722) );
  XNOR2_X1 U728 ( .A(n521), .B(n716), .ZN(n756) );
  OR2_X1 U729 ( .A1(n765), .A2(n766), .ZN(n716) );
  AND2_X1 U730 ( .A1(n767), .A2(n768), .ZN(n766) );
  AND2_X1 U731 ( .A1(n769), .A2(n770), .ZN(n765) );
  OR2_X1 U732 ( .A1(n768), .A2(n767), .ZN(n770) );
  OR2_X1 U733 ( .A1(n712), .A2(n702), .ZN(n521) );
  XNOR2_X1 U734 ( .A(n729), .B(n728), .ZN(n755) );
  OR2_X1 U735 ( .A1(n771), .A2(n772), .ZN(n728) );
  AND2_X1 U736 ( .A1(n773), .A2(n774), .ZN(n772) );
  AND2_X1 U737 ( .A1(n775), .A2(n776), .ZN(n771) );
  OR2_X1 U738 ( .A1(n774), .A2(n773), .ZN(n776) );
  OR2_X1 U739 ( .A1(n622), .A2(n713), .ZN(n729) );
  INV_X1 U740 ( .A(n527), .ZN(n537) );
  OR2_X1 U741 ( .A1(n777), .A2(n532), .ZN(n527) );
  OR2_X1 U742 ( .A1(n524), .A2(n523), .ZN(n532) );
  OR2_X1 U743 ( .A1(n778), .A2(n779), .ZN(n523) );
  AND2_X1 U744 ( .A1(n510), .A2(n509), .ZN(n779) );
  AND2_X1 U745 ( .A1(n507), .A2(n780), .ZN(n778) );
  OR2_X1 U746 ( .A1(n509), .A2(n510), .ZN(n780) );
  OR2_X1 U747 ( .A1(n661), .A2(n643), .ZN(n510) );
  OR2_X1 U748 ( .A1(n781), .A2(n782), .ZN(n509) );
  AND2_X1 U749 ( .A1(n496), .A2(n495), .ZN(n782) );
  AND2_X1 U750 ( .A1(n493), .A2(n783), .ZN(n781) );
  OR2_X1 U751 ( .A1(n495), .A2(n496), .ZN(n783) );
  OR2_X1 U752 ( .A1(n713), .A2(n643), .ZN(n496) );
  OR2_X1 U753 ( .A1(n784), .A2(n785), .ZN(n495) );
  AND2_X1 U754 ( .A1(n630), .A2(n629), .ZN(n785) );
  AND2_X1 U755 ( .A1(n627), .A2(n786), .ZN(n784) );
  OR2_X1 U756 ( .A1(n630), .A2(n629), .ZN(n786) );
  OR2_X1 U757 ( .A1(n787), .A2(n788), .ZN(n629) );
  AND2_X1 U758 ( .A1(n611), .A2(n610), .ZN(n788) );
  AND2_X1 U759 ( .A1(n608), .A2(n789), .ZN(n787) );
  OR2_X1 U760 ( .A1(n611), .A2(n610), .ZN(n789) );
  OR2_X1 U761 ( .A1(n790), .A2(n791), .ZN(n610) );
  AND2_X1 U762 ( .A1(n599), .A2(n598), .ZN(n791) );
  AND2_X1 U763 ( .A1(n596), .A2(n792), .ZN(n790) );
  OR2_X1 U764 ( .A1(n599), .A2(n598), .ZN(n792) );
  OR2_X1 U765 ( .A1(n793), .A2(n794), .ZN(n598) );
  AND2_X1 U766 ( .A1(n580), .A2(n581), .ZN(n794) );
  AND2_X1 U767 ( .A1(n578), .A2(n795), .ZN(n793) );
  OR2_X1 U768 ( .A1(n580), .A2(n581), .ZN(n795) );
  OR2_X1 U769 ( .A1(n643), .A2(n796), .ZN(n581) );
  OR2_X1 U770 ( .A1(n797), .A2(n570), .ZN(n796) );
  OR2_X1 U771 ( .A1(n640), .A2(n643), .ZN(n580) );
  XNOR2_X1 U772 ( .A(n798), .B(n799), .ZN(n578) );
  OR2_X1 U773 ( .A1(n797), .A2(n574), .ZN(n798) );
  OR2_X1 U774 ( .A1(n764), .A2(n643), .ZN(n599) );
  XNOR2_X1 U775 ( .A(n800), .B(n801), .ZN(n596) );
  XNOR2_X1 U776 ( .A(n802), .B(n803), .ZN(n800) );
  OR2_X1 U777 ( .A1(n623), .A2(n643), .ZN(n611) );
  XOR2_X1 U778 ( .A(n804), .B(n805), .Z(n608) );
  XOR2_X1 U779 ( .A(n806), .B(n807), .Z(n805) );
  OR2_X1 U780 ( .A1(n702), .A2(n643), .ZN(n630) );
  XOR2_X1 U781 ( .A(n808), .B(n809), .Z(n627) );
  XOR2_X1 U782 ( .A(n810), .B(n811), .Z(n809) );
  XOR2_X1 U783 ( .A(n812), .B(n813), .Z(n493) );
  XOR2_X1 U784 ( .A(n814), .B(n815), .Z(n813) );
  XOR2_X1 U785 ( .A(n816), .B(n817), .Z(n507) );
  XOR2_X1 U786 ( .A(n818), .B(n819), .Z(n817) );
  XOR2_X1 U787 ( .A(n820), .B(n821), .Z(n524) );
  XOR2_X1 U788 ( .A(n822), .B(n823), .Z(n821) );
  OR2_X1 U789 ( .A1(n536), .A2(n824), .ZN(n777) );
  AND2_X1 U790 ( .A1(n530), .A2(n531), .ZN(n824) );
  INV_X1 U791 ( .A(n825), .ZN(n536) );
  OR2_X1 U792 ( .A1(n530), .A2(n531), .ZN(n825) );
  OR2_X1 U793 ( .A1(n826), .A2(n827), .ZN(n531) );
  AND2_X1 U794 ( .A1(n823), .A2(n822), .ZN(n827) );
  AND2_X1 U795 ( .A1(n820), .A2(n828), .ZN(n826) );
  OR2_X1 U796 ( .A1(n822), .A2(n823), .ZN(n828) );
  OR2_X1 U797 ( .A1(n574), .A2(n661), .ZN(n823) );
  OR2_X1 U798 ( .A1(n829), .A2(n830), .ZN(n822) );
  AND2_X1 U799 ( .A1(n819), .A2(n818), .ZN(n830) );
  AND2_X1 U800 ( .A1(n816), .A2(n831), .ZN(n829) );
  OR2_X1 U801 ( .A1(n818), .A2(n819), .ZN(n831) );
  OR2_X1 U802 ( .A1(n574), .A2(n713), .ZN(n819) );
  OR2_X1 U803 ( .A1(n832), .A2(n833), .ZN(n818) );
  AND2_X1 U804 ( .A1(n815), .A2(n814), .ZN(n833) );
  AND2_X1 U805 ( .A1(n812), .A2(n834), .ZN(n832) );
  OR2_X1 U806 ( .A1(n814), .A2(n815), .ZN(n834) );
  OR2_X1 U807 ( .A1(n574), .A2(n702), .ZN(n815) );
  OR2_X1 U808 ( .A1(n835), .A2(n836), .ZN(n814) );
  AND2_X1 U809 ( .A1(n811), .A2(n810), .ZN(n836) );
  AND2_X1 U810 ( .A1(n808), .A2(n837), .ZN(n835) );
  OR2_X1 U811 ( .A1(n811), .A2(n810), .ZN(n837) );
  OR2_X1 U812 ( .A1(n838), .A2(n839), .ZN(n810) );
  AND2_X1 U813 ( .A1(n807), .A2(n806), .ZN(n839) );
  AND2_X1 U814 ( .A1(n804), .A2(n840), .ZN(n838) );
  OR2_X1 U815 ( .A1(n807), .A2(n806), .ZN(n840) );
  OR2_X1 U816 ( .A1(n841), .A2(n842), .ZN(n806) );
  AND2_X1 U817 ( .A1(n802), .A2(n803), .ZN(n842) );
  AND2_X1 U818 ( .A1(n801), .A2(n843), .ZN(n841) );
  OR2_X1 U819 ( .A1(n802), .A2(n803), .ZN(n843) );
  OR2_X1 U820 ( .A1(n570), .A2(n844), .ZN(n803) );
  OR2_X1 U821 ( .A1(n565), .A2(n574), .ZN(n570) );
  OR2_X1 U822 ( .A1(n574), .A2(n640), .ZN(n802) );
  XNOR2_X1 U823 ( .A(n845), .B(n844), .ZN(n801) );
  OR2_X1 U824 ( .A1(n797), .A2(n592), .ZN(n844) );
  OR2_X1 U825 ( .A1(n565), .A2(n748), .ZN(n845) );
  OR2_X1 U826 ( .A1(n574), .A2(n764), .ZN(n807) );
  XNOR2_X1 U827 ( .A(n846), .B(n847), .ZN(n804) );
  XNOR2_X1 U828 ( .A(n848), .B(n590), .ZN(n846) );
  OR2_X1 U829 ( .A1(n574), .A2(n623), .ZN(n811) );
  INV_X1 U830 ( .A(b_6_), .ZN(n574) );
  XOR2_X1 U831 ( .A(n849), .B(n850), .Z(n808) );
  XOR2_X1 U832 ( .A(n851), .B(n852), .Z(n850) );
  XOR2_X1 U833 ( .A(n853), .B(n854), .Z(n812) );
  XOR2_X1 U834 ( .A(n855), .B(n856), .Z(n854) );
  XOR2_X1 U835 ( .A(n857), .B(n858), .Z(n816) );
  XOR2_X1 U836 ( .A(n859), .B(n860), .Z(n858) );
  XOR2_X1 U837 ( .A(n861), .B(n862), .Z(n820) );
  XOR2_X1 U838 ( .A(n863), .B(n864), .Z(n862) );
  XOR2_X1 U839 ( .A(n743), .B(n865), .Z(n530) );
  XOR2_X1 U840 ( .A(n746), .B(n744), .Z(n865) );
  OR2_X1 U841 ( .A1(n592), .A2(n661), .ZN(n744) );
  OR2_X1 U842 ( .A1(n866), .A2(n867), .ZN(n746) );
  AND2_X1 U843 ( .A1(n864), .A2(n863), .ZN(n867) );
  AND2_X1 U844 ( .A1(n861), .A2(n868), .ZN(n866) );
  OR2_X1 U845 ( .A1(n863), .A2(n864), .ZN(n868) );
  OR2_X1 U846 ( .A1(n592), .A2(n713), .ZN(n864) );
  OR2_X1 U847 ( .A1(n869), .A2(n870), .ZN(n863) );
  AND2_X1 U848 ( .A1(n860), .A2(n859), .ZN(n870) );
  AND2_X1 U849 ( .A1(n857), .A2(n871), .ZN(n869) );
  OR2_X1 U850 ( .A1(n859), .A2(n860), .ZN(n871) );
  OR2_X1 U851 ( .A1(n592), .A2(n702), .ZN(n860) );
  OR2_X1 U852 ( .A1(n872), .A2(n873), .ZN(n859) );
  AND2_X1 U853 ( .A1(n856), .A2(n855), .ZN(n873) );
  AND2_X1 U854 ( .A1(n853), .A2(n874), .ZN(n872) );
  OR2_X1 U855 ( .A1(n855), .A2(n856), .ZN(n874) );
  OR2_X1 U856 ( .A1(n592), .A2(n623), .ZN(n856) );
  OR2_X1 U857 ( .A1(n875), .A2(n876), .ZN(n855) );
  AND2_X1 U858 ( .A1(n852), .A2(n851), .ZN(n876) );
  AND2_X1 U859 ( .A1(n849), .A2(n877), .ZN(n875) );
  OR2_X1 U860 ( .A1(n852), .A2(n851), .ZN(n877) );
  OR2_X1 U861 ( .A1(n878), .A2(n879), .ZN(n851) );
  AND2_X1 U862 ( .A1(n847), .A2(n590), .ZN(n879) );
  AND2_X1 U863 ( .A1(n880), .A2(n848), .ZN(n878) );
  OR2_X1 U864 ( .A1(n881), .A2(n882), .ZN(n848) );
  INV_X1 U865 ( .A(n883), .ZN(n882) );
  AND2_X1 U866 ( .A1(n884), .A2(n885), .ZN(n881) );
  OR2_X1 U867 ( .A1(n847), .A2(n590), .ZN(n880) );
  INV_X1 U868 ( .A(n886), .ZN(n590) );
  AND2_X1 U869 ( .A1(b_5_), .A2(a_5_), .ZN(n886) );
  OR2_X1 U870 ( .A1(n885), .A2(n799), .ZN(n847) );
  OR2_X1 U871 ( .A1(n565), .A2(n592), .ZN(n799) );
  OR2_X1 U872 ( .A1(n592), .A2(n764), .ZN(n852) );
  INV_X1 U873 ( .A(b_5_), .ZN(n592) );
  XNOR2_X1 U874 ( .A(n887), .B(n888), .ZN(n849) );
  XNOR2_X1 U875 ( .A(n889), .B(n883), .ZN(n887) );
  XNOR2_X1 U876 ( .A(n890), .B(n891), .ZN(n853) );
  XNOR2_X1 U877 ( .A(n603), .B(n892), .ZN(n890) );
  XOR2_X1 U878 ( .A(n893), .B(n894), .Z(n857) );
  XOR2_X1 U879 ( .A(n895), .B(n896), .Z(n894) );
  XOR2_X1 U880 ( .A(n897), .B(n898), .Z(n861) );
  XOR2_X1 U881 ( .A(n899), .B(n900), .Z(n898) );
  XOR2_X1 U882 ( .A(n751), .B(n901), .Z(n743) );
  XOR2_X1 U883 ( .A(n754), .B(n752), .Z(n901) );
  OR2_X1 U884 ( .A1(n748), .A2(n713), .ZN(n752) );
  OR2_X1 U885 ( .A1(n902), .A2(n903), .ZN(n754) );
  AND2_X1 U886 ( .A1(n900), .A2(n899), .ZN(n903) );
  AND2_X1 U887 ( .A1(n897), .A2(n904), .ZN(n902) );
  OR2_X1 U888 ( .A1(n899), .A2(n900), .ZN(n904) );
  OR2_X1 U889 ( .A1(n748), .A2(n702), .ZN(n900) );
  OR2_X1 U890 ( .A1(n905), .A2(n906), .ZN(n899) );
  AND2_X1 U891 ( .A1(n896), .A2(n895), .ZN(n906) );
  AND2_X1 U892 ( .A1(n893), .A2(n907), .ZN(n905) );
  OR2_X1 U893 ( .A1(n895), .A2(n896), .ZN(n907) );
  OR2_X1 U894 ( .A1(n748), .A2(n623), .ZN(n896) );
  OR2_X1 U895 ( .A1(n908), .A2(n909), .ZN(n895) );
  AND2_X1 U896 ( .A1(n892), .A2(n603), .ZN(n909) );
  AND2_X1 U897 ( .A1(n891), .A2(n910), .ZN(n908) );
  OR2_X1 U898 ( .A1(n603), .A2(n892), .ZN(n910) );
  OR2_X1 U899 ( .A1(n911), .A2(n912), .ZN(n892) );
  AND2_X1 U900 ( .A1(n888), .A2(n883), .ZN(n912) );
  AND2_X1 U901 ( .A1(n913), .A2(n889), .ZN(n911) );
  OR2_X1 U902 ( .A1(n914), .A2(n915), .ZN(n889) );
  AND2_X1 U903 ( .A1(n916), .A2(n917), .ZN(n914) );
  OR2_X1 U904 ( .A1(n888), .A2(n883), .ZN(n913) );
  OR2_X1 U905 ( .A1(n884), .A2(n885), .ZN(n883) );
  OR2_X1 U906 ( .A1(n797), .A2(n748), .ZN(n885) );
  OR2_X1 U907 ( .A1(n565), .A2(n622), .ZN(n884) );
  OR2_X1 U908 ( .A1(n640), .A2(n748), .ZN(n888) );
  OR2_X1 U909 ( .A1(n764), .A2(n748), .ZN(n603) );
  INV_X1 U910 ( .A(b_4_), .ZN(n748) );
  XOR2_X1 U911 ( .A(n918), .B(n915), .Z(n891) );
  INV_X1 U912 ( .A(n919), .ZN(n915) );
  XNOR2_X1 U913 ( .A(n920), .B(n921), .ZN(n918) );
  XNOR2_X1 U914 ( .A(n922), .B(n923), .ZN(n893) );
  XNOR2_X1 U915 ( .A(n924), .B(n925), .ZN(n922) );
  XNOR2_X1 U916 ( .A(n926), .B(n927), .ZN(n897) );
  XNOR2_X1 U917 ( .A(n635), .B(n928), .ZN(n926) );
  XNOR2_X1 U918 ( .A(n929), .B(n775), .ZN(n751) );
  XNOR2_X1 U919 ( .A(n930), .B(n769), .ZN(n775) );
  XOR2_X1 U920 ( .A(n931), .B(n760), .Z(n769) );
  OR2_X1 U921 ( .A1(n640), .A2(n703), .ZN(n760) );
  XOR2_X1 U922 ( .A(n762), .B(n761), .Z(n931) );
  OR2_X1 U923 ( .A1(n660), .A2(n764), .ZN(n761) );
  AND2_X1 U924 ( .A1(n932), .A2(n933), .ZN(n762) );
  XNOR2_X1 U925 ( .A(n768), .B(n767), .ZN(n930) );
  OR2_X1 U926 ( .A1(n934), .A2(n935), .ZN(n767) );
  AND2_X1 U927 ( .A1(n936), .A2(n937), .ZN(n935) );
  AND2_X1 U928 ( .A1(n938), .A2(n939), .ZN(n934) );
  OR2_X1 U929 ( .A1(n937), .A2(n936), .ZN(n939) );
  OR2_X1 U930 ( .A1(n712), .A2(n623), .ZN(n768) );
  XNOR2_X1 U931 ( .A(n774), .B(n773), .ZN(n929) );
  OR2_X1 U932 ( .A1(n940), .A2(n941), .ZN(n773) );
  AND2_X1 U933 ( .A1(n928), .A2(n635), .ZN(n941) );
  AND2_X1 U934 ( .A1(n927), .A2(n942), .ZN(n940) );
  OR2_X1 U935 ( .A1(n635), .A2(n928), .ZN(n942) );
  OR2_X1 U936 ( .A1(n943), .A2(n944), .ZN(n928) );
  AND2_X1 U937 ( .A1(n925), .A2(n924), .ZN(n944) );
  AND2_X1 U938 ( .A1(n923), .A2(n945), .ZN(n943) );
  OR2_X1 U939 ( .A1(n924), .A2(n925), .ZN(n945) );
  OR2_X1 U940 ( .A1(n946), .A2(n947), .ZN(n925) );
  AND2_X1 U941 ( .A1(n919), .A2(n921), .ZN(n947) );
  AND2_X1 U942 ( .A1(n948), .A2(n920), .ZN(n946) );
  OR2_X1 U943 ( .A1(n949), .A2(n950), .ZN(n920) );
  INV_X1 U944 ( .A(n951), .ZN(n950) );
  AND2_X1 U945 ( .A1(n952), .A2(n953), .ZN(n949) );
  OR2_X1 U946 ( .A1(n921), .A2(n919), .ZN(n948) );
  OR2_X1 U947 ( .A1(n916), .A2(n917), .ZN(n919) );
  OR2_X1 U948 ( .A1(n712), .A2(n565), .ZN(n917) );
  OR2_X1 U949 ( .A1(n797), .A2(n622), .ZN(n916) );
  OR2_X1 U950 ( .A1(n640), .A2(n622), .ZN(n921) );
  OR2_X1 U951 ( .A1(n764), .A2(n622), .ZN(n924) );
  XNOR2_X1 U952 ( .A(n954), .B(n955), .ZN(n923) );
  XNOR2_X1 U953 ( .A(n956), .B(n951), .ZN(n954) );
  INV_X1 U954 ( .A(n618), .ZN(n635) );
  AND2_X1 U955 ( .A1(b_3_), .A2(a_3_), .ZN(n618) );
  XOR2_X1 U956 ( .A(n938), .B(n957), .Z(n927) );
  XOR2_X1 U957 ( .A(n937), .B(n936), .Z(n957) );
  OR2_X1 U958 ( .A1(n712), .A2(n764), .ZN(n936) );
  OR2_X1 U959 ( .A1(n958), .A2(n959), .ZN(n937) );
  AND2_X1 U960 ( .A1(n955), .A2(n951), .ZN(n959) );
  AND2_X1 U961 ( .A1(n960), .A2(n956), .ZN(n958) );
  OR2_X1 U962 ( .A1(n961), .A2(n962), .ZN(n956) );
  INV_X1 U963 ( .A(n933), .ZN(n962) );
  AND2_X1 U964 ( .A1(n963), .A2(n964), .ZN(n961) );
  OR2_X1 U965 ( .A1(n951), .A2(n955), .ZN(n960) );
  OR2_X1 U966 ( .A1(n712), .A2(n640), .ZN(n955) );
  OR2_X1 U967 ( .A1(n952), .A2(n953), .ZN(n951) );
  OR2_X1 U968 ( .A1(n712), .A2(n797), .ZN(n953) );
  INV_X1 U969 ( .A(b_2_), .ZN(n712) );
  OR2_X1 U970 ( .A1(n660), .A2(n565), .ZN(n952) );
  XNOR2_X1 U971 ( .A(n965), .B(n933), .ZN(n938) );
  OR2_X1 U972 ( .A1(n964), .A2(n963), .ZN(n933) );
  OR2_X1 U973 ( .A1(n565), .A2(n703), .ZN(n963) );
  INV_X1 U974 ( .A(a_7_), .ZN(n565) );
  OR2_X1 U975 ( .A1(n660), .A2(n797), .ZN(n964) );
  OR2_X1 U976 ( .A1(n966), .A2(n967), .ZN(n965) );
  INV_X1 U977 ( .A(n932), .ZN(n967) );
  OR2_X1 U978 ( .A1(n968), .A2(n969), .ZN(n932) );
  AND2_X1 U979 ( .A1(n969), .A2(n968), .ZN(n966) );
  OR2_X1 U980 ( .A1(n660), .A2(n640), .ZN(n968) );
  INV_X1 U981 ( .A(b_1_), .ZN(n660) );
  OR2_X1 U982 ( .A1(n797), .A2(n703), .ZN(n969) );
  INV_X1 U983 ( .A(b_0_), .ZN(n703) );
  OR2_X1 U984 ( .A1(n622), .A2(n702), .ZN(n774) );
  INV_X1 U985 ( .A(b_3_), .ZN(n622) );
  INV_X1 U986 ( .A(n498), .ZN(n492) );
  OR2_X1 U987 ( .A1(n970), .A2(n513), .ZN(n498) );
  AND2_X1 U988 ( .A1(b_0_), .A2(n661), .ZN(n513) );
  AND2_X1 U989 ( .A1(n971), .A2(n972), .ZN(n970) );
  OR2_X1 U990 ( .A1(b_0_), .A2(n661), .ZN(n972) );
  INV_X1 U991 ( .A(a_0_), .ZN(n661) );
  AND2_X1 U992 ( .A1(n502), .A2(n973), .ZN(n971) );
  OR2_X1 U993 ( .A1(n974), .A2(n975), .ZN(n973) );
  OR2_X1 U994 ( .A1(n503), .A2(n976), .ZN(n975) );
  AND2_X1 U995 ( .A1(b_2_), .A2(n702), .ZN(n976) );
  AND2_X1 U996 ( .A1(n713), .A2(b_1_), .ZN(n503) );
  AND2_X1 U997 ( .A1(n977), .A2(n978), .ZN(n974) );
  OR2_X1 U998 ( .A1(b_3_), .A2(n623), .ZN(n978) );
  AND2_X1 U999 ( .A1(n979), .A2(n980), .ZN(n977) );
  OR2_X1 U1000 ( .A1(n981), .A2(n982), .ZN(n980) );
  OR2_X1 U1001 ( .A1(n983), .A2(n619), .ZN(n982) );
  AND2_X1 U1002 ( .A1(n623), .A2(b_3_), .ZN(n619) );
  INV_X1 U1003 ( .A(a_3_), .ZN(n623) );
  AND2_X1 U1004 ( .A1(n984), .A2(n985), .ZN(n983) );
  OR2_X1 U1005 ( .A1(b_5_), .A2(n640), .ZN(n985) );
  AND2_X1 U1006 ( .A1(n986), .A2(n987), .ZN(n984) );
  OR2_X1 U1007 ( .A1(n988), .A2(n989), .ZN(n987) );
  OR2_X1 U1008 ( .A1(n990), .A2(n587), .ZN(n989) );
  AND2_X1 U1009 ( .A1(n640), .A2(b_5_), .ZN(n587) );
  INV_X1 U1010 ( .A(a_5_), .ZN(n640) );
  AND2_X1 U1011 ( .A1(b_6_), .A2(n991), .ZN(n990) );
  OR2_X1 U1012 ( .A1(n992), .A2(n797), .ZN(n991) );
  AND2_X1 U1013 ( .A1(n797), .A2(n992), .ZN(n988) );
  INV_X1 U1014 ( .A(n564), .ZN(n992) );
  AND2_X1 U1015 ( .A1(n643), .A2(a_7_), .ZN(n564) );
  INV_X1 U1016 ( .A(b_7_), .ZN(n643) );
  INV_X1 U1017 ( .A(a_6_), .ZN(n797) );
  OR2_X1 U1018 ( .A1(b_4_), .A2(n764), .ZN(n986) );
  AND2_X1 U1019 ( .A1(b_4_), .A2(n764), .ZN(n981) );
  INV_X1 U1020 ( .A(a_4_), .ZN(n764) );
  OR2_X1 U1021 ( .A1(b_2_), .A2(n702), .ZN(n979) );
  INV_X1 U1022 ( .A(a_2_), .ZN(n702) );
  OR2_X1 U1023 ( .A1(b_1_), .A2(n713), .ZN(n502) );
  INV_X1 U1024 ( .A(a_1_), .ZN(n713) );
endmodule

