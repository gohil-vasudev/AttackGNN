module top ( keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880 );
input keyIn_0_0, keyIn_0_1, keyIn_0_2, keyIn_0_3, keyIn_0_4, keyIn_0_5, keyIn_0_6, keyIn_0_7, keyIn_0_8, keyIn_0_9, keyIn_0_10, keyIn_0_11, keyIn_0_12, keyIn_0_13, keyIn_0_14, keyIn_0_15, keyIn_0_16, keyIn_0_17, keyIn_0_18, keyIn_0_19, keyIn_0_20, keyIn_0_21, keyIn_0_22, keyIn_0_23, keyIn_0_24, keyIn_0_25, keyIn_0_26, keyIn_0_27, keyIn_0_28, keyIn_0_29, keyIn_0_30, keyIn_0_31, keyIn_0_32, keyIn_0_33, keyIn_0_34, keyIn_0_35, keyIn_0_36, keyIn_0_37, keyIn_0_38, keyIn_0_39, keyIn_0_40, keyIn_0_41, keyIn_0_42, keyIn_0_43, keyIn_0_44, keyIn_0_45, keyIn_0_46, keyIn_0_47, keyIn_0_48, keyIn_0_49, keyIn_0_50, keyIn_0_51, keyIn_0_52, keyIn_0_53, keyIn_0_54, keyIn_0_55, keyIn_0_56, keyIn_0_57, keyIn_0_58, keyIn_0_59, keyIn_0_60, keyIn_0_61, keyIn_0_62, keyIn_0_63, keyIn_0_64, keyIn_0_65, keyIn_0_66, keyIn_0_67, keyIn_0_68, keyIn_0_69, keyIn_0_70, keyIn_0_71, keyIn_0_72, keyIn_0_73, keyIn_0_74, keyIn_0_75, keyIn_0_76, keyIn_0_77, keyIn_0_78, keyIn_0_79, keyIn_0_80, keyIn_0_81, keyIn_0_82, keyIn_0_83, keyIn_0_84, keyIn_0_85, keyIn_0_86, keyIn_0_87, keyIn_0_88, keyIn_0_89, keyIn_0_90, keyIn_0_91, keyIn_0_92, keyIn_0_93, keyIn_0_94, keyIn_0_95, keyIn_0_96, keyIn_0_97, keyIn_0_98, keyIn_0_99, keyIn_0_100, keyIn_0_101, keyIn_0_102, keyIn_0_103, keyIn_0_104, keyIn_0_105, keyIn_0_106, keyIn_0_107, keyIn_0_108, keyIn_0_109, keyIn_0_110, keyIn_0_111, keyIn_0_112, keyIn_0_113, keyIn_0_114, keyIn_0_115, keyIn_0_116, keyIn_0_117, keyIn_0_118, keyIn_0_119, keyIn_0_120, keyIn_0_121, keyIn_0_122, keyIn_0_123, keyIn_0_124, keyIn_0_125, keyIn_0_126, keyIn_0_127, keyIn_0_128, keyIn_0_129, keyIn_0_130, keyIn_0_131, keyIn_0_132, keyIn_0_133, keyIn_0_134, keyIn_0_135, keyIn_0_136, keyIn_0_137, keyIn_0_138, keyIn_0_139, keyIn_0_140, keyIn_0_141, keyIn_0_142, keyIn_0_143, keyIn_0_144, keyIn_0_145, keyIn_0_146, keyIn_0_147, keyIn_0_148, keyIn_0_149, keyIn_0_150, keyIn_0_151, keyIn_0_152, keyIn_0_153, keyIn_0_154, keyIn_0_155, keyIn_0_156, keyIn_0_157, keyIn_0_158, keyIn_0_159, keyIn_0_160, keyIn_0_161, keyIn_0_162, keyIn_0_163, keyIn_0_164, keyIn_0_165, keyIn_0_166, keyIn_0_167, keyIn_0_168, keyIn_0_169, keyIn_0_170, keyIn_0_171, keyIn_0_172, keyIn_0_173, keyIn_0_174, keyIn_0_175, keyIn_0_176, keyIn_0_177, keyIn_0_178, keyIn_0_179, keyIn_0_180, keyIn_0_181, keyIn_0_182, keyIn_0_183, keyIn_0_184, keyIn_0_185, keyIn_0_186, keyIn_0_187, keyIn_0_188, keyIn_0_189, keyIn_0_190, keyIn_0_191, keyIn_0_192, keyIn_0_193, keyIn_0_194, keyIn_0_195, keyIn_0_196, keyIn_0_197, keyIn_0_198, keyIn_0_199, keyIn_0_200, keyIn_0_201, keyIn_0_202, keyIn_0_203, keyIn_0_204, keyIn_0_205, keyIn_0_206, keyIn_0_207, keyIn_0_208, keyIn_0_209, keyIn_0_210, keyIn_0_211, keyIn_0_212, keyIn_0_213, keyIn_0_214, keyIn_0_215, keyIn_0_216, keyIn_0_217, keyIn_0_218, keyIn_0_219, keyIn_0_220, keyIn_0_221, keyIn_0_222, keyIn_0_223, keyIn_0_224, keyIn_0_225, keyIn_0_226, keyIn_0_227, keyIn_0_228, keyIn_0_229, keyIn_0_230, keyIn_0_231, keyIn_0_232, keyIn_0_233, keyIn_0_234, keyIn_0_235, keyIn_0_236, keyIn_0_237, keyIn_0_238, keyIn_0_239, keyIn_0_240, keyIn_0_241, keyIn_0_242, keyIn_0_243, keyIn_0_244, keyIn_0_245, keyIn_0_246, keyIn_0_247, keyIn_0_248, keyIn_0_249, keyIn_0_250, keyIn_0_251, keyIn_0_252, keyIn_0_253, keyIn_0_254, keyIn_0_255, N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;
output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;
wire new_n942_, new_n595_, new_n614_, new_n895_, new_n958_, new_n445_, new_n699_, new_n976_, new_n1009_, new_n1233_, new_n479_, new_n1105_, new_n1215_, new_n1249_, new_n955_, new_n608_, new_n888_, new_n847_, new_n501_, new_n1157_, new_n798_, new_n1180_, new_n421_, new_n817_, new_n777_, new_n720_, new_n753_, new_n620_, new_n368_, new_n1048_, new_n738_, new_n941_, new_n885_, new_n439_, new_n827_, new_n390_, new_n743_, new_n366_, new_n779_, new_n1232_, new_n1025_, new_n566_, new_n641_, new_n859_, new_n386_, new_n767_, new_n401_, new_n389_, new_n1176_, new_n1207_, new_n1211_, new_n514_, new_n601_, new_n842_, new_n556_, new_n636_, new_n1057_, new_n670_, new_n1024_, new_n456_, new_n691_, new_n1125_, new_n682_, new_n1075_, new_n812_, new_n911_, new_n679_, new_n937_, new_n667_, new_n367_, new_n821_, new_n542_, new_n548_, new_n669_, new_n1237_, new_n1172_, new_n419_, new_n728_, new_n624_, new_n534_, new_n1071_, new_n1131_, new_n1120_, new_n819_, new_n637_, new_n451_, new_n489_, new_n424_, new_n804_, new_n894_, new_n853_, new_n602_, new_n1210_, new_n695_, new_n660_, new_n1060_, new_n413_, new_n526_, new_n442_, new_n677_, new_n908_, new_n642_, new_n552_, new_n678_, new_n649_, new_n706_, new_n1119_, new_n462_, new_n603_, new_n564_, new_n752_, new_n761_, new_n1213_, new_n840_, new_n735_, new_n1283_, new_n1045_, new_n500_, new_n898_, new_n1163_, new_n786_, new_n799_, new_n946_, new_n1188_, new_n344_, new_n721_, new_n504_, new_n1108_, new_n862_, new_n742_, new_n892_, new_n427_, new_n532_, new_n472_, new_n393_, new_n873_, new_n418_, new_n746_, new_n1221_, new_n1167_, new_n1264_, new_n626_, new_n959_, new_n774_, new_n716_, new_n701_, new_n1238_, new_n792_, new_n1058_, new_n953_, new_n1162_, new_n481_, new_n1265_, new_n1073_, new_n1110_, new_n1278_, new_n902_, new_n364_, new_n449_, new_n580_, new_n484_, new_n639_, new_n832_, new_n766_, new_n1262_, new_n1212_, new_n1059_, new_n634_, new_n414_, new_n1101_, new_n1250_, new_n635_, new_n685_, new_n1050_, new_n554_, new_n648_, new_n903_, new_n983_, new_n1151_, new_n844_, new_n430_, new_n822_, new_n482_, new_n1082_, new_n849_, new_n1203_, new_n1018_, new_n855_, new_n606_, new_n1037_, new_n589_, new_n796_, new_n1083_, new_n655_, new_n759_, new_n1054_, new_n630_, new_n385_, new_n1049_, new_n829_, new_n1257_, new_n988_, new_n478_, new_n694_, new_n461_, new_n1228_, new_n710_, new_n971_, new_n565_, new_n361_, new_n764_, new_n906_, new_n683_, new_n1196_, new_n511_, new_n463_, new_n510_, new_n966_, new_n1184_, new_n517_, new_n609_, new_n1285_, new_n1031_, new_n961_, new_n890_, new_n530_, new_n1216_, new_n1006_, new_n622_, new_n1281_, new_n629_, new_n702_, new_n833_, new_n1214_, new_n1005_, new_n883_, new_n999_, new_n715_, new_n811_, new_n443_, new_n1086_, new_n956_, new_n763_, new_n960_, new_n1138_, new_n486_, new_n491_, new_n549_, new_n676_, new_n466_, new_n970_, new_n995_, new_n1035_, new_n674_, new_n991_, new_n1044_, new_n497_, new_n1170_, new_n816_, new_n845_, new_n768_, new_n773_, new_n568_, new_n420_, new_n1051_, new_n876_, new_n899_, new_n1053_, new_n423_, new_n498_, new_n492_, new_n496_, new_n1046_, new_n1182_, new_n1200_, new_n650_, new_n708_, new_n750_, new_n1217_, new_n887_, new_n429_, new_n355_, new_n926_, new_n353_, new_n1222_, new_n432_, new_n734_, new_n912_, new_n1062_, new_n925_, new_n875_, new_n506_, new_n680_, new_n872_, new_n981_, new_n1226_, new_n1275_, new_n778_, new_n1277_, new_n452_, new_n1198_, new_n381_, new_n1219_, new_n920_, new_n656_, new_n1121_, new_n820_, new_n1127_, new_n771_, new_n388_, new_n979_, new_n1028_, new_n1168_, new_n508_, new_n714_, new_n483_, new_n1004_, new_n1152_, new_n1280_, new_n1007_, new_n935_, new_n1241_, new_n882_, new_n1145_, new_n657_, new_n1150_, new_n929_, new_n652_, new_n582_, new_n986_, new_n1159_, new_n1020_, new_n363_, new_n1266_, new_n1113_, new_n441_, new_n785_, new_n477_, new_n664_, new_n600_, new_n1041_, new_n917_, new_n426_, new_n1036_, new_n1133_, new_n1177_, new_n646_, new_n1132_, new_n395_, new_n538_, new_n383_, new_n343_, new_n541_, new_n458_, new_n854_, new_n447_, new_n1026_, new_n1106_, new_n473_, new_n1147_, new_n1229_, new_n790_, new_n1081_, new_n587_, new_n1247_, new_n465_, new_n739_, new_n783_, new_n969_, new_n835_, new_n1234_, new_n996_, new_n378_, new_n621_, new_n846_, new_n915_, new_n349_, new_n488_, new_n524_, new_n705_, new_n848_, new_n874_, new_n663_, new_n579_, new_n1209_, new_n347_, new_n659_, new_n1254_, new_n700_, new_n921_, new_n396_, new_n438_, new_n1003_, new_n696_, new_n939_, new_n632_, new_n1039_, new_n671_, new_n965_, new_n1239_, new_n528_, new_n952_, new_n1158_, new_n572_, new_n850_, new_n1019_, new_n436_, new_n1202_, new_n397_, new_n729_, new_n1111_, new_n975_, new_n1199_, new_n399_, new_n596_, new_n1218_, new_n870_, new_n945_, new_n805_, new_n1115_, new_n559_, new_n1201_, new_n1282_, new_n948_, new_n1231_, new_n762_, new_n1055_, new_n1193_, new_n838_, new_n923_, new_n1187_, new_n469_, new_n1154_, new_n437_, new_n1085_, new_n1253_, new_n1256_, new_n794_, new_n628_, new_n1090_, new_n457_, new_n553_, new_n1114_, new_n1084_, new_n1061_, new_n668_, new_n1128_, new_n1002_, new_n834_, new_n1169_, new_n369_, new_n448_, new_n867_, new_n954_, new_n901_, new_n1032_, new_n1171_, new_n688_, new_n1255_, new_n384_, new_n900_, new_n1161_, new_n410_, new_n985_, new_n851_, new_n932_, new_n878_, new_n543_, new_n924_, new_n775_, new_n886_, new_n509_, new_n454_, new_n1034_, new_n661_, new_n1124_, new_n1000_, new_n633_, new_n797_, new_n784_, new_n1273_, new_n724_, new_n1070_, new_n1109_, new_n860_, new_n494_, new_n672_, new_n1269_, new_n616_, new_n529_, new_n884_, new_n914_, new_n938_, new_n1160_, new_n362_, new_n1166_, new_n809_, new_n1142_, new_n654_, new_n713_, new_n880_, new_n1102_, new_n604_, new_n1104_, new_n690_, new_n416_, new_n1043_, new_n744_, new_n571_, new_n400_, new_n758_, new_n460_, new_n1175_, new_n1136_, new_n693_, new_n1267_, new_n1272_, new_n1287_, new_n505_, new_n619_, new_n471_, new_n967_, new_n577_, new_n374_, new_n1135_, new_n376_, new_n1271_, new_n380_, new_n1251_, new_n1079_, new_n747_, new_n749_, new_n861_, new_n1091_, new_n1095_, new_n1252_, new_n998_, new_n1056_, new_n352_, new_n1094_, new_n931_, new_n575_, new_n839_, new_n1030_, new_n485_, new_n525_, new_n578_, new_n944_, new_n918_, new_n940_, new_n810_, new_n808_, new_n1064_, new_n1065_, new_n1284_, new_n493_, new_n547_, new_n907_, new_n665_, new_n800_, new_n897_, new_n1012_, new_n719_, new_n869_, new_n1178_, new_n963_, new_n586_, new_n598_, new_n570_, new_n893_, new_n993_, new_n1063_, new_n1191_, new_n824_, new_n520_, new_n1001_, new_n717_, new_n403_, new_n475_, new_n868_, new_n1242_, new_n825_, new_n858_, new_n557_, new_n936_, new_n507_, new_n741_, new_n673_, new_n806_, new_n1016_, new_n605_, new_n1144_, new_n1074_, new_n748_, new_n1224_, new_n1137_, new_n1286_, new_n407_, new_n666_, new_n813_, new_n830_, new_n480_, new_n625_, new_n1107_, new_n730_, new_n1141_, new_n807_, new_n736_, new_n879_, new_n513_, new_n592_, new_n726_, new_n1263_, new_n1123_, new_n558_, new_n1080_, new_n583_, new_n617_, new_n718_, new_n1279_, new_n522_, new_n588_, new_n781_, new_n1014_, new_n428_, new_n916_, new_n487_, new_n360_, new_n675_, new_n1126_, new_n1155_, new_n546_, new_n1186_, new_n612_, new_n919_, new_n1015_, new_n755_, new_n1261_, new_n1040_, new_n1246_, new_n922_, new_n387_, new_n544_, new_n476_, new_n615_, new_n987_, new_n722_, new_n856_, new_n415_, new_n949_, new_n537_, new_n450_, new_n345_, new_n1179_, new_n499_, new_n533_, new_n1088_, new_n1130_, new_n1148_, new_n795_, new_n459_, new_n569_, new_n555_, new_n468_, new_n1122_, new_n977_, new_n1139_, new_n782_, new_n1185_, new_n1240_, new_n354_, new_n392_, new_n444_, new_n518_, new_n950_, new_n737_, new_n968_, new_n1022_, new_n1174_, new_n692_, new_n502_, new_n613_, new_n623_, new_n446_, new_n1195_, new_n590_, new_n417_, new_n658_, new_n591_, new_n826_, new_n801_, new_n837_, new_n789_, new_n515_, new_n972_, new_n1067_, new_n891_, new_n631_, new_n453_, new_n516_, new_n1227_, new_n997_, new_n519_, new_n563_, new_n662_, new_n864_, new_n910_, new_n440_, new_n733_, new_n531_, new_n1021_, new_n593_, new_n974_, new_n1076_, new_n585_, new_n1248_, new_n751_, new_n535_, new_n1038_, new_n372_, new_n725_, new_n814_, new_n503_, new_n527_, new_n772_, new_n852_, new_n1244_, new_n1181_, new_n597_, new_n978_, new_n1093_, new_n1092_, new_n408_, new_n1143_, new_n470_, new_n1072_, new_n769_, new_n1190_, new_n1097_, new_n1069_, new_n651_, new_n433_, new_n1164_, new_n871_, new_n435_, new_n1010_, new_n776_, new_n992_, new_n1098_, new_n732_, new_n687_, new_n370_, new_n1029_, new_n689_, new_n584_, new_n815_, new_n933_, new_n1052_, new_n638_, new_n523_, new_n909_, new_n857_, new_n712_, new_n1017_, new_n550_, new_n1068_, new_n512_, new_n788_, new_n841_, new_n1220_, new_n989_, new_n1204_, new_n1117_, new_n1112_, new_n711_, new_n1156_, new_n644_, new_n731_, new_n599_, new_n836_, new_n930_, new_n1116_, new_n1260_, new_n973_, new_n412_, new_n607_, new_n904_, new_n1276_, new_n645_, new_n913_, new_n1096_, new_n681_, new_n1087_, new_n723_, new_n594_, new_n561_, new_n495_, new_n756_, new_n431_, new_n823_, new_n927_, new_n1206_, new_n818_, new_n574_, new_n881_, new_n928_, new_n1268_, new_n1008_, new_n640_, new_n684_, new_n1274_, new_n707_, new_n740_, new_n957_, new_n754_, new_n1047_, new_n787_, new_n653_, new_n1134_, new_n377_, new_n539_, new_n905_, new_n1258_, new_n803_, new_n1270_, new_n727_, new_n962_, new_n760_, new_n627_, new_n1173_, new_n704_, new_n567_, new_n576_, new_n831_, new_n791_, new_n1033_, new_n1189_, new_n1153_, new_n357_, new_n1197_, new_n780_, new_n984_, new_n1183_, new_n643_, new_n474_, new_n1223_, new_n1129_, new_n467_, new_n1013_, new_n404_, new_n1194_, new_n1077_, new_n1243_, new_n560_, new_n1100_, new_n1230_, new_n865_, new_n1027_, new_n358_, new_n877_, new_n348_, new_n610_, new_n843_, new_n545_, new_n611_, new_n703_, new_n698_, new_n1011_, new_n1165_, new_n1259_, new_n425_, new_n896_, new_n802_, new_n1208_, new_n697_, new_n1099_, new_n1023_, new_n951_, new_n1236_, new_n709_, new_n373_, new_n866_, new_n1235_, new_n540_, new_n1149_, new_n1066_, new_n434_, new_n947_, new_n994_, new_n982_, new_n422_, new_n964_, new_n1078_, new_n581_, new_n686_, new_n934_, new_n551_, new_n455_, new_n770_, new_n757_, new_n618_, new_n1140_, new_n521_, new_n1225_, new_n1042_, new_n793_, new_n863_, new_n406_, new_n828_, new_n980_, new_n356_, new_n647_, new_n536_, new_n464_, new_n1089_, new_n1192_, new_n573_, new_n765_, new_n405_, new_n1103_;

not g000 ( new_n343_, N42 );
nand g001 ( new_n344_, N29, N75 );
nor g002 ( new_n345_, new_n344_, new_n343_ );
xor g003 ( N388, new_n345_, keyIn_0_5 );
not g004 ( new_n347_, N80 );
nand g005 ( new_n348_, N29, N36 );
nor g006 ( new_n349_, new_n348_, new_n347_ );
xor g007 ( N389, new_n349_, keyIn_0_6 );
nor g008 ( N390, new_n348_, new_n343_ );
not g009 ( new_n352_, keyIn_0_11 );
nand g010 ( new_n353_, N85, N86 );
nand g011 ( new_n354_, new_n353_, new_n352_ );
not g012 ( new_n355_, new_n354_ );
not g013 ( new_n356_, N86 );
nand g014 ( new_n357_, keyIn_0_11, N85 );
nor g015 ( new_n358_, new_n357_, new_n356_ );
nor g016 ( N391, new_n355_, new_n358_ );
not g017 ( new_n360_, N13 );
nand g018 ( new_n361_, N1, N8 );
nor g019 ( new_n362_, new_n361_, new_n360_ );
nand g020 ( new_n363_, new_n362_, N17 );
xor g021 ( new_n364_, new_n363_, keyIn_0_0 );
xnor g022 ( N418, new_n364_, keyIn_0_40 );
xnor g023 ( new_n366_, N390, keyIn_0_2 );
nand g024 ( new_n367_, N1, N26 );
nand g025 ( new_n368_, N13, N17 );
nor g026 ( new_n369_, new_n367_, new_n368_ );
xnor g027 ( new_n370_, new_n369_, keyIn_0_1 );
nand g028 ( N419, new_n370_, new_n366_ );
nand g029 ( new_n372_, N59, N75 );
nor g030 ( new_n373_, new_n372_, new_n347_ );
xor g031 ( new_n374_, new_n373_, keyIn_0_7 );
xnor g032 ( N420, new_n374_, keyIn_0_46 );
nand g033 ( new_n376_, N36, N59 );
nor g034 ( new_n377_, new_n376_, new_n347_ );
xnor g035 ( new_n378_, new_n377_, keyIn_0_9 );
xnor g036 ( N421, new_n378_, keyIn_0_47 );
nor g037 ( new_n380_, new_n376_, new_n343_ );
xnor g038 ( new_n381_, new_n380_, keyIn_0_10 );
xnor g039 ( N422, new_n381_, keyIn_0_48 );
not g040 ( new_n383_, N87 );
not g041 ( new_n384_, N88 );
nand g042 ( new_n385_, new_n383_, new_n384_ );
nand g043 ( new_n386_, new_n385_, keyIn_0_12 );
nor g044 ( new_n387_, keyIn_0_12, N87 );
nand g045 ( new_n388_, new_n387_, new_n384_ );
nand g046 ( new_n389_, new_n386_, new_n388_ );
nand g047 ( new_n390_, new_n389_, N90 );
xnor g048 ( N423, new_n390_, keyIn_0_50 );
xnor g049 ( new_n392_, new_n366_, keyIn_0_41 );
nand g050 ( new_n393_, new_n392_, new_n370_ );
xor g051 ( N446, new_n393_, keyIn_0_58 );
not g052 ( new_n395_, new_n367_ );
nand g053 ( new_n396_, new_n395_, N51 );
xnor g054 ( new_n397_, new_n396_, keyIn_0_43 );
xnor g055 ( N447, new_n397_, keyIn_0_60 );
nand g056 ( new_n399_, new_n362_, N55 );
nand g057 ( new_n400_, N29, N68 );
nor g058 ( new_n401_, new_n399_, new_n400_ );
xor g059 ( N448, new_n401_, keyIn_0_62 );
not g060 ( new_n403_, new_n399_ );
not g061 ( new_n404_, N74 );
nand g062 ( new_n405_, N59, N68 );
nor g063 ( new_n406_, new_n405_, new_n404_ );
nand g064 ( new_n407_, new_n403_, new_n406_ );
xnor g065 ( new_n408_, new_n407_, keyIn_0_45 );
xnor g066 ( N449, new_n408_, keyIn_0_63 );
nand g067 ( new_n410_, new_n389_, N89 );
xor g068 ( N450, new_n410_, keyIn_0_49 );
nor g069 ( new_n412_, N111, N116 );
xor g070 ( new_n413_, new_n412_, keyIn_0_17 );
nand g071 ( new_n414_, N111, N116 );
xor g072 ( new_n415_, new_n414_, keyIn_0_16 );
nand g073 ( new_n416_, new_n413_, new_n415_ );
xnor g074 ( new_n417_, new_n416_, keyIn_0_52 );
xor g075 ( new_n418_, new_n417_, keyIn_0_67 );
not g076 ( new_n419_, N121 );
not g077 ( new_n420_, N126 );
nand g078 ( new_n421_, new_n419_, new_n420_ );
nor g079 ( new_n422_, new_n421_, keyIn_0_18 );
nand g080 ( new_n423_, N121, N126 );
nand g081 ( new_n424_, new_n421_, keyIn_0_18 );
nand g082 ( new_n425_, new_n424_, new_n423_ );
nor g083 ( new_n426_, new_n425_, new_n422_ );
xor g084 ( new_n427_, new_n426_, keyIn_0_53 );
xor g085 ( new_n428_, new_n427_, keyIn_0_68 );
nand g086 ( new_n429_, new_n428_, new_n418_ );
nor g087 ( new_n430_, new_n429_, keyIn_0_78 );
nand g088 ( new_n431_, new_n429_, keyIn_0_78 );
nand g089 ( new_n432_, new_n427_, new_n417_ );
xnor g090 ( new_n433_, new_n432_, keyIn_0_69 );
nand g091 ( new_n434_, new_n431_, new_n433_ );
nor g092 ( new_n435_, new_n434_, new_n430_ );
xnor g093 ( new_n436_, new_n435_, keyIn_0_87 );
not g094 ( new_n437_, new_n436_ );
nor g095 ( new_n438_, new_n437_, N135 );
xor g096 ( new_n439_, new_n438_, keyIn_0_105 );
nand g097 ( new_n440_, new_n437_, N135 );
xor g098 ( new_n441_, new_n440_, keyIn_0_104 );
nand g099 ( new_n442_, new_n439_, new_n441_ );
xnor g100 ( new_n443_, new_n442_, keyIn_0_123 );
xnor g101 ( new_n444_, new_n443_, keyIn_0_129 );
not g102 ( new_n445_, N130 );
not g103 ( new_n446_, keyIn_0_13 );
nand g104 ( new_n447_, N91, N96 );
nand g105 ( new_n448_, new_n447_, new_n446_ );
not g106 ( new_n449_, keyIn_0_14 );
nor g107 ( new_n450_, N91, N96 );
nand g108 ( new_n451_, new_n450_, new_n449_ );
nand g109 ( new_n452_, new_n451_, new_n448_ );
not g110 ( new_n453_, new_n452_ );
nor g111 ( new_n454_, new_n450_, new_n449_ );
nor g112 ( new_n455_, new_n447_, new_n446_ );
nor g113 ( new_n456_, new_n454_, new_n455_ );
nand g114 ( new_n457_, new_n453_, new_n456_ );
xor g115 ( new_n458_, new_n457_, keyIn_0_51 );
xor g116 ( new_n459_, new_n458_, keyIn_0_64 );
not g117 ( new_n460_, keyIn_0_15 );
not g118 ( new_n461_, N101 );
not g119 ( new_n462_, N106 );
nand g120 ( new_n463_, new_n461_, new_n462_ );
nand g121 ( new_n464_, new_n463_, new_n460_ );
nor g122 ( new_n465_, new_n460_, N101 );
nand g123 ( new_n466_, new_n465_, new_n462_ );
nand g124 ( new_n467_, new_n466_, new_n464_ );
nand g125 ( new_n468_, N101, N106 );
nand g126 ( new_n469_, new_n467_, new_n468_ );
xor g127 ( new_n470_, new_n469_, keyIn_0_65 );
nand g128 ( new_n471_, new_n459_, new_n470_ );
nor g129 ( new_n472_, new_n471_, keyIn_0_77 );
nand g130 ( new_n473_, new_n471_, keyIn_0_77 );
nand g131 ( new_n474_, new_n458_, new_n469_ );
xor g132 ( new_n475_, new_n474_, keyIn_0_66 );
nand g133 ( new_n476_, new_n473_, new_n475_ );
nor g134 ( new_n477_, new_n476_, new_n472_ );
xor g135 ( new_n478_, new_n477_, keyIn_0_86 );
nand g136 ( new_n479_, new_n478_, new_n445_ );
xnor g137 ( new_n480_, new_n479_, keyIn_0_103 );
nor g138 ( new_n481_, new_n478_, new_n445_ );
xnor g139 ( new_n482_, new_n481_, keyIn_0_102 );
nand g140 ( new_n483_, new_n482_, new_n480_ );
xnor g141 ( new_n484_, new_n483_, keyIn_0_122 );
xnor g142 ( new_n485_, new_n484_, keyIn_0_128 );
nand g143 ( new_n486_, new_n444_, new_n485_ );
xnor g144 ( new_n487_, new_n486_, keyIn_0_138 );
nand g145 ( new_n488_, new_n443_, new_n484_ );
nand g146 ( new_n489_, new_n487_, new_n488_ );
xor g147 ( N767, new_n489_, keyIn_0_156 );
nand g148 ( new_n491_, N171, N177 );
nand g149 ( new_n492_, new_n491_, keyIn_0_27 );
not g150 ( new_n493_, new_n492_ );
nor g151 ( new_n494_, N171, N177 );
nor g152 ( new_n495_, new_n494_, keyIn_0_28 );
nor g153 ( new_n496_, new_n493_, new_n495_ );
nand g154 ( new_n497_, new_n494_, keyIn_0_28 );
not g155 ( new_n498_, new_n497_ );
nor g156 ( new_n499_, new_n491_, keyIn_0_27 );
nor g157 ( new_n500_, new_n498_, new_n499_ );
nand g158 ( new_n501_, new_n500_, new_n496_ );
xnor g159 ( new_n502_, new_n501_, keyIn_0_72 );
not g160 ( new_n503_, keyIn_0_25 );
nand g161 ( new_n504_, N159, N165 );
nand g162 ( new_n505_, new_n504_, new_n503_ );
not g163 ( new_n506_, keyIn_0_26 );
nor g164 ( new_n507_, N159, N165 );
nand g165 ( new_n508_, new_n507_, new_n506_ );
nand g166 ( new_n509_, new_n508_, new_n505_ );
not g167 ( new_n510_, new_n509_ );
nor g168 ( new_n511_, new_n507_, new_n506_ );
nor g169 ( new_n512_, new_n504_, new_n503_ );
nor g170 ( new_n513_, new_n511_, new_n512_ );
nand g171 ( new_n514_, new_n510_, new_n513_ );
xnor g172 ( new_n515_, new_n514_, keyIn_0_71 );
nor g173 ( new_n516_, new_n502_, new_n515_ );
xnor g174 ( new_n517_, new_n516_, keyIn_0_84 );
nand g175 ( new_n518_, new_n501_, new_n514_ );
nand g176 ( new_n519_, new_n517_, new_n518_ );
xnor g177 ( new_n520_, new_n519_, keyIn_0_101 );
nand g178 ( new_n521_, new_n520_, N130 );
xnor g179 ( new_n522_, new_n521_, keyIn_0_114 );
nor g180 ( new_n523_, new_n520_, N130 );
xnor g181 ( new_n524_, new_n523_, keyIn_0_115 );
nand g182 ( new_n525_, new_n524_, new_n522_ );
xnor g183 ( new_n526_, new_n525_, keyIn_0_136 );
not g184 ( new_n527_, N207 );
not g185 ( new_n528_, keyIn_0_30 );
nand g186 ( new_n529_, N195, N201 );
nand g187 ( new_n530_, new_n529_, new_n528_ );
not g188 ( new_n531_, keyIn_0_31 );
nor g189 ( new_n532_, N195, N201 );
nand g190 ( new_n533_, new_n532_, new_n531_ );
nand g191 ( new_n534_, new_n533_, new_n530_ );
not g192 ( new_n535_, new_n534_ );
nor g193 ( new_n536_, new_n532_, new_n531_ );
nor g194 ( new_n537_, new_n529_, new_n528_ );
nor g195 ( new_n538_, new_n536_, new_n537_ );
nand g196 ( new_n539_, new_n535_, new_n538_ );
xor g197 ( new_n540_, new_n539_, keyIn_0_57 );
xor g198 ( new_n541_, new_n540_, keyIn_0_73 );
nor g199 ( new_n542_, keyIn_0_29, N189 );
xor g200 ( new_n543_, new_n542_, keyIn_0_56 );
not g201 ( new_n544_, N183 );
nand g202 ( new_n545_, keyIn_0_29, N189 );
nand g203 ( new_n546_, new_n545_, new_n544_ );
xnor g204 ( new_n547_, new_n543_, new_n546_ );
nand g205 ( new_n548_, new_n541_, new_n547_ );
xor g206 ( new_n549_, new_n548_, keyIn_0_85 );
nor g207 ( new_n550_, new_n540_, new_n547_ );
xor g208 ( new_n551_, new_n550_, keyIn_0_74 );
nand g209 ( new_n552_, new_n549_, new_n551_ );
nor g210 ( new_n553_, new_n552_, new_n527_ );
xnor g211 ( new_n554_, new_n553_, keyIn_0_116 );
nand g212 ( new_n555_, new_n552_, new_n527_ );
nand g213 ( new_n556_, new_n554_, new_n555_ );
nor g214 ( new_n557_, new_n526_, new_n556_ );
xnor g215 ( new_n558_, new_n557_, keyIn_0_139 );
nand g216 ( new_n559_, new_n556_, new_n525_ );
xnor g217 ( new_n560_, new_n559_, keyIn_0_137 );
nand g218 ( new_n561_, new_n558_, new_n560_ );
xor g219 ( N768, new_n561_, keyIn_0_157 );
not g220 ( new_n563_, keyIn_0_215 );
not g221 ( new_n564_, N261 );
not g222 ( new_n565_, keyIn_0_135 );
not g223 ( new_n566_, keyIn_0_127 );
nand g224 ( new_n567_, new_n396_, keyIn_0_42 );
not g225 ( new_n568_, keyIn_0_42 );
not g226 ( new_n569_, N51 );
nor g227 ( new_n570_, new_n367_, new_n569_ );
nand g228 ( new_n571_, new_n570_, new_n568_ );
nand g229 ( new_n572_, new_n567_, new_n571_ );
nand g230 ( new_n573_, new_n572_, keyIn_0_59 );
not g231 ( new_n574_, keyIn_0_59 );
xnor g232 ( new_n575_, new_n570_, keyIn_0_42 );
nand g233 ( new_n576_, new_n575_, new_n574_ );
nand g234 ( new_n577_, new_n576_, new_n573_ );
nor g235 ( new_n578_, N17, N42 );
nor g236 ( new_n579_, new_n578_, keyIn_0_23 );
nand g237 ( new_n580_, N17, N42 );
nand g238 ( new_n581_, new_n580_, keyIn_0_24 );
not g239 ( new_n582_, new_n581_ );
nor g240 ( new_n583_, new_n582_, new_n579_ );
not g241 ( new_n584_, N17 );
nand g242 ( new_n585_, new_n584_, keyIn_0_23 );
nor g243 ( new_n586_, new_n585_, N42 );
nor g244 ( new_n587_, new_n580_, keyIn_0_24 );
nor g245 ( new_n588_, new_n586_, new_n587_ );
nand g246 ( new_n589_, new_n588_, new_n583_ );
nand g247 ( new_n590_, new_n589_, keyIn_0_55 );
nand g248 ( new_n591_, new_n577_, new_n590_ );
not g249 ( new_n592_, new_n591_ );
nand g250 ( new_n593_, N59, N156 );
not g251 ( new_n594_, new_n593_ );
not g252 ( new_n595_, keyIn_0_55 );
not g253 ( new_n596_, new_n585_ );
nand g254 ( new_n597_, new_n596_, new_n343_ );
nand g255 ( new_n598_, new_n597_, new_n595_ );
nor g256 ( new_n599_, new_n598_, new_n587_ );
nand g257 ( new_n600_, new_n599_, new_n583_ );
nand g258 ( new_n601_, new_n600_, new_n594_ );
not g259 ( new_n602_, new_n601_ );
nand g260 ( new_n603_, new_n592_, new_n602_ );
nand g261 ( new_n604_, new_n603_, keyIn_0_82 );
nand g262 ( new_n605_, N42, N59 );
not g263 ( new_n606_, new_n605_ );
nand g264 ( new_n607_, new_n606_, N75 );
xnor g265 ( new_n608_, new_n607_, keyIn_0_8 );
nand g266 ( new_n609_, N17, N51 );
nor g267 ( new_n610_, new_n361_, new_n609_ );
xor g268 ( new_n611_, new_n610_, keyIn_0_3 );
nand g269 ( new_n612_, new_n611_, new_n608_ );
xnor g270 ( new_n613_, new_n612_, keyIn_0_70 );
not g271 ( new_n614_, new_n579_ );
nand g272 ( new_n615_, new_n614_, new_n581_ );
not g273 ( new_n616_, new_n587_ );
nand g274 ( new_n617_, new_n597_, new_n616_ );
nor g275 ( new_n618_, new_n617_, new_n615_ );
nand g276 ( new_n619_, new_n618_, new_n595_ );
nor g277 ( new_n620_, new_n593_, keyIn_0_82 );
nand g278 ( new_n621_, new_n619_, new_n620_ );
nor g279 ( new_n622_, new_n591_, new_n621_ );
nor g280 ( new_n623_, new_n613_, new_n622_ );
nand g281 ( new_n624_, new_n604_, new_n623_ );
nand g282 ( new_n625_, new_n624_, keyIn_0_88 );
not g283 ( new_n626_, keyIn_0_88 );
not g284 ( new_n627_, keyIn_0_82 );
nor g285 ( new_n628_, new_n591_, new_n601_ );
nor g286 ( new_n629_, new_n628_, new_n627_ );
not g287 ( new_n630_, keyIn_0_70 );
xnor g288 ( new_n631_, new_n612_, new_n630_ );
not g289 ( new_n632_, new_n621_ );
nand g290 ( new_n633_, new_n592_, new_n632_ );
nand g291 ( new_n634_, new_n633_, new_n631_ );
nor g292 ( new_n635_, new_n634_, new_n629_ );
nand g293 ( new_n636_, new_n635_, new_n626_ );
nand g294 ( new_n637_, new_n636_, new_n625_ );
nand g295 ( new_n638_, new_n637_, N126 );
not g296 ( new_n639_, keyIn_0_97 );
xnor g297 ( new_n640_, new_n593_, keyIn_0_22 );
not g298 ( new_n641_, new_n640_ );
nand g299 ( new_n642_, new_n577_, new_n641_ );
nor g300 ( new_n643_, new_n642_, new_n584_ );
nand g301 ( new_n644_, new_n643_, keyIn_0_83 );
not g302 ( new_n645_, N1 );
nor g303 ( new_n646_, new_n643_, keyIn_0_83 );
nor g304 ( new_n647_, new_n646_, new_n645_ );
nand g305 ( new_n648_, new_n647_, new_n644_ );
xnor g306 ( new_n649_, new_n648_, new_n639_ );
nand g307 ( new_n650_, new_n649_, N153 );
nand g308 ( new_n651_, new_n650_, new_n638_ );
nor g309 ( new_n652_, new_n651_, new_n566_ );
not g310 ( new_n653_, new_n652_ );
not g311 ( new_n654_, N55 );
nor g312 ( new_n655_, new_n344_, new_n347_ );
nand g313 ( new_n656_, new_n577_, new_n655_ );
nor g314 ( new_n657_, new_n656_, new_n654_ );
nand g315 ( new_n658_, new_n657_, keyIn_0_81 );
xnor g316 ( new_n659_, keyIn_0_19, N268 );
xnor g317 ( new_n660_, new_n659_, keyIn_0_54 );
not g318 ( new_n661_, new_n660_ );
nor g319 ( new_n662_, new_n657_, keyIn_0_81 );
nor g320 ( new_n663_, new_n662_, new_n661_ );
nand g321 ( new_n664_, new_n663_, new_n658_ );
not g322 ( new_n665_, new_n664_ );
not g323 ( new_n666_, new_n638_ );
not g324 ( new_n667_, N153 );
nand g325 ( new_n668_, new_n648_, keyIn_0_97 );
not g326 ( new_n669_, new_n644_ );
not g327 ( new_n670_, keyIn_0_83 );
xnor g328 ( new_n671_, new_n572_, new_n574_ );
nor g329 ( new_n672_, new_n671_, new_n640_ );
nand g330 ( new_n673_, new_n672_, N17 );
nand g331 ( new_n674_, new_n673_, new_n670_ );
nand g332 ( new_n675_, new_n674_, N1 );
nor g333 ( new_n676_, new_n675_, new_n669_ );
nand g334 ( new_n677_, new_n676_, new_n639_ );
nand g335 ( new_n678_, new_n677_, new_n668_ );
nor g336 ( new_n679_, new_n678_, new_n667_ );
nor g337 ( new_n680_, new_n679_, new_n666_ );
nor g338 ( new_n681_, new_n680_, keyIn_0_127 );
nor g339 ( new_n682_, new_n681_, new_n665_ );
nand g340 ( new_n683_, new_n682_, new_n653_ );
nand g341 ( new_n684_, new_n683_, new_n565_ );
nand g342 ( new_n685_, new_n651_, new_n566_ );
nand g343 ( new_n686_, new_n685_, new_n664_ );
nor g344 ( new_n687_, new_n686_, new_n652_ );
nand g345 ( new_n688_, new_n687_, keyIn_0_135 );
nand g346 ( new_n689_, new_n684_, new_n688_ );
nor g347 ( new_n690_, new_n689_, N201 );
xnor g348 ( new_n691_, new_n690_, keyIn_0_154 );
nand g349 ( new_n692_, new_n689_, N201 );
nand g350 ( new_n693_, new_n691_, new_n692_ );
nor g351 ( new_n694_, new_n693_, new_n564_ );
xnor g352 ( new_n695_, new_n694_, keyIn_0_192 );
nand g353 ( new_n696_, new_n693_, new_n564_ );
nand g354 ( new_n697_, new_n695_, new_n696_ );
nor g355 ( new_n698_, new_n697_, keyIn_0_209 );
nand g356 ( new_n699_, new_n697_, keyIn_0_209 );
nand g357 ( new_n700_, new_n699_, N219 );
nor g358 ( new_n701_, new_n700_, new_n698_ );
nand g359 ( new_n702_, new_n701_, new_n563_ );
nor g360 ( new_n703_, new_n701_, new_n563_ );
not g361 ( new_n704_, N228 );
nor g362 ( new_n705_, new_n693_, new_n704_ );
xnor g363 ( new_n706_, new_n705_, keyIn_0_193 );
xnor g364 ( new_n707_, new_n692_, keyIn_0_172 );
nand g365 ( new_n708_, new_n707_, N237 );
xnor g366 ( new_n709_, new_n708_, keyIn_0_194 );
nand g367 ( new_n710_, new_n706_, new_n709_ );
xnor g368 ( new_n711_, new_n710_, keyIn_0_210 );
not g369 ( new_n712_, keyIn_0_155 );
nand g370 ( new_n713_, new_n689_, N246 );
nor g371 ( new_n714_, new_n713_, new_n712_ );
nand g372 ( new_n715_, new_n713_, new_n712_ );
nand g373 ( new_n716_, N255, N267 );
nand g374 ( new_n717_, new_n716_, keyIn_0_39 );
not g375 ( new_n718_, new_n717_ );
not g376 ( new_n719_, N267 );
not g377 ( new_n720_, keyIn_0_39 );
nand g378 ( new_n721_, new_n720_, N255 );
nor g379 ( new_n722_, new_n721_, new_n719_ );
nor g380 ( new_n723_, new_n722_, new_n718_ );
nand g381 ( new_n724_, new_n715_, new_n723_ );
nor g382 ( new_n725_, new_n724_, new_n714_ );
xor g383 ( new_n726_, new_n725_, keyIn_0_173 );
nand g384 ( new_n727_, N68, N72 );
nor g385 ( new_n728_, new_n605_, new_n727_ );
xor g386 ( new_n729_, new_n728_, keyIn_0_4 );
nand g387 ( new_n730_, new_n729_, new_n403_ );
xnor g388 ( new_n731_, new_n730_, keyIn_0_44 );
nand g389 ( new_n732_, new_n731_, N73 );
xnor g390 ( new_n733_, new_n732_, keyIn_0_61 );
xor g391 ( new_n734_, new_n733_, keyIn_0_76 );
nand g392 ( new_n735_, new_n734_, N201 );
nand g393 ( new_n736_, N121, N210 );
xor g394 ( new_n737_, new_n736_, keyIn_0_38 );
nand g395 ( new_n738_, new_n735_, new_n737_ );
nor g396 ( new_n739_, new_n726_, new_n738_ );
nand g397 ( new_n740_, new_n711_, new_n739_ );
nor g398 ( new_n741_, new_n703_, new_n740_ );
nand g399 ( new_n742_, new_n741_, new_n702_ );
xnor g400 ( new_n743_, new_n742_, keyIn_0_223 );
xnor g401 ( new_n744_, new_n743_, keyIn_0_229 );
xnor g402 ( N850, new_n744_, keyIn_0_234 );
not g403 ( new_n746_, keyIn_0_111 );
nand g404 ( new_n747_, new_n637_, N111 );
nor g405 ( new_n748_, new_n747_, new_n746_ );
nand g406 ( new_n749_, new_n649_, N143 );
nand g407 ( new_n750_, new_n747_, new_n746_ );
nand g408 ( new_n751_, new_n749_, new_n750_ );
nor g409 ( new_n752_, new_n751_, new_n748_ );
xor g410 ( new_n753_, new_n752_, keyIn_0_126 );
xor g411 ( new_n754_, new_n664_, keyIn_0_98 );
nand g412 ( new_n755_, new_n753_, new_n754_ );
xnor g413 ( new_n756_, new_n755_, keyIn_0_132 );
nand g414 ( new_n757_, new_n756_, new_n544_ );
xnor g415 ( new_n758_, new_n757_, keyIn_0_150 );
not g416 ( new_n759_, new_n756_ );
nand g417 ( new_n760_, new_n759_, N183 );
xor g418 ( new_n761_, new_n760_, keyIn_0_149 );
nand g419 ( new_n762_, new_n761_, new_n758_ );
xnor g420 ( new_n763_, new_n762_, keyIn_0_165 );
not g421 ( new_n764_, keyIn_0_204 );
not g422 ( new_n765_, N146 );
nor g423 ( new_n766_, new_n678_, new_n765_ );
nand g424 ( new_n767_, new_n637_, N116 );
xor g425 ( new_n768_, new_n664_, keyIn_0_99 );
nand g426 ( new_n769_, new_n768_, new_n767_ );
nor g427 ( new_n770_, new_n769_, new_n766_ );
xor g428 ( new_n771_, new_n770_, keyIn_0_133 );
not g429 ( new_n772_, new_n771_ );
nor g430 ( new_n773_, new_n772_, N189 );
not g431 ( new_n774_, new_n773_ );
not g432 ( new_n775_, N195 );
not g433 ( new_n776_, keyIn_0_134 );
nand g434 ( new_n777_, new_n649_, N149 );
nand g435 ( new_n778_, new_n777_, keyIn_0_112 );
not g436 ( new_n779_, keyIn_0_112 );
not g437 ( new_n780_, N149 );
nor g438 ( new_n781_, new_n678_, new_n780_ );
nand g439 ( new_n782_, new_n781_, new_n779_ );
nand g440 ( new_n783_, new_n778_, new_n782_ );
nand g441 ( new_n784_, new_n637_, N121 );
nor g442 ( new_n785_, new_n784_, keyIn_0_113 );
nand g443 ( new_n786_, new_n784_, keyIn_0_113 );
xnor g444 ( new_n787_, new_n664_, keyIn_0_100 );
nand g445 ( new_n788_, new_n786_, new_n787_ );
nor g446 ( new_n789_, new_n788_, new_n785_ );
nand g447 ( new_n790_, new_n783_, new_n789_ );
xnor g448 ( new_n791_, new_n790_, new_n776_ );
nand g449 ( new_n792_, new_n791_, new_n775_ );
xor g450 ( new_n793_, new_n792_, keyIn_0_152 );
nand g451 ( new_n794_, new_n691_, N261 );
nor g452 ( new_n795_, new_n794_, new_n793_ );
nand g453 ( new_n796_, new_n795_, new_n774_ );
nand g454 ( new_n797_, new_n796_, keyIn_0_176 );
not g455 ( new_n798_, keyIn_0_172 );
xnor g456 ( new_n799_, new_n692_, new_n798_ );
nor g457 ( new_n800_, new_n799_, new_n793_ );
nand g458 ( new_n801_, new_n800_, new_n774_ );
nand g459 ( new_n802_, new_n801_, keyIn_0_197 );
nand g460 ( new_n803_, new_n772_, N189 );
not g461 ( new_n804_, new_n803_ );
xnor g462 ( new_n805_, new_n790_, keyIn_0_134 );
nand g463 ( new_n806_, new_n805_, N195 );
nand g464 ( new_n807_, new_n806_, keyIn_0_169 );
not g465 ( new_n808_, keyIn_0_169 );
nor g466 ( new_n809_, new_n791_, new_n775_ );
nand g467 ( new_n810_, new_n809_, new_n808_ );
nand g468 ( new_n811_, new_n810_, new_n807_ );
nor g469 ( new_n812_, new_n811_, new_n773_ );
xnor g470 ( new_n813_, new_n812_, keyIn_0_196 );
nor g471 ( new_n814_, new_n813_, new_n804_ );
nand g472 ( new_n815_, new_n814_, new_n802_ );
not g473 ( new_n816_, keyIn_0_197 );
xnor g474 ( new_n817_, new_n792_, keyIn_0_152 );
nand g475 ( new_n818_, new_n707_, new_n817_ );
nor g476 ( new_n819_, new_n818_, new_n773_ );
nand g477 ( new_n820_, new_n819_, new_n816_ );
nor g478 ( new_n821_, new_n773_, keyIn_0_176 );
nand g479 ( new_n822_, new_n795_, new_n821_ );
nand g480 ( new_n823_, new_n822_, new_n820_ );
nor g481 ( new_n824_, new_n815_, new_n823_ );
nand g482 ( new_n825_, new_n824_, new_n797_ );
nand g483 ( new_n826_, new_n825_, new_n764_ );
not g484 ( new_n827_, new_n797_ );
nor g485 ( new_n828_, new_n819_, new_n816_ );
xnor g486 ( new_n829_, new_n806_, new_n808_ );
nand g487 ( new_n830_, new_n829_, new_n774_ );
nand g488 ( new_n831_, new_n830_, keyIn_0_196 );
not g489 ( new_n832_, keyIn_0_196 );
nand g490 ( new_n833_, new_n812_, new_n832_ );
nand g491 ( new_n834_, new_n831_, new_n833_ );
nand g492 ( new_n835_, new_n834_, new_n803_ );
nor g493 ( new_n836_, new_n828_, new_n835_ );
nor g494 ( new_n837_, new_n801_, keyIn_0_197 );
not g495 ( new_n838_, keyIn_0_154 );
xnor g496 ( new_n839_, new_n690_, new_n838_ );
nor g497 ( new_n840_, new_n839_, new_n564_ );
nand g498 ( new_n841_, new_n840_, new_n817_ );
not g499 ( new_n842_, new_n821_ );
nor g500 ( new_n843_, new_n841_, new_n842_ );
nor g501 ( new_n844_, new_n843_, new_n837_ );
nand g502 ( new_n845_, new_n844_, new_n836_ );
nor g503 ( new_n846_, new_n845_, new_n827_ );
nand g504 ( new_n847_, new_n846_, keyIn_0_204 );
nand g505 ( new_n848_, new_n847_, new_n826_ );
nor g506 ( new_n849_, new_n848_, new_n763_ );
nand g507 ( new_n850_, new_n849_, keyIn_0_211 );
not g508 ( new_n851_, new_n763_ );
not g509 ( new_n852_, new_n848_ );
nor g510 ( new_n853_, new_n852_, new_n851_ );
nor g511 ( new_n854_, new_n849_, keyIn_0_211 );
nor g512 ( new_n855_, new_n854_, new_n853_ );
nand g513 ( new_n856_, new_n855_, new_n850_ );
nor g514 ( new_n857_, new_n856_, keyIn_0_216 );
nand g515 ( new_n858_, new_n856_, keyIn_0_216 );
nand g516 ( new_n859_, new_n858_, N219 );
nor g517 ( new_n860_, new_n859_, new_n857_ );
xnor g518 ( new_n861_, new_n860_, keyIn_0_220 );
nand g519 ( new_n862_, N106, N210 );
nand g520 ( new_n863_, new_n862_, keyIn_0_34 );
not g521 ( new_n864_, new_n863_ );
not g522 ( new_n865_, N210 );
not g523 ( new_n866_, keyIn_0_34 );
nand g524 ( new_n867_, new_n866_, N106 );
nor g525 ( new_n868_, new_n867_, new_n865_ );
nor g526 ( new_n869_, new_n868_, new_n864_ );
nand g527 ( new_n870_, new_n861_, new_n869_ );
nor g528 ( new_n871_, new_n870_, keyIn_0_226 );
nand g529 ( new_n872_, new_n870_, keyIn_0_226 );
nand g530 ( new_n873_, new_n763_, N228 );
not g531 ( new_n874_, new_n761_ );
nand g532 ( new_n875_, new_n874_, N237 );
xnor g533 ( new_n876_, new_n875_, keyIn_0_186 );
nand g534 ( new_n877_, new_n873_, new_n876_ );
xnor g535 ( new_n878_, new_n877_, keyIn_0_205 );
nand g536 ( new_n879_, new_n759_, N246 );
nand g537 ( new_n880_, new_n734_, N183 );
xnor g538 ( new_n881_, new_n880_, keyIn_0_121 );
nand g539 ( new_n882_, new_n879_, new_n881_ );
xor g540 ( new_n883_, new_n882_, keyIn_0_166 );
nor g541 ( new_n884_, new_n878_, new_n883_ );
nand g542 ( new_n885_, new_n872_, new_n884_ );
nor g543 ( new_n886_, new_n885_, new_n871_ );
xnor g544 ( new_n887_, new_n886_, keyIn_0_233 );
xnor g545 ( new_n888_, new_n887_, keyIn_0_238 );
xor g546 ( N863, new_n888_, keyIn_0_245 );
not g547 ( new_n890_, keyIn_0_221 );
not g548 ( new_n891_, keyIn_0_175 );
nand g549 ( new_n892_, new_n841_, new_n891_ );
xnor g550 ( new_n893_, new_n811_, keyIn_0_189 );
nand g551 ( new_n894_, new_n892_, new_n893_ );
nand g552 ( new_n895_, new_n795_, keyIn_0_175 );
xnor g553 ( new_n896_, new_n818_, keyIn_0_195 );
nand g554 ( new_n897_, new_n896_, new_n895_ );
nor g555 ( new_n898_, new_n897_, new_n894_ );
xnor g556 ( new_n899_, new_n898_, keyIn_0_206 );
nor g557 ( new_n900_, new_n804_, new_n773_ );
xnor g558 ( new_n901_, new_n900_, keyIn_0_167 );
nor g559 ( new_n902_, new_n899_, new_n901_ );
xor g560 ( new_n903_, new_n902_, keyIn_0_212 );
nand g561 ( new_n904_, new_n899_, new_n901_ );
nand g562 ( new_n905_, new_n904_, N219 );
not g563 ( new_n906_, new_n905_ );
nand g564 ( new_n907_, new_n903_, new_n906_ );
nor g565 ( new_n908_, new_n907_, new_n890_ );
not g566 ( new_n909_, keyIn_0_35 );
nand g567 ( new_n910_, N111, N210 );
nand g568 ( new_n911_, new_n910_, new_n909_ );
nand g569 ( new_n912_, keyIn_0_35, N111 );
not g570 ( new_n913_, new_n912_ );
nand g571 ( new_n914_, new_n913_, N210 );
nand g572 ( new_n915_, new_n914_, new_n911_ );
nand g573 ( new_n916_, new_n907_, new_n890_ );
nand g574 ( new_n917_, new_n916_, new_n915_ );
nor g575 ( new_n918_, new_n917_, new_n908_ );
xor g576 ( new_n919_, new_n918_, keyIn_0_227 );
nor g577 ( new_n920_, new_n901_, new_n704_ );
xnor g578 ( new_n921_, new_n920_, keyIn_0_187 );
nand g579 ( new_n922_, new_n772_, N246 );
xnor g580 ( new_n923_, new_n922_, keyIn_0_151 );
nand g581 ( new_n924_, N255, N259 );
nand g582 ( new_n925_, new_n924_, keyIn_0_36 );
not g583 ( new_n926_, N255 );
nor g584 ( new_n927_, new_n926_, keyIn_0_36 );
nand g585 ( new_n928_, new_n927_, N259 );
nand g586 ( new_n929_, new_n928_, new_n925_ );
nand g587 ( new_n930_, new_n923_, new_n929_ );
xnor g588 ( new_n931_, new_n930_, keyIn_0_168 );
not g589 ( new_n932_, keyIn_0_188 );
nand g590 ( new_n933_, new_n804_, N237 );
nor g591 ( new_n934_, new_n933_, new_n932_ );
nand g592 ( new_n935_, new_n734_, N189 );
nand g593 ( new_n936_, new_n933_, new_n932_ );
nand g594 ( new_n937_, new_n936_, new_n935_ );
nor g595 ( new_n938_, new_n937_, new_n934_ );
nand g596 ( new_n939_, new_n931_, new_n938_ );
nor g597 ( new_n940_, new_n921_, new_n939_ );
nand g598 ( new_n941_, new_n919_, new_n940_ );
xor g599 ( new_n942_, new_n941_, keyIn_0_239 );
xnor g600 ( N864, new_n942_, keyIn_0_246 );
not g601 ( new_n944_, keyIn_0_228 );
not g602 ( new_n945_, keyIn_0_217 );
nand g603 ( new_n946_, new_n817_, new_n806_ );
xnor g604 ( new_n947_, new_n946_, keyIn_0_170 );
xnor g605 ( new_n948_, new_n794_, keyIn_0_174 );
nor g606 ( new_n949_, new_n948_, new_n707_ );
xnor g607 ( new_n950_, new_n949_, keyIn_0_207 );
nor g608 ( new_n951_, new_n950_, new_n947_ );
xnor g609 ( new_n952_, new_n951_, keyIn_0_213 );
nand g610 ( new_n953_, new_n950_, new_n947_ );
xor g611 ( new_n954_, new_n953_, keyIn_0_214 );
nand g612 ( new_n955_, new_n954_, new_n952_ );
nor g613 ( new_n956_, new_n955_, new_n945_ );
nand g614 ( new_n957_, new_n955_, new_n945_ );
nand g615 ( new_n958_, new_n957_, N219 );
nor g616 ( new_n959_, new_n958_, new_n956_ );
xor g617 ( new_n960_, new_n959_, keyIn_0_222 );
nand g618 ( new_n961_, N116, N210 );
nand g619 ( new_n962_, new_n960_, new_n961_ );
nor g620 ( new_n963_, new_n962_, new_n944_ );
nand g621 ( new_n964_, new_n962_, new_n944_ );
nand g622 ( new_n965_, new_n947_, N228 );
nor g623 ( new_n966_, new_n965_, keyIn_0_190 );
nand g624 ( new_n967_, new_n829_, N237 );
xnor g625 ( new_n968_, new_n967_, keyIn_0_191 );
nand g626 ( new_n969_, new_n965_, keyIn_0_190 );
nand g627 ( new_n970_, new_n969_, new_n968_ );
nor g628 ( new_n971_, new_n970_, new_n966_ );
xnor g629 ( new_n972_, new_n971_, keyIn_0_208 );
nand g630 ( new_n973_, new_n734_, N195 );
nand g631 ( new_n974_, new_n805_, N246 );
xnor g632 ( new_n975_, new_n974_, keyIn_0_153 );
not g633 ( new_n976_, keyIn_0_37 );
nand g634 ( new_n977_, N255, N260 );
nand g635 ( new_n978_, new_n977_, new_n976_ );
nand g636 ( new_n979_, keyIn_0_37, N255 );
not g637 ( new_n980_, new_n979_ );
nand g638 ( new_n981_, new_n980_, N260 );
nand g639 ( new_n982_, new_n981_, new_n978_ );
nand g640 ( new_n983_, new_n975_, new_n982_ );
xor g641 ( new_n984_, new_n983_, keyIn_0_171 );
nand g642 ( new_n985_, new_n984_, new_n973_ );
nor g643 ( new_n986_, new_n972_, new_n985_ );
nand g644 ( new_n987_, new_n964_, new_n986_ );
nor g645 ( new_n988_, new_n987_, new_n963_ );
xnor g646 ( new_n989_, new_n988_, keyIn_0_240 );
xnor g647 ( N865, new_n989_, keyIn_0_247 );
not g648 ( new_n991_, keyIn_0_235 );
nor g649 ( new_n992_, new_n642_, new_n654_ );
xnor g650 ( new_n993_, new_n992_, keyIn_0_79 );
nand g651 ( new_n994_, new_n993_, N146 );
xnor g652 ( new_n995_, new_n994_, keyIn_0_91 );
nor g653 ( new_n996_, new_n656_, new_n584_ );
not g654 ( new_n997_, new_n996_ );
nor g655 ( new_n998_, new_n997_, keyIn_0_80 );
nand g656 ( new_n999_, new_n997_, keyIn_0_80 );
nand g657 ( new_n1000_, new_n999_, new_n659_ );
nor g658 ( new_n1001_, new_n1000_, new_n998_ );
xnor g659 ( new_n1002_, new_n1001_, keyIn_0_92 );
nand g660 ( new_n1003_, new_n1002_, new_n995_ );
xnor g661 ( new_n1004_, new_n1003_, keyIn_0_107 );
nand g662 ( new_n1005_, new_n637_, N96 );
nor g663 ( new_n1006_, new_n1005_, keyIn_0_106 );
nand g664 ( new_n1007_, new_n1005_, keyIn_0_106 );
nand g665 ( new_n1008_, N51, N138 );
xnor g666 ( new_n1009_, new_n1008_, keyIn_0_20 );
nand g667 ( new_n1010_, new_n1007_, new_n1009_ );
nor g668 ( new_n1011_, new_n1010_, new_n1006_ );
nand g669 ( new_n1012_, new_n1004_, new_n1011_ );
xnor g670 ( new_n1013_, new_n1012_, keyIn_0_130 );
nor g671 ( new_n1014_, new_n1013_, N165 );
xnor g672 ( new_n1015_, new_n1014_, keyIn_0_144 );
not g673 ( new_n1016_, new_n1015_ );
not g674 ( new_n1017_, N171 );
nand g675 ( new_n1018_, new_n993_, N149 );
xnor g676 ( new_n1019_, new_n1018_, keyIn_0_93 );
xnor g677 ( new_n1020_, new_n1001_, keyIn_0_94 );
nand g678 ( new_n1021_, new_n1020_, new_n1019_ );
xor g679 ( new_n1022_, new_n1021_, keyIn_0_108 );
nand g680 ( new_n1023_, new_n637_, N101 );
not g681 ( new_n1024_, keyIn_0_21 );
nand g682 ( new_n1025_, N17, N138 );
nand g683 ( new_n1026_, new_n1025_, new_n1024_ );
nand g684 ( new_n1027_, keyIn_0_21, N17 );
not g685 ( new_n1028_, new_n1027_ );
nand g686 ( new_n1029_, new_n1028_, N138 );
nand g687 ( new_n1030_, new_n1029_, new_n1026_ );
nand g688 ( new_n1031_, new_n1023_, new_n1030_ );
xnor g689 ( new_n1032_, new_n1031_, keyIn_0_124 );
nand g690 ( new_n1033_, new_n1022_, new_n1032_ );
xor g691 ( new_n1034_, new_n1033_, keyIn_0_131 );
not g692 ( new_n1035_, new_n1034_ );
nand g693 ( new_n1036_, new_n1035_, new_n1017_ );
xor g694 ( new_n1037_, new_n1036_, keyIn_0_145 );
nor g695 ( new_n1038_, new_n1037_, new_n1016_ );
not g696 ( new_n1039_, new_n1038_ );
nand g697 ( new_n1040_, new_n848_, new_n758_ );
xor g698 ( new_n1041_, new_n761_, keyIn_0_185 );
nand g699 ( new_n1042_, new_n1040_, new_n1041_ );
not g700 ( new_n1043_, keyIn_0_95 );
not g701 ( new_n1044_, new_n993_ );
nor g702 ( new_n1045_, new_n1044_, new_n667_ );
not g703 ( new_n1046_, new_n1045_ );
nand g704 ( new_n1047_, new_n1046_, new_n1043_ );
not g705 ( new_n1048_, keyIn_0_96 );
not g706 ( new_n1049_, new_n1001_ );
nand g707 ( new_n1050_, new_n1049_, new_n1048_ );
nand g708 ( new_n1051_, new_n1047_, new_n1050_ );
nand g709 ( new_n1052_, new_n1001_, keyIn_0_96 );
nand g710 ( new_n1053_, new_n1045_, keyIn_0_95 );
nand g711 ( new_n1054_, new_n1053_, new_n1052_ );
nor g712 ( new_n1055_, new_n1051_, new_n1054_ );
xor g713 ( new_n1056_, new_n1055_, keyIn_0_110 );
nand g714 ( new_n1057_, new_n637_, N106 );
xor g715 ( new_n1058_, new_n1057_, keyIn_0_109 );
nand g716 ( new_n1059_, N138, N152 );
nand g717 ( new_n1060_, new_n1058_, new_n1059_ );
xnor g718 ( new_n1061_, new_n1060_, keyIn_0_125 );
nand g719 ( new_n1062_, new_n1061_, new_n1056_ );
nor g720 ( new_n1063_, new_n1062_, N177 );
xor g721 ( new_n1064_, new_n1063_, keyIn_0_147 );
nand g722 ( new_n1065_, new_n1042_, new_n1064_ );
nor g723 ( new_n1066_, new_n1065_, new_n1039_ );
xnor g724 ( new_n1067_, new_n1066_, keyIn_0_225 );
nand g725 ( new_n1068_, new_n1062_, N177 );
xnor g726 ( new_n1069_, new_n1068_, keyIn_0_146 );
xnor g727 ( new_n1070_, new_n1069_, keyIn_0_162 );
not g728 ( new_n1071_, new_n1070_ );
nor g729 ( new_n1072_, new_n1039_, new_n1071_ );
not g730 ( new_n1073_, new_n1072_ );
nor g731 ( new_n1074_, new_n1073_, keyIn_0_200 );
nand g732 ( new_n1075_, new_n1073_, keyIn_0_200 );
nor g733 ( new_n1076_, new_n1035_, new_n1017_ );
not g734 ( new_n1077_, new_n1076_ );
nor g735 ( new_n1078_, new_n1016_, new_n1077_ );
not g736 ( new_n1079_, new_n1078_ );
nor g737 ( new_n1080_, new_n1079_, keyIn_0_199 );
nand g738 ( new_n1081_, new_n1079_, keyIn_0_199 );
nand g739 ( new_n1082_, new_n1013_, N165 );
xnor g740 ( new_n1083_, new_n1082_, keyIn_0_143 );
xnor g741 ( new_n1084_, new_n1083_, keyIn_0_179 );
nand g742 ( new_n1085_, new_n1081_, new_n1084_ );
nor g743 ( new_n1086_, new_n1085_, new_n1080_ );
nand g744 ( new_n1087_, new_n1075_, new_n1086_ );
nor g745 ( new_n1088_, new_n1087_, new_n1074_ );
nand g746 ( new_n1089_, new_n1067_, new_n1088_ );
not g747 ( new_n1090_, N159 );
nand g748 ( new_n1091_, new_n993_, N143 );
nor g749 ( new_n1092_, new_n1091_, keyIn_0_89 );
nand g750 ( new_n1093_, new_n1091_, keyIn_0_89 );
not g751 ( new_n1094_, keyIn_0_90 );
nand g752 ( new_n1095_, new_n1049_, new_n1094_ );
nand g753 ( new_n1096_, new_n1095_, new_n1093_ );
nor g754 ( new_n1097_, new_n1096_, new_n1092_ );
not g755 ( new_n1098_, new_n1097_ );
nand g756 ( new_n1099_, new_n637_, N91 );
nor g757 ( new_n1100_, new_n1049_, new_n1094_ );
nand g758 ( new_n1101_, N8, N138 );
not g759 ( new_n1102_, new_n1101_ );
nor g760 ( new_n1103_, new_n1100_, new_n1102_ );
nand g761 ( new_n1104_, new_n1103_, new_n1099_ );
nor g762 ( new_n1105_, new_n1098_, new_n1104_ );
nand g763 ( new_n1106_, new_n1105_, new_n1090_ );
xor g764 ( new_n1107_, new_n1106_, keyIn_0_141 );
nand g765 ( new_n1108_, new_n1089_, new_n1107_ );
nor g766 ( new_n1109_, new_n1108_, new_n991_ );
not g767 ( new_n1110_, new_n1105_ );
nand g768 ( new_n1111_, new_n1110_, N159 );
xor g769 ( new_n1112_, new_n1111_, keyIn_0_140 );
xnor g770 ( new_n1113_, new_n1112_, keyIn_0_177 );
nand g771 ( new_n1114_, new_n1108_, new_n991_ );
nand g772 ( new_n1115_, new_n1114_, new_n1113_ );
nor g773 ( new_n1116_, new_n1115_, new_n1109_ );
xnor g774 ( new_n1117_, new_n1116_, keyIn_0_241 );
xnor g775 ( N866, new_n1117_, keyIn_0_248 );
nand g776 ( new_n1119_, new_n1064_, new_n1069_ );
xor g777 ( new_n1120_, new_n1119_, keyIn_0_163 );
nand g778 ( new_n1121_, new_n1042_, new_n1120_ );
xor g779 ( new_n1122_, new_n1121_, keyIn_0_219 );
nor g780 ( new_n1123_, new_n1042_, new_n1120_ );
nor g781 ( new_n1124_, new_n1123_, keyIn_0_218 );
nand g782 ( new_n1125_, new_n1123_, keyIn_0_218 );
nand g783 ( new_n1126_, new_n1125_, N219 );
nor g784 ( new_n1127_, new_n1126_, new_n1124_ );
nand g785 ( new_n1128_, new_n1127_, new_n1122_ );
nand g786 ( new_n1129_, new_n1120_, N228 );
xor g787 ( new_n1130_, new_n1129_, keyIn_0_184 );
nand g788 ( new_n1131_, new_n1070_, N237 );
nand g789 ( new_n1132_, new_n1062_, N246 );
xor g790 ( new_n1133_, new_n1132_, keyIn_0_148 );
nand g791 ( new_n1134_, new_n734_, N177 );
xor g792 ( new_n1135_, new_n1134_, keyIn_0_120 );
nor g793 ( new_n1136_, new_n1133_, new_n1135_ );
nor g794 ( new_n1137_, new_n1136_, keyIn_0_164 );
nand g795 ( new_n1138_, N101, N210 );
nand g796 ( new_n1139_, new_n1136_, keyIn_0_164 );
nand g797 ( new_n1140_, new_n1139_, new_n1138_ );
nor g798 ( new_n1141_, new_n1140_, new_n1137_ );
nand g799 ( new_n1142_, new_n1141_, new_n1131_ );
nor g800 ( new_n1143_, new_n1130_, new_n1142_ );
nand g801 ( new_n1144_, new_n1128_, new_n1143_ );
xnor g802 ( new_n1145_, new_n1144_, keyIn_0_244 );
xnor g803 ( N874, new_n1145_, keyIn_0_253 );
not g804 ( new_n1147_, keyIn_0_251 );
not g805 ( new_n1148_, keyIn_0_249 );
not g806 ( new_n1149_, new_n1107_ );
not g807 ( new_n1150_, new_n1112_ );
nor g808 ( new_n1151_, new_n1150_, new_n1149_ );
xor g809 ( new_n1152_, new_n1151_, keyIn_0_158 );
not g810 ( new_n1153_, new_n1152_ );
nand g811 ( new_n1154_, new_n1089_, new_n1153_ );
nand g812 ( new_n1155_, new_n1154_, keyIn_0_230 );
not g813 ( new_n1156_, keyIn_0_230 );
not g814 ( new_n1157_, keyIn_0_225 );
xnor g815 ( new_n1158_, new_n1066_, new_n1157_ );
not g816 ( new_n1159_, new_n1088_ );
nor g817 ( new_n1160_, new_n1158_, new_n1159_ );
nor g818 ( new_n1161_, new_n1160_, new_n1152_ );
nand g819 ( new_n1162_, new_n1161_, new_n1156_ );
nand g820 ( new_n1163_, new_n1162_, new_n1155_ );
nor g821 ( new_n1164_, new_n1089_, new_n1153_ );
not g822 ( new_n1165_, new_n1164_ );
nand g823 ( new_n1166_, new_n1163_, new_n1165_ );
nor g824 ( new_n1167_, new_n1166_, keyIn_0_236 );
not g825 ( new_n1168_, new_n1167_ );
nand g826 ( new_n1169_, new_n1166_, keyIn_0_236 );
nand g827 ( new_n1170_, new_n1169_, N219 );
not g828 ( new_n1171_, new_n1170_ );
nand g829 ( new_n1172_, new_n1171_, new_n1168_ );
nand g830 ( new_n1173_, new_n661_, N210 );
xnor g831 ( new_n1174_, new_n1173_, keyIn_0_75 );
nand g832 ( new_n1175_, new_n1172_, new_n1174_ );
nand g833 ( new_n1176_, new_n1175_, new_n1148_ );
nor g834 ( new_n1177_, new_n1170_, new_n1167_ );
not g835 ( new_n1178_, new_n1174_ );
nor g836 ( new_n1179_, new_n1177_, new_n1178_ );
nand g837 ( new_n1180_, new_n1179_, keyIn_0_249 );
nand g838 ( new_n1181_, new_n1176_, new_n1180_ );
nor g839 ( new_n1182_, new_n1152_, new_n704_ );
xnor g840 ( new_n1183_, new_n1182_, keyIn_0_178 );
nand g841 ( new_n1184_, new_n1150_, N237 );
nand g842 ( new_n1185_, new_n1183_, new_n1184_ );
xor g843 ( new_n1186_, new_n1185_, keyIn_0_201 );
nand g844 ( new_n1187_, new_n1110_, N246 );
xor g845 ( new_n1188_, new_n1187_, keyIn_0_142 );
nand g846 ( new_n1189_, new_n734_, N159 );
xor g847 ( new_n1190_, new_n1189_, keyIn_0_117 );
nor g848 ( new_n1191_, new_n1188_, new_n1190_ );
not g849 ( new_n1192_, new_n1191_ );
nor g850 ( new_n1193_, new_n1186_, new_n1192_ );
nand g851 ( new_n1194_, new_n1181_, new_n1193_ );
nand g852 ( new_n1195_, new_n1194_, new_n1147_ );
xnor g853 ( new_n1196_, new_n1179_, new_n1148_ );
not g854 ( new_n1197_, new_n1193_ );
nor g855 ( new_n1198_, new_n1196_, new_n1197_ );
nand g856 ( new_n1199_, new_n1198_, keyIn_0_251 );
nand g857 ( new_n1200_, new_n1199_, new_n1195_ );
nand g858 ( new_n1201_, new_n1200_, keyIn_0_254 );
not g859 ( new_n1202_, keyIn_0_254 );
xnor g860 ( new_n1203_, new_n1194_, keyIn_0_251 );
nand g861 ( new_n1204_, new_n1203_, new_n1202_ );
nand g862 ( N878, new_n1204_, new_n1201_ );
nor g863 ( new_n1206_, new_n1065_, new_n1037_ );
nand g864 ( new_n1207_, new_n1206_, keyIn_0_224 );
nor g865 ( new_n1208_, new_n1206_, keyIn_0_224 );
nor g866 ( new_n1209_, new_n1071_, new_n1037_ );
xnor g867 ( new_n1210_, new_n1209_, keyIn_0_198 );
xor g868 ( new_n1211_, new_n1076_, keyIn_0_181 );
nand g869 ( new_n1212_, new_n1210_, new_n1211_ );
nor g870 ( new_n1213_, new_n1208_, new_n1212_ );
nand g871 ( new_n1214_, new_n1213_, new_n1207_ );
nor g872 ( new_n1215_, new_n1016_, new_n1083_ );
xor g873 ( new_n1216_, new_n1215_, keyIn_0_159 );
nor g874 ( new_n1217_, new_n1214_, new_n1216_ );
nand g875 ( new_n1218_, new_n1214_, new_n1216_ );
nand g876 ( new_n1219_, new_n1218_, N219 );
nor g877 ( new_n1220_, new_n1219_, new_n1217_ );
xnor g878 ( new_n1221_, new_n1220_, keyIn_0_242 );
not g879 ( new_n1222_, keyIn_0_32 );
nand g880 ( new_n1223_, N91, N210 );
nand g881 ( new_n1224_, new_n1223_, new_n1222_ );
not g882 ( new_n1225_, new_n1224_ );
nand g883 ( new_n1226_, keyIn_0_32, N91 );
nor g884 ( new_n1227_, new_n1226_, new_n865_ );
nor g885 ( new_n1228_, new_n1225_, new_n1227_ );
nor g886 ( new_n1229_, new_n1221_, new_n1228_ );
xnor g887 ( new_n1230_, new_n1229_, keyIn_0_250 );
not g888 ( new_n1231_, keyIn_0_180 );
nand g889 ( new_n1232_, new_n1216_, N228 );
nor g890 ( new_n1233_, new_n1232_, new_n1231_ );
nand g891 ( new_n1234_, new_n1083_, N237 );
nand g892 ( new_n1235_, new_n1232_, new_n1231_ );
nand g893 ( new_n1236_, new_n1235_, new_n1234_ );
nor g894 ( new_n1237_, new_n1236_, new_n1233_ );
xnor g895 ( new_n1238_, new_n1237_, keyIn_0_202 );
nand g896 ( new_n1239_, new_n1013_, N246 );
nand g897 ( new_n1240_, new_n734_, N165 );
xnor g898 ( new_n1241_, new_n1240_, keyIn_0_118 );
nand g899 ( new_n1242_, new_n1239_, new_n1241_ );
nor g900 ( new_n1243_, new_n1238_, new_n1242_ );
nand g901 ( new_n1244_, new_n1230_, new_n1243_ );
xor g902 ( N879, new_n1244_, keyIn_0_255 );
not g903 ( new_n1246_, new_n1037_ );
nand g904 ( new_n1247_, new_n1246_, new_n1077_ );
xnor g905 ( new_n1248_, new_n1247_, keyIn_0_160 );
not g906 ( new_n1249_, new_n1248_ );
xnor g907 ( new_n1250_, new_n1070_, keyIn_0_183 );
nand g908 ( new_n1251_, new_n1065_, new_n1250_ );
nor g909 ( new_n1252_, new_n1251_, new_n1249_ );
xnor g910 ( new_n1253_, new_n1252_, keyIn_0_231 );
nand g911 ( new_n1254_, new_n1251_, new_n1249_ );
xnor g912 ( new_n1255_, new_n1254_, keyIn_0_232 );
nor g913 ( new_n1256_, new_n1253_, new_n1255_ );
nand g914 ( new_n1257_, new_n1256_, keyIn_0_237 );
not g915 ( new_n1258_, N219 );
nor g916 ( new_n1259_, new_n1256_, keyIn_0_237 );
nor g917 ( new_n1260_, new_n1259_, new_n1258_ );
nand g918 ( new_n1261_, new_n1260_, new_n1257_ );
nor g919 ( new_n1262_, new_n1261_, keyIn_0_243 );
nand g920 ( new_n1263_, new_n1261_, keyIn_0_243 );
not g921 ( new_n1264_, keyIn_0_203 );
nor g922 ( new_n1265_, new_n1248_, new_n704_ );
nand g923 ( new_n1266_, new_n1076_, N237 );
xnor g924 ( new_n1267_, new_n1266_, keyIn_0_182 );
not g925 ( new_n1268_, new_n1267_ );
nor g926 ( new_n1269_, new_n1265_, new_n1268_ );
not g927 ( new_n1270_, new_n1269_ );
nor g928 ( new_n1271_, new_n1270_, new_n1264_ );
nand g929 ( new_n1272_, new_n1270_, new_n1264_ );
not g930 ( new_n1273_, keyIn_0_161 );
nand g931 ( new_n1274_, new_n1034_, N246 );
nand g932 ( new_n1275_, new_n734_, N171 );
xnor g933 ( new_n1276_, new_n1275_, keyIn_0_119 );
nand g934 ( new_n1277_, new_n1274_, new_n1276_ );
nor g935 ( new_n1278_, new_n1277_, new_n1273_ );
nand g936 ( new_n1279_, new_n1277_, new_n1273_ );
nand g937 ( new_n1280_, N96, N210 );
xor g938 ( new_n1281_, new_n1280_, keyIn_0_33 );
nand g939 ( new_n1282_, new_n1279_, new_n1281_ );
nor g940 ( new_n1283_, new_n1282_, new_n1278_ );
nand g941 ( new_n1284_, new_n1272_, new_n1283_ );
nor g942 ( new_n1285_, new_n1284_, new_n1271_ );
nand g943 ( new_n1286_, new_n1263_, new_n1285_ );
nor g944 ( new_n1287_, new_n1286_, new_n1262_ );
xor g945 ( N880, new_n1287_, keyIn_0_252 );
endmodule