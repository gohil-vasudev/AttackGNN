module locked_c2670 (  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,  G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225  );
  input  G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire new_n359_, new_n368_, new_n369_, new_n370_, new_n371_, new_n373_, new_n374_, new_n376_, new_n378_, new_n380_, new_n381_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n396_, new_n397_, new_n398_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n500_, new_n501_, new_n503_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_, new_n977_, new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n990_, new_n991_;
  XOR2_X1 g000 ( .A(G44), .B(KEYINPUT3), .Z(new_n359_) );
  INV_X1 g001 ( .A(new_n359_), .ZN(G218) );
  INV_X1 g002 ( .A(G132), .ZN(G219) );
  INV_X1 g003 ( .A(G82), .ZN(G220) );
  INV_X1 g004 ( .A(G96), .ZN(G221) );
  INV_X1 g005 ( .A(G69), .ZN(G235) );
  INV_X1 g006 ( .A(G120), .ZN(G236) );
  INV_X1 g007 ( .A(G57), .ZN(G237) );
  INV_X1 g008 ( .A(G108), .ZN(G238) );
  NAND2_X1 g009 ( .A1(G2078), .A2(G2084), .ZN(new_n368_) );
  XOR2_X1 g010 ( .A(new_n368_), .B(KEYINPUT20), .Z(new_n369_) );
  NAND2_X1 g011 ( .A1(new_n369_), .A2(G2090), .ZN(new_n370_) );
  XNOR2_X1 g012 ( .A(new_n370_), .B(KEYINPUT21), .ZN(new_n371_) );
  NAND2_X1 g013 ( .A1(new_n371_), .A2(G2072), .ZN(G158) );
  NAND2_X1 g014 ( .A1(G2), .A2(G15), .ZN(new_n373_) );
  INV_X1 g015 ( .A(new_n373_), .ZN(new_n374_) );
  NAND2_X1 g016 ( .A1(new_n374_), .A2(G661), .ZN(G259) );
  NAND2_X1 g017 ( .A1(G94), .A2(G452), .ZN(new_n376_) );
  INV_X1 g018 ( .A(new_n376_), .ZN(G173) );
  NAND2_X1 g019 ( .A1(G7), .A2(G661), .ZN(new_n378_) );
  XNOR2_X1 g020 ( .A(new_n378_), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 g021 ( .A(G223), .ZN(new_n380_) );
  NAND2_X1 g022 ( .A1(new_n380_), .A2(G567), .ZN(new_n381_) );
  XOR2_X1 g023 ( .A(new_n381_), .B(KEYINPUT11), .Z(G234) );
  NAND2_X1 g024 ( .A1(new_n380_), .A2(G2106), .ZN(G217) );
  NAND2_X1 g025 ( .A1(G82), .A2(G132), .ZN(new_n384_) );
  XNOR2_X1 g026 ( .A(new_n384_), .B(KEYINPUT22), .ZN(new_n385_) );
  NOR2_X1 g027 ( .A1(G218), .A2(G221), .ZN(new_n386_) );
  INV_X1 g028 ( .A(new_n386_), .ZN(new_n387_) );
  NOR2_X1 g029 ( .A1(new_n387_), .A2(new_n385_), .ZN(new_n388_) );
  INV_X1 g030 ( .A(new_n388_), .ZN(new_n389_) );
  NAND2_X1 g031 ( .A1(G57), .A2(G69), .ZN(new_n390_) );
  NAND2_X1 g032 ( .A1(G108), .A2(G120), .ZN(new_n391_) );
  NOR2_X1 g033 ( .A1(new_n390_), .A2(new_n391_), .ZN(new_n392_) );
  INV_X1 g034 ( .A(new_n392_), .ZN(new_n393_) );
  NOR2_X1 g035 ( .A1(new_n389_), .A2(new_n393_), .ZN(G325) );
  INV_X1 g036 ( .A(G325), .ZN(G261) );
  NAND2_X1 g037 ( .A1(new_n389_), .A2(G2106), .ZN(new_n396_) );
  NAND2_X1 g038 ( .A1(new_n393_), .A2(G567), .ZN(new_n397_) );
  NAND2_X1 g039 ( .A1(new_n396_), .A2(new_n397_), .ZN(new_n398_) );
  INV_X1 g040 ( .A(new_n398_), .ZN(G319) );
  NAND2_X1 g041 ( .A1(G101), .A2(G2104), .ZN(new_n400_) );
  NOR2_X1 g042 ( .A1(new_n400_), .A2(G2105), .ZN(new_n401_) );
  XOR2_X1 g043 ( .A(new_n401_), .B(KEYINPUT23), .Z(new_n402_) );
  INV_X1 g044 ( .A(G2105), .ZN(new_n403_) );
  INV_X1 g045 ( .A(G2104), .ZN(new_n404_) );
  NAND2_X1 g046 ( .A1(new_n404_), .A2(G125), .ZN(new_n405_) );
  NOR2_X1 g047 ( .A1(new_n405_), .A2(new_n403_), .ZN(new_n406_) );
  INV_X1 g048 ( .A(G113), .ZN(new_n407_) );
  NAND2_X1 g049 ( .A1(G2104), .A2(G2105), .ZN(new_n408_) );
  NOR2_X1 g050 ( .A1(new_n408_), .A2(new_n407_), .ZN(new_n409_) );
  NOR2_X1 g051 ( .A1(new_n406_), .A2(new_n409_), .ZN(new_n410_) );
  NAND2_X1 g052 ( .A1(new_n404_), .A2(new_n403_), .ZN(new_n411_) );
  NAND2_X1 g053 ( .A1(new_n411_), .A2(KEYINPUT17), .ZN(new_n412_) );
  INV_X1 g054 ( .A(KEYINPUT17), .ZN(new_n413_) );
  NOR2_X1 g055 ( .A1(G2104), .A2(G2105), .ZN(new_n414_) );
  NAND2_X1 g056 ( .A1(new_n414_), .A2(new_n413_), .ZN(new_n415_) );
  NAND2_X1 g057 ( .A1(new_n412_), .A2(new_n415_), .ZN(new_n416_) );
  NAND2_X1 g058 ( .A1(new_n416_), .A2(G137), .ZN(new_n417_) );
  NAND2_X1 g059 ( .A1(new_n417_), .A2(new_n410_), .ZN(new_n418_) );
  NOR2_X1 g060 ( .A1(new_n418_), .A2(new_n402_), .ZN(G160) );
  INV_X1 g061 ( .A(G136), .ZN(new_n420_) );
  XNOR2_X1 g062 ( .A(new_n414_), .B(KEYINPUT17), .ZN(new_n421_) );
  NOR2_X1 g063 ( .A1(new_n421_), .A2(new_n420_), .ZN(new_n422_) );
  NOR2_X1 g064 ( .A1(new_n403_), .A2(G2104), .ZN(new_n423_) );
  NAND2_X1 g065 ( .A1(new_n423_), .A2(G124), .ZN(new_n424_) );
  XNOR2_X1 g066 ( .A(new_n424_), .B(KEYINPUT44), .ZN(new_n425_) );
  INV_X1 g067 ( .A(G100), .ZN(new_n426_) );
  NOR2_X1 g068 ( .A1(new_n404_), .A2(G2105), .ZN(new_n427_) );
  INV_X1 g069 ( .A(new_n427_), .ZN(new_n428_) );
  NOR2_X1 g070 ( .A1(new_n428_), .A2(new_n426_), .ZN(new_n429_) );
  INV_X1 g071 ( .A(G112), .ZN(new_n430_) );
  NOR2_X1 g072 ( .A1(new_n408_), .A2(new_n430_), .ZN(new_n431_) );
  NOR2_X1 g073 ( .A1(new_n429_), .A2(new_n431_), .ZN(new_n432_) );
  NAND2_X1 g074 ( .A1(new_n425_), .A2(new_n432_), .ZN(new_n433_) );
  NOR2_X1 g075 ( .A1(new_n433_), .A2(new_n422_), .ZN(G162) );
  NAND2_X1 g076 ( .A1(new_n416_), .A2(G138), .ZN(new_n435_) );
  INV_X1 g077 ( .A(G114), .ZN(new_n436_) );
  NOR2_X1 g078 ( .A1(new_n408_), .A2(new_n436_), .ZN(new_n437_) );
  NAND2_X1 g079 ( .A1(G102), .A2(G2104), .ZN(new_n438_) );
  NOR2_X1 g080 ( .A1(new_n438_), .A2(G2105), .ZN(new_n439_) );
  INV_X1 g081 ( .A(new_n439_), .ZN(new_n440_) );
  NAND2_X1 g082 ( .A1(new_n423_), .A2(G126), .ZN(new_n441_) );
  NAND2_X1 g083 ( .A1(new_n440_), .A2(new_n441_), .ZN(new_n442_) );
  NOR2_X1 g084 ( .A1(new_n442_), .A2(new_n437_), .ZN(new_n443_) );
  NAND2_X1 g085 ( .A1(new_n443_), .A2(new_n435_), .ZN(new_n444_) );
  INV_X1 g086 ( .A(new_n444_), .ZN(G164) );
  NOR2_X1 g087 ( .A1(G543), .A2(G651), .ZN(new_n446_) );
  NAND2_X1 g088 ( .A1(new_n446_), .A2(G88), .ZN(new_n447_) );
  INV_X1 g089 ( .A(G543), .ZN(new_n448_) );
  NAND2_X1 g090 ( .A1(new_n448_), .A2(G651), .ZN(new_n449_) );
  XNOR2_X1 g091 ( .A(new_n449_), .B(KEYINPUT1), .ZN(new_n450_) );
  NAND2_X1 g092 ( .A1(new_n450_), .A2(G62), .ZN(new_n451_) );
  NAND2_X1 g093 ( .A1(new_n451_), .A2(new_n447_), .ZN(new_n452_) );
  XOR2_X1 g094 ( .A(G543), .B(KEYINPUT0), .Z(new_n453_) );
  NOR2_X1 g095 ( .A1(new_n453_), .A2(G651), .ZN(new_n454_) );
  NAND2_X1 g096 ( .A1(new_n454_), .A2(G50), .ZN(new_n455_) );
  INV_X1 g097 ( .A(G651), .ZN(new_n456_) );
  NOR2_X1 g098 ( .A1(new_n453_), .A2(new_n456_), .ZN(new_n457_) );
  NAND2_X1 g099 ( .A1(new_n457_), .A2(G75), .ZN(new_n458_) );
  NAND2_X1 g100 ( .A1(new_n455_), .A2(new_n458_), .ZN(new_n459_) );
  NOR2_X1 g101 ( .A1(new_n459_), .A2(new_n452_), .ZN(G166) );
  NAND2_X1 g102 ( .A1(new_n454_), .A2(G51), .ZN(new_n461_) );
  NAND2_X1 g103 ( .A1(new_n450_), .A2(G63), .ZN(new_n462_) );
  NAND2_X1 g104 ( .A1(new_n461_), .A2(new_n462_), .ZN(new_n463_) );
  XOR2_X1 g105 ( .A(new_n463_), .B(KEYINPUT6), .Z(new_n464_) );
  NAND2_X1 g106 ( .A1(new_n446_), .A2(G89), .ZN(new_n465_) );
  XNOR2_X1 g107 ( .A(new_n465_), .B(KEYINPUT4), .ZN(new_n466_) );
  NAND2_X1 g108 ( .A1(new_n457_), .A2(G76), .ZN(new_n467_) );
  NAND2_X1 g109 ( .A1(new_n467_), .A2(new_n466_), .ZN(new_n468_) );
  XNOR2_X1 g110 ( .A(new_n468_), .B(KEYINPUT5), .ZN(new_n469_) );
  NAND2_X1 g111 ( .A1(new_n464_), .A2(new_n469_), .ZN(new_n470_) );
  XNOR2_X1 g112 ( .A(new_n470_), .B(KEYINPUT7), .ZN(G168) );
  INV_X1 g113 ( .A(KEYINPUT9), .ZN(new_n472_) );
  NAND2_X1 g114 ( .A1(new_n457_), .A2(G77), .ZN(new_n473_) );
  NAND2_X1 g115 ( .A1(new_n446_), .A2(G90), .ZN(new_n474_) );
  NAND2_X1 g116 ( .A1(new_n473_), .A2(new_n474_), .ZN(new_n475_) );
  NOR2_X1 g117 ( .A1(new_n475_), .A2(new_n472_), .ZN(new_n476_) );
  NAND2_X1 g118 ( .A1(new_n475_), .A2(new_n472_), .ZN(new_n477_) );
  INV_X1 g119 ( .A(new_n477_), .ZN(new_n478_) );
  NAND2_X1 g120 ( .A1(new_n454_), .A2(G52), .ZN(new_n479_) );
  NAND2_X1 g121 ( .A1(new_n450_), .A2(G64), .ZN(new_n480_) );
  NAND2_X1 g122 ( .A1(new_n479_), .A2(new_n480_), .ZN(new_n481_) );
  NOR2_X1 g123 ( .A1(new_n478_), .A2(new_n481_), .ZN(new_n482_) );
  INV_X1 g124 ( .A(new_n482_), .ZN(new_n483_) );
  NOR2_X1 g125 ( .A1(new_n483_), .A2(new_n476_), .ZN(G171) );
  NAND2_X1 g126 ( .A1(new_n446_), .A2(G81), .ZN(new_n485_) );
  XNOR2_X1 g127 ( .A(new_n485_), .B(KEYINPUT12), .ZN(new_n486_) );
  NAND2_X1 g128 ( .A1(new_n457_), .A2(G68), .ZN(new_n487_) );
  NAND2_X1 g129 ( .A1(new_n487_), .A2(new_n486_), .ZN(new_n488_) );
  XOR2_X1 g130 ( .A(new_n488_), .B(KEYINPUT13), .Z(new_n489_) );
  INV_X1 g131 ( .A(KEYINPUT14), .ZN(new_n490_) );
  NAND2_X1 g132 ( .A1(new_n450_), .A2(G56), .ZN(new_n491_) );
  NOR2_X1 g133 ( .A1(new_n491_), .A2(new_n490_), .ZN(new_n492_) );
  NAND2_X1 g134 ( .A1(new_n454_), .A2(G43), .ZN(new_n493_) );
  NAND2_X1 g135 ( .A1(new_n491_), .A2(new_n490_), .ZN(new_n494_) );
  NAND2_X1 g136 ( .A1(new_n494_), .A2(new_n493_), .ZN(new_n495_) );
  NOR2_X1 g137 ( .A1(new_n495_), .A2(new_n492_), .ZN(new_n496_) );
  INV_X1 g138 ( .A(new_n496_), .ZN(new_n497_) );
  NOR2_X1 g139 ( .A1(new_n489_), .A2(new_n497_), .ZN(new_n498_) );
  NAND2_X1 g140 ( .A1(new_n498_), .A2(G860), .ZN(G153) );
  NAND2_X1 g141 ( .A1(G483), .A2(G661), .ZN(new_n500_) );
  NOR2_X1 g142 ( .A1(new_n398_), .A2(new_n500_), .ZN(new_n501_) );
  NAND2_X1 g143 ( .A1(new_n501_), .A2(G36), .ZN(G176) );
  NAND2_X1 g144 ( .A1(G1), .A2(G3), .ZN(new_n503_) );
  NAND2_X1 g145 ( .A1(new_n501_), .A2(new_n503_), .ZN(G188) );
  NAND2_X1 g146 ( .A1(new_n446_), .A2(G91), .ZN(new_n505_) );
  NAND2_X1 g147 ( .A1(new_n450_), .A2(G65), .ZN(new_n506_) );
  NAND2_X1 g148 ( .A1(new_n506_), .A2(new_n505_), .ZN(new_n507_) );
  NAND2_X1 g149 ( .A1(new_n454_), .A2(G53), .ZN(new_n508_) );
  NAND2_X1 g150 ( .A1(new_n457_), .A2(G78), .ZN(new_n509_) );
  NAND2_X1 g151 ( .A1(new_n508_), .A2(new_n509_), .ZN(new_n510_) );
  NOR2_X1 g152 ( .A1(new_n510_), .A2(new_n507_), .ZN(new_n511_) );
  INV_X1 g153 ( .A(new_n511_), .ZN(G299) );
  INV_X1 g154 ( .A(G171), .ZN(G301) );
  XOR2_X1 g155 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 g156 ( .A(G166), .ZN(G303) );
  NAND2_X1 g157 ( .A1(new_n454_), .A2(G49), .ZN(new_n516_) );
  NAND2_X1 g158 ( .A1(new_n453_), .A2(G87), .ZN(new_n517_) );
  INV_X1 g159 ( .A(new_n517_), .ZN(new_n518_) );
  INV_X1 g160 ( .A(new_n450_), .ZN(new_n519_) );
  NAND2_X1 g161 ( .A1(G74), .A2(G651), .ZN(new_n520_) );
  NAND2_X1 g162 ( .A1(new_n519_), .A2(new_n520_), .ZN(new_n521_) );
  NOR2_X1 g163 ( .A1(new_n521_), .A2(new_n518_), .ZN(new_n522_) );
  NAND2_X1 g164 ( .A1(new_n522_), .A2(new_n516_), .ZN(G288) );
  NAND2_X1 g165 ( .A1(new_n457_), .A2(G73), .ZN(new_n524_) );
  XNOR2_X1 g166 ( .A(new_n524_), .B(KEYINPUT2), .ZN(new_n525_) );
  INV_X1 g167 ( .A(G61), .ZN(new_n526_) );
  NOR2_X1 g168 ( .A1(new_n519_), .A2(new_n526_), .ZN(new_n527_) );
  NAND2_X1 g169 ( .A1(new_n446_), .A2(G86), .ZN(new_n528_) );
  NAND2_X1 g170 ( .A1(new_n454_), .A2(G48), .ZN(new_n529_) );
  NAND2_X1 g171 ( .A1(new_n529_), .A2(new_n528_), .ZN(new_n530_) );
  NOR2_X1 g172 ( .A1(new_n530_), .A2(new_n527_), .ZN(new_n531_) );
  NAND2_X1 g173 ( .A1(new_n525_), .A2(new_n531_), .ZN(G305) );
  NAND2_X1 g174 ( .A1(new_n446_), .A2(G85), .ZN(new_n533_) );
  NAND2_X1 g175 ( .A1(new_n450_), .A2(G60), .ZN(new_n534_) );
  NAND2_X1 g176 ( .A1(new_n534_), .A2(new_n533_), .ZN(new_n535_) );
  NAND2_X1 g177 ( .A1(new_n454_), .A2(G47), .ZN(new_n536_) );
  NAND2_X1 g178 ( .A1(new_n457_), .A2(G72), .ZN(new_n537_) );
  NAND2_X1 g179 ( .A1(new_n536_), .A2(new_n537_), .ZN(new_n538_) );
  NOR2_X1 g180 ( .A1(new_n538_), .A2(new_n535_), .ZN(new_n539_) );
  INV_X1 g181 ( .A(new_n539_), .ZN(G290) );
  INV_X1 g182 ( .A(G868), .ZN(new_n541_) );
  NAND2_X1 g183 ( .A1(new_n446_), .A2(G92), .ZN(new_n542_) );
  NAND2_X1 g184 ( .A1(new_n450_), .A2(G66), .ZN(new_n543_) );
  NAND2_X1 g185 ( .A1(new_n543_), .A2(new_n542_), .ZN(new_n544_) );
  NAND2_X1 g186 ( .A1(new_n457_), .A2(G79), .ZN(new_n545_) );
  NAND2_X1 g187 ( .A1(new_n454_), .A2(G54), .ZN(new_n546_) );
  NAND2_X1 g188 ( .A1(new_n545_), .A2(new_n546_), .ZN(new_n547_) );
  NOR2_X1 g189 ( .A1(new_n547_), .A2(new_n544_), .ZN(new_n548_) );
  XNOR2_X1 g190 ( .A(new_n548_), .B(KEYINPUT15), .ZN(new_n549_) );
  NAND2_X1 g191 ( .A1(new_n549_), .A2(new_n541_), .ZN(new_n550_) );
  NAND2_X1 g192 ( .A1(G301), .A2(G868), .ZN(new_n551_) );
  NAND2_X1 g193 ( .A1(new_n551_), .A2(new_n550_), .ZN(G284) );
  INV_X1 g194 ( .A(G286), .ZN(new_n553_) );
  NAND2_X1 g195 ( .A1(new_n553_), .A2(G868), .ZN(new_n554_) );
  NAND2_X1 g196 ( .A1(new_n511_), .A2(new_n541_), .ZN(new_n555_) );
  NAND2_X1 g197 ( .A1(new_n554_), .A2(new_n555_), .ZN(new_n556_) );
  INV_X1 g198 ( .A(new_n556_), .ZN(G297) );
  INV_X1 g199 ( .A(new_n549_), .ZN(new_n558_) );
  INV_X1 g200 ( .A(G860), .ZN(new_n559_) );
  NAND2_X1 g201 ( .A1(new_n559_), .A2(G559), .ZN(new_n560_) );
  NAND2_X1 g202 ( .A1(new_n558_), .A2(new_n560_), .ZN(new_n561_) );
  XNOR2_X1 g203 ( .A(new_n561_), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 g204 ( .A(new_n498_), .ZN(new_n563_) );
  NOR2_X1 g205 ( .A1(new_n563_), .A2(G868), .ZN(new_n564_) );
  INV_X1 g206 ( .A(G559), .ZN(new_n565_) );
  NAND2_X1 g207 ( .A1(new_n565_), .A2(G868), .ZN(new_n566_) );
  NOR2_X1 g208 ( .A1(new_n549_), .A2(new_n566_), .ZN(new_n567_) );
  NOR2_X1 g209 ( .A1(new_n564_), .A2(new_n567_), .ZN(G282) );
  INV_X1 g210 ( .A(G2100), .ZN(new_n569_) );
  INV_X1 g211 ( .A(G135), .ZN(new_n570_) );
  NOR2_X1 g212 ( .A1(new_n421_), .A2(new_n570_), .ZN(new_n571_) );
  NAND2_X1 g213 ( .A1(new_n423_), .A2(G123), .ZN(new_n572_) );
  XNOR2_X1 g214 ( .A(new_n572_), .B(KEYINPUT18), .ZN(new_n573_) );
  INV_X1 g215 ( .A(G111), .ZN(new_n574_) );
  NOR2_X1 g216 ( .A1(new_n408_), .A2(new_n574_), .ZN(new_n575_) );
  INV_X1 g217 ( .A(G99), .ZN(new_n576_) );
  NOR2_X1 g218 ( .A1(new_n428_), .A2(new_n576_), .ZN(new_n577_) );
  NOR2_X1 g219 ( .A1(new_n577_), .A2(new_n575_), .ZN(new_n578_) );
  NAND2_X1 g220 ( .A1(new_n573_), .A2(new_n578_), .ZN(new_n579_) );
  NOR2_X1 g221 ( .A1(new_n579_), .A2(new_n571_), .ZN(new_n580_) );
  XNOR2_X1 g222 ( .A(new_n580_), .B(G2096), .ZN(new_n581_) );
  NAND2_X1 g223 ( .A1(new_n581_), .A2(new_n569_), .ZN(G156) );
  INV_X1 g224 ( .A(G14), .ZN(new_n583_) );
  XOR2_X1 g225 ( .A(G2430), .B(G2454), .Z(new_n584_) );
  XNOR2_X1 g226 ( .A(G1341), .B(G1348), .ZN(new_n585_) );
  XNOR2_X1 g227 ( .A(new_n584_), .B(new_n585_), .ZN(new_n586_) );
  XOR2_X1 g228 ( .A(G2435), .B(G2438), .Z(new_n587_) );
  XNOR2_X1 g229 ( .A(new_n586_), .B(new_n587_), .ZN(new_n588_) );
  XOR2_X1 g230 ( .A(G2446), .B(G2451), .Z(new_n589_) );
  XNOR2_X1 g231 ( .A(G2427), .B(G2443), .ZN(new_n590_) );
  XNOR2_X1 g232 ( .A(new_n589_), .B(new_n590_), .ZN(new_n591_) );
  XNOR2_X1 g233 ( .A(new_n588_), .B(new_n591_), .ZN(new_n592_) );
  NOR2_X1 g234 ( .A1(new_n592_), .A2(new_n583_), .ZN(G401) );
  XOR2_X1 g235 ( .A(G2090), .B(KEYINPUT42), .Z(new_n594_) );
  XNOR2_X1 g236 ( .A(G2067), .B(G2072), .ZN(new_n595_) );
  XNOR2_X1 g237 ( .A(new_n594_), .B(new_n595_), .ZN(new_n596_) );
  XNOR2_X1 g238 ( .A(G2096), .B(G2100), .ZN(new_n597_) );
  XNOR2_X1 g239 ( .A(G2678), .B(KEYINPUT43), .ZN(new_n598_) );
  XNOR2_X1 g240 ( .A(new_n597_), .B(new_n598_), .ZN(new_n599_) );
  XNOR2_X1 g241 ( .A(new_n596_), .B(new_n599_), .ZN(new_n600_) );
  XNOR2_X1 g242 ( .A(G2078), .B(G2084), .ZN(new_n601_) );
  XNOR2_X1 g243 ( .A(new_n600_), .B(new_n601_), .ZN(G227) );
  XOR2_X1 g244 ( .A(G1976), .B(G1981), .Z(new_n603_) );
  XNOR2_X1 g245 ( .A(G1956), .B(G1966), .ZN(new_n604_) );
  XNOR2_X1 g246 ( .A(new_n603_), .B(new_n604_), .ZN(new_n605_) );
  XNOR2_X1 g247 ( .A(new_n605_), .B(G2474), .ZN(new_n606_) );
  XNOR2_X1 g248 ( .A(G1991), .B(G1996), .ZN(new_n607_) );
  XNOR2_X1 g249 ( .A(new_n606_), .B(new_n607_), .ZN(new_n608_) );
  XOR2_X1 g250 ( .A(G1971), .B(KEYINPUT41), .Z(new_n609_) );
  XNOR2_X1 g251 ( .A(G1961), .B(G1986), .ZN(new_n610_) );
  XNOR2_X1 g252 ( .A(new_n609_), .B(new_n610_), .ZN(new_n611_) );
  XNOR2_X1 g253 ( .A(new_n608_), .B(new_n611_), .ZN(new_n612_) );
  INV_X1 g254 ( .A(new_n612_), .ZN(G229) );
  INV_X1 g255 ( .A(KEYINPUT55), .ZN(new_n614_) );
  INV_X1 g256 ( .A(KEYINPUT50), .ZN(new_n615_) );
  INV_X1 g257 ( .A(KEYINPUT47), .ZN(new_n616_) );
  NAND2_X1 g258 ( .A1(new_n423_), .A2(G127), .ZN(new_n617_) );
  INV_X1 g259 ( .A(new_n408_), .ZN(new_n618_) );
  NAND2_X1 g260 ( .A1(new_n618_), .A2(G115), .ZN(new_n619_) );
  NAND2_X1 g261 ( .A1(new_n617_), .A2(new_n619_), .ZN(new_n620_) );
  NOR2_X1 g262 ( .A1(new_n620_), .A2(new_n616_), .ZN(new_n621_) );
  NAND2_X1 g263 ( .A1(new_n427_), .A2(G103), .ZN(new_n622_) );
  INV_X1 g264 ( .A(new_n622_), .ZN(new_n623_) );
  NOR2_X1 g265 ( .A1(new_n621_), .A2(new_n623_), .ZN(new_n624_) );
  INV_X1 g266 ( .A(new_n624_), .ZN(new_n625_) );
  NAND2_X1 g267 ( .A1(new_n620_), .A2(new_n616_), .ZN(new_n626_) );
  NAND2_X1 g268 ( .A1(new_n416_), .A2(G139), .ZN(new_n627_) );
  NAND2_X1 g269 ( .A1(new_n626_), .A2(new_n627_), .ZN(new_n628_) );
  NOR2_X1 g270 ( .A1(new_n625_), .A2(new_n628_), .ZN(new_n629_) );
  INV_X1 g271 ( .A(new_n629_), .ZN(new_n630_) );
  NOR2_X1 g272 ( .A1(new_n630_), .A2(G2072), .ZN(new_n631_) );
  NAND2_X1 g273 ( .A1(new_n630_), .A2(G2072), .ZN(new_n632_) );
  INV_X1 g274 ( .A(new_n632_), .ZN(new_n633_) );
  XNOR2_X1 g275 ( .A(new_n444_), .B(G2078), .ZN(new_n634_) );
  NOR2_X1 g276 ( .A1(new_n633_), .A2(new_n634_), .ZN(new_n635_) );
  INV_X1 g277 ( .A(new_n635_), .ZN(new_n636_) );
  NOR2_X1 g278 ( .A1(new_n636_), .A2(new_n631_), .ZN(new_n637_) );
  NAND2_X1 g279 ( .A1(new_n637_), .A2(new_n615_), .ZN(new_n638_) );
  INV_X1 g280 ( .A(G1996), .ZN(new_n639_) );
  NAND2_X1 g281 ( .A1(new_n416_), .A2(G141), .ZN(new_n640_) );
  INV_X1 g282 ( .A(KEYINPUT38), .ZN(new_n641_) );
  NAND2_X1 g283 ( .A1(new_n427_), .A2(G105), .ZN(new_n642_) );
  NOR2_X1 g284 ( .A1(new_n642_), .A2(new_n641_), .ZN(new_n643_) );
  NAND2_X1 g285 ( .A1(new_n642_), .A2(new_n641_), .ZN(new_n644_) );
  INV_X1 g286 ( .A(new_n644_), .ZN(new_n645_) );
  NAND2_X1 g287 ( .A1(new_n618_), .A2(G117), .ZN(new_n646_) );
  NAND2_X1 g288 ( .A1(new_n423_), .A2(G129), .ZN(new_n647_) );
  NAND2_X1 g289 ( .A1(new_n647_), .A2(new_n646_), .ZN(new_n648_) );
  NOR2_X1 g290 ( .A1(new_n645_), .A2(new_n648_), .ZN(new_n649_) );
  INV_X1 g291 ( .A(new_n649_), .ZN(new_n650_) );
  NOR2_X1 g292 ( .A1(new_n650_), .A2(new_n643_), .ZN(new_n651_) );
  NAND2_X1 g293 ( .A1(new_n651_), .A2(new_n640_), .ZN(new_n652_) );
  INV_X1 g294 ( .A(new_n652_), .ZN(new_n653_) );
  NAND2_X1 g295 ( .A1(new_n653_), .A2(new_n639_), .ZN(new_n654_) );
  XNOR2_X1 g296 ( .A(G162), .B(G2090), .ZN(new_n655_) );
  NAND2_X1 g297 ( .A1(new_n654_), .A2(new_n655_), .ZN(new_n656_) );
  XNOR2_X1 g298 ( .A(new_n656_), .B(KEYINPUT51), .ZN(new_n657_) );
  NAND2_X1 g299 ( .A1(new_n638_), .A2(new_n657_), .ZN(new_n658_) );
  NAND2_X1 g300 ( .A1(new_n416_), .A2(G140), .ZN(new_n659_) );
  NAND2_X1 g301 ( .A1(new_n427_), .A2(G104), .ZN(new_n660_) );
  NAND2_X1 g302 ( .A1(new_n659_), .A2(new_n660_), .ZN(new_n661_) );
  NOR2_X1 g303 ( .A1(new_n661_), .A2(KEYINPUT34), .ZN(new_n662_) );
  NAND2_X1 g304 ( .A1(new_n661_), .A2(KEYINPUT34), .ZN(new_n663_) );
  NAND2_X1 g305 ( .A1(new_n423_), .A2(G128), .ZN(new_n664_) );
  NAND2_X1 g306 ( .A1(new_n618_), .A2(G116), .ZN(new_n665_) );
  NAND2_X1 g307 ( .A1(new_n664_), .A2(new_n665_), .ZN(new_n666_) );
  XNOR2_X1 g308 ( .A(new_n666_), .B(KEYINPUT35), .ZN(new_n667_) );
  NAND2_X1 g309 ( .A1(new_n663_), .A2(new_n667_), .ZN(new_n668_) );
  NOR2_X1 g310 ( .A1(new_n668_), .A2(new_n662_), .ZN(new_n669_) );
  XOR2_X1 g311 ( .A(new_n669_), .B(KEYINPUT36), .Z(new_n670_) );
  INV_X1 g312 ( .A(new_n670_), .ZN(new_n671_) );
  XNOR2_X1 g313 ( .A(G2067), .B(KEYINPUT37), .ZN(new_n672_) );
  NAND2_X1 g314 ( .A1(new_n671_), .A2(new_n672_), .ZN(new_n673_) );
  NOR2_X1 g315 ( .A1(new_n671_), .A2(new_n672_), .ZN(new_n674_) );
  INV_X1 g316 ( .A(new_n637_), .ZN(new_n675_) );
  NAND2_X1 g317 ( .A1(new_n675_), .A2(KEYINPUT50), .ZN(new_n676_) );
  NAND2_X1 g318 ( .A1(new_n416_), .A2(G131), .ZN(new_n677_) );
  NAND2_X1 g319 ( .A1(new_n423_), .A2(G119), .ZN(new_n678_) );
  INV_X1 g320 ( .A(new_n678_), .ZN(new_n679_) );
  NAND2_X1 g321 ( .A1(new_n618_), .A2(G107), .ZN(new_n680_) );
  NAND2_X1 g322 ( .A1(new_n427_), .A2(G95), .ZN(new_n681_) );
  NAND2_X1 g323 ( .A1(new_n681_), .A2(new_n680_), .ZN(new_n682_) );
  NOR2_X1 g324 ( .A1(new_n682_), .A2(new_n679_), .ZN(new_n683_) );
  NAND2_X1 g325 ( .A1(new_n683_), .A2(new_n677_), .ZN(new_n684_) );
  NAND2_X1 g326 ( .A1(new_n684_), .A2(G1991), .ZN(new_n685_) );
  NAND2_X1 g327 ( .A1(new_n652_), .A2(G1996), .ZN(new_n686_) );
  NAND2_X1 g328 ( .A1(new_n686_), .A2(new_n685_), .ZN(new_n687_) );
  XNOR2_X1 g329 ( .A(G160), .B(G2084), .ZN(new_n688_) );
  NOR2_X1 g330 ( .A1(new_n684_), .A2(G1991), .ZN(new_n689_) );
  NOR2_X1 g331 ( .A1(new_n580_), .A2(new_n689_), .ZN(new_n690_) );
  NAND2_X1 g332 ( .A1(new_n688_), .A2(new_n690_), .ZN(new_n691_) );
  NOR2_X1 g333 ( .A1(new_n687_), .A2(new_n691_), .ZN(new_n692_) );
  NAND2_X1 g334 ( .A1(new_n676_), .A2(new_n692_), .ZN(new_n693_) );
  NOR2_X1 g335 ( .A1(new_n693_), .A2(new_n674_), .ZN(new_n694_) );
  NAND2_X1 g336 ( .A1(new_n694_), .A2(new_n673_), .ZN(new_n695_) );
  NOR2_X1 g337 ( .A1(new_n695_), .A2(new_n658_), .ZN(new_n696_) );
  XNOR2_X1 g338 ( .A(new_n696_), .B(KEYINPUT52), .ZN(new_n697_) );
  NAND2_X1 g339 ( .A1(new_n697_), .A2(new_n614_), .ZN(new_n698_) );
  NAND2_X1 g340 ( .A1(new_n698_), .A2(G29), .ZN(new_n699_) );
  INV_X1 g341 ( .A(G1966), .ZN(new_n700_) );
  XNOR2_X1 g342 ( .A(G168), .B(new_n700_), .ZN(new_n701_) );
  XOR2_X1 g343 ( .A(G305), .B(G1981), .Z(new_n702_) );
  INV_X1 g344 ( .A(new_n702_), .ZN(new_n703_) );
  NOR2_X1 g345 ( .A1(new_n701_), .A2(new_n703_), .ZN(new_n704_) );
  XNOR2_X1 g346 ( .A(new_n704_), .B(KEYINPUT57), .ZN(new_n705_) );
  XOR2_X1 g347 ( .A(new_n511_), .B(G1956), .Z(new_n706_) );
  NAND2_X1 g348 ( .A1(G303), .A2(G1971), .ZN(new_n707_) );
  INV_X1 g349 ( .A(G1976), .ZN(new_n708_) );
  INV_X1 g350 ( .A(G288), .ZN(new_n709_) );
  NOR2_X1 g351 ( .A1(new_n709_), .A2(new_n708_), .ZN(new_n710_) );
  INV_X1 g352 ( .A(new_n710_), .ZN(new_n711_) );
  NAND2_X1 g353 ( .A1(new_n711_), .A2(new_n707_), .ZN(new_n712_) );
  NOR2_X1 g354 ( .A1(new_n712_), .A2(new_n706_), .ZN(new_n713_) );
  INV_X1 g355 ( .A(G1986), .ZN(new_n714_) );
  XNOR2_X1 g356 ( .A(new_n539_), .B(new_n714_), .ZN(new_n715_) );
  NOR2_X1 g357 ( .A1(G303), .A2(G1971), .ZN(new_n716_) );
  NOR2_X1 g358 ( .A1(G288), .A2(G1976), .ZN(new_n717_) );
  NOR2_X1 g359 ( .A1(new_n716_), .A2(new_n717_), .ZN(new_n718_) );
  INV_X1 g360 ( .A(new_n718_), .ZN(new_n719_) );
  NOR2_X1 g361 ( .A1(new_n719_), .A2(new_n715_), .ZN(new_n720_) );
  NAND2_X1 g362 ( .A1(new_n713_), .A2(new_n720_), .ZN(new_n721_) );
  XNOR2_X1 g363 ( .A(new_n549_), .B(G1348), .ZN(new_n722_) );
  NOR2_X1 g364 ( .A1(new_n721_), .A2(new_n722_), .ZN(new_n723_) );
  INV_X1 g365 ( .A(G1961), .ZN(new_n724_) );
  XNOR2_X1 g366 ( .A(G171), .B(new_n724_), .ZN(new_n725_) );
  INV_X1 g367 ( .A(G1341), .ZN(new_n726_) );
  XNOR2_X1 g368 ( .A(new_n498_), .B(new_n726_), .ZN(new_n727_) );
  NOR2_X1 g369 ( .A1(new_n725_), .A2(new_n727_), .ZN(new_n728_) );
  NAND2_X1 g370 ( .A1(new_n723_), .A2(new_n728_), .ZN(new_n729_) );
  NOR2_X1 g371 ( .A1(new_n705_), .A2(new_n729_), .ZN(new_n730_) );
  XOR2_X1 g372 ( .A(G16), .B(KEYINPUT56), .Z(new_n731_) );
  NOR2_X1 g373 ( .A1(new_n730_), .A2(new_n731_), .ZN(new_n732_) );
  INV_X1 g374 ( .A(G29), .ZN(new_n733_) );
  INV_X1 g375 ( .A(KEYINPUT53), .ZN(new_n734_) );
  XNOR2_X1 g376 ( .A(G26), .B(G2067), .ZN(new_n735_) );
  NAND2_X1 g377 ( .A1(G32), .A2(G1996), .ZN(new_n736_) );
  NAND2_X1 g378 ( .A1(new_n736_), .A2(G28), .ZN(new_n737_) );
  INV_X1 g379 ( .A(new_n737_), .ZN(new_n738_) );
  NOR2_X1 g380 ( .A1(G32), .A2(G1996), .ZN(new_n739_) );
  NOR2_X1 g381 ( .A1(G33), .A2(G2072), .ZN(new_n740_) );
  NOR2_X1 g382 ( .A1(new_n739_), .A2(new_n740_), .ZN(new_n741_) );
  NAND2_X1 g383 ( .A1(new_n738_), .A2(new_n741_), .ZN(new_n742_) );
  NOR2_X1 g384 ( .A1(new_n742_), .A2(new_n735_), .ZN(new_n743_) );
  INV_X1 g385 ( .A(G27), .ZN(new_n744_) );
  XNOR2_X1 g386 ( .A(G2078), .B(KEYINPUT25), .ZN(new_n745_) );
  NOR2_X1 g387 ( .A1(new_n745_), .A2(new_n744_), .ZN(new_n746_) );
  NAND2_X1 g388 ( .A1(new_n745_), .A2(new_n744_), .ZN(new_n747_) );
  NOR2_X1 g389 ( .A1(G25), .A2(G1991), .ZN(new_n748_) );
  NAND2_X1 g390 ( .A1(G33), .A2(G2072), .ZN(new_n749_) );
  NAND2_X1 g391 ( .A1(G25), .A2(G1991), .ZN(new_n750_) );
  NAND2_X1 g392 ( .A1(new_n749_), .A2(new_n750_), .ZN(new_n751_) );
  NOR2_X1 g393 ( .A1(new_n751_), .A2(new_n748_), .ZN(new_n752_) );
  NAND2_X1 g394 ( .A1(new_n747_), .A2(new_n752_), .ZN(new_n753_) );
  NOR2_X1 g395 ( .A1(new_n753_), .A2(new_n746_), .ZN(new_n754_) );
  NAND2_X1 g396 ( .A1(new_n754_), .A2(new_n743_), .ZN(new_n755_) );
  NAND2_X1 g397 ( .A1(new_n755_), .A2(new_n734_), .ZN(new_n756_) );
  NOR2_X1 g398 ( .A1(new_n755_), .A2(new_n734_), .ZN(new_n757_) );
  XOR2_X1 g399 ( .A(G35), .B(G2090), .Z(new_n758_) );
  XOR2_X1 g400 ( .A(G2084), .B(KEYINPUT54), .Z(new_n759_) );
  XNOR2_X1 g401 ( .A(new_n759_), .B(G34), .ZN(new_n760_) );
  NAND2_X1 g402 ( .A1(new_n760_), .A2(new_n758_), .ZN(new_n761_) );
  NOR2_X1 g403 ( .A1(new_n757_), .A2(new_n761_), .ZN(new_n762_) );
  NAND2_X1 g404 ( .A1(new_n762_), .A2(new_n756_), .ZN(new_n763_) );
  XNOR2_X1 g405 ( .A(new_n763_), .B(new_n614_), .ZN(new_n764_) );
  NAND2_X1 g406 ( .A1(new_n764_), .A2(new_n733_), .ZN(new_n765_) );
  INV_X1 g407 ( .A(G16), .ZN(new_n766_) );
  XOR2_X1 g408 ( .A(G22), .B(G1971), .Z(new_n767_) );
  XNOR2_X1 g409 ( .A(G23), .B(G1976), .ZN(new_n768_) );
  XNOR2_X1 g410 ( .A(G24), .B(G1986), .ZN(new_n769_) );
  NOR2_X1 g411 ( .A1(new_n768_), .A2(new_n769_), .ZN(new_n770_) );
  NAND2_X1 g412 ( .A1(new_n770_), .A2(new_n767_), .ZN(new_n771_) );
  NOR2_X1 g413 ( .A1(new_n771_), .A2(KEYINPUT58), .ZN(new_n772_) );
  NAND2_X1 g414 ( .A1(new_n771_), .A2(KEYINPUT58), .ZN(new_n773_) );
  XNOR2_X1 g415 ( .A(G21), .B(G1966), .ZN(new_n774_) );
  XNOR2_X1 g416 ( .A(G5), .B(G1961), .ZN(new_n775_) );
  NOR2_X1 g417 ( .A1(new_n774_), .A2(new_n775_), .ZN(new_n776_) );
  NAND2_X1 g418 ( .A1(new_n773_), .A2(new_n776_), .ZN(new_n777_) );
  NOR2_X1 g419 ( .A1(new_n777_), .A2(new_n772_), .ZN(new_n778_) );
  XOR2_X1 g420 ( .A(G1348), .B(KEYINPUT59), .Z(new_n779_) );
  XNOR2_X1 g421 ( .A(new_n779_), .B(G4), .ZN(new_n780_) );
  XOR2_X1 g422 ( .A(G20), .B(G1956), .Z(new_n781_) );
  XNOR2_X1 g423 ( .A(G6), .B(G1981), .ZN(new_n782_) );
  XNOR2_X1 g424 ( .A(G19), .B(G1341), .ZN(new_n783_) );
  NOR2_X1 g425 ( .A1(new_n782_), .A2(new_n783_), .ZN(new_n784_) );
  NAND2_X1 g426 ( .A1(new_n784_), .A2(new_n781_), .ZN(new_n785_) );
  NOR2_X1 g427 ( .A1(new_n780_), .A2(new_n785_), .ZN(new_n786_) );
  XNOR2_X1 g428 ( .A(new_n786_), .B(KEYINPUT60), .ZN(new_n787_) );
  NAND2_X1 g429 ( .A1(new_n787_), .A2(new_n778_), .ZN(new_n788_) );
  XOR2_X1 g430 ( .A(new_n788_), .B(KEYINPUT61), .Z(new_n789_) );
  NAND2_X1 g431 ( .A1(new_n789_), .A2(new_n766_), .ZN(new_n790_) );
  NAND2_X1 g432 ( .A1(new_n790_), .A2(G11), .ZN(new_n791_) );
  INV_X1 g433 ( .A(new_n791_), .ZN(new_n792_) );
  NAND2_X1 g434 ( .A1(new_n792_), .A2(new_n765_), .ZN(new_n793_) );
  NOR2_X1 g435 ( .A1(new_n732_), .A2(new_n793_), .ZN(new_n794_) );
  NAND2_X1 g436 ( .A1(new_n699_), .A2(new_n794_), .ZN(new_n795_) );
  XOR2_X1 g437 ( .A(new_n795_), .B(KEYINPUT62), .Z(G311) );
  INV_X1 g438 ( .A(G311), .ZN(G150) );
  NAND2_X1 g439 ( .A1(new_n558_), .A2(G559), .ZN(new_n798_) );
  NOR2_X1 g440 ( .A1(new_n798_), .A2(new_n563_), .ZN(new_n799_) );
  NAND2_X1 g441 ( .A1(new_n798_), .A2(new_n563_), .ZN(new_n800_) );
  NAND2_X1 g442 ( .A1(new_n800_), .A2(new_n559_), .ZN(new_n801_) );
  NOR2_X1 g443 ( .A1(new_n801_), .A2(new_n799_), .ZN(new_n802_) );
  NAND2_X1 g444 ( .A1(new_n446_), .A2(G93), .ZN(new_n803_) );
  NAND2_X1 g445 ( .A1(new_n450_), .A2(G67), .ZN(new_n804_) );
  NAND2_X1 g446 ( .A1(new_n804_), .A2(new_n803_), .ZN(new_n805_) );
  INV_X1 g447 ( .A(new_n805_), .ZN(new_n806_) );
  INV_X1 g448 ( .A(G55), .ZN(new_n807_) );
  INV_X1 g449 ( .A(new_n454_), .ZN(new_n808_) );
  NOR2_X1 g450 ( .A1(new_n808_), .A2(new_n807_), .ZN(new_n809_) );
  INV_X1 g451 ( .A(G80), .ZN(new_n810_) );
  INV_X1 g452 ( .A(new_n457_), .ZN(new_n811_) );
  NOR2_X1 g453 ( .A1(new_n811_), .A2(new_n810_), .ZN(new_n812_) );
  NOR2_X1 g454 ( .A1(new_n809_), .A2(new_n812_), .ZN(new_n813_) );
  NAND2_X1 g455 ( .A1(new_n813_), .A2(new_n806_), .ZN(new_n814_) );
  XOR2_X1 g456 ( .A(new_n802_), .B(new_n814_), .Z(G145) );
  INV_X1 g457 ( .A(KEYINPUT45), .ZN(new_n816_) );
  NAND2_X1 g458 ( .A1(new_n416_), .A2(G142), .ZN(new_n817_) );
  NAND2_X1 g459 ( .A1(new_n427_), .A2(G106), .ZN(new_n818_) );
  NAND2_X1 g460 ( .A1(new_n817_), .A2(new_n818_), .ZN(new_n819_) );
  NOR2_X1 g461 ( .A1(new_n819_), .A2(new_n816_), .ZN(new_n820_) );
  NAND2_X1 g462 ( .A1(new_n819_), .A2(new_n816_), .ZN(new_n821_) );
  INV_X1 g463 ( .A(G118), .ZN(new_n822_) );
  NOR2_X1 g464 ( .A1(new_n408_), .A2(new_n822_), .ZN(new_n823_) );
  INV_X1 g465 ( .A(G130), .ZN(new_n824_) );
  INV_X1 g466 ( .A(new_n423_), .ZN(new_n825_) );
  NOR2_X1 g467 ( .A1(new_n825_), .A2(new_n824_), .ZN(new_n826_) );
  NOR2_X1 g468 ( .A1(new_n826_), .A2(new_n823_), .ZN(new_n827_) );
  NAND2_X1 g469 ( .A1(new_n821_), .A2(new_n827_), .ZN(new_n828_) );
  NOR2_X1 g470 ( .A1(new_n828_), .A2(new_n820_), .ZN(new_n829_) );
  XNOR2_X1 g471 ( .A(new_n829_), .B(new_n652_), .ZN(new_n830_) );
  XNOR2_X1 g472 ( .A(new_n830_), .B(G162), .ZN(new_n831_) );
  INV_X1 g473 ( .A(G160), .ZN(new_n832_) );
  XNOR2_X1 g474 ( .A(new_n629_), .B(new_n832_), .ZN(new_n833_) );
  XNOR2_X1 g475 ( .A(new_n670_), .B(new_n833_), .ZN(new_n834_) );
  XNOR2_X1 g476 ( .A(new_n834_), .B(new_n831_), .ZN(new_n835_) );
  INV_X1 g477 ( .A(new_n835_), .ZN(new_n836_) );
  XNOR2_X1 g478 ( .A(new_n580_), .B(new_n684_), .ZN(new_n837_) );
  XNOR2_X1 g479 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(new_n838_) );
  XNOR2_X1 g480 ( .A(new_n837_), .B(new_n838_), .ZN(new_n839_) );
  XNOR2_X1 g481 ( .A(new_n839_), .B(new_n444_), .ZN(new_n840_) );
  NOR2_X1 g482 ( .A1(new_n836_), .A2(new_n840_), .ZN(new_n841_) );
  INV_X1 g483 ( .A(G37), .ZN(new_n842_) );
  NAND2_X1 g484 ( .A1(new_n836_), .A2(new_n840_), .ZN(new_n843_) );
  NAND2_X1 g485 ( .A1(new_n843_), .A2(new_n842_), .ZN(new_n844_) );
  NOR2_X1 g486 ( .A1(new_n844_), .A2(new_n841_), .ZN(G395) );
  XNOR2_X1 g487 ( .A(new_n498_), .B(new_n539_), .ZN(new_n846_) );
  XNOR2_X1 g488 ( .A(new_n846_), .B(G288), .ZN(new_n847_) );
  XOR2_X1 g489 ( .A(new_n511_), .B(KEYINPUT19), .Z(new_n848_) );
  XNOR2_X1 g490 ( .A(new_n848_), .B(G305), .ZN(new_n849_) );
  XNOR2_X1 g491 ( .A(new_n847_), .B(new_n849_), .ZN(new_n850_) );
  XNOR2_X1 g492 ( .A(new_n814_), .B(G303), .ZN(new_n851_) );
  XNOR2_X1 g493 ( .A(new_n850_), .B(new_n851_), .ZN(new_n852_) );
  XOR2_X1 g494 ( .A(new_n852_), .B(new_n798_), .Z(new_n853_) );
  NAND2_X1 g495 ( .A1(new_n853_), .A2(G868), .ZN(new_n854_) );
  NAND2_X1 g496 ( .A1(new_n814_), .A2(new_n541_), .ZN(new_n855_) );
  NAND2_X1 g497 ( .A1(new_n854_), .A2(new_n855_), .ZN(G295) );
  XNOR2_X1 g498 ( .A(G286), .B(new_n558_), .ZN(new_n857_) );
  XNOR2_X1 g499 ( .A(new_n852_), .B(new_n857_), .ZN(new_n858_) );
  INV_X1 g500 ( .A(new_n858_), .ZN(new_n859_) );
  NOR2_X1 g501 ( .A1(new_n859_), .A2(G301), .ZN(new_n860_) );
  NOR2_X1 g502 ( .A1(new_n858_), .A2(G171), .ZN(new_n861_) );
  NOR2_X1 g503 ( .A1(new_n861_), .A2(G37), .ZN(new_n862_) );
  INV_X1 g504 ( .A(new_n862_), .ZN(new_n863_) );
  NOR2_X1 g505 ( .A1(new_n863_), .A2(new_n860_), .ZN(G397) );
  INV_X1 g506 ( .A(KEYINPUT33), .ZN(new_n865_) );
  INV_X1 g507 ( .A(KEYINPUT29), .ZN(new_n866_) );
  INV_X1 g508 ( .A(KEYINPUT26), .ZN(new_n867_) );
  INV_X1 g509 ( .A(G1384), .ZN(new_n868_) );
  NAND2_X1 g510 ( .A1(new_n444_), .A2(new_n868_), .ZN(new_n869_) );
  NAND2_X1 g511 ( .A1(G160), .A2(G40), .ZN(new_n870_) );
  NOR2_X1 g512 ( .A1(new_n870_), .A2(new_n869_), .ZN(new_n871_) );
  NAND2_X1 g513 ( .A1(new_n871_), .A2(G1996), .ZN(new_n872_) );
  XNOR2_X1 g514 ( .A(new_n872_), .B(new_n867_), .ZN(new_n873_) );
  NOR2_X1 g515 ( .A1(new_n871_), .A2(new_n726_), .ZN(new_n874_) );
  INV_X1 g516 ( .A(new_n874_), .ZN(new_n875_) );
  NAND2_X1 g517 ( .A1(new_n875_), .A2(new_n498_), .ZN(new_n876_) );
  NOR2_X1 g518 ( .A1(new_n873_), .A2(new_n876_), .ZN(new_n877_) );
  NAND2_X1 g519 ( .A1(new_n877_), .A2(new_n558_), .ZN(new_n878_) );
  INV_X1 g520 ( .A(new_n871_), .ZN(new_n879_) );
  NAND2_X1 g521 ( .A1(new_n879_), .A2(G1348), .ZN(new_n880_) );
  NAND2_X1 g522 ( .A1(new_n871_), .A2(G2067), .ZN(new_n881_) );
  NAND2_X1 g523 ( .A1(new_n880_), .A2(new_n881_), .ZN(new_n882_) );
  NAND2_X1 g524 ( .A1(new_n878_), .A2(new_n882_), .ZN(new_n883_) );
  INV_X1 g525 ( .A(new_n877_), .ZN(new_n884_) );
  NAND2_X1 g526 ( .A1(new_n884_), .A2(new_n549_), .ZN(new_n885_) );
  NAND2_X1 g527 ( .A1(new_n883_), .A2(new_n885_), .ZN(new_n886_) );
  NAND2_X1 g528 ( .A1(new_n871_), .A2(G2072), .ZN(new_n887_) );
  NOR2_X1 g529 ( .A1(new_n887_), .A2(KEYINPUT27), .ZN(new_n888_) );
  NAND2_X1 g530 ( .A1(new_n879_), .A2(G1956), .ZN(new_n889_) );
  NAND2_X1 g531 ( .A1(new_n887_), .A2(KEYINPUT27), .ZN(new_n890_) );
  NAND2_X1 g532 ( .A1(new_n890_), .A2(new_n889_), .ZN(new_n891_) );
  NOR2_X1 g533 ( .A1(new_n891_), .A2(new_n888_), .ZN(new_n892_) );
  NAND2_X1 g534 ( .A1(new_n892_), .A2(new_n511_), .ZN(new_n893_) );
  NAND2_X1 g535 ( .A1(new_n886_), .A2(new_n893_), .ZN(new_n894_) );
  NOR2_X1 g536 ( .A1(new_n892_), .A2(new_n511_), .ZN(new_n895_) );
  XOR2_X1 g537 ( .A(new_n895_), .B(KEYINPUT28), .Z(new_n896_) );
  NAND2_X1 g538 ( .A1(new_n894_), .A2(new_n896_), .ZN(new_n897_) );
  XNOR2_X1 g539 ( .A(new_n897_), .B(new_n866_), .ZN(new_n898_) );
  NAND2_X1 g540 ( .A1(new_n879_), .A2(new_n724_), .ZN(new_n899_) );
  NAND2_X1 g541 ( .A1(new_n871_), .A2(new_n745_), .ZN(new_n900_) );
  NAND2_X1 g542 ( .A1(new_n899_), .A2(new_n900_), .ZN(new_n901_) );
  NAND2_X1 g543 ( .A1(new_n901_), .A2(G171), .ZN(new_n902_) );
  NAND2_X1 g544 ( .A1(new_n898_), .A2(new_n902_), .ZN(new_n903_) );
  INV_X1 g545 ( .A(G8), .ZN(new_n904_) );
  NOR2_X1 g546 ( .A1(new_n871_), .A2(new_n904_), .ZN(new_n905_) );
  NAND2_X1 g547 ( .A1(new_n905_), .A2(new_n700_), .ZN(new_n906_) );
  INV_X1 g548 ( .A(G2084), .ZN(new_n907_) );
  NAND2_X1 g549 ( .A1(new_n871_), .A2(new_n907_), .ZN(new_n908_) );
  NAND2_X1 g550 ( .A1(new_n908_), .A2(G8), .ZN(new_n909_) );
  INV_X1 g551 ( .A(new_n909_), .ZN(new_n910_) );
  NAND2_X1 g552 ( .A1(new_n910_), .A2(new_n906_), .ZN(new_n911_) );
  NOR2_X1 g553 ( .A1(new_n911_), .A2(KEYINPUT30), .ZN(new_n912_) );
  INV_X1 g554 ( .A(G168), .ZN(new_n913_) );
  NAND2_X1 g555 ( .A1(new_n911_), .A2(KEYINPUT30), .ZN(new_n914_) );
  NAND2_X1 g556 ( .A1(new_n914_), .A2(new_n913_), .ZN(new_n915_) );
  NOR2_X1 g557 ( .A1(new_n915_), .A2(new_n912_), .ZN(new_n916_) );
  NOR2_X1 g558 ( .A1(new_n901_), .A2(G171), .ZN(new_n917_) );
  NOR2_X1 g559 ( .A1(new_n916_), .A2(new_n917_), .ZN(new_n918_) );
  XOR2_X1 g560 ( .A(new_n918_), .B(KEYINPUT31), .Z(new_n919_) );
  NAND2_X1 g561 ( .A1(new_n903_), .A2(new_n919_), .ZN(new_n920_) );
  NAND2_X1 g562 ( .A1(new_n920_), .A2(G286), .ZN(new_n921_) );
  INV_X1 g563 ( .A(G1971), .ZN(new_n922_) );
  NAND2_X1 g564 ( .A1(new_n905_), .A2(new_n922_), .ZN(new_n923_) );
  INV_X1 g565 ( .A(G2090), .ZN(new_n924_) );
  NAND2_X1 g566 ( .A1(new_n871_), .A2(new_n924_), .ZN(new_n925_) );
  NAND2_X1 g567 ( .A1(new_n925_), .A2(G303), .ZN(new_n926_) );
  INV_X1 g568 ( .A(new_n926_), .ZN(new_n927_) );
  NAND2_X1 g569 ( .A1(new_n927_), .A2(new_n923_), .ZN(new_n928_) );
  NAND2_X1 g570 ( .A1(new_n921_), .A2(new_n928_), .ZN(new_n929_) );
  NAND2_X1 g571 ( .A1(new_n929_), .A2(G8), .ZN(new_n930_) );
  XNOR2_X1 g572 ( .A(new_n930_), .B(KEYINPUT32), .ZN(new_n931_) );
  INV_X1 g573 ( .A(new_n906_), .ZN(new_n932_) );
  NOR2_X1 g574 ( .A1(new_n908_), .A2(new_n904_), .ZN(new_n933_) );
  NOR2_X1 g575 ( .A1(new_n932_), .A2(new_n933_), .ZN(new_n934_) );
  NAND2_X1 g576 ( .A1(new_n920_), .A2(new_n934_), .ZN(new_n935_) );
  NAND2_X1 g577 ( .A1(new_n931_), .A2(new_n935_), .ZN(new_n936_) );
  NAND2_X1 g578 ( .A1(new_n936_), .A2(new_n718_), .ZN(new_n937_) );
  INV_X1 g579 ( .A(new_n905_), .ZN(new_n938_) );
  NOR2_X1 g580 ( .A1(new_n938_), .A2(new_n710_), .ZN(new_n939_) );
  NAND2_X1 g581 ( .A1(new_n937_), .A2(new_n939_), .ZN(new_n940_) );
  NAND2_X1 g582 ( .A1(new_n940_), .A2(new_n865_), .ZN(new_n941_) );
  NAND2_X1 g583 ( .A1(new_n717_), .A2(KEYINPUT33), .ZN(new_n942_) );
  NOR2_X1 g584 ( .A1(new_n938_), .A2(new_n942_), .ZN(new_n943_) );
  NOR2_X1 g585 ( .A1(new_n703_), .A2(new_n943_), .ZN(new_n944_) );
  NAND2_X1 g586 ( .A1(new_n941_), .A2(new_n944_), .ZN(new_n945_) );
  NOR2_X1 g587 ( .A1(new_n904_), .A2(G2090), .ZN(new_n946_) );
  NAND2_X1 g588 ( .A1(G166), .A2(new_n946_), .ZN(new_n947_) );
  NAND2_X1 g589 ( .A1(new_n936_), .A2(new_n947_), .ZN(new_n948_) );
  NAND2_X1 g590 ( .A1(new_n948_), .A2(new_n938_), .ZN(new_n949_) );
  INV_X1 g591 ( .A(KEYINPUT24), .ZN(new_n950_) );
  NOR2_X1 g592 ( .A1(G305), .A2(G1981), .ZN(new_n951_) );
  NAND2_X1 g593 ( .A1(new_n951_), .A2(new_n950_), .ZN(new_n952_) );
  NOR2_X1 g594 ( .A1(new_n951_), .A2(new_n950_), .ZN(new_n953_) );
  NOR2_X1 g595 ( .A1(new_n953_), .A2(new_n938_), .ZN(new_n954_) );
  NAND2_X1 g596 ( .A1(new_n954_), .A2(new_n952_), .ZN(new_n955_) );
  NAND2_X1 g597 ( .A1(new_n949_), .A2(new_n955_), .ZN(new_n956_) );
  INV_X1 g598 ( .A(new_n956_), .ZN(new_n957_) );
  NAND2_X1 g599 ( .A1(new_n945_), .A2(new_n957_), .ZN(new_n958_) );
  INV_X1 g600 ( .A(new_n869_), .ZN(new_n959_) );
  NOR2_X1 g601 ( .A1(new_n870_), .A2(new_n959_), .ZN(new_n960_) );
  NAND2_X1 g602 ( .A1(new_n674_), .A2(new_n960_), .ZN(new_n961_) );
  INV_X1 g603 ( .A(new_n961_), .ZN(new_n962_) );
  NAND2_X1 g604 ( .A1(new_n687_), .A2(new_n960_), .ZN(new_n963_) );
  NAND2_X1 g605 ( .A1(new_n715_), .A2(new_n960_), .ZN(new_n964_) );
  NAND2_X1 g606 ( .A1(new_n963_), .A2(new_n964_), .ZN(new_n965_) );
  NOR2_X1 g607 ( .A1(new_n962_), .A2(new_n965_), .ZN(new_n966_) );
  NAND2_X1 g608 ( .A1(new_n958_), .A2(new_n966_), .ZN(new_n967_) );
  INV_X1 g609 ( .A(new_n689_), .ZN(new_n968_) );
  NAND2_X1 g610 ( .A1(new_n539_), .A2(new_n714_), .ZN(new_n969_) );
  NAND2_X1 g611 ( .A1(new_n969_), .A2(new_n968_), .ZN(new_n970_) );
  NAND2_X1 g612 ( .A1(new_n963_), .A2(new_n970_), .ZN(new_n971_) );
  NAND2_X1 g613 ( .A1(new_n971_), .A2(new_n654_), .ZN(new_n972_) );
  XOR2_X1 g614 ( .A(new_n972_), .B(KEYINPUT39), .Z(new_n973_) );
  NAND2_X1 g615 ( .A1(new_n973_), .A2(new_n961_), .ZN(new_n974_) );
  NAND2_X1 g616 ( .A1(new_n974_), .A2(new_n673_), .ZN(new_n975_) );
  NAND2_X1 g617 ( .A1(new_n975_), .A2(new_n960_), .ZN(new_n976_) );
  NAND2_X1 g618 ( .A1(new_n967_), .A2(new_n976_), .ZN(new_n977_) );
  XNOR2_X1 g619 ( .A(new_n977_), .B(KEYINPUT40), .ZN(G329) );
  NOR2_X1 g620 ( .A1(G229), .A2(G227), .ZN(new_n980_) );
  NOR2_X1 g621 ( .A1(new_n980_), .A2(KEYINPUT49), .ZN(new_n981_) );
  NAND2_X1 g622 ( .A1(new_n980_), .A2(KEYINPUT49), .ZN(new_n982_) );
  INV_X1 g623 ( .A(new_n982_), .ZN(new_n983_) );
  INV_X1 g624 ( .A(G401), .ZN(new_n984_) );
  NAND2_X1 g625 ( .A1(new_n984_), .A2(G319), .ZN(new_n985_) );
  NOR2_X1 g626 ( .A1(new_n983_), .A2(new_n985_), .ZN(new_n986_) );
  INV_X1 g627 ( .A(new_n986_), .ZN(new_n987_) );
  NOR2_X1 g628 ( .A1(new_n987_), .A2(new_n981_), .ZN(new_n988_) );
  INV_X1 g629 ( .A(new_n988_), .ZN(new_n989_) );
  NOR2_X1 g630 ( .A1(G395), .A2(new_n989_), .ZN(new_n990_) );
  INV_X1 g631 ( .A(new_n990_), .ZN(new_n991_) );
  NOR2_X1 g632 ( .A1(G397), .A2(new_n991_), .ZN(G308) );
  INV_X1 g633 ( .A(G308), .ZN(G225) );
  assign   G231 = 1'b0;
  BUF_X1 g634 ( .A(G452), .Z(G350) );
  BUF_X1 g635 ( .A(G452), .Z(G335) );
  BUF_X1 g636 ( .A(G452), .Z(G409) );
  BUF_X1 g637 ( .A(G1083), .Z(G369) );
  BUF_X1 g638 ( .A(G1083), .Z(G367) );
  BUF_X1 g639 ( .A(G2066), .Z(G411) );
  BUF_X1 g640 ( .A(G2066), .Z(G337) );
  BUF_X1 g641 ( .A(G2066), .Z(G384) );
  BUF_X1 g642 ( .A(G452), .Z(G391) );
  NAND2_X1 g643 ( .A1(new_n551_), .A2(new_n550_), .ZN(G321) );
  INV_X1 g644 ( .A(new_n556_), .ZN(G280) );
  NOR2_X1 g645 ( .A1(new_n564_), .A2(new_n567_), .ZN(G323) );
  NAND2_X1 g646 ( .A1(new_n854_), .A2(new_n855_), .ZN(G331) );
endmodule


