module add_mul_mix_8_bit ( a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, 
        b_0_, b_1_, b_2_, b_3_, b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, 
        c_4_, c_5_, c_6_, c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_, 
        Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_, 
        Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_, 
        Result_12_, Result_13_, Result_14_, Result_15_ );
  input a_0_, a_1_, a_2_, a_3_, a_4_, a_5_, a_6_, a_7_, b_0_, b_1_, b_2_, b_3_,
         b_4_, b_5_, b_6_, b_7_, c_0_, c_1_, c_2_, c_3_, c_4_, c_5_, c_6_,
         c_7_, d_0_, d_1_, d_2_, d_3_, d_4_, d_5_, d_6_, d_7_;
  output Result_0_, Result_1_, Result_2_, Result_3_, Result_4_, Result_5_,
         Result_6_, Result_7_, Result_8_, Result_9_, Result_10_, Result_11_,
         Result_12_, Result_13_, Result_14_, Result_15_;
  wire   n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968;

  XNOR2_X1 U472 ( .A(n456), .B(n457), .ZN(Result_9_) );
  XNOR2_X1 U473 ( .A(n458), .B(n459), .ZN(n457) );
  XNOR2_X1 U474 ( .A(n460), .B(n461), .ZN(Result_8_) );
  XNOR2_X1 U475 ( .A(n462), .B(n463), .ZN(n461) );
  XOR2_X1 U476 ( .A(n464), .B(n465), .Z(Result_7_) );
  NOR2_X1 U477 ( .A1(n466), .A2(n467), .ZN(Result_6_) );
  NOR2_X1 U478 ( .A1(n468), .A2(n469), .ZN(n467) );
  XNOR2_X1 U479 ( .A(n466), .B(n470), .ZN(Result_5_) );
  NAND2_X1 U480 ( .A1(n471), .A2(n472), .ZN(n470) );
  NAND2_X1 U481 ( .A1(n473), .A2(n474), .ZN(n472) );
  INV_X1 U482 ( .A(n475), .ZN(n474) );
  NAND2_X1 U483 ( .A1(n476), .A2(n477), .ZN(n473) );
  XOR2_X1 U484 ( .A(n478), .B(n479), .Z(Result_4_) );
  XNOR2_X1 U485 ( .A(n480), .B(n481), .ZN(Result_3_) );
  NAND2_X1 U486 ( .A1(n482), .A2(n483), .ZN(n481) );
  XNOR2_X1 U487 ( .A(n484), .B(n485), .ZN(Result_2_) );
  NAND2_X1 U488 ( .A1(n486), .A2(n487), .ZN(n484) );
  XOR2_X1 U489 ( .A(n488), .B(n489), .Z(Result_1_) );
  NAND2_X1 U490 ( .A1(n490), .A2(n491), .ZN(n488) );
  XOR2_X1 U491 ( .A(n492), .B(n493), .Z(Result_14_) );
  NOR2_X1 U492 ( .A1(n494), .A2(n495), .ZN(n493) );
  XNOR2_X1 U493 ( .A(n496), .B(n497), .ZN(Result_13_) );
  NAND2_X1 U494 ( .A1(n498), .A2(n499), .ZN(n496) );
  XOR2_X1 U495 ( .A(n500), .B(n501), .Z(Result_12_) );
  NOR2_X1 U496 ( .A1(n502), .A2(n503), .ZN(n500) );
  INV_X1 U497 ( .A(n504), .ZN(n503) );
  NOR2_X1 U498 ( .A1(n505), .A2(n506), .ZN(n502) );
  NOR2_X1 U499 ( .A1(n495), .A2(n507), .ZN(n505) );
  XNOR2_X1 U500 ( .A(n508), .B(n509), .ZN(Result_11_) );
  XOR2_X1 U501 ( .A(n510), .B(n511), .Z(n509) );
  NAND2_X1 U502 ( .A1(n512), .A2(n513), .ZN(n511) );
  XOR2_X1 U503 ( .A(n514), .B(n515), .Z(Result_10_) );
  XOR2_X1 U504 ( .A(n516), .B(n517), .Z(n515) );
  NAND2_X1 U505 ( .A1(n518), .A2(n519), .ZN(Result_0_) );
  NAND2_X1 U506 ( .A1(n520), .A2(n521), .ZN(n519) );
  NOR2_X1 U507 ( .A1(n522), .A2(n523), .ZN(n518) );
  NOR2_X1 U508 ( .A1(n489), .A2(n524), .ZN(n523) );
  INV_X1 U509 ( .A(n491), .ZN(n524) );
  NAND2_X1 U510 ( .A1(n525), .A2(n526), .ZN(n491) );
  NAND2_X1 U511 ( .A1(n527), .A2(n528), .ZN(n526) );
  XOR2_X1 U512 ( .A(n521), .B(n529), .Z(n525) );
  AND2_X1 U513 ( .A1(n486), .A2(n530), .ZN(n489) );
  NAND2_X1 U514 ( .A1(n487), .A2(n485), .ZN(n530) );
  NAND2_X1 U515 ( .A1(n482), .A2(n531), .ZN(n485) );
  NAND2_X1 U516 ( .A1(n480), .A2(n483), .ZN(n531) );
  NAND2_X1 U517 ( .A1(n532), .A2(n533), .ZN(n483) );
  OR2_X1 U518 ( .A1(n534), .A2(n535), .ZN(n533) );
  XNOR2_X1 U519 ( .A(n536), .B(n537), .ZN(n532) );
  AND2_X1 U520 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U521 ( .A1(n538), .A2(n539), .ZN(n478) );
  NAND2_X1 U522 ( .A1(n466), .A2(n475), .ZN(n539) );
  AND2_X1 U523 ( .A1(n468), .A2(n469), .ZN(n466) );
  XOR2_X1 U524 ( .A(n477), .B(n476), .Z(n469) );
  NOR2_X1 U525 ( .A1(n464), .A2(n465), .ZN(n468) );
  XOR2_X1 U526 ( .A(n540), .B(n541), .Z(n465) );
  XOR2_X1 U527 ( .A(n542), .B(n543), .Z(n541) );
  NAND2_X1 U528 ( .A1(n520), .A2(n544), .ZN(n543) );
  AND2_X1 U529 ( .A1(n545), .A2(n546), .ZN(n464) );
  NAND2_X1 U530 ( .A1(n463), .A2(n547), .ZN(n546) );
  OR2_X1 U531 ( .A1(n462), .A2(n460), .ZN(n547) );
  NOR2_X1 U532 ( .A1(n548), .A2(n495), .ZN(n463) );
  NAND2_X1 U533 ( .A1(n460), .A2(n462), .ZN(n545) );
  NAND2_X1 U534 ( .A1(n549), .A2(n550), .ZN(n462) );
  NAND2_X1 U535 ( .A1(n459), .A2(n551), .ZN(n550) );
  NAND2_X1 U536 ( .A1(n458), .A2(n456), .ZN(n551) );
  NOR2_X1 U537 ( .A1(n552), .A2(n495), .ZN(n459) );
  OR2_X1 U538 ( .A1(n456), .A2(n458), .ZN(n549) );
  AND2_X1 U539 ( .A1(n553), .A2(n554), .ZN(n458) );
  NAND2_X1 U540 ( .A1(n517), .A2(n555), .ZN(n554) );
  OR2_X1 U541 ( .A1(n516), .A2(n514), .ZN(n555) );
  NOR2_X1 U542 ( .A1(n556), .A2(n495), .ZN(n517) );
  NAND2_X1 U543 ( .A1(n514), .A2(n516), .ZN(n553) );
  NAND2_X1 U544 ( .A1(n557), .A2(n558), .ZN(n516) );
  NAND2_X1 U545 ( .A1(n559), .A2(n512), .ZN(n558) );
  NOR2_X1 U546 ( .A1(n560), .A2(n495), .ZN(n559) );
  NOR2_X1 U547 ( .A1(n508), .A2(n510), .ZN(n560) );
  NAND2_X1 U548 ( .A1(n508), .A2(n510), .ZN(n557) );
  NAND2_X1 U549 ( .A1(n504), .A2(n561), .ZN(n510) );
  NAND2_X1 U550 ( .A1(n501), .A2(n562), .ZN(n561) );
  NAND2_X1 U551 ( .A1(n563), .A2(n564), .ZN(n562) );
  NAND2_X1 U552 ( .A1(n565), .A2(n513), .ZN(n564) );
  INV_X1 U553 ( .A(n506), .ZN(n563) );
  XOR2_X1 U554 ( .A(n566), .B(n567), .Z(n501) );
  XNOR2_X1 U555 ( .A(n568), .B(n569), .ZN(n567) );
  NAND2_X1 U556 ( .A1(n570), .A2(n544), .ZN(n569) );
  NAND2_X1 U557 ( .A1(n565), .A2(n506), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n498), .A2(n571), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n497), .A2(n499), .ZN(n571) );
  NAND2_X1 U560 ( .A1(n572), .A2(n573), .ZN(n499) );
  NAND2_X1 U561 ( .A1(n570), .A2(n513), .ZN(n572) );
  INV_X1 U562 ( .A(n495), .ZN(n513) );
  XOR2_X1 U563 ( .A(n574), .B(n575), .Z(n497) );
  NOR2_X1 U564 ( .A1(n576), .A2(n577), .ZN(n575) );
  OR2_X1 U565 ( .A1(n573), .A2(n578), .ZN(n498) );
  NAND2_X1 U566 ( .A1(Result_15_), .A2(n574), .ZN(n573) );
  NOR2_X1 U567 ( .A1(n579), .A2(n494), .ZN(n574) );
  NOR2_X1 U568 ( .A1(n495), .A2(n576), .ZN(Result_15_) );
  XOR2_X1 U569 ( .A(n580), .B(d_7_), .Z(n495) );
  XOR2_X1 U570 ( .A(n581), .B(n582), .Z(n508) );
  XOR2_X1 U571 ( .A(n583), .B(n584), .Z(n581) );
  XOR2_X1 U572 ( .A(n585), .B(n586), .Z(n514) );
  XOR2_X1 U573 ( .A(n587), .B(n588), .Z(n585) );
  NOR2_X1 U574 ( .A1(n579), .A2(n589), .ZN(n588) );
  XNOR2_X1 U575 ( .A(n590), .B(n591), .ZN(n456) );
  XOR2_X1 U576 ( .A(n592), .B(n593), .Z(n590) );
  NOR2_X1 U577 ( .A1(n579), .A2(n556), .ZN(n593) );
  XNOR2_X1 U578 ( .A(n594), .B(n595), .ZN(n460) );
  XOR2_X1 U579 ( .A(n596), .B(n597), .Z(n595) );
  NAND2_X1 U580 ( .A1(n598), .A2(n544), .ZN(n597) );
  INV_X1 U581 ( .A(n579), .ZN(n544) );
  NOR2_X1 U582 ( .A1(n599), .A2(n600), .ZN(n538) );
  INV_X1 U583 ( .A(n471), .ZN(n599) );
  NAND2_X1 U584 ( .A1(n601), .A2(n475), .ZN(n471) );
  NOR2_X1 U585 ( .A1(n600), .A2(n602), .ZN(n475) );
  AND2_X1 U586 ( .A1(n603), .A2(n604), .ZN(n602) );
  NOR2_X1 U587 ( .A1(n604), .A2(n603), .ZN(n600) );
  AND2_X1 U588 ( .A1(n605), .A2(n606), .ZN(n603) );
  NAND2_X1 U589 ( .A1(n607), .A2(n608), .ZN(n606) );
  NOR2_X1 U590 ( .A1(n609), .A2(n548), .ZN(n607) );
  NOR2_X1 U591 ( .A1(n610), .A2(n611), .ZN(n609) );
  NAND2_X1 U592 ( .A1(n611), .A2(n610), .ZN(n605) );
  XNOR2_X1 U593 ( .A(n612), .B(n613), .ZN(n604) );
  XNOR2_X1 U594 ( .A(n614), .B(n615), .ZN(n613) );
  AND2_X1 U595 ( .A1(n477), .A2(n476), .ZN(n601) );
  XOR2_X1 U596 ( .A(n616), .B(n611), .Z(n476) );
  XOR2_X1 U597 ( .A(n617), .B(n618), .Z(n611) );
  XOR2_X1 U598 ( .A(n619), .B(n620), .Z(n617) );
  NOR2_X1 U599 ( .A1(n621), .A2(n552), .ZN(n620) );
  XNOR2_X1 U600 ( .A(n622), .B(n610), .ZN(n616) );
  NAND2_X1 U601 ( .A1(n623), .A2(n624), .ZN(n610) );
  NAND2_X1 U602 ( .A1(n625), .A2(n598), .ZN(n624) );
  NOR2_X1 U603 ( .A1(n626), .A2(n577), .ZN(n625) );
  NOR2_X1 U604 ( .A1(n627), .A2(n628), .ZN(n626) );
  NAND2_X1 U605 ( .A1(n628), .A2(n627), .ZN(n623) );
  NAND2_X1 U606 ( .A1(n608), .A2(n520), .ZN(n622) );
  NAND2_X1 U607 ( .A1(n629), .A2(n630), .ZN(n477) );
  NAND2_X1 U608 ( .A1(n631), .A2(n520), .ZN(n630) );
  NOR2_X1 U609 ( .A1(n632), .A2(n579), .ZN(n631) );
  NOR2_X1 U610 ( .A1(n540), .A2(n542), .ZN(n632) );
  NAND2_X1 U611 ( .A1(n540), .A2(n542), .ZN(n629) );
  NAND2_X1 U612 ( .A1(n633), .A2(n634), .ZN(n542) );
  NAND2_X1 U613 ( .A1(n635), .A2(n598), .ZN(n634) );
  NOR2_X1 U614 ( .A1(n636), .A2(n579), .ZN(n635) );
  NOR2_X1 U615 ( .A1(n596), .A2(n594), .ZN(n636) );
  NAND2_X1 U616 ( .A1(n594), .A2(n596), .ZN(n633) );
  NAND2_X1 U617 ( .A1(n637), .A2(n638), .ZN(n596) );
  NAND2_X1 U618 ( .A1(n639), .A2(n640), .ZN(n638) );
  NOR2_X1 U619 ( .A1(n641), .A2(n579), .ZN(n639) );
  NOR2_X1 U620 ( .A1(n592), .A2(n591), .ZN(n641) );
  NAND2_X1 U621 ( .A1(n591), .A2(n592), .ZN(n637) );
  NAND2_X1 U622 ( .A1(n642), .A2(n643), .ZN(n592) );
  NAND2_X1 U623 ( .A1(n644), .A2(n512), .ZN(n643) );
  NOR2_X1 U624 ( .A1(n645), .A2(n579), .ZN(n644) );
  NOR2_X1 U625 ( .A1(n586), .A2(n587), .ZN(n645) );
  NAND2_X1 U626 ( .A1(n586), .A2(n587), .ZN(n642) );
  NAND2_X1 U627 ( .A1(n646), .A2(n647), .ZN(n587) );
  NAND2_X1 U628 ( .A1(n584), .A2(n648), .ZN(n647) );
  OR2_X1 U629 ( .A1(n583), .A2(n582), .ZN(n648) );
  NOR2_X1 U630 ( .A1(n507), .A2(n579), .ZN(n584) );
  NAND2_X1 U631 ( .A1(n582), .A2(n583), .ZN(n646) );
  NAND2_X1 U632 ( .A1(n649), .A2(n650), .ZN(n583) );
  NAND2_X1 U633 ( .A1(n651), .A2(n570), .ZN(n650) );
  NOR2_X1 U634 ( .A1(n652), .A2(n579), .ZN(n651) );
  NOR2_X1 U635 ( .A1(n568), .A2(n566), .ZN(n652) );
  NAND2_X1 U636 ( .A1(n568), .A2(n566), .ZN(n649) );
  XOR2_X1 U637 ( .A(n653), .B(n654), .Z(n566) );
  AND2_X1 U638 ( .A1(n492), .A2(n654), .ZN(n568) );
  NOR2_X1 U639 ( .A1(n579), .A2(n576), .ZN(n492) );
  XOR2_X1 U640 ( .A(n655), .B(n656), .Z(n579) );
  XOR2_X1 U641 ( .A(d_6_), .B(c_6_), .Z(n656) );
  NAND2_X1 U642 ( .A1(d_7_), .A2(c_7_), .ZN(n655) );
  XNOR2_X1 U643 ( .A(n657), .B(n658), .ZN(n582) );
  XOR2_X1 U644 ( .A(n659), .B(n660), .Z(n658) );
  NAND2_X1 U645 ( .A1(n608), .A2(n570), .ZN(n657) );
  XOR2_X1 U646 ( .A(n661), .B(n662), .Z(n586) );
  NOR2_X1 U647 ( .A1(n663), .A2(n664), .ZN(n662) );
  NOR2_X1 U648 ( .A1(n665), .A2(n666), .ZN(n663) );
  NOR2_X1 U649 ( .A1(n507), .A2(n577), .ZN(n665) );
  XNOR2_X1 U650 ( .A(n667), .B(n668), .ZN(n591) );
  XNOR2_X1 U651 ( .A(n669), .B(n670), .ZN(n667) );
  XNOR2_X1 U652 ( .A(n671), .B(n672), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n673), .A2(n674), .ZN(n671) );
  XNOR2_X1 U654 ( .A(n628), .B(n675), .ZN(n540) );
  XOR2_X1 U655 ( .A(n627), .B(n676), .Z(n675) );
  NAND2_X1 U656 ( .A1(n598), .A2(n608), .ZN(n676) );
  NAND2_X1 U657 ( .A1(n673), .A2(n677), .ZN(n627) );
  NAND2_X1 U658 ( .A1(n672), .A2(n674), .ZN(n677) );
  NAND2_X1 U659 ( .A1(n678), .A2(n679), .ZN(n674) );
  NAND2_X1 U660 ( .A1(n640), .A2(n608), .ZN(n679) );
  INV_X1 U661 ( .A(n680), .ZN(n678) );
  XNOR2_X1 U662 ( .A(n681), .B(n682), .ZN(n672) );
  XOR2_X1 U663 ( .A(n683), .B(n684), .Z(n682) );
  NAND2_X1 U664 ( .A1(n640), .A2(n680), .ZN(n673) );
  NAND2_X1 U665 ( .A1(n685), .A2(n686), .ZN(n680) );
  NAND2_X1 U666 ( .A1(n670), .A2(n687), .ZN(n686) );
  NAND2_X1 U667 ( .A1(n669), .A2(n668), .ZN(n687) );
  NOR2_X1 U668 ( .A1(n589), .A2(n577), .ZN(n670) );
  OR2_X1 U669 ( .A1(n668), .A2(n669), .ZN(n685) );
  NOR2_X1 U670 ( .A1(n664), .A2(n688), .ZN(n669) );
  AND2_X1 U671 ( .A1(n661), .A2(n689), .ZN(n688) );
  NAND2_X1 U672 ( .A1(n690), .A2(n691), .ZN(n689) );
  NAND2_X1 U673 ( .A1(n608), .A2(n565), .ZN(n691) );
  XOR2_X1 U674 ( .A(n692), .B(n693), .Z(n661) );
  XOR2_X1 U675 ( .A(n694), .B(n695), .Z(n693) );
  NAND2_X1 U676 ( .A1(n696), .A2(n570), .ZN(n695) );
  NOR2_X1 U677 ( .A1(n507), .A2(n690), .ZN(n664) );
  INV_X1 U678 ( .A(n666), .ZN(n690) );
  NAND2_X1 U679 ( .A1(n697), .A2(n698), .ZN(n666) );
  NAND2_X1 U680 ( .A1(n699), .A2(n608), .ZN(n698) );
  NOR2_X1 U681 ( .A1(n700), .A2(n578), .ZN(n699) );
  NOR2_X1 U682 ( .A1(n660), .A2(n659), .ZN(n700) );
  NAND2_X1 U683 ( .A1(n659), .A2(n660), .ZN(n697) );
  AND2_X1 U684 ( .A1(n694), .A2(n701), .ZN(n660) );
  NAND2_X1 U685 ( .A1(n702), .A2(n703), .ZN(n701) );
  OR2_X1 U686 ( .A1(n704), .A2(n576), .ZN(n703) );
  NAND2_X1 U687 ( .A1(n696), .A2(n705), .ZN(n702) );
  AND2_X1 U688 ( .A1(n654), .A2(n653), .ZN(n659) );
  NOR2_X1 U689 ( .A1(n577), .A2(n494), .ZN(n654) );
  INV_X1 U690 ( .A(n608), .ZN(n577) );
  XOR2_X1 U691 ( .A(n706), .B(n707), .Z(n608) );
  XOR2_X1 U692 ( .A(d_5_), .B(c_5_), .Z(n707) );
  XOR2_X1 U693 ( .A(n708), .B(n709), .Z(n668) );
  XOR2_X1 U694 ( .A(n710), .B(n711), .Z(n708) );
  XOR2_X1 U695 ( .A(n712), .B(n713), .Z(n628) );
  NOR2_X1 U696 ( .A1(n714), .A2(n715), .ZN(n713) );
  INV_X1 U697 ( .A(n716), .ZN(n715) );
  NOR2_X1 U698 ( .A1(n717), .A2(n718), .ZN(n714) );
  NOR2_X1 U699 ( .A1(n621), .A2(n556), .ZN(n718) );
  XOR2_X1 U700 ( .A(n534), .B(n535), .Z(n479) );
  NAND2_X1 U701 ( .A1(n719), .A2(n720), .ZN(n482) );
  XOR2_X1 U702 ( .A(n537), .B(n536), .Z(n720) );
  NOR2_X1 U703 ( .A1(n534), .A2(n535), .ZN(n719) );
  XNOR2_X1 U704 ( .A(n721), .B(n722), .ZN(n535) );
  NOR2_X1 U705 ( .A1(n723), .A2(n724), .ZN(n722) );
  NOR2_X1 U706 ( .A1(n725), .A2(n726), .ZN(n723) );
  NOR2_X1 U707 ( .A1(n548), .A2(n704), .ZN(n726) );
  INV_X1 U708 ( .A(n727), .ZN(n725) );
  NAND2_X1 U709 ( .A1(n728), .A2(n729), .ZN(n534) );
  NAND2_X1 U710 ( .A1(n614), .A2(n730), .ZN(n729) );
  OR2_X1 U711 ( .A1(n612), .A2(n615), .ZN(n730) );
  AND2_X1 U712 ( .A1(n731), .A2(n732), .ZN(n614) );
  NAND2_X1 U713 ( .A1(n733), .A2(n598), .ZN(n732) );
  NOR2_X1 U714 ( .A1(n734), .A2(n621), .ZN(n733) );
  NOR2_X1 U715 ( .A1(n618), .A2(n619), .ZN(n734) );
  NAND2_X1 U716 ( .A1(n618), .A2(n619), .ZN(n731) );
  NAND2_X1 U717 ( .A1(n716), .A2(n735), .ZN(n619) );
  NAND2_X1 U718 ( .A1(n712), .A2(n736), .ZN(n735) );
  NAND2_X1 U719 ( .A1(n737), .A2(n738), .ZN(n736) );
  NAND2_X1 U720 ( .A1(n640), .A2(n696), .ZN(n738) );
  XOR2_X1 U721 ( .A(n739), .B(n740), .Z(n712) );
  XNOR2_X1 U722 ( .A(n741), .B(n742), .ZN(n740) );
  NAND2_X1 U723 ( .A1(n717), .A2(n640), .ZN(n716) );
  INV_X1 U724 ( .A(n737), .ZN(n717) );
  NAND2_X1 U725 ( .A1(n743), .A2(n744), .ZN(n737) );
  NAND2_X1 U726 ( .A1(n681), .A2(n745), .ZN(n744) );
  OR2_X1 U727 ( .A1(n684), .A2(n683), .ZN(n745) );
  XOR2_X1 U728 ( .A(n746), .B(n747), .Z(n681) );
  NAND2_X1 U729 ( .A1(n748), .A2(n749), .ZN(n746) );
  NAND2_X1 U730 ( .A1(n684), .A2(n683), .ZN(n743) );
  NAND2_X1 U731 ( .A1(n750), .A2(n751), .ZN(n683) );
  NAND2_X1 U732 ( .A1(n709), .A2(n752), .ZN(n751) );
  NAND2_X1 U733 ( .A1(n711), .A2(n710), .ZN(n752) );
  XOR2_X1 U734 ( .A(n753), .B(n754), .Z(n709) );
  XOR2_X1 U735 ( .A(n755), .B(n756), .Z(n754) );
  NAND2_X1 U736 ( .A1(n757), .A2(n570), .ZN(n753) );
  OR2_X1 U737 ( .A1(n710), .A2(n711), .ZN(n750) );
  NOR2_X1 U738 ( .A1(n507), .A2(n621), .ZN(n711) );
  NAND2_X1 U739 ( .A1(n758), .A2(n759), .ZN(n710) );
  NAND2_X1 U740 ( .A1(n760), .A2(n696), .ZN(n759) );
  NOR2_X1 U741 ( .A1(n761), .A2(n578), .ZN(n760) );
  NOR2_X1 U742 ( .A1(n762), .A2(n692), .ZN(n761) );
  NAND2_X1 U743 ( .A1(n762), .A2(n692), .ZN(n758) );
  XOR2_X1 U744 ( .A(n763), .B(n764), .Z(n692) );
  INV_X1 U745 ( .A(n694), .ZN(n762) );
  NAND2_X1 U746 ( .A1(n653), .A2(n763), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n621), .A2(n576), .ZN(n653) );
  INV_X1 U748 ( .A(n696), .ZN(n621) );
  NAND2_X1 U749 ( .A1(n512), .A2(n696), .ZN(n684) );
  XOR2_X1 U750 ( .A(n765), .B(n766), .Z(n618) );
  XNOR2_X1 U751 ( .A(n767), .B(n768), .ZN(n766) );
  NAND2_X1 U752 ( .A1(n640), .A2(n757), .ZN(n768) );
  NAND2_X1 U753 ( .A1(n612), .A2(n615), .ZN(n728) );
  NAND2_X1 U754 ( .A1(n696), .A2(n520), .ZN(n615) );
  XOR2_X1 U755 ( .A(n769), .B(n770), .Z(n696) );
  XOR2_X1 U756 ( .A(d_4_), .B(c_4_), .Z(n770) );
  XNOR2_X1 U757 ( .A(n771), .B(n772), .ZN(n612) );
  XNOR2_X1 U758 ( .A(n773), .B(n774), .ZN(n771) );
  NAND2_X1 U759 ( .A1(n775), .A2(n776), .ZN(n487) );
  OR2_X1 U760 ( .A1(n537), .A2(n536), .ZN(n776) );
  XNOR2_X1 U761 ( .A(n528), .B(n527), .ZN(n775) );
  NAND2_X1 U762 ( .A1(n777), .A2(n778), .ZN(n486) );
  XOR2_X1 U763 ( .A(n528), .B(n527), .Z(n778) );
  NOR2_X1 U764 ( .A1(n536), .A2(n537), .ZN(n777) );
  XNOR2_X1 U765 ( .A(n779), .B(n780), .ZN(n537) );
  XOR2_X1 U766 ( .A(n781), .B(n782), .Z(n779) );
  NOR2_X1 U767 ( .A1(n548), .A2(n783), .ZN(n782) );
  NOR2_X1 U768 ( .A1(n724), .A2(n784), .ZN(n536) );
  AND2_X1 U769 ( .A1(n721), .A2(n785), .ZN(n784) );
  NAND2_X1 U770 ( .A1(n727), .A2(n786), .ZN(n785) );
  NAND2_X1 U771 ( .A1(n757), .A2(n520), .ZN(n786) );
  XNOR2_X1 U772 ( .A(n787), .B(n788), .ZN(n721) );
  NAND2_X1 U773 ( .A1(n789), .A2(n790), .ZN(n787) );
  NOR2_X1 U774 ( .A1(n727), .A2(n548), .ZN(n724) );
  NAND2_X1 U775 ( .A1(n791), .A2(n792), .ZN(n727) );
  NAND2_X1 U776 ( .A1(n774), .A2(n793), .ZN(n792) );
  NAND2_X1 U777 ( .A1(n773), .A2(n772), .ZN(n793) );
  AND2_X1 U778 ( .A1(n794), .A2(n795), .ZN(n774) );
  NAND2_X1 U779 ( .A1(n796), .A2(n640), .ZN(n795) );
  NOR2_X1 U780 ( .A1(n797), .A2(n704), .ZN(n796) );
  NOR2_X1 U781 ( .A1(n767), .A2(n765), .ZN(n797) );
  NAND2_X1 U782 ( .A1(n765), .A2(n767), .ZN(n794) );
  AND2_X1 U783 ( .A1(n798), .A2(n799), .ZN(n767) );
  NAND2_X1 U784 ( .A1(n741), .A2(n800), .ZN(n799) );
  OR2_X1 U785 ( .A1(n739), .A2(n742), .ZN(n800) );
  AND2_X1 U786 ( .A1(n748), .A2(n801), .ZN(n741) );
  NAND2_X1 U787 ( .A1(n747), .A2(n749), .ZN(n801) );
  NAND2_X1 U788 ( .A1(n802), .A2(n803), .ZN(n749) );
  NAND2_X1 U789 ( .A1(n565), .A2(n757), .ZN(n803) );
  INV_X1 U790 ( .A(n804), .ZN(n802) );
  XOR2_X1 U791 ( .A(n805), .B(n806), .Z(n747) );
  XNOR2_X1 U792 ( .A(n807), .B(n808), .ZN(n806) );
  NAND2_X1 U793 ( .A1(n809), .A2(n570), .ZN(n808) );
  NAND2_X1 U794 ( .A1(n565), .A2(n804), .ZN(n748) );
  NAND2_X1 U795 ( .A1(n810), .A2(n811), .ZN(n804) );
  NAND2_X1 U796 ( .A1(n812), .A2(n757), .ZN(n811) );
  NOR2_X1 U797 ( .A1(n813), .A2(n578), .ZN(n812) );
  NOR2_X1 U798 ( .A1(n755), .A2(n756), .ZN(n813) );
  NAND2_X1 U799 ( .A1(n756), .A2(n755), .ZN(n810) );
  AND2_X1 U800 ( .A1(n764), .A2(n763), .ZN(n755) );
  NOR2_X1 U801 ( .A1(n704), .A2(n494), .ZN(n763) );
  NOR2_X1 U802 ( .A1(n576), .A2(n783), .ZN(n764) );
  NOR2_X1 U803 ( .A1(n807), .A2(n814), .ZN(n756) );
  AND2_X1 U804 ( .A1(n815), .A2(n816), .ZN(n814) );
  NAND2_X1 U805 ( .A1(n739), .A2(n742), .ZN(n798) );
  NAND2_X1 U806 ( .A1(n512), .A2(n757), .ZN(n742) );
  XNOR2_X1 U807 ( .A(n817), .B(n818), .ZN(n739) );
  XOR2_X1 U808 ( .A(n819), .B(n820), .Z(n817) );
  XNOR2_X1 U809 ( .A(n821), .B(n822), .ZN(n765) );
  NAND2_X1 U810 ( .A1(n823), .A2(n824), .ZN(n821) );
  OR2_X1 U811 ( .A1(n772), .A2(n773), .ZN(n791) );
  NOR2_X1 U812 ( .A1(n552), .A2(n704), .ZN(n773) );
  INV_X1 U813 ( .A(n757), .ZN(n704) );
  XOR2_X1 U814 ( .A(n825), .B(n826), .Z(n757) );
  XOR2_X1 U815 ( .A(d_3_), .B(c_3_), .Z(n826) );
  XOR2_X1 U816 ( .A(n827), .B(n828), .Z(n772) );
  XOR2_X1 U817 ( .A(n829), .B(n830), .Z(n827) );
  NOR2_X1 U818 ( .A1(n783), .A2(n556), .ZN(n830) );
  INV_X1 U819 ( .A(n490), .ZN(n522) );
  NAND2_X1 U820 ( .A1(n831), .A2(n832), .ZN(n490) );
  AND2_X1 U821 ( .A1(n528), .A2(n527), .ZN(n832) );
  XOR2_X1 U822 ( .A(n833), .B(n834), .Z(n527) );
  NOR2_X1 U823 ( .A1(n835), .A2(n836), .ZN(n834) );
  INV_X1 U824 ( .A(n837), .ZN(n836) );
  NOR2_X1 U825 ( .A1(n838), .A2(n839), .ZN(n835) );
  NAND2_X1 U826 ( .A1(n840), .A2(n841), .ZN(n528) );
  NAND2_X1 U827 ( .A1(n842), .A2(n809), .ZN(n841) );
  NOR2_X1 U828 ( .A1(n843), .A2(n548), .ZN(n842) );
  NOR2_X1 U829 ( .A1(n780), .A2(n781), .ZN(n843) );
  NAND2_X1 U830 ( .A1(n780), .A2(n781), .ZN(n840) );
  NAND2_X1 U831 ( .A1(n789), .A2(n844), .ZN(n781) );
  NAND2_X1 U832 ( .A1(n788), .A2(n790), .ZN(n844) );
  NAND2_X1 U833 ( .A1(n845), .A2(n846), .ZN(n790) );
  NAND2_X1 U834 ( .A1(n598), .A2(n809), .ZN(n846) );
  INV_X1 U835 ( .A(n847), .ZN(n845) );
  XOR2_X1 U836 ( .A(n848), .B(n849), .Z(n788) );
  XOR2_X1 U837 ( .A(n850), .B(n851), .Z(n848) );
  NAND2_X1 U838 ( .A1(n598), .A2(n847), .ZN(n789) );
  NAND2_X1 U839 ( .A1(n852), .A2(n853), .ZN(n847) );
  NAND2_X1 U840 ( .A1(n854), .A2(n640), .ZN(n853) );
  NOR2_X1 U841 ( .A1(n855), .A2(n783), .ZN(n854) );
  NOR2_X1 U842 ( .A1(n828), .A2(n829), .ZN(n855) );
  NAND2_X1 U843 ( .A1(n828), .A2(n829), .ZN(n852) );
  NAND2_X1 U844 ( .A1(n823), .A2(n856), .ZN(n829) );
  NAND2_X1 U845 ( .A1(n822), .A2(n824), .ZN(n856) );
  NAND2_X1 U846 ( .A1(n857), .A2(n858), .ZN(n824) );
  NAND2_X1 U847 ( .A1(n512), .A2(n809), .ZN(n858) );
  INV_X1 U848 ( .A(n859), .ZN(n857) );
  XOR2_X1 U849 ( .A(n860), .B(n861), .Z(n822) );
  NOR2_X1 U850 ( .A1(n862), .A2(n578), .ZN(n861) );
  XOR2_X1 U851 ( .A(n863), .B(n864), .Z(n860) );
  NAND2_X1 U852 ( .A1(n512), .A2(n859), .ZN(n823) );
  NAND2_X1 U853 ( .A1(n865), .A2(n866), .ZN(n859) );
  NAND2_X1 U854 ( .A1(n820), .A2(n867), .ZN(n866) );
  OR2_X1 U855 ( .A1(n818), .A2(n819), .ZN(n867) );
  NOR2_X1 U856 ( .A1(n507), .A2(n783), .ZN(n820) );
  INV_X1 U857 ( .A(n809), .ZN(n783) );
  NAND2_X1 U858 ( .A1(n818), .A2(n819), .ZN(n865) );
  NAND2_X1 U859 ( .A1(n868), .A2(n869), .ZN(n819) );
  NAND2_X1 U860 ( .A1(n870), .A2(n809), .ZN(n869) );
  NOR2_X1 U861 ( .A1(n871), .A2(n578), .ZN(n870) );
  NOR2_X1 U862 ( .A1(n807), .A2(n805), .ZN(n871) );
  NAND2_X1 U863 ( .A1(n807), .A2(n805), .ZN(n868) );
  XNOR2_X1 U864 ( .A(n872), .B(n873), .ZN(n805) );
  NOR2_X1 U865 ( .A1(n576), .A2(n862), .ZN(n873) );
  OR2_X1 U866 ( .A1(n874), .A2(n494), .ZN(n872) );
  NOR2_X1 U867 ( .A1(n816), .A2(n815), .ZN(n807) );
  INV_X1 U868 ( .A(n875), .ZN(n815) );
  NAND2_X1 U869 ( .A1(n809), .A2(n705), .ZN(n816) );
  INV_X1 U870 ( .A(n494), .ZN(n705) );
  XOR2_X1 U871 ( .A(n876), .B(n877), .Z(n809) );
  XOR2_X1 U872 ( .A(d_2_), .B(c_2_), .Z(n877) );
  XNOR2_X1 U873 ( .A(n878), .B(n879), .ZN(n818) );
  NAND2_X1 U874 ( .A1(n880), .A2(n881), .ZN(n878) );
  XOR2_X1 U875 ( .A(n882), .B(n883), .Z(n828) );
  NOR2_X1 U876 ( .A1(n884), .A2(n885), .ZN(n883) );
  INV_X1 U877 ( .A(n886), .ZN(n885) );
  NOR2_X1 U878 ( .A1(n887), .A2(n888), .ZN(n884) );
  XOR2_X1 U879 ( .A(n889), .B(n890), .Z(n780) );
  XNOR2_X1 U880 ( .A(n891), .B(n892), .ZN(n890) );
  NAND2_X1 U881 ( .A1(n640), .A2(n893), .ZN(n889) );
  NOR2_X1 U882 ( .A1(n521), .A2(n529), .ZN(n831) );
  NAND2_X1 U883 ( .A1(n520), .A2(n893), .ZN(n529) );
  INV_X1 U884 ( .A(n862), .ZN(n893) );
  NAND2_X1 U885 ( .A1(n837), .A2(n894), .ZN(n521) );
  NAND2_X1 U886 ( .A1(n895), .A2(n833), .ZN(n894) );
  NAND2_X1 U887 ( .A1(n896), .A2(n897), .ZN(n833) );
  NAND2_X1 U888 ( .A1(n898), .A2(n640), .ZN(n897) );
  NOR2_X1 U889 ( .A1(n899), .A2(n862), .ZN(n898) );
  NOR2_X1 U890 ( .A1(n892), .A2(n891), .ZN(n899) );
  NAND2_X1 U891 ( .A1(n892), .A2(n891), .ZN(n896) );
  NAND2_X1 U892 ( .A1(n900), .A2(n901), .ZN(n891) );
  NAND2_X1 U893 ( .A1(n849), .A2(n902), .ZN(n901) );
  OR2_X1 U894 ( .A1(n850), .A2(n851), .ZN(n902) );
  NOR2_X1 U895 ( .A1(n556), .A2(n874), .ZN(n849) );
  INV_X1 U896 ( .A(n640), .ZN(n556) );
  XOR2_X1 U897 ( .A(n903), .B(n904), .Z(n640) );
  XOR2_X1 U898 ( .A(b_2_), .B(a_2_), .Z(n904) );
  NAND2_X1 U899 ( .A1(n851), .A2(n850), .ZN(n900) );
  NAND2_X1 U900 ( .A1(n886), .A2(n905), .ZN(n850) );
  NAND2_X1 U901 ( .A1(n906), .A2(n882), .ZN(n905) );
  NAND2_X1 U902 ( .A1(n907), .A2(n908), .ZN(n882) );
  NAND2_X1 U903 ( .A1(n909), .A2(n570), .ZN(n908) );
  NOR2_X1 U904 ( .A1(n910), .A2(n862), .ZN(n909) );
  NOR2_X1 U905 ( .A1(n864), .A2(n863), .ZN(n910) );
  NAND2_X1 U906 ( .A1(n864), .A2(n863), .ZN(n907) );
  NAND2_X1 U907 ( .A1(n911), .A2(n881), .ZN(n863) );
  NAND2_X1 U908 ( .A1(n880), .A2(n875), .ZN(n881) );
  NOR2_X1 U909 ( .A1(n874), .A2(n576), .ZN(n875) );
  XOR2_X1 U910 ( .A(n912), .B(b_7_), .Z(n576) );
  NAND2_X1 U911 ( .A1(n879), .A2(n880), .ZN(n911) );
  NOR2_X1 U912 ( .A1(n862), .A2(n494), .ZN(n880) );
  XOR2_X1 U913 ( .A(n913), .B(n914), .Z(n494) );
  XOR2_X1 U914 ( .A(b_6_), .B(a_6_), .Z(n914) );
  NAND2_X1 U915 ( .A1(b_7_), .A2(a_7_), .ZN(n913) );
  NOR2_X1 U916 ( .A1(n874), .A2(n578), .ZN(n879) );
  INV_X1 U917 ( .A(n570), .ZN(n578) );
  XOR2_X1 U918 ( .A(n915), .B(n916), .Z(n570) );
  XOR2_X1 U919 ( .A(b_5_), .B(a_5_), .Z(n916) );
  NOR2_X1 U920 ( .A1(n507), .A2(n874), .ZN(n864) );
  OR2_X1 U921 ( .A1(n512), .A2(n887), .ZN(n906) );
  NAND2_X1 U922 ( .A1(n888), .A2(n887), .ZN(n886) );
  NOR2_X1 U923 ( .A1(n507), .A2(n862), .ZN(n887) );
  INV_X1 U924 ( .A(n565), .ZN(n507) );
  XOR2_X1 U925 ( .A(n917), .B(n918), .Z(n565) );
  XOR2_X1 U926 ( .A(b_4_), .B(a_4_), .Z(n918) );
  NOR2_X1 U927 ( .A1(n874), .A2(n589), .ZN(n888) );
  NOR2_X1 U928 ( .A1(n589), .A2(n862), .ZN(n851) );
  INV_X1 U929 ( .A(n512), .ZN(n589) );
  XOR2_X1 U930 ( .A(n919), .B(n920), .Z(n512) );
  XOR2_X1 U931 ( .A(b_3_), .B(a_3_), .Z(n920) );
  NOR2_X1 U932 ( .A1(n552), .A2(n874), .ZN(n892) );
  OR2_X1 U933 ( .A1(n520), .A2(n838), .ZN(n895) );
  INV_X1 U934 ( .A(n548), .ZN(n520) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n837) );
  NOR2_X1 U936 ( .A1(n552), .A2(n862), .ZN(n838) );
  XOR2_X1 U937 ( .A(n921), .B(n922), .Z(n862) );
  XOR2_X1 U938 ( .A(d_0_), .B(c_0_), .Z(n922) );
  NAND2_X1 U939 ( .A1(n923), .A2(n924), .ZN(n921) );
  NAND2_X1 U940 ( .A1(n925), .A2(n926), .ZN(n924) );
  INV_X1 U941 ( .A(d_1_), .ZN(n926) );
  NAND2_X1 U942 ( .A1(c_1_), .A2(n927), .ZN(n925) );
  OR2_X1 U943 ( .A1(n927), .A2(c_1_), .ZN(n923) );
  INV_X1 U944 ( .A(n598), .ZN(n552) );
  XOR2_X1 U945 ( .A(n928), .B(n929), .Z(n598) );
  XOR2_X1 U946 ( .A(b_1_), .B(a_1_), .Z(n929) );
  NOR2_X1 U947 ( .A1(n548), .A2(n874), .ZN(n839) );
  XNOR2_X1 U948 ( .A(n927), .B(n930), .ZN(n874) );
  XOR2_X1 U949 ( .A(d_1_), .B(c_1_), .Z(n930) );
  NAND2_X1 U950 ( .A1(n931), .A2(n932), .ZN(n927) );
  NAND2_X1 U951 ( .A1(d_2_), .A2(n933), .ZN(n932) );
  OR2_X1 U952 ( .A1(n876), .A2(c_2_), .ZN(n933) );
  NAND2_X1 U953 ( .A1(c_2_), .A2(n876), .ZN(n931) );
  NAND2_X1 U954 ( .A1(n934), .A2(n935), .ZN(n876) );
  NAND2_X1 U955 ( .A1(d_3_), .A2(n936), .ZN(n935) );
  OR2_X1 U956 ( .A1(n825), .A2(c_3_), .ZN(n936) );
  NAND2_X1 U957 ( .A1(c_3_), .A2(n825), .ZN(n934) );
  NAND2_X1 U958 ( .A1(n937), .A2(n938), .ZN(n825) );
  NAND2_X1 U959 ( .A1(d_4_), .A2(n939), .ZN(n938) );
  OR2_X1 U960 ( .A1(n769), .A2(c_4_), .ZN(n939) );
  NAND2_X1 U961 ( .A1(c_4_), .A2(n769), .ZN(n937) );
  NAND2_X1 U962 ( .A1(n940), .A2(n941), .ZN(n769) );
  NAND2_X1 U963 ( .A1(d_5_), .A2(n942), .ZN(n941) );
  OR2_X1 U964 ( .A1(n706), .A2(c_5_), .ZN(n942) );
  NAND2_X1 U965 ( .A1(c_5_), .A2(n706), .ZN(n940) );
  NAND2_X1 U966 ( .A1(n943), .A2(n944), .ZN(n706) );
  NAND2_X1 U967 ( .A1(n945), .A2(d_7_), .ZN(n944) );
  NOR2_X1 U968 ( .A1(n946), .A2(n580), .ZN(n945) );
  INV_X1 U969 ( .A(c_7_), .ZN(n580) );
  NOR2_X1 U970 ( .A1(c_6_), .A2(d_6_), .ZN(n946) );
  NAND2_X1 U971 ( .A1(d_6_), .A2(c_6_), .ZN(n943) );
  XOR2_X1 U972 ( .A(n947), .B(n948), .Z(n548) );
  XOR2_X1 U973 ( .A(b_0_), .B(a_0_), .Z(n948) );
  NAND2_X1 U974 ( .A1(n949), .A2(n950), .ZN(n947) );
  NAND2_X1 U975 ( .A1(n951), .A2(n952), .ZN(n950) );
  INV_X1 U976 ( .A(b_1_), .ZN(n952) );
  NAND2_X1 U977 ( .A1(a_1_), .A2(n928), .ZN(n951) );
  OR2_X1 U978 ( .A1(n928), .A2(a_1_), .ZN(n949) );
  NAND2_X1 U979 ( .A1(n953), .A2(n954), .ZN(n928) );
  NAND2_X1 U980 ( .A1(b_2_), .A2(n955), .ZN(n954) );
  OR2_X1 U981 ( .A1(n903), .A2(a_2_), .ZN(n955) );
  NAND2_X1 U982 ( .A1(a_2_), .A2(n903), .ZN(n953) );
  NAND2_X1 U983 ( .A1(n956), .A2(n957), .ZN(n903) );
  NAND2_X1 U984 ( .A1(b_3_), .A2(n958), .ZN(n957) );
  OR2_X1 U985 ( .A1(n919), .A2(a_3_), .ZN(n958) );
  NAND2_X1 U986 ( .A1(a_3_), .A2(n919), .ZN(n956) );
  NAND2_X1 U987 ( .A1(n959), .A2(n960), .ZN(n919) );
  NAND2_X1 U988 ( .A1(b_4_), .A2(n961), .ZN(n960) );
  OR2_X1 U989 ( .A1(n917), .A2(a_4_), .ZN(n961) );
  NAND2_X1 U990 ( .A1(a_4_), .A2(n917), .ZN(n959) );
  NAND2_X1 U991 ( .A1(n962), .A2(n963), .ZN(n917) );
  NAND2_X1 U992 ( .A1(b_5_), .A2(n964), .ZN(n963) );
  OR2_X1 U993 ( .A1(n915), .A2(a_5_), .ZN(n964) );
  NAND2_X1 U994 ( .A1(a_5_), .A2(n915), .ZN(n962) );
  NAND2_X1 U995 ( .A1(n965), .A2(n966), .ZN(n915) );
  NAND2_X1 U996 ( .A1(n967), .A2(b_7_), .ZN(n966) );
  NOR2_X1 U997 ( .A1(n968), .A2(n912), .ZN(n967) );
  INV_X1 U998 ( .A(a_7_), .ZN(n912) );
  NOR2_X1 U999 ( .A1(a_6_), .A2(b_6_), .ZN(n968) );
  NAND2_X1 U1000 ( .A1(b_6_), .A2(a_6_), .ZN(n965) );
endmodule

